Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_22x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A7: buffer std_logic
);
end x25_22x;

architecture x25_22x_behav of x25_22x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2196a,a2197a,a2198a,a2199a,a2200a,a2201a,a2202a,a2203a,a2204a,a2205a,a2206a,a2207a,a2208a,a2209a,a2210a,a2211a,a2212a,a2213a,a2214a,a2215a,a2216a,a2217a,a2218a,a2219a,a2220a,a2221a,a2222a,a2223a,a2224a,a2225a,a2226a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2237a,a2238a,a2239a,a2240a,a2241a,a2242a,a2243a,a2244a,a2245a,a2246a,a2247a,a2248a,a2249a,a2250a,a2251a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2258a,a2259a,a2260a,a2261a,a2262a,a2263a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2271a,a2272a,a2273a,a2274a,a2275a,a2276a,a2277a,a2278a,a2279a,a2280a,a2281a,a2282a,a2283a,a2284a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2297a,a2298a,a2299a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2306a,a2307a,a2308a,a2309a,a2310a,a2311a,a2312a,a2313a,a2314a,a2315a,a2316a,a2317a,a2318a,a2319a,a2320a,a2321a,a2322a,a2323a,a2324a,a2325a,a2326a,a2327a,a2328a,a2329a,a2330a,a2331a,a2332a,a2333a,a2334a,a2335a,a2336a,a2337a,a2338a,a2339a,a2340a,a2341a,a2342a,a2343a,a2344a,a2345a,a2346a,a2347a,a2348a,a2349a,a2350a,a2351a,a2352a,a2353a,a2354a,a2355a,a2356a,a2357a,a2358a,a2359a,a2360a,a2361a,a2362a,a2363a,a2364a,a2365a,a2366a,a2367a,a2368a,a2369a,a2370a,a2371a,a2372a,a2373a,a2374a,a2375a,a2376a,a2377a,a2378a,a2379a,a2380a,a2381a,a2382a,a2383a,a2384a,a2385a,a2386a,a2387a,a2388a,a2389a,a2390a,a2391a,a2392a,a2393a,a2394a,a2395a,a2396a,a2397a,a2398a,a2399a,a2400a,a2401a,a2402a,a2403a,a2404a,a2405a,a2406a,a2407a,a2408a,a2409a,a2410a,a2411a,a2412a,a2413a,a2414a,a2415a,a2416a,a2417a,a2418a,a2419a,a2420a,a2421a,a2422a,a2423a,a2424a,a2425a,a2426a,a2427a,a2428a,a2429a,a2430a,a2431a,a2432a,a2433a,a2434a,a2435a,a2436a,a2437a,a2438a,a2439a,a2440a,a2441a,a2442a,a2443a,a2444a,a2445a,a2446a,a2447a,a2448a,a2449a,a2450a,a2451a,a2452a,a2453a,a2454a,a2455a,a2456a,a2457a,a2458a,a2459a,a2460a,a2461a,a2462a,a2463a,a2464a,a2465a,a2466a,a2467a,a2468a,a2469a,a2470a,a2471a,a2472a,a2473a,a2474a,a2475a,a2476a,a2477a,a2478a,a2479a,a2480a,a2481a,a2482a,a2483a,a2484a,a2485a,a2486a,a2487a,a2488a,a2489a,a2490a,a2491a,a2492a,a2493a,a2494a,a2495a,a2496a,a2497a,a2498a,a2499a,a2500a,a2501a,a2502a,a2503a,a2504a,a2505a,a2506a,a2507a,a2508a,a2509a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2516a,a2517a,a2518a,a2519a,a2520a,a2521a,a2522a,a2523a,a2524a,a2525a,a2526a,a2527a,a2528a,a2529a,a2530a,a2531a,a2532a,a2533a,a2534a,a2535a,a2536a,a2537a,a2538a,a2539a,a2540a,a2541a,a2542a,a2543a,a2544a,a2545a,a2546a,a2547a,a2548a,a2549a,a2550a,a2551a,a2552a,a2553a,a2554a,a2555a,a2556a,a2557a,a2558a,a2559a,a2560a,a2561a,a2562a,a2563a,a2564a,a2565a,a2566a,a2567a,a2568a,a2569a,a2570a,a2571a,a2572a,a2573a,a2574a,a2575a,a2576a,a2577a,a2578a,a2579a,a2580a,a2581a,a2582a,a2583a,a2584a,a2585a,a2586a,a2587a,a2588a,a2589a,a2590a,a2591a,a2592a,a2593a,a2594a,a2595a,a2596a,a2597a,a2598a,a2599a,a2600a,a2601a,a2602a,a2603a,a2604a,a2605a,a2606a,a2607a,a2608a,a2609a,a2610a,a2611a,a2612a,a2613a,a2614a,a2615a,a2616a,a2617a,a2618a,a2619a,a2620a,a2621a,a2622a,a2623a,a2624a,a2625a,a2626a,a2627a,a2628a,a2629a,a2630a,a2631a,a2632a,a2633a,a2634a,a2635a,a2636a,a2637a,a2638a,a2639a,a2640a,a2641a,a2642a,a2643a,a2644a,a2645a,a2646a,a2647a,a2648a,a2649a,a2650a,a2651a,a2652a,a2653a,a2654a,a2655a,a2656a,a2657a,a2658a,a2659a,a2660a,a2661a,a2662a,a2663a,a2664a,a2665a,a2666a,a2667a,a2668a,a2669a,a2670a,a2671a,a2672a,a2673a,a2674a,a2675a,a2676a,a2677a,a2678a,a2679a,a2680a,a2681a,a2682a,a2683a,a2684a,a2685a,a2686a,a2687a,a2688a,a2689a,a2690a,a2691a,a2692a,a2693a,a2694a,a2695a,a2696a,a2697a,a2698a,a2699a,a2700a,a2701a,a2702a,a2703a,a2704a,a2705a,a2706a,a2707a,a2708a,a2709a,a2710a,a2711a,a2712a,a2713a,a2714a,a2715a,a2716a,a2717a,a2718a,a2719a,a2720a,a2721a,a2722a,a2723a,a2724a,a2725a,a2726a,a2727a,a2728a,a2729a,a2730a,a2731a,a2732a,a2733a,a2734a,a2735a,a2736a,a2737a,a2738a,a2739a,a2740a,a2741a,a2742a,a2743a,a2744a,a2745a,a2746a,a2747a,a2748a,a2749a,a2750a,a2751a,a2752a,a2753a,a2754a,a2755a,a2756a,a2757a,a2758a,a2759a,a2760a,a2761a,a2762a,a2763a,a2764a,a2765a,a2766a,a2767a,a2768a,a2769a,a2770a,a2771a,a2772a,a2773a,a2774a,a2775a,a2776a,a2777a,a2778a,a2779a,a2780a,a2781a,a2782a,a2783a,a2784a,a2785a,a2786a,a2787a,a2788a,a2789a,a2790a,a2791a,a2792a,a2793a,a2794a,a2795a,a2796a,a2797a,a2798a,a2799a,a2800a,a2801a,a2802a,a2803a,a2804a,a2805a,a2806a,a2807a,a2808a,a2809a,a2810a,a2811a,a2812a,a2813a,a2814a,a2815a,a2816a,a2817a,a2818a,a2819a,a2820a,a2821a,a2822a,a2823a,a2824a,a2825a,a2826a,a2827a,a2828a,a2829a,a2830a,a2831a,a2832a,a2833a,a2834a,a2835a,a2836a,a2837a,a2838a,a2839a,a2840a,a2841a,a2842a,a2843a,a2844a,a2845a,a2846a,a2847a,a2848a,a2849a,a2850a,a2851a,a2852a,a2853a,a2854a,a2855a,a2856a,a2857a,a2858a,a2859a,a2860a,a2861a,a2862a,a2863a,a2864a,a2865a,a2866a,a2867a,a2868a,a2869a,a2870a,a2871a,a2872a,a2873a,a2874a,a2875a,a2876a,a2877a,a2878a,a2879a,a2880a,a2881a,a2882a,a2883a,a2884a,a2885a,a2886a,a2887a,a2888a,a2889a,a2890a,a2891a,a2892a,a2893a,a2894a,a2895a,a2896a,a2897a,a2898a,a2899a,a2900a,a2901a,a2902a,a2903a,a2904a,a2905a,a2906a,a2907a,a2908a,a2909a,a2910a,a2911a,a2912a,a2913a,a2914a,a2915a,a2916a,a2917a,a2918a,a2919a,a2920a,a2921a,a2922a,a2923a,a2924a,a2925a,a2926a,a2927a,a2928a,a2929a,a2930a,a2931a,a2932a,a2933a,a2934a,a2935a,a2936a,a2937a,a2938a,a2939a,a2940a,a2941a,a2942a,a2943a,a2944a,a2945a,a2946a,a2947a,a2948a,a2949a,a2950a,a2951a,a2952a,a2953a,a2954a,a2955a,a2956a,a2957a,a2958a,a2959a,a2960a,a2961a,a2962a,a2963a,a2964a,a2965a,a2966a,a2967a,a2968a,a2969a,a2970a,a2971a,a2972a,a2973a,a2974a,a2975a,a2976a,a2977a,a2978a,a2979a,a2980a,a2981a,a2982a,a2983a,a2984a,a2985a,a2986a,a2987a,a2988a,a2989a,a2990a,a2991a,a2992a,a2993a,a2994a,a2995a,a2996a,a2997a,a2998a,a2999a,a3000a,a3001a,a3002a,a3003a,a3004a,a3005a,a3006a,a3007a,a3008a,a3009a,a3010a,a3011a,a3012a,a3013a,a3014a,a3015a,a3016a,a3017a,a3018a,a3019a,a3020a,a3021a,a3022a,a3023a,a3024a,a3025a,a3026a,a3027a,a3028a,a3029a,a3030a,a3031a,a3032a,a3033a,a3034a,a3035a,a3036a,a3037a,a3038a,a3039a,a3040a,a3041a,a3042a,a3043a,a3044a,a3045a,a3046a,a3047a,a3048a,a3049a,a3050a,a3051a,a3052a,a3053a,a3054a,a3055a,a3056a,a3057a,a3058a,a3059a,a3060a,a3061a,a3062a,a3063a,a3064a,a3065a,a3066a,a3067a,a3068a,a3069a,a3070a,a3071a,a3072a,a3073a,a3074a,a3075a,a3076a,a3077a,a3078a,a3079a,a3080a,a3081a,a3082a,a3083a,a3084a,a3085a,a3086a,a3087a,a3088a,a3089a,a3090a,a3091a,a3092a,a3093a,a3094a,a3095a,a3096a,a3097a,a3098a,a3099a,a3100a,a3101a,a3102a,a3103a,a3104a,a3105a,a3106a,a3107a,a3108a,a3109a,a3110a,a3111a,a3112a,a3113a,a3114a,a3115a,a3116a,a3117a,a3118a,a3119a,a3120a,a3121a,a3122a,a3123a,a3124a,a3125a,a3126a,a3127a,a3128a,a3129a,a3130a,a3131a,a3132a,a3133a,a3134a,a3135a,a3136a,a3137a,a3138a,a3139a,a3140a,a3141a,a3142a,a3143a,a3144a,a3145a,a3146a,a3147a,a3148a,a3149a,a3150a,a3151a,a3152a,a3153a,a3154a,a3155a,a3156a,a3157a,a3158a,a3159a,a3160a,a3161a,a3162a,a3163a,a3164a,a3165a,a3166a,a3167a,a3168a,a3169a,a3170a,a3171a,a3172a,a3173a,a3174a,a3175a,a3176a,a3177a,a3178a,a3179a,a3180a,a3181a,a3182a,a3183a,a3184a,a3185a,a3186a,a3187a,a3188a,a3189a,a3190a,a3191a,a3192a,a3193a,a3194a,a3195a,a3196a,a3197a,a3198a,a3199a,a3200a,a3201a,a3202a,a3203a,a3204a,a3205a,a3206a,a3207a,a3208a,a3209a,a3210a,a3211a,a3212a,a3213a,a3214a,a3215a,a3216a,a3217a,a3218a,a3219a,a3220a,a3221a,a3222a,a3223a,a3224a,a3225a,a3226a,a3227a,a3228a,a3229a,a3230a,a3231a,a3232a,a3233a,a3234a,a3235a,a3236a,a3237a,a3238a,a3239a,a3240a,a3241a,a3242a,a3243a,a3244a,a3245a,a3246a,a3247a,a3248a,a3249a,a3250a,a3251a,a3252a,a3253a,a3254a,a3255a,a3256a,a3257a,a3258a,a3259a,a3260a,a3261a,a3262a,a3263a,a3264a,a3265a,a3266a,a3267a,a3268a,a3269a,a3270a,a3271a,a3272a,a3273a,a3274a,a3275a,a3276a,a3277a,a3278a,a3279a,a3280a,a3281a,a3282a,a3283a,a3284a,a3285a,a3286a,a3287a,a3288a,a3289a,a3290a,a3291a,a3292a,a3293a,a3294a,a3295a,a3296a,a3297a,a3298a,a3299a,a3300a,a3301a,a3302a,a3303a,a3304a,a3305a,a3306a,a3307a,a3308a,a3309a,a3310a,a3311a,a3312a,a3313a,a3314a,a3315a,a3316a,a3317a,a3318a,a3319a,a3320a,a3321a,a3322a,a3323a,a3324a,a3325a,a3326a,a3327a,a3328a,a3329a,a3330a,a3331a,a3332a,a3333a,a3334a,a3335a,a3336a,a3337a,a3338a,a3339a,a3340a,a3341a,a3342a,a3343a,a3344a,a3345a,a3346a,a3347a,a3348a,a3349a,a3350a,a3351a,a3352a,a3353a,a3354a,a3355a,a3356a,a3357a,a3358a,a3359a,a3360a,a3361a,a3362a,a3363a,a3364a,a3365a,a3366a,a3367a,a3368a,a3369a,a3370a,a3371a,a3372a,a3373a,a3374a,a3375a,a3376a,a3377a,a3378a,a3379a,a3380a,a3381a,a3382a,a3383a,a3384a,a3385a,a3386a,a3387a,a3388a,a3389a,a3390a,a3391a,a3392a,a3393a,a3394a,a3395a,a3396a,a3397a,a3398a,a3399a,a3400a,a3401a,a3402a,a3403a,a3404a,a3405a,a3406a,a3407a,a3408a,a3409a,a3410a,a3411a,a3412a,a3413a,a3414a,a3415a,a3416a,a3417a,a3418a,a3419a,a3420a,a3421a,a3422a,a3423a,a3424a,a3425a,a3426a,a3427a,a3428a,a3429a,a3430a,a3431a,a3432a,a3433a,a3434a,a3435a,a3436a,a3437a,a3438a,a3439a,a3440a,a3441a,a3442a,a3443a,a3444a,a3445a,a3446a,a3447a,a3448a,a3449a,a3450a,a3451a,a3452a,a3453a,a3454a,a3455a,a3456a,a3457a,a3458a,a3459a,a3460a,a3461a,a3462a,a3463a,a3464a,a3465a,a3466a,a3467a,a3468a,a3469a,a3470a,a3471a,a3472a,a3473a,a3474a,a3475a,a3476a,a3477a,a3478a,a3479a,a3480a,a3481a,a3482a,a3483a,a3484a,a3485a,a3486a,a3487a,a3488a,a3489a,a3490a,a3491a,a3492a,a3493a,a3494a,a3495a,a3496a,a3497a,a3498a,a3499a,a3500a,a3501a,a3502a,a3503a,a3504a,a3505a,a3506a,a3507a,a3508a,a3509a,a3510a,a3511a,a3512a,a3513a,a3514a,a3515a,a3516a,a3517a,a3518a,a3519a,a3520a,a3521a,a3522a,a3523a,a3524a,a3525a,a3526a,a3527a,a3528a,a3529a,a3530a,a3531a,a3532a,a3533a,a3534a,a3535a,a3536a,a3537a,a3538a,a3539a,a3540a,a3541a,a3542a,a3543a,a3544a,a3545a,a3546a,a3547a,a3548a,a3549a,a3550a,a3551a,a3552a,a3553a,a3554a,a3555a,a3556a,a3557a,a3558a,a3559a,a3560a,a3561a,a3562a,a3563a,a3564a,a3565a,a3566a,a3567a,a3568a,a3569a,a3570a,a3571a,a3572a,a3573a,a3574a,a3575a,a3576a,a3577a,a3578a,a3579a,a3580a,a3581a,a3582a,a3583a,a3584a,a3585a,a3586a,a3587a,a3588a,a3589a,a3590a,a3591a,a3592a,a3593a,a3594a,a3595a,a3596a,a3597a,a3598a,a3599a,a3600a,a3601a,a3602a,a3603a,a3604a,a3605a,a3606a,a3607a,a3608a,a3609a,a3610a,a3611a,a3612a,a3613a,a3614a,a3615a,a3616a,a3617a,a3618a,a3619a,a3620a,a3621a,a3622a,a3623a,a3624a,a3625a,a3626a,a3627a,a3628a,a3629a,a3630a,a3631a,a3632a,a3633a,a3634a,a3635a,a3636a,a3637a,a3638a,a3639a,a3640a,a3641a,a3642a,a3643a,a3644a,a3645a,a3646a,a3647a,a3648a,a3649a,a3650a,a3651a,a3652a,a3653a,a3654a,a3655a,a3656a,a3657a,a3658a,a3659a,a3660a,a3661a,a3662a,a3663a,a3664a,a3665a,a3666a,a3667a,a3668a,a3669a,a3670a,a3671a,a3672a,a3673a,a3674a,a3675a,a3676a,a3677a,a3678a,a3679a,a3680a,a3681a,a3682a,a3683a,a3684a,a3685a,a3686a,a3687a,a3688a,a3689a,a3690a,a3691a,a3692a,a3693a,a3694a,a3695a,a3696a,a3697a,a3698a,a3699a,a3700a,a3701a,a3702a,a3703a,a3704a,a3705a,a3706a,a3707a,a3708a,a3709a,a3710a,a3711a,a3712a,a3713a,a3714a,a3715a,a3716a,a3717a,a3718a,a3719a,a3720a,a3721a,a3722a,a3723a,a3724a,a3725a,a3726a,a3727a,a3728a,a3729a,a3730a,a3731a,a3732a,a3733a,a3734a,a3735a,a3736a,a3737a,a3738a,a3739a,a3740a,a3741a,a3742a,a3743a,a3744a,a3745a,a3746a,a3747a,a3748a,a3749a,a3750a,a3751a,a3752a,a3753a,a3754a,a3755a,a3756a,a3757a,a3758a,a3759a,a3760a,a3761a,a3762a,a3763a,a3764a,a3765a,a3766a,a3767a,a3768a,a3769a,a3770a,a3771a,a3772a,a3773a,a3774a,a3775a,a3776a,a3777a,a3778a,a3779a,a3780a,a3781a,a3782a,a3783a,a3784a,a3785a,a3786a,a3787a,a3788a,a3789a,a3790a,a3791a,a3792a,a3793a,a3794a,a3795a,a3796a,a3797a,a3798a,a3799a,a3800a,a3801a,a3802a,a3803a,a3804a,a3805a,a3806a,a3807a,a3808a,a3809a,a3810a,a3811a,a3812a,a3813a,a3814a,a3815a,a3816a,a3817a,a3818a,a3819a,a3820a,a3821a,a3822a,a3823a,a3824a,a3825a,a3826a,a3827a,a3828a,a3829a,a3830a,a3831a,a3832a,a3833a,a3834a,a3835a,a3836a,a3837a,a3838a,a3842a,a3843a,a3846a,a3849a,a3850a,a3851a,a3855a,a3856a,a3859a,a3862a,a3863a,a3864a,a3865a,a3869a,a3870a,a3873a,a3876a,a3877a,a3878a,a3881a,a3884a,a3885a,a3888a,a3891a,a3892a,a3893a,a3894a,a3895a,a3899a,a3900a,a3903a,a3906a,a3907a,a3908a,a3911a,a3914a,a3915a,a3918a,a3921a,a3922a,a3923a,a3924a,a3928a,a3929a,a3932a,a3935a,a3936a,a3937a,a3940a,a3943a,a3944a,a3947a,a3950a,a3951a,a3952a,a3953a,a3954a,a3955a,a3959a,a3960a,a3963a,a3966a,a3967a,a3968a,a3971a,a3974a,a3975a,a3978a,a3981a,a3982a,a3983a,a3984a,a3988a,a3989a,a3992a,a3995a,a3996a,a3997a,a4000a,a4003a,a4004a,a4007a,a4010a,a4011a,a4012a,a4013a,a4014a,a4018a,a4019a,a4022a,a4025a,a4026a,a4027a,a4030a,a4033a,a4034a,a4037a,a4040a,a4041a,a4042a,a4043a,a4047a,a4048a,a4051a,a4054a,a4055a,a4056a,a4059a,a4062a,a4063a,a4066a,a4069a,a4070a,a4071a,a4072a,a4073a,a4074a,a4075a,a4079a,a4080a,a4083a,a4086a,a4087a,a4088a,a4091a,a4094a,a4095a,a4098a,a4101a,a4102a,a4103a,a4104a,a4108a,a4109a,a4112a,a4115a,a4116a,a4117a,a4120a,a4123a,a4124a,a4127a,a4130a,a4131a,a4132a,a4133a,a4134a,a4138a,a4139a,a4142a,a4145a,a4146a,a4147a,a4150a,a4153a,a4154a,a4157a,a4160a,a4161a,a4162a,a4163a,a4167a,a4168a,a4171a,a4174a,a4175a,a4176a,a4179a,a4182a,a4183a,a4186a,a4189a,a4190a,a4191a,a4192a,a4193a,a4194a,a4198a,a4199a,a4202a,a4205a,a4206a,a4207a,a4210a,a4213a,a4214a,a4217a,a4220a,a4221a,a4222a,a4223a,a4227a,a4228a,a4231a,a4234a,a4235a,a4236a,a4239a,a4242a,a4243a,a4246a,a4249a,a4250a,a4251a,a4252a,a4253a,a4257a,a4258a,a4261a,a4264a,a4265a,a4266a,a4269a,a4272a,a4273a,a4276a,a4279a,a4280a,a4281a,a4282a,a4286a,a4287a,a4290a,a4293a,a4294a,a4295a,a4298a,a4301a,a4302a,a4305a,a4308a,a4309a,a4310a,a4311a,a4312a,a4313a,a4314a,a4315a,a4319a,a4320a,a4323a,a4326a,a4327a,a4328a,a4331a,a4334a,a4335a,a4338a,a4341a,a4342a,a4343a,a4344a,a4348a,a4349a,a4352a,a4355a,a4356a,a4357a,a4360a,a4363a,a4364a,a4367a,a4370a,a4371a,a4372a,a4373a,a4374a,a4378a,a4379a,a4382a,a4385a,a4386a,a4387a,a4390a,a4393a,a4394a,a4397a,a4400a,a4401a,a4402a,a4403a,a4407a,a4408a,a4411a,a4414a,a4415a,a4416a,a4419a,a4422a,a4423a,a4426a,a4429a,a4430a,a4431a,a4432a,a4433a,a4434a,a4438a,a4439a,a4442a,a4445a,a4446a,a4447a,a4450a,a4453a,a4454a,a4457a,a4460a,a4461a,a4462a,a4463a,a4467a,a4468a,a4471a,a4474a,a4475a,a4476a,a4479a,a4482a,a4483a,a4486a,a4489a,a4490a,a4491a,a4492a,a4493a,a4497a,a4498a,a4501a,a4504a,a4505a,a4506a,a4509a,a4512a,a4513a,a4516a,a4519a,a4520a,a4521a,a4522a,a4526a,a4527a,a4530a,a4533a,a4534a,a4535a,a4538a,a4541a,a4542a,a4545a,a4548a,a4549a,a4550a,a4551a,a4552a,a4553a,a4554a,a4558a,a4559a,a4562a,a4565a,a4566a,a4567a,a4570a,a4573a,a4574a,a4577a,a4580a,a4581a,a4582a,a4583a,a4587a,a4588a,a4591a,a4594a,a4595a,a4596a,a4599a,a4602a,a4603a,a4606a,a4609a,a4610a,a4611a,a4612a,a4613a,a4617a,a4618a,a4621a,a4624a,a4625a,a4626a,a4629a,a4632a,a4633a,a4636a,a4639a,a4640a,a4641a,a4642a,a4646a,a4647a,a4650a,a4653a,a4654a,a4655a,a4658a,a4661a,a4662a,a4665a,a4668a,a4669a,a4670a,a4671a,a4672a,a4673a,a4677a,a4678a,a4681a,a4684a,a4685a,a4686a,a4689a,a4692a,a4693a,a4696a,a4699a,a4700a,a4701a,a4702a,a4706a,a4707a,a4710a,a4713a,a4714a,a4715a,a4718a,a4721a,a4722a,a4725a,a4728a,a4729a,a4730a,a4731a,a4732a,a4736a,a4737a,a4740a,a4743a,a4744a,a4745a,a4748a,a4751a,a4752a,a4755a,a4758a,a4759a,a4760a,a4761a,a4765a,a4766a,a4769a,a4772a,a4773a,a4774a,a4777a,a4780a,a4781a,a4784a,a4787a,a4788a,a4789a,a4790a,a4791a,a4792a,a4793a,a4794a,a4795a,a4799a,a4800a,a4803a,a4806a,a4807a,a4808a,a4811a,a4814a,a4815a,a4818a,a4821a,a4822a,a4823a,a4824a,a4828a,a4829a,a4832a,a4835a,a4836a,a4837a,a4840a,a4843a,a4844a,a4847a,a4850a,a4851a,a4852a,a4853a,a4854a,a4858a,a4859a,a4862a,a4865a,a4866a,a4867a,a4870a,a4873a,a4874a,a4877a,a4880a,a4881a,a4882a,a4883a,a4887a,a4888a,a4891a,a4894a,a4895a,a4896a,a4899a,a4902a,a4903a,a4906a,a4909a,a4910a,a4911a,a4912a,a4913a,a4914a,a4918a,a4919a,a4922a,a4925a,a4926a,a4927a,a4930a,a4933a,a4934a,a4937a,a4940a,a4941a,a4942a,a4943a,a4947a,a4948a,a4951a,a4954a,a4955a,a4956a,a4959a,a4962a,a4963a,a4966a,a4969a,a4970a,a4971a,a4972a,a4973a,a4977a,a4978a,a4981a,a4984a,a4985a,a4986a,a4989a,a4992a,a4993a,a4996a,a4999a,a5000a,a5001a,a5002a,a5006a,a5007a,a5010a,a5013a,a5014a,a5015a,a5018a,a5021a,a5022a,a5025a,a5028a,a5029a,a5030a,a5031a,a5032a,a5033a,a5034a,a5038a,a5039a,a5042a,a5045a,a5046a,a5047a,a5050a,a5053a,a5054a,a5057a,a5060a,a5061a,a5062a,a5063a,a5067a,a5068a,a5071a,a5074a,a5075a,a5076a,a5079a,a5082a,a5083a,a5086a,a5089a,a5090a,a5091a,a5092a,a5093a,a5097a,a5098a,a5101a,a5104a,a5105a,a5106a,a5109a,a5112a,a5113a,a5116a,a5119a,a5120a,a5121a,a5122a,a5126a,a5127a,a5130a,a5133a,a5134a,a5135a,a5138a,a5141a,a5142a,a5145a,a5148a,a5149a,a5150a,a5151a,a5152a,a5153a,a5157a,a5158a,a5161a,a5164a,a5165a,a5166a,a5169a,a5172a,a5173a,a5176a,a5179a,a5180a,a5181a,a5182a,a5186a,a5187a,a5190a,a5193a,a5194a,a5195a,a5198a,a5201a,a5202a,a5205a,a5208a,a5209a,a5210a,a5211a,a5212a,a5216a,a5217a,a5220a,a5223a,a5224a,a5225a,a5228a,a5231a,a5232a,a5235a,a5238a,a5239a,a5240a,a5241a,a5245a,a5246a,a5249a,a5252a,a5253a,a5254a,a5257a,a5260a,a5261a,a5264a,a5267a,a5268a,a5269a,a5270a,a5271a,a5272a,a5273a,a5274a,a5278a,a5279a,a5282a,a5285a,a5286a,a5287a,a5290a,a5293a,a5294a,a5297a,a5300a,a5301a,a5302a,a5303a,a5307a,a5308a,a5311a,a5314a,a5315a,a5316a,a5319a,a5322a,a5323a,a5326a,a5329a,a5330a,a5331a,a5332a,a5333a,a5337a,a5338a,a5341a,a5344a,a5345a,a5346a,a5349a,a5352a,a5353a,a5356a,a5359a,a5360a,a5361a,a5362a,a5366a,a5367a,a5370a,a5373a,a5374a,a5375a,a5378a,a5381a,a5382a,a5385a,a5388a,a5389a,a5390a,a5391a,a5392a,a5393a,a5397a,a5398a,a5401a,a5404a,a5405a,a5406a,a5409a,a5412a,a5413a,a5416a,a5419a,a5420a,a5421a,a5422a,a5426a,a5427a,a5430a,a5433a,a5434a,a5435a,a5438a,a5441a,a5442a,a5445a,a5448a,a5449a,a5450a,a5451a,a5452a,a5456a,a5457a,a5460a,a5463a,a5464a,a5465a,a5468a,a5471a,a5472a,a5475a,a5478a,a5479a,a5480a,a5481a,a5485a,a5486a,a5489a,a5492a,a5493a,a5494a,a5497a,a5500a,a5501a,a5504a,a5507a,a5508a,a5509a,a5510a,a5511a,a5512a,a5513a,a5517a,a5518a,a5521a,a5524a,a5525a,a5526a,a5529a,a5532a,a5533a,a5536a,a5539a,a5540a,a5541a,a5542a,a5546a,a5547a,a5550a,a5553a,a5554a,a5555a,a5558a,a5561a,a5562a,a5565a,a5568a,a5569a,a5570a,a5571a,a5572a,a5576a,a5577a,a5580a,a5583a,a5584a,a5585a,a5588a,a5591a,a5592a,a5595a,a5598a,a5599a,a5600a,a5601a,a5605a,a5606a,a5609a,a5612a,a5613a,a5614a,a5617a,a5620a,a5621a,a5624a,a5627a,a5628a,a5629a,a5630a,a5631a,a5632a,a5636a,a5637a,a5640a,a5643a,a5644a,a5645a,a5648a,a5651a,a5652a,a5655a,a5658a,a5659a,a5660a,a5661a,a5665a,a5666a,a5669a,a5672a,a5673a,a5674a,a5677a,a5680a,a5681a,a5684a,a5687a,a5688a,a5689a,a5690a,a5691a,a5695a,a5696a,a5699a,a5702a,a5703a,a5704a,a5707a,a5710a,a5711a,a5714a,a5717a,a5718a,a5719a,a5720a,a5724a,a5725a,a5728a,a5731a,a5732a,a5733a,a5736a,a5739a,a5740a,a5743a,a5746a,a5747a,a5748a,a5749a,a5750a,a5751a,a5752a,a5753a,a5754a,a5755a,a5759a,a5760a,a5763a,a5766a,a5767a,a5768a,a5771a,a5774a,a5775a,a5778a,a5781a,a5782a,a5783a,a5784a,a5788a,a5789a,a5792a,a5795a,a5796a,a5797a,a5800a,a5803a,a5804a,a5807a,a5810a,a5811a,a5812a,a5813a,a5814a,a5818a,a5819a,a5822a,a5825a,a5826a,a5827a,a5830a,a5833a,a5834a,a5837a,a5840a,a5841a,a5842a,a5843a,a5847a,a5848a,a5851a,a5854a,a5855a,a5856a,a5859a,a5862a,a5863a,a5866a,a5869a,a5870a,a5871a,a5872a,a5873a,a5874a,a5878a,a5879a,a5882a,a5885a,a5886a,a5887a,a5890a,a5893a,a5894a,a5897a,a5900a,a5901a,a5902a,a5903a,a5907a,a5908a,a5911a,a5914a,a5915a,a5916a,a5919a,a5922a,a5923a,a5926a,a5929a,a5930a,a5931a,a5932a,a5933a,a5937a,a5938a,a5941a,a5944a,a5945a,a5946a,a5949a,a5952a,a5953a,a5956a,a5959a,a5960a,a5961a,a5962a,a5966a,a5967a,a5970a,a5973a,a5974a,a5975a,a5978a,a5981a,a5982a,a5985a,a5988a,a5989a,a5990a,a5991a,a5992a,a5993a,a5994a,a5998a,a5999a,a6002a,a6005a,a6006a,a6007a,a6010a,a6013a,a6014a,a6017a,a6020a,a6021a,a6022a,a6023a,a6027a,a6028a,a6031a,a6034a,a6035a,a6036a,a6039a,a6042a,a6043a,a6046a,a6049a,a6050a,a6051a,a6052a,a6053a,a6057a,a6058a,a6061a,a6064a,a6065a,a6066a,a6069a,a6072a,a6073a,a6076a,a6079a,a6080a,a6081a,a6082a,a6086a,a6087a,a6090a,a6093a,a6094a,a6095a,a6098a,a6101a,a6102a,a6105a,a6108a,a6109a,a6110a,a6111a,a6112a,a6113a,a6117a,a6118a,a6121a,a6124a,a6125a,a6126a,a6129a,a6132a,a6133a,a6136a,a6139a,a6140a,a6141a,a6142a,a6146a,a6147a,a6150a,a6153a,a6154a,a6155a,a6158a,a6161a,a6162a,a6165a,a6168a,a6169a,a6170a,a6171a,a6172a,a6176a,a6177a,a6180a,a6183a,a6184a,a6185a,a6188a,a6191a,a6192a,a6195a,a6198a,a6199a,a6200a,a6201a,a6205a,a6206a,a6209a,a6212a,a6213a,a6214a,a6217a,a6220a,a6221a,a6224a,a6227a,a6228a,a6229a,a6230a,a6231a,a6232a,a6233a,a6234a,a6238a,a6239a,a6242a,a6245a,a6246a,a6247a,a6250a,a6253a,a6254a,a6257a,a6260a,a6261a,a6262a,a6263a,a6267a,a6268a,a6271a,a6274a,a6275a,a6276a,a6279a,a6282a,a6283a,a6286a,a6289a,a6290a,a6291a,a6292a,a6293a,a6297a,a6298a,a6301a,a6304a,a6305a,a6306a,a6309a,a6312a,a6313a,a6316a,a6319a,a6320a,a6321a,a6322a,a6326a,a6327a,a6330a,a6333a,a6334a,a6335a,a6338a,a6341a,a6342a,a6345a,a6348a,a6349a,a6350a,a6351a,a6352a,a6353a,a6357a,a6358a,a6361a,a6364a,a6365a,a6366a,a6369a,a6372a,a6373a,a6376a,a6379a,a6380a,a6381a,a6382a,a6386a,a6387a,a6390a,a6393a,a6394a,a6395a,a6398a,a6401a,a6402a,a6405a,a6408a,a6409a,a6410a,a6411a,a6412a,a6416a,a6417a,a6420a,a6423a,a6424a,a6425a,a6428a,a6431a,a6432a,a6435a,a6438a,a6439a,a6440a,a6441a,a6445a,a6446a,a6449a,a6452a,a6453a,a6454a,a6457a,a6460a,a6461a,a6464a,a6467a,a6468a,a6469a,a6470a,a6471a,a6472a,a6473a,a6477a,a6478a,a6481a,a6484a,a6485a,a6486a,a6489a,a6492a,a6493a,a6496a,a6499a,a6500a,a6501a,a6502a,a6506a,a6507a,a6510a,a6513a,a6514a,a6515a,a6518a,a6521a,a6522a,a6525a,a6528a,a6529a,a6530a,a6531a,a6532a,a6536a,a6537a,a6540a,a6543a,a6544a,a6545a,a6548a,a6551a,a6552a,a6555a,a6558a,a6559a,a6560a,a6561a,a6565a,a6566a,a6569a,a6572a,a6573a,a6574a,a6577a,a6580a,a6581a,a6584a,a6587a,a6588a,a6589a,a6590a,a6591a,a6592a,a6596a,a6597a,a6600a,a6603a,a6604a,a6605a,a6608a,a6611a,a6612a,a6615a,a6618a,a6619a,a6620a,a6621a,a6625a,a6626a,a6629a,a6632a,a6633a,a6634a,a6637a,a6640a,a6641a,a6644a,a6647a,a6648a,a6649a,a6650a,a6651a,a6655a,a6656a,a6659a,a6662a,a6663a,a6664a,a6667a,a6670a,a6671a,a6674a,a6677a,a6678a,a6679a,a6680a,a6684a,a6685a,a6688a,a6691a,a6692a,a6693a,a6696a,a6699a,a6700a,a6703a,a6706a,a6707a,a6708a,a6709a,a6710a,a6711a,a6712a,a6713a,a6714a,a6718a,a6719a,a6722a,a6725a,a6726a,a6727a,a6730a,a6733a,a6734a,a6737a,a6740a,a6741a,a6742a,a6743a,a6747a,a6748a,a6751a,a6754a,a6755a,a6756a,a6759a,a6762a,a6763a,a6766a,a6769a,a6770a,a6771a,a6772a,a6773a,a6777a,a6778a,a6781a,a6784a,a6785a,a6786a,a6789a,a6792a,a6793a,a6796a,a6799a,a6800a,a6801a,a6802a,a6806a,a6807a,a6810a,a6813a,a6814a,a6815a,a6818a,a6821a,a6822a,a6825a,a6828a,a6829a,a6830a,a6831a,a6832a,a6833a,a6837a,a6838a,a6841a,a6844a,a6845a,a6846a,a6849a,a6852a,a6853a,a6856a,a6859a,a6860a,a6861a,a6862a,a6866a,a6867a,a6870a,a6873a,a6874a,a6875a,a6878a,a6881a,a6882a,a6885a,a6888a,a6889a,a6890a,a6891a,a6892a,a6896a,a6897a,a6900a,a6903a,a6904a,a6905a,a6908a,a6911a,a6912a,a6915a,a6918a,a6919a,a6920a,a6921a,a6925a,a6926a,a6929a,a6932a,a6933a,a6934a,a6937a,a6940a,a6941a,a6944a,a6947a,a6948a,a6949a,a6950a,a6951a,a6952a,a6953a,a6957a,a6958a,a6961a,a6964a,a6965a,a6966a,a6969a,a6972a,a6973a,a6976a,a6979a,a6980a,a6981a,a6982a,a6986a,a6987a,a6990a,a6993a,a6994a,a6995a,a6998a,a7001a,a7002a,a7005a,a7008a,a7009a,a7010a,a7011a,a7012a,a7016a,a7017a,a7020a,a7023a,a7024a,a7025a,a7028a,a7031a,a7032a,a7035a,a7038a,a7039a,a7040a,a7041a,a7045a,a7046a,a7049a,a7052a,a7053a,a7054a,a7057a,a7060a,a7061a,a7064a,a7067a,a7068a,a7069a,a7070a,a7071a,a7072a,a7076a,a7077a,a7080a,a7083a,a7084a,a7085a,a7088a,a7091a,a7092a,a7095a,a7098a,a7099a,a7100a,a7101a,a7105a,a7106a,a7109a,a7112a,a7113a,a7114a,a7117a,a7120a,a7121a,a7124a,a7127a,a7128a,a7129a,a7130a,a7131a,a7135a,a7136a,a7139a,a7142a,a7143a,a7144a,a7147a,a7150a,a7151a,a7154a,a7157a,a7158a,a7159a,a7160a,a7164a,a7165a,a7168a,a7171a,a7172a,a7173a,a7176a,a7179a,a7180a,a7183a,a7186a,a7187a,a7188a,a7189a,a7190a,a7191a,a7192a,a7193a,a7197a,a7198a,a7201a,a7204a,a7205a,a7206a,a7209a,a7212a,a7213a,a7216a,a7219a,a7220a,a7221a,a7222a,a7226a,a7227a,a7230a,a7233a,a7234a,a7235a,a7238a,a7241a,a7242a,a7245a,a7248a,a7249a,a7250a,a7251a,a7252a,a7256a,a7257a,a7260a,a7263a,a7264a,a7265a,a7268a,a7271a,a7272a,a7275a,a7278a,a7279a,a7280a,a7281a,a7285a,a7286a,a7289a,a7292a,a7293a,a7294a,a7297a,a7300a,a7301a,a7304a,a7307a,a7308a,a7309a,a7310a,a7311a,a7312a,a7316a,a7317a,a7320a,a7323a,a7324a,a7325a,a7328a,a7331a,a7332a,a7335a,a7338a,a7339a,a7340a,a7341a,a7345a,a7346a,a7349a,a7352a,a7353a,a7354a,a7357a,a7360a,a7361a,a7364a,a7367a,a7368a,a7369a,a7370a,a7371a,a7375a,a7376a,a7379a,a7382a,a7383a,a7384a,a7387a,a7390a,a7391a,a7394a,a7397a,a7398a,a7399a,a7400a,a7404a,a7405a,a7408a,a7411a,a7412a,a7413a,a7416a,a7419a,a7420a,a7423a,a7426a,a7427a,a7428a,a7429a,a7430a,a7431a,a7432a,a7436a,a7437a,a7440a,a7443a,a7444a,a7445a,a7448a,a7451a,a7452a,a7455a,a7458a,a7459a,a7460a,a7461a,a7465a,a7466a,a7469a,a7472a,a7473a,a7474a,a7477a,a7480a,a7481a,a7484a,a7487a,a7488a,a7489a,a7490a,a7491a,a7495a,a7496a,a7499a,a7502a,a7503a,a7504a,a7507a,a7510a,a7511a,a7514a,a7517a,a7518a,a7519a,a7520a,a7524a,a7525a,a7528a,a7531a,a7532a,a7533a,a7536a,a7539a,a7540a,a7543a,a7546a,a7547a,a7548a,a7549a,a7550a,a7551a,a7555a,a7556a,a7559a,a7562a,a7563a,a7564a,a7567a,a7570a,a7571a,a7574a,a7577a,a7578a,a7579a,a7580a,a7584a,a7585a,a7588a,a7591a,a7592a,a7593a,a7596a,a7599a,a7600a,a7603a,a7606a,a7607a,a7608a,a7609a,a7610a,a7614a,a7615a,a7618a,a7621a,a7622a,a7623a,a7626a,a7629a,a7630a,a7633a,a7636a,a7637a,a7638a,a7639a,a7643a,a7644a,a7647a,a7650a,a7651a,a7652a,a7655a,a7658a,a7659a,a7662a,a7665a,a7666a,a7667a,a7668a,a7669a,a7670a,a7671a,a7672a,a7673a,a7674a,a7675a,a7679a,a7680a,a7683a,a7686a,a7687a,a7688a,a7692a,a7693a,a7696a,a7699a,a7700a,a7701a,a7702a,a7706a,a7707a,a7710a,a7713a,a7714a,a7715a,a7718a,a7721a,a7722a,a7725a,a7728a,a7729a,a7730a,a7731a,a7732a,a7736a,a7737a,a7740a,a7743a,a7744a,a7745a,a7748a,a7751a,a7752a,a7755a,a7758a,a7759a,a7760a,a7761a,a7765a,a7766a,a7769a,a7772a,a7773a,a7774a,a7777a,a7780a,a7781a,a7784a,a7787a,a7788a,a7789a,a7790a,a7791a,a7792a,a7796a,a7797a,a7800a,a7803a,a7804a,a7805a,a7808a,a7811a,a7812a,a7815a,a7818a,a7819a,a7820a,a7821a,a7825a,a7826a,a7829a,a7832a,a7833a,a7834a,a7837a,a7840a,a7841a,a7844a,a7847a,a7848a,a7849a,a7850a,a7851a,a7855a,a7856a,a7859a,a7862a,a7863a,a7864a,a7867a,a7870a,a7871a,a7874a,a7877a,a7878a,a7879a,a7880a,a7884a,a7885a,a7888a,a7891a,a7892a,a7893a,a7896a,a7899a,a7900a,a7903a,a7906a,a7907a,a7908a,a7909a,a7910a,a7911a,a7912a,a7916a,a7917a,a7920a,a7923a,a7924a,a7925a,a7928a,a7931a,a7932a,a7935a,a7938a,a7939a,a7940a,a7941a,a7945a,a7946a,a7949a,a7952a,a7953a,a7954a,a7957a,a7960a,a7961a,a7964a,a7967a,a7968a,a7969a,a7970a,a7971a,a7975a,a7976a,a7979a,a7982a,a7983a,a7984a,a7987a,a7990a,a7991a,a7994a,a7997a,a7998a,a7999a,a8000a,a8004a,a8005a,a8008a,a8011a,a8012a,a8013a,a8016a,a8019a,a8020a,a8023a,a8026a,a8027a,a8028a,a8029a,a8030a,a8031a,a8035a,a8036a,a8039a,a8042a,a8043a,a8044a,a8047a,a8050a,a8051a,a8054a,a8057a,a8058a,a8059a,a8060a,a8064a,a8065a,a8068a,a8071a,a8072a,a8073a,a8076a,a8079a,a8080a,a8083a,a8086a,a8087a,a8088a,a8089a,a8090a,a8094a,a8095a,a8098a,a8101a,a8102a,a8103a,a8106a,a8109a,a8110a,a8113a,a8116a,a8117a,a8118a,a8119a,a8123a,a8124a,a8127a,a8130a,a8131a,a8132a,a8135a,a8138a,a8139a,a8142a,a8145a,a8146a,a8147a,a8148a,a8149a,a8150a,a8151a,a8152a,a8156a,a8157a,a8160a,a8163a,a8164a,a8165a,a8168a,a8171a,a8172a,a8175a,a8178a,a8179a,a8180a,a8181a,a8185a,a8186a,a8189a,a8192a,a8193a,a8194a,a8197a,a8200a,a8201a,a8204a,a8207a,a8208a,a8209a,a8210a,a8211a,a8215a,a8216a,a8219a,a8222a,a8223a,a8224a,a8227a,a8230a,a8231a,a8234a,a8237a,a8238a,a8239a,a8240a,a8244a,a8245a,a8248a,a8251a,a8252a,a8253a,a8256a,a8259a,a8260a,a8263a,a8266a,a8267a,a8268a,a8269a,a8270a,a8271a,a8275a,a8276a,a8279a,a8282a,a8283a,a8284a,a8287a,a8290a,a8291a,a8294a,a8297a,a8298a,a8299a,a8300a,a8304a,a8305a,a8308a,a8311a,a8312a,a8313a,a8316a,a8319a,a8320a,a8323a,a8326a,a8327a,a8328a,a8329a,a8330a,a8334a,a8335a,a8338a,a8341a,a8342a,a8343a,a8346a,a8349a,a8350a,a8353a,a8356a,a8357a,a8358a,a8359a,a8363a,a8364a,a8367a,a8370a,a8371a,a8372a,a8375a,a8378a,a8379a,a8382a,a8385a,a8386a,a8387a,a8388a,a8389a,a8390a,a8391a,a8395a,a8396a,a8399a,a8402a,a8403a,a8404a,a8407a,a8410a,a8411a,a8414a,a8417a,a8418a,a8419a,a8420a,a8424a,a8425a,a8428a,a8431a,a8432a,a8433a,a8436a,a8439a,a8440a,a8443a,a8446a,a8447a,a8448a,a8449a,a8450a,a8454a,a8455a,a8458a,a8461a,a8462a,a8463a,a8466a,a8469a,a8470a,a8473a,a8476a,a8477a,a8478a,a8479a,a8483a,a8484a,a8487a,a8490a,a8491a,a8492a,a8495a,a8498a,a8499a,a8502a,a8505a,a8506a,a8507a,a8508a,a8509a,a8510a,a8514a,a8515a,a8518a,a8521a,a8522a,a8523a,a8526a,a8529a,a8530a,a8533a,a8536a,a8537a,a8538a,a8539a,a8543a,a8544a,a8547a,a8550a,a8551a,a8552a,a8555a,a8558a,a8559a,a8562a,a8565a,a8566a,a8567a,a8568a,a8569a,a8573a,a8574a,a8577a,a8580a,a8581a,a8582a,a8585a,a8588a,a8589a,a8592a,a8595a,a8596a,a8597a,a8598a,a8602a,a8603a,a8606a,a8609a,a8610a,a8611a,a8614a,a8617a,a8618a,a8621a,a8624a,a8625a,a8626a,a8627a,a8628a,a8629a,a8630a,a8631a,a8632a,a8636a,a8637a,a8640a,a8643a,a8644a,a8645a,a8648a,a8651a,a8652a,a8655a,a8658a,a8659a,a8660a,a8661a,a8665a,a8666a,a8669a,a8672a,a8673a,a8674a,a8677a,a8680a,a8681a,a8684a,a8687a,a8688a,a8689a,a8690a,a8691a,a8695a,a8696a,a8699a,a8702a,a8703a,a8704a,a8707a,a8710a,a8711a,a8714a,a8717a,a8718a,a8719a,a8720a,a8724a,a8725a,a8728a,a8731a,a8732a,a8733a,a8736a,a8739a,a8740a,a8743a,a8746a,a8747a,a8748a,a8749a,a8750a,a8751a,a8755a,a8756a,a8759a,a8762a,a8763a,a8764a,a8767a,a8770a,a8771a,a8774a,a8777a,a8778a,a8779a,a8780a,a8784a,a8785a,a8788a,a8791a,a8792a,a8793a,a8796a,a8799a,a8800a,a8803a,a8806a,a8807a,a8808a,a8809a,a8810a,a8814a,a8815a,a8818a,a8821a,a8822a,a8823a,a8826a,a8829a,a8830a,a8833a,a8836a,a8837a,a8838a,a8839a,a8843a,a8844a,a8847a,a8850a,a8851a,a8852a,a8855a,a8858a,a8859a,a8862a,a8865a,a8866a,a8867a,a8868a,a8869a,a8870a,a8871a,a8875a,a8876a,a8879a,a8882a,a8883a,a8884a,a8887a,a8890a,a8891a,a8894a,a8897a,a8898a,a8899a,a8900a,a8904a,a8905a,a8908a,a8911a,a8912a,a8913a,a8916a,a8919a,a8920a,a8923a,a8926a,a8927a,a8928a,a8929a,a8930a,a8934a,a8935a,a8938a,a8941a,a8942a,a8943a,a8946a,a8949a,a8950a,a8953a,a8956a,a8957a,a8958a,a8959a,a8963a,a8964a,a8967a,a8970a,a8971a,a8972a,a8975a,a8978a,a8979a,a8982a,a8985a,a8986a,a8987a,a8988a,a8989a,a8990a,a8994a,a8995a,a8998a,a9001a,a9002a,a9003a,a9006a,a9009a,a9010a,a9013a,a9016a,a9017a,a9018a,a9019a,a9023a,a9024a,a9027a,a9030a,a9031a,a9032a,a9035a,a9038a,a9039a,a9042a,a9045a,a9046a,a9047a,a9048a,a9049a,a9053a,a9054a,a9057a,a9060a,a9061a,a9062a,a9065a,a9068a,a9069a,a9072a,a9075a,a9076a,a9077a,a9078a,a9082a,a9083a,a9086a,a9089a,a9090a,a9091a,a9094a,a9097a,a9098a,a9101a,a9104a,a9105a,a9106a,a9107a,a9108a,a9109a,a9110a,a9111a,a9115a,a9116a,a9119a,a9122a,a9123a,a9124a,a9127a,a9130a,a9131a,a9134a,a9137a,a9138a,a9139a,a9140a,a9144a,a9145a,a9148a,a9151a,a9152a,a9153a,a9156a,a9159a,a9160a,a9163a,a9166a,a9167a,a9168a,a9169a,a9170a,a9174a,a9175a,a9178a,a9181a,a9182a,a9183a,a9186a,a9189a,a9190a,a9193a,a9196a,a9197a,a9198a,a9199a,a9203a,a9204a,a9207a,a9210a,a9211a,a9212a,a9215a,a9218a,a9219a,a9222a,a9225a,a9226a,a9227a,a9228a,a9229a,a9230a,a9234a,a9235a,a9238a,a9241a,a9242a,a9243a,a9246a,a9249a,a9250a,a9253a,a9256a,a9257a,a9258a,a9259a,a9263a,a9264a,a9267a,a9270a,a9271a,a9272a,a9275a,a9278a,a9279a,a9282a,a9285a,a9286a,a9287a,a9288a,a9289a,a9293a,a9294a,a9297a,a9300a,a9301a,a9302a,a9305a,a9308a,a9309a,a9312a,a9315a,a9316a,a9317a,a9318a,a9322a,a9323a,a9326a,a9329a,a9330a,a9331a,a9334a,a9337a,a9338a,a9341a,a9344a,a9345a,a9346a,a9347a,a9348a,a9349a,a9350a,a9354a,a9355a,a9358a,a9361a,a9362a,a9363a,a9366a,a9369a,a9370a,a9373a,a9376a,a9377a,a9378a,a9379a,a9383a,a9384a,a9387a,a9390a,a9391a,a9392a,a9395a,a9398a,a9399a,a9402a,a9405a,a9406a,a9407a,a9408a,a9409a,a9413a,a9414a,a9417a,a9420a,a9421a,a9422a,a9425a,a9428a,a9429a,a9432a,a9435a,a9436a,a9437a,a9438a,a9442a,a9443a,a9446a,a9449a,a9450a,a9451a,a9454a,a9457a,a9458a,a9461a,a9464a,a9465a,a9466a,a9467a,a9468a,a9469a,a9473a,a9474a,a9477a,a9480a,a9481a,a9482a,a9485a,a9488a,a9489a,a9492a,a9495a,a9496a,a9497a,a9498a,a9502a,a9503a,a9506a,a9509a,a9510a,a9511a,a9514a,a9517a,a9518a,a9521a,a9524a,a9525a,a9526a,a9527a,a9528a,a9532a,a9533a,a9536a,a9539a,a9540a,a9541a,a9544a,a9547a,a9548a,a9551a,a9554a,a9555a,a9556a,a9557a,a9561a,a9562a,a9565a,a9568a,a9569a,a9570a,a9573a,a9576a,a9577a,a9580a,a9583a,a9584a,a9585a,a9586a,a9587a,a9588a,a9589a,a9590a,a9591a,a9592a,a9596a,a9597a,a9600a,a9603a,a9604a,a9605a,a9608a,a9611a,a9612a,a9615a,a9618a,a9619a,a9620a,a9621a,a9625a,a9626a,a9629a,a9632a,a9633a,a9634a,a9637a,a9640a,a9641a,a9644a,a9647a,a9648a,a9649a,a9650a,a9651a,a9655a,a9656a,a9659a,a9662a,a9663a,a9664a,a9667a,a9670a,a9671a,a9674a,a9677a,a9678a,a9679a,a9680a,a9684a,a9685a,a9688a,a9691a,a9692a,a9693a,a9696a,a9699a,a9700a,a9703a,a9706a,a9707a,a9708a,a9709a,a9710a,a9711a,a9715a,a9716a,a9719a,a9722a,a9723a,a9724a,a9727a,a9730a,a9731a,a9734a,a9737a,a9738a,a9739a,a9740a,a9744a,a9745a,a9748a,a9751a,a9752a,a9753a,a9756a,a9759a,a9760a,a9763a,a9766a,a9767a,a9768a,a9769a,a9770a,a9774a,a9775a,a9778a,a9781a,a9782a,a9783a,a9786a,a9789a,a9790a,a9793a,a9796a,a9797a,a9798a,a9799a,a9803a,a9804a,a9807a,a9810a,a9811a,a9812a,a9815a,a9818a,a9819a,a9822a,a9825a,a9826a,a9827a,a9828a,a9829a,a9830a,a9831a,a9835a,a9836a,a9839a,a9842a,a9843a,a9844a,a9847a,a9850a,a9851a,a9854a,a9857a,a9858a,a9859a,a9860a,a9864a,a9865a,a9868a,a9871a,a9872a,a9873a,a9876a,a9879a,a9880a,a9883a,a9886a,a9887a,a9888a,a9889a,a9890a,a9894a,a9895a,a9898a,a9901a,a9902a,a9903a,a9906a,a9909a,a9910a,a9913a,a9916a,a9917a,a9918a,a9919a,a9923a,a9924a,a9927a,a9930a,a9931a,a9932a,a9935a,a9938a,a9939a,a9942a,a9945a,a9946a,a9947a,a9948a,a9949a,a9950a,a9954a,a9955a,a9958a,a9961a,a9962a,a9963a,a9966a,a9969a,a9970a,a9973a,a9976a,a9977a,a9978a,a9979a,a9983a,a9984a,a9987a,a9990a,a9991a,a9992a,a9995a,a9998a,a9999a,a10002a,a10005a,a10006a,a10007a,a10008a,a10009a,a10013a,a10014a,a10017a,a10020a,a10021a,a10022a,a10025a,a10028a,a10029a,a10032a,a10035a,a10036a,a10037a,a10038a,a10042a,a10043a,a10046a,a10049a,a10050a,a10051a,a10054a,a10057a,a10058a,a10061a,a10064a,a10065a,a10066a,a10067a,a10068a,a10069a,a10070a,a10071a,a10075a,a10076a,a10079a,a10082a,a10083a,a10084a,a10087a,a10090a,a10091a,a10094a,a10097a,a10098a,a10099a,a10100a,a10104a,a10105a,a10108a,a10111a,a10112a,a10113a,a10116a,a10119a,a10120a,a10123a,a10126a,a10127a,a10128a,a10129a,a10130a,a10134a,a10135a,a10138a,a10141a,a10142a,a10143a,a10146a,a10149a,a10150a,a10153a,a10156a,a10157a,a10158a,a10159a,a10163a,a10164a,a10167a,a10170a,a10171a,a10172a,a10175a,a10178a,a10179a,a10182a,a10185a,a10186a,a10187a,a10188a,a10189a,a10190a,a10194a,a10195a,a10198a,a10201a,a10202a,a10203a,a10206a,a10209a,a10210a,a10213a,a10216a,a10217a,a10218a,a10219a,a10223a,a10224a,a10227a,a10230a,a10231a,a10232a,a10235a,a10238a,a10239a,a10242a,a10245a,a10246a,a10247a,a10248a,a10249a,a10253a,a10254a,a10257a,a10260a,a10261a,a10262a,a10265a,a10268a,a10269a,a10272a,a10275a,a10276a,a10277a,a10278a,a10282a,a10283a,a10286a,a10289a,a10290a,a10291a,a10294a,a10297a,a10298a,a10301a,a10304a,a10305a,a10306a,a10307a,a10308a,a10309a,a10310a,a10314a,a10315a,a10318a,a10321a,a10322a,a10323a,a10326a,a10329a,a10330a,a10333a,a10336a,a10337a,a10338a,a10339a,a10343a,a10344a,a10347a,a10350a,a10351a,a10352a,a10355a,a10358a,a10359a,a10362a,a10365a,a10366a,a10367a,a10368a,a10369a,a10373a,a10374a,a10377a,a10380a,a10381a,a10382a,a10385a,a10388a,a10389a,a10392a,a10395a,a10396a,a10397a,a10398a,a10402a,a10403a,a10406a,a10409a,a10410a,a10411a,a10414a,a10417a,a10418a,a10421a,a10424a,a10425a,a10426a,a10427a,a10428a,a10429a,a10433a,a10434a,a10437a,a10440a,a10441a,a10442a,a10445a,a10448a,a10449a,a10452a,a10455a,a10456a,a10457a,a10458a,a10462a,a10463a,a10466a,a10469a,a10470a,a10471a,a10474a,a10477a,a10478a,a10481a,a10484a,a10485a,a10486a,a10487a,a10488a,a10492a,a10493a,a10496a,a10499a,a10500a,a10501a,a10504a,a10507a,a10508a,a10511a,a10514a,a10515a,a10516a,a10517a,a10521a,a10522a,a10525a,a10528a,a10529a,a10530a,a10533a,a10536a,a10537a,a10540a,a10543a,a10544a,a10545a,a10546a,a10547a,a10548a,a10549a,a10550a,a10551a,a10555a,a10556a,a10559a,a10562a,a10563a,a10564a,a10567a,a10570a,a10571a,a10574a,a10577a,a10578a,a10579a,a10580a,a10584a,a10585a,a10588a,a10591a,a10592a,a10593a,a10596a,a10599a,a10600a,a10603a,a10606a,a10607a,a10608a,a10609a,a10610a,a10614a,a10615a,a10618a,a10621a,a10622a,a10623a,a10626a,a10629a,a10630a,a10633a,a10636a,a10637a,a10638a,a10639a,a10643a,a10644a,a10647a,a10650a,a10651a,a10652a,a10655a,a10658a,a10659a,a10662a,a10665a,a10666a,a10667a,a10668a,a10669a,a10670a,a10674a,a10675a,a10678a,a10681a,a10682a,a10683a,a10686a,a10689a,a10690a,a10693a,a10696a,a10697a,a10698a,a10699a,a10703a,a10704a,a10707a,a10710a,a10711a,a10712a,a10715a,a10718a,a10719a,a10722a,a10725a,a10726a,a10727a,a10728a,a10729a,a10733a,a10734a,a10737a,a10740a,a10741a,a10742a,a10745a,a10748a,a10749a,a10752a,a10755a,a10756a,a10757a,a10758a,a10762a,a10763a,a10766a,a10769a,a10770a,a10771a,a10774a,a10777a,a10778a,a10781a,a10784a,a10785a,a10786a,a10787a,a10788a,a10789a,a10790a,a10794a,a10795a,a10798a,a10801a,a10802a,a10803a,a10806a,a10809a,a10810a,a10813a,a10816a,a10817a,a10818a,a10819a,a10823a,a10824a,a10827a,a10830a,a10831a,a10832a,a10835a,a10838a,a10839a,a10842a,a10845a,a10846a,a10847a,a10848a,a10849a,a10853a,a10854a,a10857a,a10860a,a10861a,a10862a,a10865a,a10868a,a10869a,a10872a,a10875a,a10876a,a10877a,a10878a,a10882a,a10883a,a10886a,a10889a,a10890a,a10891a,a10894a,a10897a,a10898a,a10901a,a10904a,a10905a,a10906a,a10907a,a10908a,a10909a,a10913a,a10914a,a10917a,a10920a,a10921a,a10922a,a10925a,a10928a,a10929a,a10932a,a10935a,a10936a,a10937a,a10938a,a10942a,a10943a,a10946a,a10949a,a10950a,a10951a,a10954a,a10957a,a10958a,a10961a,a10964a,a10965a,a10966a,a10967a,a10968a,a10972a,a10973a,a10976a,a10979a,a10980a,a10981a,a10984a,a10987a,a10988a,a10991a,a10994a,a10995a,a10996a,a10997a,a11001a,a11002a,a11005a,a11008a,a11009a,a11010a,a11013a,a11016a,a11017a,a11020a,a11023a,a11024a,a11025a,a11026a,a11027a,a11028a,a11029a,a11030a,a11034a,a11035a,a11038a,a11041a,a11042a,a11043a,a11046a,a11049a,a11050a,a11053a,a11056a,a11057a,a11058a,a11059a,a11063a,a11064a,a11067a,a11070a,a11071a,a11072a,a11075a,a11078a,a11079a,a11082a,a11085a,a11086a,a11087a,a11088a,a11089a,a11093a,a11094a,a11097a,a11100a,a11101a,a11102a,a11105a,a11108a,a11109a,a11112a,a11115a,a11116a,a11117a,a11118a,a11122a,a11123a,a11126a,a11129a,a11130a,a11131a,a11134a,a11137a,a11138a,a11141a,a11144a,a11145a,a11146a,a11147a,a11148a,a11149a,a11153a,a11154a,a11157a,a11160a,a11161a,a11162a,a11165a,a11168a,a11169a,a11172a,a11175a,a11176a,a11177a,a11178a,a11182a,a11183a,a11186a,a11189a,a11190a,a11191a,a11194a,a11197a,a11198a,a11201a,a11204a,a11205a,a11206a,a11207a,a11208a,a11212a,a11213a,a11216a,a11219a,a11220a,a11221a,a11224a,a11227a,a11228a,a11231a,a11234a,a11235a,a11236a,a11237a,a11241a,a11242a,a11245a,a11248a,a11249a,a11250a,a11253a,a11256a,a11257a,a11260a,a11263a,a11264a,a11265a,a11266a,a11267a,a11268a,a11269a,a11273a,a11274a,a11277a,a11280a,a11281a,a11282a,a11285a,a11288a,a11289a,a11292a,a11295a,a11296a,a11297a,a11298a,a11302a,a11303a,a11306a,a11309a,a11310a,a11311a,a11314a,a11317a,a11318a,a11321a,a11324a,a11325a,a11326a,a11327a,a11328a,a11332a,a11333a,a11336a,a11339a,a11340a,a11341a,a11344a,a11347a,a11348a,a11351a,a11354a,a11355a,a11356a,a11357a,a11361a,a11362a,a11365a,a11368a,a11369a,a11370a,a11373a,a11376a,a11377a,a11380a,a11383a,a11384a,a11385a,a11386a,a11387a,a11388a,a11392a,a11393a,a11396a,a11399a,a11400a,a11401a,a11404a,a11407a,a11408a,a11411a,a11414a,a11415a,a11416a,a11417a,a11421a,a11422a,a11425a,a11428a,a11429a,a11430a,a11433a,a11436a,a11437a,a11440a,a11443a,a11444a,a11445a,a11446a,a11447a,a11451a,a11452a,a11455a,a11458a,a11459a,a11460a,a11463a,a11466a,a11467a,a11470a,a11473a,a11474a,a11475a,a11476a,a11480a,a11481a,a11484a,a11487a,a11488a,a11489a,a11492a,a11495a,a11496a,a11499a,a11502a,a11503a,a11504a,a11505a,a11506a,a11507a,a11508a,a11509a,a11510a,a11511a,a11512a,a11515a,a11518a,a11519a,a11522a,a11525a,a11526a,a11529a,a11532a,a11533a,a11536a,a11539a,a11540a,a11543a,a11546a,a11547a,a11550a,a11553a,a11554a,a11557a,a11560a,a11561a,a11564a,a11567a,a11568a,a11571a,a11574a,a11575a,a11578a,a11581a,a11582a,a11585a,a11588a,a11589a,a11592a,a11595a,a11596a,a11599a,a11602a,a11603a,a11606a,a11609a,a11610a,a11613a,a11616a,a11617a,a11620a,a11623a,a11624a,a11627a,a11630a,a11631a,a11634a,a11637a,a11638a,a11641a,a11644a,a11645a,a11648a,a11651a,a11652a,a11655a,a11658a,a11659a,a11662a,a11665a,a11666a,a11669a,a11672a,a11673a,a11676a,a11679a,a11680a,a11683a,a11686a,a11687a,a11690a,a11693a,a11694a,a11697a,a11700a,a11701a,a11704a,a11707a,a11708a,a11711a,a11714a,a11715a,a11718a,a11721a,a11722a,a11725a,a11728a,a11729a,a11732a,a11735a,a11736a,a11739a,a11742a,a11743a,a11746a,a11749a,a11750a,a11753a,a11756a,a11757a,a11760a,a11763a,a11764a,a11767a,a11770a,a11771a,a11774a,a11777a,a11778a,a11781a,a11784a,a11785a,a11788a,a11791a,a11792a,a11795a,a11798a,a11799a,a11802a,a11805a,a11806a,a11809a,a11812a,a11813a,a11816a,a11819a,a11820a,a11823a,a11826a,a11827a,a11830a,a11833a,a11834a,a11837a,a11840a,a11841a,a11844a,a11847a,a11848a,a11851a,a11854a,a11855a,a11858a,a11861a,a11862a,a11865a,a11868a,a11869a,a11872a,a11875a,a11876a,a11879a,a11882a,a11883a,a11886a,a11889a,a11890a,a11893a,a11896a,a11897a,a11900a,a11903a,a11904a,a11907a,a11910a,a11911a,a11914a,a11917a,a11918a,a11921a,a11924a,a11925a,a11928a,a11931a,a11932a,a11935a,a11938a,a11939a,a11942a,a11945a,a11946a,a11949a,a11952a,a11953a,a11956a,a11959a,a11960a,a11963a,a11966a,a11967a,a11970a,a11974a,a11975a,a11976a,a11979a,a11982a,a11983a,a11986a,a11990a,a11991a,a11992a,a11995a,a11998a,a11999a,a12002a,a12006a,a12007a,a12008a,a12011a,a12014a,a12015a,a12018a,a12022a,a12023a,a12024a,a12027a,a12030a,a12031a,a12034a,a12038a,a12039a,a12040a,a12043a,a12046a,a12047a,a12050a,a12054a,a12055a,a12056a,a12059a,a12062a,a12063a,a12066a,a12070a,a12071a,a12072a,a12075a,a12078a,a12079a,a12082a,a12086a,a12087a,a12088a,a12091a,a12094a,a12095a,a12098a,a12102a,a12103a,a12104a,a12107a,a12110a,a12111a,a12114a,a12118a,a12119a,a12120a,a12123a,a12126a,a12127a,a12130a,a12134a,a12135a,a12136a,a12139a,a12142a,a12143a,a12146a,a12150a,a12151a,a12152a,a12155a,a12158a,a12159a,a12162a,a12166a,a12167a,a12168a,a12171a,a12174a,a12175a,a12178a,a12182a,a12183a,a12184a,a12187a,a12190a,a12191a,a12194a,a12198a,a12199a,a12200a,a12203a,a12206a,a12207a,a12210a,a12214a,a12215a,a12216a,a12219a,a12222a,a12223a,a12226a,a12230a,a12231a,a12232a,a12235a,a12238a,a12239a,a12242a,a12246a,a12247a,a12248a,a12251a,a12254a,a12255a,a12258a,a12262a,a12263a,a12264a,a12267a,a12270a,a12271a,a12274a,a12278a,a12279a,a12280a,a12283a,a12286a,a12287a,a12290a,a12294a,a12295a,a12296a,a12299a,a12302a,a12303a,a12306a,a12310a,a12311a,a12312a,a12315a,a12318a,a12319a,a12322a,a12326a,a12327a,a12328a,a12331a,a12334a,a12335a,a12338a,a12342a,a12343a,a12344a,a12347a,a12351a,a12352a,a12353a,a12356a,a12360a,a12361a,a12362a,a12365a,a12369a,a12370a,a12371a,a12374a,a12378a,a12379a,a12380a,a12383a,a12387a,a12388a,a12389a,a12392a,a12396a,a12397a,a12398a,a12401a,a12405a,a12406a,a12407a,a12410a,a12414a,a12415a,a12416a,a12419a,a12423a,a12424a,a12425a,a12428a,a12432a,a12433a,a12434a,a12437a,a12441a,a12442a,a12443a,a12446a,a12450a,a12451a,a12452a,a12455a,a12459a,a12460a,a12461a,a12464a,a12468a,a12469a,a12470a,a12473a,a12477a,a12478a,a12479a,a12482a,a12486a,a12487a,a12488a,a12491a,a12495a,a12496a,a12497a,a12500a,a12504a,a12505a,a12506a,a12509a,a12513a,a12514a,a12515a,a12518a,a12522a,a12523a,a12524a,a12527a,a12531a,a12532a,a12533a,a12536a,a12540a,a12541a,a12542a,a12545a,a12549a,a12550a,a12551a,a12554a,a12558a,a12559a,a12560a,a12563a,a12567a,a12568a,a12569a,a12572a,a12576a,a12577a,a12578a,a12581a,a12585a,a12586a,a12587a,a12590a,a12594a,a12595a,a12596a,a12599a,a12603a,a12604a,a12605a,a12608a,a12612a,a12613a,a12614a,a12617a,a12621a,a12622a,a12623a,a12626a,a12630a,a12631a,a12632a,a12635a,a12639a,a12640a,a12641a,a12644a,a12648a,a12649a,a12650a,a12653a,a12657a,a12658a,a12659a,a12662a,a12666a,a12667a,a12668a,a12671a,a12675a,a12676a,a12677a,a12680a,a12684a,a12685a,a12686a,a12689a,a12693a,a12694a,a12695a,a12698a,a12702a,a12703a,a12704a,a12707a,a12711a,a12712a,a12713a,a12716a,a12720a,a12721a,a12722a,a12725a,a12729a,a12730a,a12731a,a12734a,a12738a,a12739a,a12740a,a12743a,a12747a,a12748a,a12749a,a12752a,a12756a,a12757a,a12758a,a12761a,a12765a,a12766a,a12767a,a12770a,a12774a,a12775a,a12776a,a12779a,a12783a,a12784a,a12785a,a12788a,a12792a,a12793a,a12794a,a12797a,a12801a,a12802a,a12803a,a12806a,a12810a,a12811a,a12812a,a12815a,a12819a,a12820a,a12821a,a12824a,a12828a,a12829a,a12830a,a12833a,a12837a,a12838a,a12839a,a12842a,a12846a,a12847a,a12848a,a12851a,a12855a,a12856a,a12857a,a12860a,a12864a,a12865a,a12866a,a12869a,a12873a,a12874a,a12875a,a12878a,a12882a,a12883a,a12884a,a12887a,a12891a,a12892a,a12893a,a12896a,a12900a,a12901a,a12902a,a12905a,a12909a,a12910a,a12911a,a12914a,a12918a,a12919a,a12920a,a12923a,a12927a,a12928a,a12929a,a12932a,a12936a,a12937a,a12938a,a12941a,a12945a,a12946a,a12947a,a12950a,a12954a,a12955a,a12956a,a12959a,a12963a,a12964a,a12965a,a12968a,a12972a,a12973a,a12974a,a12977a,a12981a,a12982a,a12983a,a12986a,a12990a,a12991a,a12992a,a12995a,a12999a,a13000a,a13001a,a13004a,a13008a,a13009a,a13010a,a13013a,a13017a,a13018a,a13019a,a13022a,a13026a,a13027a,a13028a,a13031a,a13035a,a13036a,a13037a,a13040a,a13044a,a13045a,a13046a,a13049a,a13053a,a13054a,a13055a,a13058a,a13062a,a13063a,a13064a,a13067a,a13071a,a13072a,a13073a,a13076a,a13080a,a13081a,a13082a,a13085a,a13089a,a13090a,a13091a,a13094a,a13098a,a13099a,a13100a,a13103a,a13107a,a13108a,a13109a,a13112a,a13116a,a13117a,a13118a,a13121a,a13125a,a13126a,a13127a,a13130a,a13134a,a13135a,a13136a,a13139a,a13143a,a13144a,a13145a,a13148a,a13152a,a13153a,a13154a,a13157a,a13161a,a13162a,a13163a,a13166a,a13170a,a13171a,a13172a,a13175a,a13179a,a13180a,a13181a,a13184a,a13188a,a13189a,a13190a,a13193a,a13197a,a13198a,a13199a,a13202a,a13206a,a13207a,a13208a,a13211a,a13215a,a13216a,a13217a,a13220a,a13224a,a13225a,a13226a,a13229a,a13233a,a13234a,a13235a,a13238a,a13242a,a13243a,a13244a,a13247a,a13251a,a13252a,a13253a,a13256a,a13260a,a13261a,a13262a,a13265a,a13269a,a13270a,a13271a,a13274a,a13278a,a13279a,a13280a,a13283a,a13287a,a13288a,a13289a,a13292a,a13296a,a13297a,a13298a,a13301a,a13305a,a13306a,a13307a,a13310a,a13314a,a13315a,a13316a,a13319a,a13323a,a13324a,a13325a,a13328a,a13332a,a13333a,a13334a,a13337a,a13341a,a13342a,a13343a,a13346a,a13350a,a13351a,a13352a,a13355a,a13359a,a13360a,a13361a,a13364a,a13368a,a13369a,a13370a,a13373a,a13377a,a13378a,a13379a,a13382a,a13386a,a13387a,a13388a,a13391a,a13395a,a13396a,a13397a,a13400a,a13404a,a13405a,a13406a,a13409a,a13413a,a13414a,a13415a,a13418a,a13422a,a13423a,a13424a,a13427a,a13431a,a13432a,a13433a,a13436a,a13440a,a13441a,a13442a,a13445a,a13449a,a13450a,a13451a,a13454a,a13458a,a13459a,a13460a,a13463a,a13467a,a13468a,a13469a,a13472a,a13476a,a13477a,a13478a,a13481a,a13485a,a13486a,a13487a,a13490a,a13494a,a13495a,a13496a,a13499a,a13503a,a13504a,a13505a,a13508a,a13512a,a13513a,a13514a,a13517a,a13521a,a13522a,a13523a,a13526a,a13530a,a13531a,a13532a,a13535a,a13539a,a13540a,a13541a,a13544a,a13548a,a13549a,a13550a,a13553a,a13557a,a13558a,a13559a,a13562a,a13566a,a13567a,a13568a,a13571a,a13575a,a13576a,a13577a,a13580a,a13584a,a13585a,a13586a,a13589a,a13593a,a13594a,a13595a,a13598a,a13602a,a13603a,a13604a,a13607a,a13611a,a13612a,a13613a,a13616a,a13620a,a13621a,a13622a,a13625a,a13629a,a13630a,a13631a,a13634a,a13638a,a13639a,a13640a,a13643a,a13647a,a13648a,a13649a,a13652a,a13656a,a13657a,a13658a,a13661a,a13665a,a13666a,a13667a,a13670a,a13674a,a13675a,a13676a,a13679a,a13683a,a13684a,a13685a,a13688a,a13692a,a13693a,a13694a,a13697a,a13701a,a13702a,a13703a,a13706a,a13710a,a13711a,a13712a,a13715a,a13719a,a13720a,a13721a,a13724a,a13728a,a13729a,a13730a,a13733a,a13737a,a13738a,a13739a,a13742a,a13746a,a13747a,a13748a,a13751a,a13755a,a13756a,a13757a,a13760a,a13764a,a13765a,a13766a,a13769a,a13773a,a13774a,a13775a,a13778a,a13782a,a13783a,a13784a,a13787a,a13791a,a13792a,a13793a,a13796a,a13800a,a13801a,a13802a,a13805a,a13809a,a13810a,a13811a,a13814a,a13818a,a13819a,a13820a,a13823a,a13827a,a13828a,a13829a,a13832a,a13836a,a13837a,a13838a,a13841a,a13845a,a13846a,a13847a,a13850a,a13854a,a13855a,a13856a,a13859a,a13863a,a13864a,a13865a,a13868a,a13872a,a13873a,a13874a,a13877a,a13881a,a13882a,a13883a,a13886a,a13890a,a13891a,a13892a,a13895a,a13899a,a13900a,a13901a,a13904a,a13908a,a13909a,a13910a,a13913a,a13917a,a13918a,a13919a,a13922a,a13926a,a13927a,a13928a,a13931a,a13935a,a13936a,a13937a,a13940a,a13944a,a13945a,a13946a,a13949a,a13953a,a13954a,a13955a,a13958a,a13962a,a13963a,a13964a,a13967a,a13971a,a13972a,a13973a,a13976a,a13980a,a13981a,a13982a,a13985a,a13989a,a13990a,a13991a,a13994a,a13998a,a13999a,a14000a,a14003a,a14007a,a14008a,a14009a,a14012a,a14016a,a14017a,a14018a,a14021a,a14025a,a14026a,a14027a,a14030a,a14034a,a14035a,a14036a,a14039a,a14043a,a14044a,a14045a,a14048a,a14052a,a14053a,a14054a,a14057a,a14061a,a14062a,a14063a,a14066a,a14070a,a14071a,a14072a,a14075a,a14079a,a14080a,a14081a,a14084a,a14088a,a14089a,a14090a,a14093a,a14097a,a14098a,a14099a,a14102a,a14106a,a14107a,a14108a,a14111a,a14115a,a14116a,a14117a,a14120a,a14124a,a14125a,a14126a,a14129a,a14133a,a14134a,a14135a,a14138a,a14142a,a14143a,a14144a,a14147a,a14151a,a14152a,a14153a,a14156a,a14160a,a14161a,a14162a,a14165a,a14169a,a14170a,a14171a,a14174a,a14178a,a14179a,a14180a,a14183a,a14187a,a14188a,a14189a,a14192a,a14196a,a14197a,a14198a,a14201a,a14205a,a14206a,a14207a,a14210a,a14214a,a14215a,a14216a,a14219a,a14223a,a14224a,a14225a,a14228a,a14232a,a14233a,a14234a,a14237a,a14241a,a14242a,a14243a,a14246a,a14250a,a14251a,a14252a,a14255a,a14259a,a14260a,a14261a,a14264a,a14268a,a14269a,a14270a,a14273a,a14277a,a14278a,a14279a,a14282a,a14286a,a14287a,a14288a,a14291a,a14295a,a14296a,a14297a,a14300a,a14304a,a14305a,a14306a,a14309a,a14313a,a14314a,a14315a,a14318a,a14322a,a14323a,a14324a,a14327a,a14331a,a14332a,a14333a,a14336a,a14340a,a14341a,a14342a,a14345a,a14349a,a14350a,a14351a,a14354a,a14358a,a14359a,a14360a,a14363a,a14367a,a14368a,a14369a,a14372a,a14376a,a14377a,a14378a,a14381a,a14385a,a14386a,a14387a,a14390a,a14394a,a14395a,a14396a,a14399a,a14403a,a14404a,a14405a,a14408a,a14412a,a14413a,a14414a,a14417a,a14421a,a14422a,a14423a,a14426a,a14430a,a14431a,a14432a,a14435a,a14439a,a14440a,a14441a,a14444a,a14448a,a14449a,a14450a,a14453a,a14457a,a14458a,a14459a,a14462a,a14466a,a14467a,a14468a,a14471a,a14475a,a14476a,a14477a,a14480a,a14484a,a14485a,a14486a,a14489a,a14493a,a14494a,a14495a,a14498a,a14502a,a14503a,a14504a,a14507a,a14511a,a14512a,a14513a,a14516a,a14520a,a14521a,a14522a,a14525a,a14529a,a14530a,a14531a,a14534a,a14538a,a14539a,a14540a,a14543a,a14547a,a14548a,a14549a,a14552a,a14556a,a14557a,a14558a,a14561a,a14565a,a14566a,a14567a,a14570a,a14574a,a14575a,a14576a,a14579a,a14583a,a14584a,a14585a,a14588a,a14592a,a14593a,a14594a,a14597a,a14601a,a14602a,a14603a,a14606a,a14610a,a14611a,a14612a,a14615a,a14619a,a14620a,a14621a,a14624a,a14628a,a14629a,a14630a,a14633a,a14637a,a14638a,a14639a,a14642a,a14646a,a14647a,a14648a,a14651a,a14655a,a14656a,a14657a,a14660a,a14664a,a14665a,a14666a,a14669a,a14673a,a14674a,a14675a,a14678a,a14682a,a14683a,a14684a,a14687a,a14691a,a14692a,a14693a,a14696a,a14700a,a14701a,a14702a,a14705a,a14709a,a14710a,a14711a,a14714a,a14718a,a14719a,a14720a,a14723a,a14727a,a14728a,a14729a,a14732a,a14736a,a14737a,a14738a,a14741a,a14745a,a14746a,a14747a,a14750a,a14754a,a14755a,a14756a,a14759a,a14763a,a14764a,a14765a,a14768a,a14772a,a14773a,a14774a,a14777a,a14781a,a14782a,a14783a,a14786a,a14790a,a14791a,a14792a,a14795a,a14799a,a14800a,a14801a,a14804a,a14808a,a14809a,a14810a,a14813a,a14817a,a14818a,a14819a,a14822a,a14826a,a14827a,a14828a,a14831a,a14835a,a14836a,a14837a,a14840a,a14844a,a14845a,a14846a,a14849a,a14853a,a14854a,a14855a,a14858a,a14862a,a14863a,a14864a,a14867a,a14871a,a14872a,a14873a,a14876a,a14880a,a14881a,a14882a,a14885a,a14889a,a14890a,a14891a,a14894a,a14898a,a14899a,a14900a,a14903a,a14907a,a14908a,a14909a,a14912a,a14916a,a14917a,a14918a,a14921a,a14925a,a14926a,a14927a,a14930a,a14934a,a14935a,a14936a,a14939a,a14943a,a14944a,a14945a,a14948a,a14952a,a14953a,a14954a,a14957a,a14961a,a14962a,a14963a,a14966a,a14970a,a14971a,a14972a,a14975a,a14979a,a14980a,a14981a,a14984a,a14988a,a14989a,a14990a,a14993a,a14997a,a14998a,a14999a,a15002a,a15006a,a15007a,a15008a,a15011a,a15015a,a15016a,a15017a,a15020a,a15024a,a15025a,a15026a,a15029a,a15033a,a15034a,a15035a,a15038a,a15042a,a15043a,a15044a,a15047a,a15051a,a15052a,a15053a,a15056a,a15060a,a15061a,a15062a,a15065a,a15069a,a15070a,a15071a,a15074a,a15078a,a15079a,a15080a,a15083a,a15087a,a15088a,a15089a,a15092a,a15096a,a15097a,a15098a,a15101a,a15105a,a15106a,a15107a,a15110a,a15114a,a15115a,a15116a,a15119a,a15123a,a15124a,a15125a,a15128a,a15132a,a15133a,a15134a,a15137a,a15141a,a15142a,a15143a,a15146a,a15150a,a15151a,a15152a,a15155a,a15159a,a15160a,a15161a,a15164a,a15168a,a15169a,a15170a,a15173a,a15177a,a15178a,a15179a,a15182a,a15186a,a15187a,a15188a,a15191a,a15195a,a15196a,a15197a,a15200a,a15204a,a15205a,a15206a,a15209a,a15213a,a15214a,a15215a,a15218a,a15222a,a15223a,a15224a,a15227a,a15231a,a15232a,a15233a,a15236a,a15240a,a15241a,a15242a,a15245a,a15249a,a15250a,a15251a,a15254a,a15258a,a15259a,a15260a,a15263a,a15267a,a15268a,a15269a,a15272a,a15276a,a15277a,a15278a,a15281a,a15285a,a15286a,a15287a,a15290a,a15294a,a15295a,a15296a,a15299a,a15303a,a15304a,a15305a,a15308a,a15312a,a15313a,a15314a,a15317a,a15321a,a15322a,a15323a,a15326a,a15330a,a15331a,a15332a,a15335a,a15339a,a15340a,a15341a,a15344a,a15348a,a15349a,a15350a,a15353a,a15357a,a15358a,a15359a,a15362a,a15366a,a15367a,a15368a,a15371a,a15375a,a15376a,a15377a,a15380a,a15384a,a15385a,a15386a,a15389a,a15393a,a15394a,a15395a,a15398a,a15402a,a15403a,a15404a,a15407a,a15411a,a15412a,a15413a,a15416a,a15420a,a15421a,a15422a,a15425a,a15429a,a15430a,a15431a,a15434a,a15438a,a15439a,a15440a,a15443a,a15447a,a15448a,a15449a,a15452a,a15456a,a15457a,a15458a,a15461a,a15465a,a15466a,a15467a,a15470a,a15474a,a15475a,a15476a,a15479a,a15483a,a15484a,a15485a,a15488a,a15492a,a15493a,a15494a,a15497a,a15501a,a15502a,a15503a,a15506a,a15510a,a15511a,a15512a,a15515a,a15519a,a15520a,a15521a,a15524a,a15528a,a15529a,a15530a,a15533a,a15537a,a15538a,a15539a,a15542a,a15546a,a15547a,a15548a,a15551a,a15555a,a15556a,a15557a,a15560a,a15564a,a15565a,a15566a,a15569a,a15573a,a15574a,a15575a,a15578a,a15582a,a15583a,a15584a,a15587a,a15591a,a15592a,a15593a,a15596a,a15600a,a15601a,a15602a,a15605a,a15609a,a15610a,a15611a,a15614a,a15618a,a15619a,a15620a,a15623a,a15627a,a15628a,a15629a,a15632a,a15636a,a15637a,a15638a,a15641a,a15645a,a15646a,a15647a,a15650a,a15654a,a15655a,a15656a,a15659a,a15663a,a15664a,a15665a,a15668a,a15672a,a15673a,a15674a,a15677a,a15681a,a15682a,a15683a,a15686a,a15690a,a15691a,a15692a,a15695a,a15699a,a15700a,a15701a,a15704a,a15708a,a15709a,a15710a,a15713a,a15717a,a15718a,a15719a,a15722a,a15726a,a15727a,a15728a,a15731a,a15735a,a15736a,a15737a,a15740a,a15744a,a15745a,a15746a,a15749a,a15753a,a15754a,a15755a,a15758a,a15762a,a15763a,a15764a,a15767a,a15771a,a15772a,a15773a,a15776a,a15780a,a15781a,a15782a,a15785a,a15789a,a15790a,a15791a,a15794a,a15798a,a15799a,a15800a,a15803a,a15807a,a15808a,a15809a,a15812a,a15816a,a15817a,a15818a,a15821a,a15825a,a15826a,a15827a,a15830a,a15834a,a15835a,a15836a,a15839a,a15843a,a15844a,a15845a,a15848a,a15852a,a15853a,a15854a,a15857a,a15861a,a15862a,a15863a,a15866a,a15870a,a15871a,a15872a,a15875a,a15879a,a15880a,a15881a,a15884a,a15888a,a15889a,a15890a,a15893a,a15897a,a15898a,a15899a,a15902a,a15906a,a15907a,a15908a,a15911a,a15915a,a15916a,a15917a,a15920a,a15924a,a15925a,a15926a,a15929a,a15933a,a15934a,a15935a,a15938a,a15942a,a15943a,a15944a,a15947a,a15951a,a15952a,a15953a,a15956a,a15960a,a15961a,a15962a,a15965a,a15969a,a15970a,a15971a,a15974a,a15978a,a15979a,a15980a,a15983a,a15987a,a15988a,a15989a,a15992a,a15996a,a15997a,a15998a,a16001a,a16005a,a16006a,a16007a,a16010a,a16014a,a16015a,a16016a,a16019a,a16023a,a16024a,a16025a,a16028a,a16032a,a16033a,a16034a,a16037a,a16041a,a16042a,a16043a,a16046a,a16050a,a16051a,a16052a,a16055a,a16059a,a16060a,a16061a,a16064a,a16068a,a16069a,a16070a,a16073a,a16077a,a16078a,a16079a,a16082a,a16086a,a16087a,a16088a,a16091a,a16095a,a16096a,a16097a,a16100a,a16104a,a16105a,a16106a,a16109a,a16113a,a16114a,a16115a,a16118a,a16122a,a16123a,a16124a,a16127a,a16131a,a16132a,a16133a,a16136a,a16140a,a16141a,a16142a,a16145a,a16149a,a16150a,a16151a,a16154a,a16158a,a16159a,a16160a,a16163a,a16167a,a16168a,a16169a,a16172a,a16176a,a16177a,a16178a,a16181a,a16185a,a16186a,a16187a,a16190a,a16194a,a16195a,a16196a,a16199a,a16203a,a16204a,a16205a,a16208a,a16212a,a16213a,a16214a,a16217a,a16221a,a16222a,a16223a,a16226a,a16230a,a16231a,a16232a,a16235a,a16239a,a16240a,a16241a,a16244a,a16248a,a16249a,a16250a,a16253a,a16257a,a16258a,a16259a,a16262a,a16266a,a16267a,a16268a,a16271a,a16275a,a16276a,a16277a,a16280a,a16284a,a16285a,a16286a,a16289a,a16293a,a16294a,a16295a,a16298a,a16302a,a16303a,a16304a,a16307a,a16311a,a16312a,a16313a,a16316a,a16320a,a16321a,a16322a,a16325a,a16329a,a16330a,a16331a,a16334a,a16338a,a16339a,a16340a,a16343a,a16347a,a16348a,a16349a,a16352a,a16356a,a16357a,a16358a,a16361a,a16365a,a16366a,a16367a,a16370a,a16374a,a16375a,a16376a,a16379a,a16383a,a16384a,a16385a,a16388a,a16392a,a16393a,a16394a,a16397a,a16401a,a16402a,a16403a,a16406a,a16410a,a16411a,a16412a,a16415a,a16419a,a16420a,a16421a,a16424a,a16428a,a16429a,a16430a,a16433a,a16437a,a16438a,a16439a,a16442a,a16446a,a16447a,a16448a,a16451a,a16455a,a16456a,a16457a,a16460a,a16464a,a16465a,a16466a,a16469a,a16473a,a16474a,a16475a,a16478a,a16482a,a16483a,a16484a,a16487a,a16491a,a16492a,a16493a,a16496a,a16500a,a16501a,a16502a,a16505a,a16509a,a16510a,a16511a,a16514a,a16518a,a16519a,a16520a,a16523a,a16527a,a16528a,a16529a,a16532a,a16536a,a16537a,a16538a,a16541a,a16545a,a16546a,a16547a,a16550a,a16554a,a16555a,a16556a,a16559a,a16563a,a16564a,a16565a,a16568a,a16572a,a16573a,a16574a,a16577a,a16581a,a16582a,a16583a,a16586a,a16590a,a16591a,a16592a,a16595a,a16599a,a16600a,a16601a,a16604a,a16608a,a16609a,a16610a,a16613a,a16617a,a16618a,a16619a,a16622a,a16626a,a16627a,a16628a,a16631a,a16635a,a16636a,a16637a,a16640a,a16644a,a16645a,a16646a,a16649a,a16653a,a16654a,a16655a,a16658a,a16662a,a16663a,a16664a,a16667a,a16671a,a16672a,a16673a,a16676a,a16680a,a16681a,a16682a,a16685a,a16689a,a16690a,a16691a,a16694a,a16698a,a16699a,a16700a,a16703a,a16707a,a16708a,a16709a,a16712a,a16716a,a16717a,a16718a,a16721a,a16725a,a16726a,a16727a,a16730a,a16734a,a16735a,a16736a,a16739a,a16743a,a16744a,a16745a,a16748a,a16752a,a16753a,a16754a,a16757a,a16761a,a16762a,a16763a,a16766a,a16770a,a16771a,a16772a,a16775a,a16779a,a16780a,a16781a,a16784a,a16788a,a16789a,a16790a,a16793a,a16797a,a16798a,a16799a,a16802a,a16806a,a16807a,a16808a,a16811a,a16815a,a16816a,a16817a,a16820a,a16824a,a16825a,a16826a,a16829a,a16833a,a16834a,a16835a,a16838a,a16842a,a16843a,a16844a,a16847a,a16851a,a16852a,a16853a,a16856a,a16860a,a16861a,a16862a,a16865a,a16869a,a16870a,a16871a,a16874a,a16878a,a16879a,a16880a,a16883a,a16887a,a16888a,a16889a,a16892a,a16896a,a16897a,a16898a,a16901a,a16905a,a16906a,a16907a,a16910a,a16914a,a16915a,a16916a,a16919a,a16923a,a16924a,a16925a,a16928a,a16932a,a16933a,a16934a,a16937a,a16941a,a16942a,a16943a,a16946a,a16950a,a16951a,a16952a,a16955a,a16959a,a16960a,a16961a,a16964a,a16968a,a16969a,a16970a,a16973a,a16977a,a16978a,a16979a,a16982a,a16986a,a16987a,a16988a,a16991a,a16995a,a16996a,a16997a,a17000a,a17004a,a17005a,a17006a,a17009a,a17013a,a17014a,a17015a,a17018a,a17022a,a17023a,a17024a,a17027a,a17031a,a17032a,a17033a,a17036a,a17040a,a17041a,a17042a,a17045a,a17049a,a17050a,a17051a,a17054a,a17058a,a17059a,a17060a,a17063a,a17067a,a17068a,a17069a,a17072a,a17076a,a17077a,a17078a,a17081a,a17085a,a17086a,a17087a,a17090a,a17094a,a17095a,a17096a,a17099a,a17103a,a17104a,a17105a,a17108a,a17112a,a17113a,a17114a,a17117a,a17121a,a17122a,a17123a,a17126a,a17130a,a17131a,a17132a,a17135a,a17139a,a17140a,a17141a,a17144a,a17148a,a17149a,a17150a,a17153a,a17157a,a17158a,a17159a,a17162a,a17166a,a17167a,a17168a,a17171a,a17175a,a17176a,a17177a,a17180a,a17184a,a17185a,a17186a,a17189a,a17193a,a17194a,a17195a,a17198a,a17202a,a17203a,a17204a,a17207a,a17211a,a17212a,a17213a,a17216a,a17220a,a17221a,a17222a,a17225a,a17229a,a17230a,a17231a,a17234a,a17238a,a17239a,a17240a,a17243a,a17247a,a17248a,a17249a,a17252a,a17256a,a17257a,a17258a,a17261a,a17265a,a17266a,a17267a,a17270a,a17274a,a17275a,a17276a,a17279a,a17283a,a17284a,a17285a,a17288a,a17292a,a17293a,a17294a,a17297a,a17301a,a17302a,a17303a,a17306a,a17310a,a17311a,a17312a,a17315a,a17319a,a17320a,a17321a,a17324a,a17328a,a17329a,a17330a,a17333a,a17337a,a17338a,a17339a,a17342a,a17346a,a17347a,a17348a,a17351a,a17355a,a17356a,a17357a,a17360a,a17364a,a17365a,a17366a,a17369a,a17373a,a17374a,a17375a,a17378a,a17382a,a17383a,a17384a,a17387a,a17391a,a17392a,a17393a,a17396a,a17400a,a17401a,a17402a,a17405a,a17409a,a17410a,a17411a,a17414a,a17418a,a17419a,a17420a,a17423a,a17427a,a17428a,a17429a,a17432a,a17436a,a17437a,a17438a,a17441a,a17445a,a17446a,a17447a,a17450a,a17454a,a17455a,a17456a,a17459a,a17463a,a17464a,a17465a,a17469a,a17470a,a17474a,a17475a,a17476a,a17479a,a17483a,a17484a,a17485a,a17489a,a17490a,a17494a,a17495a,a17496a,a17499a,a17503a,a17504a,a17505a,a17509a,a17510a,a17514a,a17515a,a17516a,a17519a,a17523a,a17524a,a17525a,a17529a,a17530a,a17534a,a17535a,a17536a,a17539a,a17543a,a17544a,a17545a,a17549a,a17550a,a17554a,a17555a,a17556a,a17559a,a17563a,a17564a,a17565a,a17569a,a17570a,a17574a,a17575a,a17576a,a17579a,a17583a,a17584a,a17585a,a17589a,a17590a,a17594a,a17595a,a17596a,a17599a,a17603a,a17604a,a17605a,a17609a,a17610a,a17614a,a17615a,a17616a,a17619a,a17623a,a17624a,a17625a,a17629a,a17630a,a17634a,a17635a,a17636a,a17639a,a17643a,a17644a,a17645a,a17649a,a17650a,a17654a,a17655a,a17656a,a17659a,a17663a,a17664a,a17665a,a17669a,a17670a,a17674a,a17675a,a17676a,a17679a,a17683a,a17684a,a17685a,a17689a,a17690a,a17694a,a17695a,a17696a,a17699a,a17703a,a17704a,a17705a,a17709a,a17710a,a17714a,a17715a,a17716a,a17719a,a17723a,a17724a,a17725a,a17729a,a17730a,a17734a,a17735a,a17736a,a17739a,a17743a,a17744a,a17745a,a17749a,a17750a,a17754a,a17755a,a17756a,a17759a,a17763a,a17764a,a17765a,a17769a,a17770a,a17774a,a17775a,a17776a,a17779a,a17783a,a17784a,a17785a,a17789a,a17790a,a17794a,a17795a,a17796a,a17799a,a17803a,a17804a,a17805a,a17809a,a17810a,a17814a,a17815a,a17816a,a17819a,a17823a,a17824a,a17825a,a17829a,a17830a,a17834a,a17835a,a17836a,a17839a,a17843a,a17844a,a17845a,a17849a,a17850a,a17854a,a17855a,a17856a,a17859a,a17863a,a17864a,a17865a,a17869a,a17870a,a17874a,a17875a,a17876a,a17879a,a17883a,a17884a,a17885a,a17889a,a17890a,a17894a,a17895a,a17896a,a17899a,a17903a,a17904a,a17905a,a17909a,a17910a,a17914a,a17915a,a17916a,a17919a,a17923a,a17924a,a17925a,a17929a,a17930a,a17934a,a17935a,a17936a,a17939a,a17943a,a17944a,a17945a,a17949a,a17950a,a17954a,a17955a,a17956a,a17959a,a17963a,a17964a,a17965a,a17969a,a17970a,a17974a,a17975a,a17976a,a17979a,a17983a,a17984a,a17985a,a17989a,a17990a,a17994a,a17995a,a17996a,a17999a,a18003a,a18004a,a18005a,a18009a,a18010a,a18014a,a18015a,a18016a,a18019a,a18023a,a18024a,a18025a,a18029a,a18030a,a18034a,a18035a,a18036a,a18039a,a18043a,a18044a,a18045a,a18049a,a18050a,a18054a,a18055a,a18056a,a18059a,a18063a,a18064a,a18065a,a18069a,a18070a,a18074a,a18075a,a18076a,a18079a,a18083a,a18084a,a18085a,a18089a,a18090a,a18094a,a18095a,a18096a,a18099a,a18103a,a18104a,a18105a,a18109a,a18110a,a18114a,a18115a,a18116a,a18119a,a18123a,a18124a,a18125a,a18129a,a18130a,a18134a,a18135a,a18136a,a18139a,a18143a,a18144a,a18145a,a18149a,a18150a,a18154a,a18155a,a18156a,a18159a,a18163a,a18164a,a18165a,a18169a,a18170a,a18174a,a18175a,a18176a,a18179a,a18183a,a18184a,a18185a,a18189a,a18190a,a18194a,a18195a,a18196a,a18199a,a18203a,a18204a,a18205a,a18209a,a18210a,a18214a,a18215a,a18216a,a18219a,a18223a,a18224a,a18225a,a18229a,a18230a,a18234a,a18235a,a18236a,a18239a,a18243a,a18244a,a18245a,a18249a,a18250a,a18254a,a18255a,a18256a,a18259a,a18263a,a18264a,a18265a,a18269a,a18270a,a18274a,a18275a,a18276a,a18279a,a18283a,a18284a,a18285a,a18289a,a18290a,a18294a,a18295a,a18296a,a18299a,a18303a,a18304a,a18305a,a18309a,a18310a,a18314a,a18315a,a18316a,a18319a,a18323a,a18324a,a18325a,a18329a,a18330a,a18334a,a18335a,a18336a,a18339a,a18343a,a18344a,a18345a,a18349a,a18350a,a18354a,a18355a,a18356a,a18359a,a18363a,a18364a,a18365a,a18369a,a18370a,a18374a,a18375a,a18376a,a18379a,a18383a,a18384a,a18385a,a18389a,a18390a,a18394a,a18395a,a18396a,a18399a,a18403a,a18404a,a18405a,a18409a,a18410a,a18414a,a18415a,a18416a,a18419a,a18423a,a18424a,a18425a,a18429a,a18430a,a18434a,a18435a,a18436a,a18439a,a18443a,a18444a,a18445a,a18449a,a18450a,a18454a,a18455a,a18456a,a18459a,a18463a,a18464a,a18465a,a18469a,a18470a,a18474a,a18475a,a18476a,a18479a,a18483a,a18484a,a18485a,a18489a,a18490a,a18494a,a18495a,a18496a,a18499a,a18503a,a18504a,a18505a,a18509a,a18510a,a18514a,a18515a,a18516a,a18519a,a18523a,a18524a,a18525a,a18529a,a18530a,a18534a,a18535a,a18536a,a18539a,a18543a,a18544a,a18545a,a18549a,a18550a,a18554a,a18555a,a18556a,a18559a,a18563a,a18564a,a18565a,a18569a,a18570a,a18574a,a18575a,a18576a,a18579a,a18583a,a18584a,a18585a,a18589a,a18590a,a18594a,a18595a,a18596a,a18599a,a18603a,a18604a,a18605a,a18609a,a18610a,a18614a,a18615a,a18616a,a18619a,a18623a,a18624a,a18625a,a18629a,a18630a,a18634a,a18635a,a18636a,a18639a,a18643a,a18644a,a18645a,a18649a,a18650a,a18654a,a18655a,a18656a,a18659a,a18663a,a18664a,a18665a,a18669a,a18670a,a18674a,a18675a,a18676a,a18679a,a18683a,a18684a,a18685a,a18689a,a18690a,a18694a,a18695a,a18696a,a18699a,a18703a,a18704a,a18705a,a18709a,a18710a,a18714a,a18715a,a18716a,a18719a,a18723a,a18724a,a18725a,a18729a,a18730a,a18734a,a18735a,a18736a,a18739a,a18743a,a18744a,a18745a,a18749a,a18750a,a18754a,a18755a,a18756a,a18759a,a18763a,a18764a,a18765a,a18769a,a18770a,a18774a,a18775a,a18776a,a18779a,a18783a,a18784a,a18785a,a18789a,a18790a,a18794a,a18795a,a18796a,a18799a,a18803a,a18804a,a18805a,a18809a,a18810a,a18814a,a18815a,a18816a,a18819a,a18823a,a18824a,a18825a,a18829a,a18830a,a18834a,a18835a,a18836a,a18839a,a18843a,a18844a,a18845a,a18849a,a18850a,a18854a,a18855a,a18856a,a18859a,a18863a,a18864a,a18865a,a18869a,a18870a,a18874a,a18875a,a18876a,a18879a,a18883a,a18884a,a18885a,a18889a,a18890a,a18894a,a18895a,a18896a,a18899a,a18903a,a18904a,a18905a,a18909a,a18910a,a18914a,a18915a,a18916a,a18919a,a18923a,a18924a,a18925a,a18929a,a18930a,a18934a,a18935a,a18936a,a18939a,a18943a,a18944a,a18945a,a18949a,a18950a,a18954a,a18955a,a18956a,a18959a,a18963a,a18964a,a18965a,a18969a,a18970a,a18974a,a18975a,a18976a,a18979a,a18983a,a18984a,a18985a,a18989a,a18990a,a18994a,a18995a,a18996a,a18999a,a19003a,a19004a,a19005a,a19009a,a19010a,a19014a,a19015a,a19016a,a19019a,a19023a,a19024a,a19025a,a19029a,a19030a,a19034a,a19035a,a19036a,a19039a,a19043a,a19044a,a19045a,a19049a,a19050a,a19054a,a19055a,a19056a,a19059a,a19063a,a19064a,a19065a,a19069a,a19070a,a19074a,a19075a,a19076a,a19079a,a19083a,a19084a,a19085a,a19089a,a19090a,a19094a,a19095a,a19096a,a19099a,a19103a,a19104a,a19105a,a19109a,a19110a,a19114a,a19115a,a19116a,a19119a,a19123a,a19124a,a19125a,a19129a,a19130a,a19134a,a19135a,a19136a,a19139a,a19143a,a19144a,a19145a,a19149a,a19150a,a19154a,a19155a,a19156a,a19159a,a19163a,a19164a,a19165a,a19169a,a19170a,a19174a,a19175a,a19176a,a19179a,a19183a,a19184a,a19185a,a19189a,a19190a,a19194a,a19195a,a19196a,a19199a,a19203a,a19204a,a19205a,a19209a,a19210a,a19214a,a19215a,a19216a,a19219a,a19223a,a19224a,a19225a,a19229a,a19230a,a19234a,a19235a,a19236a,a19239a,a19243a,a19244a,a19245a,a19249a,a19250a,a19254a,a19255a,a19256a,a19259a,a19263a,a19264a,a19265a,a19269a,a19270a,a19274a,a19275a,a19276a,a19279a,a19283a,a19284a,a19285a,a19289a,a19290a,a19294a,a19295a,a19296a,a19299a,a19303a,a19304a,a19305a,a19309a,a19310a,a19314a,a19315a,a19316a,a19319a,a19323a,a19324a,a19325a,a19329a,a19330a,a19334a,a19335a,a19336a,a19339a,a19343a,a19344a,a19345a,a19349a,a19350a,a19354a,a19355a,a19356a,a19359a,a19363a,a19364a,a19365a,a19369a,a19370a,a19374a,a19375a,a19376a,a19379a,a19383a,a19384a,a19385a,a19389a,a19390a,a19394a,a19395a,a19396a,a19399a,a19403a,a19404a,a19405a,a19409a,a19410a,a19414a,a19415a,a19416a,a19419a,a19423a,a19424a,a19425a,a19429a,a19430a,a19434a,a19435a,a19436a,a19439a,a19443a,a19444a,a19445a,a19449a,a19450a,a19454a,a19455a,a19456a,a19459a,a19463a,a19464a,a19465a,a19469a,a19470a,a19474a,a19475a,a19476a,a19479a,a19483a,a19484a,a19485a,a19489a,a19490a,a19494a,a19495a,a19496a,a19499a,a19503a,a19504a,a19505a,a19509a,a19510a,a19514a,a19515a,a19516a,a19519a,a19523a,a19524a,a19525a,a19529a,a19530a,a19534a,a19535a,a19536a,a19539a,a19543a,a19544a,a19545a,a19549a,a19550a,a19554a,a19555a,a19556a,a19559a,a19563a,a19564a,a19565a,a19569a,a19570a,a19574a,a19575a,a19576a,a19579a,a19583a,a19584a,a19585a,a19589a,a19590a,a19594a,a19595a,a19596a,a19599a,a19603a,a19604a,a19605a,a19609a,a19610a,a19614a,a19615a,a19616a,a19619a,a19623a,a19624a,a19625a,a19629a,a19630a,a19634a,a19635a,a19636a,a19639a,a19643a,a19644a,a19645a,a19649a,a19650a,a19654a,a19655a,a19656a,a19659a,a19663a,a19664a,a19665a,a19669a,a19670a,a19674a,a19675a,a19676a,a19679a,a19683a,a19684a,a19685a,a19689a,a19690a,a19694a,a19695a,a19696a,a19699a,a19703a,a19704a,a19705a,a19709a,a19710a,a19714a,a19715a,a19716a,a19719a,a19723a,a19724a,a19725a,a19729a,a19730a,a19734a,a19735a,a19736a,a19739a,a19743a,a19744a,a19745a,a19749a,a19750a,a19754a,a19755a,a19756a,a19759a,a19763a,a19764a,a19765a,a19769a,a19770a,a19774a,a19775a,a19776a,a19779a,a19783a,a19784a,a19785a,a19789a,a19790a,a19794a,a19795a,a19796a,a19799a,a19803a,a19804a,a19805a,a19809a,a19810a,a19814a,a19815a,a19816a,a19819a,a19823a,a19824a,a19825a,a19829a,a19830a,a19834a,a19835a,a19836a,a19839a,a19843a,a19844a,a19845a,a19849a,a19850a,a19854a,a19855a,a19856a,a19859a,a19863a,a19864a,a19865a,a19869a,a19870a,a19874a,a19875a,a19876a,a19879a,a19883a,a19884a,a19885a,a19889a,a19890a,a19894a,a19895a,a19896a,a19899a,a19903a,a19904a,a19905a,a19909a,a19910a,a19914a,a19915a,a19916a,a19919a,a19923a,a19924a,a19925a,a19929a,a19930a,a19934a,a19935a,a19936a,a19939a,a19943a,a19944a,a19945a,a19949a,a19950a,a19954a,a19955a,a19956a,a19959a,a19963a,a19964a,a19965a,a19969a,a19970a,a19974a,a19975a,a19976a,a19979a,a19983a,a19984a,a19985a,a19989a,a19990a,a19994a,a19995a,a19996a,a19999a,a20003a,a20004a,a20005a,a20009a,a20010a,a20014a,a20015a,a20016a,a20019a,a20023a,a20024a,a20025a,a20029a,a20030a,a20034a,a20035a,a20036a,a20039a,a20043a,a20044a,a20045a,a20049a,a20050a,a20054a,a20055a,a20056a,a20059a,a20063a,a20064a,a20065a,a20069a,a20070a,a20074a,a20075a,a20076a,a20079a,a20083a,a20084a,a20085a,a20089a,a20090a,a20094a,a20095a,a20096a,a20099a,a20103a,a20104a,a20105a,a20109a,a20110a,a20114a,a20115a,a20116a,a20119a,a20123a,a20124a,a20125a,a20129a,a20130a,a20134a,a20135a,a20136a,a20139a,a20143a,a20144a,a20145a,a20149a,a20150a,a20154a,a20155a,a20156a,a20159a,a20163a,a20164a,a20165a,a20169a,a20170a,a20174a,a20175a,a20176a,a20179a,a20183a,a20184a,a20185a,a20189a,a20190a,a20194a,a20195a,a20196a,a20199a,a20203a,a20204a,a20205a,a20209a,a20210a,a20214a,a20215a,a20216a,a20219a,a20223a,a20224a,a20225a,a20229a,a20230a,a20234a,a20235a,a20236a,a20239a,a20243a,a20244a,a20245a,a20249a,a20250a,a20254a,a20255a,a20256a,a20259a,a20263a,a20264a,a20265a,a20269a,a20270a,a20274a,a20275a,a20276a,a20279a,a20283a,a20284a,a20285a,a20289a,a20290a,a20294a,a20295a,a20296a,a20299a,a20303a,a20304a,a20305a,a20309a,a20310a,a20314a,a20315a,a20316a,a20319a,a20323a,a20324a,a20325a,a20329a,a20330a,a20334a,a20335a,a20336a,a20339a,a20343a,a20344a,a20345a,a20349a,a20350a,a20354a,a20355a,a20356a,a20359a,a20363a,a20364a,a20365a,a20369a,a20370a,a20374a,a20375a,a20376a,a20379a,a20383a,a20384a,a20385a,a20389a,a20390a,a20394a,a20395a,a20396a,a20399a,a20403a,a20404a,a20405a,a20409a,a20410a,a20414a,a20415a,a20416a,a20419a,a20423a,a20424a,a20425a,a20429a,a20430a,a20434a,a20435a,a20436a,a20439a,a20443a,a20444a,a20445a,a20449a,a20450a,a20454a,a20455a,a20456a,a20459a,a20463a,a20464a,a20465a,a20469a,a20470a,a20474a,a20475a,a20476a,a20479a,a20483a,a20484a,a20485a,a20489a,a20490a,a20494a,a20495a,a20496a,a20499a,a20503a,a20504a,a20505a,a20509a,a20510a,a20514a,a20515a,a20516a,a20519a,a20523a,a20524a,a20525a,a20529a,a20530a,a20534a,a20535a,a20536a,a20539a,a20543a,a20544a,a20545a,a20549a,a20550a,a20554a,a20555a,a20556a,a20559a,a20563a,a20564a,a20565a,a20569a,a20570a,a20574a,a20575a,a20576a,a20579a,a20583a,a20584a,a20585a,a20589a,a20590a,a20594a,a20595a,a20596a,a20599a,a20603a,a20604a,a20605a,a20609a,a20610a,a20614a,a20615a,a20616a,a20619a,a20623a,a20624a,a20625a,a20629a,a20630a,a20634a,a20635a,a20636a,a20639a,a20643a,a20644a,a20645a,a20649a,a20650a,a20654a,a20655a,a20656a,a20659a,a20663a,a20664a,a20665a,a20669a,a20670a,a20674a,a20675a,a20676a,a20679a,a20683a,a20684a,a20685a,a20689a,a20690a,a20694a,a20695a,a20696a,a20699a,a20703a,a20704a,a20705a,a20709a,a20710a,a20714a,a20715a,a20716a,a20719a,a20723a,a20724a,a20725a,a20729a,a20730a,a20734a,a20735a,a20736a,a20739a,a20743a,a20744a,a20745a,a20749a,a20750a,a20754a,a20755a,a20756a,a20759a,a20763a,a20764a,a20765a,a20769a,a20770a,a20774a,a20775a,a20776a,a20779a,a20783a,a20784a,a20785a,a20789a,a20790a,a20794a,a20795a,a20796a,a20799a,a20803a,a20804a,a20805a,a20809a,a20810a,a20814a,a20815a,a20816a,a20819a,a20823a,a20824a,a20825a,a20829a,a20830a,a20834a,a20835a,a20836a,a20839a,a20843a,a20844a,a20845a,a20849a,a20850a,a20854a,a20855a,a20856a,a20859a,a20863a,a20864a,a20865a,a20869a,a20870a,a20874a,a20875a,a20876a,a20879a,a20883a,a20884a,a20885a,a20889a,a20890a,a20894a,a20895a,a20896a,a20899a,a20903a,a20904a,a20905a,a20909a,a20910a,a20914a,a20915a,a20916a,a20919a,a20923a,a20924a,a20925a,a20929a,a20930a,a20934a,a20935a,a20936a,a20939a,a20943a,a20944a,a20945a,a20949a,a20950a,a20954a,a20955a,a20956a,a20959a,a20963a,a20964a,a20965a,a20969a,a20970a,a20974a,a20975a,a20976a,a20979a,a20983a,a20984a,a20985a,a20989a,a20990a,a20994a,a20995a,a20996a,a20999a,a21003a,a21004a,a21005a,a21009a,a21010a,a21014a,a21015a,a21016a,a21019a,a21023a,a21024a,a21025a,a21029a,a21030a,a21034a,a21035a,a21036a,a21039a,a21043a,a21044a,a21045a,a21049a,a21050a,a21054a,a21055a,a21056a,a21059a,a21063a,a21064a,a21065a,a21069a,a21070a,a21074a,a21075a,a21076a,a21079a,a21083a,a21084a,a21085a,a21089a,a21090a,a21094a,a21095a,a21096a,a21099a,a21103a,a21104a,a21105a,a21109a,a21110a,a21114a,a21115a,a21116a,a21119a,a21123a,a21124a,a21125a,a21129a,a21130a,a21134a,a21135a,a21136a,a21139a,a21143a,a21144a,a21145a,a21149a,a21150a,a21154a,a21155a,a21156a,a21159a,a21163a,a21164a,a21165a,a21169a,a21170a,a21174a,a21175a,a21176a,a21179a,a21183a,a21184a,a21185a,a21189a,a21190a,a21194a,a21195a,a21196a,a21199a,a21203a,a21204a,a21205a,a21209a,a21210a,a21214a,a21215a,a21216a,a21219a,a21223a,a21224a,a21225a,a21229a,a21230a,a21234a,a21235a,a21236a,a21239a,a21243a,a21244a,a21245a,a21249a,a21250a,a21254a,a21255a,a21256a,a21259a,a21263a,a21264a,a21265a,a21269a,a21270a,a21274a,a21275a,a21276a,a21279a,a21283a,a21284a,a21285a,a21289a,a21290a,a21294a,a21295a,a21296a,a21299a,a21303a,a21304a,a21305a,a21309a,a21310a,a21314a,a21315a,a21316a,a21319a,a21323a,a21324a,a21325a,a21329a,a21330a,a21334a,a21335a,a21336a,a21339a,a21343a,a21344a,a21345a,a21349a,a21350a,a21354a,a21355a,a21356a,a21359a,a21363a,a21364a,a21365a,a21369a,a21370a,a21374a,a21375a,a21376a,a21379a,a21383a,a21384a,a21385a,a21389a,a21390a,a21394a,a21395a,a21396a,a21399a,a21403a,a21404a,a21405a,a21409a,a21410a,a21414a,a21415a,a21416a,a21419a,a21423a,a21424a,a21425a,a21429a,a21430a,a21434a,a21435a,a21436a,a21439a,a21443a,a21444a,a21445a,a21449a,a21450a,a21454a,a21455a,a21456a,a21459a,a21463a,a21464a,a21465a,a21469a,a21470a,a21474a,a21475a,a21476a,a21479a,a21483a,a21484a,a21485a,a21489a,a21490a,a21494a,a21495a,a21496a,a21499a,a21503a,a21504a,a21505a,a21509a,a21510a,a21514a,a21515a,a21516a,a21519a,a21523a,a21524a,a21525a,a21529a,a21530a,a21534a,a21535a,a21536a,a21539a,a21543a,a21544a,a21545a,a21549a,a21550a,a21554a,a21555a,a21556a,a21559a,a21563a,a21564a,a21565a,a21569a,a21570a,a21574a,a21575a,a21576a,a21579a,a21583a,a21584a,a21585a,a21589a,a21590a,a21594a,a21595a,a21596a,a21599a,a21603a,a21604a,a21605a,a21609a,a21610a,a21614a,a21615a,a21616a,a21619a,a21623a,a21624a,a21625a,a21629a,a21630a,a21634a,a21635a,a21636a,a21639a,a21643a,a21644a,a21645a,a21649a,a21650a,a21654a,a21655a,a21656a,a21659a,a21663a,a21664a,a21665a,a21669a,a21670a,a21674a,a21675a,a21676a,a21679a,a21683a,a21684a,a21685a,a21689a,a21690a,a21694a,a21695a,a21696a,a21699a,a21703a,a21704a,a21705a,a21709a,a21710a,a21714a,a21715a,a21716a,a21719a,a21723a,a21724a,a21725a,a21729a,a21730a,a21734a,a21735a,a21736a,a21739a,a21743a,a21744a,a21745a,a21749a,a21750a,a21754a,a21755a,a21756a,a21759a,a21763a,a21764a,a21765a,a21769a,a21770a,a21774a,a21775a,a21776a,a21779a,a21783a,a21784a,a21785a,a21789a,a21790a,a21794a,a21795a,a21796a,a21799a,a21803a,a21804a,a21805a,a21809a,a21810a,a21814a,a21815a,a21816a,a21819a,a21823a,a21824a,a21825a,a21829a,a21830a,a21834a,a21835a,a21836a,a21839a,a21843a,a21844a,a21845a,a21849a,a21850a,a21854a,a21855a,a21856a,a21859a,a21863a,a21864a,a21865a,a21869a,a21870a,a21874a,a21875a,a21876a,a21879a,a21883a,a21884a,a21885a,a21889a,a21890a,a21894a,a21895a,a21896a,a21899a,a21903a,a21904a,a21905a,a21909a,a21910a,a21914a,a21915a,a21916a,a21919a,a21923a,a21924a,a21925a,a21929a,a21930a,a21934a,a21935a,a21936a,a21939a,a21943a,a21944a,a21945a,a21949a,a21950a,a21954a,a21955a,a21956a,a21959a,a21963a,a21964a,a21965a,a21969a,a21970a,a21974a,a21975a,a21976a,a21979a,a21983a,a21984a,a21985a,a21989a,a21990a,a21994a,a21995a,a21996a,a21999a,a22003a,a22004a,a22005a,a22009a,a22010a,a22014a,a22015a,a22016a,a22019a,a22023a,a22024a,a22025a,a22029a,a22030a,a22034a,a22035a,a22036a,a22039a,a22043a,a22044a,a22045a,a22049a,a22050a,a22054a,a22055a,a22056a,a22059a,a22063a,a22064a,a22065a,a22069a,a22070a,a22074a,a22075a,a22076a,a22079a,a22083a,a22084a,a22085a,a22089a,a22090a,a22094a,a22095a,a22096a,a22099a,a22103a,a22104a,a22105a,a22109a,a22110a,a22114a,a22115a,a22116a,a22119a,a22123a,a22124a,a22125a,a22129a,a22130a,a22134a,a22135a,a22136a,a22139a,a22143a,a22144a,a22145a,a22149a,a22150a,a22154a,a22155a,a22156a,a22159a,a22163a,a22164a,a22165a,a22169a,a22170a,a22174a,a22175a,a22176a,a22179a,a22183a,a22184a,a22185a,a22189a,a22190a,a22194a,a22195a,a22196a,a22199a,a22203a,a22204a,a22205a,a22209a,a22210a,a22214a,a22215a,a22216a,a22219a,a22223a,a22224a,a22225a,a22229a,a22230a,a22234a,a22235a,a22236a,a22239a,a22243a,a22244a,a22245a,a22249a,a22250a,a22254a,a22255a,a22256a,a22259a,a22263a,a22264a,a22265a,a22269a,a22270a,a22274a,a22275a,a22276a,a22279a,a22283a,a22284a,a22285a,a22289a,a22290a,a22294a,a22295a,a22296a,a22299a,a22303a,a22304a,a22305a,a22309a,a22310a,a22314a,a22315a,a22316a,a22319a,a22323a,a22324a,a22325a,a22329a,a22330a,a22334a,a22335a,a22336a,a22339a,a22343a,a22344a,a22345a,a22349a,a22350a,a22354a,a22355a,a22356a,a22359a,a22363a,a22364a,a22365a,a22369a,a22370a,a22374a,a22375a,a22376a,a22379a,a22383a,a22384a,a22385a,a22389a,a22390a,a22394a,a22395a,a22396a,a22399a,a22403a,a22404a,a22405a,a22409a,a22410a,a22414a,a22415a,a22416a,a22419a,a22423a,a22424a,a22425a,a22429a,a22430a,a22434a,a22435a,a22436a,a22439a,a22443a,a22444a,a22445a,a22449a,a22450a,a22454a,a22455a,a22456a,a22459a,a22463a,a22464a,a22465a,a22469a,a22470a,a22474a,a22475a,a22476a,a22479a,a22483a,a22484a,a22485a,a22489a,a22490a,a22494a,a22495a,a22496a,a22499a,a22503a,a22504a,a22505a,a22509a,a22510a,a22514a,a22515a,a22516a,a22519a,a22523a,a22524a,a22525a,a22529a,a22530a,a22534a,a22535a,a22536a,a22539a,a22543a,a22544a,a22545a,a22549a,a22550a,a22554a,a22555a,a22556a,a22559a,a22563a,a22564a,a22565a,a22569a,a22570a,a22574a,a22575a,a22576a,a22579a,a22583a,a22584a,a22585a,a22589a,a22590a,a22594a,a22595a,a22596a,a22599a,a22603a,a22604a,a22605a,a22609a,a22610a,a22614a,a22615a,a22616a,a22619a,a22623a,a22624a,a22625a,a22629a,a22630a,a22634a,a22635a,a22636a,a22639a,a22643a,a22644a,a22645a,a22649a,a22650a,a22654a,a22655a,a22656a,a22659a,a22663a,a22664a,a22665a,a22669a,a22670a,a22674a,a22675a,a22676a,a22679a,a22683a,a22684a,a22685a,a22689a,a22690a,a22694a,a22695a,a22696a,a22699a,a22703a,a22704a,a22705a,a22709a,a22710a,a22714a,a22715a,a22716a,a22719a,a22723a,a22724a,a22725a,a22729a,a22730a,a22734a,a22735a,a22736a,a22739a,a22743a,a22744a,a22745a,a22749a,a22750a,a22754a,a22755a,a22756a,a22759a,a22763a,a22764a,a22765a,a22769a,a22770a,a22774a,a22775a,a22776a,a22779a,a22783a,a22784a,a22785a,a22789a,a22790a,a22794a,a22795a,a22796a,a22799a,a22803a,a22804a,a22805a,a22809a,a22810a,a22814a,a22815a,a22816a,a22819a,a22823a,a22824a,a22825a,a22829a,a22830a,a22834a,a22835a,a22836a,a22839a,a22843a,a22844a,a22845a,a22849a,a22850a,a22854a,a22855a,a22856a,a22859a,a22863a,a22864a,a22865a,a22869a,a22870a,a22874a,a22875a,a22876a,a22879a,a22883a,a22884a,a22885a,a22889a,a22890a,a22894a,a22895a,a22896a,a22899a,a22903a,a22904a,a22905a,a22909a,a22910a,a22914a,a22915a,a22916a,a22919a,a22923a,a22924a,a22925a,a22929a,a22930a,a22934a,a22935a,a22936a,a22939a,a22943a,a22944a,a22945a,a22949a,a22950a,a22954a,a22955a,a22956a,a22959a,a22963a,a22964a,a22965a,a22969a,a22970a,a22974a,a22975a,a22976a,a22979a,a22983a,a22984a,a22985a,a22989a,a22990a,a22994a,a22995a,a22996a,a22999a,a23003a,a23004a,a23005a,a23009a,a23010a,a23014a,a23015a,a23016a,a23019a,a23023a,a23024a,a23025a,a23029a,a23030a,a23034a,a23035a,a23036a,a23039a,a23043a,a23044a,a23045a,a23049a,a23050a,a23054a,a23055a,a23056a,a23059a,a23063a,a23064a,a23065a,a23069a,a23070a,a23074a,a23075a,a23076a,a23079a,a23083a,a23084a,a23085a,a23089a,a23090a,a23094a,a23095a,a23096a,a23099a,a23103a,a23104a,a23105a,a23109a,a23110a,a23114a,a23115a,a23116a,a23119a,a23123a,a23124a,a23125a,a23129a,a23130a,a23134a,a23135a,a23136a,a23139a,a23143a,a23144a,a23145a,a23149a,a23150a,a23154a,a23155a,a23156a,a23159a,a23163a,a23164a,a23165a,a23169a,a23170a,a23174a,a23175a,a23176a,a23179a,a23183a,a23184a,a23185a,a23189a,a23190a,a23194a,a23195a,a23196a,a23199a,a23203a,a23204a,a23205a,a23209a,a23210a,a23214a,a23215a,a23216a,a23219a,a23223a,a23224a,a23225a,a23229a,a23230a,a23234a,a23235a,a23236a,a23239a,a23243a,a23244a,a23245a,a23249a,a23250a,a23254a,a23255a,a23256a,a23259a,a23263a,a23264a,a23265a,a23269a,a23270a,a23274a,a23275a,a23276a,a23279a,a23283a,a23284a,a23285a,a23289a,a23290a,a23294a,a23295a,a23296a,a23299a,a23303a,a23304a,a23305a,a23309a,a23310a,a23314a,a23315a,a23316a,a23319a,a23323a,a23324a,a23325a,a23329a,a23330a,a23334a,a23335a,a23336a,a23339a,a23343a,a23344a,a23345a,a23349a,a23350a,a23354a,a23355a,a23356a,a23359a,a23363a,a23364a,a23365a,a23369a,a23370a,a23374a,a23375a,a23376a,a23379a,a23383a,a23384a,a23385a,a23389a,a23390a,a23394a,a23395a,a23396a,a23399a,a23403a,a23404a,a23405a,a23409a,a23410a,a23414a,a23415a,a23416a,a23419a,a23423a,a23424a,a23425a,a23429a,a23430a,a23434a,a23435a,a23436a,a23439a,a23443a,a23444a,a23445a,a23449a,a23450a,a23454a,a23455a,a23456a,a23459a,a23463a,a23464a,a23465a,a23469a,a23470a,a23474a,a23475a,a23476a,a23479a,a23483a,a23484a,a23485a,a23489a,a23490a,a23494a,a23495a,a23496a,a23499a,a23503a,a23504a,a23505a,a23509a,a23510a,a23514a,a23515a,a23516a,a23519a,a23523a,a23524a,a23525a,a23529a,a23530a,a23534a,a23535a,a23536a,a23539a,a23543a,a23544a,a23545a,a23549a,a23550a,a23554a,a23555a,a23556a,a23559a,a23563a,a23564a,a23565a,a23569a,a23570a,a23574a,a23575a,a23576a,a23579a,a23583a,a23584a,a23585a,a23589a,a23590a,a23594a,a23595a,a23596a,a23599a,a23603a,a23604a,a23605a,a23609a,a23610a,a23614a,a23615a,a23616a,a23619a,a23623a,a23624a,a23625a,a23629a,a23630a,a23634a,a23635a,a23636a,a23639a,a23643a,a23644a,a23645a,a23649a,a23650a,a23654a,a23655a,a23656a,a23659a,a23663a,a23664a,a23665a,a23669a,a23670a,a23674a,a23675a,a23676a,a23679a,a23683a,a23684a,a23685a,a23689a,a23690a,a23694a,a23695a,a23696a,a23699a,a23703a,a23704a,a23705a,a23709a,a23710a,a23714a,a23715a,a23716a,a23719a,a23723a,a23724a,a23725a,a23729a,a23730a,a23734a,a23735a,a23736a,a23739a,a23743a,a23744a,a23745a,a23749a,a23750a,a23754a,a23755a,a23756a,a23759a,a23763a,a23764a,a23765a,a23769a,a23770a,a23774a,a23775a,a23776a,a23779a,a23783a,a23784a,a23785a,a23789a,a23790a,a23794a,a23795a,a23796a,a23799a,a23803a,a23804a,a23805a,a23809a,a23810a,a23814a,a23815a,a23816a,a23819a,a23823a,a23824a,a23825a,a23829a,a23830a,a23834a,a23835a,a23836a,a23839a,a23843a,a23844a,a23845a,a23849a,a23850a,a23854a,a23855a,a23856a,a23859a,a23863a,a23864a,a23865a,a23869a,a23870a,a23874a,a23875a,a23876a,a23879a,a23883a,a23884a,a23885a,a23889a,a23890a,a23894a,a23895a,a23896a,a23899a,a23903a,a23904a,a23905a,a23909a,a23910a,a23914a,a23915a,a23916a,a23919a,a23923a,a23924a,a23925a,a23929a,a23930a,a23934a,a23935a,a23936a,a23939a,a23943a,a23944a,a23945a,a23949a,a23950a,a23954a,a23955a,a23956a,a23959a,a23963a,a23964a,a23965a,a23969a,a23970a,a23974a,a23975a,a23976a,a23979a,a23983a,a23984a,a23985a,a23989a,a23990a,a23994a,a23995a,a23996a,a23999a,a24003a,a24004a,a24005a,a24009a,a24010a,a24014a,a24015a,a24016a,a24019a,a24023a,a24024a,a24025a,a24029a,a24030a,a24034a,a24035a,a24036a,a24039a,a24043a,a24044a,a24045a,a24049a,a24050a,a24054a,a24055a,a24056a,a24059a,a24063a,a24064a,a24065a,a24069a,a24070a,a24074a,a24075a,a24076a,a24079a,a24083a,a24084a,a24085a,a24089a,a24090a,a24094a,a24095a,a24096a,a24099a,a24103a,a24104a,a24105a,a24109a,a24110a,a24114a,a24115a,a24116a,a24119a,a24123a,a24124a,a24125a,a24129a,a24130a,a24134a,a24135a,a24136a,a24139a,a24143a,a24144a,a24145a,a24149a,a24150a,a24154a,a24155a,a24156a,a24159a,a24163a,a24164a,a24165a,a24169a,a24170a,a24174a,a24175a,a24176a,a24179a,a24183a,a24184a,a24185a,a24189a,a24190a,a24194a,a24195a,a24196a,a24199a,a24203a,a24204a,a24205a,a24209a,a24210a,a24214a,a24215a,a24216a,a24219a,a24223a,a24224a,a24225a,a24229a,a24230a,a24234a,a24235a,a24236a,a24239a,a24243a,a24244a,a24245a,a24249a,a24250a,a24254a,a24255a,a24256a,a24259a,a24263a,a24264a,a24265a,a24269a,a24270a,a24274a,a24275a,a24276a,a24279a,a24283a,a24284a,a24285a,a24289a,a24290a,a24294a,a24295a,a24296a,a24299a,a24303a,a24304a,a24305a,a24309a,a24310a,a24314a,a24315a,a24316a,a24319a,a24323a,a24324a,a24325a,a24329a,a24330a,a24334a,a24335a,a24336a,a24339a,a24343a,a24344a,a24345a,a24349a,a24350a,a24354a,a24355a,a24356a,a24359a,a24363a,a24364a,a24365a,a24369a,a24370a,a24374a,a24375a,a24376a,a24379a,a24383a,a24384a,a24385a,a24389a,a24390a,a24394a,a24395a,a24396a,a24399a,a24403a,a24404a,a24405a,a24409a,a24410a,a24414a,a24415a,a24416a,a24419a,a24423a,a24424a,a24425a,a24429a,a24430a,a24434a,a24435a,a24436a,a24439a,a24443a,a24444a,a24445a,a24449a,a24450a,a24454a,a24455a,a24456a,a24459a,a24463a,a24464a,a24465a,a24469a,a24470a,a24474a,a24475a,a24476a,a24479a,a24483a,a24484a,a24485a,a24489a,a24490a,a24494a,a24495a,a24496a,a24500a,a24501a,a24505a,a24506a,a24507a,a24511a,a24512a,a24516a,a24517a,a24518a,a24522a,a24523a,a24527a,a24528a,a24529a,a24533a,a24534a,a24538a,a24539a,a24540a,a24544a,a24545a,a24549a,a24550a,a24551a,a24555a,a24556a,a24560a,a24561a,a24562a,a24566a,a24567a,a24571a,a24572a,a24573a,a24577a,a24578a,a24582a,a24583a,a24584a,a24588a,a24589a,a24593a,a24594a,a24595a,a24599a,a24600a,a24604a,a24605a,a24606a,a24610a,a24611a,a24615a,a24616a,a24617a,a24621a,a24622a,a24626a,a24627a,a24628a,a24632a,a24633a,a24637a,a24638a,a24639a,a24643a,a24644a,a24648a,a24649a,a24650a,a24654a,a24655a,a24659a,a24660a,a24661a,a24665a,a24666a,a24670a,a24671a,a24672a,a24676a,a24677a,a24681a,a24682a,a24683a,a24687a,a24688a,a24692a,a24693a,a24694a,a24698a,a24699a,a24703a,a24704a,a24705a,a24709a,a24710a,a24714a,a24715a,a24716a,a24720a,a24721a,a24725a,a24726a,a24727a,a24731a,a24732a,a24736a,a24737a,a24738a,a24742a,a24743a,a24747a,a24748a,a24749a,a24753a,a24754a,a24758a,a24759a,a24760a,a24764a,a24765a,a24769a,a24770a,a24771a,a24775a,a24776a,a24780a,a24781a,a24782a,a24786a,a24787a,a24791a,a24792a,a24793a,a24797a,a24798a,a24802a,a24803a,a24804a,a24808a,a24809a,a24813a,a24814a,a24815a,a24819a,a24820a,a24824a,a24825a,a24826a,a24830a,a24831a,a24835a,a24836a,a24837a,a24841a,a24842a,a24846a,a24847a,a24848a,a24852a,a24853a,a24857a,a24858a,a24859a,a24863a,a24864a,a24868a,a24869a,a24870a,a24874a,a24875a,a24879a,a24880a,a24881a,a24885a,a24886a,a24890a,a24891a,a24892a,a24896a,a24897a,a24901a,a24902a,a24903a,a24907a,a24908a,a24912a,a24913a,a24914a,a24918a,a24919a,a24923a,a24924a,a24925a,a24929a,a24930a,a24934a,a24935a,a24936a,a24940a,a24941a,a24945a,a24946a,a24947a,a24951a,a24952a,a24956a,a24957a,a24958a,a24962a,a24963a,a24967a,a24968a,a24969a,a24973a,a24974a,a24978a,a24979a,a24980a,a24984a,a24985a,a24989a,a24990a,a24991a,a24995a,a24996a,a25000a,a25001a,a25002a,a25006a,a25007a,a25011a,a25012a,a25013a,a25017a,a25018a,a25022a,a25023a,a25024a,a25028a,a25029a,a25033a,a25034a,a25035a,a25039a,a25040a,a25044a,a25045a,a25046a,a25050a,a25051a,a25055a,a25056a,a25057a,a25061a,a25062a,a25066a,a25067a,a25068a,a25072a,a25073a,a25077a,a25078a,a25079a,a25083a,a25084a,a25088a,a25089a,a25090a,a25094a,a25095a,a25099a,a25100a,a25101a,a25105a,a25106a,a25110a,a25111a,a25112a,a25116a,a25117a,a25121a,a25122a,a25123a,a25127a,a25128a,a25132a,a25133a,a25134a,a25138a,a25139a,a25143a,a25144a,a25145a,a25149a,a25150a,a25154a,a25155a,a25156a,a25160a,a25161a,a25165a,a25166a,a25167a,a25171a,a25172a,a25176a,a25177a,a25178a,a25182a,a25183a,a25187a,a25188a,a25189a,a25193a,a25194a,a25198a,a25199a,a25200a,a25204a,a25205a,a25209a,a25210a,a25211a,a25215a,a25216a,a25220a,a25221a,a25222a,a25226a,a25227a,a25231a,a25232a,a25233a,a25237a,a25238a,a25242a,a25243a,a25244a,a25248a,a25249a,a25253a,a25254a,a25255a,a25259a,a25260a,a25264a,a25265a,a25266a,a25270a,a25271a,a25275a,a25276a,a25277a,a25281a,a25282a,a25286a,a25287a,a25288a,a25292a,a25293a,a25297a,a25298a,a25299a,a25303a,a25304a,a25308a,a25309a,a25310a,a25314a,a25315a,a25319a,a25320a,a25321a,a25325a,a25326a,a25330a,a25331a,a25332a,a25336a,a25337a,a25341a,a25342a,a25343a,a25347a,a25348a,a25352a,a25353a,a25354a,a25358a,a25359a,a25363a,a25364a,a25365a,a25369a,a25370a,a25374a,a25375a,a25376a,a25380a,a25381a,a25385a,a25386a,a25387a,a25391a,a25392a,a25396a,a25397a,a25398a,a25402a,a25403a,a25407a,a25408a,a25409a,a25413a,a25414a,a25418a,a25419a,a25420a,a25424a,a25425a,a25429a,a25430a,a25431a,a25435a,a25436a,a25440a,a25441a,a25442a,a25446a,a25447a,a25451a,a25452a,a25453a,a25457a,a25458a,a25462a,a25463a,a25464a,a25468a,a25469a,a25473a,a25474a,a25475a,a25479a,a25480a,a25484a,a25485a,a25486a,a25490a,a25491a,a25495a,a25496a,a25497a,a25501a,a25502a,a25506a,a25507a,a25508a,a25512a,a25513a,a25517a,a25518a,a25519a,a25523a,a25524a,a25528a,a25529a,a25530a,a25534a,a25535a,a25539a,a25540a,a25541a,a25545a,a25546a,a25550a,a25551a,a25552a,a25556a,a25557a,a25561a,a25562a,a25563a,a25567a,a25568a,a25572a,a25573a,a25574a,a25578a,a25579a,a25583a,a25584a,a25585a,a25589a,a25590a,a25594a,a25595a,a25596a,a25600a,a25601a,a25605a,a25606a,a25607a,a25611a,a25612a,a25616a,a25617a,a25618a,a25622a,a25623a,a25627a,a25628a,a25629a,a25633a,a25634a,a25638a,a25639a,a25640a,a25644a,a25645a,a25649a,a25650a,a25651a,a25655a,a25656a,a25660a,a25661a,a25662a,a25666a,a25667a,a25671a,a25672a,a25673a,a25677a,a25678a,a25682a,a25683a,a25684a,a25688a,a25689a,a25693a,a25694a,a25695a,a25699a,a25700a,a25704a,a25705a,a25706a,a25710a,a25711a,a25715a,a25716a,a25717a,a25721a,a25722a,a25726a,a25727a,a25728a,a25732a,a25733a,a25737a,a25738a,a25739a,a25743a,a25744a,a25748a,a25749a,a25750a,a25754a,a25755a,a25759a,a25760a,a25761a,a25765a,a25766a,a25770a,a25771a,a25772a,a25776a,a25777a,a25781a,a25782a,a25783a,a25787a,a25788a,a25792a,a25793a,a25794a,a25798a,a25799a,a25803a,a25804a,a25805a,a25809a,a25810a,a25814a,a25815a,a25816a,a25820a,a25821a,a25825a,a25826a,a25827a,a25831a,a25832a,a25836a,a25837a,a25838a,a25842a,a25843a,a25847a,a25848a,a25849a,a25853a,a25854a,a25858a,a25859a,a25860a,a25864a,a25865a,a25869a,a25870a,a25871a,a25875a,a25876a,a25880a,a25881a,a25882a,a25886a,a25887a,a25891a,a25892a,a25893a,a25897a,a25898a,a25902a,a25903a,a25904a,a25908a,a25909a,a25913a,a25914a,a25915a,a25919a,a25920a,a25924a,a25925a,a25926a,a25930a,a25931a,a25935a,a25936a,a25937a,a25941a,a25942a,a25946a,a25947a,a25948a,a25952a,a25953a,a25957a,a25958a,a25959a,a25963a,a25964a,a25968a,a25969a,a25970a,a25974a,a25975a,a25979a,a25980a,a25981a,a25985a,a25986a,a25990a,a25991a,a25992a,a25996a,a25997a,a26001a,a26002a,a26003a,a26007a,a26008a,a26012a,a26013a,a26014a,a26018a,a26019a,a26023a,a26024a,a26025a,a26029a,a26030a,a26034a,a26035a,a26036a,a26040a,a26041a,a26045a,a26046a,a26047a,a26051a,a26052a,a26056a,a26057a,a26058a,a26062a,a26063a,a26067a,a26068a,a26069a,a26073a,a26074a,a26078a,a26079a,a26080a,a26084a,a26085a,a26089a,a26090a,a26091a,a26095a,a26096a,a26100a,a26101a,a26102a,a26106a,a26107a,a26111a,a26112a,a26113a,a26117a,a26118a,a26122a,a26123a,a26124a,a26128a,a26129a,a26133a,a26134a,a26135a,a26139a,a26140a,a26144a,a26145a,a26146a,a26150a,a26151a,a26155a,a26156a,a26157a,a26161a,a26162a,a26166a,a26167a,a26168a,a26172a,a26173a,a26177a,a26178a,a26179a,a26183a,a26184a,a26188a,a26189a,a26190a,a26194a,a26195a,a26199a,a26200a,a26201a,a26205a,a26206a,a26210a,a26211a,a26212a,a26216a,a26217a,a26221a,a26222a,a26223a,a26227a,a26228a,a26232a,a26233a,a26234a,a26238a,a26239a,a26243a,a26244a,a26245a,a26249a,a26250a,a26254a,a26255a,a26256a,a26260a,a26261a,a26265a,a26266a,a26267a,a26271a,a26272a,a26276a,a26277a,a26278a,a26282a,a26283a,a26287a,a26288a,a26289a,a26293a,a26294a,a26298a,a26299a,a26300a,a26304a,a26305a,a26309a,a26310a,a26311a,a26315a,a26316a,a26320a,a26321a,a26322a,a26326a,a26327a,a26331a,a26332a,a26333a,a26337a,a26338a,a26342a,a26343a,a26344a,a26348a,a26349a,a26353a,a26354a,a26355a,a26359a,a26360a,a26364a,a26365a,a26366a,a26370a,a26371a,a26375a,a26376a,a26377a,a26381a,a26382a,a26386a,a26387a,a26388a,a26392a,a26393a,a26397a,a26398a,a26399a,a26403a,a26404a,a26408a,a26409a,a26410a,a26414a,a26415a,a26419a,a26420a,a26421a,a26425a,a26426a,a26430a,a26431a,a26432a,a26436a,a26437a,a26441a,a26442a,a26443a,a26447a,a26448a,a26452a,a26453a,a26454a,a26458a,a26459a,a26463a,a26464a,a26465a,a26469a,a26470a,a26474a,a26475a,a26476a,a26480a,a26481a,a26485a,a26486a,a26487a,a26491a,a26492a,a26496a,a26497a,a26498a,a26502a,a26503a,a26507a,a26508a,a26509a,a26513a,a26514a,a26518a,a26519a,a26520a,a26524a,a26525a,a26529a,a26530a,a26531a,a26535a,a26536a,a26540a,a26541a,a26542a,a26546a,a26547a,a26551a,a26552a,a26553a,a26557a,a26558a,a26562a,a26563a,a26564a,a26568a,a26569a,a26573a,a26574a,a26575a,a26579a,a26580a,a26584a,a26585a,a26586a,a26590a,a26591a,a26595a,a26596a,a26597a,a26601a,a26602a,a26606a,a26607a,a26608a,a26612a,a26613a,a26617a,a26618a,a26619a,a26623a,a26624a,a26628a,a26629a,a26630a,a26634a,a26635a,a26639a,a26640a,a26641a,a26645a,a26646a,a26650a,a26651a,a26652a,a26656a,a26657a,a26661a,a26662a,a26663a,a26667a,a26668a,a26672a,a26673a,a26674a,a26678a,a26679a,a26683a,a26684a,a26685a,a26689a,a26690a,a26694a,a26695a,a26696a,a26700a,a26701a,a26705a,a26706a,a26707a,a26711a,a26712a,a26716a,a26717a,a26718a,a26722a,a26723a,a26727a,a26728a,a26729a,a26733a,a26734a,a26738a,a26739a,a26740a,a26744a,a26745a,a26749a,a26750a,a26751a,a26755a,a26756a,a26760a,a26761a,a26762a,a26766a,a26767a,a26771a,a26772a,a26773a,a26777a,a26778a,a26782a,a26783a,a26784a,a26788a,a26789a,a26793a,a26794a,a26795a,a26799a,a26800a,a26804a,a26805a,a26806a,a26810a,a26811a,a26815a,a26816a,a26817a,a26821a,a26822a,a26826a,a26827a,a26828a,a26832a,a26833a,a26837a,a26838a,a26839a,a26843a,a26844a,a26848a,a26849a,a26850a,a26854a,a26855a,a26859a,a26860a,a26861a,a26865a,a26866a,a26870a,a26871a,a26872a,a26876a,a26877a,a26881a,a26882a,a26883a,a26887a,a26888a,a26892a,a26893a,a26894a,a26898a,a26899a,a26903a,a26904a,a26905a,a26909a,a26910a,a26914a,a26915a,a26916a,a26920a,a26921a,a26925a,a26926a,a26927a,a26931a,a26932a,a26936a,a26937a,a26938a,a26942a,a26943a,a26947a,a26948a,a26949a,a26953a,a26954a,a26958a,a26959a,a26960a,a26964a,a26965a,a26969a,a26970a,a26971a,a26975a,a26976a,a26980a,a26981a,a26982a,a26986a,a26987a,a26991a,a26992a,a26993a,a26997a,a26998a,a27002a,a27003a,a27004a,a27008a,a27009a,a27013a,a27014a,a27015a,a27019a,a27020a,a27024a,a27025a,a27026a,a27030a,a27031a,a27035a,a27036a,a27037a,a27041a,a27042a,a27046a,a27047a,a27048a,a27052a,a27053a,a27057a,a27058a,a27059a,a27063a,a27064a,a27068a,a27069a,a27070a,a27074a,a27075a,a27079a,a27080a,a27081a,a27085a,a27086a,a27090a,a27091a,a27092a,a27096a,a27097a,a27101a,a27102a,a27103a,a27107a,a27108a,a27112a,a27113a,a27114a,a27118a,a27119a,a27123a,a27124a,a27125a,a27129a,a27130a,a27134a,a27135a,a27136a,a27140a,a27141a,a27145a,a27146a,a27147a,a27151a,a27152a,a27156a,a27157a,a27158a,a27162a,a27163a,a27167a,a27168a,a27169a,a27173a,a27174a,a27178a,a27179a,a27180a,a27184a,a27185a,a27189a,a27190a,a27191a,a27195a,a27196a,a27200a,a27201a,a27202a,a27206a,a27207a,a27211a,a27212a,a27213a,a27217a,a27218a,a27222a,a27223a,a27224a,a27228a,a27229a,a27233a,a27234a,a27235a,a27239a,a27240a,a27244a,a27245a,a27246a,a27250a,a27251a,a27255a,a27256a,a27257a,a27261a,a27262a,a27266a,a27267a,a27268a,a27272a,a27273a,a27277a,a27278a,a27279a,a27283a,a27284a,a27288a,a27289a,a27290a,a27294a,a27295a,a27299a,a27300a,a27301a,a27305a,a27306a,a27310a,a27311a,a27312a,a27316a,a27317a,a27321a,a27322a,a27323a,a27327a,a27328a,a27332a,a27333a,a27334a,a27338a,a27339a,a27343a,a27344a,a27345a,a27349a,a27350a,a27354a,a27355a,a27356a,a27360a,a27361a,a27365a,a27366a,a27367a,a27371a,a27372a,a27376a,a27377a,a27378a,a27382a,a27383a,a27387a,a27388a,a27389a,a27393a,a27394a,a27398a,a27399a,a27400a,a27404a,a27405a,a27409a,a27410a,a27411a,a27415a,a27416a,a27420a,a27421a,a27422a,a27426a,a27427a,a27431a,a27432a,a27433a,a27437a,a27438a,a27442a,a27443a,a27444a,a27448a,a27449a,a27453a,a27454a,a27455a,a27459a,a27460a,a27464a,a27465a,a27466a,a27470a,a27471a,a27475a,a27476a,a27477a,a27481a,a27482a,a27486a,a27487a,a27488a,a27492a,a27493a,a27497a,a27498a,a27499a,a27503a,a27504a,a27508a,a27509a,a27510a,a27514a,a27515a,a27519a,a27520a,a27521a,a27525a,a27526a,a27530a,a27531a,a27532a,a27536a,a27537a,a27541a,a27542a,a27543a,a27547a,a27548a,a27552a,a27553a,a27554a,a27558a,a27559a,a27563a,a27564a,a27565a,a27569a,a27570a,a27574a,a27575a,a27576a,a27580a,a27581a,a27585a,a27586a,a27587a,a27591a,a27592a,a27596a,a27597a,a27598a,a27602a,a27603a,a27607a,a27608a,a27609a,a27613a,a27614a,a27618a,a27619a,a27620a,a27624a,a27625a,a27629a,a27630a,a27631a,a27635a,a27636a,a27640a,a27641a,a27642a,a27646a,a27647a,a27651a,a27652a,a27653a,a27657a,a27658a,a27662a,a27663a,a27664a,a27668a,a27669a,a27673a,a27674a,a27675a,a27679a,a27680a,a27684a,a27685a,a27686a,a27690a,a27691a,a27695a,a27696a,a27697a,a27701a,a27702a,a27706a,a27707a,a27708a,a27712a,a27713a,a27717a,a27718a,a27719a,a27723a,a27724a,a27728a,a27729a,a27730a,a27734a,a27735a,a27739a,a27740a,a27741a,a27745a,a27746a,a27750a,a27751a,a27752a,a27756a,a27757a,a27761a,a27762a,a27763a,a27767a,a27768a,a27772a,a27773a,a27774a,a27778a,a27779a,a27783a,a27784a,a27785a,a27789a,a27790a,a27794a,a27795a,a27796a,a27800a,a27801a,a27805a,a27806a,a27807a,a27811a,a27812a,a27816a,a27817a,a27818a,a27822a,a27823a,a27827a,a27828a,a27829a,a27833a,a27834a,a27838a,a27839a,a27840a,a27844a,a27845a,a27849a,a27850a,a27851a,a27855a,a27856a,a27860a,a27861a,a27862a,a27866a,a27867a,a27871a,a27872a,a27873a,a27877a,a27878a,a27882a,a27883a,a27884a,a27888a,a27889a,a27893a,a27894a,a27895a,a27899a,a27900a,a27904a,a27905a,a27906a,a27910a,a27911a,a27915a,a27916a,a27917a,a27921a,a27922a,a27926a,a27927a,a27928a,a27932a,a27933a,a27937a,a27938a,a27939a,a27943a,a27944a,a27948a,a27949a,a27950a,a27954a,a27955a,a27959a,a27960a,a27961a,a27965a,a27966a,a27970a,a27971a,a27972a,a27976a,a27977a,a27981a,a27982a,a27983a,a27987a,a27988a,a27992a,a27993a,a27994a,a27998a,a27999a,a28003a,a28004a,a28005a,a28009a,a28010a,a28014a,a28015a,a28016a,a28020a,a28021a,a28025a,a28026a,a28027a,a28031a,a28032a,a28036a,a28037a,a28038a,a28042a,a28043a,a28047a,a28048a,a28049a,a28053a,a28054a,a28058a,a28059a,a28060a,a28064a,a28065a,a28069a,a28070a,a28071a,a28075a,a28076a,a28080a,a28081a,a28082a,a28086a,a28087a,a28091a,a28092a,a28093a,a28097a,a28098a,a28102a,a28103a,a28104a,a28108a,a28109a,a28113a,a28114a,a28115a,a28119a,a28120a,a28124a,a28125a,a28126a,a28130a,a28131a,a28135a,a28136a,a28137a,a28141a,a28142a,a28146a,a28147a,a28148a,a28152a,a28153a,a28157a,a28158a,a28159a,a28163a,a28164a,a28168a,a28169a,a28170a,a28174a,a28175a,a28179a,a28180a,a28181a,a28185a,a28186a,a28190a,a28191a,a28192a,a28196a,a28197a,a28201a,a28202a,a28203a,a28207a,a28208a,a28212a,a28213a,a28214a,a28218a,a28219a,a28223a,a28224a,a28225a,a28229a,a28230a,a28234a,a28235a,a28236a,a28240a,a28241a,a28245a,a28246a,a28247a,a28251a,a28252a,a28256a,a28257a,a28258a,a28262a,a28263a,a28267a,a28268a,a28269a,a28273a,a28274a,a28278a,a28279a,a28280a,a28284a,a28285a,a28289a,a28290a,a28291a,a28295a,a28296a,a28300a,a28301a,a28302a,a28306a,a28307a,a28311a,a28312a,a28313a,a28317a,a28318a,a28322a,a28323a,a28324a,a28328a,a28329a,a28333a,a28334a,a28335a,a28339a,a28340a,a28344a,a28345a,a28346a,a28350a,a28351a,a28355a,a28356a,a28357a,a28361a,a28362a,a28366a,a28367a,a28368a,a28372a,a28373a,a28377a,a28378a,a28379a,a28383a,a28384a,a28388a,a28389a,a28390a,a28394a,a28395a,a28399a,a28400a,a28401a,a28405a,a28406a,a28410a,a28411a,a28412a,a28416a,a28417a,a28421a,a28422a,a28423a,a28427a,a28428a,a28432a,a28433a,a28434a,a28438a,a28439a,a28443a,a28444a,a28445a,a28449a,a28450a,a28454a,a28455a,a28456a,a28460a,a28461a,a28465a,a28466a,a28467a,a28471a,a28472a,a28476a,a28477a,a28478a,a28482a,a28483a,a28487a,a28488a,a28489a,a28493a,a28494a,a28498a,a28499a,a28500a,a28504a,a28505a,a28509a,a28510a,a28511a,a28515a,a28516a,a28520a,a28521a,a28522a,a28526a,a28527a,a28531a,a28532a,a28533a,a28537a,a28538a,a28542a,a28543a,a28544a,a28548a,a28549a,a28553a,a28554a,a28555a,a28559a,a28560a,a28564a,a28565a,a28566a,a28570a,a28571a,a28575a,a28576a,a28577a,a28581a,a28582a,a28586a,a28587a,a28588a,a28592a,a28593a,a28597a,a28598a,a28599a,a28603a,a28604a,a28608a,a28609a,a28610a,a28614a,a28615a,a28619a,a28620a,a28621a,a28625a,a28626a,a28630a,a28631a,a28632a,a28636a,a28637a,a28641a,a28642a,a28643a,a28647a,a28648a,a28652a,a28653a,a28654a,a28658a,a28659a,a28663a,a28664a,a28665a,a28669a,a28670a,a28674a,a28675a,a28676a,a28680a,a28681a,a28685a,a28686a,a28687a,a28691a,a28692a,a28696a,a28697a,a28698a,a28702a,a28703a,a28707a,a28708a,a28709a,a28713a,a28714a,a28718a,a28719a,a28720a,a28724a,a28725a,a28729a,a28730a,a28731a,a28735a,a28736a,a28740a,a28741a,a28742a,a28746a,a28747a,a28751a,a28752a,a28753a,a28757a,a28758a,a28762a,a28763a,a28764a,a28768a,a28769a,a28773a,a28774a,a28775a,a28779a,a28780a,a28784a,a28785a,a28786a,a28790a,a28791a,a28795a,a28796a,a28797a,a28801a,a28802a,a28806a,a28807a,a28808a,a28812a,a28813a,a28817a,a28818a,a28819a,a28823a,a28824a,a28828a,a28829a,a28830a,a28834a,a28835a,a28839a,a28840a,a28841a,a28845a,a28846a,a28850a,a28851a,a28852a,a28856a,a28857a,a28861a,a28862a,a28863a,a28867a,a28868a,a28872a,a28873a,a28874a,a28878a,a28879a,a28883a,a28884a,a28885a,a28889a,a28890a,a28894a,a28895a,a28896a,a28900a,a28901a,a28905a,a28906a,a28907a,a28911a,a28912a,a28916a,a28917a,a28918a,a28922a,a28923a,a28927a,a28928a,a28929a,a28933a,a28934a,a28938a,a28939a,a28940a,a28944a,a28945a,a28949a,a28950a,a28951a,a28955a,a28956a,a28960a,a28961a,a28962a,a28966a,a28967a,a28971a,a28972a,a28973a,a28977a,a28978a,a28982a,a28983a,a28984a,a28988a,a28989a,a28993a,a28994a,a28995a,a28999a,a29000a,a29004a,a29005a,a29006a,a29010a,a29011a,a29015a,a29016a,a29017a,a29021a,a29022a,a29026a,a29027a,a29028a,a29032a,a29033a,a29037a,a29038a,a29039a,a29043a,a29044a,a29048a,a29049a,a29050a,a29054a,a29055a,a29059a,a29060a,a29061a,a29065a,a29066a,a29070a,a29071a,a29072a,a29076a,a29077a,a29081a,a29082a,a29083a,a29087a,a29088a,a29092a,a29093a,a29094a,a29098a,a29099a,a29103a,a29104a,a29105a,a29109a,a29110a,a29114a,a29115a,a29116a,a29120a,a29121a,a29125a,a29126a,a29127a,a29131a,a29132a,a29136a,a29137a,a29138a,a29142a,a29143a,a29147a,a29148a,a29149a,a29153a,a29154a,a29158a,a29159a,a29160a,a29164a,a29165a,a29169a,a29170a,a29171a,a29175a,a29176a,a29180a,a29181a,a29182a,a29186a,a29187a,a29191a,a29192a,a29193a,a29197a,a29198a,a29202a,a29203a,a29204a,a29208a,a29209a,a29213a,a29214a,a29215a,a29219a,a29220a,a29224a,a29225a,a29226a,a29230a,a29231a,a29235a,a29236a,a29237a,a29241a,a29242a,a29246a,a29247a,a29248a,a29252a,a29253a,a29257a,a29258a,a29259a,a29263a,a29264a,a29268a,a29269a,a29270a,a29274a,a29275a,a29279a,a29280a,a29281a,a29285a,a29286a,a29290a,a29291a,a29292a,a29296a,a29297a,a29301a,a29302a,a29303a,a29307a,a29308a,a29312a,a29313a,a29314a,a29318a,a29319a,a29323a,a29324a,a29325a,a29329a,a29330a,a29334a,a29335a,a29336a,a29340a,a29341a,a29345a,a29346a,a29347a,a29351a,a29352a,a29356a,a29357a,a29358a,a29362a,a29363a,a29367a,a29368a,a29369a,a29373a,a29374a,a29378a,a29379a,a29380a,a29384a,a29385a,a29389a,a29390a,a29391a,a29395a,a29396a,a29400a,a29401a,a29402a,a29406a,a29407a,a29411a,a29412a,a29413a,a29417a,a29418a,a29422a,a29423a,a29424a,a29428a,a29429a,a29433a,a29434a,a29435a,a29439a,a29440a,a29444a,a29445a,a29446a,a29450a,a29451a,a29455a,a29456a,a29457a,a29461a,a29462a,a29466a,a29467a,a29468a,a29472a,a29473a,a29477a,a29478a,a29479a,a29483a,a29484a,a29488a,a29489a,a29490a,a29494a,a29495a,a29499a,a29500a,a29501a,a29505a,a29506a,a29510a,a29511a,a29512a,a29516a,a29517a,a29521a,a29522a,a29523a,a29527a,a29528a,a29532a,a29533a,a29534a,a29538a,a29539a,a29543a,a29544a,a29545a,a29549a,a29550a,a29554a,a29555a,a29556a,a29560a,a29561a,a29565a,a29566a,a29567a,a29571a,a29572a,a29576a,a29577a,a29578a,a29582a,a29583a,a29587a,a29588a,a29589a,a29593a,a29594a,a29598a,a29599a,a29600a,a29604a,a29605a,a29609a,a29610a,a29611a,a29615a,a29616a,a29620a,a29621a,a29622a,a29626a,a29627a,a29631a,a29632a,a29633a,a29637a,a29638a,a29642a,a29643a,a29644a,a29648a,a29649a,a29653a,a29654a,a29655a,a29659a,a29660a,a29664a,a29665a,a29666a,a29670a,a29671a,a29675a,a29676a,a29677a,a29681a,a29682a,a29686a,a29687a,a29688a,a29692a,a29693a,a29697a,a29698a,a29699a,a29703a,a29704a,a29708a,a29709a,a29710a,a29714a,a29715a,a29719a,a29720a,a29721a,a29725a,a29726a,a29730a,a29731a,a29732a,a29736a,a29737a,a29741a,a29742a,a29743a,a29747a,a29748a,a29752a,a29753a,a29754a,a29758a,a29759a,a29763a,a29764a,a29765a,a29769a,a29770a,a29774a,a29775a,a29776a,a29780a,a29781a,a29785a,a29786a,a29787a,a29791a,a29792a,a29796a,a29797a,a29798a,a29802a,a29803a,a29807a,a29808a,a29809a,a29813a,a29814a,a29818a,a29819a,a29820a,a29824a,a29825a,a29829a,a29830a,a29831a,a29835a,a29836a,a29840a,a29841a,a29842a,a29846a,a29847a,a29851a,a29852a,a29853a,a29857a,a29858a,a29862a,a29863a,a29864a,a29868a,a29869a,a29873a,a29874a,a29875a,a29879a,a29880a,a29884a,a29885a,a29886a,a29890a,a29891a,a29895a,a29896a,a29897a,a29901a,a29902a,a29906a,a29907a,a29908a,a29912a,a29913a,a29917a,a29918a,a29919a,a29923a,a29924a,a29928a,a29929a,a29930a,a29934a,a29935a,a29939a,a29940a,a29941a,a29945a,a29946a,a29950a,a29951a,a29952a,a29956a,a29957a,a29961a,a29962a,a29963a,a29967a,a29968a,a29972a,a29973a,a29974a,a29978a,a29979a,a29983a,a29984a,a29985a,a29989a,a29990a,a29994a,a29995a,a29996a,a30000a,a30001a,a30005a,a30006a,a30007a,a30011a,a30012a,a30016a,a30017a,a30018a,a30022a,a30023a,a30027a,a30028a,a30029a,a30033a,a30034a,a30038a,a30039a,a30040a,a30044a,a30045a,a30049a,a30050a,a30051a,a30055a,a30056a,a30060a,a30061a,a30062a,a30066a,a30067a,a30071a,a30072a,a30073a,a30077a,a30078a,a30082a,a30083a,a30084a,a30088a,a30089a,a30093a,a30094a,a30095a,a30099a,a30100a,a30104a,a30105a,a30106a,a30110a,a30111a,a30115a,a30116a,a30117a,a30121a,a30122a,a30126a,a30127a,a30128a,a30132a,a30133a,a30137a,a30138a,a30139a,a30143a,a30144a,a30148a,a30149a,a30150a,a30154a,a30155a,a30159a,a30160a,a30161a,a30165a,a30166a,a30170a,a30171a,a30172a,a30176a,a30177a,a30181a,a30182a,a30183a,a30187a,a30188a,a30192a,a30193a,a30194a,a30198a,a30199a,a30203a,a30204a,a30205a,a30209a,a30210a,a30214a,a30215a,a30216a,a30220a,a30221a,a30225a,a30226a,a30227a,a30231a,a30232a,a30236a,a30237a,a30238a,a30242a,a30243a,a30247a,a30248a,a30249a,a30253a,a30254a,a30258a,a30259a,a30260a,a30264a,a30265a,a30269a,a30270a,a30271a,a30275a,a30276a,a30280a,a30281a,a30282a,a30286a,a30287a,a30291a,a30292a,a30293a,a30297a,a30298a,a30302a,a30303a,a30304a,a30308a,a30309a,a30313a,a30314a,a30315a,a30319a,a30320a,a30324a,a30325a,a30326a,a30330a,a30331a,a30335a,a30336a,a30337a,a30341a,a30342a,a30346a,a30347a,a30348a,a30352a,a30353a,a30357a,a30358a,a30359a,a30363a,a30364a,a30368a,a30369a,a30370a,a30374a,a30375a,a30379a,a30380a,a30381a,a30385a,a30386a,a30390a,a30391a,a30392a,a30396a,a30397a,a30401a,a30402a,a30403a,a30407a,a30408a,a30412a,a30413a,a30414a,a30418a,a30419a,a30423a,a30424a,a30425a,a30429a,a30430a,a30434a,a30435a,a30436a,a30440a,a30441a,a30445a,a30446a,a30447a,a30451a,a30452a,a30456a,a30457a,a30458a,a30462a,a30463a,a30467a,a30468a,a30469a,a30473a,a30474a,a30478a,a30479a,a30480a,a30484a,a30485a,a30489a,a30490a,a30491a,a30495a,a30496a,a30500a,a30501a,a30502a,a30506a,a30507a,a30511a,a30512a,a30513a,a30517a,a30518a,a30522a,a30523a,a30524a,a30528a,a30529a,a30533a,a30534a,a30535a,a30539a,a30540a,a30544a,a30545a,a30546a,a30550a,a30551a,a30555a,a30556a,a30557a,a30561a,a30562a,a30566a,a30567a,a30568a,a30572a,a30573a,a30577a,a30578a,a30579a,a30583a,a30584a,a30588a,a30589a,a30590a,a30594a,a30595a,a30599a,a30600a,a30601a,a30605a,a30606a,a30610a,a30611a,a30612a,a30616a,a30617a,a30621a,a30622a,a30623a,a30627a,a30628a,a30632a,a30633a,a30634a,a30638a,a30639a,a30643a,a30644a,a30645a,a30649a,a30650a,a30654a,a30655a,a30656a,a30660a,a30661a,a30665a,a30666a,a30667a,a30671a,a30672a,a30676a,a30677a,a30678a,a30682a,a30683a,a30687a,a30688a,a30689a,a30693a,a30694a,a30698a,a30699a,a30700a,a30704a,a30705a,a30709a,a30710a,a30711a,a30715a,a30716a,a30720a,a30721a,a30722a,a30726a,a30727a,a30731a,a30732a,a30733a,a30737a,a30738a,a30742a,a30743a,a30744a,a30748a,a30749a,a30753a,a30754a,a30755a,a30759a,a30760a,a30764a,a30765a,a30766a,a30770a,a30771a,a30775a,a30776a,a30777a,a30781a,a30782a,a30786a,a30787a,a30788a,a30792a,a30793a,a30797a,a30798a,a30799a,a30803a,a30804a,a30808a,a30809a,a30810a,a30814a,a30815a,a30819a,a30820a,a30821a,a30825a,a30826a,a30830a,a30831a,a30832a,a30836a,a30837a,a30841a,a30842a,a30843a,a30847a,a30848a,a30852a,a30853a,a30854a,a30858a,a30859a,a30863a,a30864a,a30865a,a30869a,a30870a,a30874a,a30875a,a30876a,a30880a,a30881a,a30885a,a30886a,a30887a,a30891a,a30892a,a30896a,a30897a,a30898a,a30902a,a30903a,a30907a,a30908a,a30909a,a30913a,a30914a,a30918a,a30919a,a30920a,a30924a,a30925a,a30929a,a30930a,a30931a,a30935a,a30936a,a30940a,a30941a,a30942a,a30946a,a30947a,a30951a,a30952a,a30953a,a30957a,a30958a,a30962a,a30963a,a30964a,a30968a,a30969a,a30973a,a30974a,a30975a,a30979a,a30980a,a30984a,a30985a,a30986a,a30990a,a30991a,a30995a,a30996a,a30997a,a31001a,a31002a,a31006a,a31007a,a31008a,a31012a,a31013a,a31017a,a31018a,a31019a,a31023a,a31024a,a31028a,a31029a,a31030a,a31034a,a31035a,a31039a,a31040a,a31041a,a31045a,a31046a,a31050a,a31051a,a31052a,a31056a,a31057a,a31061a,a31062a,a31063a,a31067a,a31068a,a31072a,a31073a,a31074a,a31078a,a31079a,a31083a,a31084a,a31085a,a31089a,a31090a,a31094a,a31095a,a31096a,a31100a,a31101a,a31105a,a31106a,a31107a,a31111a,a31112a,a31116a,a31117a,a31118a,a31122a,a31123a,a31127a,a31128a,a31129a,a31133a,a31134a,a31138a,a31139a,a31140a,a31144a,a31145a,a31149a,a31150a,a31151a,a31155a,a31156a,a31160a,a31161a,a31162a,a31166a,a31167a,a31171a,a31172a,a31173a,a31177a,a31178a,a31182a,a31183a,a31184a,a31188a,a31189a,a31193a,a31194a,a31195a,a31199a,a31200a,a31204a,a31205a,a31206a,a31210a,a31211a,a31215a,a31216a,a31217a,a31221a,a31222a,a31226a,a31227a,a31228a,a31232a,a31233a,a31237a,a31238a,a31239a,a31243a,a31244a,a31248a,a31249a,a31250a,a31254a,a31255a,a31259a,a31260a,a31261a,a31265a,a31266a,a31270a,a31271a,a31272a,a31276a,a31277a,a31281a,a31282a,a31283a,a31287a,a31288a,a31292a,a31293a,a31294a,a31298a,a31299a,a31303a,a31304a,a31305a,a31309a,a31310a,a31314a,a31315a,a31316a,a31320a,a31321a,a31325a,a31326a,a31327a,a31331a,a31332a,a31336a,a31337a,a31338a,a31342a,a31343a,a31347a,a31348a,a31349a,a31353a,a31354a,a31358a,a31359a,a31360a,a31364a,a31365a,a31369a,a31370a,a31371a,a31375a,a31376a,a31380a,a31381a,a31382a,a31386a,a31387a,a31391a,a31392a,a31393a,a31397a,a31398a,a31402a,a31403a,a31404a,a31408a,a31409a,a31413a,a31414a,a31415a,a31419a,a31420a,a31424a,a31425a,a31426a,a31430a,a31431a,a31435a,a31436a,a31437a,a31441a,a31442a,a31446a,a31447a,a31448a,a31452a,a31453a,a31457a,a31458a,a31459a,a31463a,a31464a,a31468a,a31469a,a31470a,a31474a,a31475a,a31479a,a31480a,a31481a,a31485a,a31486a,a31490a,a31491a,a31492a,a31496a,a31497a,a31501a,a31502a,a31503a,a31507a,a31508a,a31512a,a31513a,a31514a,a31518a,a31519a,a31523a,a31524a,a31525a,a31529a,a31530a,a31534a,a31535a,a31536a,a31540a,a31541a,a31545a,a31546a,a31547a,a31551a,a31552a,a31556a,a31557a,a31558a,a31562a,a31563a,a31567a,a31568a,a31569a,a31573a,a31574a,a31578a,a31579a,a31580a,a31584a,a31585a,a31589a,a31590a,a31591a,a31595a,a31596a,a31600a,a31601a,a31602a,a31606a,a31607a,a31611a,a31612a,a31613a,a31617a,a31618a,a31622a,a31623a,a31624a,a31628a,a31629a,a31633a,a31634a,a31635a,a31639a,a31640a,a31644a,a31645a,a31646a,a31650a,a31651a,a31655a,a31656a,a31657a,a31661a,a31662a,a31666a,a31667a,a31668a,a31672a,a31673a,a31677a,a31678a,a31679a,a31683a,a31684a,a31688a,a31689a,a31690a,a31694a,a31695a,a31699a,a31700a,a31701a,a31705a,a31706a,a31710a,a31711a,a31712a,a31716a,a31717a,a31721a,a31722a,a31723a,a31727a,a31728a,a31732a,a31733a,a31734a,a31738a,a31739a,a31743a,a31744a,a31745a,a31749a,a31750a,a31754a,a31755a,a31756a,a31760a,a31761a,a31765a,a31766a,a31767a,a31771a,a31772a,a31776a,a31777a,a31778a,a31782a,a31783a,a31787a,a31788a,a31789a,a31793a,a31794a,a31798a,a31799a,a31800a,a31804a,a31805a,a31809a,a31810a,a31811a,a31815a,a31816a,a31820a,a31821a,a31822a,a31826a,a31827a,a31831a,a31832a,a31833a,a31837a,a31838a,a31842a,a31843a,a31844a,a31848a,a31849a,a31853a,a31854a,a31855a,a31859a,a31860a,a31864a,a31865a,a31866a,a31870a,a31871a,a31875a,a31876a,a31877a,a31881a,a31882a,a31886a,a31887a,a31888a,a31892a,a31893a,a31897a,a31898a,a31899a,a31903a,a31904a,a31908a,a31909a,a31910a,a31914a,a31915a,a31919a,a31920a,a31921a,a31925a,a31926a,a31930a,a31931a,a31932a,a31936a,a31937a,a31941a,a31942a,a31943a,a31947a,a31948a,a31952a,a31953a,a31954a,a31958a,a31959a,a31963a,a31964a,a31965a,a31969a,a31970a,a31974a,a31975a,a31976a,a31980a,a31981a,a31985a,a31986a,a31987a,a31991a,a31992a,a31996a,a31997a,a31998a,a32002a,a32003a,a32007a,a32008a,a32009a,a32013a,a32014a,a32018a,a32019a,a32020a,a32024a,a32025a,a32029a,a32030a,a32031a,a32035a,a32036a,a32040a,a32041a,a32042a,a32046a,a32047a,a32051a,a32052a,a32053a,a32057a,a32058a,a32062a,a32063a,a32064a,a32068a,a32069a,a32073a,a32074a,a32075a,a32079a,a32080a,a32084a,a32085a,a32086a,a32090a,a32091a,a32095a,a32096a,a32097a,a32101a,a32102a,a32106a,a32107a,a32108a,a32112a,a32113a,a32117a,a32118a,a32119a,a32123a,a32124a,a32128a,a32129a,a32130a,a32134a,a32135a,a32139a,a32140a,a32141a,a32145a,a32146a,a32150a,a32151a,a32152a,a32156a,a32157a,a32161a,a32162a,a32163a,a32167a,a32168a,a32172a,a32173a,a32174a,a32178a,a32179a,a32183a,a32184a,a32185a,a32189a,a32190a,a32194a,a32195a,a32196a,a32200a,a32201a,a32205a,a32206a,a32207a,a32211a,a32212a,a32216a,a32217a,a32218a,a32222a,a32223a,a32227a,a32228a,a32229a,a32233a,a32234a,a32238a,a32239a,a32240a,a32244a,a32245a,a32249a,a32250a,a32251a,a32255a,a32256a,a32260a,a32261a,a32262a,a32266a,a32267a,a32271a,a32272a,a32273a,a32277a,a32278a,a32282a,a32283a,a32284a,a32288a,a32289a,a32293a,a32294a,a32295a,a32299a,a32300a,a32304a,a32305a,a32306a,a32310a,a32311a,a32315a,a32316a,a32317a,a32321a,a32322a,a32326a,a32327a,a32328a,a32332a,a32333a,a32337a,a32338a,a32339a,a32343a,a32344a,a32348a,a32349a,a32350a,a32354a,a32355a,a32359a,a32360a,a32361a,a32365a,a32366a,a32370a,a32371a,a32372a,a32376a,a32377a,a32381a,a32382a,a32383a,a32387a,a32388a,a32392a,a32393a,a32394a,a32398a,a32399a,a32403a,a32404a,a32405a,a32409a,a32410a,a32414a,a32415a,a32416a,a32420a,a32421a,a32425a,a32426a,a32427a,a32431a,a32432a,a32436a,a32437a,a32438a,a32442a,a32443a,a32447a,a32448a,a32449a,a32453a,a32454a,a32458a,a32459a,a32460a,a32464a,a32465a,a32469a,a32470a,a32471a,a32475a,a32476a,a32480a,a32481a,a32482a,a32486a,a32487a,a32491a,a32492a,a32493a,a32497a,a32498a,a32502a,a32503a,a32504a,a32508a,a32509a,a32513a,a32514a,a32515a,a32519a,a32520a,a32524a,a32525a,a32526a,a32530a,a32531a,a32535a,a32536a,a32537a,a32541a,a32542a,a32546a,a32547a,a32548a,a32552a,a32553a,a32557a,a32558a,a32559a,a32563a,a32564a,a32568a,a32569a,a32570a,a32574a,a32575a,a32579a,a32580a,a32581a,a32585a,a32586a,a32590a,a32591a,a32592a,a32596a,a32597a,a32601a,a32602a,a32603a,a32607a,a32608a,a32612a,a32613a,a32614a,a32618a,a32619a,a32623a,a32624a,a32625a,a32629a,a32630a,a32634a,a32635a,a32636a,a32640a,a32641a,a32645a,a32646a,a32647a,a32651a,a32652a,a32656a,a32657a,a32658a,a32662a,a32663a,a32667a,a32668a,a32669a,a32673a,a32674a,a32678a,a32679a,a32680a,a32684a,a32685a,a32689a,a32690a,a32691a,a32695a,a32696a,a32700a,a32701a,a32702a,a32706a,a32707a,a32711a,a32712a,a32713a,a32717a,a32718a,a32722a,a32723a,a32724a,a32728a,a32729a,a32733a,a32734a,a32735a,a32739a,a32740a,a32744a,a32745a,a32746a,a32750a,a32751a,a32755a,a32756a,a32757a,a32761a,a32762a,a32766a,a32767a,a32768a,a32772a,a32773a,a32777a,a32778a,a32779a,a32783a,a32784a,a32788a,a32789a,a32790a,a32794a,a32795a,a32799a,a32800a,a32801a,a32805a,a32806a,a32810a,a32811a,a32812a,a32816a,a32817a,a32821a,a32822a,a32823a,a32827a,a32828a,a32832a,a32833a,a32834a,a32838a,a32839a,a32843a,a32844a,a32845a,a32849a,a32850a,a32854a,a32855a,a32856a,a32860a,a32861a,a32865a,a32866a,a32867a,a32871a,a32872a,a32876a,a32877a,a32878a,a32882a,a32883a,a32887a,a32888a,a32889a,a32893a,a32894a,a32898a,a32899a,a32900a,a32904a,a32905a,a32909a,a32910a,a32911a,a32915a,a32916a,a32920a,a32921a,a32922a,a32926a,a32927a,a32931a,a32932a,a32933a,a32937a,a32938a,a32942a,a32943a,a32944a,a32948a,a32949a,a32953a,a32954a,a32955a,a32959a,a32960a,a32964a,a32965a,a32966a,a32970a,a32971a,a32975a,a32976a,a32977a,a32981a,a32982a,a32986a,a32987a,a32988a,a32992a,a32993a,a32997a,a32998a,a32999a,a33003a,a33004a,a33008a,a33009a,a33010a,a33014a,a33015a,a33019a,a33020a,a33021a,a33025a,a33026a,a33030a,a33031a,a33032a,a33036a,a33037a,a33041a,a33042a,a33043a,a33047a,a33048a,a33052a,a33053a,a33054a,a33058a,a33059a,a33063a,a33064a,a33065a,a33069a,a33070a,a33074a,a33075a,a33076a,a33080a,a33081a,a33085a,a33086a,a33087a,a33091a,a33092a,a33096a,a33097a,a33098a,a33102a,a33103a,a33107a,a33108a,a33109a,a33113a,a33114a,a33118a,a33119a,a33120a,a33124a,a33125a,a33129a,a33130a,a33131a,a33135a,a33136a,a33140a,a33141a,a33142a,a33146a,a33147a,a33151a,a33152a,a33153a,a33157a,a33158a,a33162a,a33163a,a33164a,a33168a,a33169a,a33173a,a33174a,a33175a,a33179a,a33180a,a33184a,a33185a,a33186a,a33190a,a33191a,a33195a,a33196a,a33197a,a33201a,a33202a,a33206a,a33207a,a33208a,a33212a,a33213a,a33217a,a33218a,a33219a,a33223a,a33224a,a33228a,a33229a,a33230a,a33234a,a33235a,a33239a,a33240a,a33241a,a33245a,a33246a,a33250a,a33251a,a33252a,a33256a,a33257a,a33261a,a33262a,a33263a,a33267a,a33268a,a33272a,a33273a,a33274a,a33278a,a33279a,a33283a,a33284a,a33285a,a33289a,a33290a,a33294a,a33295a,a33296a,a33300a,a33301a,a33305a,a33306a,a33307a,a33311a,a33312a,a33316a,a33317a,a33318a,a33322a,a33323a,a33327a,a33328a,a33329a,a33333a,a33334a,a33338a,a33339a,a33340a,a33344a,a33345a,a33349a,a33350a,a33351a,a33355a,a33356a,a33360a,a33361a,a33362a,a33366a,a33367a,a33371a,a33372a,a33373a,a33377a,a33378a,a33382a,a33383a,a33384a,a33388a,a33389a,a33393a,a33394a,a33395a,a33399a,a33400a,a33404a,a33405a,a33406a,a33410a,a33411a,a33415a,a33416a,a33417a,a33421a,a33422a,a33426a,a33427a,a33428a,a33432a,a33433a,a33437a,a33438a,a33439a,a33443a,a33444a,a33448a,a33449a,a33450a,a33454a,a33455a,a33459a,a33460a,a33461a,a33465a,a33466a,a33470a,a33471a,a33472a,a33476a,a33477a,a33481a,a33482a,a33483a,a33487a,a33488a,a33492a,a33493a,a33494a,a33498a,a33499a,a33503a,a33504a,a33505a,a33509a,a33510a,a33514a,a33515a,a33516a,a33520a,a33521a,a33525a,a33526a,a33527a,a33531a,a33532a,a33536a,a33537a,a33538a,a33542a,a33543a,a33547a,a33548a,a33549a,a33553a,a33554a,a33558a,a33559a,a33560a,a33564a,a33565a,a33569a,a33570a,a33571a,a33575a,a33576a,a33580a,a33581a,a33582a,a33586a,a33587a,a33591a,a33592a,a33593a,a33597a,a33598a,a33602a,a33603a,a33604a,a33608a,a33609a,a33613a,a33614a,a33615a,a33619a,a33620a,a33624a,a33625a,a33626a,a33630a,a33631a,a33635a,a33636a,a33637a,a33641a,a33642a,a33646a,a33647a,a33648a,a33652a,a33653a,a33657a,a33658a,a33659a,a33663a,a33664a,a33668a,a33669a,a33670a,a33674a,a33675a,a33679a,a33680a,a33681a,a33685a,a33686a,a33690a,a33691a,a33692a,a33696a,a33697a,a33701a,a33702a,a33703a,a33707a,a33708a,a33712a,a33713a,a33714a,a33718a,a33719a,a33723a,a33724a,a33725a,a33729a,a33730a,a33734a,a33735a,a33736a,a33740a,a33741a,a33745a,a33746a,a33747a,a33751a,a33752a,a33756a,a33757a,a33758a,a33762a,a33763a,a33767a,a33768a,a33769a,a33773a,a33774a,a33778a,a33779a,a33780a,a33784a,a33785a,a33789a,a33790a,a33791a,a33795a,a33796a,a33800a,a33801a,a33802a,a33806a,a33807a,a33811a,a33812a,a33813a,a33817a,a33818a,a33822a,a33823a,a33824a,a33828a,a33829a,a33833a,a33834a,a33835a,a33839a,a33840a,a33844a,a33845a,a33846a,a33850a,a33851a,a33855a,a33856a,a33857a,a33861a,a33862a,a33866a,a33867a,a33868a,a33872a,a33873a,a33877a,a33878a,a33879a,a33883a,a33884a,a33888a,a33889a,a33890a,a33894a,a33895a,a33899a,a33900a,a33901a,a33905a,a33906a,a33910a,a33911a,a33912a,a33916a,a33917a,a33921a,a33922a,a33923a,a33927a,a33928a,a33932a,a33933a,a33934a,a33938a,a33939a,a33943a,a33944a,a33945a,a33949a,a33950a,a33954a,a33955a,a33956a,a33960a,a33961a,a33965a,a33966a,a33967a,a33971a,a33972a,a33976a,a33977a,a33978a,a33982a,a33983a,a33987a,a33988a,a33989a,a33993a,a33994a,a33998a,a33999a,a34000a,a34004a,a34005a,a34009a,a34010a,a34011a,a34015a,a34016a,a34020a,a34021a,a34022a,a34026a,a34027a,a34031a,a34032a,a34033a,a34037a,a34038a,a34042a,a34043a,a34044a,a34048a,a34049a,a34053a,a34054a,a34055a,a34059a,a34060a,a34064a,a34065a,a34066a,a34070a,a34071a,a34075a,a34076a,a34077a,a34081a,a34082a,a34086a,a34087a,a34088a,a34092a,a34093a,a34097a,a34098a,a34099a,a34103a,a34104a,a34108a,a34109a,a34110a,a34114a,a34115a,a34119a,a34120a,a34121a,a34125a,a34126a,a34130a,a34131a,a34132a,a34136a,a34137a,a34141a,a34142a,a34143a,a34147a,a34148a,a34152a,a34153a,a34154a,a34158a,a34159a,a34163a,a34164a,a34165a,a34169a,a34170a,a34174a,a34175a,a34176a,a34180a,a34181a,a34185a,a34186a,a34187a,a34191a,a34192a,a34196a,a34197a,a34198a,a34202a,a34203a,a34207a,a34208a,a34209a,a34213a,a34214a,a34218a,a34219a,a34220a,a34224a,a34225a,a34229a,a34230a,a34231a,a34235a,a34236a,a34240a,a34241a,a34242a,a34246a,a34247a,a34251a,a34252a,a34253a,a34257a,a34258a,a34262a,a34263a,a34264a,a34268a,a34269a,a34273a,a34274a,a34275a,a34279a,a34280a,a34284a,a34285a,a34286a,a34290a,a34291a,a34295a,a34296a,a34297a,a34301a,a34302a,a34306a,a34307a,a34308a,a34312a,a34313a,a34317a,a34318a,a34319a,a34323a,a34324a,a34328a,a34329a,a34330a,a34334a,a34335a,a34339a,a34340a,a34341a,a34345a,a34346a,a34350a,a34351a,a34352a,a34356a,a34357a,a34361a,a34362a,a34363a,a34367a,a34368a,a34372a,a34373a,a34374a,a34378a,a34379a,a34383a,a34384a,a34385a,a34389a,a34390a,a34394a,a34395a,a34396a,a34400a,a34401a,a34405a,a34406a,a34407a,a34411a,a34412a,a34416a,a34417a,a34418a,a34422a,a34423a,a34427a,a34428a,a34429a,a34433a,a34434a,a34438a,a34439a,a34440a,a34444a,a34445a,a34449a,a34450a,a34451a,a34455a,a34456a,a34460a,a34461a,a34462a,a34466a,a34467a,a34471a,a34472a,a34473a,a34477a,a34478a,a34482a,a34483a,a34484a,a34488a,a34489a,a34493a,a34494a,a34495a,a34499a,a34500a,a34504a,a34505a,a34506a,a34510a,a34511a,a34515a,a34516a,a34517a,a34521a,a34522a,a34526a,a34527a,a34528a,a34532a,a34533a,a34537a,a34538a,a34539a,a34543a,a34544a,a34548a,a34549a,a34550a,a34554a,a34555a,a34559a,a34560a,a34561a,a34565a,a34566a,a34570a,a34571a,a34572a,a34576a,a34577a,a34581a,a34582a,a34583a,a34587a,a34588a,a34592a,a34593a,a34594a,a34598a,a34599a,a34603a,a34604a,a34605a,a34609a,a34610a,a34614a,a34615a,a34616a,a34620a,a34621a,a34625a,a34626a,a34627a,a34631a,a34632a,a34636a,a34637a,a34638a,a34642a,a34643a,a34647a,a34648a,a34649a,a34653a,a34654a,a34658a,a34659a,a34660a,a34664a,a34665a,a34669a,a34670a,a34671a,a34675a,a34676a,a34680a,a34681a,a34682a,a34686a,a34687a,a34691a,a34692a,a34693a,a34697a,a34698a,a34702a,a34703a,a34704a,a34708a,a34709a,a34713a,a34714a,a34715a,a34719a,a34720a,a34724a,a34725a,a34726a,a34730a,a34731a,a34735a,a34736a,a34737a,a34741a,a34742a,a34746a,a34747a,a34748a,a34752a,a34753a,a34757a,a34758a,a34759a,a34763a,a34764a,a34768a,a34769a,a34770a,a34774a,a34775a,a34779a,a34780a,a34781a,a34785a,a34786a,a34790a,a34791a,a34792a,a34796a,a34797a,a34801a,a34802a,a34803a,a34807a,a34808a,a34812a,a34813a,a34814a,a34818a,a34819a,a34823a,a34824a,a34825a,a34829a,a34830a,a34834a,a34835a,a34836a,a34840a,a34841a,a34845a,a34846a,a34847a,a34851a,a34852a,a34856a,a34857a,a34858a,a34862a,a34863a,a34867a,a34868a,a34869a,a34873a,a34874a,a34878a,a34879a,a34880a,a34884a,a34885a,a34889a,a34890a,a34891a,a34895a,a34896a,a34900a,a34901a,a34902a,a34906a,a34907a,a34911a,a34912a,a34913a,a34917a,a34918a,a34922a,a34923a,a34924a,a34928a,a34929a,a34933a,a34934a,a34935a,a34939a,a34940a,a34944a,a34945a,a34946a,a34950a,a34951a,a34955a,a34956a,a34957a,a34961a,a34962a,a34966a,a34967a,a34968a,a34972a,a34973a,a34977a,a34978a,a34979a,a34983a,a34984a,a34988a,a34989a,a34990a,a34994a,a34995a,a34999a,a35000a,a35001a,a35005a,a35006a,a35010a,a35011a,a35012a,a35016a,a35017a,a35021a,a35022a,a35023a,a35027a,a35028a,a35032a,a35033a,a35034a,a35038a,a35039a,a35043a,a35044a,a35045a,a35049a,a35050a,a35054a,a35055a,a35056a,a35060a,a35061a,a35065a,a35066a,a35067a,a35071a,a35072a,a35076a,a35077a,a35078a,a35082a,a35083a,a35087a,a35088a,a35089a,a35093a,a35094a,a35098a,a35099a,a35100a,a35104a,a35105a,a35109a,a35110a,a35111a,a35115a,a35116a,a35120a,a35121a,a35122a,a35126a,a35127a,a35131a,a35132a,a35133a,a35137a,a35138a,a35142a,a35143a,a35144a,a35148a,a35149a,a35153a,a35154a,a35155a,a35159a,a35160a,a35164a,a35165a,a35166a,a35170a,a35171a,a35175a,a35176a,a35177a,a35181a,a35182a,a35186a,a35187a,a35188a,a35192a,a35193a,a35197a,a35198a,a35199a,a35203a,a35204a,a35208a,a35209a,a35210a,a35214a,a35215a,a35219a,a35220a,a35221a,a35225a,a35226a,a35230a,a35231a,a35232a,a35236a,a35237a,a35241a,a35242a,a35243a,a35247a,a35248a,a35252a,a35253a,a35254a,a35258a,a35259a,a35263a,a35264a,a35265a,a35269a,a35270a,a35274a,a35275a,a35276a,a35280a,a35281a,a35285a,a35286a,a35287a,a35291a,a35292a,a35296a,a35297a,a35298a,a35302a,a35303a,a35307a,a35308a,a35309a,a35313a,a35314a,a35318a,a35319a,a35320a,a35324a,a35325a,a35329a,a35330a,a35331a,a35335a,a35336a,a35340a,a35341a,a35342a,a35346a,a35347a,a35351a,a35352a,a35353a,a35357a,a35358a,a35362a,a35363a,a35364a,a35368a,a35369a,a35373a,a35374a,a35375a,a35379a,a35380a,a35384a,a35385a,a35386a,a35390a,a35391a,a35395a,a35396a,a35397a,a35401a,a35402a,a35406a,a35407a,a35408a,a35412a,a35413a,a35417a,a35418a,a35419a,a35423a,a35424a,a35428a,a35429a,a35430a,a35434a,a35435a,a35439a,a35440a,a35441a,a35445a,a35446a,a35450a,a35451a,a35452a,a35456a,a35457a,a35461a,a35462a,a35463a,a35467a,a35468a,a35472a,a35473a,a35474a,a35478a,a35479a,a35483a,a35484a,a35485a,a35489a,a35490a,a35494a,a35495a,a35496a,a35500a,a35501a,a35505a,a35506a,a35507a,a35511a,a35512a,a35516a,a35517a,a35518a,a35522a,a35523a,a35527a,a35528a,a35529a,a35533a,a35534a,a35538a,a35539a,a35540a,a35544a,a35545a,a35549a,a35550a,a35551a,a35555a,a35556a,a35560a,a35561a,a35562a,a35566a,a35567a,a35571a,a35572a,a35573a,a35577a,a35578a,a35582a,a35583a,a35584a,a35588a,a35589a,a35593a,a35594a,a35595a,a35599a,a35600a,a35604a,a35605a,a35606a,a35610a,a35611a,a35615a,a35616a,a35617a,a35621a,a35622a,a35626a,a35627a,a35628a,a35632a,a35633a,a35637a,a35638a,a35639a,a35643a,a35644a,a35648a,a35649a,a35650a,a35654a,a35655a,a35659a,a35660a,a35661a,a35665a,a35666a,a35670a,a35671a,a35672a,a35676a,a35677a,a35681a,a35682a,a35683a,a35687a,a35688a,a35692a,a35693a,a35694a,a35698a,a35699a,a35703a,a35704a,a35705a,a35709a,a35710a,a35714a,a35715a,a35716a,a35720a,a35721a,a35725a,a35726a,a35727a,a35731a,a35732a,a35736a,a35737a,a35738a,a35742a,a35743a,a35747a,a35748a,a35749a,a35753a,a35754a,a35758a,a35759a,a35760a,a35764a,a35765a,a35769a,a35770a,a35771a,a35775a,a35776a,a35780a,a35781a,a35782a,a35786a,a35787a,a35791a,a35792a,a35793a,a35797a,a35798a,a35802a,a35803a,a35804a,a35808a,a35809a,a35813a,a35814a,a35815a,a35819a,a35820a,a35824a,a35825a,a35826a,a35830a,a35831a,a35835a,a35836a,a35837a,a35841a,a35842a,a35846a,a35847a,a35848a,a35852a,a35853a,a35857a,a35858a,a35859a,a35863a,a35864a,a35868a,a35869a,a35870a,a35874a,a35875a,a35879a,a35880a,a35881a,a35885a,a35886a,a35890a,a35891a,a35892a,a35896a,a35897a,a35901a,a35902a,a35903a,a35907a,a35908a,a35912a,a35913a,a35914a,a35918a,a35919a,a35923a,a35924a,a35925a,a35929a,a35930a,a35934a,a35935a,a35936a,a35940a,a35941a,a35945a,a35946a,a35947a,a35951a,a35952a,a35956a,a35957a,a35958a,a35962a,a35963a,a35967a,a35968a,a35969a,a35973a,a35974a,a35978a,a35979a,a35980a,a35984a,a35985a,a35989a,a35990a,a35991a,a35995a,a35996a,a36000a,a36001a,a36002a,a36006a,a36007a,a36011a,a36012a,a36013a,a36017a,a36018a,a36022a,a36023a,a36024a,a36028a,a36029a,a36033a,a36034a,a36035a,a36039a,a36040a,a36044a,a36045a,a36046a,a36050a,a36051a,a36055a,a36056a,a36057a,a36061a,a36062a,a36066a,a36067a,a36068a,a36072a,a36073a,a36077a,a36078a,a36079a,a36083a,a36084a,a36088a,a36089a,a36090a,a36094a,a36095a,a36099a,a36100a,a36101a,a36105a,a36106a,a36110a,a36111a,a36112a,a36116a,a36117a,a36121a,a36122a,a36123a,a36127a,a36128a,a36132a,a36133a,a36134a,a36138a,a36139a,a36143a,a36144a,a36145a,a36149a,a36150a,a36154a,a36155a,a36156a,a36160a,a36161a,a36165a,a36166a,a36167a,a36171a,a36172a,a36176a,a36177a,a36178a,a36182a,a36183a,a36187a,a36188a,a36189a,a36193a,a36194a,a36198a,a36199a,a36200a,a36204a,a36205a,a36209a,a36210a,a36211a,a36215a,a36216a,a36220a,a36221a,a36222a,a36226a,a36227a,a36231a,a36232a,a36233a,a36237a,a36238a,a36242a,a36243a,a36244a,a36248a,a36249a,a36253a,a36254a,a36255a,a36259a,a36260a,a36264a,a36265a,a36266a,a36270a,a36271a,a36275a,a36276a,a36277a,a36281a,a36282a,a36286a,a36287a,a36288a,a36292a,a36293a,a36297a,a36298a,a36299a,a36303a,a36304a,a36308a,a36309a,a36310a,a36314a,a36315a,a36319a,a36320a,a36321a,a36325a,a36326a,a36330a,a36331a,a36332a,a36336a,a36337a,a36341a,a36342a,a36343a,a36347a,a36348a,a36352a,a36353a,a36354a,a36358a,a36359a,a36363a,a36364a,a36365a,a36369a,a36370a,a36374a,a36375a,a36376a,a36380a,a36381a,a36385a,a36386a,a36387a,a36391a,a36392a,a36396a,a36397a,a36398a,a36402a,a36403a,a36407a,a36408a,a36409a,a36413a,a36414a,a36418a,a36419a,a36420a,a36424a,a36425a,a36429a,a36430a,a36431a,a36435a,a36436a,a36440a,a36441a,a36442a,a36446a,a36447a,a36451a,a36452a,a36453a,a36457a,a36458a,a36462a,a36463a,a36464a,a36468a,a36469a,a36473a,a36474a,a36475a,a36479a,a36480a,a36484a,a36485a,a36486a,a36490a,a36491a,a36495a,a36496a,a36497a,a36501a,a36502a,a36506a,a36507a,a36508a,a36512a,a36513a,a36517a,a36518a,a36519a,a36523a,a36524a,a36528a,a36529a,a36530a,a36534a,a36535a,a36539a,a36540a,a36541a,a36545a,a36546a,a36550a,a36551a,a36552a,a36556a,a36557a,a36561a,a36562a,a36563a,a36567a,a36568a,a36572a,a36573a,a36574a,a36578a,a36579a,a36583a,a36584a,a36585a,a36589a,a36590a,a36594a,a36595a,a36596a,a36600a,a36601a,a36605a,a36606a,a36607a,a36611a,a36612a,a36616a,a36617a,a36618a,a36622a,a36623a,a36627a,a36628a,a36629a,a36633a,a36634a,a36638a,a36639a,a36640a,a36644a,a36645a,a36649a,a36650a,a36651a,a36655a,a36656a,a36660a,a36661a,a36662a,a36666a,a36667a,a36671a,a36672a,a36673a,a36677a,a36678a,a36682a,a36683a,a36684a,a36688a,a36689a,a36693a,a36694a,a36695a,a36699a,a36700a,a36704a,a36705a,a36706a,a36710a,a36711a,a36715a,a36716a,a36717a,a36721a,a36722a,a36726a,a36727a,a36728a,a36732a,a36733a,a36737a,a36738a,a36739a,a36743a,a36744a,a36748a,a36749a,a36750a,a36754a,a36755a,a36759a,a36760a,a36761a,a36765a,a36766a,a36770a,a36771a,a36772a,a36776a,a36777a,a36781a,a36782a,a36783a,a36787a,a36788a,a36792a,a36793a,a36794a,a36798a,a36799a,a36803a,a36804a,a36805a,a36809a,a36810a,a36814a,a36815a,a36816a,a36820a,a36821a,a36825a,a36826a,a36827a,a36831a,a36832a,a36836a,a36837a,a36838a,a36842a,a36843a,a36847a,a36848a,a36849a,a36853a,a36854a,a36858a,a36859a,a36860a,a36864a,a36865a,a36869a,a36870a,a36871a,a36875a,a36876a,a36880a,a36881a,a36882a,a36886a,a36887a,a36891a,a36892a,a36893a,a36897a,a36898a,a36902a,a36903a,a36904a,a36908a,a36909a,a36913a,a36914a,a36915a,a36919a,a36920a,a36924a,a36925a,a36926a,a36930a,a36931a,a36935a,a36936a,a36937a,a36941a,a36942a,a36946a,a36947a,a36948a,a36952a,a36953a,a36957a,a36958a,a36959a,a36963a,a36964a,a36968a,a36969a,a36970a,a36974a,a36975a,a36979a,a36980a,a36981a,a36985a,a36986a,a36990a,a36991a,a36992a,a36996a,a36997a,a37001a,a37002a,a37003a,a37007a,a37008a,a37012a,a37013a,a37014a,a37018a,a37019a,a37023a,a37024a,a37025a,a37029a,a37030a,a37034a,a37035a,a37036a,a37040a,a37041a,a37045a,a37046a,a37047a,a37051a,a37052a,a37056a,a37057a,a37058a,a37062a,a37063a,a37067a,a37068a,a37069a,a37073a,a37074a,a37078a,a37079a,a37080a,a37084a,a37085a,a37089a,a37090a,a37091a,a37095a,a37096a,a37100a,a37101a,a37102a,a37106a,a37107a,a37111a,a37112a,a37113a,a37117a,a37118a,a37122a,a37123a,a37124a,a37128a,a37129a,a37133a,a37134a,a37135a,a37139a,a37140a,a37144a,a37145a,a37146a,a37150a,a37151a,a37155a,a37156a,a37157a,a37161a,a37162a,a37166a,a37167a,a37168a,a37172a,a37173a,a37177a,a37178a,a37179a,a37183a,a37184a,a37188a,a37189a,a37190a,a37194a,a37195a,a37199a,a37200a,a37201a,a37205a,a37206a,a37210a,a37211a,a37212a,a37216a,a37217a,a37221a,a37222a,a37223a,a37227a,a37228a,a37232a,a37233a,a37234a,a37238a,a37239a,a37243a,a37244a,a37245a,a37249a,a37250a,a37254a,a37255a,a37256a,a37260a,a37261a,a37265a,a37266a,a37267a,a37271a,a37272a,a37276a,a37277a,a37278a,a37282a,a37283a,a37287a,a37288a,a37289a,a37293a,a37294a,a37298a,a37299a,a37300a,a37304a,a37305a,a37309a,a37310a,a37311a,a37315a,a37316a,a37320a,a37321a,a37322a,a37326a,a37327a,a37331a,a37332a,a37333a,a37337a,a37338a,a37342a,a37343a,a37344a,a37348a,a37349a,a37353a,a37354a,a37355a,a37359a,a37360a,a37364a,a37365a,a37366a,a37370a,a37371a,a37375a,a37376a,a37377a,a37381a,a37382a,a37386a,a37387a,a37388a,a37392a,a37393a,a37397a,a37398a,a37399a,a37403a,a37404a,a37408a,a37409a,a37410a,a37414a,a37415a,a37419a,a37420a,a37421a,a37425a,a37426a,a37430a,a37431a,a37432a,a37436a,a37437a,a37441a,a37442a,a37443a,a37447a,a37448a,a37452a,a37453a,a37454a,a37458a,a37459a,a37463a,a37464a,a37465a,a37469a,a37470a,a37474a,a37475a,a37476a,a37480a,a37481a,a37485a,a37486a,a37487a,a37491a,a37492a,a37496a,a37497a,a37498a,a37502a,a37503a,a37507a,a37508a,a37509a,a37513a,a37514a,a37518a,a37519a,a37520a,a37524a,a37525a,a37529a,a37530a,a37531a,a37535a,a37536a,a37540a,a37541a,a37542a,a37546a,a37547a,a37551a,a37552a,a37553a,a37557a,a37558a,a37562a,a37563a,a37564a,a37568a,a37569a,a37573a,a37574a,a37575a,a37579a,a37580a,a37584a,a37585a,a37586a,a37590a,a37591a,a37595a,a37596a,a37597a,a37601a,a37602a,a37606a,a37607a,a37608a,a37612a,a37613a,a37617a,a37618a,a37619a,a37623a,a37624a,a37628a,a37629a,a37630a,a37634a,a37635a,a37639a,a37640a,a37641a,a37645a,a37646a,a37650a,a37651a,a37652a,a37656a,a37657a,a37661a,a37662a,a37663a,a37667a,a37668a,a37672a,a37673a,a37674a,a37678a,a37679a,a37683a,a37684a,a37685a,a37689a,a37690a,a37694a,a37695a,a37696a,a37700a,a37701a,a37705a,a37706a,a37707a,a37711a,a37712a,a37716a,a37717a,a37718a,a37722a,a37723a,a37727a,a37728a,a37729a,a37733a,a37734a,a37738a,a37739a,a37740a,a37744a,a37745a,a37749a,a37750a,a37751a,a37755a,a37756a,a37760a,a37761a,a37762a,a37766a,a37767a,a37771a,a37772a,a37773a,a37777a,a37778a,a37782a,a37783a,a37784a,a37788a,a37789a,a37793a,a37794a,a37795a,a37799a,a37800a,a37804a,a37805a,a37806a,a37810a,a37811a,a37815a,a37816a,a37817a,a37821a,a37822a,a37826a,a37827a,a37828a,a37832a,a37833a,a37837a,a37838a,a37839a,a37843a,a37844a,a37848a,a37849a,a37850a,a37854a,a37855a,a37859a,a37860a,a37861a,a37865a,a37866a,a37870a,a37871a,a37872a,a37876a,a37877a,a37881a,a37882a,a37883a,a37887a,a37888a,a37892a,a37893a,a37894a,a37898a,a37899a,a37903a,a37904a,a37905a,a37909a,a37910a,a37914a,a37915a,a37916a,a37920a,a37921a,a37925a,a37926a,a37927a,a37931a,a37932a,a37936a,a37937a,a37938a,a37942a,a37943a,a37947a,a37948a,a37949a,a37953a,a37954a,a37958a,a37959a,a37960a,a37964a,a37965a,a37969a,a37970a,a37971a,a37975a,a37976a,a37980a,a37981a,a37982a,a37986a,a37987a,a37991a,a37992a,a37993a,a37997a,a37998a,a38002a,a38003a,a38004a,a38008a,a38009a,a38013a,a38014a,a38015a,a38019a,a38020a,a38024a,a38025a,a38026a,a38030a,a38031a,a38035a,a38036a,a38037a,a38041a,a38042a,a38046a,a38047a,a38048a,a38052a,a38053a,a38057a,a38058a,a38059a,a38063a,a38064a,a38068a,a38069a,a38070a,a38074a,a38075a,a38079a,a38080a,a38081a,a38085a,a38086a,a38090a,a38091a,a38092a,a38096a,a38097a,a38101a,a38102a,a38103a,a38107a,a38108a,a38112a,a38113a,a38114a,a38118a,a38119a,a38123a,a38124a,a38125a,a38129a,a38130a,a38134a,a38135a,a38136a,a38140a,a38141a,a38145a,a38146a,a38147a,a38151a,a38152a,a38156a,a38157a,a38158a,a38162a,a38163a,a38167a,a38168a,a38169a,a38173a,a38174a,a38178a,a38179a,a38180a,a38184a,a38185a,a38189a,a38190a,a38191a,a38195a,a38196a,a38200a,a38201a,a38202a,a38206a,a38207a,a38211a,a38212a,a38213a,a38217a,a38218a,a38222a,a38223a,a38224a,a38228a,a38229a,a38233a,a38234a,a38235a,a38239a,a38240a,a38244a,a38245a,a38246a,a38250a,a38251a,a38255a,a38256a,a38257a,a38261a,a38262a,a38266a,a38267a,a38268a,a38272a,a38273a,a38277a,a38278a,a38279a,a38283a,a38284a,a38288a,a38289a,a38290a,a38294a,a38295a,a38299a,a38300a,a38301a,a38305a,a38306a,a38310a,a38311a,a38312a,a38316a,a38317a,a38321a,a38322a,a38323a,a38327a,a38328a,a38332a,a38333a,a38334a,a38338a,a38339a,a38343a,a38344a,a38345a,a38349a,a38350a,a38354a,a38355a,a38356a,a38360a,a38361a,a38365a,a38366a,a38367a,a38371a,a38372a,a38376a,a38377a,a38378a,a38382a,a38383a,a38387a,a38388a,a38389a,a38393a,a38394a,a38398a,a38399a,a38400a,a38404a,a38405a,a38409a,a38410a,a38411a,a38415a,a38416a,a38420a,a38421a,a38422a,a38426a,a38427a,a38431a,a38432a,a38433a,a38437a,a38438a,a38442a,a38443a,a38444a,a38448a,a38449a,a38453a,a38454a,a38455a,a38459a,a38460a,a38464a,a38465a,a38466a,a38470a,a38471a,a38475a,a38476a,a38477a,a38481a,a38482a,a38486a,a38487a,a38488a,a38492a,a38493a,a38497a,a38498a,a38499a,a38503a,a38504a,a38508a,a38509a,a38510a,a38514a,a38515a,a38519a,a38520a,a38521a,a38525a,a38526a,a38530a,a38531a,a38532a,a38536a,a38537a,a38541a,a38542a,a38543a,a38547a,a38548a,a38552a,a38553a,a38554a,a38558a,a38559a,a38563a,a38564a,a38565a,a38569a,a38570a,a38574a,a38575a,a38576a,a38580a,a38581a,a38585a,a38586a,a38587a,a38591a,a38592a,a38596a,a38597a,a38598a,a38602a,a38603a,a38607a,a38608a,a38609a,a38613a,a38614a,a38618a,a38619a,a38620a,a38624a,a38625a,a38629a,a38630a,a38631a,a38635a,a38636a,a38640a,a38641a,a38642a,a38646a,a38647a,a38651a,a38652a,a38653a,a38657a,a38658a,a38662a,a38663a,a38664a,a38668a,a38669a,a38673a,a38674a,a38675a,a38679a,a38680a,a38684a,a38685a,a38686a,a38690a,a38691a,a38695a,a38696a,a38697a,a38701a,a38702a,a38706a,a38707a,a38708a,a38712a,a38713a,a38717a,a38718a,a38719a,a38723a,a38724a,a38728a,a38729a,a38730a,a38734a,a38735a,a38739a,a38740a,a38741a,a38745a,a38746a,a38750a,a38751a,a38752a,a38756a,a38757a,a38761a,a38762a,a38763a,a38767a,a38768a,a38772a,a38773a,a38774a,a38778a,a38779a,a38783a,a38784a,a38785a,a38789a,a38790a,a38794a,a38795a,a38796a,a38800a,a38801a,a38805a,a38806a,a38807a,a38811a,a38812a,a38816a,a38817a,a38818a,a38822a,a38823a,a38827a,a38828a,a38829a,a38833a,a38834a,a38838a,a38839a,a38840a,a38844a,a38845a,a38849a,a38850a,a38851a,a38855a,a38856a,a38860a,a38861a,a38862a,a38866a,a38867a,a38871a,a38872a,a38873a,a38877a,a38878a,a38882a,a38883a,a38884a,a38888a,a38889a,a38893a,a38894a,a38895a,a38899a,a38900a,a38904a,a38905a,a38906a,a38910a,a38911a,a38915a,a38916a,a38917a,a38921a,a38922a,a38926a,a38927a,a38928a,a38932a,a38933a,a38937a,a38938a,a38939a,a38943a,a38944a,a38948a,a38949a,a38950a,a38954a,a38955a,a38959a,a38960a,a38961a,a38965a,a38966a,a38970a,a38971a,a38972a,a38976a,a38977a,a38981a,a38982a,a38983a,a38987a,a38988a,a38992a,a38993a,a38994a,a38998a,a38999a,a39003a,a39004a,a39005a,a39009a,a39010a,a39014a,a39015a,a39016a,a39020a,a39021a,a39025a,a39026a,a39027a,a39031a,a39032a,a39036a,a39037a,a39038a,a39042a,a39043a,a39047a,a39048a,a39049a,a39053a,a39054a,a39058a,a39059a,a39060a,a39064a,a39065a,a39069a,a39070a,a39071a,a39075a,a39076a,a39080a,a39081a,a39082a,a39086a,a39087a,a39091a,a39092a,a39093a,a39097a,a39098a,a39102a,a39103a,a39104a,a39108a,a39109a,a39113a,a39114a,a39115a,a39119a,a39120a,a39124a,a39125a,a39126a,a39130a,a39131a,a39135a,a39136a,a39137a,a39141a,a39142a,a39146a,a39147a,a39148a,a39152a,a39153a,a39157a,a39158a,a39159a,a39163a,a39164a,a39168a,a39169a,a39170a,a39174a,a39175a,a39179a,a39180a,a39181a,a39185a,a39186a,a39190a,a39191a,a39192a,a39196a,a39197a,a39201a,a39202a,a39203a,a39207a,a39208a,a39212a,a39213a,a39214a,a39218a,a39219a,a39223a,a39224a,a39225a,a39229a,a39230a,a39234a,a39235a,a39236a,a39240a,a39241a,a39245a,a39246a,a39247a,a39251a,a39252a,a39256a,a39257a,a39258a,a39262a,a39263a,a39267a,a39268a,a39269a,a39273a,a39274a,a39278a,a39279a,a39280a,a39284a,a39285a,a39289a,a39290a,a39291a,a39295a,a39296a,a39300a,a39301a,a39302a,a39306a,a39307a,a39311a,a39312a,a39313a,a39317a,a39318a,a39322a,a39323a,a39324a,a39328a,a39329a,a39333a,a39334a,a39335a,a39339a,a39340a,a39344a,a39345a,a39346a,a39350a,a39351a,a39355a,a39356a,a39357a,a39361a,a39362a,a39366a,a39367a,a39368a,a39372a,a39373a,a39377a,a39378a,a39379a,a39383a,a39384a,a39388a,a39389a,a39390a,a39394a,a39395a,a39399a,a39400a,a39401a,a39405a,a39406a,a39410a,a39411a,a39412a,a39416a,a39417a,a39421a,a39422a,a39423a,a39427a,a39428a,a39432a,a39433a,a39434a,a39438a,a39439a,a39443a,a39444a,a39445a,a39449a,a39450a,a39454a,a39455a,a39456a,a39460a,a39461a,a39465a,a39466a,a39467a,a39471a,a39472a,a39476a,a39477a,a39478a,a39482a,a39483a,a39487a,a39488a,a39489a,a39493a,a39494a,a39498a,a39499a,a39500a,a39504a,a39505a,a39509a,a39510a,a39511a,a39515a,a39516a,a39520a,a39521a,a39522a,a39526a,a39527a,a39531a,a39532a,a39533a,a39537a,a39538a,a39542a,a39543a,a39544a,a39548a,a39549a,a39553a,a39554a,a39555a,a39559a,a39560a,a39564a,a39565a,a39566a,a39570a,a39571a,a39575a,a39576a,a39577a,a39581a,a39582a,a39586a,a39587a,a39588a,a39592a,a39593a,a39597a,a39598a,a39599a,a39603a,a39604a,a39608a,a39609a,a39610a,a39614a,a39615a,a39619a,a39620a,a39621a,a39625a,a39626a,a39630a,a39631a,a39632a,a39636a,a39637a,a39641a,a39642a,a39643a,a39647a,a39648a,a39652a,a39653a,a39654a,a39658a,a39659a,a39663a,a39664a,a39665a,a39669a,a39670a,a39674a,a39675a,a39676a,a39680a,a39681a,a39685a,a39686a,a39687a,a39691a,a39692a,a39696a,a39697a,a39698a,a39702a,a39703a,a39707a,a39708a,a39709a,a39713a,a39714a,a39718a,a39719a,a39720a,a39724a,a39725a,a39729a,a39730a,a39731a,a39735a,a39736a,a39740a,a39741a,a39742a,a39746a,a39747a,a39751a,a39752a,a39753a,a39757a,a39758a,a39762a,a39763a,a39764a,a39768a,a39769a,a39773a,a39774a,a39775a,a39779a,a39780a,a39784a,a39785a,a39786a,a39790a,a39791a,a39795a,a39796a,a39797a,a39801a,a39802a,a39806a,a39807a,a39808a,a39812a,a39813a,a39817a,a39818a,a39819a,a39823a,a39824a,a39828a,a39829a,a39830a,a39834a,a39835a,a39839a,a39840a,a39841a,a39845a,a39846a,a39850a,a39851a,a39852a,a39856a,a39857a,a39861a,a39862a,a39863a,a39867a,a39868a,a39872a,a39873a,a39874a,a39878a,a39879a,a39883a,a39884a,a39885a,a39889a,a39890a,a39894a,a39895a,a39896a,a39900a,a39901a,a39905a,a39906a,a39907a,a39911a,a39912a,a39916a,a39917a,a39918a,a39922a,a39923a,a39927a,a39928a,a39929a,a39933a,a39934a,a39938a,a39939a,a39940a,a39944a,a39945a,a39949a,a39950a,a39951a,a39955a,a39956a,a39960a,a39961a,a39962a,a39966a,a39967a,a39971a,a39972a,a39973a,a39977a,a39978a,a39982a,a39983a,a39984a,a39988a,a39989a,a39993a,a39994a,a39995a,a39999a,a40000a,a40004a,a40005a,a40006a,a40010a,a40011a,a40015a,a40016a,a40017a,a40021a,a40022a,a40026a,a40027a,a40028a,a40032a,a40033a,a40037a,a40038a,a40039a,a40043a,a40044a,a40048a,a40049a,a40050a,a40054a,a40055a,a40059a,a40060a,a40061a,a40065a,a40066a,a40070a,a40071a,a40072a,a40076a,a40077a,a40081a,a40082a,a40083a,a40087a,a40088a,a40092a,a40093a,a40094a,a40098a,a40099a,a40103a,a40104a,a40105a,a40109a,a40110a,a40114a,a40115a,a40116a,a40120a,a40121a,a40125a,a40126a,a40127a,a40131a,a40132a,a40136a,a40137a,a40138a,a40142a,a40143a,a40147a,a40148a,a40149a,a40153a,a40154a,a40158a,a40159a,a40160a,a40164a,a40165a,a40169a,a40170a,a40171a,a40175a,a40176a,a40180a,a40181a,a40182a,a40186a,a40187a,a40191a,a40192a,a40193a,a40197a,a40198a,a40202a,a40203a,a40204a,a40208a,a40209a,a40213a,a40214a,a40215a,a40219a,a40220a,a40224a,a40225a,a40226a,a40230a,a40231a,a40235a,a40236a,a40237a,a40241a,a40242a,a40246a,a40247a,a40248a,a40252a,a40253a,a40257a,a40258a,a40259a,a40263a,a40264a,a40268a,a40269a,a40270a,a40274a,a40275a,a40279a,a40280a,a40281a,a40285a,a40286a,a40290a,a40291a,a40292a,a40296a,a40297a,a40301a,a40302a,a40303a,a40307a,a40308a,a40312a,a40313a,a40314a,a40318a,a40319a,a40323a,a40324a,a40325a,a40329a,a40330a,a40334a,a40335a,a40336a,a40340a,a40341a,a40345a,a40346a,a40347a,a40351a,a40352a,a40355a,a40358a,a40359a,a40360a,a40364a,a40365a,a40369a,a40370a,a40371a,a40375a,a40376a,a40379a,a40382a,a40383a,a40384a,a40388a,a40389a,a40393a,a40394a,a40395a,a40399a,a40400a,a40403a,a40406a,a40407a,a40408a,a40412a,a40413a,a40417a,a40418a,a40419a,a40423a,a40424a,a40427a,a40430a,a40431a,a40432a,a40436a,a40437a,a40441a,a40442a,a40443a,a40447a,a40448a,a40451a,a40454a,a40455a,a40456a,a40460a,a40461a,a40465a,a40466a,a40467a,a40471a,a40472a,a40475a,a40478a,a40479a,a40480a,a40484a,a40485a,a40489a,a40490a,a40491a,a40495a,a40496a,a40499a,a40502a,a40503a,a40504a,a40508a,a40509a,a40513a,a40514a,a40515a,a40519a,a40520a,a40523a,a40526a,a40527a,a40528a,a40532a,a40533a,a40537a,a40538a,a40539a,a40543a,a40544a,a40547a,a40550a,a40551a,a40552a,a40556a,a40557a,a40561a,a40562a,a40563a,a40567a,a40568a,a40571a,a40574a,a40575a,a40576a,a40580a,a40581a,a40585a,a40586a,a40587a,a40591a,a40592a,a40595a,a40598a,a40599a,a40600a,a40604a,a40605a,a40609a,a40610a,a40611a,a40615a,a40616a,a40619a,a40622a,a40623a,a40624a,a40628a,a40629a,a40633a,a40634a,a40635a,a40639a,a40640a,a40643a,a40646a,a40647a,a40648a,a40652a,a40653a,a40657a,a40658a,a40659a,a40663a,a40664a,a40667a,a40670a,a40671a,a40672a,a40676a,a40677a,a40681a,a40682a,a40683a,a40687a,a40688a,a40691a,a40694a,a40695a,a40696a,a40700a,a40701a,a40705a,a40706a,a40707a,a40711a,a40712a,a40715a,a40718a,a40719a,a40720a,a40724a,a40725a,a40729a,a40730a,a40731a,a40735a,a40736a,a40739a,a40742a,a40743a,a40744a,a40748a,a40749a,a40753a,a40754a,a40755a,a40759a,a40760a,a40763a,a40766a,a40767a,a40768a,a40772a,a40773a,a40777a,a40778a,a40779a,a40783a,a40784a,a40787a,a40790a,a40791a,a40792a,a40796a,a40797a,a40801a,a40802a,a40803a,a40807a,a40808a,a40811a,a40814a,a40815a,a40816a,a40820a,a40821a,a40825a,a40826a,a40827a,a40831a,a40832a,a40835a,a40838a,a40839a,a40840a,a40844a,a40845a,a40849a,a40850a,a40851a,a40855a,a40856a,a40859a,a40862a,a40863a,a40864a,a40868a,a40869a,a40873a,a40874a,a40875a,a40879a,a40880a,a40883a,a40886a,a40887a,a40888a,a40892a,a40893a,a40897a,a40898a,a40899a,a40903a,a40904a,a40907a,a40910a,a40911a,a40912a,a40916a,a40917a,a40921a,a40922a,a40923a,a40927a,a40928a,a40931a,a40934a,a40935a,a40936a,a40940a,a40941a,a40945a,a40946a,a40947a,a40951a,a40952a,a40955a,a40958a,a40959a,a40960a,a40964a,a40965a,a40969a,a40970a,a40971a,a40975a,a40976a,a40979a,a40982a,a40983a,a40984a,a40988a,a40989a,a40993a,a40994a,a40995a,a40999a,a41000a,a41003a,a41006a,a41007a,a41008a,a41012a,a41013a,a41017a,a41018a,a41019a,a41023a,a41024a,a41027a,a41030a,a41031a,a41032a,a41036a,a41037a,a41041a,a41042a,a41043a,a41047a,a41048a,a41051a,a41054a,a41055a,a41056a,a41060a,a41061a,a41065a,a41066a,a41067a,a41071a,a41072a,a41075a,a41078a,a41079a,a41080a,a41084a,a41085a,a41089a,a41090a,a41091a,a41095a,a41096a,a41099a,a41102a,a41103a,a41104a,a41108a,a41109a,a41113a,a41114a,a41115a,a41119a,a41120a,a41123a,a41126a,a41127a,a41128a,a41132a,a41133a,a41137a,a41138a,a41139a,a41143a,a41144a,a41147a,a41150a,a41151a,a41152a,a41156a,a41157a,a41161a,a41162a,a41163a,a41167a,a41168a,a41171a,a41174a,a41175a,a41176a,a41180a,a41181a,a41185a,a41186a,a41187a,a41191a,a41192a,a41195a,a41198a,a41199a,a41200a,a41204a,a41205a,a41209a,a41210a,a41211a,a41215a,a41216a,a41219a,a41222a,a41223a,a41224a,a41228a,a41229a,a41233a,a41234a,a41235a,a41239a,a41240a,a41243a,a41246a,a41247a,a41248a,a41252a,a41253a,a41257a,a41258a,a41259a,a41263a,a41264a,a41267a,a41270a,a41271a,a41272a,a41276a,a41277a,a41281a,a41282a,a41283a,a41287a,a41288a,a41291a,a41294a,a41295a,a41296a,a41300a,a41301a,a41305a,a41306a,a41307a,a41311a,a41312a,a41315a,a41318a,a41319a,a41320a,a41324a,a41325a,a41329a,a41330a,a41331a,a41335a,a41336a,a41339a,a41342a,a41343a,a41344a,a41348a,a41349a,a41353a,a41354a,a41355a,a41359a,a41360a,a41363a,a41366a,a41367a,a41368a,a41372a,a41373a,a41377a,a41378a,a41379a,a41383a,a41384a,a41387a,a41390a,a41391a,a41392a,a41396a,a41397a,a41401a,a41402a,a41403a,a41407a,a41408a,a41411a,a41414a,a41415a,a41416a,a41420a,a41421a,a41425a,a41426a,a41427a,a41431a,a41432a,a41435a,a41438a,a41439a,a41440a,a41444a,a41445a,a41449a,a41450a,a41451a,a41455a,a41456a,a41459a,a41462a,a41463a,a41464a,a41468a,a41469a,a41473a,a41474a,a41475a,a41479a,a41480a,a41483a,a41486a,a41487a,a41488a,a41492a,a41493a,a41497a,a41498a,a41499a,a41503a,a41504a,a41507a,a41510a,a41511a,a41512a,a41516a,a41517a,a41521a,a41522a,a41523a,a41527a,a41528a,a41531a,a41534a,a41535a,a41536a,a41540a,a41541a,a41545a,a41546a,a41547a,a41551a,a41552a,a41555a,a41558a,a41559a,a41560a,a41564a,a41565a,a41569a,a41570a,a41571a,a41575a,a41576a,a41579a,a41582a,a41583a,a41584a,a41588a,a41589a,a41593a,a41594a,a41595a,a41599a,a41600a,a41603a,a41606a,a41607a,a41608a,a41612a,a41613a,a41617a,a41618a,a41619a,a41623a,a41624a,a41627a,a41630a,a41631a,a41632a,a41636a,a41637a,a41641a,a41642a,a41643a,a41647a,a41648a,a41651a,a41654a,a41655a,a41656a,a41660a,a41661a,a41665a,a41666a,a41667a,a41671a,a41672a,a41675a,a41678a,a41679a,a41680a,a41684a,a41685a,a41689a,a41690a,a41691a,a41695a,a41696a,a41699a,a41702a,a41703a,a41704a,a41708a,a41709a,a41713a,a41714a,a41715a,a41719a,a41720a,a41723a,a41726a,a41727a,a41728a,a41732a,a41733a,a41737a,a41738a,a41739a,a41743a,a41744a,a41747a,a41750a,a41751a,a41752a,a41756a,a41757a,a41761a,a41762a,a41763a,a41767a,a41768a,a41771a,a41774a,a41775a,a41776a,a41780a,a41781a,a41785a,a41786a,a41787a,a41791a,a41792a,a41795a,a41798a,a41799a,a41800a,a41804a,a41805a,a41809a,a41810a,a41811a,a41815a,a41816a,a41819a,a41822a,a41823a,a41824a,a41828a,a41829a,a41833a,a41834a,a41835a,a41839a,a41840a,a41843a,a41846a,a41847a,a41848a,a41852a,a41853a,a41857a,a41858a,a41859a,a41863a,a41864a,a41867a,a41870a,a41871a,a41872a,a41876a,a41877a,a41881a,a41882a,a41883a,a41887a,a41888a,a41891a,a41894a,a41895a,a41896a,a41900a,a41901a,a41905a,a41906a,a41907a,a41911a,a41912a,a41915a,a41918a,a41919a,a41920a,a41924a,a41925a,a41929a,a41930a,a41931a,a41935a,a41936a,a41939a,a41942a,a41943a,a41944a,a41948a,a41949a,a41953a,a41954a,a41955a,a41959a,a41960a,a41963a,a41966a,a41967a,a41968a,a41972a,a41973a,a41977a,a41978a,a41979a,a41983a,a41984a,a41987a,a41990a,a41991a,a41992a,a41996a,a41997a,a42001a,a42002a,a42003a,a42007a,a42008a,a42011a,a42014a,a42015a,a42016a,a42020a,a42021a,a42025a,a42026a,a42027a,a42031a,a42032a,a42035a,a42038a,a42039a,a42040a,a42044a,a42045a,a42049a,a42050a,a42051a,a42055a,a42056a,a42059a,a42062a,a42063a,a42064a,a42068a,a42069a,a42073a,a42074a,a42075a,a42079a,a42080a,a42083a,a42086a,a42087a,a42088a,a42092a,a42093a,a42097a,a42098a,a42099a,a42103a,a42104a,a42107a,a42110a,a42111a,a42112a,a42116a,a42117a,a42121a,a42122a,a42123a,a42127a,a42128a,a42131a,a42134a,a42135a,a42136a,a42140a,a42141a,a42145a,a42146a,a42147a,a42151a,a42152a,a42155a,a42158a,a42159a,a42160a,a42164a,a42165a,a42169a,a42170a,a42171a,a42175a,a42176a,a42179a,a42182a,a42183a,a42184a,a42188a,a42189a,a42193a,a42194a,a42195a,a42199a,a42200a,a42203a,a42206a,a42207a,a42208a,a42212a,a42213a,a42217a,a42218a,a42219a,a42223a,a42224a,a42227a,a42230a,a42231a,a42232a,a42236a,a42237a,a42241a,a42242a,a42243a,a42247a,a42248a,a42251a,a42254a,a42255a,a42256a,a42260a,a42261a,a42265a,a42266a,a42267a,a42271a,a42272a,a42275a,a42278a,a42279a,a42280a,a42284a,a42285a,a42289a,a42290a,a42291a,a42295a,a42296a,a42299a,a42302a,a42303a,a42304a,a42308a,a42309a,a42313a,a42314a,a42315a,a42319a,a42320a,a42323a,a42326a,a42327a,a42328a,a42332a,a42333a,a42337a,a42338a,a42339a,a42343a,a42344a,a42347a,a42350a,a42351a,a42352a,a42356a,a42357a,a42361a,a42362a,a42363a,a42367a,a42368a,a42371a,a42374a,a42375a,a42376a,a42380a,a42381a,a42385a,a42386a,a42387a,a42391a,a42392a,a42395a,a42398a,a42399a,a42400a,a42404a,a42405a,a42409a,a42410a,a42411a,a42415a,a42416a,a42419a,a42422a,a42423a,a42424a,a42428a,a42429a,a42433a,a42434a,a42435a,a42439a,a42440a,a42443a,a42446a,a42447a,a42448a,a42452a,a42453a,a42457a,a42458a,a42459a,a42463a,a42464a,a42467a,a42470a,a42471a,a42472a,a42476a,a42477a,a42481a,a42482a,a42483a,a42487a,a42488a,a42491a,a42494a,a42495a,a42496a,a42500a,a42501a,a42505a,a42506a,a42507a,a42511a,a42512a,a42515a,a42518a,a42519a,a42520a,a42524a,a42525a,a42529a,a42530a,a42531a,a42535a,a42536a,a42539a,a42542a,a42543a,a42544a,a42548a,a42549a,a42553a,a42554a,a42555a,a42559a,a42560a,a42563a,a42566a,a42567a,a42568a,a42572a,a42573a,a42577a,a42578a,a42579a,a42583a,a42584a,a42587a,a42590a,a42591a,a42592a,a42596a,a42597a,a42601a,a42602a,a42603a,a42607a,a42608a,a42611a,a42614a,a42615a,a42616a,a42620a,a42621a,a42625a,a42626a,a42627a,a42631a,a42632a,a42635a,a42638a,a42639a,a42640a,a42644a,a42645a,a42649a,a42650a,a42651a,a42655a,a42656a,a42659a,a42662a,a42663a,a42664a,a42668a,a42669a,a42673a,a42674a,a42675a,a42679a,a42680a,a42683a,a42686a,a42687a,a42688a,a42692a,a42693a,a42697a,a42698a,a42699a,a42703a,a42704a,a42707a,a42710a,a42711a,a42712a,a42716a,a42717a,a42721a,a42722a,a42723a,a42727a,a42728a,a42731a,a42734a,a42735a,a42736a,a42740a,a42741a,a42745a,a42746a,a42747a,a42751a,a42752a,a42755a,a42758a,a42759a,a42760a,a42764a,a42765a,a42769a,a42770a,a42771a,a42775a,a42776a,a42779a,a42782a,a42783a,a42784a,a42788a,a42789a,a42793a,a42794a,a42795a,a42799a,a42800a,a42803a,a42806a,a42807a,a42808a,a42812a,a42813a,a42817a,a42818a,a42819a,a42823a,a42824a,a42827a,a42830a,a42831a,a42832a,a42836a,a42837a,a42841a,a42842a,a42843a,a42847a,a42848a,a42851a,a42854a,a42855a,a42856a,a42860a,a42861a,a42865a,a42866a,a42867a,a42871a,a42872a,a42875a,a42878a,a42879a,a42880a,a42884a,a42885a,a42889a,a42890a,a42891a,a42895a,a42896a,a42899a,a42902a,a42903a,a42904a,a42908a,a42909a,a42913a,a42914a,a42915a,a42919a,a42920a,a42923a,a42926a,a42927a,a42928a,a42932a,a42933a,a42937a,a42938a,a42939a,a42943a,a42944a,a42947a,a42950a,a42951a,a42952a,a42956a,a42957a,a42961a,a42962a,a42963a,a42967a,a42968a,a42971a,a42974a,a42975a,a42976a,a42980a,a42981a,a42985a,a42986a,a42987a,a42991a,a42992a,a42995a,a42998a,a42999a,a43000a,a43004a,a43005a,a43009a,a43010a,a43011a,a43015a,a43016a,a43019a,a43022a,a43023a,a43024a,a43028a,a43029a,a43033a,a43034a,a43035a,a43039a,a43040a,a43043a,a43046a,a43047a,a43048a,a43052a,a43053a,a43057a,a43058a,a43059a,a43063a,a43064a,a43067a,a43070a,a43071a,a43072a,a43076a,a43077a,a43081a,a43082a,a43083a,a43087a,a43088a,a43091a,a43094a,a43095a,a43096a,a43100a,a43101a,a43105a,a43106a,a43107a,a43111a,a43112a,a43115a,a43118a,a43119a,a43120a,a43124a,a43125a,a43129a,a43130a,a43131a,a43135a,a43136a,a43139a,a43142a,a43143a,a43144a,a43148a,a43149a,a43153a,a43154a,a43155a,a43159a,a43160a,a43163a,a43166a,a43167a,a43168a,a43172a,a43173a,a43177a,a43178a,a43179a,a43183a,a43184a,a43187a,a43190a,a43191a,a43192a,a43196a,a43197a,a43201a,a43202a,a43203a,a43207a,a43208a,a43211a,a43214a,a43215a,a43216a,a43220a,a43221a,a43225a,a43226a,a43227a,a43231a,a43232a,a43235a,a43238a,a43239a,a43240a,a43244a,a43245a,a43249a,a43250a,a43251a,a43255a,a43256a,a43259a,a43262a,a43263a,a43264a,a43268a,a43269a,a43273a,a43274a,a43275a,a43279a,a43280a,a43283a,a43286a,a43287a,a43288a,a43292a,a43293a,a43297a,a43298a,a43299a,a43303a,a43304a,a43307a,a43310a,a43311a,a43312a,a43316a,a43317a,a43321a,a43322a,a43323a,a43327a,a43328a,a43331a,a43334a,a43335a,a43336a,a43340a,a43341a,a43345a,a43346a,a43347a,a43351a,a43352a,a43355a,a43358a,a43359a,a43360a,a43364a,a43365a,a43369a,a43370a,a43371a,a43375a,a43376a,a43379a,a43382a,a43383a,a43384a,a43388a,a43389a,a43393a,a43394a,a43395a,a43399a,a43400a,a43403a,a43406a,a43407a,a43408a,a43412a,a43413a,a43417a,a43418a,a43419a,a43423a,a43424a,a43427a,a43430a,a43431a,a43432a,a43436a,a43437a,a43441a,a43442a,a43443a,a43447a,a43448a,a43451a,a43454a,a43455a,a43456a,a43460a,a43461a,a43465a,a43466a,a43467a,a43471a,a43472a,a43475a,a43478a,a43479a,a43480a,a43484a,a43485a,a43489a,a43490a,a43491a,a43495a,a43496a,a43499a,a43502a,a43503a,a43504a,a43508a,a43509a,a43513a,a43514a,a43515a,a43519a,a43520a,a43523a,a43526a,a43527a,a43528a,a43532a,a43533a,a43537a,a43538a,a43539a,a43543a,a43544a,a43547a,a43550a,a43551a,a43552a,a43556a,a43557a,a43561a,a43562a,a43563a,a43567a,a43568a,a43571a,a43574a,a43575a,a43576a,a43580a,a43581a,a43585a,a43586a,a43587a,a43591a,a43592a,a43595a,a43598a,a43599a,a43600a,a43604a,a43605a,a43609a,a43610a,a43611a,a43615a,a43616a,a43619a,a43622a,a43623a,a43624a,a43628a,a43629a,a43633a,a43634a,a43635a,a43639a,a43640a,a43643a,a43646a,a43647a,a43648a,a43652a,a43653a,a43657a,a43658a,a43659a,a43663a,a43664a,a43667a,a43670a,a43671a,a43672a,a43676a,a43677a,a43681a,a43682a,a43683a,a43687a,a43688a,a43691a,a43694a,a43695a,a43696a,a43700a,a43701a,a43705a,a43706a,a43707a,a43711a,a43712a,a43715a,a43718a,a43719a,a43720a,a43724a,a43725a,a43729a,a43730a,a43731a,a43735a,a43736a,a43739a,a43742a,a43743a,a43744a,a43748a,a43749a,a43753a,a43754a,a43755a,a43759a,a43760a,a43763a,a43766a,a43767a,a43768a,a43772a,a43773a,a43777a,a43778a,a43779a,a43783a,a43784a,a43787a,a43790a,a43791a,a43792a,a43796a,a43797a,a43801a,a43802a,a43803a,a43807a,a43808a,a43811a,a43814a,a43815a,a43816a,a43820a,a43821a,a43825a,a43826a,a43827a,a43831a,a43832a,a43835a,a43838a,a43839a,a43840a,a43844a,a43845a,a43849a,a43850a,a43851a,a43855a,a43856a,a43859a,a43862a,a43863a,a43864a,a43868a,a43869a,a43873a,a43874a,a43875a,a43879a,a43880a,a43883a,a43886a,a43887a,a43888a,a43892a,a43893a,a43897a,a43898a,a43899a,a43903a,a43904a,a43907a,a43910a,a43911a,a43912a,a43916a,a43917a,a43921a,a43922a,a43923a,a43927a,a43928a,a43931a,a43934a,a43935a,a43936a,a43940a,a43941a,a43945a,a43946a,a43947a,a43951a,a43952a,a43955a,a43958a,a43959a,a43960a,a43964a,a43965a,a43969a,a43970a,a43971a,a43975a,a43976a,a43979a,a43982a,a43983a,a43984a,a43988a,a43989a,a43993a,a43994a,a43995a,a43999a,a44000a,a44003a,a44006a,a44007a,a44008a,a44012a,a44013a,a44017a,a44018a,a44019a,a44023a,a44024a,a44027a,a44030a,a44031a,a44032a,a44036a,a44037a,a44041a,a44042a,a44043a,a44047a,a44048a,a44051a,a44054a,a44055a,a44056a,a44060a,a44061a,a44065a,a44066a,a44067a,a44071a,a44072a,a44075a,a44078a,a44079a,a44080a,a44084a,a44085a,a44089a,a44090a,a44091a,a44095a,a44096a,a44099a,a44102a,a44103a,a44104a,a44108a,a44109a,a44113a,a44114a,a44115a,a44119a,a44120a,a44123a,a44126a,a44127a,a44128a,a44132a,a44133a,a44137a,a44138a,a44139a,a44143a,a44144a,a44147a,a44150a,a44151a,a44152a,a44156a,a44157a,a44161a,a44162a,a44163a,a44167a,a44168a,a44171a,a44174a,a44175a,a44176a,a44180a,a44181a,a44185a,a44186a,a44187a,a44191a,a44192a,a44195a,a44198a,a44199a,a44200a,a44204a,a44205a,a44209a,a44210a,a44211a,a44215a,a44216a,a44219a,a44222a,a44223a,a44224a,a44228a,a44229a,a44233a,a44234a,a44235a,a44239a,a44240a,a44243a,a44246a,a44247a,a44248a,a44252a,a44253a,a44257a,a44258a,a44259a,a44263a,a44264a,a44267a,a44270a,a44271a,a44272a,a44276a,a44277a,a44281a,a44282a,a44283a,a44287a,a44288a,a44291a,a44294a,a44295a,a44296a,a44300a,a44301a,a44305a,a44306a,a44307a,a44311a,a44312a,a44315a,a44318a,a44319a,a44320a,a44324a,a44325a,a44329a,a44330a,a44331a,a44335a,a44336a,a44339a,a44342a,a44343a,a44344a,a44348a,a44349a,a44353a,a44354a,a44355a,a44359a,a44360a,a44363a,a44366a,a44367a,a44368a,a44372a,a44373a,a44377a,a44378a,a44379a,a44383a,a44384a,a44387a,a44390a,a44391a,a44392a,a44396a,a44397a,a44401a,a44402a,a44403a,a44407a,a44408a,a44411a,a44414a,a44415a,a44416a,a44420a,a44421a,a44425a,a44426a,a44427a,a44431a,a44432a,a44435a,a44438a,a44439a,a44440a,a44444a,a44445a,a44449a,a44450a,a44451a,a44455a,a44456a,a44459a,a44462a,a44463a,a44464a,a44468a,a44469a,a44473a,a44474a,a44475a,a44479a,a44480a,a44483a,a44486a,a44487a,a44488a,a44492a,a44493a,a44497a,a44498a,a44499a,a44503a,a44504a,a44507a,a44510a,a44511a,a44512a,a44516a,a44517a,a44521a,a44522a,a44523a,a44527a,a44528a,a44531a,a44534a,a44535a,a44536a,a44540a,a44541a,a44545a,a44546a,a44547a,a44551a,a44552a,a44555a,a44558a,a44559a,a44560a,a44564a,a44565a,a44569a,a44570a,a44571a,a44575a,a44576a,a44579a,a44582a,a44583a,a44584a,a44588a,a44589a,a44593a,a44594a,a44595a,a44599a,a44600a,a44603a,a44606a,a44607a,a44608a,a44612a,a44613a,a44617a,a44618a,a44619a,a44623a,a44624a,a44627a,a44630a,a44631a,a44632a,a44636a,a44637a,a44641a,a44642a,a44643a,a44647a,a44648a,a44651a,a44654a,a44655a,a44656a,a44660a,a44661a,a44665a,a44666a,a44667a,a44671a,a44672a,a44675a,a44678a,a44679a,a44680a,a44684a,a44685a,a44689a,a44690a,a44691a,a44695a,a44696a,a44699a,a44702a,a44703a,a44704a,a44708a,a44709a,a44713a,a44714a,a44715a,a44719a,a44720a,a44723a,a44726a,a44727a,a44728a,a44732a,a44733a,a44737a,a44738a,a44739a,a44743a,a44744a,a44747a,a44750a,a44751a,a44752a,a44756a,a44757a,a44761a,a44762a,a44763a,a44767a,a44768a,a44771a,a44774a,a44775a,a44776a,a44780a,a44781a,a44785a,a44786a,a44787a,a44791a,a44792a,a44795a,a44798a,a44799a,a44800a,a44804a,a44805a,a44809a,a44810a,a44811a,a44815a,a44816a,a44819a,a44822a,a44823a,a44824a,a44828a,a44829a,a44833a,a44834a,a44835a,a44839a,a44840a,a44843a,a44846a,a44847a,a44848a,a44852a,a44853a,a44857a,a44858a,a44859a,a44863a,a44864a,a44867a,a44870a,a44871a,a44872a,a44876a,a44877a,a44881a,a44882a,a44883a,a44887a,a44888a,a44891a,a44894a,a44895a,a44896a,a44900a,a44901a,a44905a,a44906a,a44907a,a44911a,a44912a,a44915a,a44918a,a44919a,a44920a,a44924a,a44925a,a44929a,a44930a,a44931a,a44935a,a44936a,a44939a,a44942a,a44943a,a44944a,a44948a,a44949a,a44953a,a44954a,a44955a,a44959a,a44960a,a44963a,a44966a,a44967a,a44968a,a44972a,a44973a,a44977a,a44978a,a44979a,a44983a,a44984a,a44987a,a44990a,a44991a,a44992a,a44996a,a44997a,a45001a,a45002a,a45003a,a45007a,a45008a,a45011a,a45014a,a45015a,a45016a,a45020a,a45021a,a45025a,a45026a,a45027a,a45031a,a45032a,a45035a,a45038a,a45039a,a45040a,a45044a,a45045a,a45049a,a45050a,a45051a,a45055a,a45056a,a45059a,a45062a,a45063a,a45064a,a45068a,a45069a,a45073a,a45074a,a45075a,a45079a,a45080a,a45083a,a45086a,a45087a,a45088a,a45092a,a45093a,a45097a,a45098a,a45099a,a45103a,a45104a,a45107a,a45110a,a45111a,a45112a,a45116a,a45117a,a45121a,a45122a,a45123a,a45127a,a45128a,a45131a,a45134a,a45135a,a45136a,a45140a,a45141a,a45145a,a45146a,a45147a,a45151a,a45152a,a45155a,a45158a,a45159a,a45160a,a45164a,a45165a,a45169a,a45170a,a45171a,a45175a,a45176a,a45179a,a45182a,a45183a,a45184a,a45188a,a45189a,a45193a,a45194a,a45195a,a45199a,a45200a,a45203a,a45206a,a45207a,a45208a,a45212a,a45213a,a45217a,a45218a,a45219a,a45223a,a45224a,a45227a,a45230a,a45231a,a45232a,a45236a,a45237a,a45241a,a45242a,a45243a,a45247a,a45248a,a45251a,a45254a,a45255a,a45256a,a45260a,a45261a,a45265a,a45266a,a45267a,a45271a,a45272a,a45275a,a45278a,a45279a,a45280a,a45284a,a45285a,a45289a,a45290a,a45291a,a45295a,a45296a,a45299a,a45302a,a45303a,a45304a,a45308a,a45309a,a45313a,a45314a,a45315a,a45319a,a45320a,a45323a,a45326a,a45327a,a45328a,a45332a,a45333a,a45337a,a45338a,a45339a,a45343a,a45344a,a45347a,a45350a,a45351a,a45352a,a45356a,a45357a,a45361a,a45362a,a45363a,a45367a,a45368a,a45371a,a45374a,a45375a,a45376a,a45380a,a45381a,a45385a,a45386a,a45387a,a45391a,a45392a,a45395a,a45398a,a45399a,a45400a,a45404a,a45405a,a45409a,a45410a,a45411a,a45415a,a45416a,a45419a,a45422a,a45423a,a45424a,a45428a,a45429a,a45433a,a45434a,a45435a,a45439a,a45440a,a45443a,a45446a,a45447a,a45448a,a45452a,a45453a,a45457a,a45458a,a45459a,a45463a,a45464a,a45467a,a45470a,a45471a,a45472a,a45476a,a45477a,a45481a,a45482a,a45483a,a45487a,a45488a,a45491a,a45494a,a45495a,a45496a,a45500a,a45501a,a45505a,a45506a,a45507a,a45511a,a45512a,a45515a,a45518a,a45519a,a45520a,a45524a,a45525a,a45529a,a45530a,a45531a,a45535a,a45536a,a45539a,a45542a,a45543a,a45544a,a45548a,a45549a,a45553a,a45554a,a45555a,a45559a,a45560a,a45563a,a45566a,a45567a,a45568a,a45572a,a45573a,a45577a,a45578a,a45579a,a45583a,a45584a,a45587a,a45590a,a45591a,a45592a,a45596a,a45597a,a45601a,a45602a,a45603a,a45607a,a45608a,a45611a,a45614a,a45615a,a45616a,a45620a,a45621a,a45625a,a45626a,a45627a,a45631a,a45632a,a45635a,a45638a,a45639a,a45640a,a45644a,a45645a,a45649a,a45650a,a45651a,a45655a,a45656a,a45659a,a45662a,a45663a,a45664a,a45668a,a45669a,a45673a,a45674a,a45675a,a45679a,a45680a,a45683a,a45686a,a45687a,a45688a,a45692a,a45693a,a45697a,a45698a,a45699a,a45703a,a45704a,a45707a,a45710a,a45711a,a45712a,a45716a,a45717a,a45721a,a45722a,a45723a,a45727a,a45728a,a45731a,a45734a,a45735a,a45736a,a45740a,a45741a,a45745a,a45746a,a45747a,a45751a,a45752a,a45755a,a45758a,a45759a,a45760a,a45764a,a45765a,a45769a,a45770a,a45771a,a45775a,a45776a,a45779a,a45782a,a45783a,a45784a,a45788a,a45789a,a45793a,a45794a,a45795a,a45799a,a45800a,a45803a,a45806a,a45807a,a45808a,a45812a,a45813a,a45817a,a45818a,a45819a,a45823a,a45824a,a45827a,a45830a,a45831a,a45832a,a45836a,a45837a,a45841a,a45842a,a45843a,a45847a,a45848a,a45851a,a45854a,a45855a,a45856a,a45860a,a45861a,a45865a,a45866a,a45867a,a45871a,a45872a,a45875a,a45878a,a45879a,a45880a,a45884a,a45885a,a45889a,a45890a,a45891a,a45895a,a45896a,a45899a,a45902a,a45903a,a45904a,a45908a,a45909a,a45913a,a45914a,a45915a,a45919a,a45920a,a45923a,a45926a,a45927a,a45928a,a45932a,a45933a,a45937a,a45938a,a45939a,a45943a,a45944a,a45947a,a45950a,a45951a,a45952a,a45956a,a45957a,a45961a,a45962a,a45963a,a45967a,a45968a,a45971a,a45974a,a45975a,a45976a,a45980a,a45981a,a45985a,a45986a,a45987a,a45991a,a45992a,a45995a,a45998a,a45999a,a46000a,a46004a,a46005a,a46009a,a46010a,a46011a,a46015a,a46016a,a46019a,a46022a,a46023a,a46024a,a46028a,a46029a,a46033a,a46034a,a46035a,a46039a,a46040a,a46043a,a46046a,a46047a,a46048a,a46052a,a46053a,a46057a,a46058a,a46059a,a46063a,a46064a,a46067a,a46070a,a46071a,a46072a,a46076a,a46077a,a46081a,a46082a,a46083a,a46087a,a46088a,a46091a,a46094a,a46095a,a46096a,a46100a,a46101a,a46105a,a46106a,a46107a,a46111a,a46112a,a46115a,a46118a,a46119a,a46120a,a46124a,a46125a,a46129a,a46130a,a46131a,a46135a,a46136a,a46139a,a46142a,a46143a,a46144a,a46148a,a46149a,a46153a,a46154a,a46155a,a46159a,a46160a,a46163a,a46166a,a46167a,a46168a,a46172a,a46173a,a46177a,a46178a,a46179a,a46183a,a46184a,a46187a,a46190a,a46191a,a46192a,a46196a,a46197a,a46201a,a46202a,a46203a,a46207a,a46208a,a46211a,a46214a,a46215a,a46216a,a46220a,a46221a,a46225a,a46226a,a46227a,a46231a,a46232a,a46235a,a46238a,a46239a,a46240a,a46244a,a46245a,a46249a,a46250a,a46251a,a46255a,a46256a,a46259a,a46262a,a46263a,a46264a,a46268a,a46269a,a46273a,a46274a,a46275a,a46279a,a46280a,a46283a,a46286a,a46287a,a46288a,a46292a,a46293a,a46297a,a46298a,a46299a,a46303a,a46304a,a46307a,a46310a,a46311a,a46312a,a46316a,a46317a,a46321a,a46322a,a46323a,a46327a,a46328a,a46331a,a46334a,a46335a,a46336a,a46340a,a46341a,a46345a,a46346a,a46347a,a46351a,a46352a,a46355a,a46358a,a46359a,a46360a,a46364a,a46365a,a46369a,a46370a,a46371a,a46375a,a46376a,a46379a,a46382a,a46383a,a46384a,a46388a,a46389a,a46393a,a46394a,a46395a,a46399a,a46400a,a46403a,a46406a,a46407a,a46408a,a46412a,a46413a,a46417a,a46418a,a46419a,a46423a,a46424a,a46427a,a46430a,a46431a,a46432a,a46436a,a46437a,a46441a,a46442a,a46443a,a46447a,a46448a,a46451a,a46454a,a46455a,a46456a,a46460a,a46461a,a46465a,a46466a,a46467a,a46471a,a46472a,a46475a,a46478a,a46479a,a46480a,a46484a,a46485a,a46489a,a46490a,a46491a,a46495a,a46496a,a46499a,a46502a,a46503a,a46504a,a46508a,a46509a,a46513a,a46514a,a46515a,a46519a,a46520a,a46523a,a46526a,a46527a,a46528a,a46532a,a46533a,a46537a,a46538a,a46539a,a46543a,a46544a,a46547a,a46550a,a46551a,a46552a,a46556a,a46557a,a46561a,a46562a,a46563a,a46567a,a46568a,a46571a,a46574a,a46575a,a46576a,a46580a,a46581a,a46585a,a46586a,a46587a,a46591a,a46592a,a46595a,a46598a,a46599a,a46600a,a46604a,a46605a,a46609a,a46610a,a46611a,a46615a,a46616a,a46619a,a46622a,a46623a,a46624a,a46628a,a46629a,a46633a,a46634a,a46635a,a46639a,a46640a,a46643a,a46646a,a46647a,a46648a,a46652a,a46653a,a46657a,a46658a,a46659a,a46663a,a46664a,a46667a,a46670a,a46671a,a46672a,a46676a,a46677a,a46681a,a46682a,a46683a,a46687a,a46688a,a46691a,a46694a,a46695a,a46696a,a46700a,a46701a,a46705a,a46706a,a46707a,a46711a,a46712a,a46715a,a46718a,a46719a,a46720a,a46724a,a46725a,a46729a,a46730a,a46731a,a46735a,a46736a,a46739a,a46742a,a46743a,a46744a,a46748a,a46749a,a46753a,a46754a,a46755a,a46759a,a46760a,a46763a,a46766a,a46767a,a46768a,a46772a,a46773a,a46777a,a46778a,a46779a,a46783a,a46784a,a46787a,a46790a,a46791a,a46792a,a46796a,a46797a,a46801a,a46802a,a46803a,a46807a,a46808a,a46811a,a46814a,a46815a,a46816a,a46820a,a46821a,a46825a,a46826a,a46827a,a46831a,a46832a,a46835a,a46838a,a46839a,a46840a,a46844a,a46845a,a46849a,a46850a,a46851a,a46855a,a46856a,a46859a,a46862a,a46863a,a46864a,a46868a,a46869a,a46873a,a46874a,a46875a,a46879a,a46880a,a46883a,a46886a,a46887a,a46888a,a46892a,a46893a,a46897a,a46898a,a46899a,a46903a,a46904a,a46907a,a46910a,a46911a,a46912a,a46916a,a46917a,a46921a,a46922a,a46923a,a46927a,a46928a,a46931a,a46934a,a46935a,a46936a,a46940a,a46941a,a46945a,a46946a,a46947a,a46951a,a46952a,a46955a,a46958a,a46959a,a46960a,a46964a,a46965a,a46969a,a46970a,a46971a,a46975a,a46976a,a46979a,a46982a,a46983a,a46984a,a46988a,a46989a,a46993a,a46994a,a46995a,a46999a,a47000a,a47003a,a47006a,a47007a,a47008a,a47012a,a47013a,a47017a,a47018a,a47019a,a47023a,a47024a,a47027a,a47030a,a47031a,a47032a,a47036a,a47037a,a47041a,a47042a,a47043a,a47047a,a47048a,a47051a,a47054a,a47055a,a47056a,a47060a,a47061a,a47065a,a47066a,a47067a,a47071a,a47072a,a47075a,a47078a,a47079a,a47080a,a47084a,a47085a,a47089a,a47090a,a47091a,a47095a,a47096a,a47099a,a47102a,a47103a,a47104a,a47108a,a47109a,a47113a,a47114a,a47115a,a47119a,a47120a,a47123a,a47126a,a47127a,a47128a,a47132a,a47133a,a47137a,a47138a,a47139a,a47143a,a47144a,a47147a,a47150a,a47151a,a47152a,a47156a,a47157a,a47161a,a47162a,a47163a,a47167a,a47168a,a47171a,a47174a,a47175a,a47176a,a47180a,a47181a,a47185a,a47186a,a47187a,a47191a,a47192a,a47195a,a47198a,a47199a,a47200a,a47204a,a47205a,a47209a,a47210a,a47211a,a47215a,a47216a,a47219a,a47222a,a47223a,a47224a,a47228a,a47229a,a47233a,a47234a,a47235a,a47239a,a47240a,a47243a,a47246a,a47247a,a47248a,a47252a,a47253a,a47257a,a47258a,a47259a,a47263a,a47264a,a47267a,a47270a,a47271a,a47272a,a47276a,a47277a,a47281a,a47282a,a47283a,a47287a,a47288a,a47291a,a47294a,a47295a,a47296a,a47300a,a47301a,a47305a,a47306a,a47307a,a47311a,a47312a,a47315a,a47318a,a47319a,a47320a,a47324a,a47325a,a47329a,a47330a,a47331a,a47335a,a47336a,a47339a,a47342a,a47343a,a47344a,a47348a,a47349a,a47353a,a47354a,a47355a,a47359a,a47360a,a47363a,a47366a,a47367a,a47368a,a47372a,a47373a,a47377a,a47378a,a47379a,a47383a,a47384a,a47387a,a47390a,a47391a,a47392a,a47396a,a47397a,a47401a,a47402a,a47403a,a47407a,a47408a,a47411a,a47414a,a47415a,a47416a,a47420a,a47421a,a47425a,a47426a,a47427a,a47431a,a47432a,a47435a,a47438a,a47439a,a47440a,a47444a,a47445a,a47449a,a47450a,a47451a,a47455a,a47456a,a47459a,a47462a,a47463a,a47464a,a47468a,a47469a,a47473a,a47474a,a47475a,a47479a,a47480a,a47483a,a47486a,a47487a,a47488a,a47492a,a47493a,a47497a,a47498a,a47499a,a47503a,a47504a,a47507a,a47510a,a47511a,a47512a,a47516a,a47517a,a47521a,a47522a,a47523a,a47527a,a47528a,a47531a,a47534a,a47535a,a47536a,a47540a,a47541a,a47545a,a47546a,a47547a,a47551a,a47552a,a47555a,a47558a,a47559a,a47560a,a47564a,a47565a,a47569a,a47570a,a47571a,a47575a,a47576a,a47579a,a47582a,a47583a,a47584a,a47588a,a47589a,a47593a,a47594a,a47595a,a47599a,a47600a,a47603a,a47606a,a47607a,a47608a,a47612a,a47613a,a47617a,a47618a,a47619a,a47623a,a47624a,a47627a,a47630a,a47631a,a47632a,a47636a,a47637a,a47641a,a47642a,a47643a,a47647a,a47648a,a47651a,a47654a,a47655a,a47656a,a47660a,a47661a,a47665a,a47666a,a47667a,a47671a,a47672a,a47675a,a47678a,a47679a,a47680a,a47684a,a47685a,a47689a,a47690a,a47691a,a47695a,a47696a,a47699a,a47702a,a47703a,a47704a,a47708a,a47709a,a47713a,a47714a,a47715a,a47719a,a47720a,a47723a,a47726a,a47727a,a47728a,a47732a,a47733a,a47737a,a47738a,a47739a,a47743a,a47744a,a47747a,a47750a,a47751a,a47752a,a47756a,a47757a,a47761a,a47762a,a47763a,a47767a,a47768a,a47771a,a47774a,a47775a,a47776a,a47780a,a47781a,a47785a,a47786a,a47787a,a47791a,a47792a,a47795a,a47798a,a47799a,a47800a,a47804a,a47805a,a47809a,a47810a,a47811a,a47815a,a47816a,a47819a,a47822a,a47823a,a47824a,a47828a,a47829a,a47833a,a47834a,a47835a,a47839a,a47840a,a47843a,a47846a,a47847a,a47848a,a47852a,a47853a,a47857a,a47858a,a47859a,a47863a,a47864a,a47867a,a47870a,a47871a,a47872a,a47876a,a47877a,a47881a,a47882a,a47883a,a47887a,a47888a,a47891a,a47894a,a47895a,a47896a,a47900a,a47901a,a47905a,a47906a,a47907a,a47911a,a47912a,a47915a,a47918a,a47919a,a47920a,a47924a,a47925a,a47929a,a47930a,a47931a,a47935a,a47936a,a47939a,a47942a,a47943a,a47944a,a47948a,a47949a,a47953a,a47954a,a47955a,a47959a,a47960a,a47963a,a47966a,a47967a,a47968a,a47972a,a47973a,a47977a,a47978a,a47979a,a47983a,a47984a,a47987a,a47990a,a47991a,a47992a,a47996a,a47997a,a48001a,a48002a,a48003a,a48007a,a48008a,a48011a,a48014a,a48015a,a48016a,a48020a,a48021a,a48025a,a48026a,a48027a,a48031a,a48032a,a48035a,a48038a,a48039a,a48040a,a48044a,a48045a,a48049a,a48050a,a48051a,a48055a,a48056a,a48059a,a48062a,a48063a,a48064a,a48068a,a48069a,a48073a,a48074a,a48075a,a48079a,a48080a,a48083a,a48086a,a48087a,a48088a,a48092a,a48093a,a48097a,a48098a,a48099a,a48103a,a48104a,a48107a,a48110a,a48111a,a48112a,a48116a,a48117a,a48121a,a48122a,a48123a,a48127a,a48128a,a48131a,a48134a,a48135a,a48136a,a48140a,a48141a,a48145a,a48146a,a48147a,a48151a,a48152a,a48155a,a48158a,a48159a,a48160a,a48164a,a48165a,a48169a,a48170a,a48171a,a48175a,a48176a,a48179a,a48182a,a48183a,a48184a,a48188a,a48189a,a48193a,a48194a,a48195a,a48199a,a48200a,a48203a,a48206a,a48207a,a48208a,a48212a,a48213a,a48217a,a48218a,a48219a,a48223a,a48224a,a48227a,a48230a,a48231a,a48232a,a48236a,a48237a,a48241a,a48242a,a48243a,a48247a,a48248a,a48251a,a48254a,a48255a,a48256a,a48260a,a48261a,a48265a,a48266a,a48267a,a48271a,a48272a,a48275a,a48278a,a48279a,a48280a,a48284a,a48285a,a48289a,a48290a,a48291a,a48295a,a48296a,a48299a,a48302a,a48303a,a48304a,a48308a,a48309a,a48313a,a48314a,a48315a,a48319a,a48320a,a48323a,a48326a,a48327a,a48328a,a48332a,a48333a,a48337a,a48338a,a48339a,a48343a,a48344a,a48347a,a48350a,a48351a,a48352a,a48356a,a48357a,a48361a,a48362a,a48363a,a48367a,a48368a,a48371a,a48374a,a48375a,a48376a,a48380a,a48381a,a48385a,a48386a,a48387a,a48391a,a48392a,a48395a,a48398a,a48399a,a48400a,a48404a,a48405a,a48409a,a48410a,a48411a,a48415a,a48416a,a48419a,a48422a,a48423a,a48424a,a48428a,a48429a,a48433a,a48434a,a48435a,a48439a,a48440a,a48443a,a48446a,a48447a,a48448a,a48452a,a48453a,a48457a,a48458a,a48459a,a48463a,a48464a,a48467a,a48470a,a48471a,a48472a,a48476a,a48477a,a48481a,a48482a,a48483a,a48487a,a48488a,a48491a,a48494a,a48495a,a48496a,a48500a,a48501a,a48505a,a48506a,a48507a,a48511a,a48512a,a48515a,a48518a,a48519a,a48520a,a48524a,a48525a,a48529a,a48530a,a48531a,a48535a,a48536a,a48539a,a48542a,a48543a,a48544a,a48548a,a48549a,a48553a,a48554a,a48555a,a48559a,a48560a,a48563a,a48566a,a48567a,a48568a,a48572a,a48573a,a48577a,a48578a,a48579a,a48583a,a48584a,a48587a,a48590a,a48591a,a48592a,a48596a,a48597a,a48601a,a48602a,a48603a,a48607a,a48608a,a48611a,a48614a,a48615a,a48616a,a48620a,a48621a,a48625a,a48626a,a48627a,a48631a,a48632a,a48635a,a48638a,a48639a,a48640a,a48644a,a48645a,a48649a,a48650a,a48651a,a48655a,a48656a,a48659a,a48662a,a48663a,a48664a,a48668a,a48669a,a48673a,a48674a,a48675a,a48679a,a48680a,a48683a,a48686a,a48687a,a48688a,a48692a,a48693a,a48697a,a48698a,a48699a,a48703a,a48704a,a48707a,a48710a,a48711a,a48712a,a48716a,a48717a,a48721a,a48722a,a48723a,a48727a,a48728a,a48731a,a48734a,a48735a,a48736a,a48740a,a48741a,a48745a,a48746a,a48747a,a48751a,a48752a,a48755a,a48758a,a48759a,a48760a,a48764a,a48765a,a48769a,a48770a,a48771a,a48775a,a48776a,a48779a,a48782a,a48783a,a48784a,a48788a,a48789a,a48793a,a48794a,a48795a,a48799a,a48800a,a48803a,a48806a,a48807a,a48808a,a48812a,a48813a,a48817a,a48818a,a48819a,a48823a,a48824a,a48827a,a48830a,a48831a,a48832a,a48836a,a48837a,a48841a,a48842a,a48843a,a48847a,a48848a,a48851a,a48854a,a48855a,a48856a,a48860a,a48861a,a48865a,a48866a,a48867a,a48871a,a48872a,a48875a,a48878a,a48879a,a48880a,a48884a,a48885a,a48889a,a48890a,a48891a,a48895a,a48896a,a48899a,a48902a,a48903a,a48904a,a48908a,a48909a,a48913a,a48914a,a48915a,a48919a,a48920a,a48923a,a48926a,a48927a,a48928a,a48932a,a48933a,a48937a,a48938a,a48939a,a48943a,a48944a,a48947a,a48950a,a48951a,a48952a,a48956a,a48957a,a48961a,a48962a,a48963a,a48967a,a48968a,a48971a,a48974a,a48975a,a48976a,a48980a,a48981a,a48985a,a48986a,a48987a,a48991a,a48992a,a48995a,a48998a,a48999a,a49000a,a49004a,a49005a,a49009a,a49010a,a49011a,a49015a,a49016a,a49019a,a49022a,a49023a,a49024a,a49028a,a49029a,a49033a,a49034a,a49035a,a49039a,a49040a,a49043a,a49046a,a49047a,a49048a,a49052a,a49053a,a49057a,a49058a,a49059a,a49063a,a49064a,a49067a,a49070a,a49071a,a49072a,a49076a,a49077a,a49081a,a49082a,a49083a,a49087a,a49088a,a49091a,a49094a,a49095a,a49096a,a49100a,a49101a,a49105a,a49106a,a49107a,a49111a,a49112a,a49115a,a49118a,a49119a,a49120a,a49124a,a49125a,a49129a,a49130a,a49131a,a49135a,a49136a,a49139a,a49142a,a49143a,a49144a,a49148a,a49149a,a49153a,a49154a,a49155a,a49159a,a49160a,a49163a,a49166a,a49167a,a49168a,a49172a,a49173a,a49177a,a49178a,a49179a,a49183a,a49184a,a49187a,a49190a,a49191a,a49192a,a49196a,a49197a,a49201a,a49202a,a49203a,a49207a,a49208a,a49211a,a49214a,a49215a,a49216a,a49220a,a49221a,a49225a,a49226a,a49227a,a49231a,a49232a,a49235a,a49238a,a49239a,a49240a,a49244a,a49245a,a49249a,a49250a,a49251a,a49255a,a49256a,a49259a,a49262a,a49263a,a49264a,a49268a,a49269a,a49273a,a49274a,a49275a,a49279a,a49280a,a49283a,a49286a,a49287a,a49288a,a49292a,a49293a,a49297a,a49298a,a49299a,a49303a,a49304a,a49307a,a49310a,a49311a,a49312a,a49316a,a49317a,a49321a,a49322a,a49323a,a49327a,a49328a,a49331a,a49334a,a49335a,a49336a,a49340a,a49341a,a49345a,a49346a,a49347a,a49351a,a49352a,a49355a,a49358a,a49359a,a49360a,a49364a,a49365a,a49369a,a49370a,a49371a,a49375a,a49376a,a49379a,a49382a,a49383a,a49384a,a49388a,a49389a,a49393a,a49394a,a49395a,a49399a,a49400a,a49403a,a49406a,a49407a,a49408a,a49412a,a49413a,a49417a,a49418a,a49419a,a49423a,a49424a,a49427a,a49430a,a49431a,a49432a,a49436a,a49437a,a49441a,a49442a,a49443a,a49447a,a49448a,a49451a,a49454a,a49455a,a49456a,a49460a,a49461a,a49465a,a49466a,a49467a,a49471a,a49472a,a49475a,a49478a,a49479a,a49480a,a49484a,a49485a,a49489a,a49490a,a49491a,a49495a,a49496a,a49499a,a49502a,a49503a,a49504a,a49508a,a49509a,a49513a,a49514a,a49515a,a49519a,a49520a,a49523a,a49526a,a49527a,a49528a,a49532a,a49533a,a49537a,a49538a,a49539a,a49543a,a49544a,a49547a,a49550a,a49551a,a49552a,a49556a,a49557a,a49561a,a49562a,a49563a,a49567a,a49568a,a49571a,a49574a,a49575a,a49576a,a49580a,a49581a,a49585a,a49586a,a49587a,a49591a,a49592a,a49595a,a49598a,a49599a,a49600a,a49604a,a49605a,a49609a,a49610a,a49611a,a49615a,a49616a,a49619a,a49622a,a49623a,a49624a,a49628a,a49629a,a49633a,a49634a,a49635a,a49639a,a49640a,a49643a,a49646a,a49647a,a49648a,a49652a,a49653a,a49657a,a49658a,a49659a,a49663a,a49664a,a49667a,a49670a,a49671a,a49672a,a49676a,a49677a,a49681a,a49682a,a49683a,a49687a,a49688a,a49691a,a49694a,a49695a,a49696a,a49700a,a49701a,a49705a,a49706a,a49707a,a49711a,a49712a,a49715a,a49718a,a49719a,a49720a,a49724a,a49725a,a49729a,a49730a,a49731a,a49735a,a49736a,a49739a,a49742a,a49743a,a49744a,a49748a,a49749a,a49753a,a49754a,a49755a,a49759a,a49760a,a49763a,a49766a,a49767a,a49768a,a49772a,a49773a,a49777a,a49778a,a49779a,a49783a,a49784a,a49787a,a49790a,a49791a,a49792a,a49796a,a49797a,a49801a,a49802a,a49803a,a49807a,a49808a,a49811a,a49814a,a49815a,a49816a,a49820a,a49821a,a49825a,a49826a,a49827a,a49831a,a49832a,a49835a,a49838a,a49839a,a49840a,a49844a,a49845a,a49849a,a49850a,a49851a,a49855a,a49856a,a49859a,a49862a,a49863a,a49864a,a49868a,a49869a,a49873a,a49874a,a49875a,a49879a,a49880a,a49883a,a49886a,a49887a,a49888a,a49892a,a49893a,a49897a,a49898a,a49899a,a49903a,a49904a,a49907a,a49910a,a49911a,a49912a,a49916a,a49917a,a49921a,a49922a,a49923a,a49927a,a49928a,a49931a,a49934a,a49935a,a49936a,a49940a,a49941a,a49945a,a49946a,a49947a,a49951a,a49952a,a49955a,a49958a,a49959a,a49960a,a49964a,a49965a,a49969a,a49970a,a49971a,a49975a,a49976a,a49979a,a49982a,a49983a,a49984a,a49988a,a49989a,a49993a,a49994a,a49995a,a49999a,a50000a,a50003a,a50006a,a50007a,a50008a,a50012a,a50013a,a50017a,a50018a,a50019a,a50023a,a50024a,a50027a,a50030a,a50031a,a50032a,a50036a,a50037a,a50041a,a50042a,a50043a,a50047a,a50048a,a50051a,a50054a,a50055a,a50056a,a50060a,a50061a,a50065a,a50066a,a50067a,a50071a,a50072a,a50075a,a50078a,a50079a,a50080a,a50084a,a50085a,a50089a,a50090a,a50091a,a50095a,a50096a,a50099a,a50102a,a50103a,a50104a,a50108a,a50109a,a50113a,a50114a,a50115a,a50119a,a50120a,a50123a,a50126a,a50127a,a50128a,a50132a,a50133a,a50137a,a50138a,a50139a,a50143a,a50144a,a50147a,a50150a,a50151a,a50152a,a50156a,a50157a,a50161a,a50162a,a50163a,a50167a,a50168a,a50171a,a50174a,a50175a,a50176a,a50180a,a50181a,a50185a,a50186a,a50187a,a50191a,a50192a,a50195a,a50198a,a50199a,a50200a,a50204a,a50205a,a50209a,a50210a,a50211a,a50215a,a50216a,a50219a,a50222a,a50223a,a50224a,a50228a,a50229a,a50233a,a50234a,a50235a,a50239a,a50240a,a50243a,a50246a,a50247a,a50248a,a50252a,a50253a,a50257a,a50258a,a50259a,a50263a,a50264a,a50267a,a50270a,a50271a,a50272a,a50276a,a50277a,a50281a,a50282a,a50283a,a50287a,a50288a,a50291a,a50294a,a50295a,a50296a,a50300a,a50301a,a50305a,a50306a,a50307a,a50311a,a50312a,a50315a,a50318a,a50319a,a50320a,a50324a,a50325a,a50329a,a50330a,a50331a,a50335a,a50336a,a50339a,a50342a,a50343a,a50344a,a50348a,a50349a,a50353a,a50354a,a50355a,a50359a,a50360a,a50363a,a50366a,a50367a,a50368a,a50372a,a50373a,a50377a,a50378a,a50379a,a50383a,a50384a,a50387a,a50390a,a50391a,a50392a,a50396a,a50397a,a50401a,a50402a,a50403a,a50407a,a50408a,a50411a,a50414a,a50415a,a50416a,a50420a,a50421a,a50425a,a50426a,a50427a,a50431a,a50432a,a50435a,a50438a,a50439a,a50440a,a50444a,a50445a,a50449a,a50450a,a50451a,a50455a,a50456a,a50459a,a50462a,a50463a,a50464a,a50468a,a50469a,a50473a,a50474a,a50475a,a50479a,a50480a,a50483a,a50486a,a50487a,a50488a,a50492a,a50493a,a50497a,a50498a,a50499a,a50503a,a50504a,a50507a,a50510a,a50511a,a50512a,a50516a,a50517a,a50521a,a50522a,a50523a,a50527a,a50528a,a50531a,a50534a,a50535a,a50536a,a50540a,a50541a,a50545a,a50546a,a50547a,a50551a,a50552a,a50555a,a50558a,a50559a,a50560a,a50564a,a50565a,a50569a,a50570a,a50571a,a50575a,a50576a,a50579a,a50582a,a50583a,a50584a,a50588a,a50589a,a50593a,a50594a,a50595a,a50599a,a50600a,a50603a,a50606a,a50607a,a50608a,a50612a,a50613a,a50617a,a50618a,a50619a,a50623a,a50624a,a50627a,a50630a,a50631a,a50632a,a50636a,a50637a,a50641a,a50642a,a50643a,a50647a,a50648a,a50651a,a50654a,a50655a,a50656a,a50660a,a50661a,a50665a,a50666a,a50667a,a50671a,a50672a,a50675a,a50678a,a50679a,a50680a,a50684a,a50685a,a50689a,a50690a,a50691a,a50695a,a50696a,a50699a,a50702a,a50703a,a50704a,a50708a,a50709a,a50713a,a50714a,a50715a,a50719a,a50720a,a50723a,a50726a,a50727a,a50728a,a50732a,a50733a,a50737a,a50738a,a50739a,a50743a,a50744a,a50747a,a50750a,a50751a,a50752a,a50756a,a50757a,a50761a,a50762a,a50763a,a50767a,a50768a,a50771a,a50774a,a50775a,a50776a,a50780a,a50781a,a50785a,a50786a,a50787a,a50791a,a50792a,a50795a,a50798a,a50799a,a50800a,a50804a,a50805a,a50809a,a50810a,a50811a,a50815a,a50816a,a50819a,a50822a,a50823a,a50824a,a50828a,a50829a,a50833a,a50834a,a50835a,a50839a,a50840a,a50843a,a50846a,a50847a,a50848a,a50852a,a50853a,a50857a,a50858a,a50859a,a50863a,a50864a,a50867a,a50870a,a50871a,a50872a,a50876a,a50877a,a50881a,a50882a,a50883a,a50887a,a50888a,a50891a,a50894a,a50895a,a50896a,a50900a,a50901a,a50905a,a50906a,a50907a,a50911a,a50912a,a50915a,a50918a,a50919a,a50920a,a50924a,a50925a,a50929a,a50930a,a50931a,a50935a,a50936a,a50939a,a50942a,a50943a,a50944a,a50948a,a50949a,a50953a,a50954a,a50955a,a50959a,a50960a,a50963a,a50966a,a50967a,a50968a,a50972a,a50973a,a50977a,a50978a,a50979a,a50983a,a50984a,a50987a,a50990a,a50991a,a50992a,a50996a,a50997a,a51001a,a51002a,a51003a,a51007a,a51008a,a51011a,a51014a,a51015a,a51016a,a51020a,a51021a,a51025a,a51026a,a51027a,a51031a,a51032a,a51035a,a51038a,a51039a,a51040a,a51044a,a51045a,a51049a,a51050a,a51051a,a51055a,a51056a,a51059a,a51062a,a51063a,a51064a,a51068a,a51069a,a51073a,a51074a,a51075a,a51079a,a51080a,a51083a,a51086a,a51087a,a51088a,a51092a,a51093a,a51097a,a51098a,a51099a,a51103a,a51104a,a51107a,a51110a,a51111a,a51112a,a51116a,a51117a,a51121a,a51122a,a51123a,a51127a,a51128a,a51131a,a51134a,a51135a,a51136a,a51140a,a51141a,a51145a,a51146a,a51147a,a51151a,a51152a,a51155a,a51158a,a51159a,a51160a,a51164a,a51165a,a51169a,a51170a,a51171a,a51175a,a51176a,a51179a,a51182a,a51183a,a51184a,a51188a,a51189a,a51193a,a51194a,a51195a,a51199a,a51200a,a51203a,a51206a,a51207a,a51208a,a51212a,a51213a,a51217a,a51218a,a51219a,a51223a,a51224a,a51227a,a51230a,a51231a,a51232a,a51236a,a51237a,a51241a,a51242a,a51243a,a51247a,a51248a,a51251a,a51254a,a51255a,a51256a,a51260a,a51261a,a51265a,a51266a,a51267a,a51271a,a51272a,a51275a,a51278a,a51279a,a51280a,a51284a,a51285a,a51289a,a51290a,a51291a,a51295a,a51296a,a51299a,a51302a,a51303a,a51304a,a51308a,a51309a,a51313a,a51314a,a51315a,a51319a,a51320a,a51323a,a51326a,a51327a,a51328a,a51332a,a51333a,a51337a,a51338a,a51339a,a51343a,a51344a,a51347a,a51350a,a51351a,a51352a,a51356a,a51357a,a51361a,a51362a,a51363a,a51367a,a51368a,a51371a,a51374a,a51375a,a51376a,a51380a,a51381a,a51385a,a51386a,a51387a,a51391a,a51392a,a51395a,a51398a,a51399a,a51400a,a51404a,a51405a,a51409a,a51410a,a51411a,a51415a,a51416a,a51419a,a51422a,a51423a,a51424a,a51428a,a51429a,a51433a,a51434a,a51435a,a51439a,a51440a,a51443a,a51446a,a51447a,a51448a,a51452a,a51453a,a51457a,a51458a,a51459a,a51463a,a51464a,a51467a,a51470a,a51471a,a51472a,a51476a,a51477a,a51481a,a51482a,a51483a,a51487a,a51488a,a51491a,a51494a,a51495a,a51496a,a51500a,a51501a,a51505a,a51506a,a51507a,a51511a,a51512a,a51515a,a51518a,a51519a,a51520a,a51524a,a51525a,a51529a,a51530a,a51531a,a51535a,a51536a,a51539a,a51542a,a51543a,a51544a,a51548a,a51549a,a51553a,a51554a,a51555a,a51559a,a51560a,a51563a,a51566a,a51567a,a51568a,a51572a,a51573a,a51577a,a51578a,a51579a,a51583a,a51584a,a51587a,a51590a,a51591a,a51592a,a51596a,a51597a,a51601a,a51602a,a51603a,a51607a,a51608a,a51611a,a51614a,a51615a,a51616a,a51620a,a51621a,a51625a,a51626a,a51627a,a51631a,a51632a,a51635a,a51638a,a51639a,a51640a,a51644a,a51645a,a51649a,a51650a,a51651a,a51655a,a51656a,a51659a,a51662a,a51663a,a51664a,a51668a,a51669a,a51673a,a51674a,a51675a,a51679a,a51680a,a51683a,a51686a,a51687a,a51688a,a51692a,a51693a,a51697a,a51698a,a51699a,a51703a,a51704a,a51707a,a51710a,a51711a,a51712a,a51716a,a51717a,a51721a,a51722a,a51723a,a51727a,a51728a,a51731a,a51734a,a51735a,a51736a,a51740a,a51741a,a51745a,a51746a,a51747a,a51751a,a51752a,a51755a,a51758a,a51759a,a51760a,a51764a,a51765a,a51769a,a51770a,a51771a,a51775a,a51776a,a51779a,a51782a,a51783a,a51784a,a51788a,a51789a,a51793a,a51794a,a51795a,a51799a,a51800a,a51803a,a51806a,a51807a,a51808a,a51812a,a51813a,a51817a,a51818a,a51819a,a51823a,a51824a,a51827a,a51830a,a51831a,a51832a,a51836a,a51837a,a51841a,a51842a,a51843a,a51847a,a51848a,a51851a,a51854a,a51855a,a51856a,a51860a,a51861a,a51865a,a51866a,a51867a,a51871a,a51872a,a51875a,a51878a,a51879a,a51880a,a51884a,a51885a,a51889a,a51890a,a51891a,a51895a,a51896a,a51899a,a51902a,a51903a,a51904a,a51908a,a51909a,a51913a,a51914a,a51915a,a51919a,a51920a,a51923a,a51926a,a51927a,a51928a,a51932a,a51933a,a51937a,a51938a,a51939a,a51943a,a51944a,a51947a,a51950a,a51951a,a51952a,a51956a,a51957a,a51961a,a51962a,a51963a,a51967a,a51968a,a51971a,a51974a,a51975a,a51976a,a51980a,a51981a,a51985a,a51986a,a51987a,a51991a,a51992a,a51995a,a51998a,a51999a,a52000a,a52004a,a52005a,a52009a,a52010a,a52011a,a52015a,a52016a,a52019a,a52022a,a52023a,a52024a,a52028a,a52029a,a52033a,a52034a,a52035a,a52039a,a52040a,a52043a,a52046a,a52047a,a52048a,a52052a,a52053a,a52057a,a52058a,a52059a,a52063a,a52064a,a52067a,a52070a,a52071a,a52072a,a52076a,a52077a,a52081a,a52082a,a52083a,a52087a,a52088a,a52091a,a52094a,a52095a,a52096a,a52100a,a52101a,a52105a,a52106a,a52107a,a52111a,a52112a,a52115a,a52118a,a52119a,a52120a,a52124a,a52125a,a52129a,a52130a,a52131a,a52135a,a52136a,a52139a,a52142a,a52143a,a52144a,a52148a,a52149a,a52153a,a52154a,a52155a,a52159a,a52160a,a52163a,a52166a,a52167a,a52168a,a52172a,a52173a,a52177a,a52178a,a52179a,a52183a,a52184a,a52187a,a52190a,a52191a,a52192a,a52196a,a52197a,a52201a,a52202a,a52203a,a52207a,a52208a,a52211a,a52214a,a52215a,a52216a,a52220a,a52221a,a52225a,a52226a,a52227a,a52231a,a52232a,a52235a,a52238a,a52239a,a52240a,a52244a,a52245a,a52249a,a52250a,a52251a,a52255a,a52256a,a52259a,a52262a,a52263a,a52264a,a52268a,a52269a,a52273a,a52274a,a52275a,a52279a,a52280a,a52283a,a52286a,a52287a,a52288a,a52292a,a52293a,a52297a,a52298a,a52299a,a52303a,a52304a,a52307a,a52310a,a52311a,a52312a,a52316a,a52317a,a52321a,a52322a,a52323a,a52327a,a52328a,a52331a,a52334a,a52335a,a52336a,a52340a,a52341a,a52345a,a52346a,a52347a,a52351a,a52352a,a52355a,a52358a,a52359a,a52360a,a52364a,a52365a,a52369a,a52370a,a52371a,a52375a,a52376a,a52379a,a52382a,a52383a,a52384a,a52388a,a52389a,a52393a,a52394a,a52395a,a52399a,a52400a,a52403a,a52406a,a52407a,a52408a,a52412a,a52413a,a52417a,a52418a,a52419a,a52423a,a52424a,a52427a,a52430a,a52431a,a52432a,a52436a,a52437a,a52441a,a52442a,a52443a,a52447a,a52448a,a52451a,a52454a,a52455a,a52456a,a52460a,a52461a,a52465a,a52466a,a52467a,a52471a,a52472a,a52475a,a52478a,a52479a,a52480a,a52484a,a52485a,a52489a,a52490a,a52491a,a52495a,a52496a,a52499a,a52502a,a52503a,a52504a,a52508a,a52509a,a52513a,a52514a,a52515a,a52519a,a52520a,a52523a,a52526a,a52527a,a52528a,a52532a,a52533a,a52537a,a52538a,a52539a,a52543a,a52544a,a52547a,a52550a,a52551a,a52552a,a52556a,a52557a,a52561a,a52562a,a52563a,a52567a,a52568a,a52571a,a52574a,a52575a,a52576a,a52580a,a52581a,a52585a,a52586a,a52587a,a52591a,a52592a,a52595a,a52598a,a52599a,a52600a,a52604a,a52605a,a52609a,a52610a,a52611a,a52615a,a52616a,a52619a,a52622a,a52623a,a52624a,a52628a,a52629a,a52633a,a52634a,a52635a,a52639a,a52640a,a52643a,a52646a,a52647a,a52648a,a52652a,a52653a,a52657a,a52658a,a52659a,a52663a,a52664a,a52667a,a52670a,a52671a,a52672a,a52676a,a52677a,a52681a,a52682a,a52683a,a52687a,a52688a,a52691a,a52694a,a52695a,a52696a,a52700a,a52701a,a52705a,a52706a,a52707a,a52711a,a52712a,a52715a,a52718a,a52719a,a52720a,a52724a,a52725a,a52729a,a52730a,a52731a,a52735a,a52736a,a52739a,a52742a,a52743a,a52744a,a52748a,a52749a,a52753a,a52754a,a52755a,a52759a,a52760a,a52763a,a52766a,a52767a,a52768a,a52772a,a52773a,a52777a,a52778a,a52779a,a52783a,a52784a,a52787a,a52790a,a52791a,a52792a,a52796a,a52797a,a52801a,a52802a,a52803a,a52807a,a52808a,a52811a,a52814a,a52815a,a52816a,a52820a,a52821a,a52825a,a52826a,a52827a,a52831a,a52832a,a52835a,a52838a,a52839a,a52840a,a52844a,a52845a,a52849a,a52850a,a52851a,a52855a,a52856a,a52859a,a52862a,a52863a,a52864a,a52868a,a52869a,a52873a,a52874a,a52875a,a52879a,a52880a,a52883a,a52886a,a52887a,a52888a,a52892a,a52893a,a52897a,a52898a,a52899a,a52903a,a52904a,a52907a,a52910a,a52911a,a52912a,a52916a,a52917a,a52921a,a52922a,a52923a,a52927a,a52928a,a52931a,a52934a,a52935a,a52936a,a52940a,a52941a,a52945a,a52946a,a52947a,a52951a,a52952a,a52955a,a52958a,a52959a,a52960a,a52964a,a52965a,a52969a,a52970a,a52971a,a52975a,a52976a,a52979a,a52982a,a52983a,a52984a,a52988a,a52989a,a52993a,a52994a,a52995a,a52999a,a53000a,a53003a,a53006a,a53007a,a53008a,a53012a,a53013a,a53017a,a53018a,a53019a,a53023a,a53024a,a53027a,a53030a,a53031a,a53032a,a53036a,a53037a,a53041a,a53042a,a53043a,a53047a,a53048a,a53051a,a53054a,a53055a,a53056a,a53060a,a53061a,a53065a,a53066a,a53067a,a53071a,a53072a,a53075a,a53078a,a53079a,a53080a,a53084a,a53085a,a53089a,a53090a,a53091a,a53095a,a53096a,a53099a,a53102a,a53103a,a53104a,a53108a,a53109a,a53113a,a53114a,a53115a,a53119a,a53120a,a53123a,a53126a,a53127a,a53128a,a53132a,a53133a,a53137a,a53138a,a53139a,a53143a,a53144a,a53147a,a53150a,a53151a,a53152a,a53156a,a53157a,a53161a,a53162a,a53163a,a53167a,a53168a,a53171a,a53174a,a53175a,a53176a,a53180a,a53181a,a53185a,a53186a,a53187a,a53191a,a53192a,a53195a,a53198a,a53199a,a53200a,a53204a,a53205a,a53209a,a53210a,a53211a,a53215a,a53216a,a53219a,a53222a,a53223a,a53224a,a53228a,a53229a,a53233a,a53234a,a53235a,a53239a,a53240a,a53243a,a53246a,a53247a,a53248a,a53252a,a53253a,a53257a,a53258a,a53259a,a53263a,a53264a,a53267a,a53270a,a53271a,a53272a,a53276a,a53277a,a53281a,a53282a,a53283a,a53287a,a53288a,a53291a,a53294a,a53295a,a53296a,a53300a,a53301a,a53305a,a53306a,a53307a,a53311a,a53312a,a53315a,a53318a,a53319a,a53320a,a53324a,a53325a,a53329a,a53330a,a53331a,a53335a,a53336a,a53339a,a53342a,a53343a,a53344a,a53348a,a53349a,a53353a,a53354a,a53355a,a53359a,a53360a,a53363a,a53366a,a53367a,a53368a,a53372a,a53373a,a53377a,a53378a,a53379a,a53383a,a53384a,a53387a,a53390a,a53391a,a53392a,a53396a,a53397a,a53401a,a53402a,a53403a,a53407a,a53408a,a53411a,a53414a,a53415a,a53416a,a53420a,a53421a,a53425a,a53426a,a53427a,a53431a,a53432a,a53435a,a53438a,a53439a,a53440a,a53444a,a53445a,a53449a,a53450a,a53451a,a53455a,a53456a,a53459a,a53462a,a53463a,a53464a,a53468a,a53469a,a53473a,a53474a,a53475a,a53479a,a53480a,a53483a,a53486a,a53487a,a53488a,a53492a,a53493a,a53497a,a53498a,a53499a,a53503a,a53504a,a53507a,a53510a,a53511a,a53512a,a53516a,a53517a,a53521a,a53522a,a53523a,a53527a,a53528a,a53531a,a53534a,a53535a,a53536a,a53540a,a53541a,a53545a,a53546a,a53547a,a53551a,a53552a,a53555a,a53558a,a53559a,a53560a,a53564a,a53565a,a53569a,a53570a,a53571a,a53575a,a53576a,a53579a,a53582a,a53583a,a53584a,a53588a,a53589a,a53593a,a53594a,a53595a,a53599a,a53600a,a53603a,a53606a,a53607a,a53608a,a53612a,a53613a,a53617a,a53618a,a53619a,a53623a,a53624a,a53627a,a53630a,a53631a,a53632a,a53636a,a53637a,a53641a,a53642a,a53643a,a53647a,a53648a,a53651a,a53654a,a53655a,a53656a,a53660a,a53661a,a53665a,a53666a,a53667a,a53671a,a53672a,a53675a,a53678a,a53679a,a53680a,a53684a,a53685a,a53689a,a53690a,a53691a,a53695a,a53696a,a53699a,a53702a,a53703a,a53704a,a53708a,a53709a,a53713a,a53714a,a53715a,a53719a,a53720a,a53723a,a53726a,a53727a,a53728a,a53732a,a53733a,a53737a,a53738a,a53739a,a53743a,a53744a,a53747a,a53750a,a53751a,a53752a,a53756a,a53757a,a53761a,a53762a,a53763a,a53767a,a53768a,a53771a,a53774a,a53775a,a53776a,a53780a,a53781a,a53785a,a53786a,a53787a,a53791a,a53792a,a53795a,a53798a,a53799a,a53800a,a53804a,a53805a,a53809a,a53810a,a53811a,a53815a,a53816a,a53819a,a53822a,a53823a,a53824a,a53828a,a53829a,a53833a,a53834a,a53835a,a53839a,a53840a,a53843a,a53846a,a53847a,a53848a,a53852a,a53853a,a53857a,a53858a,a53859a,a53863a,a53864a,a53867a,a53870a,a53871a,a53872a,a53876a,a53877a,a53881a,a53882a,a53883a,a53887a,a53888a,a53891a,a53894a,a53895a,a53896a,a53900a,a53901a,a53905a,a53906a,a53907a,a53911a,a53912a,a53915a,a53918a,a53919a,a53920a,a53924a,a53925a,a53929a,a53930a,a53931a,a53935a,a53936a,a53939a,a53942a,a53943a,a53944a,a53948a,a53949a,a53953a,a53954a,a53955a,a53959a,a53960a,a53963a,a53966a,a53967a,a53968a,a53972a,a53973a,a53977a,a53978a,a53979a,a53983a,a53984a,a53987a,a53990a,a53991a,a53992a,a53996a,a53997a,a54001a,a54002a,a54003a,a54007a,a54008a,a54011a,a54014a,a54015a,a54016a,a54020a,a54021a,a54025a,a54026a,a54027a,a54031a,a54032a,a54035a,a54038a,a54039a,a54040a,a54044a,a54045a,a54049a,a54050a,a54051a,a54055a,a54056a,a54059a,a54062a,a54063a,a54064a,a54068a,a54069a,a54073a,a54074a,a54075a,a54079a,a54080a,a54083a,a54086a,a54087a,a54088a,a54092a,a54093a,a54097a,a54098a,a54099a,a54103a,a54104a,a54107a,a54110a,a54111a,a54112a,a54116a,a54117a,a54121a,a54122a,a54123a,a54127a,a54128a,a54131a,a54134a,a54135a,a54136a,a54140a,a54141a,a54145a,a54146a,a54147a,a54151a,a54152a,a54155a,a54158a,a54159a,a54160a,a54164a,a54165a,a54169a,a54170a,a54171a,a54175a,a54176a,a54179a,a54182a,a54183a,a54184a,a54188a,a54189a,a54193a,a54194a,a54195a,a54199a,a54200a,a54203a,a54206a,a54207a,a54208a,a54212a,a54213a,a54217a,a54218a,a54219a,a54223a,a54224a,a54227a,a54230a,a54231a,a54232a,a54236a,a54237a,a54241a,a54242a,a54243a,a54247a,a54248a,a54251a,a54254a,a54255a,a54256a,a54260a,a54261a,a54265a,a54266a,a54267a,a54271a,a54272a,a54275a,a54278a,a54279a,a54280a,a54284a,a54285a,a54289a,a54290a,a54291a,a54295a,a54296a,a54299a,a54302a,a54303a,a54304a,a54308a,a54309a,a54313a,a54314a,a54315a,a54319a,a54320a,a54323a,a54326a,a54327a,a54328a,a54332a,a54333a,a54337a,a54338a,a54339a,a54343a,a54344a,a54347a,a54350a,a54351a,a54352a,a54356a,a54357a,a54361a,a54362a,a54363a,a54367a,a54368a,a54371a,a54374a,a54375a,a54376a,a54380a,a54381a,a54385a,a54386a,a54387a,a54391a,a54392a,a54395a,a54398a,a54399a,a54400a,a54404a,a54405a,a54409a,a54410a,a54411a,a54415a,a54416a,a54419a,a54422a,a54423a,a54424a,a54428a,a54429a,a54433a,a54434a,a54435a,a54439a,a54440a,a54443a,a54446a,a54447a,a54448a,a54452a,a54453a,a54457a,a54458a,a54459a,a54463a,a54464a,a54467a,a54470a,a54471a,a54472a,a54476a,a54477a,a54481a,a54482a,a54483a,a54487a,a54488a,a54491a,a54494a,a54495a,a54496a,a54500a,a54501a,a54505a,a54506a,a54507a,a54511a,a54512a,a54515a,a54518a,a54519a,a54520a,a54524a,a54525a,a54529a,a54530a,a54531a,a54535a,a54536a,a54539a,a54542a,a54543a,a54544a,a54548a,a54549a,a54553a,a54554a,a54555a,a54559a,a54560a,a54563a,a54566a,a54567a,a54568a,a54572a,a54573a,a54577a,a54578a,a54579a,a54583a,a54584a,a54587a,a54590a,a54591a,a54592a,a54596a,a54597a,a54601a,a54602a,a54603a,a54607a,a54608a,a54611a,a54614a,a54615a,a54616a,a54620a,a54621a,a54625a,a54626a,a54627a,a54631a,a54632a,a54635a,a54638a,a54639a,a54640a,a54644a,a54645a,a54649a,a54650a,a54651a,a54655a,a54656a,a54659a,a54662a,a54663a,a54664a,a54668a,a54669a,a54673a,a54674a,a54675a,a54679a,a54680a,a54683a,a54686a,a54687a,a54688a,a54692a,a54693a,a54697a,a54698a,a54699a,a54703a,a54704a,a54707a,a54710a,a54711a,a54712a,a54716a,a54717a,a54721a,a54722a,a54723a,a54727a,a54728a,a54731a,a54734a,a54735a,a54736a,a54740a,a54741a,a54745a,a54746a,a54747a,a54751a,a54752a,a54755a,a54758a,a54759a,a54760a,a54764a,a54765a,a54769a,a54770a,a54771a,a54775a,a54776a,a54779a,a54782a,a54783a,a54784a,a54788a,a54789a,a54793a,a54794a,a54795a,a54799a,a54800a,a54803a,a54806a,a54807a,a54808a,a54812a,a54813a,a54817a,a54818a,a54819a,a54823a,a54824a,a54827a,a54830a,a54831a,a54832a,a54836a,a54837a,a54841a,a54842a,a54843a,a54847a,a54848a,a54851a,a54854a,a54855a,a54856a,a54860a,a54861a,a54865a,a54866a,a54867a,a54871a,a54872a,a54875a,a54878a,a54879a,a54880a,a54884a,a54885a,a54889a,a54890a,a54891a,a54895a,a54896a,a54899a,a54902a,a54903a,a54904a,a54908a,a54909a,a54913a,a54914a,a54915a,a54919a,a54920a,a54923a,a54926a,a54927a,a54928a,a54932a,a54933a,a54937a,a54938a,a54939a,a54943a,a54944a,a54947a,a54950a,a54951a,a54952a,a54956a,a54957a,a54961a,a54962a,a54963a,a54967a,a54968a,a54971a,a54974a,a54975a,a54976a,a54980a,a54981a,a54985a,a54986a,a54987a,a54991a,a54992a,a54995a,a54998a,a54999a,a55000a,a55004a,a55005a,a55009a,a55010a,a55011a,a55015a,a55016a,a55019a,a55022a,a55023a,a55024a,a55028a,a55029a,a55033a,a55034a,a55035a,a55039a,a55040a,a55043a,a55046a,a55047a,a55048a,a55052a,a55053a,a55057a,a55058a,a55059a,a55063a,a55064a,a55067a,a55070a,a55071a,a55072a,a55076a,a55077a,a55081a,a55082a,a55083a,a55087a,a55088a,a55091a,a55094a,a55095a,a55096a,a55100a,a55101a,a55105a,a55106a,a55107a,a55111a,a55112a,a55115a,a55118a,a55119a,a55120a,a55124a,a55125a,a55129a,a55130a,a55131a,a55135a,a55136a,a55139a,a55142a,a55143a,a55144a,a55148a,a55149a,a55153a,a55154a,a55155a,a55159a,a55160a,a55163a,a55166a,a55167a,a55168a,a55172a,a55173a,a55177a,a55178a,a55179a,a55183a,a55184a,a55187a,a55190a,a55191a,a55192a,a55196a,a55197a,a55201a,a55202a,a55203a,a55207a,a55208a,a55211a,a55214a,a55215a,a55216a,a55220a,a55221a,a55225a,a55226a,a55227a,a55231a,a55232a,a55235a,a55238a,a55239a,a55240a,a55244a,a55245a,a55249a,a55250a,a55251a,a55255a,a55256a,a55259a,a55262a,a55263a,a55264a,a55268a,a55269a,a55273a,a55274a,a55275a,a55279a,a55280a,a55283a,a55286a,a55287a,a55288a,a55292a,a55293a,a55297a,a55298a,a55299a,a55303a,a55304a,a55307a,a55310a,a55311a,a55312a,a55316a,a55317a,a55321a,a55322a,a55323a,a55327a,a55328a,a55331a,a55334a,a55335a,a55336a,a55340a,a55341a,a55345a,a55346a,a55347a,a55351a,a55352a,a55355a,a55358a,a55359a,a55360a,a55364a,a55365a,a55369a,a55370a,a55371a,a55375a,a55376a,a55379a,a55382a,a55383a,a55384a,a55388a,a55389a,a55393a,a55394a,a55395a,a55399a,a55400a,a55403a,a55406a,a55407a,a55408a,a55412a,a55413a,a55417a,a55418a,a55419a,a55423a,a55424a,a55427a,a55430a,a55431a,a55432a,a55436a,a55437a,a55441a,a55442a,a55443a,a55447a,a55448a,a55451a,a55454a,a55455a,a55456a,a55460a,a55461a,a55465a,a55466a,a55467a,a55471a,a55472a,a55475a,a55478a,a55479a,a55480a,a55484a,a55485a,a55489a,a55490a,a55491a,a55495a,a55496a,a55499a,a55502a,a55503a,a55504a,a55508a,a55509a,a55513a,a55514a,a55515a,a55519a,a55520a,a55523a,a55526a,a55527a,a55528a,a55532a,a55533a,a55537a,a55538a,a55539a,a55543a,a55544a,a55547a,a55550a,a55551a,a55552a,a55556a,a55557a,a55561a,a55562a,a55563a,a55567a,a55568a,a55571a,a55574a,a55575a,a55576a,a55580a,a55581a,a55585a,a55586a,a55587a,a55591a,a55592a,a55595a,a55598a,a55599a,a55600a,a55604a,a55605a,a55609a,a55610a,a55611a,a55615a,a55616a,a55619a,a55622a,a55623a,a55624a,a55628a,a55629a,a55633a,a55634a,a55635a,a55639a,a55640a,a55643a,a55646a,a55647a,a55648a,a55652a,a55653a,a55657a,a55658a,a55659a,a55663a,a55664a,a55667a,a55670a,a55671a,a55672a,a55676a,a55677a,a55681a,a55682a,a55683a,a55687a,a55688a,a55691a,a55694a,a55695a,a55696a,a55700a,a55701a,a55705a,a55706a,a55707a,a55711a,a55712a,a55715a,a55718a,a55719a,a55720a,a55724a,a55725a,a55729a,a55730a,a55731a,a55735a,a55736a,a55739a,a55742a,a55743a,a55744a,a55748a,a55749a,a55753a,a55754a,a55755a,a55759a,a55760a,a55763a,a55766a,a55767a,a55768a,a55772a,a55773a,a55777a,a55778a,a55779a,a55783a,a55784a,a55787a,a55790a,a55791a,a55792a,a55796a,a55797a,a55801a,a55802a,a55803a,a55807a,a55808a,a55811a,a55814a,a55815a,a55816a,a55820a,a55821a,a55825a,a55826a,a55827a,a55831a,a55832a,a55835a,a55838a,a55839a,a55840a,a55844a,a55845a,a55849a,a55850a,a55851a,a55855a,a55856a,a55859a,a55862a,a55863a,a55864a,a55868a,a55869a,a55873a,a55874a,a55875a,a55879a,a55880a,a55883a,a55886a,a55887a,a55888a,a55892a,a55893a,a55897a,a55898a,a55899a,a55903a,a55904a,a55907a,a55910a,a55911a,a55912a,a55916a,a55917a,a55921a,a55922a,a55923a,a55927a,a55928a,a55931a,a55934a,a55935a,a55936a,a55940a,a55941a,a55945a,a55946a,a55947a,a55951a,a55952a,a55955a,a55958a,a55959a,a55960a,a55964a,a55965a,a55969a,a55970a,a55971a,a55975a,a55976a,a55979a,a55982a,a55983a,a55984a,a55988a,a55989a,a55993a,a55994a,a55995a,a55999a,a56000a,a56003a,a56006a,a56007a,a56008a,a56012a,a56013a,a56017a,a56018a,a56019a,a56023a,a56024a,a56027a,a56030a,a56031a,a56032a,a56036a,a56037a,a56041a,a56042a,a56043a,a56047a,a56048a,a56051a,a56054a,a56055a,a56056a,a56060a,a56061a,a56065a,a56066a,a56067a,a56071a,a56072a,a56075a,a56078a,a56079a,a56080a,a56084a,a56085a,a56089a,a56090a,a56091a,a56095a,a56096a,a56099a,a56102a,a56103a,a56104a,a56108a,a56109a,a56113a,a56114a,a56115a,a56119a,a56120a,a56123a,a56126a,a56127a,a56128a,a56132a,a56133a,a56137a,a56138a,a56139a,a56143a,a56144a,a56147a,a56150a,a56151a,a56152a,a56156a,a56157a,a56161a,a56162a,a56163a,a56167a,a56168a,a56171a,a56174a,a56175a,a56176a,a56180a,a56181a,a56185a,a56186a,a56187a,a56191a,a56192a,a56195a,a56198a,a56199a,a56200a,a56204a,a56205a,a56209a,a56210a,a56211a,a56215a,a56216a,a56219a,a56222a,a56223a,a56224a,a56228a,a56229a,a56233a,a56234a,a56235a,a56239a,a56240a,a56243a,a56246a,a56247a,a56248a,a56252a,a56253a,a56257a,a56258a,a56259a,a56263a,a56264a,a56267a,a56270a,a56271a,a56272a,a56276a,a56277a,a56281a,a56282a,a56283a,a56287a,a56288a,a56291a,a56294a,a56295a,a56296a,a56300a,a56301a,a56305a,a56306a,a56307a,a56311a,a56312a,a56315a,a56318a,a56319a,a56320a,a56324a,a56325a,a56329a,a56330a,a56331a,a56335a,a56336a,a56339a,a56342a,a56343a,a56344a,a56348a,a56349a,a56353a,a56354a,a56355a,a56359a,a56360a,a56363a,a56366a,a56367a,a56368a,a56372a,a56373a,a56377a,a56378a,a56379a,a56383a,a56384a,a56387a,a56390a,a56391a,a56392a,a56396a,a56397a,a56401a,a56402a,a56403a,a56407a,a56408a,a56411a,a56414a,a56415a,a56416a,a56420a,a56421a,a56425a,a56426a,a56427a,a56431a,a56432a,a56435a,a56438a,a56439a,a56440a,a56444a,a56445a,a56449a,a56450a,a56451a,a56455a,a56456a,a56459a,a56462a,a56463a,a56464a,a56468a,a56469a,a56473a,a56474a,a56475a,a56479a,a56480a,a56483a,a56486a,a56487a,a56488a,a56492a,a56493a,a56497a,a56498a,a56499a,a56503a,a56504a,a56507a,a56510a,a56511a,a56512a,a56516a,a56517a,a56521a,a56522a,a56523a,a56527a,a56528a,a56531a,a56534a,a56535a,a56536a,a56540a,a56541a,a56545a,a56546a,a56547a,a56551a,a56552a,a56555a,a56558a,a56559a,a56560a,a56564a,a56565a,a56569a,a56570a,a56571a,a56575a,a56576a,a56579a,a56582a,a56583a,a56584a,a56588a,a56589a,a56593a,a56594a,a56595a,a56599a,a56600a,a56603a,a56606a,a56607a,a56608a,a56612a,a56613a,a56617a,a56618a,a56619a,a56623a,a56624a,a56627a,a56630a,a56631a,a56632a,a56636a,a56637a,a56641a,a56642a,a56643a,a56647a,a56648a,a56651a,a56654a,a56655a,a56656a,a56660a,a56661a,a56665a,a56666a,a56667a,a56671a,a56672a,a56675a,a56678a,a56679a,a56680a,a56684a,a56685a,a56689a,a56690a,a56691a,a56695a,a56696a,a56699a,a56702a,a56703a,a56704a,a56708a,a56709a,a56713a,a56714a,a56715a,a56719a,a56720a,a56723a,a56726a,a56727a,a56728a,a56732a,a56733a,a56737a,a56738a,a56739a,a56743a,a56744a,a56747a,a56750a,a56751a,a56752a,a56756a,a56757a,a56761a,a56762a,a56763a,a56767a,a56768a,a56771a,a56774a,a56775a,a56776a,a56780a,a56781a,a56785a,a56786a,a56787a,a56791a,a56792a,a56795a,a56798a,a56799a,a56800a,a56804a,a56805a,a56809a,a56810a,a56811a,a56815a,a56816a,a56819a,a56822a,a56823a,a56824a,a56828a,a56829a,a56833a,a56834a,a56835a,a56839a,a56840a,a56843a,a56846a,a56847a,a56848a,a56852a,a56853a,a56857a,a56858a,a56859a,a56863a,a56864a,a56867a,a56870a,a56871a,a56872a,a56876a,a56877a,a56881a,a56882a,a56883a,a56887a,a56888a,a56891a,a56894a,a56895a,a56896a,a56900a,a56901a,a56905a,a56906a,a56907a,a56911a,a56912a,a56915a,a56918a,a56919a,a56920a,a56924a,a56925a,a56929a,a56930a,a56931a,a56935a,a56936a,a56939a,a56942a,a56943a,a56944a,a56948a,a56949a,a56953a,a56954a,a56955a,a56959a,a56960a,a56963a,a56966a,a56967a,a56968a,a56972a,a56973a,a56977a,a56978a,a56979a,a56983a,a56984a,a56987a,a56990a,a56991a,a56992a,a56996a,a56997a,a57001a,a57002a,a57003a,a57007a,a57008a,a57011a,a57014a,a57015a,a57016a,a57020a,a57021a,a57025a,a57026a,a57027a,a57031a,a57032a,a57035a,a57038a,a57039a,a57040a,a57044a,a57045a,a57049a,a57050a,a57051a,a57055a,a57056a,a57059a,a57062a,a57063a,a57064a,a57068a,a57069a,a57073a,a57074a,a57075a,a57079a,a57080a,a57083a,a57086a,a57087a,a57088a,a57092a,a57093a,a57097a,a57098a,a57099a,a57103a,a57104a,a57107a,a57110a,a57111a,a57112a,a57116a,a57117a,a57121a,a57122a,a57123a,a57127a,a57128a,a57131a,a57134a,a57135a,a57136a,a57140a,a57141a,a57145a,a57146a,a57147a,a57151a,a57152a,a57155a,a57158a,a57159a,a57160a,a57164a,a57165a,a57169a,a57170a,a57171a,a57175a,a57176a,a57179a,a57182a,a57183a,a57184a,a57188a,a57189a,a57193a,a57194a,a57195a,a57199a,a57200a,a57203a,a57206a,a57207a,a57208a,a57212a,a57213a,a57217a,a57218a,a57219a,a57223a,a57224a,a57227a,a57230a,a57231a,a57232a,a57236a,a57237a,a57241a,a57242a,a57243a,a57247a,a57248a,a57251a,a57254a,a57255a,a57256a,a57260a,a57261a,a57265a,a57266a,a57267a,a57271a,a57272a,a57275a,a57278a,a57279a,a57280a,a57284a,a57285a,a57289a,a57290a,a57291a,a57295a,a57296a,a57299a,a57302a,a57303a,a57304a,a57308a,a57309a,a57313a,a57314a,a57315a,a57319a,a57320a,a57323a,a57326a,a57327a,a57328a,a57332a,a57333a,a57337a,a57338a,a57339a,a57343a,a57344a,a57347a,a57350a,a57351a,a57352a,a57356a,a57357a,a57361a,a57362a,a57363a,a57367a,a57368a,a57371a,a57374a,a57375a,a57376a,a57380a,a57381a,a57385a,a57386a,a57387a,a57391a,a57392a,a57395a,a57398a,a57399a,a57400a,a57404a,a57405a,a57409a,a57410a,a57411a,a57415a,a57416a,a57419a,a57422a,a57423a,a57424a,a57428a,a57429a,a57433a,a57434a,a57435a,a57439a,a57440a,a57443a,a57446a,a57447a,a57448a,a57452a,a57453a,a57457a,a57458a,a57459a,a57463a,a57464a,a57467a,a57470a,a57471a,a57472a,a57476a,a57477a,a57481a,a57482a,a57483a,a57487a,a57488a,a57491a,a57494a,a57495a,a57496a,a57500a,a57501a,a57505a,a57506a,a57507a,a57511a,a57512a,a57515a,a57518a,a57519a,a57520a,a57524a,a57525a,a57529a,a57530a,a57531a,a57535a,a57536a,a57539a,a57542a,a57543a,a57544a,a57548a,a57549a,a57553a,a57554a,a57555a,a57559a,a57560a,a57563a,a57566a,a57567a,a57568a,a57572a,a57573a,a57577a,a57578a,a57579a,a57583a,a57584a,a57587a,a57590a,a57591a,a57592a,a57596a,a57597a,a57601a,a57602a,a57603a,a57607a,a57608a,a57611a,a57614a,a57615a,a57616a,a57620a,a57621a,a57625a,a57626a,a57627a,a57631a,a57632a,a57635a,a57638a,a57639a,a57640a,a57644a,a57645a,a57649a,a57650a,a57651a,a57655a,a57656a,a57659a,a57662a,a57663a,a57664a,a57668a,a57669a,a57673a,a57674a,a57675a,a57679a,a57680a,a57683a,a57686a,a57687a,a57688a,a57692a,a57693a,a57697a,a57698a,a57699a,a57703a,a57704a,a57707a,a57710a,a57711a,a57712a,a57716a,a57717a,a57721a,a57722a,a57723a,a57727a,a57728a,a57731a,a57734a,a57735a,a57736a,a57740a,a57741a,a57745a,a57746a,a57747a,a57751a,a57752a,a57755a,a57758a,a57759a,a57760a,a57764a,a57765a,a57769a,a57770a,a57771a,a57775a,a57776a,a57779a,a57782a,a57783a,a57784a,a57788a,a57789a,a57793a,a57794a,a57795a,a57799a,a57800a,a57803a,a57806a,a57807a,a57808a,a57812a,a57813a,a57817a,a57818a,a57819a,a57823a,a57824a,a57827a,a57830a,a57831a,a57832a,a57836a,a57837a,a57841a,a57842a,a57843a,a57847a,a57848a,a57851a,a57854a,a57855a,a57856a,a57860a,a57861a,a57865a,a57866a,a57867a,a57871a,a57872a,a57875a,a57878a,a57879a,a57880a,a57884a,a57885a,a57889a,a57890a,a57891a,a57895a,a57896a,a57899a,a57902a,a57903a,a57904a,a57908a,a57909a,a57913a,a57914a,a57915a,a57919a,a57920a,a57923a,a57926a,a57927a,a57928a,a57932a,a57933a,a57937a,a57938a,a57939a,a57943a,a57944a,a57947a,a57950a,a57951a,a57952a,a57956a,a57957a,a57961a,a57962a,a57963a,a57967a,a57968a,a57971a,a57974a,a57975a,a57976a,a57980a,a57981a,a57985a,a57986a,a57987a,a57991a,a57992a,a57995a,a57998a,a57999a,a58000a,a58004a,a58005a,a58009a,a58010a,a58011a,a58015a,a58016a,a58019a,a58022a,a58023a,a58024a,a58028a,a58029a,a58033a,a58034a,a58035a,a58039a,a58040a,a58043a,a58046a,a58047a,a58048a,a58052a,a58053a,a58057a,a58058a,a58059a,a58063a,a58064a,a58067a,a58070a,a58071a,a58072a,a58076a,a58077a,a58081a,a58082a,a58083a,a58087a,a58088a,a58091a,a58094a,a58095a,a58096a,a58100a,a58101a,a58105a,a58106a,a58107a,a58111a,a58112a,a58115a,a58118a,a58119a,a58120a,a58124a,a58125a,a58129a,a58130a,a58131a,a58135a,a58136a,a58139a,a58142a,a58143a,a58144a,a58148a,a58149a,a58153a,a58154a,a58155a,a58159a,a58160a,a58163a,a58166a,a58167a,a58168a,a58172a,a58173a,a58177a,a58178a,a58179a,a58183a,a58184a,a58187a,a58190a,a58191a,a58192a,a58196a,a58197a,a58201a,a58202a,a58203a,a58207a,a58208a,a58211a,a58214a,a58215a,a58216a,a58220a,a58221a,a58225a,a58226a,a58227a,a58231a,a58232a,a58235a,a58238a,a58239a,a58240a,a58244a,a58245a,a58249a,a58250a,a58251a,a58255a,a58256a,a58259a,a58262a,a58263a,a58264a,a58268a,a58269a,a58273a,a58274a,a58275a,a58279a,a58280a,a58283a,a58286a,a58287a,a58288a,a58292a,a58293a,a58297a,a58298a,a58299a,a58303a,a58304a,a58307a,a58310a,a58311a,a58312a,a58316a,a58317a,a58321a,a58322a,a58323a,a58327a,a58328a,a58331a,a58334a,a58335a,a58336a,a58340a,a58341a,a58345a,a58346a,a58347a,a58351a,a58352a,a58355a,a58358a,a58359a,a58360a,a58364a,a58365a,a58369a,a58370a,a58371a,a58375a,a58376a,a58379a,a58382a,a58383a,a58384a,a58388a,a58389a,a58393a,a58394a,a58395a,a58399a,a58400a,a58403a,a58406a,a58407a,a58408a,a58412a,a58413a,a58417a,a58418a,a58419a,a58423a,a58424a,a58427a,a58430a,a58431a,a58432a,a58436a,a58437a,a58441a,a58442a,a58443a,a58447a,a58448a,a58451a,a58454a,a58455a,a58456a,a58460a,a58461a,a58465a,a58466a,a58467a,a58471a,a58472a,a58475a,a58478a,a58479a,a58480a,a58484a,a58485a,a58489a,a58490a,a58491a,a58495a,a58496a,a58499a,a58502a,a58503a,a58504a,a58508a,a58509a,a58513a,a58514a,a58515a,a58519a,a58520a,a58523a,a58526a,a58527a,a58528a,a58532a,a58533a,a58537a,a58538a,a58539a,a58543a,a58544a,a58547a,a58550a,a58551a,a58552a,a58556a,a58557a,a58561a,a58562a,a58563a,a58567a,a58568a,a58571a,a58574a,a58575a,a58576a,a58580a,a58581a,a58585a,a58586a,a58587a,a58591a,a58592a,a58595a,a58598a,a58599a,a58600a,a58604a,a58605a,a58609a,a58610a,a58611a,a58615a,a58616a,a58619a,a58622a,a58623a,a58624a,a58628a,a58629a,a58633a,a58634a,a58635a,a58639a,a58640a,a58643a,a58646a,a58647a,a58648a,a58652a,a58653a,a58657a,a58658a,a58659a,a58663a,a58664a,a58667a,a58670a,a58671a,a58672a,a58676a,a58677a,a58681a,a58682a,a58683a,a58687a,a58688a,a58691a,a58694a,a58695a,a58696a,a58700a,a58701a,a58705a,a58706a,a58707a,a58711a,a58712a,a58715a,a58718a,a58719a,a58720a,a58724a,a58725a,a58729a,a58730a,a58731a,a58735a,a58736a,a58739a,a58742a,a58743a,a58744a,a58748a,a58749a,a58753a,a58754a,a58755a,a58759a,a58760a,a58763a,a58766a,a58767a,a58768a,a58772a,a58773a,a58777a,a58778a,a58779a,a58783a,a58784a,a58787a,a58790a,a58791a,a58792a,a58796a,a58797a,a58801a,a58802a,a58803a,a58807a,a58808a,a58811a,a58814a,a58815a,a58816a,a58820a,a58821a,a58825a,a58826a,a58827a,a58831a,a58832a,a58835a,a58838a,a58839a,a58840a,a58844a,a58845a,a58849a,a58850a,a58851a,a58855a,a58856a,a58859a,a58862a,a58863a,a58864a,a58868a,a58869a,a58873a,a58874a,a58875a,a58879a,a58880a,a58883a,a58886a,a58887a,a58888a,a58892a,a58893a,a58897a,a58898a,a58899a,a58903a,a58904a,a58907a,a58910a,a58911a,a58912a,a58916a,a58917a,a58921a,a58922a,a58923a,a58927a,a58928a,a58931a,a58934a,a58935a,a58936a,a58940a,a58941a,a58945a,a58946a,a58947a,a58951a,a58952a,a58955a,a58958a,a58959a,a58960a,a58964a,a58965a,a58969a,a58970a,a58971a,a58975a,a58976a,a58979a,a58982a,a58983a,a58984a,a58988a,a58989a,a58993a,a58994a,a58995a,a58999a,a59000a,a59003a,a59006a,a59007a,a59008a,a59012a,a59013a,a59017a,a59018a,a59019a,a59023a,a59024a,a59027a,a59030a,a59031a,a59032a,a59036a,a59037a,a59041a,a59042a,a59043a,a59047a,a59048a,a59051a,a59054a,a59055a,a59056a,a59060a,a59061a,a59065a,a59066a,a59067a,a59071a,a59072a,a59075a,a59078a,a59079a,a59080a,a59084a,a59085a,a59089a,a59090a,a59091a,a59095a,a59096a,a59099a,a59102a,a59103a,a59104a,a59108a,a59109a,a59113a,a59114a,a59115a,a59119a,a59120a,a59123a,a59126a,a59127a,a59128a,a59132a,a59133a,a59137a,a59138a,a59139a,a59143a,a59144a,a59147a,a59150a,a59151a,a59152a,a59156a,a59157a,a59161a,a59162a,a59163a,a59167a,a59168a,a59171a,a59174a,a59175a,a59176a,a59180a,a59181a,a59185a,a59186a,a59187a,a59191a,a59192a,a59195a,a59198a,a59199a,a59200a,a59204a,a59205a,a59209a,a59210a,a59211a,a59215a,a59216a,a59219a,a59222a,a59223a,a59224a,a59228a,a59229a,a59233a,a59234a,a59235a,a59239a,a59240a,a59243a,a59246a,a59247a,a59248a,a59252a,a59253a,a59257a,a59258a,a59259a,a59263a,a59264a,a59267a,a59270a,a59271a,a59272a,a59276a,a59277a,a59281a,a59282a,a59283a,a59287a,a59288a,a59291a,a59294a,a59295a,a59296a,a59300a,a59301a,a59305a,a59306a,a59307a,a59311a,a59312a,a59315a,a59318a,a59319a,a59320a,a59324a,a59325a,a59329a,a59330a,a59331a,a59335a,a59336a,a59339a,a59342a,a59343a,a59344a,a59348a,a59349a,a59353a,a59354a,a59355a,a59359a,a59360a,a59363a,a59366a,a59367a,a59368a,a59372a,a59373a,a59377a,a59378a,a59379a,a59383a,a59384a,a59387a,a59390a,a59391a,a59392a,a59396a,a59397a,a59401a,a59402a,a59403a,a59407a,a59408a,a59411a,a59414a,a59415a,a59416a,a59420a,a59421a,a59425a,a59426a,a59427a,a59431a,a59432a,a59435a,a59438a,a59439a,a59440a,a59444a,a59445a,a59449a,a59450a,a59451a,a59455a,a59456a,a59459a,a59462a,a59463a,a59464a,a59468a,a59469a,a59473a,a59474a,a59475a,a59479a,a59480a,a59483a,a59486a,a59487a,a59488a,a59492a,a59493a,a59497a,a59498a,a59499a,a59503a,a59504a,a59507a,a59510a,a59511a,a59512a,a59516a,a59517a,a59521a,a59522a,a59523a,a59527a,a59528a,a59531a,a59534a,a59535a,a59536a,a59540a,a59541a,a59545a,a59546a,a59547a,a59551a,a59552a,a59555a,a59558a,a59559a,a59560a,a59564a,a59565a,a59569a,a59570a,a59571a,a59575a,a59576a,a59579a,a59582a,a59583a,a59584a,a59588a,a59589a,a59593a,a59594a,a59595a,a59599a,a59600a,a59603a,a59606a,a59607a,a59608a,a59612a,a59613a,a59617a,a59618a,a59619a,a59623a,a59624a,a59627a,a59630a,a59631a,a59632a,a59636a,a59637a,a59641a,a59642a,a59643a,a59647a,a59648a,a59651a,a59654a,a59655a,a59656a,a59660a,a59661a,a59665a,a59666a,a59667a,a59671a,a59672a,a59675a,a59678a,a59679a,a59680a,a59684a,a59685a,a59689a,a59690a,a59691a,a59695a,a59696a,a59699a,a59702a,a59703a,a59704a,a59708a,a59709a,a59713a,a59714a,a59715a,a59719a,a59720a,a59723a,a59726a,a59727a,a59728a,a59732a,a59733a,a59737a,a59738a,a59739a,a59743a,a59744a,a59747a,a59750a,a59751a,a59752a,a59756a,a59757a,a59761a,a59762a,a59763a,a59767a,a59768a,a59771a,a59774a,a59775a,a59776a,a59780a,a59781a,a59785a,a59786a,a59787a,a59791a,a59792a,a59795a,a59798a,a59799a,a59800a,a59804a,a59805a,a59809a,a59810a,a59811a,a59815a,a59816a,a59819a,a59822a,a59823a,a59824a,a59828a,a59829a,a59833a,a59834a,a59835a,a59839a,a59840a,a59843a,a59846a,a59847a,a59848a,a59852a,a59853a,a59857a,a59858a,a59859a,a59863a,a59864a,a59867a,a59870a,a59871a,a59872a,a59876a,a59877a,a59881a,a59882a,a59883a,a59887a,a59888a,a59891a,a59894a,a59895a,a59896a,a59900a,a59901a,a59905a,a59906a,a59907a,a59911a,a59912a,a59915a,a59918a,a59919a,a59920a,a59924a,a59925a,a59929a,a59930a,a59931a,a59935a,a59936a,a59939a,a59942a,a59943a,a59944a,a59948a,a59949a,a59953a,a59954a,a59955a,a59959a,a59960a,a59963a,a59966a,a59967a,a59968a,a59972a,a59973a,a59977a,a59978a,a59979a,a59983a,a59984a,a59987a,a59990a,a59991a,a59992a,a59996a,a59997a,a60001a,a60002a,a60003a,a60007a,a60008a,a60011a,a60014a,a60015a,a60016a,a60020a,a60021a,a60025a,a60026a,a60027a,a60031a,a60032a,a60035a,a60038a,a60039a,a60040a,a60044a,a60045a,a60049a,a60050a,a60051a,a60055a,a60056a,a60059a,a60062a,a60063a,a60064a,a60068a,a60069a,a60073a,a60074a,a60075a,a60079a,a60080a,a60083a,a60086a,a60087a,a60088a,a60092a,a60093a,a60097a,a60098a,a60099a,a60103a,a60104a,a60107a,a60110a,a60111a,a60112a,a60116a,a60117a,a60120a,a60123a,a60124a,a60125a,a60129a,a60130a,a60133a,a60136a,a60137a,a60138a,a60142a,a60143a,a60146a,a60149a,a60150a,a60151a,a60155a,a60156a,a60159a,a60162a,a60163a,a60164a,a60168a,a60169a,a60172a,a60175a,a60176a,a60177a,a60181a,a60182a,a60185a,a60188a,a60189a,a60190a,a60194a,a60195a,a60198a,a60201a,a60202a,a60203a,a60207a,a60208a,a60211a,a60214a,a60215a,a60216a,a60220a,a60221a,a60224a,a60227a,a60228a,a60229a,a60233a,a60234a,a60237a,a60240a,a60241a,a60242a,a60246a,a60247a,a60250a,a60253a,a60254a,a60255a,a60259a,a60260a,a60263a,a60266a,a60267a,a60268a,a60272a,a60273a,a60276a,a60279a,a60280a,a60281a,a60285a,a60286a,a60289a,a60292a,a60293a,a60294a,a60298a,a60299a,a60302a,a60305a,a60306a,a60307a,a60311a,a60312a,a60315a,a60318a,a60319a,a60320a,a60324a,a60325a,a60328a,a60331a,a60332a,a60333a,a60337a,a60338a,a60341a,a60344a,a60345a,a60346a,a60350a,a60351a,a60354a,a60357a,a60358a,a60359a,a60363a,a60364a,a60367a,a60370a,a60371a,a60372a,a60376a,a60377a,a60380a,a60383a,a60384a,a60385a,a60389a,a60390a,a60393a,a60396a,a60397a,a60398a,a60402a,a60403a,a60406a,a60409a,a60410a,a60411a,a60415a,a60416a,a60419a,a60422a,a60423a,a60424a,a60428a,a60429a,a60432a,a60435a,a60436a,a60437a,a60441a,a60442a,a60445a,a60448a,a60449a,a60450a,a60454a,a60455a,a60458a,a60461a,a60462a,a60463a,a60467a,a60468a,a60471a,a60474a,a60475a,a60476a,a60480a,a60481a,a60484a,a60487a,a60488a,a60489a,a60493a,a60494a,a60497a,a60500a,a60501a,a60502a,a60506a,a60507a,a60510a,a60513a,a60514a,a60515a,a60519a,a60520a,a60523a,a60526a,a60527a,a60528a,a60532a,a60533a,a60536a,a60539a,a60540a,a60541a,a60545a,a60546a,a60549a,a60552a,a60553a,a60554a,a60558a,a60559a,a60562a,a60565a,a60566a,a60567a,a60571a,a60572a,a60575a,a60578a,a60579a,a60580a,a60584a,a60585a,a60588a,a60591a,a60592a,a60593a,a60597a,a60598a,a60601a,a60604a,a60605a,a60606a,a60610a,a60611a,a60614a,a60617a,a60618a,a60619a,a60623a,a60624a,a60627a,a60630a,a60631a,a60632a,a60636a,a60637a,a60640a,a60643a,a60644a,a60645a,a60649a,a60650a,a60653a,a60656a,a60657a,a60658a,a60662a,a60663a,a60666a,a60669a,a60670a,a60671a,a60675a,a60676a,a60679a,a60682a,a60683a,a60684a,a60688a,a60689a,a60692a,a60695a,a60696a,a60697a,a60701a,a60702a,a60705a,a60708a,a60709a,a60710a,a60714a,a60715a,a60718a,a60721a,a60722a,a60723a,a60727a,a60728a,a60731a,a60734a,a60735a,a60736a,a60740a,a60741a,a60744a,a60747a,a60748a,a60749a,a60753a,a60754a,a60757a,a60760a,a60761a,a60762a,a60766a,a60767a,a60770a,a60773a,a60774a,a60775a,a60779a,a60780a,a60783a,a60786a,a60787a,a60788a,a60792a,a60793a,a60796a,a60799a,a60800a,a60801a,a60805a,a60806a,a60809a,a60812a,a60813a,a60814a,a60818a,a60819a,a60822a,a60825a,a60826a,a60827a,a60831a,a60832a,a60835a,a60838a,a60839a,a60840a,a60844a,a60845a,a60848a,a60851a,a60852a,a60853a,a60857a,a60858a,a60861a,a60864a,a60865a,a60866a,a60870a,a60871a,a60874a,a60877a,a60878a,a60879a,a60883a,a60884a,a60887a,a60890a,a60891a,a60892a,a60896a,a60897a,a60900a,a60903a,a60904a,a60905a,a60909a,a60910a,a60913a,a60916a,a60917a,a60918a,a60922a,a60923a,a60926a,a60929a,a60930a,a60931a,a60935a,a60936a,a60939a,a60942a,a60943a,a60944a,a60948a,a60949a,a60952a,a60955a,a60956a,a60957a,a60961a,a60962a,a60965a,a60968a,a60969a,a60970a,a60974a,a60975a,a60978a,a60981a,a60982a,a60983a,a60987a,a60988a,a60991a,a60994a,a60995a,a60996a,a61000a,a61001a,a61004a,a61007a,a61008a,a61009a,a61013a,a61014a,a61017a,a61020a,a61021a,a61022a,a61026a,a61027a,a61030a,a61033a,a61034a,a61035a,a61039a,a61040a,a61043a,a61046a,a61047a,a61048a,a61052a,a61053a,a61056a,a61059a,a61060a,a61061a,a61065a,a61066a,a61069a,a61072a,a61073a,a61074a,a61078a,a61079a,a61082a,a61085a,a61086a,a61087a,a61091a,a61092a,a61095a,a61098a,a61099a,a61100a,a61104a,a61105a,a61108a,a61111a,a61112a,a61113a,a61117a,a61118a,a61121a,a61124a,a61125a,a61126a,a61130a,a61131a,a61134a,a61137a,a61138a,a61139a,a61143a,a61144a,a61147a,a61150a,a61151a,a61152a,a61156a,a61157a,a61160a,a61163a,a61164a,a61165a,a61169a,a61170a,a61173a,a61176a,a61177a,a61178a,a61182a,a61183a,a61186a,a61189a,a61190a,a61191a,a61195a,a61196a,a61199a,a61202a,a61203a,a61204a,a61208a,a61209a,a61212a,a61215a,a61216a,a61217a,a61221a,a61222a,a61225a,a61228a,a61229a,a61230a,a61234a,a61235a,a61238a,a61241a,a61242a,a61243a,a61247a,a61248a,a61251a,a61254a,a61255a,a61256a,a61260a,a61261a,a61264a,a61267a,a61268a,a61269a,a61273a,a61274a,a61277a,a61280a,a61281a,a61282a,a61286a,a61287a,a61290a,a61293a,a61294a,a61295a,a61299a,a61300a,a61303a,a61306a,a61307a,a61308a,a61312a,a61313a,a61316a,a61319a,a61320a,a61321a,a61325a,a61326a,a61329a,a61332a,a61333a,a61334a,a61338a,a61339a,a61342a,a61345a,a61346a,a61347a,a61351a,a61352a,a61355a,a61358a,a61359a,a61360a,a61364a,a61365a,a61368a,a61371a,a61372a,a61373a,a61377a,a61378a,a61381a,a61384a,a61385a,a61386a,a61390a,a61391a,a61394a,a61397a,a61398a,a61399a,a61403a,a61404a,a61407a,a61410a,a61411a,a61412a,a61416a,a61417a,a61420a,a61423a,a61424a,a61425a,a61429a,a61430a,a61433a,a61436a,a61437a,a61438a,a61442a,a61443a,a61446a,a61449a,a61450a,a61451a,a61455a,a61456a,a61459a,a61462a,a61463a,a61464a,a61468a,a61469a,a61472a,a61475a,a61476a,a61477a,a61481a,a61482a,a61485a,a61488a,a61489a,a61490a,a61494a,a61495a,a61498a,a61501a,a61502a,a61503a,a61507a,a61508a,a61511a,a61514a,a61515a,a61516a,a61520a,a61521a,a61524a,a61527a,a61528a,a61529a,a61533a,a61534a,a61537a,a61540a,a61541a,a61542a,a61546a,a61547a,a61550a,a61553a,a61554a,a61555a,a61559a,a61560a,a61563a,a61566a,a61567a,a61568a,a61572a,a61573a,a61576a,a61579a,a61580a,a61581a,a61585a,a61586a,a61589a,a61592a,a61593a,a61594a,a61598a,a61599a,a61602a,a61605a,a61606a,a61607a,a61611a,a61612a,a61615a,a61618a,a61619a,a61620a,a61624a,a61625a,a61628a,a61631a,a61632a,a61633a,a61637a,a61638a,a61641a,a61644a,a61645a,a61646a,a61650a,a61651a,a61654a,a61657a,a61658a,a61659a,a61663a,a61664a,a61667a,a61670a,a61671a,a61672a,a61676a,a61677a,a61680a,a61683a,a61684a,a61685a,a61689a,a61690a,a61693a,a61696a,a61697a,a61698a,a61702a,a61703a,a61706a,a61709a,a61710a,a61711a,a61715a,a61716a,a61719a,a61722a,a61723a,a61724a,a61728a,a61729a,a61732a,a61735a,a61736a,a61737a,a61741a,a61742a,a61745a,a61748a,a61749a,a61750a,a61754a,a61755a,a61758a,a61761a,a61762a,a61763a,a61767a,a61768a,a61771a,a61774a,a61775a,a61776a,a61780a,a61781a,a61784a,a61787a,a61788a,a61789a,a61793a,a61794a,a61797a,a61800a,a61801a,a61802a,a61806a,a61807a,a61810a,a61813a,a61814a,a61815a,a61819a,a61820a,a61823a,a61826a,a61827a,a61828a,a61832a,a61833a,a61836a,a61839a,a61840a,a61841a,a61845a,a61846a,a61849a,a61852a,a61853a,a61854a,a61858a,a61859a,a61862a,a61865a,a61866a,a61867a,a61871a,a61872a,a61875a,a61878a,a61879a,a61880a,a61884a,a61885a,a61888a,a61891a,a61892a,a61893a,a61897a,a61898a,a61901a,a61904a,a61905a,a61906a,a61910a,a61911a,a61914a,a61917a,a61918a,a61919a,a61923a,a61924a,a61927a,a61930a,a61931a,a61932a,a61936a,a61937a,a61940a,a61943a,a61944a,a61945a,a61949a,a61950a,a61953a,a61956a,a61957a,a61958a,a61962a,a61963a,a61966a,a61969a,a61970a,a61971a,a61975a,a61976a,a61979a,a61982a,a61983a,a61984a,a61988a,a61989a,a61992a,a61995a,a61996a,a61997a,a62001a,a62002a,a62005a,a62008a,a62009a,a62010a,a62014a,a62015a,a62018a,a62021a,a62022a,a62023a,a62027a,a62028a,a62031a,a62034a,a62035a,a62036a,a62040a,a62041a,a62044a,a62047a,a62048a,a62049a,a62053a,a62054a,a62057a,a62060a,a62061a,a62062a,a62066a,a62067a,a62070a,a62073a,a62074a,a62075a,a62079a,a62080a,a62083a,a62086a,a62087a,a62088a,a62092a,a62093a,a62096a,a62099a,a62100a,a62101a,a62105a,a62106a,a62109a,a62112a,a62113a,a62114a,a62118a,a62119a,a62122a,a62125a,a62126a,a62127a,a62131a,a62132a,a62135a,a62138a,a62139a,a62140a,a62144a,a62145a,a62148a,a62151a,a62152a,a62153a,a62157a,a62158a,a62161a,a62164a,a62165a,a62166a,a62170a,a62171a,a62174a,a62177a,a62178a,a62179a,a62183a,a62184a,a62187a,a62190a,a62191a,a62192a,a62196a,a62197a,a62200a,a62203a,a62204a,a62205a,a62209a,a62210a,a62213a,a62216a,a62217a,a62218a,a62222a,a62223a,a62226a,a62229a,a62230a,a62231a,a62235a,a62236a,a62239a,a62242a,a62243a,a62244a,a62248a,a62249a,a62252a,a62255a,a62256a,a62257a,a62261a,a62262a,a62265a,a62268a,a62269a,a62270a,a62274a,a62275a,a62278a,a62281a,a62282a,a62283a,a62287a,a62288a,a62291a,a62294a,a62295a,a62296a,a62300a,a62301a,a62304a,a62307a,a62308a,a62309a,a62313a,a62314a,a62317a,a62320a,a62321a,a62322a,a62326a,a62327a,a62330a,a62333a,a62334a,a62335a,a62339a,a62340a,a62343a,a62346a,a62347a,a62348a,a62352a,a62353a,a62356a,a62359a,a62360a,a62361a,a62365a,a62366a,a62369a,a62372a,a62373a,a62374a,a62378a,a62379a,a62382a,a62385a,a62386a,a62387a,a62391a,a62392a,a62395a,a62398a,a62399a,a62400a,a62404a,a62405a,a62408a,a62411a,a62412a,a62413a,a62417a,a62418a,a62421a,a62424a,a62425a,a62426a,a62430a,a62431a,a62434a,a62437a,a62438a,a62439a,a62443a,a62444a,a62447a,a62450a,a62451a,a62452a,a62456a,a62457a,a62460a,a62463a,a62464a,a62465a,a62469a,a62470a,a62473a,a62476a,a62477a,a62478a,a62482a,a62483a,a62486a,a62489a,a62490a,a62491a,a62495a,a62496a,a62499a,a62502a,a62503a,a62504a,a62508a,a62509a,a62512a,a62515a,a62516a,a62517a,a62521a,a62522a,a62525a,a62528a,a62529a,a62530a,a62534a,a62535a,a62538a,a62541a,a62542a,a62543a,a62547a,a62548a,a62551a,a62554a,a62555a,a62556a,a62560a,a62561a,a62564a,a62567a,a62568a,a62569a,a62573a,a62574a,a62577a,a62580a,a62581a,a62582a,a62586a,a62587a,a62590a,a62593a,a62594a,a62595a,a62599a,a62600a,a62603a,a62606a,a62607a,a62608a,a62612a,a62613a,a62616a,a62619a,a62620a,a62621a,a62625a,a62626a,a62629a,a62632a,a62633a,a62634a,a62638a,a62639a,a62642a,a62645a,a62646a,a62647a,a62651a,a62652a,a62655a,a62658a,a62659a,a62660a,a62664a,a62665a,a62668a,a62671a,a62672a,a62673a,a62677a,a62678a,a62681a,a62684a,a62685a,a62686a,a62690a,a62691a,a62694a,a62697a,a62698a,a62699a,a62703a,a62704a,a62707a,a62710a,a62711a,a62712a,a62716a,a62717a,a62720a,a62723a,a62724a,a62725a,a62729a,a62730a,a62733a,a62736a,a62737a,a62738a,a62742a,a62743a,a62746a,a62749a,a62750a,a62751a,a62755a,a62756a,a62759a,a62762a,a62763a,a62764a,a62768a,a62769a,a62772a,a62775a,a62776a,a62777a,a62781a,a62782a,a62785a,a62788a,a62789a,a62790a,a62794a,a62795a,a62798a,a62801a,a62802a,a62803a,a62807a,a62808a,a62811a,a62814a,a62815a,a62816a,a62820a,a62821a,a62824a,a62827a,a62828a,a62829a,a62833a,a62834a,a62837a,a62840a,a62841a,a62842a,a62846a,a62847a,a62850a,a62853a,a62854a,a62855a,a62859a,a62860a,a62863a,a62866a,a62867a,a62868a,a62872a,a62873a,a62876a,a62879a,a62880a,a62881a,a62885a,a62886a,a62889a,a62892a,a62893a,a62894a,a62898a,a62899a,a62902a,a62905a,a62906a,a62907a,a62911a,a62912a,a62915a,a62918a,a62919a,a62920a,a62924a,a62925a,a62928a,a62931a,a62932a,a62933a,a62937a,a62938a,a62941a,a62944a,a62945a,a62946a,a62950a,a62951a,a62954a,a62957a,a62958a,a62959a,a62963a,a62964a,a62967a,a62970a,a62971a,a62972a,a62976a,a62977a,a62980a,a62983a,a62984a,a62985a,a62989a,a62990a,a62993a,a62996a,a62997a,a62998a,a63002a,a63003a,a63006a,a63009a,a63010a,a63011a,a63015a,a63016a,a63019a,a63022a,a63023a,a63024a,a63028a,a63029a,a63032a,a63035a,a63036a,a63037a,a63041a,a63042a,a63045a,a63048a,a63049a,a63050a,a63054a,a63055a,a63058a,a63061a,a63062a,a63063a,a63067a,a63068a,a63071a,a63074a,a63075a,a63076a,a63080a,a63081a,a63084a,a63087a,a63088a,a63089a,a63093a,a63094a,a63097a,a63100a,a63101a,a63102a,a63106a,a63107a,a63110a,a63113a,a63114a,a63115a,a63119a,a63120a,a63123a,a63126a,a63127a,a63128a,a63132a,a63133a,a63136a,a63139a,a63140a,a63141a,a63145a,a63146a,a63149a,a63152a,a63153a,a63154a,a63158a,a63159a,a63162a,a63165a,a63166a,a63167a,a63171a,a63172a,a63175a,a63178a,a63179a,a63180a,a63184a,a63185a,a63188a,a63191a,a63192a,a63193a,a63197a,a63198a,a63201a,a63204a,a63205a,a63206a,a63210a,a63211a,a63214a,a63217a,a63218a,a63219a,a63223a,a63224a,a63227a,a63230a,a63231a,a63232a,a63236a,a63237a,a63240a,a63243a,a63244a,a63245a,a63249a,a63250a,a63253a,a63256a,a63257a,a63258a,a63262a,a63263a,a63266a,a63269a,a63270a,a63271a,a63275a,a63276a,a63279a,a63282a,a63283a,a63284a,a63288a,a63289a,a63292a,a63295a,a63296a,a63297a,a63301a,a63302a,a63305a,a63308a,a63309a,a63310a,a63314a,a63315a,a63318a,a63321a,a63322a,a63323a,a63327a,a63328a,a63331a,a63334a,a63335a,a63336a,a63340a,a63341a,a63344a,a63347a,a63348a,a63349a,a63353a,a63354a,a63357a,a63360a,a63361a,a63362a,a63366a,a63367a,a63370a,a63373a,a63374a,a63375a,a63379a,a63380a,a63383a,a63386a,a63387a,a63388a,a63392a,a63393a,a63396a,a63399a,a63400a,a63401a,a63405a,a63406a,a63409a,a63412a,a63413a,a63414a,a63418a,a63419a,a63422a,a63425a,a63426a,a63427a,a63431a,a63432a,a63435a,a63438a,a63439a,a63440a,a63444a,a63445a,a63448a,a63451a,a63452a,a63453a,a63457a,a63458a,a63461a,a63464a,a63465a,a63466a,a63470a,a63471a,a63474a,a63477a,a63478a,a63479a,a63483a,a63484a,a63487a,a63490a,a63491a,a63492a,a63496a,a63497a,a63500a,a63503a,a63504a,a63505a,a63509a,a63510a,a63513a,a63516a,a63517a,a63518a,a63522a,a63523a,a63526a,a63529a,a63530a,a63531a,a63535a,a63536a,a63539a,a63542a,a63543a,a63544a,a63548a,a63549a,a63552a,a63555a,a63556a,a63557a,a63561a,a63562a,a63565a,a63568a,a63569a,a63570a,a63574a,a63575a,a63578a,a63581a,a63582a,a63583a,a63587a,a63588a,a63591a,a63594a,a63595a,a63596a,a63600a,a63601a,a63604a,a63607a,a63608a,a63609a,a63613a,a63614a,a63617a,a63620a,a63621a,a63622a,a63626a,a63627a,a63630a,a63633a,a63634a,a63635a,a63639a,a63640a,a63643a,a63646a,a63647a,a63648a,a63652a,a63653a,a63656a,a63659a,a63660a,a63661a,a63665a,a63666a,a63669a,a63672a,a63673a,a63674a,a63678a,a63679a,a63682a,a63685a,a63686a,a63687a,a63691a,a63692a,a63695a,a63698a,a63699a,a63700a,a63704a,a63705a,a63708a,a63711a,a63712a,a63713a,a63717a,a63718a,a63721a,a63724a,a63725a,a63726a,a63730a,a63731a,a63734a,a63737a,a63738a,a63739a,a63743a,a63744a,a63747a,a63750a,a63751a,a63752a,a63756a,a63757a,a63760a,a63763a,a63764a,a63765a,a63769a,a63770a,a63773a,a63776a,a63777a,a63778a,a63782a,a63783a,a63786a,a63789a,a63790a,a63791a,a63795a,a63796a,a63799a,a63802a,a63803a,a63804a,a63808a,a63809a,a63812a,a63815a,a63816a,a63817a,a63821a,a63822a,a63825a,a63828a,a63829a,a63830a,a63834a,a63835a,a63838a,a63841a,a63842a,a63843a,a63847a,a63848a,a63851a,a63854a,a63855a,a63856a,a63860a,a63861a,a63864a,a63867a,a63868a,a63869a,a63873a,a63874a,a63877a,a63880a,a63881a,a63882a,a63886a,a63887a,a63890a,a63893a,a63894a,a63895a,a63899a,a63900a,a63903a,a63906a,a63907a,a63908a,a63912a,a63913a,a63916a,a63919a,a63920a,a63921a,a63925a,a63926a,a63929a,a63932a,a63933a,a63934a,a63938a,a63939a,a63942a,a63945a,a63946a,a63947a,a63951a,a63952a,a63955a,a63958a,a63959a,a63960a,a63964a,a63965a,a63968a,a63971a,a63972a,a63973a,a63977a,a63978a,a63981a,a63984a,a63985a,a63986a,a63990a,a63991a,a63994a,a63997a,a63998a,a63999a,a64003a,a64004a,a64007a,a64010a,a64011a,a64012a,a64016a,a64017a,a64020a,a64023a,a64024a,a64025a,a64029a,a64030a,a64033a,a64036a,a64037a,a64038a,a64042a,a64043a,a64046a,a64049a,a64050a,a64051a,a64055a,a64056a,a64059a,a64062a,a64063a,a64064a,a64068a,a64069a,a64072a,a64075a,a64076a,a64077a,a64081a,a64082a,a64085a,a64088a,a64089a,a64090a,a64094a,a64095a,a64098a,a64101a,a64102a,a64103a,a64107a,a64108a,a64111a,a64114a,a64115a,a64116a,a64120a,a64121a,a64124a,a64127a,a64128a,a64129a,a64133a,a64134a,a64137a,a64140a,a64141a,a64142a,a64146a,a64147a,a64150a,a64153a,a64154a,a64155a,a64159a,a64160a,a64163a,a64166a,a64167a,a64168a,a64172a,a64173a,a64176a,a64179a,a64180a,a64181a,a64185a,a64186a,a64189a,a64192a,a64193a,a64194a,a64198a,a64199a,a64202a,a64205a,a64206a,a64207a,a64211a,a64212a,a64215a,a64218a,a64219a,a64220a,a64224a,a64225a,a64228a,a64231a,a64232a,a64233a,a64237a,a64238a,a64241a,a64244a,a64245a,a64246a,a64250a,a64251a,a64254a,a64257a,a64258a,a64259a,a64263a,a64264a,a64267a,a64270a,a64271a,a64272a,a64276a,a64277a,a64280a,a64283a,a64284a,a64285a,a64289a,a64290a,a64293a,a64296a,a64297a,a64298a,a64302a,a64303a,a64306a,a64309a,a64310a,a64311a,a64315a,a64316a,a64319a,a64322a,a64323a,a64324a,a64328a,a64329a,a64332a,a64335a,a64336a,a64337a,a64341a,a64342a,a64345a,a64348a,a64349a,a64350a,a64354a,a64355a,a64358a,a64361a,a64362a,a64363a,a64367a,a64368a,a64371a,a64374a,a64375a,a64376a,a64380a,a64381a,a64384a,a64387a,a64388a,a64389a,a64393a,a64394a,a64397a,a64400a,a64401a,a64402a,a64406a,a64407a,a64410a,a64413a,a64414a,a64415a,a64419a,a64420a,a64423a,a64426a,a64427a,a64428a,a64432a,a64433a,a64436a,a64439a,a64440a,a64441a,a64445a,a64446a,a64449a,a64452a,a64453a,a64454a,a64458a,a64459a,a64462a,a64465a,a64466a,a64467a,a64471a,a64472a,a64475a,a64478a,a64479a,a64480a,a64484a,a64485a,a64488a,a64491a,a64492a,a64493a,a64497a,a64498a,a64501a,a64504a,a64505a,a64506a,a64510a,a64511a,a64514a,a64517a,a64518a,a64519a,a64523a,a64524a,a64527a,a64530a,a64531a,a64532a,a64536a,a64537a,a64540a,a64543a,a64544a,a64545a,a64549a,a64550a,a64553a,a64556a,a64557a,a64558a,a64562a,a64563a,a64566a,a64569a,a64570a,a64571a,a64575a,a64576a,a64579a,a64582a,a64583a,a64584a,a64588a,a64589a,a64592a,a64595a,a64596a,a64597a,a64601a,a64602a,a64605a,a64608a,a64609a,a64610a,a64614a,a64615a,a64618a,a64621a,a64622a,a64623a,a64627a,a64628a,a64631a,a64634a,a64635a,a64636a,a64640a,a64641a,a64644a,a64647a,a64648a,a64649a,a64653a,a64654a,a64657a,a64660a,a64661a,a64662a,a64666a,a64667a,a64670a,a64673a,a64674a,a64675a,a64679a,a64680a,a64683a,a64686a,a64687a,a64688a,a64692a,a64693a,a64696a,a64699a,a64700a,a64701a,a64705a,a64706a,a64709a,a64712a,a64713a,a64714a,a64718a,a64719a,a64722a,a64725a,a64726a,a64727a,a64731a,a64732a,a64735a,a64738a,a64739a,a64740a,a64744a,a64745a,a64748a,a64751a,a64752a,a64753a,a64757a,a64758a,a64761a,a64764a,a64765a,a64766a,a64770a,a64771a,a64774a,a64777a,a64778a,a64779a,a64783a,a64784a,a64787a,a64790a,a64791a,a64792a,a64796a,a64797a,a64800a,a64803a,a64804a,a64805a,a64809a,a64810a,a64813a,a64816a,a64817a,a64818a,a64822a,a64823a,a64826a,a64829a,a64830a,a64831a,a64835a,a64836a,a64839a,a64842a,a64843a,a64844a,a64848a,a64849a,a64852a,a64855a,a64856a,a64857a,a64861a,a64862a,a64865a,a64868a,a64869a,a64870a,a64874a,a64875a,a64878a,a64881a,a64882a,a64883a,a64887a,a64888a,a64891a,a64894a,a64895a,a64896a,a64900a,a64901a,a64904a,a64907a,a64908a,a64909a,a64913a,a64914a,a64917a,a64920a,a64921a,a64922a,a64926a,a64927a,a64930a,a64933a,a64934a,a64935a,a64939a,a64940a,a64943a,a64946a,a64947a,a64948a,a64952a,a64953a,a64956a,a64959a,a64960a,a64961a,a64965a,a64966a,a64969a,a64972a,a64973a,a64974a,a64978a,a64979a,a64982a,a64985a,a64986a,a64987a,a64991a,a64992a,a64995a,a64998a,a64999a,a65000a,a65004a,a65005a,a65008a,a65011a,a65012a,a65013a,a65017a,a65018a,a65021a,a65024a,a65025a,a65026a,a65030a,a65031a,a65034a,a65037a,a65038a,a65039a,a65043a,a65044a,a65047a,a65050a,a65051a,a65052a,a65056a,a65057a,a65060a,a65063a,a65064a,a65065a,a65069a,a65070a,a65073a,a65076a,a65077a,a65078a,a65082a,a65083a,a65086a,a65089a,a65090a,a65091a,a65095a,a65096a,a65099a,a65102a,a65103a,a65104a,a65108a,a65109a,a65112a,a65115a,a65116a,a65117a,a65121a,a65122a,a65125a,a65128a,a65129a,a65130a,a65134a,a65135a,a65138a,a65141a,a65142a,a65143a,a65147a,a65148a,a65151a,a65154a,a65155a,a65156a,a65160a,a65161a,a65164a,a65167a,a65168a,a65169a,a65173a,a65174a,a65177a,a65180a,a65181a,a65182a,a65186a,a65187a,a65190a,a65193a,a65194a,a65195a,a65199a,a65200a,a65203a,a65206a,a65207a,a65208a,a65212a,a65213a,a65216a,a65219a,a65220a,a65221a,a65225a,a65226a,a65229a,a65232a,a65233a,a65234a,a65238a,a65239a,a65242a,a65245a,a65246a,a65247a,a65251a,a65252a,a65255a,a65258a,a65259a,a65260a,a65264a,a65265a,a65268a,a65271a,a65272a,a65273a,a65277a,a65278a,a65281a,a65284a,a65285a,a65286a,a65290a,a65291a,a65294a,a65297a,a65298a,a65299a,a65303a,a65304a,a65307a,a65310a,a65311a,a65312a,a65316a,a65317a,a65320a,a65323a,a65324a,a65325a,a65329a,a65330a,a65333a,a65336a,a65337a,a65338a,a65342a,a65343a,a65346a,a65349a,a65350a,a65351a,a65355a,a65356a,a65359a,a65362a,a65363a,a65364a,a65368a,a65369a,a65372a,a65375a,a65376a,a65377a,a65381a,a65382a,a65385a,a65388a,a65389a,a65390a,a65394a,a65395a,a65398a,a65401a,a65402a,a65403a,a65407a,a65408a,a65411a,a65414a,a65415a,a65416a,a65420a,a65421a,a65424a,a65427a,a65428a,a65429a,a65433a,a65434a,a65437a,a65440a,a65441a,a65442a,a65446a,a65447a,a65450a,a65453a,a65454a,a65455a,a65459a,a65460a,a65463a,a65466a,a65467a,a65468a,a65472a,a65473a,a65476a,a65479a,a65480a,a65481a,a65485a,a65486a,a65489a,a65492a,a65493a,a65494a,a65498a,a65499a,a65502a,a65505a,a65506a,a65507a,a65511a,a65512a,a65515a,a65518a,a65519a,a65520a,a65524a,a65525a,a65528a,a65531a,a65532a,a65533a,a65537a,a65538a,a65541a,a65544a,a65545a,a65546a,a65550a,a65551a,a65554a,a65557a,a65558a,a65559a,a65563a,a65564a,a65567a,a65570a,a65571a,a65572a,a65576a,a65577a,a65580a,a65583a,a65584a,a65585a,a65589a,a65590a,a65593a,a65596a,a65597a,a65598a,a65602a,a65603a,a65606a,a65609a,a65610a,a65611a,a65615a,a65616a,a65619a,a65622a,a65623a,a65624a,a65628a,a65629a,a65632a,a65635a,a65636a,a65637a,a65641a,a65642a,a65645a,a65648a,a65649a,a65650a,a65654a,a65655a,a65658a,a65661a,a65662a,a65663a,a65667a,a65668a,a65671a,a65674a,a65675a,a65676a,a65680a,a65681a,a65684a,a65687a,a65688a,a65689a,a65693a,a65694a,a65697a,a65700a,a65701a,a65702a,a65706a,a65707a,a65710a,a65713a,a65714a,a65715a,a65719a,a65720a,a65723a,a65726a,a65727a,a65728a,a65732a,a65733a,a65736a,a65739a,a65740a,a65741a,a65745a,a65746a,a65749a,a65752a,a65753a,a65754a,a65758a,a65759a,a65762a,a65765a,a65766a,a65767a,a65771a,a65772a,a65775a,a65778a,a65779a,a65780a,a65784a,a65785a,a65788a,a65791a,a65792a,a65793a,a65797a,a65798a,a65801a,a65804a,a65805a,a65806a,a65810a,a65811a,a65814a,a65817a,a65818a,a65819a,a65823a,a65824a,a65827a,a65830a,a65831a,a65832a,a65836a,a65837a,a65840a,a65843a,a65844a,a65845a,a65849a,a65850a,a65853a,a65856a,a65857a,a65858a,a65862a,a65863a,a65866a,a65869a,a65870a,a65871a,a65875a,a65876a,a65879a,a65882a,a65883a,a65884a,a65888a,a65889a,a65892a,a65895a,a65896a,a65897a,a65901a,a65902a,a65905a,a65908a,a65909a,a65910a,a65914a,a65915a,a65918a,a65921a,a65922a,a65923a,a65927a,a65928a,a65931a,a65934a,a65935a,a65936a,a65940a,a65941a,a65944a,a65947a,a65948a,a65949a,a65953a,a65954a,a65957a,a65960a,a65961a,a65962a,a65966a,a65967a,a65970a,a65973a,a65974a,a65975a,a65979a,a65980a,a65983a,a65986a,a65987a,a65988a,a65992a,a65993a,a65996a,a65999a,a66000a,a66001a,a66005a,a66006a,a66009a,a66012a,a66013a,a66014a,a66018a,a66019a,a66022a,a66025a,a66026a,a66027a,a66031a,a66032a,a66035a,a66038a,a66039a,a66040a,a66044a,a66045a,a66048a,a66051a,a66052a,a66053a,a66057a,a66058a,a66061a,a66064a,a66065a,a66066a,a66070a,a66071a,a66074a,a66077a,a66078a,a66079a,a66083a,a66084a,a66087a,a66090a,a66091a,a66092a,a66096a,a66097a,a66100a,a66103a,a66104a,a66105a,a66109a,a66110a,a66113a,a66116a,a66117a,a66118a,a66122a,a66123a,a66126a,a66129a,a66130a,a66131a,a66135a,a66136a,a66139a,a66142a,a66143a,a66144a,a66148a,a66149a,a66152a,a66155a,a66156a,a66157a,a66161a,a66162a,a66165a,a66168a,a66169a,a66170a,a66174a,a66175a,a66178a,a66181a,a66182a,a66183a,a66187a,a66188a,a66191a,a66194a,a66195a,a66196a,a66200a,a66201a,a66204a,a66207a,a66208a,a66209a,a66213a,a66214a,a66217a,a66220a,a66221a,a66222a,a66226a,a66227a,a66230a,a66233a,a66234a,a66235a,a66239a,a66240a,a66243a,a66246a,a66247a,a66248a,a66252a,a66253a,a66256a,a66259a,a66260a,a66261a,a66265a,a66266a,a66269a,a66272a,a66273a,a66274a,a66278a,a66279a,a66282a,a66285a,a66286a,a66287a,a66291a,a66292a,a66295a,a66298a,a66299a,a66300a,a66304a,a66305a,a66308a,a66311a,a66312a,a66313a,a66317a,a66318a,a66321a,a66324a,a66325a,a66326a,a66330a,a66331a,a66334a,a66337a,a66338a,a66339a,a66343a,a66344a,a66347a,a66350a,a66351a,a66352a,a66356a,a66357a,a66360a,a66363a,a66364a,a66365a,a66369a,a66370a,a66373a,a66376a,a66377a,a66378a,a66382a,a66383a,a66386a,a66389a,a66390a,a66391a,a66395a,a66396a,a66399a,a66402a,a66403a,a66404a,a66408a,a66409a,a66412a,a66415a,a66416a,a66417a,a66421a,a66422a,a66425a,a66428a,a66429a,a66430a,a66434a,a66435a,a66438a,a66441a,a66442a,a66443a,a66447a,a66448a,a66451a,a66454a,a66455a,a66456a,a66460a,a66461a,a66464a,a66467a,a66468a,a66469a,a66473a,a66474a,a66477a,a66480a,a66481a,a66482a,a66486a,a66487a,a66490a,a66493a,a66494a,a66495a,a66499a,a66500a,a66503a,a66506a,a66507a,a66508a,a66512a,a66513a,a66516a,a66519a,a66520a,a66521a,a66525a,a66526a,a66529a,a66532a,a66533a,a66534a,a66538a,a66539a,a66542a,a66545a,a66546a,a66547a,a66551a,a66552a,a66555a,a66558a,a66559a,a66560a,a66564a,a66565a,a66568a,a66571a,a66572a,a66573a,a66577a,a66578a,a66581a,a66584a,a66585a,a66586a,a66590a,a66591a,a66594a,a66597a,a66598a,a66599a,a66603a,a66604a,a66607a,a66610a,a66611a,a66612a,a66616a,a66617a,a66620a,a66623a,a66624a,a66625a,a66629a,a66630a,a66633a,a66636a,a66637a,a66638a,a66642a,a66643a,a66646a,a66649a,a66650a,a66651a,a66655a,a66656a,a66659a,a66662a,a66663a,a66664a,a66668a,a66669a,a66672a,a66675a,a66676a,a66677a,a66681a,a66682a,a66685a,a66688a,a66689a,a66690a,a66694a,a66695a,a66698a,a66701a,a66702a,a66703a,a66707a,a66708a,a66711a,a66714a,a66715a,a66716a,a66720a,a66721a,a66724a,a66727a,a66728a,a66729a,a66733a,a66734a,a66737a,a66740a,a66741a,a66742a,a66746a,a66747a,a66750a,a66753a,a66754a,a66755a,a66759a,a66760a,a66763a,a66766a,a66767a,a66768a,a66772a,a66773a,a66776a,a66779a,a66780a,a66781a,a66785a,a66786a,a66789a,a66792a,a66793a,a66794a,a66798a,a66799a,a66802a,a66805a,a66806a,a66807a,a66811a,a66812a,a66815a,a66818a,a66819a,a66820a,a66824a,a66825a,a66828a,a66831a,a66832a,a66833a,a66837a,a66838a,a66841a,a66844a,a66845a,a66846a,a66850a,a66851a,a66854a,a66857a,a66858a,a66859a,a66863a,a66864a,a66867a,a66870a,a66871a,a66872a,a66876a,a66877a,a66880a,a66883a,a66884a,a66885a,a66889a,a66890a,a66893a,a66896a,a66897a,a66898a,a66902a,a66903a,a66906a,a66909a,a66910a,a66911a,a66915a,a66916a,a66919a,a66922a,a66923a,a66924a,a66928a,a66929a,a66932a,a66935a,a66936a,a66937a,a66941a,a66942a,a66945a,a66948a,a66949a,a66950a,a66954a,a66955a,a66958a,a66961a,a66962a,a66963a,a66967a,a66968a,a66971a,a66974a,a66975a,a66976a,a66980a,a66981a,a66984a,a66987a,a66988a,a66989a,a66993a,a66994a,a66997a,a67000a,a67001a,a67002a,a67006a,a67007a,a67010a,a67013a,a67014a,a67015a,a67019a,a67020a,a67023a,a67026a,a67027a,a67028a,a67032a,a67033a,a67036a,a67039a,a67040a,a67041a,a67045a,a67046a,a67049a,a67052a,a67053a,a67054a,a67058a,a67059a,a67062a,a67065a,a67066a,a67067a,a67071a,a67072a,a67075a,a67078a,a67079a,a67080a,a67084a,a67085a,a67088a,a67091a,a67092a,a67093a,a67097a,a67098a,a67101a,a67104a,a67105a,a67106a,a67110a,a67111a,a67114a,a67117a,a67118a,a67119a,a67123a,a67124a,a67127a,a67130a,a67131a,a67132a,a67136a,a67137a,a67140a,a67143a,a67144a,a67145a,a67149a,a67150a,a67153a,a67156a,a67157a,a67158a,a67162a,a67163a,a67166a,a67169a,a67170a,a67171a,a67175a,a67176a,a67179a,a67182a,a67183a,a67184a,a67188a,a67189a,a67192a,a67195a,a67196a,a67197a,a67201a,a67202a,a67205a,a67208a,a67209a,a67210a,a67214a,a67215a,a67218a,a67221a,a67222a,a67223a,a67227a,a67228a,a67231a,a67234a,a67235a,a67236a,a67240a,a67241a,a67244a,a67247a,a67248a,a67249a,a67253a,a67254a,a67257a,a67260a,a67261a,a67262a,a67266a,a67267a,a67270a,a67273a,a67274a,a67275a,a67279a,a67280a,a67283a,a67286a,a67287a,a67288a,a67292a,a67293a,a67296a,a67299a,a67300a,a67301a,a67305a,a67306a,a67309a,a67312a,a67313a,a67314a,a67318a,a67319a,a67322a,a67325a,a67326a,a67327a,a67331a,a67332a,a67335a,a67338a,a67339a,a67340a,a67344a,a67345a,a67348a,a67351a,a67352a,a67353a,a67357a,a67358a,a67361a,a67364a,a67365a,a67366a,a67370a,a67371a,a67374a,a67377a,a67378a,a67379a,a67383a,a67384a,a67387a,a67390a,a67391a,a67392a,a67396a,a67397a,a67400a,a67403a,a67404a,a67405a,a67409a,a67410a,a67413a,a67416a,a67417a,a67418a,a67422a,a67423a,a67426a,a67429a,a67430a,a67431a,a67435a,a67436a,a67439a,a67442a,a67443a,a67444a,a67448a,a67449a,a67452a,a67455a,a67456a,a67457a,a67461a,a67462a,a67465a,a67468a,a67469a,a67470a,a67474a,a67475a,a67478a,a67481a,a67482a,a67483a,a67487a,a67488a,a67491a,a67494a,a67495a,a67496a,a67500a,a67501a,a67504a,a67507a,a67508a,a67509a,a67513a,a67514a,a67517a,a67520a,a67521a,a67522a,a67526a,a67527a,a67530a,a67533a,a67534a,a67535a,a67539a,a67540a,a67543a,a67546a,a67547a,a67548a,a67552a,a67553a,a67556a,a67559a,a67560a,a67561a,a67565a,a67566a,a67569a,a67572a,a67573a,a67574a,a67578a,a67579a,a67582a,a67585a,a67586a,a67587a,a67591a,a67592a,a67595a,a67598a,a67599a,a67600a,a67604a,a67605a,a67608a,a67611a,a67612a,a67613a,a67617a,a67618a,a67621a,a67624a,a67625a,a67626a,a67630a,a67631a,a67634a,a67637a,a67638a,a67639a,a67643a,a67644a,a67647a,a67650a,a67651a,a67652a,a67656a,a67657a,a67660a,a67663a,a67664a,a67665a,a67669a,a67670a,a67673a,a67676a,a67677a,a67678a,a67682a,a67683a,a67686a,a67689a,a67690a,a67691a,a67695a,a67696a,a67699a,a67702a,a67703a,a67704a,a67708a,a67709a,a67712a,a67715a,a67716a,a67717a,a67721a,a67722a,a67725a,a67728a,a67729a,a67730a,a67734a,a67735a,a67738a,a67741a,a67742a,a67743a,a67747a,a67748a,a67751a,a67754a,a67755a,a67756a,a67760a,a67761a,a67764a,a67767a,a67768a,a67769a,a67773a,a67774a,a67777a,a67780a,a67781a,a67782a,a67786a,a67787a,a67790a,a67793a,a67794a,a67795a,a67799a,a67800a,a67803a,a67806a,a67807a,a67808a,a67812a,a67813a,a67816a,a67819a,a67820a,a67821a,a67825a,a67826a,a67829a,a67832a,a67833a,a67834a,a67838a,a67839a,a67842a,a67845a,a67846a,a67847a,a67851a,a67852a,a67855a,a67858a,a67859a,a67860a,a67864a,a67865a,a67868a,a67871a,a67872a,a67873a,a67877a,a67878a,a67881a,a67884a,a67885a,a67886a,a67890a,a67891a,a67894a,a67897a,a67898a,a67899a,a67903a,a67904a,a67907a,a67910a,a67911a,a67912a,a67916a,a67917a,a67920a,a67923a,a67924a,a67925a,a67929a,a67930a,a67933a,a67936a,a67937a,a67938a,a67942a,a67943a,a67946a,a67949a,a67950a,a67951a,a67955a,a67956a,a67959a,a67962a,a67963a,a67964a,a67968a,a67969a,a67972a,a67975a,a67976a,a67977a,a67981a,a67982a,a67985a,a67988a,a67989a,a67990a,a67994a,a67995a,a67998a,a68001a,a68002a,a68003a,a68007a,a68008a,a68011a,a68014a,a68015a,a68016a,a68020a,a68021a,a68024a,a68027a,a68028a,a68029a,a68033a,a68034a,a68037a,a68040a,a68041a,a68042a,a68046a,a68047a,a68050a,a68053a,a68054a,a68055a,a68059a,a68060a,a68063a,a68066a,a68067a,a68068a,a68072a,a68073a,a68076a,a68079a,a68080a,a68081a,a68085a,a68086a,a68089a,a68092a,a68093a,a68094a,a68098a,a68099a,a68102a,a68105a,a68106a,a68107a,a68111a,a68112a,a68115a,a68118a,a68119a,a68120a,a68124a,a68125a,a68128a,a68131a,a68132a,a68133a,a68137a,a68138a,a68141a,a68144a,a68145a,a68146a,a68150a,a68151a,a68154a,a68157a,a68158a,a68159a,a68163a,a68164a,a68167a,a68170a,a68171a,a68172a,a68176a,a68177a,a68180a,a68183a,a68184a,a68185a,a68189a,a68190a,a68193a,a68196a,a68197a,a68198a,a68202a,a68203a,a68206a,a68209a,a68210a,a68211a,a68215a,a68216a,a68219a,a68222a,a68223a,a68224a,a68228a,a68229a,a68232a,a68235a,a68236a,a68237a,a68241a,a68242a,a68245a,a68248a,a68249a,a68250a,a68254a,a68255a,a68258a,a68261a,a68262a,a68263a,a68267a,a68268a,a68271a,a68274a,a68275a,a68276a,a68280a,a68281a,a68284a,a68287a,a68288a,a68289a,a68293a,a68294a,a68297a,a68300a,a68301a,a68302a,a68306a,a68307a,a68310a,a68313a,a68314a,a68315a,a68319a,a68320a,a68323a,a68326a,a68327a,a68328a,a68332a,a68333a,a68336a,a68339a,a68340a,a68341a,a68345a,a68346a,a68349a,a68352a,a68353a,a68354a,a68358a,a68359a,a68362a,a68365a,a68366a,a68367a,a68371a,a68372a,a68375a,a68378a,a68379a,a68380a,a68384a,a68385a,a68388a,a68391a,a68392a,a68393a,a68397a,a68398a,a68401a,a68404a,a68405a,a68406a,a68410a,a68411a,a68414a,a68417a,a68418a,a68419a,a68423a,a68424a,a68427a,a68430a,a68431a,a68432a,a68436a,a68437a,a68440a,a68443a,a68444a,a68445a,a68449a,a68450a,a68453a,a68456a,a68457a,a68458a,a68462a,a68463a,a68466a,a68469a,a68470a,a68471a,a68475a,a68476a,a68479a,a68482a,a68483a,a68484a,a68488a,a68489a,a68492a,a68495a,a68496a,a68497a,a68501a,a68502a,a68505a,a68508a,a68509a,a68510a,a68514a,a68515a,a68518a,a68521a,a68522a,a68523a,a68527a,a68528a,a68531a,a68534a,a68535a,a68536a,a68540a,a68541a,a68544a,a68547a,a68548a,a68549a,a68553a,a68554a,a68557a,a68560a,a68561a,a68562a,a68566a,a68567a,a68570a,a68573a,a68574a,a68575a,a68579a,a68580a,a68583a,a68586a,a68587a,a68588a,a68592a,a68593a,a68596a,a68599a,a68600a,a68601a,a68605a,a68606a,a68609a,a68612a,a68613a,a68614a,a68618a,a68619a,a68622a,a68625a,a68626a,a68627a,a68631a,a68632a,a68635a,a68638a,a68639a,a68640a,a68644a,a68645a,a68648a,a68651a,a68652a,a68653a,a68657a,a68658a,a68661a,a68664a,a68665a,a68666a,a68670a,a68671a,a68674a,a68677a,a68678a,a68679a,a68683a,a68684a,a68687a,a68690a,a68691a,a68692a,a68696a,a68697a,a68700a,a68703a,a68704a,a68705a,a68709a,a68710a,a68713a,a68716a,a68717a,a68718a,a68722a,a68723a,a68726a,a68729a,a68730a,a68731a,a68735a,a68736a,a68739a,a68742a,a68743a,a68744a,a68748a,a68749a,a68752a,a68755a,a68756a,a68757a,a68761a,a68762a,a68765a,a68768a,a68769a,a68770a,a68774a,a68775a,a68778a,a68781a,a68782a,a68783a,a68787a,a68788a,a68791a,a68794a,a68795a,a68796a,a68800a,a68801a,a68804a,a68807a,a68808a,a68809a,a68813a,a68814a,a68817a,a68820a,a68821a,a68822a,a68826a,a68827a,a68830a,a68833a,a68834a,a68835a,a68839a,a68840a,a68843a,a68846a,a68847a,a68848a,a68852a,a68853a,a68856a,a68859a,a68860a,a68861a,a68865a,a68866a,a68869a,a68872a,a68873a,a68874a,a68878a,a68879a,a68882a,a68885a,a68886a,a68887a,a68891a,a68892a,a68895a,a68898a,a68899a,a68900a,a68904a,a68905a,a68908a,a68911a,a68912a,a68913a,a68917a,a68918a,a68921a,a68924a,a68925a,a68926a,a68930a,a68931a,a68934a,a68937a,a68938a,a68939a,a68943a,a68944a,a68947a,a68950a,a68951a,a68952a,a68956a,a68957a,a68960a,a68963a,a68964a,a68965a,a68969a,a68970a,a68973a,a68976a,a68977a,a68978a,a68982a,a68983a,a68986a,a68989a,a68990a,a68991a,a68995a,a68996a,a68999a,a69002a,a69003a,a69004a,a69008a,a69009a,a69012a,a69015a,a69016a,a69017a,a69021a,a69022a,a69025a,a69028a,a69029a,a69030a,a69034a,a69035a,a69038a,a69041a,a69042a,a69043a,a69047a,a69048a,a69051a,a69054a,a69055a,a69056a,a69060a,a69061a,a69064a,a69067a,a69068a,a69069a,a69073a,a69074a,a69077a,a69080a,a69081a,a69082a,a69086a,a69087a,a69090a,a69093a,a69094a,a69095a,a69099a,a69100a,a69103a,a69106a,a69107a,a69108a,a69112a,a69113a,a69116a,a69119a,a69120a,a69121a,a69125a,a69126a,a69129a,a69132a,a69133a,a69134a,a69138a,a69139a,a69142a,a69145a,a69146a,a69147a,a69151a,a69152a,a69155a,a69158a,a69159a,a69160a,a69164a,a69165a,a69168a,a69171a,a69172a,a69173a,a69177a,a69178a,a69181a,a69184a,a69185a,a69186a,a69190a,a69191a,a69194a,a69197a,a69198a,a69199a,a69203a,a69204a,a69207a,a69210a,a69211a,a69212a,a69216a,a69217a,a69220a,a69223a,a69224a,a69225a,a69229a,a69230a,a69233a,a69236a,a69237a,a69238a,a69242a,a69243a,a69246a,a69249a,a69250a,a69251a,a69255a,a69256a,a69259a,a69262a,a69263a,a69264a,a69268a,a69269a,a69272a,a69275a,a69276a,a69277a,a69281a,a69282a,a69285a,a69288a,a69289a,a69290a,a69294a,a69295a,a69298a,a69301a,a69302a,a69303a,a69307a,a69308a,a69311a,a69314a,a69315a,a69316a,a69320a,a69321a,a69324a,a69327a,a69328a,a69329a,a69333a,a69334a,a69337a,a69340a,a69341a,a69342a,a69346a,a69347a,a69350a,a69353a,a69354a,a69355a,a69359a,a69360a,a69363a,a69366a,a69367a,a69368a,a69372a,a69373a,a69376a,a69379a,a69380a,a69381a,a69385a,a69386a,a69389a,a69392a,a69393a,a69394a,a69398a,a69399a,a69402a,a69405a,a69406a,a69407a,a69411a,a69412a,a69415a,a69418a,a69419a,a69420a,a69424a,a69425a,a69428a,a69431a,a69432a,a69433a,a69437a,a69438a,a69441a,a69444a,a69445a,a69446a,a69450a,a69451a,a69454a,a69457a,a69458a,a69459a,a69463a,a69464a,a69467a,a69470a,a69471a,a69472a,a69476a,a69477a,a69480a,a69483a,a69484a,a69485a,a69489a,a69490a,a69493a,a69496a,a69497a,a69498a,a69502a,a69503a,a69506a,a69509a,a69510a,a69511a,a69515a,a69516a,a69519a,a69522a,a69523a,a69524a,a69528a,a69529a,a69532a,a69535a,a69536a,a69537a,a69541a,a69542a,a69545a,a69548a,a69549a,a69550a,a69554a,a69555a,a69558a,a69561a,a69562a,a69563a,a69567a,a69568a,a69571a,a69574a,a69575a,a69576a,a69580a,a69581a,a69584a,a69587a,a69588a,a69589a,a69593a,a69594a,a69597a,a69600a,a69601a,a69602a,a69606a,a69607a,a69610a,a69613a,a69614a,a69615a,a69619a,a69620a,a69623a,a69626a,a69627a,a69628a,a69632a,a69633a,a69636a,a69639a,a69640a,a69641a,a69645a,a69646a,a69649a,a69652a,a69653a,a69654a,a69658a,a69659a,a69662a,a69665a,a69666a,a69667a,a69671a,a69672a,a69675a,a69678a,a69679a,a69680a,a69684a,a69685a,a69688a,a69691a,a69692a,a69693a,a69697a,a69698a,a69701a,a69704a,a69705a,a69706a,a69710a,a69711a,a69714a,a69717a,a69718a,a69719a,a69723a,a69724a,a69727a,a69730a,a69731a,a69732a,a69736a,a69737a,a69740a,a69743a,a69744a,a69745a,a69749a,a69750a,a69753a,a69756a,a69757a,a69758a,a69762a,a69763a,a69766a,a69769a,a69770a,a69771a,a69775a,a69776a,a69779a,a69782a,a69783a,a69784a,a69788a,a69789a,a69792a,a69795a,a69796a,a69797a,a69801a,a69802a,a69805a,a69808a,a69809a,a69810a,a69814a,a69815a,a69818a,a69821a,a69822a,a69823a,a69827a,a69828a,a69831a,a69834a,a69835a,a69836a,a69840a,a69841a,a69844a,a69847a,a69848a,a69849a,a69853a,a69854a,a69857a,a69860a,a69861a,a69862a,a69866a,a69867a,a69870a,a69873a,a69874a,a69875a,a69879a,a69880a,a69883a,a69886a,a69887a,a69888a,a69892a,a69893a,a69896a,a69899a,a69900a,a69901a,a69905a,a69906a,a69909a,a69912a,a69913a,a69914a,a69918a,a69919a,a69922a,a69925a,a69926a,a69927a,a69931a,a69932a,a69935a,a69938a,a69939a,a69940a,a69944a,a69945a,a69948a,a69951a,a69952a,a69953a,a69957a,a69958a,a69961a,a69964a,a69965a,a69966a,a69970a,a69971a,a69974a,a69977a,a69978a,a69979a,a69983a,a69984a,a69987a,a69990a,a69991a,a69992a,a69996a,a69997a,a70000a,a70003a,a70004a,a70005a,a70009a,a70010a,a70013a,a70016a,a70017a,a70018a,a70022a,a70023a,a70026a,a70029a,a70030a,a70031a,a70035a,a70036a,a70039a,a70042a,a70043a,a70044a,a70048a,a70049a,a70052a,a70055a,a70056a,a70057a,a70061a,a70062a,a70065a,a70068a,a70069a,a70070a,a70074a,a70075a,a70078a,a70081a,a70082a,a70083a,a70087a,a70088a,a70091a,a70094a,a70095a,a70096a,a70100a,a70101a,a70104a,a70107a,a70108a,a70109a,a70113a,a70114a,a70117a,a70120a,a70121a,a70122a,a70126a,a70127a,a70130a,a70133a,a70134a,a70135a,a70139a,a70140a,a70143a,a70146a,a70147a,a70148a,a70152a,a70153a,a70156a,a70159a,a70160a,a70161a,a70165a,a70166a,a70169a,a70172a,a70173a,a70174a,a70178a,a70179a,a70182a,a70185a,a70186a,a70187a,a70191a,a70192a,a70195a,a70198a,a70199a,a70200a,a70204a,a70205a,a70208a,a70211a,a70212a,a70213a,a70217a,a70218a,a70221a,a70224a,a70225a,a70226a,a70230a,a70231a,a70234a,a70237a,a70238a,a70239a,a70243a,a70244a,a70247a,a70250a,a70251a,a70252a,a70256a,a70257a,a70260a,a70263a,a70264a,a70265a,a70269a,a70270a,a70273a,a70276a,a70277a,a70278a,a70282a,a70283a,a70286a,a70289a,a70290a,a70291a,a70295a,a70296a,a70299a,a70302a,a70303a,a70304a,a70308a,a70309a,a70312a,a70315a,a70316a,a70317a,a70321a,a70322a,a70325a,a70328a,a70329a,a70330a,a70334a,a70335a,a70338a,a70341a,a70342a,a70343a,a70347a,a70348a,a70351a,a70354a,a70355a,a70356a,a70360a,a70361a,a70364a,a70367a,a70368a,a70369a,a70373a,a70374a,a70377a,a70380a,a70381a,a70382a,a70386a,a70387a,a70390a,a70393a,a70394a,a70395a,a70399a,a70400a,a70403a,a70406a,a70407a,a70408a,a70412a,a70413a,a70416a,a70419a,a70420a,a70421a,a70425a,a70426a,a70429a,a70432a,a70433a,a70434a,a70438a,a70439a,a70442a,a70445a,a70446a,a70447a,a70451a,a70452a,a70455a,a70458a,a70459a,a70460a,a70464a,a70465a,a70468a,a70471a,a70472a,a70473a,a70477a,a70478a,a70481a,a70484a,a70485a,a70486a,a70490a,a70491a,a70494a,a70497a,a70498a,a70499a,a70503a,a70504a,a70507a,a70510a,a70511a,a70512a,a70516a,a70517a,a70520a,a70523a,a70524a,a70525a,a70529a,a70530a,a70533a,a70536a,a70537a,a70538a,a70542a,a70543a,a70546a,a70549a,a70550a,a70551a,a70555a,a70556a,a70559a,a70562a,a70563a,a70564a,a70568a,a70569a,a70572a,a70575a,a70576a,a70577a,a70581a,a70582a,a70585a,a70588a,a70589a,a70590a,a70594a,a70595a,a70598a,a70601a,a70602a,a70603a,a70607a,a70608a,a70611a,a70614a,a70615a,a70616a,a70620a,a70621a,a70624a,a70627a,a70628a,a70629a,a70633a,a70634a,a70637a,a70640a,a70641a,a70642a,a70646a,a70647a,a70650a,a70653a,a70654a,a70655a,a70659a,a70660a,a70663a,a70666a,a70667a,a70668a,a70672a,a70673a,a70676a,a70679a,a70680a,a70681a,a70685a,a70686a,a70689a,a70692a,a70693a,a70694a,a70698a,a70699a,a70702a,a70705a,a70706a,a70707a,a70711a,a70712a,a70715a,a70718a,a70719a,a70720a,a70724a,a70725a,a70728a,a70731a,a70732a,a70733a,a70737a,a70738a,a70741a,a70744a,a70745a,a70746a,a70750a,a70751a,a70754a,a70757a,a70758a,a70759a,a70763a,a70764a,a70767a,a70770a,a70771a,a70772a,a70776a,a70777a,a70780a,a70783a,a70784a,a70785a,a70789a,a70790a,a70793a,a70796a,a70797a,a70798a,a70802a,a70803a,a70806a,a70809a,a70810a,a70811a,a70815a,a70816a,a70819a,a70822a,a70823a,a70824a,a70828a,a70829a,a70832a,a70835a,a70836a,a70837a,a70841a,a70842a,a70845a,a70848a,a70849a,a70850a,a70854a,a70855a,a70858a,a70861a,a70862a,a70863a,a70867a,a70868a,a70871a,a70874a,a70875a,a70876a,a70880a,a70881a,a70884a,a70887a,a70888a,a70889a,a70893a,a70894a,a70897a,a70900a,a70901a,a70902a,a70906a,a70907a,a70910a,a70913a,a70914a,a70915a,a70919a,a70920a,a70923a,a70926a,a70927a,a70928a,a70932a,a70933a,a70936a,a70939a,a70940a,a70941a,a70945a,a70946a,a70949a,a70952a,a70953a,a70954a,a70958a,a70959a,a70962a,a70965a,a70966a,a70967a,a70971a,a70972a,a70975a,a70978a,a70979a,a70980a,a70984a,a70985a,a70988a,a70991a,a70992a,a70993a,a70997a,a70998a,a71001a,a71004a,a71005a,a71006a,a71010a,a71011a,a71014a,a71017a,a71018a,a71019a,a71023a,a71024a,a71027a,a71030a,a71031a,a71032a,a71036a,a71037a,a71040a,a71043a,a71044a,a71045a,a71049a,a71050a,a71053a,a71056a,a71057a,a71058a,a71062a,a71063a,a71066a,a71069a,a71070a,a71071a,a71075a,a71076a,a71079a,a71082a,a71083a,a71084a,a71088a,a71089a,a71092a,a71095a,a71096a,a71097a,a71101a,a71102a,a71105a,a71108a,a71109a,a71110a,a71114a,a71115a,a71118a,a71121a,a71122a,a71123a,a71127a,a71128a,a71131a,a71134a,a71135a,a71136a,a71140a,a71141a,a71144a,a71147a,a71148a,a71149a,a71153a,a71154a,a71157a,a71160a,a71161a,a71162a,a71166a,a71167a,a71170a,a71173a,a71174a,a71175a,a71179a,a71180a,a71183a,a71186a,a71187a,a71188a,a71192a,a71193a,a71196a,a71199a,a71200a,a71201a,a71205a,a71206a,a71209a,a71212a,a71213a,a71214a,a71218a,a71219a,a71222a,a71225a,a71226a,a71227a,a71231a,a71232a,a71235a,a71238a,a71239a,a71240a,a71244a,a71245a,a71248a,a71251a,a71252a,a71253a,a71257a,a71258a,a71261a,a71264a,a71265a,a71266a,a71270a,a71271a,a71274a,a71277a,a71278a,a71279a,a71283a,a71284a,a71287a,a71290a,a71291a,a71292a,a71296a,a71297a,a71300a,a71303a,a71304a,a71305a,a71309a,a71310a,a71313a,a71316a,a71317a,a71318a,a71322a,a71323a,a71326a,a71329a,a71330a,a71331a,a71335a,a71336a,a71339a,a71342a,a71343a,a71344a,a71348a,a71349a,a71352a,a71355a,a71356a,a71357a,a71361a,a71362a,a71365a,a71368a,a71369a,a71370a,a71374a,a71375a,a71378a,a71381a,a71382a,a71383a,a71387a,a71388a,a71391a,a71394a,a71395a,a71396a,a71400a,a71401a,a71404a,a71407a,a71408a,a71409a,a71413a,a71414a,a71417a,a71420a,a71421a,a71422a,a71426a,a71427a,a71430a,a71433a,a71434a,a71435a,a71439a,a71440a,a71443a,a71446a,a71447a,a71448a,a71452a,a71453a,a71456a,a71459a,a71460a,a71461a,a71465a,a71466a,a71469a,a71472a,a71473a,a71474a,a71478a,a71479a,a71482a,a71485a,a71486a,a71487a,a71491a,a71492a,a71495a,a71498a,a71499a,a71500a,a71504a,a71505a,a71508a,a71511a,a71512a,a71513a,a71517a,a71518a,a71521a,a71524a,a71525a,a71526a,a71530a,a71531a,a71534a,a71537a,a71538a,a71539a,a71543a,a71544a,a71547a,a71550a,a71551a,a71552a,a71556a,a71557a,a71560a,a71563a,a71564a,a71565a,a71569a,a71570a,a71573a,a71576a,a71577a,a71578a,a71582a,a71583a,a71586a,a71589a,a71590a,a71591a,a71595a,a71596a,a71599a,a71602a,a71603a,a71604a,a71608a,a71609a,a71612a,a71615a,a71616a,a71617a,a71621a,a71622a,a71625a,a71628a,a71629a,a71630a,a71634a,a71635a,a71638a,a71641a,a71642a,a71643a,a71647a,a71648a,a71651a,a71654a,a71655a,a71656a,a71660a,a71661a,a71664a,a71667a,a71668a,a71669a,a71673a,a71674a,a71677a,a71680a,a71681a,a71682a,a71686a,a71687a,a71690a,a71693a,a71694a,a71695a,a71699a,a71700a,a71703a,a71706a,a71707a,a71708a,a71712a,a71713a,a71716a,a71719a,a71720a,a71721a,a71725a,a71726a,a71729a,a71732a,a71733a,a71734a,a71738a,a71739a,a71742a,a71745a,a71746a,a71747a,a71751a,a71752a,a71755a,a71758a,a71759a,a71760a,a71764a,a71765a,a71768a,a71771a,a71772a,a71773a,a71777a,a71778a,a71781a,a71784a,a71785a,a71786a,a71790a,a71791a,a71794a,a71797a,a71798a,a71799a,a71803a,a71804a,a71807a,a71810a,a71811a,a71812a,a71816a,a71817a,a71820a,a71823a,a71824a,a71825a,a71829a,a71830a,a71833a,a71836a,a71837a,a71838a,a71842a,a71843a,a71846a,a71849a,a71850a,a71851a,a71855a,a71856a,a71859a,a71862a,a71863a,a71864a,a71868a,a71869a,a71872a,a71875a,a71876a,a71877a,a71881a,a71882a,a71885a,a71888a,a71889a,a71890a,a71894a,a71895a,a71898a,a71901a,a71902a,a71903a,a71907a,a71908a,a71911a,a71914a,a71915a,a71916a,a71920a,a71921a,a71924a,a71927a,a71928a,a71929a,a71933a,a71934a,a71937a,a71940a,a71941a,a71942a,a71946a,a71947a,a71950a,a71953a,a71954a,a71955a,a71959a,a71960a,a71963a,a71966a,a71967a,a71968a,a71972a,a71973a,a71976a,a71979a,a71980a,a71981a,a71985a,a71986a,a71989a,a71992a,a71993a,a71994a,a71998a,a71999a,a72002a,a72005a,a72006a,a72007a,a72011a,a72012a,a72015a,a72018a,a72019a,a72020a,a72024a,a72025a,a72028a,a72031a,a72032a,a72033a,a72037a,a72038a,a72041a,a72044a,a72045a,a72046a,a72050a,a72051a,a72054a,a72057a,a72058a,a72059a,a72063a,a72064a,a72067a,a72070a,a72071a,a72072a,a72076a,a72077a,a72080a,a72083a,a72084a,a72085a,a72089a,a72090a,a72093a,a72096a,a72097a,a72098a,a72102a,a72103a,a72106a,a72109a,a72110a,a72111a,a72115a,a72116a,a72119a,a72122a,a72123a,a72124a,a72128a,a72129a,a72132a,a72135a,a72136a,a72137a,a72141a,a72142a,a72145a,a72148a,a72149a,a72150a,a72154a,a72155a,a72158a,a72161a,a72162a,a72163a,a72167a,a72168a,a72171a,a72174a,a72175a,a72176a,a72180a,a72181a,a72184a,a72187a,a72188a,a72189a,a72193a,a72194a,a72197a,a72200a,a72201a,a72202a,a72206a,a72207a,a72210a,a72213a,a72214a,a72215a,a72219a,a72220a,a72223a,a72226a,a72227a,a72228a,a72232a,a72233a,a72236a,a72239a,a72240a,a72241a,a72245a,a72246a,a72249a,a72252a,a72253a,a72254a,a72258a,a72259a,a72262a,a72265a,a72266a,a72267a,a72271a,a72272a,a72275a,a72278a,a72279a,a72280a,a72284a,a72285a,a72288a,a72291a,a72292a,a72293a,a72297a,a72298a,a72301a,a72304a,a72305a,a72306a,a72310a,a72311a,a72314a,a72317a,a72318a,a72319a,a72323a,a72324a,a72327a,a72330a,a72331a,a72332a,a72336a,a72337a,a72340a,a72343a,a72344a,a72345a,a72349a,a72350a,a72353a,a72356a,a72357a,a72358a,a72362a,a72363a,a72366a,a72369a,a72370a,a72371a,a72375a,a72376a,a72379a,a72382a,a72383a,a72384a,a72388a,a72389a,a72392a,a72395a,a72396a,a72397a,a72401a,a72402a,a72405a,a72408a,a72409a,a72410a,a72414a,a72415a,a72418a,a72421a,a72422a,a72423a,a72427a,a72428a,a72431a,a72434a,a72435a,a72436a,a72440a,a72441a,a72444a,a72447a,a72448a,a72449a,a72453a,a72454a,a72457a,a72460a,a72461a,a72462a,a72466a,a72467a,a72470a,a72473a,a72474a,a72475a,a72479a,a72480a,a72483a,a72486a,a72487a,a72488a,a72492a,a72493a,a72496a,a72499a,a72500a,a72501a,a72505a,a72506a,a72509a,a72512a,a72513a,a72514a,a72518a,a72519a,a72522a,a72525a,a72526a,a72527a,a72531a,a72532a,a72535a,a72538a,a72539a,a72540a,a72544a,a72545a,a72548a,a72551a,a72552a,a72553a,a72557a,a72558a,a72561a,a72564a,a72565a,a72566a,a72570a,a72571a,a72574a,a72577a,a72578a,a72579a,a72583a,a72584a,a72587a,a72590a,a72591a,a72592a,a72596a,a72597a,a72600a,a72603a,a72604a,a72605a,a72609a,a72610a,a72613a,a72616a,a72617a,a72618a,a72622a,a72623a,a72626a,a72629a,a72630a,a72631a,a72635a,a72636a,a72639a,a72642a,a72643a,a72644a,a72648a,a72649a,a72652a,a72655a,a72656a,a72657a,a72661a,a72662a,a72665a,a72668a,a72669a,a72670a,a72674a,a72675a,a72678a,a72681a,a72682a,a72683a,a72687a,a72688a,a72691a,a72694a,a72695a,a72696a,a72700a,a72701a,a72704a,a72707a,a72708a,a72709a,a72713a,a72714a,a72717a,a72720a,a72721a,a72722a,a72726a,a72727a,a72730a,a72733a,a72734a,a72735a,a72739a,a72740a,a72743a,a72746a,a72747a,a72748a,a72752a,a72753a,a72756a,a72759a,a72760a,a72761a,a72765a,a72766a,a72769a,a72772a,a72773a,a72774a,a72778a,a72779a,a72782a,a72785a,a72786a,a72787a,a72791a,a72792a,a72795a,a72798a,a72799a,a72800a,a72804a,a72805a,a72808a,a72811a,a72812a,a72813a,a72817a,a72818a,a72821a,a72824a,a72825a,a72826a,a72830a,a72831a,a72834a,a72837a,a72838a,a72839a,a72843a,a72844a,a72847a,a72850a,a72851a,a72852a,a72856a,a72857a,a72860a,a72863a,a72864a,a72865a,a72869a,a72870a,a72873a,a72876a,a72877a,a72878a,a72882a,a72883a,a72886a,a72889a,a72890a,a72891a,a72895a,a72896a,a72899a,a72902a,a72903a,a72904a,a72908a,a72909a,a72912a,a72915a,a72916a,a72917a,a72921a,a72922a,a72925a,a72928a,a72929a,a72930a,a72934a,a72935a,a72938a,a72941a,a72942a,a72943a,a72947a,a72948a,a72951a,a72954a,a72955a,a72956a,a72960a,a72961a,a72964a,a72967a,a72968a,a72969a,a72973a,a72974a,a72977a,a72980a,a72981a,a72982a,a72986a,a72987a,a72990a,a72993a,a72994a,a72995a,a72999a,a73000a,a73003a,a73006a,a73007a,a73008a,a73012a,a73013a,a73016a,a73019a,a73020a,a73021a,a73025a,a73026a,a73029a,a73032a,a73033a,a73034a,a73038a,a73039a,a73042a,a73045a,a73046a,a73047a,a73051a,a73052a,a73055a,a73058a,a73059a,a73060a,a73064a,a73065a,a73068a,a73071a,a73072a,a73073a,a73077a,a73078a,a73081a,a73084a,a73085a,a73086a,a73090a,a73091a,a73094a,a73097a,a73098a,a73099a,a73103a,a73104a,a73107a,a73110a,a73111a,a73112a,a73116a,a73117a,a73120a,a73123a,a73124a,a73125a,a73129a,a73130a,a73133a,a73136a,a73137a,a73138a,a73142a,a73143a,a73146a,a73149a,a73150a,a73151a,a73155a,a73156a,a73159a,a73162a,a73163a,a73164a,a73168a,a73169a,a73172a,a73175a,a73176a,a73177a,a73181a,a73182a,a73185a,a73188a,a73189a,a73190a,a73194a,a73195a,a73198a,a73201a,a73202a,a73203a,a73207a,a73208a,a73211a,a73214a,a73215a,a73216a,a73220a,a73221a,a73224a,a73227a,a73228a,a73229a,a73233a,a73234a,a73237a,a73240a,a73241a,a73242a,a73246a,a73247a,a73250a,a73253a,a73254a,a73255a,a73259a,a73260a,a73263a,a73266a,a73267a,a73268a,a73272a,a73273a,a73276a,a73279a,a73280a,a73281a,a73285a,a73286a,a73289a,a73292a,a73293a,a73294a,a73298a,a73299a,a73302a,a73305a,a73306a,a73307a,a73311a,a73312a,a73315a,a73318a,a73319a,a73320a,a73324a,a73325a,a73328a,a73331a,a73332a,a73333a,a73337a,a73338a,a73341a,a73344a,a73345a,a73346a,a73350a,a73351a,a73354a,a73357a,a73358a,a73359a,a73363a,a73364a,a73367a,a73370a,a73371a,a73372a,a73376a,a73377a,a73380a,a73383a,a73384a,a73385a,a73389a,a73390a,a73393a,a73396a,a73397a,a73398a,a73402a,a73403a,a73406a,a73409a,a73410a,a73411a,a73415a,a73416a,a73419a,a73422a,a73423a,a73424a,a73428a,a73429a,a73432a,a73435a,a73436a,a73437a,a73441a,a73442a,a73445a,a73448a,a73449a,a73450a,a73454a,a73455a,a73458a,a73461a,a73462a,a73463a,a73467a,a73468a,a73471a,a73474a,a73475a,a73476a,a73480a,a73481a,a73484a,a73487a,a73488a,a73489a,a73493a,a73494a,a73497a,a73500a,a73501a,a73502a,a73506a,a73507a,a73510a,a73513a,a73514a,a73515a,a73519a,a73520a,a73523a,a73526a,a73527a,a73528a,a73532a,a73533a,a73536a,a73539a,a73540a,a73541a,a73545a,a73546a,a73549a,a73552a,a73553a,a73554a,a73558a,a73559a,a73562a,a73565a,a73566a,a73567a,a73571a,a73572a,a73575a,a73578a,a73579a,a73580a,a73584a,a73585a,a73588a,a73591a,a73592a,a73593a,a73597a,a73598a,a73601a,a73604a,a73605a,a73606a,a73610a,a73611a,a73614a,a73617a,a73618a,a73619a,a73623a,a73624a,a73627a,a73630a,a73631a,a73632a,a73636a,a73637a,a73640a,a73643a,a73644a,a73645a,a73649a,a73650a,a73653a,a73656a,a73657a,a73658a,a73662a,a73663a,a73666a,a73669a,a73670a,a73671a,a73675a,a73676a,a73679a,a73682a,a73683a,a73684a,a73688a,a73689a,a73692a,a73695a,a73696a,a73697a,a73701a,a73702a,a73705a,a73708a,a73709a,a73710a,a73714a,a73715a,a73718a,a73721a,a73722a,a73723a,a73727a,a73728a,a73731a,a73734a,a73735a,a73736a,a73740a,a73741a,a73744a,a73747a,a73748a,a73749a,a73753a,a73754a,a73757a,a73760a,a73761a,a73762a,a73766a,a73767a,a73770a,a73773a,a73774a,a73775a,a73779a,a73780a,a73783a,a73786a,a73787a,a73788a,a73792a,a73793a,a73796a,a73799a,a73800a,a73801a,a73805a,a73806a,a73809a,a73812a,a73813a,a73814a,a73818a,a73819a,a73822a,a73825a,a73826a,a73827a,a73831a,a73832a,a73835a,a73838a,a73839a,a73840a,a73844a,a73845a,a73848a,a73851a,a73852a,a73853a,a73857a,a73858a,a73861a,a73864a,a73865a,a73866a,a73870a,a73871a,a73874a,a73877a,a73878a,a73879a,a73883a,a73884a,a73887a,a73890a,a73891a,a73892a,a73896a,a73897a,a73900a,a73903a,a73904a,a73905a,a73909a,a73910a,a73913a,a73916a,a73917a,a73918a,a73922a,a73923a,a73926a,a73929a,a73930a,a73931a,a73935a,a73936a,a73939a,a73942a,a73943a,a73944a,a73948a,a73949a,a73952a,a73955a,a73956a,a73957a,a73961a,a73962a,a73965a,a73968a,a73969a,a73970a,a73974a,a73975a,a73978a,a73981a,a73982a,a73983a,a73987a,a73988a,a73991a,a73994a,a73995a,a73996a,a74000a,a74001a,a74004a,a74007a,a74008a,a74009a,a74013a,a74014a,a74017a,a74020a,a74021a,a74022a,a74026a,a74027a,a74030a,a74033a,a74034a,a74035a,a74039a,a74040a,a74043a,a74046a,a74047a,a74048a,a74052a,a74053a,a74056a,a74059a,a74060a,a74061a,a74065a,a74066a,a74069a,a74072a,a74073a,a74074a,a74078a,a74079a,a74082a,a74085a,a74086a,a74087a,a74091a,a74092a,a74095a,a74098a,a74099a,a74100a,a74104a,a74105a,a74108a,a74111a,a74112a,a74113a,a74117a,a74118a,a74121a,a74124a,a74125a,a74126a,a74130a,a74131a,a74134a,a74137a,a74138a,a74139a,a74143a,a74144a,a74147a,a74150a,a74151a,a74152a,a74156a,a74157a,a74160a,a74163a,a74164a,a74165a,a74169a,a74170a,a74173a,a74176a,a74177a,a74178a,a74182a,a74183a,a74186a,a74189a,a74190a,a74191a,a74195a,a74196a,a74199a,a74202a,a74203a,a74204a,a74208a,a74209a,a74212a,a74215a,a74216a,a74217a,a74221a,a74222a,a74225a,a74228a,a74229a,a74230a,a74234a,a74235a,a74238a,a74241a,a74242a,a74243a,a74247a,a74248a,a74251a,a74254a,a74255a,a74256a,a74260a,a74261a,a74264a,a74267a,a74268a,a74269a,a74273a,a74274a,a74277a,a74280a,a74281a,a74282a,a74286a,a74287a,a74290a,a74293a,a74294a,a74295a,a74299a,a74300a,a74303a,a74306a,a74307a,a74308a,a74312a,a74313a,a74316a,a74319a,a74320a,a74321a,a74325a,a74326a,a74329a,a74332a,a74333a,a74334a,a74338a,a74339a,a74342a,a74345a,a74346a,a74347a,a74351a,a74352a,a74355a,a74358a,a74359a,a74360a,a74364a,a74365a,a74368a,a74371a,a74372a,a74373a,a74377a,a74378a,a74381a,a74384a,a74385a,a74386a,a74390a,a74391a,a74394a,a74397a,a74398a,a74399a,a74403a,a74404a,a74407a,a74410a,a74411a,a74412a,a74416a,a74417a,a74420a,a74423a,a74424a,a74425a,a74429a,a74430a,a74433a,a74436a,a74437a,a74438a,a74442a,a74443a,a74446a,a74449a,a74450a,a74451a,a74455a,a74456a,a74459a,a74462a,a74463a,a74464a,a74468a,a74469a,a74472a,a74475a,a74476a,a74477a,a74481a,a74482a,a74485a,a74488a,a74489a,a74490a,a74494a,a74495a,a74498a,a74501a,a74502a,a74503a,a74507a,a74508a,a74511a,a74514a,a74515a,a74516a,a74520a,a74521a,a74524a,a74527a,a74528a,a74529a,a74533a,a74534a,a74537a,a74540a,a74541a,a74542a,a74546a,a74547a,a74550a,a74553a,a74554a,a74555a,a74559a,a74560a,a74563a,a74566a,a74567a,a74568a,a74572a,a74573a,a74576a,a74579a,a74580a,a74581a,a74585a,a74586a,a74589a,a74592a,a74593a,a74594a,a74598a,a74599a,a74602a,a74605a,a74606a,a74607a,a74611a,a74612a,a74615a,a74618a,a74619a,a74620a,a74624a,a74625a,a74628a,a74631a,a74632a,a74633a,a74637a,a74638a,a74641a,a74644a,a74645a,a74646a,a74650a,a74651a,a74654a,a74657a,a74658a,a74659a,a74663a,a74664a,a74667a,a74670a,a74671a,a74672a,a74676a,a74677a,a74680a,a74683a,a74684a,a74685a,a74689a,a74690a,a74693a,a74696a,a74697a,a74698a,a74702a,a74703a,a74706a,a74709a,a74710a,a74711a,a74715a,a74716a,a74719a,a74722a,a74723a,a74724a,a74728a,a74729a,a74732a,a74735a,a74736a,a74737a,a74741a,a74742a,a74745a,a74748a,a74749a,a74750a,a74754a,a74755a,a74758a,a74761a,a74762a,a74763a,a74767a,a74768a,a74771a,a74774a,a74775a,a74776a,a74780a,a74781a,a74784a,a74787a,a74788a,a74789a,a74793a,a74794a,a74797a,a74800a,a74801a,a74802a,a74806a,a74807a,a74810a,a74813a,a74814a,a74815a,a74819a,a74820a,a74823a,a74826a,a74827a,a74828a,a74832a,a74833a,a74836a,a74839a,a74840a,a74841a,a74845a,a74846a,a74849a,a74852a,a74853a,a74854a,a74858a,a74859a,a74862a,a74865a,a74866a,a74867a,a74871a,a74872a,a74875a,a74878a,a74879a,a74880a,a74884a,a74885a,a74888a,a74891a,a74892a,a74893a,a74897a,a74898a,a74901a,a74904a,a74905a,a74906a,a74910a,a74911a,a74914a,a74917a,a74918a,a74919a,a74923a,a74924a,a74927a,a74930a,a74931a,a74932a,a74936a,a74937a,a74940a,a74943a,a74944a,a74945a,a74949a,a74950a,a74953a,a74956a,a74957a,a74958a,a74962a,a74963a,a74966a,a74969a,a74970a,a74971a,a74975a,a74976a,a74979a,a74982a,a74983a,a74984a,a74988a,a74989a,a74992a,a74995a,a74996a,a74997a,a75001a,a75002a,a75005a,a75008a,a75009a,a75010a,a75014a,a75015a,a75018a,a75021a,a75022a,a75023a,a75027a,a75028a,a75031a,a75034a,a75035a,a75036a,a75040a,a75041a,a75044a,a75047a,a75048a,a75049a,a75053a,a75054a,a75057a,a75060a,a75061a,a75062a,a75066a,a75067a,a75070a,a75073a,a75074a,a75075a,a75079a,a75080a,a75083a,a75086a,a75087a,a75088a,a75092a,a75093a,a75096a,a75099a,a75100a,a75101a,a75105a,a75106a,a75109a,a75112a,a75113a,a75114a,a75118a,a75119a,a75122a,a75125a,a75126a,a75127a,a75131a,a75132a,a75135a,a75138a,a75139a,a75140a,a75144a,a75145a,a75148a,a75151a,a75152a,a75153a,a75157a,a75158a,a75161a,a75164a,a75165a,a75166a,a75170a,a75171a,a75174a,a75177a,a75178a,a75179a,a75183a,a75184a,a75187a,a75190a,a75191a,a75192a,a75196a,a75197a,a75200a,a75203a,a75204a,a75205a,a75209a,a75210a,a75213a,a75216a,a75217a,a75218a,a75222a,a75223a,a75226a,a75229a,a75230a,a75231a,a75235a,a75236a,a75239a,a75242a,a75243a,a75244a,a75248a,a75249a,a75252a,a75255a,a75256a,a75257a,a75261a,a75262a,a75265a,a75268a,a75269a,a75270a,a75274a,a75275a,a75278a,a75281a,a75282a,a75283a,a75287a,a75288a,a75291a,a75294a,a75295a,a75296a,a75300a,a75301a,a75304a,a75307a,a75308a,a75309a,a75313a,a75314a,a75317a,a75320a,a75321a,a75322a,a75326a,a75327a,a75330a,a75333a,a75334a,a75335a,a75339a,a75340a,a75343a,a75346a,a75347a,a75348a,a75352a,a75353a,a75356a,a75359a,a75360a,a75361a,a75365a,a75366a,a75369a,a75372a,a75373a,a75374a,a75378a,a75379a,a75382a,a75385a,a75386a,a75387a,a75391a,a75392a,a75395a,a75398a,a75399a,a75400a,a75404a,a75405a,a75408a,a75411a,a75412a,a75413a,a75417a,a75418a,a75421a,a75424a,a75425a,a75426a,a75430a,a75431a,a75434a,a75437a,a75438a,a75439a,a75443a,a75444a,a75447a,a75450a,a75451a,a75452a,a75456a,a75457a,a75460a,a75463a,a75464a,a75465a,a75469a,a75470a,a75473a,a75476a,a75477a,a75478a,a75482a,a75483a,a75486a,a75489a,a75490a,a75491a,a75495a,a75496a,a75499a,a75502a,a75503a,a75504a,a75508a,a75509a,a75512a,a75515a,a75516a,a75517a,a75521a,a75522a,a75525a,a75528a,a75529a,a75530a,a75534a,a75535a,a75538a,a75541a,a75542a,a75543a,a75547a,a75548a,a75551a,a75554a,a75555a,a75556a,a75560a,a75561a,a75564a,a75567a,a75568a,a75569a,a75573a,a75574a,a75577a,a75580a,a75581a,a75582a,a75586a,a75587a,a75590a,a75593a,a75594a,a75595a,a75599a,a75600a,a75603a,a75606a,a75607a,a75608a,a75612a,a75613a,a75616a,a75619a,a75620a,a75621a,a75625a,a75626a,a75629a,a75632a,a75633a,a75634a,a75638a,a75639a,a75642a,a75645a,a75646a,a75647a,a75651a,a75652a,a75655a,a75658a,a75659a,a75660a,a75664a,a75665a,a75668a,a75671a,a75672a,a75673a,a75677a,a75678a,a75681a,a75684a,a75685a,a75686a,a75690a,a75691a,a75694a,a75697a,a75698a,a75699a,a75703a,a75704a,a75707a,a75710a,a75711a,a75712a,a75716a,a75717a,a75720a,a75723a,a75724a,a75725a,a75729a,a75730a,a75733a,a75736a,a75737a,a75738a,a75742a,a75743a,a75746a,a75749a,a75750a,a75751a,a75755a,a75756a,a75759a,a75762a,a75763a,a75764a,a75768a,a75769a,a75772a,a75775a,a75776a,a75777a,a75781a,a75782a,a75785a,a75788a,a75789a,a75790a,a75794a,a75795a,a75798a,a75801a,a75802a,a75803a,a75807a,a75808a,a75811a,a75814a,a75815a,a75816a,a75820a,a75821a,a75824a,a75827a,a75828a,a75829a,a75833a,a75834a,a75837a,a75840a,a75841a,a75842a,a75846a,a75847a,a75850a,a75853a,a75854a,a75855a,a75859a,a75860a,a75863a,a75866a,a75867a,a75868a,a75872a,a75873a,a75876a,a75879a,a75880a,a75881a,a75885a,a75886a,a75889a,a75892a,a75893a,a75894a,a75898a,a75899a,a75902a,a75905a,a75906a,a75907a,a75911a,a75912a,a75915a,a75918a,a75919a,a75920a,a75924a,a75925a,a75928a,a75931a,a75932a,a75933a,a75937a,a75938a,a75941a,a75944a,a75945a,a75946a,a75950a,a75951a,a75954a,a75957a,a75958a,a75959a,a75963a,a75964a,a75967a,a75970a,a75971a,a75972a,a75976a,a75977a,a75980a,a75983a,a75984a,a75985a,a75989a,a75990a,a75993a,a75996a,a75997a,a75998a,a76002a,a76003a,a76006a,a76009a,a76010a,a76011a,a76015a,a76016a,a76019a,a76022a,a76023a,a76024a,a76028a,a76029a,a76032a,a76035a,a76036a,a76037a,a76041a,a76042a,a76045a,a76048a,a76049a,a76050a,a76054a,a76055a,a76058a,a76061a,a76062a,a76063a,a76067a,a76068a,a76071a,a76074a,a76075a,a76076a,a76080a,a76081a,a76084a,a76087a,a76088a,a76089a,a76093a,a76094a,a76097a,a76100a,a76101a,a76102a,a76106a,a76107a,a76110a,a76113a,a76114a,a76115a,a76119a,a76120a,a76123a,a76126a,a76127a,a76128a,a76132a,a76133a,a76136a,a76139a,a76140a,a76141a,a76145a,a76146a,a76149a,a76152a,a76153a,a76154a,a76158a,a76159a,a76162a,a76165a,a76166a,a76167a,a76171a,a76172a,a76175a,a76178a,a76179a,a76180a,a76184a,a76185a,a76188a,a76191a,a76192a,a76193a,a76197a,a76198a,a76201a,a76204a,a76205a,a76206a,a76210a,a76211a,a76214a,a76217a,a76218a,a76219a,a76223a,a76224a,a76227a,a76230a,a76231a,a76232a,a76236a,a76237a,a76240a,a76243a,a76244a,a76245a,a76249a,a76250a,a76253a,a76256a,a76257a,a76258a,a76262a,a76263a,a76266a,a76269a,a76270a,a76271a,a76275a,a76276a,a76279a,a76282a,a76283a,a76284a,a76288a,a76289a,a76292a,a76295a,a76296a,a76297a,a76301a,a76302a,a76305a,a76308a,a76309a,a76310a,a76314a,a76315a,a76318a,a76321a,a76322a,a76323a,a76327a,a76328a,a76331a,a76334a,a76335a,a76336a,a76340a,a76341a,a76344a,a76347a,a76348a,a76349a,a76353a,a76354a,a76357a,a76360a,a76361a,a76362a,a76366a,a76367a,a76370a,a76373a,a76374a,a76375a,a76379a,a76380a,a76383a,a76386a,a76387a,a76388a,a76392a,a76393a,a76396a,a76399a,a76400a,a76401a,a76405a,a76406a,a76409a,a76412a,a76413a,a76414a,a76418a,a76419a,a76422a,a76425a,a76426a,a76427a,a76431a,a76432a,a76435a,a76438a,a76439a,a76440a,a76444a,a76445a,a76448a,a76451a,a76452a,a76453a,a76457a,a76458a,a76461a,a76464a,a76465a,a76466a,a76470a,a76471a,a76474a,a76477a,a76478a,a76479a,a76483a,a76484a,a76487a,a76490a,a76491a,a76492a,a76496a,a76497a,a76500a,a76503a,a76504a,a76505a,a76509a,a76510a,a76513a,a76516a,a76517a,a76518a,a76522a,a76523a,a76526a,a76529a,a76530a,a76531a,a76535a,a76536a,a76539a,a76542a,a76543a,a76544a,a76548a,a76549a,a76552a,a76555a,a76556a,a76557a,a76561a,a76562a,a76565a,a76568a,a76569a,a76570a,a76574a,a76575a,a76578a,a76581a,a76582a,a76583a,a76587a,a76588a,a76591a,a76594a,a76595a,a76596a,a76600a,a76601a,a76604a,a76607a,a76608a,a76609a,a76613a,a76614a,a76617a,a76620a,a76621a,a76622a,a76626a,a76627a,a76630a,a76633a,a76634a,a76635a,a76639a,a76640a,a76643a,a76646a,a76647a,a76648a,a76652a,a76653a,a76656a,a76659a,a76660a,a76661a,a76665a,a76666a,a76669a,a76672a,a76673a,a76674a,a76678a,a76679a,a76682a,a76685a,a76686a,a76687a,a76691a,a76692a,a76695a,a76698a,a76699a,a76700a,a76704a,a76705a,a76708a,a76711a,a76712a,a76713a,a76717a,a76718a,a76721a,a76724a,a76725a,a76726a,a76730a,a76731a,a76734a,a76737a,a76738a,a76739a,a76743a,a76744a,a76747a,a76750a,a76751a,a76752a,a76756a,a76757a,a76760a,a76763a,a76764a,a76765a,a76769a,a76770a,a76773a,a76776a,a76777a,a76778a,a76782a,a76783a,a76786a,a76789a,a76790a,a76791a,a76795a,a76796a,a76799a,a76802a,a76803a,a76804a,a76808a,a76809a,a76812a,a76815a,a76816a,a76817a,a76821a,a76822a,a76825a,a76828a,a76829a,a76830a,a76834a,a76835a,a76838a,a76841a,a76842a,a76843a,a76847a,a76848a,a76851a,a76854a,a76855a,a76856a,a76860a,a76861a,a76864a,a76867a,a76868a,a76869a,a76873a,a76874a,a76877a,a76880a,a76881a,a76882a,a76886a,a76887a,a76890a,a76893a,a76894a,a76895a,a76899a,a76900a,a76903a,a76906a,a76907a,a76908a,a76912a,a76913a,a76916a,a76919a,a76920a,a76921a,a76925a,a76926a,a76929a,a76932a,a76933a,a76934a,a76938a,a76939a,a76942a,a76945a,a76946a,a76947a,a76951a,a76952a,a76955a,a76958a,a76959a,a76960a,a76964a,a76965a,a76968a,a76971a,a76972a,a76973a,a76977a,a76978a,a76981a,a76984a,a76985a,a76986a,a76990a,a76991a,a76994a,a76997a,a76998a,a76999a,a77003a,a77004a,a77007a,a77010a,a77011a,a77012a,a77016a,a77017a,a77020a,a77023a,a77024a,a77025a,a77029a,a77030a,a77033a,a77036a,a77037a,a77038a,a77042a,a77043a,a77046a,a77049a,a77050a,a77051a,a77055a,a77056a,a77059a,a77062a,a77063a,a77064a,a77068a,a77069a,a77072a,a77075a,a77076a,a77077a,a77081a,a77082a,a77085a,a77088a,a77089a,a77090a,a77094a,a77095a,a77098a,a77101a,a77102a,a77103a,a77107a,a77108a,a77111a,a77114a,a77115a,a77116a,a77120a,a77121a,a77124a,a77127a,a77128a,a77129a,a77133a,a77134a,a77137a,a77140a,a77141a,a77142a,a77146a,a77147a,a77150a,a77153a,a77154a,a77155a,a77159a,a77160a,a77163a,a77166a,a77167a,a77168a,a77172a,a77173a,a77176a,a77179a,a77180a,a77181a,a77185a,a77186a,a77189a,a77192a,a77193a,a77194a,a77198a,a77199a,a77202a,a77205a,a77206a,a77207a,a77211a,a77212a,a77215a,a77218a,a77219a,a77220a,a77224a,a77225a,a77228a,a77231a,a77232a,a77233a,a77237a,a77238a,a77241a,a77244a,a77245a,a77246a,a77250a,a77251a,a77254a,a77257a,a77258a,a77259a,a77263a,a77264a,a77267a,a77270a,a77271a,a77272a,a77276a,a77277a,a77280a,a77283a,a77284a,a77285a,a77289a,a77290a,a77293a,a77296a,a77297a,a77298a,a77302a,a77303a,a77306a,a77309a,a77310a,a77311a,a77315a,a77316a,a77319a,a77322a,a77323a,a77324a,a77328a,a77329a,a77332a,a77335a,a77336a,a77337a,a77341a,a77342a,a77345a,a77348a,a77349a,a77350a,a77354a,a77355a,a77358a,a77361a,a77362a,a77363a,a77367a,a77368a,a77371a,a77374a,a77375a,a77376a,a77380a,a77381a,a77384a,a77387a,a77388a,a77389a,a77393a,a77394a,a77397a,a77400a,a77401a,a77402a,a77406a,a77407a,a77410a,a77413a,a77414a,a77415a,a77419a,a77420a,a77423a,a77426a,a77427a,a77428a,a77432a,a77433a,a77436a,a77439a,a77440a,a77441a,a77445a,a77446a,a77449a,a77452a,a77453a,a77454a,a77458a,a77459a,a77462a,a77465a,a77466a,a77467a,a77471a,a77472a,a77475a,a77478a,a77479a,a77480a,a77484a,a77485a,a77488a,a77491a,a77492a,a77493a,a77497a,a77498a,a77501a,a77504a,a77505a,a77506a,a77510a,a77511a,a77514a,a77517a,a77518a,a77519a,a77523a,a77524a,a77527a,a77530a,a77531a,a77532a,a77536a,a77537a,a77540a,a77543a,a77544a,a77545a,a77549a,a77550a,a77553a,a77556a,a77557a,a77558a,a77562a,a77563a,a77566a,a77569a,a77570a,a77571a,a77575a,a77576a,a77579a,a77582a,a77583a,a77584a,a77588a,a77589a,a77592a,a77595a,a77596a,a77597a,a77601a,a77602a,a77605a,a77608a,a77609a,a77610a,a77614a,a77615a,a77618a,a77621a,a77622a,a77623a,a77627a,a77628a,a77631a,a77634a,a77635a,a77636a,a77640a,a77641a,a77644a,a77647a,a77648a,a77649a,a77652a,a77655a,a77656a,a77659a,a77662a,a77663a,a77664a,a77668a,a77669a,a77672a,a77675a,a77676a,a77677a,a77680a,a77683a,a77684a,a77687a,a77690a,a77691a,a77692a,a77696a,a77697a,a77700a,a77703a,a77704a,a77705a,a77708a,a77711a,a77712a,a77715a,a77718a,a77719a,a77720a,a77724a,a77725a,a77728a,a77731a,a77732a,a77733a,a77736a,a77739a,a77740a,a77743a,a77746a,a77747a,a77748a,a77752a,a77753a,a77756a,a77759a,a77760a,a77761a,a77764a,a77767a,a77768a,a77771a,a77774a,a77775a,a77776a,a77780a,a77781a,a77784a,a77787a,a77788a,a77789a,a77792a,a77795a,a77796a,a77799a,a77802a,a77803a,a77804a,a77808a,a77809a,a77812a,a77815a,a77816a,a77817a,a77820a,a77823a,a77824a,a77827a,a77830a,a77831a,a77832a,a77836a,a77837a,a77840a,a77843a,a77844a,a77845a,a77848a,a77851a,a77852a,a77855a,a77858a,a77859a,a77860a,a77864a,a77865a,a77868a,a77871a,a77872a,a77873a,a77876a,a77879a,a77880a,a77883a,a77886a,a77887a,a77888a,a77892a,a77893a,a77896a,a77899a,a77900a,a77901a,a77904a,a77907a,a77908a,a77911a,a77914a,a77915a,a77916a,a77920a,a77921a,a77924a,a77927a,a77928a,a77929a,a77932a,a77935a,a77936a,a77939a,a77942a,a77943a,a77944a,a77948a,a77949a,a77952a,a77955a,a77956a,a77957a,a77960a,a77963a,a77964a,a77967a,a77970a,a77971a,a77972a,a77976a,a77977a,a77980a,a77983a,a77984a,a77985a,a77988a,a77991a,a77992a,a77995a,a77998a,a77999a,a78000a,a78004a,a78005a,a78008a,a78011a,a78012a,a78013a,a78016a,a78019a,a78020a,a78023a,a78026a,a78027a,a78028a,a78032a,a78033a,a78036a,a78039a,a78040a,a78041a,a78044a,a78047a,a78048a,a78051a,a78054a,a78055a,a78056a,a78060a,a78061a,a78064a,a78067a,a78068a,a78069a,a78072a,a78075a,a78076a,a78079a,a78082a,a78083a,a78084a,a78088a,a78089a,a78092a,a78095a,a78096a,a78097a,a78100a,a78103a,a78104a,a78107a,a78110a,a78111a,a78112a,a78116a,a78117a,a78120a,a78123a,a78124a,a78125a,a78128a,a78131a,a78132a,a78135a,a78138a,a78139a,a78140a,a78144a,a78145a,a78148a,a78151a,a78152a,a78153a,a78156a,a78159a,a78160a,a78163a,a78166a,a78167a,a78168a,a78172a,a78173a,a78176a,a78179a,a78180a,a78181a,a78184a,a78187a,a78188a,a78191a,a78194a,a78195a,a78196a,a78200a,a78201a,a78204a,a78207a,a78208a,a78209a,a78212a,a78215a,a78216a,a78219a,a78222a,a78223a,a78224a,a78228a,a78229a,a78232a,a78235a,a78236a,a78237a,a78240a,a78243a,a78244a,a78247a,a78250a,a78251a,a78252a,a78256a,a78257a,a78260a,a78263a,a78264a,a78265a,a78268a,a78271a,a78272a,a78275a,a78278a,a78279a,a78280a,a78284a,a78285a,a78288a,a78291a,a78292a,a78293a,a78296a,a78299a,a78300a,a78303a,a78306a,a78307a,a78308a,a78312a,a78313a,a78316a,a78319a,a78320a,a78321a,a78324a,a78327a,a78328a,a78331a,a78334a,a78335a,a78336a,a78340a,a78341a,a78344a,a78347a,a78348a,a78349a,a78352a,a78355a,a78356a,a78359a,a78362a,a78363a,a78364a,a78368a,a78369a,a78372a,a78375a,a78376a,a78377a,a78380a,a78383a,a78384a,a78387a,a78390a,a78391a,a78392a,a78396a,a78397a,a78400a,a78403a,a78404a,a78405a,a78408a,a78411a,a78412a,a78415a,a78418a,a78419a,a78420a,a78424a,a78425a,a78428a,a78431a,a78432a,a78433a,a78436a,a78439a,a78440a,a78443a,a78446a,a78447a,a78448a,a78452a,a78453a,a78456a,a78459a,a78460a,a78461a,a78464a,a78467a,a78468a,a78471a,a78474a,a78475a,a78476a,a78480a,a78481a,a78484a,a78487a,a78488a,a78489a,a78492a,a78495a,a78496a,a78499a,a78502a,a78503a,a78504a,a78508a,a78509a,a78512a,a78515a,a78516a,a78517a,a78520a,a78523a,a78524a,a78527a,a78530a,a78531a,a78532a,a78536a,a78537a,a78540a,a78543a,a78544a,a78545a,a78548a,a78551a,a78552a,a78555a,a78558a,a78559a,a78560a,a78564a,a78565a,a78568a,a78571a,a78572a,a78573a,a78576a,a78579a,a78580a,a78583a,a78586a,a78587a,a78588a,a78592a,a78593a,a78596a,a78599a,a78600a,a78601a,a78604a,a78607a,a78608a,a78611a,a78614a,a78615a,a78616a,a78620a,a78621a,a78624a,a78627a,a78628a,a78629a,a78632a,a78635a,a78636a,a78639a,a78642a,a78643a,a78644a,a78648a,a78649a,a78652a,a78655a,a78656a,a78657a,a78660a,a78663a,a78664a,a78667a,a78670a,a78671a,a78672a,a78676a,a78677a,a78680a,a78683a,a78684a,a78685a,a78688a,a78691a,a78692a,a78695a,a78698a,a78699a,a78700a,a78704a,a78705a,a78708a,a78711a,a78712a,a78713a,a78716a,a78719a,a78720a,a78723a,a78726a,a78727a,a78728a,a78732a,a78733a,a78736a,a78739a,a78740a,a78741a,a78744a,a78747a,a78748a,a78751a,a78754a,a78755a,a78756a,a78760a,a78761a,a78764a,a78767a,a78768a,a78769a,a78772a,a78775a,a78776a,a78779a,a78782a,a78783a,a78784a,a78788a,a78789a,a78792a,a78795a,a78796a,a78797a,a78800a,a78803a,a78804a,a78807a,a78810a,a78811a,a78812a,a78816a,a78817a,a78820a,a78823a,a78824a,a78825a,a78828a,a78831a,a78832a,a78835a,a78838a,a78839a,a78840a,a78844a,a78845a,a78848a,a78851a,a78852a,a78853a,a78856a,a78859a,a78860a,a78863a,a78866a,a78867a,a78868a,a78872a,a78873a,a78876a,a78879a,a78880a,a78881a,a78884a,a78887a,a78888a,a78891a,a78894a,a78895a,a78896a,a78900a,a78901a,a78904a,a78907a,a78908a,a78909a,a78912a,a78915a,a78916a,a78919a,a78922a,a78923a,a78924a,a78928a,a78929a,a78932a,a78935a,a78936a,a78937a,a78940a,a78943a,a78944a,a78947a,a78950a,a78951a,a78952a,a78956a,a78957a,a78960a,a78963a,a78964a,a78965a,a78968a,a78971a,a78972a,a78975a,a78978a,a78979a,a78980a,a78984a,a78985a,a78988a,a78991a,a78992a,a78993a,a78996a,a78999a,a79000a,a79003a,a79006a,a79007a,a79008a,a79012a,a79013a,a79016a,a79019a,a79020a,a79021a,a79024a,a79027a,a79028a,a79031a,a79034a,a79035a,a79036a,a79040a,a79041a,a79044a,a79047a,a79048a,a79049a,a79052a,a79055a,a79056a,a79059a,a79062a,a79063a,a79064a,a79068a,a79069a,a79072a,a79075a,a79076a,a79077a,a79080a,a79083a,a79084a,a79087a,a79090a,a79091a,a79092a,a79096a,a79097a,a79100a,a79103a,a79104a,a79105a,a79108a,a79111a,a79112a,a79115a,a79118a,a79119a,a79120a,a79124a,a79125a,a79128a,a79131a,a79132a,a79133a,a79136a,a79139a,a79140a,a79143a,a79146a,a79147a,a79148a,a79152a,a79153a,a79156a,a79159a,a79160a,a79161a,a79164a,a79167a,a79168a,a79171a,a79174a,a79175a,a79176a,a79180a,a79181a,a79184a,a79187a,a79188a,a79189a,a79192a,a79195a,a79196a,a79199a,a79202a,a79203a,a79204a,a79208a,a79209a,a79212a,a79215a,a79216a,a79217a,a79220a,a79223a,a79224a,a79227a,a79230a,a79231a,a79232a,a79236a,a79237a,a79240a,a79243a,a79244a,a79245a,a79248a,a79251a,a79252a,a79255a,a79258a,a79259a,a79260a,a79264a,a79265a,a79268a,a79271a,a79272a,a79273a,a79276a,a79279a,a79280a,a79283a,a79286a,a79287a,a79288a,a79292a,a79293a,a79296a,a79299a,a79300a,a79301a,a79304a,a79307a,a79308a,a79311a,a79314a,a79315a,a79316a,a79320a,a79321a,a79324a,a79327a,a79328a,a79329a,a79332a,a79335a,a79336a,a79339a,a79342a,a79343a,a79344a,a79348a,a79349a,a79352a,a79355a,a79356a,a79357a,a79360a,a79363a,a79364a,a79367a,a79370a,a79371a,a79372a,a79376a,a79377a,a79380a,a79383a,a79384a,a79385a,a79388a,a79391a,a79392a,a79395a,a79398a,a79399a,a79400a,a79404a,a79405a,a79408a,a79411a,a79412a,a79413a,a79416a,a79419a,a79420a,a79423a,a79426a,a79427a,a79428a,a79432a,a79433a,a79436a,a79439a,a79440a,a79441a,a79444a,a79447a,a79448a,a79451a,a79454a,a79455a,a79456a,a79460a,a79461a,a79464a,a79467a,a79468a,a79469a,a79472a,a79475a,a79476a,a79479a,a79482a,a79483a,a79484a,a79488a,a79489a,a79492a,a79495a,a79496a,a79497a,a79500a,a79503a,a79504a,a79507a,a79510a,a79511a,a79512a,a79516a,a79517a,a79520a,a79523a,a79524a,a79525a,a79528a,a79531a,a79532a,a79535a,a79538a,a79539a,a79540a,a79544a,a79545a,a79548a,a79551a,a79552a,a79553a,a79556a,a79559a,a79560a,a79563a,a79566a,a79567a,a79568a,a79572a,a79573a,a79576a,a79579a,a79580a,a79581a,a79584a,a79587a,a79588a,a79591a,a79594a,a79595a,a79596a,a79600a,a79601a,a79604a,a79607a,a79608a,a79609a,a79612a,a79615a,a79616a,a79619a,a79622a,a79623a,a79624a,a79628a,a79629a,a79632a,a79635a,a79636a,a79637a,a79640a,a79643a,a79644a,a79647a,a79650a,a79651a,a79652a,a79656a,a79657a,a79660a,a79663a,a79664a,a79665a,a79668a,a79671a,a79672a,a79675a,a79678a,a79679a,a79680a,a79684a,a79685a,a79688a,a79691a,a79692a,a79693a,a79696a,a79699a,a79700a,a79703a,a79706a,a79707a,a79708a,a79712a,a79713a,a79716a,a79719a,a79720a,a79721a,a79724a,a79727a,a79728a,a79731a,a79734a,a79735a,a79736a,a79740a,a79741a,a79744a,a79747a,a79748a,a79749a,a79752a,a79755a,a79756a,a79759a,a79762a,a79763a,a79764a,a79768a,a79769a,a79772a,a79775a,a79776a,a79777a,a79780a,a79783a,a79784a,a79787a,a79790a,a79791a,a79792a,a79796a,a79797a,a79800a,a79803a,a79804a,a79805a,a79808a,a79811a,a79812a,a79815a,a79818a,a79819a,a79820a,a79824a,a79825a,a79828a,a79831a,a79832a,a79833a,a79836a,a79839a,a79840a,a79843a,a79846a,a79847a,a79848a,a79852a,a79853a,a79856a,a79859a,a79860a,a79861a,a79864a,a79867a,a79868a,a79871a,a79874a,a79875a,a79876a,a79880a,a79881a,a79884a,a79887a,a79888a,a79889a,a79892a,a79895a,a79896a,a79899a,a79902a,a79903a,a79904a,a79908a,a79909a,a79912a,a79915a,a79916a,a79917a,a79920a,a79923a,a79924a,a79927a,a79930a,a79931a,a79932a,a79936a,a79937a,a79940a,a79943a,a79944a,a79945a,a79948a,a79951a,a79952a,a79955a,a79958a,a79959a,a79960a,a79964a,a79965a,a79968a,a79971a,a79972a,a79973a,a79976a,a79979a,a79980a,a79983a,a79986a,a79987a,a79988a,a79992a,a79993a,a79996a,a79999a,a80000a,a80001a,a80004a,a80007a,a80008a,a80011a,a80014a,a80015a,a80016a,a80020a,a80021a,a80024a,a80027a,a80028a,a80029a,a80032a,a80035a,a80036a,a80039a,a80042a,a80043a,a80044a,a80048a,a80049a,a80052a,a80055a,a80056a,a80057a,a80060a,a80063a,a80064a,a80067a,a80070a,a80071a,a80072a,a80076a,a80077a,a80080a,a80083a,a80084a,a80085a,a80088a,a80091a,a80092a,a80095a,a80098a,a80099a,a80100a,a80104a,a80105a,a80108a,a80111a,a80112a,a80113a,a80116a,a80119a,a80120a,a80123a,a80126a,a80127a,a80128a,a80132a,a80133a,a80136a,a80139a,a80140a,a80141a,a80144a,a80147a,a80148a,a80151a,a80154a,a80155a,a80156a,a80160a,a80161a,a80164a,a80167a,a80168a,a80169a,a80172a,a80175a,a80176a,a80179a,a80182a,a80183a,a80184a,a80188a,a80189a,a80192a,a80195a,a80196a,a80197a,a80200a,a80203a,a80204a,a80207a,a80210a,a80211a,a80212a,a80216a,a80217a,a80220a,a80223a,a80224a,a80225a,a80228a,a80231a,a80232a,a80235a,a80238a,a80239a,a80240a,a80244a,a80245a,a80248a,a80251a,a80252a,a80253a,a80256a,a80259a,a80260a,a80263a,a80266a,a80267a,a80268a,a80272a,a80273a,a80276a,a80279a,a80280a,a80281a,a80284a,a80287a,a80288a,a80291a,a80294a,a80295a,a80296a,a80300a,a80301a,a80304a,a80307a,a80308a,a80309a,a80312a,a80315a,a80316a,a80319a,a80322a,a80323a,a80324a,a80328a,a80329a,a80332a,a80335a,a80336a,a80337a,a80340a,a80343a,a80344a,a80347a,a80350a,a80351a,a80352a,a80356a,a80357a,a80360a,a80363a,a80364a,a80365a,a80368a,a80371a,a80372a,a80375a,a80378a,a80379a,a80380a,a80384a,a80385a,a80388a,a80391a,a80392a,a80393a,a80396a,a80399a,a80400a,a80403a,a80406a,a80407a,a80408a,a80412a,a80413a,a80416a,a80419a,a80420a,a80421a,a80424a,a80427a,a80428a,a80431a,a80434a,a80435a,a80436a,a80440a,a80441a,a80444a,a80447a,a80448a,a80449a,a80452a,a80455a,a80456a,a80459a,a80462a,a80463a,a80464a,a80468a,a80469a,a80472a,a80475a,a80476a,a80477a,a80480a,a80483a,a80484a,a80487a,a80490a,a80491a,a80492a,a80496a,a80497a,a80500a,a80503a,a80504a,a80505a,a80508a,a80511a,a80512a,a80515a,a80518a,a80519a,a80520a,a80524a,a80525a,a80528a,a80531a,a80532a,a80533a,a80536a,a80539a,a80540a,a80543a,a80546a,a80547a,a80548a,a80552a,a80553a,a80556a,a80559a,a80560a,a80561a,a80564a,a80567a,a80568a,a80571a,a80574a,a80575a,a80576a,a80580a,a80581a,a80584a,a80587a,a80588a,a80589a,a80592a,a80595a,a80596a,a80599a,a80602a,a80603a,a80604a,a80608a,a80609a,a80612a,a80615a,a80616a,a80617a,a80620a,a80623a,a80624a,a80627a,a80630a,a80631a,a80632a,a80636a,a80637a,a80640a,a80643a,a80644a,a80645a,a80648a,a80651a,a80652a,a80655a,a80658a,a80659a,a80660a,a80664a,a80665a,a80668a,a80671a,a80672a,a80673a,a80676a,a80679a,a80680a,a80683a,a80686a,a80687a,a80688a,a80692a,a80693a,a80696a,a80699a,a80700a,a80701a,a80704a,a80707a,a80708a,a80711a,a80714a,a80715a,a80716a,a80720a,a80721a,a80724a,a80727a,a80728a,a80729a,a80732a,a80735a,a80736a,a80739a,a80742a,a80743a,a80744a,a80748a,a80749a,a80752a,a80755a,a80756a,a80757a,a80760a,a80763a,a80764a,a80767a,a80770a,a80771a,a80772a,a80776a,a80777a,a80780a,a80783a,a80784a,a80785a,a80788a,a80791a,a80792a,a80795a,a80798a,a80799a,a80800a,a80804a,a80805a,a80808a,a80811a,a80812a,a80813a,a80816a,a80819a,a80820a,a80823a,a80826a,a80827a,a80828a,a80832a,a80833a,a80836a,a80839a,a80840a,a80841a,a80844a,a80847a,a80848a,a80851a,a80854a,a80855a,a80856a,a80860a,a80861a,a80864a,a80867a,a80868a,a80869a,a80872a,a80875a,a80876a,a80879a,a80882a,a80883a,a80884a,a80888a,a80889a,a80892a,a80895a,a80896a,a80897a,a80900a,a80903a,a80904a,a80907a,a80910a,a80911a,a80912a,a80916a,a80917a,a80920a,a80923a,a80924a,a80925a,a80928a,a80931a,a80932a,a80935a,a80938a,a80939a,a80940a,a80944a,a80945a,a80948a,a80951a,a80952a,a80953a,a80956a,a80959a,a80960a,a80963a,a80966a,a80967a,a80968a,a80972a,a80973a,a80976a,a80979a,a80980a,a80981a,a80984a,a80987a,a80988a,a80991a,a80994a,a80995a,a80996a,a81000a,a81001a,a81004a,a81007a,a81008a,a81009a,a81012a,a81015a,a81016a,a81019a,a81022a,a81023a,a81024a,a81028a,a81029a,a81032a,a81035a,a81036a,a81037a,a81040a,a81043a,a81044a,a81047a,a81050a,a81051a,a81052a,a81056a,a81057a,a81060a,a81063a,a81064a,a81065a,a81068a,a81071a,a81072a,a81075a,a81078a,a81079a,a81080a,a81084a,a81085a,a81088a,a81091a,a81092a,a81093a,a81096a,a81099a,a81100a,a81103a,a81106a,a81107a,a81108a,a81112a,a81113a,a81116a,a81119a,a81120a,a81121a,a81124a,a81127a,a81128a,a81131a,a81134a,a81135a,a81136a,a81140a,a81141a,a81144a,a81147a,a81148a,a81149a,a81152a,a81155a,a81156a,a81159a,a81162a,a81163a,a81164a,a81168a,a81169a,a81172a,a81175a,a81176a,a81177a,a81180a,a81183a,a81184a,a81187a,a81190a,a81191a,a81192a,a81196a,a81197a,a81200a,a81203a,a81204a,a81205a,a81208a,a81211a,a81212a,a81215a,a81218a,a81219a,a81220a,a81224a,a81225a,a81228a,a81231a,a81232a,a81233a,a81236a,a81239a,a81240a,a81243a,a81246a,a81247a,a81248a,a81252a,a81253a,a81256a,a81259a,a81260a,a81261a,a81264a,a81267a,a81268a,a81271a,a81274a,a81275a,a81276a,a81280a,a81281a,a81284a,a81287a,a81288a,a81289a,a81292a,a81295a,a81296a,a81299a,a81302a,a81303a,a81304a,a81308a,a81309a,a81312a,a81315a,a81316a,a81317a,a81320a,a81323a,a81324a,a81327a,a81330a,a81331a,a81332a,a81336a,a81337a,a81340a,a81343a,a81344a,a81345a,a81348a,a81351a,a81352a,a81355a,a81358a,a81359a,a81360a,a81364a,a81365a,a81368a,a81371a,a81372a,a81373a,a81376a,a81379a,a81380a,a81383a,a81386a,a81387a,a81388a,a81392a,a81393a,a81396a,a81399a,a81400a,a81401a,a81404a,a81407a,a81408a,a81411a,a81414a,a81415a,a81416a,a81420a,a81421a,a81424a,a81427a,a81428a,a81429a,a81432a,a81435a,a81436a,a81439a,a81442a,a81443a,a81444a,a81448a,a81449a,a81452a,a81455a,a81456a,a81457a,a81460a,a81463a,a81464a,a81467a,a81470a,a81471a,a81472a,a81476a,a81477a,a81480a,a81483a,a81484a,a81485a,a81488a,a81491a,a81492a,a81495a,a81498a,a81499a,a81500a,a81504a,a81505a,a81508a,a81511a,a81512a,a81513a,a81516a,a81519a,a81520a,a81523a,a81526a,a81527a,a81528a,a81532a,a81533a,a81536a,a81539a,a81540a,a81541a,a81544a,a81547a,a81548a,a81551a,a81554a,a81555a,a81556a,a81560a,a81561a,a81564a,a81567a,a81568a,a81569a,a81572a,a81575a,a81576a,a81579a,a81582a,a81583a,a81584a,a81588a,a81589a,a81592a,a81595a,a81596a,a81597a,a81600a,a81603a,a81604a,a81607a,a81610a,a81611a,a81612a,a81616a,a81617a,a81620a,a81623a,a81624a,a81625a,a81628a,a81631a,a81632a,a81635a,a81638a,a81639a,a81640a,a81644a,a81645a,a81648a,a81651a,a81652a,a81653a,a81656a,a81659a,a81660a,a81663a,a81666a,a81667a,a81668a,a81672a,a81673a,a81676a,a81679a,a81680a,a81681a,a81684a,a81687a,a81688a,a81691a,a81694a,a81695a,a81696a,a81700a,a81701a,a81704a,a81707a,a81708a,a81709a,a81712a,a81715a,a81716a,a81719a,a81722a,a81723a,a81724a,a81728a,a81729a,a81732a,a81735a,a81736a,a81737a,a81740a,a81743a,a81744a,a81747a,a81750a,a81751a,a81752a,a81756a,a81757a,a81760a,a81763a,a81764a,a81765a,a81768a,a81771a,a81772a,a81775a,a81778a,a81779a,a81780a,a81784a,a81785a,a81788a,a81791a,a81792a,a81793a,a81796a,a81799a,a81800a,a81803a,a81806a,a81807a,a81808a,a81812a,a81813a,a81816a,a81819a,a81820a,a81821a,a81824a,a81827a,a81828a,a81831a,a81834a,a81835a,a81836a,a81840a,a81841a,a81844a,a81847a,a81848a,a81849a,a81852a,a81855a,a81856a,a81859a,a81862a,a81863a,a81864a,a81868a,a81869a,a81872a,a81875a,a81876a,a81877a,a81880a,a81883a,a81884a,a81887a,a81890a,a81891a,a81892a,a81896a,a81897a,a81900a,a81903a,a81904a,a81905a,a81908a,a81911a,a81912a,a81915a,a81918a,a81919a,a81920a,a81924a,a81925a,a81928a,a81931a,a81932a,a81933a,a81936a,a81939a,a81940a,a81943a,a81946a,a81947a,a81948a,a81952a,a81953a,a81956a,a81959a,a81960a,a81961a,a81964a,a81967a,a81968a,a81971a,a81974a,a81975a,a81976a,a81980a,a81981a,a81984a,a81987a,a81988a,a81989a,a81992a,a81995a,a81996a,a81999a,a82002a,a82003a,a82004a,a82008a,a82009a,a82012a,a82015a,a82016a,a82017a,a82020a,a82023a,a82024a,a82027a,a82030a,a82031a,a82032a,a82036a,a82037a,a82040a,a82043a,a82044a,a82045a,a82048a,a82051a,a82052a,a82055a,a82058a,a82059a,a82060a,a82064a,a82065a,a82068a,a82071a,a82072a,a82073a,a82076a,a82079a,a82080a,a82083a,a82086a,a82087a,a82088a,a82092a,a82093a,a82096a,a82099a,a82100a,a82101a,a82104a,a82107a,a82108a,a82111a,a82114a,a82115a,a82116a,a82120a,a82121a,a82124a,a82127a,a82128a,a82129a,a82132a,a82135a,a82136a,a82139a,a82142a,a82143a,a82144a,a82148a,a82149a,a82152a,a82155a,a82156a,a82157a,a82160a,a82163a,a82164a,a82167a,a82170a,a82171a,a82172a,a82176a,a82177a,a82180a,a82183a,a82184a,a82185a,a82188a,a82191a,a82192a,a82195a,a82198a,a82199a,a82200a,a82204a,a82205a,a82208a,a82211a,a82212a,a82213a,a82216a,a82219a,a82220a,a82223a,a82226a,a82227a,a82228a,a82232a,a82233a,a82236a,a82239a,a82240a,a82241a,a82244a,a82247a,a82248a,a82251a,a82254a,a82255a,a82256a,a82260a,a82261a,a82264a,a82267a,a82268a,a82269a,a82272a,a82275a,a82276a,a82279a,a82282a,a82283a,a82284a,a82288a,a82289a,a82292a,a82295a,a82296a,a82297a,a82300a,a82303a,a82304a,a82307a,a82310a,a82311a,a82312a,a82316a,a82317a,a82320a,a82323a,a82324a,a82325a,a82328a,a82331a,a82332a,a82335a,a82338a,a82339a,a82340a,a82344a,a82345a,a82348a,a82351a,a82352a,a82353a,a82356a,a82359a,a82360a,a82363a,a82366a,a82367a,a82368a,a82372a,a82373a,a82376a,a82379a,a82380a,a82381a,a82384a,a82387a,a82388a,a82391a,a82394a,a82395a,a82396a,a82400a,a82401a,a82404a,a82407a,a82408a,a82409a,a82412a,a82415a,a82416a,a82419a,a82422a,a82423a,a82424a,a82428a,a82429a,a82432a,a82435a,a82436a,a82437a,a82440a,a82443a,a82444a,a82447a,a82450a,a82451a,a82452a,a82456a,a82457a,a82460a,a82463a,a82464a,a82465a,a82468a,a82471a,a82472a,a82475a,a82478a,a82479a,a82480a,a82484a,a82485a,a82488a,a82491a,a82492a,a82493a,a82496a,a82499a,a82500a,a82503a,a82506a,a82507a,a82508a,a82512a,a82513a,a82516a,a82519a,a82520a,a82521a,a82524a,a82527a,a82528a,a82531a,a82534a,a82535a,a82536a,a82540a,a82541a,a82544a,a82547a,a82548a,a82549a,a82552a,a82555a,a82556a,a82559a,a82562a,a82563a,a82564a,a82568a,a82569a,a82572a,a82575a,a82576a,a82577a,a82580a,a82583a,a82584a,a82587a,a82590a,a82591a,a82592a,a82596a,a82597a,a82600a,a82603a,a82604a,a82605a,a82608a,a82611a,a82612a,a82615a,a82618a,a82619a,a82620a,a82624a,a82625a,a82628a,a82631a,a82632a,a82633a,a82636a,a82639a,a82640a,a82643a,a82646a,a82647a,a82648a,a82652a,a82653a,a82656a,a82659a,a82660a,a82661a,a82664a,a82667a,a82668a,a82671a,a82674a,a82675a,a82676a,a82680a,a82681a,a82684a,a82687a,a82688a,a82689a,a82692a,a82695a,a82696a,a82699a,a82702a,a82703a,a82704a,a82708a,a82709a,a82712a,a82715a,a82716a,a82717a,a82720a,a82723a,a82724a,a82727a,a82730a,a82731a,a82732a,a82736a,a82737a,a82740a,a82743a,a82744a,a82745a,a82748a,a82751a,a82752a,a82755a,a82758a,a82759a,a82760a,a82764a,a82765a,a82768a,a82771a,a82772a,a82773a,a82776a,a82779a,a82780a,a82783a,a82786a,a82787a,a82788a,a82792a,a82793a,a82796a,a82799a,a82800a,a82801a,a82804a,a82807a,a82808a,a82811a,a82814a,a82815a,a82816a,a82820a,a82821a,a82824a,a82827a,a82828a,a82829a,a82832a,a82835a,a82836a,a82839a,a82842a,a82843a,a82844a,a82848a,a82849a,a82852a,a82855a,a82856a,a82857a,a82860a,a82863a,a82864a,a82867a,a82870a,a82871a,a82872a,a82876a,a82877a,a82880a,a82883a,a82884a,a82885a,a82888a,a82891a,a82892a,a82895a,a82898a,a82899a,a82900a,a82904a,a82905a,a82908a,a82911a,a82912a,a82913a,a82916a,a82919a,a82920a,a82923a,a82926a,a82927a,a82928a,a82932a,a82933a,a82936a,a82939a,a82940a,a82941a,a82944a,a82947a,a82948a,a82951a,a82954a,a82955a,a82956a,a82960a,a82961a,a82964a,a82967a,a82968a,a82969a,a82972a,a82975a,a82976a,a82979a,a82982a,a82983a,a82984a,a82988a,a82989a,a82992a,a82995a,a82996a,a82997a,a83000a,a83003a,a83004a,a83007a,a83010a,a83011a,a83012a,a83016a,a83017a,a83020a,a83023a,a83024a,a83025a,a83028a,a83031a,a83032a,a83035a,a83038a,a83039a,a83040a,a83044a,a83045a,a83048a,a83051a,a83052a,a83053a,a83056a,a83059a,a83060a,a83063a,a83066a,a83067a,a83068a,a83072a,a83073a,a83076a,a83079a,a83080a,a83081a,a83084a,a83087a,a83088a,a83091a,a83094a,a83095a,a83096a,a83100a,a83101a,a83104a,a83107a,a83108a,a83109a,a83112a,a83115a,a83116a,a83119a,a83122a,a83123a,a83124a,a83128a,a83129a,a83132a,a83135a,a83136a,a83137a,a83140a,a83143a,a83144a,a83147a,a83150a,a83151a,a83152a,a83156a,a83157a,a83160a,a83163a,a83164a,a83165a,a83168a,a83171a,a83172a,a83175a,a83178a,a83179a,a83180a,a83184a,a83185a,a83188a,a83191a,a83192a,a83193a,a83196a,a83199a,a83200a,a83203a,a83206a,a83207a,a83208a,a83212a,a83213a,a83216a,a83219a,a83220a,a83221a,a83224a,a83227a,a83228a,a83231a,a83234a,a83235a,a83236a,a83240a,a83241a,a83244a,a83247a,a83248a,a83249a,a83252a,a83255a,a83256a,a83259a,a83262a,a83263a,a83264a,a83268a,a83269a,a83272a,a83275a,a83276a,a83277a,a83280a,a83283a,a83284a,a83287a,a83290a,a83291a,a83292a,a83296a,a83297a,a83300a,a83303a,a83304a,a83305a,a83308a,a83311a,a83312a,a83315a,a83318a,a83319a,a83320a,a83324a,a83325a,a83328a,a83331a,a83332a,a83333a,a83336a,a83339a,a83340a,a83343a,a83346a,a83347a,a83348a,a83352a,a83353a,a83356a,a83359a,a83360a,a83361a,a83364a,a83367a,a83368a,a83371a,a83374a,a83375a,a83376a,a83380a,a83381a,a83384a,a83387a,a83388a,a83389a,a83392a,a83395a,a83396a,a83399a,a83402a,a83403a,a83404a,a83408a,a83409a,a83412a,a83415a,a83416a,a83417a,a83420a,a83423a,a83424a,a83427a,a83430a,a83431a,a83432a,a83436a,a83437a,a83440a,a83443a,a83444a,a83445a,a83448a,a83451a,a83452a,a83455a,a83458a,a83459a,a83460a,a83464a,a83465a,a83468a,a83471a,a83472a,a83473a,a83476a,a83479a,a83480a,a83483a,a83486a,a83487a,a83488a,a83492a,a83493a,a83496a,a83499a,a83500a,a83501a,a83504a,a83507a,a83508a,a83511a,a83514a,a83515a,a83516a,a83520a,a83521a,a83524a,a83527a,a83528a,a83529a,a83532a,a83535a,a83536a,a83539a,a83542a,a83543a,a83544a,a83548a,a83549a,a83552a,a83555a,a83556a,a83557a,a83560a,a83563a,a83564a,a83567a,a83570a,a83571a,a83572a,a83576a,a83577a,a83580a,a83583a,a83584a,a83585a,a83588a,a83591a,a83592a,a83595a,a83598a,a83599a,a83600a,a83604a,a83605a,a83608a,a83611a,a83612a,a83613a,a83616a,a83619a,a83620a,a83623a,a83626a,a83627a,a83628a,a83632a,a83633a,a83636a,a83639a,a83640a,a83641a,a83644a,a83647a,a83648a,a83651a,a83654a,a83655a,a83656a,a83660a,a83661a,a83664a,a83667a,a83668a,a83669a,a83672a,a83675a,a83676a,a83679a,a83682a,a83683a,a83684a,a83688a,a83689a,a83692a,a83695a,a83696a,a83697a,a83700a,a83703a,a83704a,a83707a,a83710a,a83711a,a83712a,a83716a,a83717a,a83720a,a83723a,a83724a,a83725a,a83728a,a83731a,a83732a,a83735a,a83738a,a83739a,a83740a,a83744a,a83745a,a83748a,a83751a,a83752a,a83753a,a83756a,a83759a,a83760a,a83763a,a83766a,a83767a,a83768a,a83772a,a83773a,a83776a,a83779a,a83780a,a83781a,a83784a,a83787a,a83788a,a83791a,a83794a,a83795a,a83796a,a83800a,a83801a,a83804a,a83807a,a83808a,a83809a,a83812a,a83815a,a83816a,a83819a,a83822a,a83823a,a83824a,a83828a,a83829a,a83832a,a83835a,a83836a,a83837a,a83840a,a83843a,a83844a,a83847a,a83850a,a83851a,a83852a,a83856a,a83857a,a83860a,a83863a,a83864a,a83865a,a83868a,a83871a,a83872a,a83875a,a83878a,a83879a,a83880a,a83884a,a83885a,a83888a,a83891a,a83892a,a83893a,a83896a,a83899a,a83900a,a83903a,a83906a,a83907a,a83908a,a83912a,a83913a,a83916a,a83919a,a83920a,a83921a,a83924a,a83927a,a83928a,a83931a,a83934a,a83935a,a83936a,a83940a,a83941a,a83944a,a83947a,a83948a,a83949a,a83952a,a83955a,a83956a,a83959a,a83962a,a83963a,a83964a,a83968a,a83969a,a83972a,a83975a,a83976a,a83977a,a83980a,a83983a,a83984a,a83987a,a83990a,a83991a,a83992a,a83996a,a83997a,a84000a,a84003a,a84004a,a84005a,a84008a,a84011a,a84012a,a84015a,a84018a,a84019a,a84020a,a84024a,a84025a,a84028a,a84031a,a84032a,a84033a,a84036a,a84039a,a84040a,a84043a,a84046a,a84047a,a84048a,a84052a,a84053a,a84056a,a84059a,a84060a,a84061a,a84064a,a84067a,a84068a,a84071a,a84074a,a84075a,a84076a,a84080a,a84081a,a84084a,a84087a,a84088a,a84089a,a84092a,a84095a,a84096a,a84099a,a84102a,a84103a,a84104a,a84108a,a84109a,a84112a,a84115a,a84116a,a84117a,a84120a,a84123a,a84124a,a84127a,a84130a,a84131a,a84132a,a84136a,a84137a,a84140a,a84143a,a84144a,a84145a,a84148a,a84151a,a84152a,a84155a,a84158a,a84159a,a84160a,a84164a,a84165a,a84168a,a84171a,a84172a,a84173a,a84176a,a84179a,a84180a,a84183a,a84186a,a84187a,a84188a,a84192a,a84193a,a84196a,a84199a,a84200a,a84201a,a84204a,a84207a,a84208a,a84211a,a84214a,a84215a,a84216a,a84220a,a84221a,a84224a,a84227a,a84228a,a84229a,a84232a,a84235a,a84236a,a84239a,a84242a,a84243a,a84244a,a84248a,a84249a,a84252a,a84255a,a84256a,a84257a,a84260a,a84263a,a84264a,a84267a,a84270a,a84271a,a84272a,a84276a,a84277a,a84280a,a84283a,a84284a,a84285a,a84288a,a84291a,a84292a,a84295a,a84298a,a84299a,a84300a,a84304a,a84305a,a84308a,a84311a,a84312a,a84313a,a84316a,a84319a,a84320a,a84323a,a84326a,a84327a,a84328a,a84332a,a84333a,a84336a,a84339a,a84340a,a84341a,a84344a,a84347a,a84348a,a84351a,a84354a,a84355a,a84356a,a84360a,a84361a,a84364a,a84367a,a84368a,a84369a,a84372a,a84375a,a84376a,a84379a,a84382a,a84383a,a84384a,a84388a,a84389a,a84392a,a84395a,a84396a,a84397a,a84400a,a84403a,a84404a,a84407a,a84410a,a84411a,a84412a,a84416a,a84417a,a84420a,a84423a,a84424a,a84425a,a84428a,a84431a,a84432a,a84435a,a84438a,a84439a,a84440a,a84444a,a84445a,a84448a,a84451a,a84452a,a84453a,a84456a,a84459a,a84460a,a84463a,a84466a,a84467a,a84468a,a84472a,a84473a,a84476a,a84479a,a84480a,a84481a,a84484a,a84487a,a84488a,a84491a,a84494a,a84495a,a84496a,a84500a,a84501a,a84504a,a84507a,a84508a,a84509a,a84512a,a84515a,a84516a,a84519a,a84522a,a84523a,a84524a,a84528a,a84529a,a84532a,a84535a,a84536a,a84537a,a84540a,a84543a,a84544a,a84547a,a84550a,a84551a,a84552a,a84556a,a84557a,a84560a,a84563a,a84564a,a84565a,a84568a,a84571a,a84572a,a84575a,a84578a,a84579a,a84580a,a84584a,a84585a,a84588a,a84591a,a84592a,a84593a,a84596a,a84599a,a84600a,a84603a,a84606a,a84607a,a84608a,a84612a,a84613a,a84616a,a84619a,a84620a,a84621a,a84624a,a84627a,a84628a,a84631a,a84634a,a84635a,a84636a,a84640a,a84641a,a84644a,a84647a,a84648a,a84649a,a84652a,a84655a,a84656a,a84659a,a84662a,a84663a,a84664a,a84668a,a84669a,a84672a,a84675a,a84676a,a84677a,a84680a,a84683a,a84684a,a84687a,a84690a,a84691a,a84692a,a84696a,a84697a,a84700a,a84703a,a84704a,a84705a,a84708a,a84711a,a84712a,a84715a,a84718a,a84719a,a84720a,a84724a,a84725a,a84728a,a84731a,a84732a,a84733a,a84736a,a84739a,a84740a,a84743a,a84746a,a84747a,a84748a,a84752a,a84753a,a84756a,a84759a,a84760a,a84761a,a84764a,a84767a,a84768a,a84771a,a84774a,a84775a,a84776a,a84780a,a84781a,a84784a,a84787a,a84788a,a84789a,a84792a,a84795a,a84796a,a84799a,a84802a,a84803a,a84804a,a84808a,a84809a,a84812a,a84815a,a84816a,a84817a,a84820a,a84823a,a84824a,a84827a,a84830a,a84831a,a84832a,a84836a,a84837a,a84840a,a84843a,a84844a,a84845a,a84848a,a84851a,a84852a,a84855a,a84858a,a84859a,a84860a,a84864a,a84865a,a84868a,a84871a,a84872a,a84873a,a84876a,a84879a,a84880a,a84883a,a84886a,a84887a,a84888a,a84892a,a84893a,a84896a,a84899a,a84900a,a84901a,a84904a,a84907a,a84908a,a84911a,a84914a,a84915a,a84916a,a84920a,a84921a,a84924a,a84927a,a84928a,a84929a,a84932a,a84935a,a84936a,a84939a,a84942a,a84943a,a84944a,a84948a,a84949a,a84952a,a84955a,a84956a,a84957a,a84960a,a84963a,a84964a,a84967a,a84970a,a84971a,a84972a,a84976a,a84977a,a84980a,a84983a,a84984a,a84985a,a84988a,a84991a,a84992a,a84995a,a84998a,a84999a,a85000a,a85004a,a85005a,a85008a,a85011a,a85012a,a85013a,a85016a,a85019a,a85020a,a85023a,a85026a,a85027a,a85028a,a85032a,a85033a,a85036a,a85039a,a85040a,a85041a,a85044a,a85047a,a85048a,a85051a,a85054a,a85055a,a85056a,a85060a,a85061a,a85064a,a85067a,a85068a,a85069a,a85072a,a85075a,a85076a,a85079a,a85082a,a85083a,a85084a,a85088a,a85089a,a85092a,a85095a,a85096a,a85097a,a85100a,a85103a,a85104a,a85107a,a85110a,a85111a,a85112a,a85116a,a85117a,a85120a,a85123a,a85124a,a85125a,a85128a,a85131a,a85132a,a85135a,a85138a,a85139a,a85140a,a85144a,a85145a,a85148a,a85151a,a85152a,a85153a,a85156a,a85159a,a85160a,a85163a,a85166a,a85167a,a85168a,a85172a,a85173a,a85176a,a85179a,a85180a,a85181a,a85184a,a85187a,a85188a,a85191a,a85194a,a85195a,a85196a,a85200a,a85201a,a85204a,a85207a,a85208a,a85209a,a85212a,a85215a,a85216a,a85219a,a85222a,a85223a,a85224a,a85228a,a85229a,a85232a,a85235a,a85236a,a85237a,a85240a,a85243a,a85244a,a85247a,a85250a,a85251a,a85252a,a85256a,a85257a,a85260a,a85263a,a85264a,a85265a,a85268a,a85271a,a85272a,a85275a,a85278a,a85279a,a85280a,a85284a,a85285a,a85288a,a85291a,a85292a,a85293a,a85296a,a85299a,a85300a,a85303a,a85306a,a85307a,a85308a,a85312a,a85313a,a85316a,a85319a,a85320a,a85321a,a85324a,a85327a,a85328a,a85331a,a85334a,a85335a,a85336a,a85340a,a85341a,a85344a,a85347a,a85348a,a85349a,a85352a,a85355a,a85356a,a85359a,a85362a,a85363a,a85364a,a85368a,a85369a,a85372a,a85375a,a85376a,a85377a,a85380a,a85383a,a85384a,a85387a,a85390a,a85391a,a85392a,a85396a,a85397a,a85400a,a85403a,a85404a,a85405a,a85408a,a85411a,a85412a,a85415a,a85418a,a85419a,a85420a,a85424a,a85425a,a85428a,a85431a,a85432a,a85433a,a85436a,a85439a,a85440a,a85443a,a85446a,a85447a,a85448a,a85452a,a85453a,a85456a,a85459a,a85460a,a85461a,a85464a,a85467a,a85468a,a85471a,a85474a,a85475a,a85476a,a85480a,a85481a,a85484a,a85487a,a85488a,a85489a,a85492a,a85495a,a85496a,a85499a,a85502a,a85503a,a85504a,a85508a,a85509a,a85512a,a85515a,a85516a,a85517a,a85520a,a85523a,a85524a,a85527a,a85530a,a85531a,a85532a,a85536a,a85537a,a85540a,a85543a,a85544a,a85545a,a85548a,a85551a,a85552a,a85555a,a85558a,a85559a,a85560a,a85564a,a85565a,a85568a,a85571a,a85572a,a85573a,a85576a,a85579a,a85580a,a85583a,a85586a,a85587a,a85588a,a85592a,a85593a,a85596a,a85599a,a85600a,a85601a,a85604a,a85607a,a85608a,a85611a,a85614a,a85615a,a85616a,a85620a,a85621a,a85624a,a85627a,a85628a,a85629a,a85632a,a85635a,a85636a,a85639a,a85642a,a85643a,a85644a,a85648a,a85649a,a85652a,a85655a,a85656a,a85657a,a85660a,a85663a,a85664a,a85667a,a85670a,a85671a,a85672a,a85676a,a85677a,a85680a,a85683a,a85684a,a85685a,a85688a,a85691a,a85692a,a85695a,a85698a,a85699a,a85700a,a85704a,a85705a,a85708a,a85711a,a85712a,a85713a,a85716a,a85719a,a85720a,a85723a,a85726a,a85727a,a85728a,a85732a,a85733a,a85736a,a85739a,a85740a,a85741a,a85744a,a85747a,a85748a,a85751a,a85754a,a85755a,a85756a,a85760a,a85761a,a85764a,a85767a,a85768a,a85769a,a85772a,a85775a,a85776a,a85779a,a85782a,a85783a,a85784a,a85788a,a85789a,a85792a,a85795a,a85796a,a85797a,a85800a,a85803a,a85804a,a85807a,a85810a,a85811a,a85812a,a85816a,a85817a,a85820a,a85823a,a85824a,a85825a,a85828a,a85831a,a85832a,a85835a,a85838a,a85839a,a85840a,a85844a,a85845a,a85848a,a85851a,a85852a,a85853a,a85856a,a85859a,a85860a,a85863a,a85866a,a85867a,a85868a,a85872a,a85873a,a85876a,a85879a,a85880a,a85881a,a85884a,a85887a,a85888a,a85891a,a85894a,a85895a,a85896a,a85900a,a85901a,a85904a,a85907a,a85908a,a85909a,a85912a,a85915a,a85916a,a85919a,a85922a,a85923a,a85924a,a85928a,a85929a,a85932a,a85935a,a85936a,a85937a,a85940a,a85943a,a85944a,a85947a,a85950a,a85951a,a85952a,a85956a,a85957a,a85960a,a85963a,a85964a,a85965a,a85968a,a85971a,a85972a,a85975a,a85978a,a85979a,a85980a,a85984a,a85985a,a85988a,a85991a,a85992a,a85993a,a85996a,a85999a,a86000a,a86003a,a86006a,a86007a,a86008a,a86012a,a86013a,a86016a,a86019a,a86020a,a86021a,a86024a,a86027a,a86028a,a86031a,a86034a,a86035a,a86036a,a86040a,a86041a,a86044a,a86047a,a86048a,a86049a,a86052a,a86055a,a86056a,a86059a,a86062a,a86063a,a86064a,a86068a,a86069a,a86072a,a86075a,a86076a,a86077a,a86080a,a86083a,a86084a,a86087a,a86090a,a86091a,a86092a,a86096a,a86097a,a86100a,a86103a,a86104a,a86105a,a86108a,a86111a,a86112a,a86115a,a86118a,a86119a,a86120a,a86124a,a86125a,a86128a,a86131a,a86132a,a86133a,a86136a,a86139a,a86140a,a86143a,a86146a,a86147a,a86148a,a86152a,a86153a,a86156a,a86159a,a86160a,a86161a,a86164a,a86167a,a86168a,a86171a,a86174a,a86175a,a86176a,a86180a,a86181a,a86184a,a86187a,a86188a,a86189a,a86192a,a86195a,a86196a,a86199a,a86202a,a86203a,a86204a,a86208a,a86209a,a86212a,a86215a,a86216a,a86217a,a86220a,a86223a,a86224a,a86227a,a86230a,a86231a,a86232a,a86236a,a86237a,a86240a,a86243a,a86244a,a86245a,a86248a,a86251a,a86252a,a86255a,a86258a,a86259a,a86260a,a86264a,a86265a,a86268a,a86271a,a86272a,a86273a,a86276a,a86279a,a86280a,a86283a,a86286a,a86287a,a86288a,a86292a,a86293a,a86296a,a86299a,a86300a,a86301a,a86304a,a86307a,a86308a,a86311a,a86314a,a86315a,a86316a,a86320a,a86321a,a86324a,a86327a,a86328a,a86329a,a86332a,a86335a,a86336a,a86339a,a86342a,a86343a,a86344a,a86348a,a86349a,a86352a,a86355a,a86356a,a86357a,a86360a,a86363a,a86364a,a86367a,a86370a,a86371a,a86372a,a86376a,a86377a,a86380a,a86383a,a86384a,a86385a,a86388a,a86391a,a86392a,a86395a,a86398a,a86399a,a86400a,a86404a,a86405a,a86408a,a86411a,a86412a,a86413a,a86416a,a86419a,a86420a,a86423a,a86426a,a86427a,a86428a,a86432a,a86433a,a86436a,a86439a,a86440a,a86441a,a86444a,a86447a,a86448a,a86451a,a86454a,a86455a,a86456a,a86460a,a86461a,a86464a,a86467a,a86468a,a86469a,a86472a,a86475a,a86476a,a86479a,a86482a,a86483a,a86484a,a86488a,a86489a,a86492a,a86495a,a86496a,a86497a,a86500a,a86503a,a86504a,a86507a,a86510a,a86511a,a86512a,a86516a,a86517a,a86520a,a86523a,a86524a,a86525a,a86528a,a86531a,a86532a,a86535a,a86538a,a86539a,a86540a,a86544a,a86545a,a86548a,a86551a,a86552a,a86553a,a86556a,a86559a,a86560a,a86563a,a86566a,a86567a,a86568a,a86572a,a86573a,a86576a,a86579a,a86580a,a86581a,a86584a,a86587a,a86588a,a86591a,a86594a,a86595a,a86596a,a86600a,a86601a,a86604a,a86607a,a86608a,a86609a,a86612a,a86615a,a86616a,a86619a,a86622a,a86623a,a86624a,a86628a,a86629a,a86632a,a86635a,a86636a,a86637a,a86640a,a86643a,a86644a,a86647a,a86650a,a86651a,a86652a,a86656a,a86657a,a86660a,a86663a,a86664a,a86665a,a86668a,a86671a,a86672a,a86675a,a86678a,a86679a,a86680a,a86684a,a86685a,a86688a,a86691a,a86692a,a86693a,a86696a,a86699a,a86700a,a86703a,a86706a,a86707a,a86708a,a86712a,a86713a,a86716a,a86719a,a86720a,a86721a,a86724a,a86727a,a86728a,a86731a,a86734a,a86735a,a86736a,a86740a,a86741a,a86744a,a86747a,a86748a,a86749a,a86752a,a86755a,a86756a,a86759a,a86762a,a86763a,a86764a,a86768a,a86769a,a86772a,a86775a,a86776a,a86777a,a86780a,a86783a,a86784a,a86787a,a86790a,a86791a,a86792a,a86796a,a86797a,a86800a,a86803a,a86804a,a86805a,a86808a,a86811a,a86812a,a86815a,a86818a,a86819a,a86820a,a86824a,a86825a,a86828a,a86831a,a86832a,a86833a,a86836a,a86839a,a86840a,a86843a,a86846a,a86847a,a86848a,a86852a,a86853a,a86856a,a86859a,a86860a,a86861a,a86864a,a86867a,a86868a,a86871a,a86874a,a86875a,a86876a,a86880a,a86881a,a86884a,a86887a,a86888a,a86889a,a86892a,a86895a,a86896a,a86899a,a86902a,a86903a,a86904a,a86908a,a86909a,a86912a,a86915a,a86916a,a86917a,a86920a,a86923a,a86924a,a86927a,a86930a,a86931a,a86932a,a86936a,a86937a,a86940a,a86943a,a86944a,a86945a,a86948a,a86951a,a86952a,a86955a,a86958a,a86959a,a86960a,a86964a,a86965a,a86968a,a86971a,a86972a,a86973a,a86976a,a86979a,a86980a,a86983a,a86986a,a86987a,a86988a,a86992a,a86993a,a86996a,a86999a,a87000a,a87001a,a87004a,a87007a,a87008a,a87011a,a87014a,a87015a,a87016a,a87020a,a87021a,a87024a,a87027a,a87028a,a87029a,a87032a,a87035a,a87036a,a87039a,a87042a,a87043a,a87044a,a87048a,a87049a,a87052a,a87055a,a87056a,a87057a,a87060a,a87063a,a87064a,a87067a,a87070a,a87071a,a87072a,a87076a,a87077a,a87080a,a87083a,a87084a,a87085a,a87088a,a87091a,a87092a,a87095a,a87098a,a87099a,a87100a,a87104a,a87105a,a87108a,a87111a,a87112a,a87113a,a87116a,a87119a,a87120a,a87123a,a87126a,a87127a,a87128a,a87132a,a87133a,a87136a,a87139a,a87140a,a87141a,a87144a,a87147a,a87148a,a87151a,a87154a,a87155a,a87156a,a87160a,a87161a,a87164a,a87167a,a87168a,a87169a,a87172a,a87175a,a87176a,a87179a,a87182a,a87183a,a87184a,a87188a,a87189a,a87192a,a87195a,a87196a,a87197a,a87200a,a87203a,a87204a,a87207a,a87210a,a87211a,a87212a,a87216a,a87217a,a87220a,a87223a,a87224a,a87225a,a87228a,a87231a,a87232a,a87235a,a87238a,a87239a,a87240a,a87244a,a87245a,a87248a,a87251a,a87252a,a87253a,a87256a,a87259a,a87260a,a87263a,a87266a,a87267a,a87268a,a87272a,a87273a,a87276a,a87279a,a87280a,a87281a,a87284a,a87287a,a87288a,a87291a,a87294a,a87295a,a87296a,a87300a,a87301a,a87304a,a87307a,a87308a,a87309a,a87312a,a87315a,a87316a,a87319a,a87322a,a87323a,a87324a,a87328a,a87329a,a87332a,a87335a,a87336a,a87337a,a87340a,a87343a,a87344a,a87347a,a87350a,a87351a,a87352a,a87356a,a87357a,a87360a,a87363a,a87364a,a87365a,a87368a,a87371a,a87372a,a87375a,a87378a,a87379a,a87380a,a87384a,a87385a,a87388a,a87391a,a87392a,a87393a,a87396a,a87399a,a87400a,a87403a,a87406a,a87407a,a87408a,a87412a,a87413a,a87416a,a87419a,a87420a,a87421a,a87424a,a87427a,a87428a,a87431a,a87434a,a87435a,a87436a,a87440a,a87441a,a87444a,a87447a,a87448a,a87449a,a87452a,a87455a,a87456a,a87459a,a87462a,a87463a,a87464a,a87468a,a87469a,a87472a,a87475a,a87476a,a87477a,a87480a,a87483a,a87484a,a87487a,a87490a,a87491a,a87492a,a87496a,a87497a,a87500a,a87503a,a87504a,a87505a,a87508a,a87511a,a87512a,a87515a,a87518a,a87519a,a87520a,a87524a,a87525a,a87528a,a87531a,a87532a,a87533a,a87536a,a87539a,a87540a,a87543a,a87546a,a87547a,a87548a,a87552a,a87553a,a87556a,a87559a,a87560a,a87561a,a87564a,a87567a,a87568a,a87571a,a87574a,a87575a,a87576a,a87580a,a87581a,a87584a,a87587a,a87588a,a87589a,a87592a,a87595a,a87596a,a87599a,a87602a,a87603a,a87604a,a87608a,a87609a,a87612a,a87615a,a87616a,a87617a,a87620a,a87623a,a87624a,a87627a,a87630a,a87631a,a87632a,a87636a,a87637a,a87640a,a87643a,a87644a,a87645a,a87648a,a87651a,a87652a,a87655a,a87658a,a87659a,a87660a,a87664a,a87665a,a87668a,a87671a,a87672a,a87673a,a87676a,a87679a,a87680a,a87683a,a87686a,a87687a,a87688a,a87692a,a87693a,a87696a,a87699a,a87700a,a87701a,a87704a,a87707a,a87708a,a87711a,a87714a,a87715a,a87716a,a87720a,a87721a,a87724a,a87727a,a87728a,a87729a,a87732a,a87735a,a87736a,a87739a,a87742a,a87743a,a87744a,a87748a,a87749a,a87752a,a87755a,a87756a,a87757a,a87760a,a87763a,a87764a,a87767a,a87770a,a87771a,a87772a,a87776a,a87777a,a87780a,a87783a,a87784a,a87785a,a87788a,a87791a,a87792a,a87795a,a87798a,a87799a,a87800a,a87804a,a87805a,a87808a,a87811a,a87812a,a87813a,a87816a,a87819a,a87820a,a87823a,a87826a,a87827a,a87828a,a87832a,a87833a,a87836a,a87839a,a87840a,a87841a,a87844a,a87847a,a87848a,a87851a,a87854a,a87855a,a87856a,a87860a,a87861a,a87864a,a87867a,a87868a,a87869a,a87872a,a87875a,a87876a,a87879a,a87882a,a87883a,a87884a,a87888a,a87889a,a87892a,a87895a,a87896a,a87897a,a87900a,a87903a,a87904a,a87907a,a87910a,a87911a,a87912a,a87916a,a87917a,a87920a,a87923a,a87924a,a87925a,a87928a,a87931a,a87932a,a87935a,a87938a,a87939a,a87940a,a87944a,a87945a,a87948a,a87951a,a87952a,a87953a,a87956a,a87959a,a87960a,a87963a,a87966a,a87967a,a87968a,a87972a,a87973a,a87976a,a87979a,a87980a,a87981a,a87984a,a87987a,a87988a,a87991a,a87994a,a87995a,a87996a,a88000a,a88001a,a88004a,a88007a,a88008a,a88009a,a88012a,a88015a,a88016a,a88019a,a88022a,a88023a,a88024a,a88028a,a88029a,a88032a,a88035a,a88036a,a88037a,a88040a,a88043a,a88044a,a88047a,a88050a,a88051a,a88052a,a88056a,a88057a,a88060a,a88063a,a88064a,a88065a,a88068a,a88071a,a88072a,a88075a,a88078a,a88079a,a88080a,a88084a,a88085a,a88088a,a88091a,a88092a,a88093a,a88096a,a88099a,a88100a,a88103a,a88106a,a88107a,a88108a,a88112a,a88113a,a88116a,a88119a,a88120a,a88121a,a88124a,a88127a,a88128a,a88131a,a88134a,a88135a,a88136a,a88140a,a88141a,a88144a,a88147a,a88148a,a88149a,a88152a,a88155a,a88156a,a88159a,a88162a,a88163a,a88164a,a88168a,a88169a,a88172a,a88175a,a88176a,a88177a,a88180a,a88183a,a88184a,a88187a,a88190a,a88191a,a88192a,a88196a,a88197a,a88200a,a88203a,a88204a,a88205a,a88208a,a88211a,a88212a,a88215a,a88218a,a88219a,a88220a,a88224a,a88225a,a88228a,a88231a,a88232a,a88233a,a88236a,a88239a,a88240a,a88243a,a88246a,a88247a,a88248a,a88252a,a88253a,a88256a,a88259a,a88260a,a88261a,a88264a,a88267a,a88268a,a88271a,a88274a,a88275a,a88276a,a88280a,a88281a,a88284a,a88287a,a88288a,a88289a,a88292a,a88295a,a88296a,a88299a,a88302a,a88303a,a88304a,a88308a,a88309a,a88312a,a88315a,a88316a,a88317a,a88320a,a88323a,a88324a,a88327a,a88330a,a88331a,a88332a,a88336a,a88337a,a88340a,a88343a,a88344a,a88345a,a88348a,a88351a,a88352a,a88355a,a88358a,a88359a,a88360a,a88364a,a88365a,a88368a,a88371a,a88372a,a88373a,a88376a,a88379a,a88380a,a88383a,a88386a,a88387a,a88388a,a88392a,a88393a,a88396a,a88399a,a88400a,a88401a,a88404a,a88407a,a88408a,a88411a,a88414a,a88415a,a88416a,a88420a,a88421a,a88424a,a88427a,a88428a,a88429a,a88432a,a88435a,a88436a,a88439a,a88442a,a88443a,a88444a,a88448a,a88449a,a88452a,a88455a,a88456a,a88457a,a88460a,a88463a,a88464a,a88467a,a88470a,a88471a,a88472a,a88476a,a88477a,a88480a,a88483a,a88484a,a88485a,a88488a,a88491a,a88492a,a88495a,a88498a,a88499a,a88500a,a88504a,a88505a,a88508a,a88511a,a88512a,a88513a,a88516a,a88519a,a88520a,a88523a,a88526a,a88527a,a88528a,a88532a,a88533a,a88536a,a88539a,a88540a,a88541a,a88544a,a88547a,a88548a,a88551a,a88554a,a88555a,a88556a,a88560a,a88561a,a88564a,a88567a,a88568a,a88569a,a88572a,a88575a,a88576a,a88579a,a88582a,a88583a,a88584a,a88588a,a88589a,a88592a,a88595a,a88596a,a88597a,a88600a,a88603a,a88604a,a88607a,a88610a,a88611a,a88612a,a88616a,a88617a,a88620a,a88623a,a88624a,a88625a,a88628a,a88631a,a88632a,a88635a,a88638a,a88639a,a88640a,a88644a,a88645a,a88648a,a88651a,a88652a,a88653a,a88656a,a88659a,a88660a,a88663a,a88666a,a88667a,a88668a,a88672a,a88673a,a88676a,a88679a,a88680a,a88681a,a88684a,a88687a,a88688a,a88691a,a88694a,a88695a,a88696a,a88700a,a88701a,a88704a,a88707a,a88708a,a88709a,a88712a,a88715a,a88716a,a88719a,a88722a,a88723a,a88724a,a88728a,a88729a,a88732a,a88735a,a88736a,a88737a,a88740a,a88743a,a88744a,a88747a,a88750a,a88751a,a88752a,a88756a,a88757a,a88760a,a88763a,a88764a,a88765a,a88768a,a88771a,a88772a,a88775a,a88778a,a88779a,a88780a,a88784a,a88785a,a88788a,a88791a,a88792a,a88793a,a88796a,a88799a,a88800a,a88803a,a88806a,a88807a,a88808a,a88812a,a88813a,a88816a,a88819a,a88820a,a88821a,a88824a,a88827a,a88828a,a88831a,a88834a,a88835a,a88836a,a88840a,a88841a,a88844a,a88847a,a88848a,a88849a,a88852a,a88855a,a88856a,a88859a,a88862a,a88863a,a88864a,a88868a,a88869a,a88872a,a88875a,a88876a,a88877a,a88880a,a88883a,a88884a,a88887a,a88890a,a88891a,a88892a,a88896a,a88897a,a88900a,a88903a,a88904a,a88905a,a88908a,a88911a,a88912a,a88915a,a88918a,a88919a,a88920a,a88924a,a88925a,a88928a,a88931a,a88932a,a88933a,a88936a,a88939a,a88940a,a88943a,a88946a,a88947a,a88948a,a88952a,a88953a,a88956a,a88959a,a88960a,a88961a,a88964a,a88967a,a88968a,a88971a,a88974a,a88975a,a88976a,a88980a,a88981a,a88984a,a88987a,a88988a,a88989a,a88992a,a88995a,a88996a,a88999a,a89002a,a89003a,a89004a,a89008a,a89009a,a89012a,a89015a,a89016a,a89017a,a89020a,a89023a,a89024a,a89027a,a89030a,a89031a,a89032a,a89036a,a89037a,a89040a,a89043a,a89044a,a89045a,a89048a,a89051a,a89052a,a89055a,a89058a,a89059a,a89060a,a89064a,a89065a,a89068a,a89071a,a89072a,a89073a,a89076a,a89079a,a89080a,a89083a,a89086a,a89087a,a89088a,a89092a,a89093a,a89096a,a89099a,a89100a,a89101a,a89104a,a89107a,a89108a,a89111a,a89114a,a89115a,a89116a,a89120a,a89121a,a89124a,a89127a,a89128a,a89129a,a89132a,a89135a,a89136a,a89139a,a89142a,a89143a,a89144a,a89148a,a89149a,a89152a,a89155a,a89156a,a89157a,a89160a,a89163a,a89164a,a89167a,a89170a,a89171a,a89172a,a89176a,a89177a,a89180a,a89183a,a89184a,a89185a,a89188a,a89191a,a89192a,a89195a,a89198a,a89199a,a89200a,a89204a,a89205a,a89208a,a89211a,a89212a,a89213a,a89216a,a89219a,a89220a,a89223a,a89226a,a89227a,a89228a,a89232a,a89233a,a89236a,a89239a,a89240a,a89241a,a89244a,a89247a,a89248a,a89251a,a89254a,a89255a,a89256a,a89260a,a89261a,a89264a,a89267a,a89268a,a89269a,a89272a,a89275a,a89276a,a89279a,a89282a,a89283a,a89284a,a89288a,a89289a,a89292a,a89295a,a89296a,a89297a,a89300a,a89303a,a89304a,a89307a,a89310a,a89311a,a89312a,a89316a,a89317a,a89320a,a89323a,a89324a,a89325a,a89328a,a89331a,a89332a,a89335a,a89338a,a89339a,a89340a,a89344a,a89345a,a89348a,a89351a,a89352a,a89353a,a89356a,a89359a,a89360a,a89363a,a89366a,a89367a,a89368a,a89372a,a89373a,a89376a,a89379a,a89380a,a89381a,a89384a,a89387a,a89388a,a89391a,a89394a,a89395a,a89396a,a89400a,a89401a,a89404a,a89407a,a89408a,a89409a,a89412a,a89415a,a89416a,a89419a,a89422a,a89423a,a89424a,a89428a,a89429a,a89432a,a89435a,a89436a,a89437a,a89440a,a89443a,a89444a,a89447a,a89450a,a89451a,a89452a,a89456a,a89457a,a89460a,a89463a,a89464a,a89465a,a89468a,a89471a,a89472a,a89475a,a89478a,a89479a,a89480a,a89484a,a89485a,a89488a,a89491a,a89492a,a89493a,a89496a,a89499a,a89500a,a89503a,a89506a,a89507a,a89508a,a89512a,a89513a,a89516a,a89519a,a89520a,a89521a,a89524a,a89527a,a89528a,a89531a,a89534a,a89535a,a89536a,a89540a,a89541a,a89544a,a89547a,a89548a,a89549a,a89552a,a89555a,a89556a,a89559a,a89562a,a89563a,a89564a,a89568a,a89569a,a89572a,a89575a,a89576a,a89577a,a89580a,a89583a,a89584a,a89587a,a89590a,a89591a,a89592a,a89596a,a89597a,a89600a,a89603a,a89604a,a89605a,a89608a,a89611a,a89612a,a89615a,a89618a,a89619a,a89620a,a89624a,a89625a,a89628a,a89631a,a89632a,a89633a,a89636a,a89639a,a89640a,a89643a,a89646a,a89647a,a89648a,a89652a,a89653a,a89656a,a89659a,a89660a,a89661a,a89664a,a89667a,a89668a,a89671a,a89674a,a89675a,a89676a,a89680a,a89681a,a89684a,a89687a,a89688a,a89689a,a89692a,a89695a,a89696a,a89699a,a89702a,a89703a,a89704a,a89708a,a89709a,a89712a,a89715a,a89716a,a89717a,a89720a,a89723a,a89724a,a89727a,a89730a,a89731a,a89732a,a89736a,a89737a,a89740a,a89743a,a89744a,a89745a,a89748a,a89751a,a89752a,a89755a,a89758a,a89759a,a89760a,a89764a,a89765a,a89768a,a89771a,a89772a,a89773a,a89776a,a89779a,a89780a,a89783a,a89786a,a89787a,a89788a,a89792a,a89793a,a89796a,a89799a,a89800a,a89801a,a89804a,a89807a,a89808a,a89811a,a89814a,a89815a,a89816a,a89820a,a89821a,a89824a,a89827a,a89828a,a89829a,a89832a,a89835a,a89836a,a89839a,a89842a,a89843a,a89844a,a89848a,a89849a,a89852a,a89855a,a89856a,a89857a,a89860a,a89863a,a89864a,a89867a,a89870a,a89871a,a89872a,a89876a,a89877a,a89880a,a89883a,a89884a,a89885a,a89888a,a89891a,a89892a,a89895a,a89898a,a89899a,a89900a,a89904a,a89905a,a89908a,a89911a,a89912a,a89913a,a89916a,a89919a,a89920a,a89923a,a89926a,a89927a,a89928a,a89932a,a89933a,a89936a,a89939a,a89940a,a89941a,a89944a,a89947a,a89948a,a89951a,a89954a,a89955a,a89956a,a89960a,a89961a,a89964a,a89967a,a89968a,a89969a,a89972a,a89975a,a89976a,a89979a,a89982a,a89983a,a89984a,a89988a,a89989a,a89992a,a89995a,a89996a,a89997a,a90000a,a90003a,a90004a,a90007a,a90010a,a90011a,a90012a,a90016a,a90017a,a90020a,a90023a,a90024a,a90025a,a90028a,a90031a,a90032a,a90035a,a90038a,a90039a,a90040a,a90044a,a90045a,a90048a,a90051a,a90052a,a90053a,a90056a,a90059a,a90060a,a90063a,a90066a,a90067a,a90068a,a90072a,a90073a,a90076a,a90079a,a90080a,a90081a,a90084a,a90087a,a90088a,a90091a,a90094a,a90095a,a90096a,a90100a,a90101a,a90104a,a90107a,a90108a,a90109a,a90112a,a90115a,a90116a,a90119a,a90122a,a90123a,a90124a,a90128a,a90129a,a90132a,a90135a,a90136a,a90137a,a90140a,a90143a,a90144a,a90147a,a90150a,a90151a,a90152a,a90156a,a90157a,a90160a,a90163a,a90164a,a90165a,a90168a,a90171a,a90172a,a90175a,a90178a,a90179a,a90180a,a90184a,a90185a,a90188a,a90191a,a90192a,a90193a,a90196a,a90199a,a90200a,a90203a,a90206a,a90207a,a90208a,a90212a,a90213a,a90216a,a90219a,a90220a,a90221a,a90224a,a90227a,a90228a,a90231a,a90234a,a90235a,a90236a,a90240a,a90241a,a90244a,a90247a,a90248a,a90249a,a90252a,a90255a,a90256a,a90259a,a90262a,a90263a,a90264a,a90268a,a90269a,a90272a,a90275a,a90276a,a90277a,a90280a,a90283a,a90284a,a90287a,a90290a,a90291a,a90292a,a90296a,a90297a,a90300a,a90303a,a90304a,a90305a,a90308a,a90311a,a90312a,a90315a,a90318a,a90319a,a90320a,a90324a,a90325a,a90328a,a90331a,a90332a,a90333a,a90336a,a90339a,a90340a,a90343a,a90346a,a90347a,a90348a,a90352a,a90353a,a90356a,a90359a,a90360a,a90361a,a90364a,a90367a,a90368a,a90371a,a90374a,a90375a,a90376a,a90380a,a90381a,a90384a,a90387a,a90388a,a90389a,a90392a,a90395a,a90396a,a90399a,a90402a,a90403a,a90404a,a90408a,a90409a,a90412a,a90415a,a90416a,a90417a,a90420a,a90423a,a90424a,a90427a,a90430a,a90431a,a90432a,a90436a,a90437a,a90440a,a90443a,a90444a,a90445a,a90448a,a90451a,a90452a,a90455a,a90458a,a90459a,a90460a,a90464a,a90465a,a90468a,a90471a,a90472a,a90473a,a90476a,a90479a,a90480a,a90483a,a90486a,a90487a,a90488a,a90492a,a90493a,a90496a,a90499a,a90500a,a90501a,a90504a,a90507a,a90508a,a90511a,a90514a,a90515a,a90516a,a90520a,a90521a,a90524a,a90527a,a90528a,a90529a,a90532a,a90535a,a90536a,a90539a,a90542a,a90543a,a90544a,a90548a,a90549a,a90552a,a90555a,a90556a,a90557a,a90560a,a90563a,a90564a,a90567a,a90570a,a90571a,a90572a,a90576a,a90577a,a90580a,a90583a,a90584a,a90585a,a90588a,a90591a,a90592a,a90595a,a90598a,a90599a,a90600a,a90604a,a90605a,a90608a,a90611a,a90612a,a90613a,a90616a,a90619a,a90620a,a90623a,a90626a,a90627a,a90628a,a90632a,a90633a,a90636a,a90639a,a90640a,a90641a,a90644a,a90647a,a90648a,a90651a,a90654a,a90655a,a90656a,a90660a,a90661a,a90664a,a90667a,a90668a,a90669a,a90672a,a90675a,a90676a,a90679a,a90682a,a90683a,a90684a,a90688a,a90689a,a90692a,a90695a,a90696a,a90697a,a90700a,a90703a,a90704a,a90707a,a90710a,a90711a,a90712a,a90716a,a90717a,a90720a,a90723a,a90724a,a90725a,a90728a,a90731a,a90732a,a90735a,a90738a,a90739a,a90740a,a90744a,a90745a,a90748a,a90751a,a90752a,a90753a,a90756a,a90759a,a90760a,a90763a,a90766a,a90767a,a90768a,a90772a,a90773a,a90776a,a90779a,a90780a,a90781a,a90784a,a90787a,a90788a,a90791a,a90794a,a90795a,a90796a,a90800a,a90801a,a90804a,a90807a,a90808a,a90809a,a90812a,a90815a,a90816a,a90819a,a90822a,a90823a,a90824a,a90828a,a90829a,a90832a,a90835a,a90836a,a90837a,a90840a,a90843a,a90844a,a90847a,a90850a,a90851a,a90852a,a90856a,a90857a,a90860a,a90863a,a90864a,a90865a,a90868a,a90871a,a90872a,a90875a,a90878a,a90879a,a90880a,a90884a,a90885a,a90888a,a90891a,a90892a,a90893a,a90896a,a90899a,a90900a,a90903a,a90906a,a90907a,a90908a,a90912a,a90913a,a90916a,a90919a,a90920a,a90921a,a90924a,a90927a,a90928a,a90931a,a90934a,a90935a,a90936a,a90940a,a90941a,a90944a,a90947a,a90948a,a90949a,a90952a,a90955a,a90956a,a90959a,a90962a,a90963a,a90964a,a90968a,a90969a,a90972a,a90975a,a90976a,a90977a,a90980a,a90983a,a90984a,a90987a,a90990a,a90991a,a90992a,a90996a,a90997a,a91000a,a91003a,a91004a,a91005a,a91008a,a91011a,a91012a,a91015a,a91018a,a91019a,a91020a,a91024a,a91025a,a91028a,a91031a,a91032a,a91033a,a91036a,a91039a,a91040a,a91043a,a91046a,a91047a,a91048a,a91052a,a91053a,a91056a,a91059a,a91060a,a91061a,a91064a,a91067a,a91068a,a91071a,a91074a,a91075a,a91076a,a91080a,a91081a,a91084a,a91087a,a91088a,a91089a,a91092a,a91095a,a91096a,a91099a,a91102a,a91103a,a91104a,a91108a,a91109a,a91112a,a91115a,a91116a,a91117a,a91120a,a91123a,a91124a,a91127a,a91130a,a91131a,a91132a,a91136a,a91137a,a91140a,a91143a,a91144a,a91145a,a91148a,a91151a,a91152a,a91155a,a91158a,a91159a,a91160a,a91164a,a91165a,a91168a,a91171a,a91172a,a91173a,a91176a,a91179a,a91180a,a91183a,a91186a,a91187a,a91188a,a91192a,a91193a,a91196a,a91199a,a91200a,a91201a,a91204a,a91207a,a91208a,a91211a,a91214a,a91215a,a91216a,a91220a,a91221a,a91224a,a91227a,a91228a,a91229a,a91232a,a91235a,a91236a,a91239a,a91242a,a91243a,a91244a,a91248a,a91249a,a91252a,a91255a,a91256a,a91257a,a91260a,a91263a,a91264a,a91267a,a91270a,a91271a,a91272a,a91276a,a91277a,a91280a,a91283a,a91284a,a91285a,a91288a,a91291a,a91292a,a91295a,a91298a,a91299a,a91300a,a91304a,a91305a,a91308a,a91311a,a91312a,a91313a,a91316a,a91319a,a91320a,a91323a,a91326a,a91327a,a91328a,a91332a,a91333a,a91336a,a91339a,a91340a,a91341a,a91344a,a91347a,a91348a,a91351a,a91354a,a91355a,a91356a,a91360a,a91361a,a91364a,a91367a,a91368a,a91369a,a91372a,a91375a,a91376a,a91379a,a91382a,a91383a,a91384a,a91388a,a91389a,a91392a,a91395a,a91396a,a91397a,a91400a,a91403a,a91404a,a91407a,a91410a,a91411a,a91412a,a91416a,a91417a,a91420a,a91423a,a91424a,a91425a,a91428a,a91431a,a91432a,a91435a,a91438a,a91439a,a91440a,a91444a,a91445a,a91448a,a91451a,a91452a,a91453a,a91456a,a91459a,a91460a,a91463a,a91466a,a91467a,a91468a,a91472a,a91473a,a91476a,a91479a,a91480a,a91481a,a91484a,a91487a,a91488a,a91491a,a91494a,a91495a,a91496a,a91500a,a91501a,a91504a,a91507a,a91508a,a91509a,a91512a,a91515a,a91516a,a91519a,a91522a,a91523a,a91524a,a91528a,a91529a,a91532a,a91535a,a91536a,a91537a,a91540a,a91543a,a91544a,a91547a,a91550a,a91551a,a91552a,a91556a,a91557a,a91560a,a91563a,a91564a,a91565a,a91568a,a91571a,a91572a,a91575a,a91578a,a91579a,a91580a,a91584a,a91585a,a91588a,a91591a,a91592a,a91593a,a91596a,a91599a,a91600a,a91603a,a91606a,a91607a,a91608a,a91612a,a91613a,a91616a,a91619a,a91620a,a91621a,a91624a,a91627a,a91628a,a91631a,a91634a,a91635a,a91636a,a91640a,a91641a,a91644a,a91647a,a91648a,a91649a,a91652a,a91655a,a91656a,a91659a,a91662a,a91663a,a91664a,a91668a,a91669a,a91672a,a91675a,a91676a,a91677a,a91680a,a91683a,a91684a,a91687a,a91690a,a91691a,a91692a,a91696a,a91697a,a91700a,a91703a,a91704a,a91705a,a91708a,a91711a,a91712a,a91715a,a91718a,a91719a,a91720a,a91724a,a91725a,a91728a,a91731a,a91732a,a91733a,a91736a,a91739a,a91740a,a91743a,a91746a,a91747a,a91748a,a91752a,a91753a,a91756a,a91759a,a91760a,a91761a,a91764a,a91767a,a91768a,a91771a,a91774a,a91775a,a91776a,a91780a,a91781a,a91784a,a91787a,a91788a,a91789a,a91792a,a91795a,a91796a,a91799a,a91802a,a91803a,a91804a,a91808a,a91809a,a91812a,a91815a,a91816a,a91817a,a91820a,a91823a,a91824a,a91827a,a91830a,a91831a,a91832a,a91836a,a91837a,a91840a,a91843a,a91844a,a91845a,a91848a,a91851a,a91852a,a91855a,a91858a,a91859a,a91860a,a91864a,a91865a,a91868a,a91871a,a91872a,a91873a,a91876a,a91879a,a91880a,a91883a,a91886a,a91887a,a91888a,a91892a,a91893a,a91896a,a91899a,a91900a,a91901a,a91904a,a91907a,a91908a,a91911a,a91914a,a91915a,a91916a,a91920a,a91921a,a91924a,a91927a,a91928a,a91929a,a91932a,a91935a,a91936a,a91939a,a91942a,a91943a,a91944a,a91948a,a91949a,a91952a,a91955a,a91956a,a91957a,a91960a,a91963a,a91964a,a91967a,a91970a,a91971a,a91972a,a91976a,a91977a,a91980a,a91983a,a91984a,a91985a,a91988a,a91991a,a91992a,a91995a,a91998a,a91999a,a92000a,a92004a,a92005a,a92008a,a92011a,a92012a,a92013a,a92016a,a92019a,a92020a,a92023a,a92026a,a92027a,a92028a,a92032a,a92033a,a92036a,a92039a,a92040a,a92041a,a92044a,a92047a,a92048a,a92051a,a92054a,a92055a,a92056a,a92060a,a92061a,a92064a,a92067a,a92068a,a92069a,a92072a,a92075a,a92076a,a92079a,a92082a,a92083a,a92084a,a92088a,a92089a,a92092a,a92095a,a92096a,a92097a,a92100a,a92103a,a92104a,a92107a,a92110a,a92111a,a92112a,a92116a,a92117a,a92120a,a92123a,a92124a,a92125a,a92128a,a92131a,a92132a,a92135a,a92138a,a92139a,a92140a,a92144a,a92145a,a92148a,a92151a,a92152a,a92153a,a92156a,a92159a,a92160a,a92163a,a92166a,a92167a,a92168a,a92172a,a92173a,a92176a,a92179a,a92180a,a92181a,a92184a,a92187a,a92188a,a92191a,a92194a,a92195a,a92196a,a92200a,a92201a,a92204a,a92207a,a92208a,a92209a,a92212a,a92215a,a92216a,a92219a,a92222a,a92223a,a92224a,a92228a,a92229a,a92232a,a92235a,a92236a,a92237a,a92240a,a92243a,a92244a,a92247a,a92250a,a92251a,a92252a,a92256a,a92257a,a92260a,a92263a,a92264a,a92265a,a92268a,a92271a,a92272a,a92275a,a92278a,a92279a,a92280a,a92284a,a92285a,a92288a,a92291a,a92292a,a92293a,a92296a,a92299a,a92300a,a92303a,a92306a,a92307a,a92308a,a92312a,a92313a,a92316a,a92319a,a92320a,a92321a,a92324a,a92327a,a92328a,a92331a,a92334a,a92335a,a92336a,a92340a,a92341a,a92344a,a92347a,a92348a,a92349a,a92352a,a92355a,a92356a,a92359a,a92362a,a92363a,a92364a,a92368a,a92369a,a92372a,a92375a,a92376a,a92377a,a92380a,a92383a,a92384a,a92387a,a92390a,a92391a,a92392a,a92396a,a92397a,a92400a,a92403a,a92404a,a92405a,a92408a,a92411a,a92412a,a92415a,a92418a,a92419a,a92420a,a92424a,a92425a,a92428a,a92431a,a92432a,a92433a,a92436a,a92439a,a92440a,a92443a,a92446a,a92447a,a92448a,a92452a,a92453a,a92456a,a92459a,a92460a,a92461a,a92464a,a92467a,a92468a,a92471a,a92474a,a92475a,a92476a,a92480a,a92481a,a92484a,a92487a,a92488a,a92489a,a92492a,a92495a,a92496a,a92499a,a92502a,a92503a,a92504a,a92508a,a92509a,a92512a,a92515a,a92516a,a92517a,a92520a,a92523a,a92524a,a92527a,a92530a,a92531a,a92532a,a92536a,a92537a,a92540a,a92543a,a92544a,a92545a,a92548a,a92551a,a92552a,a92555a,a92558a,a92559a,a92560a,a92564a,a92565a,a92568a,a92571a,a92572a,a92573a,a92576a,a92579a,a92580a,a92583a,a92586a,a92587a,a92588a,a92592a,a92593a,a92596a,a92599a,a92600a,a92601a,a92604a,a92607a,a92608a,a92611a,a92614a,a92615a,a92616a,a92620a,a92621a,a92624a,a92627a,a92628a,a92629a,a92632a,a92635a,a92636a,a92639a,a92642a,a92643a,a92644a,a92648a,a92649a,a92652a,a92655a,a92656a,a92657a,a92660a,a92663a,a92664a,a92667a,a92670a,a92671a,a92672a,a92676a,a92677a,a92680a,a92683a,a92684a,a92685a,a92688a,a92691a,a92692a,a92695a,a92698a,a92699a,a92700a,a92704a,a92705a,a92708a,a92711a,a92712a,a92713a,a92716a,a92719a,a92720a,a92723a,a92726a,a92727a,a92728a,a92732a,a92733a,a92736a,a92739a,a92740a,a92741a,a92744a,a92747a,a92748a,a92751a,a92754a,a92755a,a92756a,a92760a,a92761a,a92764a,a92767a,a92768a,a92769a,a92772a,a92775a,a92776a,a92779a,a92782a,a92783a,a92784a,a92788a,a92789a,a92792a,a92795a,a92796a,a92797a,a92800a,a92803a,a92804a,a92807a,a92810a,a92811a,a92812a,a92816a,a92817a,a92820a,a92823a,a92824a,a92825a,a92828a,a92831a,a92832a,a92835a,a92838a,a92839a,a92840a,a92844a,a92845a,a92848a,a92851a,a92852a,a92853a,a92856a,a92859a,a92860a,a92863a,a92866a,a92867a,a92868a,a92871a,a92874a,a92875a,a92878a,a92881a,a92882a,a92883a,a92886a,a92889a,a92890a,a92893a,a92896a,a92897a,a92898a,a92901a,a92904a,a92905a,a92908a,a92911a,a92912a,a92913a,a92916a,a92919a,a92920a,a92923a,a92926a,a92927a,a92928a,a92931a,a92934a,a92935a,a92938a,a92941a,a92942a,a92943a,a92946a,a92949a,a92950a,a92953a,a92956a,a92957a,a92958a,a92961a,a92964a,a92965a,a92968a,a92971a,a92972a,a92973a,a92976a,a92979a,a92980a,a92983a,a92986a,a92987a,a92988a,a92991a,a92994a,a92995a,a92998a,a93001a,a93002a,a93003a,a93006a,a93009a,a93010a,a93013a,a93016a,a93017a,a93018a,a93021a,a93024a,a93025a,a93028a,a93031a,a93032a,a93033a,a93036a,a93039a,a93040a,a93043a,a93046a,a93047a,a93048a,a93051a,a93054a,a93055a,a93058a,a93061a,a93062a,a93063a,a93066a,a93069a,a93070a,a93073a,a93076a,a93077a,a93078a,a93081a,a93084a,a93085a,a93088a,a93091a,a93092a,a93093a,a93096a,a93099a,a93100a,a93103a,a93106a,a93107a,a93108a,a93111a,a93114a,a93115a,a93118a,a93121a,a93122a,a93123a,a93126a,a93129a,a93130a,a93133a,a93136a,a93137a,a93138a,a93141a,a93144a,a93145a,a93148a,a93151a,a93152a,a93153a,a93156a,a93159a,a93160a,a93163a,a93166a,a93167a,a93168a,a93171a,a93174a,a93175a,a93178a,a93181a,a93182a,a93183a,a93186a,a93189a,a93190a,a93193a,a93196a,a93197a,a93198a,a93201a,a93204a,a93205a,a93208a,a93211a,a93212a,a93213a,a93216a,a93219a,a93220a,a93223a,a93226a,a93227a,a93228a,a93231a,a93234a,a93235a,a93238a,a93241a,a93242a,a93243a,a93246a,a93249a,a93250a,a93253a,a93256a,a93257a,a93258a,a93261a,a93264a,a93265a,a93268a,a93271a,a93272a,a93273a,a93276a,a93279a,a93280a,a93283a,a93286a,a93287a,a93288a,a93291a,a93294a,a93295a,a93298a,a93301a,a93302a,a93303a,a93306a,a93309a,a93310a,a93313a,a93316a,a93317a,a93318a,a93321a,a93324a,a93325a,a93328a,a93331a,a93332a,a93333a,a93336a,a93339a,a93340a,a93343a,a93346a,a93347a,a93348a,a93351a,a93354a,a93355a,a93358a,a93361a,a93362a,a93363a,a93366a,a93369a,a93370a,a93373a,a93376a,a93377a,a93378a,a93381a,a93384a,a93385a,a93388a,a93391a,a93392a,a93393a,a93396a,a93399a,a93400a,a93403a,a93406a,a93407a,a93408a,a93411a,a93414a,a93415a,a93418a,a93421a,a93422a,a93423a,a93426a,a93429a,a93430a,a93433a,a93436a,a93437a,a93438a,a93441a,a93444a,a93445a,a93448a,a93451a,a93452a,a93453a,a93456a,a93459a,a93460a,a93463a,a93466a,a93467a,a93468a,a93471a,a93474a,a93475a,a93478a,a93481a,a93482a,a93483a,a93486a,a93489a,a93490a,a93493a,a93496a,a93497a,a93498a,a93501a,a93504a,a93505a,a93508a,a93511a,a93512a,a93513a,a93516a,a93519a,a93520a,a93523a,a93526a,a93527a,a93528a,a93531a,a93534a,a93535a,a93538a,a93541a,a93542a,a93543a,a93546a,a93549a,a93550a,a93553a,a93556a,a93557a,a93558a,a93561a,a93564a,a93565a,a93568a,a93571a,a93572a,a93573a,a93576a,a93579a,a93580a,a93583a,a93586a,a93587a,a93588a,a93591a,a93594a,a93595a,a93598a,a93601a,a93602a,a93603a,a93606a,a93609a,a93610a,a93613a,a93616a,a93617a,a93618a,a93621a,a93624a,a93625a,a93628a,a93631a,a93632a,a93633a,a93636a,a93639a,a93640a,a93643a,a93646a,a93647a,a93648a,a93651a,a93654a,a93655a,a93658a,a93661a,a93662a,a93663a,a93666a,a93669a,a93670a,a93673a,a93676a,a93677a,a93678a,a93681a,a93684a,a93685a,a93688a,a93691a,a93692a,a93693a,a93696a,a93699a,a93700a,a93703a,a93706a,a93707a,a93708a,a93711a,a93714a,a93715a,a93718a,a93721a,a93722a,a93723a,a93726a,a93729a,a93730a,a93733a,a93736a,a93737a,a93738a,a93741a,a93744a,a93745a,a93748a,a93751a,a93752a,a93753a,a93756a,a93759a,a93760a,a93763a,a93766a,a93767a,a93768a,a93771a,a93774a,a93775a,a93778a,a93781a,a93782a,a93783a,a93786a,a93789a,a93790a,a93793a,a93796a,a93797a,a93798a,a93801a,a93804a,a93805a,a93808a,a93811a,a93812a,a93813a,a93816a,a93819a,a93820a,a93823a,a93826a,a93827a,a93828a,a93831a,a93834a,a93835a,a93838a,a93841a,a93842a,a93843a,a93846a,a93849a,a93850a,a93853a,a93856a,a93857a,a93858a,a93861a,a93864a,a93865a,a93868a,a93871a,a93872a,a93873a,a93876a,a93879a,a93880a,a93883a,a93886a,a93887a,a93888a,a93891a,a93894a,a93895a,a93898a,a93901a,a93902a,a93903a,a93906a,a93909a,a93910a,a93913a,a93916a,a93917a,a93918a,a93921a,a93924a,a93925a,a93928a,a93931a,a93932a,a93933a,a93936a,a93939a,a93940a,a93943a,a93946a,a93947a,a93948a,a93951a,a93954a,a93955a,a93958a,a93961a,a93962a,a93963a,a93966a,a93969a,a93970a,a93973a,a93976a,a93977a,a93978a,a93981a,a93984a,a93985a,a93988a,a93991a,a93992a,a93993a,a93996a,a93999a,a94000a,a94003a,a94006a,a94007a,a94008a,a94011a,a94014a,a94015a,a94018a,a94021a,a94022a,a94023a,a94026a,a94029a,a94030a,a94033a,a94036a,a94037a,a94038a,a94041a,a94044a,a94045a,a94048a,a94051a,a94052a,a94053a,a94056a,a94059a,a94060a,a94063a,a94066a,a94067a,a94068a,a94071a,a94074a,a94075a,a94078a,a94081a,a94082a,a94083a,a94086a,a94089a,a94090a,a94093a,a94096a,a94097a,a94098a,a94101a,a94104a,a94105a,a94108a,a94111a,a94112a,a94113a,a94116a,a94119a,a94120a,a94123a,a94126a,a94127a,a94128a,a94131a,a94134a,a94135a,a94138a,a94141a,a94142a,a94143a,a94146a,a94149a,a94150a,a94153a,a94156a,a94157a,a94158a,a94161a,a94164a,a94165a,a94168a,a94171a,a94172a,a94173a,a94176a,a94179a,a94180a,a94183a,a94186a,a94187a,a94188a,a94191a,a94194a,a94195a,a94198a,a94201a,a94202a,a94203a,a94206a,a94209a,a94210a,a94213a,a94216a,a94217a,a94218a,a94221a,a94224a,a94225a,a94228a,a94231a,a94232a,a94233a,a94236a,a94239a,a94240a,a94243a,a94246a,a94247a,a94248a,a94251a,a94254a,a94255a,a94258a,a94261a,a94262a,a94263a,a94266a,a94269a,a94270a,a94273a,a94276a,a94277a,a94278a,a94281a,a94284a,a94285a,a94288a,a94291a,a94292a,a94293a,a94296a,a94299a,a94300a,a94303a,a94306a,a94307a,a94308a,a94311a,a94314a,a94315a,a94318a,a94321a,a94322a,a94323a,a94326a,a94329a,a94330a,a94333a,a94336a,a94337a,a94338a,a94341a,a94344a,a94345a,a94348a,a94351a,a94352a,a94353a,a94356a,a94359a,a94360a,a94363a,a94366a,a94367a,a94368a,a94371a,a94374a,a94375a,a94378a,a94381a,a94382a,a94383a,a94386a,a94389a,a94390a,a94393a,a94396a,a94397a,a94398a,a94401a,a94404a,a94405a,a94408a,a94411a,a94412a,a94413a,a94416a,a94419a,a94420a,a94423a,a94426a,a94427a,a94428a,a94431a,a94434a,a94435a,a94438a,a94441a,a94442a,a94443a,a94446a,a94449a,a94450a,a94453a,a94456a,a94457a,a94458a,a94461a,a94464a,a94465a,a94468a,a94471a,a94472a,a94473a,a94476a,a94479a,a94480a,a94483a,a94486a,a94487a,a94488a,a94491a,a94494a,a94495a,a94498a,a94501a,a94502a,a94503a,a94506a,a94509a,a94510a,a94513a,a94516a,a94517a,a94518a,a94521a,a94524a,a94525a,a94528a,a94531a,a94532a,a94533a,a94536a,a94539a,a94540a,a94543a,a94546a,a94547a,a94548a,a94551a,a94554a,a94555a,a94558a,a94561a,a94562a,a94563a,a94566a,a94569a,a94570a,a94573a,a94576a,a94577a,a94578a,a94581a,a94584a,a94585a,a94588a,a94591a,a94592a,a94593a,a94596a,a94599a,a94600a,a94603a,a94606a,a94607a,a94608a,a94611a,a94614a,a94615a,a94618a,a94621a,a94622a,a94623a,a94626a,a94629a,a94630a,a94633a,a94636a,a94637a,a94638a,a94641a,a94644a,a94645a,a94648a,a94651a,a94652a,a94653a,a94656a,a94659a,a94660a,a94663a,a94666a,a94667a,a94668a,a94671a,a94674a,a94675a,a94678a,a94681a,a94682a,a94683a,a94686a,a94689a,a94690a,a94693a,a94696a,a94697a,a94698a,a94701a,a94704a,a94705a,a94708a,a94711a,a94712a,a94713a,a94716a,a94719a,a94720a,a94723a,a94726a,a94727a,a94728a,a94731a,a94734a,a94735a,a94738a,a94741a,a94742a,a94743a,a94746a,a94749a,a94750a,a94753a,a94756a,a94757a,a94758a,a94761a,a94764a,a94765a,a94768a,a94771a,a94772a,a94773a,a94776a,a94779a,a94780a,a94783a,a94786a,a94787a,a94788a,a94791a,a94794a,a94795a,a94798a,a94801a,a94802a,a94803a,a94806a,a94809a,a94810a,a94813a,a94816a,a94817a,a94818a,a94821a,a94824a,a94825a,a94828a,a94831a,a94832a,a94833a,a94836a,a94839a,a94840a,a94843a,a94846a,a94847a,a94848a,a94851a,a94854a,a94855a,a94858a,a94861a,a94862a,a94863a,a94866a,a94869a,a94870a,a94873a,a94876a,a94877a,a94878a,a94881a,a94884a,a94885a,a94888a,a94891a,a94892a,a94893a,a94896a,a94899a,a94900a,a94903a,a94906a,a94907a,a94908a,a94911a,a94914a,a94915a,a94918a,a94921a,a94922a,a94923a,a94926a,a94929a,a94930a,a94933a,a94936a,a94937a,a94938a,a94941a,a94944a,a94945a,a94948a,a94951a,a94952a,a94953a,a94956a,a94959a,a94960a,a94963a,a94966a,a94967a,a94968a,a94971a,a94974a,a94975a,a94978a,a94981a,a94982a,a94983a,a94986a,a94989a,a94990a,a94993a,a94996a,a94997a,a94998a,a95001a,a95004a,a95005a,a95008a,a95011a,a95012a,a95013a,a95016a,a95019a,a95020a,a95023a,a95026a,a95027a,a95028a,a95031a,a95034a,a95035a,a95038a,a95041a,a95042a,a95043a,a95046a,a95049a,a95050a,a95053a,a95056a,a95057a,a95058a,a95061a,a95064a,a95065a,a95068a,a95071a,a95072a,a95073a,a95076a,a95079a,a95080a,a95083a,a95086a,a95087a,a95088a,a95091a,a95094a,a95095a,a95098a,a95101a,a95102a,a95103a,a95106a,a95109a,a95110a,a95113a,a95116a,a95117a,a95118a,a95121a,a95124a,a95125a,a95128a,a95131a,a95132a,a95133a,a95136a,a95139a,a95140a,a95143a,a95146a,a95147a,a95148a,a95151a,a95154a,a95155a,a95158a,a95161a,a95162a,a95163a,a95166a,a95169a,a95170a,a95173a,a95176a,a95177a,a95178a,a95181a,a95184a,a95185a,a95188a,a95191a,a95192a,a95193a,a95196a,a95199a,a95200a,a95203a,a95206a,a95207a,a95208a,a95211a,a95214a,a95215a,a95218a,a95221a,a95222a,a95223a,a95226a,a95229a,a95230a,a95233a,a95236a,a95237a,a95238a,a95241a,a95244a,a95245a,a95248a,a95251a,a95252a,a95253a,a95256a,a95259a,a95260a,a95263a,a95266a,a95267a,a95268a,a95271a,a95274a,a95275a,a95278a,a95281a,a95282a,a95283a,a95286a,a95289a,a95290a,a95293a,a95296a,a95297a,a95298a,a95301a,a95304a,a95305a,a95308a,a95311a,a95312a,a95313a,a95316a,a95319a,a95320a,a95323a,a95326a,a95327a,a95328a,a95331a,a95334a,a95335a,a95338a,a95341a,a95342a,a95343a,a95346a,a95349a,a95350a,a95353a,a95356a,a95357a,a95358a,a95361a,a95364a,a95365a,a95368a,a95371a,a95372a,a95373a,a95376a,a95379a,a95380a,a95383a,a95386a,a95387a,a95388a,a95391a,a95394a,a95395a,a95398a,a95401a,a95402a,a95403a,a95406a,a95409a,a95410a,a95413a,a95416a,a95417a,a95418a,a95421a,a95424a,a95425a,a95428a,a95431a,a95432a,a95433a,a95436a,a95439a,a95440a,a95443a,a95446a,a95447a,a95448a,a95451a,a95454a,a95455a,a95458a,a95461a,a95462a,a95463a,a95466a,a95469a,a95470a,a95473a,a95476a,a95477a,a95478a,a95481a,a95484a,a95485a,a95488a,a95491a,a95492a,a95493a,a95496a,a95499a,a95500a,a95503a,a95506a,a95507a,a95508a,a95511a,a95514a,a95515a,a95518a,a95521a,a95522a,a95523a,a95526a,a95529a,a95530a,a95533a,a95536a,a95537a,a95538a,a95541a,a95544a,a95545a,a95548a,a95551a,a95552a,a95553a,a95556a,a95559a,a95560a,a95563a,a95566a,a95567a,a95568a,a95571a,a95574a,a95575a,a95578a,a95581a,a95582a,a95583a,a95586a,a95589a,a95590a,a95593a,a95596a,a95597a,a95598a,a95601a,a95604a,a95605a,a95608a,a95611a,a95612a,a95613a,a95616a,a95619a,a95620a,a95623a,a95626a,a95627a,a95628a,a95631a,a95634a,a95635a,a95638a,a95641a,a95642a,a95643a,a95646a,a95649a,a95650a,a95653a,a95656a,a95657a,a95658a,a95661a,a95664a,a95665a,a95668a,a95671a,a95672a,a95673a,a95676a,a95679a,a95680a,a95683a,a95686a,a95687a,a95688a,a95691a,a95694a,a95695a,a95698a,a95701a,a95702a,a95703a,a95706a,a95709a,a95710a,a95713a,a95716a,a95717a,a95718a,a95721a,a95724a,a95725a,a95728a,a95731a,a95732a,a95733a,a95736a,a95739a,a95740a,a95743a,a95746a,a95747a,a95748a,a95751a,a95754a,a95755a,a95758a,a95761a,a95762a,a95763a,a95766a,a95769a,a95770a,a95773a,a95776a,a95777a,a95778a,a95781a,a95784a,a95785a,a95788a,a95791a,a95792a,a95793a,a95796a,a95799a,a95800a,a95803a,a95806a,a95807a,a95808a,a95811a,a95814a,a95815a,a95818a,a95821a,a95822a,a95823a,a95826a,a95829a,a95830a,a95833a,a95836a,a95837a,a95838a,a95841a,a95844a,a95845a,a95848a,a95851a,a95852a,a95853a,a95856a,a95859a,a95860a,a95863a,a95866a,a95867a,a95868a,a95871a,a95874a,a95875a,a95878a,a95881a,a95882a,a95883a,a95886a,a95889a,a95890a,a95893a,a95896a,a95897a,a95898a,a95901a,a95904a,a95905a,a95908a,a95911a,a95912a,a95913a,a95916a,a95919a,a95920a,a95923a,a95926a,a95927a,a95928a,a95931a,a95934a,a95935a,a95938a,a95941a,a95942a,a95943a,a95946a,a95949a,a95950a,a95953a,a95956a,a95957a,a95958a,a95961a,a95964a,a95965a,a95968a,a95971a,a95972a,a95973a,a95976a,a95979a,a95980a,a95983a,a95986a,a95987a,a95988a,a95991a,a95994a,a95995a,a95998a,a96001a,a96002a,a96003a,a96006a,a96009a,a96010a,a96013a,a96016a,a96017a,a96018a,a96021a,a96024a,a96025a,a96028a,a96031a,a96032a,a96033a,a96036a,a96039a,a96040a,a96043a,a96046a,a96047a,a96048a,a96051a,a96054a,a96055a,a96058a,a96061a,a96062a,a96063a,a96066a,a96069a,a96070a,a96073a,a96076a,a96077a,a96078a,a96081a,a96084a,a96085a,a96088a,a96091a,a96092a,a96093a,a96096a,a96099a,a96100a,a96103a,a96106a,a96107a,a96108a,a96111a,a96114a,a96115a,a96118a,a96121a,a96122a,a96123a,a96126a,a96129a,a96130a,a96133a,a96136a,a96137a,a96138a,a96141a,a96144a,a96145a,a96148a,a96151a,a96152a,a96153a,a96156a,a96159a,a96160a,a96163a,a96166a,a96167a,a96168a,a96171a,a96174a,a96175a,a96178a,a96181a,a96182a,a96183a,a96186a,a96189a,a96190a,a96193a,a96196a,a96197a,a96198a,a96201a,a96204a,a96205a,a96208a,a96211a,a96212a,a96213a,a96216a,a96219a,a96220a,a96223a,a96226a,a96227a,a96228a,a96231a,a96234a,a96235a,a96238a,a96241a,a96242a,a96243a,a96246a,a96249a,a96250a,a96253a,a96256a,a96257a,a96258a,a96261a,a96264a,a96265a,a96268a,a96271a,a96272a,a96273a,a96276a,a96279a,a96280a,a96283a,a96286a,a96287a,a96288a,a96291a,a96294a,a96295a,a96298a,a96301a,a96302a,a96303a,a96306a,a96309a,a96310a,a96313a,a96316a,a96317a,a96318a,a96321a,a96324a,a96325a,a96328a,a96331a,a96332a,a96333a,a96336a,a96339a,a96340a,a96343a,a96346a,a96347a,a96348a,a96351a,a96354a,a96355a,a96358a,a96361a,a96362a,a96363a,a96366a,a96369a,a96370a,a96373a,a96376a,a96377a,a96378a,a96381a,a96384a,a96385a,a96388a,a96391a,a96392a,a96393a,a96396a,a96399a,a96400a,a96403a,a96406a,a96407a,a96408a,a96411a,a96414a,a96415a,a96418a,a96421a,a96422a,a96423a,a96426a,a96429a,a96430a,a96433a,a96436a,a96437a,a96438a,a96441a,a96444a,a96445a,a96448a,a96451a,a96452a,a96453a,a96456a,a96459a,a96460a,a96463a,a96466a,a96467a,a96468a,a96471a,a96474a,a96475a,a96478a,a96481a,a96482a,a96483a,a96486a,a96489a,a96490a,a96493a,a96496a,a96497a,a96498a,a96501a,a96504a,a96505a,a96508a,a96511a,a96512a,a96513a,a96516a,a96519a,a96520a,a96523a,a96526a,a96527a,a96528a,a96531a,a96534a,a96535a,a96538a,a96541a,a96542a,a96543a,a96546a,a96549a,a96550a,a96553a,a96556a,a96557a,a96558a,a96561a,a96564a,a96565a,a96568a,a96571a,a96572a,a96573a,a96576a,a96579a,a96580a,a96583a,a96586a,a96587a,a96588a,a96591a,a96594a,a96595a,a96598a,a96601a,a96602a,a96603a,a96606a,a96609a,a96610a,a96613a,a96616a,a96617a,a96618a,a96621a,a96624a,a96625a,a96628a,a96631a,a96632a,a96633a,a96636a,a96639a,a96640a,a96643a,a96646a,a96647a,a96648a,a96651a,a96654a,a96655a,a96658a,a96661a,a96662a,a96663a,a96666a,a96669a,a96670a,a96673a,a96676a,a96677a,a96678a,a96681a,a96684a,a96685a,a96688a,a96691a,a96692a,a96693a,a96696a,a96699a,a96700a,a96703a,a96706a,a96707a,a96708a,a96711a,a96714a,a96715a,a96718a,a96721a,a96722a,a96723a,a96726a,a96729a,a96730a,a96733a,a96736a,a96737a,a96738a,a96741a,a96744a,a96745a,a96748a,a96751a,a96752a,a96753a,a96756a,a96759a,a96760a,a96763a,a96766a,a96767a,a96768a,a96771a,a96774a,a96775a,a96778a,a96781a,a96782a,a96783a,a96786a,a96789a,a96790a,a96793a,a96796a,a96797a,a96798a,a96801a,a96804a,a96805a,a96808a,a96811a,a96812a,a96813a,a96816a,a96819a,a96820a,a96823a,a96826a,a96827a,a96828a,a96831a,a96834a,a96835a,a96838a,a96841a,a96842a,a96843a,a96846a,a96849a,a96850a,a96853a,a96856a,a96857a,a96858a,a96861a,a96864a,a96865a,a96868a,a96871a,a96872a,a96873a,a96876a,a96879a,a96880a,a96883a,a96886a,a96887a,a96888a,a96891a,a96894a,a96895a,a96898a,a96901a,a96902a,a96903a,a96906a,a96909a,a96910a,a96913a,a96916a,a96917a,a96918a,a96921a,a96924a,a96925a,a96928a,a96931a,a96932a,a96933a,a96936a,a96939a,a96940a,a96943a,a96946a,a96947a,a96948a,a96951a,a96954a,a96955a,a96958a,a96961a,a96962a,a96963a,a96966a,a96969a,a96970a,a96973a,a96976a,a96977a,a96978a,a96981a,a96984a,a96985a,a96988a,a96991a,a96992a,a96993a,a96996a,a96999a,a97000a,a97003a,a97006a,a97007a,a97008a,a97011a,a97014a,a97015a,a97018a,a97021a,a97022a,a97023a,a97026a,a97029a,a97030a,a97033a,a97036a,a97037a,a97038a,a97041a,a97044a,a97045a,a97048a,a97051a,a97052a,a97053a,a97056a,a97059a,a97060a,a97063a,a97066a,a97067a,a97068a,a97071a,a97074a,a97075a,a97078a,a97081a,a97082a,a97083a,a97086a,a97089a,a97090a,a97093a,a97096a,a97097a,a97098a,a97101a,a97104a,a97105a,a97108a,a97111a,a97112a,a97113a,a97116a,a97119a,a97120a,a97123a,a97126a,a97127a,a97128a,a97131a,a97134a,a97135a,a97138a,a97141a,a97142a,a97143a,a97146a,a97149a,a97150a,a97153a,a97156a,a97157a,a97158a,a97161a,a97164a,a97165a,a97168a,a97171a,a97172a,a97173a,a97176a,a97179a,a97180a,a97183a,a97186a,a97187a,a97188a,a97191a,a97194a,a97195a,a97198a,a97201a,a97202a,a97203a,a97206a,a97209a,a97210a,a97213a,a97216a,a97217a,a97218a,a97221a,a97224a,a97225a,a97228a,a97231a,a97232a,a97233a,a97236a,a97239a,a97240a,a97243a,a97246a,a97247a,a97248a,a97251a,a97254a,a97255a,a97258a,a97261a,a97262a,a97263a,a97266a,a97269a,a97270a,a97273a,a97276a,a97277a,a97278a,a97281a,a97284a,a97285a,a97288a,a97291a,a97292a,a97293a,a97296a,a97299a,a97300a,a97303a,a97306a,a97307a,a97308a,a97311a,a97314a,a97315a,a97318a,a97321a,a97322a,a97323a,a97326a,a97329a,a97330a,a97333a,a97336a,a97337a,a97338a,a97341a,a97344a,a97345a,a97348a,a97351a,a97352a,a97353a,a97356a,a97359a,a97360a,a97363a,a97366a,a97367a,a97368a,a97371a,a97374a,a97375a,a97378a,a97381a,a97382a,a97383a,a97386a,a97389a,a97390a,a97393a,a97396a,a97397a,a97398a,a97401a,a97404a,a97405a,a97408a,a97411a,a97412a,a97413a,a97416a,a97419a,a97420a,a97423a,a97426a,a97427a,a97428a,a97431a,a97434a,a97435a,a97438a,a97441a,a97442a,a97443a,a97446a,a97449a,a97450a,a97453a,a97456a,a97457a,a97458a,a97461a,a97464a,a97465a,a97468a,a97471a,a97472a,a97473a,a97476a,a97479a,a97480a,a97483a,a97486a,a97487a,a97488a,a97491a,a97494a,a97495a,a97498a,a97501a,a97502a,a97503a,a97506a,a97509a,a97510a,a97513a,a97516a,a97517a,a97518a,a97521a,a97524a,a97525a,a97528a,a97531a,a97532a,a97533a,a97536a,a97539a,a97540a,a97543a,a97546a,a97547a,a97548a,a97551a,a97554a,a97555a,a97558a,a97561a,a97562a,a97563a,a97566a,a97569a,a97570a,a97573a,a97576a,a97577a,a97578a,a97581a,a97584a,a97585a,a97588a,a97591a,a97592a,a97593a,a97596a,a97599a,a97600a,a97603a,a97606a,a97607a,a97608a,a97611a,a97614a,a97615a,a97618a,a97621a,a97622a,a97623a,a97626a,a97629a,a97630a,a97633a,a97636a,a97637a,a97638a,a97641a,a97644a,a97645a,a97648a,a97651a,a97652a,a97653a,a97656a,a97659a,a97660a,a97663a,a97666a,a97667a,a97668a,a97671a,a97674a,a97675a,a97678a,a97681a,a97682a,a97683a,a97686a,a97689a,a97690a,a97693a,a97696a,a97697a,a97698a,a97701a,a97704a,a97705a,a97708a,a97711a,a97712a,a97713a,a97716a,a97719a,a97720a,a97723a,a97726a,a97727a,a97728a,a97731a,a97734a,a97735a,a97738a,a97741a,a97742a,a97743a,a97746a,a97749a,a97750a,a97753a,a97756a,a97757a,a97758a,a97761a,a97764a,a97765a,a97768a,a97771a,a97772a,a97773a,a97776a,a97779a,a97780a,a97783a,a97786a,a97787a,a97788a,a97791a,a97794a,a97795a,a97798a,a97801a,a97802a,a97803a,a97806a,a97809a,a97810a,a97813a,a97816a,a97817a,a97818a,a97821a,a97824a,a97825a,a97828a,a97831a,a97832a,a97833a,a97836a,a97839a,a97840a,a97843a,a97846a,a97847a,a97848a,a97851a,a97854a,a97855a,a97858a,a97861a,a97862a,a97863a,a97866a,a97869a,a97870a,a97873a,a97876a,a97877a,a97878a,a97881a,a97884a,a97885a,a97888a,a97891a,a97892a,a97893a,a97896a,a97899a,a97900a,a97903a,a97906a,a97907a,a97908a,a97911a,a97914a,a97915a,a97918a,a97921a,a97922a,a97923a,a97926a,a97929a,a97930a,a97933a,a97936a,a97937a,a97938a,a97941a,a97944a,a97945a,a97948a,a97951a,a97952a,a97953a,a97956a,a97959a,a97960a,a97963a,a97966a,a97967a,a97968a,a97971a,a97974a,a97975a,a97978a,a97981a,a97982a,a97983a,a97986a,a97989a,a97990a,a97993a,a97996a,a97997a,a97998a,a98001a,a98004a,a98005a,a98008a,a98011a,a98012a,a98013a,a98016a,a98019a,a98020a,a98023a,a98026a,a98027a,a98028a,a98031a,a98034a,a98035a,a98038a,a98041a,a98042a,a98043a,a98046a,a98049a,a98050a,a98053a,a98056a,a98057a,a98058a,a98061a,a98064a,a98065a,a98068a,a98071a,a98072a,a98073a,a98076a,a98079a,a98080a,a98083a,a98086a,a98087a,a98088a,a98091a,a98094a,a98095a,a98098a,a98101a,a98102a,a98103a,a98106a,a98109a,a98110a,a98113a,a98116a,a98117a,a98118a,a98121a,a98124a,a98125a,a98128a,a98131a,a98132a,a98133a,a98136a,a98139a,a98140a,a98143a,a98146a,a98147a,a98148a,a98151a,a98154a,a98155a,a98158a,a98161a,a98162a,a98163a,a98166a,a98169a,a98170a,a98173a,a98176a,a98177a,a98178a,a98181a,a98184a,a98185a,a98188a,a98191a,a98192a,a98193a,a98196a,a98199a,a98200a,a98203a,a98206a,a98207a,a98208a,a98211a,a98214a,a98215a,a98218a,a98221a,a98222a,a98223a,a98226a,a98229a,a98230a,a98233a,a98236a,a98237a,a98238a,a98241a,a98244a,a98245a,a98248a,a98251a,a98252a,a98253a,a98256a,a98259a,a98260a,a98263a,a98266a,a98267a,a98268a,a98271a,a98274a,a98275a,a98278a,a98281a,a98282a,a98283a,a98286a,a98289a,a98290a,a98293a,a98296a,a98297a,a98298a,a98301a,a98304a,a98305a,a98308a,a98311a,a98312a,a98313a,a98316a,a98319a,a98320a,a98323a,a98326a,a98327a,a98328a,a98331a,a98334a,a98335a,a98338a,a98341a,a98342a,a98343a,a98346a,a98349a,a98350a,a98353a,a98356a,a98357a,a98358a,a98361a,a98364a,a98365a,a98368a,a98371a,a98372a,a98373a,a98376a,a98379a,a98380a,a98383a,a98386a,a98387a,a98388a,a98391a,a98394a,a98395a,a98398a,a98401a,a98402a,a98403a,a98406a,a98409a,a98410a,a98413a,a98416a,a98417a,a98418a,a98421a,a98424a,a98425a,a98428a,a98431a,a98432a,a98433a,a98436a,a98439a,a98440a,a98443a,a98446a,a98447a,a98448a,a98451a,a98454a,a98455a,a98458a,a98461a,a98462a,a98463a,a98466a,a98469a,a98470a,a98473a,a98476a,a98477a,a98478a,a98481a,a98484a,a98485a,a98488a,a98491a,a98492a,a98493a,a98496a,a98499a,a98500a,a98503a,a98506a,a98507a,a98508a,a98511a,a98514a,a98515a,a98518a,a98521a,a98522a,a98523a,a98526a,a98529a,a98530a,a98533a,a98536a,a98537a,a98538a,a98541a,a98544a,a98545a,a98548a,a98551a,a98552a,a98553a,a98556a,a98559a,a98560a,a98563a,a98566a,a98567a,a98568a,a98571a,a98574a,a98575a,a98578a,a98581a,a98582a,a98583a,a98586a,a98589a,a98590a,a98593a,a98596a,a98597a,a98598a,a98601a,a98604a,a98605a,a98608a,a98611a,a98612a,a98613a,a98616a,a98619a,a98620a,a98623a,a98626a,a98627a,a98628a,a98631a,a98634a,a98635a,a98638a,a98641a,a98642a,a98643a,a98646a,a98649a,a98650a,a98653a,a98656a,a98657a,a98658a,a98661a,a98664a,a98665a,a98668a,a98671a,a98672a,a98673a,a98676a,a98679a,a98680a,a98683a,a98686a,a98687a,a98688a,a98691a,a98694a,a98695a,a98698a,a98701a,a98702a,a98703a,a98706a,a98709a,a98710a,a98713a,a98716a,a98717a,a98718a,a98721a,a98724a,a98725a,a98728a,a98731a,a98732a,a98733a,a98736a,a98739a,a98740a,a98743a,a98746a,a98747a,a98748a,a98751a,a98754a,a98755a,a98758a,a98761a,a98762a,a98763a,a98766a,a98769a,a98770a,a98773a,a98776a,a98777a,a98778a,a98781a,a98784a,a98785a,a98788a,a98791a,a98792a,a98793a,a98796a,a98799a,a98800a,a98803a,a98806a,a98807a,a98808a,a98811a,a98814a,a98815a,a98818a,a98821a,a98822a,a98823a,a98826a,a98829a,a98830a,a98833a,a98836a,a98837a,a98838a,a98841a,a98844a,a98845a,a98848a,a98851a,a98852a,a98853a,a98856a,a98859a,a98860a,a98863a,a98866a,a98867a,a98868a,a98871a,a98874a,a98875a,a98878a,a98881a,a98882a,a98883a,a98886a,a98889a,a98890a,a98893a,a98896a,a98897a,a98898a,a98901a,a98904a,a98905a,a98908a,a98911a,a98912a,a98913a,a98916a,a98919a,a98920a,a98923a,a98926a,a98927a,a98928a,a98931a,a98934a,a98935a,a98938a,a98941a,a98942a,a98943a,a98946a,a98949a,a98950a,a98953a,a98956a,a98957a,a98958a,a98961a,a98964a,a98965a,a98968a,a98971a,a98972a,a98973a,a98976a,a98979a,a98980a,a98983a,a98986a,a98987a,a98988a,a98991a,a98994a,a98995a,a98998a,a99001a,a99002a,a99003a,a99006a,a99009a,a99010a,a99013a,a99016a,a99017a,a99018a,a99021a,a99024a,a99025a,a99028a,a99031a,a99032a,a99033a,a99036a,a99039a,a99040a,a99043a,a99046a,a99047a,a99048a,a99051a,a99054a,a99055a,a99058a,a99061a,a99062a,a99063a,a99066a,a99069a,a99070a,a99073a,a99076a,a99077a,a99078a,a99081a,a99084a,a99085a,a99088a,a99091a,a99092a,a99093a,a99096a,a99099a,a99100a,a99103a,a99106a,a99107a,a99108a,a99111a,a99114a,a99115a,a99118a,a99121a,a99122a,a99123a,a99126a,a99129a,a99130a,a99133a,a99136a,a99137a,a99138a,a99141a,a99144a,a99145a,a99148a,a99151a,a99152a,a99153a,a99156a,a99159a,a99160a,a99163a,a99166a,a99167a,a99168a,a99171a,a99174a,a99175a,a99178a,a99181a,a99182a,a99183a,a99186a,a99189a,a99190a,a99193a,a99196a,a99197a,a99198a,a99201a,a99204a,a99205a,a99208a,a99211a,a99212a,a99213a,a99216a,a99219a,a99220a,a99223a,a99226a,a99227a,a99228a,a99231a,a99234a,a99235a,a99238a,a99241a,a99242a,a99243a,a99246a,a99249a,a99250a,a99253a,a99256a,a99257a,a99258a,a99261a,a99264a,a99265a,a99268a,a99271a,a99272a,a99273a,a99276a,a99279a,a99280a,a99283a,a99286a,a99287a,a99288a,a99291a,a99294a,a99295a,a99298a,a99301a,a99302a,a99303a,a99306a,a99309a,a99310a,a99313a,a99316a,a99317a,a99318a,a99321a,a99324a,a99325a,a99328a,a99331a,a99332a,a99333a,a99336a,a99339a,a99340a,a99343a,a99346a,a99347a,a99348a,a99351a,a99354a,a99355a,a99358a,a99361a,a99362a,a99363a,a99366a,a99369a,a99370a,a99373a,a99376a,a99377a,a99378a,a99381a,a99384a,a99385a,a99388a,a99391a,a99392a,a99393a,a99396a,a99399a,a99400a,a99403a,a99406a,a99407a,a99408a,a99411a,a99414a,a99415a,a99418a,a99421a,a99422a,a99423a,a99426a,a99429a,a99430a,a99433a,a99436a,a99437a,a99438a,a99441a,a99444a,a99445a,a99448a,a99451a,a99452a,a99453a,a99456a,a99459a,a99460a,a99463a,a99466a,a99467a,a99468a,a99471a,a99474a,a99475a,a99478a,a99481a,a99482a,a99483a,a99486a,a99489a,a99490a,a99493a,a99496a,a99497a,a99498a,a99501a,a99504a,a99505a,a99508a,a99511a,a99512a,a99513a,a99516a,a99519a,a99520a,a99523a,a99526a,a99527a,a99528a,a99531a,a99534a,a99535a,a99538a,a99541a,a99542a,a99543a,a99546a,a99549a,a99550a,a99553a,a99556a,a99557a,a99558a,a99561a,a99564a,a99565a,a99568a,a99571a,a99572a,a99573a,a99576a,a99579a,a99580a,a99583a,a99586a,a99587a,a99588a,a99591a,a99594a,a99595a,a99598a,a99601a,a99602a,a99603a,a99606a,a99609a,a99610a,a99613a,a99616a,a99617a,a99618a,a99621a,a99624a,a99625a,a99628a,a99631a,a99632a,a99633a,a99636a,a99639a,a99640a,a99643a,a99646a,a99647a,a99648a,a99651a,a99654a,a99655a,a99658a,a99661a,a99662a,a99663a,a99666a,a99669a,a99670a,a99673a,a99676a,a99677a,a99678a,a99681a,a99684a,a99685a,a99688a,a99691a,a99692a,a99693a,a99696a,a99699a,a99700a,a99703a,a99706a,a99707a,a99708a,a99711a,a99714a,a99715a,a99718a,a99721a,a99722a,a99723a,a99726a,a99729a,a99730a,a99733a,a99736a,a99737a,a99738a,a99741a,a99744a,a99745a,a99748a,a99751a,a99752a,a99753a,a99756a,a99759a,a99760a,a99763a,a99766a,a99767a,a99768a,a99771a,a99774a,a99775a,a99778a,a99781a,a99782a,a99783a,a99786a,a99789a,a99790a,a99793a,a99796a,a99797a,a99798a,a99801a,a99804a,a99805a,a99808a,a99811a,a99812a,a99813a,a99816a,a99819a,a99820a,a99823a,a99826a,a99827a,a99828a,a99831a,a99834a,a99835a,a99838a,a99841a,a99842a,a99843a,a99846a,a99849a,a99850a,a99853a,a99856a,a99857a,a99858a,a99861a,a99864a,a99865a,a99868a,a99871a,a99872a,a99873a,a99876a,a99879a,a99880a,a99883a,a99886a,a99887a,a99888a,a99891a,a99894a,a99895a,a99898a,a99901a,a99902a,a99903a,a99906a,a99909a,a99910a,a99913a,a99916a,a99917a,a99918a,a99921a,a99924a,a99925a,a99928a,a99931a,a99932a,a99933a,a99936a,a99939a,a99940a,a99943a,a99946a,a99947a,a99948a,a99951a,a99954a,a99955a,a99958a,a99961a,a99962a,a99963a,a99966a,a99969a,a99970a,a99973a,a99976a,a99977a,a99978a,a99981a,a99984a,a99985a,a99988a,a99991a,a99992a,a99993a,a99996a,a99999a,a100000a,a100003a,a100006a,a100007a,a100008a,a100011a,a100014a,a100015a,a100018a,a100021a,a100022a,a100023a,a100026a,a100029a,a100030a,a100033a,a100036a,a100037a,a100038a,a100041a,a100044a,a100045a,a100048a,a100051a,a100052a,a100053a,a100056a,a100059a,a100060a,a100063a,a100066a,a100067a,a100068a,a100071a,a100074a,a100075a,a100078a,a100081a,a100082a,a100083a,a100086a,a100089a,a100090a,a100093a,a100096a,a100097a,a100098a,a100101a,a100104a,a100105a,a100108a,a100111a,a100112a,a100113a,a100116a,a100119a,a100120a,a100123a,a100126a,a100127a,a100128a,a100131a,a100134a,a100135a,a100138a,a100141a,a100142a,a100143a,a100146a,a100149a,a100150a,a100153a,a100156a,a100157a,a100158a,a100161a,a100164a,a100165a,a100168a,a100171a,a100172a,a100173a,a100176a,a100179a,a100180a,a100183a,a100186a,a100187a,a100188a,a100191a,a100194a,a100195a,a100198a,a100201a,a100202a,a100203a,a100206a,a100209a,a100210a,a100213a,a100216a,a100217a,a100218a,a100221a,a100224a,a100225a,a100228a,a100231a,a100232a,a100233a,a100236a,a100239a,a100240a,a100243a,a100246a,a100247a,a100248a,a100251a,a100254a,a100255a,a100258a,a100261a,a100262a,a100263a,a100266a,a100269a,a100270a,a100273a,a100276a,a100277a,a100278a,a100281a,a100284a,a100285a,a100288a,a100291a,a100292a,a100293a,a100296a,a100299a,a100300a,a100303a,a100306a,a100307a,a100308a,a100311a,a100314a,a100315a,a100318a,a100321a,a100322a,a100323a,a100326a,a100329a,a100330a,a100333a,a100336a,a100337a,a100338a,a100341a,a100344a,a100345a,a100348a,a100351a,a100352a,a100353a,a100356a,a100359a,a100360a,a100363a,a100366a,a100367a,a100368a,a100371a,a100374a,a100375a,a100378a,a100381a,a100382a,a100383a,a100386a,a100389a,a100390a,a100393a,a100396a,a100397a,a100398a,a100401a,a100404a,a100405a,a100408a,a100411a,a100412a,a100413a,a100416a,a100419a,a100420a,a100423a,a100426a,a100427a,a100428a,a100431a,a100434a,a100435a,a100438a,a100441a,a100442a,a100443a,a100446a,a100449a,a100450a,a100453a,a100456a,a100457a,a100458a,a100461a,a100464a,a100465a,a100468a,a100471a,a100472a,a100473a,a100476a,a100479a,a100480a,a100483a,a100486a,a100487a,a100488a,a100491a,a100494a,a100495a,a100498a,a100501a,a100502a,a100503a,a100506a,a100509a,a100510a,a100513a,a100516a,a100517a,a100518a,a100521a,a100524a,a100525a,a100528a,a100531a,a100532a,a100533a,a100536a,a100539a,a100540a,a100543a,a100546a,a100547a,a100548a,a100551a,a100554a,a100555a,a100558a,a100561a,a100562a,a100563a,a100566a,a100569a,a100570a,a100573a,a100576a,a100577a,a100578a,a100581a,a100584a,a100585a,a100588a,a100591a,a100592a,a100593a,a100596a,a100599a,a100600a,a100603a,a100606a,a100607a,a100608a,a100611a,a100614a,a100615a,a100618a,a100621a,a100622a,a100623a,a100626a,a100629a,a100630a,a100633a,a100636a,a100637a,a100638a,a100641a,a100644a,a100645a,a100648a,a100651a,a100652a,a100653a,a100656a,a100659a,a100660a,a100663a,a100666a,a100667a,a100668a,a100671a,a100674a,a100675a,a100678a,a100681a,a100682a,a100683a,a100686a,a100689a,a100690a,a100693a,a100696a,a100697a,a100698a,a100701a,a100704a,a100705a,a100708a,a100711a,a100712a,a100713a,a100716a,a100719a,a100720a,a100723a,a100726a,a100727a,a100728a,a100731a,a100734a,a100735a,a100738a,a100741a,a100742a,a100743a,a100746a,a100749a,a100750a,a100753a,a100756a,a100757a,a100758a,a100761a,a100764a,a100765a,a100768a,a100771a,a100772a,a100773a,a100776a,a100779a,a100780a,a100783a,a100786a,a100787a,a100788a,a100791a,a100794a,a100795a,a100798a,a100801a,a100802a,a100803a,a100806a,a100809a,a100810a,a100813a,a100816a,a100817a,a100818a,a100821a,a100824a,a100825a,a100828a,a100831a,a100832a,a100833a,a100836a,a100839a,a100840a,a100843a,a100846a,a100847a,a100848a,a100851a,a100854a,a100855a,a100858a,a100861a,a100862a,a100863a,a100866a,a100869a,a100870a,a100873a,a100876a,a100877a,a100878a,a100881a,a100884a,a100885a,a100888a,a100891a,a100892a,a100893a,a100896a,a100899a,a100900a,a100903a,a100906a,a100907a,a100908a,a100911a,a100914a,a100915a,a100918a,a100921a,a100922a,a100923a,a100926a,a100929a,a100930a,a100933a,a100936a,a100937a,a100938a,a100941a,a100944a,a100945a,a100948a,a100951a,a100952a,a100953a,a100956a,a100959a,a100960a,a100963a,a100966a,a100967a,a100968a,a100971a,a100974a,a100975a,a100978a,a100981a,a100982a,a100983a,a100986a,a100989a,a100990a,a100993a,a100996a,a100997a,a100998a,a101001a,a101004a,a101005a,a101008a,a101011a,a101012a,a101013a,a101016a,a101019a,a101020a,a101023a,a101026a,a101027a,a101028a,a101031a,a101034a,a101035a,a101038a,a101041a,a101042a,a101043a,a101046a,a101049a,a101050a,a101053a,a101056a,a101057a,a101058a,a101061a,a101064a,a101065a,a101068a,a101071a,a101072a,a101073a,a101076a,a101079a,a101080a,a101083a,a101086a,a101087a,a101088a,a101091a,a101094a,a101095a,a101098a,a101101a,a101102a,a101103a,a101106a,a101109a,a101110a,a101113a,a101116a,a101117a,a101118a,a101121a,a101124a,a101125a,a101128a,a101131a,a101132a,a101133a,a101136a,a101139a,a101140a,a101143a,a101146a,a101147a,a101148a,a101151a,a101154a,a101155a,a101158a,a101161a,a101162a,a101163a,a101166a,a101169a,a101170a,a101173a,a101176a,a101177a,a101178a,a101181a,a101184a,a101185a,a101188a,a101191a,a101192a,a101193a,a101196a,a101199a,a101200a,a101203a,a101206a,a101207a,a101208a,a101211a,a101214a,a101215a,a101218a,a101221a,a101222a,a101223a,a101226a,a101229a,a101230a,a101233a,a101236a,a101237a,a101238a,a101241a,a101244a,a101245a,a101248a,a101251a,a101252a,a101253a,a101256a,a101259a,a101260a,a101263a,a101266a,a101267a,a101268a,a101271a,a101274a,a101275a,a101278a,a101281a,a101282a,a101283a,a101286a,a101289a,a101290a,a101293a,a101296a,a101297a,a101298a,a101301a,a101304a,a101305a,a101308a,a101311a,a101312a,a101313a,a101316a,a101319a,a101320a,a101323a,a101326a,a101327a,a101328a,a101331a,a101334a,a101335a,a101338a,a101341a,a101342a,a101343a,a101346a,a101349a,a101350a,a101353a,a101356a,a101357a,a101358a,a101361a,a101364a,a101365a,a101368a,a101371a,a101372a,a101373a,a101376a,a101379a,a101380a,a101383a,a101386a,a101387a,a101388a,a101391a,a101394a,a101395a,a101398a,a101401a,a101402a,a101403a,a101406a,a101409a,a101410a,a101413a,a101416a,a101417a,a101418a,a101421a,a101424a,a101425a,a101428a,a101431a,a101432a,a101433a,a101436a,a101439a,a101440a,a101443a,a101446a,a101447a,a101448a,a101451a,a101454a,a101455a,a101458a,a101461a,a101462a,a101463a,a101466a,a101469a,a101470a,a101473a,a101476a,a101477a,a101478a,a101481a,a101484a,a101485a,a101488a,a101491a,a101492a,a101493a,a101496a,a101499a,a101500a,a101503a,a101506a,a101507a,a101508a,a101511a,a101514a,a101515a,a101518a,a101521a,a101522a,a101523a,a101526a,a101529a,a101530a,a101533a,a101536a,a101537a,a101538a,a101541a,a101544a,a101545a,a101548a,a101551a,a101552a,a101553a,a101556a,a101559a,a101560a,a101563a,a101566a,a101567a,a101568a,a101571a,a101574a,a101575a,a101578a,a101581a,a101582a,a101583a,a101586a,a101589a,a101590a,a101593a,a101596a,a101597a,a101598a,a101601a,a101604a,a101605a,a101608a,a101611a,a101612a,a101613a,a101616a,a101619a,a101620a,a101623a,a101626a,a101627a,a101628a,a101631a,a101634a,a101635a,a101638a,a101641a,a101642a,a101643a,a101646a,a101649a,a101650a,a101653a,a101656a,a101657a,a101658a,a101661a,a101664a,a101665a,a101668a,a101671a,a101672a,a101673a,a101676a,a101679a,a101680a,a101683a,a101686a,a101687a,a101688a,a101691a,a101694a,a101695a,a101698a,a101701a,a101702a,a101703a,a101706a,a101709a,a101710a,a101713a,a101716a,a101717a,a101718a,a101721a,a101724a,a101725a,a101728a,a101731a,a101732a,a101733a,a101736a,a101739a,a101740a,a101743a,a101746a,a101747a,a101748a,a101751a,a101754a,a101755a,a101758a,a101761a,a101762a,a101763a,a101766a,a101769a,a101770a,a101773a,a101777a,a101778a,a101779a,a101780a,a101783a,a101786a,a101787a,a101790a,a101793a,a101794a,a101795a,a101798a,a101801a,a101802a,a101805a,a101809a,a101810a,a101811a,a101812a,a101815a,a101818a,a101819a,a101822a,a101825a,a101826a,a101827a,a101830a,a101833a,a101834a,a101837a,a101841a,a101842a,a101843a,a101844a,a101847a,a101850a,a101851a,a101854a,a101857a,a101858a,a101859a,a101862a,a101865a,a101866a,a101869a,a101873a,a101874a,a101875a,a101876a,a101879a,a101882a,a101883a,a101886a,a101889a,a101890a,a101891a,a101894a,a101897a,a101898a,a101901a,a101905a,a101906a,a101907a,a101908a,a101911a,a101914a,a101915a,a101918a,a101921a,a101922a,a101923a,a101926a,a101929a,a101930a,a101933a,a101937a,a101938a,a101939a,a101940a,a101943a,a101946a,a101947a,a101950a,a101953a,a101954a,a101955a,a101958a,a101961a,a101962a,a101965a,a101969a,a101970a,a101971a,a101972a,a101975a,a101978a,a101979a,a101982a,a101985a,a101986a,a101987a,a101990a,a101993a,a101994a,a101997a,a102001a,a102002a,a102003a,a102004a,a102007a,a102010a,a102011a,a102014a,a102017a,a102018a,a102019a,a102022a,a102025a,a102026a,a102029a,a102033a,a102034a,a102035a,a102036a,a102039a,a102042a,a102043a,a102046a,a102049a,a102050a,a102051a,a102054a,a102057a,a102058a,a102061a,a102065a,a102066a,a102067a,a102068a,a102071a,a102074a,a102075a,a102078a,a102081a,a102082a,a102083a,a102086a,a102089a,a102090a,a102093a,a102097a,a102098a,a102099a,a102100a,a102103a,a102106a,a102107a,a102110a,a102113a,a102114a,a102115a,a102118a,a102121a,a102122a,a102125a,a102129a,a102130a,a102131a,a102132a,a102135a,a102138a,a102139a,a102142a,a102145a,a102146a,a102147a,a102150a,a102153a,a102154a,a102157a,a102161a,a102162a,a102163a,a102164a,a102167a,a102170a,a102171a,a102174a,a102177a,a102178a,a102179a,a102182a,a102185a,a102186a,a102189a,a102193a,a102194a,a102195a,a102196a,a102199a,a102202a,a102203a,a102206a,a102209a,a102210a,a102211a,a102214a,a102217a,a102218a,a102221a,a102225a,a102226a,a102227a,a102228a,a102231a,a102234a,a102235a,a102238a,a102241a,a102242a,a102243a,a102246a,a102249a,a102250a,a102253a,a102257a,a102258a,a102259a,a102260a,a102263a,a102266a,a102267a,a102270a,a102273a,a102274a,a102275a,a102278a,a102281a,a102282a,a102285a,a102289a,a102290a,a102291a,a102292a,a102295a,a102298a,a102299a,a102302a,a102305a,a102306a,a102307a,a102310a,a102313a,a102314a,a102317a,a102321a,a102322a,a102323a,a102324a,a102327a,a102330a,a102331a,a102334a,a102337a,a102338a,a102339a,a102342a,a102345a,a102346a,a102349a,a102353a,a102354a,a102355a,a102356a,a102359a,a102362a,a102363a,a102366a,a102369a,a102370a,a102371a,a102374a,a102377a,a102378a,a102381a,a102385a,a102386a,a102387a,a102388a,a102391a,a102394a,a102395a,a102398a,a102401a,a102402a,a102403a,a102406a,a102409a,a102410a,a102413a,a102417a,a102418a,a102419a,a102420a,a102423a,a102426a,a102427a,a102430a,a102433a,a102434a,a102435a,a102438a,a102441a,a102442a,a102445a,a102449a,a102450a,a102451a,a102452a,a102455a,a102458a,a102459a,a102462a,a102465a,a102466a,a102467a,a102470a,a102473a,a102474a,a102477a,a102481a,a102482a,a102483a,a102484a,a102487a,a102490a,a102491a,a102494a,a102497a,a102498a,a102499a,a102502a,a102505a,a102506a,a102509a,a102513a,a102514a,a102515a,a102516a,a102519a,a102522a,a102523a,a102526a,a102529a,a102530a,a102531a,a102534a,a102537a,a102538a,a102541a,a102545a,a102546a,a102547a,a102548a,a102551a,a102554a,a102555a,a102558a,a102561a,a102562a,a102563a,a102566a,a102569a,a102570a,a102573a,a102577a,a102578a,a102579a,a102580a,a102583a,a102586a,a102587a,a102590a,a102593a,a102594a,a102595a,a102598a,a102601a,a102602a,a102605a,a102609a,a102610a,a102611a,a102612a,a102615a,a102618a,a102619a,a102622a,a102625a,a102626a,a102627a,a102630a,a102633a,a102634a,a102637a,a102641a,a102642a,a102643a,a102644a,a102647a,a102650a,a102651a,a102654a,a102657a,a102658a,a102659a,a102662a,a102665a,a102666a,a102669a,a102673a,a102674a,a102675a,a102676a,a102679a,a102682a,a102683a,a102686a,a102689a,a102690a,a102691a,a102694a,a102697a,a102698a,a102701a,a102705a,a102706a,a102707a,a102708a,a102711a,a102714a,a102715a,a102718a,a102721a,a102722a,a102723a,a102726a,a102729a,a102730a,a102733a,a102737a,a102738a,a102739a,a102740a,a102743a,a102746a,a102747a,a102750a,a102753a,a102754a,a102755a,a102758a,a102761a,a102762a,a102765a,a102769a,a102770a,a102771a,a102772a,a102775a,a102778a,a102779a,a102782a,a102785a,a102786a,a102787a,a102790a,a102793a,a102794a,a102797a,a102801a,a102802a,a102803a,a102804a,a102807a,a102810a,a102811a,a102814a,a102817a,a102818a,a102819a,a102822a,a102825a,a102826a,a102829a,a102833a,a102834a,a102835a,a102836a,a102839a,a102842a,a102843a,a102846a,a102849a,a102850a,a102851a,a102854a,a102857a,a102858a,a102861a,a102865a,a102866a,a102867a,a102868a,a102871a,a102874a,a102875a,a102878a,a102881a,a102882a,a102883a,a102886a,a102889a,a102890a,a102893a,a102897a,a102898a,a102899a,a102900a,a102903a,a102906a,a102907a,a102910a,a102913a,a102914a,a102915a,a102918a,a102921a,a102922a,a102925a,a102929a,a102930a,a102931a,a102932a,a102935a,a102938a,a102939a,a102942a,a102945a,a102946a,a102947a,a102950a,a102953a,a102954a,a102957a,a102961a,a102962a,a102963a,a102964a,a102967a,a102970a,a102971a,a102974a,a102977a,a102978a,a102979a,a102982a,a102985a,a102986a,a102989a,a102993a,a102994a,a102995a,a102996a,a102999a,a103002a,a103003a,a103006a,a103009a,a103010a,a103011a,a103014a,a103017a,a103018a,a103021a,a103025a,a103026a,a103027a,a103028a,a103031a,a103034a,a103035a,a103038a,a103041a,a103042a,a103043a,a103046a,a103049a,a103050a,a103053a,a103057a,a103058a,a103059a,a103060a,a103063a,a103066a,a103067a,a103070a,a103073a,a103074a,a103075a,a103078a,a103081a,a103082a,a103085a,a103089a,a103090a,a103091a,a103092a,a103095a,a103098a,a103099a,a103102a,a103105a,a103106a,a103107a,a103110a,a103113a,a103114a,a103117a,a103121a,a103122a,a103123a,a103124a,a103127a,a103130a,a103131a,a103134a,a103137a,a103138a,a103139a,a103142a,a103145a,a103146a,a103149a,a103153a,a103154a,a103155a,a103156a,a103159a,a103162a,a103163a,a103166a,a103169a,a103170a,a103171a,a103174a,a103177a,a103178a,a103181a,a103185a,a103186a,a103187a,a103188a,a103191a,a103194a,a103195a,a103198a,a103201a,a103202a,a103203a,a103206a,a103209a,a103210a,a103213a,a103217a,a103218a,a103219a,a103220a,a103223a,a103226a,a103227a,a103230a,a103233a,a103234a,a103235a,a103238a,a103241a,a103242a,a103245a,a103249a,a103250a,a103251a,a103252a,a103255a,a103258a,a103259a,a103262a,a103265a,a103266a,a103267a,a103270a,a103273a,a103274a,a103277a,a103281a,a103282a,a103283a,a103284a,a103287a,a103290a,a103291a,a103294a,a103297a,a103298a,a103299a,a103302a,a103305a,a103306a,a103309a,a103313a,a103314a,a103315a,a103316a,a103319a,a103322a,a103323a,a103326a,a103329a,a103330a,a103331a,a103334a,a103337a,a103338a,a103341a,a103345a,a103346a,a103347a,a103348a,a103351a,a103354a,a103355a,a103358a,a103361a,a103362a,a103363a,a103366a,a103369a,a103370a,a103373a,a103377a,a103378a,a103379a,a103380a,a103383a,a103386a,a103387a,a103390a,a103393a,a103394a,a103395a,a103398a,a103401a,a103402a,a103405a,a103409a,a103410a,a103411a,a103412a,a103415a,a103418a,a103419a,a103422a,a103425a,a103426a,a103427a,a103430a,a103433a,a103434a,a103437a,a103441a,a103442a,a103443a,a103444a,a103447a,a103450a,a103451a,a103454a,a103457a,a103458a,a103459a,a103462a,a103465a,a103466a,a103469a,a103473a,a103474a,a103475a,a103476a,a103479a,a103482a,a103483a,a103486a,a103489a,a103490a,a103491a,a103494a,a103497a,a103498a,a103501a,a103505a,a103506a,a103507a,a103508a,a103511a,a103514a,a103515a,a103518a,a103521a,a103522a,a103523a,a103526a,a103529a,a103530a,a103533a,a103537a,a103538a,a103539a,a103540a,a103543a,a103546a,a103547a,a103550a,a103553a,a103554a,a103555a,a103558a,a103561a,a103562a,a103565a,a103569a,a103570a,a103571a,a103572a,a103575a,a103578a,a103579a,a103582a,a103585a,a103586a,a103587a,a103590a,a103593a,a103594a,a103597a,a103601a,a103602a,a103603a,a103604a,a103607a,a103610a,a103611a,a103614a,a103617a,a103618a,a103619a,a103622a,a103625a,a103626a,a103629a,a103633a,a103634a,a103635a,a103636a,a103639a,a103642a,a103643a,a103646a,a103649a,a103650a,a103651a,a103654a,a103657a,a103658a,a103661a,a103665a,a103666a,a103667a,a103668a,a103671a,a103674a,a103675a,a103678a,a103681a,a103682a,a103683a,a103686a,a103689a,a103690a,a103693a,a103697a,a103698a,a103699a,a103700a,a103703a,a103706a,a103707a,a103710a,a103713a,a103714a,a103715a,a103718a,a103721a,a103722a,a103725a,a103729a,a103730a,a103731a,a103732a,a103735a,a103738a,a103739a,a103742a,a103745a,a103746a,a103747a,a103750a,a103753a,a103754a,a103757a,a103761a,a103762a,a103763a,a103764a,a103767a,a103770a,a103771a,a103774a,a103777a,a103778a,a103779a,a103782a,a103785a,a103786a,a103789a,a103793a,a103794a,a103795a,a103796a,a103799a,a103802a,a103803a,a103806a,a103809a,a103810a,a103811a,a103814a,a103817a,a103818a,a103821a,a103825a,a103826a,a103827a,a103828a,a103831a,a103834a,a103835a,a103838a,a103841a,a103842a,a103843a,a103846a,a103849a,a103850a,a103853a,a103857a,a103858a,a103859a,a103860a,a103863a,a103866a,a103867a,a103870a,a103873a,a103874a,a103875a,a103878a,a103881a,a103882a,a103885a,a103889a,a103890a,a103891a,a103892a,a103895a,a103898a,a103899a,a103902a,a103905a,a103906a,a103907a,a103910a,a103913a,a103914a,a103917a,a103921a,a103922a,a103923a,a103924a,a103927a,a103930a,a103931a,a103934a,a103937a,a103938a,a103939a,a103942a,a103945a,a103946a,a103949a,a103953a,a103954a,a103955a,a103956a,a103959a,a103962a,a103963a,a103966a,a103969a,a103970a,a103971a,a103974a,a103977a,a103978a,a103981a,a103985a,a103986a,a103987a,a103988a,a103991a,a103994a,a103995a,a103998a,a104001a,a104002a,a104003a,a104006a,a104009a,a104010a,a104013a,a104017a,a104018a,a104019a,a104020a,a104023a,a104026a,a104027a,a104030a,a104033a,a104034a,a104035a,a104038a,a104041a,a104042a,a104045a,a104049a,a104050a,a104051a,a104052a,a104055a,a104058a,a104059a,a104062a,a104065a,a104066a,a104067a,a104070a,a104073a,a104074a,a104077a,a104081a,a104082a,a104083a,a104084a,a104087a,a104090a,a104091a,a104094a,a104097a,a104098a,a104099a,a104102a,a104105a,a104106a,a104109a,a104113a,a104114a,a104115a,a104116a,a104119a,a104122a,a104123a,a104126a,a104129a,a104130a,a104131a,a104134a,a104137a,a104138a,a104141a,a104145a,a104146a,a104147a,a104148a,a104151a,a104154a,a104155a,a104158a,a104161a,a104162a,a104163a,a104166a,a104169a,a104170a,a104173a,a104177a,a104178a,a104179a,a104180a,a104183a,a104186a,a104187a,a104190a,a104193a,a104194a,a104195a,a104198a,a104201a,a104202a,a104205a,a104209a,a104210a,a104211a,a104212a,a104215a,a104218a,a104219a,a104222a,a104225a,a104226a,a104227a,a104230a,a104233a,a104234a,a104237a,a104241a,a104242a,a104243a,a104244a,a104247a,a104250a,a104251a,a104254a,a104257a,a104258a,a104259a,a104262a,a104265a,a104266a,a104269a,a104273a,a104274a,a104275a,a104276a,a104279a,a104282a,a104283a,a104286a,a104289a,a104290a,a104291a,a104294a,a104297a,a104298a,a104301a,a104305a,a104306a,a104307a,a104308a,a104311a,a104314a,a104315a,a104318a,a104322a,a104323a,a104324a,a104325a,a104328a,a104331a,a104332a,a104335a,a104339a,a104340a,a104341a,a104342a,a104345a,a104348a,a104349a,a104352a,a104356a,a104357a,a104358a,a104359a,a104362a,a104365a,a104366a,a104369a,a104373a,a104374a,a104375a,a104376a,a104379a,a104382a,a104383a,a104386a,a104390a,a104391a,a104392a,a104393a,a104396a,a104399a,a104400a,a104403a,a104407a,a104408a,a104409a,a104410a,a104413a,a104416a,a104417a,a104420a,a104424a,a104425a,a104426a,a104427a,a104430a,a104433a,a104434a,a104437a,a104441a,a104442a,a104443a,a104444a,a104447a,a104450a,a104451a,a104454a,a104458a,a104459a,a104460a,a104461a,a104464a,a104467a,a104468a,a104471a,a104475a,a104476a,a104477a,a104478a,a104481a,a104484a,a104485a,a104488a,a104492a,a104493a,a104494a,a104495a,a104498a,a104501a,a104502a,a104505a,a104509a,a104510a,a104511a,a104512a,a104515a,a104518a,a104519a,a104522a,a104526a,a104527a,a104528a,a104529a,a104532a,a104535a,a104536a,a104539a,a104543a,a104544a,a104545a,a104546a,a104549a,a104552a,a104553a,a104556a,a104560a,a104561a,a104562a,a104563a,a104566a,a104569a,a104570a,a104573a,a104577a,a104578a,a104579a,a104580a: std_logic;
begin

A7 <=( a11512a ) or ( a7675a );
 a1a <=( a104580a  and  a104563a );
 a2a <=( a104546a  and  a104529a );
 a3a <=( a104512a  and  a104495a );
 a4a <=( a104478a  and  a104461a );
 a5a <=( a104444a  and  a104427a );
 a6a <=( a104410a  and  a104393a );
 a7a <=( a104376a  and  a104359a );
 a8a <=( a104342a  and  a104325a );
 a9a <=( a104308a  and  a104291a );
 a10a <=( a104276a  and  a104259a );
 a11a <=( a104244a  and  a104227a );
 a12a <=( a104212a  and  a104195a );
 a13a <=( a104180a  and  a104163a );
 a14a <=( a104148a  and  a104131a );
 a15a <=( a104116a  and  a104099a );
 a16a <=( a104084a  and  a104067a );
 a17a <=( a104052a  and  a104035a );
 a18a <=( a104020a  and  a104003a );
 a19a <=( a103988a  and  a103971a );
 a20a <=( a103956a  and  a103939a );
 a21a <=( a103924a  and  a103907a );
 a22a <=( a103892a  and  a103875a );
 a23a <=( a103860a  and  a103843a );
 a24a <=( a103828a  and  a103811a );
 a25a <=( a103796a  and  a103779a );
 a26a <=( a103764a  and  a103747a );
 a27a <=( a103732a  and  a103715a );
 a28a <=( a103700a  and  a103683a );
 a29a <=( a103668a  and  a103651a );
 a30a <=( a103636a  and  a103619a );
 a31a <=( a103604a  and  a103587a );
 a32a <=( a103572a  and  a103555a );
 a33a <=( a103540a  and  a103523a );
 a34a <=( a103508a  and  a103491a );
 a35a <=( a103476a  and  a103459a );
 a36a <=( a103444a  and  a103427a );
 a37a <=( a103412a  and  a103395a );
 a38a <=( a103380a  and  a103363a );
 a39a <=( a103348a  and  a103331a );
 a40a <=( a103316a  and  a103299a );
 a41a <=( a103284a  and  a103267a );
 a42a <=( a103252a  and  a103235a );
 a43a <=( a103220a  and  a103203a );
 a44a <=( a103188a  and  a103171a );
 a45a <=( a103156a  and  a103139a );
 a46a <=( a103124a  and  a103107a );
 a47a <=( a103092a  and  a103075a );
 a48a <=( a103060a  and  a103043a );
 a49a <=( a103028a  and  a103011a );
 a50a <=( a102996a  and  a102979a );
 a51a <=( a102964a  and  a102947a );
 a52a <=( a102932a  and  a102915a );
 a53a <=( a102900a  and  a102883a );
 a54a <=( a102868a  and  a102851a );
 a55a <=( a102836a  and  a102819a );
 a56a <=( a102804a  and  a102787a );
 a57a <=( a102772a  and  a102755a );
 a58a <=( a102740a  and  a102723a );
 a59a <=( a102708a  and  a102691a );
 a60a <=( a102676a  and  a102659a );
 a61a <=( a102644a  and  a102627a );
 a62a <=( a102612a  and  a102595a );
 a63a <=( a102580a  and  a102563a );
 a64a <=( a102548a  and  a102531a );
 a65a <=( a102516a  and  a102499a );
 a66a <=( a102484a  and  a102467a );
 a67a <=( a102452a  and  a102435a );
 a68a <=( a102420a  and  a102403a );
 a69a <=( a102388a  and  a102371a );
 a70a <=( a102356a  and  a102339a );
 a71a <=( a102324a  and  a102307a );
 a72a <=( a102292a  and  a102275a );
 a73a <=( a102260a  and  a102243a );
 a74a <=( a102228a  and  a102211a );
 a75a <=( a102196a  and  a102179a );
 a76a <=( a102164a  and  a102147a );
 a77a <=( a102132a  and  a102115a );
 a78a <=( a102100a  and  a102083a );
 a79a <=( a102068a  and  a102051a );
 a80a <=( a102036a  and  a102019a );
 a81a <=( a102004a  and  a101987a );
 a82a <=( a101972a  and  a101955a );
 a83a <=( a101940a  and  a101923a );
 a84a <=( a101908a  and  a101891a );
 a85a <=( a101876a  and  a101859a );
 a86a <=( a101844a  and  a101827a );
 a87a <=( a101812a  and  a101795a );
 a88a <=( a101780a  and  a101763a );
 a89a <=( a101748a  and  a101733a );
 a90a <=( a101718a  and  a101703a );
 a91a <=( a101688a  and  a101673a );
 a92a <=( a101658a  and  a101643a );
 a93a <=( a101628a  and  a101613a );
 a94a <=( a101598a  and  a101583a );
 a95a <=( a101568a  and  a101553a );
 a96a <=( a101538a  and  a101523a );
 a97a <=( a101508a  and  a101493a );
 a98a <=( a101478a  and  a101463a );
 a99a <=( a101448a  and  a101433a );
 a100a <=( a101418a  and  a101403a );
 a101a <=( a101388a  and  a101373a );
 a102a <=( a101358a  and  a101343a );
 a103a <=( a101328a  and  a101313a );
 a104a <=( a101298a  and  a101283a );
 a105a <=( a101268a  and  a101253a );
 a106a <=( a101238a  and  a101223a );
 a107a <=( a101208a  and  a101193a );
 a108a <=( a101178a  and  a101163a );
 a109a <=( a101148a  and  a101133a );
 a110a <=( a101118a  and  a101103a );
 a111a <=( a101088a  and  a101073a );
 a112a <=( a101058a  and  a101043a );
 a113a <=( a101028a  and  a101013a );
 a114a <=( a100998a  and  a100983a );
 a115a <=( a100968a  and  a100953a );
 a116a <=( a100938a  and  a100923a );
 a117a <=( a100908a  and  a100893a );
 a118a <=( a100878a  and  a100863a );
 a119a <=( a100848a  and  a100833a );
 a120a <=( a100818a  and  a100803a );
 a121a <=( a100788a  and  a100773a );
 a122a <=( a100758a  and  a100743a );
 a123a <=( a100728a  and  a100713a );
 a124a <=( a100698a  and  a100683a );
 a125a <=( a100668a  and  a100653a );
 a126a <=( a100638a  and  a100623a );
 a127a <=( a100608a  and  a100593a );
 a128a <=( a100578a  and  a100563a );
 a129a <=( a100548a  and  a100533a );
 a130a <=( a100518a  and  a100503a );
 a131a <=( a100488a  and  a100473a );
 a132a <=( a100458a  and  a100443a );
 a133a <=( a100428a  and  a100413a );
 a134a <=( a100398a  and  a100383a );
 a135a <=( a100368a  and  a100353a );
 a136a <=( a100338a  and  a100323a );
 a137a <=( a100308a  and  a100293a );
 a138a <=( a100278a  and  a100263a );
 a139a <=( a100248a  and  a100233a );
 a140a <=( a100218a  and  a100203a );
 a141a <=( a100188a  and  a100173a );
 a142a <=( a100158a  and  a100143a );
 a143a <=( a100128a  and  a100113a );
 a144a <=( a100098a  and  a100083a );
 a145a <=( a100068a  and  a100053a );
 a146a <=( a100038a  and  a100023a );
 a147a <=( a100008a  and  a99993a );
 a148a <=( a99978a  and  a99963a );
 a149a <=( a99948a  and  a99933a );
 a150a <=( a99918a  and  a99903a );
 a151a <=( a99888a  and  a99873a );
 a152a <=( a99858a  and  a99843a );
 a153a <=( a99828a  and  a99813a );
 a154a <=( a99798a  and  a99783a );
 a155a <=( a99768a  and  a99753a );
 a156a <=( a99738a  and  a99723a );
 a157a <=( a99708a  and  a99693a );
 a158a <=( a99678a  and  a99663a );
 a159a <=( a99648a  and  a99633a );
 a160a <=( a99618a  and  a99603a );
 a161a <=( a99588a  and  a99573a );
 a162a <=( a99558a  and  a99543a );
 a163a <=( a99528a  and  a99513a );
 a164a <=( a99498a  and  a99483a );
 a165a <=( a99468a  and  a99453a );
 a166a <=( a99438a  and  a99423a );
 a167a <=( a99408a  and  a99393a );
 a168a <=( a99378a  and  a99363a );
 a169a <=( a99348a  and  a99333a );
 a170a <=( a99318a  and  a99303a );
 a171a <=( a99288a  and  a99273a );
 a172a <=( a99258a  and  a99243a );
 a173a <=( a99228a  and  a99213a );
 a174a <=( a99198a  and  a99183a );
 a175a <=( a99168a  and  a99153a );
 a176a <=( a99138a  and  a99123a );
 a177a <=( a99108a  and  a99093a );
 a178a <=( a99078a  and  a99063a );
 a179a <=( a99048a  and  a99033a );
 a180a <=( a99018a  and  a99003a );
 a181a <=( a98988a  and  a98973a );
 a182a <=( a98958a  and  a98943a );
 a183a <=( a98928a  and  a98913a );
 a184a <=( a98898a  and  a98883a );
 a185a <=( a98868a  and  a98853a );
 a186a <=( a98838a  and  a98823a );
 a187a <=( a98808a  and  a98793a );
 a188a <=( a98778a  and  a98763a );
 a189a <=( a98748a  and  a98733a );
 a190a <=( a98718a  and  a98703a );
 a191a <=( a98688a  and  a98673a );
 a192a <=( a98658a  and  a98643a );
 a193a <=( a98628a  and  a98613a );
 a194a <=( a98598a  and  a98583a );
 a195a <=( a98568a  and  a98553a );
 a196a <=( a98538a  and  a98523a );
 a197a <=( a98508a  and  a98493a );
 a198a <=( a98478a  and  a98463a );
 a199a <=( a98448a  and  a98433a );
 a200a <=( a98418a  and  a98403a );
 a201a <=( a98388a  and  a98373a );
 a202a <=( a98358a  and  a98343a );
 a203a <=( a98328a  and  a98313a );
 a204a <=( a98298a  and  a98283a );
 a205a <=( a98268a  and  a98253a );
 a206a <=( a98238a  and  a98223a );
 a207a <=( a98208a  and  a98193a );
 a208a <=( a98178a  and  a98163a );
 a209a <=( a98148a  and  a98133a );
 a210a <=( a98118a  and  a98103a );
 a211a <=( a98088a  and  a98073a );
 a212a <=( a98058a  and  a98043a );
 a213a <=( a98028a  and  a98013a );
 a214a <=( a97998a  and  a97983a );
 a215a <=( a97968a  and  a97953a );
 a216a <=( a97938a  and  a97923a );
 a217a <=( a97908a  and  a97893a );
 a218a <=( a97878a  and  a97863a );
 a219a <=( a97848a  and  a97833a );
 a220a <=( a97818a  and  a97803a );
 a221a <=( a97788a  and  a97773a );
 a222a <=( a97758a  and  a97743a );
 a223a <=( a97728a  and  a97713a );
 a224a <=( a97698a  and  a97683a );
 a225a <=( a97668a  and  a97653a );
 a226a <=( a97638a  and  a97623a );
 a227a <=( a97608a  and  a97593a );
 a228a <=( a97578a  and  a97563a );
 a229a <=( a97548a  and  a97533a );
 a230a <=( a97518a  and  a97503a );
 a231a <=( a97488a  and  a97473a );
 a232a <=( a97458a  and  a97443a );
 a233a <=( a97428a  and  a97413a );
 a234a <=( a97398a  and  a97383a );
 a235a <=( a97368a  and  a97353a );
 a236a <=( a97338a  and  a97323a );
 a237a <=( a97308a  and  a97293a );
 a238a <=( a97278a  and  a97263a );
 a239a <=( a97248a  and  a97233a );
 a240a <=( a97218a  and  a97203a );
 a241a <=( a97188a  and  a97173a );
 a242a <=( a97158a  and  a97143a );
 a243a <=( a97128a  and  a97113a );
 a244a <=( a97098a  and  a97083a );
 a245a <=( a97068a  and  a97053a );
 a246a <=( a97038a  and  a97023a );
 a247a <=( a97008a  and  a96993a );
 a248a <=( a96978a  and  a96963a );
 a249a <=( a96948a  and  a96933a );
 a250a <=( a96918a  and  a96903a );
 a251a <=( a96888a  and  a96873a );
 a252a <=( a96858a  and  a96843a );
 a253a <=( a96828a  and  a96813a );
 a254a <=( a96798a  and  a96783a );
 a255a <=( a96768a  and  a96753a );
 a256a <=( a96738a  and  a96723a );
 a257a <=( a96708a  and  a96693a );
 a258a <=( a96678a  and  a96663a );
 a259a <=( a96648a  and  a96633a );
 a260a <=( a96618a  and  a96603a );
 a261a <=( a96588a  and  a96573a );
 a262a <=( a96558a  and  a96543a );
 a263a <=( a96528a  and  a96513a );
 a264a <=( a96498a  and  a96483a );
 a265a <=( a96468a  and  a96453a );
 a266a <=( a96438a  and  a96423a );
 a267a <=( a96408a  and  a96393a );
 a268a <=( a96378a  and  a96363a );
 a269a <=( a96348a  and  a96333a );
 a270a <=( a96318a  and  a96303a );
 a271a <=( a96288a  and  a96273a );
 a272a <=( a96258a  and  a96243a );
 a273a <=( a96228a  and  a96213a );
 a274a <=( a96198a  and  a96183a );
 a275a <=( a96168a  and  a96153a );
 a276a <=( a96138a  and  a96123a );
 a277a <=( a96108a  and  a96093a );
 a278a <=( a96078a  and  a96063a );
 a279a <=( a96048a  and  a96033a );
 a280a <=( a96018a  and  a96003a );
 a281a <=( a95988a  and  a95973a );
 a282a <=( a95958a  and  a95943a );
 a283a <=( a95928a  and  a95913a );
 a284a <=( a95898a  and  a95883a );
 a285a <=( a95868a  and  a95853a );
 a286a <=( a95838a  and  a95823a );
 a287a <=( a95808a  and  a95793a );
 a288a <=( a95778a  and  a95763a );
 a289a <=( a95748a  and  a95733a );
 a290a <=( a95718a  and  a95703a );
 a291a <=( a95688a  and  a95673a );
 a292a <=( a95658a  and  a95643a );
 a293a <=( a95628a  and  a95613a );
 a294a <=( a95598a  and  a95583a );
 a295a <=( a95568a  and  a95553a );
 a296a <=( a95538a  and  a95523a );
 a297a <=( a95508a  and  a95493a );
 a298a <=( a95478a  and  a95463a );
 a299a <=( a95448a  and  a95433a );
 a300a <=( a95418a  and  a95403a );
 a301a <=( a95388a  and  a95373a );
 a302a <=( a95358a  and  a95343a );
 a303a <=( a95328a  and  a95313a );
 a304a <=( a95298a  and  a95283a );
 a305a <=( a95268a  and  a95253a );
 a306a <=( a95238a  and  a95223a );
 a307a <=( a95208a  and  a95193a );
 a308a <=( a95178a  and  a95163a );
 a309a <=( a95148a  and  a95133a );
 a310a <=( a95118a  and  a95103a );
 a311a <=( a95088a  and  a95073a );
 a312a <=( a95058a  and  a95043a );
 a313a <=( a95028a  and  a95013a );
 a314a <=( a94998a  and  a94983a );
 a315a <=( a94968a  and  a94953a );
 a316a <=( a94938a  and  a94923a );
 a317a <=( a94908a  and  a94893a );
 a318a <=( a94878a  and  a94863a );
 a319a <=( a94848a  and  a94833a );
 a320a <=( a94818a  and  a94803a );
 a321a <=( a94788a  and  a94773a );
 a322a <=( a94758a  and  a94743a );
 a323a <=( a94728a  and  a94713a );
 a324a <=( a94698a  and  a94683a );
 a325a <=( a94668a  and  a94653a );
 a326a <=( a94638a  and  a94623a );
 a327a <=( a94608a  and  a94593a );
 a328a <=( a94578a  and  a94563a );
 a329a <=( a94548a  and  a94533a );
 a330a <=( a94518a  and  a94503a );
 a331a <=( a94488a  and  a94473a );
 a332a <=( a94458a  and  a94443a );
 a333a <=( a94428a  and  a94413a );
 a334a <=( a94398a  and  a94383a );
 a335a <=( a94368a  and  a94353a );
 a336a <=( a94338a  and  a94323a );
 a337a <=( a94308a  and  a94293a );
 a338a <=( a94278a  and  a94263a );
 a339a <=( a94248a  and  a94233a );
 a340a <=( a94218a  and  a94203a );
 a341a <=( a94188a  and  a94173a );
 a342a <=( a94158a  and  a94143a );
 a343a <=( a94128a  and  a94113a );
 a344a <=( a94098a  and  a94083a );
 a345a <=( a94068a  and  a94053a );
 a346a <=( a94038a  and  a94023a );
 a347a <=( a94008a  and  a93993a );
 a348a <=( a93978a  and  a93963a );
 a349a <=( a93948a  and  a93933a );
 a350a <=( a93918a  and  a93903a );
 a351a <=( a93888a  and  a93873a );
 a352a <=( a93858a  and  a93843a );
 a353a <=( a93828a  and  a93813a );
 a354a <=( a93798a  and  a93783a );
 a355a <=( a93768a  and  a93753a );
 a356a <=( a93738a  and  a93723a );
 a357a <=( a93708a  and  a93693a );
 a358a <=( a93678a  and  a93663a );
 a359a <=( a93648a  and  a93633a );
 a360a <=( a93618a  and  a93603a );
 a361a <=( a93588a  and  a93573a );
 a362a <=( a93558a  and  a93543a );
 a363a <=( a93528a  and  a93513a );
 a364a <=( a93498a  and  a93483a );
 a365a <=( a93468a  and  a93453a );
 a366a <=( a93438a  and  a93423a );
 a367a <=( a93408a  and  a93393a );
 a368a <=( a93378a  and  a93363a );
 a369a <=( a93348a  and  a93333a );
 a370a <=( a93318a  and  a93303a );
 a371a <=( a93288a  and  a93273a );
 a372a <=( a93258a  and  a93243a );
 a373a <=( a93228a  and  a93213a );
 a374a <=( a93198a  and  a93183a );
 a375a <=( a93168a  and  a93153a );
 a376a <=( a93138a  and  a93123a );
 a377a <=( a93108a  and  a93093a );
 a378a <=( a93078a  and  a93063a );
 a379a <=( a93048a  and  a93033a );
 a380a <=( a93018a  and  a93003a );
 a381a <=( a92988a  and  a92973a );
 a382a <=( a92958a  and  a92943a );
 a383a <=( a92928a  and  a92913a );
 a384a <=( a92898a  and  a92883a );
 a385a <=( a92868a  and  a92853a );
 a386a <=( a92840a  and  a92825a );
 a387a <=( a92812a  and  a92797a );
 a388a <=( a92784a  and  a92769a );
 a389a <=( a92756a  and  a92741a );
 a390a <=( a92728a  and  a92713a );
 a391a <=( a92700a  and  a92685a );
 a392a <=( a92672a  and  a92657a );
 a393a <=( a92644a  and  a92629a );
 a394a <=( a92616a  and  a92601a );
 a395a <=( a92588a  and  a92573a );
 a396a <=( a92560a  and  a92545a );
 a397a <=( a92532a  and  a92517a );
 a398a <=( a92504a  and  a92489a );
 a399a <=( a92476a  and  a92461a );
 a400a <=( a92448a  and  a92433a );
 a401a <=( a92420a  and  a92405a );
 a402a <=( a92392a  and  a92377a );
 a403a <=( a92364a  and  a92349a );
 a404a <=( a92336a  and  a92321a );
 a405a <=( a92308a  and  a92293a );
 a406a <=( a92280a  and  a92265a );
 a407a <=( a92252a  and  a92237a );
 a408a <=( a92224a  and  a92209a );
 a409a <=( a92196a  and  a92181a );
 a410a <=( a92168a  and  a92153a );
 a411a <=( a92140a  and  a92125a );
 a412a <=( a92112a  and  a92097a );
 a413a <=( a92084a  and  a92069a );
 a414a <=( a92056a  and  a92041a );
 a415a <=( a92028a  and  a92013a );
 a416a <=( a92000a  and  a91985a );
 a417a <=( a91972a  and  a91957a );
 a418a <=( a91944a  and  a91929a );
 a419a <=( a91916a  and  a91901a );
 a420a <=( a91888a  and  a91873a );
 a421a <=( a91860a  and  a91845a );
 a422a <=( a91832a  and  a91817a );
 a423a <=( a91804a  and  a91789a );
 a424a <=( a91776a  and  a91761a );
 a425a <=( a91748a  and  a91733a );
 a426a <=( a91720a  and  a91705a );
 a427a <=( a91692a  and  a91677a );
 a428a <=( a91664a  and  a91649a );
 a429a <=( a91636a  and  a91621a );
 a430a <=( a91608a  and  a91593a );
 a431a <=( a91580a  and  a91565a );
 a432a <=( a91552a  and  a91537a );
 a433a <=( a91524a  and  a91509a );
 a434a <=( a91496a  and  a91481a );
 a435a <=( a91468a  and  a91453a );
 a436a <=( a91440a  and  a91425a );
 a437a <=( a91412a  and  a91397a );
 a438a <=( a91384a  and  a91369a );
 a439a <=( a91356a  and  a91341a );
 a440a <=( a91328a  and  a91313a );
 a441a <=( a91300a  and  a91285a );
 a442a <=( a91272a  and  a91257a );
 a443a <=( a91244a  and  a91229a );
 a444a <=( a91216a  and  a91201a );
 a445a <=( a91188a  and  a91173a );
 a446a <=( a91160a  and  a91145a );
 a447a <=( a91132a  and  a91117a );
 a448a <=( a91104a  and  a91089a );
 a449a <=( a91076a  and  a91061a );
 a450a <=( a91048a  and  a91033a );
 a451a <=( a91020a  and  a91005a );
 a452a <=( a90992a  and  a90977a );
 a453a <=( a90964a  and  a90949a );
 a454a <=( a90936a  and  a90921a );
 a455a <=( a90908a  and  a90893a );
 a456a <=( a90880a  and  a90865a );
 a457a <=( a90852a  and  a90837a );
 a458a <=( a90824a  and  a90809a );
 a459a <=( a90796a  and  a90781a );
 a460a <=( a90768a  and  a90753a );
 a461a <=( a90740a  and  a90725a );
 a462a <=( a90712a  and  a90697a );
 a463a <=( a90684a  and  a90669a );
 a464a <=( a90656a  and  a90641a );
 a465a <=( a90628a  and  a90613a );
 a466a <=( a90600a  and  a90585a );
 a467a <=( a90572a  and  a90557a );
 a468a <=( a90544a  and  a90529a );
 a469a <=( a90516a  and  a90501a );
 a470a <=( a90488a  and  a90473a );
 a471a <=( a90460a  and  a90445a );
 a472a <=( a90432a  and  a90417a );
 a473a <=( a90404a  and  a90389a );
 a474a <=( a90376a  and  a90361a );
 a475a <=( a90348a  and  a90333a );
 a476a <=( a90320a  and  a90305a );
 a477a <=( a90292a  and  a90277a );
 a478a <=( a90264a  and  a90249a );
 a479a <=( a90236a  and  a90221a );
 a480a <=( a90208a  and  a90193a );
 a481a <=( a90180a  and  a90165a );
 a482a <=( a90152a  and  a90137a );
 a483a <=( a90124a  and  a90109a );
 a484a <=( a90096a  and  a90081a );
 a485a <=( a90068a  and  a90053a );
 a486a <=( a90040a  and  a90025a );
 a487a <=( a90012a  and  a89997a );
 a488a <=( a89984a  and  a89969a );
 a489a <=( a89956a  and  a89941a );
 a490a <=( a89928a  and  a89913a );
 a491a <=( a89900a  and  a89885a );
 a492a <=( a89872a  and  a89857a );
 a493a <=( a89844a  and  a89829a );
 a494a <=( a89816a  and  a89801a );
 a495a <=( a89788a  and  a89773a );
 a496a <=( a89760a  and  a89745a );
 a497a <=( a89732a  and  a89717a );
 a498a <=( a89704a  and  a89689a );
 a499a <=( a89676a  and  a89661a );
 a500a <=( a89648a  and  a89633a );
 a501a <=( a89620a  and  a89605a );
 a502a <=( a89592a  and  a89577a );
 a503a <=( a89564a  and  a89549a );
 a504a <=( a89536a  and  a89521a );
 a505a <=( a89508a  and  a89493a );
 a506a <=( a89480a  and  a89465a );
 a507a <=( a89452a  and  a89437a );
 a508a <=( a89424a  and  a89409a );
 a509a <=( a89396a  and  a89381a );
 a510a <=( a89368a  and  a89353a );
 a511a <=( a89340a  and  a89325a );
 a512a <=( a89312a  and  a89297a );
 a513a <=( a89284a  and  a89269a );
 a514a <=( a89256a  and  a89241a );
 a515a <=( a89228a  and  a89213a );
 a516a <=( a89200a  and  a89185a );
 a517a <=( a89172a  and  a89157a );
 a518a <=( a89144a  and  a89129a );
 a519a <=( a89116a  and  a89101a );
 a520a <=( a89088a  and  a89073a );
 a521a <=( a89060a  and  a89045a );
 a522a <=( a89032a  and  a89017a );
 a523a <=( a89004a  and  a88989a );
 a524a <=( a88976a  and  a88961a );
 a525a <=( a88948a  and  a88933a );
 a526a <=( a88920a  and  a88905a );
 a527a <=( a88892a  and  a88877a );
 a528a <=( a88864a  and  a88849a );
 a529a <=( a88836a  and  a88821a );
 a530a <=( a88808a  and  a88793a );
 a531a <=( a88780a  and  a88765a );
 a532a <=( a88752a  and  a88737a );
 a533a <=( a88724a  and  a88709a );
 a534a <=( a88696a  and  a88681a );
 a535a <=( a88668a  and  a88653a );
 a536a <=( a88640a  and  a88625a );
 a537a <=( a88612a  and  a88597a );
 a538a <=( a88584a  and  a88569a );
 a539a <=( a88556a  and  a88541a );
 a540a <=( a88528a  and  a88513a );
 a541a <=( a88500a  and  a88485a );
 a542a <=( a88472a  and  a88457a );
 a543a <=( a88444a  and  a88429a );
 a544a <=( a88416a  and  a88401a );
 a545a <=( a88388a  and  a88373a );
 a546a <=( a88360a  and  a88345a );
 a547a <=( a88332a  and  a88317a );
 a548a <=( a88304a  and  a88289a );
 a549a <=( a88276a  and  a88261a );
 a550a <=( a88248a  and  a88233a );
 a551a <=( a88220a  and  a88205a );
 a552a <=( a88192a  and  a88177a );
 a553a <=( a88164a  and  a88149a );
 a554a <=( a88136a  and  a88121a );
 a555a <=( a88108a  and  a88093a );
 a556a <=( a88080a  and  a88065a );
 a557a <=( a88052a  and  a88037a );
 a558a <=( a88024a  and  a88009a );
 a559a <=( a87996a  and  a87981a );
 a560a <=( a87968a  and  a87953a );
 a561a <=( a87940a  and  a87925a );
 a562a <=( a87912a  and  a87897a );
 a563a <=( a87884a  and  a87869a );
 a564a <=( a87856a  and  a87841a );
 a565a <=( a87828a  and  a87813a );
 a566a <=( a87800a  and  a87785a );
 a567a <=( a87772a  and  a87757a );
 a568a <=( a87744a  and  a87729a );
 a569a <=( a87716a  and  a87701a );
 a570a <=( a87688a  and  a87673a );
 a571a <=( a87660a  and  a87645a );
 a572a <=( a87632a  and  a87617a );
 a573a <=( a87604a  and  a87589a );
 a574a <=( a87576a  and  a87561a );
 a575a <=( a87548a  and  a87533a );
 a576a <=( a87520a  and  a87505a );
 a577a <=( a87492a  and  a87477a );
 a578a <=( a87464a  and  a87449a );
 a579a <=( a87436a  and  a87421a );
 a580a <=( a87408a  and  a87393a );
 a581a <=( a87380a  and  a87365a );
 a582a <=( a87352a  and  a87337a );
 a583a <=( a87324a  and  a87309a );
 a584a <=( a87296a  and  a87281a );
 a585a <=( a87268a  and  a87253a );
 a586a <=( a87240a  and  a87225a );
 a587a <=( a87212a  and  a87197a );
 a588a <=( a87184a  and  a87169a );
 a589a <=( a87156a  and  a87141a );
 a590a <=( a87128a  and  a87113a );
 a591a <=( a87100a  and  a87085a );
 a592a <=( a87072a  and  a87057a );
 a593a <=( a87044a  and  a87029a );
 a594a <=( a87016a  and  a87001a );
 a595a <=( a86988a  and  a86973a );
 a596a <=( a86960a  and  a86945a );
 a597a <=( a86932a  and  a86917a );
 a598a <=( a86904a  and  a86889a );
 a599a <=( a86876a  and  a86861a );
 a600a <=( a86848a  and  a86833a );
 a601a <=( a86820a  and  a86805a );
 a602a <=( a86792a  and  a86777a );
 a603a <=( a86764a  and  a86749a );
 a604a <=( a86736a  and  a86721a );
 a605a <=( a86708a  and  a86693a );
 a606a <=( a86680a  and  a86665a );
 a607a <=( a86652a  and  a86637a );
 a608a <=( a86624a  and  a86609a );
 a609a <=( a86596a  and  a86581a );
 a610a <=( a86568a  and  a86553a );
 a611a <=( a86540a  and  a86525a );
 a612a <=( a86512a  and  a86497a );
 a613a <=( a86484a  and  a86469a );
 a614a <=( a86456a  and  a86441a );
 a615a <=( a86428a  and  a86413a );
 a616a <=( a86400a  and  a86385a );
 a617a <=( a86372a  and  a86357a );
 a618a <=( a86344a  and  a86329a );
 a619a <=( a86316a  and  a86301a );
 a620a <=( a86288a  and  a86273a );
 a621a <=( a86260a  and  a86245a );
 a622a <=( a86232a  and  a86217a );
 a623a <=( a86204a  and  a86189a );
 a624a <=( a86176a  and  a86161a );
 a625a <=( a86148a  and  a86133a );
 a626a <=( a86120a  and  a86105a );
 a627a <=( a86092a  and  a86077a );
 a628a <=( a86064a  and  a86049a );
 a629a <=( a86036a  and  a86021a );
 a630a <=( a86008a  and  a85993a );
 a631a <=( a85980a  and  a85965a );
 a632a <=( a85952a  and  a85937a );
 a633a <=( a85924a  and  a85909a );
 a634a <=( a85896a  and  a85881a );
 a635a <=( a85868a  and  a85853a );
 a636a <=( a85840a  and  a85825a );
 a637a <=( a85812a  and  a85797a );
 a638a <=( a85784a  and  a85769a );
 a639a <=( a85756a  and  a85741a );
 a640a <=( a85728a  and  a85713a );
 a641a <=( a85700a  and  a85685a );
 a642a <=( a85672a  and  a85657a );
 a643a <=( a85644a  and  a85629a );
 a644a <=( a85616a  and  a85601a );
 a645a <=( a85588a  and  a85573a );
 a646a <=( a85560a  and  a85545a );
 a647a <=( a85532a  and  a85517a );
 a648a <=( a85504a  and  a85489a );
 a649a <=( a85476a  and  a85461a );
 a650a <=( a85448a  and  a85433a );
 a651a <=( a85420a  and  a85405a );
 a652a <=( a85392a  and  a85377a );
 a653a <=( a85364a  and  a85349a );
 a654a <=( a85336a  and  a85321a );
 a655a <=( a85308a  and  a85293a );
 a656a <=( a85280a  and  a85265a );
 a657a <=( a85252a  and  a85237a );
 a658a <=( a85224a  and  a85209a );
 a659a <=( a85196a  and  a85181a );
 a660a <=( a85168a  and  a85153a );
 a661a <=( a85140a  and  a85125a );
 a662a <=( a85112a  and  a85097a );
 a663a <=( a85084a  and  a85069a );
 a664a <=( a85056a  and  a85041a );
 a665a <=( a85028a  and  a85013a );
 a666a <=( a85000a  and  a84985a );
 a667a <=( a84972a  and  a84957a );
 a668a <=( a84944a  and  a84929a );
 a669a <=( a84916a  and  a84901a );
 a670a <=( a84888a  and  a84873a );
 a671a <=( a84860a  and  a84845a );
 a672a <=( a84832a  and  a84817a );
 a673a <=( a84804a  and  a84789a );
 a674a <=( a84776a  and  a84761a );
 a675a <=( a84748a  and  a84733a );
 a676a <=( a84720a  and  a84705a );
 a677a <=( a84692a  and  a84677a );
 a678a <=( a84664a  and  a84649a );
 a679a <=( a84636a  and  a84621a );
 a680a <=( a84608a  and  a84593a );
 a681a <=( a84580a  and  a84565a );
 a682a <=( a84552a  and  a84537a );
 a683a <=( a84524a  and  a84509a );
 a684a <=( a84496a  and  a84481a );
 a685a <=( a84468a  and  a84453a );
 a686a <=( a84440a  and  a84425a );
 a687a <=( a84412a  and  a84397a );
 a688a <=( a84384a  and  a84369a );
 a689a <=( a84356a  and  a84341a );
 a690a <=( a84328a  and  a84313a );
 a691a <=( a84300a  and  a84285a );
 a692a <=( a84272a  and  a84257a );
 a693a <=( a84244a  and  a84229a );
 a694a <=( a84216a  and  a84201a );
 a695a <=( a84188a  and  a84173a );
 a696a <=( a84160a  and  a84145a );
 a697a <=( a84132a  and  a84117a );
 a698a <=( a84104a  and  a84089a );
 a699a <=( a84076a  and  a84061a );
 a700a <=( a84048a  and  a84033a );
 a701a <=( a84020a  and  a84005a );
 a702a <=( a83992a  and  a83977a );
 a703a <=( a83964a  and  a83949a );
 a704a <=( a83936a  and  a83921a );
 a705a <=( a83908a  and  a83893a );
 a706a <=( a83880a  and  a83865a );
 a707a <=( a83852a  and  a83837a );
 a708a <=( a83824a  and  a83809a );
 a709a <=( a83796a  and  a83781a );
 a710a <=( a83768a  and  a83753a );
 a711a <=( a83740a  and  a83725a );
 a712a <=( a83712a  and  a83697a );
 a713a <=( a83684a  and  a83669a );
 a714a <=( a83656a  and  a83641a );
 a715a <=( a83628a  and  a83613a );
 a716a <=( a83600a  and  a83585a );
 a717a <=( a83572a  and  a83557a );
 a718a <=( a83544a  and  a83529a );
 a719a <=( a83516a  and  a83501a );
 a720a <=( a83488a  and  a83473a );
 a721a <=( a83460a  and  a83445a );
 a722a <=( a83432a  and  a83417a );
 a723a <=( a83404a  and  a83389a );
 a724a <=( a83376a  and  a83361a );
 a725a <=( a83348a  and  a83333a );
 a726a <=( a83320a  and  a83305a );
 a727a <=( a83292a  and  a83277a );
 a728a <=( a83264a  and  a83249a );
 a729a <=( a83236a  and  a83221a );
 a730a <=( a83208a  and  a83193a );
 a731a <=( a83180a  and  a83165a );
 a732a <=( a83152a  and  a83137a );
 a733a <=( a83124a  and  a83109a );
 a734a <=( a83096a  and  a83081a );
 a735a <=( a83068a  and  a83053a );
 a736a <=( a83040a  and  a83025a );
 a737a <=( a83012a  and  a82997a );
 a738a <=( a82984a  and  a82969a );
 a739a <=( a82956a  and  a82941a );
 a740a <=( a82928a  and  a82913a );
 a741a <=( a82900a  and  a82885a );
 a742a <=( a82872a  and  a82857a );
 a743a <=( a82844a  and  a82829a );
 a744a <=( a82816a  and  a82801a );
 a745a <=( a82788a  and  a82773a );
 a746a <=( a82760a  and  a82745a );
 a747a <=( a82732a  and  a82717a );
 a748a <=( a82704a  and  a82689a );
 a749a <=( a82676a  and  a82661a );
 a750a <=( a82648a  and  a82633a );
 a751a <=( a82620a  and  a82605a );
 a752a <=( a82592a  and  a82577a );
 a753a <=( a82564a  and  a82549a );
 a754a <=( a82536a  and  a82521a );
 a755a <=( a82508a  and  a82493a );
 a756a <=( a82480a  and  a82465a );
 a757a <=( a82452a  and  a82437a );
 a758a <=( a82424a  and  a82409a );
 a759a <=( a82396a  and  a82381a );
 a760a <=( a82368a  and  a82353a );
 a761a <=( a82340a  and  a82325a );
 a762a <=( a82312a  and  a82297a );
 a763a <=( a82284a  and  a82269a );
 a764a <=( a82256a  and  a82241a );
 a765a <=( a82228a  and  a82213a );
 a766a <=( a82200a  and  a82185a );
 a767a <=( a82172a  and  a82157a );
 a768a <=( a82144a  and  a82129a );
 a769a <=( a82116a  and  a82101a );
 a770a <=( a82088a  and  a82073a );
 a771a <=( a82060a  and  a82045a );
 a772a <=( a82032a  and  a82017a );
 a773a <=( a82004a  and  a81989a );
 a774a <=( a81976a  and  a81961a );
 a775a <=( a81948a  and  a81933a );
 a776a <=( a81920a  and  a81905a );
 a777a <=( a81892a  and  a81877a );
 a778a <=( a81864a  and  a81849a );
 a779a <=( a81836a  and  a81821a );
 a780a <=( a81808a  and  a81793a );
 a781a <=( a81780a  and  a81765a );
 a782a <=( a81752a  and  a81737a );
 a783a <=( a81724a  and  a81709a );
 a784a <=( a81696a  and  a81681a );
 a785a <=( a81668a  and  a81653a );
 a786a <=( a81640a  and  a81625a );
 a787a <=( a81612a  and  a81597a );
 a788a <=( a81584a  and  a81569a );
 a789a <=( a81556a  and  a81541a );
 a790a <=( a81528a  and  a81513a );
 a791a <=( a81500a  and  a81485a );
 a792a <=( a81472a  and  a81457a );
 a793a <=( a81444a  and  a81429a );
 a794a <=( a81416a  and  a81401a );
 a795a <=( a81388a  and  a81373a );
 a796a <=( a81360a  and  a81345a );
 a797a <=( a81332a  and  a81317a );
 a798a <=( a81304a  and  a81289a );
 a799a <=( a81276a  and  a81261a );
 a800a <=( a81248a  and  a81233a );
 a801a <=( a81220a  and  a81205a );
 a802a <=( a81192a  and  a81177a );
 a803a <=( a81164a  and  a81149a );
 a804a <=( a81136a  and  a81121a );
 a805a <=( a81108a  and  a81093a );
 a806a <=( a81080a  and  a81065a );
 a807a <=( a81052a  and  a81037a );
 a808a <=( a81024a  and  a81009a );
 a809a <=( a80996a  and  a80981a );
 a810a <=( a80968a  and  a80953a );
 a811a <=( a80940a  and  a80925a );
 a812a <=( a80912a  and  a80897a );
 a813a <=( a80884a  and  a80869a );
 a814a <=( a80856a  and  a80841a );
 a815a <=( a80828a  and  a80813a );
 a816a <=( a80800a  and  a80785a );
 a817a <=( a80772a  and  a80757a );
 a818a <=( a80744a  and  a80729a );
 a819a <=( a80716a  and  a80701a );
 a820a <=( a80688a  and  a80673a );
 a821a <=( a80660a  and  a80645a );
 a822a <=( a80632a  and  a80617a );
 a823a <=( a80604a  and  a80589a );
 a824a <=( a80576a  and  a80561a );
 a825a <=( a80548a  and  a80533a );
 a826a <=( a80520a  and  a80505a );
 a827a <=( a80492a  and  a80477a );
 a828a <=( a80464a  and  a80449a );
 a829a <=( a80436a  and  a80421a );
 a830a <=( a80408a  and  a80393a );
 a831a <=( a80380a  and  a80365a );
 a832a <=( a80352a  and  a80337a );
 a833a <=( a80324a  and  a80309a );
 a834a <=( a80296a  and  a80281a );
 a835a <=( a80268a  and  a80253a );
 a836a <=( a80240a  and  a80225a );
 a837a <=( a80212a  and  a80197a );
 a838a <=( a80184a  and  a80169a );
 a839a <=( a80156a  and  a80141a );
 a840a <=( a80128a  and  a80113a );
 a841a <=( a80100a  and  a80085a );
 a842a <=( a80072a  and  a80057a );
 a843a <=( a80044a  and  a80029a );
 a844a <=( a80016a  and  a80001a );
 a845a <=( a79988a  and  a79973a );
 a846a <=( a79960a  and  a79945a );
 a847a <=( a79932a  and  a79917a );
 a848a <=( a79904a  and  a79889a );
 a849a <=( a79876a  and  a79861a );
 a850a <=( a79848a  and  a79833a );
 a851a <=( a79820a  and  a79805a );
 a852a <=( a79792a  and  a79777a );
 a853a <=( a79764a  and  a79749a );
 a854a <=( a79736a  and  a79721a );
 a855a <=( a79708a  and  a79693a );
 a856a <=( a79680a  and  a79665a );
 a857a <=( a79652a  and  a79637a );
 a858a <=( a79624a  and  a79609a );
 a859a <=( a79596a  and  a79581a );
 a860a <=( a79568a  and  a79553a );
 a861a <=( a79540a  and  a79525a );
 a862a <=( a79512a  and  a79497a );
 a863a <=( a79484a  and  a79469a );
 a864a <=( a79456a  and  a79441a );
 a865a <=( a79428a  and  a79413a );
 a866a <=( a79400a  and  a79385a );
 a867a <=( a79372a  and  a79357a );
 a868a <=( a79344a  and  a79329a );
 a869a <=( a79316a  and  a79301a );
 a870a <=( a79288a  and  a79273a );
 a871a <=( a79260a  and  a79245a );
 a872a <=( a79232a  and  a79217a );
 a873a <=( a79204a  and  a79189a );
 a874a <=( a79176a  and  a79161a );
 a875a <=( a79148a  and  a79133a );
 a876a <=( a79120a  and  a79105a );
 a877a <=( a79092a  and  a79077a );
 a878a <=( a79064a  and  a79049a );
 a879a <=( a79036a  and  a79021a );
 a880a <=( a79008a  and  a78993a );
 a881a <=( a78980a  and  a78965a );
 a882a <=( a78952a  and  a78937a );
 a883a <=( a78924a  and  a78909a );
 a884a <=( a78896a  and  a78881a );
 a885a <=( a78868a  and  a78853a );
 a886a <=( a78840a  and  a78825a );
 a887a <=( a78812a  and  a78797a );
 a888a <=( a78784a  and  a78769a );
 a889a <=( a78756a  and  a78741a );
 a890a <=( a78728a  and  a78713a );
 a891a <=( a78700a  and  a78685a );
 a892a <=( a78672a  and  a78657a );
 a893a <=( a78644a  and  a78629a );
 a894a <=( a78616a  and  a78601a );
 a895a <=( a78588a  and  a78573a );
 a896a <=( a78560a  and  a78545a );
 a897a <=( a78532a  and  a78517a );
 a898a <=( a78504a  and  a78489a );
 a899a <=( a78476a  and  a78461a );
 a900a <=( a78448a  and  a78433a );
 a901a <=( a78420a  and  a78405a );
 a902a <=( a78392a  and  a78377a );
 a903a <=( a78364a  and  a78349a );
 a904a <=( a78336a  and  a78321a );
 a905a <=( a78308a  and  a78293a );
 a906a <=( a78280a  and  a78265a );
 a907a <=( a78252a  and  a78237a );
 a908a <=( a78224a  and  a78209a );
 a909a <=( a78196a  and  a78181a );
 a910a <=( a78168a  and  a78153a );
 a911a <=( a78140a  and  a78125a );
 a912a <=( a78112a  and  a78097a );
 a913a <=( a78084a  and  a78069a );
 a914a <=( a78056a  and  a78041a );
 a915a <=( a78028a  and  a78013a );
 a916a <=( a78000a  and  a77985a );
 a917a <=( a77972a  and  a77957a );
 a918a <=( a77944a  and  a77929a );
 a919a <=( a77916a  and  a77901a );
 a920a <=( a77888a  and  a77873a );
 a921a <=( a77860a  and  a77845a );
 a922a <=( a77832a  and  a77817a );
 a923a <=( a77804a  and  a77789a );
 a924a <=( a77776a  and  a77761a );
 a925a <=( a77748a  and  a77733a );
 a926a <=( a77720a  and  a77705a );
 a927a <=( a77692a  and  a77677a );
 a928a <=( a77664a  and  a77649a );
 a929a <=( a77636a  and  a77623a );
 a930a <=( a77610a  and  a77597a );
 a931a <=( a77584a  and  a77571a );
 a932a <=( a77558a  and  a77545a );
 a933a <=( a77532a  and  a77519a );
 a934a <=( a77506a  and  a77493a );
 a935a <=( a77480a  and  a77467a );
 a936a <=( a77454a  and  a77441a );
 a937a <=( a77428a  and  a77415a );
 a938a <=( a77402a  and  a77389a );
 a939a <=( a77376a  and  a77363a );
 a940a <=( a77350a  and  a77337a );
 a941a <=( a77324a  and  a77311a );
 a942a <=( a77298a  and  a77285a );
 a943a <=( a77272a  and  a77259a );
 a944a <=( a77246a  and  a77233a );
 a945a <=( a77220a  and  a77207a );
 a946a <=( a77194a  and  a77181a );
 a947a <=( a77168a  and  a77155a );
 a948a <=( a77142a  and  a77129a );
 a949a <=( a77116a  and  a77103a );
 a950a <=( a77090a  and  a77077a );
 a951a <=( a77064a  and  a77051a );
 a952a <=( a77038a  and  a77025a );
 a953a <=( a77012a  and  a76999a );
 a954a <=( a76986a  and  a76973a );
 a955a <=( a76960a  and  a76947a );
 a956a <=( a76934a  and  a76921a );
 a957a <=( a76908a  and  a76895a );
 a958a <=( a76882a  and  a76869a );
 a959a <=( a76856a  and  a76843a );
 a960a <=( a76830a  and  a76817a );
 a961a <=( a76804a  and  a76791a );
 a962a <=( a76778a  and  a76765a );
 a963a <=( a76752a  and  a76739a );
 a964a <=( a76726a  and  a76713a );
 a965a <=( a76700a  and  a76687a );
 a966a <=( a76674a  and  a76661a );
 a967a <=( a76648a  and  a76635a );
 a968a <=( a76622a  and  a76609a );
 a969a <=( a76596a  and  a76583a );
 a970a <=( a76570a  and  a76557a );
 a971a <=( a76544a  and  a76531a );
 a972a <=( a76518a  and  a76505a );
 a973a <=( a76492a  and  a76479a );
 a974a <=( a76466a  and  a76453a );
 a975a <=( a76440a  and  a76427a );
 a976a <=( a76414a  and  a76401a );
 a977a <=( a76388a  and  a76375a );
 a978a <=( a76362a  and  a76349a );
 a979a <=( a76336a  and  a76323a );
 a980a <=( a76310a  and  a76297a );
 a981a <=( a76284a  and  a76271a );
 a982a <=( a76258a  and  a76245a );
 a983a <=( a76232a  and  a76219a );
 a984a <=( a76206a  and  a76193a );
 a985a <=( a76180a  and  a76167a );
 a986a <=( a76154a  and  a76141a );
 a987a <=( a76128a  and  a76115a );
 a988a <=( a76102a  and  a76089a );
 a989a <=( a76076a  and  a76063a );
 a990a <=( a76050a  and  a76037a );
 a991a <=( a76024a  and  a76011a );
 a992a <=( a75998a  and  a75985a );
 a993a <=( a75972a  and  a75959a );
 a994a <=( a75946a  and  a75933a );
 a995a <=( a75920a  and  a75907a );
 a996a <=( a75894a  and  a75881a );
 a997a <=( a75868a  and  a75855a );
 a998a <=( a75842a  and  a75829a );
 a999a <=( a75816a  and  a75803a );
 a1000a <=( a75790a  and  a75777a );
 a1001a <=( a75764a  and  a75751a );
 a1002a <=( a75738a  and  a75725a );
 a1003a <=( a75712a  and  a75699a );
 a1004a <=( a75686a  and  a75673a );
 a1005a <=( a75660a  and  a75647a );
 a1006a <=( a75634a  and  a75621a );
 a1007a <=( a75608a  and  a75595a );
 a1008a <=( a75582a  and  a75569a );
 a1009a <=( a75556a  and  a75543a );
 a1010a <=( a75530a  and  a75517a );
 a1011a <=( a75504a  and  a75491a );
 a1012a <=( a75478a  and  a75465a );
 a1013a <=( a75452a  and  a75439a );
 a1014a <=( a75426a  and  a75413a );
 a1015a <=( a75400a  and  a75387a );
 a1016a <=( a75374a  and  a75361a );
 a1017a <=( a75348a  and  a75335a );
 a1018a <=( a75322a  and  a75309a );
 a1019a <=( a75296a  and  a75283a );
 a1020a <=( a75270a  and  a75257a );
 a1021a <=( a75244a  and  a75231a );
 a1022a <=( a75218a  and  a75205a );
 a1023a <=( a75192a  and  a75179a );
 a1024a <=( a75166a  and  a75153a );
 a1025a <=( a75140a  and  a75127a );
 a1026a <=( a75114a  and  a75101a );
 a1027a <=( a75088a  and  a75075a );
 a1028a <=( a75062a  and  a75049a );
 a1029a <=( a75036a  and  a75023a );
 a1030a <=( a75010a  and  a74997a );
 a1031a <=( a74984a  and  a74971a );
 a1032a <=( a74958a  and  a74945a );
 a1033a <=( a74932a  and  a74919a );
 a1034a <=( a74906a  and  a74893a );
 a1035a <=( a74880a  and  a74867a );
 a1036a <=( a74854a  and  a74841a );
 a1037a <=( a74828a  and  a74815a );
 a1038a <=( a74802a  and  a74789a );
 a1039a <=( a74776a  and  a74763a );
 a1040a <=( a74750a  and  a74737a );
 a1041a <=( a74724a  and  a74711a );
 a1042a <=( a74698a  and  a74685a );
 a1043a <=( a74672a  and  a74659a );
 a1044a <=( a74646a  and  a74633a );
 a1045a <=( a74620a  and  a74607a );
 a1046a <=( a74594a  and  a74581a );
 a1047a <=( a74568a  and  a74555a );
 a1048a <=( a74542a  and  a74529a );
 a1049a <=( a74516a  and  a74503a );
 a1050a <=( a74490a  and  a74477a );
 a1051a <=( a74464a  and  a74451a );
 a1052a <=( a74438a  and  a74425a );
 a1053a <=( a74412a  and  a74399a );
 a1054a <=( a74386a  and  a74373a );
 a1055a <=( a74360a  and  a74347a );
 a1056a <=( a74334a  and  a74321a );
 a1057a <=( a74308a  and  a74295a );
 a1058a <=( a74282a  and  a74269a );
 a1059a <=( a74256a  and  a74243a );
 a1060a <=( a74230a  and  a74217a );
 a1061a <=( a74204a  and  a74191a );
 a1062a <=( a74178a  and  a74165a );
 a1063a <=( a74152a  and  a74139a );
 a1064a <=( a74126a  and  a74113a );
 a1065a <=( a74100a  and  a74087a );
 a1066a <=( a74074a  and  a74061a );
 a1067a <=( a74048a  and  a74035a );
 a1068a <=( a74022a  and  a74009a );
 a1069a <=( a73996a  and  a73983a );
 a1070a <=( a73970a  and  a73957a );
 a1071a <=( a73944a  and  a73931a );
 a1072a <=( a73918a  and  a73905a );
 a1073a <=( a73892a  and  a73879a );
 a1074a <=( a73866a  and  a73853a );
 a1075a <=( a73840a  and  a73827a );
 a1076a <=( a73814a  and  a73801a );
 a1077a <=( a73788a  and  a73775a );
 a1078a <=( a73762a  and  a73749a );
 a1079a <=( a73736a  and  a73723a );
 a1080a <=( a73710a  and  a73697a );
 a1081a <=( a73684a  and  a73671a );
 a1082a <=( a73658a  and  a73645a );
 a1083a <=( a73632a  and  a73619a );
 a1084a <=( a73606a  and  a73593a );
 a1085a <=( a73580a  and  a73567a );
 a1086a <=( a73554a  and  a73541a );
 a1087a <=( a73528a  and  a73515a );
 a1088a <=( a73502a  and  a73489a );
 a1089a <=( a73476a  and  a73463a );
 a1090a <=( a73450a  and  a73437a );
 a1091a <=( a73424a  and  a73411a );
 a1092a <=( a73398a  and  a73385a );
 a1093a <=( a73372a  and  a73359a );
 a1094a <=( a73346a  and  a73333a );
 a1095a <=( a73320a  and  a73307a );
 a1096a <=( a73294a  and  a73281a );
 a1097a <=( a73268a  and  a73255a );
 a1098a <=( a73242a  and  a73229a );
 a1099a <=( a73216a  and  a73203a );
 a1100a <=( a73190a  and  a73177a );
 a1101a <=( a73164a  and  a73151a );
 a1102a <=( a73138a  and  a73125a );
 a1103a <=( a73112a  and  a73099a );
 a1104a <=( a73086a  and  a73073a );
 a1105a <=( a73060a  and  a73047a );
 a1106a <=( a73034a  and  a73021a );
 a1107a <=( a73008a  and  a72995a );
 a1108a <=( a72982a  and  a72969a );
 a1109a <=( a72956a  and  a72943a );
 a1110a <=( a72930a  and  a72917a );
 a1111a <=( a72904a  and  a72891a );
 a1112a <=( a72878a  and  a72865a );
 a1113a <=( a72852a  and  a72839a );
 a1114a <=( a72826a  and  a72813a );
 a1115a <=( a72800a  and  a72787a );
 a1116a <=( a72774a  and  a72761a );
 a1117a <=( a72748a  and  a72735a );
 a1118a <=( a72722a  and  a72709a );
 a1119a <=( a72696a  and  a72683a );
 a1120a <=( a72670a  and  a72657a );
 a1121a <=( a72644a  and  a72631a );
 a1122a <=( a72618a  and  a72605a );
 a1123a <=( a72592a  and  a72579a );
 a1124a <=( a72566a  and  a72553a );
 a1125a <=( a72540a  and  a72527a );
 a1126a <=( a72514a  and  a72501a );
 a1127a <=( a72488a  and  a72475a );
 a1128a <=( a72462a  and  a72449a );
 a1129a <=( a72436a  and  a72423a );
 a1130a <=( a72410a  and  a72397a );
 a1131a <=( a72384a  and  a72371a );
 a1132a <=( a72358a  and  a72345a );
 a1133a <=( a72332a  and  a72319a );
 a1134a <=( a72306a  and  a72293a );
 a1135a <=( a72280a  and  a72267a );
 a1136a <=( a72254a  and  a72241a );
 a1137a <=( a72228a  and  a72215a );
 a1138a <=( a72202a  and  a72189a );
 a1139a <=( a72176a  and  a72163a );
 a1140a <=( a72150a  and  a72137a );
 a1141a <=( a72124a  and  a72111a );
 a1142a <=( a72098a  and  a72085a );
 a1143a <=( a72072a  and  a72059a );
 a1144a <=( a72046a  and  a72033a );
 a1145a <=( a72020a  and  a72007a );
 a1146a <=( a71994a  and  a71981a );
 a1147a <=( a71968a  and  a71955a );
 a1148a <=( a71942a  and  a71929a );
 a1149a <=( a71916a  and  a71903a );
 a1150a <=( a71890a  and  a71877a );
 a1151a <=( a71864a  and  a71851a );
 a1152a <=( a71838a  and  a71825a );
 a1153a <=( a71812a  and  a71799a );
 a1154a <=( a71786a  and  a71773a );
 a1155a <=( a71760a  and  a71747a );
 a1156a <=( a71734a  and  a71721a );
 a1157a <=( a71708a  and  a71695a );
 a1158a <=( a71682a  and  a71669a );
 a1159a <=( a71656a  and  a71643a );
 a1160a <=( a71630a  and  a71617a );
 a1161a <=( a71604a  and  a71591a );
 a1162a <=( a71578a  and  a71565a );
 a1163a <=( a71552a  and  a71539a );
 a1164a <=( a71526a  and  a71513a );
 a1165a <=( a71500a  and  a71487a );
 a1166a <=( a71474a  and  a71461a );
 a1167a <=( a71448a  and  a71435a );
 a1168a <=( a71422a  and  a71409a );
 a1169a <=( a71396a  and  a71383a );
 a1170a <=( a71370a  and  a71357a );
 a1171a <=( a71344a  and  a71331a );
 a1172a <=( a71318a  and  a71305a );
 a1173a <=( a71292a  and  a71279a );
 a1174a <=( a71266a  and  a71253a );
 a1175a <=( a71240a  and  a71227a );
 a1176a <=( a71214a  and  a71201a );
 a1177a <=( a71188a  and  a71175a );
 a1178a <=( a71162a  and  a71149a );
 a1179a <=( a71136a  and  a71123a );
 a1180a <=( a71110a  and  a71097a );
 a1181a <=( a71084a  and  a71071a );
 a1182a <=( a71058a  and  a71045a );
 a1183a <=( a71032a  and  a71019a );
 a1184a <=( a71006a  and  a70993a );
 a1185a <=( a70980a  and  a70967a );
 a1186a <=( a70954a  and  a70941a );
 a1187a <=( a70928a  and  a70915a );
 a1188a <=( a70902a  and  a70889a );
 a1189a <=( a70876a  and  a70863a );
 a1190a <=( a70850a  and  a70837a );
 a1191a <=( a70824a  and  a70811a );
 a1192a <=( a70798a  and  a70785a );
 a1193a <=( a70772a  and  a70759a );
 a1194a <=( a70746a  and  a70733a );
 a1195a <=( a70720a  and  a70707a );
 a1196a <=( a70694a  and  a70681a );
 a1197a <=( a70668a  and  a70655a );
 a1198a <=( a70642a  and  a70629a );
 a1199a <=( a70616a  and  a70603a );
 a1200a <=( a70590a  and  a70577a );
 a1201a <=( a70564a  and  a70551a );
 a1202a <=( a70538a  and  a70525a );
 a1203a <=( a70512a  and  a70499a );
 a1204a <=( a70486a  and  a70473a );
 a1205a <=( a70460a  and  a70447a );
 a1206a <=( a70434a  and  a70421a );
 a1207a <=( a70408a  and  a70395a );
 a1208a <=( a70382a  and  a70369a );
 a1209a <=( a70356a  and  a70343a );
 a1210a <=( a70330a  and  a70317a );
 a1211a <=( a70304a  and  a70291a );
 a1212a <=( a70278a  and  a70265a );
 a1213a <=( a70252a  and  a70239a );
 a1214a <=( a70226a  and  a70213a );
 a1215a <=( a70200a  and  a70187a );
 a1216a <=( a70174a  and  a70161a );
 a1217a <=( a70148a  and  a70135a );
 a1218a <=( a70122a  and  a70109a );
 a1219a <=( a70096a  and  a70083a );
 a1220a <=( a70070a  and  a70057a );
 a1221a <=( a70044a  and  a70031a );
 a1222a <=( a70018a  and  a70005a );
 a1223a <=( a69992a  and  a69979a );
 a1224a <=( a69966a  and  a69953a );
 a1225a <=( a69940a  and  a69927a );
 a1226a <=( a69914a  and  a69901a );
 a1227a <=( a69888a  and  a69875a );
 a1228a <=( a69862a  and  a69849a );
 a1229a <=( a69836a  and  a69823a );
 a1230a <=( a69810a  and  a69797a );
 a1231a <=( a69784a  and  a69771a );
 a1232a <=( a69758a  and  a69745a );
 a1233a <=( a69732a  and  a69719a );
 a1234a <=( a69706a  and  a69693a );
 a1235a <=( a69680a  and  a69667a );
 a1236a <=( a69654a  and  a69641a );
 a1237a <=( a69628a  and  a69615a );
 a1238a <=( a69602a  and  a69589a );
 a1239a <=( a69576a  and  a69563a );
 a1240a <=( a69550a  and  a69537a );
 a1241a <=( a69524a  and  a69511a );
 a1242a <=( a69498a  and  a69485a );
 a1243a <=( a69472a  and  a69459a );
 a1244a <=( a69446a  and  a69433a );
 a1245a <=( a69420a  and  a69407a );
 a1246a <=( a69394a  and  a69381a );
 a1247a <=( a69368a  and  a69355a );
 a1248a <=( a69342a  and  a69329a );
 a1249a <=( a69316a  and  a69303a );
 a1250a <=( a69290a  and  a69277a );
 a1251a <=( a69264a  and  a69251a );
 a1252a <=( a69238a  and  a69225a );
 a1253a <=( a69212a  and  a69199a );
 a1254a <=( a69186a  and  a69173a );
 a1255a <=( a69160a  and  a69147a );
 a1256a <=( a69134a  and  a69121a );
 a1257a <=( a69108a  and  a69095a );
 a1258a <=( a69082a  and  a69069a );
 a1259a <=( a69056a  and  a69043a );
 a1260a <=( a69030a  and  a69017a );
 a1261a <=( a69004a  and  a68991a );
 a1262a <=( a68978a  and  a68965a );
 a1263a <=( a68952a  and  a68939a );
 a1264a <=( a68926a  and  a68913a );
 a1265a <=( a68900a  and  a68887a );
 a1266a <=( a68874a  and  a68861a );
 a1267a <=( a68848a  and  a68835a );
 a1268a <=( a68822a  and  a68809a );
 a1269a <=( a68796a  and  a68783a );
 a1270a <=( a68770a  and  a68757a );
 a1271a <=( a68744a  and  a68731a );
 a1272a <=( a68718a  and  a68705a );
 a1273a <=( a68692a  and  a68679a );
 a1274a <=( a68666a  and  a68653a );
 a1275a <=( a68640a  and  a68627a );
 a1276a <=( a68614a  and  a68601a );
 a1277a <=( a68588a  and  a68575a );
 a1278a <=( a68562a  and  a68549a );
 a1279a <=( a68536a  and  a68523a );
 a1280a <=( a68510a  and  a68497a );
 a1281a <=( a68484a  and  a68471a );
 a1282a <=( a68458a  and  a68445a );
 a1283a <=( a68432a  and  a68419a );
 a1284a <=( a68406a  and  a68393a );
 a1285a <=( a68380a  and  a68367a );
 a1286a <=( a68354a  and  a68341a );
 a1287a <=( a68328a  and  a68315a );
 a1288a <=( a68302a  and  a68289a );
 a1289a <=( a68276a  and  a68263a );
 a1290a <=( a68250a  and  a68237a );
 a1291a <=( a68224a  and  a68211a );
 a1292a <=( a68198a  and  a68185a );
 a1293a <=( a68172a  and  a68159a );
 a1294a <=( a68146a  and  a68133a );
 a1295a <=( a68120a  and  a68107a );
 a1296a <=( a68094a  and  a68081a );
 a1297a <=( a68068a  and  a68055a );
 a1298a <=( a68042a  and  a68029a );
 a1299a <=( a68016a  and  a68003a );
 a1300a <=( a67990a  and  a67977a );
 a1301a <=( a67964a  and  a67951a );
 a1302a <=( a67938a  and  a67925a );
 a1303a <=( a67912a  and  a67899a );
 a1304a <=( a67886a  and  a67873a );
 a1305a <=( a67860a  and  a67847a );
 a1306a <=( a67834a  and  a67821a );
 a1307a <=( a67808a  and  a67795a );
 a1308a <=( a67782a  and  a67769a );
 a1309a <=( a67756a  and  a67743a );
 a1310a <=( a67730a  and  a67717a );
 a1311a <=( a67704a  and  a67691a );
 a1312a <=( a67678a  and  a67665a );
 a1313a <=( a67652a  and  a67639a );
 a1314a <=( a67626a  and  a67613a );
 a1315a <=( a67600a  and  a67587a );
 a1316a <=( a67574a  and  a67561a );
 a1317a <=( a67548a  and  a67535a );
 a1318a <=( a67522a  and  a67509a );
 a1319a <=( a67496a  and  a67483a );
 a1320a <=( a67470a  and  a67457a );
 a1321a <=( a67444a  and  a67431a );
 a1322a <=( a67418a  and  a67405a );
 a1323a <=( a67392a  and  a67379a );
 a1324a <=( a67366a  and  a67353a );
 a1325a <=( a67340a  and  a67327a );
 a1326a <=( a67314a  and  a67301a );
 a1327a <=( a67288a  and  a67275a );
 a1328a <=( a67262a  and  a67249a );
 a1329a <=( a67236a  and  a67223a );
 a1330a <=( a67210a  and  a67197a );
 a1331a <=( a67184a  and  a67171a );
 a1332a <=( a67158a  and  a67145a );
 a1333a <=( a67132a  and  a67119a );
 a1334a <=( a67106a  and  a67093a );
 a1335a <=( a67080a  and  a67067a );
 a1336a <=( a67054a  and  a67041a );
 a1337a <=( a67028a  and  a67015a );
 a1338a <=( a67002a  and  a66989a );
 a1339a <=( a66976a  and  a66963a );
 a1340a <=( a66950a  and  a66937a );
 a1341a <=( a66924a  and  a66911a );
 a1342a <=( a66898a  and  a66885a );
 a1343a <=( a66872a  and  a66859a );
 a1344a <=( a66846a  and  a66833a );
 a1345a <=( a66820a  and  a66807a );
 a1346a <=( a66794a  and  a66781a );
 a1347a <=( a66768a  and  a66755a );
 a1348a <=( a66742a  and  a66729a );
 a1349a <=( a66716a  and  a66703a );
 a1350a <=( a66690a  and  a66677a );
 a1351a <=( a66664a  and  a66651a );
 a1352a <=( a66638a  and  a66625a );
 a1353a <=( a66612a  and  a66599a );
 a1354a <=( a66586a  and  a66573a );
 a1355a <=( a66560a  and  a66547a );
 a1356a <=( a66534a  and  a66521a );
 a1357a <=( a66508a  and  a66495a );
 a1358a <=( a66482a  and  a66469a );
 a1359a <=( a66456a  and  a66443a );
 a1360a <=( a66430a  and  a66417a );
 a1361a <=( a66404a  and  a66391a );
 a1362a <=( a66378a  and  a66365a );
 a1363a <=( a66352a  and  a66339a );
 a1364a <=( a66326a  and  a66313a );
 a1365a <=( a66300a  and  a66287a );
 a1366a <=( a66274a  and  a66261a );
 a1367a <=( a66248a  and  a66235a );
 a1368a <=( a66222a  and  a66209a );
 a1369a <=( a66196a  and  a66183a );
 a1370a <=( a66170a  and  a66157a );
 a1371a <=( a66144a  and  a66131a );
 a1372a <=( a66118a  and  a66105a );
 a1373a <=( a66092a  and  a66079a );
 a1374a <=( a66066a  and  a66053a );
 a1375a <=( a66040a  and  a66027a );
 a1376a <=( a66014a  and  a66001a );
 a1377a <=( a65988a  and  a65975a );
 a1378a <=( a65962a  and  a65949a );
 a1379a <=( a65936a  and  a65923a );
 a1380a <=( a65910a  and  a65897a );
 a1381a <=( a65884a  and  a65871a );
 a1382a <=( a65858a  and  a65845a );
 a1383a <=( a65832a  and  a65819a );
 a1384a <=( a65806a  and  a65793a );
 a1385a <=( a65780a  and  a65767a );
 a1386a <=( a65754a  and  a65741a );
 a1387a <=( a65728a  and  a65715a );
 a1388a <=( a65702a  and  a65689a );
 a1389a <=( a65676a  and  a65663a );
 a1390a <=( a65650a  and  a65637a );
 a1391a <=( a65624a  and  a65611a );
 a1392a <=( a65598a  and  a65585a );
 a1393a <=( a65572a  and  a65559a );
 a1394a <=( a65546a  and  a65533a );
 a1395a <=( a65520a  and  a65507a );
 a1396a <=( a65494a  and  a65481a );
 a1397a <=( a65468a  and  a65455a );
 a1398a <=( a65442a  and  a65429a );
 a1399a <=( a65416a  and  a65403a );
 a1400a <=( a65390a  and  a65377a );
 a1401a <=( a65364a  and  a65351a );
 a1402a <=( a65338a  and  a65325a );
 a1403a <=( a65312a  and  a65299a );
 a1404a <=( a65286a  and  a65273a );
 a1405a <=( a65260a  and  a65247a );
 a1406a <=( a65234a  and  a65221a );
 a1407a <=( a65208a  and  a65195a );
 a1408a <=( a65182a  and  a65169a );
 a1409a <=( a65156a  and  a65143a );
 a1410a <=( a65130a  and  a65117a );
 a1411a <=( a65104a  and  a65091a );
 a1412a <=( a65078a  and  a65065a );
 a1413a <=( a65052a  and  a65039a );
 a1414a <=( a65026a  and  a65013a );
 a1415a <=( a65000a  and  a64987a );
 a1416a <=( a64974a  and  a64961a );
 a1417a <=( a64948a  and  a64935a );
 a1418a <=( a64922a  and  a64909a );
 a1419a <=( a64896a  and  a64883a );
 a1420a <=( a64870a  and  a64857a );
 a1421a <=( a64844a  and  a64831a );
 a1422a <=( a64818a  and  a64805a );
 a1423a <=( a64792a  and  a64779a );
 a1424a <=( a64766a  and  a64753a );
 a1425a <=( a64740a  and  a64727a );
 a1426a <=( a64714a  and  a64701a );
 a1427a <=( a64688a  and  a64675a );
 a1428a <=( a64662a  and  a64649a );
 a1429a <=( a64636a  and  a64623a );
 a1430a <=( a64610a  and  a64597a );
 a1431a <=( a64584a  and  a64571a );
 a1432a <=( a64558a  and  a64545a );
 a1433a <=( a64532a  and  a64519a );
 a1434a <=( a64506a  and  a64493a );
 a1435a <=( a64480a  and  a64467a );
 a1436a <=( a64454a  and  a64441a );
 a1437a <=( a64428a  and  a64415a );
 a1438a <=( a64402a  and  a64389a );
 a1439a <=( a64376a  and  a64363a );
 a1440a <=( a64350a  and  a64337a );
 a1441a <=( a64324a  and  a64311a );
 a1442a <=( a64298a  and  a64285a );
 a1443a <=( a64272a  and  a64259a );
 a1444a <=( a64246a  and  a64233a );
 a1445a <=( a64220a  and  a64207a );
 a1446a <=( a64194a  and  a64181a );
 a1447a <=( a64168a  and  a64155a );
 a1448a <=( a64142a  and  a64129a );
 a1449a <=( a64116a  and  a64103a );
 a1450a <=( a64090a  and  a64077a );
 a1451a <=( a64064a  and  a64051a );
 a1452a <=( a64038a  and  a64025a );
 a1453a <=( a64012a  and  a63999a );
 a1454a <=( a63986a  and  a63973a );
 a1455a <=( a63960a  and  a63947a );
 a1456a <=( a63934a  and  a63921a );
 a1457a <=( a63908a  and  a63895a );
 a1458a <=( a63882a  and  a63869a );
 a1459a <=( a63856a  and  a63843a );
 a1460a <=( a63830a  and  a63817a );
 a1461a <=( a63804a  and  a63791a );
 a1462a <=( a63778a  and  a63765a );
 a1463a <=( a63752a  and  a63739a );
 a1464a <=( a63726a  and  a63713a );
 a1465a <=( a63700a  and  a63687a );
 a1466a <=( a63674a  and  a63661a );
 a1467a <=( a63648a  and  a63635a );
 a1468a <=( a63622a  and  a63609a );
 a1469a <=( a63596a  and  a63583a );
 a1470a <=( a63570a  and  a63557a );
 a1471a <=( a63544a  and  a63531a );
 a1472a <=( a63518a  and  a63505a );
 a1473a <=( a63492a  and  a63479a );
 a1474a <=( a63466a  and  a63453a );
 a1475a <=( a63440a  and  a63427a );
 a1476a <=( a63414a  and  a63401a );
 a1477a <=( a63388a  and  a63375a );
 a1478a <=( a63362a  and  a63349a );
 a1479a <=( a63336a  and  a63323a );
 a1480a <=( a63310a  and  a63297a );
 a1481a <=( a63284a  and  a63271a );
 a1482a <=( a63258a  and  a63245a );
 a1483a <=( a63232a  and  a63219a );
 a1484a <=( a63206a  and  a63193a );
 a1485a <=( a63180a  and  a63167a );
 a1486a <=( a63154a  and  a63141a );
 a1487a <=( a63128a  and  a63115a );
 a1488a <=( a63102a  and  a63089a );
 a1489a <=( a63076a  and  a63063a );
 a1490a <=( a63050a  and  a63037a );
 a1491a <=( a63024a  and  a63011a );
 a1492a <=( a62998a  and  a62985a );
 a1493a <=( a62972a  and  a62959a );
 a1494a <=( a62946a  and  a62933a );
 a1495a <=( a62920a  and  a62907a );
 a1496a <=( a62894a  and  a62881a );
 a1497a <=( a62868a  and  a62855a );
 a1498a <=( a62842a  and  a62829a );
 a1499a <=( a62816a  and  a62803a );
 a1500a <=( a62790a  and  a62777a );
 a1501a <=( a62764a  and  a62751a );
 a1502a <=( a62738a  and  a62725a );
 a1503a <=( a62712a  and  a62699a );
 a1504a <=( a62686a  and  a62673a );
 a1505a <=( a62660a  and  a62647a );
 a1506a <=( a62634a  and  a62621a );
 a1507a <=( a62608a  and  a62595a );
 a1508a <=( a62582a  and  a62569a );
 a1509a <=( a62556a  and  a62543a );
 a1510a <=( a62530a  and  a62517a );
 a1511a <=( a62504a  and  a62491a );
 a1512a <=( a62478a  and  a62465a );
 a1513a <=( a62452a  and  a62439a );
 a1514a <=( a62426a  and  a62413a );
 a1515a <=( a62400a  and  a62387a );
 a1516a <=( a62374a  and  a62361a );
 a1517a <=( a62348a  and  a62335a );
 a1518a <=( a62322a  and  a62309a );
 a1519a <=( a62296a  and  a62283a );
 a1520a <=( a62270a  and  a62257a );
 a1521a <=( a62244a  and  a62231a );
 a1522a <=( a62218a  and  a62205a );
 a1523a <=( a62192a  and  a62179a );
 a1524a <=( a62166a  and  a62153a );
 a1525a <=( a62140a  and  a62127a );
 a1526a <=( a62114a  and  a62101a );
 a1527a <=( a62088a  and  a62075a );
 a1528a <=( a62062a  and  a62049a );
 a1529a <=( a62036a  and  a62023a );
 a1530a <=( a62010a  and  a61997a );
 a1531a <=( a61984a  and  a61971a );
 a1532a <=( a61958a  and  a61945a );
 a1533a <=( a61932a  and  a61919a );
 a1534a <=( a61906a  and  a61893a );
 a1535a <=( a61880a  and  a61867a );
 a1536a <=( a61854a  and  a61841a );
 a1537a <=( a61828a  and  a61815a );
 a1538a <=( a61802a  and  a61789a );
 a1539a <=( a61776a  and  a61763a );
 a1540a <=( a61750a  and  a61737a );
 a1541a <=( a61724a  and  a61711a );
 a1542a <=( a61698a  and  a61685a );
 a1543a <=( a61672a  and  a61659a );
 a1544a <=( a61646a  and  a61633a );
 a1545a <=( a61620a  and  a61607a );
 a1546a <=( a61594a  and  a61581a );
 a1547a <=( a61568a  and  a61555a );
 a1548a <=( a61542a  and  a61529a );
 a1549a <=( a61516a  and  a61503a );
 a1550a <=( a61490a  and  a61477a );
 a1551a <=( a61464a  and  a61451a );
 a1552a <=( a61438a  and  a61425a );
 a1553a <=( a61412a  and  a61399a );
 a1554a <=( a61386a  and  a61373a );
 a1555a <=( a61360a  and  a61347a );
 a1556a <=( a61334a  and  a61321a );
 a1557a <=( a61308a  and  a61295a );
 a1558a <=( a61282a  and  a61269a );
 a1559a <=( a61256a  and  a61243a );
 a1560a <=( a61230a  and  a61217a );
 a1561a <=( a61204a  and  a61191a );
 a1562a <=( a61178a  and  a61165a );
 a1563a <=( a61152a  and  a61139a );
 a1564a <=( a61126a  and  a61113a );
 a1565a <=( a61100a  and  a61087a );
 a1566a <=( a61074a  and  a61061a );
 a1567a <=( a61048a  and  a61035a );
 a1568a <=( a61022a  and  a61009a );
 a1569a <=( a60996a  and  a60983a );
 a1570a <=( a60970a  and  a60957a );
 a1571a <=( a60944a  and  a60931a );
 a1572a <=( a60918a  and  a60905a );
 a1573a <=( a60892a  and  a60879a );
 a1574a <=( a60866a  and  a60853a );
 a1575a <=( a60840a  and  a60827a );
 a1576a <=( a60814a  and  a60801a );
 a1577a <=( a60788a  and  a60775a );
 a1578a <=( a60762a  and  a60749a );
 a1579a <=( a60736a  and  a60723a );
 a1580a <=( a60710a  and  a60697a );
 a1581a <=( a60684a  and  a60671a );
 a1582a <=( a60658a  and  a60645a );
 a1583a <=( a60632a  and  a60619a );
 a1584a <=( a60606a  and  a60593a );
 a1585a <=( a60580a  and  a60567a );
 a1586a <=( a60554a  and  a60541a );
 a1587a <=( a60528a  and  a60515a );
 a1588a <=( a60502a  and  a60489a );
 a1589a <=( a60476a  and  a60463a );
 a1590a <=( a60450a  and  a60437a );
 a1591a <=( a60424a  and  a60411a );
 a1592a <=( a60398a  and  a60385a );
 a1593a <=( a60372a  and  a60359a );
 a1594a <=( a60346a  and  a60333a );
 a1595a <=( a60320a  and  a60307a );
 a1596a <=( a60294a  and  a60281a );
 a1597a <=( a60268a  and  a60255a );
 a1598a <=( a60242a  and  a60229a );
 a1599a <=( a60216a  and  a60203a );
 a1600a <=( a60190a  and  a60177a );
 a1601a <=( a60164a  and  a60151a );
 a1602a <=( a60138a  and  a60125a );
 a1603a <=( a60112a  and  a60099a );
 a1604a <=( a60088a  and  a60075a );
 a1605a <=( a60064a  and  a60051a );
 a1606a <=( a60040a  and  a60027a );
 a1607a <=( a60016a  and  a60003a );
 a1608a <=( a59992a  and  a59979a );
 a1609a <=( a59968a  and  a59955a );
 a1610a <=( a59944a  and  a59931a );
 a1611a <=( a59920a  and  a59907a );
 a1612a <=( a59896a  and  a59883a );
 a1613a <=( a59872a  and  a59859a );
 a1614a <=( a59848a  and  a59835a );
 a1615a <=( a59824a  and  a59811a );
 a1616a <=( a59800a  and  a59787a );
 a1617a <=( a59776a  and  a59763a );
 a1618a <=( a59752a  and  a59739a );
 a1619a <=( a59728a  and  a59715a );
 a1620a <=( a59704a  and  a59691a );
 a1621a <=( a59680a  and  a59667a );
 a1622a <=( a59656a  and  a59643a );
 a1623a <=( a59632a  and  a59619a );
 a1624a <=( a59608a  and  a59595a );
 a1625a <=( a59584a  and  a59571a );
 a1626a <=( a59560a  and  a59547a );
 a1627a <=( a59536a  and  a59523a );
 a1628a <=( a59512a  and  a59499a );
 a1629a <=( a59488a  and  a59475a );
 a1630a <=( a59464a  and  a59451a );
 a1631a <=( a59440a  and  a59427a );
 a1632a <=( a59416a  and  a59403a );
 a1633a <=( a59392a  and  a59379a );
 a1634a <=( a59368a  and  a59355a );
 a1635a <=( a59344a  and  a59331a );
 a1636a <=( a59320a  and  a59307a );
 a1637a <=( a59296a  and  a59283a );
 a1638a <=( a59272a  and  a59259a );
 a1639a <=( a59248a  and  a59235a );
 a1640a <=( a59224a  and  a59211a );
 a1641a <=( a59200a  and  a59187a );
 a1642a <=( a59176a  and  a59163a );
 a1643a <=( a59152a  and  a59139a );
 a1644a <=( a59128a  and  a59115a );
 a1645a <=( a59104a  and  a59091a );
 a1646a <=( a59080a  and  a59067a );
 a1647a <=( a59056a  and  a59043a );
 a1648a <=( a59032a  and  a59019a );
 a1649a <=( a59008a  and  a58995a );
 a1650a <=( a58984a  and  a58971a );
 a1651a <=( a58960a  and  a58947a );
 a1652a <=( a58936a  and  a58923a );
 a1653a <=( a58912a  and  a58899a );
 a1654a <=( a58888a  and  a58875a );
 a1655a <=( a58864a  and  a58851a );
 a1656a <=( a58840a  and  a58827a );
 a1657a <=( a58816a  and  a58803a );
 a1658a <=( a58792a  and  a58779a );
 a1659a <=( a58768a  and  a58755a );
 a1660a <=( a58744a  and  a58731a );
 a1661a <=( a58720a  and  a58707a );
 a1662a <=( a58696a  and  a58683a );
 a1663a <=( a58672a  and  a58659a );
 a1664a <=( a58648a  and  a58635a );
 a1665a <=( a58624a  and  a58611a );
 a1666a <=( a58600a  and  a58587a );
 a1667a <=( a58576a  and  a58563a );
 a1668a <=( a58552a  and  a58539a );
 a1669a <=( a58528a  and  a58515a );
 a1670a <=( a58504a  and  a58491a );
 a1671a <=( a58480a  and  a58467a );
 a1672a <=( a58456a  and  a58443a );
 a1673a <=( a58432a  and  a58419a );
 a1674a <=( a58408a  and  a58395a );
 a1675a <=( a58384a  and  a58371a );
 a1676a <=( a58360a  and  a58347a );
 a1677a <=( a58336a  and  a58323a );
 a1678a <=( a58312a  and  a58299a );
 a1679a <=( a58288a  and  a58275a );
 a1680a <=( a58264a  and  a58251a );
 a1681a <=( a58240a  and  a58227a );
 a1682a <=( a58216a  and  a58203a );
 a1683a <=( a58192a  and  a58179a );
 a1684a <=( a58168a  and  a58155a );
 a1685a <=( a58144a  and  a58131a );
 a1686a <=( a58120a  and  a58107a );
 a1687a <=( a58096a  and  a58083a );
 a1688a <=( a58072a  and  a58059a );
 a1689a <=( a58048a  and  a58035a );
 a1690a <=( a58024a  and  a58011a );
 a1691a <=( a58000a  and  a57987a );
 a1692a <=( a57976a  and  a57963a );
 a1693a <=( a57952a  and  a57939a );
 a1694a <=( a57928a  and  a57915a );
 a1695a <=( a57904a  and  a57891a );
 a1696a <=( a57880a  and  a57867a );
 a1697a <=( a57856a  and  a57843a );
 a1698a <=( a57832a  and  a57819a );
 a1699a <=( a57808a  and  a57795a );
 a1700a <=( a57784a  and  a57771a );
 a1701a <=( a57760a  and  a57747a );
 a1702a <=( a57736a  and  a57723a );
 a1703a <=( a57712a  and  a57699a );
 a1704a <=( a57688a  and  a57675a );
 a1705a <=( a57664a  and  a57651a );
 a1706a <=( a57640a  and  a57627a );
 a1707a <=( a57616a  and  a57603a );
 a1708a <=( a57592a  and  a57579a );
 a1709a <=( a57568a  and  a57555a );
 a1710a <=( a57544a  and  a57531a );
 a1711a <=( a57520a  and  a57507a );
 a1712a <=( a57496a  and  a57483a );
 a1713a <=( a57472a  and  a57459a );
 a1714a <=( a57448a  and  a57435a );
 a1715a <=( a57424a  and  a57411a );
 a1716a <=( a57400a  and  a57387a );
 a1717a <=( a57376a  and  a57363a );
 a1718a <=( a57352a  and  a57339a );
 a1719a <=( a57328a  and  a57315a );
 a1720a <=( a57304a  and  a57291a );
 a1721a <=( a57280a  and  a57267a );
 a1722a <=( a57256a  and  a57243a );
 a1723a <=( a57232a  and  a57219a );
 a1724a <=( a57208a  and  a57195a );
 a1725a <=( a57184a  and  a57171a );
 a1726a <=( a57160a  and  a57147a );
 a1727a <=( a57136a  and  a57123a );
 a1728a <=( a57112a  and  a57099a );
 a1729a <=( a57088a  and  a57075a );
 a1730a <=( a57064a  and  a57051a );
 a1731a <=( a57040a  and  a57027a );
 a1732a <=( a57016a  and  a57003a );
 a1733a <=( a56992a  and  a56979a );
 a1734a <=( a56968a  and  a56955a );
 a1735a <=( a56944a  and  a56931a );
 a1736a <=( a56920a  and  a56907a );
 a1737a <=( a56896a  and  a56883a );
 a1738a <=( a56872a  and  a56859a );
 a1739a <=( a56848a  and  a56835a );
 a1740a <=( a56824a  and  a56811a );
 a1741a <=( a56800a  and  a56787a );
 a1742a <=( a56776a  and  a56763a );
 a1743a <=( a56752a  and  a56739a );
 a1744a <=( a56728a  and  a56715a );
 a1745a <=( a56704a  and  a56691a );
 a1746a <=( a56680a  and  a56667a );
 a1747a <=( a56656a  and  a56643a );
 a1748a <=( a56632a  and  a56619a );
 a1749a <=( a56608a  and  a56595a );
 a1750a <=( a56584a  and  a56571a );
 a1751a <=( a56560a  and  a56547a );
 a1752a <=( a56536a  and  a56523a );
 a1753a <=( a56512a  and  a56499a );
 a1754a <=( a56488a  and  a56475a );
 a1755a <=( a56464a  and  a56451a );
 a1756a <=( a56440a  and  a56427a );
 a1757a <=( a56416a  and  a56403a );
 a1758a <=( a56392a  and  a56379a );
 a1759a <=( a56368a  and  a56355a );
 a1760a <=( a56344a  and  a56331a );
 a1761a <=( a56320a  and  a56307a );
 a1762a <=( a56296a  and  a56283a );
 a1763a <=( a56272a  and  a56259a );
 a1764a <=( a56248a  and  a56235a );
 a1765a <=( a56224a  and  a56211a );
 a1766a <=( a56200a  and  a56187a );
 a1767a <=( a56176a  and  a56163a );
 a1768a <=( a56152a  and  a56139a );
 a1769a <=( a56128a  and  a56115a );
 a1770a <=( a56104a  and  a56091a );
 a1771a <=( a56080a  and  a56067a );
 a1772a <=( a56056a  and  a56043a );
 a1773a <=( a56032a  and  a56019a );
 a1774a <=( a56008a  and  a55995a );
 a1775a <=( a55984a  and  a55971a );
 a1776a <=( a55960a  and  a55947a );
 a1777a <=( a55936a  and  a55923a );
 a1778a <=( a55912a  and  a55899a );
 a1779a <=( a55888a  and  a55875a );
 a1780a <=( a55864a  and  a55851a );
 a1781a <=( a55840a  and  a55827a );
 a1782a <=( a55816a  and  a55803a );
 a1783a <=( a55792a  and  a55779a );
 a1784a <=( a55768a  and  a55755a );
 a1785a <=( a55744a  and  a55731a );
 a1786a <=( a55720a  and  a55707a );
 a1787a <=( a55696a  and  a55683a );
 a1788a <=( a55672a  and  a55659a );
 a1789a <=( a55648a  and  a55635a );
 a1790a <=( a55624a  and  a55611a );
 a1791a <=( a55600a  and  a55587a );
 a1792a <=( a55576a  and  a55563a );
 a1793a <=( a55552a  and  a55539a );
 a1794a <=( a55528a  and  a55515a );
 a1795a <=( a55504a  and  a55491a );
 a1796a <=( a55480a  and  a55467a );
 a1797a <=( a55456a  and  a55443a );
 a1798a <=( a55432a  and  a55419a );
 a1799a <=( a55408a  and  a55395a );
 a1800a <=( a55384a  and  a55371a );
 a1801a <=( a55360a  and  a55347a );
 a1802a <=( a55336a  and  a55323a );
 a1803a <=( a55312a  and  a55299a );
 a1804a <=( a55288a  and  a55275a );
 a1805a <=( a55264a  and  a55251a );
 a1806a <=( a55240a  and  a55227a );
 a1807a <=( a55216a  and  a55203a );
 a1808a <=( a55192a  and  a55179a );
 a1809a <=( a55168a  and  a55155a );
 a1810a <=( a55144a  and  a55131a );
 a1811a <=( a55120a  and  a55107a );
 a1812a <=( a55096a  and  a55083a );
 a1813a <=( a55072a  and  a55059a );
 a1814a <=( a55048a  and  a55035a );
 a1815a <=( a55024a  and  a55011a );
 a1816a <=( a55000a  and  a54987a );
 a1817a <=( a54976a  and  a54963a );
 a1818a <=( a54952a  and  a54939a );
 a1819a <=( a54928a  and  a54915a );
 a1820a <=( a54904a  and  a54891a );
 a1821a <=( a54880a  and  a54867a );
 a1822a <=( a54856a  and  a54843a );
 a1823a <=( a54832a  and  a54819a );
 a1824a <=( a54808a  and  a54795a );
 a1825a <=( a54784a  and  a54771a );
 a1826a <=( a54760a  and  a54747a );
 a1827a <=( a54736a  and  a54723a );
 a1828a <=( a54712a  and  a54699a );
 a1829a <=( a54688a  and  a54675a );
 a1830a <=( a54664a  and  a54651a );
 a1831a <=( a54640a  and  a54627a );
 a1832a <=( a54616a  and  a54603a );
 a1833a <=( a54592a  and  a54579a );
 a1834a <=( a54568a  and  a54555a );
 a1835a <=( a54544a  and  a54531a );
 a1836a <=( a54520a  and  a54507a );
 a1837a <=( a54496a  and  a54483a );
 a1838a <=( a54472a  and  a54459a );
 a1839a <=( a54448a  and  a54435a );
 a1840a <=( a54424a  and  a54411a );
 a1841a <=( a54400a  and  a54387a );
 a1842a <=( a54376a  and  a54363a );
 a1843a <=( a54352a  and  a54339a );
 a1844a <=( a54328a  and  a54315a );
 a1845a <=( a54304a  and  a54291a );
 a1846a <=( a54280a  and  a54267a );
 a1847a <=( a54256a  and  a54243a );
 a1848a <=( a54232a  and  a54219a );
 a1849a <=( a54208a  and  a54195a );
 a1850a <=( a54184a  and  a54171a );
 a1851a <=( a54160a  and  a54147a );
 a1852a <=( a54136a  and  a54123a );
 a1853a <=( a54112a  and  a54099a );
 a1854a <=( a54088a  and  a54075a );
 a1855a <=( a54064a  and  a54051a );
 a1856a <=( a54040a  and  a54027a );
 a1857a <=( a54016a  and  a54003a );
 a1858a <=( a53992a  and  a53979a );
 a1859a <=( a53968a  and  a53955a );
 a1860a <=( a53944a  and  a53931a );
 a1861a <=( a53920a  and  a53907a );
 a1862a <=( a53896a  and  a53883a );
 a1863a <=( a53872a  and  a53859a );
 a1864a <=( a53848a  and  a53835a );
 a1865a <=( a53824a  and  a53811a );
 a1866a <=( a53800a  and  a53787a );
 a1867a <=( a53776a  and  a53763a );
 a1868a <=( a53752a  and  a53739a );
 a1869a <=( a53728a  and  a53715a );
 a1870a <=( a53704a  and  a53691a );
 a1871a <=( a53680a  and  a53667a );
 a1872a <=( a53656a  and  a53643a );
 a1873a <=( a53632a  and  a53619a );
 a1874a <=( a53608a  and  a53595a );
 a1875a <=( a53584a  and  a53571a );
 a1876a <=( a53560a  and  a53547a );
 a1877a <=( a53536a  and  a53523a );
 a1878a <=( a53512a  and  a53499a );
 a1879a <=( a53488a  and  a53475a );
 a1880a <=( a53464a  and  a53451a );
 a1881a <=( a53440a  and  a53427a );
 a1882a <=( a53416a  and  a53403a );
 a1883a <=( a53392a  and  a53379a );
 a1884a <=( a53368a  and  a53355a );
 a1885a <=( a53344a  and  a53331a );
 a1886a <=( a53320a  and  a53307a );
 a1887a <=( a53296a  and  a53283a );
 a1888a <=( a53272a  and  a53259a );
 a1889a <=( a53248a  and  a53235a );
 a1890a <=( a53224a  and  a53211a );
 a1891a <=( a53200a  and  a53187a );
 a1892a <=( a53176a  and  a53163a );
 a1893a <=( a53152a  and  a53139a );
 a1894a <=( a53128a  and  a53115a );
 a1895a <=( a53104a  and  a53091a );
 a1896a <=( a53080a  and  a53067a );
 a1897a <=( a53056a  and  a53043a );
 a1898a <=( a53032a  and  a53019a );
 a1899a <=( a53008a  and  a52995a );
 a1900a <=( a52984a  and  a52971a );
 a1901a <=( a52960a  and  a52947a );
 a1902a <=( a52936a  and  a52923a );
 a1903a <=( a52912a  and  a52899a );
 a1904a <=( a52888a  and  a52875a );
 a1905a <=( a52864a  and  a52851a );
 a1906a <=( a52840a  and  a52827a );
 a1907a <=( a52816a  and  a52803a );
 a1908a <=( a52792a  and  a52779a );
 a1909a <=( a52768a  and  a52755a );
 a1910a <=( a52744a  and  a52731a );
 a1911a <=( a52720a  and  a52707a );
 a1912a <=( a52696a  and  a52683a );
 a1913a <=( a52672a  and  a52659a );
 a1914a <=( a52648a  and  a52635a );
 a1915a <=( a52624a  and  a52611a );
 a1916a <=( a52600a  and  a52587a );
 a1917a <=( a52576a  and  a52563a );
 a1918a <=( a52552a  and  a52539a );
 a1919a <=( a52528a  and  a52515a );
 a1920a <=( a52504a  and  a52491a );
 a1921a <=( a52480a  and  a52467a );
 a1922a <=( a52456a  and  a52443a );
 a1923a <=( a52432a  and  a52419a );
 a1924a <=( a52408a  and  a52395a );
 a1925a <=( a52384a  and  a52371a );
 a1926a <=( a52360a  and  a52347a );
 a1927a <=( a52336a  and  a52323a );
 a1928a <=( a52312a  and  a52299a );
 a1929a <=( a52288a  and  a52275a );
 a1930a <=( a52264a  and  a52251a );
 a1931a <=( a52240a  and  a52227a );
 a1932a <=( a52216a  and  a52203a );
 a1933a <=( a52192a  and  a52179a );
 a1934a <=( a52168a  and  a52155a );
 a1935a <=( a52144a  and  a52131a );
 a1936a <=( a52120a  and  a52107a );
 a1937a <=( a52096a  and  a52083a );
 a1938a <=( a52072a  and  a52059a );
 a1939a <=( a52048a  and  a52035a );
 a1940a <=( a52024a  and  a52011a );
 a1941a <=( a52000a  and  a51987a );
 a1942a <=( a51976a  and  a51963a );
 a1943a <=( a51952a  and  a51939a );
 a1944a <=( a51928a  and  a51915a );
 a1945a <=( a51904a  and  a51891a );
 a1946a <=( a51880a  and  a51867a );
 a1947a <=( a51856a  and  a51843a );
 a1948a <=( a51832a  and  a51819a );
 a1949a <=( a51808a  and  a51795a );
 a1950a <=( a51784a  and  a51771a );
 a1951a <=( a51760a  and  a51747a );
 a1952a <=( a51736a  and  a51723a );
 a1953a <=( a51712a  and  a51699a );
 a1954a <=( a51688a  and  a51675a );
 a1955a <=( a51664a  and  a51651a );
 a1956a <=( a51640a  and  a51627a );
 a1957a <=( a51616a  and  a51603a );
 a1958a <=( a51592a  and  a51579a );
 a1959a <=( a51568a  and  a51555a );
 a1960a <=( a51544a  and  a51531a );
 a1961a <=( a51520a  and  a51507a );
 a1962a <=( a51496a  and  a51483a );
 a1963a <=( a51472a  and  a51459a );
 a1964a <=( a51448a  and  a51435a );
 a1965a <=( a51424a  and  a51411a );
 a1966a <=( a51400a  and  a51387a );
 a1967a <=( a51376a  and  a51363a );
 a1968a <=( a51352a  and  a51339a );
 a1969a <=( a51328a  and  a51315a );
 a1970a <=( a51304a  and  a51291a );
 a1971a <=( a51280a  and  a51267a );
 a1972a <=( a51256a  and  a51243a );
 a1973a <=( a51232a  and  a51219a );
 a1974a <=( a51208a  and  a51195a );
 a1975a <=( a51184a  and  a51171a );
 a1976a <=( a51160a  and  a51147a );
 a1977a <=( a51136a  and  a51123a );
 a1978a <=( a51112a  and  a51099a );
 a1979a <=( a51088a  and  a51075a );
 a1980a <=( a51064a  and  a51051a );
 a1981a <=( a51040a  and  a51027a );
 a1982a <=( a51016a  and  a51003a );
 a1983a <=( a50992a  and  a50979a );
 a1984a <=( a50968a  and  a50955a );
 a1985a <=( a50944a  and  a50931a );
 a1986a <=( a50920a  and  a50907a );
 a1987a <=( a50896a  and  a50883a );
 a1988a <=( a50872a  and  a50859a );
 a1989a <=( a50848a  and  a50835a );
 a1990a <=( a50824a  and  a50811a );
 a1991a <=( a50800a  and  a50787a );
 a1992a <=( a50776a  and  a50763a );
 a1993a <=( a50752a  and  a50739a );
 a1994a <=( a50728a  and  a50715a );
 a1995a <=( a50704a  and  a50691a );
 a1996a <=( a50680a  and  a50667a );
 a1997a <=( a50656a  and  a50643a );
 a1998a <=( a50632a  and  a50619a );
 a1999a <=( a50608a  and  a50595a );
 a2000a <=( a50584a  and  a50571a );
 a2001a <=( a50560a  and  a50547a );
 a2002a <=( a50536a  and  a50523a );
 a2003a <=( a50512a  and  a50499a );
 a2004a <=( a50488a  and  a50475a );
 a2005a <=( a50464a  and  a50451a );
 a2006a <=( a50440a  and  a50427a );
 a2007a <=( a50416a  and  a50403a );
 a2008a <=( a50392a  and  a50379a );
 a2009a <=( a50368a  and  a50355a );
 a2010a <=( a50344a  and  a50331a );
 a2011a <=( a50320a  and  a50307a );
 a2012a <=( a50296a  and  a50283a );
 a2013a <=( a50272a  and  a50259a );
 a2014a <=( a50248a  and  a50235a );
 a2015a <=( a50224a  and  a50211a );
 a2016a <=( a50200a  and  a50187a );
 a2017a <=( a50176a  and  a50163a );
 a2018a <=( a50152a  and  a50139a );
 a2019a <=( a50128a  and  a50115a );
 a2020a <=( a50104a  and  a50091a );
 a2021a <=( a50080a  and  a50067a );
 a2022a <=( a50056a  and  a50043a );
 a2023a <=( a50032a  and  a50019a );
 a2024a <=( a50008a  and  a49995a );
 a2025a <=( a49984a  and  a49971a );
 a2026a <=( a49960a  and  a49947a );
 a2027a <=( a49936a  and  a49923a );
 a2028a <=( a49912a  and  a49899a );
 a2029a <=( a49888a  and  a49875a );
 a2030a <=( a49864a  and  a49851a );
 a2031a <=( a49840a  and  a49827a );
 a2032a <=( a49816a  and  a49803a );
 a2033a <=( a49792a  and  a49779a );
 a2034a <=( a49768a  and  a49755a );
 a2035a <=( a49744a  and  a49731a );
 a2036a <=( a49720a  and  a49707a );
 a2037a <=( a49696a  and  a49683a );
 a2038a <=( a49672a  and  a49659a );
 a2039a <=( a49648a  and  a49635a );
 a2040a <=( a49624a  and  a49611a );
 a2041a <=( a49600a  and  a49587a );
 a2042a <=( a49576a  and  a49563a );
 a2043a <=( a49552a  and  a49539a );
 a2044a <=( a49528a  and  a49515a );
 a2045a <=( a49504a  and  a49491a );
 a2046a <=( a49480a  and  a49467a );
 a2047a <=( a49456a  and  a49443a );
 a2048a <=( a49432a  and  a49419a );
 a2049a <=( a49408a  and  a49395a );
 a2050a <=( a49384a  and  a49371a );
 a2051a <=( a49360a  and  a49347a );
 a2052a <=( a49336a  and  a49323a );
 a2053a <=( a49312a  and  a49299a );
 a2054a <=( a49288a  and  a49275a );
 a2055a <=( a49264a  and  a49251a );
 a2056a <=( a49240a  and  a49227a );
 a2057a <=( a49216a  and  a49203a );
 a2058a <=( a49192a  and  a49179a );
 a2059a <=( a49168a  and  a49155a );
 a2060a <=( a49144a  and  a49131a );
 a2061a <=( a49120a  and  a49107a );
 a2062a <=( a49096a  and  a49083a );
 a2063a <=( a49072a  and  a49059a );
 a2064a <=( a49048a  and  a49035a );
 a2065a <=( a49024a  and  a49011a );
 a2066a <=( a49000a  and  a48987a );
 a2067a <=( a48976a  and  a48963a );
 a2068a <=( a48952a  and  a48939a );
 a2069a <=( a48928a  and  a48915a );
 a2070a <=( a48904a  and  a48891a );
 a2071a <=( a48880a  and  a48867a );
 a2072a <=( a48856a  and  a48843a );
 a2073a <=( a48832a  and  a48819a );
 a2074a <=( a48808a  and  a48795a );
 a2075a <=( a48784a  and  a48771a );
 a2076a <=( a48760a  and  a48747a );
 a2077a <=( a48736a  and  a48723a );
 a2078a <=( a48712a  and  a48699a );
 a2079a <=( a48688a  and  a48675a );
 a2080a <=( a48664a  and  a48651a );
 a2081a <=( a48640a  and  a48627a );
 a2082a <=( a48616a  and  a48603a );
 a2083a <=( a48592a  and  a48579a );
 a2084a <=( a48568a  and  a48555a );
 a2085a <=( a48544a  and  a48531a );
 a2086a <=( a48520a  and  a48507a );
 a2087a <=( a48496a  and  a48483a );
 a2088a <=( a48472a  and  a48459a );
 a2089a <=( a48448a  and  a48435a );
 a2090a <=( a48424a  and  a48411a );
 a2091a <=( a48400a  and  a48387a );
 a2092a <=( a48376a  and  a48363a );
 a2093a <=( a48352a  and  a48339a );
 a2094a <=( a48328a  and  a48315a );
 a2095a <=( a48304a  and  a48291a );
 a2096a <=( a48280a  and  a48267a );
 a2097a <=( a48256a  and  a48243a );
 a2098a <=( a48232a  and  a48219a );
 a2099a <=( a48208a  and  a48195a );
 a2100a <=( a48184a  and  a48171a );
 a2101a <=( a48160a  and  a48147a );
 a2102a <=( a48136a  and  a48123a );
 a2103a <=( a48112a  and  a48099a );
 a2104a <=( a48088a  and  a48075a );
 a2105a <=( a48064a  and  a48051a );
 a2106a <=( a48040a  and  a48027a );
 a2107a <=( a48016a  and  a48003a );
 a2108a <=( a47992a  and  a47979a );
 a2109a <=( a47968a  and  a47955a );
 a2110a <=( a47944a  and  a47931a );
 a2111a <=( a47920a  and  a47907a );
 a2112a <=( a47896a  and  a47883a );
 a2113a <=( a47872a  and  a47859a );
 a2114a <=( a47848a  and  a47835a );
 a2115a <=( a47824a  and  a47811a );
 a2116a <=( a47800a  and  a47787a );
 a2117a <=( a47776a  and  a47763a );
 a2118a <=( a47752a  and  a47739a );
 a2119a <=( a47728a  and  a47715a );
 a2120a <=( a47704a  and  a47691a );
 a2121a <=( a47680a  and  a47667a );
 a2122a <=( a47656a  and  a47643a );
 a2123a <=( a47632a  and  a47619a );
 a2124a <=( a47608a  and  a47595a );
 a2125a <=( a47584a  and  a47571a );
 a2126a <=( a47560a  and  a47547a );
 a2127a <=( a47536a  and  a47523a );
 a2128a <=( a47512a  and  a47499a );
 a2129a <=( a47488a  and  a47475a );
 a2130a <=( a47464a  and  a47451a );
 a2131a <=( a47440a  and  a47427a );
 a2132a <=( a47416a  and  a47403a );
 a2133a <=( a47392a  and  a47379a );
 a2134a <=( a47368a  and  a47355a );
 a2135a <=( a47344a  and  a47331a );
 a2136a <=( a47320a  and  a47307a );
 a2137a <=( a47296a  and  a47283a );
 a2138a <=( a47272a  and  a47259a );
 a2139a <=( a47248a  and  a47235a );
 a2140a <=( a47224a  and  a47211a );
 a2141a <=( a47200a  and  a47187a );
 a2142a <=( a47176a  and  a47163a );
 a2143a <=( a47152a  and  a47139a );
 a2144a <=( a47128a  and  a47115a );
 a2145a <=( a47104a  and  a47091a );
 a2146a <=( a47080a  and  a47067a );
 a2147a <=( a47056a  and  a47043a );
 a2148a <=( a47032a  and  a47019a );
 a2149a <=( a47008a  and  a46995a );
 a2150a <=( a46984a  and  a46971a );
 a2151a <=( a46960a  and  a46947a );
 a2152a <=( a46936a  and  a46923a );
 a2153a <=( a46912a  and  a46899a );
 a2154a <=( a46888a  and  a46875a );
 a2155a <=( a46864a  and  a46851a );
 a2156a <=( a46840a  and  a46827a );
 a2157a <=( a46816a  and  a46803a );
 a2158a <=( a46792a  and  a46779a );
 a2159a <=( a46768a  and  a46755a );
 a2160a <=( a46744a  and  a46731a );
 a2161a <=( a46720a  and  a46707a );
 a2162a <=( a46696a  and  a46683a );
 a2163a <=( a46672a  and  a46659a );
 a2164a <=( a46648a  and  a46635a );
 a2165a <=( a46624a  and  a46611a );
 a2166a <=( a46600a  and  a46587a );
 a2167a <=( a46576a  and  a46563a );
 a2168a <=( a46552a  and  a46539a );
 a2169a <=( a46528a  and  a46515a );
 a2170a <=( a46504a  and  a46491a );
 a2171a <=( a46480a  and  a46467a );
 a2172a <=( a46456a  and  a46443a );
 a2173a <=( a46432a  and  a46419a );
 a2174a <=( a46408a  and  a46395a );
 a2175a <=( a46384a  and  a46371a );
 a2176a <=( a46360a  and  a46347a );
 a2177a <=( a46336a  and  a46323a );
 a2178a <=( a46312a  and  a46299a );
 a2179a <=( a46288a  and  a46275a );
 a2180a <=( a46264a  and  a46251a );
 a2181a <=( a46240a  and  a46227a );
 a2182a <=( a46216a  and  a46203a );
 a2183a <=( a46192a  and  a46179a );
 a2184a <=( a46168a  and  a46155a );
 a2185a <=( a46144a  and  a46131a );
 a2186a <=( a46120a  and  a46107a );
 a2187a <=( a46096a  and  a46083a );
 a2188a <=( a46072a  and  a46059a );
 a2189a <=( a46048a  and  a46035a );
 a2190a <=( a46024a  and  a46011a );
 a2191a <=( a46000a  and  a45987a );
 a2192a <=( a45976a  and  a45963a );
 a2193a <=( a45952a  and  a45939a );
 a2194a <=( a45928a  and  a45915a );
 a2195a <=( a45904a  and  a45891a );
 a2196a <=( a45880a  and  a45867a );
 a2197a <=( a45856a  and  a45843a );
 a2198a <=( a45832a  and  a45819a );
 a2199a <=( a45808a  and  a45795a );
 a2200a <=( a45784a  and  a45771a );
 a2201a <=( a45760a  and  a45747a );
 a2202a <=( a45736a  and  a45723a );
 a2203a <=( a45712a  and  a45699a );
 a2204a <=( a45688a  and  a45675a );
 a2205a <=( a45664a  and  a45651a );
 a2206a <=( a45640a  and  a45627a );
 a2207a <=( a45616a  and  a45603a );
 a2208a <=( a45592a  and  a45579a );
 a2209a <=( a45568a  and  a45555a );
 a2210a <=( a45544a  and  a45531a );
 a2211a <=( a45520a  and  a45507a );
 a2212a <=( a45496a  and  a45483a );
 a2213a <=( a45472a  and  a45459a );
 a2214a <=( a45448a  and  a45435a );
 a2215a <=( a45424a  and  a45411a );
 a2216a <=( a45400a  and  a45387a );
 a2217a <=( a45376a  and  a45363a );
 a2218a <=( a45352a  and  a45339a );
 a2219a <=( a45328a  and  a45315a );
 a2220a <=( a45304a  and  a45291a );
 a2221a <=( a45280a  and  a45267a );
 a2222a <=( a45256a  and  a45243a );
 a2223a <=( a45232a  and  a45219a );
 a2224a <=( a45208a  and  a45195a );
 a2225a <=( a45184a  and  a45171a );
 a2226a <=( a45160a  and  a45147a );
 a2227a <=( a45136a  and  a45123a );
 a2228a <=( a45112a  and  a45099a );
 a2229a <=( a45088a  and  a45075a );
 a2230a <=( a45064a  and  a45051a );
 a2231a <=( a45040a  and  a45027a );
 a2232a <=( a45016a  and  a45003a );
 a2233a <=( a44992a  and  a44979a );
 a2234a <=( a44968a  and  a44955a );
 a2235a <=( a44944a  and  a44931a );
 a2236a <=( a44920a  and  a44907a );
 a2237a <=( a44896a  and  a44883a );
 a2238a <=( a44872a  and  a44859a );
 a2239a <=( a44848a  and  a44835a );
 a2240a <=( a44824a  and  a44811a );
 a2241a <=( a44800a  and  a44787a );
 a2242a <=( a44776a  and  a44763a );
 a2243a <=( a44752a  and  a44739a );
 a2244a <=( a44728a  and  a44715a );
 a2245a <=( a44704a  and  a44691a );
 a2246a <=( a44680a  and  a44667a );
 a2247a <=( a44656a  and  a44643a );
 a2248a <=( a44632a  and  a44619a );
 a2249a <=( a44608a  and  a44595a );
 a2250a <=( a44584a  and  a44571a );
 a2251a <=( a44560a  and  a44547a );
 a2252a <=( a44536a  and  a44523a );
 a2253a <=( a44512a  and  a44499a );
 a2254a <=( a44488a  and  a44475a );
 a2255a <=( a44464a  and  a44451a );
 a2256a <=( a44440a  and  a44427a );
 a2257a <=( a44416a  and  a44403a );
 a2258a <=( a44392a  and  a44379a );
 a2259a <=( a44368a  and  a44355a );
 a2260a <=( a44344a  and  a44331a );
 a2261a <=( a44320a  and  a44307a );
 a2262a <=( a44296a  and  a44283a );
 a2263a <=( a44272a  and  a44259a );
 a2264a <=( a44248a  and  a44235a );
 a2265a <=( a44224a  and  a44211a );
 a2266a <=( a44200a  and  a44187a );
 a2267a <=( a44176a  and  a44163a );
 a2268a <=( a44152a  and  a44139a );
 a2269a <=( a44128a  and  a44115a );
 a2270a <=( a44104a  and  a44091a );
 a2271a <=( a44080a  and  a44067a );
 a2272a <=( a44056a  and  a44043a );
 a2273a <=( a44032a  and  a44019a );
 a2274a <=( a44008a  and  a43995a );
 a2275a <=( a43984a  and  a43971a );
 a2276a <=( a43960a  and  a43947a );
 a2277a <=( a43936a  and  a43923a );
 a2278a <=( a43912a  and  a43899a );
 a2279a <=( a43888a  and  a43875a );
 a2280a <=( a43864a  and  a43851a );
 a2281a <=( a43840a  and  a43827a );
 a2282a <=( a43816a  and  a43803a );
 a2283a <=( a43792a  and  a43779a );
 a2284a <=( a43768a  and  a43755a );
 a2285a <=( a43744a  and  a43731a );
 a2286a <=( a43720a  and  a43707a );
 a2287a <=( a43696a  and  a43683a );
 a2288a <=( a43672a  and  a43659a );
 a2289a <=( a43648a  and  a43635a );
 a2290a <=( a43624a  and  a43611a );
 a2291a <=( a43600a  and  a43587a );
 a2292a <=( a43576a  and  a43563a );
 a2293a <=( a43552a  and  a43539a );
 a2294a <=( a43528a  and  a43515a );
 a2295a <=( a43504a  and  a43491a );
 a2296a <=( a43480a  and  a43467a );
 a2297a <=( a43456a  and  a43443a );
 a2298a <=( a43432a  and  a43419a );
 a2299a <=( a43408a  and  a43395a );
 a2300a <=( a43384a  and  a43371a );
 a2301a <=( a43360a  and  a43347a );
 a2302a <=( a43336a  and  a43323a );
 a2303a <=( a43312a  and  a43299a );
 a2304a <=( a43288a  and  a43275a );
 a2305a <=( a43264a  and  a43251a );
 a2306a <=( a43240a  and  a43227a );
 a2307a <=( a43216a  and  a43203a );
 a2308a <=( a43192a  and  a43179a );
 a2309a <=( a43168a  and  a43155a );
 a2310a <=( a43144a  and  a43131a );
 a2311a <=( a43120a  and  a43107a );
 a2312a <=( a43096a  and  a43083a );
 a2313a <=( a43072a  and  a43059a );
 a2314a <=( a43048a  and  a43035a );
 a2315a <=( a43024a  and  a43011a );
 a2316a <=( a43000a  and  a42987a );
 a2317a <=( a42976a  and  a42963a );
 a2318a <=( a42952a  and  a42939a );
 a2319a <=( a42928a  and  a42915a );
 a2320a <=( a42904a  and  a42891a );
 a2321a <=( a42880a  and  a42867a );
 a2322a <=( a42856a  and  a42843a );
 a2323a <=( a42832a  and  a42819a );
 a2324a <=( a42808a  and  a42795a );
 a2325a <=( a42784a  and  a42771a );
 a2326a <=( a42760a  and  a42747a );
 a2327a <=( a42736a  and  a42723a );
 a2328a <=( a42712a  and  a42699a );
 a2329a <=( a42688a  and  a42675a );
 a2330a <=( a42664a  and  a42651a );
 a2331a <=( a42640a  and  a42627a );
 a2332a <=( a42616a  and  a42603a );
 a2333a <=( a42592a  and  a42579a );
 a2334a <=( a42568a  and  a42555a );
 a2335a <=( a42544a  and  a42531a );
 a2336a <=( a42520a  and  a42507a );
 a2337a <=( a42496a  and  a42483a );
 a2338a <=( a42472a  and  a42459a );
 a2339a <=( a42448a  and  a42435a );
 a2340a <=( a42424a  and  a42411a );
 a2341a <=( a42400a  and  a42387a );
 a2342a <=( a42376a  and  a42363a );
 a2343a <=( a42352a  and  a42339a );
 a2344a <=( a42328a  and  a42315a );
 a2345a <=( a42304a  and  a42291a );
 a2346a <=( a42280a  and  a42267a );
 a2347a <=( a42256a  and  a42243a );
 a2348a <=( a42232a  and  a42219a );
 a2349a <=( a42208a  and  a42195a );
 a2350a <=( a42184a  and  a42171a );
 a2351a <=( a42160a  and  a42147a );
 a2352a <=( a42136a  and  a42123a );
 a2353a <=( a42112a  and  a42099a );
 a2354a <=( a42088a  and  a42075a );
 a2355a <=( a42064a  and  a42051a );
 a2356a <=( a42040a  and  a42027a );
 a2357a <=( a42016a  and  a42003a );
 a2358a <=( a41992a  and  a41979a );
 a2359a <=( a41968a  and  a41955a );
 a2360a <=( a41944a  and  a41931a );
 a2361a <=( a41920a  and  a41907a );
 a2362a <=( a41896a  and  a41883a );
 a2363a <=( a41872a  and  a41859a );
 a2364a <=( a41848a  and  a41835a );
 a2365a <=( a41824a  and  a41811a );
 a2366a <=( a41800a  and  a41787a );
 a2367a <=( a41776a  and  a41763a );
 a2368a <=( a41752a  and  a41739a );
 a2369a <=( a41728a  and  a41715a );
 a2370a <=( a41704a  and  a41691a );
 a2371a <=( a41680a  and  a41667a );
 a2372a <=( a41656a  and  a41643a );
 a2373a <=( a41632a  and  a41619a );
 a2374a <=( a41608a  and  a41595a );
 a2375a <=( a41584a  and  a41571a );
 a2376a <=( a41560a  and  a41547a );
 a2377a <=( a41536a  and  a41523a );
 a2378a <=( a41512a  and  a41499a );
 a2379a <=( a41488a  and  a41475a );
 a2380a <=( a41464a  and  a41451a );
 a2381a <=( a41440a  and  a41427a );
 a2382a <=( a41416a  and  a41403a );
 a2383a <=( a41392a  and  a41379a );
 a2384a <=( a41368a  and  a41355a );
 a2385a <=( a41344a  and  a41331a );
 a2386a <=( a41320a  and  a41307a );
 a2387a <=( a41296a  and  a41283a );
 a2388a <=( a41272a  and  a41259a );
 a2389a <=( a41248a  and  a41235a );
 a2390a <=( a41224a  and  a41211a );
 a2391a <=( a41200a  and  a41187a );
 a2392a <=( a41176a  and  a41163a );
 a2393a <=( a41152a  and  a41139a );
 a2394a <=( a41128a  and  a41115a );
 a2395a <=( a41104a  and  a41091a );
 a2396a <=( a41080a  and  a41067a );
 a2397a <=( a41056a  and  a41043a );
 a2398a <=( a41032a  and  a41019a );
 a2399a <=( a41008a  and  a40995a );
 a2400a <=( a40984a  and  a40971a );
 a2401a <=( a40960a  and  a40947a );
 a2402a <=( a40936a  and  a40923a );
 a2403a <=( a40912a  and  a40899a );
 a2404a <=( a40888a  and  a40875a );
 a2405a <=( a40864a  and  a40851a );
 a2406a <=( a40840a  and  a40827a );
 a2407a <=( a40816a  and  a40803a );
 a2408a <=( a40792a  and  a40779a );
 a2409a <=( a40768a  and  a40755a );
 a2410a <=( a40744a  and  a40731a );
 a2411a <=( a40720a  and  a40707a );
 a2412a <=( a40696a  and  a40683a );
 a2413a <=( a40672a  and  a40659a );
 a2414a <=( a40648a  and  a40635a );
 a2415a <=( a40624a  and  a40611a );
 a2416a <=( a40600a  and  a40587a );
 a2417a <=( a40576a  and  a40563a );
 a2418a <=( a40552a  and  a40539a );
 a2419a <=( a40528a  and  a40515a );
 a2420a <=( a40504a  and  a40491a );
 a2421a <=( a40480a  and  a40467a );
 a2422a <=( a40456a  and  a40443a );
 a2423a <=( a40432a  and  a40419a );
 a2424a <=( a40408a  and  a40395a );
 a2425a <=( a40384a  and  a40371a );
 a2426a <=( a40360a  and  a40347a );
 a2427a <=( a40336a  and  a40325a );
 a2428a <=( a40314a  and  a40303a );
 a2429a <=( a40292a  and  a40281a );
 a2430a <=( a40270a  and  a40259a );
 a2431a <=( a40248a  and  a40237a );
 a2432a <=( a40226a  and  a40215a );
 a2433a <=( a40204a  and  a40193a );
 a2434a <=( a40182a  and  a40171a );
 a2435a <=( a40160a  and  a40149a );
 a2436a <=( a40138a  and  a40127a );
 a2437a <=( a40116a  and  a40105a );
 a2438a <=( a40094a  and  a40083a );
 a2439a <=( a40072a  and  a40061a );
 a2440a <=( a40050a  and  a40039a );
 a2441a <=( a40028a  and  a40017a );
 a2442a <=( a40006a  and  a39995a );
 a2443a <=( a39984a  and  a39973a );
 a2444a <=( a39962a  and  a39951a );
 a2445a <=( a39940a  and  a39929a );
 a2446a <=( a39918a  and  a39907a );
 a2447a <=( a39896a  and  a39885a );
 a2448a <=( a39874a  and  a39863a );
 a2449a <=( a39852a  and  a39841a );
 a2450a <=( a39830a  and  a39819a );
 a2451a <=( a39808a  and  a39797a );
 a2452a <=( a39786a  and  a39775a );
 a2453a <=( a39764a  and  a39753a );
 a2454a <=( a39742a  and  a39731a );
 a2455a <=( a39720a  and  a39709a );
 a2456a <=( a39698a  and  a39687a );
 a2457a <=( a39676a  and  a39665a );
 a2458a <=( a39654a  and  a39643a );
 a2459a <=( a39632a  and  a39621a );
 a2460a <=( a39610a  and  a39599a );
 a2461a <=( a39588a  and  a39577a );
 a2462a <=( a39566a  and  a39555a );
 a2463a <=( a39544a  and  a39533a );
 a2464a <=( a39522a  and  a39511a );
 a2465a <=( a39500a  and  a39489a );
 a2466a <=( a39478a  and  a39467a );
 a2467a <=( a39456a  and  a39445a );
 a2468a <=( a39434a  and  a39423a );
 a2469a <=( a39412a  and  a39401a );
 a2470a <=( a39390a  and  a39379a );
 a2471a <=( a39368a  and  a39357a );
 a2472a <=( a39346a  and  a39335a );
 a2473a <=( a39324a  and  a39313a );
 a2474a <=( a39302a  and  a39291a );
 a2475a <=( a39280a  and  a39269a );
 a2476a <=( a39258a  and  a39247a );
 a2477a <=( a39236a  and  a39225a );
 a2478a <=( a39214a  and  a39203a );
 a2479a <=( a39192a  and  a39181a );
 a2480a <=( a39170a  and  a39159a );
 a2481a <=( a39148a  and  a39137a );
 a2482a <=( a39126a  and  a39115a );
 a2483a <=( a39104a  and  a39093a );
 a2484a <=( a39082a  and  a39071a );
 a2485a <=( a39060a  and  a39049a );
 a2486a <=( a39038a  and  a39027a );
 a2487a <=( a39016a  and  a39005a );
 a2488a <=( a38994a  and  a38983a );
 a2489a <=( a38972a  and  a38961a );
 a2490a <=( a38950a  and  a38939a );
 a2491a <=( a38928a  and  a38917a );
 a2492a <=( a38906a  and  a38895a );
 a2493a <=( a38884a  and  a38873a );
 a2494a <=( a38862a  and  a38851a );
 a2495a <=( a38840a  and  a38829a );
 a2496a <=( a38818a  and  a38807a );
 a2497a <=( a38796a  and  a38785a );
 a2498a <=( a38774a  and  a38763a );
 a2499a <=( a38752a  and  a38741a );
 a2500a <=( a38730a  and  a38719a );
 a2501a <=( a38708a  and  a38697a );
 a2502a <=( a38686a  and  a38675a );
 a2503a <=( a38664a  and  a38653a );
 a2504a <=( a38642a  and  a38631a );
 a2505a <=( a38620a  and  a38609a );
 a2506a <=( a38598a  and  a38587a );
 a2507a <=( a38576a  and  a38565a );
 a2508a <=( a38554a  and  a38543a );
 a2509a <=( a38532a  and  a38521a );
 a2510a <=( a38510a  and  a38499a );
 a2511a <=( a38488a  and  a38477a );
 a2512a <=( a38466a  and  a38455a );
 a2513a <=( a38444a  and  a38433a );
 a2514a <=( a38422a  and  a38411a );
 a2515a <=( a38400a  and  a38389a );
 a2516a <=( a38378a  and  a38367a );
 a2517a <=( a38356a  and  a38345a );
 a2518a <=( a38334a  and  a38323a );
 a2519a <=( a38312a  and  a38301a );
 a2520a <=( a38290a  and  a38279a );
 a2521a <=( a38268a  and  a38257a );
 a2522a <=( a38246a  and  a38235a );
 a2523a <=( a38224a  and  a38213a );
 a2524a <=( a38202a  and  a38191a );
 a2525a <=( a38180a  and  a38169a );
 a2526a <=( a38158a  and  a38147a );
 a2527a <=( a38136a  and  a38125a );
 a2528a <=( a38114a  and  a38103a );
 a2529a <=( a38092a  and  a38081a );
 a2530a <=( a38070a  and  a38059a );
 a2531a <=( a38048a  and  a38037a );
 a2532a <=( a38026a  and  a38015a );
 a2533a <=( a38004a  and  a37993a );
 a2534a <=( a37982a  and  a37971a );
 a2535a <=( a37960a  and  a37949a );
 a2536a <=( a37938a  and  a37927a );
 a2537a <=( a37916a  and  a37905a );
 a2538a <=( a37894a  and  a37883a );
 a2539a <=( a37872a  and  a37861a );
 a2540a <=( a37850a  and  a37839a );
 a2541a <=( a37828a  and  a37817a );
 a2542a <=( a37806a  and  a37795a );
 a2543a <=( a37784a  and  a37773a );
 a2544a <=( a37762a  and  a37751a );
 a2545a <=( a37740a  and  a37729a );
 a2546a <=( a37718a  and  a37707a );
 a2547a <=( a37696a  and  a37685a );
 a2548a <=( a37674a  and  a37663a );
 a2549a <=( a37652a  and  a37641a );
 a2550a <=( a37630a  and  a37619a );
 a2551a <=( a37608a  and  a37597a );
 a2552a <=( a37586a  and  a37575a );
 a2553a <=( a37564a  and  a37553a );
 a2554a <=( a37542a  and  a37531a );
 a2555a <=( a37520a  and  a37509a );
 a2556a <=( a37498a  and  a37487a );
 a2557a <=( a37476a  and  a37465a );
 a2558a <=( a37454a  and  a37443a );
 a2559a <=( a37432a  and  a37421a );
 a2560a <=( a37410a  and  a37399a );
 a2561a <=( a37388a  and  a37377a );
 a2562a <=( a37366a  and  a37355a );
 a2563a <=( a37344a  and  a37333a );
 a2564a <=( a37322a  and  a37311a );
 a2565a <=( a37300a  and  a37289a );
 a2566a <=( a37278a  and  a37267a );
 a2567a <=( a37256a  and  a37245a );
 a2568a <=( a37234a  and  a37223a );
 a2569a <=( a37212a  and  a37201a );
 a2570a <=( a37190a  and  a37179a );
 a2571a <=( a37168a  and  a37157a );
 a2572a <=( a37146a  and  a37135a );
 a2573a <=( a37124a  and  a37113a );
 a2574a <=( a37102a  and  a37091a );
 a2575a <=( a37080a  and  a37069a );
 a2576a <=( a37058a  and  a37047a );
 a2577a <=( a37036a  and  a37025a );
 a2578a <=( a37014a  and  a37003a );
 a2579a <=( a36992a  and  a36981a );
 a2580a <=( a36970a  and  a36959a );
 a2581a <=( a36948a  and  a36937a );
 a2582a <=( a36926a  and  a36915a );
 a2583a <=( a36904a  and  a36893a );
 a2584a <=( a36882a  and  a36871a );
 a2585a <=( a36860a  and  a36849a );
 a2586a <=( a36838a  and  a36827a );
 a2587a <=( a36816a  and  a36805a );
 a2588a <=( a36794a  and  a36783a );
 a2589a <=( a36772a  and  a36761a );
 a2590a <=( a36750a  and  a36739a );
 a2591a <=( a36728a  and  a36717a );
 a2592a <=( a36706a  and  a36695a );
 a2593a <=( a36684a  and  a36673a );
 a2594a <=( a36662a  and  a36651a );
 a2595a <=( a36640a  and  a36629a );
 a2596a <=( a36618a  and  a36607a );
 a2597a <=( a36596a  and  a36585a );
 a2598a <=( a36574a  and  a36563a );
 a2599a <=( a36552a  and  a36541a );
 a2600a <=( a36530a  and  a36519a );
 a2601a <=( a36508a  and  a36497a );
 a2602a <=( a36486a  and  a36475a );
 a2603a <=( a36464a  and  a36453a );
 a2604a <=( a36442a  and  a36431a );
 a2605a <=( a36420a  and  a36409a );
 a2606a <=( a36398a  and  a36387a );
 a2607a <=( a36376a  and  a36365a );
 a2608a <=( a36354a  and  a36343a );
 a2609a <=( a36332a  and  a36321a );
 a2610a <=( a36310a  and  a36299a );
 a2611a <=( a36288a  and  a36277a );
 a2612a <=( a36266a  and  a36255a );
 a2613a <=( a36244a  and  a36233a );
 a2614a <=( a36222a  and  a36211a );
 a2615a <=( a36200a  and  a36189a );
 a2616a <=( a36178a  and  a36167a );
 a2617a <=( a36156a  and  a36145a );
 a2618a <=( a36134a  and  a36123a );
 a2619a <=( a36112a  and  a36101a );
 a2620a <=( a36090a  and  a36079a );
 a2621a <=( a36068a  and  a36057a );
 a2622a <=( a36046a  and  a36035a );
 a2623a <=( a36024a  and  a36013a );
 a2624a <=( a36002a  and  a35991a );
 a2625a <=( a35980a  and  a35969a );
 a2626a <=( a35958a  and  a35947a );
 a2627a <=( a35936a  and  a35925a );
 a2628a <=( a35914a  and  a35903a );
 a2629a <=( a35892a  and  a35881a );
 a2630a <=( a35870a  and  a35859a );
 a2631a <=( a35848a  and  a35837a );
 a2632a <=( a35826a  and  a35815a );
 a2633a <=( a35804a  and  a35793a );
 a2634a <=( a35782a  and  a35771a );
 a2635a <=( a35760a  and  a35749a );
 a2636a <=( a35738a  and  a35727a );
 a2637a <=( a35716a  and  a35705a );
 a2638a <=( a35694a  and  a35683a );
 a2639a <=( a35672a  and  a35661a );
 a2640a <=( a35650a  and  a35639a );
 a2641a <=( a35628a  and  a35617a );
 a2642a <=( a35606a  and  a35595a );
 a2643a <=( a35584a  and  a35573a );
 a2644a <=( a35562a  and  a35551a );
 a2645a <=( a35540a  and  a35529a );
 a2646a <=( a35518a  and  a35507a );
 a2647a <=( a35496a  and  a35485a );
 a2648a <=( a35474a  and  a35463a );
 a2649a <=( a35452a  and  a35441a );
 a2650a <=( a35430a  and  a35419a );
 a2651a <=( a35408a  and  a35397a );
 a2652a <=( a35386a  and  a35375a );
 a2653a <=( a35364a  and  a35353a );
 a2654a <=( a35342a  and  a35331a );
 a2655a <=( a35320a  and  a35309a );
 a2656a <=( a35298a  and  a35287a );
 a2657a <=( a35276a  and  a35265a );
 a2658a <=( a35254a  and  a35243a );
 a2659a <=( a35232a  and  a35221a );
 a2660a <=( a35210a  and  a35199a );
 a2661a <=( a35188a  and  a35177a );
 a2662a <=( a35166a  and  a35155a );
 a2663a <=( a35144a  and  a35133a );
 a2664a <=( a35122a  and  a35111a );
 a2665a <=( a35100a  and  a35089a );
 a2666a <=( a35078a  and  a35067a );
 a2667a <=( a35056a  and  a35045a );
 a2668a <=( a35034a  and  a35023a );
 a2669a <=( a35012a  and  a35001a );
 a2670a <=( a34990a  and  a34979a );
 a2671a <=( a34968a  and  a34957a );
 a2672a <=( a34946a  and  a34935a );
 a2673a <=( a34924a  and  a34913a );
 a2674a <=( a34902a  and  a34891a );
 a2675a <=( a34880a  and  a34869a );
 a2676a <=( a34858a  and  a34847a );
 a2677a <=( a34836a  and  a34825a );
 a2678a <=( a34814a  and  a34803a );
 a2679a <=( a34792a  and  a34781a );
 a2680a <=( a34770a  and  a34759a );
 a2681a <=( a34748a  and  a34737a );
 a2682a <=( a34726a  and  a34715a );
 a2683a <=( a34704a  and  a34693a );
 a2684a <=( a34682a  and  a34671a );
 a2685a <=( a34660a  and  a34649a );
 a2686a <=( a34638a  and  a34627a );
 a2687a <=( a34616a  and  a34605a );
 a2688a <=( a34594a  and  a34583a );
 a2689a <=( a34572a  and  a34561a );
 a2690a <=( a34550a  and  a34539a );
 a2691a <=( a34528a  and  a34517a );
 a2692a <=( a34506a  and  a34495a );
 a2693a <=( a34484a  and  a34473a );
 a2694a <=( a34462a  and  a34451a );
 a2695a <=( a34440a  and  a34429a );
 a2696a <=( a34418a  and  a34407a );
 a2697a <=( a34396a  and  a34385a );
 a2698a <=( a34374a  and  a34363a );
 a2699a <=( a34352a  and  a34341a );
 a2700a <=( a34330a  and  a34319a );
 a2701a <=( a34308a  and  a34297a );
 a2702a <=( a34286a  and  a34275a );
 a2703a <=( a34264a  and  a34253a );
 a2704a <=( a34242a  and  a34231a );
 a2705a <=( a34220a  and  a34209a );
 a2706a <=( a34198a  and  a34187a );
 a2707a <=( a34176a  and  a34165a );
 a2708a <=( a34154a  and  a34143a );
 a2709a <=( a34132a  and  a34121a );
 a2710a <=( a34110a  and  a34099a );
 a2711a <=( a34088a  and  a34077a );
 a2712a <=( a34066a  and  a34055a );
 a2713a <=( a34044a  and  a34033a );
 a2714a <=( a34022a  and  a34011a );
 a2715a <=( a34000a  and  a33989a );
 a2716a <=( a33978a  and  a33967a );
 a2717a <=( a33956a  and  a33945a );
 a2718a <=( a33934a  and  a33923a );
 a2719a <=( a33912a  and  a33901a );
 a2720a <=( a33890a  and  a33879a );
 a2721a <=( a33868a  and  a33857a );
 a2722a <=( a33846a  and  a33835a );
 a2723a <=( a33824a  and  a33813a );
 a2724a <=( a33802a  and  a33791a );
 a2725a <=( a33780a  and  a33769a );
 a2726a <=( a33758a  and  a33747a );
 a2727a <=( a33736a  and  a33725a );
 a2728a <=( a33714a  and  a33703a );
 a2729a <=( a33692a  and  a33681a );
 a2730a <=( a33670a  and  a33659a );
 a2731a <=( a33648a  and  a33637a );
 a2732a <=( a33626a  and  a33615a );
 a2733a <=( a33604a  and  a33593a );
 a2734a <=( a33582a  and  a33571a );
 a2735a <=( a33560a  and  a33549a );
 a2736a <=( a33538a  and  a33527a );
 a2737a <=( a33516a  and  a33505a );
 a2738a <=( a33494a  and  a33483a );
 a2739a <=( a33472a  and  a33461a );
 a2740a <=( a33450a  and  a33439a );
 a2741a <=( a33428a  and  a33417a );
 a2742a <=( a33406a  and  a33395a );
 a2743a <=( a33384a  and  a33373a );
 a2744a <=( a33362a  and  a33351a );
 a2745a <=( a33340a  and  a33329a );
 a2746a <=( a33318a  and  a33307a );
 a2747a <=( a33296a  and  a33285a );
 a2748a <=( a33274a  and  a33263a );
 a2749a <=( a33252a  and  a33241a );
 a2750a <=( a33230a  and  a33219a );
 a2751a <=( a33208a  and  a33197a );
 a2752a <=( a33186a  and  a33175a );
 a2753a <=( a33164a  and  a33153a );
 a2754a <=( a33142a  and  a33131a );
 a2755a <=( a33120a  and  a33109a );
 a2756a <=( a33098a  and  a33087a );
 a2757a <=( a33076a  and  a33065a );
 a2758a <=( a33054a  and  a33043a );
 a2759a <=( a33032a  and  a33021a );
 a2760a <=( a33010a  and  a32999a );
 a2761a <=( a32988a  and  a32977a );
 a2762a <=( a32966a  and  a32955a );
 a2763a <=( a32944a  and  a32933a );
 a2764a <=( a32922a  and  a32911a );
 a2765a <=( a32900a  and  a32889a );
 a2766a <=( a32878a  and  a32867a );
 a2767a <=( a32856a  and  a32845a );
 a2768a <=( a32834a  and  a32823a );
 a2769a <=( a32812a  and  a32801a );
 a2770a <=( a32790a  and  a32779a );
 a2771a <=( a32768a  and  a32757a );
 a2772a <=( a32746a  and  a32735a );
 a2773a <=( a32724a  and  a32713a );
 a2774a <=( a32702a  and  a32691a );
 a2775a <=( a32680a  and  a32669a );
 a2776a <=( a32658a  and  a32647a );
 a2777a <=( a32636a  and  a32625a );
 a2778a <=( a32614a  and  a32603a );
 a2779a <=( a32592a  and  a32581a );
 a2780a <=( a32570a  and  a32559a );
 a2781a <=( a32548a  and  a32537a );
 a2782a <=( a32526a  and  a32515a );
 a2783a <=( a32504a  and  a32493a );
 a2784a <=( a32482a  and  a32471a );
 a2785a <=( a32460a  and  a32449a );
 a2786a <=( a32438a  and  a32427a );
 a2787a <=( a32416a  and  a32405a );
 a2788a <=( a32394a  and  a32383a );
 a2789a <=( a32372a  and  a32361a );
 a2790a <=( a32350a  and  a32339a );
 a2791a <=( a32328a  and  a32317a );
 a2792a <=( a32306a  and  a32295a );
 a2793a <=( a32284a  and  a32273a );
 a2794a <=( a32262a  and  a32251a );
 a2795a <=( a32240a  and  a32229a );
 a2796a <=( a32218a  and  a32207a );
 a2797a <=( a32196a  and  a32185a );
 a2798a <=( a32174a  and  a32163a );
 a2799a <=( a32152a  and  a32141a );
 a2800a <=( a32130a  and  a32119a );
 a2801a <=( a32108a  and  a32097a );
 a2802a <=( a32086a  and  a32075a );
 a2803a <=( a32064a  and  a32053a );
 a2804a <=( a32042a  and  a32031a );
 a2805a <=( a32020a  and  a32009a );
 a2806a <=( a31998a  and  a31987a );
 a2807a <=( a31976a  and  a31965a );
 a2808a <=( a31954a  and  a31943a );
 a2809a <=( a31932a  and  a31921a );
 a2810a <=( a31910a  and  a31899a );
 a2811a <=( a31888a  and  a31877a );
 a2812a <=( a31866a  and  a31855a );
 a2813a <=( a31844a  and  a31833a );
 a2814a <=( a31822a  and  a31811a );
 a2815a <=( a31800a  and  a31789a );
 a2816a <=( a31778a  and  a31767a );
 a2817a <=( a31756a  and  a31745a );
 a2818a <=( a31734a  and  a31723a );
 a2819a <=( a31712a  and  a31701a );
 a2820a <=( a31690a  and  a31679a );
 a2821a <=( a31668a  and  a31657a );
 a2822a <=( a31646a  and  a31635a );
 a2823a <=( a31624a  and  a31613a );
 a2824a <=( a31602a  and  a31591a );
 a2825a <=( a31580a  and  a31569a );
 a2826a <=( a31558a  and  a31547a );
 a2827a <=( a31536a  and  a31525a );
 a2828a <=( a31514a  and  a31503a );
 a2829a <=( a31492a  and  a31481a );
 a2830a <=( a31470a  and  a31459a );
 a2831a <=( a31448a  and  a31437a );
 a2832a <=( a31426a  and  a31415a );
 a2833a <=( a31404a  and  a31393a );
 a2834a <=( a31382a  and  a31371a );
 a2835a <=( a31360a  and  a31349a );
 a2836a <=( a31338a  and  a31327a );
 a2837a <=( a31316a  and  a31305a );
 a2838a <=( a31294a  and  a31283a );
 a2839a <=( a31272a  and  a31261a );
 a2840a <=( a31250a  and  a31239a );
 a2841a <=( a31228a  and  a31217a );
 a2842a <=( a31206a  and  a31195a );
 a2843a <=( a31184a  and  a31173a );
 a2844a <=( a31162a  and  a31151a );
 a2845a <=( a31140a  and  a31129a );
 a2846a <=( a31118a  and  a31107a );
 a2847a <=( a31096a  and  a31085a );
 a2848a <=( a31074a  and  a31063a );
 a2849a <=( a31052a  and  a31041a );
 a2850a <=( a31030a  and  a31019a );
 a2851a <=( a31008a  and  a30997a );
 a2852a <=( a30986a  and  a30975a );
 a2853a <=( a30964a  and  a30953a );
 a2854a <=( a30942a  and  a30931a );
 a2855a <=( a30920a  and  a30909a );
 a2856a <=( a30898a  and  a30887a );
 a2857a <=( a30876a  and  a30865a );
 a2858a <=( a30854a  and  a30843a );
 a2859a <=( a30832a  and  a30821a );
 a2860a <=( a30810a  and  a30799a );
 a2861a <=( a30788a  and  a30777a );
 a2862a <=( a30766a  and  a30755a );
 a2863a <=( a30744a  and  a30733a );
 a2864a <=( a30722a  and  a30711a );
 a2865a <=( a30700a  and  a30689a );
 a2866a <=( a30678a  and  a30667a );
 a2867a <=( a30656a  and  a30645a );
 a2868a <=( a30634a  and  a30623a );
 a2869a <=( a30612a  and  a30601a );
 a2870a <=( a30590a  and  a30579a );
 a2871a <=( a30568a  and  a30557a );
 a2872a <=( a30546a  and  a30535a );
 a2873a <=( a30524a  and  a30513a );
 a2874a <=( a30502a  and  a30491a );
 a2875a <=( a30480a  and  a30469a );
 a2876a <=( a30458a  and  a30447a );
 a2877a <=( a30436a  and  a30425a );
 a2878a <=( a30414a  and  a30403a );
 a2879a <=( a30392a  and  a30381a );
 a2880a <=( a30370a  and  a30359a );
 a2881a <=( a30348a  and  a30337a );
 a2882a <=( a30326a  and  a30315a );
 a2883a <=( a30304a  and  a30293a );
 a2884a <=( a30282a  and  a30271a );
 a2885a <=( a30260a  and  a30249a );
 a2886a <=( a30238a  and  a30227a );
 a2887a <=( a30216a  and  a30205a );
 a2888a <=( a30194a  and  a30183a );
 a2889a <=( a30172a  and  a30161a );
 a2890a <=( a30150a  and  a30139a );
 a2891a <=( a30128a  and  a30117a );
 a2892a <=( a30106a  and  a30095a );
 a2893a <=( a30084a  and  a30073a );
 a2894a <=( a30062a  and  a30051a );
 a2895a <=( a30040a  and  a30029a );
 a2896a <=( a30018a  and  a30007a );
 a2897a <=( a29996a  and  a29985a );
 a2898a <=( a29974a  and  a29963a );
 a2899a <=( a29952a  and  a29941a );
 a2900a <=( a29930a  and  a29919a );
 a2901a <=( a29908a  and  a29897a );
 a2902a <=( a29886a  and  a29875a );
 a2903a <=( a29864a  and  a29853a );
 a2904a <=( a29842a  and  a29831a );
 a2905a <=( a29820a  and  a29809a );
 a2906a <=( a29798a  and  a29787a );
 a2907a <=( a29776a  and  a29765a );
 a2908a <=( a29754a  and  a29743a );
 a2909a <=( a29732a  and  a29721a );
 a2910a <=( a29710a  and  a29699a );
 a2911a <=( a29688a  and  a29677a );
 a2912a <=( a29666a  and  a29655a );
 a2913a <=( a29644a  and  a29633a );
 a2914a <=( a29622a  and  a29611a );
 a2915a <=( a29600a  and  a29589a );
 a2916a <=( a29578a  and  a29567a );
 a2917a <=( a29556a  and  a29545a );
 a2918a <=( a29534a  and  a29523a );
 a2919a <=( a29512a  and  a29501a );
 a2920a <=( a29490a  and  a29479a );
 a2921a <=( a29468a  and  a29457a );
 a2922a <=( a29446a  and  a29435a );
 a2923a <=( a29424a  and  a29413a );
 a2924a <=( a29402a  and  a29391a );
 a2925a <=( a29380a  and  a29369a );
 a2926a <=( a29358a  and  a29347a );
 a2927a <=( a29336a  and  a29325a );
 a2928a <=( a29314a  and  a29303a );
 a2929a <=( a29292a  and  a29281a );
 a2930a <=( a29270a  and  a29259a );
 a2931a <=( a29248a  and  a29237a );
 a2932a <=( a29226a  and  a29215a );
 a2933a <=( a29204a  and  a29193a );
 a2934a <=( a29182a  and  a29171a );
 a2935a <=( a29160a  and  a29149a );
 a2936a <=( a29138a  and  a29127a );
 a2937a <=( a29116a  and  a29105a );
 a2938a <=( a29094a  and  a29083a );
 a2939a <=( a29072a  and  a29061a );
 a2940a <=( a29050a  and  a29039a );
 a2941a <=( a29028a  and  a29017a );
 a2942a <=( a29006a  and  a28995a );
 a2943a <=( a28984a  and  a28973a );
 a2944a <=( a28962a  and  a28951a );
 a2945a <=( a28940a  and  a28929a );
 a2946a <=( a28918a  and  a28907a );
 a2947a <=( a28896a  and  a28885a );
 a2948a <=( a28874a  and  a28863a );
 a2949a <=( a28852a  and  a28841a );
 a2950a <=( a28830a  and  a28819a );
 a2951a <=( a28808a  and  a28797a );
 a2952a <=( a28786a  and  a28775a );
 a2953a <=( a28764a  and  a28753a );
 a2954a <=( a28742a  and  a28731a );
 a2955a <=( a28720a  and  a28709a );
 a2956a <=( a28698a  and  a28687a );
 a2957a <=( a28676a  and  a28665a );
 a2958a <=( a28654a  and  a28643a );
 a2959a <=( a28632a  and  a28621a );
 a2960a <=( a28610a  and  a28599a );
 a2961a <=( a28588a  and  a28577a );
 a2962a <=( a28566a  and  a28555a );
 a2963a <=( a28544a  and  a28533a );
 a2964a <=( a28522a  and  a28511a );
 a2965a <=( a28500a  and  a28489a );
 a2966a <=( a28478a  and  a28467a );
 a2967a <=( a28456a  and  a28445a );
 a2968a <=( a28434a  and  a28423a );
 a2969a <=( a28412a  and  a28401a );
 a2970a <=( a28390a  and  a28379a );
 a2971a <=( a28368a  and  a28357a );
 a2972a <=( a28346a  and  a28335a );
 a2973a <=( a28324a  and  a28313a );
 a2974a <=( a28302a  and  a28291a );
 a2975a <=( a28280a  and  a28269a );
 a2976a <=( a28258a  and  a28247a );
 a2977a <=( a28236a  and  a28225a );
 a2978a <=( a28214a  and  a28203a );
 a2979a <=( a28192a  and  a28181a );
 a2980a <=( a28170a  and  a28159a );
 a2981a <=( a28148a  and  a28137a );
 a2982a <=( a28126a  and  a28115a );
 a2983a <=( a28104a  and  a28093a );
 a2984a <=( a28082a  and  a28071a );
 a2985a <=( a28060a  and  a28049a );
 a2986a <=( a28038a  and  a28027a );
 a2987a <=( a28016a  and  a28005a );
 a2988a <=( a27994a  and  a27983a );
 a2989a <=( a27972a  and  a27961a );
 a2990a <=( a27950a  and  a27939a );
 a2991a <=( a27928a  and  a27917a );
 a2992a <=( a27906a  and  a27895a );
 a2993a <=( a27884a  and  a27873a );
 a2994a <=( a27862a  and  a27851a );
 a2995a <=( a27840a  and  a27829a );
 a2996a <=( a27818a  and  a27807a );
 a2997a <=( a27796a  and  a27785a );
 a2998a <=( a27774a  and  a27763a );
 a2999a <=( a27752a  and  a27741a );
 a3000a <=( a27730a  and  a27719a );
 a3001a <=( a27708a  and  a27697a );
 a3002a <=( a27686a  and  a27675a );
 a3003a <=( a27664a  and  a27653a );
 a3004a <=( a27642a  and  a27631a );
 a3005a <=( a27620a  and  a27609a );
 a3006a <=( a27598a  and  a27587a );
 a3007a <=( a27576a  and  a27565a );
 a3008a <=( a27554a  and  a27543a );
 a3009a <=( a27532a  and  a27521a );
 a3010a <=( a27510a  and  a27499a );
 a3011a <=( a27488a  and  a27477a );
 a3012a <=( a27466a  and  a27455a );
 a3013a <=( a27444a  and  a27433a );
 a3014a <=( a27422a  and  a27411a );
 a3015a <=( a27400a  and  a27389a );
 a3016a <=( a27378a  and  a27367a );
 a3017a <=( a27356a  and  a27345a );
 a3018a <=( a27334a  and  a27323a );
 a3019a <=( a27312a  and  a27301a );
 a3020a <=( a27290a  and  a27279a );
 a3021a <=( a27268a  and  a27257a );
 a3022a <=( a27246a  and  a27235a );
 a3023a <=( a27224a  and  a27213a );
 a3024a <=( a27202a  and  a27191a );
 a3025a <=( a27180a  and  a27169a );
 a3026a <=( a27158a  and  a27147a );
 a3027a <=( a27136a  and  a27125a );
 a3028a <=( a27114a  and  a27103a );
 a3029a <=( a27092a  and  a27081a );
 a3030a <=( a27070a  and  a27059a );
 a3031a <=( a27048a  and  a27037a );
 a3032a <=( a27026a  and  a27015a );
 a3033a <=( a27004a  and  a26993a );
 a3034a <=( a26982a  and  a26971a );
 a3035a <=( a26960a  and  a26949a );
 a3036a <=( a26938a  and  a26927a );
 a3037a <=( a26916a  and  a26905a );
 a3038a <=( a26894a  and  a26883a );
 a3039a <=( a26872a  and  a26861a );
 a3040a <=( a26850a  and  a26839a );
 a3041a <=( a26828a  and  a26817a );
 a3042a <=( a26806a  and  a26795a );
 a3043a <=( a26784a  and  a26773a );
 a3044a <=( a26762a  and  a26751a );
 a3045a <=( a26740a  and  a26729a );
 a3046a <=( a26718a  and  a26707a );
 a3047a <=( a26696a  and  a26685a );
 a3048a <=( a26674a  and  a26663a );
 a3049a <=( a26652a  and  a26641a );
 a3050a <=( a26630a  and  a26619a );
 a3051a <=( a26608a  and  a26597a );
 a3052a <=( a26586a  and  a26575a );
 a3053a <=( a26564a  and  a26553a );
 a3054a <=( a26542a  and  a26531a );
 a3055a <=( a26520a  and  a26509a );
 a3056a <=( a26498a  and  a26487a );
 a3057a <=( a26476a  and  a26465a );
 a3058a <=( a26454a  and  a26443a );
 a3059a <=( a26432a  and  a26421a );
 a3060a <=( a26410a  and  a26399a );
 a3061a <=( a26388a  and  a26377a );
 a3062a <=( a26366a  and  a26355a );
 a3063a <=( a26344a  and  a26333a );
 a3064a <=( a26322a  and  a26311a );
 a3065a <=( a26300a  and  a26289a );
 a3066a <=( a26278a  and  a26267a );
 a3067a <=( a26256a  and  a26245a );
 a3068a <=( a26234a  and  a26223a );
 a3069a <=( a26212a  and  a26201a );
 a3070a <=( a26190a  and  a26179a );
 a3071a <=( a26168a  and  a26157a );
 a3072a <=( a26146a  and  a26135a );
 a3073a <=( a26124a  and  a26113a );
 a3074a <=( a26102a  and  a26091a );
 a3075a <=( a26080a  and  a26069a );
 a3076a <=( a26058a  and  a26047a );
 a3077a <=( a26036a  and  a26025a );
 a3078a <=( a26014a  and  a26003a );
 a3079a <=( a25992a  and  a25981a );
 a3080a <=( a25970a  and  a25959a );
 a3081a <=( a25948a  and  a25937a );
 a3082a <=( a25926a  and  a25915a );
 a3083a <=( a25904a  and  a25893a );
 a3084a <=( a25882a  and  a25871a );
 a3085a <=( a25860a  and  a25849a );
 a3086a <=( a25838a  and  a25827a );
 a3087a <=( a25816a  and  a25805a );
 a3088a <=( a25794a  and  a25783a );
 a3089a <=( a25772a  and  a25761a );
 a3090a <=( a25750a  and  a25739a );
 a3091a <=( a25728a  and  a25717a );
 a3092a <=( a25706a  and  a25695a );
 a3093a <=( a25684a  and  a25673a );
 a3094a <=( a25662a  and  a25651a );
 a3095a <=( a25640a  and  a25629a );
 a3096a <=( a25618a  and  a25607a );
 a3097a <=( a25596a  and  a25585a );
 a3098a <=( a25574a  and  a25563a );
 a3099a <=( a25552a  and  a25541a );
 a3100a <=( a25530a  and  a25519a );
 a3101a <=( a25508a  and  a25497a );
 a3102a <=( a25486a  and  a25475a );
 a3103a <=( a25464a  and  a25453a );
 a3104a <=( a25442a  and  a25431a );
 a3105a <=( a25420a  and  a25409a );
 a3106a <=( a25398a  and  a25387a );
 a3107a <=( a25376a  and  a25365a );
 a3108a <=( a25354a  and  a25343a );
 a3109a <=( a25332a  and  a25321a );
 a3110a <=( a25310a  and  a25299a );
 a3111a <=( a25288a  and  a25277a );
 a3112a <=( a25266a  and  a25255a );
 a3113a <=( a25244a  and  a25233a );
 a3114a <=( a25222a  and  a25211a );
 a3115a <=( a25200a  and  a25189a );
 a3116a <=( a25178a  and  a25167a );
 a3117a <=( a25156a  and  a25145a );
 a3118a <=( a25134a  and  a25123a );
 a3119a <=( a25112a  and  a25101a );
 a3120a <=( a25090a  and  a25079a );
 a3121a <=( a25068a  and  a25057a );
 a3122a <=( a25046a  and  a25035a );
 a3123a <=( a25024a  and  a25013a );
 a3124a <=( a25002a  and  a24991a );
 a3125a <=( a24980a  and  a24969a );
 a3126a <=( a24958a  and  a24947a );
 a3127a <=( a24936a  and  a24925a );
 a3128a <=( a24914a  and  a24903a );
 a3129a <=( a24892a  and  a24881a );
 a3130a <=( a24870a  and  a24859a );
 a3131a <=( a24848a  and  a24837a );
 a3132a <=( a24826a  and  a24815a );
 a3133a <=( a24804a  and  a24793a );
 a3134a <=( a24782a  and  a24771a );
 a3135a <=( a24760a  and  a24749a );
 a3136a <=( a24738a  and  a24727a );
 a3137a <=( a24716a  and  a24705a );
 a3138a <=( a24694a  and  a24683a );
 a3139a <=( a24672a  and  a24661a );
 a3140a <=( a24650a  and  a24639a );
 a3141a <=( a24628a  and  a24617a );
 a3142a <=( a24606a  and  a24595a );
 a3143a <=( a24584a  and  a24573a );
 a3144a <=( a24562a  and  a24551a );
 a3145a <=( a24540a  and  a24529a );
 a3146a <=( a24518a  and  a24507a );
 a3147a <=( a24496a  and  a24485a );
 a3148a <=( a24476a  and  a24465a );
 a3149a <=( a24456a  and  a24445a );
 a3150a <=( a24436a  and  a24425a );
 a3151a <=( a24416a  and  a24405a );
 a3152a <=( a24396a  and  a24385a );
 a3153a <=( a24376a  and  a24365a );
 a3154a <=( a24356a  and  a24345a );
 a3155a <=( a24336a  and  a24325a );
 a3156a <=( a24316a  and  a24305a );
 a3157a <=( a24296a  and  a24285a );
 a3158a <=( a24276a  and  a24265a );
 a3159a <=( a24256a  and  a24245a );
 a3160a <=( a24236a  and  a24225a );
 a3161a <=( a24216a  and  a24205a );
 a3162a <=( a24196a  and  a24185a );
 a3163a <=( a24176a  and  a24165a );
 a3164a <=( a24156a  and  a24145a );
 a3165a <=( a24136a  and  a24125a );
 a3166a <=( a24116a  and  a24105a );
 a3167a <=( a24096a  and  a24085a );
 a3168a <=( a24076a  and  a24065a );
 a3169a <=( a24056a  and  a24045a );
 a3170a <=( a24036a  and  a24025a );
 a3171a <=( a24016a  and  a24005a );
 a3172a <=( a23996a  and  a23985a );
 a3173a <=( a23976a  and  a23965a );
 a3174a <=( a23956a  and  a23945a );
 a3175a <=( a23936a  and  a23925a );
 a3176a <=( a23916a  and  a23905a );
 a3177a <=( a23896a  and  a23885a );
 a3178a <=( a23876a  and  a23865a );
 a3179a <=( a23856a  and  a23845a );
 a3180a <=( a23836a  and  a23825a );
 a3181a <=( a23816a  and  a23805a );
 a3182a <=( a23796a  and  a23785a );
 a3183a <=( a23776a  and  a23765a );
 a3184a <=( a23756a  and  a23745a );
 a3185a <=( a23736a  and  a23725a );
 a3186a <=( a23716a  and  a23705a );
 a3187a <=( a23696a  and  a23685a );
 a3188a <=( a23676a  and  a23665a );
 a3189a <=( a23656a  and  a23645a );
 a3190a <=( a23636a  and  a23625a );
 a3191a <=( a23616a  and  a23605a );
 a3192a <=( a23596a  and  a23585a );
 a3193a <=( a23576a  and  a23565a );
 a3194a <=( a23556a  and  a23545a );
 a3195a <=( a23536a  and  a23525a );
 a3196a <=( a23516a  and  a23505a );
 a3197a <=( a23496a  and  a23485a );
 a3198a <=( a23476a  and  a23465a );
 a3199a <=( a23456a  and  a23445a );
 a3200a <=( a23436a  and  a23425a );
 a3201a <=( a23416a  and  a23405a );
 a3202a <=( a23396a  and  a23385a );
 a3203a <=( a23376a  and  a23365a );
 a3204a <=( a23356a  and  a23345a );
 a3205a <=( a23336a  and  a23325a );
 a3206a <=( a23316a  and  a23305a );
 a3207a <=( a23296a  and  a23285a );
 a3208a <=( a23276a  and  a23265a );
 a3209a <=( a23256a  and  a23245a );
 a3210a <=( a23236a  and  a23225a );
 a3211a <=( a23216a  and  a23205a );
 a3212a <=( a23196a  and  a23185a );
 a3213a <=( a23176a  and  a23165a );
 a3214a <=( a23156a  and  a23145a );
 a3215a <=( a23136a  and  a23125a );
 a3216a <=( a23116a  and  a23105a );
 a3217a <=( a23096a  and  a23085a );
 a3218a <=( a23076a  and  a23065a );
 a3219a <=( a23056a  and  a23045a );
 a3220a <=( a23036a  and  a23025a );
 a3221a <=( a23016a  and  a23005a );
 a3222a <=( a22996a  and  a22985a );
 a3223a <=( a22976a  and  a22965a );
 a3224a <=( a22956a  and  a22945a );
 a3225a <=( a22936a  and  a22925a );
 a3226a <=( a22916a  and  a22905a );
 a3227a <=( a22896a  and  a22885a );
 a3228a <=( a22876a  and  a22865a );
 a3229a <=( a22856a  and  a22845a );
 a3230a <=( a22836a  and  a22825a );
 a3231a <=( a22816a  and  a22805a );
 a3232a <=( a22796a  and  a22785a );
 a3233a <=( a22776a  and  a22765a );
 a3234a <=( a22756a  and  a22745a );
 a3235a <=( a22736a  and  a22725a );
 a3236a <=( a22716a  and  a22705a );
 a3237a <=( a22696a  and  a22685a );
 a3238a <=( a22676a  and  a22665a );
 a3239a <=( a22656a  and  a22645a );
 a3240a <=( a22636a  and  a22625a );
 a3241a <=( a22616a  and  a22605a );
 a3242a <=( a22596a  and  a22585a );
 a3243a <=( a22576a  and  a22565a );
 a3244a <=( a22556a  and  a22545a );
 a3245a <=( a22536a  and  a22525a );
 a3246a <=( a22516a  and  a22505a );
 a3247a <=( a22496a  and  a22485a );
 a3248a <=( a22476a  and  a22465a );
 a3249a <=( a22456a  and  a22445a );
 a3250a <=( a22436a  and  a22425a );
 a3251a <=( a22416a  and  a22405a );
 a3252a <=( a22396a  and  a22385a );
 a3253a <=( a22376a  and  a22365a );
 a3254a <=( a22356a  and  a22345a );
 a3255a <=( a22336a  and  a22325a );
 a3256a <=( a22316a  and  a22305a );
 a3257a <=( a22296a  and  a22285a );
 a3258a <=( a22276a  and  a22265a );
 a3259a <=( a22256a  and  a22245a );
 a3260a <=( a22236a  and  a22225a );
 a3261a <=( a22216a  and  a22205a );
 a3262a <=( a22196a  and  a22185a );
 a3263a <=( a22176a  and  a22165a );
 a3264a <=( a22156a  and  a22145a );
 a3265a <=( a22136a  and  a22125a );
 a3266a <=( a22116a  and  a22105a );
 a3267a <=( a22096a  and  a22085a );
 a3268a <=( a22076a  and  a22065a );
 a3269a <=( a22056a  and  a22045a );
 a3270a <=( a22036a  and  a22025a );
 a3271a <=( a22016a  and  a22005a );
 a3272a <=( a21996a  and  a21985a );
 a3273a <=( a21976a  and  a21965a );
 a3274a <=( a21956a  and  a21945a );
 a3275a <=( a21936a  and  a21925a );
 a3276a <=( a21916a  and  a21905a );
 a3277a <=( a21896a  and  a21885a );
 a3278a <=( a21876a  and  a21865a );
 a3279a <=( a21856a  and  a21845a );
 a3280a <=( a21836a  and  a21825a );
 a3281a <=( a21816a  and  a21805a );
 a3282a <=( a21796a  and  a21785a );
 a3283a <=( a21776a  and  a21765a );
 a3284a <=( a21756a  and  a21745a );
 a3285a <=( a21736a  and  a21725a );
 a3286a <=( a21716a  and  a21705a );
 a3287a <=( a21696a  and  a21685a );
 a3288a <=( a21676a  and  a21665a );
 a3289a <=( a21656a  and  a21645a );
 a3290a <=( a21636a  and  a21625a );
 a3291a <=( a21616a  and  a21605a );
 a3292a <=( a21596a  and  a21585a );
 a3293a <=( a21576a  and  a21565a );
 a3294a <=( a21556a  and  a21545a );
 a3295a <=( a21536a  and  a21525a );
 a3296a <=( a21516a  and  a21505a );
 a3297a <=( a21496a  and  a21485a );
 a3298a <=( a21476a  and  a21465a );
 a3299a <=( a21456a  and  a21445a );
 a3300a <=( a21436a  and  a21425a );
 a3301a <=( a21416a  and  a21405a );
 a3302a <=( a21396a  and  a21385a );
 a3303a <=( a21376a  and  a21365a );
 a3304a <=( a21356a  and  a21345a );
 a3305a <=( a21336a  and  a21325a );
 a3306a <=( a21316a  and  a21305a );
 a3307a <=( a21296a  and  a21285a );
 a3308a <=( a21276a  and  a21265a );
 a3309a <=( a21256a  and  a21245a );
 a3310a <=( a21236a  and  a21225a );
 a3311a <=( a21216a  and  a21205a );
 a3312a <=( a21196a  and  a21185a );
 a3313a <=( a21176a  and  a21165a );
 a3314a <=( a21156a  and  a21145a );
 a3315a <=( a21136a  and  a21125a );
 a3316a <=( a21116a  and  a21105a );
 a3317a <=( a21096a  and  a21085a );
 a3318a <=( a21076a  and  a21065a );
 a3319a <=( a21056a  and  a21045a );
 a3320a <=( a21036a  and  a21025a );
 a3321a <=( a21016a  and  a21005a );
 a3322a <=( a20996a  and  a20985a );
 a3323a <=( a20976a  and  a20965a );
 a3324a <=( a20956a  and  a20945a );
 a3325a <=( a20936a  and  a20925a );
 a3326a <=( a20916a  and  a20905a );
 a3327a <=( a20896a  and  a20885a );
 a3328a <=( a20876a  and  a20865a );
 a3329a <=( a20856a  and  a20845a );
 a3330a <=( a20836a  and  a20825a );
 a3331a <=( a20816a  and  a20805a );
 a3332a <=( a20796a  and  a20785a );
 a3333a <=( a20776a  and  a20765a );
 a3334a <=( a20756a  and  a20745a );
 a3335a <=( a20736a  and  a20725a );
 a3336a <=( a20716a  and  a20705a );
 a3337a <=( a20696a  and  a20685a );
 a3338a <=( a20676a  and  a20665a );
 a3339a <=( a20656a  and  a20645a );
 a3340a <=( a20636a  and  a20625a );
 a3341a <=( a20616a  and  a20605a );
 a3342a <=( a20596a  and  a20585a );
 a3343a <=( a20576a  and  a20565a );
 a3344a <=( a20556a  and  a20545a );
 a3345a <=( a20536a  and  a20525a );
 a3346a <=( a20516a  and  a20505a );
 a3347a <=( a20496a  and  a20485a );
 a3348a <=( a20476a  and  a20465a );
 a3349a <=( a20456a  and  a20445a );
 a3350a <=( a20436a  and  a20425a );
 a3351a <=( a20416a  and  a20405a );
 a3352a <=( a20396a  and  a20385a );
 a3353a <=( a20376a  and  a20365a );
 a3354a <=( a20356a  and  a20345a );
 a3355a <=( a20336a  and  a20325a );
 a3356a <=( a20316a  and  a20305a );
 a3357a <=( a20296a  and  a20285a );
 a3358a <=( a20276a  and  a20265a );
 a3359a <=( a20256a  and  a20245a );
 a3360a <=( a20236a  and  a20225a );
 a3361a <=( a20216a  and  a20205a );
 a3362a <=( a20196a  and  a20185a );
 a3363a <=( a20176a  and  a20165a );
 a3364a <=( a20156a  and  a20145a );
 a3365a <=( a20136a  and  a20125a );
 a3366a <=( a20116a  and  a20105a );
 a3367a <=( a20096a  and  a20085a );
 a3368a <=( a20076a  and  a20065a );
 a3369a <=( a20056a  and  a20045a );
 a3370a <=( a20036a  and  a20025a );
 a3371a <=( a20016a  and  a20005a );
 a3372a <=( a19996a  and  a19985a );
 a3373a <=( a19976a  and  a19965a );
 a3374a <=( a19956a  and  a19945a );
 a3375a <=( a19936a  and  a19925a );
 a3376a <=( a19916a  and  a19905a );
 a3377a <=( a19896a  and  a19885a );
 a3378a <=( a19876a  and  a19865a );
 a3379a <=( a19856a  and  a19845a );
 a3380a <=( a19836a  and  a19825a );
 a3381a <=( a19816a  and  a19805a );
 a3382a <=( a19796a  and  a19785a );
 a3383a <=( a19776a  and  a19765a );
 a3384a <=( a19756a  and  a19745a );
 a3385a <=( a19736a  and  a19725a );
 a3386a <=( a19716a  and  a19705a );
 a3387a <=( a19696a  and  a19685a );
 a3388a <=( a19676a  and  a19665a );
 a3389a <=( a19656a  and  a19645a );
 a3390a <=( a19636a  and  a19625a );
 a3391a <=( a19616a  and  a19605a );
 a3392a <=( a19596a  and  a19585a );
 a3393a <=( a19576a  and  a19565a );
 a3394a <=( a19556a  and  a19545a );
 a3395a <=( a19536a  and  a19525a );
 a3396a <=( a19516a  and  a19505a );
 a3397a <=( a19496a  and  a19485a );
 a3398a <=( a19476a  and  a19465a );
 a3399a <=( a19456a  and  a19445a );
 a3400a <=( a19436a  and  a19425a );
 a3401a <=( a19416a  and  a19405a );
 a3402a <=( a19396a  and  a19385a );
 a3403a <=( a19376a  and  a19365a );
 a3404a <=( a19356a  and  a19345a );
 a3405a <=( a19336a  and  a19325a );
 a3406a <=( a19316a  and  a19305a );
 a3407a <=( a19296a  and  a19285a );
 a3408a <=( a19276a  and  a19265a );
 a3409a <=( a19256a  and  a19245a );
 a3410a <=( a19236a  and  a19225a );
 a3411a <=( a19216a  and  a19205a );
 a3412a <=( a19196a  and  a19185a );
 a3413a <=( a19176a  and  a19165a );
 a3414a <=( a19156a  and  a19145a );
 a3415a <=( a19136a  and  a19125a );
 a3416a <=( a19116a  and  a19105a );
 a3417a <=( a19096a  and  a19085a );
 a3418a <=( a19076a  and  a19065a );
 a3419a <=( a19056a  and  a19045a );
 a3420a <=( a19036a  and  a19025a );
 a3421a <=( a19016a  and  a19005a );
 a3422a <=( a18996a  and  a18985a );
 a3423a <=( a18976a  and  a18965a );
 a3424a <=( a18956a  and  a18945a );
 a3425a <=( a18936a  and  a18925a );
 a3426a <=( a18916a  and  a18905a );
 a3427a <=( a18896a  and  a18885a );
 a3428a <=( a18876a  and  a18865a );
 a3429a <=( a18856a  and  a18845a );
 a3430a <=( a18836a  and  a18825a );
 a3431a <=( a18816a  and  a18805a );
 a3432a <=( a18796a  and  a18785a );
 a3433a <=( a18776a  and  a18765a );
 a3434a <=( a18756a  and  a18745a );
 a3435a <=( a18736a  and  a18725a );
 a3436a <=( a18716a  and  a18705a );
 a3437a <=( a18696a  and  a18685a );
 a3438a <=( a18676a  and  a18665a );
 a3439a <=( a18656a  and  a18645a );
 a3440a <=( a18636a  and  a18625a );
 a3441a <=( a18616a  and  a18605a );
 a3442a <=( a18596a  and  a18585a );
 a3443a <=( a18576a  and  a18565a );
 a3444a <=( a18556a  and  a18545a );
 a3445a <=( a18536a  and  a18525a );
 a3446a <=( a18516a  and  a18505a );
 a3447a <=( a18496a  and  a18485a );
 a3448a <=( a18476a  and  a18465a );
 a3449a <=( a18456a  and  a18445a );
 a3450a <=( a18436a  and  a18425a );
 a3451a <=( a18416a  and  a18405a );
 a3452a <=( a18396a  and  a18385a );
 a3453a <=( a18376a  and  a18365a );
 a3454a <=( a18356a  and  a18345a );
 a3455a <=( a18336a  and  a18325a );
 a3456a <=( a18316a  and  a18305a );
 a3457a <=( a18296a  and  a18285a );
 a3458a <=( a18276a  and  a18265a );
 a3459a <=( a18256a  and  a18245a );
 a3460a <=( a18236a  and  a18225a );
 a3461a <=( a18216a  and  a18205a );
 a3462a <=( a18196a  and  a18185a );
 a3463a <=( a18176a  and  a18165a );
 a3464a <=( a18156a  and  a18145a );
 a3465a <=( a18136a  and  a18125a );
 a3466a <=( a18116a  and  a18105a );
 a3467a <=( a18096a  and  a18085a );
 a3468a <=( a18076a  and  a18065a );
 a3469a <=( a18056a  and  a18045a );
 a3470a <=( a18036a  and  a18025a );
 a3471a <=( a18016a  and  a18005a );
 a3472a <=( a17996a  and  a17985a );
 a3473a <=( a17976a  and  a17965a );
 a3474a <=( a17956a  and  a17945a );
 a3475a <=( a17936a  and  a17925a );
 a3476a <=( a17916a  and  a17905a );
 a3477a <=( a17896a  and  a17885a );
 a3478a <=( a17876a  and  a17865a );
 a3479a <=( a17856a  and  a17845a );
 a3480a <=( a17836a  and  a17825a );
 a3481a <=( a17816a  and  a17805a );
 a3482a <=( a17796a  and  a17785a );
 a3483a <=( a17776a  and  a17765a );
 a3484a <=( a17756a  and  a17745a );
 a3485a <=( a17736a  and  a17725a );
 a3486a <=( a17716a  and  a17705a );
 a3487a <=( a17696a  and  a17685a );
 a3488a <=( a17676a  and  a17665a );
 a3489a <=( a17656a  and  a17645a );
 a3490a <=( a17636a  and  a17625a );
 a3491a <=( a17616a  and  a17605a );
 a3492a <=( a17596a  and  a17585a );
 a3493a <=( a17576a  and  a17565a );
 a3494a <=( a17556a  and  a17545a );
 a3495a <=( a17536a  and  a17525a );
 a3496a <=( a17516a  and  a17505a );
 a3497a <=( a17496a  and  a17485a );
 a3498a <=( a17476a  and  a17465a );
 a3499a <=( a17456a  and  a17447a );
 a3500a <=( a17438a  and  a17429a );
 a3501a <=( a17420a  and  a17411a );
 a3502a <=( a17402a  and  a17393a );
 a3503a <=( a17384a  and  a17375a );
 a3504a <=( a17366a  and  a17357a );
 a3505a <=( a17348a  and  a17339a );
 a3506a <=( a17330a  and  a17321a );
 a3507a <=( a17312a  and  a17303a );
 a3508a <=( a17294a  and  a17285a );
 a3509a <=( a17276a  and  a17267a );
 a3510a <=( a17258a  and  a17249a );
 a3511a <=( a17240a  and  a17231a );
 a3512a <=( a17222a  and  a17213a );
 a3513a <=( a17204a  and  a17195a );
 a3514a <=( a17186a  and  a17177a );
 a3515a <=( a17168a  and  a17159a );
 a3516a <=( a17150a  and  a17141a );
 a3517a <=( a17132a  and  a17123a );
 a3518a <=( a17114a  and  a17105a );
 a3519a <=( a17096a  and  a17087a );
 a3520a <=( a17078a  and  a17069a );
 a3521a <=( a17060a  and  a17051a );
 a3522a <=( a17042a  and  a17033a );
 a3523a <=( a17024a  and  a17015a );
 a3524a <=( a17006a  and  a16997a );
 a3525a <=( a16988a  and  a16979a );
 a3526a <=( a16970a  and  a16961a );
 a3527a <=( a16952a  and  a16943a );
 a3528a <=( a16934a  and  a16925a );
 a3529a <=( a16916a  and  a16907a );
 a3530a <=( a16898a  and  a16889a );
 a3531a <=( a16880a  and  a16871a );
 a3532a <=( a16862a  and  a16853a );
 a3533a <=( a16844a  and  a16835a );
 a3534a <=( a16826a  and  a16817a );
 a3535a <=( a16808a  and  a16799a );
 a3536a <=( a16790a  and  a16781a );
 a3537a <=( a16772a  and  a16763a );
 a3538a <=( a16754a  and  a16745a );
 a3539a <=( a16736a  and  a16727a );
 a3540a <=( a16718a  and  a16709a );
 a3541a <=( a16700a  and  a16691a );
 a3542a <=( a16682a  and  a16673a );
 a3543a <=( a16664a  and  a16655a );
 a3544a <=( a16646a  and  a16637a );
 a3545a <=( a16628a  and  a16619a );
 a3546a <=( a16610a  and  a16601a );
 a3547a <=( a16592a  and  a16583a );
 a3548a <=( a16574a  and  a16565a );
 a3549a <=( a16556a  and  a16547a );
 a3550a <=( a16538a  and  a16529a );
 a3551a <=( a16520a  and  a16511a );
 a3552a <=( a16502a  and  a16493a );
 a3553a <=( a16484a  and  a16475a );
 a3554a <=( a16466a  and  a16457a );
 a3555a <=( a16448a  and  a16439a );
 a3556a <=( a16430a  and  a16421a );
 a3557a <=( a16412a  and  a16403a );
 a3558a <=( a16394a  and  a16385a );
 a3559a <=( a16376a  and  a16367a );
 a3560a <=( a16358a  and  a16349a );
 a3561a <=( a16340a  and  a16331a );
 a3562a <=( a16322a  and  a16313a );
 a3563a <=( a16304a  and  a16295a );
 a3564a <=( a16286a  and  a16277a );
 a3565a <=( a16268a  and  a16259a );
 a3566a <=( a16250a  and  a16241a );
 a3567a <=( a16232a  and  a16223a );
 a3568a <=( a16214a  and  a16205a );
 a3569a <=( a16196a  and  a16187a );
 a3570a <=( a16178a  and  a16169a );
 a3571a <=( a16160a  and  a16151a );
 a3572a <=( a16142a  and  a16133a );
 a3573a <=( a16124a  and  a16115a );
 a3574a <=( a16106a  and  a16097a );
 a3575a <=( a16088a  and  a16079a );
 a3576a <=( a16070a  and  a16061a );
 a3577a <=( a16052a  and  a16043a );
 a3578a <=( a16034a  and  a16025a );
 a3579a <=( a16016a  and  a16007a );
 a3580a <=( a15998a  and  a15989a );
 a3581a <=( a15980a  and  a15971a );
 a3582a <=( a15962a  and  a15953a );
 a3583a <=( a15944a  and  a15935a );
 a3584a <=( a15926a  and  a15917a );
 a3585a <=( a15908a  and  a15899a );
 a3586a <=( a15890a  and  a15881a );
 a3587a <=( a15872a  and  a15863a );
 a3588a <=( a15854a  and  a15845a );
 a3589a <=( a15836a  and  a15827a );
 a3590a <=( a15818a  and  a15809a );
 a3591a <=( a15800a  and  a15791a );
 a3592a <=( a15782a  and  a15773a );
 a3593a <=( a15764a  and  a15755a );
 a3594a <=( a15746a  and  a15737a );
 a3595a <=( a15728a  and  a15719a );
 a3596a <=( a15710a  and  a15701a );
 a3597a <=( a15692a  and  a15683a );
 a3598a <=( a15674a  and  a15665a );
 a3599a <=( a15656a  and  a15647a );
 a3600a <=( a15638a  and  a15629a );
 a3601a <=( a15620a  and  a15611a );
 a3602a <=( a15602a  and  a15593a );
 a3603a <=( a15584a  and  a15575a );
 a3604a <=( a15566a  and  a15557a );
 a3605a <=( a15548a  and  a15539a );
 a3606a <=( a15530a  and  a15521a );
 a3607a <=( a15512a  and  a15503a );
 a3608a <=( a15494a  and  a15485a );
 a3609a <=( a15476a  and  a15467a );
 a3610a <=( a15458a  and  a15449a );
 a3611a <=( a15440a  and  a15431a );
 a3612a <=( a15422a  and  a15413a );
 a3613a <=( a15404a  and  a15395a );
 a3614a <=( a15386a  and  a15377a );
 a3615a <=( a15368a  and  a15359a );
 a3616a <=( a15350a  and  a15341a );
 a3617a <=( a15332a  and  a15323a );
 a3618a <=( a15314a  and  a15305a );
 a3619a <=( a15296a  and  a15287a );
 a3620a <=( a15278a  and  a15269a );
 a3621a <=( a15260a  and  a15251a );
 a3622a <=( a15242a  and  a15233a );
 a3623a <=( a15224a  and  a15215a );
 a3624a <=( a15206a  and  a15197a );
 a3625a <=( a15188a  and  a15179a );
 a3626a <=( a15170a  and  a15161a );
 a3627a <=( a15152a  and  a15143a );
 a3628a <=( a15134a  and  a15125a );
 a3629a <=( a15116a  and  a15107a );
 a3630a <=( a15098a  and  a15089a );
 a3631a <=( a15080a  and  a15071a );
 a3632a <=( a15062a  and  a15053a );
 a3633a <=( a15044a  and  a15035a );
 a3634a <=( a15026a  and  a15017a );
 a3635a <=( a15008a  and  a14999a );
 a3636a <=( a14990a  and  a14981a );
 a3637a <=( a14972a  and  a14963a );
 a3638a <=( a14954a  and  a14945a );
 a3639a <=( a14936a  and  a14927a );
 a3640a <=( a14918a  and  a14909a );
 a3641a <=( a14900a  and  a14891a );
 a3642a <=( a14882a  and  a14873a );
 a3643a <=( a14864a  and  a14855a );
 a3644a <=( a14846a  and  a14837a );
 a3645a <=( a14828a  and  a14819a );
 a3646a <=( a14810a  and  a14801a );
 a3647a <=( a14792a  and  a14783a );
 a3648a <=( a14774a  and  a14765a );
 a3649a <=( a14756a  and  a14747a );
 a3650a <=( a14738a  and  a14729a );
 a3651a <=( a14720a  and  a14711a );
 a3652a <=( a14702a  and  a14693a );
 a3653a <=( a14684a  and  a14675a );
 a3654a <=( a14666a  and  a14657a );
 a3655a <=( a14648a  and  a14639a );
 a3656a <=( a14630a  and  a14621a );
 a3657a <=( a14612a  and  a14603a );
 a3658a <=( a14594a  and  a14585a );
 a3659a <=( a14576a  and  a14567a );
 a3660a <=( a14558a  and  a14549a );
 a3661a <=( a14540a  and  a14531a );
 a3662a <=( a14522a  and  a14513a );
 a3663a <=( a14504a  and  a14495a );
 a3664a <=( a14486a  and  a14477a );
 a3665a <=( a14468a  and  a14459a );
 a3666a <=( a14450a  and  a14441a );
 a3667a <=( a14432a  and  a14423a );
 a3668a <=( a14414a  and  a14405a );
 a3669a <=( a14396a  and  a14387a );
 a3670a <=( a14378a  and  a14369a );
 a3671a <=( a14360a  and  a14351a );
 a3672a <=( a14342a  and  a14333a );
 a3673a <=( a14324a  and  a14315a );
 a3674a <=( a14306a  and  a14297a );
 a3675a <=( a14288a  and  a14279a );
 a3676a <=( a14270a  and  a14261a );
 a3677a <=( a14252a  and  a14243a );
 a3678a <=( a14234a  and  a14225a );
 a3679a <=( a14216a  and  a14207a );
 a3680a <=( a14198a  and  a14189a );
 a3681a <=( a14180a  and  a14171a );
 a3682a <=( a14162a  and  a14153a );
 a3683a <=( a14144a  and  a14135a );
 a3684a <=( a14126a  and  a14117a );
 a3685a <=( a14108a  and  a14099a );
 a3686a <=( a14090a  and  a14081a );
 a3687a <=( a14072a  and  a14063a );
 a3688a <=( a14054a  and  a14045a );
 a3689a <=( a14036a  and  a14027a );
 a3690a <=( a14018a  and  a14009a );
 a3691a <=( a14000a  and  a13991a );
 a3692a <=( a13982a  and  a13973a );
 a3693a <=( a13964a  and  a13955a );
 a3694a <=( a13946a  and  a13937a );
 a3695a <=( a13928a  and  a13919a );
 a3696a <=( a13910a  and  a13901a );
 a3697a <=( a13892a  and  a13883a );
 a3698a <=( a13874a  and  a13865a );
 a3699a <=( a13856a  and  a13847a );
 a3700a <=( a13838a  and  a13829a );
 a3701a <=( a13820a  and  a13811a );
 a3702a <=( a13802a  and  a13793a );
 a3703a <=( a13784a  and  a13775a );
 a3704a <=( a13766a  and  a13757a );
 a3705a <=( a13748a  and  a13739a );
 a3706a <=( a13730a  and  a13721a );
 a3707a <=( a13712a  and  a13703a );
 a3708a <=( a13694a  and  a13685a );
 a3709a <=( a13676a  and  a13667a );
 a3710a <=( a13658a  and  a13649a );
 a3711a <=( a13640a  and  a13631a );
 a3712a <=( a13622a  and  a13613a );
 a3713a <=( a13604a  and  a13595a );
 a3714a <=( a13586a  and  a13577a );
 a3715a <=( a13568a  and  a13559a );
 a3716a <=( a13550a  and  a13541a );
 a3717a <=( a13532a  and  a13523a );
 a3718a <=( a13514a  and  a13505a );
 a3719a <=( a13496a  and  a13487a );
 a3720a <=( a13478a  and  a13469a );
 a3721a <=( a13460a  and  a13451a );
 a3722a <=( a13442a  and  a13433a );
 a3723a <=( a13424a  and  a13415a );
 a3724a <=( a13406a  and  a13397a );
 a3725a <=( a13388a  and  a13379a );
 a3726a <=( a13370a  and  a13361a );
 a3727a <=( a13352a  and  a13343a );
 a3728a <=( a13334a  and  a13325a );
 a3729a <=( a13316a  and  a13307a );
 a3730a <=( a13298a  and  a13289a );
 a3731a <=( a13280a  and  a13271a );
 a3732a <=( a13262a  and  a13253a );
 a3733a <=( a13244a  and  a13235a );
 a3734a <=( a13226a  and  a13217a );
 a3735a <=( a13208a  and  a13199a );
 a3736a <=( a13190a  and  a13181a );
 a3737a <=( a13172a  and  a13163a );
 a3738a <=( a13154a  and  a13145a );
 a3739a <=( a13136a  and  a13127a );
 a3740a <=( a13118a  and  a13109a );
 a3741a <=( a13100a  and  a13091a );
 a3742a <=( a13082a  and  a13073a );
 a3743a <=( a13064a  and  a13055a );
 a3744a <=( a13046a  and  a13037a );
 a3745a <=( a13028a  and  a13019a );
 a3746a <=( a13010a  and  a13001a );
 a3747a <=( a12992a  and  a12983a );
 a3748a <=( a12974a  and  a12965a );
 a3749a <=( a12956a  and  a12947a );
 a3750a <=( a12938a  and  a12929a );
 a3751a <=( a12920a  and  a12911a );
 a3752a <=( a12902a  and  a12893a );
 a3753a <=( a12884a  and  a12875a );
 a3754a <=( a12866a  and  a12857a );
 a3755a <=( a12848a  and  a12839a );
 a3756a <=( a12830a  and  a12821a );
 a3757a <=( a12812a  and  a12803a );
 a3758a <=( a12794a  and  a12785a );
 a3759a <=( a12776a  and  a12767a );
 a3760a <=( a12758a  and  a12749a );
 a3761a <=( a12740a  and  a12731a );
 a3762a <=( a12722a  and  a12713a );
 a3763a <=( a12704a  and  a12695a );
 a3764a <=( a12686a  and  a12677a );
 a3765a <=( a12668a  and  a12659a );
 a3766a <=( a12650a  and  a12641a );
 a3767a <=( a12632a  and  a12623a );
 a3768a <=( a12614a  and  a12605a );
 a3769a <=( a12596a  and  a12587a );
 a3770a <=( a12578a  and  a12569a );
 a3771a <=( a12560a  and  a12551a );
 a3772a <=( a12542a  and  a12533a );
 a3773a <=( a12524a  and  a12515a );
 a3774a <=( a12506a  and  a12497a );
 a3775a <=( a12488a  and  a12479a );
 a3776a <=( a12470a  and  a12461a );
 a3777a <=( a12452a  and  a12443a );
 a3778a <=( a12434a  and  a12425a );
 a3779a <=( a12416a  and  a12407a );
 a3780a <=( a12398a  and  a12389a );
 a3781a <=( a12380a  and  a12371a );
 a3782a <=( a12362a  and  a12353a );
 a3783a <=( a12344a  and  a12335a );
 a3784a <=( a12328a  and  a12319a );
 a3785a <=( a12312a  and  a12303a );
 a3786a <=( a12296a  and  a12287a );
 a3787a <=( a12280a  and  a12271a );
 a3788a <=( a12264a  and  a12255a );
 a3789a <=( a12248a  and  a12239a );
 a3790a <=( a12232a  and  a12223a );
 a3791a <=( a12216a  and  a12207a );
 a3792a <=( a12200a  and  a12191a );
 a3793a <=( a12184a  and  a12175a );
 a3794a <=( a12168a  and  a12159a );
 a3795a <=( a12152a  and  a12143a );
 a3796a <=( a12136a  and  a12127a );
 a3797a <=( a12120a  and  a12111a );
 a3798a <=( a12104a  and  a12095a );
 a3799a <=( a12088a  and  a12079a );
 a3800a <=( a12072a  and  a12063a );
 a3801a <=( a12056a  and  a12047a );
 a3802a <=( a12040a  and  a12031a );
 a3803a <=( a12024a  and  a12015a );
 a3804a <=( a12008a  and  a11999a );
 a3805a <=( a11992a  and  a11983a );
 a3806a <=( a11976a  and  a11967a );
 a3807a <=( a11960a  and  a11953a );
 a3808a <=( a11946a  and  a11939a );
 a3809a <=( a11932a  and  a11925a );
 a3810a <=( a11918a  and  a11911a );
 a3811a <=( a11904a  and  a11897a );
 a3812a <=( a11890a  and  a11883a );
 a3813a <=( a11876a  and  a11869a );
 a3814a <=( a11862a  and  a11855a );
 a3815a <=( a11848a  and  a11841a );
 a3816a <=( a11834a  and  a11827a );
 a3817a <=( a11820a  and  a11813a );
 a3818a <=( a11806a  and  a11799a );
 a3819a <=( a11792a  and  a11785a );
 a3820a <=( a11778a  and  a11771a );
 a3821a <=( a11764a  and  a11757a );
 a3822a <=( a11750a  and  a11743a );
 a3823a <=( a11736a  and  a11729a );
 a3824a <=( a11722a  and  a11715a );
 a3825a <=( a11708a  and  a11701a );
 a3826a <=( a11694a  and  a11687a );
 a3827a <=( a11680a  and  a11673a );
 a3828a <=( a11666a  and  a11659a );
 a3829a <=( a11652a  and  a11645a );
 a3830a <=( a11638a  and  a11631a );
 a3831a <=( a11624a  and  a11617a );
 a3832a <=( a11610a  and  a11603a );
 a3833a <=( a11596a  and  a11589a );
 a3834a <=( a11582a  and  a11575a );
 a3835a <=( a11568a  and  a11561a );
 a3836a <=( a11554a  and  a11547a );
 a3837a <=( a11540a  and  a11533a );
 a3838a <=( a11526a  and  a11519a );
 a3842a <=( a3836a ) or ( a3837a );
 a3843a <=( a3838a ) or ( a3842a );
 a3846a <=( a3834a ) or ( a3835a );
 a3849a <=( a3832a ) or ( a3833a );
 a3850a <=( a3849a ) or ( a3846a );
 a3851a <=( a3850a ) or ( a3843a );
 a3855a <=( a3829a ) or ( a3830a );
 a3856a <=( a3831a ) or ( a3855a );
 a3859a <=( a3827a ) or ( a3828a );
 a3862a <=( a3825a ) or ( a3826a );
 a3863a <=( a3862a ) or ( a3859a );
 a3864a <=( a3863a ) or ( a3856a );
 a3865a <=( a3864a ) or ( a3851a );
 a3869a <=( a3822a ) or ( a3823a );
 a3870a <=( a3824a ) or ( a3869a );
 a3873a <=( a3820a ) or ( a3821a );
 a3876a <=( a3818a ) or ( a3819a );
 a3877a <=( a3876a ) or ( a3873a );
 a3878a <=( a3877a ) or ( a3870a );
 a3881a <=( a3816a ) or ( a3817a );
 a3884a <=( a3814a ) or ( a3815a );
 a3885a <=( a3884a ) or ( a3881a );
 a3888a <=( a3812a ) or ( a3813a );
 a3891a <=( a3810a ) or ( a3811a );
 a3892a <=( a3891a ) or ( a3888a );
 a3893a <=( a3892a ) or ( a3885a );
 a3894a <=( a3893a ) or ( a3878a );
 a3895a <=( a3894a ) or ( a3865a );
 a3899a <=( a3807a ) or ( a3808a );
 a3900a <=( a3809a ) or ( a3899a );
 a3903a <=( a3805a ) or ( a3806a );
 a3906a <=( a3803a ) or ( a3804a );
 a3907a <=( a3906a ) or ( a3903a );
 a3908a <=( a3907a ) or ( a3900a );
 a3911a <=( a3801a ) or ( a3802a );
 a3914a <=( a3799a ) or ( a3800a );
 a3915a <=( a3914a ) or ( a3911a );
 a3918a <=( a3797a ) or ( a3798a );
 a3921a <=( a3795a ) or ( a3796a );
 a3922a <=( a3921a ) or ( a3918a );
 a3923a <=( a3922a ) or ( a3915a );
 a3924a <=( a3923a ) or ( a3908a );
 a3928a <=( a3792a ) or ( a3793a );
 a3929a <=( a3794a ) or ( a3928a );
 a3932a <=( a3790a ) or ( a3791a );
 a3935a <=( a3788a ) or ( a3789a );
 a3936a <=( a3935a ) or ( a3932a );
 a3937a <=( a3936a ) or ( a3929a );
 a3940a <=( a3786a ) or ( a3787a );
 a3943a <=( a3784a ) or ( a3785a );
 a3944a <=( a3943a ) or ( a3940a );
 a3947a <=( a3782a ) or ( a3783a );
 a3950a <=( a3780a ) or ( a3781a );
 a3951a <=( a3950a ) or ( a3947a );
 a3952a <=( a3951a ) or ( a3944a );
 a3953a <=( a3952a ) or ( a3937a );
 a3954a <=( a3953a ) or ( a3924a );
 a3955a <=( a3954a ) or ( a3895a );
 a3959a <=( a3777a ) or ( a3778a );
 a3960a <=( a3779a ) or ( a3959a );
 a3963a <=( a3775a ) or ( a3776a );
 a3966a <=( a3773a ) or ( a3774a );
 a3967a <=( a3966a ) or ( a3963a );
 a3968a <=( a3967a ) or ( a3960a );
 a3971a <=( a3771a ) or ( a3772a );
 a3974a <=( a3769a ) or ( a3770a );
 a3975a <=( a3974a ) or ( a3971a );
 a3978a <=( a3767a ) or ( a3768a );
 a3981a <=( a3765a ) or ( a3766a );
 a3982a <=( a3981a ) or ( a3978a );
 a3983a <=( a3982a ) or ( a3975a );
 a3984a <=( a3983a ) or ( a3968a );
 a3988a <=( a3762a ) or ( a3763a );
 a3989a <=( a3764a ) or ( a3988a );
 a3992a <=( a3760a ) or ( a3761a );
 a3995a <=( a3758a ) or ( a3759a );
 a3996a <=( a3995a ) or ( a3992a );
 a3997a <=( a3996a ) or ( a3989a );
 a4000a <=( a3756a ) or ( a3757a );
 a4003a <=( a3754a ) or ( a3755a );
 a4004a <=( a4003a ) or ( a4000a );
 a4007a <=( a3752a ) or ( a3753a );
 a4010a <=( a3750a ) or ( a3751a );
 a4011a <=( a4010a ) or ( a4007a );
 a4012a <=( a4011a ) or ( a4004a );
 a4013a <=( a4012a ) or ( a3997a );
 a4014a <=( a4013a ) or ( a3984a );
 a4018a <=( a3747a ) or ( a3748a );
 a4019a <=( a3749a ) or ( a4018a );
 a4022a <=( a3745a ) or ( a3746a );
 a4025a <=( a3743a ) or ( a3744a );
 a4026a <=( a4025a ) or ( a4022a );
 a4027a <=( a4026a ) or ( a4019a );
 a4030a <=( a3741a ) or ( a3742a );
 a4033a <=( a3739a ) or ( a3740a );
 a4034a <=( a4033a ) or ( a4030a );
 a4037a <=( a3737a ) or ( a3738a );
 a4040a <=( a3735a ) or ( a3736a );
 a4041a <=( a4040a ) or ( a4037a );
 a4042a <=( a4041a ) or ( a4034a );
 a4043a <=( a4042a ) or ( a4027a );
 a4047a <=( a3732a ) or ( a3733a );
 a4048a <=( a3734a ) or ( a4047a );
 a4051a <=( a3730a ) or ( a3731a );
 a4054a <=( a3728a ) or ( a3729a );
 a4055a <=( a4054a ) or ( a4051a );
 a4056a <=( a4055a ) or ( a4048a );
 a4059a <=( a3726a ) or ( a3727a );
 a4062a <=( a3724a ) or ( a3725a );
 a4063a <=( a4062a ) or ( a4059a );
 a4066a <=( a3722a ) or ( a3723a );
 a4069a <=( a3720a ) or ( a3721a );
 a4070a <=( a4069a ) or ( a4066a );
 a4071a <=( a4070a ) or ( a4063a );
 a4072a <=( a4071a ) or ( a4056a );
 a4073a <=( a4072a ) or ( a4043a );
 a4074a <=( a4073a ) or ( a4014a );
 a4075a <=( a4074a ) or ( a3955a );
 a4079a <=( a3717a ) or ( a3718a );
 a4080a <=( a3719a ) or ( a4079a );
 a4083a <=( a3715a ) or ( a3716a );
 a4086a <=( a3713a ) or ( a3714a );
 a4087a <=( a4086a ) or ( a4083a );
 a4088a <=( a4087a ) or ( a4080a );
 a4091a <=( a3711a ) or ( a3712a );
 a4094a <=( a3709a ) or ( a3710a );
 a4095a <=( a4094a ) or ( a4091a );
 a4098a <=( a3707a ) or ( a3708a );
 a4101a <=( a3705a ) or ( a3706a );
 a4102a <=( a4101a ) or ( a4098a );
 a4103a <=( a4102a ) or ( a4095a );
 a4104a <=( a4103a ) or ( a4088a );
 a4108a <=( a3702a ) or ( a3703a );
 a4109a <=( a3704a ) or ( a4108a );
 a4112a <=( a3700a ) or ( a3701a );
 a4115a <=( a3698a ) or ( a3699a );
 a4116a <=( a4115a ) or ( a4112a );
 a4117a <=( a4116a ) or ( a4109a );
 a4120a <=( a3696a ) or ( a3697a );
 a4123a <=( a3694a ) or ( a3695a );
 a4124a <=( a4123a ) or ( a4120a );
 a4127a <=( a3692a ) or ( a3693a );
 a4130a <=( a3690a ) or ( a3691a );
 a4131a <=( a4130a ) or ( a4127a );
 a4132a <=( a4131a ) or ( a4124a );
 a4133a <=( a4132a ) or ( a4117a );
 a4134a <=( a4133a ) or ( a4104a );
 a4138a <=( a3687a ) or ( a3688a );
 a4139a <=( a3689a ) or ( a4138a );
 a4142a <=( a3685a ) or ( a3686a );
 a4145a <=( a3683a ) or ( a3684a );
 a4146a <=( a4145a ) or ( a4142a );
 a4147a <=( a4146a ) or ( a4139a );
 a4150a <=( a3681a ) or ( a3682a );
 a4153a <=( a3679a ) or ( a3680a );
 a4154a <=( a4153a ) or ( a4150a );
 a4157a <=( a3677a ) or ( a3678a );
 a4160a <=( a3675a ) or ( a3676a );
 a4161a <=( a4160a ) or ( a4157a );
 a4162a <=( a4161a ) or ( a4154a );
 a4163a <=( a4162a ) or ( a4147a );
 a4167a <=( a3672a ) or ( a3673a );
 a4168a <=( a3674a ) or ( a4167a );
 a4171a <=( a3670a ) or ( a3671a );
 a4174a <=( a3668a ) or ( a3669a );
 a4175a <=( a4174a ) or ( a4171a );
 a4176a <=( a4175a ) or ( a4168a );
 a4179a <=( a3666a ) or ( a3667a );
 a4182a <=( a3664a ) or ( a3665a );
 a4183a <=( a4182a ) or ( a4179a );
 a4186a <=( a3662a ) or ( a3663a );
 a4189a <=( a3660a ) or ( a3661a );
 a4190a <=( a4189a ) or ( a4186a );
 a4191a <=( a4190a ) or ( a4183a );
 a4192a <=( a4191a ) or ( a4176a );
 a4193a <=( a4192a ) or ( a4163a );
 a4194a <=( a4193a ) or ( a4134a );
 a4198a <=( a3657a ) or ( a3658a );
 a4199a <=( a3659a ) or ( a4198a );
 a4202a <=( a3655a ) or ( a3656a );
 a4205a <=( a3653a ) or ( a3654a );
 a4206a <=( a4205a ) or ( a4202a );
 a4207a <=( a4206a ) or ( a4199a );
 a4210a <=( a3651a ) or ( a3652a );
 a4213a <=( a3649a ) or ( a3650a );
 a4214a <=( a4213a ) or ( a4210a );
 a4217a <=( a3647a ) or ( a3648a );
 a4220a <=( a3645a ) or ( a3646a );
 a4221a <=( a4220a ) or ( a4217a );
 a4222a <=( a4221a ) or ( a4214a );
 a4223a <=( a4222a ) or ( a4207a );
 a4227a <=( a3642a ) or ( a3643a );
 a4228a <=( a3644a ) or ( a4227a );
 a4231a <=( a3640a ) or ( a3641a );
 a4234a <=( a3638a ) or ( a3639a );
 a4235a <=( a4234a ) or ( a4231a );
 a4236a <=( a4235a ) or ( a4228a );
 a4239a <=( a3636a ) or ( a3637a );
 a4242a <=( a3634a ) or ( a3635a );
 a4243a <=( a4242a ) or ( a4239a );
 a4246a <=( a3632a ) or ( a3633a );
 a4249a <=( a3630a ) or ( a3631a );
 a4250a <=( a4249a ) or ( a4246a );
 a4251a <=( a4250a ) or ( a4243a );
 a4252a <=( a4251a ) or ( a4236a );
 a4253a <=( a4252a ) or ( a4223a );
 a4257a <=( a3627a ) or ( a3628a );
 a4258a <=( a3629a ) or ( a4257a );
 a4261a <=( a3625a ) or ( a3626a );
 a4264a <=( a3623a ) or ( a3624a );
 a4265a <=( a4264a ) or ( a4261a );
 a4266a <=( a4265a ) or ( a4258a );
 a4269a <=( a3621a ) or ( a3622a );
 a4272a <=( a3619a ) or ( a3620a );
 a4273a <=( a4272a ) or ( a4269a );
 a4276a <=( a3617a ) or ( a3618a );
 a4279a <=( a3615a ) or ( a3616a );
 a4280a <=( a4279a ) or ( a4276a );
 a4281a <=( a4280a ) or ( a4273a );
 a4282a <=( a4281a ) or ( a4266a );
 a4286a <=( a3612a ) or ( a3613a );
 a4287a <=( a3614a ) or ( a4286a );
 a4290a <=( a3610a ) or ( a3611a );
 a4293a <=( a3608a ) or ( a3609a );
 a4294a <=( a4293a ) or ( a4290a );
 a4295a <=( a4294a ) or ( a4287a );
 a4298a <=( a3606a ) or ( a3607a );
 a4301a <=( a3604a ) or ( a3605a );
 a4302a <=( a4301a ) or ( a4298a );
 a4305a <=( a3602a ) or ( a3603a );
 a4308a <=( a3600a ) or ( a3601a );
 a4309a <=( a4308a ) or ( a4305a );
 a4310a <=( a4309a ) or ( a4302a );
 a4311a <=( a4310a ) or ( a4295a );
 a4312a <=( a4311a ) or ( a4282a );
 a4313a <=( a4312a ) or ( a4253a );
 a4314a <=( a4313a ) or ( a4194a );
 a4315a <=( a4314a ) or ( a4075a );
 a4319a <=( a3597a ) or ( a3598a );
 a4320a <=( a3599a ) or ( a4319a );
 a4323a <=( a3595a ) or ( a3596a );
 a4326a <=( a3593a ) or ( a3594a );
 a4327a <=( a4326a ) or ( a4323a );
 a4328a <=( a4327a ) or ( a4320a );
 a4331a <=( a3591a ) or ( a3592a );
 a4334a <=( a3589a ) or ( a3590a );
 a4335a <=( a4334a ) or ( a4331a );
 a4338a <=( a3587a ) or ( a3588a );
 a4341a <=( a3585a ) or ( a3586a );
 a4342a <=( a4341a ) or ( a4338a );
 a4343a <=( a4342a ) or ( a4335a );
 a4344a <=( a4343a ) or ( a4328a );
 a4348a <=( a3582a ) or ( a3583a );
 a4349a <=( a3584a ) or ( a4348a );
 a4352a <=( a3580a ) or ( a3581a );
 a4355a <=( a3578a ) or ( a3579a );
 a4356a <=( a4355a ) or ( a4352a );
 a4357a <=( a4356a ) or ( a4349a );
 a4360a <=( a3576a ) or ( a3577a );
 a4363a <=( a3574a ) or ( a3575a );
 a4364a <=( a4363a ) or ( a4360a );
 a4367a <=( a3572a ) or ( a3573a );
 a4370a <=( a3570a ) or ( a3571a );
 a4371a <=( a4370a ) or ( a4367a );
 a4372a <=( a4371a ) or ( a4364a );
 a4373a <=( a4372a ) or ( a4357a );
 a4374a <=( a4373a ) or ( a4344a );
 a4378a <=( a3567a ) or ( a3568a );
 a4379a <=( a3569a ) or ( a4378a );
 a4382a <=( a3565a ) or ( a3566a );
 a4385a <=( a3563a ) or ( a3564a );
 a4386a <=( a4385a ) or ( a4382a );
 a4387a <=( a4386a ) or ( a4379a );
 a4390a <=( a3561a ) or ( a3562a );
 a4393a <=( a3559a ) or ( a3560a );
 a4394a <=( a4393a ) or ( a4390a );
 a4397a <=( a3557a ) or ( a3558a );
 a4400a <=( a3555a ) or ( a3556a );
 a4401a <=( a4400a ) or ( a4397a );
 a4402a <=( a4401a ) or ( a4394a );
 a4403a <=( a4402a ) or ( a4387a );
 a4407a <=( a3552a ) or ( a3553a );
 a4408a <=( a3554a ) or ( a4407a );
 a4411a <=( a3550a ) or ( a3551a );
 a4414a <=( a3548a ) or ( a3549a );
 a4415a <=( a4414a ) or ( a4411a );
 a4416a <=( a4415a ) or ( a4408a );
 a4419a <=( a3546a ) or ( a3547a );
 a4422a <=( a3544a ) or ( a3545a );
 a4423a <=( a4422a ) or ( a4419a );
 a4426a <=( a3542a ) or ( a3543a );
 a4429a <=( a3540a ) or ( a3541a );
 a4430a <=( a4429a ) or ( a4426a );
 a4431a <=( a4430a ) or ( a4423a );
 a4432a <=( a4431a ) or ( a4416a );
 a4433a <=( a4432a ) or ( a4403a );
 a4434a <=( a4433a ) or ( a4374a );
 a4438a <=( a3537a ) or ( a3538a );
 a4439a <=( a3539a ) or ( a4438a );
 a4442a <=( a3535a ) or ( a3536a );
 a4445a <=( a3533a ) or ( a3534a );
 a4446a <=( a4445a ) or ( a4442a );
 a4447a <=( a4446a ) or ( a4439a );
 a4450a <=( a3531a ) or ( a3532a );
 a4453a <=( a3529a ) or ( a3530a );
 a4454a <=( a4453a ) or ( a4450a );
 a4457a <=( a3527a ) or ( a3528a );
 a4460a <=( a3525a ) or ( a3526a );
 a4461a <=( a4460a ) or ( a4457a );
 a4462a <=( a4461a ) or ( a4454a );
 a4463a <=( a4462a ) or ( a4447a );
 a4467a <=( a3522a ) or ( a3523a );
 a4468a <=( a3524a ) or ( a4467a );
 a4471a <=( a3520a ) or ( a3521a );
 a4474a <=( a3518a ) or ( a3519a );
 a4475a <=( a4474a ) or ( a4471a );
 a4476a <=( a4475a ) or ( a4468a );
 a4479a <=( a3516a ) or ( a3517a );
 a4482a <=( a3514a ) or ( a3515a );
 a4483a <=( a4482a ) or ( a4479a );
 a4486a <=( a3512a ) or ( a3513a );
 a4489a <=( a3510a ) or ( a3511a );
 a4490a <=( a4489a ) or ( a4486a );
 a4491a <=( a4490a ) or ( a4483a );
 a4492a <=( a4491a ) or ( a4476a );
 a4493a <=( a4492a ) or ( a4463a );
 a4497a <=( a3507a ) or ( a3508a );
 a4498a <=( a3509a ) or ( a4497a );
 a4501a <=( a3505a ) or ( a3506a );
 a4504a <=( a3503a ) or ( a3504a );
 a4505a <=( a4504a ) or ( a4501a );
 a4506a <=( a4505a ) or ( a4498a );
 a4509a <=( a3501a ) or ( a3502a );
 a4512a <=( a3499a ) or ( a3500a );
 a4513a <=( a4512a ) or ( a4509a );
 a4516a <=( a3497a ) or ( a3498a );
 a4519a <=( a3495a ) or ( a3496a );
 a4520a <=( a4519a ) or ( a4516a );
 a4521a <=( a4520a ) or ( a4513a );
 a4522a <=( a4521a ) or ( a4506a );
 a4526a <=( a3492a ) or ( a3493a );
 a4527a <=( a3494a ) or ( a4526a );
 a4530a <=( a3490a ) or ( a3491a );
 a4533a <=( a3488a ) or ( a3489a );
 a4534a <=( a4533a ) or ( a4530a );
 a4535a <=( a4534a ) or ( a4527a );
 a4538a <=( a3486a ) or ( a3487a );
 a4541a <=( a3484a ) or ( a3485a );
 a4542a <=( a4541a ) or ( a4538a );
 a4545a <=( a3482a ) or ( a3483a );
 a4548a <=( a3480a ) or ( a3481a );
 a4549a <=( a4548a ) or ( a4545a );
 a4550a <=( a4549a ) or ( a4542a );
 a4551a <=( a4550a ) or ( a4535a );
 a4552a <=( a4551a ) or ( a4522a );
 a4553a <=( a4552a ) or ( a4493a );
 a4554a <=( a4553a ) or ( a4434a );
 a4558a <=( a3477a ) or ( a3478a );
 a4559a <=( a3479a ) or ( a4558a );
 a4562a <=( a3475a ) or ( a3476a );
 a4565a <=( a3473a ) or ( a3474a );
 a4566a <=( a4565a ) or ( a4562a );
 a4567a <=( a4566a ) or ( a4559a );
 a4570a <=( a3471a ) or ( a3472a );
 a4573a <=( a3469a ) or ( a3470a );
 a4574a <=( a4573a ) or ( a4570a );
 a4577a <=( a3467a ) or ( a3468a );
 a4580a <=( a3465a ) or ( a3466a );
 a4581a <=( a4580a ) or ( a4577a );
 a4582a <=( a4581a ) or ( a4574a );
 a4583a <=( a4582a ) or ( a4567a );
 a4587a <=( a3462a ) or ( a3463a );
 a4588a <=( a3464a ) or ( a4587a );
 a4591a <=( a3460a ) or ( a3461a );
 a4594a <=( a3458a ) or ( a3459a );
 a4595a <=( a4594a ) or ( a4591a );
 a4596a <=( a4595a ) or ( a4588a );
 a4599a <=( a3456a ) or ( a3457a );
 a4602a <=( a3454a ) or ( a3455a );
 a4603a <=( a4602a ) or ( a4599a );
 a4606a <=( a3452a ) or ( a3453a );
 a4609a <=( a3450a ) or ( a3451a );
 a4610a <=( a4609a ) or ( a4606a );
 a4611a <=( a4610a ) or ( a4603a );
 a4612a <=( a4611a ) or ( a4596a );
 a4613a <=( a4612a ) or ( a4583a );
 a4617a <=( a3447a ) or ( a3448a );
 a4618a <=( a3449a ) or ( a4617a );
 a4621a <=( a3445a ) or ( a3446a );
 a4624a <=( a3443a ) or ( a3444a );
 a4625a <=( a4624a ) or ( a4621a );
 a4626a <=( a4625a ) or ( a4618a );
 a4629a <=( a3441a ) or ( a3442a );
 a4632a <=( a3439a ) or ( a3440a );
 a4633a <=( a4632a ) or ( a4629a );
 a4636a <=( a3437a ) or ( a3438a );
 a4639a <=( a3435a ) or ( a3436a );
 a4640a <=( a4639a ) or ( a4636a );
 a4641a <=( a4640a ) or ( a4633a );
 a4642a <=( a4641a ) or ( a4626a );
 a4646a <=( a3432a ) or ( a3433a );
 a4647a <=( a3434a ) or ( a4646a );
 a4650a <=( a3430a ) or ( a3431a );
 a4653a <=( a3428a ) or ( a3429a );
 a4654a <=( a4653a ) or ( a4650a );
 a4655a <=( a4654a ) or ( a4647a );
 a4658a <=( a3426a ) or ( a3427a );
 a4661a <=( a3424a ) or ( a3425a );
 a4662a <=( a4661a ) or ( a4658a );
 a4665a <=( a3422a ) or ( a3423a );
 a4668a <=( a3420a ) or ( a3421a );
 a4669a <=( a4668a ) or ( a4665a );
 a4670a <=( a4669a ) or ( a4662a );
 a4671a <=( a4670a ) or ( a4655a );
 a4672a <=( a4671a ) or ( a4642a );
 a4673a <=( a4672a ) or ( a4613a );
 a4677a <=( a3417a ) or ( a3418a );
 a4678a <=( a3419a ) or ( a4677a );
 a4681a <=( a3415a ) or ( a3416a );
 a4684a <=( a3413a ) or ( a3414a );
 a4685a <=( a4684a ) or ( a4681a );
 a4686a <=( a4685a ) or ( a4678a );
 a4689a <=( a3411a ) or ( a3412a );
 a4692a <=( a3409a ) or ( a3410a );
 a4693a <=( a4692a ) or ( a4689a );
 a4696a <=( a3407a ) or ( a3408a );
 a4699a <=( a3405a ) or ( a3406a );
 a4700a <=( a4699a ) or ( a4696a );
 a4701a <=( a4700a ) or ( a4693a );
 a4702a <=( a4701a ) or ( a4686a );
 a4706a <=( a3402a ) or ( a3403a );
 a4707a <=( a3404a ) or ( a4706a );
 a4710a <=( a3400a ) or ( a3401a );
 a4713a <=( a3398a ) or ( a3399a );
 a4714a <=( a4713a ) or ( a4710a );
 a4715a <=( a4714a ) or ( a4707a );
 a4718a <=( a3396a ) or ( a3397a );
 a4721a <=( a3394a ) or ( a3395a );
 a4722a <=( a4721a ) or ( a4718a );
 a4725a <=( a3392a ) or ( a3393a );
 a4728a <=( a3390a ) or ( a3391a );
 a4729a <=( a4728a ) or ( a4725a );
 a4730a <=( a4729a ) or ( a4722a );
 a4731a <=( a4730a ) or ( a4715a );
 a4732a <=( a4731a ) or ( a4702a );
 a4736a <=( a3387a ) or ( a3388a );
 a4737a <=( a3389a ) or ( a4736a );
 a4740a <=( a3385a ) or ( a3386a );
 a4743a <=( a3383a ) or ( a3384a );
 a4744a <=( a4743a ) or ( a4740a );
 a4745a <=( a4744a ) or ( a4737a );
 a4748a <=( a3381a ) or ( a3382a );
 a4751a <=( a3379a ) or ( a3380a );
 a4752a <=( a4751a ) or ( a4748a );
 a4755a <=( a3377a ) or ( a3378a );
 a4758a <=( a3375a ) or ( a3376a );
 a4759a <=( a4758a ) or ( a4755a );
 a4760a <=( a4759a ) or ( a4752a );
 a4761a <=( a4760a ) or ( a4745a );
 a4765a <=( a3372a ) or ( a3373a );
 a4766a <=( a3374a ) or ( a4765a );
 a4769a <=( a3370a ) or ( a3371a );
 a4772a <=( a3368a ) or ( a3369a );
 a4773a <=( a4772a ) or ( a4769a );
 a4774a <=( a4773a ) or ( a4766a );
 a4777a <=( a3366a ) or ( a3367a );
 a4780a <=( a3364a ) or ( a3365a );
 a4781a <=( a4780a ) or ( a4777a );
 a4784a <=( a3362a ) or ( a3363a );
 a4787a <=( a3360a ) or ( a3361a );
 a4788a <=( a4787a ) or ( a4784a );
 a4789a <=( a4788a ) or ( a4781a );
 a4790a <=( a4789a ) or ( a4774a );
 a4791a <=( a4790a ) or ( a4761a );
 a4792a <=( a4791a ) or ( a4732a );
 a4793a <=( a4792a ) or ( a4673a );
 a4794a <=( a4793a ) or ( a4554a );
 a4795a <=( a4794a ) or ( a4315a );
 a4799a <=( a3357a ) or ( a3358a );
 a4800a <=( a3359a ) or ( a4799a );
 a4803a <=( a3355a ) or ( a3356a );
 a4806a <=( a3353a ) or ( a3354a );
 a4807a <=( a4806a ) or ( a4803a );
 a4808a <=( a4807a ) or ( a4800a );
 a4811a <=( a3351a ) or ( a3352a );
 a4814a <=( a3349a ) or ( a3350a );
 a4815a <=( a4814a ) or ( a4811a );
 a4818a <=( a3347a ) or ( a3348a );
 a4821a <=( a3345a ) or ( a3346a );
 a4822a <=( a4821a ) or ( a4818a );
 a4823a <=( a4822a ) or ( a4815a );
 a4824a <=( a4823a ) or ( a4808a );
 a4828a <=( a3342a ) or ( a3343a );
 a4829a <=( a3344a ) or ( a4828a );
 a4832a <=( a3340a ) or ( a3341a );
 a4835a <=( a3338a ) or ( a3339a );
 a4836a <=( a4835a ) or ( a4832a );
 a4837a <=( a4836a ) or ( a4829a );
 a4840a <=( a3336a ) or ( a3337a );
 a4843a <=( a3334a ) or ( a3335a );
 a4844a <=( a4843a ) or ( a4840a );
 a4847a <=( a3332a ) or ( a3333a );
 a4850a <=( a3330a ) or ( a3331a );
 a4851a <=( a4850a ) or ( a4847a );
 a4852a <=( a4851a ) or ( a4844a );
 a4853a <=( a4852a ) or ( a4837a );
 a4854a <=( a4853a ) or ( a4824a );
 a4858a <=( a3327a ) or ( a3328a );
 a4859a <=( a3329a ) or ( a4858a );
 a4862a <=( a3325a ) or ( a3326a );
 a4865a <=( a3323a ) or ( a3324a );
 a4866a <=( a4865a ) or ( a4862a );
 a4867a <=( a4866a ) or ( a4859a );
 a4870a <=( a3321a ) or ( a3322a );
 a4873a <=( a3319a ) or ( a3320a );
 a4874a <=( a4873a ) or ( a4870a );
 a4877a <=( a3317a ) or ( a3318a );
 a4880a <=( a3315a ) or ( a3316a );
 a4881a <=( a4880a ) or ( a4877a );
 a4882a <=( a4881a ) or ( a4874a );
 a4883a <=( a4882a ) or ( a4867a );
 a4887a <=( a3312a ) or ( a3313a );
 a4888a <=( a3314a ) or ( a4887a );
 a4891a <=( a3310a ) or ( a3311a );
 a4894a <=( a3308a ) or ( a3309a );
 a4895a <=( a4894a ) or ( a4891a );
 a4896a <=( a4895a ) or ( a4888a );
 a4899a <=( a3306a ) or ( a3307a );
 a4902a <=( a3304a ) or ( a3305a );
 a4903a <=( a4902a ) or ( a4899a );
 a4906a <=( a3302a ) or ( a3303a );
 a4909a <=( a3300a ) or ( a3301a );
 a4910a <=( a4909a ) or ( a4906a );
 a4911a <=( a4910a ) or ( a4903a );
 a4912a <=( a4911a ) or ( a4896a );
 a4913a <=( a4912a ) or ( a4883a );
 a4914a <=( a4913a ) or ( a4854a );
 a4918a <=( a3297a ) or ( a3298a );
 a4919a <=( a3299a ) or ( a4918a );
 a4922a <=( a3295a ) or ( a3296a );
 a4925a <=( a3293a ) or ( a3294a );
 a4926a <=( a4925a ) or ( a4922a );
 a4927a <=( a4926a ) or ( a4919a );
 a4930a <=( a3291a ) or ( a3292a );
 a4933a <=( a3289a ) or ( a3290a );
 a4934a <=( a4933a ) or ( a4930a );
 a4937a <=( a3287a ) or ( a3288a );
 a4940a <=( a3285a ) or ( a3286a );
 a4941a <=( a4940a ) or ( a4937a );
 a4942a <=( a4941a ) or ( a4934a );
 a4943a <=( a4942a ) or ( a4927a );
 a4947a <=( a3282a ) or ( a3283a );
 a4948a <=( a3284a ) or ( a4947a );
 a4951a <=( a3280a ) or ( a3281a );
 a4954a <=( a3278a ) or ( a3279a );
 a4955a <=( a4954a ) or ( a4951a );
 a4956a <=( a4955a ) or ( a4948a );
 a4959a <=( a3276a ) or ( a3277a );
 a4962a <=( a3274a ) or ( a3275a );
 a4963a <=( a4962a ) or ( a4959a );
 a4966a <=( a3272a ) or ( a3273a );
 a4969a <=( a3270a ) or ( a3271a );
 a4970a <=( a4969a ) or ( a4966a );
 a4971a <=( a4970a ) or ( a4963a );
 a4972a <=( a4971a ) or ( a4956a );
 a4973a <=( a4972a ) or ( a4943a );
 a4977a <=( a3267a ) or ( a3268a );
 a4978a <=( a3269a ) or ( a4977a );
 a4981a <=( a3265a ) or ( a3266a );
 a4984a <=( a3263a ) or ( a3264a );
 a4985a <=( a4984a ) or ( a4981a );
 a4986a <=( a4985a ) or ( a4978a );
 a4989a <=( a3261a ) or ( a3262a );
 a4992a <=( a3259a ) or ( a3260a );
 a4993a <=( a4992a ) or ( a4989a );
 a4996a <=( a3257a ) or ( a3258a );
 a4999a <=( a3255a ) or ( a3256a );
 a5000a <=( a4999a ) or ( a4996a );
 a5001a <=( a5000a ) or ( a4993a );
 a5002a <=( a5001a ) or ( a4986a );
 a5006a <=( a3252a ) or ( a3253a );
 a5007a <=( a3254a ) or ( a5006a );
 a5010a <=( a3250a ) or ( a3251a );
 a5013a <=( a3248a ) or ( a3249a );
 a5014a <=( a5013a ) or ( a5010a );
 a5015a <=( a5014a ) or ( a5007a );
 a5018a <=( a3246a ) or ( a3247a );
 a5021a <=( a3244a ) or ( a3245a );
 a5022a <=( a5021a ) or ( a5018a );
 a5025a <=( a3242a ) or ( a3243a );
 a5028a <=( a3240a ) or ( a3241a );
 a5029a <=( a5028a ) or ( a5025a );
 a5030a <=( a5029a ) or ( a5022a );
 a5031a <=( a5030a ) or ( a5015a );
 a5032a <=( a5031a ) or ( a5002a );
 a5033a <=( a5032a ) or ( a4973a );
 a5034a <=( a5033a ) or ( a4914a );
 a5038a <=( a3237a ) or ( a3238a );
 a5039a <=( a3239a ) or ( a5038a );
 a5042a <=( a3235a ) or ( a3236a );
 a5045a <=( a3233a ) or ( a3234a );
 a5046a <=( a5045a ) or ( a5042a );
 a5047a <=( a5046a ) or ( a5039a );
 a5050a <=( a3231a ) or ( a3232a );
 a5053a <=( a3229a ) or ( a3230a );
 a5054a <=( a5053a ) or ( a5050a );
 a5057a <=( a3227a ) or ( a3228a );
 a5060a <=( a3225a ) or ( a3226a );
 a5061a <=( a5060a ) or ( a5057a );
 a5062a <=( a5061a ) or ( a5054a );
 a5063a <=( a5062a ) or ( a5047a );
 a5067a <=( a3222a ) or ( a3223a );
 a5068a <=( a3224a ) or ( a5067a );
 a5071a <=( a3220a ) or ( a3221a );
 a5074a <=( a3218a ) or ( a3219a );
 a5075a <=( a5074a ) or ( a5071a );
 a5076a <=( a5075a ) or ( a5068a );
 a5079a <=( a3216a ) or ( a3217a );
 a5082a <=( a3214a ) or ( a3215a );
 a5083a <=( a5082a ) or ( a5079a );
 a5086a <=( a3212a ) or ( a3213a );
 a5089a <=( a3210a ) or ( a3211a );
 a5090a <=( a5089a ) or ( a5086a );
 a5091a <=( a5090a ) or ( a5083a );
 a5092a <=( a5091a ) or ( a5076a );
 a5093a <=( a5092a ) or ( a5063a );
 a5097a <=( a3207a ) or ( a3208a );
 a5098a <=( a3209a ) or ( a5097a );
 a5101a <=( a3205a ) or ( a3206a );
 a5104a <=( a3203a ) or ( a3204a );
 a5105a <=( a5104a ) or ( a5101a );
 a5106a <=( a5105a ) or ( a5098a );
 a5109a <=( a3201a ) or ( a3202a );
 a5112a <=( a3199a ) or ( a3200a );
 a5113a <=( a5112a ) or ( a5109a );
 a5116a <=( a3197a ) or ( a3198a );
 a5119a <=( a3195a ) or ( a3196a );
 a5120a <=( a5119a ) or ( a5116a );
 a5121a <=( a5120a ) or ( a5113a );
 a5122a <=( a5121a ) or ( a5106a );
 a5126a <=( a3192a ) or ( a3193a );
 a5127a <=( a3194a ) or ( a5126a );
 a5130a <=( a3190a ) or ( a3191a );
 a5133a <=( a3188a ) or ( a3189a );
 a5134a <=( a5133a ) or ( a5130a );
 a5135a <=( a5134a ) or ( a5127a );
 a5138a <=( a3186a ) or ( a3187a );
 a5141a <=( a3184a ) or ( a3185a );
 a5142a <=( a5141a ) or ( a5138a );
 a5145a <=( a3182a ) or ( a3183a );
 a5148a <=( a3180a ) or ( a3181a );
 a5149a <=( a5148a ) or ( a5145a );
 a5150a <=( a5149a ) or ( a5142a );
 a5151a <=( a5150a ) or ( a5135a );
 a5152a <=( a5151a ) or ( a5122a );
 a5153a <=( a5152a ) or ( a5093a );
 a5157a <=( a3177a ) or ( a3178a );
 a5158a <=( a3179a ) or ( a5157a );
 a5161a <=( a3175a ) or ( a3176a );
 a5164a <=( a3173a ) or ( a3174a );
 a5165a <=( a5164a ) or ( a5161a );
 a5166a <=( a5165a ) or ( a5158a );
 a5169a <=( a3171a ) or ( a3172a );
 a5172a <=( a3169a ) or ( a3170a );
 a5173a <=( a5172a ) or ( a5169a );
 a5176a <=( a3167a ) or ( a3168a );
 a5179a <=( a3165a ) or ( a3166a );
 a5180a <=( a5179a ) or ( a5176a );
 a5181a <=( a5180a ) or ( a5173a );
 a5182a <=( a5181a ) or ( a5166a );
 a5186a <=( a3162a ) or ( a3163a );
 a5187a <=( a3164a ) or ( a5186a );
 a5190a <=( a3160a ) or ( a3161a );
 a5193a <=( a3158a ) or ( a3159a );
 a5194a <=( a5193a ) or ( a5190a );
 a5195a <=( a5194a ) or ( a5187a );
 a5198a <=( a3156a ) or ( a3157a );
 a5201a <=( a3154a ) or ( a3155a );
 a5202a <=( a5201a ) or ( a5198a );
 a5205a <=( a3152a ) or ( a3153a );
 a5208a <=( a3150a ) or ( a3151a );
 a5209a <=( a5208a ) or ( a5205a );
 a5210a <=( a5209a ) or ( a5202a );
 a5211a <=( a5210a ) or ( a5195a );
 a5212a <=( a5211a ) or ( a5182a );
 a5216a <=( a3147a ) or ( a3148a );
 a5217a <=( a3149a ) or ( a5216a );
 a5220a <=( a3145a ) or ( a3146a );
 a5223a <=( a3143a ) or ( a3144a );
 a5224a <=( a5223a ) or ( a5220a );
 a5225a <=( a5224a ) or ( a5217a );
 a5228a <=( a3141a ) or ( a3142a );
 a5231a <=( a3139a ) or ( a3140a );
 a5232a <=( a5231a ) or ( a5228a );
 a5235a <=( a3137a ) or ( a3138a );
 a5238a <=( a3135a ) or ( a3136a );
 a5239a <=( a5238a ) or ( a5235a );
 a5240a <=( a5239a ) or ( a5232a );
 a5241a <=( a5240a ) or ( a5225a );
 a5245a <=( a3132a ) or ( a3133a );
 a5246a <=( a3134a ) or ( a5245a );
 a5249a <=( a3130a ) or ( a3131a );
 a5252a <=( a3128a ) or ( a3129a );
 a5253a <=( a5252a ) or ( a5249a );
 a5254a <=( a5253a ) or ( a5246a );
 a5257a <=( a3126a ) or ( a3127a );
 a5260a <=( a3124a ) or ( a3125a );
 a5261a <=( a5260a ) or ( a5257a );
 a5264a <=( a3122a ) or ( a3123a );
 a5267a <=( a3120a ) or ( a3121a );
 a5268a <=( a5267a ) or ( a5264a );
 a5269a <=( a5268a ) or ( a5261a );
 a5270a <=( a5269a ) or ( a5254a );
 a5271a <=( a5270a ) or ( a5241a );
 a5272a <=( a5271a ) or ( a5212a );
 a5273a <=( a5272a ) or ( a5153a );
 a5274a <=( a5273a ) or ( a5034a );
 a5278a <=( a3117a ) or ( a3118a );
 a5279a <=( a3119a ) or ( a5278a );
 a5282a <=( a3115a ) or ( a3116a );
 a5285a <=( a3113a ) or ( a3114a );
 a5286a <=( a5285a ) or ( a5282a );
 a5287a <=( a5286a ) or ( a5279a );
 a5290a <=( a3111a ) or ( a3112a );
 a5293a <=( a3109a ) or ( a3110a );
 a5294a <=( a5293a ) or ( a5290a );
 a5297a <=( a3107a ) or ( a3108a );
 a5300a <=( a3105a ) or ( a3106a );
 a5301a <=( a5300a ) or ( a5297a );
 a5302a <=( a5301a ) or ( a5294a );
 a5303a <=( a5302a ) or ( a5287a );
 a5307a <=( a3102a ) or ( a3103a );
 a5308a <=( a3104a ) or ( a5307a );
 a5311a <=( a3100a ) or ( a3101a );
 a5314a <=( a3098a ) or ( a3099a );
 a5315a <=( a5314a ) or ( a5311a );
 a5316a <=( a5315a ) or ( a5308a );
 a5319a <=( a3096a ) or ( a3097a );
 a5322a <=( a3094a ) or ( a3095a );
 a5323a <=( a5322a ) or ( a5319a );
 a5326a <=( a3092a ) or ( a3093a );
 a5329a <=( a3090a ) or ( a3091a );
 a5330a <=( a5329a ) or ( a5326a );
 a5331a <=( a5330a ) or ( a5323a );
 a5332a <=( a5331a ) or ( a5316a );
 a5333a <=( a5332a ) or ( a5303a );
 a5337a <=( a3087a ) or ( a3088a );
 a5338a <=( a3089a ) or ( a5337a );
 a5341a <=( a3085a ) or ( a3086a );
 a5344a <=( a3083a ) or ( a3084a );
 a5345a <=( a5344a ) or ( a5341a );
 a5346a <=( a5345a ) or ( a5338a );
 a5349a <=( a3081a ) or ( a3082a );
 a5352a <=( a3079a ) or ( a3080a );
 a5353a <=( a5352a ) or ( a5349a );
 a5356a <=( a3077a ) or ( a3078a );
 a5359a <=( a3075a ) or ( a3076a );
 a5360a <=( a5359a ) or ( a5356a );
 a5361a <=( a5360a ) or ( a5353a );
 a5362a <=( a5361a ) or ( a5346a );
 a5366a <=( a3072a ) or ( a3073a );
 a5367a <=( a3074a ) or ( a5366a );
 a5370a <=( a3070a ) or ( a3071a );
 a5373a <=( a3068a ) or ( a3069a );
 a5374a <=( a5373a ) or ( a5370a );
 a5375a <=( a5374a ) or ( a5367a );
 a5378a <=( a3066a ) or ( a3067a );
 a5381a <=( a3064a ) or ( a3065a );
 a5382a <=( a5381a ) or ( a5378a );
 a5385a <=( a3062a ) or ( a3063a );
 a5388a <=( a3060a ) or ( a3061a );
 a5389a <=( a5388a ) or ( a5385a );
 a5390a <=( a5389a ) or ( a5382a );
 a5391a <=( a5390a ) or ( a5375a );
 a5392a <=( a5391a ) or ( a5362a );
 a5393a <=( a5392a ) or ( a5333a );
 a5397a <=( a3057a ) or ( a3058a );
 a5398a <=( a3059a ) or ( a5397a );
 a5401a <=( a3055a ) or ( a3056a );
 a5404a <=( a3053a ) or ( a3054a );
 a5405a <=( a5404a ) or ( a5401a );
 a5406a <=( a5405a ) or ( a5398a );
 a5409a <=( a3051a ) or ( a3052a );
 a5412a <=( a3049a ) or ( a3050a );
 a5413a <=( a5412a ) or ( a5409a );
 a5416a <=( a3047a ) or ( a3048a );
 a5419a <=( a3045a ) or ( a3046a );
 a5420a <=( a5419a ) or ( a5416a );
 a5421a <=( a5420a ) or ( a5413a );
 a5422a <=( a5421a ) or ( a5406a );
 a5426a <=( a3042a ) or ( a3043a );
 a5427a <=( a3044a ) or ( a5426a );
 a5430a <=( a3040a ) or ( a3041a );
 a5433a <=( a3038a ) or ( a3039a );
 a5434a <=( a5433a ) or ( a5430a );
 a5435a <=( a5434a ) or ( a5427a );
 a5438a <=( a3036a ) or ( a3037a );
 a5441a <=( a3034a ) or ( a3035a );
 a5442a <=( a5441a ) or ( a5438a );
 a5445a <=( a3032a ) or ( a3033a );
 a5448a <=( a3030a ) or ( a3031a );
 a5449a <=( a5448a ) or ( a5445a );
 a5450a <=( a5449a ) or ( a5442a );
 a5451a <=( a5450a ) or ( a5435a );
 a5452a <=( a5451a ) or ( a5422a );
 a5456a <=( a3027a ) or ( a3028a );
 a5457a <=( a3029a ) or ( a5456a );
 a5460a <=( a3025a ) or ( a3026a );
 a5463a <=( a3023a ) or ( a3024a );
 a5464a <=( a5463a ) or ( a5460a );
 a5465a <=( a5464a ) or ( a5457a );
 a5468a <=( a3021a ) or ( a3022a );
 a5471a <=( a3019a ) or ( a3020a );
 a5472a <=( a5471a ) or ( a5468a );
 a5475a <=( a3017a ) or ( a3018a );
 a5478a <=( a3015a ) or ( a3016a );
 a5479a <=( a5478a ) or ( a5475a );
 a5480a <=( a5479a ) or ( a5472a );
 a5481a <=( a5480a ) or ( a5465a );
 a5485a <=( a3012a ) or ( a3013a );
 a5486a <=( a3014a ) or ( a5485a );
 a5489a <=( a3010a ) or ( a3011a );
 a5492a <=( a3008a ) or ( a3009a );
 a5493a <=( a5492a ) or ( a5489a );
 a5494a <=( a5493a ) or ( a5486a );
 a5497a <=( a3006a ) or ( a3007a );
 a5500a <=( a3004a ) or ( a3005a );
 a5501a <=( a5500a ) or ( a5497a );
 a5504a <=( a3002a ) or ( a3003a );
 a5507a <=( a3000a ) or ( a3001a );
 a5508a <=( a5507a ) or ( a5504a );
 a5509a <=( a5508a ) or ( a5501a );
 a5510a <=( a5509a ) or ( a5494a );
 a5511a <=( a5510a ) or ( a5481a );
 a5512a <=( a5511a ) or ( a5452a );
 a5513a <=( a5512a ) or ( a5393a );
 a5517a <=( a2997a ) or ( a2998a );
 a5518a <=( a2999a ) or ( a5517a );
 a5521a <=( a2995a ) or ( a2996a );
 a5524a <=( a2993a ) or ( a2994a );
 a5525a <=( a5524a ) or ( a5521a );
 a5526a <=( a5525a ) or ( a5518a );
 a5529a <=( a2991a ) or ( a2992a );
 a5532a <=( a2989a ) or ( a2990a );
 a5533a <=( a5532a ) or ( a5529a );
 a5536a <=( a2987a ) or ( a2988a );
 a5539a <=( a2985a ) or ( a2986a );
 a5540a <=( a5539a ) or ( a5536a );
 a5541a <=( a5540a ) or ( a5533a );
 a5542a <=( a5541a ) or ( a5526a );
 a5546a <=( a2982a ) or ( a2983a );
 a5547a <=( a2984a ) or ( a5546a );
 a5550a <=( a2980a ) or ( a2981a );
 a5553a <=( a2978a ) or ( a2979a );
 a5554a <=( a5553a ) or ( a5550a );
 a5555a <=( a5554a ) or ( a5547a );
 a5558a <=( a2976a ) or ( a2977a );
 a5561a <=( a2974a ) or ( a2975a );
 a5562a <=( a5561a ) or ( a5558a );
 a5565a <=( a2972a ) or ( a2973a );
 a5568a <=( a2970a ) or ( a2971a );
 a5569a <=( a5568a ) or ( a5565a );
 a5570a <=( a5569a ) or ( a5562a );
 a5571a <=( a5570a ) or ( a5555a );
 a5572a <=( a5571a ) or ( a5542a );
 a5576a <=( a2967a ) or ( a2968a );
 a5577a <=( a2969a ) or ( a5576a );
 a5580a <=( a2965a ) or ( a2966a );
 a5583a <=( a2963a ) or ( a2964a );
 a5584a <=( a5583a ) or ( a5580a );
 a5585a <=( a5584a ) or ( a5577a );
 a5588a <=( a2961a ) or ( a2962a );
 a5591a <=( a2959a ) or ( a2960a );
 a5592a <=( a5591a ) or ( a5588a );
 a5595a <=( a2957a ) or ( a2958a );
 a5598a <=( a2955a ) or ( a2956a );
 a5599a <=( a5598a ) or ( a5595a );
 a5600a <=( a5599a ) or ( a5592a );
 a5601a <=( a5600a ) or ( a5585a );
 a5605a <=( a2952a ) or ( a2953a );
 a5606a <=( a2954a ) or ( a5605a );
 a5609a <=( a2950a ) or ( a2951a );
 a5612a <=( a2948a ) or ( a2949a );
 a5613a <=( a5612a ) or ( a5609a );
 a5614a <=( a5613a ) or ( a5606a );
 a5617a <=( a2946a ) or ( a2947a );
 a5620a <=( a2944a ) or ( a2945a );
 a5621a <=( a5620a ) or ( a5617a );
 a5624a <=( a2942a ) or ( a2943a );
 a5627a <=( a2940a ) or ( a2941a );
 a5628a <=( a5627a ) or ( a5624a );
 a5629a <=( a5628a ) or ( a5621a );
 a5630a <=( a5629a ) or ( a5614a );
 a5631a <=( a5630a ) or ( a5601a );
 a5632a <=( a5631a ) or ( a5572a );
 a5636a <=( a2937a ) or ( a2938a );
 a5637a <=( a2939a ) or ( a5636a );
 a5640a <=( a2935a ) or ( a2936a );
 a5643a <=( a2933a ) or ( a2934a );
 a5644a <=( a5643a ) or ( a5640a );
 a5645a <=( a5644a ) or ( a5637a );
 a5648a <=( a2931a ) or ( a2932a );
 a5651a <=( a2929a ) or ( a2930a );
 a5652a <=( a5651a ) or ( a5648a );
 a5655a <=( a2927a ) or ( a2928a );
 a5658a <=( a2925a ) or ( a2926a );
 a5659a <=( a5658a ) or ( a5655a );
 a5660a <=( a5659a ) or ( a5652a );
 a5661a <=( a5660a ) or ( a5645a );
 a5665a <=( a2922a ) or ( a2923a );
 a5666a <=( a2924a ) or ( a5665a );
 a5669a <=( a2920a ) or ( a2921a );
 a5672a <=( a2918a ) or ( a2919a );
 a5673a <=( a5672a ) or ( a5669a );
 a5674a <=( a5673a ) or ( a5666a );
 a5677a <=( a2916a ) or ( a2917a );
 a5680a <=( a2914a ) or ( a2915a );
 a5681a <=( a5680a ) or ( a5677a );
 a5684a <=( a2912a ) or ( a2913a );
 a5687a <=( a2910a ) or ( a2911a );
 a5688a <=( a5687a ) or ( a5684a );
 a5689a <=( a5688a ) or ( a5681a );
 a5690a <=( a5689a ) or ( a5674a );
 a5691a <=( a5690a ) or ( a5661a );
 a5695a <=( a2907a ) or ( a2908a );
 a5696a <=( a2909a ) or ( a5695a );
 a5699a <=( a2905a ) or ( a2906a );
 a5702a <=( a2903a ) or ( a2904a );
 a5703a <=( a5702a ) or ( a5699a );
 a5704a <=( a5703a ) or ( a5696a );
 a5707a <=( a2901a ) or ( a2902a );
 a5710a <=( a2899a ) or ( a2900a );
 a5711a <=( a5710a ) or ( a5707a );
 a5714a <=( a2897a ) or ( a2898a );
 a5717a <=( a2895a ) or ( a2896a );
 a5718a <=( a5717a ) or ( a5714a );
 a5719a <=( a5718a ) or ( a5711a );
 a5720a <=( a5719a ) or ( a5704a );
 a5724a <=( a2892a ) or ( a2893a );
 a5725a <=( a2894a ) or ( a5724a );
 a5728a <=( a2890a ) or ( a2891a );
 a5731a <=( a2888a ) or ( a2889a );
 a5732a <=( a5731a ) or ( a5728a );
 a5733a <=( a5732a ) or ( a5725a );
 a5736a <=( a2886a ) or ( a2887a );
 a5739a <=( a2884a ) or ( a2885a );
 a5740a <=( a5739a ) or ( a5736a );
 a5743a <=( a2882a ) or ( a2883a );
 a5746a <=( a2880a ) or ( a2881a );
 a5747a <=( a5746a ) or ( a5743a );
 a5748a <=( a5747a ) or ( a5740a );
 a5749a <=( a5748a ) or ( a5733a );
 a5750a <=( a5749a ) or ( a5720a );
 a5751a <=( a5750a ) or ( a5691a );
 a5752a <=( a5751a ) or ( a5632a );
 a5753a <=( a5752a ) or ( a5513a );
 a5754a <=( a5753a ) or ( a5274a );
 a5755a <=( a5754a ) or ( a4795a );
 a5759a <=( a2877a ) or ( a2878a );
 a5760a <=( a2879a ) or ( a5759a );
 a5763a <=( a2875a ) or ( a2876a );
 a5766a <=( a2873a ) or ( a2874a );
 a5767a <=( a5766a ) or ( a5763a );
 a5768a <=( a5767a ) or ( a5760a );
 a5771a <=( a2871a ) or ( a2872a );
 a5774a <=( a2869a ) or ( a2870a );
 a5775a <=( a5774a ) or ( a5771a );
 a5778a <=( a2867a ) or ( a2868a );
 a5781a <=( a2865a ) or ( a2866a );
 a5782a <=( a5781a ) or ( a5778a );
 a5783a <=( a5782a ) or ( a5775a );
 a5784a <=( a5783a ) or ( a5768a );
 a5788a <=( a2862a ) or ( a2863a );
 a5789a <=( a2864a ) or ( a5788a );
 a5792a <=( a2860a ) or ( a2861a );
 a5795a <=( a2858a ) or ( a2859a );
 a5796a <=( a5795a ) or ( a5792a );
 a5797a <=( a5796a ) or ( a5789a );
 a5800a <=( a2856a ) or ( a2857a );
 a5803a <=( a2854a ) or ( a2855a );
 a5804a <=( a5803a ) or ( a5800a );
 a5807a <=( a2852a ) or ( a2853a );
 a5810a <=( a2850a ) or ( a2851a );
 a5811a <=( a5810a ) or ( a5807a );
 a5812a <=( a5811a ) or ( a5804a );
 a5813a <=( a5812a ) or ( a5797a );
 a5814a <=( a5813a ) or ( a5784a );
 a5818a <=( a2847a ) or ( a2848a );
 a5819a <=( a2849a ) or ( a5818a );
 a5822a <=( a2845a ) or ( a2846a );
 a5825a <=( a2843a ) or ( a2844a );
 a5826a <=( a5825a ) or ( a5822a );
 a5827a <=( a5826a ) or ( a5819a );
 a5830a <=( a2841a ) or ( a2842a );
 a5833a <=( a2839a ) or ( a2840a );
 a5834a <=( a5833a ) or ( a5830a );
 a5837a <=( a2837a ) or ( a2838a );
 a5840a <=( a2835a ) or ( a2836a );
 a5841a <=( a5840a ) or ( a5837a );
 a5842a <=( a5841a ) or ( a5834a );
 a5843a <=( a5842a ) or ( a5827a );
 a5847a <=( a2832a ) or ( a2833a );
 a5848a <=( a2834a ) or ( a5847a );
 a5851a <=( a2830a ) or ( a2831a );
 a5854a <=( a2828a ) or ( a2829a );
 a5855a <=( a5854a ) or ( a5851a );
 a5856a <=( a5855a ) or ( a5848a );
 a5859a <=( a2826a ) or ( a2827a );
 a5862a <=( a2824a ) or ( a2825a );
 a5863a <=( a5862a ) or ( a5859a );
 a5866a <=( a2822a ) or ( a2823a );
 a5869a <=( a2820a ) or ( a2821a );
 a5870a <=( a5869a ) or ( a5866a );
 a5871a <=( a5870a ) or ( a5863a );
 a5872a <=( a5871a ) or ( a5856a );
 a5873a <=( a5872a ) or ( a5843a );
 a5874a <=( a5873a ) or ( a5814a );
 a5878a <=( a2817a ) or ( a2818a );
 a5879a <=( a2819a ) or ( a5878a );
 a5882a <=( a2815a ) or ( a2816a );
 a5885a <=( a2813a ) or ( a2814a );
 a5886a <=( a5885a ) or ( a5882a );
 a5887a <=( a5886a ) or ( a5879a );
 a5890a <=( a2811a ) or ( a2812a );
 a5893a <=( a2809a ) or ( a2810a );
 a5894a <=( a5893a ) or ( a5890a );
 a5897a <=( a2807a ) or ( a2808a );
 a5900a <=( a2805a ) or ( a2806a );
 a5901a <=( a5900a ) or ( a5897a );
 a5902a <=( a5901a ) or ( a5894a );
 a5903a <=( a5902a ) or ( a5887a );
 a5907a <=( a2802a ) or ( a2803a );
 a5908a <=( a2804a ) or ( a5907a );
 a5911a <=( a2800a ) or ( a2801a );
 a5914a <=( a2798a ) or ( a2799a );
 a5915a <=( a5914a ) or ( a5911a );
 a5916a <=( a5915a ) or ( a5908a );
 a5919a <=( a2796a ) or ( a2797a );
 a5922a <=( a2794a ) or ( a2795a );
 a5923a <=( a5922a ) or ( a5919a );
 a5926a <=( a2792a ) or ( a2793a );
 a5929a <=( a2790a ) or ( a2791a );
 a5930a <=( a5929a ) or ( a5926a );
 a5931a <=( a5930a ) or ( a5923a );
 a5932a <=( a5931a ) or ( a5916a );
 a5933a <=( a5932a ) or ( a5903a );
 a5937a <=( a2787a ) or ( a2788a );
 a5938a <=( a2789a ) or ( a5937a );
 a5941a <=( a2785a ) or ( a2786a );
 a5944a <=( a2783a ) or ( a2784a );
 a5945a <=( a5944a ) or ( a5941a );
 a5946a <=( a5945a ) or ( a5938a );
 a5949a <=( a2781a ) or ( a2782a );
 a5952a <=( a2779a ) or ( a2780a );
 a5953a <=( a5952a ) or ( a5949a );
 a5956a <=( a2777a ) or ( a2778a );
 a5959a <=( a2775a ) or ( a2776a );
 a5960a <=( a5959a ) or ( a5956a );
 a5961a <=( a5960a ) or ( a5953a );
 a5962a <=( a5961a ) or ( a5946a );
 a5966a <=( a2772a ) or ( a2773a );
 a5967a <=( a2774a ) or ( a5966a );
 a5970a <=( a2770a ) or ( a2771a );
 a5973a <=( a2768a ) or ( a2769a );
 a5974a <=( a5973a ) or ( a5970a );
 a5975a <=( a5974a ) or ( a5967a );
 a5978a <=( a2766a ) or ( a2767a );
 a5981a <=( a2764a ) or ( a2765a );
 a5982a <=( a5981a ) or ( a5978a );
 a5985a <=( a2762a ) or ( a2763a );
 a5988a <=( a2760a ) or ( a2761a );
 a5989a <=( a5988a ) or ( a5985a );
 a5990a <=( a5989a ) or ( a5982a );
 a5991a <=( a5990a ) or ( a5975a );
 a5992a <=( a5991a ) or ( a5962a );
 a5993a <=( a5992a ) or ( a5933a );
 a5994a <=( a5993a ) or ( a5874a );
 a5998a <=( a2757a ) or ( a2758a );
 a5999a <=( a2759a ) or ( a5998a );
 a6002a <=( a2755a ) or ( a2756a );
 a6005a <=( a2753a ) or ( a2754a );
 a6006a <=( a6005a ) or ( a6002a );
 a6007a <=( a6006a ) or ( a5999a );
 a6010a <=( a2751a ) or ( a2752a );
 a6013a <=( a2749a ) or ( a2750a );
 a6014a <=( a6013a ) or ( a6010a );
 a6017a <=( a2747a ) or ( a2748a );
 a6020a <=( a2745a ) or ( a2746a );
 a6021a <=( a6020a ) or ( a6017a );
 a6022a <=( a6021a ) or ( a6014a );
 a6023a <=( a6022a ) or ( a6007a );
 a6027a <=( a2742a ) or ( a2743a );
 a6028a <=( a2744a ) or ( a6027a );
 a6031a <=( a2740a ) or ( a2741a );
 a6034a <=( a2738a ) or ( a2739a );
 a6035a <=( a6034a ) or ( a6031a );
 a6036a <=( a6035a ) or ( a6028a );
 a6039a <=( a2736a ) or ( a2737a );
 a6042a <=( a2734a ) or ( a2735a );
 a6043a <=( a6042a ) or ( a6039a );
 a6046a <=( a2732a ) or ( a2733a );
 a6049a <=( a2730a ) or ( a2731a );
 a6050a <=( a6049a ) or ( a6046a );
 a6051a <=( a6050a ) or ( a6043a );
 a6052a <=( a6051a ) or ( a6036a );
 a6053a <=( a6052a ) or ( a6023a );
 a6057a <=( a2727a ) or ( a2728a );
 a6058a <=( a2729a ) or ( a6057a );
 a6061a <=( a2725a ) or ( a2726a );
 a6064a <=( a2723a ) or ( a2724a );
 a6065a <=( a6064a ) or ( a6061a );
 a6066a <=( a6065a ) or ( a6058a );
 a6069a <=( a2721a ) or ( a2722a );
 a6072a <=( a2719a ) or ( a2720a );
 a6073a <=( a6072a ) or ( a6069a );
 a6076a <=( a2717a ) or ( a2718a );
 a6079a <=( a2715a ) or ( a2716a );
 a6080a <=( a6079a ) or ( a6076a );
 a6081a <=( a6080a ) or ( a6073a );
 a6082a <=( a6081a ) or ( a6066a );
 a6086a <=( a2712a ) or ( a2713a );
 a6087a <=( a2714a ) or ( a6086a );
 a6090a <=( a2710a ) or ( a2711a );
 a6093a <=( a2708a ) or ( a2709a );
 a6094a <=( a6093a ) or ( a6090a );
 a6095a <=( a6094a ) or ( a6087a );
 a6098a <=( a2706a ) or ( a2707a );
 a6101a <=( a2704a ) or ( a2705a );
 a6102a <=( a6101a ) or ( a6098a );
 a6105a <=( a2702a ) or ( a2703a );
 a6108a <=( a2700a ) or ( a2701a );
 a6109a <=( a6108a ) or ( a6105a );
 a6110a <=( a6109a ) or ( a6102a );
 a6111a <=( a6110a ) or ( a6095a );
 a6112a <=( a6111a ) or ( a6082a );
 a6113a <=( a6112a ) or ( a6053a );
 a6117a <=( a2697a ) or ( a2698a );
 a6118a <=( a2699a ) or ( a6117a );
 a6121a <=( a2695a ) or ( a2696a );
 a6124a <=( a2693a ) or ( a2694a );
 a6125a <=( a6124a ) or ( a6121a );
 a6126a <=( a6125a ) or ( a6118a );
 a6129a <=( a2691a ) or ( a2692a );
 a6132a <=( a2689a ) or ( a2690a );
 a6133a <=( a6132a ) or ( a6129a );
 a6136a <=( a2687a ) or ( a2688a );
 a6139a <=( a2685a ) or ( a2686a );
 a6140a <=( a6139a ) or ( a6136a );
 a6141a <=( a6140a ) or ( a6133a );
 a6142a <=( a6141a ) or ( a6126a );
 a6146a <=( a2682a ) or ( a2683a );
 a6147a <=( a2684a ) or ( a6146a );
 a6150a <=( a2680a ) or ( a2681a );
 a6153a <=( a2678a ) or ( a2679a );
 a6154a <=( a6153a ) or ( a6150a );
 a6155a <=( a6154a ) or ( a6147a );
 a6158a <=( a2676a ) or ( a2677a );
 a6161a <=( a2674a ) or ( a2675a );
 a6162a <=( a6161a ) or ( a6158a );
 a6165a <=( a2672a ) or ( a2673a );
 a6168a <=( a2670a ) or ( a2671a );
 a6169a <=( a6168a ) or ( a6165a );
 a6170a <=( a6169a ) or ( a6162a );
 a6171a <=( a6170a ) or ( a6155a );
 a6172a <=( a6171a ) or ( a6142a );
 a6176a <=( a2667a ) or ( a2668a );
 a6177a <=( a2669a ) or ( a6176a );
 a6180a <=( a2665a ) or ( a2666a );
 a6183a <=( a2663a ) or ( a2664a );
 a6184a <=( a6183a ) or ( a6180a );
 a6185a <=( a6184a ) or ( a6177a );
 a6188a <=( a2661a ) or ( a2662a );
 a6191a <=( a2659a ) or ( a2660a );
 a6192a <=( a6191a ) or ( a6188a );
 a6195a <=( a2657a ) or ( a2658a );
 a6198a <=( a2655a ) or ( a2656a );
 a6199a <=( a6198a ) or ( a6195a );
 a6200a <=( a6199a ) or ( a6192a );
 a6201a <=( a6200a ) or ( a6185a );
 a6205a <=( a2652a ) or ( a2653a );
 a6206a <=( a2654a ) or ( a6205a );
 a6209a <=( a2650a ) or ( a2651a );
 a6212a <=( a2648a ) or ( a2649a );
 a6213a <=( a6212a ) or ( a6209a );
 a6214a <=( a6213a ) or ( a6206a );
 a6217a <=( a2646a ) or ( a2647a );
 a6220a <=( a2644a ) or ( a2645a );
 a6221a <=( a6220a ) or ( a6217a );
 a6224a <=( a2642a ) or ( a2643a );
 a6227a <=( a2640a ) or ( a2641a );
 a6228a <=( a6227a ) or ( a6224a );
 a6229a <=( a6228a ) or ( a6221a );
 a6230a <=( a6229a ) or ( a6214a );
 a6231a <=( a6230a ) or ( a6201a );
 a6232a <=( a6231a ) or ( a6172a );
 a6233a <=( a6232a ) or ( a6113a );
 a6234a <=( a6233a ) or ( a5994a );
 a6238a <=( a2637a ) or ( a2638a );
 a6239a <=( a2639a ) or ( a6238a );
 a6242a <=( a2635a ) or ( a2636a );
 a6245a <=( a2633a ) or ( a2634a );
 a6246a <=( a6245a ) or ( a6242a );
 a6247a <=( a6246a ) or ( a6239a );
 a6250a <=( a2631a ) or ( a2632a );
 a6253a <=( a2629a ) or ( a2630a );
 a6254a <=( a6253a ) or ( a6250a );
 a6257a <=( a2627a ) or ( a2628a );
 a6260a <=( a2625a ) or ( a2626a );
 a6261a <=( a6260a ) or ( a6257a );
 a6262a <=( a6261a ) or ( a6254a );
 a6263a <=( a6262a ) or ( a6247a );
 a6267a <=( a2622a ) or ( a2623a );
 a6268a <=( a2624a ) or ( a6267a );
 a6271a <=( a2620a ) or ( a2621a );
 a6274a <=( a2618a ) or ( a2619a );
 a6275a <=( a6274a ) or ( a6271a );
 a6276a <=( a6275a ) or ( a6268a );
 a6279a <=( a2616a ) or ( a2617a );
 a6282a <=( a2614a ) or ( a2615a );
 a6283a <=( a6282a ) or ( a6279a );
 a6286a <=( a2612a ) or ( a2613a );
 a6289a <=( a2610a ) or ( a2611a );
 a6290a <=( a6289a ) or ( a6286a );
 a6291a <=( a6290a ) or ( a6283a );
 a6292a <=( a6291a ) or ( a6276a );
 a6293a <=( a6292a ) or ( a6263a );
 a6297a <=( a2607a ) or ( a2608a );
 a6298a <=( a2609a ) or ( a6297a );
 a6301a <=( a2605a ) or ( a2606a );
 a6304a <=( a2603a ) or ( a2604a );
 a6305a <=( a6304a ) or ( a6301a );
 a6306a <=( a6305a ) or ( a6298a );
 a6309a <=( a2601a ) or ( a2602a );
 a6312a <=( a2599a ) or ( a2600a );
 a6313a <=( a6312a ) or ( a6309a );
 a6316a <=( a2597a ) or ( a2598a );
 a6319a <=( a2595a ) or ( a2596a );
 a6320a <=( a6319a ) or ( a6316a );
 a6321a <=( a6320a ) or ( a6313a );
 a6322a <=( a6321a ) or ( a6306a );
 a6326a <=( a2592a ) or ( a2593a );
 a6327a <=( a2594a ) or ( a6326a );
 a6330a <=( a2590a ) or ( a2591a );
 a6333a <=( a2588a ) or ( a2589a );
 a6334a <=( a6333a ) or ( a6330a );
 a6335a <=( a6334a ) or ( a6327a );
 a6338a <=( a2586a ) or ( a2587a );
 a6341a <=( a2584a ) or ( a2585a );
 a6342a <=( a6341a ) or ( a6338a );
 a6345a <=( a2582a ) or ( a2583a );
 a6348a <=( a2580a ) or ( a2581a );
 a6349a <=( a6348a ) or ( a6345a );
 a6350a <=( a6349a ) or ( a6342a );
 a6351a <=( a6350a ) or ( a6335a );
 a6352a <=( a6351a ) or ( a6322a );
 a6353a <=( a6352a ) or ( a6293a );
 a6357a <=( a2577a ) or ( a2578a );
 a6358a <=( a2579a ) or ( a6357a );
 a6361a <=( a2575a ) or ( a2576a );
 a6364a <=( a2573a ) or ( a2574a );
 a6365a <=( a6364a ) or ( a6361a );
 a6366a <=( a6365a ) or ( a6358a );
 a6369a <=( a2571a ) or ( a2572a );
 a6372a <=( a2569a ) or ( a2570a );
 a6373a <=( a6372a ) or ( a6369a );
 a6376a <=( a2567a ) or ( a2568a );
 a6379a <=( a2565a ) or ( a2566a );
 a6380a <=( a6379a ) or ( a6376a );
 a6381a <=( a6380a ) or ( a6373a );
 a6382a <=( a6381a ) or ( a6366a );
 a6386a <=( a2562a ) or ( a2563a );
 a6387a <=( a2564a ) or ( a6386a );
 a6390a <=( a2560a ) or ( a2561a );
 a6393a <=( a2558a ) or ( a2559a );
 a6394a <=( a6393a ) or ( a6390a );
 a6395a <=( a6394a ) or ( a6387a );
 a6398a <=( a2556a ) or ( a2557a );
 a6401a <=( a2554a ) or ( a2555a );
 a6402a <=( a6401a ) or ( a6398a );
 a6405a <=( a2552a ) or ( a2553a );
 a6408a <=( a2550a ) or ( a2551a );
 a6409a <=( a6408a ) or ( a6405a );
 a6410a <=( a6409a ) or ( a6402a );
 a6411a <=( a6410a ) or ( a6395a );
 a6412a <=( a6411a ) or ( a6382a );
 a6416a <=( a2547a ) or ( a2548a );
 a6417a <=( a2549a ) or ( a6416a );
 a6420a <=( a2545a ) or ( a2546a );
 a6423a <=( a2543a ) or ( a2544a );
 a6424a <=( a6423a ) or ( a6420a );
 a6425a <=( a6424a ) or ( a6417a );
 a6428a <=( a2541a ) or ( a2542a );
 a6431a <=( a2539a ) or ( a2540a );
 a6432a <=( a6431a ) or ( a6428a );
 a6435a <=( a2537a ) or ( a2538a );
 a6438a <=( a2535a ) or ( a2536a );
 a6439a <=( a6438a ) or ( a6435a );
 a6440a <=( a6439a ) or ( a6432a );
 a6441a <=( a6440a ) or ( a6425a );
 a6445a <=( a2532a ) or ( a2533a );
 a6446a <=( a2534a ) or ( a6445a );
 a6449a <=( a2530a ) or ( a2531a );
 a6452a <=( a2528a ) or ( a2529a );
 a6453a <=( a6452a ) or ( a6449a );
 a6454a <=( a6453a ) or ( a6446a );
 a6457a <=( a2526a ) or ( a2527a );
 a6460a <=( a2524a ) or ( a2525a );
 a6461a <=( a6460a ) or ( a6457a );
 a6464a <=( a2522a ) or ( a2523a );
 a6467a <=( a2520a ) or ( a2521a );
 a6468a <=( a6467a ) or ( a6464a );
 a6469a <=( a6468a ) or ( a6461a );
 a6470a <=( a6469a ) or ( a6454a );
 a6471a <=( a6470a ) or ( a6441a );
 a6472a <=( a6471a ) or ( a6412a );
 a6473a <=( a6472a ) or ( a6353a );
 a6477a <=( a2517a ) or ( a2518a );
 a6478a <=( a2519a ) or ( a6477a );
 a6481a <=( a2515a ) or ( a2516a );
 a6484a <=( a2513a ) or ( a2514a );
 a6485a <=( a6484a ) or ( a6481a );
 a6486a <=( a6485a ) or ( a6478a );
 a6489a <=( a2511a ) or ( a2512a );
 a6492a <=( a2509a ) or ( a2510a );
 a6493a <=( a6492a ) or ( a6489a );
 a6496a <=( a2507a ) or ( a2508a );
 a6499a <=( a2505a ) or ( a2506a );
 a6500a <=( a6499a ) or ( a6496a );
 a6501a <=( a6500a ) or ( a6493a );
 a6502a <=( a6501a ) or ( a6486a );
 a6506a <=( a2502a ) or ( a2503a );
 a6507a <=( a2504a ) or ( a6506a );
 a6510a <=( a2500a ) or ( a2501a );
 a6513a <=( a2498a ) or ( a2499a );
 a6514a <=( a6513a ) or ( a6510a );
 a6515a <=( a6514a ) or ( a6507a );
 a6518a <=( a2496a ) or ( a2497a );
 a6521a <=( a2494a ) or ( a2495a );
 a6522a <=( a6521a ) or ( a6518a );
 a6525a <=( a2492a ) or ( a2493a );
 a6528a <=( a2490a ) or ( a2491a );
 a6529a <=( a6528a ) or ( a6525a );
 a6530a <=( a6529a ) or ( a6522a );
 a6531a <=( a6530a ) or ( a6515a );
 a6532a <=( a6531a ) or ( a6502a );
 a6536a <=( a2487a ) or ( a2488a );
 a6537a <=( a2489a ) or ( a6536a );
 a6540a <=( a2485a ) or ( a2486a );
 a6543a <=( a2483a ) or ( a2484a );
 a6544a <=( a6543a ) or ( a6540a );
 a6545a <=( a6544a ) or ( a6537a );
 a6548a <=( a2481a ) or ( a2482a );
 a6551a <=( a2479a ) or ( a2480a );
 a6552a <=( a6551a ) or ( a6548a );
 a6555a <=( a2477a ) or ( a2478a );
 a6558a <=( a2475a ) or ( a2476a );
 a6559a <=( a6558a ) or ( a6555a );
 a6560a <=( a6559a ) or ( a6552a );
 a6561a <=( a6560a ) or ( a6545a );
 a6565a <=( a2472a ) or ( a2473a );
 a6566a <=( a2474a ) or ( a6565a );
 a6569a <=( a2470a ) or ( a2471a );
 a6572a <=( a2468a ) or ( a2469a );
 a6573a <=( a6572a ) or ( a6569a );
 a6574a <=( a6573a ) or ( a6566a );
 a6577a <=( a2466a ) or ( a2467a );
 a6580a <=( a2464a ) or ( a2465a );
 a6581a <=( a6580a ) or ( a6577a );
 a6584a <=( a2462a ) or ( a2463a );
 a6587a <=( a2460a ) or ( a2461a );
 a6588a <=( a6587a ) or ( a6584a );
 a6589a <=( a6588a ) or ( a6581a );
 a6590a <=( a6589a ) or ( a6574a );
 a6591a <=( a6590a ) or ( a6561a );
 a6592a <=( a6591a ) or ( a6532a );
 a6596a <=( a2457a ) or ( a2458a );
 a6597a <=( a2459a ) or ( a6596a );
 a6600a <=( a2455a ) or ( a2456a );
 a6603a <=( a2453a ) or ( a2454a );
 a6604a <=( a6603a ) or ( a6600a );
 a6605a <=( a6604a ) or ( a6597a );
 a6608a <=( a2451a ) or ( a2452a );
 a6611a <=( a2449a ) or ( a2450a );
 a6612a <=( a6611a ) or ( a6608a );
 a6615a <=( a2447a ) or ( a2448a );
 a6618a <=( a2445a ) or ( a2446a );
 a6619a <=( a6618a ) or ( a6615a );
 a6620a <=( a6619a ) or ( a6612a );
 a6621a <=( a6620a ) or ( a6605a );
 a6625a <=( a2442a ) or ( a2443a );
 a6626a <=( a2444a ) or ( a6625a );
 a6629a <=( a2440a ) or ( a2441a );
 a6632a <=( a2438a ) or ( a2439a );
 a6633a <=( a6632a ) or ( a6629a );
 a6634a <=( a6633a ) or ( a6626a );
 a6637a <=( a2436a ) or ( a2437a );
 a6640a <=( a2434a ) or ( a2435a );
 a6641a <=( a6640a ) or ( a6637a );
 a6644a <=( a2432a ) or ( a2433a );
 a6647a <=( a2430a ) or ( a2431a );
 a6648a <=( a6647a ) or ( a6644a );
 a6649a <=( a6648a ) or ( a6641a );
 a6650a <=( a6649a ) or ( a6634a );
 a6651a <=( a6650a ) or ( a6621a );
 a6655a <=( a2427a ) or ( a2428a );
 a6656a <=( a2429a ) or ( a6655a );
 a6659a <=( a2425a ) or ( a2426a );
 a6662a <=( a2423a ) or ( a2424a );
 a6663a <=( a6662a ) or ( a6659a );
 a6664a <=( a6663a ) or ( a6656a );
 a6667a <=( a2421a ) or ( a2422a );
 a6670a <=( a2419a ) or ( a2420a );
 a6671a <=( a6670a ) or ( a6667a );
 a6674a <=( a2417a ) or ( a2418a );
 a6677a <=( a2415a ) or ( a2416a );
 a6678a <=( a6677a ) or ( a6674a );
 a6679a <=( a6678a ) or ( a6671a );
 a6680a <=( a6679a ) or ( a6664a );
 a6684a <=( a2412a ) or ( a2413a );
 a6685a <=( a2414a ) or ( a6684a );
 a6688a <=( a2410a ) or ( a2411a );
 a6691a <=( a2408a ) or ( a2409a );
 a6692a <=( a6691a ) or ( a6688a );
 a6693a <=( a6692a ) or ( a6685a );
 a6696a <=( a2406a ) or ( a2407a );
 a6699a <=( a2404a ) or ( a2405a );
 a6700a <=( a6699a ) or ( a6696a );
 a6703a <=( a2402a ) or ( a2403a );
 a6706a <=( a2400a ) or ( a2401a );
 a6707a <=( a6706a ) or ( a6703a );
 a6708a <=( a6707a ) or ( a6700a );
 a6709a <=( a6708a ) or ( a6693a );
 a6710a <=( a6709a ) or ( a6680a );
 a6711a <=( a6710a ) or ( a6651a );
 a6712a <=( a6711a ) or ( a6592a );
 a6713a <=( a6712a ) or ( a6473a );
 a6714a <=( a6713a ) or ( a6234a );
 a6718a <=( a2397a ) or ( a2398a );
 a6719a <=( a2399a ) or ( a6718a );
 a6722a <=( a2395a ) or ( a2396a );
 a6725a <=( a2393a ) or ( a2394a );
 a6726a <=( a6725a ) or ( a6722a );
 a6727a <=( a6726a ) or ( a6719a );
 a6730a <=( a2391a ) or ( a2392a );
 a6733a <=( a2389a ) or ( a2390a );
 a6734a <=( a6733a ) or ( a6730a );
 a6737a <=( a2387a ) or ( a2388a );
 a6740a <=( a2385a ) or ( a2386a );
 a6741a <=( a6740a ) or ( a6737a );
 a6742a <=( a6741a ) or ( a6734a );
 a6743a <=( a6742a ) or ( a6727a );
 a6747a <=( a2382a ) or ( a2383a );
 a6748a <=( a2384a ) or ( a6747a );
 a6751a <=( a2380a ) or ( a2381a );
 a6754a <=( a2378a ) or ( a2379a );
 a6755a <=( a6754a ) or ( a6751a );
 a6756a <=( a6755a ) or ( a6748a );
 a6759a <=( a2376a ) or ( a2377a );
 a6762a <=( a2374a ) or ( a2375a );
 a6763a <=( a6762a ) or ( a6759a );
 a6766a <=( a2372a ) or ( a2373a );
 a6769a <=( a2370a ) or ( a2371a );
 a6770a <=( a6769a ) or ( a6766a );
 a6771a <=( a6770a ) or ( a6763a );
 a6772a <=( a6771a ) or ( a6756a );
 a6773a <=( a6772a ) or ( a6743a );
 a6777a <=( a2367a ) or ( a2368a );
 a6778a <=( a2369a ) or ( a6777a );
 a6781a <=( a2365a ) or ( a2366a );
 a6784a <=( a2363a ) or ( a2364a );
 a6785a <=( a6784a ) or ( a6781a );
 a6786a <=( a6785a ) or ( a6778a );
 a6789a <=( a2361a ) or ( a2362a );
 a6792a <=( a2359a ) or ( a2360a );
 a6793a <=( a6792a ) or ( a6789a );
 a6796a <=( a2357a ) or ( a2358a );
 a6799a <=( a2355a ) or ( a2356a );
 a6800a <=( a6799a ) or ( a6796a );
 a6801a <=( a6800a ) or ( a6793a );
 a6802a <=( a6801a ) or ( a6786a );
 a6806a <=( a2352a ) or ( a2353a );
 a6807a <=( a2354a ) or ( a6806a );
 a6810a <=( a2350a ) or ( a2351a );
 a6813a <=( a2348a ) or ( a2349a );
 a6814a <=( a6813a ) or ( a6810a );
 a6815a <=( a6814a ) or ( a6807a );
 a6818a <=( a2346a ) or ( a2347a );
 a6821a <=( a2344a ) or ( a2345a );
 a6822a <=( a6821a ) or ( a6818a );
 a6825a <=( a2342a ) or ( a2343a );
 a6828a <=( a2340a ) or ( a2341a );
 a6829a <=( a6828a ) or ( a6825a );
 a6830a <=( a6829a ) or ( a6822a );
 a6831a <=( a6830a ) or ( a6815a );
 a6832a <=( a6831a ) or ( a6802a );
 a6833a <=( a6832a ) or ( a6773a );
 a6837a <=( a2337a ) or ( a2338a );
 a6838a <=( a2339a ) or ( a6837a );
 a6841a <=( a2335a ) or ( a2336a );
 a6844a <=( a2333a ) or ( a2334a );
 a6845a <=( a6844a ) or ( a6841a );
 a6846a <=( a6845a ) or ( a6838a );
 a6849a <=( a2331a ) or ( a2332a );
 a6852a <=( a2329a ) or ( a2330a );
 a6853a <=( a6852a ) or ( a6849a );
 a6856a <=( a2327a ) or ( a2328a );
 a6859a <=( a2325a ) or ( a2326a );
 a6860a <=( a6859a ) or ( a6856a );
 a6861a <=( a6860a ) or ( a6853a );
 a6862a <=( a6861a ) or ( a6846a );
 a6866a <=( a2322a ) or ( a2323a );
 a6867a <=( a2324a ) or ( a6866a );
 a6870a <=( a2320a ) or ( a2321a );
 a6873a <=( a2318a ) or ( a2319a );
 a6874a <=( a6873a ) or ( a6870a );
 a6875a <=( a6874a ) or ( a6867a );
 a6878a <=( a2316a ) or ( a2317a );
 a6881a <=( a2314a ) or ( a2315a );
 a6882a <=( a6881a ) or ( a6878a );
 a6885a <=( a2312a ) or ( a2313a );
 a6888a <=( a2310a ) or ( a2311a );
 a6889a <=( a6888a ) or ( a6885a );
 a6890a <=( a6889a ) or ( a6882a );
 a6891a <=( a6890a ) or ( a6875a );
 a6892a <=( a6891a ) or ( a6862a );
 a6896a <=( a2307a ) or ( a2308a );
 a6897a <=( a2309a ) or ( a6896a );
 a6900a <=( a2305a ) or ( a2306a );
 a6903a <=( a2303a ) or ( a2304a );
 a6904a <=( a6903a ) or ( a6900a );
 a6905a <=( a6904a ) or ( a6897a );
 a6908a <=( a2301a ) or ( a2302a );
 a6911a <=( a2299a ) or ( a2300a );
 a6912a <=( a6911a ) or ( a6908a );
 a6915a <=( a2297a ) or ( a2298a );
 a6918a <=( a2295a ) or ( a2296a );
 a6919a <=( a6918a ) or ( a6915a );
 a6920a <=( a6919a ) or ( a6912a );
 a6921a <=( a6920a ) or ( a6905a );
 a6925a <=( a2292a ) or ( a2293a );
 a6926a <=( a2294a ) or ( a6925a );
 a6929a <=( a2290a ) or ( a2291a );
 a6932a <=( a2288a ) or ( a2289a );
 a6933a <=( a6932a ) or ( a6929a );
 a6934a <=( a6933a ) or ( a6926a );
 a6937a <=( a2286a ) or ( a2287a );
 a6940a <=( a2284a ) or ( a2285a );
 a6941a <=( a6940a ) or ( a6937a );
 a6944a <=( a2282a ) or ( a2283a );
 a6947a <=( a2280a ) or ( a2281a );
 a6948a <=( a6947a ) or ( a6944a );
 a6949a <=( a6948a ) or ( a6941a );
 a6950a <=( a6949a ) or ( a6934a );
 a6951a <=( a6950a ) or ( a6921a );
 a6952a <=( a6951a ) or ( a6892a );
 a6953a <=( a6952a ) or ( a6833a );
 a6957a <=( a2277a ) or ( a2278a );
 a6958a <=( a2279a ) or ( a6957a );
 a6961a <=( a2275a ) or ( a2276a );
 a6964a <=( a2273a ) or ( a2274a );
 a6965a <=( a6964a ) or ( a6961a );
 a6966a <=( a6965a ) or ( a6958a );
 a6969a <=( a2271a ) or ( a2272a );
 a6972a <=( a2269a ) or ( a2270a );
 a6973a <=( a6972a ) or ( a6969a );
 a6976a <=( a2267a ) or ( a2268a );
 a6979a <=( a2265a ) or ( a2266a );
 a6980a <=( a6979a ) or ( a6976a );
 a6981a <=( a6980a ) or ( a6973a );
 a6982a <=( a6981a ) or ( a6966a );
 a6986a <=( a2262a ) or ( a2263a );
 a6987a <=( a2264a ) or ( a6986a );
 a6990a <=( a2260a ) or ( a2261a );
 a6993a <=( a2258a ) or ( a2259a );
 a6994a <=( a6993a ) or ( a6990a );
 a6995a <=( a6994a ) or ( a6987a );
 a6998a <=( a2256a ) or ( a2257a );
 a7001a <=( a2254a ) or ( a2255a );
 a7002a <=( a7001a ) or ( a6998a );
 a7005a <=( a2252a ) or ( a2253a );
 a7008a <=( a2250a ) or ( a2251a );
 a7009a <=( a7008a ) or ( a7005a );
 a7010a <=( a7009a ) or ( a7002a );
 a7011a <=( a7010a ) or ( a6995a );
 a7012a <=( a7011a ) or ( a6982a );
 a7016a <=( a2247a ) or ( a2248a );
 a7017a <=( a2249a ) or ( a7016a );
 a7020a <=( a2245a ) or ( a2246a );
 a7023a <=( a2243a ) or ( a2244a );
 a7024a <=( a7023a ) or ( a7020a );
 a7025a <=( a7024a ) or ( a7017a );
 a7028a <=( a2241a ) or ( a2242a );
 a7031a <=( a2239a ) or ( a2240a );
 a7032a <=( a7031a ) or ( a7028a );
 a7035a <=( a2237a ) or ( a2238a );
 a7038a <=( a2235a ) or ( a2236a );
 a7039a <=( a7038a ) or ( a7035a );
 a7040a <=( a7039a ) or ( a7032a );
 a7041a <=( a7040a ) or ( a7025a );
 a7045a <=( a2232a ) or ( a2233a );
 a7046a <=( a2234a ) or ( a7045a );
 a7049a <=( a2230a ) or ( a2231a );
 a7052a <=( a2228a ) or ( a2229a );
 a7053a <=( a7052a ) or ( a7049a );
 a7054a <=( a7053a ) or ( a7046a );
 a7057a <=( a2226a ) or ( a2227a );
 a7060a <=( a2224a ) or ( a2225a );
 a7061a <=( a7060a ) or ( a7057a );
 a7064a <=( a2222a ) or ( a2223a );
 a7067a <=( a2220a ) or ( a2221a );
 a7068a <=( a7067a ) or ( a7064a );
 a7069a <=( a7068a ) or ( a7061a );
 a7070a <=( a7069a ) or ( a7054a );
 a7071a <=( a7070a ) or ( a7041a );
 a7072a <=( a7071a ) or ( a7012a );
 a7076a <=( a2217a ) or ( a2218a );
 a7077a <=( a2219a ) or ( a7076a );
 a7080a <=( a2215a ) or ( a2216a );
 a7083a <=( a2213a ) or ( a2214a );
 a7084a <=( a7083a ) or ( a7080a );
 a7085a <=( a7084a ) or ( a7077a );
 a7088a <=( a2211a ) or ( a2212a );
 a7091a <=( a2209a ) or ( a2210a );
 a7092a <=( a7091a ) or ( a7088a );
 a7095a <=( a2207a ) or ( a2208a );
 a7098a <=( a2205a ) or ( a2206a );
 a7099a <=( a7098a ) or ( a7095a );
 a7100a <=( a7099a ) or ( a7092a );
 a7101a <=( a7100a ) or ( a7085a );
 a7105a <=( a2202a ) or ( a2203a );
 a7106a <=( a2204a ) or ( a7105a );
 a7109a <=( a2200a ) or ( a2201a );
 a7112a <=( a2198a ) or ( a2199a );
 a7113a <=( a7112a ) or ( a7109a );
 a7114a <=( a7113a ) or ( a7106a );
 a7117a <=( a2196a ) or ( a2197a );
 a7120a <=( a2194a ) or ( a2195a );
 a7121a <=( a7120a ) or ( a7117a );
 a7124a <=( a2192a ) or ( a2193a );
 a7127a <=( a2190a ) or ( a2191a );
 a7128a <=( a7127a ) or ( a7124a );
 a7129a <=( a7128a ) or ( a7121a );
 a7130a <=( a7129a ) or ( a7114a );
 a7131a <=( a7130a ) or ( a7101a );
 a7135a <=( a2187a ) or ( a2188a );
 a7136a <=( a2189a ) or ( a7135a );
 a7139a <=( a2185a ) or ( a2186a );
 a7142a <=( a2183a ) or ( a2184a );
 a7143a <=( a7142a ) or ( a7139a );
 a7144a <=( a7143a ) or ( a7136a );
 a7147a <=( a2181a ) or ( a2182a );
 a7150a <=( a2179a ) or ( a2180a );
 a7151a <=( a7150a ) or ( a7147a );
 a7154a <=( a2177a ) or ( a2178a );
 a7157a <=( a2175a ) or ( a2176a );
 a7158a <=( a7157a ) or ( a7154a );
 a7159a <=( a7158a ) or ( a7151a );
 a7160a <=( a7159a ) or ( a7144a );
 a7164a <=( a2172a ) or ( a2173a );
 a7165a <=( a2174a ) or ( a7164a );
 a7168a <=( a2170a ) or ( a2171a );
 a7171a <=( a2168a ) or ( a2169a );
 a7172a <=( a7171a ) or ( a7168a );
 a7173a <=( a7172a ) or ( a7165a );
 a7176a <=( a2166a ) or ( a2167a );
 a7179a <=( a2164a ) or ( a2165a );
 a7180a <=( a7179a ) or ( a7176a );
 a7183a <=( a2162a ) or ( a2163a );
 a7186a <=( a2160a ) or ( a2161a );
 a7187a <=( a7186a ) or ( a7183a );
 a7188a <=( a7187a ) or ( a7180a );
 a7189a <=( a7188a ) or ( a7173a );
 a7190a <=( a7189a ) or ( a7160a );
 a7191a <=( a7190a ) or ( a7131a );
 a7192a <=( a7191a ) or ( a7072a );
 a7193a <=( a7192a ) or ( a6953a );
 a7197a <=( a2157a ) or ( a2158a );
 a7198a <=( a2159a ) or ( a7197a );
 a7201a <=( a2155a ) or ( a2156a );
 a7204a <=( a2153a ) or ( a2154a );
 a7205a <=( a7204a ) or ( a7201a );
 a7206a <=( a7205a ) or ( a7198a );
 a7209a <=( a2151a ) or ( a2152a );
 a7212a <=( a2149a ) or ( a2150a );
 a7213a <=( a7212a ) or ( a7209a );
 a7216a <=( a2147a ) or ( a2148a );
 a7219a <=( a2145a ) or ( a2146a );
 a7220a <=( a7219a ) or ( a7216a );
 a7221a <=( a7220a ) or ( a7213a );
 a7222a <=( a7221a ) or ( a7206a );
 a7226a <=( a2142a ) or ( a2143a );
 a7227a <=( a2144a ) or ( a7226a );
 a7230a <=( a2140a ) or ( a2141a );
 a7233a <=( a2138a ) or ( a2139a );
 a7234a <=( a7233a ) or ( a7230a );
 a7235a <=( a7234a ) or ( a7227a );
 a7238a <=( a2136a ) or ( a2137a );
 a7241a <=( a2134a ) or ( a2135a );
 a7242a <=( a7241a ) or ( a7238a );
 a7245a <=( a2132a ) or ( a2133a );
 a7248a <=( a2130a ) or ( a2131a );
 a7249a <=( a7248a ) or ( a7245a );
 a7250a <=( a7249a ) or ( a7242a );
 a7251a <=( a7250a ) or ( a7235a );
 a7252a <=( a7251a ) or ( a7222a );
 a7256a <=( a2127a ) or ( a2128a );
 a7257a <=( a2129a ) or ( a7256a );
 a7260a <=( a2125a ) or ( a2126a );
 a7263a <=( a2123a ) or ( a2124a );
 a7264a <=( a7263a ) or ( a7260a );
 a7265a <=( a7264a ) or ( a7257a );
 a7268a <=( a2121a ) or ( a2122a );
 a7271a <=( a2119a ) or ( a2120a );
 a7272a <=( a7271a ) or ( a7268a );
 a7275a <=( a2117a ) or ( a2118a );
 a7278a <=( a2115a ) or ( a2116a );
 a7279a <=( a7278a ) or ( a7275a );
 a7280a <=( a7279a ) or ( a7272a );
 a7281a <=( a7280a ) or ( a7265a );
 a7285a <=( a2112a ) or ( a2113a );
 a7286a <=( a2114a ) or ( a7285a );
 a7289a <=( a2110a ) or ( a2111a );
 a7292a <=( a2108a ) or ( a2109a );
 a7293a <=( a7292a ) or ( a7289a );
 a7294a <=( a7293a ) or ( a7286a );
 a7297a <=( a2106a ) or ( a2107a );
 a7300a <=( a2104a ) or ( a2105a );
 a7301a <=( a7300a ) or ( a7297a );
 a7304a <=( a2102a ) or ( a2103a );
 a7307a <=( a2100a ) or ( a2101a );
 a7308a <=( a7307a ) or ( a7304a );
 a7309a <=( a7308a ) or ( a7301a );
 a7310a <=( a7309a ) or ( a7294a );
 a7311a <=( a7310a ) or ( a7281a );
 a7312a <=( a7311a ) or ( a7252a );
 a7316a <=( a2097a ) or ( a2098a );
 a7317a <=( a2099a ) or ( a7316a );
 a7320a <=( a2095a ) or ( a2096a );
 a7323a <=( a2093a ) or ( a2094a );
 a7324a <=( a7323a ) or ( a7320a );
 a7325a <=( a7324a ) or ( a7317a );
 a7328a <=( a2091a ) or ( a2092a );
 a7331a <=( a2089a ) or ( a2090a );
 a7332a <=( a7331a ) or ( a7328a );
 a7335a <=( a2087a ) or ( a2088a );
 a7338a <=( a2085a ) or ( a2086a );
 a7339a <=( a7338a ) or ( a7335a );
 a7340a <=( a7339a ) or ( a7332a );
 a7341a <=( a7340a ) or ( a7325a );
 a7345a <=( a2082a ) or ( a2083a );
 a7346a <=( a2084a ) or ( a7345a );
 a7349a <=( a2080a ) or ( a2081a );
 a7352a <=( a2078a ) or ( a2079a );
 a7353a <=( a7352a ) or ( a7349a );
 a7354a <=( a7353a ) or ( a7346a );
 a7357a <=( a2076a ) or ( a2077a );
 a7360a <=( a2074a ) or ( a2075a );
 a7361a <=( a7360a ) or ( a7357a );
 a7364a <=( a2072a ) or ( a2073a );
 a7367a <=( a2070a ) or ( a2071a );
 a7368a <=( a7367a ) or ( a7364a );
 a7369a <=( a7368a ) or ( a7361a );
 a7370a <=( a7369a ) or ( a7354a );
 a7371a <=( a7370a ) or ( a7341a );
 a7375a <=( a2067a ) or ( a2068a );
 a7376a <=( a2069a ) or ( a7375a );
 a7379a <=( a2065a ) or ( a2066a );
 a7382a <=( a2063a ) or ( a2064a );
 a7383a <=( a7382a ) or ( a7379a );
 a7384a <=( a7383a ) or ( a7376a );
 a7387a <=( a2061a ) or ( a2062a );
 a7390a <=( a2059a ) or ( a2060a );
 a7391a <=( a7390a ) or ( a7387a );
 a7394a <=( a2057a ) or ( a2058a );
 a7397a <=( a2055a ) or ( a2056a );
 a7398a <=( a7397a ) or ( a7394a );
 a7399a <=( a7398a ) or ( a7391a );
 a7400a <=( a7399a ) or ( a7384a );
 a7404a <=( a2052a ) or ( a2053a );
 a7405a <=( a2054a ) or ( a7404a );
 a7408a <=( a2050a ) or ( a2051a );
 a7411a <=( a2048a ) or ( a2049a );
 a7412a <=( a7411a ) or ( a7408a );
 a7413a <=( a7412a ) or ( a7405a );
 a7416a <=( a2046a ) or ( a2047a );
 a7419a <=( a2044a ) or ( a2045a );
 a7420a <=( a7419a ) or ( a7416a );
 a7423a <=( a2042a ) or ( a2043a );
 a7426a <=( a2040a ) or ( a2041a );
 a7427a <=( a7426a ) or ( a7423a );
 a7428a <=( a7427a ) or ( a7420a );
 a7429a <=( a7428a ) or ( a7413a );
 a7430a <=( a7429a ) or ( a7400a );
 a7431a <=( a7430a ) or ( a7371a );
 a7432a <=( a7431a ) or ( a7312a );
 a7436a <=( a2037a ) or ( a2038a );
 a7437a <=( a2039a ) or ( a7436a );
 a7440a <=( a2035a ) or ( a2036a );
 a7443a <=( a2033a ) or ( a2034a );
 a7444a <=( a7443a ) or ( a7440a );
 a7445a <=( a7444a ) or ( a7437a );
 a7448a <=( a2031a ) or ( a2032a );
 a7451a <=( a2029a ) or ( a2030a );
 a7452a <=( a7451a ) or ( a7448a );
 a7455a <=( a2027a ) or ( a2028a );
 a7458a <=( a2025a ) or ( a2026a );
 a7459a <=( a7458a ) or ( a7455a );
 a7460a <=( a7459a ) or ( a7452a );
 a7461a <=( a7460a ) or ( a7445a );
 a7465a <=( a2022a ) or ( a2023a );
 a7466a <=( a2024a ) or ( a7465a );
 a7469a <=( a2020a ) or ( a2021a );
 a7472a <=( a2018a ) or ( a2019a );
 a7473a <=( a7472a ) or ( a7469a );
 a7474a <=( a7473a ) or ( a7466a );
 a7477a <=( a2016a ) or ( a2017a );
 a7480a <=( a2014a ) or ( a2015a );
 a7481a <=( a7480a ) or ( a7477a );
 a7484a <=( a2012a ) or ( a2013a );
 a7487a <=( a2010a ) or ( a2011a );
 a7488a <=( a7487a ) or ( a7484a );
 a7489a <=( a7488a ) or ( a7481a );
 a7490a <=( a7489a ) or ( a7474a );
 a7491a <=( a7490a ) or ( a7461a );
 a7495a <=( a2007a ) or ( a2008a );
 a7496a <=( a2009a ) or ( a7495a );
 a7499a <=( a2005a ) or ( a2006a );
 a7502a <=( a2003a ) or ( a2004a );
 a7503a <=( a7502a ) or ( a7499a );
 a7504a <=( a7503a ) or ( a7496a );
 a7507a <=( a2001a ) or ( a2002a );
 a7510a <=( a1999a ) or ( a2000a );
 a7511a <=( a7510a ) or ( a7507a );
 a7514a <=( a1997a ) or ( a1998a );
 a7517a <=( a1995a ) or ( a1996a );
 a7518a <=( a7517a ) or ( a7514a );
 a7519a <=( a7518a ) or ( a7511a );
 a7520a <=( a7519a ) or ( a7504a );
 a7524a <=( a1992a ) or ( a1993a );
 a7525a <=( a1994a ) or ( a7524a );
 a7528a <=( a1990a ) or ( a1991a );
 a7531a <=( a1988a ) or ( a1989a );
 a7532a <=( a7531a ) or ( a7528a );
 a7533a <=( a7532a ) or ( a7525a );
 a7536a <=( a1986a ) or ( a1987a );
 a7539a <=( a1984a ) or ( a1985a );
 a7540a <=( a7539a ) or ( a7536a );
 a7543a <=( a1982a ) or ( a1983a );
 a7546a <=( a1980a ) or ( a1981a );
 a7547a <=( a7546a ) or ( a7543a );
 a7548a <=( a7547a ) or ( a7540a );
 a7549a <=( a7548a ) or ( a7533a );
 a7550a <=( a7549a ) or ( a7520a );
 a7551a <=( a7550a ) or ( a7491a );
 a7555a <=( a1977a ) or ( a1978a );
 a7556a <=( a1979a ) or ( a7555a );
 a7559a <=( a1975a ) or ( a1976a );
 a7562a <=( a1973a ) or ( a1974a );
 a7563a <=( a7562a ) or ( a7559a );
 a7564a <=( a7563a ) or ( a7556a );
 a7567a <=( a1971a ) or ( a1972a );
 a7570a <=( a1969a ) or ( a1970a );
 a7571a <=( a7570a ) or ( a7567a );
 a7574a <=( a1967a ) or ( a1968a );
 a7577a <=( a1965a ) or ( a1966a );
 a7578a <=( a7577a ) or ( a7574a );
 a7579a <=( a7578a ) or ( a7571a );
 a7580a <=( a7579a ) or ( a7564a );
 a7584a <=( a1962a ) or ( a1963a );
 a7585a <=( a1964a ) or ( a7584a );
 a7588a <=( a1960a ) or ( a1961a );
 a7591a <=( a1958a ) or ( a1959a );
 a7592a <=( a7591a ) or ( a7588a );
 a7593a <=( a7592a ) or ( a7585a );
 a7596a <=( a1956a ) or ( a1957a );
 a7599a <=( a1954a ) or ( a1955a );
 a7600a <=( a7599a ) or ( a7596a );
 a7603a <=( a1952a ) or ( a1953a );
 a7606a <=( a1950a ) or ( a1951a );
 a7607a <=( a7606a ) or ( a7603a );
 a7608a <=( a7607a ) or ( a7600a );
 a7609a <=( a7608a ) or ( a7593a );
 a7610a <=( a7609a ) or ( a7580a );
 a7614a <=( a1947a ) or ( a1948a );
 a7615a <=( a1949a ) or ( a7614a );
 a7618a <=( a1945a ) or ( a1946a );
 a7621a <=( a1943a ) or ( a1944a );
 a7622a <=( a7621a ) or ( a7618a );
 a7623a <=( a7622a ) or ( a7615a );
 a7626a <=( a1941a ) or ( a1942a );
 a7629a <=( a1939a ) or ( a1940a );
 a7630a <=( a7629a ) or ( a7626a );
 a7633a <=( a1937a ) or ( a1938a );
 a7636a <=( a1935a ) or ( a1936a );
 a7637a <=( a7636a ) or ( a7633a );
 a7638a <=( a7637a ) or ( a7630a );
 a7639a <=( a7638a ) or ( a7623a );
 a7643a <=( a1932a ) or ( a1933a );
 a7644a <=( a1934a ) or ( a7643a );
 a7647a <=( a1930a ) or ( a1931a );
 a7650a <=( a1928a ) or ( a1929a );
 a7651a <=( a7650a ) or ( a7647a );
 a7652a <=( a7651a ) or ( a7644a );
 a7655a <=( a1926a ) or ( a1927a );
 a7658a <=( a1924a ) or ( a1925a );
 a7659a <=( a7658a ) or ( a7655a );
 a7662a <=( a1922a ) or ( a1923a );
 a7665a <=( a1920a ) or ( a1921a );
 a7666a <=( a7665a ) or ( a7662a );
 a7667a <=( a7666a ) or ( a7659a );
 a7668a <=( a7667a ) or ( a7652a );
 a7669a <=( a7668a ) or ( a7639a );
 a7670a <=( a7669a ) or ( a7610a );
 a7671a <=( a7670a ) or ( a7551a );
 a7672a <=( a7671a ) or ( a7432a );
 a7673a <=( a7672a ) or ( a7193a );
 a7674a <=( a7673a ) or ( a6714a );
 a7675a <=( a7674a ) or ( a5755a );
 a7679a <=( a1917a ) or ( a1918a );
 a7680a <=( a1919a ) or ( a7679a );
 a7683a <=( a1915a ) or ( a1916a );
 a7686a <=( a1913a ) or ( a1914a );
 a7687a <=( a7686a ) or ( a7683a );
 a7688a <=( a7687a ) or ( a7680a );
 a7692a <=( a1910a ) or ( a1911a );
 a7693a <=( a1912a ) or ( a7692a );
 a7696a <=( a1908a ) or ( a1909a );
 a7699a <=( a1906a ) or ( a1907a );
 a7700a <=( a7699a ) or ( a7696a );
 a7701a <=( a7700a ) or ( a7693a );
 a7702a <=( a7701a ) or ( a7688a );
 a7706a <=( a1903a ) or ( a1904a );
 a7707a <=( a1905a ) or ( a7706a );
 a7710a <=( a1901a ) or ( a1902a );
 a7713a <=( a1899a ) or ( a1900a );
 a7714a <=( a7713a ) or ( a7710a );
 a7715a <=( a7714a ) or ( a7707a );
 a7718a <=( a1897a ) or ( a1898a );
 a7721a <=( a1895a ) or ( a1896a );
 a7722a <=( a7721a ) or ( a7718a );
 a7725a <=( a1893a ) or ( a1894a );
 a7728a <=( a1891a ) or ( a1892a );
 a7729a <=( a7728a ) or ( a7725a );
 a7730a <=( a7729a ) or ( a7722a );
 a7731a <=( a7730a ) or ( a7715a );
 a7732a <=( a7731a ) or ( a7702a );
 a7736a <=( a1888a ) or ( a1889a );
 a7737a <=( a1890a ) or ( a7736a );
 a7740a <=( a1886a ) or ( a1887a );
 a7743a <=( a1884a ) or ( a1885a );
 a7744a <=( a7743a ) or ( a7740a );
 a7745a <=( a7744a ) or ( a7737a );
 a7748a <=( a1882a ) or ( a1883a );
 a7751a <=( a1880a ) or ( a1881a );
 a7752a <=( a7751a ) or ( a7748a );
 a7755a <=( a1878a ) or ( a1879a );
 a7758a <=( a1876a ) or ( a1877a );
 a7759a <=( a7758a ) or ( a7755a );
 a7760a <=( a7759a ) or ( a7752a );
 a7761a <=( a7760a ) or ( a7745a );
 a7765a <=( a1873a ) or ( a1874a );
 a7766a <=( a1875a ) or ( a7765a );
 a7769a <=( a1871a ) or ( a1872a );
 a7772a <=( a1869a ) or ( a1870a );
 a7773a <=( a7772a ) or ( a7769a );
 a7774a <=( a7773a ) or ( a7766a );
 a7777a <=( a1867a ) or ( a1868a );
 a7780a <=( a1865a ) or ( a1866a );
 a7781a <=( a7780a ) or ( a7777a );
 a7784a <=( a1863a ) or ( a1864a );
 a7787a <=( a1861a ) or ( a1862a );
 a7788a <=( a7787a ) or ( a7784a );
 a7789a <=( a7788a ) or ( a7781a );
 a7790a <=( a7789a ) or ( a7774a );
 a7791a <=( a7790a ) or ( a7761a );
 a7792a <=( a7791a ) or ( a7732a );
 a7796a <=( a1858a ) or ( a1859a );
 a7797a <=( a1860a ) or ( a7796a );
 a7800a <=( a1856a ) or ( a1857a );
 a7803a <=( a1854a ) or ( a1855a );
 a7804a <=( a7803a ) or ( a7800a );
 a7805a <=( a7804a ) or ( a7797a );
 a7808a <=( a1852a ) or ( a1853a );
 a7811a <=( a1850a ) or ( a1851a );
 a7812a <=( a7811a ) or ( a7808a );
 a7815a <=( a1848a ) or ( a1849a );
 a7818a <=( a1846a ) or ( a1847a );
 a7819a <=( a7818a ) or ( a7815a );
 a7820a <=( a7819a ) or ( a7812a );
 a7821a <=( a7820a ) or ( a7805a );
 a7825a <=( a1843a ) or ( a1844a );
 a7826a <=( a1845a ) or ( a7825a );
 a7829a <=( a1841a ) or ( a1842a );
 a7832a <=( a1839a ) or ( a1840a );
 a7833a <=( a7832a ) or ( a7829a );
 a7834a <=( a7833a ) or ( a7826a );
 a7837a <=( a1837a ) or ( a1838a );
 a7840a <=( a1835a ) or ( a1836a );
 a7841a <=( a7840a ) or ( a7837a );
 a7844a <=( a1833a ) or ( a1834a );
 a7847a <=( a1831a ) or ( a1832a );
 a7848a <=( a7847a ) or ( a7844a );
 a7849a <=( a7848a ) or ( a7841a );
 a7850a <=( a7849a ) or ( a7834a );
 a7851a <=( a7850a ) or ( a7821a );
 a7855a <=( a1828a ) or ( a1829a );
 a7856a <=( a1830a ) or ( a7855a );
 a7859a <=( a1826a ) or ( a1827a );
 a7862a <=( a1824a ) or ( a1825a );
 a7863a <=( a7862a ) or ( a7859a );
 a7864a <=( a7863a ) or ( a7856a );
 a7867a <=( a1822a ) or ( a1823a );
 a7870a <=( a1820a ) or ( a1821a );
 a7871a <=( a7870a ) or ( a7867a );
 a7874a <=( a1818a ) or ( a1819a );
 a7877a <=( a1816a ) or ( a1817a );
 a7878a <=( a7877a ) or ( a7874a );
 a7879a <=( a7878a ) or ( a7871a );
 a7880a <=( a7879a ) or ( a7864a );
 a7884a <=( a1813a ) or ( a1814a );
 a7885a <=( a1815a ) or ( a7884a );
 a7888a <=( a1811a ) or ( a1812a );
 a7891a <=( a1809a ) or ( a1810a );
 a7892a <=( a7891a ) or ( a7888a );
 a7893a <=( a7892a ) or ( a7885a );
 a7896a <=( a1807a ) or ( a1808a );
 a7899a <=( a1805a ) or ( a1806a );
 a7900a <=( a7899a ) or ( a7896a );
 a7903a <=( a1803a ) or ( a1804a );
 a7906a <=( a1801a ) or ( a1802a );
 a7907a <=( a7906a ) or ( a7903a );
 a7908a <=( a7907a ) or ( a7900a );
 a7909a <=( a7908a ) or ( a7893a );
 a7910a <=( a7909a ) or ( a7880a );
 a7911a <=( a7910a ) or ( a7851a );
 a7912a <=( a7911a ) or ( a7792a );
 a7916a <=( a1798a ) or ( a1799a );
 a7917a <=( a1800a ) or ( a7916a );
 a7920a <=( a1796a ) or ( a1797a );
 a7923a <=( a1794a ) or ( a1795a );
 a7924a <=( a7923a ) or ( a7920a );
 a7925a <=( a7924a ) or ( a7917a );
 a7928a <=( a1792a ) or ( a1793a );
 a7931a <=( a1790a ) or ( a1791a );
 a7932a <=( a7931a ) or ( a7928a );
 a7935a <=( a1788a ) or ( a1789a );
 a7938a <=( a1786a ) or ( a1787a );
 a7939a <=( a7938a ) or ( a7935a );
 a7940a <=( a7939a ) or ( a7932a );
 a7941a <=( a7940a ) or ( a7925a );
 a7945a <=( a1783a ) or ( a1784a );
 a7946a <=( a1785a ) or ( a7945a );
 a7949a <=( a1781a ) or ( a1782a );
 a7952a <=( a1779a ) or ( a1780a );
 a7953a <=( a7952a ) or ( a7949a );
 a7954a <=( a7953a ) or ( a7946a );
 a7957a <=( a1777a ) or ( a1778a );
 a7960a <=( a1775a ) or ( a1776a );
 a7961a <=( a7960a ) or ( a7957a );
 a7964a <=( a1773a ) or ( a1774a );
 a7967a <=( a1771a ) or ( a1772a );
 a7968a <=( a7967a ) or ( a7964a );
 a7969a <=( a7968a ) or ( a7961a );
 a7970a <=( a7969a ) or ( a7954a );
 a7971a <=( a7970a ) or ( a7941a );
 a7975a <=( a1768a ) or ( a1769a );
 a7976a <=( a1770a ) or ( a7975a );
 a7979a <=( a1766a ) or ( a1767a );
 a7982a <=( a1764a ) or ( a1765a );
 a7983a <=( a7982a ) or ( a7979a );
 a7984a <=( a7983a ) or ( a7976a );
 a7987a <=( a1762a ) or ( a1763a );
 a7990a <=( a1760a ) or ( a1761a );
 a7991a <=( a7990a ) or ( a7987a );
 a7994a <=( a1758a ) or ( a1759a );
 a7997a <=( a1756a ) or ( a1757a );
 a7998a <=( a7997a ) or ( a7994a );
 a7999a <=( a7998a ) or ( a7991a );
 a8000a <=( a7999a ) or ( a7984a );
 a8004a <=( a1753a ) or ( a1754a );
 a8005a <=( a1755a ) or ( a8004a );
 a8008a <=( a1751a ) or ( a1752a );
 a8011a <=( a1749a ) or ( a1750a );
 a8012a <=( a8011a ) or ( a8008a );
 a8013a <=( a8012a ) or ( a8005a );
 a8016a <=( a1747a ) or ( a1748a );
 a8019a <=( a1745a ) or ( a1746a );
 a8020a <=( a8019a ) or ( a8016a );
 a8023a <=( a1743a ) or ( a1744a );
 a8026a <=( a1741a ) or ( a1742a );
 a8027a <=( a8026a ) or ( a8023a );
 a8028a <=( a8027a ) or ( a8020a );
 a8029a <=( a8028a ) or ( a8013a );
 a8030a <=( a8029a ) or ( a8000a );
 a8031a <=( a8030a ) or ( a7971a );
 a8035a <=( a1738a ) or ( a1739a );
 a8036a <=( a1740a ) or ( a8035a );
 a8039a <=( a1736a ) or ( a1737a );
 a8042a <=( a1734a ) or ( a1735a );
 a8043a <=( a8042a ) or ( a8039a );
 a8044a <=( a8043a ) or ( a8036a );
 a8047a <=( a1732a ) or ( a1733a );
 a8050a <=( a1730a ) or ( a1731a );
 a8051a <=( a8050a ) or ( a8047a );
 a8054a <=( a1728a ) or ( a1729a );
 a8057a <=( a1726a ) or ( a1727a );
 a8058a <=( a8057a ) or ( a8054a );
 a8059a <=( a8058a ) or ( a8051a );
 a8060a <=( a8059a ) or ( a8044a );
 a8064a <=( a1723a ) or ( a1724a );
 a8065a <=( a1725a ) or ( a8064a );
 a8068a <=( a1721a ) or ( a1722a );
 a8071a <=( a1719a ) or ( a1720a );
 a8072a <=( a8071a ) or ( a8068a );
 a8073a <=( a8072a ) or ( a8065a );
 a8076a <=( a1717a ) or ( a1718a );
 a8079a <=( a1715a ) or ( a1716a );
 a8080a <=( a8079a ) or ( a8076a );
 a8083a <=( a1713a ) or ( a1714a );
 a8086a <=( a1711a ) or ( a1712a );
 a8087a <=( a8086a ) or ( a8083a );
 a8088a <=( a8087a ) or ( a8080a );
 a8089a <=( a8088a ) or ( a8073a );
 a8090a <=( a8089a ) or ( a8060a );
 a8094a <=( a1708a ) or ( a1709a );
 a8095a <=( a1710a ) or ( a8094a );
 a8098a <=( a1706a ) or ( a1707a );
 a8101a <=( a1704a ) or ( a1705a );
 a8102a <=( a8101a ) or ( a8098a );
 a8103a <=( a8102a ) or ( a8095a );
 a8106a <=( a1702a ) or ( a1703a );
 a8109a <=( a1700a ) or ( a1701a );
 a8110a <=( a8109a ) or ( a8106a );
 a8113a <=( a1698a ) or ( a1699a );
 a8116a <=( a1696a ) or ( a1697a );
 a8117a <=( a8116a ) or ( a8113a );
 a8118a <=( a8117a ) or ( a8110a );
 a8119a <=( a8118a ) or ( a8103a );
 a8123a <=( a1693a ) or ( a1694a );
 a8124a <=( a1695a ) or ( a8123a );
 a8127a <=( a1691a ) or ( a1692a );
 a8130a <=( a1689a ) or ( a1690a );
 a8131a <=( a8130a ) or ( a8127a );
 a8132a <=( a8131a ) or ( a8124a );
 a8135a <=( a1687a ) or ( a1688a );
 a8138a <=( a1685a ) or ( a1686a );
 a8139a <=( a8138a ) or ( a8135a );
 a8142a <=( a1683a ) or ( a1684a );
 a8145a <=( a1681a ) or ( a1682a );
 a8146a <=( a8145a ) or ( a8142a );
 a8147a <=( a8146a ) or ( a8139a );
 a8148a <=( a8147a ) or ( a8132a );
 a8149a <=( a8148a ) or ( a8119a );
 a8150a <=( a8149a ) or ( a8090a );
 a8151a <=( a8150a ) or ( a8031a );
 a8152a <=( a8151a ) or ( a7912a );
 a8156a <=( a1678a ) or ( a1679a );
 a8157a <=( a1680a ) or ( a8156a );
 a8160a <=( a1676a ) or ( a1677a );
 a8163a <=( a1674a ) or ( a1675a );
 a8164a <=( a8163a ) or ( a8160a );
 a8165a <=( a8164a ) or ( a8157a );
 a8168a <=( a1672a ) or ( a1673a );
 a8171a <=( a1670a ) or ( a1671a );
 a8172a <=( a8171a ) or ( a8168a );
 a8175a <=( a1668a ) or ( a1669a );
 a8178a <=( a1666a ) or ( a1667a );
 a8179a <=( a8178a ) or ( a8175a );
 a8180a <=( a8179a ) or ( a8172a );
 a8181a <=( a8180a ) or ( a8165a );
 a8185a <=( a1663a ) or ( a1664a );
 a8186a <=( a1665a ) or ( a8185a );
 a8189a <=( a1661a ) or ( a1662a );
 a8192a <=( a1659a ) or ( a1660a );
 a8193a <=( a8192a ) or ( a8189a );
 a8194a <=( a8193a ) or ( a8186a );
 a8197a <=( a1657a ) or ( a1658a );
 a8200a <=( a1655a ) or ( a1656a );
 a8201a <=( a8200a ) or ( a8197a );
 a8204a <=( a1653a ) or ( a1654a );
 a8207a <=( a1651a ) or ( a1652a );
 a8208a <=( a8207a ) or ( a8204a );
 a8209a <=( a8208a ) or ( a8201a );
 a8210a <=( a8209a ) or ( a8194a );
 a8211a <=( a8210a ) or ( a8181a );
 a8215a <=( a1648a ) or ( a1649a );
 a8216a <=( a1650a ) or ( a8215a );
 a8219a <=( a1646a ) or ( a1647a );
 a8222a <=( a1644a ) or ( a1645a );
 a8223a <=( a8222a ) or ( a8219a );
 a8224a <=( a8223a ) or ( a8216a );
 a8227a <=( a1642a ) or ( a1643a );
 a8230a <=( a1640a ) or ( a1641a );
 a8231a <=( a8230a ) or ( a8227a );
 a8234a <=( a1638a ) or ( a1639a );
 a8237a <=( a1636a ) or ( a1637a );
 a8238a <=( a8237a ) or ( a8234a );
 a8239a <=( a8238a ) or ( a8231a );
 a8240a <=( a8239a ) or ( a8224a );
 a8244a <=( a1633a ) or ( a1634a );
 a8245a <=( a1635a ) or ( a8244a );
 a8248a <=( a1631a ) or ( a1632a );
 a8251a <=( a1629a ) or ( a1630a );
 a8252a <=( a8251a ) or ( a8248a );
 a8253a <=( a8252a ) or ( a8245a );
 a8256a <=( a1627a ) or ( a1628a );
 a8259a <=( a1625a ) or ( a1626a );
 a8260a <=( a8259a ) or ( a8256a );
 a8263a <=( a1623a ) or ( a1624a );
 a8266a <=( a1621a ) or ( a1622a );
 a8267a <=( a8266a ) or ( a8263a );
 a8268a <=( a8267a ) or ( a8260a );
 a8269a <=( a8268a ) or ( a8253a );
 a8270a <=( a8269a ) or ( a8240a );
 a8271a <=( a8270a ) or ( a8211a );
 a8275a <=( a1618a ) or ( a1619a );
 a8276a <=( a1620a ) or ( a8275a );
 a8279a <=( a1616a ) or ( a1617a );
 a8282a <=( a1614a ) or ( a1615a );
 a8283a <=( a8282a ) or ( a8279a );
 a8284a <=( a8283a ) or ( a8276a );
 a8287a <=( a1612a ) or ( a1613a );
 a8290a <=( a1610a ) or ( a1611a );
 a8291a <=( a8290a ) or ( a8287a );
 a8294a <=( a1608a ) or ( a1609a );
 a8297a <=( a1606a ) or ( a1607a );
 a8298a <=( a8297a ) or ( a8294a );
 a8299a <=( a8298a ) or ( a8291a );
 a8300a <=( a8299a ) or ( a8284a );
 a8304a <=( a1603a ) or ( a1604a );
 a8305a <=( a1605a ) or ( a8304a );
 a8308a <=( a1601a ) or ( a1602a );
 a8311a <=( a1599a ) or ( a1600a );
 a8312a <=( a8311a ) or ( a8308a );
 a8313a <=( a8312a ) or ( a8305a );
 a8316a <=( a1597a ) or ( a1598a );
 a8319a <=( a1595a ) or ( a1596a );
 a8320a <=( a8319a ) or ( a8316a );
 a8323a <=( a1593a ) or ( a1594a );
 a8326a <=( a1591a ) or ( a1592a );
 a8327a <=( a8326a ) or ( a8323a );
 a8328a <=( a8327a ) or ( a8320a );
 a8329a <=( a8328a ) or ( a8313a );
 a8330a <=( a8329a ) or ( a8300a );
 a8334a <=( a1588a ) or ( a1589a );
 a8335a <=( a1590a ) or ( a8334a );
 a8338a <=( a1586a ) or ( a1587a );
 a8341a <=( a1584a ) or ( a1585a );
 a8342a <=( a8341a ) or ( a8338a );
 a8343a <=( a8342a ) or ( a8335a );
 a8346a <=( a1582a ) or ( a1583a );
 a8349a <=( a1580a ) or ( a1581a );
 a8350a <=( a8349a ) or ( a8346a );
 a8353a <=( a1578a ) or ( a1579a );
 a8356a <=( a1576a ) or ( a1577a );
 a8357a <=( a8356a ) or ( a8353a );
 a8358a <=( a8357a ) or ( a8350a );
 a8359a <=( a8358a ) or ( a8343a );
 a8363a <=( a1573a ) or ( a1574a );
 a8364a <=( a1575a ) or ( a8363a );
 a8367a <=( a1571a ) or ( a1572a );
 a8370a <=( a1569a ) or ( a1570a );
 a8371a <=( a8370a ) or ( a8367a );
 a8372a <=( a8371a ) or ( a8364a );
 a8375a <=( a1567a ) or ( a1568a );
 a8378a <=( a1565a ) or ( a1566a );
 a8379a <=( a8378a ) or ( a8375a );
 a8382a <=( a1563a ) or ( a1564a );
 a8385a <=( a1561a ) or ( a1562a );
 a8386a <=( a8385a ) or ( a8382a );
 a8387a <=( a8386a ) or ( a8379a );
 a8388a <=( a8387a ) or ( a8372a );
 a8389a <=( a8388a ) or ( a8359a );
 a8390a <=( a8389a ) or ( a8330a );
 a8391a <=( a8390a ) or ( a8271a );
 a8395a <=( a1558a ) or ( a1559a );
 a8396a <=( a1560a ) or ( a8395a );
 a8399a <=( a1556a ) or ( a1557a );
 a8402a <=( a1554a ) or ( a1555a );
 a8403a <=( a8402a ) or ( a8399a );
 a8404a <=( a8403a ) or ( a8396a );
 a8407a <=( a1552a ) or ( a1553a );
 a8410a <=( a1550a ) or ( a1551a );
 a8411a <=( a8410a ) or ( a8407a );
 a8414a <=( a1548a ) or ( a1549a );
 a8417a <=( a1546a ) or ( a1547a );
 a8418a <=( a8417a ) or ( a8414a );
 a8419a <=( a8418a ) or ( a8411a );
 a8420a <=( a8419a ) or ( a8404a );
 a8424a <=( a1543a ) or ( a1544a );
 a8425a <=( a1545a ) or ( a8424a );
 a8428a <=( a1541a ) or ( a1542a );
 a8431a <=( a1539a ) or ( a1540a );
 a8432a <=( a8431a ) or ( a8428a );
 a8433a <=( a8432a ) or ( a8425a );
 a8436a <=( a1537a ) or ( a1538a );
 a8439a <=( a1535a ) or ( a1536a );
 a8440a <=( a8439a ) or ( a8436a );
 a8443a <=( a1533a ) or ( a1534a );
 a8446a <=( a1531a ) or ( a1532a );
 a8447a <=( a8446a ) or ( a8443a );
 a8448a <=( a8447a ) or ( a8440a );
 a8449a <=( a8448a ) or ( a8433a );
 a8450a <=( a8449a ) or ( a8420a );
 a8454a <=( a1528a ) or ( a1529a );
 a8455a <=( a1530a ) or ( a8454a );
 a8458a <=( a1526a ) or ( a1527a );
 a8461a <=( a1524a ) or ( a1525a );
 a8462a <=( a8461a ) or ( a8458a );
 a8463a <=( a8462a ) or ( a8455a );
 a8466a <=( a1522a ) or ( a1523a );
 a8469a <=( a1520a ) or ( a1521a );
 a8470a <=( a8469a ) or ( a8466a );
 a8473a <=( a1518a ) or ( a1519a );
 a8476a <=( a1516a ) or ( a1517a );
 a8477a <=( a8476a ) or ( a8473a );
 a8478a <=( a8477a ) or ( a8470a );
 a8479a <=( a8478a ) or ( a8463a );
 a8483a <=( a1513a ) or ( a1514a );
 a8484a <=( a1515a ) or ( a8483a );
 a8487a <=( a1511a ) or ( a1512a );
 a8490a <=( a1509a ) or ( a1510a );
 a8491a <=( a8490a ) or ( a8487a );
 a8492a <=( a8491a ) or ( a8484a );
 a8495a <=( a1507a ) or ( a1508a );
 a8498a <=( a1505a ) or ( a1506a );
 a8499a <=( a8498a ) or ( a8495a );
 a8502a <=( a1503a ) or ( a1504a );
 a8505a <=( a1501a ) or ( a1502a );
 a8506a <=( a8505a ) or ( a8502a );
 a8507a <=( a8506a ) or ( a8499a );
 a8508a <=( a8507a ) or ( a8492a );
 a8509a <=( a8508a ) or ( a8479a );
 a8510a <=( a8509a ) or ( a8450a );
 a8514a <=( a1498a ) or ( a1499a );
 a8515a <=( a1500a ) or ( a8514a );
 a8518a <=( a1496a ) or ( a1497a );
 a8521a <=( a1494a ) or ( a1495a );
 a8522a <=( a8521a ) or ( a8518a );
 a8523a <=( a8522a ) or ( a8515a );
 a8526a <=( a1492a ) or ( a1493a );
 a8529a <=( a1490a ) or ( a1491a );
 a8530a <=( a8529a ) or ( a8526a );
 a8533a <=( a1488a ) or ( a1489a );
 a8536a <=( a1486a ) or ( a1487a );
 a8537a <=( a8536a ) or ( a8533a );
 a8538a <=( a8537a ) or ( a8530a );
 a8539a <=( a8538a ) or ( a8523a );
 a8543a <=( a1483a ) or ( a1484a );
 a8544a <=( a1485a ) or ( a8543a );
 a8547a <=( a1481a ) or ( a1482a );
 a8550a <=( a1479a ) or ( a1480a );
 a8551a <=( a8550a ) or ( a8547a );
 a8552a <=( a8551a ) or ( a8544a );
 a8555a <=( a1477a ) or ( a1478a );
 a8558a <=( a1475a ) or ( a1476a );
 a8559a <=( a8558a ) or ( a8555a );
 a8562a <=( a1473a ) or ( a1474a );
 a8565a <=( a1471a ) or ( a1472a );
 a8566a <=( a8565a ) or ( a8562a );
 a8567a <=( a8566a ) or ( a8559a );
 a8568a <=( a8567a ) or ( a8552a );
 a8569a <=( a8568a ) or ( a8539a );
 a8573a <=( a1468a ) or ( a1469a );
 a8574a <=( a1470a ) or ( a8573a );
 a8577a <=( a1466a ) or ( a1467a );
 a8580a <=( a1464a ) or ( a1465a );
 a8581a <=( a8580a ) or ( a8577a );
 a8582a <=( a8581a ) or ( a8574a );
 a8585a <=( a1462a ) or ( a1463a );
 a8588a <=( a1460a ) or ( a1461a );
 a8589a <=( a8588a ) or ( a8585a );
 a8592a <=( a1458a ) or ( a1459a );
 a8595a <=( a1456a ) or ( a1457a );
 a8596a <=( a8595a ) or ( a8592a );
 a8597a <=( a8596a ) or ( a8589a );
 a8598a <=( a8597a ) or ( a8582a );
 a8602a <=( a1453a ) or ( a1454a );
 a8603a <=( a1455a ) or ( a8602a );
 a8606a <=( a1451a ) or ( a1452a );
 a8609a <=( a1449a ) or ( a1450a );
 a8610a <=( a8609a ) or ( a8606a );
 a8611a <=( a8610a ) or ( a8603a );
 a8614a <=( a1447a ) or ( a1448a );
 a8617a <=( a1445a ) or ( a1446a );
 a8618a <=( a8617a ) or ( a8614a );
 a8621a <=( a1443a ) or ( a1444a );
 a8624a <=( a1441a ) or ( a1442a );
 a8625a <=( a8624a ) or ( a8621a );
 a8626a <=( a8625a ) or ( a8618a );
 a8627a <=( a8626a ) or ( a8611a );
 a8628a <=( a8627a ) or ( a8598a );
 a8629a <=( a8628a ) or ( a8569a );
 a8630a <=( a8629a ) or ( a8510a );
 a8631a <=( a8630a ) or ( a8391a );
 a8632a <=( a8631a ) or ( a8152a );
 a8636a <=( a1438a ) or ( a1439a );
 a8637a <=( a1440a ) or ( a8636a );
 a8640a <=( a1436a ) or ( a1437a );
 a8643a <=( a1434a ) or ( a1435a );
 a8644a <=( a8643a ) or ( a8640a );
 a8645a <=( a8644a ) or ( a8637a );
 a8648a <=( a1432a ) or ( a1433a );
 a8651a <=( a1430a ) or ( a1431a );
 a8652a <=( a8651a ) or ( a8648a );
 a8655a <=( a1428a ) or ( a1429a );
 a8658a <=( a1426a ) or ( a1427a );
 a8659a <=( a8658a ) or ( a8655a );
 a8660a <=( a8659a ) or ( a8652a );
 a8661a <=( a8660a ) or ( a8645a );
 a8665a <=( a1423a ) or ( a1424a );
 a8666a <=( a1425a ) or ( a8665a );
 a8669a <=( a1421a ) or ( a1422a );
 a8672a <=( a1419a ) or ( a1420a );
 a8673a <=( a8672a ) or ( a8669a );
 a8674a <=( a8673a ) or ( a8666a );
 a8677a <=( a1417a ) or ( a1418a );
 a8680a <=( a1415a ) or ( a1416a );
 a8681a <=( a8680a ) or ( a8677a );
 a8684a <=( a1413a ) or ( a1414a );
 a8687a <=( a1411a ) or ( a1412a );
 a8688a <=( a8687a ) or ( a8684a );
 a8689a <=( a8688a ) or ( a8681a );
 a8690a <=( a8689a ) or ( a8674a );
 a8691a <=( a8690a ) or ( a8661a );
 a8695a <=( a1408a ) or ( a1409a );
 a8696a <=( a1410a ) or ( a8695a );
 a8699a <=( a1406a ) or ( a1407a );
 a8702a <=( a1404a ) or ( a1405a );
 a8703a <=( a8702a ) or ( a8699a );
 a8704a <=( a8703a ) or ( a8696a );
 a8707a <=( a1402a ) or ( a1403a );
 a8710a <=( a1400a ) or ( a1401a );
 a8711a <=( a8710a ) or ( a8707a );
 a8714a <=( a1398a ) or ( a1399a );
 a8717a <=( a1396a ) or ( a1397a );
 a8718a <=( a8717a ) or ( a8714a );
 a8719a <=( a8718a ) or ( a8711a );
 a8720a <=( a8719a ) or ( a8704a );
 a8724a <=( a1393a ) or ( a1394a );
 a8725a <=( a1395a ) or ( a8724a );
 a8728a <=( a1391a ) or ( a1392a );
 a8731a <=( a1389a ) or ( a1390a );
 a8732a <=( a8731a ) or ( a8728a );
 a8733a <=( a8732a ) or ( a8725a );
 a8736a <=( a1387a ) or ( a1388a );
 a8739a <=( a1385a ) or ( a1386a );
 a8740a <=( a8739a ) or ( a8736a );
 a8743a <=( a1383a ) or ( a1384a );
 a8746a <=( a1381a ) or ( a1382a );
 a8747a <=( a8746a ) or ( a8743a );
 a8748a <=( a8747a ) or ( a8740a );
 a8749a <=( a8748a ) or ( a8733a );
 a8750a <=( a8749a ) or ( a8720a );
 a8751a <=( a8750a ) or ( a8691a );
 a8755a <=( a1378a ) or ( a1379a );
 a8756a <=( a1380a ) or ( a8755a );
 a8759a <=( a1376a ) or ( a1377a );
 a8762a <=( a1374a ) or ( a1375a );
 a8763a <=( a8762a ) or ( a8759a );
 a8764a <=( a8763a ) or ( a8756a );
 a8767a <=( a1372a ) or ( a1373a );
 a8770a <=( a1370a ) or ( a1371a );
 a8771a <=( a8770a ) or ( a8767a );
 a8774a <=( a1368a ) or ( a1369a );
 a8777a <=( a1366a ) or ( a1367a );
 a8778a <=( a8777a ) or ( a8774a );
 a8779a <=( a8778a ) or ( a8771a );
 a8780a <=( a8779a ) or ( a8764a );
 a8784a <=( a1363a ) or ( a1364a );
 a8785a <=( a1365a ) or ( a8784a );
 a8788a <=( a1361a ) or ( a1362a );
 a8791a <=( a1359a ) or ( a1360a );
 a8792a <=( a8791a ) or ( a8788a );
 a8793a <=( a8792a ) or ( a8785a );
 a8796a <=( a1357a ) or ( a1358a );
 a8799a <=( a1355a ) or ( a1356a );
 a8800a <=( a8799a ) or ( a8796a );
 a8803a <=( a1353a ) or ( a1354a );
 a8806a <=( a1351a ) or ( a1352a );
 a8807a <=( a8806a ) or ( a8803a );
 a8808a <=( a8807a ) or ( a8800a );
 a8809a <=( a8808a ) or ( a8793a );
 a8810a <=( a8809a ) or ( a8780a );
 a8814a <=( a1348a ) or ( a1349a );
 a8815a <=( a1350a ) or ( a8814a );
 a8818a <=( a1346a ) or ( a1347a );
 a8821a <=( a1344a ) or ( a1345a );
 a8822a <=( a8821a ) or ( a8818a );
 a8823a <=( a8822a ) or ( a8815a );
 a8826a <=( a1342a ) or ( a1343a );
 a8829a <=( a1340a ) or ( a1341a );
 a8830a <=( a8829a ) or ( a8826a );
 a8833a <=( a1338a ) or ( a1339a );
 a8836a <=( a1336a ) or ( a1337a );
 a8837a <=( a8836a ) or ( a8833a );
 a8838a <=( a8837a ) or ( a8830a );
 a8839a <=( a8838a ) or ( a8823a );
 a8843a <=( a1333a ) or ( a1334a );
 a8844a <=( a1335a ) or ( a8843a );
 a8847a <=( a1331a ) or ( a1332a );
 a8850a <=( a1329a ) or ( a1330a );
 a8851a <=( a8850a ) or ( a8847a );
 a8852a <=( a8851a ) or ( a8844a );
 a8855a <=( a1327a ) or ( a1328a );
 a8858a <=( a1325a ) or ( a1326a );
 a8859a <=( a8858a ) or ( a8855a );
 a8862a <=( a1323a ) or ( a1324a );
 a8865a <=( a1321a ) or ( a1322a );
 a8866a <=( a8865a ) or ( a8862a );
 a8867a <=( a8866a ) or ( a8859a );
 a8868a <=( a8867a ) or ( a8852a );
 a8869a <=( a8868a ) or ( a8839a );
 a8870a <=( a8869a ) or ( a8810a );
 a8871a <=( a8870a ) or ( a8751a );
 a8875a <=( a1318a ) or ( a1319a );
 a8876a <=( a1320a ) or ( a8875a );
 a8879a <=( a1316a ) or ( a1317a );
 a8882a <=( a1314a ) or ( a1315a );
 a8883a <=( a8882a ) or ( a8879a );
 a8884a <=( a8883a ) or ( a8876a );
 a8887a <=( a1312a ) or ( a1313a );
 a8890a <=( a1310a ) or ( a1311a );
 a8891a <=( a8890a ) or ( a8887a );
 a8894a <=( a1308a ) or ( a1309a );
 a8897a <=( a1306a ) or ( a1307a );
 a8898a <=( a8897a ) or ( a8894a );
 a8899a <=( a8898a ) or ( a8891a );
 a8900a <=( a8899a ) or ( a8884a );
 a8904a <=( a1303a ) or ( a1304a );
 a8905a <=( a1305a ) or ( a8904a );
 a8908a <=( a1301a ) or ( a1302a );
 a8911a <=( a1299a ) or ( a1300a );
 a8912a <=( a8911a ) or ( a8908a );
 a8913a <=( a8912a ) or ( a8905a );
 a8916a <=( a1297a ) or ( a1298a );
 a8919a <=( a1295a ) or ( a1296a );
 a8920a <=( a8919a ) or ( a8916a );
 a8923a <=( a1293a ) or ( a1294a );
 a8926a <=( a1291a ) or ( a1292a );
 a8927a <=( a8926a ) or ( a8923a );
 a8928a <=( a8927a ) or ( a8920a );
 a8929a <=( a8928a ) or ( a8913a );
 a8930a <=( a8929a ) or ( a8900a );
 a8934a <=( a1288a ) or ( a1289a );
 a8935a <=( a1290a ) or ( a8934a );
 a8938a <=( a1286a ) or ( a1287a );
 a8941a <=( a1284a ) or ( a1285a );
 a8942a <=( a8941a ) or ( a8938a );
 a8943a <=( a8942a ) or ( a8935a );
 a8946a <=( a1282a ) or ( a1283a );
 a8949a <=( a1280a ) or ( a1281a );
 a8950a <=( a8949a ) or ( a8946a );
 a8953a <=( a1278a ) or ( a1279a );
 a8956a <=( a1276a ) or ( a1277a );
 a8957a <=( a8956a ) or ( a8953a );
 a8958a <=( a8957a ) or ( a8950a );
 a8959a <=( a8958a ) or ( a8943a );
 a8963a <=( a1273a ) or ( a1274a );
 a8964a <=( a1275a ) or ( a8963a );
 a8967a <=( a1271a ) or ( a1272a );
 a8970a <=( a1269a ) or ( a1270a );
 a8971a <=( a8970a ) or ( a8967a );
 a8972a <=( a8971a ) or ( a8964a );
 a8975a <=( a1267a ) or ( a1268a );
 a8978a <=( a1265a ) or ( a1266a );
 a8979a <=( a8978a ) or ( a8975a );
 a8982a <=( a1263a ) or ( a1264a );
 a8985a <=( a1261a ) or ( a1262a );
 a8986a <=( a8985a ) or ( a8982a );
 a8987a <=( a8986a ) or ( a8979a );
 a8988a <=( a8987a ) or ( a8972a );
 a8989a <=( a8988a ) or ( a8959a );
 a8990a <=( a8989a ) or ( a8930a );
 a8994a <=( a1258a ) or ( a1259a );
 a8995a <=( a1260a ) or ( a8994a );
 a8998a <=( a1256a ) or ( a1257a );
 a9001a <=( a1254a ) or ( a1255a );
 a9002a <=( a9001a ) or ( a8998a );
 a9003a <=( a9002a ) or ( a8995a );
 a9006a <=( a1252a ) or ( a1253a );
 a9009a <=( a1250a ) or ( a1251a );
 a9010a <=( a9009a ) or ( a9006a );
 a9013a <=( a1248a ) or ( a1249a );
 a9016a <=( a1246a ) or ( a1247a );
 a9017a <=( a9016a ) or ( a9013a );
 a9018a <=( a9017a ) or ( a9010a );
 a9019a <=( a9018a ) or ( a9003a );
 a9023a <=( a1243a ) or ( a1244a );
 a9024a <=( a1245a ) or ( a9023a );
 a9027a <=( a1241a ) or ( a1242a );
 a9030a <=( a1239a ) or ( a1240a );
 a9031a <=( a9030a ) or ( a9027a );
 a9032a <=( a9031a ) or ( a9024a );
 a9035a <=( a1237a ) or ( a1238a );
 a9038a <=( a1235a ) or ( a1236a );
 a9039a <=( a9038a ) or ( a9035a );
 a9042a <=( a1233a ) or ( a1234a );
 a9045a <=( a1231a ) or ( a1232a );
 a9046a <=( a9045a ) or ( a9042a );
 a9047a <=( a9046a ) or ( a9039a );
 a9048a <=( a9047a ) or ( a9032a );
 a9049a <=( a9048a ) or ( a9019a );
 a9053a <=( a1228a ) or ( a1229a );
 a9054a <=( a1230a ) or ( a9053a );
 a9057a <=( a1226a ) or ( a1227a );
 a9060a <=( a1224a ) or ( a1225a );
 a9061a <=( a9060a ) or ( a9057a );
 a9062a <=( a9061a ) or ( a9054a );
 a9065a <=( a1222a ) or ( a1223a );
 a9068a <=( a1220a ) or ( a1221a );
 a9069a <=( a9068a ) or ( a9065a );
 a9072a <=( a1218a ) or ( a1219a );
 a9075a <=( a1216a ) or ( a1217a );
 a9076a <=( a9075a ) or ( a9072a );
 a9077a <=( a9076a ) or ( a9069a );
 a9078a <=( a9077a ) or ( a9062a );
 a9082a <=( a1213a ) or ( a1214a );
 a9083a <=( a1215a ) or ( a9082a );
 a9086a <=( a1211a ) or ( a1212a );
 a9089a <=( a1209a ) or ( a1210a );
 a9090a <=( a9089a ) or ( a9086a );
 a9091a <=( a9090a ) or ( a9083a );
 a9094a <=( a1207a ) or ( a1208a );
 a9097a <=( a1205a ) or ( a1206a );
 a9098a <=( a9097a ) or ( a9094a );
 a9101a <=( a1203a ) or ( a1204a );
 a9104a <=( a1201a ) or ( a1202a );
 a9105a <=( a9104a ) or ( a9101a );
 a9106a <=( a9105a ) or ( a9098a );
 a9107a <=( a9106a ) or ( a9091a );
 a9108a <=( a9107a ) or ( a9078a );
 a9109a <=( a9108a ) or ( a9049a );
 a9110a <=( a9109a ) or ( a8990a );
 a9111a <=( a9110a ) or ( a8871a );
 a9115a <=( a1198a ) or ( a1199a );
 a9116a <=( a1200a ) or ( a9115a );
 a9119a <=( a1196a ) or ( a1197a );
 a9122a <=( a1194a ) or ( a1195a );
 a9123a <=( a9122a ) or ( a9119a );
 a9124a <=( a9123a ) or ( a9116a );
 a9127a <=( a1192a ) or ( a1193a );
 a9130a <=( a1190a ) or ( a1191a );
 a9131a <=( a9130a ) or ( a9127a );
 a9134a <=( a1188a ) or ( a1189a );
 a9137a <=( a1186a ) or ( a1187a );
 a9138a <=( a9137a ) or ( a9134a );
 a9139a <=( a9138a ) or ( a9131a );
 a9140a <=( a9139a ) or ( a9124a );
 a9144a <=( a1183a ) or ( a1184a );
 a9145a <=( a1185a ) or ( a9144a );
 a9148a <=( a1181a ) or ( a1182a );
 a9151a <=( a1179a ) or ( a1180a );
 a9152a <=( a9151a ) or ( a9148a );
 a9153a <=( a9152a ) or ( a9145a );
 a9156a <=( a1177a ) or ( a1178a );
 a9159a <=( a1175a ) or ( a1176a );
 a9160a <=( a9159a ) or ( a9156a );
 a9163a <=( a1173a ) or ( a1174a );
 a9166a <=( a1171a ) or ( a1172a );
 a9167a <=( a9166a ) or ( a9163a );
 a9168a <=( a9167a ) or ( a9160a );
 a9169a <=( a9168a ) or ( a9153a );
 a9170a <=( a9169a ) or ( a9140a );
 a9174a <=( a1168a ) or ( a1169a );
 a9175a <=( a1170a ) or ( a9174a );
 a9178a <=( a1166a ) or ( a1167a );
 a9181a <=( a1164a ) or ( a1165a );
 a9182a <=( a9181a ) or ( a9178a );
 a9183a <=( a9182a ) or ( a9175a );
 a9186a <=( a1162a ) or ( a1163a );
 a9189a <=( a1160a ) or ( a1161a );
 a9190a <=( a9189a ) or ( a9186a );
 a9193a <=( a1158a ) or ( a1159a );
 a9196a <=( a1156a ) or ( a1157a );
 a9197a <=( a9196a ) or ( a9193a );
 a9198a <=( a9197a ) or ( a9190a );
 a9199a <=( a9198a ) or ( a9183a );
 a9203a <=( a1153a ) or ( a1154a );
 a9204a <=( a1155a ) or ( a9203a );
 a9207a <=( a1151a ) or ( a1152a );
 a9210a <=( a1149a ) or ( a1150a );
 a9211a <=( a9210a ) or ( a9207a );
 a9212a <=( a9211a ) or ( a9204a );
 a9215a <=( a1147a ) or ( a1148a );
 a9218a <=( a1145a ) or ( a1146a );
 a9219a <=( a9218a ) or ( a9215a );
 a9222a <=( a1143a ) or ( a1144a );
 a9225a <=( a1141a ) or ( a1142a );
 a9226a <=( a9225a ) or ( a9222a );
 a9227a <=( a9226a ) or ( a9219a );
 a9228a <=( a9227a ) or ( a9212a );
 a9229a <=( a9228a ) or ( a9199a );
 a9230a <=( a9229a ) or ( a9170a );
 a9234a <=( a1138a ) or ( a1139a );
 a9235a <=( a1140a ) or ( a9234a );
 a9238a <=( a1136a ) or ( a1137a );
 a9241a <=( a1134a ) or ( a1135a );
 a9242a <=( a9241a ) or ( a9238a );
 a9243a <=( a9242a ) or ( a9235a );
 a9246a <=( a1132a ) or ( a1133a );
 a9249a <=( a1130a ) or ( a1131a );
 a9250a <=( a9249a ) or ( a9246a );
 a9253a <=( a1128a ) or ( a1129a );
 a9256a <=( a1126a ) or ( a1127a );
 a9257a <=( a9256a ) or ( a9253a );
 a9258a <=( a9257a ) or ( a9250a );
 a9259a <=( a9258a ) or ( a9243a );
 a9263a <=( a1123a ) or ( a1124a );
 a9264a <=( a1125a ) or ( a9263a );
 a9267a <=( a1121a ) or ( a1122a );
 a9270a <=( a1119a ) or ( a1120a );
 a9271a <=( a9270a ) or ( a9267a );
 a9272a <=( a9271a ) or ( a9264a );
 a9275a <=( a1117a ) or ( a1118a );
 a9278a <=( a1115a ) or ( a1116a );
 a9279a <=( a9278a ) or ( a9275a );
 a9282a <=( a1113a ) or ( a1114a );
 a9285a <=( a1111a ) or ( a1112a );
 a9286a <=( a9285a ) or ( a9282a );
 a9287a <=( a9286a ) or ( a9279a );
 a9288a <=( a9287a ) or ( a9272a );
 a9289a <=( a9288a ) or ( a9259a );
 a9293a <=( a1108a ) or ( a1109a );
 a9294a <=( a1110a ) or ( a9293a );
 a9297a <=( a1106a ) or ( a1107a );
 a9300a <=( a1104a ) or ( a1105a );
 a9301a <=( a9300a ) or ( a9297a );
 a9302a <=( a9301a ) or ( a9294a );
 a9305a <=( a1102a ) or ( a1103a );
 a9308a <=( a1100a ) or ( a1101a );
 a9309a <=( a9308a ) or ( a9305a );
 a9312a <=( a1098a ) or ( a1099a );
 a9315a <=( a1096a ) or ( a1097a );
 a9316a <=( a9315a ) or ( a9312a );
 a9317a <=( a9316a ) or ( a9309a );
 a9318a <=( a9317a ) or ( a9302a );
 a9322a <=( a1093a ) or ( a1094a );
 a9323a <=( a1095a ) or ( a9322a );
 a9326a <=( a1091a ) or ( a1092a );
 a9329a <=( a1089a ) or ( a1090a );
 a9330a <=( a9329a ) or ( a9326a );
 a9331a <=( a9330a ) or ( a9323a );
 a9334a <=( a1087a ) or ( a1088a );
 a9337a <=( a1085a ) or ( a1086a );
 a9338a <=( a9337a ) or ( a9334a );
 a9341a <=( a1083a ) or ( a1084a );
 a9344a <=( a1081a ) or ( a1082a );
 a9345a <=( a9344a ) or ( a9341a );
 a9346a <=( a9345a ) or ( a9338a );
 a9347a <=( a9346a ) or ( a9331a );
 a9348a <=( a9347a ) or ( a9318a );
 a9349a <=( a9348a ) or ( a9289a );
 a9350a <=( a9349a ) or ( a9230a );
 a9354a <=( a1078a ) or ( a1079a );
 a9355a <=( a1080a ) or ( a9354a );
 a9358a <=( a1076a ) or ( a1077a );
 a9361a <=( a1074a ) or ( a1075a );
 a9362a <=( a9361a ) or ( a9358a );
 a9363a <=( a9362a ) or ( a9355a );
 a9366a <=( a1072a ) or ( a1073a );
 a9369a <=( a1070a ) or ( a1071a );
 a9370a <=( a9369a ) or ( a9366a );
 a9373a <=( a1068a ) or ( a1069a );
 a9376a <=( a1066a ) or ( a1067a );
 a9377a <=( a9376a ) or ( a9373a );
 a9378a <=( a9377a ) or ( a9370a );
 a9379a <=( a9378a ) or ( a9363a );
 a9383a <=( a1063a ) or ( a1064a );
 a9384a <=( a1065a ) or ( a9383a );
 a9387a <=( a1061a ) or ( a1062a );
 a9390a <=( a1059a ) or ( a1060a );
 a9391a <=( a9390a ) or ( a9387a );
 a9392a <=( a9391a ) or ( a9384a );
 a9395a <=( a1057a ) or ( a1058a );
 a9398a <=( a1055a ) or ( a1056a );
 a9399a <=( a9398a ) or ( a9395a );
 a9402a <=( a1053a ) or ( a1054a );
 a9405a <=( a1051a ) or ( a1052a );
 a9406a <=( a9405a ) or ( a9402a );
 a9407a <=( a9406a ) or ( a9399a );
 a9408a <=( a9407a ) or ( a9392a );
 a9409a <=( a9408a ) or ( a9379a );
 a9413a <=( a1048a ) or ( a1049a );
 a9414a <=( a1050a ) or ( a9413a );
 a9417a <=( a1046a ) or ( a1047a );
 a9420a <=( a1044a ) or ( a1045a );
 a9421a <=( a9420a ) or ( a9417a );
 a9422a <=( a9421a ) or ( a9414a );
 a9425a <=( a1042a ) or ( a1043a );
 a9428a <=( a1040a ) or ( a1041a );
 a9429a <=( a9428a ) or ( a9425a );
 a9432a <=( a1038a ) or ( a1039a );
 a9435a <=( a1036a ) or ( a1037a );
 a9436a <=( a9435a ) or ( a9432a );
 a9437a <=( a9436a ) or ( a9429a );
 a9438a <=( a9437a ) or ( a9422a );
 a9442a <=( a1033a ) or ( a1034a );
 a9443a <=( a1035a ) or ( a9442a );
 a9446a <=( a1031a ) or ( a1032a );
 a9449a <=( a1029a ) or ( a1030a );
 a9450a <=( a9449a ) or ( a9446a );
 a9451a <=( a9450a ) or ( a9443a );
 a9454a <=( a1027a ) or ( a1028a );
 a9457a <=( a1025a ) or ( a1026a );
 a9458a <=( a9457a ) or ( a9454a );
 a9461a <=( a1023a ) or ( a1024a );
 a9464a <=( a1021a ) or ( a1022a );
 a9465a <=( a9464a ) or ( a9461a );
 a9466a <=( a9465a ) or ( a9458a );
 a9467a <=( a9466a ) or ( a9451a );
 a9468a <=( a9467a ) or ( a9438a );
 a9469a <=( a9468a ) or ( a9409a );
 a9473a <=( a1018a ) or ( a1019a );
 a9474a <=( a1020a ) or ( a9473a );
 a9477a <=( a1016a ) or ( a1017a );
 a9480a <=( a1014a ) or ( a1015a );
 a9481a <=( a9480a ) or ( a9477a );
 a9482a <=( a9481a ) or ( a9474a );
 a9485a <=( a1012a ) or ( a1013a );
 a9488a <=( a1010a ) or ( a1011a );
 a9489a <=( a9488a ) or ( a9485a );
 a9492a <=( a1008a ) or ( a1009a );
 a9495a <=( a1006a ) or ( a1007a );
 a9496a <=( a9495a ) or ( a9492a );
 a9497a <=( a9496a ) or ( a9489a );
 a9498a <=( a9497a ) or ( a9482a );
 a9502a <=( a1003a ) or ( a1004a );
 a9503a <=( a1005a ) or ( a9502a );
 a9506a <=( a1001a ) or ( a1002a );
 a9509a <=( a999a ) or ( a1000a );
 a9510a <=( a9509a ) or ( a9506a );
 a9511a <=( a9510a ) or ( a9503a );
 a9514a <=( a997a ) or ( a998a );
 a9517a <=( a995a ) or ( a996a );
 a9518a <=( a9517a ) or ( a9514a );
 a9521a <=( a993a ) or ( a994a );
 a9524a <=( a991a ) or ( a992a );
 a9525a <=( a9524a ) or ( a9521a );
 a9526a <=( a9525a ) or ( a9518a );
 a9527a <=( a9526a ) or ( a9511a );
 a9528a <=( a9527a ) or ( a9498a );
 a9532a <=( a988a ) or ( a989a );
 a9533a <=( a990a ) or ( a9532a );
 a9536a <=( a986a ) or ( a987a );
 a9539a <=( a984a ) or ( a985a );
 a9540a <=( a9539a ) or ( a9536a );
 a9541a <=( a9540a ) or ( a9533a );
 a9544a <=( a982a ) or ( a983a );
 a9547a <=( a980a ) or ( a981a );
 a9548a <=( a9547a ) or ( a9544a );
 a9551a <=( a978a ) or ( a979a );
 a9554a <=( a976a ) or ( a977a );
 a9555a <=( a9554a ) or ( a9551a );
 a9556a <=( a9555a ) or ( a9548a );
 a9557a <=( a9556a ) or ( a9541a );
 a9561a <=( a973a ) or ( a974a );
 a9562a <=( a975a ) or ( a9561a );
 a9565a <=( a971a ) or ( a972a );
 a9568a <=( a969a ) or ( a970a );
 a9569a <=( a9568a ) or ( a9565a );
 a9570a <=( a9569a ) or ( a9562a );
 a9573a <=( a967a ) or ( a968a );
 a9576a <=( a965a ) or ( a966a );
 a9577a <=( a9576a ) or ( a9573a );
 a9580a <=( a963a ) or ( a964a );
 a9583a <=( a961a ) or ( a962a );
 a9584a <=( a9583a ) or ( a9580a );
 a9585a <=( a9584a ) or ( a9577a );
 a9586a <=( a9585a ) or ( a9570a );
 a9587a <=( a9586a ) or ( a9557a );
 a9588a <=( a9587a ) or ( a9528a );
 a9589a <=( a9588a ) or ( a9469a );
 a9590a <=( a9589a ) or ( a9350a );
 a9591a <=( a9590a ) or ( a9111a );
 a9592a <=( a9591a ) or ( a8632a );
 a9596a <=( a958a ) or ( a959a );
 a9597a <=( a960a ) or ( a9596a );
 a9600a <=( a956a ) or ( a957a );
 a9603a <=( a954a ) or ( a955a );
 a9604a <=( a9603a ) or ( a9600a );
 a9605a <=( a9604a ) or ( a9597a );
 a9608a <=( a952a ) or ( a953a );
 a9611a <=( a950a ) or ( a951a );
 a9612a <=( a9611a ) or ( a9608a );
 a9615a <=( a948a ) or ( a949a );
 a9618a <=( a946a ) or ( a947a );
 a9619a <=( a9618a ) or ( a9615a );
 a9620a <=( a9619a ) or ( a9612a );
 a9621a <=( a9620a ) or ( a9605a );
 a9625a <=( a943a ) or ( a944a );
 a9626a <=( a945a ) or ( a9625a );
 a9629a <=( a941a ) or ( a942a );
 a9632a <=( a939a ) or ( a940a );
 a9633a <=( a9632a ) or ( a9629a );
 a9634a <=( a9633a ) or ( a9626a );
 a9637a <=( a937a ) or ( a938a );
 a9640a <=( a935a ) or ( a936a );
 a9641a <=( a9640a ) or ( a9637a );
 a9644a <=( a933a ) or ( a934a );
 a9647a <=( a931a ) or ( a932a );
 a9648a <=( a9647a ) or ( a9644a );
 a9649a <=( a9648a ) or ( a9641a );
 a9650a <=( a9649a ) or ( a9634a );
 a9651a <=( a9650a ) or ( a9621a );
 a9655a <=( a928a ) or ( a929a );
 a9656a <=( a930a ) or ( a9655a );
 a9659a <=( a926a ) or ( a927a );
 a9662a <=( a924a ) or ( a925a );
 a9663a <=( a9662a ) or ( a9659a );
 a9664a <=( a9663a ) or ( a9656a );
 a9667a <=( a922a ) or ( a923a );
 a9670a <=( a920a ) or ( a921a );
 a9671a <=( a9670a ) or ( a9667a );
 a9674a <=( a918a ) or ( a919a );
 a9677a <=( a916a ) or ( a917a );
 a9678a <=( a9677a ) or ( a9674a );
 a9679a <=( a9678a ) or ( a9671a );
 a9680a <=( a9679a ) or ( a9664a );
 a9684a <=( a913a ) or ( a914a );
 a9685a <=( a915a ) or ( a9684a );
 a9688a <=( a911a ) or ( a912a );
 a9691a <=( a909a ) or ( a910a );
 a9692a <=( a9691a ) or ( a9688a );
 a9693a <=( a9692a ) or ( a9685a );
 a9696a <=( a907a ) or ( a908a );
 a9699a <=( a905a ) or ( a906a );
 a9700a <=( a9699a ) or ( a9696a );
 a9703a <=( a903a ) or ( a904a );
 a9706a <=( a901a ) or ( a902a );
 a9707a <=( a9706a ) or ( a9703a );
 a9708a <=( a9707a ) or ( a9700a );
 a9709a <=( a9708a ) or ( a9693a );
 a9710a <=( a9709a ) or ( a9680a );
 a9711a <=( a9710a ) or ( a9651a );
 a9715a <=( a898a ) or ( a899a );
 a9716a <=( a900a ) or ( a9715a );
 a9719a <=( a896a ) or ( a897a );
 a9722a <=( a894a ) or ( a895a );
 a9723a <=( a9722a ) or ( a9719a );
 a9724a <=( a9723a ) or ( a9716a );
 a9727a <=( a892a ) or ( a893a );
 a9730a <=( a890a ) or ( a891a );
 a9731a <=( a9730a ) or ( a9727a );
 a9734a <=( a888a ) or ( a889a );
 a9737a <=( a886a ) or ( a887a );
 a9738a <=( a9737a ) or ( a9734a );
 a9739a <=( a9738a ) or ( a9731a );
 a9740a <=( a9739a ) or ( a9724a );
 a9744a <=( a883a ) or ( a884a );
 a9745a <=( a885a ) or ( a9744a );
 a9748a <=( a881a ) or ( a882a );
 a9751a <=( a879a ) or ( a880a );
 a9752a <=( a9751a ) or ( a9748a );
 a9753a <=( a9752a ) or ( a9745a );
 a9756a <=( a877a ) or ( a878a );
 a9759a <=( a875a ) or ( a876a );
 a9760a <=( a9759a ) or ( a9756a );
 a9763a <=( a873a ) or ( a874a );
 a9766a <=( a871a ) or ( a872a );
 a9767a <=( a9766a ) or ( a9763a );
 a9768a <=( a9767a ) or ( a9760a );
 a9769a <=( a9768a ) or ( a9753a );
 a9770a <=( a9769a ) or ( a9740a );
 a9774a <=( a868a ) or ( a869a );
 a9775a <=( a870a ) or ( a9774a );
 a9778a <=( a866a ) or ( a867a );
 a9781a <=( a864a ) or ( a865a );
 a9782a <=( a9781a ) or ( a9778a );
 a9783a <=( a9782a ) or ( a9775a );
 a9786a <=( a862a ) or ( a863a );
 a9789a <=( a860a ) or ( a861a );
 a9790a <=( a9789a ) or ( a9786a );
 a9793a <=( a858a ) or ( a859a );
 a9796a <=( a856a ) or ( a857a );
 a9797a <=( a9796a ) or ( a9793a );
 a9798a <=( a9797a ) or ( a9790a );
 a9799a <=( a9798a ) or ( a9783a );
 a9803a <=( a853a ) or ( a854a );
 a9804a <=( a855a ) or ( a9803a );
 a9807a <=( a851a ) or ( a852a );
 a9810a <=( a849a ) or ( a850a );
 a9811a <=( a9810a ) or ( a9807a );
 a9812a <=( a9811a ) or ( a9804a );
 a9815a <=( a847a ) or ( a848a );
 a9818a <=( a845a ) or ( a846a );
 a9819a <=( a9818a ) or ( a9815a );
 a9822a <=( a843a ) or ( a844a );
 a9825a <=( a841a ) or ( a842a );
 a9826a <=( a9825a ) or ( a9822a );
 a9827a <=( a9826a ) or ( a9819a );
 a9828a <=( a9827a ) or ( a9812a );
 a9829a <=( a9828a ) or ( a9799a );
 a9830a <=( a9829a ) or ( a9770a );
 a9831a <=( a9830a ) or ( a9711a );
 a9835a <=( a838a ) or ( a839a );
 a9836a <=( a840a ) or ( a9835a );
 a9839a <=( a836a ) or ( a837a );
 a9842a <=( a834a ) or ( a835a );
 a9843a <=( a9842a ) or ( a9839a );
 a9844a <=( a9843a ) or ( a9836a );
 a9847a <=( a832a ) or ( a833a );
 a9850a <=( a830a ) or ( a831a );
 a9851a <=( a9850a ) or ( a9847a );
 a9854a <=( a828a ) or ( a829a );
 a9857a <=( a826a ) or ( a827a );
 a9858a <=( a9857a ) or ( a9854a );
 a9859a <=( a9858a ) or ( a9851a );
 a9860a <=( a9859a ) or ( a9844a );
 a9864a <=( a823a ) or ( a824a );
 a9865a <=( a825a ) or ( a9864a );
 a9868a <=( a821a ) or ( a822a );
 a9871a <=( a819a ) or ( a820a );
 a9872a <=( a9871a ) or ( a9868a );
 a9873a <=( a9872a ) or ( a9865a );
 a9876a <=( a817a ) or ( a818a );
 a9879a <=( a815a ) or ( a816a );
 a9880a <=( a9879a ) or ( a9876a );
 a9883a <=( a813a ) or ( a814a );
 a9886a <=( a811a ) or ( a812a );
 a9887a <=( a9886a ) or ( a9883a );
 a9888a <=( a9887a ) or ( a9880a );
 a9889a <=( a9888a ) or ( a9873a );
 a9890a <=( a9889a ) or ( a9860a );
 a9894a <=( a808a ) or ( a809a );
 a9895a <=( a810a ) or ( a9894a );
 a9898a <=( a806a ) or ( a807a );
 a9901a <=( a804a ) or ( a805a );
 a9902a <=( a9901a ) or ( a9898a );
 a9903a <=( a9902a ) or ( a9895a );
 a9906a <=( a802a ) or ( a803a );
 a9909a <=( a800a ) or ( a801a );
 a9910a <=( a9909a ) or ( a9906a );
 a9913a <=( a798a ) or ( a799a );
 a9916a <=( a796a ) or ( a797a );
 a9917a <=( a9916a ) or ( a9913a );
 a9918a <=( a9917a ) or ( a9910a );
 a9919a <=( a9918a ) or ( a9903a );
 a9923a <=( a793a ) or ( a794a );
 a9924a <=( a795a ) or ( a9923a );
 a9927a <=( a791a ) or ( a792a );
 a9930a <=( a789a ) or ( a790a );
 a9931a <=( a9930a ) or ( a9927a );
 a9932a <=( a9931a ) or ( a9924a );
 a9935a <=( a787a ) or ( a788a );
 a9938a <=( a785a ) or ( a786a );
 a9939a <=( a9938a ) or ( a9935a );
 a9942a <=( a783a ) or ( a784a );
 a9945a <=( a781a ) or ( a782a );
 a9946a <=( a9945a ) or ( a9942a );
 a9947a <=( a9946a ) or ( a9939a );
 a9948a <=( a9947a ) or ( a9932a );
 a9949a <=( a9948a ) or ( a9919a );
 a9950a <=( a9949a ) or ( a9890a );
 a9954a <=( a778a ) or ( a779a );
 a9955a <=( a780a ) or ( a9954a );
 a9958a <=( a776a ) or ( a777a );
 a9961a <=( a774a ) or ( a775a );
 a9962a <=( a9961a ) or ( a9958a );
 a9963a <=( a9962a ) or ( a9955a );
 a9966a <=( a772a ) or ( a773a );
 a9969a <=( a770a ) or ( a771a );
 a9970a <=( a9969a ) or ( a9966a );
 a9973a <=( a768a ) or ( a769a );
 a9976a <=( a766a ) or ( a767a );
 a9977a <=( a9976a ) or ( a9973a );
 a9978a <=( a9977a ) or ( a9970a );
 a9979a <=( a9978a ) or ( a9963a );
 a9983a <=( a763a ) or ( a764a );
 a9984a <=( a765a ) or ( a9983a );
 a9987a <=( a761a ) or ( a762a );
 a9990a <=( a759a ) or ( a760a );
 a9991a <=( a9990a ) or ( a9987a );
 a9992a <=( a9991a ) or ( a9984a );
 a9995a <=( a757a ) or ( a758a );
 a9998a <=( a755a ) or ( a756a );
 a9999a <=( a9998a ) or ( a9995a );
 a10002a <=( a753a ) or ( a754a );
 a10005a <=( a751a ) or ( a752a );
 a10006a <=( a10005a ) or ( a10002a );
 a10007a <=( a10006a ) or ( a9999a );
 a10008a <=( a10007a ) or ( a9992a );
 a10009a <=( a10008a ) or ( a9979a );
 a10013a <=( a748a ) or ( a749a );
 a10014a <=( a750a ) or ( a10013a );
 a10017a <=( a746a ) or ( a747a );
 a10020a <=( a744a ) or ( a745a );
 a10021a <=( a10020a ) or ( a10017a );
 a10022a <=( a10021a ) or ( a10014a );
 a10025a <=( a742a ) or ( a743a );
 a10028a <=( a740a ) or ( a741a );
 a10029a <=( a10028a ) or ( a10025a );
 a10032a <=( a738a ) or ( a739a );
 a10035a <=( a736a ) or ( a737a );
 a10036a <=( a10035a ) or ( a10032a );
 a10037a <=( a10036a ) or ( a10029a );
 a10038a <=( a10037a ) or ( a10022a );
 a10042a <=( a733a ) or ( a734a );
 a10043a <=( a735a ) or ( a10042a );
 a10046a <=( a731a ) or ( a732a );
 a10049a <=( a729a ) or ( a730a );
 a10050a <=( a10049a ) or ( a10046a );
 a10051a <=( a10050a ) or ( a10043a );
 a10054a <=( a727a ) or ( a728a );
 a10057a <=( a725a ) or ( a726a );
 a10058a <=( a10057a ) or ( a10054a );
 a10061a <=( a723a ) or ( a724a );
 a10064a <=( a721a ) or ( a722a );
 a10065a <=( a10064a ) or ( a10061a );
 a10066a <=( a10065a ) or ( a10058a );
 a10067a <=( a10066a ) or ( a10051a );
 a10068a <=( a10067a ) or ( a10038a );
 a10069a <=( a10068a ) or ( a10009a );
 a10070a <=( a10069a ) or ( a9950a );
 a10071a <=( a10070a ) or ( a9831a );
 a10075a <=( a718a ) or ( a719a );
 a10076a <=( a720a ) or ( a10075a );
 a10079a <=( a716a ) or ( a717a );
 a10082a <=( a714a ) or ( a715a );
 a10083a <=( a10082a ) or ( a10079a );
 a10084a <=( a10083a ) or ( a10076a );
 a10087a <=( a712a ) or ( a713a );
 a10090a <=( a710a ) or ( a711a );
 a10091a <=( a10090a ) or ( a10087a );
 a10094a <=( a708a ) or ( a709a );
 a10097a <=( a706a ) or ( a707a );
 a10098a <=( a10097a ) or ( a10094a );
 a10099a <=( a10098a ) or ( a10091a );
 a10100a <=( a10099a ) or ( a10084a );
 a10104a <=( a703a ) or ( a704a );
 a10105a <=( a705a ) or ( a10104a );
 a10108a <=( a701a ) or ( a702a );
 a10111a <=( a699a ) or ( a700a );
 a10112a <=( a10111a ) or ( a10108a );
 a10113a <=( a10112a ) or ( a10105a );
 a10116a <=( a697a ) or ( a698a );
 a10119a <=( a695a ) or ( a696a );
 a10120a <=( a10119a ) or ( a10116a );
 a10123a <=( a693a ) or ( a694a );
 a10126a <=( a691a ) or ( a692a );
 a10127a <=( a10126a ) or ( a10123a );
 a10128a <=( a10127a ) or ( a10120a );
 a10129a <=( a10128a ) or ( a10113a );
 a10130a <=( a10129a ) or ( a10100a );
 a10134a <=( a688a ) or ( a689a );
 a10135a <=( a690a ) or ( a10134a );
 a10138a <=( a686a ) or ( a687a );
 a10141a <=( a684a ) or ( a685a );
 a10142a <=( a10141a ) or ( a10138a );
 a10143a <=( a10142a ) or ( a10135a );
 a10146a <=( a682a ) or ( a683a );
 a10149a <=( a680a ) or ( a681a );
 a10150a <=( a10149a ) or ( a10146a );
 a10153a <=( a678a ) or ( a679a );
 a10156a <=( a676a ) or ( a677a );
 a10157a <=( a10156a ) or ( a10153a );
 a10158a <=( a10157a ) or ( a10150a );
 a10159a <=( a10158a ) or ( a10143a );
 a10163a <=( a673a ) or ( a674a );
 a10164a <=( a675a ) or ( a10163a );
 a10167a <=( a671a ) or ( a672a );
 a10170a <=( a669a ) or ( a670a );
 a10171a <=( a10170a ) or ( a10167a );
 a10172a <=( a10171a ) or ( a10164a );
 a10175a <=( a667a ) or ( a668a );
 a10178a <=( a665a ) or ( a666a );
 a10179a <=( a10178a ) or ( a10175a );
 a10182a <=( a663a ) or ( a664a );
 a10185a <=( a661a ) or ( a662a );
 a10186a <=( a10185a ) or ( a10182a );
 a10187a <=( a10186a ) or ( a10179a );
 a10188a <=( a10187a ) or ( a10172a );
 a10189a <=( a10188a ) or ( a10159a );
 a10190a <=( a10189a ) or ( a10130a );
 a10194a <=( a658a ) or ( a659a );
 a10195a <=( a660a ) or ( a10194a );
 a10198a <=( a656a ) or ( a657a );
 a10201a <=( a654a ) or ( a655a );
 a10202a <=( a10201a ) or ( a10198a );
 a10203a <=( a10202a ) or ( a10195a );
 a10206a <=( a652a ) or ( a653a );
 a10209a <=( a650a ) or ( a651a );
 a10210a <=( a10209a ) or ( a10206a );
 a10213a <=( a648a ) or ( a649a );
 a10216a <=( a646a ) or ( a647a );
 a10217a <=( a10216a ) or ( a10213a );
 a10218a <=( a10217a ) or ( a10210a );
 a10219a <=( a10218a ) or ( a10203a );
 a10223a <=( a643a ) or ( a644a );
 a10224a <=( a645a ) or ( a10223a );
 a10227a <=( a641a ) or ( a642a );
 a10230a <=( a639a ) or ( a640a );
 a10231a <=( a10230a ) or ( a10227a );
 a10232a <=( a10231a ) or ( a10224a );
 a10235a <=( a637a ) or ( a638a );
 a10238a <=( a635a ) or ( a636a );
 a10239a <=( a10238a ) or ( a10235a );
 a10242a <=( a633a ) or ( a634a );
 a10245a <=( a631a ) or ( a632a );
 a10246a <=( a10245a ) or ( a10242a );
 a10247a <=( a10246a ) or ( a10239a );
 a10248a <=( a10247a ) or ( a10232a );
 a10249a <=( a10248a ) or ( a10219a );
 a10253a <=( a628a ) or ( a629a );
 a10254a <=( a630a ) or ( a10253a );
 a10257a <=( a626a ) or ( a627a );
 a10260a <=( a624a ) or ( a625a );
 a10261a <=( a10260a ) or ( a10257a );
 a10262a <=( a10261a ) or ( a10254a );
 a10265a <=( a622a ) or ( a623a );
 a10268a <=( a620a ) or ( a621a );
 a10269a <=( a10268a ) or ( a10265a );
 a10272a <=( a618a ) or ( a619a );
 a10275a <=( a616a ) or ( a617a );
 a10276a <=( a10275a ) or ( a10272a );
 a10277a <=( a10276a ) or ( a10269a );
 a10278a <=( a10277a ) or ( a10262a );
 a10282a <=( a613a ) or ( a614a );
 a10283a <=( a615a ) or ( a10282a );
 a10286a <=( a611a ) or ( a612a );
 a10289a <=( a609a ) or ( a610a );
 a10290a <=( a10289a ) or ( a10286a );
 a10291a <=( a10290a ) or ( a10283a );
 a10294a <=( a607a ) or ( a608a );
 a10297a <=( a605a ) or ( a606a );
 a10298a <=( a10297a ) or ( a10294a );
 a10301a <=( a603a ) or ( a604a );
 a10304a <=( a601a ) or ( a602a );
 a10305a <=( a10304a ) or ( a10301a );
 a10306a <=( a10305a ) or ( a10298a );
 a10307a <=( a10306a ) or ( a10291a );
 a10308a <=( a10307a ) or ( a10278a );
 a10309a <=( a10308a ) or ( a10249a );
 a10310a <=( a10309a ) or ( a10190a );
 a10314a <=( a598a ) or ( a599a );
 a10315a <=( a600a ) or ( a10314a );
 a10318a <=( a596a ) or ( a597a );
 a10321a <=( a594a ) or ( a595a );
 a10322a <=( a10321a ) or ( a10318a );
 a10323a <=( a10322a ) or ( a10315a );
 a10326a <=( a592a ) or ( a593a );
 a10329a <=( a590a ) or ( a591a );
 a10330a <=( a10329a ) or ( a10326a );
 a10333a <=( a588a ) or ( a589a );
 a10336a <=( a586a ) or ( a587a );
 a10337a <=( a10336a ) or ( a10333a );
 a10338a <=( a10337a ) or ( a10330a );
 a10339a <=( a10338a ) or ( a10323a );
 a10343a <=( a583a ) or ( a584a );
 a10344a <=( a585a ) or ( a10343a );
 a10347a <=( a581a ) or ( a582a );
 a10350a <=( a579a ) or ( a580a );
 a10351a <=( a10350a ) or ( a10347a );
 a10352a <=( a10351a ) or ( a10344a );
 a10355a <=( a577a ) or ( a578a );
 a10358a <=( a575a ) or ( a576a );
 a10359a <=( a10358a ) or ( a10355a );
 a10362a <=( a573a ) or ( a574a );
 a10365a <=( a571a ) or ( a572a );
 a10366a <=( a10365a ) or ( a10362a );
 a10367a <=( a10366a ) or ( a10359a );
 a10368a <=( a10367a ) or ( a10352a );
 a10369a <=( a10368a ) or ( a10339a );
 a10373a <=( a568a ) or ( a569a );
 a10374a <=( a570a ) or ( a10373a );
 a10377a <=( a566a ) or ( a567a );
 a10380a <=( a564a ) or ( a565a );
 a10381a <=( a10380a ) or ( a10377a );
 a10382a <=( a10381a ) or ( a10374a );
 a10385a <=( a562a ) or ( a563a );
 a10388a <=( a560a ) or ( a561a );
 a10389a <=( a10388a ) or ( a10385a );
 a10392a <=( a558a ) or ( a559a );
 a10395a <=( a556a ) or ( a557a );
 a10396a <=( a10395a ) or ( a10392a );
 a10397a <=( a10396a ) or ( a10389a );
 a10398a <=( a10397a ) or ( a10382a );
 a10402a <=( a553a ) or ( a554a );
 a10403a <=( a555a ) or ( a10402a );
 a10406a <=( a551a ) or ( a552a );
 a10409a <=( a549a ) or ( a550a );
 a10410a <=( a10409a ) or ( a10406a );
 a10411a <=( a10410a ) or ( a10403a );
 a10414a <=( a547a ) or ( a548a );
 a10417a <=( a545a ) or ( a546a );
 a10418a <=( a10417a ) or ( a10414a );
 a10421a <=( a543a ) or ( a544a );
 a10424a <=( a541a ) or ( a542a );
 a10425a <=( a10424a ) or ( a10421a );
 a10426a <=( a10425a ) or ( a10418a );
 a10427a <=( a10426a ) or ( a10411a );
 a10428a <=( a10427a ) or ( a10398a );
 a10429a <=( a10428a ) or ( a10369a );
 a10433a <=( a538a ) or ( a539a );
 a10434a <=( a540a ) or ( a10433a );
 a10437a <=( a536a ) or ( a537a );
 a10440a <=( a534a ) or ( a535a );
 a10441a <=( a10440a ) or ( a10437a );
 a10442a <=( a10441a ) or ( a10434a );
 a10445a <=( a532a ) or ( a533a );
 a10448a <=( a530a ) or ( a531a );
 a10449a <=( a10448a ) or ( a10445a );
 a10452a <=( a528a ) or ( a529a );
 a10455a <=( a526a ) or ( a527a );
 a10456a <=( a10455a ) or ( a10452a );
 a10457a <=( a10456a ) or ( a10449a );
 a10458a <=( a10457a ) or ( a10442a );
 a10462a <=( a523a ) or ( a524a );
 a10463a <=( a525a ) or ( a10462a );
 a10466a <=( a521a ) or ( a522a );
 a10469a <=( a519a ) or ( a520a );
 a10470a <=( a10469a ) or ( a10466a );
 a10471a <=( a10470a ) or ( a10463a );
 a10474a <=( a517a ) or ( a518a );
 a10477a <=( a515a ) or ( a516a );
 a10478a <=( a10477a ) or ( a10474a );
 a10481a <=( a513a ) or ( a514a );
 a10484a <=( a511a ) or ( a512a );
 a10485a <=( a10484a ) or ( a10481a );
 a10486a <=( a10485a ) or ( a10478a );
 a10487a <=( a10486a ) or ( a10471a );
 a10488a <=( a10487a ) or ( a10458a );
 a10492a <=( a508a ) or ( a509a );
 a10493a <=( a510a ) or ( a10492a );
 a10496a <=( a506a ) or ( a507a );
 a10499a <=( a504a ) or ( a505a );
 a10500a <=( a10499a ) or ( a10496a );
 a10501a <=( a10500a ) or ( a10493a );
 a10504a <=( a502a ) or ( a503a );
 a10507a <=( a500a ) or ( a501a );
 a10508a <=( a10507a ) or ( a10504a );
 a10511a <=( a498a ) or ( a499a );
 a10514a <=( a496a ) or ( a497a );
 a10515a <=( a10514a ) or ( a10511a );
 a10516a <=( a10515a ) or ( a10508a );
 a10517a <=( a10516a ) or ( a10501a );
 a10521a <=( a493a ) or ( a494a );
 a10522a <=( a495a ) or ( a10521a );
 a10525a <=( a491a ) or ( a492a );
 a10528a <=( a489a ) or ( a490a );
 a10529a <=( a10528a ) or ( a10525a );
 a10530a <=( a10529a ) or ( a10522a );
 a10533a <=( a487a ) or ( a488a );
 a10536a <=( a485a ) or ( a486a );
 a10537a <=( a10536a ) or ( a10533a );
 a10540a <=( a483a ) or ( a484a );
 a10543a <=( a481a ) or ( a482a );
 a10544a <=( a10543a ) or ( a10540a );
 a10545a <=( a10544a ) or ( a10537a );
 a10546a <=( a10545a ) or ( a10530a );
 a10547a <=( a10546a ) or ( a10517a );
 a10548a <=( a10547a ) or ( a10488a );
 a10549a <=( a10548a ) or ( a10429a );
 a10550a <=( a10549a ) or ( a10310a );
 a10551a <=( a10550a ) or ( a10071a );
 a10555a <=( a478a ) or ( a479a );
 a10556a <=( a480a ) or ( a10555a );
 a10559a <=( a476a ) or ( a477a );
 a10562a <=( a474a ) or ( a475a );
 a10563a <=( a10562a ) or ( a10559a );
 a10564a <=( a10563a ) or ( a10556a );
 a10567a <=( a472a ) or ( a473a );
 a10570a <=( a470a ) or ( a471a );
 a10571a <=( a10570a ) or ( a10567a );
 a10574a <=( a468a ) or ( a469a );
 a10577a <=( a466a ) or ( a467a );
 a10578a <=( a10577a ) or ( a10574a );
 a10579a <=( a10578a ) or ( a10571a );
 a10580a <=( a10579a ) or ( a10564a );
 a10584a <=( a463a ) or ( a464a );
 a10585a <=( a465a ) or ( a10584a );
 a10588a <=( a461a ) or ( a462a );
 a10591a <=( a459a ) or ( a460a );
 a10592a <=( a10591a ) or ( a10588a );
 a10593a <=( a10592a ) or ( a10585a );
 a10596a <=( a457a ) or ( a458a );
 a10599a <=( a455a ) or ( a456a );
 a10600a <=( a10599a ) or ( a10596a );
 a10603a <=( a453a ) or ( a454a );
 a10606a <=( a451a ) or ( a452a );
 a10607a <=( a10606a ) or ( a10603a );
 a10608a <=( a10607a ) or ( a10600a );
 a10609a <=( a10608a ) or ( a10593a );
 a10610a <=( a10609a ) or ( a10580a );
 a10614a <=( a448a ) or ( a449a );
 a10615a <=( a450a ) or ( a10614a );
 a10618a <=( a446a ) or ( a447a );
 a10621a <=( a444a ) or ( a445a );
 a10622a <=( a10621a ) or ( a10618a );
 a10623a <=( a10622a ) or ( a10615a );
 a10626a <=( a442a ) or ( a443a );
 a10629a <=( a440a ) or ( a441a );
 a10630a <=( a10629a ) or ( a10626a );
 a10633a <=( a438a ) or ( a439a );
 a10636a <=( a436a ) or ( a437a );
 a10637a <=( a10636a ) or ( a10633a );
 a10638a <=( a10637a ) or ( a10630a );
 a10639a <=( a10638a ) or ( a10623a );
 a10643a <=( a433a ) or ( a434a );
 a10644a <=( a435a ) or ( a10643a );
 a10647a <=( a431a ) or ( a432a );
 a10650a <=( a429a ) or ( a430a );
 a10651a <=( a10650a ) or ( a10647a );
 a10652a <=( a10651a ) or ( a10644a );
 a10655a <=( a427a ) or ( a428a );
 a10658a <=( a425a ) or ( a426a );
 a10659a <=( a10658a ) or ( a10655a );
 a10662a <=( a423a ) or ( a424a );
 a10665a <=( a421a ) or ( a422a );
 a10666a <=( a10665a ) or ( a10662a );
 a10667a <=( a10666a ) or ( a10659a );
 a10668a <=( a10667a ) or ( a10652a );
 a10669a <=( a10668a ) or ( a10639a );
 a10670a <=( a10669a ) or ( a10610a );
 a10674a <=( a418a ) or ( a419a );
 a10675a <=( a420a ) or ( a10674a );
 a10678a <=( a416a ) or ( a417a );
 a10681a <=( a414a ) or ( a415a );
 a10682a <=( a10681a ) or ( a10678a );
 a10683a <=( a10682a ) or ( a10675a );
 a10686a <=( a412a ) or ( a413a );
 a10689a <=( a410a ) or ( a411a );
 a10690a <=( a10689a ) or ( a10686a );
 a10693a <=( a408a ) or ( a409a );
 a10696a <=( a406a ) or ( a407a );
 a10697a <=( a10696a ) or ( a10693a );
 a10698a <=( a10697a ) or ( a10690a );
 a10699a <=( a10698a ) or ( a10683a );
 a10703a <=( a403a ) or ( a404a );
 a10704a <=( a405a ) or ( a10703a );
 a10707a <=( a401a ) or ( a402a );
 a10710a <=( a399a ) or ( a400a );
 a10711a <=( a10710a ) or ( a10707a );
 a10712a <=( a10711a ) or ( a10704a );
 a10715a <=( a397a ) or ( a398a );
 a10718a <=( a395a ) or ( a396a );
 a10719a <=( a10718a ) or ( a10715a );
 a10722a <=( a393a ) or ( a394a );
 a10725a <=( a391a ) or ( a392a );
 a10726a <=( a10725a ) or ( a10722a );
 a10727a <=( a10726a ) or ( a10719a );
 a10728a <=( a10727a ) or ( a10712a );
 a10729a <=( a10728a ) or ( a10699a );
 a10733a <=( a388a ) or ( a389a );
 a10734a <=( a390a ) or ( a10733a );
 a10737a <=( a386a ) or ( a387a );
 a10740a <=( a384a ) or ( a385a );
 a10741a <=( a10740a ) or ( a10737a );
 a10742a <=( a10741a ) or ( a10734a );
 a10745a <=( a382a ) or ( a383a );
 a10748a <=( a380a ) or ( a381a );
 a10749a <=( a10748a ) or ( a10745a );
 a10752a <=( a378a ) or ( a379a );
 a10755a <=( a376a ) or ( a377a );
 a10756a <=( a10755a ) or ( a10752a );
 a10757a <=( a10756a ) or ( a10749a );
 a10758a <=( a10757a ) or ( a10742a );
 a10762a <=( a373a ) or ( a374a );
 a10763a <=( a375a ) or ( a10762a );
 a10766a <=( a371a ) or ( a372a );
 a10769a <=( a369a ) or ( a370a );
 a10770a <=( a10769a ) or ( a10766a );
 a10771a <=( a10770a ) or ( a10763a );
 a10774a <=( a367a ) or ( a368a );
 a10777a <=( a365a ) or ( a366a );
 a10778a <=( a10777a ) or ( a10774a );
 a10781a <=( a363a ) or ( a364a );
 a10784a <=( a361a ) or ( a362a );
 a10785a <=( a10784a ) or ( a10781a );
 a10786a <=( a10785a ) or ( a10778a );
 a10787a <=( a10786a ) or ( a10771a );
 a10788a <=( a10787a ) or ( a10758a );
 a10789a <=( a10788a ) or ( a10729a );
 a10790a <=( a10789a ) or ( a10670a );
 a10794a <=( a358a ) or ( a359a );
 a10795a <=( a360a ) or ( a10794a );
 a10798a <=( a356a ) or ( a357a );
 a10801a <=( a354a ) or ( a355a );
 a10802a <=( a10801a ) or ( a10798a );
 a10803a <=( a10802a ) or ( a10795a );
 a10806a <=( a352a ) or ( a353a );
 a10809a <=( a350a ) or ( a351a );
 a10810a <=( a10809a ) or ( a10806a );
 a10813a <=( a348a ) or ( a349a );
 a10816a <=( a346a ) or ( a347a );
 a10817a <=( a10816a ) or ( a10813a );
 a10818a <=( a10817a ) or ( a10810a );
 a10819a <=( a10818a ) or ( a10803a );
 a10823a <=( a343a ) or ( a344a );
 a10824a <=( a345a ) or ( a10823a );
 a10827a <=( a341a ) or ( a342a );
 a10830a <=( a339a ) or ( a340a );
 a10831a <=( a10830a ) or ( a10827a );
 a10832a <=( a10831a ) or ( a10824a );
 a10835a <=( a337a ) or ( a338a );
 a10838a <=( a335a ) or ( a336a );
 a10839a <=( a10838a ) or ( a10835a );
 a10842a <=( a333a ) or ( a334a );
 a10845a <=( a331a ) or ( a332a );
 a10846a <=( a10845a ) or ( a10842a );
 a10847a <=( a10846a ) or ( a10839a );
 a10848a <=( a10847a ) or ( a10832a );
 a10849a <=( a10848a ) or ( a10819a );
 a10853a <=( a328a ) or ( a329a );
 a10854a <=( a330a ) or ( a10853a );
 a10857a <=( a326a ) or ( a327a );
 a10860a <=( a324a ) or ( a325a );
 a10861a <=( a10860a ) or ( a10857a );
 a10862a <=( a10861a ) or ( a10854a );
 a10865a <=( a322a ) or ( a323a );
 a10868a <=( a320a ) or ( a321a );
 a10869a <=( a10868a ) or ( a10865a );
 a10872a <=( a318a ) or ( a319a );
 a10875a <=( a316a ) or ( a317a );
 a10876a <=( a10875a ) or ( a10872a );
 a10877a <=( a10876a ) or ( a10869a );
 a10878a <=( a10877a ) or ( a10862a );
 a10882a <=( a313a ) or ( a314a );
 a10883a <=( a315a ) or ( a10882a );
 a10886a <=( a311a ) or ( a312a );
 a10889a <=( a309a ) or ( a310a );
 a10890a <=( a10889a ) or ( a10886a );
 a10891a <=( a10890a ) or ( a10883a );
 a10894a <=( a307a ) or ( a308a );
 a10897a <=( a305a ) or ( a306a );
 a10898a <=( a10897a ) or ( a10894a );
 a10901a <=( a303a ) or ( a304a );
 a10904a <=( a301a ) or ( a302a );
 a10905a <=( a10904a ) or ( a10901a );
 a10906a <=( a10905a ) or ( a10898a );
 a10907a <=( a10906a ) or ( a10891a );
 a10908a <=( a10907a ) or ( a10878a );
 a10909a <=( a10908a ) or ( a10849a );
 a10913a <=( a298a ) or ( a299a );
 a10914a <=( a300a ) or ( a10913a );
 a10917a <=( a296a ) or ( a297a );
 a10920a <=( a294a ) or ( a295a );
 a10921a <=( a10920a ) or ( a10917a );
 a10922a <=( a10921a ) or ( a10914a );
 a10925a <=( a292a ) or ( a293a );
 a10928a <=( a290a ) or ( a291a );
 a10929a <=( a10928a ) or ( a10925a );
 a10932a <=( a288a ) or ( a289a );
 a10935a <=( a286a ) or ( a287a );
 a10936a <=( a10935a ) or ( a10932a );
 a10937a <=( a10936a ) or ( a10929a );
 a10938a <=( a10937a ) or ( a10922a );
 a10942a <=( a283a ) or ( a284a );
 a10943a <=( a285a ) or ( a10942a );
 a10946a <=( a281a ) or ( a282a );
 a10949a <=( a279a ) or ( a280a );
 a10950a <=( a10949a ) or ( a10946a );
 a10951a <=( a10950a ) or ( a10943a );
 a10954a <=( a277a ) or ( a278a );
 a10957a <=( a275a ) or ( a276a );
 a10958a <=( a10957a ) or ( a10954a );
 a10961a <=( a273a ) or ( a274a );
 a10964a <=( a271a ) or ( a272a );
 a10965a <=( a10964a ) or ( a10961a );
 a10966a <=( a10965a ) or ( a10958a );
 a10967a <=( a10966a ) or ( a10951a );
 a10968a <=( a10967a ) or ( a10938a );
 a10972a <=( a268a ) or ( a269a );
 a10973a <=( a270a ) or ( a10972a );
 a10976a <=( a266a ) or ( a267a );
 a10979a <=( a264a ) or ( a265a );
 a10980a <=( a10979a ) or ( a10976a );
 a10981a <=( a10980a ) or ( a10973a );
 a10984a <=( a262a ) or ( a263a );
 a10987a <=( a260a ) or ( a261a );
 a10988a <=( a10987a ) or ( a10984a );
 a10991a <=( a258a ) or ( a259a );
 a10994a <=( a256a ) or ( a257a );
 a10995a <=( a10994a ) or ( a10991a );
 a10996a <=( a10995a ) or ( a10988a );
 a10997a <=( a10996a ) or ( a10981a );
 a11001a <=( a253a ) or ( a254a );
 a11002a <=( a255a ) or ( a11001a );
 a11005a <=( a251a ) or ( a252a );
 a11008a <=( a249a ) or ( a250a );
 a11009a <=( a11008a ) or ( a11005a );
 a11010a <=( a11009a ) or ( a11002a );
 a11013a <=( a247a ) or ( a248a );
 a11016a <=( a245a ) or ( a246a );
 a11017a <=( a11016a ) or ( a11013a );
 a11020a <=( a243a ) or ( a244a );
 a11023a <=( a241a ) or ( a242a );
 a11024a <=( a11023a ) or ( a11020a );
 a11025a <=( a11024a ) or ( a11017a );
 a11026a <=( a11025a ) or ( a11010a );
 a11027a <=( a11026a ) or ( a10997a );
 a11028a <=( a11027a ) or ( a10968a );
 a11029a <=( a11028a ) or ( a10909a );
 a11030a <=( a11029a ) or ( a10790a );
 a11034a <=( a238a ) or ( a239a );
 a11035a <=( a240a ) or ( a11034a );
 a11038a <=( a236a ) or ( a237a );
 a11041a <=( a234a ) or ( a235a );
 a11042a <=( a11041a ) or ( a11038a );
 a11043a <=( a11042a ) or ( a11035a );
 a11046a <=( a232a ) or ( a233a );
 a11049a <=( a230a ) or ( a231a );
 a11050a <=( a11049a ) or ( a11046a );
 a11053a <=( a228a ) or ( a229a );
 a11056a <=( a226a ) or ( a227a );
 a11057a <=( a11056a ) or ( a11053a );
 a11058a <=( a11057a ) or ( a11050a );
 a11059a <=( a11058a ) or ( a11043a );
 a11063a <=( a223a ) or ( a224a );
 a11064a <=( a225a ) or ( a11063a );
 a11067a <=( a221a ) or ( a222a );
 a11070a <=( a219a ) or ( a220a );
 a11071a <=( a11070a ) or ( a11067a );
 a11072a <=( a11071a ) or ( a11064a );
 a11075a <=( a217a ) or ( a218a );
 a11078a <=( a215a ) or ( a216a );
 a11079a <=( a11078a ) or ( a11075a );
 a11082a <=( a213a ) or ( a214a );
 a11085a <=( a211a ) or ( a212a );
 a11086a <=( a11085a ) or ( a11082a );
 a11087a <=( a11086a ) or ( a11079a );
 a11088a <=( a11087a ) or ( a11072a );
 a11089a <=( a11088a ) or ( a11059a );
 a11093a <=( a208a ) or ( a209a );
 a11094a <=( a210a ) or ( a11093a );
 a11097a <=( a206a ) or ( a207a );
 a11100a <=( a204a ) or ( a205a );
 a11101a <=( a11100a ) or ( a11097a );
 a11102a <=( a11101a ) or ( a11094a );
 a11105a <=( a202a ) or ( a203a );
 a11108a <=( a200a ) or ( a201a );
 a11109a <=( a11108a ) or ( a11105a );
 a11112a <=( a198a ) or ( a199a );
 a11115a <=( a196a ) or ( a197a );
 a11116a <=( a11115a ) or ( a11112a );
 a11117a <=( a11116a ) or ( a11109a );
 a11118a <=( a11117a ) or ( a11102a );
 a11122a <=( a193a ) or ( a194a );
 a11123a <=( a195a ) or ( a11122a );
 a11126a <=( a191a ) or ( a192a );
 a11129a <=( a189a ) or ( a190a );
 a11130a <=( a11129a ) or ( a11126a );
 a11131a <=( a11130a ) or ( a11123a );
 a11134a <=( a187a ) or ( a188a );
 a11137a <=( a185a ) or ( a186a );
 a11138a <=( a11137a ) or ( a11134a );
 a11141a <=( a183a ) or ( a184a );
 a11144a <=( a181a ) or ( a182a );
 a11145a <=( a11144a ) or ( a11141a );
 a11146a <=( a11145a ) or ( a11138a );
 a11147a <=( a11146a ) or ( a11131a );
 a11148a <=( a11147a ) or ( a11118a );
 a11149a <=( a11148a ) or ( a11089a );
 a11153a <=( a178a ) or ( a179a );
 a11154a <=( a180a ) or ( a11153a );
 a11157a <=( a176a ) or ( a177a );
 a11160a <=( a174a ) or ( a175a );
 a11161a <=( a11160a ) or ( a11157a );
 a11162a <=( a11161a ) or ( a11154a );
 a11165a <=( a172a ) or ( a173a );
 a11168a <=( a170a ) or ( a171a );
 a11169a <=( a11168a ) or ( a11165a );
 a11172a <=( a168a ) or ( a169a );
 a11175a <=( a166a ) or ( a167a );
 a11176a <=( a11175a ) or ( a11172a );
 a11177a <=( a11176a ) or ( a11169a );
 a11178a <=( a11177a ) or ( a11162a );
 a11182a <=( a163a ) or ( a164a );
 a11183a <=( a165a ) or ( a11182a );
 a11186a <=( a161a ) or ( a162a );
 a11189a <=( a159a ) or ( a160a );
 a11190a <=( a11189a ) or ( a11186a );
 a11191a <=( a11190a ) or ( a11183a );
 a11194a <=( a157a ) or ( a158a );
 a11197a <=( a155a ) or ( a156a );
 a11198a <=( a11197a ) or ( a11194a );
 a11201a <=( a153a ) or ( a154a );
 a11204a <=( a151a ) or ( a152a );
 a11205a <=( a11204a ) or ( a11201a );
 a11206a <=( a11205a ) or ( a11198a );
 a11207a <=( a11206a ) or ( a11191a );
 a11208a <=( a11207a ) or ( a11178a );
 a11212a <=( a148a ) or ( a149a );
 a11213a <=( a150a ) or ( a11212a );
 a11216a <=( a146a ) or ( a147a );
 a11219a <=( a144a ) or ( a145a );
 a11220a <=( a11219a ) or ( a11216a );
 a11221a <=( a11220a ) or ( a11213a );
 a11224a <=( a142a ) or ( a143a );
 a11227a <=( a140a ) or ( a141a );
 a11228a <=( a11227a ) or ( a11224a );
 a11231a <=( a138a ) or ( a139a );
 a11234a <=( a136a ) or ( a137a );
 a11235a <=( a11234a ) or ( a11231a );
 a11236a <=( a11235a ) or ( a11228a );
 a11237a <=( a11236a ) or ( a11221a );
 a11241a <=( a133a ) or ( a134a );
 a11242a <=( a135a ) or ( a11241a );
 a11245a <=( a131a ) or ( a132a );
 a11248a <=( a129a ) or ( a130a );
 a11249a <=( a11248a ) or ( a11245a );
 a11250a <=( a11249a ) or ( a11242a );
 a11253a <=( a127a ) or ( a128a );
 a11256a <=( a125a ) or ( a126a );
 a11257a <=( a11256a ) or ( a11253a );
 a11260a <=( a123a ) or ( a124a );
 a11263a <=( a121a ) or ( a122a );
 a11264a <=( a11263a ) or ( a11260a );
 a11265a <=( a11264a ) or ( a11257a );
 a11266a <=( a11265a ) or ( a11250a );
 a11267a <=( a11266a ) or ( a11237a );
 a11268a <=( a11267a ) or ( a11208a );
 a11269a <=( a11268a ) or ( a11149a );
 a11273a <=( a118a ) or ( a119a );
 a11274a <=( a120a ) or ( a11273a );
 a11277a <=( a116a ) or ( a117a );
 a11280a <=( a114a ) or ( a115a );
 a11281a <=( a11280a ) or ( a11277a );
 a11282a <=( a11281a ) or ( a11274a );
 a11285a <=( a112a ) or ( a113a );
 a11288a <=( a110a ) or ( a111a );
 a11289a <=( a11288a ) or ( a11285a );
 a11292a <=( a108a ) or ( a109a );
 a11295a <=( a106a ) or ( a107a );
 a11296a <=( a11295a ) or ( a11292a );
 a11297a <=( a11296a ) or ( a11289a );
 a11298a <=( a11297a ) or ( a11282a );
 a11302a <=( a103a ) or ( a104a );
 a11303a <=( a105a ) or ( a11302a );
 a11306a <=( a101a ) or ( a102a );
 a11309a <=( a99a ) or ( a100a );
 a11310a <=( a11309a ) or ( a11306a );
 a11311a <=( a11310a ) or ( a11303a );
 a11314a <=( a97a ) or ( a98a );
 a11317a <=( a95a ) or ( a96a );
 a11318a <=( a11317a ) or ( a11314a );
 a11321a <=( a93a ) or ( a94a );
 a11324a <=( a91a ) or ( a92a );
 a11325a <=( a11324a ) or ( a11321a );
 a11326a <=( a11325a ) or ( a11318a );
 a11327a <=( a11326a ) or ( a11311a );
 a11328a <=( a11327a ) or ( a11298a );
 a11332a <=( a88a ) or ( a89a );
 a11333a <=( a90a ) or ( a11332a );
 a11336a <=( a86a ) or ( a87a );
 a11339a <=( a84a ) or ( a85a );
 a11340a <=( a11339a ) or ( a11336a );
 a11341a <=( a11340a ) or ( a11333a );
 a11344a <=( a82a ) or ( a83a );
 a11347a <=( a80a ) or ( a81a );
 a11348a <=( a11347a ) or ( a11344a );
 a11351a <=( a78a ) or ( a79a );
 a11354a <=( a76a ) or ( a77a );
 a11355a <=( a11354a ) or ( a11351a );
 a11356a <=( a11355a ) or ( a11348a );
 a11357a <=( a11356a ) or ( a11341a );
 a11361a <=( a73a ) or ( a74a );
 a11362a <=( a75a ) or ( a11361a );
 a11365a <=( a71a ) or ( a72a );
 a11368a <=( a69a ) or ( a70a );
 a11369a <=( a11368a ) or ( a11365a );
 a11370a <=( a11369a ) or ( a11362a );
 a11373a <=( a67a ) or ( a68a );
 a11376a <=( a65a ) or ( a66a );
 a11377a <=( a11376a ) or ( a11373a );
 a11380a <=( a63a ) or ( a64a );
 a11383a <=( a61a ) or ( a62a );
 a11384a <=( a11383a ) or ( a11380a );
 a11385a <=( a11384a ) or ( a11377a );
 a11386a <=( a11385a ) or ( a11370a );
 a11387a <=( a11386a ) or ( a11357a );
 a11388a <=( a11387a ) or ( a11328a );
 a11392a <=( a58a ) or ( a59a );
 a11393a <=( a60a ) or ( a11392a );
 a11396a <=( a56a ) or ( a57a );
 a11399a <=( a54a ) or ( a55a );
 a11400a <=( a11399a ) or ( a11396a );
 a11401a <=( a11400a ) or ( a11393a );
 a11404a <=( a52a ) or ( a53a );
 a11407a <=( a50a ) or ( a51a );
 a11408a <=( a11407a ) or ( a11404a );
 a11411a <=( a48a ) or ( a49a );
 a11414a <=( a46a ) or ( a47a );
 a11415a <=( a11414a ) or ( a11411a );
 a11416a <=( a11415a ) or ( a11408a );
 a11417a <=( a11416a ) or ( a11401a );
 a11421a <=( a43a ) or ( a44a );
 a11422a <=( a45a ) or ( a11421a );
 a11425a <=( a41a ) or ( a42a );
 a11428a <=( a39a ) or ( a40a );
 a11429a <=( a11428a ) or ( a11425a );
 a11430a <=( a11429a ) or ( a11422a );
 a11433a <=( a37a ) or ( a38a );
 a11436a <=( a35a ) or ( a36a );
 a11437a <=( a11436a ) or ( a11433a );
 a11440a <=( a33a ) or ( a34a );
 a11443a <=( a31a ) or ( a32a );
 a11444a <=( a11443a ) or ( a11440a );
 a11445a <=( a11444a ) or ( a11437a );
 a11446a <=( a11445a ) or ( a11430a );
 a11447a <=( a11446a ) or ( a11417a );
 a11451a <=( a28a ) or ( a29a );
 a11452a <=( a30a ) or ( a11451a );
 a11455a <=( a26a ) or ( a27a );
 a11458a <=( a24a ) or ( a25a );
 a11459a <=( a11458a ) or ( a11455a );
 a11460a <=( a11459a ) or ( a11452a );
 a11463a <=( a22a ) or ( a23a );
 a11466a <=( a20a ) or ( a21a );
 a11467a <=( a11466a ) or ( a11463a );
 a11470a <=( a18a ) or ( a19a );
 a11473a <=( a16a ) or ( a17a );
 a11474a <=( a11473a ) or ( a11470a );
 a11475a <=( a11474a ) or ( a11467a );
 a11476a <=( a11475a ) or ( a11460a );
 a11480a <=( a13a ) or ( a14a );
 a11481a <=( a15a ) or ( a11480a );
 a11484a <=( a11a ) or ( a12a );
 a11487a <=( a9a ) or ( a10a );
 a11488a <=( a11487a ) or ( a11484a );
 a11489a <=( a11488a ) or ( a11481a );
 a11492a <=( a7a ) or ( a8a );
 a11495a <=( a5a ) or ( a6a );
 a11496a <=( a11495a ) or ( a11492a );
 a11499a <=( a3a ) or ( a4a );
 a11502a <=( a1a ) or ( a2a );
 a11503a <=( a11502a ) or ( a11499a );
 a11504a <=( a11503a ) or ( a11496a );
 a11505a <=( a11504a ) or ( a11489a );
 a11506a <=( a11505a ) or ( a11476a );
 a11507a <=( a11506a ) or ( a11447a );
 a11508a <=( a11507a ) or ( a11388a );
 a11509a <=( a11508a ) or ( a11269a );
 a11510a <=( a11509a ) or ( a11030a );
 a11511a <=( a11510a ) or ( a10551a );
 a11512a <=( a11511a ) or ( a9592a );
 a11515a <=( A233  and  (not A232) );
 a11518a <=( A235  and  A234 );
 a11519a <=( a11518a  and  a11515a );
 a11522a <=( (not A299)  and  A298 );
 a11525a <=( A301  and  A300 );
 a11526a <=( a11525a  and  a11522a );
 a11529a <=( A233  and  (not A232) );
 a11532a <=( A235  and  A234 );
 a11533a <=( a11532a  and  a11529a );
 a11536a <=( (not A299)  and  A298 );
 a11539a <=( (not A302)  and  A300 );
 a11540a <=( a11539a  and  a11536a );
 a11543a <=( A233  and  (not A232) );
 a11546a <=( A235  and  A234 );
 a11547a <=( a11546a  and  a11543a );
 a11550a <=( A299  and  (not A298) );
 a11553a <=( A301  and  A300 );
 a11554a <=( a11553a  and  a11550a );
 a11557a <=( A233  and  (not A232) );
 a11560a <=( A235  and  A234 );
 a11561a <=( a11560a  and  a11557a );
 a11564a <=( A299  and  (not A298) );
 a11567a <=( (not A302)  and  A300 );
 a11568a <=( a11567a  and  a11564a );
 a11571a <=( A233  and  (not A232) );
 a11574a <=( A235  and  A234 );
 a11575a <=( a11574a  and  a11571a );
 a11578a <=( A266  and  (not A265) );
 a11581a <=( A268  and  A267 );
 a11582a <=( a11581a  and  a11578a );
 a11585a <=( A233  and  (not A232) );
 a11588a <=( A235  and  A234 );
 a11589a <=( a11588a  and  a11585a );
 a11592a <=( A266  and  (not A265) );
 a11595a <=( (not A269)  and  A267 );
 a11596a <=( a11595a  and  a11592a );
 a11599a <=( A233  and  (not A232) );
 a11602a <=( A235  and  A234 );
 a11603a <=( a11602a  and  a11599a );
 a11606a <=( (not A266)  and  A265 );
 a11609a <=( A268  and  A267 );
 a11610a <=( a11609a  and  a11606a );
 a11613a <=( A233  and  (not A232) );
 a11616a <=( A235  and  A234 );
 a11617a <=( a11616a  and  a11613a );
 a11620a <=( (not A266)  and  A265 );
 a11623a <=( (not A269)  and  A267 );
 a11624a <=( a11623a  and  a11620a );
 a11627a <=( A233  and  (not A232) );
 a11630a <=( (not A236)  and  A234 );
 a11631a <=( a11630a  and  a11627a );
 a11634a <=( (not A299)  and  A298 );
 a11637a <=( A301  and  A300 );
 a11638a <=( a11637a  and  a11634a );
 a11641a <=( A233  and  (not A232) );
 a11644a <=( (not A236)  and  A234 );
 a11645a <=( a11644a  and  a11641a );
 a11648a <=( (not A299)  and  A298 );
 a11651a <=( (not A302)  and  A300 );
 a11652a <=( a11651a  and  a11648a );
 a11655a <=( A233  and  (not A232) );
 a11658a <=( (not A236)  and  A234 );
 a11659a <=( a11658a  and  a11655a );
 a11662a <=( A299  and  (not A298) );
 a11665a <=( A301  and  A300 );
 a11666a <=( a11665a  and  a11662a );
 a11669a <=( A233  and  (not A232) );
 a11672a <=( (not A236)  and  A234 );
 a11673a <=( a11672a  and  a11669a );
 a11676a <=( A299  and  (not A298) );
 a11679a <=( (not A302)  and  A300 );
 a11680a <=( a11679a  and  a11676a );
 a11683a <=( A233  and  (not A232) );
 a11686a <=( (not A236)  and  A234 );
 a11687a <=( a11686a  and  a11683a );
 a11690a <=( A266  and  (not A265) );
 a11693a <=( A268  and  A267 );
 a11694a <=( a11693a  and  a11690a );
 a11697a <=( A233  and  (not A232) );
 a11700a <=( (not A236)  and  A234 );
 a11701a <=( a11700a  and  a11697a );
 a11704a <=( A266  and  (not A265) );
 a11707a <=( (not A269)  and  A267 );
 a11708a <=( a11707a  and  a11704a );
 a11711a <=( A233  and  (not A232) );
 a11714a <=( (not A236)  and  A234 );
 a11715a <=( a11714a  and  a11711a );
 a11718a <=( (not A266)  and  A265 );
 a11721a <=( A268  and  A267 );
 a11722a <=( a11721a  and  a11718a );
 a11725a <=( A233  and  (not A232) );
 a11728a <=( (not A236)  and  A234 );
 a11729a <=( a11728a  and  a11725a );
 a11732a <=( (not A266)  and  A265 );
 a11735a <=( (not A269)  and  A267 );
 a11736a <=( a11735a  and  a11732a );
 a11739a <=( (not A233)  and  A232 );
 a11742a <=( A235  and  A234 );
 a11743a <=( a11742a  and  a11739a );
 a11746a <=( (not A299)  and  A298 );
 a11749a <=( A301  and  A300 );
 a11750a <=( a11749a  and  a11746a );
 a11753a <=( (not A233)  and  A232 );
 a11756a <=( A235  and  A234 );
 a11757a <=( a11756a  and  a11753a );
 a11760a <=( (not A299)  and  A298 );
 a11763a <=( (not A302)  and  A300 );
 a11764a <=( a11763a  and  a11760a );
 a11767a <=( (not A233)  and  A232 );
 a11770a <=( A235  and  A234 );
 a11771a <=( a11770a  and  a11767a );
 a11774a <=( A299  and  (not A298) );
 a11777a <=( A301  and  A300 );
 a11778a <=( a11777a  and  a11774a );
 a11781a <=( (not A233)  and  A232 );
 a11784a <=( A235  and  A234 );
 a11785a <=( a11784a  and  a11781a );
 a11788a <=( A299  and  (not A298) );
 a11791a <=( (not A302)  and  A300 );
 a11792a <=( a11791a  and  a11788a );
 a11795a <=( (not A233)  and  A232 );
 a11798a <=( A235  and  A234 );
 a11799a <=( a11798a  and  a11795a );
 a11802a <=( A266  and  (not A265) );
 a11805a <=( A268  and  A267 );
 a11806a <=( a11805a  and  a11802a );
 a11809a <=( (not A233)  and  A232 );
 a11812a <=( A235  and  A234 );
 a11813a <=( a11812a  and  a11809a );
 a11816a <=( A266  and  (not A265) );
 a11819a <=( (not A269)  and  A267 );
 a11820a <=( a11819a  and  a11816a );
 a11823a <=( (not A233)  and  A232 );
 a11826a <=( A235  and  A234 );
 a11827a <=( a11826a  and  a11823a );
 a11830a <=( (not A266)  and  A265 );
 a11833a <=( A268  and  A267 );
 a11834a <=( a11833a  and  a11830a );
 a11837a <=( (not A233)  and  A232 );
 a11840a <=( A235  and  A234 );
 a11841a <=( a11840a  and  a11837a );
 a11844a <=( (not A266)  and  A265 );
 a11847a <=( (not A269)  and  A267 );
 a11848a <=( a11847a  and  a11844a );
 a11851a <=( (not A233)  and  A232 );
 a11854a <=( (not A236)  and  A234 );
 a11855a <=( a11854a  and  a11851a );
 a11858a <=( (not A299)  and  A298 );
 a11861a <=( A301  and  A300 );
 a11862a <=( a11861a  and  a11858a );
 a11865a <=( (not A233)  and  A232 );
 a11868a <=( (not A236)  and  A234 );
 a11869a <=( a11868a  and  a11865a );
 a11872a <=( (not A299)  and  A298 );
 a11875a <=( (not A302)  and  A300 );
 a11876a <=( a11875a  and  a11872a );
 a11879a <=( (not A233)  and  A232 );
 a11882a <=( (not A236)  and  A234 );
 a11883a <=( a11882a  and  a11879a );
 a11886a <=( A299  and  (not A298) );
 a11889a <=( A301  and  A300 );
 a11890a <=( a11889a  and  a11886a );
 a11893a <=( (not A233)  and  A232 );
 a11896a <=( (not A236)  and  A234 );
 a11897a <=( a11896a  and  a11893a );
 a11900a <=( A299  and  (not A298) );
 a11903a <=( (not A302)  and  A300 );
 a11904a <=( a11903a  and  a11900a );
 a11907a <=( (not A233)  and  A232 );
 a11910a <=( (not A236)  and  A234 );
 a11911a <=( a11910a  and  a11907a );
 a11914a <=( A266  and  (not A265) );
 a11917a <=( A268  and  A267 );
 a11918a <=( a11917a  and  a11914a );
 a11921a <=( (not A233)  and  A232 );
 a11924a <=( (not A236)  and  A234 );
 a11925a <=( a11924a  and  a11921a );
 a11928a <=( A266  and  (not A265) );
 a11931a <=( (not A269)  and  A267 );
 a11932a <=( a11931a  and  a11928a );
 a11935a <=( (not A233)  and  A232 );
 a11938a <=( (not A236)  and  A234 );
 a11939a <=( a11938a  and  a11935a );
 a11942a <=( (not A266)  and  A265 );
 a11945a <=( A268  and  A267 );
 a11946a <=( a11945a  and  a11942a );
 a11949a <=( (not A233)  and  A232 );
 a11952a <=( (not A236)  and  A234 );
 a11953a <=( a11952a  and  a11949a );
 a11956a <=( (not A266)  and  A265 );
 a11959a <=( (not A269)  and  A267 );
 a11960a <=( a11959a  and  a11956a );
 a11963a <=( A233  and  (not A232) );
 a11966a <=( A235  and  A234 );
 a11967a <=( a11966a  and  a11963a );
 a11970a <=( (not A299)  and  A298 );
 a11974a <=( A302  and  (not A301) );
 a11975a <=( (not A300)  and  a11974a );
 a11976a <=( a11975a  and  a11970a );
 a11979a <=( A233  and  (not A232) );
 a11982a <=( A235  and  A234 );
 a11983a <=( a11982a  and  a11979a );
 a11986a <=( A299  and  (not A298) );
 a11990a <=( A302  and  (not A301) );
 a11991a <=( (not A300)  and  a11990a );
 a11992a <=( a11991a  and  a11986a );
 a11995a <=( A233  and  (not A232) );
 a11998a <=( (not A236)  and  A234 );
 a11999a <=( a11998a  and  a11995a );
 a12002a <=( (not A299)  and  A298 );
 a12006a <=( A302  and  (not A301) );
 a12007a <=( (not A300)  and  a12006a );
 a12008a <=( a12007a  and  a12002a );
 a12011a <=( A233  and  (not A232) );
 a12014a <=( (not A236)  and  A234 );
 a12015a <=( a12014a  and  a12011a );
 a12018a <=( A299  and  (not A298) );
 a12022a <=( A302  and  (not A301) );
 a12023a <=( (not A300)  and  a12022a );
 a12024a <=( a12023a  and  a12018a );
 a12027a <=( A233  and  (not A232) );
 a12030a <=( (not A235)  and  (not A234) );
 a12031a <=( a12030a  and  a12027a );
 a12034a <=( A298  and  A236 );
 a12038a <=( A301  and  A300 );
 a12039a <=( (not A299)  and  a12038a );
 a12040a <=( a12039a  and  a12034a );
 a12043a <=( A233  and  (not A232) );
 a12046a <=( (not A235)  and  (not A234) );
 a12047a <=( a12046a  and  a12043a );
 a12050a <=( A298  and  A236 );
 a12054a <=( (not A302)  and  A300 );
 a12055a <=( (not A299)  and  a12054a );
 a12056a <=( a12055a  and  a12050a );
 a12059a <=( A233  and  (not A232) );
 a12062a <=( (not A235)  and  (not A234) );
 a12063a <=( a12062a  and  a12059a );
 a12066a <=( (not A298)  and  A236 );
 a12070a <=( A301  and  A300 );
 a12071a <=( A299  and  a12070a );
 a12072a <=( a12071a  and  a12066a );
 a12075a <=( A233  and  (not A232) );
 a12078a <=( (not A235)  and  (not A234) );
 a12079a <=( a12078a  and  a12075a );
 a12082a <=( (not A298)  and  A236 );
 a12086a <=( (not A302)  and  A300 );
 a12087a <=( A299  and  a12086a );
 a12088a <=( a12087a  and  a12082a );
 a12091a <=( A233  and  (not A232) );
 a12094a <=( (not A235)  and  (not A234) );
 a12095a <=( a12094a  and  a12091a );
 a12098a <=( (not A265)  and  A236 );
 a12102a <=( A268  and  A267 );
 a12103a <=( A266  and  a12102a );
 a12104a <=( a12103a  and  a12098a );
 a12107a <=( A233  and  (not A232) );
 a12110a <=( (not A235)  and  (not A234) );
 a12111a <=( a12110a  and  a12107a );
 a12114a <=( (not A265)  and  A236 );
 a12118a <=( (not A269)  and  A267 );
 a12119a <=( A266  and  a12118a );
 a12120a <=( a12119a  and  a12114a );
 a12123a <=( A233  and  (not A232) );
 a12126a <=( (not A235)  and  (not A234) );
 a12127a <=( a12126a  and  a12123a );
 a12130a <=( A265  and  A236 );
 a12134a <=( A268  and  A267 );
 a12135a <=( (not A266)  and  a12134a );
 a12136a <=( a12135a  and  a12130a );
 a12139a <=( A233  and  (not A232) );
 a12142a <=( (not A235)  and  (not A234) );
 a12143a <=( a12142a  and  a12139a );
 a12146a <=( A265  and  A236 );
 a12150a <=( (not A269)  and  A267 );
 a12151a <=( (not A266)  and  a12150a );
 a12152a <=( a12151a  and  a12146a );
 a12155a <=( (not A233)  and  A232 );
 a12158a <=( A235  and  A234 );
 a12159a <=( a12158a  and  a12155a );
 a12162a <=( (not A299)  and  A298 );
 a12166a <=( A302  and  (not A301) );
 a12167a <=( (not A300)  and  a12166a );
 a12168a <=( a12167a  and  a12162a );
 a12171a <=( (not A233)  and  A232 );
 a12174a <=( A235  and  A234 );
 a12175a <=( a12174a  and  a12171a );
 a12178a <=( A299  and  (not A298) );
 a12182a <=( A302  and  (not A301) );
 a12183a <=( (not A300)  and  a12182a );
 a12184a <=( a12183a  and  a12178a );
 a12187a <=( (not A233)  and  A232 );
 a12190a <=( (not A236)  and  A234 );
 a12191a <=( a12190a  and  a12187a );
 a12194a <=( (not A299)  and  A298 );
 a12198a <=( A302  and  (not A301) );
 a12199a <=( (not A300)  and  a12198a );
 a12200a <=( a12199a  and  a12194a );
 a12203a <=( (not A233)  and  A232 );
 a12206a <=( (not A236)  and  A234 );
 a12207a <=( a12206a  and  a12203a );
 a12210a <=( A299  and  (not A298) );
 a12214a <=( A302  and  (not A301) );
 a12215a <=( (not A300)  and  a12214a );
 a12216a <=( a12215a  and  a12210a );
 a12219a <=( (not A233)  and  A232 );
 a12222a <=( (not A235)  and  (not A234) );
 a12223a <=( a12222a  and  a12219a );
 a12226a <=( A298  and  A236 );
 a12230a <=( A301  and  A300 );
 a12231a <=( (not A299)  and  a12230a );
 a12232a <=( a12231a  and  a12226a );
 a12235a <=( (not A233)  and  A232 );
 a12238a <=( (not A235)  and  (not A234) );
 a12239a <=( a12238a  and  a12235a );
 a12242a <=( A298  and  A236 );
 a12246a <=( (not A302)  and  A300 );
 a12247a <=( (not A299)  and  a12246a );
 a12248a <=( a12247a  and  a12242a );
 a12251a <=( (not A233)  and  A232 );
 a12254a <=( (not A235)  and  (not A234) );
 a12255a <=( a12254a  and  a12251a );
 a12258a <=( (not A298)  and  A236 );
 a12262a <=( A301  and  A300 );
 a12263a <=( A299  and  a12262a );
 a12264a <=( a12263a  and  a12258a );
 a12267a <=( (not A233)  and  A232 );
 a12270a <=( (not A235)  and  (not A234) );
 a12271a <=( a12270a  and  a12267a );
 a12274a <=( (not A298)  and  A236 );
 a12278a <=( (not A302)  and  A300 );
 a12279a <=( A299  and  a12278a );
 a12280a <=( a12279a  and  a12274a );
 a12283a <=( (not A233)  and  A232 );
 a12286a <=( (not A235)  and  (not A234) );
 a12287a <=( a12286a  and  a12283a );
 a12290a <=( (not A265)  and  A236 );
 a12294a <=( A268  and  A267 );
 a12295a <=( A266  and  a12294a );
 a12296a <=( a12295a  and  a12290a );
 a12299a <=( (not A233)  and  A232 );
 a12302a <=( (not A235)  and  (not A234) );
 a12303a <=( a12302a  and  a12299a );
 a12306a <=( (not A265)  and  A236 );
 a12310a <=( (not A269)  and  A267 );
 a12311a <=( A266  and  a12310a );
 a12312a <=( a12311a  and  a12306a );
 a12315a <=( (not A233)  and  A232 );
 a12318a <=( (not A235)  and  (not A234) );
 a12319a <=( a12318a  and  a12315a );
 a12322a <=( A265  and  A236 );
 a12326a <=( A268  and  A267 );
 a12327a <=( (not A266)  and  a12326a );
 a12328a <=( a12327a  and  a12322a );
 a12331a <=( (not A233)  and  A232 );
 a12334a <=( (not A235)  and  (not A234) );
 a12335a <=( a12334a  and  a12331a );
 a12338a <=( A265  and  A236 );
 a12342a <=( (not A269)  and  A267 );
 a12343a <=( (not A266)  and  a12342a );
 a12344a <=( a12343a  and  a12338a );
 a12347a <=( A233  and  (not A232) );
 a12351a <=( (not A265)  and  A235 );
 a12352a <=( A234  and  a12351a );
 a12353a <=( a12352a  and  a12347a );
 a12356a <=( (not A267)  and  A266 );
 a12360a <=( A300  and  A269 );
 a12361a <=( (not A268)  and  a12360a );
 a12362a <=( a12361a  and  a12356a );
 a12365a <=( A233  and  (not A232) );
 a12369a <=( A265  and  A235 );
 a12370a <=( A234  and  a12369a );
 a12371a <=( a12370a  and  a12365a );
 a12374a <=( (not A267)  and  (not A266) );
 a12378a <=( A300  and  A269 );
 a12379a <=( (not A268)  and  a12378a );
 a12380a <=( a12379a  and  a12374a );
 a12383a <=( A233  and  (not A232) );
 a12387a <=( (not A265)  and  (not A236) );
 a12388a <=( A234  and  a12387a );
 a12389a <=( a12388a  and  a12383a );
 a12392a <=( (not A267)  and  A266 );
 a12396a <=( A300  and  A269 );
 a12397a <=( (not A268)  and  a12396a );
 a12398a <=( a12397a  and  a12392a );
 a12401a <=( A233  and  (not A232) );
 a12405a <=( A265  and  (not A236) );
 a12406a <=( A234  and  a12405a );
 a12407a <=( a12406a  and  a12401a );
 a12410a <=( (not A267)  and  (not A266) );
 a12414a <=( A300  and  A269 );
 a12415a <=( (not A268)  and  a12414a );
 a12416a <=( a12415a  and  a12410a );
 a12419a <=( A233  and  (not A232) );
 a12423a <=( A236  and  (not A235) );
 a12424a <=( (not A234)  and  a12423a );
 a12425a <=( a12424a  and  a12419a );
 a12428a <=( (not A299)  and  A298 );
 a12432a <=( A302  and  (not A301) );
 a12433a <=( (not A300)  and  a12432a );
 a12434a <=( a12433a  and  a12428a );
 a12437a <=( A233  and  (not A232) );
 a12441a <=( A236  and  (not A235) );
 a12442a <=( (not A234)  and  a12441a );
 a12443a <=( a12442a  and  a12437a );
 a12446a <=( A299  and  (not A298) );
 a12450a <=( A302  and  (not A301) );
 a12451a <=( (not A300)  and  a12450a );
 a12452a <=( a12451a  and  a12446a );
 a12455a <=( (not A233)  and  A232 );
 a12459a <=( (not A265)  and  A235 );
 a12460a <=( A234  and  a12459a );
 a12461a <=( a12460a  and  a12455a );
 a12464a <=( (not A267)  and  A266 );
 a12468a <=( A300  and  A269 );
 a12469a <=( (not A268)  and  a12468a );
 a12470a <=( a12469a  and  a12464a );
 a12473a <=( (not A233)  and  A232 );
 a12477a <=( A265  and  A235 );
 a12478a <=( A234  and  a12477a );
 a12479a <=( a12478a  and  a12473a );
 a12482a <=( (not A267)  and  (not A266) );
 a12486a <=( A300  and  A269 );
 a12487a <=( (not A268)  and  a12486a );
 a12488a <=( a12487a  and  a12482a );
 a12491a <=( (not A233)  and  A232 );
 a12495a <=( (not A265)  and  (not A236) );
 a12496a <=( A234  and  a12495a );
 a12497a <=( a12496a  and  a12491a );
 a12500a <=( (not A267)  and  A266 );
 a12504a <=( A300  and  A269 );
 a12505a <=( (not A268)  and  a12504a );
 a12506a <=( a12505a  and  a12500a );
 a12509a <=( (not A233)  and  A232 );
 a12513a <=( A265  and  (not A236) );
 a12514a <=( A234  and  a12513a );
 a12515a <=( a12514a  and  a12509a );
 a12518a <=( (not A267)  and  (not A266) );
 a12522a <=( A300  and  A269 );
 a12523a <=( (not A268)  and  a12522a );
 a12524a <=( a12523a  and  a12518a );
 a12527a <=( (not A233)  and  A232 );
 a12531a <=( A236  and  (not A235) );
 a12532a <=( (not A234)  and  a12531a );
 a12533a <=( a12532a  and  a12527a );
 a12536a <=( (not A299)  and  A298 );
 a12540a <=( A302  and  (not A301) );
 a12541a <=( (not A300)  and  a12540a );
 a12542a <=( a12541a  and  a12536a );
 a12545a <=( (not A233)  and  A232 );
 a12549a <=( A236  and  (not A235) );
 a12550a <=( (not A234)  and  a12549a );
 a12551a <=( a12550a  and  a12545a );
 a12554a <=( A299  and  (not A298) );
 a12558a <=( A302  and  (not A301) );
 a12559a <=( (not A300)  and  a12558a );
 a12560a <=( a12559a  and  a12554a );
 a12563a <=( (not A232)  and  (not A201) );
 a12567a <=( A235  and  A234 );
 a12568a <=( A233  and  a12567a );
 a12569a <=( a12568a  and  a12563a );
 a12572a <=( A266  and  (not A265) );
 a12576a <=( A269  and  (not A268) );
 a12577a <=( (not A267)  and  a12576a );
 a12578a <=( a12577a  and  a12572a );
 a12581a <=( (not A232)  and  (not A201) );
 a12585a <=( A235  and  A234 );
 a12586a <=( A233  and  a12585a );
 a12587a <=( a12586a  and  a12581a );
 a12590a <=( (not A266)  and  A265 );
 a12594a <=( A269  and  (not A268) );
 a12595a <=( (not A267)  and  a12594a );
 a12596a <=( a12595a  and  a12590a );
 a12599a <=( (not A232)  and  (not A201) );
 a12603a <=( (not A236)  and  A234 );
 a12604a <=( A233  and  a12603a );
 a12605a <=( a12604a  and  a12599a );
 a12608a <=( A266  and  (not A265) );
 a12612a <=( A269  and  (not A268) );
 a12613a <=( (not A267)  and  a12612a );
 a12614a <=( a12613a  and  a12608a );
 a12617a <=( (not A232)  and  (not A201) );
 a12621a <=( (not A236)  and  A234 );
 a12622a <=( A233  and  a12621a );
 a12623a <=( a12622a  and  a12617a );
 a12626a <=( (not A266)  and  A265 );
 a12630a <=( A269  and  (not A268) );
 a12631a <=( (not A267)  and  a12630a );
 a12632a <=( a12631a  and  a12626a );
 a12635a <=( A232  and  (not A201) );
 a12639a <=( A235  and  A234 );
 a12640a <=( (not A233)  and  a12639a );
 a12641a <=( a12640a  and  a12635a );
 a12644a <=( A266  and  (not A265) );
 a12648a <=( A269  and  (not A268) );
 a12649a <=( (not A267)  and  a12648a );
 a12650a <=( a12649a  and  a12644a );
 a12653a <=( A232  and  (not A201) );
 a12657a <=( A235  and  A234 );
 a12658a <=( (not A233)  and  a12657a );
 a12659a <=( a12658a  and  a12653a );
 a12662a <=( (not A266)  and  A265 );
 a12666a <=( A269  and  (not A268) );
 a12667a <=( (not A267)  and  a12666a );
 a12668a <=( a12667a  and  a12662a );
 a12671a <=( A232  and  (not A201) );
 a12675a <=( (not A236)  and  A234 );
 a12676a <=( (not A233)  and  a12675a );
 a12677a <=( a12676a  and  a12671a );
 a12680a <=( A266  and  (not A265) );
 a12684a <=( A269  and  (not A268) );
 a12685a <=( (not A267)  and  a12684a );
 a12686a <=( a12685a  and  a12680a );
 a12689a <=( A232  and  (not A201) );
 a12693a <=( (not A236)  and  A234 );
 a12694a <=( (not A233)  and  a12693a );
 a12695a <=( a12694a  and  a12689a );
 a12698a <=( (not A266)  and  A265 );
 a12702a <=( A269  and  (not A268) );
 a12703a <=( (not A267)  and  a12702a );
 a12704a <=( a12703a  and  a12698a );
 a12707a <=( A166  and  A167 );
 a12711a <=( A201  and  A200 );
 a12712a <=( (not A199)  and  a12711a );
 a12713a <=( a12712a  and  a12707a );
 a12716a <=( (not A267)  and  A202 );
 a12720a <=( A301  and  (not A300) );
 a12721a <=( A268  and  a12720a );
 a12722a <=( a12721a  and  a12716a );
 a12725a <=( A166  and  A167 );
 a12729a <=( A201  and  A200 );
 a12730a <=( (not A199)  and  a12729a );
 a12731a <=( a12730a  and  a12725a );
 a12734a <=( (not A267)  and  A202 );
 a12738a <=( (not A302)  and  (not A300) );
 a12739a <=( A268  and  a12738a );
 a12740a <=( a12739a  and  a12734a );
 a12743a <=( A166  and  A167 );
 a12747a <=( A201  and  A200 );
 a12748a <=( (not A199)  and  a12747a );
 a12749a <=( a12748a  and  a12743a );
 a12752a <=( (not A267)  and  A202 );
 a12756a <=( A299  and  A298 );
 a12757a <=( A268  and  a12756a );
 a12758a <=( a12757a  and  a12752a );
 a12761a <=( A166  and  A167 );
 a12765a <=( A201  and  A200 );
 a12766a <=( (not A199)  and  a12765a );
 a12767a <=( a12766a  and  a12761a );
 a12770a <=( (not A267)  and  A202 );
 a12774a <=( (not A299)  and  (not A298) );
 a12775a <=( A268  and  a12774a );
 a12776a <=( a12775a  and  a12770a );
 a12779a <=( A166  and  A167 );
 a12783a <=( A201  and  A200 );
 a12784a <=( (not A199)  and  a12783a );
 a12785a <=( a12784a  and  a12779a );
 a12788a <=( (not A267)  and  A202 );
 a12792a <=( A301  and  (not A300) );
 a12793a <=( (not A269)  and  a12792a );
 a12794a <=( a12793a  and  a12788a );
 a12797a <=( A166  and  A167 );
 a12801a <=( A201  and  A200 );
 a12802a <=( (not A199)  and  a12801a );
 a12803a <=( a12802a  and  a12797a );
 a12806a <=( (not A267)  and  A202 );
 a12810a <=( (not A302)  and  (not A300) );
 a12811a <=( (not A269)  and  a12810a );
 a12812a <=( a12811a  and  a12806a );
 a12815a <=( A166  and  A167 );
 a12819a <=( A201  and  A200 );
 a12820a <=( (not A199)  and  a12819a );
 a12821a <=( a12820a  and  a12815a );
 a12824a <=( (not A267)  and  A202 );
 a12828a <=( A299  and  A298 );
 a12829a <=( (not A269)  and  a12828a );
 a12830a <=( a12829a  and  a12824a );
 a12833a <=( A166  and  A167 );
 a12837a <=( A201  and  A200 );
 a12838a <=( (not A199)  and  a12837a );
 a12839a <=( a12838a  and  a12833a );
 a12842a <=( (not A267)  and  A202 );
 a12846a <=( (not A299)  and  (not A298) );
 a12847a <=( (not A269)  and  a12846a );
 a12848a <=( a12847a  and  a12842a );
 a12851a <=( A166  and  A167 );
 a12855a <=( A201  and  A200 );
 a12856a <=( (not A199)  and  a12855a );
 a12857a <=( a12856a  and  a12851a );
 a12860a <=( A265  and  A202 );
 a12864a <=( A301  and  (not A300) );
 a12865a <=( A266  and  a12864a );
 a12866a <=( a12865a  and  a12860a );
 a12869a <=( A166  and  A167 );
 a12873a <=( A201  and  A200 );
 a12874a <=( (not A199)  and  a12873a );
 a12875a <=( a12874a  and  a12869a );
 a12878a <=( A265  and  A202 );
 a12882a <=( (not A302)  and  (not A300) );
 a12883a <=( A266  and  a12882a );
 a12884a <=( a12883a  and  a12878a );
 a12887a <=( A166  and  A167 );
 a12891a <=( A201  and  A200 );
 a12892a <=( (not A199)  and  a12891a );
 a12893a <=( a12892a  and  a12887a );
 a12896a <=( A265  and  A202 );
 a12900a <=( A299  and  A298 );
 a12901a <=( A266  and  a12900a );
 a12902a <=( a12901a  and  a12896a );
 a12905a <=( A166  and  A167 );
 a12909a <=( A201  and  A200 );
 a12910a <=( (not A199)  and  a12909a );
 a12911a <=( a12910a  and  a12905a );
 a12914a <=( A265  and  A202 );
 a12918a <=( (not A299)  and  (not A298) );
 a12919a <=( A266  and  a12918a );
 a12920a <=( a12919a  and  a12914a );
 a12923a <=( A166  and  A167 );
 a12927a <=( A201  and  A200 );
 a12928a <=( (not A199)  and  a12927a );
 a12929a <=( a12928a  and  a12923a );
 a12932a <=( (not A265)  and  A202 );
 a12936a <=( A301  and  (not A300) );
 a12937a <=( (not A266)  and  a12936a );
 a12938a <=( a12937a  and  a12932a );
 a12941a <=( A166  and  A167 );
 a12945a <=( A201  and  A200 );
 a12946a <=( (not A199)  and  a12945a );
 a12947a <=( a12946a  and  a12941a );
 a12950a <=( (not A265)  and  A202 );
 a12954a <=( (not A302)  and  (not A300) );
 a12955a <=( (not A266)  and  a12954a );
 a12956a <=( a12955a  and  a12950a );
 a12959a <=( A166  and  A167 );
 a12963a <=( A201  and  A200 );
 a12964a <=( (not A199)  and  a12963a );
 a12965a <=( a12964a  and  a12959a );
 a12968a <=( (not A265)  and  A202 );
 a12972a <=( A299  and  A298 );
 a12973a <=( (not A266)  and  a12972a );
 a12974a <=( a12973a  and  a12968a );
 a12977a <=( A166  and  A167 );
 a12981a <=( A201  and  A200 );
 a12982a <=( (not A199)  and  a12981a );
 a12983a <=( a12982a  and  a12977a );
 a12986a <=( (not A265)  and  A202 );
 a12990a <=( (not A299)  and  (not A298) );
 a12991a <=( (not A266)  and  a12990a );
 a12992a <=( a12991a  and  a12986a );
 a12995a <=( A166  and  A167 );
 a12999a <=( A201  and  A200 );
 a13000a <=( (not A199)  and  a12999a );
 a13001a <=( a13000a  and  a12995a );
 a13004a <=( (not A267)  and  (not A203) );
 a13008a <=( A301  and  (not A300) );
 a13009a <=( A268  and  a13008a );
 a13010a <=( a13009a  and  a13004a );
 a13013a <=( A166  and  A167 );
 a13017a <=( A201  and  A200 );
 a13018a <=( (not A199)  and  a13017a );
 a13019a <=( a13018a  and  a13013a );
 a13022a <=( (not A267)  and  (not A203) );
 a13026a <=( (not A302)  and  (not A300) );
 a13027a <=( A268  and  a13026a );
 a13028a <=( a13027a  and  a13022a );
 a13031a <=( A166  and  A167 );
 a13035a <=( A201  and  A200 );
 a13036a <=( (not A199)  and  a13035a );
 a13037a <=( a13036a  and  a13031a );
 a13040a <=( (not A267)  and  (not A203) );
 a13044a <=( A299  and  A298 );
 a13045a <=( A268  and  a13044a );
 a13046a <=( a13045a  and  a13040a );
 a13049a <=( A166  and  A167 );
 a13053a <=( A201  and  A200 );
 a13054a <=( (not A199)  and  a13053a );
 a13055a <=( a13054a  and  a13049a );
 a13058a <=( (not A267)  and  (not A203) );
 a13062a <=( (not A299)  and  (not A298) );
 a13063a <=( A268  and  a13062a );
 a13064a <=( a13063a  and  a13058a );
 a13067a <=( A166  and  A167 );
 a13071a <=( A201  and  A200 );
 a13072a <=( (not A199)  and  a13071a );
 a13073a <=( a13072a  and  a13067a );
 a13076a <=( (not A267)  and  (not A203) );
 a13080a <=( A301  and  (not A300) );
 a13081a <=( (not A269)  and  a13080a );
 a13082a <=( a13081a  and  a13076a );
 a13085a <=( A166  and  A167 );
 a13089a <=( A201  and  A200 );
 a13090a <=( (not A199)  and  a13089a );
 a13091a <=( a13090a  and  a13085a );
 a13094a <=( (not A267)  and  (not A203) );
 a13098a <=( (not A302)  and  (not A300) );
 a13099a <=( (not A269)  and  a13098a );
 a13100a <=( a13099a  and  a13094a );
 a13103a <=( A166  and  A167 );
 a13107a <=( A201  and  A200 );
 a13108a <=( (not A199)  and  a13107a );
 a13109a <=( a13108a  and  a13103a );
 a13112a <=( (not A267)  and  (not A203) );
 a13116a <=( A299  and  A298 );
 a13117a <=( (not A269)  and  a13116a );
 a13118a <=( a13117a  and  a13112a );
 a13121a <=( A166  and  A167 );
 a13125a <=( A201  and  A200 );
 a13126a <=( (not A199)  and  a13125a );
 a13127a <=( a13126a  and  a13121a );
 a13130a <=( (not A267)  and  (not A203) );
 a13134a <=( (not A299)  and  (not A298) );
 a13135a <=( (not A269)  and  a13134a );
 a13136a <=( a13135a  and  a13130a );
 a13139a <=( A166  and  A167 );
 a13143a <=( A201  and  A200 );
 a13144a <=( (not A199)  and  a13143a );
 a13145a <=( a13144a  and  a13139a );
 a13148a <=( A265  and  (not A203) );
 a13152a <=( A301  and  (not A300) );
 a13153a <=( A266  and  a13152a );
 a13154a <=( a13153a  and  a13148a );
 a13157a <=( A166  and  A167 );
 a13161a <=( A201  and  A200 );
 a13162a <=( (not A199)  and  a13161a );
 a13163a <=( a13162a  and  a13157a );
 a13166a <=( A265  and  (not A203) );
 a13170a <=( (not A302)  and  (not A300) );
 a13171a <=( A266  and  a13170a );
 a13172a <=( a13171a  and  a13166a );
 a13175a <=( A166  and  A167 );
 a13179a <=( A201  and  A200 );
 a13180a <=( (not A199)  and  a13179a );
 a13181a <=( a13180a  and  a13175a );
 a13184a <=( A265  and  (not A203) );
 a13188a <=( A299  and  A298 );
 a13189a <=( A266  and  a13188a );
 a13190a <=( a13189a  and  a13184a );
 a13193a <=( A166  and  A167 );
 a13197a <=( A201  and  A200 );
 a13198a <=( (not A199)  and  a13197a );
 a13199a <=( a13198a  and  a13193a );
 a13202a <=( A265  and  (not A203) );
 a13206a <=( (not A299)  and  (not A298) );
 a13207a <=( A266  and  a13206a );
 a13208a <=( a13207a  and  a13202a );
 a13211a <=( A166  and  A167 );
 a13215a <=( A201  and  A200 );
 a13216a <=( (not A199)  and  a13215a );
 a13217a <=( a13216a  and  a13211a );
 a13220a <=( (not A265)  and  (not A203) );
 a13224a <=( A301  and  (not A300) );
 a13225a <=( (not A266)  and  a13224a );
 a13226a <=( a13225a  and  a13220a );
 a13229a <=( A166  and  A167 );
 a13233a <=( A201  and  A200 );
 a13234a <=( (not A199)  and  a13233a );
 a13235a <=( a13234a  and  a13229a );
 a13238a <=( (not A265)  and  (not A203) );
 a13242a <=( (not A302)  and  (not A300) );
 a13243a <=( (not A266)  and  a13242a );
 a13244a <=( a13243a  and  a13238a );
 a13247a <=( A166  and  A167 );
 a13251a <=( A201  and  A200 );
 a13252a <=( (not A199)  and  a13251a );
 a13253a <=( a13252a  and  a13247a );
 a13256a <=( (not A265)  and  (not A203) );
 a13260a <=( A299  and  A298 );
 a13261a <=( (not A266)  and  a13260a );
 a13262a <=( a13261a  and  a13256a );
 a13265a <=( A166  and  A167 );
 a13269a <=( A201  and  A200 );
 a13270a <=( (not A199)  and  a13269a );
 a13271a <=( a13270a  and  a13265a );
 a13274a <=( (not A265)  and  (not A203) );
 a13278a <=( (not A299)  and  (not A298) );
 a13279a <=( (not A266)  and  a13278a );
 a13280a <=( a13279a  and  a13274a );
 a13283a <=( A166  and  A167 );
 a13287a <=( A201  and  (not A200) );
 a13288a <=( A199  and  a13287a );
 a13289a <=( a13288a  and  a13283a );
 a13292a <=( (not A267)  and  A202 );
 a13296a <=( A301  and  (not A300) );
 a13297a <=( A268  and  a13296a );
 a13298a <=( a13297a  and  a13292a );
 a13301a <=( A166  and  A167 );
 a13305a <=( A201  and  (not A200) );
 a13306a <=( A199  and  a13305a );
 a13307a <=( a13306a  and  a13301a );
 a13310a <=( (not A267)  and  A202 );
 a13314a <=( (not A302)  and  (not A300) );
 a13315a <=( A268  and  a13314a );
 a13316a <=( a13315a  and  a13310a );
 a13319a <=( A166  and  A167 );
 a13323a <=( A201  and  (not A200) );
 a13324a <=( A199  and  a13323a );
 a13325a <=( a13324a  and  a13319a );
 a13328a <=( (not A267)  and  A202 );
 a13332a <=( A299  and  A298 );
 a13333a <=( A268  and  a13332a );
 a13334a <=( a13333a  and  a13328a );
 a13337a <=( A166  and  A167 );
 a13341a <=( A201  and  (not A200) );
 a13342a <=( A199  and  a13341a );
 a13343a <=( a13342a  and  a13337a );
 a13346a <=( (not A267)  and  A202 );
 a13350a <=( (not A299)  and  (not A298) );
 a13351a <=( A268  and  a13350a );
 a13352a <=( a13351a  and  a13346a );
 a13355a <=( A166  and  A167 );
 a13359a <=( A201  and  (not A200) );
 a13360a <=( A199  and  a13359a );
 a13361a <=( a13360a  and  a13355a );
 a13364a <=( (not A267)  and  A202 );
 a13368a <=( A301  and  (not A300) );
 a13369a <=( (not A269)  and  a13368a );
 a13370a <=( a13369a  and  a13364a );
 a13373a <=( A166  and  A167 );
 a13377a <=( A201  and  (not A200) );
 a13378a <=( A199  and  a13377a );
 a13379a <=( a13378a  and  a13373a );
 a13382a <=( (not A267)  and  A202 );
 a13386a <=( (not A302)  and  (not A300) );
 a13387a <=( (not A269)  and  a13386a );
 a13388a <=( a13387a  and  a13382a );
 a13391a <=( A166  and  A167 );
 a13395a <=( A201  and  (not A200) );
 a13396a <=( A199  and  a13395a );
 a13397a <=( a13396a  and  a13391a );
 a13400a <=( (not A267)  and  A202 );
 a13404a <=( A299  and  A298 );
 a13405a <=( (not A269)  and  a13404a );
 a13406a <=( a13405a  and  a13400a );
 a13409a <=( A166  and  A167 );
 a13413a <=( A201  and  (not A200) );
 a13414a <=( A199  and  a13413a );
 a13415a <=( a13414a  and  a13409a );
 a13418a <=( (not A267)  and  A202 );
 a13422a <=( (not A299)  and  (not A298) );
 a13423a <=( (not A269)  and  a13422a );
 a13424a <=( a13423a  and  a13418a );
 a13427a <=( A166  and  A167 );
 a13431a <=( A201  and  (not A200) );
 a13432a <=( A199  and  a13431a );
 a13433a <=( a13432a  and  a13427a );
 a13436a <=( A265  and  A202 );
 a13440a <=( A301  and  (not A300) );
 a13441a <=( A266  and  a13440a );
 a13442a <=( a13441a  and  a13436a );
 a13445a <=( A166  and  A167 );
 a13449a <=( A201  and  (not A200) );
 a13450a <=( A199  and  a13449a );
 a13451a <=( a13450a  and  a13445a );
 a13454a <=( A265  and  A202 );
 a13458a <=( (not A302)  and  (not A300) );
 a13459a <=( A266  and  a13458a );
 a13460a <=( a13459a  and  a13454a );
 a13463a <=( A166  and  A167 );
 a13467a <=( A201  and  (not A200) );
 a13468a <=( A199  and  a13467a );
 a13469a <=( a13468a  and  a13463a );
 a13472a <=( A265  and  A202 );
 a13476a <=( A299  and  A298 );
 a13477a <=( A266  and  a13476a );
 a13478a <=( a13477a  and  a13472a );
 a13481a <=( A166  and  A167 );
 a13485a <=( A201  and  (not A200) );
 a13486a <=( A199  and  a13485a );
 a13487a <=( a13486a  and  a13481a );
 a13490a <=( A265  and  A202 );
 a13494a <=( (not A299)  and  (not A298) );
 a13495a <=( A266  and  a13494a );
 a13496a <=( a13495a  and  a13490a );
 a13499a <=( A166  and  A167 );
 a13503a <=( A201  and  (not A200) );
 a13504a <=( A199  and  a13503a );
 a13505a <=( a13504a  and  a13499a );
 a13508a <=( (not A265)  and  A202 );
 a13512a <=( A301  and  (not A300) );
 a13513a <=( (not A266)  and  a13512a );
 a13514a <=( a13513a  and  a13508a );
 a13517a <=( A166  and  A167 );
 a13521a <=( A201  and  (not A200) );
 a13522a <=( A199  and  a13521a );
 a13523a <=( a13522a  and  a13517a );
 a13526a <=( (not A265)  and  A202 );
 a13530a <=( (not A302)  and  (not A300) );
 a13531a <=( (not A266)  and  a13530a );
 a13532a <=( a13531a  and  a13526a );
 a13535a <=( A166  and  A167 );
 a13539a <=( A201  and  (not A200) );
 a13540a <=( A199  and  a13539a );
 a13541a <=( a13540a  and  a13535a );
 a13544a <=( (not A265)  and  A202 );
 a13548a <=( A299  and  A298 );
 a13549a <=( (not A266)  and  a13548a );
 a13550a <=( a13549a  and  a13544a );
 a13553a <=( A166  and  A167 );
 a13557a <=( A201  and  (not A200) );
 a13558a <=( A199  and  a13557a );
 a13559a <=( a13558a  and  a13553a );
 a13562a <=( (not A265)  and  A202 );
 a13566a <=( (not A299)  and  (not A298) );
 a13567a <=( (not A266)  and  a13566a );
 a13568a <=( a13567a  and  a13562a );
 a13571a <=( A166  and  A167 );
 a13575a <=( A201  and  (not A200) );
 a13576a <=( A199  and  a13575a );
 a13577a <=( a13576a  and  a13571a );
 a13580a <=( (not A267)  and  (not A203) );
 a13584a <=( A301  and  (not A300) );
 a13585a <=( A268  and  a13584a );
 a13586a <=( a13585a  and  a13580a );
 a13589a <=( A166  and  A167 );
 a13593a <=( A201  and  (not A200) );
 a13594a <=( A199  and  a13593a );
 a13595a <=( a13594a  and  a13589a );
 a13598a <=( (not A267)  and  (not A203) );
 a13602a <=( (not A302)  and  (not A300) );
 a13603a <=( A268  and  a13602a );
 a13604a <=( a13603a  and  a13598a );
 a13607a <=( A166  and  A167 );
 a13611a <=( A201  and  (not A200) );
 a13612a <=( A199  and  a13611a );
 a13613a <=( a13612a  and  a13607a );
 a13616a <=( (not A267)  and  (not A203) );
 a13620a <=( A299  and  A298 );
 a13621a <=( A268  and  a13620a );
 a13622a <=( a13621a  and  a13616a );
 a13625a <=( A166  and  A167 );
 a13629a <=( A201  and  (not A200) );
 a13630a <=( A199  and  a13629a );
 a13631a <=( a13630a  and  a13625a );
 a13634a <=( (not A267)  and  (not A203) );
 a13638a <=( (not A299)  and  (not A298) );
 a13639a <=( A268  and  a13638a );
 a13640a <=( a13639a  and  a13634a );
 a13643a <=( A166  and  A167 );
 a13647a <=( A201  and  (not A200) );
 a13648a <=( A199  and  a13647a );
 a13649a <=( a13648a  and  a13643a );
 a13652a <=( (not A267)  and  (not A203) );
 a13656a <=( A301  and  (not A300) );
 a13657a <=( (not A269)  and  a13656a );
 a13658a <=( a13657a  and  a13652a );
 a13661a <=( A166  and  A167 );
 a13665a <=( A201  and  (not A200) );
 a13666a <=( A199  and  a13665a );
 a13667a <=( a13666a  and  a13661a );
 a13670a <=( (not A267)  and  (not A203) );
 a13674a <=( (not A302)  and  (not A300) );
 a13675a <=( (not A269)  and  a13674a );
 a13676a <=( a13675a  and  a13670a );
 a13679a <=( A166  and  A167 );
 a13683a <=( A201  and  (not A200) );
 a13684a <=( A199  and  a13683a );
 a13685a <=( a13684a  and  a13679a );
 a13688a <=( (not A267)  and  (not A203) );
 a13692a <=( A299  and  A298 );
 a13693a <=( (not A269)  and  a13692a );
 a13694a <=( a13693a  and  a13688a );
 a13697a <=( A166  and  A167 );
 a13701a <=( A201  and  (not A200) );
 a13702a <=( A199  and  a13701a );
 a13703a <=( a13702a  and  a13697a );
 a13706a <=( (not A267)  and  (not A203) );
 a13710a <=( (not A299)  and  (not A298) );
 a13711a <=( (not A269)  and  a13710a );
 a13712a <=( a13711a  and  a13706a );
 a13715a <=( A166  and  A167 );
 a13719a <=( A201  and  (not A200) );
 a13720a <=( A199  and  a13719a );
 a13721a <=( a13720a  and  a13715a );
 a13724a <=( A265  and  (not A203) );
 a13728a <=( A301  and  (not A300) );
 a13729a <=( A266  and  a13728a );
 a13730a <=( a13729a  and  a13724a );
 a13733a <=( A166  and  A167 );
 a13737a <=( A201  and  (not A200) );
 a13738a <=( A199  and  a13737a );
 a13739a <=( a13738a  and  a13733a );
 a13742a <=( A265  and  (not A203) );
 a13746a <=( (not A302)  and  (not A300) );
 a13747a <=( A266  and  a13746a );
 a13748a <=( a13747a  and  a13742a );
 a13751a <=( A166  and  A167 );
 a13755a <=( A201  and  (not A200) );
 a13756a <=( A199  and  a13755a );
 a13757a <=( a13756a  and  a13751a );
 a13760a <=( A265  and  (not A203) );
 a13764a <=( A299  and  A298 );
 a13765a <=( A266  and  a13764a );
 a13766a <=( a13765a  and  a13760a );
 a13769a <=( A166  and  A167 );
 a13773a <=( A201  and  (not A200) );
 a13774a <=( A199  and  a13773a );
 a13775a <=( a13774a  and  a13769a );
 a13778a <=( A265  and  (not A203) );
 a13782a <=( (not A299)  and  (not A298) );
 a13783a <=( A266  and  a13782a );
 a13784a <=( a13783a  and  a13778a );
 a13787a <=( A166  and  A167 );
 a13791a <=( A201  and  (not A200) );
 a13792a <=( A199  and  a13791a );
 a13793a <=( a13792a  and  a13787a );
 a13796a <=( (not A265)  and  (not A203) );
 a13800a <=( A301  and  (not A300) );
 a13801a <=( (not A266)  and  a13800a );
 a13802a <=( a13801a  and  a13796a );
 a13805a <=( A166  and  A167 );
 a13809a <=( A201  and  (not A200) );
 a13810a <=( A199  and  a13809a );
 a13811a <=( a13810a  and  a13805a );
 a13814a <=( (not A265)  and  (not A203) );
 a13818a <=( (not A302)  and  (not A300) );
 a13819a <=( (not A266)  and  a13818a );
 a13820a <=( a13819a  and  a13814a );
 a13823a <=( A166  and  A167 );
 a13827a <=( A201  and  (not A200) );
 a13828a <=( A199  and  a13827a );
 a13829a <=( a13828a  and  a13823a );
 a13832a <=( (not A265)  and  (not A203) );
 a13836a <=( A299  and  A298 );
 a13837a <=( (not A266)  and  a13836a );
 a13838a <=( a13837a  and  a13832a );
 a13841a <=( A166  and  A167 );
 a13845a <=( A201  and  (not A200) );
 a13846a <=( A199  and  a13845a );
 a13847a <=( a13846a  and  a13841a );
 a13850a <=( (not A265)  and  (not A203) );
 a13854a <=( (not A299)  and  (not A298) );
 a13855a <=( (not A266)  and  a13854a );
 a13856a <=( a13855a  and  a13850a );
 a13859a <=( (not A166)  and  (not A167) );
 a13863a <=( A201  and  A200 );
 a13864a <=( (not A199)  and  a13863a );
 a13865a <=( a13864a  and  a13859a );
 a13868a <=( (not A267)  and  A202 );
 a13872a <=( A301  and  (not A300) );
 a13873a <=( A268  and  a13872a );
 a13874a <=( a13873a  and  a13868a );
 a13877a <=( (not A166)  and  (not A167) );
 a13881a <=( A201  and  A200 );
 a13882a <=( (not A199)  and  a13881a );
 a13883a <=( a13882a  and  a13877a );
 a13886a <=( (not A267)  and  A202 );
 a13890a <=( (not A302)  and  (not A300) );
 a13891a <=( A268  and  a13890a );
 a13892a <=( a13891a  and  a13886a );
 a13895a <=( (not A166)  and  (not A167) );
 a13899a <=( A201  and  A200 );
 a13900a <=( (not A199)  and  a13899a );
 a13901a <=( a13900a  and  a13895a );
 a13904a <=( (not A267)  and  A202 );
 a13908a <=( A299  and  A298 );
 a13909a <=( A268  and  a13908a );
 a13910a <=( a13909a  and  a13904a );
 a13913a <=( (not A166)  and  (not A167) );
 a13917a <=( A201  and  A200 );
 a13918a <=( (not A199)  and  a13917a );
 a13919a <=( a13918a  and  a13913a );
 a13922a <=( (not A267)  and  A202 );
 a13926a <=( (not A299)  and  (not A298) );
 a13927a <=( A268  and  a13926a );
 a13928a <=( a13927a  and  a13922a );
 a13931a <=( (not A166)  and  (not A167) );
 a13935a <=( A201  and  A200 );
 a13936a <=( (not A199)  and  a13935a );
 a13937a <=( a13936a  and  a13931a );
 a13940a <=( (not A267)  and  A202 );
 a13944a <=( A301  and  (not A300) );
 a13945a <=( (not A269)  and  a13944a );
 a13946a <=( a13945a  and  a13940a );
 a13949a <=( (not A166)  and  (not A167) );
 a13953a <=( A201  and  A200 );
 a13954a <=( (not A199)  and  a13953a );
 a13955a <=( a13954a  and  a13949a );
 a13958a <=( (not A267)  and  A202 );
 a13962a <=( (not A302)  and  (not A300) );
 a13963a <=( (not A269)  and  a13962a );
 a13964a <=( a13963a  and  a13958a );
 a13967a <=( (not A166)  and  (not A167) );
 a13971a <=( A201  and  A200 );
 a13972a <=( (not A199)  and  a13971a );
 a13973a <=( a13972a  and  a13967a );
 a13976a <=( (not A267)  and  A202 );
 a13980a <=( A299  and  A298 );
 a13981a <=( (not A269)  and  a13980a );
 a13982a <=( a13981a  and  a13976a );
 a13985a <=( (not A166)  and  (not A167) );
 a13989a <=( A201  and  A200 );
 a13990a <=( (not A199)  and  a13989a );
 a13991a <=( a13990a  and  a13985a );
 a13994a <=( (not A267)  and  A202 );
 a13998a <=( (not A299)  and  (not A298) );
 a13999a <=( (not A269)  and  a13998a );
 a14000a <=( a13999a  and  a13994a );
 a14003a <=( (not A166)  and  (not A167) );
 a14007a <=( A201  and  A200 );
 a14008a <=( (not A199)  and  a14007a );
 a14009a <=( a14008a  and  a14003a );
 a14012a <=( A265  and  A202 );
 a14016a <=( A301  and  (not A300) );
 a14017a <=( A266  and  a14016a );
 a14018a <=( a14017a  and  a14012a );
 a14021a <=( (not A166)  and  (not A167) );
 a14025a <=( A201  and  A200 );
 a14026a <=( (not A199)  and  a14025a );
 a14027a <=( a14026a  and  a14021a );
 a14030a <=( A265  and  A202 );
 a14034a <=( (not A302)  and  (not A300) );
 a14035a <=( A266  and  a14034a );
 a14036a <=( a14035a  and  a14030a );
 a14039a <=( (not A166)  and  (not A167) );
 a14043a <=( A201  and  A200 );
 a14044a <=( (not A199)  and  a14043a );
 a14045a <=( a14044a  and  a14039a );
 a14048a <=( A265  and  A202 );
 a14052a <=( A299  and  A298 );
 a14053a <=( A266  and  a14052a );
 a14054a <=( a14053a  and  a14048a );
 a14057a <=( (not A166)  and  (not A167) );
 a14061a <=( A201  and  A200 );
 a14062a <=( (not A199)  and  a14061a );
 a14063a <=( a14062a  and  a14057a );
 a14066a <=( A265  and  A202 );
 a14070a <=( (not A299)  and  (not A298) );
 a14071a <=( A266  and  a14070a );
 a14072a <=( a14071a  and  a14066a );
 a14075a <=( (not A166)  and  (not A167) );
 a14079a <=( A201  and  A200 );
 a14080a <=( (not A199)  and  a14079a );
 a14081a <=( a14080a  and  a14075a );
 a14084a <=( (not A265)  and  A202 );
 a14088a <=( A301  and  (not A300) );
 a14089a <=( (not A266)  and  a14088a );
 a14090a <=( a14089a  and  a14084a );
 a14093a <=( (not A166)  and  (not A167) );
 a14097a <=( A201  and  A200 );
 a14098a <=( (not A199)  and  a14097a );
 a14099a <=( a14098a  and  a14093a );
 a14102a <=( (not A265)  and  A202 );
 a14106a <=( (not A302)  and  (not A300) );
 a14107a <=( (not A266)  and  a14106a );
 a14108a <=( a14107a  and  a14102a );
 a14111a <=( (not A166)  and  (not A167) );
 a14115a <=( A201  and  A200 );
 a14116a <=( (not A199)  and  a14115a );
 a14117a <=( a14116a  and  a14111a );
 a14120a <=( (not A265)  and  A202 );
 a14124a <=( A299  and  A298 );
 a14125a <=( (not A266)  and  a14124a );
 a14126a <=( a14125a  and  a14120a );
 a14129a <=( (not A166)  and  (not A167) );
 a14133a <=( A201  and  A200 );
 a14134a <=( (not A199)  and  a14133a );
 a14135a <=( a14134a  and  a14129a );
 a14138a <=( (not A265)  and  A202 );
 a14142a <=( (not A299)  and  (not A298) );
 a14143a <=( (not A266)  and  a14142a );
 a14144a <=( a14143a  and  a14138a );
 a14147a <=( (not A166)  and  (not A167) );
 a14151a <=( A201  and  A200 );
 a14152a <=( (not A199)  and  a14151a );
 a14153a <=( a14152a  and  a14147a );
 a14156a <=( (not A267)  and  (not A203) );
 a14160a <=( A301  and  (not A300) );
 a14161a <=( A268  and  a14160a );
 a14162a <=( a14161a  and  a14156a );
 a14165a <=( (not A166)  and  (not A167) );
 a14169a <=( A201  and  A200 );
 a14170a <=( (not A199)  and  a14169a );
 a14171a <=( a14170a  and  a14165a );
 a14174a <=( (not A267)  and  (not A203) );
 a14178a <=( (not A302)  and  (not A300) );
 a14179a <=( A268  and  a14178a );
 a14180a <=( a14179a  and  a14174a );
 a14183a <=( (not A166)  and  (not A167) );
 a14187a <=( A201  and  A200 );
 a14188a <=( (not A199)  and  a14187a );
 a14189a <=( a14188a  and  a14183a );
 a14192a <=( (not A267)  and  (not A203) );
 a14196a <=( A299  and  A298 );
 a14197a <=( A268  and  a14196a );
 a14198a <=( a14197a  and  a14192a );
 a14201a <=( (not A166)  and  (not A167) );
 a14205a <=( A201  and  A200 );
 a14206a <=( (not A199)  and  a14205a );
 a14207a <=( a14206a  and  a14201a );
 a14210a <=( (not A267)  and  (not A203) );
 a14214a <=( (not A299)  and  (not A298) );
 a14215a <=( A268  and  a14214a );
 a14216a <=( a14215a  and  a14210a );
 a14219a <=( (not A166)  and  (not A167) );
 a14223a <=( A201  and  A200 );
 a14224a <=( (not A199)  and  a14223a );
 a14225a <=( a14224a  and  a14219a );
 a14228a <=( (not A267)  and  (not A203) );
 a14232a <=( A301  and  (not A300) );
 a14233a <=( (not A269)  and  a14232a );
 a14234a <=( a14233a  and  a14228a );
 a14237a <=( (not A166)  and  (not A167) );
 a14241a <=( A201  and  A200 );
 a14242a <=( (not A199)  and  a14241a );
 a14243a <=( a14242a  and  a14237a );
 a14246a <=( (not A267)  and  (not A203) );
 a14250a <=( (not A302)  and  (not A300) );
 a14251a <=( (not A269)  and  a14250a );
 a14252a <=( a14251a  and  a14246a );
 a14255a <=( (not A166)  and  (not A167) );
 a14259a <=( A201  and  A200 );
 a14260a <=( (not A199)  and  a14259a );
 a14261a <=( a14260a  and  a14255a );
 a14264a <=( (not A267)  and  (not A203) );
 a14268a <=( A299  and  A298 );
 a14269a <=( (not A269)  and  a14268a );
 a14270a <=( a14269a  and  a14264a );
 a14273a <=( (not A166)  and  (not A167) );
 a14277a <=( A201  and  A200 );
 a14278a <=( (not A199)  and  a14277a );
 a14279a <=( a14278a  and  a14273a );
 a14282a <=( (not A267)  and  (not A203) );
 a14286a <=( (not A299)  and  (not A298) );
 a14287a <=( (not A269)  and  a14286a );
 a14288a <=( a14287a  and  a14282a );
 a14291a <=( (not A166)  and  (not A167) );
 a14295a <=( A201  and  A200 );
 a14296a <=( (not A199)  and  a14295a );
 a14297a <=( a14296a  and  a14291a );
 a14300a <=( A265  and  (not A203) );
 a14304a <=( A301  and  (not A300) );
 a14305a <=( A266  and  a14304a );
 a14306a <=( a14305a  and  a14300a );
 a14309a <=( (not A166)  and  (not A167) );
 a14313a <=( A201  and  A200 );
 a14314a <=( (not A199)  and  a14313a );
 a14315a <=( a14314a  and  a14309a );
 a14318a <=( A265  and  (not A203) );
 a14322a <=( (not A302)  and  (not A300) );
 a14323a <=( A266  and  a14322a );
 a14324a <=( a14323a  and  a14318a );
 a14327a <=( (not A166)  and  (not A167) );
 a14331a <=( A201  and  A200 );
 a14332a <=( (not A199)  and  a14331a );
 a14333a <=( a14332a  and  a14327a );
 a14336a <=( A265  and  (not A203) );
 a14340a <=( A299  and  A298 );
 a14341a <=( A266  and  a14340a );
 a14342a <=( a14341a  and  a14336a );
 a14345a <=( (not A166)  and  (not A167) );
 a14349a <=( A201  and  A200 );
 a14350a <=( (not A199)  and  a14349a );
 a14351a <=( a14350a  and  a14345a );
 a14354a <=( A265  and  (not A203) );
 a14358a <=( (not A299)  and  (not A298) );
 a14359a <=( A266  and  a14358a );
 a14360a <=( a14359a  and  a14354a );
 a14363a <=( (not A166)  and  (not A167) );
 a14367a <=( A201  and  A200 );
 a14368a <=( (not A199)  and  a14367a );
 a14369a <=( a14368a  and  a14363a );
 a14372a <=( (not A265)  and  (not A203) );
 a14376a <=( A301  and  (not A300) );
 a14377a <=( (not A266)  and  a14376a );
 a14378a <=( a14377a  and  a14372a );
 a14381a <=( (not A166)  and  (not A167) );
 a14385a <=( A201  and  A200 );
 a14386a <=( (not A199)  and  a14385a );
 a14387a <=( a14386a  and  a14381a );
 a14390a <=( (not A265)  and  (not A203) );
 a14394a <=( (not A302)  and  (not A300) );
 a14395a <=( (not A266)  and  a14394a );
 a14396a <=( a14395a  and  a14390a );
 a14399a <=( (not A166)  and  (not A167) );
 a14403a <=( A201  and  A200 );
 a14404a <=( (not A199)  and  a14403a );
 a14405a <=( a14404a  and  a14399a );
 a14408a <=( (not A265)  and  (not A203) );
 a14412a <=( A299  and  A298 );
 a14413a <=( (not A266)  and  a14412a );
 a14414a <=( a14413a  and  a14408a );
 a14417a <=( (not A166)  and  (not A167) );
 a14421a <=( A201  and  A200 );
 a14422a <=( (not A199)  and  a14421a );
 a14423a <=( a14422a  and  a14417a );
 a14426a <=( (not A265)  and  (not A203) );
 a14430a <=( (not A299)  and  (not A298) );
 a14431a <=( (not A266)  and  a14430a );
 a14432a <=( a14431a  and  a14426a );
 a14435a <=( (not A166)  and  (not A167) );
 a14439a <=( A201  and  (not A200) );
 a14440a <=( A199  and  a14439a );
 a14441a <=( a14440a  and  a14435a );
 a14444a <=( (not A267)  and  A202 );
 a14448a <=( A301  and  (not A300) );
 a14449a <=( A268  and  a14448a );
 a14450a <=( a14449a  and  a14444a );
 a14453a <=( (not A166)  and  (not A167) );
 a14457a <=( A201  and  (not A200) );
 a14458a <=( A199  and  a14457a );
 a14459a <=( a14458a  and  a14453a );
 a14462a <=( (not A267)  and  A202 );
 a14466a <=( (not A302)  and  (not A300) );
 a14467a <=( A268  and  a14466a );
 a14468a <=( a14467a  and  a14462a );
 a14471a <=( (not A166)  and  (not A167) );
 a14475a <=( A201  and  (not A200) );
 a14476a <=( A199  and  a14475a );
 a14477a <=( a14476a  and  a14471a );
 a14480a <=( (not A267)  and  A202 );
 a14484a <=( A299  and  A298 );
 a14485a <=( A268  and  a14484a );
 a14486a <=( a14485a  and  a14480a );
 a14489a <=( (not A166)  and  (not A167) );
 a14493a <=( A201  and  (not A200) );
 a14494a <=( A199  and  a14493a );
 a14495a <=( a14494a  and  a14489a );
 a14498a <=( (not A267)  and  A202 );
 a14502a <=( (not A299)  and  (not A298) );
 a14503a <=( A268  and  a14502a );
 a14504a <=( a14503a  and  a14498a );
 a14507a <=( (not A166)  and  (not A167) );
 a14511a <=( A201  and  (not A200) );
 a14512a <=( A199  and  a14511a );
 a14513a <=( a14512a  and  a14507a );
 a14516a <=( (not A267)  and  A202 );
 a14520a <=( A301  and  (not A300) );
 a14521a <=( (not A269)  and  a14520a );
 a14522a <=( a14521a  and  a14516a );
 a14525a <=( (not A166)  and  (not A167) );
 a14529a <=( A201  and  (not A200) );
 a14530a <=( A199  and  a14529a );
 a14531a <=( a14530a  and  a14525a );
 a14534a <=( (not A267)  and  A202 );
 a14538a <=( (not A302)  and  (not A300) );
 a14539a <=( (not A269)  and  a14538a );
 a14540a <=( a14539a  and  a14534a );
 a14543a <=( (not A166)  and  (not A167) );
 a14547a <=( A201  and  (not A200) );
 a14548a <=( A199  and  a14547a );
 a14549a <=( a14548a  and  a14543a );
 a14552a <=( (not A267)  and  A202 );
 a14556a <=( A299  and  A298 );
 a14557a <=( (not A269)  and  a14556a );
 a14558a <=( a14557a  and  a14552a );
 a14561a <=( (not A166)  and  (not A167) );
 a14565a <=( A201  and  (not A200) );
 a14566a <=( A199  and  a14565a );
 a14567a <=( a14566a  and  a14561a );
 a14570a <=( (not A267)  and  A202 );
 a14574a <=( (not A299)  and  (not A298) );
 a14575a <=( (not A269)  and  a14574a );
 a14576a <=( a14575a  and  a14570a );
 a14579a <=( (not A166)  and  (not A167) );
 a14583a <=( A201  and  (not A200) );
 a14584a <=( A199  and  a14583a );
 a14585a <=( a14584a  and  a14579a );
 a14588a <=( A265  and  A202 );
 a14592a <=( A301  and  (not A300) );
 a14593a <=( A266  and  a14592a );
 a14594a <=( a14593a  and  a14588a );
 a14597a <=( (not A166)  and  (not A167) );
 a14601a <=( A201  and  (not A200) );
 a14602a <=( A199  and  a14601a );
 a14603a <=( a14602a  and  a14597a );
 a14606a <=( A265  and  A202 );
 a14610a <=( (not A302)  and  (not A300) );
 a14611a <=( A266  and  a14610a );
 a14612a <=( a14611a  and  a14606a );
 a14615a <=( (not A166)  and  (not A167) );
 a14619a <=( A201  and  (not A200) );
 a14620a <=( A199  and  a14619a );
 a14621a <=( a14620a  and  a14615a );
 a14624a <=( A265  and  A202 );
 a14628a <=( A299  and  A298 );
 a14629a <=( A266  and  a14628a );
 a14630a <=( a14629a  and  a14624a );
 a14633a <=( (not A166)  and  (not A167) );
 a14637a <=( A201  and  (not A200) );
 a14638a <=( A199  and  a14637a );
 a14639a <=( a14638a  and  a14633a );
 a14642a <=( A265  and  A202 );
 a14646a <=( (not A299)  and  (not A298) );
 a14647a <=( A266  and  a14646a );
 a14648a <=( a14647a  and  a14642a );
 a14651a <=( (not A166)  and  (not A167) );
 a14655a <=( A201  and  (not A200) );
 a14656a <=( A199  and  a14655a );
 a14657a <=( a14656a  and  a14651a );
 a14660a <=( (not A265)  and  A202 );
 a14664a <=( A301  and  (not A300) );
 a14665a <=( (not A266)  and  a14664a );
 a14666a <=( a14665a  and  a14660a );
 a14669a <=( (not A166)  and  (not A167) );
 a14673a <=( A201  and  (not A200) );
 a14674a <=( A199  and  a14673a );
 a14675a <=( a14674a  and  a14669a );
 a14678a <=( (not A265)  and  A202 );
 a14682a <=( (not A302)  and  (not A300) );
 a14683a <=( (not A266)  and  a14682a );
 a14684a <=( a14683a  and  a14678a );
 a14687a <=( (not A166)  and  (not A167) );
 a14691a <=( A201  and  (not A200) );
 a14692a <=( A199  and  a14691a );
 a14693a <=( a14692a  and  a14687a );
 a14696a <=( (not A265)  and  A202 );
 a14700a <=( A299  and  A298 );
 a14701a <=( (not A266)  and  a14700a );
 a14702a <=( a14701a  and  a14696a );
 a14705a <=( (not A166)  and  (not A167) );
 a14709a <=( A201  and  (not A200) );
 a14710a <=( A199  and  a14709a );
 a14711a <=( a14710a  and  a14705a );
 a14714a <=( (not A265)  and  A202 );
 a14718a <=( (not A299)  and  (not A298) );
 a14719a <=( (not A266)  and  a14718a );
 a14720a <=( a14719a  and  a14714a );
 a14723a <=( (not A166)  and  (not A167) );
 a14727a <=( A201  and  (not A200) );
 a14728a <=( A199  and  a14727a );
 a14729a <=( a14728a  and  a14723a );
 a14732a <=( (not A267)  and  (not A203) );
 a14736a <=( A301  and  (not A300) );
 a14737a <=( A268  and  a14736a );
 a14738a <=( a14737a  and  a14732a );
 a14741a <=( (not A166)  and  (not A167) );
 a14745a <=( A201  and  (not A200) );
 a14746a <=( A199  and  a14745a );
 a14747a <=( a14746a  and  a14741a );
 a14750a <=( (not A267)  and  (not A203) );
 a14754a <=( (not A302)  and  (not A300) );
 a14755a <=( A268  and  a14754a );
 a14756a <=( a14755a  and  a14750a );
 a14759a <=( (not A166)  and  (not A167) );
 a14763a <=( A201  and  (not A200) );
 a14764a <=( A199  and  a14763a );
 a14765a <=( a14764a  and  a14759a );
 a14768a <=( (not A267)  and  (not A203) );
 a14772a <=( A299  and  A298 );
 a14773a <=( A268  and  a14772a );
 a14774a <=( a14773a  and  a14768a );
 a14777a <=( (not A166)  and  (not A167) );
 a14781a <=( A201  and  (not A200) );
 a14782a <=( A199  and  a14781a );
 a14783a <=( a14782a  and  a14777a );
 a14786a <=( (not A267)  and  (not A203) );
 a14790a <=( (not A299)  and  (not A298) );
 a14791a <=( A268  and  a14790a );
 a14792a <=( a14791a  and  a14786a );
 a14795a <=( (not A166)  and  (not A167) );
 a14799a <=( A201  and  (not A200) );
 a14800a <=( A199  and  a14799a );
 a14801a <=( a14800a  and  a14795a );
 a14804a <=( (not A267)  and  (not A203) );
 a14808a <=( A301  and  (not A300) );
 a14809a <=( (not A269)  and  a14808a );
 a14810a <=( a14809a  and  a14804a );
 a14813a <=( (not A166)  and  (not A167) );
 a14817a <=( A201  and  (not A200) );
 a14818a <=( A199  and  a14817a );
 a14819a <=( a14818a  and  a14813a );
 a14822a <=( (not A267)  and  (not A203) );
 a14826a <=( (not A302)  and  (not A300) );
 a14827a <=( (not A269)  and  a14826a );
 a14828a <=( a14827a  and  a14822a );
 a14831a <=( (not A166)  and  (not A167) );
 a14835a <=( A201  and  (not A200) );
 a14836a <=( A199  and  a14835a );
 a14837a <=( a14836a  and  a14831a );
 a14840a <=( (not A267)  and  (not A203) );
 a14844a <=( A299  and  A298 );
 a14845a <=( (not A269)  and  a14844a );
 a14846a <=( a14845a  and  a14840a );
 a14849a <=( (not A166)  and  (not A167) );
 a14853a <=( A201  and  (not A200) );
 a14854a <=( A199  and  a14853a );
 a14855a <=( a14854a  and  a14849a );
 a14858a <=( (not A267)  and  (not A203) );
 a14862a <=( (not A299)  and  (not A298) );
 a14863a <=( (not A269)  and  a14862a );
 a14864a <=( a14863a  and  a14858a );
 a14867a <=( (not A166)  and  (not A167) );
 a14871a <=( A201  and  (not A200) );
 a14872a <=( A199  and  a14871a );
 a14873a <=( a14872a  and  a14867a );
 a14876a <=( A265  and  (not A203) );
 a14880a <=( A301  and  (not A300) );
 a14881a <=( A266  and  a14880a );
 a14882a <=( a14881a  and  a14876a );
 a14885a <=( (not A166)  and  (not A167) );
 a14889a <=( A201  and  (not A200) );
 a14890a <=( A199  and  a14889a );
 a14891a <=( a14890a  and  a14885a );
 a14894a <=( A265  and  (not A203) );
 a14898a <=( (not A302)  and  (not A300) );
 a14899a <=( A266  and  a14898a );
 a14900a <=( a14899a  and  a14894a );
 a14903a <=( (not A166)  and  (not A167) );
 a14907a <=( A201  and  (not A200) );
 a14908a <=( A199  and  a14907a );
 a14909a <=( a14908a  and  a14903a );
 a14912a <=( A265  and  (not A203) );
 a14916a <=( A299  and  A298 );
 a14917a <=( A266  and  a14916a );
 a14918a <=( a14917a  and  a14912a );
 a14921a <=( (not A166)  and  (not A167) );
 a14925a <=( A201  and  (not A200) );
 a14926a <=( A199  and  a14925a );
 a14927a <=( a14926a  and  a14921a );
 a14930a <=( A265  and  (not A203) );
 a14934a <=( (not A299)  and  (not A298) );
 a14935a <=( A266  and  a14934a );
 a14936a <=( a14935a  and  a14930a );
 a14939a <=( (not A166)  and  (not A167) );
 a14943a <=( A201  and  (not A200) );
 a14944a <=( A199  and  a14943a );
 a14945a <=( a14944a  and  a14939a );
 a14948a <=( (not A265)  and  (not A203) );
 a14952a <=( A301  and  (not A300) );
 a14953a <=( (not A266)  and  a14952a );
 a14954a <=( a14953a  and  a14948a );
 a14957a <=( (not A166)  and  (not A167) );
 a14961a <=( A201  and  (not A200) );
 a14962a <=( A199  and  a14961a );
 a14963a <=( a14962a  and  a14957a );
 a14966a <=( (not A265)  and  (not A203) );
 a14970a <=( (not A302)  and  (not A300) );
 a14971a <=( (not A266)  and  a14970a );
 a14972a <=( a14971a  and  a14966a );
 a14975a <=( (not A166)  and  (not A167) );
 a14979a <=( A201  and  (not A200) );
 a14980a <=( A199  and  a14979a );
 a14981a <=( a14980a  and  a14975a );
 a14984a <=( (not A265)  and  (not A203) );
 a14988a <=( A299  and  A298 );
 a14989a <=( (not A266)  and  a14988a );
 a14990a <=( a14989a  and  a14984a );
 a14993a <=( (not A166)  and  (not A167) );
 a14997a <=( A201  and  (not A200) );
 a14998a <=( A199  and  a14997a );
 a14999a <=( a14998a  and  a14993a );
 a15002a <=( (not A265)  and  (not A203) );
 a15006a <=( (not A299)  and  (not A298) );
 a15007a <=( (not A266)  and  a15006a );
 a15008a <=( a15007a  and  a15002a );
 a15011a <=( (not A232)  and  (not A168) );
 a15015a <=( A235  and  A234 );
 a15016a <=( A233  and  a15015a );
 a15017a <=( a15016a  and  a15011a );
 a15020a <=( A266  and  (not A265) );
 a15024a <=( A269  and  (not A268) );
 a15025a <=( (not A267)  and  a15024a );
 a15026a <=( a15025a  and  a15020a );
 a15029a <=( (not A232)  and  (not A168) );
 a15033a <=( A235  and  A234 );
 a15034a <=( A233  and  a15033a );
 a15035a <=( a15034a  and  a15029a );
 a15038a <=( (not A266)  and  A265 );
 a15042a <=( A269  and  (not A268) );
 a15043a <=( (not A267)  and  a15042a );
 a15044a <=( a15043a  and  a15038a );
 a15047a <=( (not A232)  and  (not A168) );
 a15051a <=( (not A236)  and  A234 );
 a15052a <=( A233  and  a15051a );
 a15053a <=( a15052a  and  a15047a );
 a15056a <=( A266  and  (not A265) );
 a15060a <=( A269  and  (not A268) );
 a15061a <=( (not A267)  and  a15060a );
 a15062a <=( a15061a  and  a15056a );
 a15065a <=( (not A232)  and  (not A168) );
 a15069a <=( (not A236)  and  A234 );
 a15070a <=( A233  and  a15069a );
 a15071a <=( a15070a  and  a15065a );
 a15074a <=( (not A266)  and  A265 );
 a15078a <=( A269  and  (not A268) );
 a15079a <=( (not A267)  and  a15078a );
 a15080a <=( a15079a  and  a15074a );
 a15083a <=( A232  and  (not A168) );
 a15087a <=( A235  and  A234 );
 a15088a <=( (not A233)  and  a15087a );
 a15089a <=( a15088a  and  a15083a );
 a15092a <=( A266  and  (not A265) );
 a15096a <=( A269  and  (not A268) );
 a15097a <=( (not A267)  and  a15096a );
 a15098a <=( a15097a  and  a15092a );
 a15101a <=( A232  and  (not A168) );
 a15105a <=( A235  and  A234 );
 a15106a <=( (not A233)  and  a15105a );
 a15107a <=( a15106a  and  a15101a );
 a15110a <=( (not A266)  and  A265 );
 a15114a <=( A269  and  (not A268) );
 a15115a <=( (not A267)  and  a15114a );
 a15116a <=( a15115a  and  a15110a );
 a15119a <=( A232  and  (not A168) );
 a15123a <=( (not A236)  and  A234 );
 a15124a <=( (not A233)  and  a15123a );
 a15125a <=( a15124a  and  a15119a );
 a15128a <=( A266  and  (not A265) );
 a15132a <=( A269  and  (not A268) );
 a15133a <=( (not A267)  and  a15132a );
 a15134a <=( a15133a  and  a15128a );
 a15137a <=( A232  and  (not A168) );
 a15141a <=( (not A236)  and  A234 );
 a15142a <=( (not A233)  and  a15141a );
 a15143a <=( a15142a  and  a15137a );
 a15146a <=( (not A266)  and  A265 );
 a15150a <=( A269  and  (not A268) );
 a15151a <=( (not A267)  and  a15150a );
 a15152a <=( a15151a  and  a15146a );
 a15155a <=( (not A168)  and  A170 );
 a15159a <=( A201  and  A200 );
 a15160a <=( (not A199)  and  a15159a );
 a15161a <=( a15160a  and  a15155a );
 a15164a <=( (not A267)  and  A202 );
 a15168a <=( A301  and  (not A300) );
 a15169a <=( A268  and  a15168a );
 a15170a <=( a15169a  and  a15164a );
 a15173a <=( (not A168)  and  A170 );
 a15177a <=( A201  and  A200 );
 a15178a <=( (not A199)  and  a15177a );
 a15179a <=( a15178a  and  a15173a );
 a15182a <=( (not A267)  and  A202 );
 a15186a <=( (not A302)  and  (not A300) );
 a15187a <=( A268  and  a15186a );
 a15188a <=( a15187a  and  a15182a );
 a15191a <=( (not A168)  and  A170 );
 a15195a <=( A201  and  A200 );
 a15196a <=( (not A199)  and  a15195a );
 a15197a <=( a15196a  and  a15191a );
 a15200a <=( (not A267)  and  A202 );
 a15204a <=( A299  and  A298 );
 a15205a <=( A268  and  a15204a );
 a15206a <=( a15205a  and  a15200a );
 a15209a <=( (not A168)  and  A170 );
 a15213a <=( A201  and  A200 );
 a15214a <=( (not A199)  and  a15213a );
 a15215a <=( a15214a  and  a15209a );
 a15218a <=( (not A267)  and  A202 );
 a15222a <=( (not A299)  and  (not A298) );
 a15223a <=( A268  and  a15222a );
 a15224a <=( a15223a  and  a15218a );
 a15227a <=( (not A168)  and  A170 );
 a15231a <=( A201  and  A200 );
 a15232a <=( (not A199)  and  a15231a );
 a15233a <=( a15232a  and  a15227a );
 a15236a <=( (not A267)  and  A202 );
 a15240a <=( A301  and  (not A300) );
 a15241a <=( (not A269)  and  a15240a );
 a15242a <=( a15241a  and  a15236a );
 a15245a <=( (not A168)  and  A170 );
 a15249a <=( A201  and  A200 );
 a15250a <=( (not A199)  and  a15249a );
 a15251a <=( a15250a  and  a15245a );
 a15254a <=( (not A267)  and  A202 );
 a15258a <=( (not A302)  and  (not A300) );
 a15259a <=( (not A269)  and  a15258a );
 a15260a <=( a15259a  and  a15254a );
 a15263a <=( (not A168)  and  A170 );
 a15267a <=( A201  and  A200 );
 a15268a <=( (not A199)  and  a15267a );
 a15269a <=( a15268a  and  a15263a );
 a15272a <=( (not A267)  and  A202 );
 a15276a <=( A299  and  A298 );
 a15277a <=( (not A269)  and  a15276a );
 a15278a <=( a15277a  and  a15272a );
 a15281a <=( (not A168)  and  A170 );
 a15285a <=( A201  and  A200 );
 a15286a <=( (not A199)  and  a15285a );
 a15287a <=( a15286a  and  a15281a );
 a15290a <=( (not A267)  and  A202 );
 a15294a <=( (not A299)  and  (not A298) );
 a15295a <=( (not A269)  and  a15294a );
 a15296a <=( a15295a  and  a15290a );
 a15299a <=( (not A168)  and  A170 );
 a15303a <=( A201  and  A200 );
 a15304a <=( (not A199)  and  a15303a );
 a15305a <=( a15304a  and  a15299a );
 a15308a <=( A265  and  A202 );
 a15312a <=( A301  and  (not A300) );
 a15313a <=( A266  and  a15312a );
 a15314a <=( a15313a  and  a15308a );
 a15317a <=( (not A168)  and  A170 );
 a15321a <=( A201  and  A200 );
 a15322a <=( (not A199)  and  a15321a );
 a15323a <=( a15322a  and  a15317a );
 a15326a <=( A265  and  A202 );
 a15330a <=( (not A302)  and  (not A300) );
 a15331a <=( A266  and  a15330a );
 a15332a <=( a15331a  and  a15326a );
 a15335a <=( (not A168)  and  A170 );
 a15339a <=( A201  and  A200 );
 a15340a <=( (not A199)  and  a15339a );
 a15341a <=( a15340a  and  a15335a );
 a15344a <=( A265  and  A202 );
 a15348a <=( A299  and  A298 );
 a15349a <=( A266  and  a15348a );
 a15350a <=( a15349a  and  a15344a );
 a15353a <=( (not A168)  and  A170 );
 a15357a <=( A201  and  A200 );
 a15358a <=( (not A199)  and  a15357a );
 a15359a <=( a15358a  and  a15353a );
 a15362a <=( A265  and  A202 );
 a15366a <=( (not A299)  and  (not A298) );
 a15367a <=( A266  and  a15366a );
 a15368a <=( a15367a  and  a15362a );
 a15371a <=( (not A168)  and  A170 );
 a15375a <=( A201  and  A200 );
 a15376a <=( (not A199)  and  a15375a );
 a15377a <=( a15376a  and  a15371a );
 a15380a <=( (not A265)  and  A202 );
 a15384a <=( A301  and  (not A300) );
 a15385a <=( (not A266)  and  a15384a );
 a15386a <=( a15385a  and  a15380a );
 a15389a <=( (not A168)  and  A170 );
 a15393a <=( A201  and  A200 );
 a15394a <=( (not A199)  and  a15393a );
 a15395a <=( a15394a  and  a15389a );
 a15398a <=( (not A265)  and  A202 );
 a15402a <=( (not A302)  and  (not A300) );
 a15403a <=( (not A266)  and  a15402a );
 a15404a <=( a15403a  and  a15398a );
 a15407a <=( (not A168)  and  A170 );
 a15411a <=( A201  and  A200 );
 a15412a <=( (not A199)  and  a15411a );
 a15413a <=( a15412a  and  a15407a );
 a15416a <=( (not A265)  and  A202 );
 a15420a <=( A299  and  A298 );
 a15421a <=( (not A266)  and  a15420a );
 a15422a <=( a15421a  and  a15416a );
 a15425a <=( (not A168)  and  A170 );
 a15429a <=( A201  and  A200 );
 a15430a <=( (not A199)  and  a15429a );
 a15431a <=( a15430a  and  a15425a );
 a15434a <=( (not A265)  and  A202 );
 a15438a <=( (not A299)  and  (not A298) );
 a15439a <=( (not A266)  and  a15438a );
 a15440a <=( a15439a  and  a15434a );
 a15443a <=( (not A168)  and  A170 );
 a15447a <=( A201  and  A200 );
 a15448a <=( (not A199)  and  a15447a );
 a15449a <=( a15448a  and  a15443a );
 a15452a <=( (not A267)  and  (not A203) );
 a15456a <=( A301  and  (not A300) );
 a15457a <=( A268  and  a15456a );
 a15458a <=( a15457a  and  a15452a );
 a15461a <=( (not A168)  and  A170 );
 a15465a <=( A201  and  A200 );
 a15466a <=( (not A199)  and  a15465a );
 a15467a <=( a15466a  and  a15461a );
 a15470a <=( (not A267)  and  (not A203) );
 a15474a <=( (not A302)  and  (not A300) );
 a15475a <=( A268  and  a15474a );
 a15476a <=( a15475a  and  a15470a );
 a15479a <=( (not A168)  and  A170 );
 a15483a <=( A201  and  A200 );
 a15484a <=( (not A199)  and  a15483a );
 a15485a <=( a15484a  and  a15479a );
 a15488a <=( (not A267)  and  (not A203) );
 a15492a <=( A299  and  A298 );
 a15493a <=( A268  and  a15492a );
 a15494a <=( a15493a  and  a15488a );
 a15497a <=( (not A168)  and  A170 );
 a15501a <=( A201  and  A200 );
 a15502a <=( (not A199)  and  a15501a );
 a15503a <=( a15502a  and  a15497a );
 a15506a <=( (not A267)  and  (not A203) );
 a15510a <=( (not A299)  and  (not A298) );
 a15511a <=( A268  and  a15510a );
 a15512a <=( a15511a  and  a15506a );
 a15515a <=( (not A168)  and  A170 );
 a15519a <=( A201  and  A200 );
 a15520a <=( (not A199)  and  a15519a );
 a15521a <=( a15520a  and  a15515a );
 a15524a <=( (not A267)  and  (not A203) );
 a15528a <=( A301  and  (not A300) );
 a15529a <=( (not A269)  and  a15528a );
 a15530a <=( a15529a  and  a15524a );
 a15533a <=( (not A168)  and  A170 );
 a15537a <=( A201  and  A200 );
 a15538a <=( (not A199)  and  a15537a );
 a15539a <=( a15538a  and  a15533a );
 a15542a <=( (not A267)  and  (not A203) );
 a15546a <=( (not A302)  and  (not A300) );
 a15547a <=( (not A269)  and  a15546a );
 a15548a <=( a15547a  and  a15542a );
 a15551a <=( (not A168)  and  A170 );
 a15555a <=( A201  and  A200 );
 a15556a <=( (not A199)  and  a15555a );
 a15557a <=( a15556a  and  a15551a );
 a15560a <=( (not A267)  and  (not A203) );
 a15564a <=( A299  and  A298 );
 a15565a <=( (not A269)  and  a15564a );
 a15566a <=( a15565a  and  a15560a );
 a15569a <=( (not A168)  and  A170 );
 a15573a <=( A201  and  A200 );
 a15574a <=( (not A199)  and  a15573a );
 a15575a <=( a15574a  and  a15569a );
 a15578a <=( (not A267)  and  (not A203) );
 a15582a <=( (not A299)  and  (not A298) );
 a15583a <=( (not A269)  and  a15582a );
 a15584a <=( a15583a  and  a15578a );
 a15587a <=( (not A168)  and  A170 );
 a15591a <=( A201  and  A200 );
 a15592a <=( (not A199)  and  a15591a );
 a15593a <=( a15592a  and  a15587a );
 a15596a <=( A265  and  (not A203) );
 a15600a <=( A301  and  (not A300) );
 a15601a <=( A266  and  a15600a );
 a15602a <=( a15601a  and  a15596a );
 a15605a <=( (not A168)  and  A170 );
 a15609a <=( A201  and  A200 );
 a15610a <=( (not A199)  and  a15609a );
 a15611a <=( a15610a  and  a15605a );
 a15614a <=( A265  and  (not A203) );
 a15618a <=( (not A302)  and  (not A300) );
 a15619a <=( A266  and  a15618a );
 a15620a <=( a15619a  and  a15614a );
 a15623a <=( (not A168)  and  A170 );
 a15627a <=( A201  and  A200 );
 a15628a <=( (not A199)  and  a15627a );
 a15629a <=( a15628a  and  a15623a );
 a15632a <=( A265  and  (not A203) );
 a15636a <=( A299  and  A298 );
 a15637a <=( A266  and  a15636a );
 a15638a <=( a15637a  and  a15632a );
 a15641a <=( (not A168)  and  A170 );
 a15645a <=( A201  and  A200 );
 a15646a <=( (not A199)  and  a15645a );
 a15647a <=( a15646a  and  a15641a );
 a15650a <=( A265  and  (not A203) );
 a15654a <=( (not A299)  and  (not A298) );
 a15655a <=( A266  and  a15654a );
 a15656a <=( a15655a  and  a15650a );
 a15659a <=( (not A168)  and  A170 );
 a15663a <=( A201  and  A200 );
 a15664a <=( (not A199)  and  a15663a );
 a15665a <=( a15664a  and  a15659a );
 a15668a <=( (not A265)  and  (not A203) );
 a15672a <=( A301  and  (not A300) );
 a15673a <=( (not A266)  and  a15672a );
 a15674a <=( a15673a  and  a15668a );
 a15677a <=( (not A168)  and  A170 );
 a15681a <=( A201  and  A200 );
 a15682a <=( (not A199)  and  a15681a );
 a15683a <=( a15682a  and  a15677a );
 a15686a <=( (not A265)  and  (not A203) );
 a15690a <=( (not A302)  and  (not A300) );
 a15691a <=( (not A266)  and  a15690a );
 a15692a <=( a15691a  and  a15686a );
 a15695a <=( (not A168)  and  A170 );
 a15699a <=( A201  and  A200 );
 a15700a <=( (not A199)  and  a15699a );
 a15701a <=( a15700a  and  a15695a );
 a15704a <=( (not A265)  and  (not A203) );
 a15708a <=( A299  and  A298 );
 a15709a <=( (not A266)  and  a15708a );
 a15710a <=( a15709a  and  a15704a );
 a15713a <=( (not A168)  and  A170 );
 a15717a <=( A201  and  A200 );
 a15718a <=( (not A199)  and  a15717a );
 a15719a <=( a15718a  and  a15713a );
 a15722a <=( (not A265)  and  (not A203) );
 a15726a <=( (not A299)  and  (not A298) );
 a15727a <=( (not A266)  and  a15726a );
 a15728a <=( a15727a  and  a15722a );
 a15731a <=( (not A168)  and  A170 );
 a15735a <=( A201  and  (not A200) );
 a15736a <=( A199  and  a15735a );
 a15737a <=( a15736a  and  a15731a );
 a15740a <=( (not A267)  and  A202 );
 a15744a <=( A301  and  (not A300) );
 a15745a <=( A268  and  a15744a );
 a15746a <=( a15745a  and  a15740a );
 a15749a <=( (not A168)  and  A170 );
 a15753a <=( A201  and  (not A200) );
 a15754a <=( A199  and  a15753a );
 a15755a <=( a15754a  and  a15749a );
 a15758a <=( (not A267)  and  A202 );
 a15762a <=( (not A302)  and  (not A300) );
 a15763a <=( A268  and  a15762a );
 a15764a <=( a15763a  and  a15758a );
 a15767a <=( (not A168)  and  A170 );
 a15771a <=( A201  and  (not A200) );
 a15772a <=( A199  and  a15771a );
 a15773a <=( a15772a  and  a15767a );
 a15776a <=( (not A267)  and  A202 );
 a15780a <=( A299  and  A298 );
 a15781a <=( A268  and  a15780a );
 a15782a <=( a15781a  and  a15776a );
 a15785a <=( (not A168)  and  A170 );
 a15789a <=( A201  and  (not A200) );
 a15790a <=( A199  and  a15789a );
 a15791a <=( a15790a  and  a15785a );
 a15794a <=( (not A267)  and  A202 );
 a15798a <=( (not A299)  and  (not A298) );
 a15799a <=( A268  and  a15798a );
 a15800a <=( a15799a  and  a15794a );
 a15803a <=( (not A168)  and  A170 );
 a15807a <=( A201  and  (not A200) );
 a15808a <=( A199  and  a15807a );
 a15809a <=( a15808a  and  a15803a );
 a15812a <=( (not A267)  and  A202 );
 a15816a <=( A301  and  (not A300) );
 a15817a <=( (not A269)  and  a15816a );
 a15818a <=( a15817a  and  a15812a );
 a15821a <=( (not A168)  and  A170 );
 a15825a <=( A201  and  (not A200) );
 a15826a <=( A199  and  a15825a );
 a15827a <=( a15826a  and  a15821a );
 a15830a <=( (not A267)  and  A202 );
 a15834a <=( (not A302)  and  (not A300) );
 a15835a <=( (not A269)  and  a15834a );
 a15836a <=( a15835a  and  a15830a );
 a15839a <=( (not A168)  and  A170 );
 a15843a <=( A201  and  (not A200) );
 a15844a <=( A199  and  a15843a );
 a15845a <=( a15844a  and  a15839a );
 a15848a <=( (not A267)  and  A202 );
 a15852a <=( A299  and  A298 );
 a15853a <=( (not A269)  and  a15852a );
 a15854a <=( a15853a  and  a15848a );
 a15857a <=( (not A168)  and  A170 );
 a15861a <=( A201  and  (not A200) );
 a15862a <=( A199  and  a15861a );
 a15863a <=( a15862a  and  a15857a );
 a15866a <=( (not A267)  and  A202 );
 a15870a <=( (not A299)  and  (not A298) );
 a15871a <=( (not A269)  and  a15870a );
 a15872a <=( a15871a  and  a15866a );
 a15875a <=( (not A168)  and  A170 );
 a15879a <=( A201  and  (not A200) );
 a15880a <=( A199  and  a15879a );
 a15881a <=( a15880a  and  a15875a );
 a15884a <=( A265  and  A202 );
 a15888a <=( A301  and  (not A300) );
 a15889a <=( A266  and  a15888a );
 a15890a <=( a15889a  and  a15884a );
 a15893a <=( (not A168)  and  A170 );
 a15897a <=( A201  and  (not A200) );
 a15898a <=( A199  and  a15897a );
 a15899a <=( a15898a  and  a15893a );
 a15902a <=( A265  and  A202 );
 a15906a <=( (not A302)  and  (not A300) );
 a15907a <=( A266  and  a15906a );
 a15908a <=( a15907a  and  a15902a );
 a15911a <=( (not A168)  and  A170 );
 a15915a <=( A201  and  (not A200) );
 a15916a <=( A199  and  a15915a );
 a15917a <=( a15916a  and  a15911a );
 a15920a <=( A265  and  A202 );
 a15924a <=( A299  and  A298 );
 a15925a <=( A266  and  a15924a );
 a15926a <=( a15925a  and  a15920a );
 a15929a <=( (not A168)  and  A170 );
 a15933a <=( A201  and  (not A200) );
 a15934a <=( A199  and  a15933a );
 a15935a <=( a15934a  and  a15929a );
 a15938a <=( A265  and  A202 );
 a15942a <=( (not A299)  and  (not A298) );
 a15943a <=( A266  and  a15942a );
 a15944a <=( a15943a  and  a15938a );
 a15947a <=( (not A168)  and  A170 );
 a15951a <=( A201  and  (not A200) );
 a15952a <=( A199  and  a15951a );
 a15953a <=( a15952a  and  a15947a );
 a15956a <=( (not A265)  and  A202 );
 a15960a <=( A301  and  (not A300) );
 a15961a <=( (not A266)  and  a15960a );
 a15962a <=( a15961a  and  a15956a );
 a15965a <=( (not A168)  and  A170 );
 a15969a <=( A201  and  (not A200) );
 a15970a <=( A199  and  a15969a );
 a15971a <=( a15970a  and  a15965a );
 a15974a <=( (not A265)  and  A202 );
 a15978a <=( (not A302)  and  (not A300) );
 a15979a <=( (not A266)  and  a15978a );
 a15980a <=( a15979a  and  a15974a );
 a15983a <=( (not A168)  and  A170 );
 a15987a <=( A201  and  (not A200) );
 a15988a <=( A199  and  a15987a );
 a15989a <=( a15988a  and  a15983a );
 a15992a <=( (not A265)  and  A202 );
 a15996a <=( A299  and  A298 );
 a15997a <=( (not A266)  and  a15996a );
 a15998a <=( a15997a  and  a15992a );
 a16001a <=( (not A168)  and  A170 );
 a16005a <=( A201  and  (not A200) );
 a16006a <=( A199  and  a16005a );
 a16007a <=( a16006a  and  a16001a );
 a16010a <=( (not A265)  and  A202 );
 a16014a <=( (not A299)  and  (not A298) );
 a16015a <=( (not A266)  and  a16014a );
 a16016a <=( a16015a  and  a16010a );
 a16019a <=( (not A168)  and  A170 );
 a16023a <=( A201  and  (not A200) );
 a16024a <=( A199  and  a16023a );
 a16025a <=( a16024a  and  a16019a );
 a16028a <=( (not A267)  and  (not A203) );
 a16032a <=( A301  and  (not A300) );
 a16033a <=( A268  and  a16032a );
 a16034a <=( a16033a  and  a16028a );
 a16037a <=( (not A168)  and  A170 );
 a16041a <=( A201  and  (not A200) );
 a16042a <=( A199  and  a16041a );
 a16043a <=( a16042a  and  a16037a );
 a16046a <=( (not A267)  and  (not A203) );
 a16050a <=( (not A302)  and  (not A300) );
 a16051a <=( A268  and  a16050a );
 a16052a <=( a16051a  and  a16046a );
 a16055a <=( (not A168)  and  A170 );
 a16059a <=( A201  and  (not A200) );
 a16060a <=( A199  and  a16059a );
 a16061a <=( a16060a  and  a16055a );
 a16064a <=( (not A267)  and  (not A203) );
 a16068a <=( A299  and  A298 );
 a16069a <=( A268  and  a16068a );
 a16070a <=( a16069a  and  a16064a );
 a16073a <=( (not A168)  and  A170 );
 a16077a <=( A201  and  (not A200) );
 a16078a <=( A199  and  a16077a );
 a16079a <=( a16078a  and  a16073a );
 a16082a <=( (not A267)  and  (not A203) );
 a16086a <=( (not A299)  and  (not A298) );
 a16087a <=( A268  and  a16086a );
 a16088a <=( a16087a  and  a16082a );
 a16091a <=( (not A168)  and  A170 );
 a16095a <=( A201  and  (not A200) );
 a16096a <=( A199  and  a16095a );
 a16097a <=( a16096a  and  a16091a );
 a16100a <=( (not A267)  and  (not A203) );
 a16104a <=( A301  and  (not A300) );
 a16105a <=( (not A269)  and  a16104a );
 a16106a <=( a16105a  and  a16100a );
 a16109a <=( (not A168)  and  A170 );
 a16113a <=( A201  and  (not A200) );
 a16114a <=( A199  and  a16113a );
 a16115a <=( a16114a  and  a16109a );
 a16118a <=( (not A267)  and  (not A203) );
 a16122a <=( (not A302)  and  (not A300) );
 a16123a <=( (not A269)  and  a16122a );
 a16124a <=( a16123a  and  a16118a );
 a16127a <=( (not A168)  and  A170 );
 a16131a <=( A201  and  (not A200) );
 a16132a <=( A199  and  a16131a );
 a16133a <=( a16132a  and  a16127a );
 a16136a <=( (not A267)  and  (not A203) );
 a16140a <=( A299  and  A298 );
 a16141a <=( (not A269)  and  a16140a );
 a16142a <=( a16141a  and  a16136a );
 a16145a <=( (not A168)  and  A170 );
 a16149a <=( A201  and  (not A200) );
 a16150a <=( A199  and  a16149a );
 a16151a <=( a16150a  and  a16145a );
 a16154a <=( (not A267)  and  (not A203) );
 a16158a <=( (not A299)  and  (not A298) );
 a16159a <=( (not A269)  and  a16158a );
 a16160a <=( a16159a  and  a16154a );
 a16163a <=( (not A168)  and  A170 );
 a16167a <=( A201  and  (not A200) );
 a16168a <=( A199  and  a16167a );
 a16169a <=( a16168a  and  a16163a );
 a16172a <=( A265  and  (not A203) );
 a16176a <=( A301  and  (not A300) );
 a16177a <=( A266  and  a16176a );
 a16178a <=( a16177a  and  a16172a );
 a16181a <=( (not A168)  and  A170 );
 a16185a <=( A201  and  (not A200) );
 a16186a <=( A199  and  a16185a );
 a16187a <=( a16186a  and  a16181a );
 a16190a <=( A265  and  (not A203) );
 a16194a <=( (not A302)  and  (not A300) );
 a16195a <=( A266  and  a16194a );
 a16196a <=( a16195a  and  a16190a );
 a16199a <=( (not A168)  and  A170 );
 a16203a <=( A201  and  (not A200) );
 a16204a <=( A199  and  a16203a );
 a16205a <=( a16204a  and  a16199a );
 a16208a <=( A265  and  (not A203) );
 a16212a <=( A299  and  A298 );
 a16213a <=( A266  and  a16212a );
 a16214a <=( a16213a  and  a16208a );
 a16217a <=( (not A168)  and  A170 );
 a16221a <=( A201  and  (not A200) );
 a16222a <=( A199  and  a16221a );
 a16223a <=( a16222a  and  a16217a );
 a16226a <=( A265  and  (not A203) );
 a16230a <=( (not A299)  and  (not A298) );
 a16231a <=( A266  and  a16230a );
 a16232a <=( a16231a  and  a16226a );
 a16235a <=( (not A168)  and  A170 );
 a16239a <=( A201  and  (not A200) );
 a16240a <=( A199  and  a16239a );
 a16241a <=( a16240a  and  a16235a );
 a16244a <=( (not A265)  and  (not A203) );
 a16248a <=( A301  and  (not A300) );
 a16249a <=( (not A266)  and  a16248a );
 a16250a <=( a16249a  and  a16244a );
 a16253a <=( (not A168)  and  A170 );
 a16257a <=( A201  and  (not A200) );
 a16258a <=( A199  and  a16257a );
 a16259a <=( a16258a  and  a16253a );
 a16262a <=( (not A265)  and  (not A203) );
 a16266a <=( (not A302)  and  (not A300) );
 a16267a <=( (not A266)  and  a16266a );
 a16268a <=( a16267a  and  a16262a );
 a16271a <=( (not A168)  and  A170 );
 a16275a <=( A201  and  (not A200) );
 a16276a <=( A199  and  a16275a );
 a16277a <=( a16276a  and  a16271a );
 a16280a <=( (not A265)  and  (not A203) );
 a16284a <=( A299  and  A298 );
 a16285a <=( (not A266)  and  a16284a );
 a16286a <=( a16285a  and  a16280a );
 a16289a <=( (not A168)  and  A170 );
 a16293a <=( A201  and  (not A200) );
 a16294a <=( A199  and  a16293a );
 a16295a <=( a16294a  and  a16289a );
 a16298a <=( (not A265)  and  (not A203) );
 a16302a <=( (not A299)  and  (not A298) );
 a16303a <=( (not A266)  and  a16302a );
 a16304a <=( a16303a  and  a16298a );
 a16307a <=( (not A168)  and  A169 );
 a16311a <=( A201  and  A200 );
 a16312a <=( (not A199)  and  a16311a );
 a16313a <=( a16312a  and  a16307a );
 a16316a <=( (not A267)  and  A202 );
 a16320a <=( A301  and  (not A300) );
 a16321a <=( A268  and  a16320a );
 a16322a <=( a16321a  and  a16316a );
 a16325a <=( (not A168)  and  A169 );
 a16329a <=( A201  and  A200 );
 a16330a <=( (not A199)  and  a16329a );
 a16331a <=( a16330a  and  a16325a );
 a16334a <=( (not A267)  and  A202 );
 a16338a <=( (not A302)  and  (not A300) );
 a16339a <=( A268  and  a16338a );
 a16340a <=( a16339a  and  a16334a );
 a16343a <=( (not A168)  and  A169 );
 a16347a <=( A201  and  A200 );
 a16348a <=( (not A199)  and  a16347a );
 a16349a <=( a16348a  and  a16343a );
 a16352a <=( (not A267)  and  A202 );
 a16356a <=( A299  and  A298 );
 a16357a <=( A268  and  a16356a );
 a16358a <=( a16357a  and  a16352a );
 a16361a <=( (not A168)  and  A169 );
 a16365a <=( A201  and  A200 );
 a16366a <=( (not A199)  and  a16365a );
 a16367a <=( a16366a  and  a16361a );
 a16370a <=( (not A267)  and  A202 );
 a16374a <=( (not A299)  and  (not A298) );
 a16375a <=( A268  and  a16374a );
 a16376a <=( a16375a  and  a16370a );
 a16379a <=( (not A168)  and  A169 );
 a16383a <=( A201  and  A200 );
 a16384a <=( (not A199)  and  a16383a );
 a16385a <=( a16384a  and  a16379a );
 a16388a <=( (not A267)  and  A202 );
 a16392a <=( A301  and  (not A300) );
 a16393a <=( (not A269)  and  a16392a );
 a16394a <=( a16393a  and  a16388a );
 a16397a <=( (not A168)  and  A169 );
 a16401a <=( A201  and  A200 );
 a16402a <=( (not A199)  and  a16401a );
 a16403a <=( a16402a  and  a16397a );
 a16406a <=( (not A267)  and  A202 );
 a16410a <=( (not A302)  and  (not A300) );
 a16411a <=( (not A269)  and  a16410a );
 a16412a <=( a16411a  and  a16406a );
 a16415a <=( (not A168)  and  A169 );
 a16419a <=( A201  and  A200 );
 a16420a <=( (not A199)  and  a16419a );
 a16421a <=( a16420a  and  a16415a );
 a16424a <=( (not A267)  and  A202 );
 a16428a <=( A299  and  A298 );
 a16429a <=( (not A269)  and  a16428a );
 a16430a <=( a16429a  and  a16424a );
 a16433a <=( (not A168)  and  A169 );
 a16437a <=( A201  and  A200 );
 a16438a <=( (not A199)  and  a16437a );
 a16439a <=( a16438a  and  a16433a );
 a16442a <=( (not A267)  and  A202 );
 a16446a <=( (not A299)  and  (not A298) );
 a16447a <=( (not A269)  and  a16446a );
 a16448a <=( a16447a  and  a16442a );
 a16451a <=( (not A168)  and  A169 );
 a16455a <=( A201  and  A200 );
 a16456a <=( (not A199)  and  a16455a );
 a16457a <=( a16456a  and  a16451a );
 a16460a <=( A265  and  A202 );
 a16464a <=( A301  and  (not A300) );
 a16465a <=( A266  and  a16464a );
 a16466a <=( a16465a  and  a16460a );
 a16469a <=( (not A168)  and  A169 );
 a16473a <=( A201  and  A200 );
 a16474a <=( (not A199)  and  a16473a );
 a16475a <=( a16474a  and  a16469a );
 a16478a <=( A265  and  A202 );
 a16482a <=( (not A302)  and  (not A300) );
 a16483a <=( A266  and  a16482a );
 a16484a <=( a16483a  and  a16478a );
 a16487a <=( (not A168)  and  A169 );
 a16491a <=( A201  and  A200 );
 a16492a <=( (not A199)  and  a16491a );
 a16493a <=( a16492a  and  a16487a );
 a16496a <=( A265  and  A202 );
 a16500a <=( A299  and  A298 );
 a16501a <=( A266  and  a16500a );
 a16502a <=( a16501a  and  a16496a );
 a16505a <=( (not A168)  and  A169 );
 a16509a <=( A201  and  A200 );
 a16510a <=( (not A199)  and  a16509a );
 a16511a <=( a16510a  and  a16505a );
 a16514a <=( A265  and  A202 );
 a16518a <=( (not A299)  and  (not A298) );
 a16519a <=( A266  and  a16518a );
 a16520a <=( a16519a  and  a16514a );
 a16523a <=( (not A168)  and  A169 );
 a16527a <=( A201  and  A200 );
 a16528a <=( (not A199)  and  a16527a );
 a16529a <=( a16528a  and  a16523a );
 a16532a <=( (not A265)  and  A202 );
 a16536a <=( A301  and  (not A300) );
 a16537a <=( (not A266)  and  a16536a );
 a16538a <=( a16537a  and  a16532a );
 a16541a <=( (not A168)  and  A169 );
 a16545a <=( A201  and  A200 );
 a16546a <=( (not A199)  and  a16545a );
 a16547a <=( a16546a  and  a16541a );
 a16550a <=( (not A265)  and  A202 );
 a16554a <=( (not A302)  and  (not A300) );
 a16555a <=( (not A266)  and  a16554a );
 a16556a <=( a16555a  and  a16550a );
 a16559a <=( (not A168)  and  A169 );
 a16563a <=( A201  and  A200 );
 a16564a <=( (not A199)  and  a16563a );
 a16565a <=( a16564a  and  a16559a );
 a16568a <=( (not A265)  and  A202 );
 a16572a <=( A299  and  A298 );
 a16573a <=( (not A266)  and  a16572a );
 a16574a <=( a16573a  and  a16568a );
 a16577a <=( (not A168)  and  A169 );
 a16581a <=( A201  and  A200 );
 a16582a <=( (not A199)  and  a16581a );
 a16583a <=( a16582a  and  a16577a );
 a16586a <=( (not A265)  and  A202 );
 a16590a <=( (not A299)  and  (not A298) );
 a16591a <=( (not A266)  and  a16590a );
 a16592a <=( a16591a  and  a16586a );
 a16595a <=( (not A168)  and  A169 );
 a16599a <=( A201  and  A200 );
 a16600a <=( (not A199)  and  a16599a );
 a16601a <=( a16600a  and  a16595a );
 a16604a <=( (not A267)  and  (not A203) );
 a16608a <=( A301  and  (not A300) );
 a16609a <=( A268  and  a16608a );
 a16610a <=( a16609a  and  a16604a );
 a16613a <=( (not A168)  and  A169 );
 a16617a <=( A201  and  A200 );
 a16618a <=( (not A199)  and  a16617a );
 a16619a <=( a16618a  and  a16613a );
 a16622a <=( (not A267)  and  (not A203) );
 a16626a <=( (not A302)  and  (not A300) );
 a16627a <=( A268  and  a16626a );
 a16628a <=( a16627a  and  a16622a );
 a16631a <=( (not A168)  and  A169 );
 a16635a <=( A201  and  A200 );
 a16636a <=( (not A199)  and  a16635a );
 a16637a <=( a16636a  and  a16631a );
 a16640a <=( (not A267)  and  (not A203) );
 a16644a <=( A299  and  A298 );
 a16645a <=( A268  and  a16644a );
 a16646a <=( a16645a  and  a16640a );
 a16649a <=( (not A168)  and  A169 );
 a16653a <=( A201  and  A200 );
 a16654a <=( (not A199)  and  a16653a );
 a16655a <=( a16654a  and  a16649a );
 a16658a <=( (not A267)  and  (not A203) );
 a16662a <=( (not A299)  and  (not A298) );
 a16663a <=( A268  and  a16662a );
 a16664a <=( a16663a  and  a16658a );
 a16667a <=( (not A168)  and  A169 );
 a16671a <=( A201  and  A200 );
 a16672a <=( (not A199)  and  a16671a );
 a16673a <=( a16672a  and  a16667a );
 a16676a <=( (not A267)  and  (not A203) );
 a16680a <=( A301  and  (not A300) );
 a16681a <=( (not A269)  and  a16680a );
 a16682a <=( a16681a  and  a16676a );
 a16685a <=( (not A168)  and  A169 );
 a16689a <=( A201  and  A200 );
 a16690a <=( (not A199)  and  a16689a );
 a16691a <=( a16690a  and  a16685a );
 a16694a <=( (not A267)  and  (not A203) );
 a16698a <=( (not A302)  and  (not A300) );
 a16699a <=( (not A269)  and  a16698a );
 a16700a <=( a16699a  and  a16694a );
 a16703a <=( (not A168)  and  A169 );
 a16707a <=( A201  and  A200 );
 a16708a <=( (not A199)  and  a16707a );
 a16709a <=( a16708a  and  a16703a );
 a16712a <=( (not A267)  and  (not A203) );
 a16716a <=( A299  and  A298 );
 a16717a <=( (not A269)  and  a16716a );
 a16718a <=( a16717a  and  a16712a );
 a16721a <=( (not A168)  and  A169 );
 a16725a <=( A201  and  A200 );
 a16726a <=( (not A199)  and  a16725a );
 a16727a <=( a16726a  and  a16721a );
 a16730a <=( (not A267)  and  (not A203) );
 a16734a <=( (not A299)  and  (not A298) );
 a16735a <=( (not A269)  and  a16734a );
 a16736a <=( a16735a  and  a16730a );
 a16739a <=( (not A168)  and  A169 );
 a16743a <=( A201  and  A200 );
 a16744a <=( (not A199)  and  a16743a );
 a16745a <=( a16744a  and  a16739a );
 a16748a <=( A265  and  (not A203) );
 a16752a <=( A301  and  (not A300) );
 a16753a <=( A266  and  a16752a );
 a16754a <=( a16753a  and  a16748a );
 a16757a <=( (not A168)  and  A169 );
 a16761a <=( A201  and  A200 );
 a16762a <=( (not A199)  and  a16761a );
 a16763a <=( a16762a  and  a16757a );
 a16766a <=( A265  and  (not A203) );
 a16770a <=( (not A302)  and  (not A300) );
 a16771a <=( A266  and  a16770a );
 a16772a <=( a16771a  and  a16766a );
 a16775a <=( (not A168)  and  A169 );
 a16779a <=( A201  and  A200 );
 a16780a <=( (not A199)  and  a16779a );
 a16781a <=( a16780a  and  a16775a );
 a16784a <=( A265  and  (not A203) );
 a16788a <=( A299  and  A298 );
 a16789a <=( A266  and  a16788a );
 a16790a <=( a16789a  and  a16784a );
 a16793a <=( (not A168)  and  A169 );
 a16797a <=( A201  and  A200 );
 a16798a <=( (not A199)  and  a16797a );
 a16799a <=( a16798a  and  a16793a );
 a16802a <=( A265  and  (not A203) );
 a16806a <=( (not A299)  and  (not A298) );
 a16807a <=( A266  and  a16806a );
 a16808a <=( a16807a  and  a16802a );
 a16811a <=( (not A168)  and  A169 );
 a16815a <=( A201  and  A200 );
 a16816a <=( (not A199)  and  a16815a );
 a16817a <=( a16816a  and  a16811a );
 a16820a <=( (not A265)  and  (not A203) );
 a16824a <=( A301  and  (not A300) );
 a16825a <=( (not A266)  and  a16824a );
 a16826a <=( a16825a  and  a16820a );
 a16829a <=( (not A168)  and  A169 );
 a16833a <=( A201  and  A200 );
 a16834a <=( (not A199)  and  a16833a );
 a16835a <=( a16834a  and  a16829a );
 a16838a <=( (not A265)  and  (not A203) );
 a16842a <=( (not A302)  and  (not A300) );
 a16843a <=( (not A266)  and  a16842a );
 a16844a <=( a16843a  and  a16838a );
 a16847a <=( (not A168)  and  A169 );
 a16851a <=( A201  and  A200 );
 a16852a <=( (not A199)  and  a16851a );
 a16853a <=( a16852a  and  a16847a );
 a16856a <=( (not A265)  and  (not A203) );
 a16860a <=( A299  and  A298 );
 a16861a <=( (not A266)  and  a16860a );
 a16862a <=( a16861a  and  a16856a );
 a16865a <=( (not A168)  and  A169 );
 a16869a <=( A201  and  A200 );
 a16870a <=( (not A199)  and  a16869a );
 a16871a <=( a16870a  and  a16865a );
 a16874a <=( (not A265)  and  (not A203) );
 a16878a <=( (not A299)  and  (not A298) );
 a16879a <=( (not A266)  and  a16878a );
 a16880a <=( a16879a  and  a16874a );
 a16883a <=( (not A168)  and  A169 );
 a16887a <=( A201  and  (not A200) );
 a16888a <=( A199  and  a16887a );
 a16889a <=( a16888a  and  a16883a );
 a16892a <=( (not A267)  and  A202 );
 a16896a <=( A301  and  (not A300) );
 a16897a <=( A268  and  a16896a );
 a16898a <=( a16897a  and  a16892a );
 a16901a <=( (not A168)  and  A169 );
 a16905a <=( A201  and  (not A200) );
 a16906a <=( A199  and  a16905a );
 a16907a <=( a16906a  and  a16901a );
 a16910a <=( (not A267)  and  A202 );
 a16914a <=( (not A302)  and  (not A300) );
 a16915a <=( A268  and  a16914a );
 a16916a <=( a16915a  and  a16910a );
 a16919a <=( (not A168)  and  A169 );
 a16923a <=( A201  and  (not A200) );
 a16924a <=( A199  and  a16923a );
 a16925a <=( a16924a  and  a16919a );
 a16928a <=( (not A267)  and  A202 );
 a16932a <=( A299  and  A298 );
 a16933a <=( A268  and  a16932a );
 a16934a <=( a16933a  and  a16928a );
 a16937a <=( (not A168)  and  A169 );
 a16941a <=( A201  and  (not A200) );
 a16942a <=( A199  and  a16941a );
 a16943a <=( a16942a  and  a16937a );
 a16946a <=( (not A267)  and  A202 );
 a16950a <=( (not A299)  and  (not A298) );
 a16951a <=( A268  and  a16950a );
 a16952a <=( a16951a  and  a16946a );
 a16955a <=( (not A168)  and  A169 );
 a16959a <=( A201  and  (not A200) );
 a16960a <=( A199  and  a16959a );
 a16961a <=( a16960a  and  a16955a );
 a16964a <=( (not A267)  and  A202 );
 a16968a <=( A301  and  (not A300) );
 a16969a <=( (not A269)  and  a16968a );
 a16970a <=( a16969a  and  a16964a );
 a16973a <=( (not A168)  and  A169 );
 a16977a <=( A201  and  (not A200) );
 a16978a <=( A199  and  a16977a );
 a16979a <=( a16978a  and  a16973a );
 a16982a <=( (not A267)  and  A202 );
 a16986a <=( (not A302)  and  (not A300) );
 a16987a <=( (not A269)  and  a16986a );
 a16988a <=( a16987a  and  a16982a );
 a16991a <=( (not A168)  and  A169 );
 a16995a <=( A201  and  (not A200) );
 a16996a <=( A199  and  a16995a );
 a16997a <=( a16996a  and  a16991a );
 a17000a <=( (not A267)  and  A202 );
 a17004a <=( A299  and  A298 );
 a17005a <=( (not A269)  and  a17004a );
 a17006a <=( a17005a  and  a17000a );
 a17009a <=( (not A168)  and  A169 );
 a17013a <=( A201  and  (not A200) );
 a17014a <=( A199  and  a17013a );
 a17015a <=( a17014a  and  a17009a );
 a17018a <=( (not A267)  and  A202 );
 a17022a <=( (not A299)  and  (not A298) );
 a17023a <=( (not A269)  and  a17022a );
 a17024a <=( a17023a  and  a17018a );
 a17027a <=( (not A168)  and  A169 );
 a17031a <=( A201  and  (not A200) );
 a17032a <=( A199  and  a17031a );
 a17033a <=( a17032a  and  a17027a );
 a17036a <=( A265  and  A202 );
 a17040a <=( A301  and  (not A300) );
 a17041a <=( A266  and  a17040a );
 a17042a <=( a17041a  and  a17036a );
 a17045a <=( (not A168)  and  A169 );
 a17049a <=( A201  and  (not A200) );
 a17050a <=( A199  and  a17049a );
 a17051a <=( a17050a  and  a17045a );
 a17054a <=( A265  and  A202 );
 a17058a <=( (not A302)  and  (not A300) );
 a17059a <=( A266  and  a17058a );
 a17060a <=( a17059a  and  a17054a );
 a17063a <=( (not A168)  and  A169 );
 a17067a <=( A201  and  (not A200) );
 a17068a <=( A199  and  a17067a );
 a17069a <=( a17068a  and  a17063a );
 a17072a <=( A265  and  A202 );
 a17076a <=( A299  and  A298 );
 a17077a <=( A266  and  a17076a );
 a17078a <=( a17077a  and  a17072a );
 a17081a <=( (not A168)  and  A169 );
 a17085a <=( A201  and  (not A200) );
 a17086a <=( A199  and  a17085a );
 a17087a <=( a17086a  and  a17081a );
 a17090a <=( A265  and  A202 );
 a17094a <=( (not A299)  and  (not A298) );
 a17095a <=( A266  and  a17094a );
 a17096a <=( a17095a  and  a17090a );
 a17099a <=( (not A168)  and  A169 );
 a17103a <=( A201  and  (not A200) );
 a17104a <=( A199  and  a17103a );
 a17105a <=( a17104a  and  a17099a );
 a17108a <=( (not A265)  and  A202 );
 a17112a <=( A301  and  (not A300) );
 a17113a <=( (not A266)  and  a17112a );
 a17114a <=( a17113a  and  a17108a );
 a17117a <=( (not A168)  and  A169 );
 a17121a <=( A201  and  (not A200) );
 a17122a <=( A199  and  a17121a );
 a17123a <=( a17122a  and  a17117a );
 a17126a <=( (not A265)  and  A202 );
 a17130a <=( (not A302)  and  (not A300) );
 a17131a <=( (not A266)  and  a17130a );
 a17132a <=( a17131a  and  a17126a );
 a17135a <=( (not A168)  and  A169 );
 a17139a <=( A201  and  (not A200) );
 a17140a <=( A199  and  a17139a );
 a17141a <=( a17140a  and  a17135a );
 a17144a <=( (not A265)  and  A202 );
 a17148a <=( A299  and  A298 );
 a17149a <=( (not A266)  and  a17148a );
 a17150a <=( a17149a  and  a17144a );
 a17153a <=( (not A168)  and  A169 );
 a17157a <=( A201  and  (not A200) );
 a17158a <=( A199  and  a17157a );
 a17159a <=( a17158a  and  a17153a );
 a17162a <=( (not A265)  and  A202 );
 a17166a <=( (not A299)  and  (not A298) );
 a17167a <=( (not A266)  and  a17166a );
 a17168a <=( a17167a  and  a17162a );
 a17171a <=( (not A168)  and  A169 );
 a17175a <=( A201  and  (not A200) );
 a17176a <=( A199  and  a17175a );
 a17177a <=( a17176a  and  a17171a );
 a17180a <=( (not A267)  and  (not A203) );
 a17184a <=( A301  and  (not A300) );
 a17185a <=( A268  and  a17184a );
 a17186a <=( a17185a  and  a17180a );
 a17189a <=( (not A168)  and  A169 );
 a17193a <=( A201  and  (not A200) );
 a17194a <=( A199  and  a17193a );
 a17195a <=( a17194a  and  a17189a );
 a17198a <=( (not A267)  and  (not A203) );
 a17202a <=( (not A302)  and  (not A300) );
 a17203a <=( A268  and  a17202a );
 a17204a <=( a17203a  and  a17198a );
 a17207a <=( (not A168)  and  A169 );
 a17211a <=( A201  and  (not A200) );
 a17212a <=( A199  and  a17211a );
 a17213a <=( a17212a  and  a17207a );
 a17216a <=( (not A267)  and  (not A203) );
 a17220a <=( A299  and  A298 );
 a17221a <=( A268  and  a17220a );
 a17222a <=( a17221a  and  a17216a );
 a17225a <=( (not A168)  and  A169 );
 a17229a <=( A201  and  (not A200) );
 a17230a <=( A199  and  a17229a );
 a17231a <=( a17230a  and  a17225a );
 a17234a <=( (not A267)  and  (not A203) );
 a17238a <=( (not A299)  and  (not A298) );
 a17239a <=( A268  and  a17238a );
 a17240a <=( a17239a  and  a17234a );
 a17243a <=( (not A168)  and  A169 );
 a17247a <=( A201  and  (not A200) );
 a17248a <=( A199  and  a17247a );
 a17249a <=( a17248a  and  a17243a );
 a17252a <=( (not A267)  and  (not A203) );
 a17256a <=( A301  and  (not A300) );
 a17257a <=( (not A269)  and  a17256a );
 a17258a <=( a17257a  and  a17252a );
 a17261a <=( (not A168)  and  A169 );
 a17265a <=( A201  and  (not A200) );
 a17266a <=( A199  and  a17265a );
 a17267a <=( a17266a  and  a17261a );
 a17270a <=( (not A267)  and  (not A203) );
 a17274a <=( (not A302)  and  (not A300) );
 a17275a <=( (not A269)  and  a17274a );
 a17276a <=( a17275a  and  a17270a );
 a17279a <=( (not A168)  and  A169 );
 a17283a <=( A201  and  (not A200) );
 a17284a <=( A199  and  a17283a );
 a17285a <=( a17284a  and  a17279a );
 a17288a <=( (not A267)  and  (not A203) );
 a17292a <=( A299  and  A298 );
 a17293a <=( (not A269)  and  a17292a );
 a17294a <=( a17293a  and  a17288a );
 a17297a <=( (not A168)  and  A169 );
 a17301a <=( A201  and  (not A200) );
 a17302a <=( A199  and  a17301a );
 a17303a <=( a17302a  and  a17297a );
 a17306a <=( (not A267)  and  (not A203) );
 a17310a <=( (not A299)  and  (not A298) );
 a17311a <=( (not A269)  and  a17310a );
 a17312a <=( a17311a  and  a17306a );
 a17315a <=( (not A168)  and  A169 );
 a17319a <=( A201  and  (not A200) );
 a17320a <=( A199  and  a17319a );
 a17321a <=( a17320a  and  a17315a );
 a17324a <=( A265  and  (not A203) );
 a17328a <=( A301  and  (not A300) );
 a17329a <=( A266  and  a17328a );
 a17330a <=( a17329a  and  a17324a );
 a17333a <=( (not A168)  and  A169 );
 a17337a <=( A201  and  (not A200) );
 a17338a <=( A199  and  a17337a );
 a17339a <=( a17338a  and  a17333a );
 a17342a <=( A265  and  (not A203) );
 a17346a <=( (not A302)  and  (not A300) );
 a17347a <=( A266  and  a17346a );
 a17348a <=( a17347a  and  a17342a );
 a17351a <=( (not A168)  and  A169 );
 a17355a <=( A201  and  (not A200) );
 a17356a <=( A199  and  a17355a );
 a17357a <=( a17356a  and  a17351a );
 a17360a <=( A265  and  (not A203) );
 a17364a <=( A299  and  A298 );
 a17365a <=( A266  and  a17364a );
 a17366a <=( a17365a  and  a17360a );
 a17369a <=( (not A168)  and  A169 );
 a17373a <=( A201  and  (not A200) );
 a17374a <=( A199  and  a17373a );
 a17375a <=( a17374a  and  a17369a );
 a17378a <=( A265  and  (not A203) );
 a17382a <=( (not A299)  and  (not A298) );
 a17383a <=( A266  and  a17382a );
 a17384a <=( a17383a  and  a17378a );
 a17387a <=( (not A168)  and  A169 );
 a17391a <=( A201  and  (not A200) );
 a17392a <=( A199  and  a17391a );
 a17393a <=( a17392a  and  a17387a );
 a17396a <=( (not A265)  and  (not A203) );
 a17400a <=( A301  and  (not A300) );
 a17401a <=( (not A266)  and  a17400a );
 a17402a <=( a17401a  and  a17396a );
 a17405a <=( (not A168)  and  A169 );
 a17409a <=( A201  and  (not A200) );
 a17410a <=( A199  and  a17409a );
 a17411a <=( a17410a  and  a17405a );
 a17414a <=( (not A265)  and  (not A203) );
 a17418a <=( (not A302)  and  (not A300) );
 a17419a <=( (not A266)  and  a17418a );
 a17420a <=( a17419a  and  a17414a );
 a17423a <=( (not A168)  and  A169 );
 a17427a <=( A201  and  (not A200) );
 a17428a <=( A199  and  a17427a );
 a17429a <=( a17428a  and  a17423a );
 a17432a <=( (not A265)  and  (not A203) );
 a17436a <=( A299  and  A298 );
 a17437a <=( (not A266)  and  a17436a );
 a17438a <=( a17437a  and  a17432a );
 a17441a <=( (not A168)  and  A169 );
 a17445a <=( A201  and  (not A200) );
 a17446a <=( A199  and  a17445a );
 a17447a <=( a17446a  and  a17441a );
 a17450a <=( (not A265)  and  (not A203) );
 a17454a <=( (not A299)  and  (not A298) );
 a17455a <=( (not A266)  and  a17454a );
 a17456a <=( a17455a  and  a17450a );
 a17459a <=( A233  and  (not A232) );
 a17463a <=( A236  and  (not A235) );
 a17464a <=( (not A234)  and  a17463a );
 a17465a <=( a17464a  and  a17459a );
 a17469a <=( (not A267)  and  A266 );
 a17470a <=( (not A265)  and  a17469a );
 a17474a <=( A300  and  A269 );
 a17475a <=( (not A268)  and  a17474a );
 a17476a <=( a17475a  and  a17470a );
 a17479a <=( A233  and  (not A232) );
 a17483a <=( A236  and  (not A235) );
 a17484a <=( (not A234)  and  a17483a );
 a17485a <=( a17484a  and  a17479a );
 a17489a <=( (not A267)  and  (not A266) );
 a17490a <=( A265  and  a17489a );
 a17494a <=( A300  and  A269 );
 a17495a <=( (not A268)  and  a17494a );
 a17496a <=( a17495a  and  a17490a );
 a17499a <=( (not A233)  and  A232 );
 a17503a <=( A236  and  (not A235) );
 a17504a <=( (not A234)  and  a17503a );
 a17505a <=( a17504a  and  a17499a );
 a17509a <=( (not A267)  and  A266 );
 a17510a <=( (not A265)  and  a17509a );
 a17514a <=( A300  and  A269 );
 a17515a <=( (not A268)  and  a17514a );
 a17516a <=( a17515a  and  a17510a );
 a17519a <=( (not A233)  and  A232 );
 a17523a <=( A236  and  (not A235) );
 a17524a <=( (not A234)  and  a17523a );
 a17525a <=( a17524a  and  a17519a );
 a17529a <=( (not A267)  and  (not A266) );
 a17530a <=( A265  and  a17529a );
 a17534a <=( A300  and  A269 );
 a17535a <=( (not A268)  and  a17534a );
 a17536a <=( a17535a  and  a17530a );
 a17539a <=( (not A232)  and  (not A201) );
 a17543a <=( (not A235)  and  (not A234) );
 a17544a <=( A233  and  a17543a );
 a17545a <=( a17544a  and  a17539a );
 a17549a <=( A266  and  (not A265) );
 a17550a <=( A236  and  a17549a );
 a17554a <=( A269  and  (not A268) );
 a17555a <=( (not A267)  and  a17554a );
 a17556a <=( a17555a  and  a17550a );
 a17559a <=( (not A232)  and  (not A201) );
 a17563a <=( (not A235)  and  (not A234) );
 a17564a <=( A233  and  a17563a );
 a17565a <=( a17564a  and  a17559a );
 a17569a <=( (not A266)  and  A265 );
 a17570a <=( A236  and  a17569a );
 a17574a <=( A269  and  (not A268) );
 a17575a <=( (not A267)  and  a17574a );
 a17576a <=( a17575a  and  a17570a );
 a17579a <=( A232  and  (not A201) );
 a17583a <=( (not A235)  and  (not A234) );
 a17584a <=( (not A233)  and  a17583a );
 a17585a <=( a17584a  and  a17579a );
 a17589a <=( A266  and  (not A265) );
 a17590a <=( A236  and  a17589a );
 a17594a <=( A269  and  (not A268) );
 a17595a <=( (not A267)  and  a17594a );
 a17596a <=( a17595a  and  a17590a );
 a17599a <=( A232  and  (not A201) );
 a17603a <=( (not A235)  and  (not A234) );
 a17604a <=( (not A233)  and  a17603a );
 a17605a <=( a17604a  and  a17599a );
 a17609a <=( (not A266)  and  A265 );
 a17610a <=( A236  and  a17609a );
 a17614a <=( A269  and  (not A268) );
 a17615a <=( (not A267)  and  a17614a );
 a17616a <=( a17615a  and  a17610a );
 a17619a <=( A166  and  A167 );
 a17623a <=( A234  and  A233 );
 a17624a <=( (not A232)  and  a17623a );
 a17625a <=( a17624a  and  a17619a );
 a17629a <=( A266  and  (not A265) );
 a17630a <=( A235  and  a17629a );
 a17634a <=( A269  and  (not A268) );
 a17635a <=( (not A267)  and  a17634a );
 a17636a <=( a17635a  and  a17630a );
 a17639a <=( A166  and  A167 );
 a17643a <=( A234  and  A233 );
 a17644a <=( (not A232)  and  a17643a );
 a17645a <=( a17644a  and  a17639a );
 a17649a <=( (not A266)  and  A265 );
 a17650a <=( A235  and  a17649a );
 a17654a <=( A269  and  (not A268) );
 a17655a <=( (not A267)  and  a17654a );
 a17656a <=( a17655a  and  a17650a );
 a17659a <=( A166  and  A167 );
 a17663a <=( A234  and  A233 );
 a17664a <=( (not A232)  and  a17663a );
 a17665a <=( a17664a  and  a17659a );
 a17669a <=( A266  and  (not A265) );
 a17670a <=( (not A236)  and  a17669a );
 a17674a <=( A269  and  (not A268) );
 a17675a <=( (not A267)  and  a17674a );
 a17676a <=( a17675a  and  a17670a );
 a17679a <=( A166  and  A167 );
 a17683a <=( A234  and  A233 );
 a17684a <=( (not A232)  and  a17683a );
 a17685a <=( a17684a  and  a17679a );
 a17689a <=( (not A266)  and  A265 );
 a17690a <=( (not A236)  and  a17689a );
 a17694a <=( A269  and  (not A268) );
 a17695a <=( (not A267)  and  a17694a );
 a17696a <=( a17695a  and  a17690a );
 a17699a <=( A166  and  A167 );
 a17703a <=( A234  and  (not A233) );
 a17704a <=( A232  and  a17703a );
 a17705a <=( a17704a  and  a17699a );
 a17709a <=( A266  and  (not A265) );
 a17710a <=( A235  and  a17709a );
 a17714a <=( A269  and  (not A268) );
 a17715a <=( (not A267)  and  a17714a );
 a17716a <=( a17715a  and  a17710a );
 a17719a <=( A166  and  A167 );
 a17723a <=( A234  and  (not A233) );
 a17724a <=( A232  and  a17723a );
 a17725a <=( a17724a  and  a17719a );
 a17729a <=( (not A266)  and  A265 );
 a17730a <=( A235  and  a17729a );
 a17734a <=( A269  and  (not A268) );
 a17735a <=( (not A267)  and  a17734a );
 a17736a <=( a17735a  and  a17730a );
 a17739a <=( A166  and  A167 );
 a17743a <=( A234  and  (not A233) );
 a17744a <=( A232  and  a17743a );
 a17745a <=( a17744a  and  a17739a );
 a17749a <=( A266  and  (not A265) );
 a17750a <=( (not A236)  and  a17749a );
 a17754a <=( A269  and  (not A268) );
 a17755a <=( (not A267)  and  a17754a );
 a17756a <=( a17755a  and  a17750a );
 a17759a <=( A166  and  A167 );
 a17763a <=( A234  and  (not A233) );
 a17764a <=( A232  and  a17763a );
 a17765a <=( a17764a  and  a17759a );
 a17769a <=( (not A266)  and  A265 );
 a17770a <=( (not A236)  and  a17769a );
 a17774a <=( A269  and  (not A268) );
 a17775a <=( (not A267)  and  a17774a );
 a17776a <=( a17775a  and  a17770a );
 a17779a <=( A166  and  A167 );
 a17783a <=( A201  and  A200 );
 a17784a <=( (not A199)  and  a17783a );
 a17785a <=( a17784a  and  a17779a );
 a17789a <=( (not A268)  and  A267 );
 a17790a <=( A202  and  a17789a );
 a17794a <=( A301  and  (not A300) );
 a17795a <=( A269  and  a17794a );
 a17796a <=( a17795a  and  a17790a );
 a17799a <=( A166  and  A167 );
 a17803a <=( A201  and  A200 );
 a17804a <=( (not A199)  and  a17803a );
 a17805a <=( a17804a  and  a17799a );
 a17809a <=( (not A268)  and  A267 );
 a17810a <=( A202  and  a17809a );
 a17814a <=( (not A302)  and  (not A300) );
 a17815a <=( A269  and  a17814a );
 a17816a <=( a17815a  and  a17810a );
 a17819a <=( A166  and  A167 );
 a17823a <=( A201  and  A200 );
 a17824a <=( (not A199)  and  a17823a );
 a17825a <=( a17824a  and  a17819a );
 a17829a <=( (not A268)  and  A267 );
 a17830a <=( A202  and  a17829a );
 a17834a <=( A299  and  A298 );
 a17835a <=( A269  and  a17834a );
 a17836a <=( a17835a  and  a17830a );
 a17839a <=( A166  and  A167 );
 a17843a <=( A201  and  A200 );
 a17844a <=( (not A199)  and  a17843a );
 a17845a <=( a17844a  and  a17839a );
 a17849a <=( (not A268)  and  A267 );
 a17850a <=( A202  and  a17849a );
 a17854a <=( (not A299)  and  (not A298) );
 a17855a <=( A269  and  a17854a );
 a17856a <=( a17855a  and  a17850a );
 a17859a <=( A166  and  A167 );
 a17863a <=( A201  and  A200 );
 a17864a <=( (not A199)  and  a17863a );
 a17865a <=( a17864a  and  a17859a );
 a17869a <=( A268  and  (not A267) );
 a17870a <=( A202  and  a17869a );
 a17874a <=( A302  and  (not A301) );
 a17875a <=( A300  and  a17874a );
 a17876a <=( a17875a  and  a17870a );
 a17879a <=( A166  and  A167 );
 a17883a <=( A201  and  A200 );
 a17884a <=( (not A199)  and  a17883a );
 a17885a <=( a17884a  and  a17879a );
 a17889a <=( (not A269)  and  (not A267) );
 a17890a <=( A202  and  a17889a );
 a17894a <=( A302  and  (not A301) );
 a17895a <=( A300  and  a17894a );
 a17896a <=( a17895a  and  a17890a );
 a17899a <=( A166  and  A167 );
 a17903a <=( A201  and  A200 );
 a17904a <=( (not A199)  and  a17903a );
 a17905a <=( a17904a  and  a17899a );
 a17909a <=( A266  and  A265 );
 a17910a <=( A202  and  a17909a );
 a17914a <=( A302  and  (not A301) );
 a17915a <=( A300  and  a17914a );
 a17916a <=( a17915a  and  a17910a );
 a17919a <=( A166  and  A167 );
 a17923a <=( A201  and  A200 );
 a17924a <=( (not A199)  and  a17923a );
 a17925a <=( a17924a  and  a17919a );
 a17929a <=( (not A266)  and  (not A265) );
 a17930a <=( A202  and  a17929a );
 a17934a <=( A302  and  (not A301) );
 a17935a <=( A300  and  a17934a );
 a17936a <=( a17935a  and  a17930a );
 a17939a <=( A166  and  A167 );
 a17943a <=( A201  and  A200 );
 a17944a <=( (not A199)  and  a17943a );
 a17945a <=( a17944a  and  a17939a );
 a17949a <=( (not A268)  and  A267 );
 a17950a <=( (not A203)  and  a17949a );
 a17954a <=( A301  and  (not A300) );
 a17955a <=( A269  and  a17954a );
 a17956a <=( a17955a  and  a17950a );
 a17959a <=( A166  and  A167 );
 a17963a <=( A201  and  A200 );
 a17964a <=( (not A199)  and  a17963a );
 a17965a <=( a17964a  and  a17959a );
 a17969a <=( (not A268)  and  A267 );
 a17970a <=( (not A203)  and  a17969a );
 a17974a <=( (not A302)  and  (not A300) );
 a17975a <=( A269  and  a17974a );
 a17976a <=( a17975a  and  a17970a );
 a17979a <=( A166  and  A167 );
 a17983a <=( A201  and  A200 );
 a17984a <=( (not A199)  and  a17983a );
 a17985a <=( a17984a  and  a17979a );
 a17989a <=( (not A268)  and  A267 );
 a17990a <=( (not A203)  and  a17989a );
 a17994a <=( A299  and  A298 );
 a17995a <=( A269  and  a17994a );
 a17996a <=( a17995a  and  a17990a );
 a17999a <=( A166  and  A167 );
 a18003a <=( A201  and  A200 );
 a18004a <=( (not A199)  and  a18003a );
 a18005a <=( a18004a  and  a17999a );
 a18009a <=( (not A268)  and  A267 );
 a18010a <=( (not A203)  and  a18009a );
 a18014a <=( (not A299)  and  (not A298) );
 a18015a <=( A269  and  a18014a );
 a18016a <=( a18015a  and  a18010a );
 a18019a <=( A166  and  A167 );
 a18023a <=( A201  and  A200 );
 a18024a <=( (not A199)  and  a18023a );
 a18025a <=( a18024a  and  a18019a );
 a18029a <=( A268  and  (not A267) );
 a18030a <=( (not A203)  and  a18029a );
 a18034a <=( A302  and  (not A301) );
 a18035a <=( A300  and  a18034a );
 a18036a <=( a18035a  and  a18030a );
 a18039a <=( A166  and  A167 );
 a18043a <=( A201  and  A200 );
 a18044a <=( (not A199)  and  a18043a );
 a18045a <=( a18044a  and  a18039a );
 a18049a <=( (not A269)  and  (not A267) );
 a18050a <=( (not A203)  and  a18049a );
 a18054a <=( A302  and  (not A301) );
 a18055a <=( A300  and  a18054a );
 a18056a <=( a18055a  and  a18050a );
 a18059a <=( A166  and  A167 );
 a18063a <=( A201  and  A200 );
 a18064a <=( (not A199)  and  a18063a );
 a18065a <=( a18064a  and  a18059a );
 a18069a <=( A266  and  A265 );
 a18070a <=( (not A203)  and  a18069a );
 a18074a <=( A302  and  (not A301) );
 a18075a <=( A300  and  a18074a );
 a18076a <=( a18075a  and  a18070a );
 a18079a <=( A166  and  A167 );
 a18083a <=( A201  and  A200 );
 a18084a <=( (not A199)  and  a18083a );
 a18085a <=( a18084a  and  a18079a );
 a18089a <=( (not A266)  and  (not A265) );
 a18090a <=( (not A203)  and  a18089a );
 a18094a <=( A302  and  (not A301) );
 a18095a <=( A300  and  a18094a );
 a18096a <=( a18095a  and  a18090a );
 a18099a <=( A166  and  A167 );
 a18103a <=( (not A201)  and  A200 );
 a18104a <=( (not A199)  and  a18103a );
 a18105a <=( a18104a  and  a18099a );
 a18109a <=( (not A267)  and  A203 );
 a18110a <=( (not A202)  and  a18109a );
 a18114a <=( A301  and  (not A300) );
 a18115a <=( A268  and  a18114a );
 a18116a <=( a18115a  and  a18110a );
 a18119a <=( A166  and  A167 );
 a18123a <=( (not A201)  and  A200 );
 a18124a <=( (not A199)  and  a18123a );
 a18125a <=( a18124a  and  a18119a );
 a18129a <=( (not A267)  and  A203 );
 a18130a <=( (not A202)  and  a18129a );
 a18134a <=( (not A302)  and  (not A300) );
 a18135a <=( A268  and  a18134a );
 a18136a <=( a18135a  and  a18130a );
 a18139a <=( A166  and  A167 );
 a18143a <=( (not A201)  and  A200 );
 a18144a <=( (not A199)  and  a18143a );
 a18145a <=( a18144a  and  a18139a );
 a18149a <=( (not A267)  and  A203 );
 a18150a <=( (not A202)  and  a18149a );
 a18154a <=( A299  and  A298 );
 a18155a <=( A268  and  a18154a );
 a18156a <=( a18155a  and  a18150a );
 a18159a <=( A166  and  A167 );
 a18163a <=( (not A201)  and  A200 );
 a18164a <=( (not A199)  and  a18163a );
 a18165a <=( a18164a  and  a18159a );
 a18169a <=( (not A267)  and  A203 );
 a18170a <=( (not A202)  and  a18169a );
 a18174a <=( (not A299)  and  (not A298) );
 a18175a <=( A268  and  a18174a );
 a18176a <=( a18175a  and  a18170a );
 a18179a <=( A166  and  A167 );
 a18183a <=( (not A201)  and  A200 );
 a18184a <=( (not A199)  and  a18183a );
 a18185a <=( a18184a  and  a18179a );
 a18189a <=( (not A267)  and  A203 );
 a18190a <=( (not A202)  and  a18189a );
 a18194a <=( A301  and  (not A300) );
 a18195a <=( (not A269)  and  a18194a );
 a18196a <=( a18195a  and  a18190a );
 a18199a <=( A166  and  A167 );
 a18203a <=( (not A201)  and  A200 );
 a18204a <=( (not A199)  and  a18203a );
 a18205a <=( a18204a  and  a18199a );
 a18209a <=( (not A267)  and  A203 );
 a18210a <=( (not A202)  and  a18209a );
 a18214a <=( (not A302)  and  (not A300) );
 a18215a <=( (not A269)  and  a18214a );
 a18216a <=( a18215a  and  a18210a );
 a18219a <=( A166  and  A167 );
 a18223a <=( (not A201)  and  A200 );
 a18224a <=( (not A199)  and  a18223a );
 a18225a <=( a18224a  and  a18219a );
 a18229a <=( (not A267)  and  A203 );
 a18230a <=( (not A202)  and  a18229a );
 a18234a <=( A299  and  A298 );
 a18235a <=( (not A269)  and  a18234a );
 a18236a <=( a18235a  and  a18230a );
 a18239a <=( A166  and  A167 );
 a18243a <=( (not A201)  and  A200 );
 a18244a <=( (not A199)  and  a18243a );
 a18245a <=( a18244a  and  a18239a );
 a18249a <=( (not A267)  and  A203 );
 a18250a <=( (not A202)  and  a18249a );
 a18254a <=( (not A299)  and  (not A298) );
 a18255a <=( (not A269)  and  a18254a );
 a18256a <=( a18255a  and  a18250a );
 a18259a <=( A166  and  A167 );
 a18263a <=( (not A201)  and  A200 );
 a18264a <=( (not A199)  and  a18263a );
 a18265a <=( a18264a  and  a18259a );
 a18269a <=( A265  and  A203 );
 a18270a <=( (not A202)  and  a18269a );
 a18274a <=( A301  and  (not A300) );
 a18275a <=( A266  and  a18274a );
 a18276a <=( a18275a  and  a18270a );
 a18279a <=( A166  and  A167 );
 a18283a <=( (not A201)  and  A200 );
 a18284a <=( (not A199)  and  a18283a );
 a18285a <=( a18284a  and  a18279a );
 a18289a <=( A265  and  A203 );
 a18290a <=( (not A202)  and  a18289a );
 a18294a <=( (not A302)  and  (not A300) );
 a18295a <=( A266  and  a18294a );
 a18296a <=( a18295a  and  a18290a );
 a18299a <=( A166  and  A167 );
 a18303a <=( (not A201)  and  A200 );
 a18304a <=( (not A199)  and  a18303a );
 a18305a <=( a18304a  and  a18299a );
 a18309a <=( A265  and  A203 );
 a18310a <=( (not A202)  and  a18309a );
 a18314a <=( A299  and  A298 );
 a18315a <=( A266  and  a18314a );
 a18316a <=( a18315a  and  a18310a );
 a18319a <=( A166  and  A167 );
 a18323a <=( (not A201)  and  A200 );
 a18324a <=( (not A199)  and  a18323a );
 a18325a <=( a18324a  and  a18319a );
 a18329a <=( A265  and  A203 );
 a18330a <=( (not A202)  and  a18329a );
 a18334a <=( (not A299)  and  (not A298) );
 a18335a <=( A266  and  a18334a );
 a18336a <=( a18335a  and  a18330a );
 a18339a <=( A166  and  A167 );
 a18343a <=( (not A201)  and  A200 );
 a18344a <=( (not A199)  and  a18343a );
 a18345a <=( a18344a  and  a18339a );
 a18349a <=( (not A265)  and  A203 );
 a18350a <=( (not A202)  and  a18349a );
 a18354a <=( A301  and  (not A300) );
 a18355a <=( (not A266)  and  a18354a );
 a18356a <=( a18355a  and  a18350a );
 a18359a <=( A166  and  A167 );
 a18363a <=( (not A201)  and  A200 );
 a18364a <=( (not A199)  and  a18363a );
 a18365a <=( a18364a  and  a18359a );
 a18369a <=( (not A265)  and  A203 );
 a18370a <=( (not A202)  and  a18369a );
 a18374a <=( (not A302)  and  (not A300) );
 a18375a <=( (not A266)  and  a18374a );
 a18376a <=( a18375a  and  a18370a );
 a18379a <=( A166  and  A167 );
 a18383a <=( (not A201)  and  A200 );
 a18384a <=( (not A199)  and  a18383a );
 a18385a <=( a18384a  and  a18379a );
 a18389a <=( (not A265)  and  A203 );
 a18390a <=( (not A202)  and  a18389a );
 a18394a <=( A299  and  A298 );
 a18395a <=( (not A266)  and  a18394a );
 a18396a <=( a18395a  and  a18390a );
 a18399a <=( A166  and  A167 );
 a18403a <=( (not A201)  and  A200 );
 a18404a <=( (not A199)  and  a18403a );
 a18405a <=( a18404a  and  a18399a );
 a18409a <=( (not A265)  and  A203 );
 a18410a <=( (not A202)  and  a18409a );
 a18414a <=( (not A299)  and  (not A298) );
 a18415a <=( (not A266)  and  a18414a );
 a18416a <=( a18415a  and  a18410a );
 a18419a <=( A166  and  A167 );
 a18423a <=( A201  and  (not A200) );
 a18424a <=( A199  and  a18423a );
 a18425a <=( a18424a  and  a18419a );
 a18429a <=( (not A268)  and  A267 );
 a18430a <=( A202  and  a18429a );
 a18434a <=( A301  and  (not A300) );
 a18435a <=( A269  and  a18434a );
 a18436a <=( a18435a  and  a18430a );
 a18439a <=( A166  and  A167 );
 a18443a <=( A201  and  (not A200) );
 a18444a <=( A199  and  a18443a );
 a18445a <=( a18444a  and  a18439a );
 a18449a <=( (not A268)  and  A267 );
 a18450a <=( A202  and  a18449a );
 a18454a <=( (not A302)  and  (not A300) );
 a18455a <=( A269  and  a18454a );
 a18456a <=( a18455a  and  a18450a );
 a18459a <=( A166  and  A167 );
 a18463a <=( A201  and  (not A200) );
 a18464a <=( A199  and  a18463a );
 a18465a <=( a18464a  and  a18459a );
 a18469a <=( (not A268)  and  A267 );
 a18470a <=( A202  and  a18469a );
 a18474a <=( A299  and  A298 );
 a18475a <=( A269  and  a18474a );
 a18476a <=( a18475a  and  a18470a );
 a18479a <=( A166  and  A167 );
 a18483a <=( A201  and  (not A200) );
 a18484a <=( A199  and  a18483a );
 a18485a <=( a18484a  and  a18479a );
 a18489a <=( (not A268)  and  A267 );
 a18490a <=( A202  and  a18489a );
 a18494a <=( (not A299)  and  (not A298) );
 a18495a <=( A269  and  a18494a );
 a18496a <=( a18495a  and  a18490a );
 a18499a <=( A166  and  A167 );
 a18503a <=( A201  and  (not A200) );
 a18504a <=( A199  and  a18503a );
 a18505a <=( a18504a  and  a18499a );
 a18509a <=( A268  and  (not A267) );
 a18510a <=( A202  and  a18509a );
 a18514a <=( A302  and  (not A301) );
 a18515a <=( A300  and  a18514a );
 a18516a <=( a18515a  and  a18510a );
 a18519a <=( A166  and  A167 );
 a18523a <=( A201  and  (not A200) );
 a18524a <=( A199  and  a18523a );
 a18525a <=( a18524a  and  a18519a );
 a18529a <=( (not A269)  and  (not A267) );
 a18530a <=( A202  and  a18529a );
 a18534a <=( A302  and  (not A301) );
 a18535a <=( A300  and  a18534a );
 a18536a <=( a18535a  and  a18530a );
 a18539a <=( A166  and  A167 );
 a18543a <=( A201  and  (not A200) );
 a18544a <=( A199  and  a18543a );
 a18545a <=( a18544a  and  a18539a );
 a18549a <=( A266  and  A265 );
 a18550a <=( A202  and  a18549a );
 a18554a <=( A302  and  (not A301) );
 a18555a <=( A300  and  a18554a );
 a18556a <=( a18555a  and  a18550a );
 a18559a <=( A166  and  A167 );
 a18563a <=( A201  and  (not A200) );
 a18564a <=( A199  and  a18563a );
 a18565a <=( a18564a  and  a18559a );
 a18569a <=( (not A266)  and  (not A265) );
 a18570a <=( A202  and  a18569a );
 a18574a <=( A302  and  (not A301) );
 a18575a <=( A300  and  a18574a );
 a18576a <=( a18575a  and  a18570a );
 a18579a <=( A166  and  A167 );
 a18583a <=( A201  and  (not A200) );
 a18584a <=( A199  and  a18583a );
 a18585a <=( a18584a  and  a18579a );
 a18589a <=( (not A268)  and  A267 );
 a18590a <=( (not A203)  and  a18589a );
 a18594a <=( A301  and  (not A300) );
 a18595a <=( A269  and  a18594a );
 a18596a <=( a18595a  and  a18590a );
 a18599a <=( A166  and  A167 );
 a18603a <=( A201  and  (not A200) );
 a18604a <=( A199  and  a18603a );
 a18605a <=( a18604a  and  a18599a );
 a18609a <=( (not A268)  and  A267 );
 a18610a <=( (not A203)  and  a18609a );
 a18614a <=( (not A302)  and  (not A300) );
 a18615a <=( A269  and  a18614a );
 a18616a <=( a18615a  and  a18610a );
 a18619a <=( A166  and  A167 );
 a18623a <=( A201  and  (not A200) );
 a18624a <=( A199  and  a18623a );
 a18625a <=( a18624a  and  a18619a );
 a18629a <=( (not A268)  and  A267 );
 a18630a <=( (not A203)  and  a18629a );
 a18634a <=( A299  and  A298 );
 a18635a <=( A269  and  a18634a );
 a18636a <=( a18635a  and  a18630a );
 a18639a <=( A166  and  A167 );
 a18643a <=( A201  and  (not A200) );
 a18644a <=( A199  and  a18643a );
 a18645a <=( a18644a  and  a18639a );
 a18649a <=( (not A268)  and  A267 );
 a18650a <=( (not A203)  and  a18649a );
 a18654a <=( (not A299)  and  (not A298) );
 a18655a <=( A269  and  a18654a );
 a18656a <=( a18655a  and  a18650a );
 a18659a <=( A166  and  A167 );
 a18663a <=( A201  and  (not A200) );
 a18664a <=( A199  and  a18663a );
 a18665a <=( a18664a  and  a18659a );
 a18669a <=( A268  and  (not A267) );
 a18670a <=( (not A203)  and  a18669a );
 a18674a <=( A302  and  (not A301) );
 a18675a <=( A300  and  a18674a );
 a18676a <=( a18675a  and  a18670a );
 a18679a <=( A166  and  A167 );
 a18683a <=( A201  and  (not A200) );
 a18684a <=( A199  and  a18683a );
 a18685a <=( a18684a  and  a18679a );
 a18689a <=( (not A269)  and  (not A267) );
 a18690a <=( (not A203)  and  a18689a );
 a18694a <=( A302  and  (not A301) );
 a18695a <=( A300  and  a18694a );
 a18696a <=( a18695a  and  a18690a );
 a18699a <=( A166  and  A167 );
 a18703a <=( A201  and  (not A200) );
 a18704a <=( A199  and  a18703a );
 a18705a <=( a18704a  and  a18699a );
 a18709a <=( A266  and  A265 );
 a18710a <=( (not A203)  and  a18709a );
 a18714a <=( A302  and  (not A301) );
 a18715a <=( A300  and  a18714a );
 a18716a <=( a18715a  and  a18710a );
 a18719a <=( A166  and  A167 );
 a18723a <=( A201  and  (not A200) );
 a18724a <=( A199  and  a18723a );
 a18725a <=( a18724a  and  a18719a );
 a18729a <=( (not A266)  and  (not A265) );
 a18730a <=( (not A203)  and  a18729a );
 a18734a <=( A302  and  (not A301) );
 a18735a <=( A300  and  a18734a );
 a18736a <=( a18735a  and  a18730a );
 a18739a <=( A166  and  A167 );
 a18743a <=( (not A201)  and  (not A200) );
 a18744a <=( A199  and  a18743a );
 a18745a <=( a18744a  and  a18739a );
 a18749a <=( (not A267)  and  A203 );
 a18750a <=( (not A202)  and  a18749a );
 a18754a <=( A301  and  (not A300) );
 a18755a <=( A268  and  a18754a );
 a18756a <=( a18755a  and  a18750a );
 a18759a <=( A166  and  A167 );
 a18763a <=( (not A201)  and  (not A200) );
 a18764a <=( A199  and  a18763a );
 a18765a <=( a18764a  and  a18759a );
 a18769a <=( (not A267)  and  A203 );
 a18770a <=( (not A202)  and  a18769a );
 a18774a <=( (not A302)  and  (not A300) );
 a18775a <=( A268  and  a18774a );
 a18776a <=( a18775a  and  a18770a );
 a18779a <=( A166  and  A167 );
 a18783a <=( (not A201)  and  (not A200) );
 a18784a <=( A199  and  a18783a );
 a18785a <=( a18784a  and  a18779a );
 a18789a <=( (not A267)  and  A203 );
 a18790a <=( (not A202)  and  a18789a );
 a18794a <=( A299  and  A298 );
 a18795a <=( A268  and  a18794a );
 a18796a <=( a18795a  and  a18790a );
 a18799a <=( A166  and  A167 );
 a18803a <=( (not A201)  and  (not A200) );
 a18804a <=( A199  and  a18803a );
 a18805a <=( a18804a  and  a18799a );
 a18809a <=( (not A267)  and  A203 );
 a18810a <=( (not A202)  and  a18809a );
 a18814a <=( (not A299)  and  (not A298) );
 a18815a <=( A268  and  a18814a );
 a18816a <=( a18815a  and  a18810a );
 a18819a <=( A166  and  A167 );
 a18823a <=( (not A201)  and  (not A200) );
 a18824a <=( A199  and  a18823a );
 a18825a <=( a18824a  and  a18819a );
 a18829a <=( (not A267)  and  A203 );
 a18830a <=( (not A202)  and  a18829a );
 a18834a <=( A301  and  (not A300) );
 a18835a <=( (not A269)  and  a18834a );
 a18836a <=( a18835a  and  a18830a );
 a18839a <=( A166  and  A167 );
 a18843a <=( (not A201)  and  (not A200) );
 a18844a <=( A199  and  a18843a );
 a18845a <=( a18844a  and  a18839a );
 a18849a <=( (not A267)  and  A203 );
 a18850a <=( (not A202)  and  a18849a );
 a18854a <=( (not A302)  and  (not A300) );
 a18855a <=( (not A269)  and  a18854a );
 a18856a <=( a18855a  and  a18850a );
 a18859a <=( A166  and  A167 );
 a18863a <=( (not A201)  and  (not A200) );
 a18864a <=( A199  and  a18863a );
 a18865a <=( a18864a  and  a18859a );
 a18869a <=( (not A267)  and  A203 );
 a18870a <=( (not A202)  and  a18869a );
 a18874a <=( A299  and  A298 );
 a18875a <=( (not A269)  and  a18874a );
 a18876a <=( a18875a  and  a18870a );
 a18879a <=( A166  and  A167 );
 a18883a <=( (not A201)  and  (not A200) );
 a18884a <=( A199  and  a18883a );
 a18885a <=( a18884a  and  a18879a );
 a18889a <=( (not A267)  and  A203 );
 a18890a <=( (not A202)  and  a18889a );
 a18894a <=( (not A299)  and  (not A298) );
 a18895a <=( (not A269)  and  a18894a );
 a18896a <=( a18895a  and  a18890a );
 a18899a <=( A166  and  A167 );
 a18903a <=( (not A201)  and  (not A200) );
 a18904a <=( A199  and  a18903a );
 a18905a <=( a18904a  and  a18899a );
 a18909a <=( A265  and  A203 );
 a18910a <=( (not A202)  and  a18909a );
 a18914a <=( A301  and  (not A300) );
 a18915a <=( A266  and  a18914a );
 a18916a <=( a18915a  and  a18910a );
 a18919a <=( A166  and  A167 );
 a18923a <=( (not A201)  and  (not A200) );
 a18924a <=( A199  and  a18923a );
 a18925a <=( a18924a  and  a18919a );
 a18929a <=( A265  and  A203 );
 a18930a <=( (not A202)  and  a18929a );
 a18934a <=( (not A302)  and  (not A300) );
 a18935a <=( A266  and  a18934a );
 a18936a <=( a18935a  and  a18930a );
 a18939a <=( A166  and  A167 );
 a18943a <=( (not A201)  and  (not A200) );
 a18944a <=( A199  and  a18943a );
 a18945a <=( a18944a  and  a18939a );
 a18949a <=( A265  and  A203 );
 a18950a <=( (not A202)  and  a18949a );
 a18954a <=( A299  and  A298 );
 a18955a <=( A266  and  a18954a );
 a18956a <=( a18955a  and  a18950a );
 a18959a <=( A166  and  A167 );
 a18963a <=( (not A201)  and  (not A200) );
 a18964a <=( A199  and  a18963a );
 a18965a <=( a18964a  and  a18959a );
 a18969a <=( A265  and  A203 );
 a18970a <=( (not A202)  and  a18969a );
 a18974a <=( (not A299)  and  (not A298) );
 a18975a <=( A266  and  a18974a );
 a18976a <=( a18975a  and  a18970a );
 a18979a <=( A166  and  A167 );
 a18983a <=( (not A201)  and  (not A200) );
 a18984a <=( A199  and  a18983a );
 a18985a <=( a18984a  and  a18979a );
 a18989a <=( (not A265)  and  A203 );
 a18990a <=( (not A202)  and  a18989a );
 a18994a <=( A301  and  (not A300) );
 a18995a <=( (not A266)  and  a18994a );
 a18996a <=( a18995a  and  a18990a );
 a18999a <=( A166  and  A167 );
 a19003a <=( (not A201)  and  (not A200) );
 a19004a <=( A199  and  a19003a );
 a19005a <=( a19004a  and  a18999a );
 a19009a <=( (not A265)  and  A203 );
 a19010a <=( (not A202)  and  a19009a );
 a19014a <=( (not A302)  and  (not A300) );
 a19015a <=( (not A266)  and  a19014a );
 a19016a <=( a19015a  and  a19010a );
 a19019a <=( A166  and  A167 );
 a19023a <=( (not A201)  and  (not A200) );
 a19024a <=( A199  and  a19023a );
 a19025a <=( a19024a  and  a19019a );
 a19029a <=( (not A265)  and  A203 );
 a19030a <=( (not A202)  and  a19029a );
 a19034a <=( A299  and  A298 );
 a19035a <=( (not A266)  and  a19034a );
 a19036a <=( a19035a  and  a19030a );
 a19039a <=( A166  and  A167 );
 a19043a <=( (not A201)  and  (not A200) );
 a19044a <=( A199  and  a19043a );
 a19045a <=( a19044a  and  a19039a );
 a19049a <=( (not A265)  and  A203 );
 a19050a <=( (not A202)  and  a19049a );
 a19054a <=( (not A299)  and  (not A298) );
 a19055a <=( (not A266)  and  a19054a );
 a19056a <=( a19055a  and  a19050a );
 a19059a <=( (not A166)  and  (not A167) );
 a19063a <=( A234  and  A233 );
 a19064a <=( (not A232)  and  a19063a );
 a19065a <=( a19064a  and  a19059a );
 a19069a <=( A266  and  (not A265) );
 a19070a <=( A235  and  a19069a );
 a19074a <=( A269  and  (not A268) );
 a19075a <=( (not A267)  and  a19074a );
 a19076a <=( a19075a  and  a19070a );
 a19079a <=( (not A166)  and  (not A167) );
 a19083a <=( A234  and  A233 );
 a19084a <=( (not A232)  and  a19083a );
 a19085a <=( a19084a  and  a19079a );
 a19089a <=( (not A266)  and  A265 );
 a19090a <=( A235  and  a19089a );
 a19094a <=( A269  and  (not A268) );
 a19095a <=( (not A267)  and  a19094a );
 a19096a <=( a19095a  and  a19090a );
 a19099a <=( (not A166)  and  (not A167) );
 a19103a <=( A234  and  A233 );
 a19104a <=( (not A232)  and  a19103a );
 a19105a <=( a19104a  and  a19099a );
 a19109a <=( A266  and  (not A265) );
 a19110a <=( (not A236)  and  a19109a );
 a19114a <=( A269  and  (not A268) );
 a19115a <=( (not A267)  and  a19114a );
 a19116a <=( a19115a  and  a19110a );
 a19119a <=( (not A166)  and  (not A167) );
 a19123a <=( A234  and  A233 );
 a19124a <=( (not A232)  and  a19123a );
 a19125a <=( a19124a  and  a19119a );
 a19129a <=( (not A266)  and  A265 );
 a19130a <=( (not A236)  and  a19129a );
 a19134a <=( A269  and  (not A268) );
 a19135a <=( (not A267)  and  a19134a );
 a19136a <=( a19135a  and  a19130a );
 a19139a <=( (not A166)  and  (not A167) );
 a19143a <=( A234  and  (not A233) );
 a19144a <=( A232  and  a19143a );
 a19145a <=( a19144a  and  a19139a );
 a19149a <=( A266  and  (not A265) );
 a19150a <=( A235  and  a19149a );
 a19154a <=( A269  and  (not A268) );
 a19155a <=( (not A267)  and  a19154a );
 a19156a <=( a19155a  and  a19150a );
 a19159a <=( (not A166)  and  (not A167) );
 a19163a <=( A234  and  (not A233) );
 a19164a <=( A232  and  a19163a );
 a19165a <=( a19164a  and  a19159a );
 a19169a <=( (not A266)  and  A265 );
 a19170a <=( A235  and  a19169a );
 a19174a <=( A269  and  (not A268) );
 a19175a <=( (not A267)  and  a19174a );
 a19176a <=( a19175a  and  a19170a );
 a19179a <=( (not A166)  and  (not A167) );
 a19183a <=( A234  and  (not A233) );
 a19184a <=( A232  and  a19183a );
 a19185a <=( a19184a  and  a19179a );
 a19189a <=( A266  and  (not A265) );
 a19190a <=( (not A236)  and  a19189a );
 a19194a <=( A269  and  (not A268) );
 a19195a <=( (not A267)  and  a19194a );
 a19196a <=( a19195a  and  a19190a );
 a19199a <=( (not A166)  and  (not A167) );
 a19203a <=( A234  and  (not A233) );
 a19204a <=( A232  and  a19203a );
 a19205a <=( a19204a  and  a19199a );
 a19209a <=( (not A266)  and  A265 );
 a19210a <=( (not A236)  and  a19209a );
 a19214a <=( A269  and  (not A268) );
 a19215a <=( (not A267)  and  a19214a );
 a19216a <=( a19215a  and  a19210a );
 a19219a <=( (not A166)  and  (not A167) );
 a19223a <=( A201  and  A200 );
 a19224a <=( (not A199)  and  a19223a );
 a19225a <=( a19224a  and  a19219a );
 a19229a <=( (not A268)  and  A267 );
 a19230a <=( A202  and  a19229a );
 a19234a <=( A301  and  (not A300) );
 a19235a <=( A269  and  a19234a );
 a19236a <=( a19235a  and  a19230a );
 a19239a <=( (not A166)  and  (not A167) );
 a19243a <=( A201  and  A200 );
 a19244a <=( (not A199)  and  a19243a );
 a19245a <=( a19244a  and  a19239a );
 a19249a <=( (not A268)  and  A267 );
 a19250a <=( A202  and  a19249a );
 a19254a <=( (not A302)  and  (not A300) );
 a19255a <=( A269  and  a19254a );
 a19256a <=( a19255a  and  a19250a );
 a19259a <=( (not A166)  and  (not A167) );
 a19263a <=( A201  and  A200 );
 a19264a <=( (not A199)  and  a19263a );
 a19265a <=( a19264a  and  a19259a );
 a19269a <=( (not A268)  and  A267 );
 a19270a <=( A202  and  a19269a );
 a19274a <=( A299  and  A298 );
 a19275a <=( A269  and  a19274a );
 a19276a <=( a19275a  and  a19270a );
 a19279a <=( (not A166)  and  (not A167) );
 a19283a <=( A201  and  A200 );
 a19284a <=( (not A199)  and  a19283a );
 a19285a <=( a19284a  and  a19279a );
 a19289a <=( (not A268)  and  A267 );
 a19290a <=( A202  and  a19289a );
 a19294a <=( (not A299)  and  (not A298) );
 a19295a <=( A269  and  a19294a );
 a19296a <=( a19295a  and  a19290a );
 a19299a <=( (not A166)  and  (not A167) );
 a19303a <=( A201  and  A200 );
 a19304a <=( (not A199)  and  a19303a );
 a19305a <=( a19304a  and  a19299a );
 a19309a <=( A268  and  (not A267) );
 a19310a <=( A202  and  a19309a );
 a19314a <=( A302  and  (not A301) );
 a19315a <=( A300  and  a19314a );
 a19316a <=( a19315a  and  a19310a );
 a19319a <=( (not A166)  and  (not A167) );
 a19323a <=( A201  and  A200 );
 a19324a <=( (not A199)  and  a19323a );
 a19325a <=( a19324a  and  a19319a );
 a19329a <=( (not A269)  and  (not A267) );
 a19330a <=( A202  and  a19329a );
 a19334a <=( A302  and  (not A301) );
 a19335a <=( A300  and  a19334a );
 a19336a <=( a19335a  and  a19330a );
 a19339a <=( (not A166)  and  (not A167) );
 a19343a <=( A201  and  A200 );
 a19344a <=( (not A199)  and  a19343a );
 a19345a <=( a19344a  and  a19339a );
 a19349a <=( A266  and  A265 );
 a19350a <=( A202  and  a19349a );
 a19354a <=( A302  and  (not A301) );
 a19355a <=( A300  and  a19354a );
 a19356a <=( a19355a  and  a19350a );
 a19359a <=( (not A166)  and  (not A167) );
 a19363a <=( A201  and  A200 );
 a19364a <=( (not A199)  and  a19363a );
 a19365a <=( a19364a  and  a19359a );
 a19369a <=( (not A266)  and  (not A265) );
 a19370a <=( A202  and  a19369a );
 a19374a <=( A302  and  (not A301) );
 a19375a <=( A300  and  a19374a );
 a19376a <=( a19375a  and  a19370a );
 a19379a <=( (not A166)  and  (not A167) );
 a19383a <=( A201  and  A200 );
 a19384a <=( (not A199)  and  a19383a );
 a19385a <=( a19384a  and  a19379a );
 a19389a <=( (not A268)  and  A267 );
 a19390a <=( (not A203)  and  a19389a );
 a19394a <=( A301  and  (not A300) );
 a19395a <=( A269  and  a19394a );
 a19396a <=( a19395a  and  a19390a );
 a19399a <=( (not A166)  and  (not A167) );
 a19403a <=( A201  and  A200 );
 a19404a <=( (not A199)  and  a19403a );
 a19405a <=( a19404a  and  a19399a );
 a19409a <=( (not A268)  and  A267 );
 a19410a <=( (not A203)  and  a19409a );
 a19414a <=( (not A302)  and  (not A300) );
 a19415a <=( A269  and  a19414a );
 a19416a <=( a19415a  and  a19410a );
 a19419a <=( (not A166)  and  (not A167) );
 a19423a <=( A201  and  A200 );
 a19424a <=( (not A199)  and  a19423a );
 a19425a <=( a19424a  and  a19419a );
 a19429a <=( (not A268)  and  A267 );
 a19430a <=( (not A203)  and  a19429a );
 a19434a <=( A299  and  A298 );
 a19435a <=( A269  and  a19434a );
 a19436a <=( a19435a  and  a19430a );
 a19439a <=( (not A166)  and  (not A167) );
 a19443a <=( A201  and  A200 );
 a19444a <=( (not A199)  and  a19443a );
 a19445a <=( a19444a  and  a19439a );
 a19449a <=( (not A268)  and  A267 );
 a19450a <=( (not A203)  and  a19449a );
 a19454a <=( (not A299)  and  (not A298) );
 a19455a <=( A269  and  a19454a );
 a19456a <=( a19455a  and  a19450a );
 a19459a <=( (not A166)  and  (not A167) );
 a19463a <=( A201  and  A200 );
 a19464a <=( (not A199)  and  a19463a );
 a19465a <=( a19464a  and  a19459a );
 a19469a <=( A268  and  (not A267) );
 a19470a <=( (not A203)  and  a19469a );
 a19474a <=( A302  and  (not A301) );
 a19475a <=( A300  and  a19474a );
 a19476a <=( a19475a  and  a19470a );
 a19479a <=( (not A166)  and  (not A167) );
 a19483a <=( A201  and  A200 );
 a19484a <=( (not A199)  and  a19483a );
 a19485a <=( a19484a  and  a19479a );
 a19489a <=( (not A269)  and  (not A267) );
 a19490a <=( (not A203)  and  a19489a );
 a19494a <=( A302  and  (not A301) );
 a19495a <=( A300  and  a19494a );
 a19496a <=( a19495a  and  a19490a );
 a19499a <=( (not A166)  and  (not A167) );
 a19503a <=( A201  and  A200 );
 a19504a <=( (not A199)  and  a19503a );
 a19505a <=( a19504a  and  a19499a );
 a19509a <=( A266  and  A265 );
 a19510a <=( (not A203)  and  a19509a );
 a19514a <=( A302  and  (not A301) );
 a19515a <=( A300  and  a19514a );
 a19516a <=( a19515a  and  a19510a );
 a19519a <=( (not A166)  and  (not A167) );
 a19523a <=( A201  and  A200 );
 a19524a <=( (not A199)  and  a19523a );
 a19525a <=( a19524a  and  a19519a );
 a19529a <=( (not A266)  and  (not A265) );
 a19530a <=( (not A203)  and  a19529a );
 a19534a <=( A302  and  (not A301) );
 a19535a <=( A300  and  a19534a );
 a19536a <=( a19535a  and  a19530a );
 a19539a <=( (not A166)  and  (not A167) );
 a19543a <=( (not A201)  and  A200 );
 a19544a <=( (not A199)  and  a19543a );
 a19545a <=( a19544a  and  a19539a );
 a19549a <=( (not A267)  and  A203 );
 a19550a <=( (not A202)  and  a19549a );
 a19554a <=( A301  and  (not A300) );
 a19555a <=( A268  and  a19554a );
 a19556a <=( a19555a  and  a19550a );
 a19559a <=( (not A166)  and  (not A167) );
 a19563a <=( (not A201)  and  A200 );
 a19564a <=( (not A199)  and  a19563a );
 a19565a <=( a19564a  and  a19559a );
 a19569a <=( (not A267)  and  A203 );
 a19570a <=( (not A202)  and  a19569a );
 a19574a <=( (not A302)  and  (not A300) );
 a19575a <=( A268  and  a19574a );
 a19576a <=( a19575a  and  a19570a );
 a19579a <=( (not A166)  and  (not A167) );
 a19583a <=( (not A201)  and  A200 );
 a19584a <=( (not A199)  and  a19583a );
 a19585a <=( a19584a  and  a19579a );
 a19589a <=( (not A267)  and  A203 );
 a19590a <=( (not A202)  and  a19589a );
 a19594a <=( A299  and  A298 );
 a19595a <=( A268  and  a19594a );
 a19596a <=( a19595a  and  a19590a );
 a19599a <=( (not A166)  and  (not A167) );
 a19603a <=( (not A201)  and  A200 );
 a19604a <=( (not A199)  and  a19603a );
 a19605a <=( a19604a  and  a19599a );
 a19609a <=( (not A267)  and  A203 );
 a19610a <=( (not A202)  and  a19609a );
 a19614a <=( (not A299)  and  (not A298) );
 a19615a <=( A268  and  a19614a );
 a19616a <=( a19615a  and  a19610a );
 a19619a <=( (not A166)  and  (not A167) );
 a19623a <=( (not A201)  and  A200 );
 a19624a <=( (not A199)  and  a19623a );
 a19625a <=( a19624a  and  a19619a );
 a19629a <=( (not A267)  and  A203 );
 a19630a <=( (not A202)  and  a19629a );
 a19634a <=( A301  and  (not A300) );
 a19635a <=( (not A269)  and  a19634a );
 a19636a <=( a19635a  and  a19630a );
 a19639a <=( (not A166)  and  (not A167) );
 a19643a <=( (not A201)  and  A200 );
 a19644a <=( (not A199)  and  a19643a );
 a19645a <=( a19644a  and  a19639a );
 a19649a <=( (not A267)  and  A203 );
 a19650a <=( (not A202)  and  a19649a );
 a19654a <=( (not A302)  and  (not A300) );
 a19655a <=( (not A269)  and  a19654a );
 a19656a <=( a19655a  and  a19650a );
 a19659a <=( (not A166)  and  (not A167) );
 a19663a <=( (not A201)  and  A200 );
 a19664a <=( (not A199)  and  a19663a );
 a19665a <=( a19664a  and  a19659a );
 a19669a <=( (not A267)  and  A203 );
 a19670a <=( (not A202)  and  a19669a );
 a19674a <=( A299  and  A298 );
 a19675a <=( (not A269)  and  a19674a );
 a19676a <=( a19675a  and  a19670a );
 a19679a <=( (not A166)  and  (not A167) );
 a19683a <=( (not A201)  and  A200 );
 a19684a <=( (not A199)  and  a19683a );
 a19685a <=( a19684a  and  a19679a );
 a19689a <=( (not A267)  and  A203 );
 a19690a <=( (not A202)  and  a19689a );
 a19694a <=( (not A299)  and  (not A298) );
 a19695a <=( (not A269)  and  a19694a );
 a19696a <=( a19695a  and  a19690a );
 a19699a <=( (not A166)  and  (not A167) );
 a19703a <=( (not A201)  and  A200 );
 a19704a <=( (not A199)  and  a19703a );
 a19705a <=( a19704a  and  a19699a );
 a19709a <=( A265  and  A203 );
 a19710a <=( (not A202)  and  a19709a );
 a19714a <=( A301  and  (not A300) );
 a19715a <=( A266  and  a19714a );
 a19716a <=( a19715a  and  a19710a );
 a19719a <=( (not A166)  and  (not A167) );
 a19723a <=( (not A201)  and  A200 );
 a19724a <=( (not A199)  and  a19723a );
 a19725a <=( a19724a  and  a19719a );
 a19729a <=( A265  and  A203 );
 a19730a <=( (not A202)  and  a19729a );
 a19734a <=( (not A302)  and  (not A300) );
 a19735a <=( A266  and  a19734a );
 a19736a <=( a19735a  and  a19730a );
 a19739a <=( (not A166)  and  (not A167) );
 a19743a <=( (not A201)  and  A200 );
 a19744a <=( (not A199)  and  a19743a );
 a19745a <=( a19744a  and  a19739a );
 a19749a <=( A265  and  A203 );
 a19750a <=( (not A202)  and  a19749a );
 a19754a <=( A299  and  A298 );
 a19755a <=( A266  and  a19754a );
 a19756a <=( a19755a  and  a19750a );
 a19759a <=( (not A166)  and  (not A167) );
 a19763a <=( (not A201)  and  A200 );
 a19764a <=( (not A199)  and  a19763a );
 a19765a <=( a19764a  and  a19759a );
 a19769a <=( A265  and  A203 );
 a19770a <=( (not A202)  and  a19769a );
 a19774a <=( (not A299)  and  (not A298) );
 a19775a <=( A266  and  a19774a );
 a19776a <=( a19775a  and  a19770a );
 a19779a <=( (not A166)  and  (not A167) );
 a19783a <=( (not A201)  and  A200 );
 a19784a <=( (not A199)  and  a19783a );
 a19785a <=( a19784a  and  a19779a );
 a19789a <=( (not A265)  and  A203 );
 a19790a <=( (not A202)  and  a19789a );
 a19794a <=( A301  and  (not A300) );
 a19795a <=( (not A266)  and  a19794a );
 a19796a <=( a19795a  and  a19790a );
 a19799a <=( (not A166)  and  (not A167) );
 a19803a <=( (not A201)  and  A200 );
 a19804a <=( (not A199)  and  a19803a );
 a19805a <=( a19804a  and  a19799a );
 a19809a <=( (not A265)  and  A203 );
 a19810a <=( (not A202)  and  a19809a );
 a19814a <=( (not A302)  and  (not A300) );
 a19815a <=( (not A266)  and  a19814a );
 a19816a <=( a19815a  and  a19810a );
 a19819a <=( (not A166)  and  (not A167) );
 a19823a <=( (not A201)  and  A200 );
 a19824a <=( (not A199)  and  a19823a );
 a19825a <=( a19824a  and  a19819a );
 a19829a <=( (not A265)  and  A203 );
 a19830a <=( (not A202)  and  a19829a );
 a19834a <=( A299  and  A298 );
 a19835a <=( (not A266)  and  a19834a );
 a19836a <=( a19835a  and  a19830a );
 a19839a <=( (not A166)  and  (not A167) );
 a19843a <=( (not A201)  and  A200 );
 a19844a <=( (not A199)  and  a19843a );
 a19845a <=( a19844a  and  a19839a );
 a19849a <=( (not A265)  and  A203 );
 a19850a <=( (not A202)  and  a19849a );
 a19854a <=( (not A299)  and  (not A298) );
 a19855a <=( (not A266)  and  a19854a );
 a19856a <=( a19855a  and  a19850a );
 a19859a <=( (not A166)  and  (not A167) );
 a19863a <=( A201  and  (not A200) );
 a19864a <=( A199  and  a19863a );
 a19865a <=( a19864a  and  a19859a );
 a19869a <=( (not A268)  and  A267 );
 a19870a <=( A202  and  a19869a );
 a19874a <=( A301  and  (not A300) );
 a19875a <=( A269  and  a19874a );
 a19876a <=( a19875a  and  a19870a );
 a19879a <=( (not A166)  and  (not A167) );
 a19883a <=( A201  and  (not A200) );
 a19884a <=( A199  and  a19883a );
 a19885a <=( a19884a  and  a19879a );
 a19889a <=( (not A268)  and  A267 );
 a19890a <=( A202  and  a19889a );
 a19894a <=( (not A302)  and  (not A300) );
 a19895a <=( A269  and  a19894a );
 a19896a <=( a19895a  and  a19890a );
 a19899a <=( (not A166)  and  (not A167) );
 a19903a <=( A201  and  (not A200) );
 a19904a <=( A199  and  a19903a );
 a19905a <=( a19904a  and  a19899a );
 a19909a <=( (not A268)  and  A267 );
 a19910a <=( A202  and  a19909a );
 a19914a <=( A299  and  A298 );
 a19915a <=( A269  and  a19914a );
 a19916a <=( a19915a  and  a19910a );
 a19919a <=( (not A166)  and  (not A167) );
 a19923a <=( A201  and  (not A200) );
 a19924a <=( A199  and  a19923a );
 a19925a <=( a19924a  and  a19919a );
 a19929a <=( (not A268)  and  A267 );
 a19930a <=( A202  and  a19929a );
 a19934a <=( (not A299)  and  (not A298) );
 a19935a <=( A269  and  a19934a );
 a19936a <=( a19935a  and  a19930a );
 a19939a <=( (not A166)  and  (not A167) );
 a19943a <=( A201  and  (not A200) );
 a19944a <=( A199  and  a19943a );
 a19945a <=( a19944a  and  a19939a );
 a19949a <=( A268  and  (not A267) );
 a19950a <=( A202  and  a19949a );
 a19954a <=( A302  and  (not A301) );
 a19955a <=( A300  and  a19954a );
 a19956a <=( a19955a  and  a19950a );
 a19959a <=( (not A166)  and  (not A167) );
 a19963a <=( A201  and  (not A200) );
 a19964a <=( A199  and  a19963a );
 a19965a <=( a19964a  and  a19959a );
 a19969a <=( (not A269)  and  (not A267) );
 a19970a <=( A202  and  a19969a );
 a19974a <=( A302  and  (not A301) );
 a19975a <=( A300  and  a19974a );
 a19976a <=( a19975a  and  a19970a );
 a19979a <=( (not A166)  and  (not A167) );
 a19983a <=( A201  and  (not A200) );
 a19984a <=( A199  and  a19983a );
 a19985a <=( a19984a  and  a19979a );
 a19989a <=( A266  and  A265 );
 a19990a <=( A202  and  a19989a );
 a19994a <=( A302  and  (not A301) );
 a19995a <=( A300  and  a19994a );
 a19996a <=( a19995a  and  a19990a );
 a19999a <=( (not A166)  and  (not A167) );
 a20003a <=( A201  and  (not A200) );
 a20004a <=( A199  and  a20003a );
 a20005a <=( a20004a  and  a19999a );
 a20009a <=( (not A266)  and  (not A265) );
 a20010a <=( A202  and  a20009a );
 a20014a <=( A302  and  (not A301) );
 a20015a <=( A300  and  a20014a );
 a20016a <=( a20015a  and  a20010a );
 a20019a <=( (not A166)  and  (not A167) );
 a20023a <=( A201  and  (not A200) );
 a20024a <=( A199  and  a20023a );
 a20025a <=( a20024a  and  a20019a );
 a20029a <=( (not A268)  and  A267 );
 a20030a <=( (not A203)  and  a20029a );
 a20034a <=( A301  and  (not A300) );
 a20035a <=( A269  and  a20034a );
 a20036a <=( a20035a  and  a20030a );
 a20039a <=( (not A166)  and  (not A167) );
 a20043a <=( A201  and  (not A200) );
 a20044a <=( A199  and  a20043a );
 a20045a <=( a20044a  and  a20039a );
 a20049a <=( (not A268)  and  A267 );
 a20050a <=( (not A203)  and  a20049a );
 a20054a <=( (not A302)  and  (not A300) );
 a20055a <=( A269  and  a20054a );
 a20056a <=( a20055a  and  a20050a );
 a20059a <=( (not A166)  and  (not A167) );
 a20063a <=( A201  and  (not A200) );
 a20064a <=( A199  and  a20063a );
 a20065a <=( a20064a  and  a20059a );
 a20069a <=( (not A268)  and  A267 );
 a20070a <=( (not A203)  and  a20069a );
 a20074a <=( A299  and  A298 );
 a20075a <=( A269  and  a20074a );
 a20076a <=( a20075a  and  a20070a );
 a20079a <=( (not A166)  and  (not A167) );
 a20083a <=( A201  and  (not A200) );
 a20084a <=( A199  and  a20083a );
 a20085a <=( a20084a  and  a20079a );
 a20089a <=( (not A268)  and  A267 );
 a20090a <=( (not A203)  and  a20089a );
 a20094a <=( (not A299)  and  (not A298) );
 a20095a <=( A269  and  a20094a );
 a20096a <=( a20095a  and  a20090a );
 a20099a <=( (not A166)  and  (not A167) );
 a20103a <=( A201  and  (not A200) );
 a20104a <=( A199  and  a20103a );
 a20105a <=( a20104a  and  a20099a );
 a20109a <=( A268  and  (not A267) );
 a20110a <=( (not A203)  and  a20109a );
 a20114a <=( A302  and  (not A301) );
 a20115a <=( A300  and  a20114a );
 a20116a <=( a20115a  and  a20110a );
 a20119a <=( (not A166)  and  (not A167) );
 a20123a <=( A201  and  (not A200) );
 a20124a <=( A199  and  a20123a );
 a20125a <=( a20124a  and  a20119a );
 a20129a <=( (not A269)  and  (not A267) );
 a20130a <=( (not A203)  and  a20129a );
 a20134a <=( A302  and  (not A301) );
 a20135a <=( A300  and  a20134a );
 a20136a <=( a20135a  and  a20130a );
 a20139a <=( (not A166)  and  (not A167) );
 a20143a <=( A201  and  (not A200) );
 a20144a <=( A199  and  a20143a );
 a20145a <=( a20144a  and  a20139a );
 a20149a <=( A266  and  A265 );
 a20150a <=( (not A203)  and  a20149a );
 a20154a <=( A302  and  (not A301) );
 a20155a <=( A300  and  a20154a );
 a20156a <=( a20155a  and  a20150a );
 a20159a <=( (not A166)  and  (not A167) );
 a20163a <=( A201  and  (not A200) );
 a20164a <=( A199  and  a20163a );
 a20165a <=( a20164a  and  a20159a );
 a20169a <=( (not A266)  and  (not A265) );
 a20170a <=( (not A203)  and  a20169a );
 a20174a <=( A302  and  (not A301) );
 a20175a <=( A300  and  a20174a );
 a20176a <=( a20175a  and  a20170a );
 a20179a <=( (not A166)  and  (not A167) );
 a20183a <=( (not A201)  and  (not A200) );
 a20184a <=( A199  and  a20183a );
 a20185a <=( a20184a  and  a20179a );
 a20189a <=( (not A267)  and  A203 );
 a20190a <=( (not A202)  and  a20189a );
 a20194a <=( A301  and  (not A300) );
 a20195a <=( A268  and  a20194a );
 a20196a <=( a20195a  and  a20190a );
 a20199a <=( (not A166)  and  (not A167) );
 a20203a <=( (not A201)  and  (not A200) );
 a20204a <=( A199  and  a20203a );
 a20205a <=( a20204a  and  a20199a );
 a20209a <=( (not A267)  and  A203 );
 a20210a <=( (not A202)  and  a20209a );
 a20214a <=( (not A302)  and  (not A300) );
 a20215a <=( A268  and  a20214a );
 a20216a <=( a20215a  and  a20210a );
 a20219a <=( (not A166)  and  (not A167) );
 a20223a <=( (not A201)  and  (not A200) );
 a20224a <=( A199  and  a20223a );
 a20225a <=( a20224a  and  a20219a );
 a20229a <=( (not A267)  and  A203 );
 a20230a <=( (not A202)  and  a20229a );
 a20234a <=( A299  and  A298 );
 a20235a <=( A268  and  a20234a );
 a20236a <=( a20235a  and  a20230a );
 a20239a <=( (not A166)  and  (not A167) );
 a20243a <=( (not A201)  and  (not A200) );
 a20244a <=( A199  and  a20243a );
 a20245a <=( a20244a  and  a20239a );
 a20249a <=( (not A267)  and  A203 );
 a20250a <=( (not A202)  and  a20249a );
 a20254a <=( (not A299)  and  (not A298) );
 a20255a <=( A268  and  a20254a );
 a20256a <=( a20255a  and  a20250a );
 a20259a <=( (not A166)  and  (not A167) );
 a20263a <=( (not A201)  and  (not A200) );
 a20264a <=( A199  and  a20263a );
 a20265a <=( a20264a  and  a20259a );
 a20269a <=( (not A267)  and  A203 );
 a20270a <=( (not A202)  and  a20269a );
 a20274a <=( A301  and  (not A300) );
 a20275a <=( (not A269)  and  a20274a );
 a20276a <=( a20275a  and  a20270a );
 a20279a <=( (not A166)  and  (not A167) );
 a20283a <=( (not A201)  and  (not A200) );
 a20284a <=( A199  and  a20283a );
 a20285a <=( a20284a  and  a20279a );
 a20289a <=( (not A267)  and  A203 );
 a20290a <=( (not A202)  and  a20289a );
 a20294a <=( (not A302)  and  (not A300) );
 a20295a <=( (not A269)  and  a20294a );
 a20296a <=( a20295a  and  a20290a );
 a20299a <=( (not A166)  and  (not A167) );
 a20303a <=( (not A201)  and  (not A200) );
 a20304a <=( A199  and  a20303a );
 a20305a <=( a20304a  and  a20299a );
 a20309a <=( (not A267)  and  A203 );
 a20310a <=( (not A202)  and  a20309a );
 a20314a <=( A299  and  A298 );
 a20315a <=( (not A269)  and  a20314a );
 a20316a <=( a20315a  and  a20310a );
 a20319a <=( (not A166)  and  (not A167) );
 a20323a <=( (not A201)  and  (not A200) );
 a20324a <=( A199  and  a20323a );
 a20325a <=( a20324a  and  a20319a );
 a20329a <=( (not A267)  and  A203 );
 a20330a <=( (not A202)  and  a20329a );
 a20334a <=( (not A299)  and  (not A298) );
 a20335a <=( (not A269)  and  a20334a );
 a20336a <=( a20335a  and  a20330a );
 a20339a <=( (not A166)  and  (not A167) );
 a20343a <=( (not A201)  and  (not A200) );
 a20344a <=( A199  and  a20343a );
 a20345a <=( a20344a  and  a20339a );
 a20349a <=( A265  and  A203 );
 a20350a <=( (not A202)  and  a20349a );
 a20354a <=( A301  and  (not A300) );
 a20355a <=( A266  and  a20354a );
 a20356a <=( a20355a  and  a20350a );
 a20359a <=( (not A166)  and  (not A167) );
 a20363a <=( (not A201)  and  (not A200) );
 a20364a <=( A199  and  a20363a );
 a20365a <=( a20364a  and  a20359a );
 a20369a <=( A265  and  A203 );
 a20370a <=( (not A202)  and  a20369a );
 a20374a <=( (not A302)  and  (not A300) );
 a20375a <=( A266  and  a20374a );
 a20376a <=( a20375a  and  a20370a );
 a20379a <=( (not A166)  and  (not A167) );
 a20383a <=( (not A201)  and  (not A200) );
 a20384a <=( A199  and  a20383a );
 a20385a <=( a20384a  and  a20379a );
 a20389a <=( A265  and  A203 );
 a20390a <=( (not A202)  and  a20389a );
 a20394a <=( A299  and  A298 );
 a20395a <=( A266  and  a20394a );
 a20396a <=( a20395a  and  a20390a );
 a20399a <=( (not A166)  and  (not A167) );
 a20403a <=( (not A201)  and  (not A200) );
 a20404a <=( A199  and  a20403a );
 a20405a <=( a20404a  and  a20399a );
 a20409a <=( A265  and  A203 );
 a20410a <=( (not A202)  and  a20409a );
 a20414a <=( (not A299)  and  (not A298) );
 a20415a <=( A266  and  a20414a );
 a20416a <=( a20415a  and  a20410a );
 a20419a <=( (not A166)  and  (not A167) );
 a20423a <=( (not A201)  and  (not A200) );
 a20424a <=( A199  and  a20423a );
 a20425a <=( a20424a  and  a20419a );
 a20429a <=( (not A265)  and  A203 );
 a20430a <=( (not A202)  and  a20429a );
 a20434a <=( A301  and  (not A300) );
 a20435a <=( (not A266)  and  a20434a );
 a20436a <=( a20435a  and  a20430a );
 a20439a <=( (not A166)  and  (not A167) );
 a20443a <=( (not A201)  and  (not A200) );
 a20444a <=( A199  and  a20443a );
 a20445a <=( a20444a  and  a20439a );
 a20449a <=( (not A265)  and  A203 );
 a20450a <=( (not A202)  and  a20449a );
 a20454a <=( (not A302)  and  (not A300) );
 a20455a <=( (not A266)  and  a20454a );
 a20456a <=( a20455a  and  a20450a );
 a20459a <=( (not A166)  and  (not A167) );
 a20463a <=( (not A201)  and  (not A200) );
 a20464a <=( A199  and  a20463a );
 a20465a <=( a20464a  and  a20459a );
 a20469a <=( (not A265)  and  A203 );
 a20470a <=( (not A202)  and  a20469a );
 a20474a <=( A299  and  A298 );
 a20475a <=( (not A266)  and  a20474a );
 a20476a <=( a20475a  and  a20470a );
 a20479a <=( (not A166)  and  (not A167) );
 a20483a <=( (not A201)  and  (not A200) );
 a20484a <=( A199  and  a20483a );
 a20485a <=( a20484a  and  a20479a );
 a20489a <=( (not A265)  and  A203 );
 a20490a <=( (not A202)  and  a20489a );
 a20494a <=( (not A299)  and  (not A298) );
 a20495a <=( (not A266)  and  a20494a );
 a20496a <=( a20495a  and  a20490a );
 a20499a <=( (not A168)  and  A170 );
 a20503a <=( A201  and  A200 );
 a20504a <=( (not A199)  and  a20503a );
 a20505a <=( a20504a  and  a20499a );
 a20509a <=( (not A268)  and  A267 );
 a20510a <=( A202  and  a20509a );
 a20514a <=( A301  and  (not A300) );
 a20515a <=( A269  and  a20514a );
 a20516a <=( a20515a  and  a20510a );
 a20519a <=( (not A168)  and  A170 );
 a20523a <=( A201  and  A200 );
 a20524a <=( (not A199)  and  a20523a );
 a20525a <=( a20524a  and  a20519a );
 a20529a <=( (not A268)  and  A267 );
 a20530a <=( A202  and  a20529a );
 a20534a <=( (not A302)  and  (not A300) );
 a20535a <=( A269  and  a20534a );
 a20536a <=( a20535a  and  a20530a );
 a20539a <=( (not A168)  and  A170 );
 a20543a <=( A201  and  A200 );
 a20544a <=( (not A199)  and  a20543a );
 a20545a <=( a20544a  and  a20539a );
 a20549a <=( (not A268)  and  A267 );
 a20550a <=( A202  and  a20549a );
 a20554a <=( A299  and  A298 );
 a20555a <=( A269  and  a20554a );
 a20556a <=( a20555a  and  a20550a );
 a20559a <=( (not A168)  and  A170 );
 a20563a <=( A201  and  A200 );
 a20564a <=( (not A199)  and  a20563a );
 a20565a <=( a20564a  and  a20559a );
 a20569a <=( (not A268)  and  A267 );
 a20570a <=( A202  and  a20569a );
 a20574a <=( (not A299)  and  (not A298) );
 a20575a <=( A269  and  a20574a );
 a20576a <=( a20575a  and  a20570a );
 a20579a <=( (not A168)  and  A170 );
 a20583a <=( A201  and  A200 );
 a20584a <=( (not A199)  and  a20583a );
 a20585a <=( a20584a  and  a20579a );
 a20589a <=( A268  and  (not A267) );
 a20590a <=( A202  and  a20589a );
 a20594a <=( A302  and  (not A301) );
 a20595a <=( A300  and  a20594a );
 a20596a <=( a20595a  and  a20590a );
 a20599a <=( (not A168)  and  A170 );
 a20603a <=( A201  and  A200 );
 a20604a <=( (not A199)  and  a20603a );
 a20605a <=( a20604a  and  a20599a );
 a20609a <=( (not A269)  and  (not A267) );
 a20610a <=( A202  and  a20609a );
 a20614a <=( A302  and  (not A301) );
 a20615a <=( A300  and  a20614a );
 a20616a <=( a20615a  and  a20610a );
 a20619a <=( (not A168)  and  A170 );
 a20623a <=( A201  and  A200 );
 a20624a <=( (not A199)  and  a20623a );
 a20625a <=( a20624a  and  a20619a );
 a20629a <=( A266  and  A265 );
 a20630a <=( A202  and  a20629a );
 a20634a <=( A302  and  (not A301) );
 a20635a <=( A300  and  a20634a );
 a20636a <=( a20635a  and  a20630a );
 a20639a <=( (not A168)  and  A170 );
 a20643a <=( A201  and  A200 );
 a20644a <=( (not A199)  and  a20643a );
 a20645a <=( a20644a  and  a20639a );
 a20649a <=( (not A266)  and  (not A265) );
 a20650a <=( A202  and  a20649a );
 a20654a <=( A302  and  (not A301) );
 a20655a <=( A300  and  a20654a );
 a20656a <=( a20655a  and  a20650a );
 a20659a <=( (not A168)  and  A170 );
 a20663a <=( A201  and  A200 );
 a20664a <=( (not A199)  and  a20663a );
 a20665a <=( a20664a  and  a20659a );
 a20669a <=( (not A268)  and  A267 );
 a20670a <=( (not A203)  and  a20669a );
 a20674a <=( A301  and  (not A300) );
 a20675a <=( A269  and  a20674a );
 a20676a <=( a20675a  and  a20670a );
 a20679a <=( (not A168)  and  A170 );
 a20683a <=( A201  and  A200 );
 a20684a <=( (not A199)  and  a20683a );
 a20685a <=( a20684a  and  a20679a );
 a20689a <=( (not A268)  and  A267 );
 a20690a <=( (not A203)  and  a20689a );
 a20694a <=( (not A302)  and  (not A300) );
 a20695a <=( A269  and  a20694a );
 a20696a <=( a20695a  and  a20690a );
 a20699a <=( (not A168)  and  A170 );
 a20703a <=( A201  and  A200 );
 a20704a <=( (not A199)  and  a20703a );
 a20705a <=( a20704a  and  a20699a );
 a20709a <=( (not A268)  and  A267 );
 a20710a <=( (not A203)  and  a20709a );
 a20714a <=( A299  and  A298 );
 a20715a <=( A269  and  a20714a );
 a20716a <=( a20715a  and  a20710a );
 a20719a <=( (not A168)  and  A170 );
 a20723a <=( A201  and  A200 );
 a20724a <=( (not A199)  and  a20723a );
 a20725a <=( a20724a  and  a20719a );
 a20729a <=( (not A268)  and  A267 );
 a20730a <=( (not A203)  and  a20729a );
 a20734a <=( (not A299)  and  (not A298) );
 a20735a <=( A269  and  a20734a );
 a20736a <=( a20735a  and  a20730a );
 a20739a <=( (not A168)  and  A170 );
 a20743a <=( A201  and  A200 );
 a20744a <=( (not A199)  and  a20743a );
 a20745a <=( a20744a  and  a20739a );
 a20749a <=( A268  and  (not A267) );
 a20750a <=( (not A203)  and  a20749a );
 a20754a <=( A302  and  (not A301) );
 a20755a <=( A300  and  a20754a );
 a20756a <=( a20755a  and  a20750a );
 a20759a <=( (not A168)  and  A170 );
 a20763a <=( A201  and  A200 );
 a20764a <=( (not A199)  and  a20763a );
 a20765a <=( a20764a  and  a20759a );
 a20769a <=( (not A269)  and  (not A267) );
 a20770a <=( (not A203)  and  a20769a );
 a20774a <=( A302  and  (not A301) );
 a20775a <=( A300  and  a20774a );
 a20776a <=( a20775a  and  a20770a );
 a20779a <=( (not A168)  and  A170 );
 a20783a <=( A201  and  A200 );
 a20784a <=( (not A199)  and  a20783a );
 a20785a <=( a20784a  and  a20779a );
 a20789a <=( A266  and  A265 );
 a20790a <=( (not A203)  and  a20789a );
 a20794a <=( A302  and  (not A301) );
 a20795a <=( A300  and  a20794a );
 a20796a <=( a20795a  and  a20790a );
 a20799a <=( (not A168)  and  A170 );
 a20803a <=( A201  and  A200 );
 a20804a <=( (not A199)  and  a20803a );
 a20805a <=( a20804a  and  a20799a );
 a20809a <=( (not A266)  and  (not A265) );
 a20810a <=( (not A203)  and  a20809a );
 a20814a <=( A302  and  (not A301) );
 a20815a <=( A300  and  a20814a );
 a20816a <=( a20815a  and  a20810a );
 a20819a <=( (not A168)  and  A170 );
 a20823a <=( (not A201)  and  A200 );
 a20824a <=( (not A199)  and  a20823a );
 a20825a <=( a20824a  and  a20819a );
 a20829a <=( (not A267)  and  A203 );
 a20830a <=( (not A202)  and  a20829a );
 a20834a <=( A301  and  (not A300) );
 a20835a <=( A268  and  a20834a );
 a20836a <=( a20835a  and  a20830a );
 a20839a <=( (not A168)  and  A170 );
 a20843a <=( (not A201)  and  A200 );
 a20844a <=( (not A199)  and  a20843a );
 a20845a <=( a20844a  and  a20839a );
 a20849a <=( (not A267)  and  A203 );
 a20850a <=( (not A202)  and  a20849a );
 a20854a <=( (not A302)  and  (not A300) );
 a20855a <=( A268  and  a20854a );
 a20856a <=( a20855a  and  a20850a );
 a20859a <=( (not A168)  and  A170 );
 a20863a <=( (not A201)  and  A200 );
 a20864a <=( (not A199)  and  a20863a );
 a20865a <=( a20864a  and  a20859a );
 a20869a <=( (not A267)  and  A203 );
 a20870a <=( (not A202)  and  a20869a );
 a20874a <=( A299  and  A298 );
 a20875a <=( A268  and  a20874a );
 a20876a <=( a20875a  and  a20870a );
 a20879a <=( (not A168)  and  A170 );
 a20883a <=( (not A201)  and  A200 );
 a20884a <=( (not A199)  and  a20883a );
 a20885a <=( a20884a  and  a20879a );
 a20889a <=( (not A267)  and  A203 );
 a20890a <=( (not A202)  and  a20889a );
 a20894a <=( (not A299)  and  (not A298) );
 a20895a <=( A268  and  a20894a );
 a20896a <=( a20895a  and  a20890a );
 a20899a <=( (not A168)  and  A170 );
 a20903a <=( (not A201)  and  A200 );
 a20904a <=( (not A199)  and  a20903a );
 a20905a <=( a20904a  and  a20899a );
 a20909a <=( (not A267)  and  A203 );
 a20910a <=( (not A202)  and  a20909a );
 a20914a <=( A301  and  (not A300) );
 a20915a <=( (not A269)  and  a20914a );
 a20916a <=( a20915a  and  a20910a );
 a20919a <=( (not A168)  and  A170 );
 a20923a <=( (not A201)  and  A200 );
 a20924a <=( (not A199)  and  a20923a );
 a20925a <=( a20924a  and  a20919a );
 a20929a <=( (not A267)  and  A203 );
 a20930a <=( (not A202)  and  a20929a );
 a20934a <=( (not A302)  and  (not A300) );
 a20935a <=( (not A269)  and  a20934a );
 a20936a <=( a20935a  and  a20930a );
 a20939a <=( (not A168)  and  A170 );
 a20943a <=( (not A201)  and  A200 );
 a20944a <=( (not A199)  and  a20943a );
 a20945a <=( a20944a  and  a20939a );
 a20949a <=( (not A267)  and  A203 );
 a20950a <=( (not A202)  and  a20949a );
 a20954a <=( A299  and  A298 );
 a20955a <=( (not A269)  and  a20954a );
 a20956a <=( a20955a  and  a20950a );
 a20959a <=( (not A168)  and  A170 );
 a20963a <=( (not A201)  and  A200 );
 a20964a <=( (not A199)  and  a20963a );
 a20965a <=( a20964a  and  a20959a );
 a20969a <=( (not A267)  and  A203 );
 a20970a <=( (not A202)  and  a20969a );
 a20974a <=( (not A299)  and  (not A298) );
 a20975a <=( (not A269)  and  a20974a );
 a20976a <=( a20975a  and  a20970a );
 a20979a <=( (not A168)  and  A170 );
 a20983a <=( (not A201)  and  A200 );
 a20984a <=( (not A199)  and  a20983a );
 a20985a <=( a20984a  and  a20979a );
 a20989a <=( A265  and  A203 );
 a20990a <=( (not A202)  and  a20989a );
 a20994a <=( A301  and  (not A300) );
 a20995a <=( A266  and  a20994a );
 a20996a <=( a20995a  and  a20990a );
 a20999a <=( (not A168)  and  A170 );
 a21003a <=( (not A201)  and  A200 );
 a21004a <=( (not A199)  and  a21003a );
 a21005a <=( a21004a  and  a20999a );
 a21009a <=( A265  and  A203 );
 a21010a <=( (not A202)  and  a21009a );
 a21014a <=( (not A302)  and  (not A300) );
 a21015a <=( A266  and  a21014a );
 a21016a <=( a21015a  and  a21010a );
 a21019a <=( (not A168)  and  A170 );
 a21023a <=( (not A201)  and  A200 );
 a21024a <=( (not A199)  and  a21023a );
 a21025a <=( a21024a  and  a21019a );
 a21029a <=( A265  and  A203 );
 a21030a <=( (not A202)  and  a21029a );
 a21034a <=( A299  and  A298 );
 a21035a <=( A266  and  a21034a );
 a21036a <=( a21035a  and  a21030a );
 a21039a <=( (not A168)  and  A170 );
 a21043a <=( (not A201)  and  A200 );
 a21044a <=( (not A199)  and  a21043a );
 a21045a <=( a21044a  and  a21039a );
 a21049a <=( A265  and  A203 );
 a21050a <=( (not A202)  and  a21049a );
 a21054a <=( (not A299)  and  (not A298) );
 a21055a <=( A266  and  a21054a );
 a21056a <=( a21055a  and  a21050a );
 a21059a <=( (not A168)  and  A170 );
 a21063a <=( (not A201)  and  A200 );
 a21064a <=( (not A199)  and  a21063a );
 a21065a <=( a21064a  and  a21059a );
 a21069a <=( (not A265)  and  A203 );
 a21070a <=( (not A202)  and  a21069a );
 a21074a <=( A301  and  (not A300) );
 a21075a <=( (not A266)  and  a21074a );
 a21076a <=( a21075a  and  a21070a );
 a21079a <=( (not A168)  and  A170 );
 a21083a <=( (not A201)  and  A200 );
 a21084a <=( (not A199)  and  a21083a );
 a21085a <=( a21084a  and  a21079a );
 a21089a <=( (not A265)  and  A203 );
 a21090a <=( (not A202)  and  a21089a );
 a21094a <=( (not A302)  and  (not A300) );
 a21095a <=( (not A266)  and  a21094a );
 a21096a <=( a21095a  and  a21090a );
 a21099a <=( (not A168)  and  A170 );
 a21103a <=( (not A201)  and  A200 );
 a21104a <=( (not A199)  and  a21103a );
 a21105a <=( a21104a  and  a21099a );
 a21109a <=( (not A265)  and  A203 );
 a21110a <=( (not A202)  and  a21109a );
 a21114a <=( A299  and  A298 );
 a21115a <=( (not A266)  and  a21114a );
 a21116a <=( a21115a  and  a21110a );
 a21119a <=( (not A168)  and  A170 );
 a21123a <=( (not A201)  and  A200 );
 a21124a <=( (not A199)  and  a21123a );
 a21125a <=( a21124a  and  a21119a );
 a21129a <=( (not A265)  and  A203 );
 a21130a <=( (not A202)  and  a21129a );
 a21134a <=( (not A299)  and  (not A298) );
 a21135a <=( (not A266)  and  a21134a );
 a21136a <=( a21135a  and  a21130a );
 a21139a <=( (not A168)  and  A170 );
 a21143a <=( A201  and  (not A200) );
 a21144a <=( A199  and  a21143a );
 a21145a <=( a21144a  and  a21139a );
 a21149a <=( (not A268)  and  A267 );
 a21150a <=( A202  and  a21149a );
 a21154a <=( A301  and  (not A300) );
 a21155a <=( A269  and  a21154a );
 a21156a <=( a21155a  and  a21150a );
 a21159a <=( (not A168)  and  A170 );
 a21163a <=( A201  and  (not A200) );
 a21164a <=( A199  and  a21163a );
 a21165a <=( a21164a  and  a21159a );
 a21169a <=( (not A268)  and  A267 );
 a21170a <=( A202  and  a21169a );
 a21174a <=( (not A302)  and  (not A300) );
 a21175a <=( A269  and  a21174a );
 a21176a <=( a21175a  and  a21170a );
 a21179a <=( (not A168)  and  A170 );
 a21183a <=( A201  and  (not A200) );
 a21184a <=( A199  and  a21183a );
 a21185a <=( a21184a  and  a21179a );
 a21189a <=( (not A268)  and  A267 );
 a21190a <=( A202  and  a21189a );
 a21194a <=( A299  and  A298 );
 a21195a <=( A269  and  a21194a );
 a21196a <=( a21195a  and  a21190a );
 a21199a <=( (not A168)  and  A170 );
 a21203a <=( A201  and  (not A200) );
 a21204a <=( A199  and  a21203a );
 a21205a <=( a21204a  and  a21199a );
 a21209a <=( (not A268)  and  A267 );
 a21210a <=( A202  and  a21209a );
 a21214a <=( (not A299)  and  (not A298) );
 a21215a <=( A269  and  a21214a );
 a21216a <=( a21215a  and  a21210a );
 a21219a <=( (not A168)  and  A170 );
 a21223a <=( A201  and  (not A200) );
 a21224a <=( A199  and  a21223a );
 a21225a <=( a21224a  and  a21219a );
 a21229a <=( A268  and  (not A267) );
 a21230a <=( A202  and  a21229a );
 a21234a <=( A302  and  (not A301) );
 a21235a <=( A300  and  a21234a );
 a21236a <=( a21235a  and  a21230a );
 a21239a <=( (not A168)  and  A170 );
 a21243a <=( A201  and  (not A200) );
 a21244a <=( A199  and  a21243a );
 a21245a <=( a21244a  and  a21239a );
 a21249a <=( (not A269)  and  (not A267) );
 a21250a <=( A202  and  a21249a );
 a21254a <=( A302  and  (not A301) );
 a21255a <=( A300  and  a21254a );
 a21256a <=( a21255a  and  a21250a );
 a21259a <=( (not A168)  and  A170 );
 a21263a <=( A201  and  (not A200) );
 a21264a <=( A199  and  a21263a );
 a21265a <=( a21264a  and  a21259a );
 a21269a <=( A266  and  A265 );
 a21270a <=( A202  and  a21269a );
 a21274a <=( A302  and  (not A301) );
 a21275a <=( A300  and  a21274a );
 a21276a <=( a21275a  and  a21270a );
 a21279a <=( (not A168)  and  A170 );
 a21283a <=( A201  and  (not A200) );
 a21284a <=( A199  and  a21283a );
 a21285a <=( a21284a  and  a21279a );
 a21289a <=( (not A266)  and  (not A265) );
 a21290a <=( A202  and  a21289a );
 a21294a <=( A302  and  (not A301) );
 a21295a <=( A300  and  a21294a );
 a21296a <=( a21295a  and  a21290a );
 a21299a <=( (not A168)  and  A170 );
 a21303a <=( A201  and  (not A200) );
 a21304a <=( A199  and  a21303a );
 a21305a <=( a21304a  and  a21299a );
 a21309a <=( (not A268)  and  A267 );
 a21310a <=( (not A203)  and  a21309a );
 a21314a <=( A301  and  (not A300) );
 a21315a <=( A269  and  a21314a );
 a21316a <=( a21315a  and  a21310a );
 a21319a <=( (not A168)  and  A170 );
 a21323a <=( A201  and  (not A200) );
 a21324a <=( A199  and  a21323a );
 a21325a <=( a21324a  and  a21319a );
 a21329a <=( (not A268)  and  A267 );
 a21330a <=( (not A203)  and  a21329a );
 a21334a <=( (not A302)  and  (not A300) );
 a21335a <=( A269  and  a21334a );
 a21336a <=( a21335a  and  a21330a );
 a21339a <=( (not A168)  and  A170 );
 a21343a <=( A201  and  (not A200) );
 a21344a <=( A199  and  a21343a );
 a21345a <=( a21344a  and  a21339a );
 a21349a <=( (not A268)  and  A267 );
 a21350a <=( (not A203)  and  a21349a );
 a21354a <=( A299  and  A298 );
 a21355a <=( A269  and  a21354a );
 a21356a <=( a21355a  and  a21350a );
 a21359a <=( (not A168)  and  A170 );
 a21363a <=( A201  and  (not A200) );
 a21364a <=( A199  and  a21363a );
 a21365a <=( a21364a  and  a21359a );
 a21369a <=( (not A268)  and  A267 );
 a21370a <=( (not A203)  and  a21369a );
 a21374a <=( (not A299)  and  (not A298) );
 a21375a <=( A269  and  a21374a );
 a21376a <=( a21375a  and  a21370a );
 a21379a <=( (not A168)  and  A170 );
 a21383a <=( A201  and  (not A200) );
 a21384a <=( A199  and  a21383a );
 a21385a <=( a21384a  and  a21379a );
 a21389a <=( A268  and  (not A267) );
 a21390a <=( (not A203)  and  a21389a );
 a21394a <=( A302  and  (not A301) );
 a21395a <=( A300  and  a21394a );
 a21396a <=( a21395a  and  a21390a );
 a21399a <=( (not A168)  and  A170 );
 a21403a <=( A201  and  (not A200) );
 a21404a <=( A199  and  a21403a );
 a21405a <=( a21404a  and  a21399a );
 a21409a <=( (not A269)  and  (not A267) );
 a21410a <=( (not A203)  and  a21409a );
 a21414a <=( A302  and  (not A301) );
 a21415a <=( A300  and  a21414a );
 a21416a <=( a21415a  and  a21410a );
 a21419a <=( (not A168)  and  A170 );
 a21423a <=( A201  and  (not A200) );
 a21424a <=( A199  and  a21423a );
 a21425a <=( a21424a  and  a21419a );
 a21429a <=( A266  and  A265 );
 a21430a <=( (not A203)  and  a21429a );
 a21434a <=( A302  and  (not A301) );
 a21435a <=( A300  and  a21434a );
 a21436a <=( a21435a  and  a21430a );
 a21439a <=( (not A168)  and  A170 );
 a21443a <=( A201  and  (not A200) );
 a21444a <=( A199  and  a21443a );
 a21445a <=( a21444a  and  a21439a );
 a21449a <=( (not A266)  and  (not A265) );
 a21450a <=( (not A203)  and  a21449a );
 a21454a <=( A302  and  (not A301) );
 a21455a <=( A300  and  a21454a );
 a21456a <=( a21455a  and  a21450a );
 a21459a <=( (not A168)  and  A170 );
 a21463a <=( (not A201)  and  (not A200) );
 a21464a <=( A199  and  a21463a );
 a21465a <=( a21464a  and  a21459a );
 a21469a <=( (not A267)  and  A203 );
 a21470a <=( (not A202)  and  a21469a );
 a21474a <=( A301  and  (not A300) );
 a21475a <=( A268  and  a21474a );
 a21476a <=( a21475a  and  a21470a );
 a21479a <=( (not A168)  and  A170 );
 a21483a <=( (not A201)  and  (not A200) );
 a21484a <=( A199  and  a21483a );
 a21485a <=( a21484a  and  a21479a );
 a21489a <=( (not A267)  and  A203 );
 a21490a <=( (not A202)  and  a21489a );
 a21494a <=( (not A302)  and  (not A300) );
 a21495a <=( A268  and  a21494a );
 a21496a <=( a21495a  and  a21490a );
 a21499a <=( (not A168)  and  A170 );
 a21503a <=( (not A201)  and  (not A200) );
 a21504a <=( A199  and  a21503a );
 a21505a <=( a21504a  and  a21499a );
 a21509a <=( (not A267)  and  A203 );
 a21510a <=( (not A202)  and  a21509a );
 a21514a <=( A299  and  A298 );
 a21515a <=( A268  and  a21514a );
 a21516a <=( a21515a  and  a21510a );
 a21519a <=( (not A168)  and  A170 );
 a21523a <=( (not A201)  and  (not A200) );
 a21524a <=( A199  and  a21523a );
 a21525a <=( a21524a  and  a21519a );
 a21529a <=( (not A267)  and  A203 );
 a21530a <=( (not A202)  and  a21529a );
 a21534a <=( (not A299)  and  (not A298) );
 a21535a <=( A268  and  a21534a );
 a21536a <=( a21535a  and  a21530a );
 a21539a <=( (not A168)  and  A170 );
 a21543a <=( (not A201)  and  (not A200) );
 a21544a <=( A199  and  a21543a );
 a21545a <=( a21544a  and  a21539a );
 a21549a <=( (not A267)  and  A203 );
 a21550a <=( (not A202)  and  a21549a );
 a21554a <=( A301  and  (not A300) );
 a21555a <=( (not A269)  and  a21554a );
 a21556a <=( a21555a  and  a21550a );
 a21559a <=( (not A168)  and  A170 );
 a21563a <=( (not A201)  and  (not A200) );
 a21564a <=( A199  and  a21563a );
 a21565a <=( a21564a  and  a21559a );
 a21569a <=( (not A267)  and  A203 );
 a21570a <=( (not A202)  and  a21569a );
 a21574a <=( (not A302)  and  (not A300) );
 a21575a <=( (not A269)  and  a21574a );
 a21576a <=( a21575a  and  a21570a );
 a21579a <=( (not A168)  and  A170 );
 a21583a <=( (not A201)  and  (not A200) );
 a21584a <=( A199  and  a21583a );
 a21585a <=( a21584a  and  a21579a );
 a21589a <=( (not A267)  and  A203 );
 a21590a <=( (not A202)  and  a21589a );
 a21594a <=( A299  and  A298 );
 a21595a <=( (not A269)  and  a21594a );
 a21596a <=( a21595a  and  a21590a );
 a21599a <=( (not A168)  and  A170 );
 a21603a <=( (not A201)  and  (not A200) );
 a21604a <=( A199  and  a21603a );
 a21605a <=( a21604a  and  a21599a );
 a21609a <=( (not A267)  and  A203 );
 a21610a <=( (not A202)  and  a21609a );
 a21614a <=( (not A299)  and  (not A298) );
 a21615a <=( (not A269)  and  a21614a );
 a21616a <=( a21615a  and  a21610a );
 a21619a <=( (not A168)  and  A170 );
 a21623a <=( (not A201)  and  (not A200) );
 a21624a <=( A199  and  a21623a );
 a21625a <=( a21624a  and  a21619a );
 a21629a <=( A265  and  A203 );
 a21630a <=( (not A202)  and  a21629a );
 a21634a <=( A301  and  (not A300) );
 a21635a <=( A266  and  a21634a );
 a21636a <=( a21635a  and  a21630a );
 a21639a <=( (not A168)  and  A170 );
 a21643a <=( (not A201)  and  (not A200) );
 a21644a <=( A199  and  a21643a );
 a21645a <=( a21644a  and  a21639a );
 a21649a <=( A265  and  A203 );
 a21650a <=( (not A202)  and  a21649a );
 a21654a <=( (not A302)  and  (not A300) );
 a21655a <=( A266  and  a21654a );
 a21656a <=( a21655a  and  a21650a );
 a21659a <=( (not A168)  and  A170 );
 a21663a <=( (not A201)  and  (not A200) );
 a21664a <=( A199  and  a21663a );
 a21665a <=( a21664a  and  a21659a );
 a21669a <=( A265  and  A203 );
 a21670a <=( (not A202)  and  a21669a );
 a21674a <=( A299  and  A298 );
 a21675a <=( A266  and  a21674a );
 a21676a <=( a21675a  and  a21670a );
 a21679a <=( (not A168)  and  A170 );
 a21683a <=( (not A201)  and  (not A200) );
 a21684a <=( A199  and  a21683a );
 a21685a <=( a21684a  and  a21679a );
 a21689a <=( A265  and  A203 );
 a21690a <=( (not A202)  and  a21689a );
 a21694a <=( (not A299)  and  (not A298) );
 a21695a <=( A266  and  a21694a );
 a21696a <=( a21695a  and  a21690a );
 a21699a <=( (not A168)  and  A170 );
 a21703a <=( (not A201)  and  (not A200) );
 a21704a <=( A199  and  a21703a );
 a21705a <=( a21704a  and  a21699a );
 a21709a <=( (not A265)  and  A203 );
 a21710a <=( (not A202)  and  a21709a );
 a21714a <=( A301  and  (not A300) );
 a21715a <=( (not A266)  and  a21714a );
 a21716a <=( a21715a  and  a21710a );
 a21719a <=( (not A168)  and  A170 );
 a21723a <=( (not A201)  and  (not A200) );
 a21724a <=( A199  and  a21723a );
 a21725a <=( a21724a  and  a21719a );
 a21729a <=( (not A265)  and  A203 );
 a21730a <=( (not A202)  and  a21729a );
 a21734a <=( (not A302)  and  (not A300) );
 a21735a <=( (not A266)  and  a21734a );
 a21736a <=( a21735a  and  a21730a );
 a21739a <=( (not A168)  and  A170 );
 a21743a <=( (not A201)  and  (not A200) );
 a21744a <=( A199  and  a21743a );
 a21745a <=( a21744a  and  a21739a );
 a21749a <=( (not A265)  and  A203 );
 a21750a <=( (not A202)  and  a21749a );
 a21754a <=( A299  and  A298 );
 a21755a <=( (not A266)  and  a21754a );
 a21756a <=( a21755a  and  a21750a );
 a21759a <=( (not A168)  and  A170 );
 a21763a <=( (not A201)  and  (not A200) );
 a21764a <=( A199  and  a21763a );
 a21765a <=( a21764a  and  a21759a );
 a21769a <=( (not A265)  and  A203 );
 a21770a <=( (not A202)  and  a21769a );
 a21774a <=( (not A299)  and  (not A298) );
 a21775a <=( (not A266)  and  a21774a );
 a21776a <=( a21775a  and  a21770a );
 a21779a <=( (not A168)  and  A169 );
 a21783a <=( A201  and  A200 );
 a21784a <=( (not A199)  and  a21783a );
 a21785a <=( a21784a  and  a21779a );
 a21789a <=( (not A268)  and  A267 );
 a21790a <=( A202  and  a21789a );
 a21794a <=( A301  and  (not A300) );
 a21795a <=( A269  and  a21794a );
 a21796a <=( a21795a  and  a21790a );
 a21799a <=( (not A168)  and  A169 );
 a21803a <=( A201  and  A200 );
 a21804a <=( (not A199)  and  a21803a );
 a21805a <=( a21804a  and  a21799a );
 a21809a <=( (not A268)  and  A267 );
 a21810a <=( A202  and  a21809a );
 a21814a <=( (not A302)  and  (not A300) );
 a21815a <=( A269  and  a21814a );
 a21816a <=( a21815a  and  a21810a );
 a21819a <=( (not A168)  and  A169 );
 a21823a <=( A201  and  A200 );
 a21824a <=( (not A199)  and  a21823a );
 a21825a <=( a21824a  and  a21819a );
 a21829a <=( (not A268)  and  A267 );
 a21830a <=( A202  and  a21829a );
 a21834a <=( A299  and  A298 );
 a21835a <=( A269  and  a21834a );
 a21836a <=( a21835a  and  a21830a );
 a21839a <=( (not A168)  and  A169 );
 a21843a <=( A201  and  A200 );
 a21844a <=( (not A199)  and  a21843a );
 a21845a <=( a21844a  and  a21839a );
 a21849a <=( (not A268)  and  A267 );
 a21850a <=( A202  and  a21849a );
 a21854a <=( (not A299)  and  (not A298) );
 a21855a <=( A269  and  a21854a );
 a21856a <=( a21855a  and  a21850a );
 a21859a <=( (not A168)  and  A169 );
 a21863a <=( A201  and  A200 );
 a21864a <=( (not A199)  and  a21863a );
 a21865a <=( a21864a  and  a21859a );
 a21869a <=( A268  and  (not A267) );
 a21870a <=( A202  and  a21869a );
 a21874a <=( A302  and  (not A301) );
 a21875a <=( A300  and  a21874a );
 a21876a <=( a21875a  and  a21870a );
 a21879a <=( (not A168)  and  A169 );
 a21883a <=( A201  and  A200 );
 a21884a <=( (not A199)  and  a21883a );
 a21885a <=( a21884a  and  a21879a );
 a21889a <=( (not A269)  and  (not A267) );
 a21890a <=( A202  and  a21889a );
 a21894a <=( A302  and  (not A301) );
 a21895a <=( A300  and  a21894a );
 a21896a <=( a21895a  and  a21890a );
 a21899a <=( (not A168)  and  A169 );
 a21903a <=( A201  and  A200 );
 a21904a <=( (not A199)  and  a21903a );
 a21905a <=( a21904a  and  a21899a );
 a21909a <=( A266  and  A265 );
 a21910a <=( A202  and  a21909a );
 a21914a <=( A302  and  (not A301) );
 a21915a <=( A300  and  a21914a );
 a21916a <=( a21915a  and  a21910a );
 a21919a <=( (not A168)  and  A169 );
 a21923a <=( A201  and  A200 );
 a21924a <=( (not A199)  and  a21923a );
 a21925a <=( a21924a  and  a21919a );
 a21929a <=( (not A266)  and  (not A265) );
 a21930a <=( A202  and  a21929a );
 a21934a <=( A302  and  (not A301) );
 a21935a <=( A300  and  a21934a );
 a21936a <=( a21935a  and  a21930a );
 a21939a <=( (not A168)  and  A169 );
 a21943a <=( A201  and  A200 );
 a21944a <=( (not A199)  and  a21943a );
 a21945a <=( a21944a  and  a21939a );
 a21949a <=( (not A268)  and  A267 );
 a21950a <=( (not A203)  and  a21949a );
 a21954a <=( A301  and  (not A300) );
 a21955a <=( A269  and  a21954a );
 a21956a <=( a21955a  and  a21950a );
 a21959a <=( (not A168)  and  A169 );
 a21963a <=( A201  and  A200 );
 a21964a <=( (not A199)  and  a21963a );
 a21965a <=( a21964a  and  a21959a );
 a21969a <=( (not A268)  and  A267 );
 a21970a <=( (not A203)  and  a21969a );
 a21974a <=( (not A302)  and  (not A300) );
 a21975a <=( A269  and  a21974a );
 a21976a <=( a21975a  and  a21970a );
 a21979a <=( (not A168)  and  A169 );
 a21983a <=( A201  and  A200 );
 a21984a <=( (not A199)  and  a21983a );
 a21985a <=( a21984a  and  a21979a );
 a21989a <=( (not A268)  and  A267 );
 a21990a <=( (not A203)  and  a21989a );
 a21994a <=( A299  and  A298 );
 a21995a <=( A269  and  a21994a );
 a21996a <=( a21995a  and  a21990a );
 a21999a <=( (not A168)  and  A169 );
 a22003a <=( A201  and  A200 );
 a22004a <=( (not A199)  and  a22003a );
 a22005a <=( a22004a  and  a21999a );
 a22009a <=( (not A268)  and  A267 );
 a22010a <=( (not A203)  and  a22009a );
 a22014a <=( (not A299)  and  (not A298) );
 a22015a <=( A269  and  a22014a );
 a22016a <=( a22015a  and  a22010a );
 a22019a <=( (not A168)  and  A169 );
 a22023a <=( A201  and  A200 );
 a22024a <=( (not A199)  and  a22023a );
 a22025a <=( a22024a  and  a22019a );
 a22029a <=( A268  and  (not A267) );
 a22030a <=( (not A203)  and  a22029a );
 a22034a <=( A302  and  (not A301) );
 a22035a <=( A300  and  a22034a );
 a22036a <=( a22035a  and  a22030a );
 a22039a <=( (not A168)  and  A169 );
 a22043a <=( A201  and  A200 );
 a22044a <=( (not A199)  and  a22043a );
 a22045a <=( a22044a  and  a22039a );
 a22049a <=( (not A269)  and  (not A267) );
 a22050a <=( (not A203)  and  a22049a );
 a22054a <=( A302  and  (not A301) );
 a22055a <=( A300  and  a22054a );
 a22056a <=( a22055a  and  a22050a );
 a22059a <=( (not A168)  and  A169 );
 a22063a <=( A201  and  A200 );
 a22064a <=( (not A199)  and  a22063a );
 a22065a <=( a22064a  and  a22059a );
 a22069a <=( A266  and  A265 );
 a22070a <=( (not A203)  and  a22069a );
 a22074a <=( A302  and  (not A301) );
 a22075a <=( A300  and  a22074a );
 a22076a <=( a22075a  and  a22070a );
 a22079a <=( (not A168)  and  A169 );
 a22083a <=( A201  and  A200 );
 a22084a <=( (not A199)  and  a22083a );
 a22085a <=( a22084a  and  a22079a );
 a22089a <=( (not A266)  and  (not A265) );
 a22090a <=( (not A203)  and  a22089a );
 a22094a <=( A302  and  (not A301) );
 a22095a <=( A300  and  a22094a );
 a22096a <=( a22095a  and  a22090a );
 a22099a <=( (not A168)  and  A169 );
 a22103a <=( (not A201)  and  A200 );
 a22104a <=( (not A199)  and  a22103a );
 a22105a <=( a22104a  and  a22099a );
 a22109a <=( (not A267)  and  A203 );
 a22110a <=( (not A202)  and  a22109a );
 a22114a <=( A301  and  (not A300) );
 a22115a <=( A268  and  a22114a );
 a22116a <=( a22115a  and  a22110a );
 a22119a <=( (not A168)  and  A169 );
 a22123a <=( (not A201)  and  A200 );
 a22124a <=( (not A199)  and  a22123a );
 a22125a <=( a22124a  and  a22119a );
 a22129a <=( (not A267)  and  A203 );
 a22130a <=( (not A202)  and  a22129a );
 a22134a <=( (not A302)  and  (not A300) );
 a22135a <=( A268  and  a22134a );
 a22136a <=( a22135a  and  a22130a );
 a22139a <=( (not A168)  and  A169 );
 a22143a <=( (not A201)  and  A200 );
 a22144a <=( (not A199)  and  a22143a );
 a22145a <=( a22144a  and  a22139a );
 a22149a <=( (not A267)  and  A203 );
 a22150a <=( (not A202)  and  a22149a );
 a22154a <=( A299  and  A298 );
 a22155a <=( A268  and  a22154a );
 a22156a <=( a22155a  and  a22150a );
 a22159a <=( (not A168)  and  A169 );
 a22163a <=( (not A201)  and  A200 );
 a22164a <=( (not A199)  and  a22163a );
 a22165a <=( a22164a  and  a22159a );
 a22169a <=( (not A267)  and  A203 );
 a22170a <=( (not A202)  and  a22169a );
 a22174a <=( (not A299)  and  (not A298) );
 a22175a <=( A268  and  a22174a );
 a22176a <=( a22175a  and  a22170a );
 a22179a <=( (not A168)  and  A169 );
 a22183a <=( (not A201)  and  A200 );
 a22184a <=( (not A199)  and  a22183a );
 a22185a <=( a22184a  and  a22179a );
 a22189a <=( (not A267)  and  A203 );
 a22190a <=( (not A202)  and  a22189a );
 a22194a <=( A301  and  (not A300) );
 a22195a <=( (not A269)  and  a22194a );
 a22196a <=( a22195a  and  a22190a );
 a22199a <=( (not A168)  and  A169 );
 a22203a <=( (not A201)  and  A200 );
 a22204a <=( (not A199)  and  a22203a );
 a22205a <=( a22204a  and  a22199a );
 a22209a <=( (not A267)  and  A203 );
 a22210a <=( (not A202)  and  a22209a );
 a22214a <=( (not A302)  and  (not A300) );
 a22215a <=( (not A269)  and  a22214a );
 a22216a <=( a22215a  and  a22210a );
 a22219a <=( (not A168)  and  A169 );
 a22223a <=( (not A201)  and  A200 );
 a22224a <=( (not A199)  and  a22223a );
 a22225a <=( a22224a  and  a22219a );
 a22229a <=( (not A267)  and  A203 );
 a22230a <=( (not A202)  and  a22229a );
 a22234a <=( A299  and  A298 );
 a22235a <=( (not A269)  and  a22234a );
 a22236a <=( a22235a  and  a22230a );
 a22239a <=( (not A168)  and  A169 );
 a22243a <=( (not A201)  and  A200 );
 a22244a <=( (not A199)  and  a22243a );
 a22245a <=( a22244a  and  a22239a );
 a22249a <=( (not A267)  and  A203 );
 a22250a <=( (not A202)  and  a22249a );
 a22254a <=( (not A299)  and  (not A298) );
 a22255a <=( (not A269)  and  a22254a );
 a22256a <=( a22255a  and  a22250a );
 a22259a <=( (not A168)  and  A169 );
 a22263a <=( (not A201)  and  A200 );
 a22264a <=( (not A199)  and  a22263a );
 a22265a <=( a22264a  and  a22259a );
 a22269a <=( A265  and  A203 );
 a22270a <=( (not A202)  and  a22269a );
 a22274a <=( A301  and  (not A300) );
 a22275a <=( A266  and  a22274a );
 a22276a <=( a22275a  and  a22270a );
 a22279a <=( (not A168)  and  A169 );
 a22283a <=( (not A201)  and  A200 );
 a22284a <=( (not A199)  and  a22283a );
 a22285a <=( a22284a  and  a22279a );
 a22289a <=( A265  and  A203 );
 a22290a <=( (not A202)  and  a22289a );
 a22294a <=( (not A302)  and  (not A300) );
 a22295a <=( A266  and  a22294a );
 a22296a <=( a22295a  and  a22290a );
 a22299a <=( (not A168)  and  A169 );
 a22303a <=( (not A201)  and  A200 );
 a22304a <=( (not A199)  and  a22303a );
 a22305a <=( a22304a  and  a22299a );
 a22309a <=( A265  and  A203 );
 a22310a <=( (not A202)  and  a22309a );
 a22314a <=( A299  and  A298 );
 a22315a <=( A266  and  a22314a );
 a22316a <=( a22315a  and  a22310a );
 a22319a <=( (not A168)  and  A169 );
 a22323a <=( (not A201)  and  A200 );
 a22324a <=( (not A199)  and  a22323a );
 a22325a <=( a22324a  and  a22319a );
 a22329a <=( A265  and  A203 );
 a22330a <=( (not A202)  and  a22329a );
 a22334a <=( (not A299)  and  (not A298) );
 a22335a <=( A266  and  a22334a );
 a22336a <=( a22335a  and  a22330a );
 a22339a <=( (not A168)  and  A169 );
 a22343a <=( (not A201)  and  A200 );
 a22344a <=( (not A199)  and  a22343a );
 a22345a <=( a22344a  and  a22339a );
 a22349a <=( (not A265)  and  A203 );
 a22350a <=( (not A202)  and  a22349a );
 a22354a <=( A301  and  (not A300) );
 a22355a <=( (not A266)  and  a22354a );
 a22356a <=( a22355a  and  a22350a );
 a22359a <=( (not A168)  and  A169 );
 a22363a <=( (not A201)  and  A200 );
 a22364a <=( (not A199)  and  a22363a );
 a22365a <=( a22364a  and  a22359a );
 a22369a <=( (not A265)  and  A203 );
 a22370a <=( (not A202)  and  a22369a );
 a22374a <=( (not A302)  and  (not A300) );
 a22375a <=( (not A266)  and  a22374a );
 a22376a <=( a22375a  and  a22370a );
 a22379a <=( (not A168)  and  A169 );
 a22383a <=( (not A201)  and  A200 );
 a22384a <=( (not A199)  and  a22383a );
 a22385a <=( a22384a  and  a22379a );
 a22389a <=( (not A265)  and  A203 );
 a22390a <=( (not A202)  and  a22389a );
 a22394a <=( A299  and  A298 );
 a22395a <=( (not A266)  and  a22394a );
 a22396a <=( a22395a  and  a22390a );
 a22399a <=( (not A168)  and  A169 );
 a22403a <=( (not A201)  and  A200 );
 a22404a <=( (not A199)  and  a22403a );
 a22405a <=( a22404a  and  a22399a );
 a22409a <=( (not A265)  and  A203 );
 a22410a <=( (not A202)  and  a22409a );
 a22414a <=( (not A299)  and  (not A298) );
 a22415a <=( (not A266)  and  a22414a );
 a22416a <=( a22415a  and  a22410a );
 a22419a <=( (not A168)  and  A169 );
 a22423a <=( A201  and  (not A200) );
 a22424a <=( A199  and  a22423a );
 a22425a <=( a22424a  and  a22419a );
 a22429a <=( (not A268)  and  A267 );
 a22430a <=( A202  and  a22429a );
 a22434a <=( A301  and  (not A300) );
 a22435a <=( A269  and  a22434a );
 a22436a <=( a22435a  and  a22430a );
 a22439a <=( (not A168)  and  A169 );
 a22443a <=( A201  and  (not A200) );
 a22444a <=( A199  and  a22443a );
 a22445a <=( a22444a  and  a22439a );
 a22449a <=( (not A268)  and  A267 );
 a22450a <=( A202  and  a22449a );
 a22454a <=( (not A302)  and  (not A300) );
 a22455a <=( A269  and  a22454a );
 a22456a <=( a22455a  and  a22450a );
 a22459a <=( (not A168)  and  A169 );
 a22463a <=( A201  and  (not A200) );
 a22464a <=( A199  and  a22463a );
 a22465a <=( a22464a  and  a22459a );
 a22469a <=( (not A268)  and  A267 );
 a22470a <=( A202  and  a22469a );
 a22474a <=( A299  and  A298 );
 a22475a <=( A269  and  a22474a );
 a22476a <=( a22475a  and  a22470a );
 a22479a <=( (not A168)  and  A169 );
 a22483a <=( A201  and  (not A200) );
 a22484a <=( A199  and  a22483a );
 a22485a <=( a22484a  and  a22479a );
 a22489a <=( (not A268)  and  A267 );
 a22490a <=( A202  and  a22489a );
 a22494a <=( (not A299)  and  (not A298) );
 a22495a <=( A269  and  a22494a );
 a22496a <=( a22495a  and  a22490a );
 a22499a <=( (not A168)  and  A169 );
 a22503a <=( A201  and  (not A200) );
 a22504a <=( A199  and  a22503a );
 a22505a <=( a22504a  and  a22499a );
 a22509a <=( A268  and  (not A267) );
 a22510a <=( A202  and  a22509a );
 a22514a <=( A302  and  (not A301) );
 a22515a <=( A300  and  a22514a );
 a22516a <=( a22515a  and  a22510a );
 a22519a <=( (not A168)  and  A169 );
 a22523a <=( A201  and  (not A200) );
 a22524a <=( A199  and  a22523a );
 a22525a <=( a22524a  and  a22519a );
 a22529a <=( (not A269)  and  (not A267) );
 a22530a <=( A202  and  a22529a );
 a22534a <=( A302  and  (not A301) );
 a22535a <=( A300  and  a22534a );
 a22536a <=( a22535a  and  a22530a );
 a22539a <=( (not A168)  and  A169 );
 a22543a <=( A201  and  (not A200) );
 a22544a <=( A199  and  a22543a );
 a22545a <=( a22544a  and  a22539a );
 a22549a <=( A266  and  A265 );
 a22550a <=( A202  and  a22549a );
 a22554a <=( A302  and  (not A301) );
 a22555a <=( A300  and  a22554a );
 a22556a <=( a22555a  and  a22550a );
 a22559a <=( (not A168)  and  A169 );
 a22563a <=( A201  and  (not A200) );
 a22564a <=( A199  and  a22563a );
 a22565a <=( a22564a  and  a22559a );
 a22569a <=( (not A266)  and  (not A265) );
 a22570a <=( A202  and  a22569a );
 a22574a <=( A302  and  (not A301) );
 a22575a <=( A300  and  a22574a );
 a22576a <=( a22575a  and  a22570a );
 a22579a <=( (not A168)  and  A169 );
 a22583a <=( A201  and  (not A200) );
 a22584a <=( A199  and  a22583a );
 a22585a <=( a22584a  and  a22579a );
 a22589a <=( (not A268)  and  A267 );
 a22590a <=( (not A203)  and  a22589a );
 a22594a <=( A301  and  (not A300) );
 a22595a <=( A269  and  a22594a );
 a22596a <=( a22595a  and  a22590a );
 a22599a <=( (not A168)  and  A169 );
 a22603a <=( A201  and  (not A200) );
 a22604a <=( A199  and  a22603a );
 a22605a <=( a22604a  and  a22599a );
 a22609a <=( (not A268)  and  A267 );
 a22610a <=( (not A203)  and  a22609a );
 a22614a <=( (not A302)  and  (not A300) );
 a22615a <=( A269  and  a22614a );
 a22616a <=( a22615a  and  a22610a );
 a22619a <=( (not A168)  and  A169 );
 a22623a <=( A201  and  (not A200) );
 a22624a <=( A199  and  a22623a );
 a22625a <=( a22624a  and  a22619a );
 a22629a <=( (not A268)  and  A267 );
 a22630a <=( (not A203)  and  a22629a );
 a22634a <=( A299  and  A298 );
 a22635a <=( A269  and  a22634a );
 a22636a <=( a22635a  and  a22630a );
 a22639a <=( (not A168)  and  A169 );
 a22643a <=( A201  and  (not A200) );
 a22644a <=( A199  and  a22643a );
 a22645a <=( a22644a  and  a22639a );
 a22649a <=( (not A268)  and  A267 );
 a22650a <=( (not A203)  and  a22649a );
 a22654a <=( (not A299)  and  (not A298) );
 a22655a <=( A269  and  a22654a );
 a22656a <=( a22655a  and  a22650a );
 a22659a <=( (not A168)  and  A169 );
 a22663a <=( A201  and  (not A200) );
 a22664a <=( A199  and  a22663a );
 a22665a <=( a22664a  and  a22659a );
 a22669a <=( A268  and  (not A267) );
 a22670a <=( (not A203)  and  a22669a );
 a22674a <=( A302  and  (not A301) );
 a22675a <=( A300  and  a22674a );
 a22676a <=( a22675a  and  a22670a );
 a22679a <=( (not A168)  and  A169 );
 a22683a <=( A201  and  (not A200) );
 a22684a <=( A199  and  a22683a );
 a22685a <=( a22684a  and  a22679a );
 a22689a <=( (not A269)  and  (not A267) );
 a22690a <=( (not A203)  and  a22689a );
 a22694a <=( A302  and  (not A301) );
 a22695a <=( A300  and  a22694a );
 a22696a <=( a22695a  and  a22690a );
 a22699a <=( (not A168)  and  A169 );
 a22703a <=( A201  and  (not A200) );
 a22704a <=( A199  and  a22703a );
 a22705a <=( a22704a  and  a22699a );
 a22709a <=( A266  and  A265 );
 a22710a <=( (not A203)  and  a22709a );
 a22714a <=( A302  and  (not A301) );
 a22715a <=( A300  and  a22714a );
 a22716a <=( a22715a  and  a22710a );
 a22719a <=( (not A168)  and  A169 );
 a22723a <=( A201  and  (not A200) );
 a22724a <=( A199  and  a22723a );
 a22725a <=( a22724a  and  a22719a );
 a22729a <=( (not A266)  and  (not A265) );
 a22730a <=( (not A203)  and  a22729a );
 a22734a <=( A302  and  (not A301) );
 a22735a <=( A300  and  a22734a );
 a22736a <=( a22735a  and  a22730a );
 a22739a <=( (not A168)  and  A169 );
 a22743a <=( (not A201)  and  (not A200) );
 a22744a <=( A199  and  a22743a );
 a22745a <=( a22744a  and  a22739a );
 a22749a <=( (not A267)  and  A203 );
 a22750a <=( (not A202)  and  a22749a );
 a22754a <=( A301  and  (not A300) );
 a22755a <=( A268  and  a22754a );
 a22756a <=( a22755a  and  a22750a );
 a22759a <=( (not A168)  and  A169 );
 a22763a <=( (not A201)  and  (not A200) );
 a22764a <=( A199  and  a22763a );
 a22765a <=( a22764a  and  a22759a );
 a22769a <=( (not A267)  and  A203 );
 a22770a <=( (not A202)  and  a22769a );
 a22774a <=( (not A302)  and  (not A300) );
 a22775a <=( A268  and  a22774a );
 a22776a <=( a22775a  and  a22770a );
 a22779a <=( (not A168)  and  A169 );
 a22783a <=( (not A201)  and  (not A200) );
 a22784a <=( A199  and  a22783a );
 a22785a <=( a22784a  and  a22779a );
 a22789a <=( (not A267)  and  A203 );
 a22790a <=( (not A202)  and  a22789a );
 a22794a <=( A299  and  A298 );
 a22795a <=( A268  and  a22794a );
 a22796a <=( a22795a  and  a22790a );
 a22799a <=( (not A168)  and  A169 );
 a22803a <=( (not A201)  and  (not A200) );
 a22804a <=( A199  and  a22803a );
 a22805a <=( a22804a  and  a22799a );
 a22809a <=( (not A267)  and  A203 );
 a22810a <=( (not A202)  and  a22809a );
 a22814a <=( (not A299)  and  (not A298) );
 a22815a <=( A268  and  a22814a );
 a22816a <=( a22815a  and  a22810a );
 a22819a <=( (not A168)  and  A169 );
 a22823a <=( (not A201)  and  (not A200) );
 a22824a <=( A199  and  a22823a );
 a22825a <=( a22824a  and  a22819a );
 a22829a <=( (not A267)  and  A203 );
 a22830a <=( (not A202)  and  a22829a );
 a22834a <=( A301  and  (not A300) );
 a22835a <=( (not A269)  and  a22834a );
 a22836a <=( a22835a  and  a22830a );
 a22839a <=( (not A168)  and  A169 );
 a22843a <=( (not A201)  and  (not A200) );
 a22844a <=( A199  and  a22843a );
 a22845a <=( a22844a  and  a22839a );
 a22849a <=( (not A267)  and  A203 );
 a22850a <=( (not A202)  and  a22849a );
 a22854a <=( (not A302)  and  (not A300) );
 a22855a <=( (not A269)  and  a22854a );
 a22856a <=( a22855a  and  a22850a );
 a22859a <=( (not A168)  and  A169 );
 a22863a <=( (not A201)  and  (not A200) );
 a22864a <=( A199  and  a22863a );
 a22865a <=( a22864a  and  a22859a );
 a22869a <=( (not A267)  and  A203 );
 a22870a <=( (not A202)  and  a22869a );
 a22874a <=( A299  and  A298 );
 a22875a <=( (not A269)  and  a22874a );
 a22876a <=( a22875a  and  a22870a );
 a22879a <=( (not A168)  and  A169 );
 a22883a <=( (not A201)  and  (not A200) );
 a22884a <=( A199  and  a22883a );
 a22885a <=( a22884a  and  a22879a );
 a22889a <=( (not A267)  and  A203 );
 a22890a <=( (not A202)  and  a22889a );
 a22894a <=( (not A299)  and  (not A298) );
 a22895a <=( (not A269)  and  a22894a );
 a22896a <=( a22895a  and  a22890a );
 a22899a <=( (not A168)  and  A169 );
 a22903a <=( (not A201)  and  (not A200) );
 a22904a <=( A199  and  a22903a );
 a22905a <=( a22904a  and  a22899a );
 a22909a <=( A265  and  A203 );
 a22910a <=( (not A202)  and  a22909a );
 a22914a <=( A301  and  (not A300) );
 a22915a <=( A266  and  a22914a );
 a22916a <=( a22915a  and  a22910a );
 a22919a <=( (not A168)  and  A169 );
 a22923a <=( (not A201)  and  (not A200) );
 a22924a <=( A199  and  a22923a );
 a22925a <=( a22924a  and  a22919a );
 a22929a <=( A265  and  A203 );
 a22930a <=( (not A202)  and  a22929a );
 a22934a <=( (not A302)  and  (not A300) );
 a22935a <=( A266  and  a22934a );
 a22936a <=( a22935a  and  a22930a );
 a22939a <=( (not A168)  and  A169 );
 a22943a <=( (not A201)  and  (not A200) );
 a22944a <=( A199  and  a22943a );
 a22945a <=( a22944a  and  a22939a );
 a22949a <=( A265  and  A203 );
 a22950a <=( (not A202)  and  a22949a );
 a22954a <=( A299  and  A298 );
 a22955a <=( A266  and  a22954a );
 a22956a <=( a22955a  and  a22950a );
 a22959a <=( (not A168)  and  A169 );
 a22963a <=( (not A201)  and  (not A200) );
 a22964a <=( A199  and  a22963a );
 a22965a <=( a22964a  and  a22959a );
 a22969a <=( A265  and  A203 );
 a22970a <=( (not A202)  and  a22969a );
 a22974a <=( (not A299)  and  (not A298) );
 a22975a <=( A266  and  a22974a );
 a22976a <=( a22975a  and  a22970a );
 a22979a <=( (not A168)  and  A169 );
 a22983a <=( (not A201)  and  (not A200) );
 a22984a <=( A199  and  a22983a );
 a22985a <=( a22984a  and  a22979a );
 a22989a <=( (not A265)  and  A203 );
 a22990a <=( (not A202)  and  a22989a );
 a22994a <=( A301  and  (not A300) );
 a22995a <=( (not A266)  and  a22994a );
 a22996a <=( a22995a  and  a22990a );
 a22999a <=( (not A168)  and  A169 );
 a23003a <=( (not A201)  and  (not A200) );
 a23004a <=( A199  and  a23003a );
 a23005a <=( a23004a  and  a22999a );
 a23009a <=( (not A265)  and  A203 );
 a23010a <=( (not A202)  and  a23009a );
 a23014a <=( (not A302)  and  (not A300) );
 a23015a <=( (not A266)  and  a23014a );
 a23016a <=( a23015a  and  a23010a );
 a23019a <=( (not A168)  and  A169 );
 a23023a <=( (not A201)  and  (not A200) );
 a23024a <=( A199  and  a23023a );
 a23025a <=( a23024a  and  a23019a );
 a23029a <=( (not A265)  and  A203 );
 a23030a <=( (not A202)  and  a23029a );
 a23034a <=( A299  and  A298 );
 a23035a <=( (not A266)  and  a23034a );
 a23036a <=( a23035a  and  a23030a );
 a23039a <=( (not A168)  and  A169 );
 a23043a <=( (not A201)  and  (not A200) );
 a23044a <=( A199  and  a23043a );
 a23045a <=( a23044a  and  a23039a );
 a23049a <=( (not A265)  and  A203 );
 a23050a <=( (not A202)  and  a23049a );
 a23054a <=( (not A299)  and  (not A298) );
 a23055a <=( (not A266)  and  a23054a );
 a23056a <=( a23055a  and  a23050a );
 a23059a <=( (not A169)  and  (not A170) );
 a23063a <=( A234  and  A233 );
 a23064a <=( (not A232)  and  a23063a );
 a23065a <=( a23064a  and  a23059a );
 a23069a <=( A266  and  (not A265) );
 a23070a <=( A235  and  a23069a );
 a23074a <=( A269  and  (not A268) );
 a23075a <=( (not A267)  and  a23074a );
 a23076a <=( a23075a  and  a23070a );
 a23079a <=( (not A169)  and  (not A170) );
 a23083a <=( A234  and  A233 );
 a23084a <=( (not A232)  and  a23083a );
 a23085a <=( a23084a  and  a23079a );
 a23089a <=( (not A266)  and  A265 );
 a23090a <=( A235  and  a23089a );
 a23094a <=( A269  and  (not A268) );
 a23095a <=( (not A267)  and  a23094a );
 a23096a <=( a23095a  and  a23090a );
 a23099a <=( (not A169)  and  (not A170) );
 a23103a <=( A234  and  A233 );
 a23104a <=( (not A232)  and  a23103a );
 a23105a <=( a23104a  and  a23099a );
 a23109a <=( A266  and  (not A265) );
 a23110a <=( (not A236)  and  a23109a );
 a23114a <=( A269  and  (not A268) );
 a23115a <=( (not A267)  and  a23114a );
 a23116a <=( a23115a  and  a23110a );
 a23119a <=( (not A169)  and  (not A170) );
 a23123a <=( A234  and  A233 );
 a23124a <=( (not A232)  and  a23123a );
 a23125a <=( a23124a  and  a23119a );
 a23129a <=( (not A266)  and  A265 );
 a23130a <=( (not A236)  and  a23129a );
 a23134a <=( A269  and  (not A268) );
 a23135a <=( (not A267)  and  a23134a );
 a23136a <=( a23135a  and  a23130a );
 a23139a <=( (not A169)  and  (not A170) );
 a23143a <=( A234  and  (not A233) );
 a23144a <=( A232  and  a23143a );
 a23145a <=( a23144a  and  a23139a );
 a23149a <=( A266  and  (not A265) );
 a23150a <=( A235  and  a23149a );
 a23154a <=( A269  and  (not A268) );
 a23155a <=( (not A267)  and  a23154a );
 a23156a <=( a23155a  and  a23150a );
 a23159a <=( (not A169)  and  (not A170) );
 a23163a <=( A234  and  (not A233) );
 a23164a <=( A232  and  a23163a );
 a23165a <=( a23164a  and  a23159a );
 a23169a <=( (not A266)  and  A265 );
 a23170a <=( A235  and  a23169a );
 a23174a <=( A269  and  (not A268) );
 a23175a <=( (not A267)  and  a23174a );
 a23176a <=( a23175a  and  a23170a );
 a23179a <=( (not A169)  and  (not A170) );
 a23183a <=( A234  and  (not A233) );
 a23184a <=( A232  and  a23183a );
 a23185a <=( a23184a  and  a23179a );
 a23189a <=( A266  and  (not A265) );
 a23190a <=( (not A236)  and  a23189a );
 a23194a <=( A269  and  (not A268) );
 a23195a <=( (not A267)  and  a23194a );
 a23196a <=( a23195a  and  a23190a );
 a23199a <=( (not A169)  and  (not A170) );
 a23203a <=( A234  and  (not A233) );
 a23204a <=( A232  and  a23203a );
 a23205a <=( a23204a  and  a23199a );
 a23209a <=( (not A266)  and  A265 );
 a23210a <=( (not A236)  and  a23209a );
 a23214a <=( A269  and  (not A268) );
 a23215a <=( (not A267)  and  a23214a );
 a23216a <=( a23215a  and  a23210a );
 a23219a <=( (not A169)  and  (not A170) );
 a23223a <=( A200  and  (not A199) );
 a23224a <=( A168  and  a23223a );
 a23225a <=( a23224a  and  a23219a );
 a23229a <=( (not A267)  and  A202 );
 a23230a <=( A201  and  a23229a );
 a23234a <=( A301  and  (not A300) );
 a23235a <=( A268  and  a23234a );
 a23236a <=( a23235a  and  a23230a );
 a23239a <=( (not A169)  and  (not A170) );
 a23243a <=( A200  and  (not A199) );
 a23244a <=( A168  and  a23243a );
 a23245a <=( a23244a  and  a23239a );
 a23249a <=( (not A267)  and  A202 );
 a23250a <=( A201  and  a23249a );
 a23254a <=( (not A302)  and  (not A300) );
 a23255a <=( A268  and  a23254a );
 a23256a <=( a23255a  and  a23250a );
 a23259a <=( (not A169)  and  (not A170) );
 a23263a <=( A200  and  (not A199) );
 a23264a <=( A168  and  a23263a );
 a23265a <=( a23264a  and  a23259a );
 a23269a <=( (not A267)  and  A202 );
 a23270a <=( A201  and  a23269a );
 a23274a <=( A299  and  A298 );
 a23275a <=( A268  and  a23274a );
 a23276a <=( a23275a  and  a23270a );
 a23279a <=( (not A169)  and  (not A170) );
 a23283a <=( A200  and  (not A199) );
 a23284a <=( A168  and  a23283a );
 a23285a <=( a23284a  and  a23279a );
 a23289a <=( (not A267)  and  A202 );
 a23290a <=( A201  and  a23289a );
 a23294a <=( (not A299)  and  (not A298) );
 a23295a <=( A268  and  a23294a );
 a23296a <=( a23295a  and  a23290a );
 a23299a <=( (not A169)  and  (not A170) );
 a23303a <=( A200  and  (not A199) );
 a23304a <=( A168  and  a23303a );
 a23305a <=( a23304a  and  a23299a );
 a23309a <=( (not A267)  and  A202 );
 a23310a <=( A201  and  a23309a );
 a23314a <=( A301  and  (not A300) );
 a23315a <=( (not A269)  and  a23314a );
 a23316a <=( a23315a  and  a23310a );
 a23319a <=( (not A169)  and  (not A170) );
 a23323a <=( A200  and  (not A199) );
 a23324a <=( A168  and  a23323a );
 a23325a <=( a23324a  and  a23319a );
 a23329a <=( (not A267)  and  A202 );
 a23330a <=( A201  and  a23329a );
 a23334a <=( (not A302)  and  (not A300) );
 a23335a <=( (not A269)  and  a23334a );
 a23336a <=( a23335a  and  a23330a );
 a23339a <=( (not A169)  and  (not A170) );
 a23343a <=( A200  and  (not A199) );
 a23344a <=( A168  and  a23343a );
 a23345a <=( a23344a  and  a23339a );
 a23349a <=( (not A267)  and  A202 );
 a23350a <=( A201  and  a23349a );
 a23354a <=( A299  and  A298 );
 a23355a <=( (not A269)  and  a23354a );
 a23356a <=( a23355a  and  a23350a );
 a23359a <=( (not A169)  and  (not A170) );
 a23363a <=( A200  and  (not A199) );
 a23364a <=( A168  and  a23363a );
 a23365a <=( a23364a  and  a23359a );
 a23369a <=( (not A267)  and  A202 );
 a23370a <=( A201  and  a23369a );
 a23374a <=( (not A299)  and  (not A298) );
 a23375a <=( (not A269)  and  a23374a );
 a23376a <=( a23375a  and  a23370a );
 a23379a <=( (not A169)  and  (not A170) );
 a23383a <=( A200  and  (not A199) );
 a23384a <=( A168  and  a23383a );
 a23385a <=( a23384a  and  a23379a );
 a23389a <=( A265  and  A202 );
 a23390a <=( A201  and  a23389a );
 a23394a <=( A301  and  (not A300) );
 a23395a <=( A266  and  a23394a );
 a23396a <=( a23395a  and  a23390a );
 a23399a <=( (not A169)  and  (not A170) );
 a23403a <=( A200  and  (not A199) );
 a23404a <=( A168  and  a23403a );
 a23405a <=( a23404a  and  a23399a );
 a23409a <=( A265  and  A202 );
 a23410a <=( A201  and  a23409a );
 a23414a <=( (not A302)  and  (not A300) );
 a23415a <=( A266  and  a23414a );
 a23416a <=( a23415a  and  a23410a );
 a23419a <=( (not A169)  and  (not A170) );
 a23423a <=( A200  and  (not A199) );
 a23424a <=( A168  and  a23423a );
 a23425a <=( a23424a  and  a23419a );
 a23429a <=( A265  and  A202 );
 a23430a <=( A201  and  a23429a );
 a23434a <=( A299  and  A298 );
 a23435a <=( A266  and  a23434a );
 a23436a <=( a23435a  and  a23430a );
 a23439a <=( (not A169)  and  (not A170) );
 a23443a <=( A200  and  (not A199) );
 a23444a <=( A168  and  a23443a );
 a23445a <=( a23444a  and  a23439a );
 a23449a <=( A265  and  A202 );
 a23450a <=( A201  and  a23449a );
 a23454a <=( (not A299)  and  (not A298) );
 a23455a <=( A266  and  a23454a );
 a23456a <=( a23455a  and  a23450a );
 a23459a <=( (not A169)  and  (not A170) );
 a23463a <=( A200  and  (not A199) );
 a23464a <=( A168  and  a23463a );
 a23465a <=( a23464a  and  a23459a );
 a23469a <=( (not A265)  and  A202 );
 a23470a <=( A201  and  a23469a );
 a23474a <=( A301  and  (not A300) );
 a23475a <=( (not A266)  and  a23474a );
 a23476a <=( a23475a  and  a23470a );
 a23479a <=( (not A169)  and  (not A170) );
 a23483a <=( A200  and  (not A199) );
 a23484a <=( A168  and  a23483a );
 a23485a <=( a23484a  and  a23479a );
 a23489a <=( (not A265)  and  A202 );
 a23490a <=( A201  and  a23489a );
 a23494a <=( (not A302)  and  (not A300) );
 a23495a <=( (not A266)  and  a23494a );
 a23496a <=( a23495a  and  a23490a );
 a23499a <=( (not A169)  and  (not A170) );
 a23503a <=( A200  and  (not A199) );
 a23504a <=( A168  and  a23503a );
 a23505a <=( a23504a  and  a23499a );
 a23509a <=( (not A265)  and  A202 );
 a23510a <=( A201  and  a23509a );
 a23514a <=( A299  and  A298 );
 a23515a <=( (not A266)  and  a23514a );
 a23516a <=( a23515a  and  a23510a );
 a23519a <=( (not A169)  and  (not A170) );
 a23523a <=( A200  and  (not A199) );
 a23524a <=( A168  and  a23523a );
 a23525a <=( a23524a  and  a23519a );
 a23529a <=( (not A265)  and  A202 );
 a23530a <=( A201  and  a23529a );
 a23534a <=( (not A299)  and  (not A298) );
 a23535a <=( (not A266)  and  a23534a );
 a23536a <=( a23535a  and  a23530a );
 a23539a <=( (not A169)  and  (not A170) );
 a23543a <=( A200  and  (not A199) );
 a23544a <=( A168  and  a23543a );
 a23545a <=( a23544a  and  a23539a );
 a23549a <=( (not A267)  and  (not A203) );
 a23550a <=( A201  and  a23549a );
 a23554a <=( A301  and  (not A300) );
 a23555a <=( A268  and  a23554a );
 a23556a <=( a23555a  and  a23550a );
 a23559a <=( (not A169)  and  (not A170) );
 a23563a <=( A200  and  (not A199) );
 a23564a <=( A168  and  a23563a );
 a23565a <=( a23564a  and  a23559a );
 a23569a <=( (not A267)  and  (not A203) );
 a23570a <=( A201  and  a23569a );
 a23574a <=( (not A302)  and  (not A300) );
 a23575a <=( A268  and  a23574a );
 a23576a <=( a23575a  and  a23570a );
 a23579a <=( (not A169)  and  (not A170) );
 a23583a <=( A200  and  (not A199) );
 a23584a <=( A168  and  a23583a );
 a23585a <=( a23584a  and  a23579a );
 a23589a <=( (not A267)  and  (not A203) );
 a23590a <=( A201  and  a23589a );
 a23594a <=( A299  and  A298 );
 a23595a <=( A268  and  a23594a );
 a23596a <=( a23595a  and  a23590a );
 a23599a <=( (not A169)  and  (not A170) );
 a23603a <=( A200  and  (not A199) );
 a23604a <=( A168  and  a23603a );
 a23605a <=( a23604a  and  a23599a );
 a23609a <=( (not A267)  and  (not A203) );
 a23610a <=( A201  and  a23609a );
 a23614a <=( (not A299)  and  (not A298) );
 a23615a <=( A268  and  a23614a );
 a23616a <=( a23615a  and  a23610a );
 a23619a <=( (not A169)  and  (not A170) );
 a23623a <=( A200  and  (not A199) );
 a23624a <=( A168  and  a23623a );
 a23625a <=( a23624a  and  a23619a );
 a23629a <=( (not A267)  and  (not A203) );
 a23630a <=( A201  and  a23629a );
 a23634a <=( A301  and  (not A300) );
 a23635a <=( (not A269)  and  a23634a );
 a23636a <=( a23635a  and  a23630a );
 a23639a <=( (not A169)  and  (not A170) );
 a23643a <=( A200  and  (not A199) );
 a23644a <=( A168  and  a23643a );
 a23645a <=( a23644a  and  a23639a );
 a23649a <=( (not A267)  and  (not A203) );
 a23650a <=( A201  and  a23649a );
 a23654a <=( (not A302)  and  (not A300) );
 a23655a <=( (not A269)  and  a23654a );
 a23656a <=( a23655a  and  a23650a );
 a23659a <=( (not A169)  and  (not A170) );
 a23663a <=( A200  and  (not A199) );
 a23664a <=( A168  and  a23663a );
 a23665a <=( a23664a  and  a23659a );
 a23669a <=( (not A267)  and  (not A203) );
 a23670a <=( A201  and  a23669a );
 a23674a <=( A299  and  A298 );
 a23675a <=( (not A269)  and  a23674a );
 a23676a <=( a23675a  and  a23670a );
 a23679a <=( (not A169)  and  (not A170) );
 a23683a <=( A200  and  (not A199) );
 a23684a <=( A168  and  a23683a );
 a23685a <=( a23684a  and  a23679a );
 a23689a <=( (not A267)  and  (not A203) );
 a23690a <=( A201  and  a23689a );
 a23694a <=( (not A299)  and  (not A298) );
 a23695a <=( (not A269)  and  a23694a );
 a23696a <=( a23695a  and  a23690a );
 a23699a <=( (not A169)  and  (not A170) );
 a23703a <=( A200  and  (not A199) );
 a23704a <=( A168  and  a23703a );
 a23705a <=( a23704a  and  a23699a );
 a23709a <=( A265  and  (not A203) );
 a23710a <=( A201  and  a23709a );
 a23714a <=( A301  and  (not A300) );
 a23715a <=( A266  and  a23714a );
 a23716a <=( a23715a  and  a23710a );
 a23719a <=( (not A169)  and  (not A170) );
 a23723a <=( A200  and  (not A199) );
 a23724a <=( A168  and  a23723a );
 a23725a <=( a23724a  and  a23719a );
 a23729a <=( A265  and  (not A203) );
 a23730a <=( A201  and  a23729a );
 a23734a <=( (not A302)  and  (not A300) );
 a23735a <=( A266  and  a23734a );
 a23736a <=( a23735a  and  a23730a );
 a23739a <=( (not A169)  and  (not A170) );
 a23743a <=( A200  and  (not A199) );
 a23744a <=( A168  and  a23743a );
 a23745a <=( a23744a  and  a23739a );
 a23749a <=( A265  and  (not A203) );
 a23750a <=( A201  and  a23749a );
 a23754a <=( A299  and  A298 );
 a23755a <=( A266  and  a23754a );
 a23756a <=( a23755a  and  a23750a );
 a23759a <=( (not A169)  and  (not A170) );
 a23763a <=( A200  and  (not A199) );
 a23764a <=( A168  and  a23763a );
 a23765a <=( a23764a  and  a23759a );
 a23769a <=( A265  and  (not A203) );
 a23770a <=( A201  and  a23769a );
 a23774a <=( (not A299)  and  (not A298) );
 a23775a <=( A266  and  a23774a );
 a23776a <=( a23775a  and  a23770a );
 a23779a <=( (not A169)  and  (not A170) );
 a23783a <=( A200  and  (not A199) );
 a23784a <=( A168  and  a23783a );
 a23785a <=( a23784a  and  a23779a );
 a23789a <=( (not A265)  and  (not A203) );
 a23790a <=( A201  and  a23789a );
 a23794a <=( A301  and  (not A300) );
 a23795a <=( (not A266)  and  a23794a );
 a23796a <=( a23795a  and  a23790a );
 a23799a <=( (not A169)  and  (not A170) );
 a23803a <=( A200  and  (not A199) );
 a23804a <=( A168  and  a23803a );
 a23805a <=( a23804a  and  a23799a );
 a23809a <=( (not A265)  and  (not A203) );
 a23810a <=( A201  and  a23809a );
 a23814a <=( (not A302)  and  (not A300) );
 a23815a <=( (not A266)  and  a23814a );
 a23816a <=( a23815a  and  a23810a );
 a23819a <=( (not A169)  and  (not A170) );
 a23823a <=( A200  and  (not A199) );
 a23824a <=( A168  and  a23823a );
 a23825a <=( a23824a  and  a23819a );
 a23829a <=( (not A265)  and  (not A203) );
 a23830a <=( A201  and  a23829a );
 a23834a <=( A299  and  A298 );
 a23835a <=( (not A266)  and  a23834a );
 a23836a <=( a23835a  and  a23830a );
 a23839a <=( (not A169)  and  (not A170) );
 a23843a <=( A200  and  (not A199) );
 a23844a <=( A168  and  a23843a );
 a23845a <=( a23844a  and  a23839a );
 a23849a <=( (not A265)  and  (not A203) );
 a23850a <=( A201  and  a23849a );
 a23854a <=( (not A299)  and  (not A298) );
 a23855a <=( (not A266)  and  a23854a );
 a23856a <=( a23855a  and  a23850a );
 a23859a <=( (not A169)  and  (not A170) );
 a23863a <=( (not A200)  and  A199 );
 a23864a <=( A168  and  a23863a );
 a23865a <=( a23864a  and  a23859a );
 a23869a <=( (not A267)  and  A202 );
 a23870a <=( A201  and  a23869a );
 a23874a <=( A301  and  (not A300) );
 a23875a <=( A268  and  a23874a );
 a23876a <=( a23875a  and  a23870a );
 a23879a <=( (not A169)  and  (not A170) );
 a23883a <=( (not A200)  and  A199 );
 a23884a <=( A168  and  a23883a );
 a23885a <=( a23884a  and  a23879a );
 a23889a <=( (not A267)  and  A202 );
 a23890a <=( A201  and  a23889a );
 a23894a <=( (not A302)  and  (not A300) );
 a23895a <=( A268  and  a23894a );
 a23896a <=( a23895a  and  a23890a );
 a23899a <=( (not A169)  and  (not A170) );
 a23903a <=( (not A200)  and  A199 );
 a23904a <=( A168  and  a23903a );
 a23905a <=( a23904a  and  a23899a );
 a23909a <=( (not A267)  and  A202 );
 a23910a <=( A201  and  a23909a );
 a23914a <=( A299  and  A298 );
 a23915a <=( A268  and  a23914a );
 a23916a <=( a23915a  and  a23910a );
 a23919a <=( (not A169)  and  (not A170) );
 a23923a <=( (not A200)  and  A199 );
 a23924a <=( A168  and  a23923a );
 a23925a <=( a23924a  and  a23919a );
 a23929a <=( (not A267)  and  A202 );
 a23930a <=( A201  and  a23929a );
 a23934a <=( (not A299)  and  (not A298) );
 a23935a <=( A268  and  a23934a );
 a23936a <=( a23935a  and  a23930a );
 a23939a <=( (not A169)  and  (not A170) );
 a23943a <=( (not A200)  and  A199 );
 a23944a <=( A168  and  a23943a );
 a23945a <=( a23944a  and  a23939a );
 a23949a <=( (not A267)  and  A202 );
 a23950a <=( A201  and  a23949a );
 a23954a <=( A301  and  (not A300) );
 a23955a <=( (not A269)  and  a23954a );
 a23956a <=( a23955a  and  a23950a );
 a23959a <=( (not A169)  and  (not A170) );
 a23963a <=( (not A200)  and  A199 );
 a23964a <=( A168  and  a23963a );
 a23965a <=( a23964a  and  a23959a );
 a23969a <=( (not A267)  and  A202 );
 a23970a <=( A201  and  a23969a );
 a23974a <=( (not A302)  and  (not A300) );
 a23975a <=( (not A269)  and  a23974a );
 a23976a <=( a23975a  and  a23970a );
 a23979a <=( (not A169)  and  (not A170) );
 a23983a <=( (not A200)  and  A199 );
 a23984a <=( A168  and  a23983a );
 a23985a <=( a23984a  and  a23979a );
 a23989a <=( (not A267)  and  A202 );
 a23990a <=( A201  and  a23989a );
 a23994a <=( A299  and  A298 );
 a23995a <=( (not A269)  and  a23994a );
 a23996a <=( a23995a  and  a23990a );
 a23999a <=( (not A169)  and  (not A170) );
 a24003a <=( (not A200)  and  A199 );
 a24004a <=( A168  and  a24003a );
 a24005a <=( a24004a  and  a23999a );
 a24009a <=( (not A267)  and  A202 );
 a24010a <=( A201  and  a24009a );
 a24014a <=( (not A299)  and  (not A298) );
 a24015a <=( (not A269)  and  a24014a );
 a24016a <=( a24015a  and  a24010a );
 a24019a <=( (not A169)  and  (not A170) );
 a24023a <=( (not A200)  and  A199 );
 a24024a <=( A168  and  a24023a );
 a24025a <=( a24024a  and  a24019a );
 a24029a <=( A265  and  A202 );
 a24030a <=( A201  and  a24029a );
 a24034a <=( A301  and  (not A300) );
 a24035a <=( A266  and  a24034a );
 a24036a <=( a24035a  and  a24030a );
 a24039a <=( (not A169)  and  (not A170) );
 a24043a <=( (not A200)  and  A199 );
 a24044a <=( A168  and  a24043a );
 a24045a <=( a24044a  and  a24039a );
 a24049a <=( A265  and  A202 );
 a24050a <=( A201  and  a24049a );
 a24054a <=( (not A302)  and  (not A300) );
 a24055a <=( A266  and  a24054a );
 a24056a <=( a24055a  and  a24050a );
 a24059a <=( (not A169)  and  (not A170) );
 a24063a <=( (not A200)  and  A199 );
 a24064a <=( A168  and  a24063a );
 a24065a <=( a24064a  and  a24059a );
 a24069a <=( A265  and  A202 );
 a24070a <=( A201  and  a24069a );
 a24074a <=( A299  and  A298 );
 a24075a <=( A266  and  a24074a );
 a24076a <=( a24075a  and  a24070a );
 a24079a <=( (not A169)  and  (not A170) );
 a24083a <=( (not A200)  and  A199 );
 a24084a <=( A168  and  a24083a );
 a24085a <=( a24084a  and  a24079a );
 a24089a <=( A265  and  A202 );
 a24090a <=( A201  and  a24089a );
 a24094a <=( (not A299)  and  (not A298) );
 a24095a <=( A266  and  a24094a );
 a24096a <=( a24095a  and  a24090a );
 a24099a <=( (not A169)  and  (not A170) );
 a24103a <=( (not A200)  and  A199 );
 a24104a <=( A168  and  a24103a );
 a24105a <=( a24104a  and  a24099a );
 a24109a <=( (not A265)  and  A202 );
 a24110a <=( A201  and  a24109a );
 a24114a <=( A301  and  (not A300) );
 a24115a <=( (not A266)  and  a24114a );
 a24116a <=( a24115a  and  a24110a );
 a24119a <=( (not A169)  and  (not A170) );
 a24123a <=( (not A200)  and  A199 );
 a24124a <=( A168  and  a24123a );
 a24125a <=( a24124a  and  a24119a );
 a24129a <=( (not A265)  and  A202 );
 a24130a <=( A201  and  a24129a );
 a24134a <=( (not A302)  and  (not A300) );
 a24135a <=( (not A266)  and  a24134a );
 a24136a <=( a24135a  and  a24130a );
 a24139a <=( (not A169)  and  (not A170) );
 a24143a <=( (not A200)  and  A199 );
 a24144a <=( A168  and  a24143a );
 a24145a <=( a24144a  and  a24139a );
 a24149a <=( (not A265)  and  A202 );
 a24150a <=( A201  and  a24149a );
 a24154a <=( A299  and  A298 );
 a24155a <=( (not A266)  and  a24154a );
 a24156a <=( a24155a  and  a24150a );
 a24159a <=( (not A169)  and  (not A170) );
 a24163a <=( (not A200)  and  A199 );
 a24164a <=( A168  and  a24163a );
 a24165a <=( a24164a  and  a24159a );
 a24169a <=( (not A265)  and  A202 );
 a24170a <=( A201  and  a24169a );
 a24174a <=( (not A299)  and  (not A298) );
 a24175a <=( (not A266)  and  a24174a );
 a24176a <=( a24175a  and  a24170a );
 a24179a <=( (not A169)  and  (not A170) );
 a24183a <=( (not A200)  and  A199 );
 a24184a <=( A168  and  a24183a );
 a24185a <=( a24184a  and  a24179a );
 a24189a <=( (not A267)  and  (not A203) );
 a24190a <=( A201  and  a24189a );
 a24194a <=( A301  and  (not A300) );
 a24195a <=( A268  and  a24194a );
 a24196a <=( a24195a  and  a24190a );
 a24199a <=( (not A169)  and  (not A170) );
 a24203a <=( (not A200)  and  A199 );
 a24204a <=( A168  and  a24203a );
 a24205a <=( a24204a  and  a24199a );
 a24209a <=( (not A267)  and  (not A203) );
 a24210a <=( A201  and  a24209a );
 a24214a <=( (not A302)  and  (not A300) );
 a24215a <=( A268  and  a24214a );
 a24216a <=( a24215a  and  a24210a );
 a24219a <=( (not A169)  and  (not A170) );
 a24223a <=( (not A200)  and  A199 );
 a24224a <=( A168  and  a24223a );
 a24225a <=( a24224a  and  a24219a );
 a24229a <=( (not A267)  and  (not A203) );
 a24230a <=( A201  and  a24229a );
 a24234a <=( A299  and  A298 );
 a24235a <=( A268  and  a24234a );
 a24236a <=( a24235a  and  a24230a );
 a24239a <=( (not A169)  and  (not A170) );
 a24243a <=( (not A200)  and  A199 );
 a24244a <=( A168  and  a24243a );
 a24245a <=( a24244a  and  a24239a );
 a24249a <=( (not A267)  and  (not A203) );
 a24250a <=( A201  and  a24249a );
 a24254a <=( (not A299)  and  (not A298) );
 a24255a <=( A268  and  a24254a );
 a24256a <=( a24255a  and  a24250a );
 a24259a <=( (not A169)  and  (not A170) );
 a24263a <=( (not A200)  and  A199 );
 a24264a <=( A168  and  a24263a );
 a24265a <=( a24264a  and  a24259a );
 a24269a <=( (not A267)  and  (not A203) );
 a24270a <=( A201  and  a24269a );
 a24274a <=( A301  and  (not A300) );
 a24275a <=( (not A269)  and  a24274a );
 a24276a <=( a24275a  and  a24270a );
 a24279a <=( (not A169)  and  (not A170) );
 a24283a <=( (not A200)  and  A199 );
 a24284a <=( A168  and  a24283a );
 a24285a <=( a24284a  and  a24279a );
 a24289a <=( (not A267)  and  (not A203) );
 a24290a <=( A201  and  a24289a );
 a24294a <=( (not A302)  and  (not A300) );
 a24295a <=( (not A269)  and  a24294a );
 a24296a <=( a24295a  and  a24290a );
 a24299a <=( (not A169)  and  (not A170) );
 a24303a <=( (not A200)  and  A199 );
 a24304a <=( A168  and  a24303a );
 a24305a <=( a24304a  and  a24299a );
 a24309a <=( (not A267)  and  (not A203) );
 a24310a <=( A201  and  a24309a );
 a24314a <=( A299  and  A298 );
 a24315a <=( (not A269)  and  a24314a );
 a24316a <=( a24315a  and  a24310a );
 a24319a <=( (not A169)  and  (not A170) );
 a24323a <=( (not A200)  and  A199 );
 a24324a <=( A168  and  a24323a );
 a24325a <=( a24324a  and  a24319a );
 a24329a <=( (not A267)  and  (not A203) );
 a24330a <=( A201  and  a24329a );
 a24334a <=( (not A299)  and  (not A298) );
 a24335a <=( (not A269)  and  a24334a );
 a24336a <=( a24335a  and  a24330a );
 a24339a <=( (not A169)  and  (not A170) );
 a24343a <=( (not A200)  and  A199 );
 a24344a <=( A168  and  a24343a );
 a24345a <=( a24344a  and  a24339a );
 a24349a <=( A265  and  (not A203) );
 a24350a <=( A201  and  a24349a );
 a24354a <=( A301  and  (not A300) );
 a24355a <=( A266  and  a24354a );
 a24356a <=( a24355a  and  a24350a );
 a24359a <=( (not A169)  and  (not A170) );
 a24363a <=( (not A200)  and  A199 );
 a24364a <=( A168  and  a24363a );
 a24365a <=( a24364a  and  a24359a );
 a24369a <=( A265  and  (not A203) );
 a24370a <=( A201  and  a24369a );
 a24374a <=( (not A302)  and  (not A300) );
 a24375a <=( A266  and  a24374a );
 a24376a <=( a24375a  and  a24370a );
 a24379a <=( (not A169)  and  (not A170) );
 a24383a <=( (not A200)  and  A199 );
 a24384a <=( A168  and  a24383a );
 a24385a <=( a24384a  and  a24379a );
 a24389a <=( A265  and  (not A203) );
 a24390a <=( A201  and  a24389a );
 a24394a <=( A299  and  A298 );
 a24395a <=( A266  and  a24394a );
 a24396a <=( a24395a  and  a24390a );
 a24399a <=( (not A169)  and  (not A170) );
 a24403a <=( (not A200)  and  A199 );
 a24404a <=( A168  and  a24403a );
 a24405a <=( a24404a  and  a24399a );
 a24409a <=( A265  and  (not A203) );
 a24410a <=( A201  and  a24409a );
 a24414a <=( (not A299)  and  (not A298) );
 a24415a <=( A266  and  a24414a );
 a24416a <=( a24415a  and  a24410a );
 a24419a <=( (not A169)  and  (not A170) );
 a24423a <=( (not A200)  and  A199 );
 a24424a <=( A168  and  a24423a );
 a24425a <=( a24424a  and  a24419a );
 a24429a <=( (not A265)  and  (not A203) );
 a24430a <=( A201  and  a24429a );
 a24434a <=( A301  and  (not A300) );
 a24435a <=( (not A266)  and  a24434a );
 a24436a <=( a24435a  and  a24430a );
 a24439a <=( (not A169)  and  (not A170) );
 a24443a <=( (not A200)  and  A199 );
 a24444a <=( A168  and  a24443a );
 a24445a <=( a24444a  and  a24439a );
 a24449a <=( (not A265)  and  (not A203) );
 a24450a <=( A201  and  a24449a );
 a24454a <=( (not A302)  and  (not A300) );
 a24455a <=( (not A266)  and  a24454a );
 a24456a <=( a24455a  and  a24450a );
 a24459a <=( (not A169)  and  (not A170) );
 a24463a <=( (not A200)  and  A199 );
 a24464a <=( A168  and  a24463a );
 a24465a <=( a24464a  and  a24459a );
 a24469a <=( (not A265)  and  (not A203) );
 a24470a <=( A201  and  a24469a );
 a24474a <=( A299  and  A298 );
 a24475a <=( (not A266)  and  a24474a );
 a24476a <=( a24475a  and  a24470a );
 a24479a <=( (not A169)  and  (not A170) );
 a24483a <=( (not A200)  and  A199 );
 a24484a <=( A168  and  a24483a );
 a24485a <=( a24484a  and  a24479a );
 a24489a <=( (not A265)  and  (not A203) );
 a24490a <=( A201  and  a24489a );
 a24494a <=( (not A299)  and  (not A298) );
 a24495a <=( (not A266)  and  a24494a );
 a24496a <=( a24495a  and  a24490a );
 a24500a <=( A202  and  A200 );
 a24501a <=( (not A199)  and  a24500a );
 a24505a <=( A234  and  A233 );
 a24506a <=( (not A232)  and  a24505a );
 a24507a <=( a24506a  and  a24501a );
 a24511a <=( A266  and  (not A265) );
 a24512a <=( A235  and  a24511a );
 a24516a <=( A269  and  (not A268) );
 a24517a <=( (not A267)  and  a24516a );
 a24518a <=( a24517a  and  a24512a );
 a24522a <=( A202  and  A200 );
 a24523a <=( (not A199)  and  a24522a );
 a24527a <=( A234  and  A233 );
 a24528a <=( (not A232)  and  a24527a );
 a24529a <=( a24528a  and  a24523a );
 a24533a <=( (not A266)  and  A265 );
 a24534a <=( A235  and  a24533a );
 a24538a <=( A269  and  (not A268) );
 a24539a <=( (not A267)  and  a24538a );
 a24540a <=( a24539a  and  a24534a );
 a24544a <=( A202  and  A200 );
 a24545a <=( (not A199)  and  a24544a );
 a24549a <=( A234  and  A233 );
 a24550a <=( (not A232)  and  a24549a );
 a24551a <=( a24550a  and  a24545a );
 a24555a <=( A266  and  (not A265) );
 a24556a <=( (not A236)  and  a24555a );
 a24560a <=( A269  and  (not A268) );
 a24561a <=( (not A267)  and  a24560a );
 a24562a <=( a24561a  and  a24556a );
 a24566a <=( A202  and  A200 );
 a24567a <=( (not A199)  and  a24566a );
 a24571a <=( A234  and  A233 );
 a24572a <=( (not A232)  and  a24571a );
 a24573a <=( a24572a  and  a24567a );
 a24577a <=( (not A266)  and  A265 );
 a24578a <=( (not A236)  and  a24577a );
 a24582a <=( A269  and  (not A268) );
 a24583a <=( (not A267)  and  a24582a );
 a24584a <=( a24583a  and  a24578a );
 a24588a <=( A202  and  A200 );
 a24589a <=( (not A199)  and  a24588a );
 a24593a <=( A234  and  (not A233) );
 a24594a <=( A232  and  a24593a );
 a24595a <=( a24594a  and  a24589a );
 a24599a <=( A266  and  (not A265) );
 a24600a <=( A235  and  a24599a );
 a24604a <=( A269  and  (not A268) );
 a24605a <=( (not A267)  and  a24604a );
 a24606a <=( a24605a  and  a24600a );
 a24610a <=( A202  and  A200 );
 a24611a <=( (not A199)  and  a24610a );
 a24615a <=( A234  and  (not A233) );
 a24616a <=( A232  and  a24615a );
 a24617a <=( a24616a  and  a24611a );
 a24621a <=( (not A266)  and  A265 );
 a24622a <=( A235  and  a24621a );
 a24626a <=( A269  and  (not A268) );
 a24627a <=( (not A267)  and  a24626a );
 a24628a <=( a24627a  and  a24622a );
 a24632a <=( A202  and  A200 );
 a24633a <=( (not A199)  and  a24632a );
 a24637a <=( A234  and  (not A233) );
 a24638a <=( A232  and  a24637a );
 a24639a <=( a24638a  and  a24633a );
 a24643a <=( A266  and  (not A265) );
 a24644a <=( (not A236)  and  a24643a );
 a24648a <=( A269  and  (not A268) );
 a24649a <=( (not A267)  and  a24648a );
 a24650a <=( a24649a  and  a24644a );
 a24654a <=( A202  and  A200 );
 a24655a <=( (not A199)  and  a24654a );
 a24659a <=( A234  and  (not A233) );
 a24660a <=( A232  and  a24659a );
 a24661a <=( a24660a  and  a24655a );
 a24665a <=( (not A266)  and  A265 );
 a24666a <=( (not A236)  and  a24665a );
 a24670a <=( A269  and  (not A268) );
 a24671a <=( (not A267)  and  a24670a );
 a24672a <=( a24671a  and  a24666a );
 a24676a <=( (not A203)  and  A200 );
 a24677a <=( (not A199)  and  a24676a );
 a24681a <=( A234  and  A233 );
 a24682a <=( (not A232)  and  a24681a );
 a24683a <=( a24682a  and  a24677a );
 a24687a <=( A266  and  (not A265) );
 a24688a <=( A235  and  a24687a );
 a24692a <=( A269  and  (not A268) );
 a24693a <=( (not A267)  and  a24692a );
 a24694a <=( a24693a  and  a24688a );
 a24698a <=( (not A203)  and  A200 );
 a24699a <=( (not A199)  and  a24698a );
 a24703a <=( A234  and  A233 );
 a24704a <=( (not A232)  and  a24703a );
 a24705a <=( a24704a  and  a24699a );
 a24709a <=( (not A266)  and  A265 );
 a24710a <=( A235  and  a24709a );
 a24714a <=( A269  and  (not A268) );
 a24715a <=( (not A267)  and  a24714a );
 a24716a <=( a24715a  and  a24710a );
 a24720a <=( (not A203)  and  A200 );
 a24721a <=( (not A199)  and  a24720a );
 a24725a <=( A234  and  A233 );
 a24726a <=( (not A232)  and  a24725a );
 a24727a <=( a24726a  and  a24721a );
 a24731a <=( A266  and  (not A265) );
 a24732a <=( (not A236)  and  a24731a );
 a24736a <=( A269  and  (not A268) );
 a24737a <=( (not A267)  and  a24736a );
 a24738a <=( a24737a  and  a24732a );
 a24742a <=( (not A203)  and  A200 );
 a24743a <=( (not A199)  and  a24742a );
 a24747a <=( A234  and  A233 );
 a24748a <=( (not A232)  and  a24747a );
 a24749a <=( a24748a  and  a24743a );
 a24753a <=( (not A266)  and  A265 );
 a24754a <=( (not A236)  and  a24753a );
 a24758a <=( A269  and  (not A268) );
 a24759a <=( (not A267)  and  a24758a );
 a24760a <=( a24759a  and  a24754a );
 a24764a <=( (not A203)  and  A200 );
 a24765a <=( (not A199)  and  a24764a );
 a24769a <=( A234  and  (not A233) );
 a24770a <=( A232  and  a24769a );
 a24771a <=( a24770a  and  a24765a );
 a24775a <=( A266  and  (not A265) );
 a24776a <=( A235  and  a24775a );
 a24780a <=( A269  and  (not A268) );
 a24781a <=( (not A267)  and  a24780a );
 a24782a <=( a24781a  and  a24776a );
 a24786a <=( (not A203)  and  A200 );
 a24787a <=( (not A199)  and  a24786a );
 a24791a <=( A234  and  (not A233) );
 a24792a <=( A232  and  a24791a );
 a24793a <=( a24792a  and  a24787a );
 a24797a <=( (not A266)  and  A265 );
 a24798a <=( A235  and  a24797a );
 a24802a <=( A269  and  (not A268) );
 a24803a <=( (not A267)  and  a24802a );
 a24804a <=( a24803a  and  a24798a );
 a24808a <=( (not A203)  and  A200 );
 a24809a <=( (not A199)  and  a24808a );
 a24813a <=( A234  and  (not A233) );
 a24814a <=( A232  and  a24813a );
 a24815a <=( a24814a  and  a24809a );
 a24819a <=( A266  and  (not A265) );
 a24820a <=( (not A236)  and  a24819a );
 a24824a <=( A269  and  (not A268) );
 a24825a <=( (not A267)  and  a24824a );
 a24826a <=( a24825a  and  a24820a );
 a24830a <=( (not A203)  and  A200 );
 a24831a <=( (not A199)  and  a24830a );
 a24835a <=( A234  and  (not A233) );
 a24836a <=( A232  and  a24835a );
 a24837a <=( a24836a  and  a24831a );
 a24841a <=( (not A266)  and  A265 );
 a24842a <=( (not A236)  and  a24841a );
 a24846a <=( A269  and  (not A268) );
 a24847a <=( (not A267)  and  a24846a );
 a24848a <=( a24847a  and  a24842a );
 a24852a <=( A202  and  (not A200) );
 a24853a <=( A199  and  a24852a );
 a24857a <=( A234  and  A233 );
 a24858a <=( (not A232)  and  a24857a );
 a24859a <=( a24858a  and  a24853a );
 a24863a <=( A266  and  (not A265) );
 a24864a <=( A235  and  a24863a );
 a24868a <=( A269  and  (not A268) );
 a24869a <=( (not A267)  and  a24868a );
 a24870a <=( a24869a  and  a24864a );
 a24874a <=( A202  and  (not A200) );
 a24875a <=( A199  and  a24874a );
 a24879a <=( A234  and  A233 );
 a24880a <=( (not A232)  and  a24879a );
 a24881a <=( a24880a  and  a24875a );
 a24885a <=( (not A266)  and  A265 );
 a24886a <=( A235  and  a24885a );
 a24890a <=( A269  and  (not A268) );
 a24891a <=( (not A267)  and  a24890a );
 a24892a <=( a24891a  and  a24886a );
 a24896a <=( A202  and  (not A200) );
 a24897a <=( A199  and  a24896a );
 a24901a <=( A234  and  A233 );
 a24902a <=( (not A232)  and  a24901a );
 a24903a <=( a24902a  and  a24897a );
 a24907a <=( A266  and  (not A265) );
 a24908a <=( (not A236)  and  a24907a );
 a24912a <=( A269  and  (not A268) );
 a24913a <=( (not A267)  and  a24912a );
 a24914a <=( a24913a  and  a24908a );
 a24918a <=( A202  and  (not A200) );
 a24919a <=( A199  and  a24918a );
 a24923a <=( A234  and  A233 );
 a24924a <=( (not A232)  and  a24923a );
 a24925a <=( a24924a  and  a24919a );
 a24929a <=( (not A266)  and  A265 );
 a24930a <=( (not A236)  and  a24929a );
 a24934a <=( A269  and  (not A268) );
 a24935a <=( (not A267)  and  a24934a );
 a24936a <=( a24935a  and  a24930a );
 a24940a <=( A202  and  (not A200) );
 a24941a <=( A199  and  a24940a );
 a24945a <=( A234  and  (not A233) );
 a24946a <=( A232  and  a24945a );
 a24947a <=( a24946a  and  a24941a );
 a24951a <=( A266  and  (not A265) );
 a24952a <=( A235  and  a24951a );
 a24956a <=( A269  and  (not A268) );
 a24957a <=( (not A267)  and  a24956a );
 a24958a <=( a24957a  and  a24952a );
 a24962a <=( A202  and  (not A200) );
 a24963a <=( A199  and  a24962a );
 a24967a <=( A234  and  (not A233) );
 a24968a <=( A232  and  a24967a );
 a24969a <=( a24968a  and  a24963a );
 a24973a <=( (not A266)  and  A265 );
 a24974a <=( A235  and  a24973a );
 a24978a <=( A269  and  (not A268) );
 a24979a <=( (not A267)  and  a24978a );
 a24980a <=( a24979a  and  a24974a );
 a24984a <=( A202  and  (not A200) );
 a24985a <=( A199  and  a24984a );
 a24989a <=( A234  and  (not A233) );
 a24990a <=( A232  and  a24989a );
 a24991a <=( a24990a  and  a24985a );
 a24995a <=( A266  and  (not A265) );
 a24996a <=( (not A236)  and  a24995a );
 a25000a <=( A269  and  (not A268) );
 a25001a <=( (not A267)  and  a25000a );
 a25002a <=( a25001a  and  a24996a );
 a25006a <=( A202  and  (not A200) );
 a25007a <=( A199  and  a25006a );
 a25011a <=( A234  and  (not A233) );
 a25012a <=( A232  and  a25011a );
 a25013a <=( a25012a  and  a25007a );
 a25017a <=( (not A266)  and  A265 );
 a25018a <=( (not A236)  and  a25017a );
 a25022a <=( A269  and  (not A268) );
 a25023a <=( (not A267)  and  a25022a );
 a25024a <=( a25023a  and  a25018a );
 a25028a <=( (not A203)  and  (not A200) );
 a25029a <=( A199  and  a25028a );
 a25033a <=( A234  and  A233 );
 a25034a <=( (not A232)  and  a25033a );
 a25035a <=( a25034a  and  a25029a );
 a25039a <=( A266  and  (not A265) );
 a25040a <=( A235  and  a25039a );
 a25044a <=( A269  and  (not A268) );
 a25045a <=( (not A267)  and  a25044a );
 a25046a <=( a25045a  and  a25040a );
 a25050a <=( (not A203)  and  (not A200) );
 a25051a <=( A199  and  a25050a );
 a25055a <=( A234  and  A233 );
 a25056a <=( (not A232)  and  a25055a );
 a25057a <=( a25056a  and  a25051a );
 a25061a <=( (not A266)  and  A265 );
 a25062a <=( A235  and  a25061a );
 a25066a <=( A269  and  (not A268) );
 a25067a <=( (not A267)  and  a25066a );
 a25068a <=( a25067a  and  a25062a );
 a25072a <=( (not A203)  and  (not A200) );
 a25073a <=( A199  and  a25072a );
 a25077a <=( A234  and  A233 );
 a25078a <=( (not A232)  and  a25077a );
 a25079a <=( a25078a  and  a25073a );
 a25083a <=( A266  and  (not A265) );
 a25084a <=( (not A236)  and  a25083a );
 a25088a <=( A269  and  (not A268) );
 a25089a <=( (not A267)  and  a25088a );
 a25090a <=( a25089a  and  a25084a );
 a25094a <=( (not A203)  and  (not A200) );
 a25095a <=( A199  and  a25094a );
 a25099a <=( A234  and  A233 );
 a25100a <=( (not A232)  and  a25099a );
 a25101a <=( a25100a  and  a25095a );
 a25105a <=( (not A266)  and  A265 );
 a25106a <=( (not A236)  and  a25105a );
 a25110a <=( A269  and  (not A268) );
 a25111a <=( (not A267)  and  a25110a );
 a25112a <=( a25111a  and  a25106a );
 a25116a <=( (not A203)  and  (not A200) );
 a25117a <=( A199  and  a25116a );
 a25121a <=( A234  and  (not A233) );
 a25122a <=( A232  and  a25121a );
 a25123a <=( a25122a  and  a25117a );
 a25127a <=( A266  and  (not A265) );
 a25128a <=( A235  and  a25127a );
 a25132a <=( A269  and  (not A268) );
 a25133a <=( (not A267)  and  a25132a );
 a25134a <=( a25133a  and  a25128a );
 a25138a <=( (not A203)  and  (not A200) );
 a25139a <=( A199  and  a25138a );
 a25143a <=( A234  and  (not A233) );
 a25144a <=( A232  and  a25143a );
 a25145a <=( a25144a  and  a25139a );
 a25149a <=( (not A266)  and  A265 );
 a25150a <=( A235  and  a25149a );
 a25154a <=( A269  and  (not A268) );
 a25155a <=( (not A267)  and  a25154a );
 a25156a <=( a25155a  and  a25150a );
 a25160a <=( (not A203)  and  (not A200) );
 a25161a <=( A199  and  a25160a );
 a25165a <=( A234  and  (not A233) );
 a25166a <=( A232  and  a25165a );
 a25167a <=( a25166a  and  a25161a );
 a25171a <=( A266  and  (not A265) );
 a25172a <=( (not A236)  and  a25171a );
 a25176a <=( A269  and  (not A268) );
 a25177a <=( (not A267)  and  a25176a );
 a25178a <=( a25177a  and  a25172a );
 a25182a <=( (not A203)  and  (not A200) );
 a25183a <=( A199  and  a25182a );
 a25187a <=( A234  and  (not A233) );
 a25188a <=( A232  and  a25187a );
 a25189a <=( a25188a  and  a25183a );
 a25193a <=( (not A266)  and  A265 );
 a25194a <=( (not A236)  and  a25193a );
 a25198a <=( A269  and  (not A268) );
 a25199a <=( (not A267)  and  a25198a );
 a25200a <=( a25199a  and  a25194a );
 a25204a <=( (not A232)  and  A166 );
 a25205a <=( A167  and  a25204a );
 a25209a <=( (not A235)  and  (not A234) );
 a25210a <=( A233  and  a25209a );
 a25211a <=( a25210a  and  a25205a );
 a25215a <=( A266  and  (not A265) );
 a25216a <=( A236  and  a25215a );
 a25220a <=( A269  and  (not A268) );
 a25221a <=( (not A267)  and  a25220a );
 a25222a <=( a25221a  and  a25216a );
 a25226a <=( (not A232)  and  A166 );
 a25227a <=( A167  and  a25226a );
 a25231a <=( (not A235)  and  (not A234) );
 a25232a <=( A233  and  a25231a );
 a25233a <=( a25232a  and  a25227a );
 a25237a <=( (not A266)  and  A265 );
 a25238a <=( A236  and  a25237a );
 a25242a <=( A269  and  (not A268) );
 a25243a <=( (not A267)  and  a25242a );
 a25244a <=( a25243a  and  a25238a );
 a25248a <=( A232  and  A166 );
 a25249a <=( A167  and  a25248a );
 a25253a <=( (not A235)  and  (not A234) );
 a25254a <=( (not A233)  and  a25253a );
 a25255a <=( a25254a  and  a25249a );
 a25259a <=( A266  and  (not A265) );
 a25260a <=( A236  and  a25259a );
 a25264a <=( A269  and  (not A268) );
 a25265a <=( (not A267)  and  a25264a );
 a25266a <=( a25265a  and  a25260a );
 a25270a <=( A232  and  A166 );
 a25271a <=( A167  and  a25270a );
 a25275a <=( (not A235)  and  (not A234) );
 a25276a <=( (not A233)  and  a25275a );
 a25277a <=( a25276a  and  a25271a );
 a25281a <=( (not A266)  and  A265 );
 a25282a <=( A236  and  a25281a );
 a25286a <=( A269  and  (not A268) );
 a25287a <=( (not A267)  and  a25286a );
 a25288a <=( a25287a  and  a25282a );
 a25292a <=( (not A199)  and  A166 );
 a25293a <=( A167  and  a25292a );
 a25297a <=( A202  and  A201 );
 a25298a <=( A200  and  a25297a );
 a25299a <=( a25298a  and  a25293a );
 a25303a <=( A269  and  (not A268) );
 a25304a <=( A267  and  a25303a );
 a25308a <=( A302  and  (not A301) );
 a25309a <=( A300  and  a25308a );
 a25310a <=( a25309a  and  a25304a );
 a25314a <=( (not A199)  and  A166 );
 a25315a <=( A167  and  a25314a );
 a25319a <=( (not A203)  and  A201 );
 a25320a <=( A200  and  a25319a );
 a25321a <=( a25320a  and  a25315a );
 a25325a <=( A269  and  (not A268) );
 a25326a <=( A267  and  a25325a );
 a25330a <=( A302  and  (not A301) );
 a25331a <=( A300  and  a25330a );
 a25332a <=( a25331a  and  a25326a );
 a25336a <=( (not A199)  and  A166 );
 a25337a <=( A167  and  a25336a );
 a25341a <=( (not A202)  and  (not A201) );
 a25342a <=( A200  and  a25341a );
 a25343a <=( a25342a  and  a25337a );
 a25347a <=( (not A268)  and  A267 );
 a25348a <=( A203  and  a25347a );
 a25352a <=( A301  and  (not A300) );
 a25353a <=( A269  and  a25352a );
 a25354a <=( a25353a  and  a25348a );
 a25358a <=( (not A199)  and  A166 );
 a25359a <=( A167  and  a25358a );
 a25363a <=( (not A202)  and  (not A201) );
 a25364a <=( A200  and  a25363a );
 a25365a <=( a25364a  and  a25359a );
 a25369a <=( (not A268)  and  A267 );
 a25370a <=( A203  and  a25369a );
 a25374a <=( (not A302)  and  (not A300) );
 a25375a <=( A269  and  a25374a );
 a25376a <=( a25375a  and  a25370a );
 a25380a <=( (not A199)  and  A166 );
 a25381a <=( A167  and  a25380a );
 a25385a <=( (not A202)  and  (not A201) );
 a25386a <=( A200  and  a25385a );
 a25387a <=( a25386a  and  a25381a );
 a25391a <=( (not A268)  and  A267 );
 a25392a <=( A203  and  a25391a );
 a25396a <=( A299  and  A298 );
 a25397a <=( A269  and  a25396a );
 a25398a <=( a25397a  and  a25392a );
 a25402a <=( (not A199)  and  A166 );
 a25403a <=( A167  and  a25402a );
 a25407a <=( (not A202)  and  (not A201) );
 a25408a <=( A200  and  a25407a );
 a25409a <=( a25408a  and  a25403a );
 a25413a <=( (not A268)  and  A267 );
 a25414a <=( A203  and  a25413a );
 a25418a <=( (not A299)  and  (not A298) );
 a25419a <=( A269  and  a25418a );
 a25420a <=( a25419a  and  a25414a );
 a25424a <=( (not A199)  and  A166 );
 a25425a <=( A167  and  a25424a );
 a25429a <=( (not A202)  and  (not A201) );
 a25430a <=( A200  and  a25429a );
 a25431a <=( a25430a  and  a25425a );
 a25435a <=( A268  and  (not A267) );
 a25436a <=( A203  and  a25435a );
 a25440a <=( A302  and  (not A301) );
 a25441a <=( A300  and  a25440a );
 a25442a <=( a25441a  and  a25436a );
 a25446a <=( (not A199)  and  A166 );
 a25447a <=( A167  and  a25446a );
 a25451a <=( (not A202)  and  (not A201) );
 a25452a <=( A200  and  a25451a );
 a25453a <=( a25452a  and  a25447a );
 a25457a <=( (not A269)  and  (not A267) );
 a25458a <=( A203  and  a25457a );
 a25462a <=( A302  and  (not A301) );
 a25463a <=( A300  and  a25462a );
 a25464a <=( a25463a  and  a25458a );
 a25468a <=( (not A199)  and  A166 );
 a25469a <=( A167  and  a25468a );
 a25473a <=( (not A202)  and  (not A201) );
 a25474a <=( A200  and  a25473a );
 a25475a <=( a25474a  and  a25469a );
 a25479a <=( A266  and  A265 );
 a25480a <=( A203  and  a25479a );
 a25484a <=( A302  and  (not A301) );
 a25485a <=( A300  and  a25484a );
 a25486a <=( a25485a  and  a25480a );
 a25490a <=( (not A199)  and  A166 );
 a25491a <=( A167  and  a25490a );
 a25495a <=( (not A202)  and  (not A201) );
 a25496a <=( A200  and  a25495a );
 a25497a <=( a25496a  and  a25491a );
 a25501a <=( (not A266)  and  (not A265) );
 a25502a <=( A203  and  a25501a );
 a25506a <=( A302  and  (not A301) );
 a25507a <=( A300  and  a25506a );
 a25508a <=( a25507a  and  a25502a );
 a25512a <=( A199  and  A166 );
 a25513a <=( A167  and  a25512a );
 a25517a <=( A202  and  A201 );
 a25518a <=( (not A200)  and  a25517a );
 a25519a <=( a25518a  and  a25513a );
 a25523a <=( A269  and  (not A268) );
 a25524a <=( A267  and  a25523a );
 a25528a <=( A302  and  (not A301) );
 a25529a <=( A300  and  a25528a );
 a25530a <=( a25529a  and  a25524a );
 a25534a <=( A199  and  A166 );
 a25535a <=( A167  and  a25534a );
 a25539a <=( (not A203)  and  A201 );
 a25540a <=( (not A200)  and  a25539a );
 a25541a <=( a25540a  and  a25535a );
 a25545a <=( A269  and  (not A268) );
 a25546a <=( A267  and  a25545a );
 a25550a <=( A302  and  (not A301) );
 a25551a <=( A300  and  a25550a );
 a25552a <=( a25551a  and  a25546a );
 a25556a <=( A199  and  A166 );
 a25557a <=( A167  and  a25556a );
 a25561a <=( (not A202)  and  (not A201) );
 a25562a <=( (not A200)  and  a25561a );
 a25563a <=( a25562a  and  a25557a );
 a25567a <=( (not A268)  and  A267 );
 a25568a <=( A203  and  a25567a );
 a25572a <=( A301  and  (not A300) );
 a25573a <=( A269  and  a25572a );
 a25574a <=( a25573a  and  a25568a );
 a25578a <=( A199  and  A166 );
 a25579a <=( A167  and  a25578a );
 a25583a <=( (not A202)  and  (not A201) );
 a25584a <=( (not A200)  and  a25583a );
 a25585a <=( a25584a  and  a25579a );
 a25589a <=( (not A268)  and  A267 );
 a25590a <=( A203  and  a25589a );
 a25594a <=( (not A302)  and  (not A300) );
 a25595a <=( A269  and  a25594a );
 a25596a <=( a25595a  and  a25590a );
 a25600a <=( A199  and  A166 );
 a25601a <=( A167  and  a25600a );
 a25605a <=( (not A202)  and  (not A201) );
 a25606a <=( (not A200)  and  a25605a );
 a25607a <=( a25606a  and  a25601a );
 a25611a <=( (not A268)  and  A267 );
 a25612a <=( A203  and  a25611a );
 a25616a <=( A299  and  A298 );
 a25617a <=( A269  and  a25616a );
 a25618a <=( a25617a  and  a25612a );
 a25622a <=( A199  and  A166 );
 a25623a <=( A167  and  a25622a );
 a25627a <=( (not A202)  and  (not A201) );
 a25628a <=( (not A200)  and  a25627a );
 a25629a <=( a25628a  and  a25623a );
 a25633a <=( (not A268)  and  A267 );
 a25634a <=( A203  and  a25633a );
 a25638a <=( (not A299)  and  (not A298) );
 a25639a <=( A269  and  a25638a );
 a25640a <=( a25639a  and  a25634a );
 a25644a <=( A199  and  A166 );
 a25645a <=( A167  and  a25644a );
 a25649a <=( (not A202)  and  (not A201) );
 a25650a <=( (not A200)  and  a25649a );
 a25651a <=( a25650a  and  a25645a );
 a25655a <=( A268  and  (not A267) );
 a25656a <=( A203  and  a25655a );
 a25660a <=( A302  and  (not A301) );
 a25661a <=( A300  and  a25660a );
 a25662a <=( a25661a  and  a25656a );
 a25666a <=( A199  and  A166 );
 a25667a <=( A167  and  a25666a );
 a25671a <=( (not A202)  and  (not A201) );
 a25672a <=( (not A200)  and  a25671a );
 a25673a <=( a25672a  and  a25667a );
 a25677a <=( (not A269)  and  (not A267) );
 a25678a <=( A203  and  a25677a );
 a25682a <=( A302  and  (not A301) );
 a25683a <=( A300  and  a25682a );
 a25684a <=( a25683a  and  a25678a );
 a25688a <=( A199  and  A166 );
 a25689a <=( A167  and  a25688a );
 a25693a <=( (not A202)  and  (not A201) );
 a25694a <=( (not A200)  and  a25693a );
 a25695a <=( a25694a  and  a25689a );
 a25699a <=( A266  and  A265 );
 a25700a <=( A203  and  a25699a );
 a25704a <=( A302  and  (not A301) );
 a25705a <=( A300  and  a25704a );
 a25706a <=( a25705a  and  a25700a );
 a25710a <=( A199  and  A166 );
 a25711a <=( A167  and  a25710a );
 a25715a <=( (not A202)  and  (not A201) );
 a25716a <=( (not A200)  and  a25715a );
 a25717a <=( a25716a  and  a25711a );
 a25721a <=( (not A266)  and  (not A265) );
 a25722a <=( A203  and  a25721a );
 a25726a <=( A302  and  (not A301) );
 a25727a <=( A300  and  a25726a );
 a25728a <=( a25727a  and  a25722a );
 a25732a <=( (not A232)  and  (not A166) );
 a25733a <=( (not A167)  and  a25732a );
 a25737a <=( (not A235)  and  (not A234) );
 a25738a <=( A233  and  a25737a );
 a25739a <=( a25738a  and  a25733a );
 a25743a <=( A266  and  (not A265) );
 a25744a <=( A236  and  a25743a );
 a25748a <=( A269  and  (not A268) );
 a25749a <=( (not A267)  and  a25748a );
 a25750a <=( a25749a  and  a25744a );
 a25754a <=( (not A232)  and  (not A166) );
 a25755a <=( (not A167)  and  a25754a );
 a25759a <=( (not A235)  and  (not A234) );
 a25760a <=( A233  and  a25759a );
 a25761a <=( a25760a  and  a25755a );
 a25765a <=( (not A266)  and  A265 );
 a25766a <=( A236  and  a25765a );
 a25770a <=( A269  and  (not A268) );
 a25771a <=( (not A267)  and  a25770a );
 a25772a <=( a25771a  and  a25766a );
 a25776a <=( A232  and  (not A166) );
 a25777a <=( (not A167)  and  a25776a );
 a25781a <=( (not A235)  and  (not A234) );
 a25782a <=( (not A233)  and  a25781a );
 a25783a <=( a25782a  and  a25777a );
 a25787a <=( A266  and  (not A265) );
 a25788a <=( A236  and  a25787a );
 a25792a <=( A269  and  (not A268) );
 a25793a <=( (not A267)  and  a25792a );
 a25794a <=( a25793a  and  a25788a );
 a25798a <=( A232  and  (not A166) );
 a25799a <=( (not A167)  and  a25798a );
 a25803a <=( (not A235)  and  (not A234) );
 a25804a <=( (not A233)  and  a25803a );
 a25805a <=( a25804a  and  a25799a );
 a25809a <=( (not A266)  and  A265 );
 a25810a <=( A236  and  a25809a );
 a25814a <=( A269  and  (not A268) );
 a25815a <=( (not A267)  and  a25814a );
 a25816a <=( a25815a  and  a25810a );
 a25820a <=( (not A199)  and  (not A166) );
 a25821a <=( (not A167)  and  a25820a );
 a25825a <=( A202  and  A201 );
 a25826a <=( A200  and  a25825a );
 a25827a <=( a25826a  and  a25821a );
 a25831a <=( A269  and  (not A268) );
 a25832a <=( A267  and  a25831a );
 a25836a <=( A302  and  (not A301) );
 a25837a <=( A300  and  a25836a );
 a25838a <=( a25837a  and  a25832a );
 a25842a <=( (not A199)  and  (not A166) );
 a25843a <=( (not A167)  and  a25842a );
 a25847a <=( (not A203)  and  A201 );
 a25848a <=( A200  and  a25847a );
 a25849a <=( a25848a  and  a25843a );
 a25853a <=( A269  and  (not A268) );
 a25854a <=( A267  and  a25853a );
 a25858a <=( A302  and  (not A301) );
 a25859a <=( A300  and  a25858a );
 a25860a <=( a25859a  and  a25854a );
 a25864a <=( (not A199)  and  (not A166) );
 a25865a <=( (not A167)  and  a25864a );
 a25869a <=( (not A202)  and  (not A201) );
 a25870a <=( A200  and  a25869a );
 a25871a <=( a25870a  and  a25865a );
 a25875a <=( (not A268)  and  A267 );
 a25876a <=( A203  and  a25875a );
 a25880a <=( A301  and  (not A300) );
 a25881a <=( A269  and  a25880a );
 a25882a <=( a25881a  and  a25876a );
 a25886a <=( (not A199)  and  (not A166) );
 a25887a <=( (not A167)  and  a25886a );
 a25891a <=( (not A202)  and  (not A201) );
 a25892a <=( A200  and  a25891a );
 a25893a <=( a25892a  and  a25887a );
 a25897a <=( (not A268)  and  A267 );
 a25898a <=( A203  and  a25897a );
 a25902a <=( (not A302)  and  (not A300) );
 a25903a <=( A269  and  a25902a );
 a25904a <=( a25903a  and  a25898a );
 a25908a <=( (not A199)  and  (not A166) );
 a25909a <=( (not A167)  and  a25908a );
 a25913a <=( (not A202)  and  (not A201) );
 a25914a <=( A200  and  a25913a );
 a25915a <=( a25914a  and  a25909a );
 a25919a <=( (not A268)  and  A267 );
 a25920a <=( A203  and  a25919a );
 a25924a <=( A299  and  A298 );
 a25925a <=( A269  and  a25924a );
 a25926a <=( a25925a  and  a25920a );
 a25930a <=( (not A199)  and  (not A166) );
 a25931a <=( (not A167)  and  a25930a );
 a25935a <=( (not A202)  and  (not A201) );
 a25936a <=( A200  and  a25935a );
 a25937a <=( a25936a  and  a25931a );
 a25941a <=( (not A268)  and  A267 );
 a25942a <=( A203  and  a25941a );
 a25946a <=( (not A299)  and  (not A298) );
 a25947a <=( A269  and  a25946a );
 a25948a <=( a25947a  and  a25942a );
 a25952a <=( (not A199)  and  (not A166) );
 a25953a <=( (not A167)  and  a25952a );
 a25957a <=( (not A202)  and  (not A201) );
 a25958a <=( A200  and  a25957a );
 a25959a <=( a25958a  and  a25953a );
 a25963a <=( A268  and  (not A267) );
 a25964a <=( A203  and  a25963a );
 a25968a <=( A302  and  (not A301) );
 a25969a <=( A300  and  a25968a );
 a25970a <=( a25969a  and  a25964a );
 a25974a <=( (not A199)  and  (not A166) );
 a25975a <=( (not A167)  and  a25974a );
 a25979a <=( (not A202)  and  (not A201) );
 a25980a <=( A200  and  a25979a );
 a25981a <=( a25980a  and  a25975a );
 a25985a <=( (not A269)  and  (not A267) );
 a25986a <=( A203  and  a25985a );
 a25990a <=( A302  and  (not A301) );
 a25991a <=( A300  and  a25990a );
 a25992a <=( a25991a  and  a25986a );
 a25996a <=( (not A199)  and  (not A166) );
 a25997a <=( (not A167)  and  a25996a );
 a26001a <=( (not A202)  and  (not A201) );
 a26002a <=( A200  and  a26001a );
 a26003a <=( a26002a  and  a25997a );
 a26007a <=( A266  and  A265 );
 a26008a <=( A203  and  a26007a );
 a26012a <=( A302  and  (not A301) );
 a26013a <=( A300  and  a26012a );
 a26014a <=( a26013a  and  a26008a );
 a26018a <=( (not A199)  and  (not A166) );
 a26019a <=( (not A167)  and  a26018a );
 a26023a <=( (not A202)  and  (not A201) );
 a26024a <=( A200  and  a26023a );
 a26025a <=( a26024a  and  a26019a );
 a26029a <=( (not A266)  and  (not A265) );
 a26030a <=( A203  and  a26029a );
 a26034a <=( A302  and  (not A301) );
 a26035a <=( A300  and  a26034a );
 a26036a <=( a26035a  and  a26030a );
 a26040a <=( A199  and  (not A166) );
 a26041a <=( (not A167)  and  a26040a );
 a26045a <=( A202  and  A201 );
 a26046a <=( (not A200)  and  a26045a );
 a26047a <=( a26046a  and  a26041a );
 a26051a <=( A269  and  (not A268) );
 a26052a <=( A267  and  a26051a );
 a26056a <=( A302  and  (not A301) );
 a26057a <=( A300  and  a26056a );
 a26058a <=( a26057a  and  a26052a );
 a26062a <=( A199  and  (not A166) );
 a26063a <=( (not A167)  and  a26062a );
 a26067a <=( (not A203)  and  A201 );
 a26068a <=( (not A200)  and  a26067a );
 a26069a <=( a26068a  and  a26063a );
 a26073a <=( A269  and  (not A268) );
 a26074a <=( A267  and  a26073a );
 a26078a <=( A302  and  (not A301) );
 a26079a <=( A300  and  a26078a );
 a26080a <=( a26079a  and  a26074a );
 a26084a <=( A199  and  (not A166) );
 a26085a <=( (not A167)  and  a26084a );
 a26089a <=( (not A202)  and  (not A201) );
 a26090a <=( (not A200)  and  a26089a );
 a26091a <=( a26090a  and  a26085a );
 a26095a <=( (not A268)  and  A267 );
 a26096a <=( A203  and  a26095a );
 a26100a <=( A301  and  (not A300) );
 a26101a <=( A269  and  a26100a );
 a26102a <=( a26101a  and  a26096a );
 a26106a <=( A199  and  (not A166) );
 a26107a <=( (not A167)  and  a26106a );
 a26111a <=( (not A202)  and  (not A201) );
 a26112a <=( (not A200)  and  a26111a );
 a26113a <=( a26112a  and  a26107a );
 a26117a <=( (not A268)  and  A267 );
 a26118a <=( A203  and  a26117a );
 a26122a <=( (not A302)  and  (not A300) );
 a26123a <=( A269  and  a26122a );
 a26124a <=( a26123a  and  a26118a );
 a26128a <=( A199  and  (not A166) );
 a26129a <=( (not A167)  and  a26128a );
 a26133a <=( (not A202)  and  (not A201) );
 a26134a <=( (not A200)  and  a26133a );
 a26135a <=( a26134a  and  a26129a );
 a26139a <=( (not A268)  and  A267 );
 a26140a <=( A203  and  a26139a );
 a26144a <=( A299  and  A298 );
 a26145a <=( A269  and  a26144a );
 a26146a <=( a26145a  and  a26140a );
 a26150a <=( A199  and  (not A166) );
 a26151a <=( (not A167)  and  a26150a );
 a26155a <=( (not A202)  and  (not A201) );
 a26156a <=( (not A200)  and  a26155a );
 a26157a <=( a26156a  and  a26151a );
 a26161a <=( (not A268)  and  A267 );
 a26162a <=( A203  and  a26161a );
 a26166a <=( (not A299)  and  (not A298) );
 a26167a <=( A269  and  a26166a );
 a26168a <=( a26167a  and  a26162a );
 a26172a <=( A199  and  (not A166) );
 a26173a <=( (not A167)  and  a26172a );
 a26177a <=( (not A202)  and  (not A201) );
 a26178a <=( (not A200)  and  a26177a );
 a26179a <=( a26178a  and  a26173a );
 a26183a <=( A268  and  (not A267) );
 a26184a <=( A203  and  a26183a );
 a26188a <=( A302  and  (not A301) );
 a26189a <=( A300  and  a26188a );
 a26190a <=( a26189a  and  a26184a );
 a26194a <=( A199  and  (not A166) );
 a26195a <=( (not A167)  and  a26194a );
 a26199a <=( (not A202)  and  (not A201) );
 a26200a <=( (not A200)  and  a26199a );
 a26201a <=( a26200a  and  a26195a );
 a26205a <=( (not A269)  and  (not A267) );
 a26206a <=( A203  and  a26205a );
 a26210a <=( A302  and  (not A301) );
 a26211a <=( A300  and  a26210a );
 a26212a <=( a26211a  and  a26206a );
 a26216a <=( A199  and  (not A166) );
 a26217a <=( (not A167)  and  a26216a );
 a26221a <=( (not A202)  and  (not A201) );
 a26222a <=( (not A200)  and  a26221a );
 a26223a <=( a26222a  and  a26217a );
 a26227a <=( A266  and  A265 );
 a26228a <=( A203  and  a26227a );
 a26232a <=( A302  and  (not A301) );
 a26233a <=( A300  and  a26232a );
 a26234a <=( a26233a  and  a26228a );
 a26238a <=( A199  and  (not A166) );
 a26239a <=( (not A167)  and  a26238a );
 a26243a <=( (not A202)  and  (not A201) );
 a26244a <=( (not A200)  and  a26243a );
 a26245a <=( a26244a  and  a26239a );
 a26249a <=( (not A266)  and  (not A265) );
 a26250a <=( A203  and  a26249a );
 a26254a <=( A302  and  (not A301) );
 a26255a <=( A300  and  a26254a );
 a26256a <=( a26255a  and  a26250a );
 a26260a <=( A200  and  (not A199) );
 a26261a <=( A170  and  a26260a );
 a26265a <=( A234  and  A233 );
 a26266a <=( (not A232)  and  a26265a );
 a26267a <=( a26266a  and  a26261a );
 a26271a <=( A266  and  (not A265) );
 a26272a <=( A235  and  a26271a );
 a26276a <=( A269  and  (not A268) );
 a26277a <=( (not A267)  and  a26276a );
 a26278a <=( a26277a  and  a26272a );
 a26282a <=( A200  and  (not A199) );
 a26283a <=( A170  and  a26282a );
 a26287a <=( A234  and  A233 );
 a26288a <=( (not A232)  and  a26287a );
 a26289a <=( a26288a  and  a26283a );
 a26293a <=( (not A266)  and  A265 );
 a26294a <=( A235  and  a26293a );
 a26298a <=( A269  and  (not A268) );
 a26299a <=( (not A267)  and  a26298a );
 a26300a <=( a26299a  and  a26294a );
 a26304a <=( A200  and  (not A199) );
 a26305a <=( A170  and  a26304a );
 a26309a <=( A234  and  A233 );
 a26310a <=( (not A232)  and  a26309a );
 a26311a <=( a26310a  and  a26305a );
 a26315a <=( A266  and  (not A265) );
 a26316a <=( (not A236)  and  a26315a );
 a26320a <=( A269  and  (not A268) );
 a26321a <=( (not A267)  and  a26320a );
 a26322a <=( a26321a  and  a26316a );
 a26326a <=( A200  and  (not A199) );
 a26327a <=( A170  and  a26326a );
 a26331a <=( A234  and  A233 );
 a26332a <=( (not A232)  and  a26331a );
 a26333a <=( a26332a  and  a26327a );
 a26337a <=( (not A266)  and  A265 );
 a26338a <=( (not A236)  and  a26337a );
 a26342a <=( A269  and  (not A268) );
 a26343a <=( (not A267)  and  a26342a );
 a26344a <=( a26343a  and  a26338a );
 a26348a <=( A200  and  (not A199) );
 a26349a <=( A170  and  a26348a );
 a26353a <=( A234  and  (not A233) );
 a26354a <=( A232  and  a26353a );
 a26355a <=( a26354a  and  a26349a );
 a26359a <=( A266  and  (not A265) );
 a26360a <=( A235  and  a26359a );
 a26364a <=( A269  and  (not A268) );
 a26365a <=( (not A267)  and  a26364a );
 a26366a <=( a26365a  and  a26360a );
 a26370a <=( A200  and  (not A199) );
 a26371a <=( A170  and  a26370a );
 a26375a <=( A234  and  (not A233) );
 a26376a <=( A232  and  a26375a );
 a26377a <=( a26376a  and  a26371a );
 a26381a <=( (not A266)  and  A265 );
 a26382a <=( A235  and  a26381a );
 a26386a <=( A269  and  (not A268) );
 a26387a <=( (not A267)  and  a26386a );
 a26388a <=( a26387a  and  a26382a );
 a26392a <=( A200  and  (not A199) );
 a26393a <=( A170  and  a26392a );
 a26397a <=( A234  and  (not A233) );
 a26398a <=( A232  and  a26397a );
 a26399a <=( a26398a  and  a26393a );
 a26403a <=( A266  and  (not A265) );
 a26404a <=( (not A236)  and  a26403a );
 a26408a <=( A269  and  (not A268) );
 a26409a <=( (not A267)  and  a26408a );
 a26410a <=( a26409a  and  a26404a );
 a26414a <=( A200  and  (not A199) );
 a26415a <=( A170  and  a26414a );
 a26419a <=( A234  and  (not A233) );
 a26420a <=( A232  and  a26419a );
 a26421a <=( a26420a  and  a26415a );
 a26425a <=( (not A266)  and  A265 );
 a26426a <=( (not A236)  and  a26425a );
 a26430a <=( A269  and  (not A268) );
 a26431a <=( (not A267)  and  a26430a );
 a26432a <=( a26431a  and  a26426a );
 a26436a <=( (not A200)  and  A199 );
 a26437a <=( A170  and  a26436a );
 a26441a <=( A234  and  A233 );
 a26442a <=( (not A232)  and  a26441a );
 a26443a <=( a26442a  and  a26437a );
 a26447a <=( A266  and  (not A265) );
 a26448a <=( A235  and  a26447a );
 a26452a <=( A269  and  (not A268) );
 a26453a <=( (not A267)  and  a26452a );
 a26454a <=( a26453a  and  a26448a );
 a26458a <=( (not A200)  and  A199 );
 a26459a <=( A170  and  a26458a );
 a26463a <=( A234  and  A233 );
 a26464a <=( (not A232)  and  a26463a );
 a26465a <=( a26464a  and  a26459a );
 a26469a <=( (not A266)  and  A265 );
 a26470a <=( A235  and  a26469a );
 a26474a <=( A269  and  (not A268) );
 a26475a <=( (not A267)  and  a26474a );
 a26476a <=( a26475a  and  a26470a );
 a26480a <=( (not A200)  and  A199 );
 a26481a <=( A170  and  a26480a );
 a26485a <=( A234  and  A233 );
 a26486a <=( (not A232)  and  a26485a );
 a26487a <=( a26486a  and  a26481a );
 a26491a <=( A266  and  (not A265) );
 a26492a <=( (not A236)  and  a26491a );
 a26496a <=( A269  and  (not A268) );
 a26497a <=( (not A267)  and  a26496a );
 a26498a <=( a26497a  and  a26492a );
 a26502a <=( (not A200)  and  A199 );
 a26503a <=( A170  and  a26502a );
 a26507a <=( A234  and  A233 );
 a26508a <=( (not A232)  and  a26507a );
 a26509a <=( a26508a  and  a26503a );
 a26513a <=( (not A266)  and  A265 );
 a26514a <=( (not A236)  and  a26513a );
 a26518a <=( A269  and  (not A268) );
 a26519a <=( (not A267)  and  a26518a );
 a26520a <=( a26519a  and  a26514a );
 a26524a <=( (not A200)  and  A199 );
 a26525a <=( A170  and  a26524a );
 a26529a <=( A234  and  (not A233) );
 a26530a <=( A232  and  a26529a );
 a26531a <=( a26530a  and  a26525a );
 a26535a <=( A266  and  (not A265) );
 a26536a <=( A235  and  a26535a );
 a26540a <=( A269  and  (not A268) );
 a26541a <=( (not A267)  and  a26540a );
 a26542a <=( a26541a  and  a26536a );
 a26546a <=( (not A200)  and  A199 );
 a26547a <=( A170  and  a26546a );
 a26551a <=( A234  and  (not A233) );
 a26552a <=( A232  and  a26551a );
 a26553a <=( a26552a  and  a26547a );
 a26557a <=( (not A266)  and  A265 );
 a26558a <=( A235  and  a26557a );
 a26562a <=( A269  and  (not A268) );
 a26563a <=( (not A267)  and  a26562a );
 a26564a <=( a26563a  and  a26558a );
 a26568a <=( (not A200)  and  A199 );
 a26569a <=( A170  and  a26568a );
 a26573a <=( A234  and  (not A233) );
 a26574a <=( A232  and  a26573a );
 a26575a <=( a26574a  and  a26569a );
 a26579a <=( A266  and  (not A265) );
 a26580a <=( (not A236)  and  a26579a );
 a26584a <=( A269  and  (not A268) );
 a26585a <=( (not A267)  and  a26584a );
 a26586a <=( a26585a  and  a26580a );
 a26590a <=( (not A200)  and  A199 );
 a26591a <=( A170  and  a26590a );
 a26595a <=( A234  and  (not A233) );
 a26596a <=( A232  and  a26595a );
 a26597a <=( a26596a  and  a26591a );
 a26601a <=( (not A266)  and  A265 );
 a26602a <=( (not A236)  and  a26601a );
 a26606a <=( A269  and  (not A268) );
 a26607a <=( (not A267)  and  a26606a );
 a26608a <=( a26607a  and  a26602a );
 a26612a <=( A167  and  A168 );
 a26613a <=( A170  and  a26612a );
 a26617a <=( A202  and  (not A201) );
 a26618a <=( (not A166)  and  a26617a );
 a26619a <=( a26618a  and  a26613a );
 a26623a <=( A298  and  A268 );
 a26624a <=( (not A267)  and  a26623a );
 a26628a <=( A301  and  A300 );
 a26629a <=( (not A299)  and  a26628a );
 a26630a <=( a26629a  and  a26624a );
 a26634a <=( A167  and  A168 );
 a26635a <=( A170  and  a26634a );
 a26639a <=( A202  and  (not A201) );
 a26640a <=( (not A166)  and  a26639a );
 a26641a <=( a26640a  and  a26635a );
 a26645a <=( A298  and  A268 );
 a26646a <=( (not A267)  and  a26645a );
 a26650a <=( (not A302)  and  A300 );
 a26651a <=( (not A299)  and  a26650a );
 a26652a <=( a26651a  and  a26646a );
 a26656a <=( A167  and  A168 );
 a26657a <=( A170  and  a26656a );
 a26661a <=( A202  and  (not A201) );
 a26662a <=( (not A166)  and  a26661a );
 a26663a <=( a26662a  and  a26657a );
 a26667a <=( (not A298)  and  A268 );
 a26668a <=( (not A267)  and  a26667a );
 a26672a <=( A301  and  A300 );
 a26673a <=( A299  and  a26672a );
 a26674a <=( a26673a  and  a26668a );
 a26678a <=( A167  and  A168 );
 a26679a <=( A170  and  a26678a );
 a26683a <=( A202  and  (not A201) );
 a26684a <=( (not A166)  and  a26683a );
 a26685a <=( a26684a  and  a26679a );
 a26689a <=( (not A298)  and  A268 );
 a26690a <=( (not A267)  and  a26689a );
 a26694a <=( (not A302)  and  A300 );
 a26695a <=( A299  and  a26694a );
 a26696a <=( a26695a  and  a26690a );
 a26700a <=( A167  and  A168 );
 a26701a <=( A170  and  a26700a );
 a26705a <=( A202  and  (not A201) );
 a26706a <=( (not A166)  and  a26705a );
 a26707a <=( a26706a  and  a26701a );
 a26711a <=( A298  and  (not A269) );
 a26712a <=( (not A267)  and  a26711a );
 a26716a <=( A301  and  A300 );
 a26717a <=( (not A299)  and  a26716a );
 a26718a <=( a26717a  and  a26712a );
 a26722a <=( A167  and  A168 );
 a26723a <=( A170  and  a26722a );
 a26727a <=( A202  and  (not A201) );
 a26728a <=( (not A166)  and  a26727a );
 a26729a <=( a26728a  and  a26723a );
 a26733a <=( A298  and  (not A269) );
 a26734a <=( (not A267)  and  a26733a );
 a26738a <=( (not A302)  and  A300 );
 a26739a <=( (not A299)  and  a26738a );
 a26740a <=( a26739a  and  a26734a );
 a26744a <=( A167  and  A168 );
 a26745a <=( A170  and  a26744a );
 a26749a <=( A202  and  (not A201) );
 a26750a <=( (not A166)  and  a26749a );
 a26751a <=( a26750a  and  a26745a );
 a26755a <=( (not A298)  and  (not A269) );
 a26756a <=( (not A267)  and  a26755a );
 a26760a <=( A301  and  A300 );
 a26761a <=( A299  and  a26760a );
 a26762a <=( a26761a  and  a26756a );
 a26766a <=( A167  and  A168 );
 a26767a <=( A170  and  a26766a );
 a26771a <=( A202  and  (not A201) );
 a26772a <=( (not A166)  and  a26771a );
 a26773a <=( a26772a  and  a26767a );
 a26777a <=( (not A298)  and  (not A269) );
 a26778a <=( (not A267)  and  a26777a );
 a26782a <=( (not A302)  and  A300 );
 a26783a <=( A299  and  a26782a );
 a26784a <=( a26783a  and  a26778a );
 a26788a <=( A167  and  A168 );
 a26789a <=( A170  and  a26788a );
 a26793a <=( A202  and  (not A201) );
 a26794a <=( (not A166)  and  a26793a );
 a26795a <=( a26794a  and  a26789a );
 a26799a <=( A298  and  A266 );
 a26800a <=( A265  and  a26799a );
 a26804a <=( A301  and  A300 );
 a26805a <=( (not A299)  and  a26804a );
 a26806a <=( a26805a  and  a26800a );
 a26810a <=( A167  and  A168 );
 a26811a <=( A170  and  a26810a );
 a26815a <=( A202  and  (not A201) );
 a26816a <=( (not A166)  and  a26815a );
 a26817a <=( a26816a  and  a26811a );
 a26821a <=( A298  and  A266 );
 a26822a <=( A265  and  a26821a );
 a26826a <=( (not A302)  and  A300 );
 a26827a <=( (not A299)  and  a26826a );
 a26828a <=( a26827a  and  a26822a );
 a26832a <=( A167  and  A168 );
 a26833a <=( A170  and  a26832a );
 a26837a <=( A202  and  (not A201) );
 a26838a <=( (not A166)  and  a26837a );
 a26839a <=( a26838a  and  a26833a );
 a26843a <=( (not A298)  and  A266 );
 a26844a <=( A265  and  a26843a );
 a26848a <=( A301  and  A300 );
 a26849a <=( A299  and  a26848a );
 a26850a <=( a26849a  and  a26844a );
 a26854a <=( A167  and  A168 );
 a26855a <=( A170  and  a26854a );
 a26859a <=( A202  and  (not A201) );
 a26860a <=( (not A166)  and  a26859a );
 a26861a <=( a26860a  and  a26855a );
 a26865a <=( (not A298)  and  A266 );
 a26866a <=( A265  and  a26865a );
 a26870a <=( (not A302)  and  A300 );
 a26871a <=( A299  and  a26870a );
 a26872a <=( a26871a  and  a26866a );
 a26876a <=( A167  and  A168 );
 a26877a <=( A170  and  a26876a );
 a26881a <=( A202  and  (not A201) );
 a26882a <=( (not A166)  and  a26881a );
 a26883a <=( a26882a  and  a26877a );
 a26887a <=( A267  and  A266 );
 a26888a <=( (not A265)  and  a26887a );
 a26892a <=( A301  and  (not A300) );
 a26893a <=( A268  and  a26892a );
 a26894a <=( a26893a  and  a26888a );
 a26898a <=( A167  and  A168 );
 a26899a <=( A170  and  a26898a );
 a26903a <=( A202  and  (not A201) );
 a26904a <=( (not A166)  and  a26903a );
 a26905a <=( a26904a  and  a26899a );
 a26909a <=( A267  and  A266 );
 a26910a <=( (not A265)  and  a26909a );
 a26914a <=( (not A302)  and  (not A300) );
 a26915a <=( A268  and  a26914a );
 a26916a <=( a26915a  and  a26910a );
 a26920a <=( A167  and  A168 );
 a26921a <=( A170  and  a26920a );
 a26925a <=( A202  and  (not A201) );
 a26926a <=( (not A166)  and  a26925a );
 a26927a <=( a26926a  and  a26921a );
 a26931a <=( A267  and  A266 );
 a26932a <=( (not A265)  and  a26931a );
 a26936a <=( A299  and  A298 );
 a26937a <=( A268  and  a26936a );
 a26938a <=( a26937a  and  a26932a );
 a26942a <=( A167  and  A168 );
 a26943a <=( A170  and  a26942a );
 a26947a <=( A202  and  (not A201) );
 a26948a <=( (not A166)  and  a26947a );
 a26949a <=( a26948a  and  a26943a );
 a26953a <=( A267  and  A266 );
 a26954a <=( (not A265)  and  a26953a );
 a26958a <=( (not A299)  and  (not A298) );
 a26959a <=( A268  and  a26958a );
 a26960a <=( a26959a  and  a26954a );
 a26964a <=( A167  and  A168 );
 a26965a <=( A170  and  a26964a );
 a26969a <=( A202  and  (not A201) );
 a26970a <=( (not A166)  and  a26969a );
 a26971a <=( a26970a  and  a26965a );
 a26975a <=( A267  and  A266 );
 a26976a <=( (not A265)  and  a26975a );
 a26980a <=( A301  and  (not A300) );
 a26981a <=( (not A269)  and  a26980a );
 a26982a <=( a26981a  and  a26976a );
 a26986a <=( A167  and  A168 );
 a26987a <=( A170  and  a26986a );
 a26991a <=( A202  and  (not A201) );
 a26992a <=( (not A166)  and  a26991a );
 a26993a <=( a26992a  and  a26987a );
 a26997a <=( A267  and  A266 );
 a26998a <=( (not A265)  and  a26997a );
 a27002a <=( (not A302)  and  (not A300) );
 a27003a <=( (not A269)  and  a27002a );
 a27004a <=( a27003a  and  a26998a );
 a27008a <=( A167  and  A168 );
 a27009a <=( A170  and  a27008a );
 a27013a <=( A202  and  (not A201) );
 a27014a <=( (not A166)  and  a27013a );
 a27015a <=( a27014a  and  a27009a );
 a27019a <=( A267  and  A266 );
 a27020a <=( (not A265)  and  a27019a );
 a27024a <=( A299  and  A298 );
 a27025a <=( (not A269)  and  a27024a );
 a27026a <=( a27025a  and  a27020a );
 a27030a <=( A167  and  A168 );
 a27031a <=( A170  and  a27030a );
 a27035a <=( A202  and  (not A201) );
 a27036a <=( (not A166)  and  a27035a );
 a27037a <=( a27036a  and  a27031a );
 a27041a <=( A267  and  A266 );
 a27042a <=( (not A265)  and  a27041a );
 a27046a <=( (not A299)  and  (not A298) );
 a27047a <=( (not A269)  and  a27046a );
 a27048a <=( a27047a  and  a27042a );
 a27052a <=( A167  and  A168 );
 a27053a <=( A170  and  a27052a );
 a27057a <=( A202  and  (not A201) );
 a27058a <=( (not A166)  and  a27057a );
 a27059a <=( a27058a  and  a27053a );
 a27063a <=( A267  and  (not A266) );
 a27064a <=( A265  and  a27063a );
 a27068a <=( A301  and  (not A300) );
 a27069a <=( A268  and  a27068a );
 a27070a <=( a27069a  and  a27064a );
 a27074a <=( A167  and  A168 );
 a27075a <=( A170  and  a27074a );
 a27079a <=( A202  and  (not A201) );
 a27080a <=( (not A166)  and  a27079a );
 a27081a <=( a27080a  and  a27075a );
 a27085a <=( A267  and  (not A266) );
 a27086a <=( A265  and  a27085a );
 a27090a <=( (not A302)  and  (not A300) );
 a27091a <=( A268  and  a27090a );
 a27092a <=( a27091a  and  a27086a );
 a27096a <=( A167  and  A168 );
 a27097a <=( A170  and  a27096a );
 a27101a <=( A202  and  (not A201) );
 a27102a <=( (not A166)  and  a27101a );
 a27103a <=( a27102a  and  a27097a );
 a27107a <=( A267  and  (not A266) );
 a27108a <=( A265  and  a27107a );
 a27112a <=( A299  and  A298 );
 a27113a <=( A268  and  a27112a );
 a27114a <=( a27113a  and  a27108a );
 a27118a <=( A167  and  A168 );
 a27119a <=( A170  and  a27118a );
 a27123a <=( A202  and  (not A201) );
 a27124a <=( (not A166)  and  a27123a );
 a27125a <=( a27124a  and  a27119a );
 a27129a <=( A267  and  (not A266) );
 a27130a <=( A265  and  a27129a );
 a27134a <=( (not A299)  and  (not A298) );
 a27135a <=( A268  and  a27134a );
 a27136a <=( a27135a  and  a27130a );
 a27140a <=( A167  and  A168 );
 a27141a <=( A170  and  a27140a );
 a27145a <=( A202  and  (not A201) );
 a27146a <=( (not A166)  and  a27145a );
 a27147a <=( a27146a  and  a27141a );
 a27151a <=( A267  and  (not A266) );
 a27152a <=( A265  and  a27151a );
 a27156a <=( A301  and  (not A300) );
 a27157a <=( (not A269)  and  a27156a );
 a27158a <=( a27157a  and  a27152a );
 a27162a <=( A167  and  A168 );
 a27163a <=( A170  and  a27162a );
 a27167a <=( A202  and  (not A201) );
 a27168a <=( (not A166)  and  a27167a );
 a27169a <=( a27168a  and  a27163a );
 a27173a <=( A267  and  (not A266) );
 a27174a <=( A265  and  a27173a );
 a27178a <=( (not A302)  and  (not A300) );
 a27179a <=( (not A269)  and  a27178a );
 a27180a <=( a27179a  and  a27174a );
 a27184a <=( A167  and  A168 );
 a27185a <=( A170  and  a27184a );
 a27189a <=( A202  and  (not A201) );
 a27190a <=( (not A166)  and  a27189a );
 a27191a <=( a27190a  and  a27185a );
 a27195a <=( A267  and  (not A266) );
 a27196a <=( A265  and  a27195a );
 a27200a <=( A299  and  A298 );
 a27201a <=( (not A269)  and  a27200a );
 a27202a <=( a27201a  and  a27196a );
 a27206a <=( A167  and  A168 );
 a27207a <=( A170  and  a27206a );
 a27211a <=( A202  and  (not A201) );
 a27212a <=( (not A166)  and  a27211a );
 a27213a <=( a27212a  and  a27207a );
 a27217a <=( A267  and  (not A266) );
 a27218a <=( A265  and  a27217a );
 a27222a <=( (not A299)  and  (not A298) );
 a27223a <=( (not A269)  and  a27222a );
 a27224a <=( a27223a  and  a27218a );
 a27228a <=( A167  and  A168 );
 a27229a <=( A170  and  a27228a );
 a27233a <=( A202  and  (not A201) );
 a27234a <=( (not A166)  and  a27233a );
 a27235a <=( a27234a  and  a27229a );
 a27239a <=( A298  and  (not A266) );
 a27240a <=( (not A265)  and  a27239a );
 a27244a <=( A301  and  A300 );
 a27245a <=( (not A299)  and  a27244a );
 a27246a <=( a27245a  and  a27240a );
 a27250a <=( A167  and  A168 );
 a27251a <=( A170  and  a27250a );
 a27255a <=( A202  and  (not A201) );
 a27256a <=( (not A166)  and  a27255a );
 a27257a <=( a27256a  and  a27251a );
 a27261a <=( A298  and  (not A266) );
 a27262a <=( (not A265)  and  a27261a );
 a27266a <=( (not A302)  and  A300 );
 a27267a <=( (not A299)  and  a27266a );
 a27268a <=( a27267a  and  a27262a );
 a27272a <=( A167  and  A168 );
 a27273a <=( A170  and  a27272a );
 a27277a <=( A202  and  (not A201) );
 a27278a <=( (not A166)  and  a27277a );
 a27279a <=( a27278a  and  a27273a );
 a27283a <=( (not A298)  and  (not A266) );
 a27284a <=( (not A265)  and  a27283a );
 a27288a <=( A301  and  A300 );
 a27289a <=( A299  and  a27288a );
 a27290a <=( a27289a  and  a27284a );
 a27294a <=( A167  and  A168 );
 a27295a <=( A170  and  a27294a );
 a27299a <=( A202  and  (not A201) );
 a27300a <=( (not A166)  and  a27299a );
 a27301a <=( a27300a  and  a27295a );
 a27305a <=( (not A298)  and  (not A266) );
 a27306a <=( (not A265)  and  a27305a );
 a27310a <=( (not A302)  and  A300 );
 a27311a <=( A299  and  a27310a );
 a27312a <=( a27311a  and  a27306a );
 a27316a <=( A167  and  A168 );
 a27317a <=( A170  and  a27316a );
 a27321a <=( (not A203)  and  (not A201) );
 a27322a <=( (not A166)  and  a27321a );
 a27323a <=( a27322a  and  a27317a );
 a27327a <=( A298  and  A268 );
 a27328a <=( (not A267)  and  a27327a );
 a27332a <=( A301  and  A300 );
 a27333a <=( (not A299)  and  a27332a );
 a27334a <=( a27333a  and  a27328a );
 a27338a <=( A167  and  A168 );
 a27339a <=( A170  and  a27338a );
 a27343a <=( (not A203)  and  (not A201) );
 a27344a <=( (not A166)  and  a27343a );
 a27345a <=( a27344a  and  a27339a );
 a27349a <=( A298  and  A268 );
 a27350a <=( (not A267)  and  a27349a );
 a27354a <=( (not A302)  and  A300 );
 a27355a <=( (not A299)  and  a27354a );
 a27356a <=( a27355a  and  a27350a );
 a27360a <=( A167  and  A168 );
 a27361a <=( A170  and  a27360a );
 a27365a <=( (not A203)  and  (not A201) );
 a27366a <=( (not A166)  and  a27365a );
 a27367a <=( a27366a  and  a27361a );
 a27371a <=( (not A298)  and  A268 );
 a27372a <=( (not A267)  and  a27371a );
 a27376a <=( A301  and  A300 );
 a27377a <=( A299  and  a27376a );
 a27378a <=( a27377a  and  a27372a );
 a27382a <=( A167  and  A168 );
 a27383a <=( A170  and  a27382a );
 a27387a <=( (not A203)  and  (not A201) );
 a27388a <=( (not A166)  and  a27387a );
 a27389a <=( a27388a  and  a27383a );
 a27393a <=( (not A298)  and  A268 );
 a27394a <=( (not A267)  and  a27393a );
 a27398a <=( (not A302)  and  A300 );
 a27399a <=( A299  and  a27398a );
 a27400a <=( a27399a  and  a27394a );
 a27404a <=( A167  and  A168 );
 a27405a <=( A170  and  a27404a );
 a27409a <=( (not A203)  and  (not A201) );
 a27410a <=( (not A166)  and  a27409a );
 a27411a <=( a27410a  and  a27405a );
 a27415a <=( A298  and  (not A269) );
 a27416a <=( (not A267)  and  a27415a );
 a27420a <=( A301  and  A300 );
 a27421a <=( (not A299)  and  a27420a );
 a27422a <=( a27421a  and  a27416a );
 a27426a <=( A167  and  A168 );
 a27427a <=( A170  and  a27426a );
 a27431a <=( (not A203)  and  (not A201) );
 a27432a <=( (not A166)  and  a27431a );
 a27433a <=( a27432a  and  a27427a );
 a27437a <=( A298  and  (not A269) );
 a27438a <=( (not A267)  and  a27437a );
 a27442a <=( (not A302)  and  A300 );
 a27443a <=( (not A299)  and  a27442a );
 a27444a <=( a27443a  and  a27438a );
 a27448a <=( A167  and  A168 );
 a27449a <=( A170  and  a27448a );
 a27453a <=( (not A203)  and  (not A201) );
 a27454a <=( (not A166)  and  a27453a );
 a27455a <=( a27454a  and  a27449a );
 a27459a <=( (not A298)  and  (not A269) );
 a27460a <=( (not A267)  and  a27459a );
 a27464a <=( A301  and  A300 );
 a27465a <=( A299  and  a27464a );
 a27466a <=( a27465a  and  a27460a );
 a27470a <=( A167  and  A168 );
 a27471a <=( A170  and  a27470a );
 a27475a <=( (not A203)  and  (not A201) );
 a27476a <=( (not A166)  and  a27475a );
 a27477a <=( a27476a  and  a27471a );
 a27481a <=( (not A298)  and  (not A269) );
 a27482a <=( (not A267)  and  a27481a );
 a27486a <=( (not A302)  and  A300 );
 a27487a <=( A299  and  a27486a );
 a27488a <=( a27487a  and  a27482a );
 a27492a <=( A167  and  A168 );
 a27493a <=( A170  and  a27492a );
 a27497a <=( (not A203)  and  (not A201) );
 a27498a <=( (not A166)  and  a27497a );
 a27499a <=( a27498a  and  a27493a );
 a27503a <=( A298  and  A266 );
 a27504a <=( A265  and  a27503a );
 a27508a <=( A301  and  A300 );
 a27509a <=( (not A299)  and  a27508a );
 a27510a <=( a27509a  and  a27504a );
 a27514a <=( A167  and  A168 );
 a27515a <=( A170  and  a27514a );
 a27519a <=( (not A203)  and  (not A201) );
 a27520a <=( (not A166)  and  a27519a );
 a27521a <=( a27520a  and  a27515a );
 a27525a <=( A298  and  A266 );
 a27526a <=( A265  and  a27525a );
 a27530a <=( (not A302)  and  A300 );
 a27531a <=( (not A299)  and  a27530a );
 a27532a <=( a27531a  and  a27526a );
 a27536a <=( A167  and  A168 );
 a27537a <=( A170  and  a27536a );
 a27541a <=( (not A203)  and  (not A201) );
 a27542a <=( (not A166)  and  a27541a );
 a27543a <=( a27542a  and  a27537a );
 a27547a <=( (not A298)  and  A266 );
 a27548a <=( A265  and  a27547a );
 a27552a <=( A301  and  A300 );
 a27553a <=( A299  and  a27552a );
 a27554a <=( a27553a  and  a27548a );
 a27558a <=( A167  and  A168 );
 a27559a <=( A170  and  a27558a );
 a27563a <=( (not A203)  and  (not A201) );
 a27564a <=( (not A166)  and  a27563a );
 a27565a <=( a27564a  and  a27559a );
 a27569a <=( (not A298)  and  A266 );
 a27570a <=( A265  and  a27569a );
 a27574a <=( (not A302)  and  A300 );
 a27575a <=( A299  and  a27574a );
 a27576a <=( a27575a  and  a27570a );
 a27580a <=( A167  and  A168 );
 a27581a <=( A170  and  a27580a );
 a27585a <=( (not A203)  and  (not A201) );
 a27586a <=( (not A166)  and  a27585a );
 a27587a <=( a27586a  and  a27581a );
 a27591a <=( A267  and  A266 );
 a27592a <=( (not A265)  and  a27591a );
 a27596a <=( A301  and  (not A300) );
 a27597a <=( A268  and  a27596a );
 a27598a <=( a27597a  and  a27592a );
 a27602a <=( A167  and  A168 );
 a27603a <=( A170  and  a27602a );
 a27607a <=( (not A203)  and  (not A201) );
 a27608a <=( (not A166)  and  a27607a );
 a27609a <=( a27608a  and  a27603a );
 a27613a <=( A267  and  A266 );
 a27614a <=( (not A265)  and  a27613a );
 a27618a <=( (not A302)  and  (not A300) );
 a27619a <=( A268  and  a27618a );
 a27620a <=( a27619a  and  a27614a );
 a27624a <=( A167  and  A168 );
 a27625a <=( A170  and  a27624a );
 a27629a <=( (not A203)  and  (not A201) );
 a27630a <=( (not A166)  and  a27629a );
 a27631a <=( a27630a  and  a27625a );
 a27635a <=( A267  and  A266 );
 a27636a <=( (not A265)  and  a27635a );
 a27640a <=( A299  and  A298 );
 a27641a <=( A268  and  a27640a );
 a27642a <=( a27641a  and  a27636a );
 a27646a <=( A167  and  A168 );
 a27647a <=( A170  and  a27646a );
 a27651a <=( (not A203)  and  (not A201) );
 a27652a <=( (not A166)  and  a27651a );
 a27653a <=( a27652a  and  a27647a );
 a27657a <=( A267  and  A266 );
 a27658a <=( (not A265)  and  a27657a );
 a27662a <=( (not A299)  and  (not A298) );
 a27663a <=( A268  and  a27662a );
 a27664a <=( a27663a  and  a27658a );
 a27668a <=( A167  and  A168 );
 a27669a <=( A170  and  a27668a );
 a27673a <=( (not A203)  and  (not A201) );
 a27674a <=( (not A166)  and  a27673a );
 a27675a <=( a27674a  and  a27669a );
 a27679a <=( A267  and  A266 );
 a27680a <=( (not A265)  and  a27679a );
 a27684a <=( A301  and  (not A300) );
 a27685a <=( (not A269)  and  a27684a );
 a27686a <=( a27685a  and  a27680a );
 a27690a <=( A167  and  A168 );
 a27691a <=( A170  and  a27690a );
 a27695a <=( (not A203)  and  (not A201) );
 a27696a <=( (not A166)  and  a27695a );
 a27697a <=( a27696a  and  a27691a );
 a27701a <=( A267  and  A266 );
 a27702a <=( (not A265)  and  a27701a );
 a27706a <=( (not A302)  and  (not A300) );
 a27707a <=( (not A269)  and  a27706a );
 a27708a <=( a27707a  and  a27702a );
 a27712a <=( A167  and  A168 );
 a27713a <=( A170  and  a27712a );
 a27717a <=( (not A203)  and  (not A201) );
 a27718a <=( (not A166)  and  a27717a );
 a27719a <=( a27718a  and  a27713a );
 a27723a <=( A267  and  A266 );
 a27724a <=( (not A265)  and  a27723a );
 a27728a <=( A299  and  A298 );
 a27729a <=( (not A269)  and  a27728a );
 a27730a <=( a27729a  and  a27724a );
 a27734a <=( A167  and  A168 );
 a27735a <=( A170  and  a27734a );
 a27739a <=( (not A203)  and  (not A201) );
 a27740a <=( (not A166)  and  a27739a );
 a27741a <=( a27740a  and  a27735a );
 a27745a <=( A267  and  A266 );
 a27746a <=( (not A265)  and  a27745a );
 a27750a <=( (not A299)  and  (not A298) );
 a27751a <=( (not A269)  and  a27750a );
 a27752a <=( a27751a  and  a27746a );
 a27756a <=( A167  and  A168 );
 a27757a <=( A170  and  a27756a );
 a27761a <=( (not A203)  and  (not A201) );
 a27762a <=( (not A166)  and  a27761a );
 a27763a <=( a27762a  and  a27757a );
 a27767a <=( A267  and  (not A266) );
 a27768a <=( A265  and  a27767a );
 a27772a <=( A301  and  (not A300) );
 a27773a <=( A268  and  a27772a );
 a27774a <=( a27773a  and  a27768a );
 a27778a <=( A167  and  A168 );
 a27779a <=( A170  and  a27778a );
 a27783a <=( (not A203)  and  (not A201) );
 a27784a <=( (not A166)  and  a27783a );
 a27785a <=( a27784a  and  a27779a );
 a27789a <=( A267  and  (not A266) );
 a27790a <=( A265  and  a27789a );
 a27794a <=( (not A302)  and  (not A300) );
 a27795a <=( A268  and  a27794a );
 a27796a <=( a27795a  and  a27790a );
 a27800a <=( A167  and  A168 );
 a27801a <=( A170  and  a27800a );
 a27805a <=( (not A203)  and  (not A201) );
 a27806a <=( (not A166)  and  a27805a );
 a27807a <=( a27806a  and  a27801a );
 a27811a <=( A267  and  (not A266) );
 a27812a <=( A265  and  a27811a );
 a27816a <=( A299  and  A298 );
 a27817a <=( A268  and  a27816a );
 a27818a <=( a27817a  and  a27812a );
 a27822a <=( A167  and  A168 );
 a27823a <=( A170  and  a27822a );
 a27827a <=( (not A203)  and  (not A201) );
 a27828a <=( (not A166)  and  a27827a );
 a27829a <=( a27828a  and  a27823a );
 a27833a <=( A267  and  (not A266) );
 a27834a <=( A265  and  a27833a );
 a27838a <=( (not A299)  and  (not A298) );
 a27839a <=( A268  and  a27838a );
 a27840a <=( a27839a  and  a27834a );
 a27844a <=( A167  and  A168 );
 a27845a <=( A170  and  a27844a );
 a27849a <=( (not A203)  and  (not A201) );
 a27850a <=( (not A166)  and  a27849a );
 a27851a <=( a27850a  and  a27845a );
 a27855a <=( A267  and  (not A266) );
 a27856a <=( A265  and  a27855a );
 a27860a <=( A301  and  (not A300) );
 a27861a <=( (not A269)  and  a27860a );
 a27862a <=( a27861a  and  a27856a );
 a27866a <=( A167  and  A168 );
 a27867a <=( A170  and  a27866a );
 a27871a <=( (not A203)  and  (not A201) );
 a27872a <=( (not A166)  and  a27871a );
 a27873a <=( a27872a  and  a27867a );
 a27877a <=( A267  and  (not A266) );
 a27878a <=( A265  and  a27877a );
 a27882a <=( (not A302)  and  (not A300) );
 a27883a <=( (not A269)  and  a27882a );
 a27884a <=( a27883a  and  a27878a );
 a27888a <=( A167  and  A168 );
 a27889a <=( A170  and  a27888a );
 a27893a <=( (not A203)  and  (not A201) );
 a27894a <=( (not A166)  and  a27893a );
 a27895a <=( a27894a  and  a27889a );
 a27899a <=( A267  and  (not A266) );
 a27900a <=( A265  and  a27899a );
 a27904a <=( A299  and  A298 );
 a27905a <=( (not A269)  and  a27904a );
 a27906a <=( a27905a  and  a27900a );
 a27910a <=( A167  and  A168 );
 a27911a <=( A170  and  a27910a );
 a27915a <=( (not A203)  and  (not A201) );
 a27916a <=( (not A166)  and  a27915a );
 a27917a <=( a27916a  and  a27911a );
 a27921a <=( A267  and  (not A266) );
 a27922a <=( A265  and  a27921a );
 a27926a <=( (not A299)  and  (not A298) );
 a27927a <=( (not A269)  and  a27926a );
 a27928a <=( a27927a  and  a27922a );
 a27932a <=( A167  and  A168 );
 a27933a <=( A170  and  a27932a );
 a27937a <=( (not A203)  and  (not A201) );
 a27938a <=( (not A166)  and  a27937a );
 a27939a <=( a27938a  and  a27933a );
 a27943a <=( A298  and  (not A266) );
 a27944a <=( (not A265)  and  a27943a );
 a27948a <=( A301  and  A300 );
 a27949a <=( (not A299)  and  a27948a );
 a27950a <=( a27949a  and  a27944a );
 a27954a <=( A167  and  A168 );
 a27955a <=( A170  and  a27954a );
 a27959a <=( (not A203)  and  (not A201) );
 a27960a <=( (not A166)  and  a27959a );
 a27961a <=( a27960a  and  a27955a );
 a27965a <=( A298  and  (not A266) );
 a27966a <=( (not A265)  and  a27965a );
 a27970a <=( (not A302)  and  A300 );
 a27971a <=( (not A299)  and  a27970a );
 a27972a <=( a27971a  and  a27966a );
 a27976a <=( A167  and  A168 );
 a27977a <=( A170  and  a27976a );
 a27981a <=( (not A203)  and  (not A201) );
 a27982a <=( (not A166)  and  a27981a );
 a27983a <=( a27982a  and  a27977a );
 a27987a <=( (not A298)  and  (not A266) );
 a27988a <=( (not A265)  and  a27987a );
 a27992a <=( A301  and  A300 );
 a27993a <=( A299  and  a27992a );
 a27994a <=( a27993a  and  a27988a );
 a27998a <=( A167  and  A168 );
 a27999a <=( A170  and  a27998a );
 a28003a <=( (not A203)  and  (not A201) );
 a28004a <=( (not A166)  and  a28003a );
 a28005a <=( a28004a  and  a27999a );
 a28009a <=( (not A298)  and  (not A266) );
 a28010a <=( (not A265)  and  a28009a );
 a28014a <=( (not A302)  and  A300 );
 a28015a <=( A299  and  a28014a );
 a28016a <=( a28015a  and  a28010a );
 a28020a <=( A167  and  A168 );
 a28021a <=( A170  and  a28020a );
 a28025a <=( A200  and  A199 );
 a28026a <=( (not A166)  and  a28025a );
 a28027a <=( a28026a  and  a28021a );
 a28031a <=( A298  and  A268 );
 a28032a <=( (not A267)  and  a28031a );
 a28036a <=( A301  and  A300 );
 a28037a <=( (not A299)  and  a28036a );
 a28038a <=( a28037a  and  a28032a );
 a28042a <=( A167  and  A168 );
 a28043a <=( A170  and  a28042a );
 a28047a <=( A200  and  A199 );
 a28048a <=( (not A166)  and  a28047a );
 a28049a <=( a28048a  and  a28043a );
 a28053a <=( A298  and  A268 );
 a28054a <=( (not A267)  and  a28053a );
 a28058a <=( (not A302)  and  A300 );
 a28059a <=( (not A299)  and  a28058a );
 a28060a <=( a28059a  and  a28054a );
 a28064a <=( A167  and  A168 );
 a28065a <=( A170  and  a28064a );
 a28069a <=( A200  and  A199 );
 a28070a <=( (not A166)  and  a28069a );
 a28071a <=( a28070a  and  a28065a );
 a28075a <=( (not A298)  and  A268 );
 a28076a <=( (not A267)  and  a28075a );
 a28080a <=( A301  and  A300 );
 a28081a <=( A299  and  a28080a );
 a28082a <=( a28081a  and  a28076a );
 a28086a <=( A167  and  A168 );
 a28087a <=( A170  and  a28086a );
 a28091a <=( A200  and  A199 );
 a28092a <=( (not A166)  and  a28091a );
 a28093a <=( a28092a  and  a28087a );
 a28097a <=( (not A298)  and  A268 );
 a28098a <=( (not A267)  and  a28097a );
 a28102a <=( (not A302)  and  A300 );
 a28103a <=( A299  and  a28102a );
 a28104a <=( a28103a  and  a28098a );
 a28108a <=( A167  and  A168 );
 a28109a <=( A170  and  a28108a );
 a28113a <=( A200  and  A199 );
 a28114a <=( (not A166)  and  a28113a );
 a28115a <=( a28114a  and  a28109a );
 a28119a <=( A298  and  (not A269) );
 a28120a <=( (not A267)  and  a28119a );
 a28124a <=( A301  and  A300 );
 a28125a <=( (not A299)  and  a28124a );
 a28126a <=( a28125a  and  a28120a );
 a28130a <=( A167  and  A168 );
 a28131a <=( A170  and  a28130a );
 a28135a <=( A200  and  A199 );
 a28136a <=( (not A166)  and  a28135a );
 a28137a <=( a28136a  and  a28131a );
 a28141a <=( A298  and  (not A269) );
 a28142a <=( (not A267)  and  a28141a );
 a28146a <=( (not A302)  and  A300 );
 a28147a <=( (not A299)  and  a28146a );
 a28148a <=( a28147a  and  a28142a );
 a28152a <=( A167  and  A168 );
 a28153a <=( A170  and  a28152a );
 a28157a <=( A200  and  A199 );
 a28158a <=( (not A166)  and  a28157a );
 a28159a <=( a28158a  and  a28153a );
 a28163a <=( (not A298)  and  (not A269) );
 a28164a <=( (not A267)  and  a28163a );
 a28168a <=( A301  and  A300 );
 a28169a <=( A299  and  a28168a );
 a28170a <=( a28169a  and  a28164a );
 a28174a <=( A167  and  A168 );
 a28175a <=( A170  and  a28174a );
 a28179a <=( A200  and  A199 );
 a28180a <=( (not A166)  and  a28179a );
 a28181a <=( a28180a  and  a28175a );
 a28185a <=( (not A298)  and  (not A269) );
 a28186a <=( (not A267)  and  a28185a );
 a28190a <=( (not A302)  and  A300 );
 a28191a <=( A299  and  a28190a );
 a28192a <=( a28191a  and  a28186a );
 a28196a <=( A167  and  A168 );
 a28197a <=( A170  and  a28196a );
 a28201a <=( A200  and  A199 );
 a28202a <=( (not A166)  and  a28201a );
 a28203a <=( a28202a  and  a28197a );
 a28207a <=( A298  and  A266 );
 a28208a <=( A265  and  a28207a );
 a28212a <=( A301  and  A300 );
 a28213a <=( (not A299)  and  a28212a );
 a28214a <=( a28213a  and  a28208a );
 a28218a <=( A167  and  A168 );
 a28219a <=( A170  and  a28218a );
 a28223a <=( A200  and  A199 );
 a28224a <=( (not A166)  and  a28223a );
 a28225a <=( a28224a  and  a28219a );
 a28229a <=( A298  and  A266 );
 a28230a <=( A265  and  a28229a );
 a28234a <=( (not A302)  and  A300 );
 a28235a <=( (not A299)  and  a28234a );
 a28236a <=( a28235a  and  a28230a );
 a28240a <=( A167  and  A168 );
 a28241a <=( A170  and  a28240a );
 a28245a <=( A200  and  A199 );
 a28246a <=( (not A166)  and  a28245a );
 a28247a <=( a28246a  and  a28241a );
 a28251a <=( (not A298)  and  A266 );
 a28252a <=( A265  and  a28251a );
 a28256a <=( A301  and  A300 );
 a28257a <=( A299  and  a28256a );
 a28258a <=( a28257a  and  a28252a );
 a28262a <=( A167  and  A168 );
 a28263a <=( A170  and  a28262a );
 a28267a <=( A200  and  A199 );
 a28268a <=( (not A166)  and  a28267a );
 a28269a <=( a28268a  and  a28263a );
 a28273a <=( (not A298)  and  A266 );
 a28274a <=( A265  and  a28273a );
 a28278a <=( (not A302)  and  A300 );
 a28279a <=( A299  and  a28278a );
 a28280a <=( a28279a  and  a28274a );
 a28284a <=( A167  and  A168 );
 a28285a <=( A170  and  a28284a );
 a28289a <=( A200  and  A199 );
 a28290a <=( (not A166)  and  a28289a );
 a28291a <=( a28290a  and  a28285a );
 a28295a <=( A267  and  A266 );
 a28296a <=( (not A265)  and  a28295a );
 a28300a <=( A301  and  (not A300) );
 a28301a <=( A268  and  a28300a );
 a28302a <=( a28301a  and  a28296a );
 a28306a <=( A167  and  A168 );
 a28307a <=( A170  and  a28306a );
 a28311a <=( A200  and  A199 );
 a28312a <=( (not A166)  and  a28311a );
 a28313a <=( a28312a  and  a28307a );
 a28317a <=( A267  and  A266 );
 a28318a <=( (not A265)  and  a28317a );
 a28322a <=( (not A302)  and  (not A300) );
 a28323a <=( A268  and  a28322a );
 a28324a <=( a28323a  and  a28318a );
 a28328a <=( A167  and  A168 );
 a28329a <=( A170  and  a28328a );
 a28333a <=( A200  and  A199 );
 a28334a <=( (not A166)  and  a28333a );
 a28335a <=( a28334a  and  a28329a );
 a28339a <=( A267  and  A266 );
 a28340a <=( (not A265)  and  a28339a );
 a28344a <=( A299  and  A298 );
 a28345a <=( A268  and  a28344a );
 a28346a <=( a28345a  and  a28340a );
 a28350a <=( A167  and  A168 );
 a28351a <=( A170  and  a28350a );
 a28355a <=( A200  and  A199 );
 a28356a <=( (not A166)  and  a28355a );
 a28357a <=( a28356a  and  a28351a );
 a28361a <=( A267  and  A266 );
 a28362a <=( (not A265)  and  a28361a );
 a28366a <=( (not A299)  and  (not A298) );
 a28367a <=( A268  and  a28366a );
 a28368a <=( a28367a  and  a28362a );
 a28372a <=( A167  and  A168 );
 a28373a <=( A170  and  a28372a );
 a28377a <=( A200  and  A199 );
 a28378a <=( (not A166)  and  a28377a );
 a28379a <=( a28378a  and  a28373a );
 a28383a <=( A267  and  A266 );
 a28384a <=( (not A265)  and  a28383a );
 a28388a <=( A301  and  (not A300) );
 a28389a <=( (not A269)  and  a28388a );
 a28390a <=( a28389a  and  a28384a );
 a28394a <=( A167  and  A168 );
 a28395a <=( A170  and  a28394a );
 a28399a <=( A200  and  A199 );
 a28400a <=( (not A166)  and  a28399a );
 a28401a <=( a28400a  and  a28395a );
 a28405a <=( A267  and  A266 );
 a28406a <=( (not A265)  and  a28405a );
 a28410a <=( (not A302)  and  (not A300) );
 a28411a <=( (not A269)  and  a28410a );
 a28412a <=( a28411a  and  a28406a );
 a28416a <=( A167  and  A168 );
 a28417a <=( A170  and  a28416a );
 a28421a <=( A200  and  A199 );
 a28422a <=( (not A166)  and  a28421a );
 a28423a <=( a28422a  and  a28417a );
 a28427a <=( A267  and  A266 );
 a28428a <=( (not A265)  and  a28427a );
 a28432a <=( A299  and  A298 );
 a28433a <=( (not A269)  and  a28432a );
 a28434a <=( a28433a  and  a28428a );
 a28438a <=( A167  and  A168 );
 a28439a <=( A170  and  a28438a );
 a28443a <=( A200  and  A199 );
 a28444a <=( (not A166)  and  a28443a );
 a28445a <=( a28444a  and  a28439a );
 a28449a <=( A267  and  A266 );
 a28450a <=( (not A265)  and  a28449a );
 a28454a <=( (not A299)  and  (not A298) );
 a28455a <=( (not A269)  and  a28454a );
 a28456a <=( a28455a  and  a28450a );
 a28460a <=( A167  and  A168 );
 a28461a <=( A170  and  a28460a );
 a28465a <=( A200  and  A199 );
 a28466a <=( (not A166)  and  a28465a );
 a28467a <=( a28466a  and  a28461a );
 a28471a <=( A267  and  (not A266) );
 a28472a <=( A265  and  a28471a );
 a28476a <=( A301  and  (not A300) );
 a28477a <=( A268  and  a28476a );
 a28478a <=( a28477a  and  a28472a );
 a28482a <=( A167  and  A168 );
 a28483a <=( A170  and  a28482a );
 a28487a <=( A200  and  A199 );
 a28488a <=( (not A166)  and  a28487a );
 a28489a <=( a28488a  and  a28483a );
 a28493a <=( A267  and  (not A266) );
 a28494a <=( A265  and  a28493a );
 a28498a <=( (not A302)  and  (not A300) );
 a28499a <=( A268  and  a28498a );
 a28500a <=( a28499a  and  a28494a );
 a28504a <=( A167  and  A168 );
 a28505a <=( A170  and  a28504a );
 a28509a <=( A200  and  A199 );
 a28510a <=( (not A166)  and  a28509a );
 a28511a <=( a28510a  and  a28505a );
 a28515a <=( A267  and  (not A266) );
 a28516a <=( A265  and  a28515a );
 a28520a <=( A299  and  A298 );
 a28521a <=( A268  and  a28520a );
 a28522a <=( a28521a  and  a28516a );
 a28526a <=( A167  and  A168 );
 a28527a <=( A170  and  a28526a );
 a28531a <=( A200  and  A199 );
 a28532a <=( (not A166)  and  a28531a );
 a28533a <=( a28532a  and  a28527a );
 a28537a <=( A267  and  (not A266) );
 a28538a <=( A265  and  a28537a );
 a28542a <=( (not A299)  and  (not A298) );
 a28543a <=( A268  and  a28542a );
 a28544a <=( a28543a  and  a28538a );
 a28548a <=( A167  and  A168 );
 a28549a <=( A170  and  a28548a );
 a28553a <=( A200  and  A199 );
 a28554a <=( (not A166)  and  a28553a );
 a28555a <=( a28554a  and  a28549a );
 a28559a <=( A267  and  (not A266) );
 a28560a <=( A265  and  a28559a );
 a28564a <=( A301  and  (not A300) );
 a28565a <=( (not A269)  and  a28564a );
 a28566a <=( a28565a  and  a28560a );
 a28570a <=( A167  and  A168 );
 a28571a <=( A170  and  a28570a );
 a28575a <=( A200  and  A199 );
 a28576a <=( (not A166)  and  a28575a );
 a28577a <=( a28576a  and  a28571a );
 a28581a <=( A267  and  (not A266) );
 a28582a <=( A265  and  a28581a );
 a28586a <=( (not A302)  and  (not A300) );
 a28587a <=( (not A269)  and  a28586a );
 a28588a <=( a28587a  and  a28582a );
 a28592a <=( A167  and  A168 );
 a28593a <=( A170  and  a28592a );
 a28597a <=( A200  and  A199 );
 a28598a <=( (not A166)  and  a28597a );
 a28599a <=( a28598a  and  a28593a );
 a28603a <=( A267  and  (not A266) );
 a28604a <=( A265  and  a28603a );
 a28608a <=( A299  and  A298 );
 a28609a <=( (not A269)  and  a28608a );
 a28610a <=( a28609a  and  a28604a );
 a28614a <=( A167  and  A168 );
 a28615a <=( A170  and  a28614a );
 a28619a <=( A200  and  A199 );
 a28620a <=( (not A166)  and  a28619a );
 a28621a <=( a28620a  and  a28615a );
 a28625a <=( A267  and  (not A266) );
 a28626a <=( A265  and  a28625a );
 a28630a <=( (not A299)  and  (not A298) );
 a28631a <=( (not A269)  and  a28630a );
 a28632a <=( a28631a  and  a28626a );
 a28636a <=( A167  and  A168 );
 a28637a <=( A170  and  a28636a );
 a28641a <=( A200  and  A199 );
 a28642a <=( (not A166)  and  a28641a );
 a28643a <=( a28642a  and  a28637a );
 a28647a <=( A298  and  (not A266) );
 a28648a <=( (not A265)  and  a28647a );
 a28652a <=( A301  and  A300 );
 a28653a <=( (not A299)  and  a28652a );
 a28654a <=( a28653a  and  a28648a );
 a28658a <=( A167  and  A168 );
 a28659a <=( A170  and  a28658a );
 a28663a <=( A200  and  A199 );
 a28664a <=( (not A166)  and  a28663a );
 a28665a <=( a28664a  and  a28659a );
 a28669a <=( A298  and  (not A266) );
 a28670a <=( (not A265)  and  a28669a );
 a28674a <=( (not A302)  and  A300 );
 a28675a <=( (not A299)  and  a28674a );
 a28676a <=( a28675a  and  a28670a );
 a28680a <=( A167  and  A168 );
 a28681a <=( A170  and  a28680a );
 a28685a <=( A200  and  A199 );
 a28686a <=( (not A166)  and  a28685a );
 a28687a <=( a28686a  and  a28681a );
 a28691a <=( (not A298)  and  (not A266) );
 a28692a <=( (not A265)  and  a28691a );
 a28696a <=( A301  and  A300 );
 a28697a <=( A299  and  a28696a );
 a28698a <=( a28697a  and  a28692a );
 a28702a <=( A167  and  A168 );
 a28703a <=( A170  and  a28702a );
 a28707a <=( A200  and  A199 );
 a28708a <=( (not A166)  and  a28707a );
 a28709a <=( a28708a  and  a28703a );
 a28713a <=( (not A298)  and  (not A266) );
 a28714a <=( (not A265)  and  a28713a );
 a28718a <=( (not A302)  and  A300 );
 a28719a <=( A299  and  a28718a );
 a28720a <=( a28719a  and  a28714a );
 a28724a <=( A167  and  A168 );
 a28725a <=( A170  and  a28724a );
 a28729a <=( (not A200)  and  (not A199) );
 a28730a <=( (not A166)  and  a28729a );
 a28731a <=( a28730a  and  a28725a );
 a28735a <=( A298  and  A268 );
 a28736a <=( (not A267)  and  a28735a );
 a28740a <=( A301  and  A300 );
 a28741a <=( (not A299)  and  a28740a );
 a28742a <=( a28741a  and  a28736a );
 a28746a <=( A167  and  A168 );
 a28747a <=( A170  and  a28746a );
 a28751a <=( (not A200)  and  (not A199) );
 a28752a <=( (not A166)  and  a28751a );
 a28753a <=( a28752a  and  a28747a );
 a28757a <=( A298  and  A268 );
 a28758a <=( (not A267)  and  a28757a );
 a28762a <=( (not A302)  and  A300 );
 a28763a <=( (not A299)  and  a28762a );
 a28764a <=( a28763a  and  a28758a );
 a28768a <=( A167  and  A168 );
 a28769a <=( A170  and  a28768a );
 a28773a <=( (not A200)  and  (not A199) );
 a28774a <=( (not A166)  and  a28773a );
 a28775a <=( a28774a  and  a28769a );
 a28779a <=( (not A298)  and  A268 );
 a28780a <=( (not A267)  and  a28779a );
 a28784a <=( A301  and  A300 );
 a28785a <=( A299  and  a28784a );
 a28786a <=( a28785a  and  a28780a );
 a28790a <=( A167  and  A168 );
 a28791a <=( A170  and  a28790a );
 a28795a <=( (not A200)  and  (not A199) );
 a28796a <=( (not A166)  and  a28795a );
 a28797a <=( a28796a  and  a28791a );
 a28801a <=( (not A298)  and  A268 );
 a28802a <=( (not A267)  and  a28801a );
 a28806a <=( (not A302)  and  A300 );
 a28807a <=( A299  and  a28806a );
 a28808a <=( a28807a  and  a28802a );
 a28812a <=( A167  and  A168 );
 a28813a <=( A170  and  a28812a );
 a28817a <=( (not A200)  and  (not A199) );
 a28818a <=( (not A166)  and  a28817a );
 a28819a <=( a28818a  and  a28813a );
 a28823a <=( A298  and  (not A269) );
 a28824a <=( (not A267)  and  a28823a );
 a28828a <=( A301  and  A300 );
 a28829a <=( (not A299)  and  a28828a );
 a28830a <=( a28829a  and  a28824a );
 a28834a <=( A167  and  A168 );
 a28835a <=( A170  and  a28834a );
 a28839a <=( (not A200)  and  (not A199) );
 a28840a <=( (not A166)  and  a28839a );
 a28841a <=( a28840a  and  a28835a );
 a28845a <=( A298  and  (not A269) );
 a28846a <=( (not A267)  and  a28845a );
 a28850a <=( (not A302)  and  A300 );
 a28851a <=( (not A299)  and  a28850a );
 a28852a <=( a28851a  and  a28846a );
 a28856a <=( A167  and  A168 );
 a28857a <=( A170  and  a28856a );
 a28861a <=( (not A200)  and  (not A199) );
 a28862a <=( (not A166)  and  a28861a );
 a28863a <=( a28862a  and  a28857a );
 a28867a <=( (not A298)  and  (not A269) );
 a28868a <=( (not A267)  and  a28867a );
 a28872a <=( A301  and  A300 );
 a28873a <=( A299  and  a28872a );
 a28874a <=( a28873a  and  a28868a );
 a28878a <=( A167  and  A168 );
 a28879a <=( A170  and  a28878a );
 a28883a <=( (not A200)  and  (not A199) );
 a28884a <=( (not A166)  and  a28883a );
 a28885a <=( a28884a  and  a28879a );
 a28889a <=( (not A298)  and  (not A269) );
 a28890a <=( (not A267)  and  a28889a );
 a28894a <=( (not A302)  and  A300 );
 a28895a <=( A299  and  a28894a );
 a28896a <=( a28895a  and  a28890a );
 a28900a <=( A167  and  A168 );
 a28901a <=( A170  and  a28900a );
 a28905a <=( (not A200)  and  (not A199) );
 a28906a <=( (not A166)  and  a28905a );
 a28907a <=( a28906a  and  a28901a );
 a28911a <=( A298  and  A266 );
 a28912a <=( A265  and  a28911a );
 a28916a <=( A301  and  A300 );
 a28917a <=( (not A299)  and  a28916a );
 a28918a <=( a28917a  and  a28912a );
 a28922a <=( A167  and  A168 );
 a28923a <=( A170  and  a28922a );
 a28927a <=( (not A200)  and  (not A199) );
 a28928a <=( (not A166)  and  a28927a );
 a28929a <=( a28928a  and  a28923a );
 a28933a <=( A298  and  A266 );
 a28934a <=( A265  and  a28933a );
 a28938a <=( (not A302)  and  A300 );
 a28939a <=( (not A299)  and  a28938a );
 a28940a <=( a28939a  and  a28934a );
 a28944a <=( A167  and  A168 );
 a28945a <=( A170  and  a28944a );
 a28949a <=( (not A200)  and  (not A199) );
 a28950a <=( (not A166)  and  a28949a );
 a28951a <=( a28950a  and  a28945a );
 a28955a <=( (not A298)  and  A266 );
 a28956a <=( A265  and  a28955a );
 a28960a <=( A301  and  A300 );
 a28961a <=( A299  and  a28960a );
 a28962a <=( a28961a  and  a28956a );
 a28966a <=( A167  and  A168 );
 a28967a <=( A170  and  a28966a );
 a28971a <=( (not A200)  and  (not A199) );
 a28972a <=( (not A166)  and  a28971a );
 a28973a <=( a28972a  and  a28967a );
 a28977a <=( (not A298)  and  A266 );
 a28978a <=( A265  and  a28977a );
 a28982a <=( (not A302)  and  A300 );
 a28983a <=( A299  and  a28982a );
 a28984a <=( a28983a  and  a28978a );
 a28988a <=( A167  and  A168 );
 a28989a <=( A170  and  a28988a );
 a28993a <=( (not A200)  and  (not A199) );
 a28994a <=( (not A166)  and  a28993a );
 a28995a <=( a28994a  and  a28989a );
 a28999a <=( A267  and  A266 );
 a29000a <=( (not A265)  and  a28999a );
 a29004a <=( A301  and  (not A300) );
 a29005a <=( A268  and  a29004a );
 a29006a <=( a29005a  and  a29000a );
 a29010a <=( A167  and  A168 );
 a29011a <=( A170  and  a29010a );
 a29015a <=( (not A200)  and  (not A199) );
 a29016a <=( (not A166)  and  a29015a );
 a29017a <=( a29016a  and  a29011a );
 a29021a <=( A267  and  A266 );
 a29022a <=( (not A265)  and  a29021a );
 a29026a <=( (not A302)  and  (not A300) );
 a29027a <=( A268  and  a29026a );
 a29028a <=( a29027a  and  a29022a );
 a29032a <=( A167  and  A168 );
 a29033a <=( A170  and  a29032a );
 a29037a <=( (not A200)  and  (not A199) );
 a29038a <=( (not A166)  and  a29037a );
 a29039a <=( a29038a  and  a29033a );
 a29043a <=( A267  and  A266 );
 a29044a <=( (not A265)  and  a29043a );
 a29048a <=( A299  and  A298 );
 a29049a <=( A268  and  a29048a );
 a29050a <=( a29049a  and  a29044a );
 a29054a <=( A167  and  A168 );
 a29055a <=( A170  and  a29054a );
 a29059a <=( (not A200)  and  (not A199) );
 a29060a <=( (not A166)  and  a29059a );
 a29061a <=( a29060a  and  a29055a );
 a29065a <=( A267  and  A266 );
 a29066a <=( (not A265)  and  a29065a );
 a29070a <=( (not A299)  and  (not A298) );
 a29071a <=( A268  and  a29070a );
 a29072a <=( a29071a  and  a29066a );
 a29076a <=( A167  and  A168 );
 a29077a <=( A170  and  a29076a );
 a29081a <=( (not A200)  and  (not A199) );
 a29082a <=( (not A166)  and  a29081a );
 a29083a <=( a29082a  and  a29077a );
 a29087a <=( A267  and  A266 );
 a29088a <=( (not A265)  and  a29087a );
 a29092a <=( A301  and  (not A300) );
 a29093a <=( (not A269)  and  a29092a );
 a29094a <=( a29093a  and  a29088a );
 a29098a <=( A167  and  A168 );
 a29099a <=( A170  and  a29098a );
 a29103a <=( (not A200)  and  (not A199) );
 a29104a <=( (not A166)  and  a29103a );
 a29105a <=( a29104a  and  a29099a );
 a29109a <=( A267  and  A266 );
 a29110a <=( (not A265)  and  a29109a );
 a29114a <=( (not A302)  and  (not A300) );
 a29115a <=( (not A269)  and  a29114a );
 a29116a <=( a29115a  and  a29110a );
 a29120a <=( A167  and  A168 );
 a29121a <=( A170  and  a29120a );
 a29125a <=( (not A200)  and  (not A199) );
 a29126a <=( (not A166)  and  a29125a );
 a29127a <=( a29126a  and  a29121a );
 a29131a <=( A267  and  A266 );
 a29132a <=( (not A265)  and  a29131a );
 a29136a <=( A299  and  A298 );
 a29137a <=( (not A269)  and  a29136a );
 a29138a <=( a29137a  and  a29132a );
 a29142a <=( A167  and  A168 );
 a29143a <=( A170  and  a29142a );
 a29147a <=( (not A200)  and  (not A199) );
 a29148a <=( (not A166)  and  a29147a );
 a29149a <=( a29148a  and  a29143a );
 a29153a <=( A267  and  A266 );
 a29154a <=( (not A265)  and  a29153a );
 a29158a <=( (not A299)  and  (not A298) );
 a29159a <=( (not A269)  and  a29158a );
 a29160a <=( a29159a  and  a29154a );
 a29164a <=( A167  and  A168 );
 a29165a <=( A170  and  a29164a );
 a29169a <=( (not A200)  and  (not A199) );
 a29170a <=( (not A166)  and  a29169a );
 a29171a <=( a29170a  and  a29165a );
 a29175a <=( A267  and  (not A266) );
 a29176a <=( A265  and  a29175a );
 a29180a <=( A301  and  (not A300) );
 a29181a <=( A268  and  a29180a );
 a29182a <=( a29181a  and  a29176a );
 a29186a <=( A167  and  A168 );
 a29187a <=( A170  and  a29186a );
 a29191a <=( (not A200)  and  (not A199) );
 a29192a <=( (not A166)  and  a29191a );
 a29193a <=( a29192a  and  a29187a );
 a29197a <=( A267  and  (not A266) );
 a29198a <=( A265  and  a29197a );
 a29202a <=( (not A302)  and  (not A300) );
 a29203a <=( A268  and  a29202a );
 a29204a <=( a29203a  and  a29198a );
 a29208a <=( A167  and  A168 );
 a29209a <=( A170  and  a29208a );
 a29213a <=( (not A200)  and  (not A199) );
 a29214a <=( (not A166)  and  a29213a );
 a29215a <=( a29214a  and  a29209a );
 a29219a <=( A267  and  (not A266) );
 a29220a <=( A265  and  a29219a );
 a29224a <=( A299  and  A298 );
 a29225a <=( A268  and  a29224a );
 a29226a <=( a29225a  and  a29220a );
 a29230a <=( A167  and  A168 );
 a29231a <=( A170  and  a29230a );
 a29235a <=( (not A200)  and  (not A199) );
 a29236a <=( (not A166)  and  a29235a );
 a29237a <=( a29236a  and  a29231a );
 a29241a <=( A267  and  (not A266) );
 a29242a <=( A265  and  a29241a );
 a29246a <=( (not A299)  and  (not A298) );
 a29247a <=( A268  and  a29246a );
 a29248a <=( a29247a  and  a29242a );
 a29252a <=( A167  and  A168 );
 a29253a <=( A170  and  a29252a );
 a29257a <=( (not A200)  and  (not A199) );
 a29258a <=( (not A166)  and  a29257a );
 a29259a <=( a29258a  and  a29253a );
 a29263a <=( A267  and  (not A266) );
 a29264a <=( A265  and  a29263a );
 a29268a <=( A301  and  (not A300) );
 a29269a <=( (not A269)  and  a29268a );
 a29270a <=( a29269a  and  a29264a );
 a29274a <=( A167  and  A168 );
 a29275a <=( A170  and  a29274a );
 a29279a <=( (not A200)  and  (not A199) );
 a29280a <=( (not A166)  and  a29279a );
 a29281a <=( a29280a  and  a29275a );
 a29285a <=( A267  and  (not A266) );
 a29286a <=( A265  and  a29285a );
 a29290a <=( (not A302)  and  (not A300) );
 a29291a <=( (not A269)  and  a29290a );
 a29292a <=( a29291a  and  a29286a );
 a29296a <=( A167  and  A168 );
 a29297a <=( A170  and  a29296a );
 a29301a <=( (not A200)  and  (not A199) );
 a29302a <=( (not A166)  and  a29301a );
 a29303a <=( a29302a  and  a29297a );
 a29307a <=( A267  and  (not A266) );
 a29308a <=( A265  and  a29307a );
 a29312a <=( A299  and  A298 );
 a29313a <=( (not A269)  and  a29312a );
 a29314a <=( a29313a  and  a29308a );
 a29318a <=( A167  and  A168 );
 a29319a <=( A170  and  a29318a );
 a29323a <=( (not A200)  and  (not A199) );
 a29324a <=( (not A166)  and  a29323a );
 a29325a <=( a29324a  and  a29319a );
 a29329a <=( A267  and  (not A266) );
 a29330a <=( A265  and  a29329a );
 a29334a <=( (not A299)  and  (not A298) );
 a29335a <=( (not A269)  and  a29334a );
 a29336a <=( a29335a  and  a29330a );
 a29340a <=( A167  and  A168 );
 a29341a <=( A170  and  a29340a );
 a29345a <=( (not A200)  and  (not A199) );
 a29346a <=( (not A166)  and  a29345a );
 a29347a <=( a29346a  and  a29341a );
 a29351a <=( A298  and  (not A266) );
 a29352a <=( (not A265)  and  a29351a );
 a29356a <=( A301  and  A300 );
 a29357a <=( (not A299)  and  a29356a );
 a29358a <=( a29357a  and  a29352a );
 a29362a <=( A167  and  A168 );
 a29363a <=( A170  and  a29362a );
 a29367a <=( (not A200)  and  (not A199) );
 a29368a <=( (not A166)  and  a29367a );
 a29369a <=( a29368a  and  a29363a );
 a29373a <=( A298  and  (not A266) );
 a29374a <=( (not A265)  and  a29373a );
 a29378a <=( (not A302)  and  A300 );
 a29379a <=( (not A299)  and  a29378a );
 a29380a <=( a29379a  and  a29374a );
 a29384a <=( A167  and  A168 );
 a29385a <=( A170  and  a29384a );
 a29389a <=( (not A200)  and  (not A199) );
 a29390a <=( (not A166)  and  a29389a );
 a29391a <=( a29390a  and  a29385a );
 a29395a <=( (not A298)  and  (not A266) );
 a29396a <=( (not A265)  and  a29395a );
 a29400a <=( A301  and  A300 );
 a29401a <=( A299  and  a29400a );
 a29402a <=( a29401a  and  a29396a );
 a29406a <=( A167  and  A168 );
 a29407a <=( A170  and  a29406a );
 a29411a <=( (not A200)  and  (not A199) );
 a29412a <=( (not A166)  and  a29411a );
 a29413a <=( a29412a  and  a29407a );
 a29417a <=( (not A298)  and  (not A266) );
 a29418a <=( (not A265)  and  a29417a );
 a29422a <=( (not A302)  and  A300 );
 a29423a <=( A299  and  a29422a );
 a29424a <=( a29423a  and  a29418a );
 a29428a <=( (not A167)  and  A168 );
 a29429a <=( A170  and  a29428a );
 a29433a <=( A202  and  (not A201) );
 a29434a <=( A166  and  a29433a );
 a29435a <=( a29434a  and  a29429a );
 a29439a <=( A298  and  A268 );
 a29440a <=( (not A267)  and  a29439a );
 a29444a <=( A301  and  A300 );
 a29445a <=( (not A299)  and  a29444a );
 a29446a <=( a29445a  and  a29440a );
 a29450a <=( (not A167)  and  A168 );
 a29451a <=( A170  and  a29450a );
 a29455a <=( A202  and  (not A201) );
 a29456a <=( A166  and  a29455a );
 a29457a <=( a29456a  and  a29451a );
 a29461a <=( A298  and  A268 );
 a29462a <=( (not A267)  and  a29461a );
 a29466a <=( (not A302)  and  A300 );
 a29467a <=( (not A299)  and  a29466a );
 a29468a <=( a29467a  and  a29462a );
 a29472a <=( (not A167)  and  A168 );
 a29473a <=( A170  and  a29472a );
 a29477a <=( A202  and  (not A201) );
 a29478a <=( A166  and  a29477a );
 a29479a <=( a29478a  and  a29473a );
 a29483a <=( (not A298)  and  A268 );
 a29484a <=( (not A267)  and  a29483a );
 a29488a <=( A301  and  A300 );
 a29489a <=( A299  and  a29488a );
 a29490a <=( a29489a  and  a29484a );
 a29494a <=( (not A167)  and  A168 );
 a29495a <=( A170  and  a29494a );
 a29499a <=( A202  and  (not A201) );
 a29500a <=( A166  and  a29499a );
 a29501a <=( a29500a  and  a29495a );
 a29505a <=( (not A298)  and  A268 );
 a29506a <=( (not A267)  and  a29505a );
 a29510a <=( (not A302)  and  A300 );
 a29511a <=( A299  and  a29510a );
 a29512a <=( a29511a  and  a29506a );
 a29516a <=( (not A167)  and  A168 );
 a29517a <=( A170  and  a29516a );
 a29521a <=( A202  and  (not A201) );
 a29522a <=( A166  and  a29521a );
 a29523a <=( a29522a  and  a29517a );
 a29527a <=( A298  and  (not A269) );
 a29528a <=( (not A267)  and  a29527a );
 a29532a <=( A301  and  A300 );
 a29533a <=( (not A299)  and  a29532a );
 a29534a <=( a29533a  and  a29528a );
 a29538a <=( (not A167)  and  A168 );
 a29539a <=( A170  and  a29538a );
 a29543a <=( A202  and  (not A201) );
 a29544a <=( A166  and  a29543a );
 a29545a <=( a29544a  and  a29539a );
 a29549a <=( A298  and  (not A269) );
 a29550a <=( (not A267)  and  a29549a );
 a29554a <=( (not A302)  and  A300 );
 a29555a <=( (not A299)  and  a29554a );
 a29556a <=( a29555a  and  a29550a );
 a29560a <=( (not A167)  and  A168 );
 a29561a <=( A170  and  a29560a );
 a29565a <=( A202  and  (not A201) );
 a29566a <=( A166  and  a29565a );
 a29567a <=( a29566a  and  a29561a );
 a29571a <=( (not A298)  and  (not A269) );
 a29572a <=( (not A267)  and  a29571a );
 a29576a <=( A301  and  A300 );
 a29577a <=( A299  and  a29576a );
 a29578a <=( a29577a  and  a29572a );
 a29582a <=( (not A167)  and  A168 );
 a29583a <=( A170  and  a29582a );
 a29587a <=( A202  and  (not A201) );
 a29588a <=( A166  and  a29587a );
 a29589a <=( a29588a  and  a29583a );
 a29593a <=( (not A298)  and  (not A269) );
 a29594a <=( (not A267)  and  a29593a );
 a29598a <=( (not A302)  and  A300 );
 a29599a <=( A299  and  a29598a );
 a29600a <=( a29599a  and  a29594a );
 a29604a <=( (not A167)  and  A168 );
 a29605a <=( A170  and  a29604a );
 a29609a <=( A202  and  (not A201) );
 a29610a <=( A166  and  a29609a );
 a29611a <=( a29610a  and  a29605a );
 a29615a <=( A298  and  A266 );
 a29616a <=( A265  and  a29615a );
 a29620a <=( A301  and  A300 );
 a29621a <=( (not A299)  and  a29620a );
 a29622a <=( a29621a  and  a29616a );
 a29626a <=( (not A167)  and  A168 );
 a29627a <=( A170  and  a29626a );
 a29631a <=( A202  and  (not A201) );
 a29632a <=( A166  and  a29631a );
 a29633a <=( a29632a  and  a29627a );
 a29637a <=( A298  and  A266 );
 a29638a <=( A265  and  a29637a );
 a29642a <=( (not A302)  and  A300 );
 a29643a <=( (not A299)  and  a29642a );
 a29644a <=( a29643a  and  a29638a );
 a29648a <=( (not A167)  and  A168 );
 a29649a <=( A170  and  a29648a );
 a29653a <=( A202  and  (not A201) );
 a29654a <=( A166  and  a29653a );
 a29655a <=( a29654a  and  a29649a );
 a29659a <=( (not A298)  and  A266 );
 a29660a <=( A265  and  a29659a );
 a29664a <=( A301  and  A300 );
 a29665a <=( A299  and  a29664a );
 a29666a <=( a29665a  and  a29660a );
 a29670a <=( (not A167)  and  A168 );
 a29671a <=( A170  and  a29670a );
 a29675a <=( A202  and  (not A201) );
 a29676a <=( A166  and  a29675a );
 a29677a <=( a29676a  and  a29671a );
 a29681a <=( (not A298)  and  A266 );
 a29682a <=( A265  and  a29681a );
 a29686a <=( (not A302)  and  A300 );
 a29687a <=( A299  and  a29686a );
 a29688a <=( a29687a  and  a29682a );
 a29692a <=( (not A167)  and  A168 );
 a29693a <=( A170  and  a29692a );
 a29697a <=( A202  and  (not A201) );
 a29698a <=( A166  and  a29697a );
 a29699a <=( a29698a  and  a29693a );
 a29703a <=( A267  and  A266 );
 a29704a <=( (not A265)  and  a29703a );
 a29708a <=( A301  and  (not A300) );
 a29709a <=( A268  and  a29708a );
 a29710a <=( a29709a  and  a29704a );
 a29714a <=( (not A167)  and  A168 );
 a29715a <=( A170  and  a29714a );
 a29719a <=( A202  and  (not A201) );
 a29720a <=( A166  and  a29719a );
 a29721a <=( a29720a  and  a29715a );
 a29725a <=( A267  and  A266 );
 a29726a <=( (not A265)  and  a29725a );
 a29730a <=( (not A302)  and  (not A300) );
 a29731a <=( A268  and  a29730a );
 a29732a <=( a29731a  and  a29726a );
 a29736a <=( (not A167)  and  A168 );
 a29737a <=( A170  and  a29736a );
 a29741a <=( A202  and  (not A201) );
 a29742a <=( A166  and  a29741a );
 a29743a <=( a29742a  and  a29737a );
 a29747a <=( A267  and  A266 );
 a29748a <=( (not A265)  and  a29747a );
 a29752a <=( A299  and  A298 );
 a29753a <=( A268  and  a29752a );
 a29754a <=( a29753a  and  a29748a );
 a29758a <=( (not A167)  and  A168 );
 a29759a <=( A170  and  a29758a );
 a29763a <=( A202  and  (not A201) );
 a29764a <=( A166  and  a29763a );
 a29765a <=( a29764a  and  a29759a );
 a29769a <=( A267  and  A266 );
 a29770a <=( (not A265)  and  a29769a );
 a29774a <=( (not A299)  and  (not A298) );
 a29775a <=( A268  and  a29774a );
 a29776a <=( a29775a  and  a29770a );
 a29780a <=( (not A167)  and  A168 );
 a29781a <=( A170  and  a29780a );
 a29785a <=( A202  and  (not A201) );
 a29786a <=( A166  and  a29785a );
 a29787a <=( a29786a  and  a29781a );
 a29791a <=( A267  and  A266 );
 a29792a <=( (not A265)  and  a29791a );
 a29796a <=( A301  and  (not A300) );
 a29797a <=( (not A269)  and  a29796a );
 a29798a <=( a29797a  and  a29792a );
 a29802a <=( (not A167)  and  A168 );
 a29803a <=( A170  and  a29802a );
 a29807a <=( A202  and  (not A201) );
 a29808a <=( A166  and  a29807a );
 a29809a <=( a29808a  and  a29803a );
 a29813a <=( A267  and  A266 );
 a29814a <=( (not A265)  and  a29813a );
 a29818a <=( (not A302)  and  (not A300) );
 a29819a <=( (not A269)  and  a29818a );
 a29820a <=( a29819a  and  a29814a );
 a29824a <=( (not A167)  and  A168 );
 a29825a <=( A170  and  a29824a );
 a29829a <=( A202  and  (not A201) );
 a29830a <=( A166  and  a29829a );
 a29831a <=( a29830a  and  a29825a );
 a29835a <=( A267  and  A266 );
 a29836a <=( (not A265)  and  a29835a );
 a29840a <=( A299  and  A298 );
 a29841a <=( (not A269)  and  a29840a );
 a29842a <=( a29841a  and  a29836a );
 a29846a <=( (not A167)  and  A168 );
 a29847a <=( A170  and  a29846a );
 a29851a <=( A202  and  (not A201) );
 a29852a <=( A166  and  a29851a );
 a29853a <=( a29852a  and  a29847a );
 a29857a <=( A267  and  A266 );
 a29858a <=( (not A265)  and  a29857a );
 a29862a <=( (not A299)  and  (not A298) );
 a29863a <=( (not A269)  and  a29862a );
 a29864a <=( a29863a  and  a29858a );
 a29868a <=( (not A167)  and  A168 );
 a29869a <=( A170  and  a29868a );
 a29873a <=( A202  and  (not A201) );
 a29874a <=( A166  and  a29873a );
 a29875a <=( a29874a  and  a29869a );
 a29879a <=( A267  and  (not A266) );
 a29880a <=( A265  and  a29879a );
 a29884a <=( A301  and  (not A300) );
 a29885a <=( A268  and  a29884a );
 a29886a <=( a29885a  and  a29880a );
 a29890a <=( (not A167)  and  A168 );
 a29891a <=( A170  and  a29890a );
 a29895a <=( A202  and  (not A201) );
 a29896a <=( A166  and  a29895a );
 a29897a <=( a29896a  and  a29891a );
 a29901a <=( A267  and  (not A266) );
 a29902a <=( A265  and  a29901a );
 a29906a <=( (not A302)  and  (not A300) );
 a29907a <=( A268  and  a29906a );
 a29908a <=( a29907a  and  a29902a );
 a29912a <=( (not A167)  and  A168 );
 a29913a <=( A170  and  a29912a );
 a29917a <=( A202  and  (not A201) );
 a29918a <=( A166  and  a29917a );
 a29919a <=( a29918a  and  a29913a );
 a29923a <=( A267  and  (not A266) );
 a29924a <=( A265  and  a29923a );
 a29928a <=( A299  and  A298 );
 a29929a <=( A268  and  a29928a );
 a29930a <=( a29929a  and  a29924a );
 a29934a <=( (not A167)  and  A168 );
 a29935a <=( A170  and  a29934a );
 a29939a <=( A202  and  (not A201) );
 a29940a <=( A166  and  a29939a );
 a29941a <=( a29940a  and  a29935a );
 a29945a <=( A267  and  (not A266) );
 a29946a <=( A265  and  a29945a );
 a29950a <=( (not A299)  and  (not A298) );
 a29951a <=( A268  and  a29950a );
 a29952a <=( a29951a  and  a29946a );
 a29956a <=( (not A167)  and  A168 );
 a29957a <=( A170  and  a29956a );
 a29961a <=( A202  and  (not A201) );
 a29962a <=( A166  and  a29961a );
 a29963a <=( a29962a  and  a29957a );
 a29967a <=( A267  and  (not A266) );
 a29968a <=( A265  and  a29967a );
 a29972a <=( A301  and  (not A300) );
 a29973a <=( (not A269)  and  a29972a );
 a29974a <=( a29973a  and  a29968a );
 a29978a <=( (not A167)  and  A168 );
 a29979a <=( A170  and  a29978a );
 a29983a <=( A202  and  (not A201) );
 a29984a <=( A166  and  a29983a );
 a29985a <=( a29984a  and  a29979a );
 a29989a <=( A267  and  (not A266) );
 a29990a <=( A265  and  a29989a );
 a29994a <=( (not A302)  and  (not A300) );
 a29995a <=( (not A269)  and  a29994a );
 a29996a <=( a29995a  and  a29990a );
 a30000a <=( (not A167)  and  A168 );
 a30001a <=( A170  and  a30000a );
 a30005a <=( A202  and  (not A201) );
 a30006a <=( A166  and  a30005a );
 a30007a <=( a30006a  and  a30001a );
 a30011a <=( A267  and  (not A266) );
 a30012a <=( A265  and  a30011a );
 a30016a <=( A299  and  A298 );
 a30017a <=( (not A269)  and  a30016a );
 a30018a <=( a30017a  and  a30012a );
 a30022a <=( (not A167)  and  A168 );
 a30023a <=( A170  and  a30022a );
 a30027a <=( A202  and  (not A201) );
 a30028a <=( A166  and  a30027a );
 a30029a <=( a30028a  and  a30023a );
 a30033a <=( A267  and  (not A266) );
 a30034a <=( A265  and  a30033a );
 a30038a <=( (not A299)  and  (not A298) );
 a30039a <=( (not A269)  and  a30038a );
 a30040a <=( a30039a  and  a30034a );
 a30044a <=( (not A167)  and  A168 );
 a30045a <=( A170  and  a30044a );
 a30049a <=( A202  and  (not A201) );
 a30050a <=( A166  and  a30049a );
 a30051a <=( a30050a  and  a30045a );
 a30055a <=( A298  and  (not A266) );
 a30056a <=( (not A265)  and  a30055a );
 a30060a <=( A301  and  A300 );
 a30061a <=( (not A299)  and  a30060a );
 a30062a <=( a30061a  and  a30056a );
 a30066a <=( (not A167)  and  A168 );
 a30067a <=( A170  and  a30066a );
 a30071a <=( A202  and  (not A201) );
 a30072a <=( A166  and  a30071a );
 a30073a <=( a30072a  and  a30067a );
 a30077a <=( A298  and  (not A266) );
 a30078a <=( (not A265)  and  a30077a );
 a30082a <=( (not A302)  and  A300 );
 a30083a <=( (not A299)  and  a30082a );
 a30084a <=( a30083a  and  a30078a );
 a30088a <=( (not A167)  and  A168 );
 a30089a <=( A170  and  a30088a );
 a30093a <=( A202  and  (not A201) );
 a30094a <=( A166  and  a30093a );
 a30095a <=( a30094a  and  a30089a );
 a30099a <=( (not A298)  and  (not A266) );
 a30100a <=( (not A265)  and  a30099a );
 a30104a <=( A301  and  A300 );
 a30105a <=( A299  and  a30104a );
 a30106a <=( a30105a  and  a30100a );
 a30110a <=( (not A167)  and  A168 );
 a30111a <=( A170  and  a30110a );
 a30115a <=( A202  and  (not A201) );
 a30116a <=( A166  and  a30115a );
 a30117a <=( a30116a  and  a30111a );
 a30121a <=( (not A298)  and  (not A266) );
 a30122a <=( (not A265)  and  a30121a );
 a30126a <=( (not A302)  and  A300 );
 a30127a <=( A299  and  a30126a );
 a30128a <=( a30127a  and  a30122a );
 a30132a <=( (not A167)  and  A168 );
 a30133a <=( A170  and  a30132a );
 a30137a <=( (not A203)  and  (not A201) );
 a30138a <=( A166  and  a30137a );
 a30139a <=( a30138a  and  a30133a );
 a30143a <=( A298  and  A268 );
 a30144a <=( (not A267)  and  a30143a );
 a30148a <=( A301  and  A300 );
 a30149a <=( (not A299)  and  a30148a );
 a30150a <=( a30149a  and  a30144a );
 a30154a <=( (not A167)  and  A168 );
 a30155a <=( A170  and  a30154a );
 a30159a <=( (not A203)  and  (not A201) );
 a30160a <=( A166  and  a30159a );
 a30161a <=( a30160a  and  a30155a );
 a30165a <=( A298  and  A268 );
 a30166a <=( (not A267)  and  a30165a );
 a30170a <=( (not A302)  and  A300 );
 a30171a <=( (not A299)  and  a30170a );
 a30172a <=( a30171a  and  a30166a );
 a30176a <=( (not A167)  and  A168 );
 a30177a <=( A170  and  a30176a );
 a30181a <=( (not A203)  and  (not A201) );
 a30182a <=( A166  and  a30181a );
 a30183a <=( a30182a  and  a30177a );
 a30187a <=( (not A298)  and  A268 );
 a30188a <=( (not A267)  and  a30187a );
 a30192a <=( A301  and  A300 );
 a30193a <=( A299  and  a30192a );
 a30194a <=( a30193a  and  a30188a );
 a30198a <=( (not A167)  and  A168 );
 a30199a <=( A170  and  a30198a );
 a30203a <=( (not A203)  and  (not A201) );
 a30204a <=( A166  and  a30203a );
 a30205a <=( a30204a  and  a30199a );
 a30209a <=( (not A298)  and  A268 );
 a30210a <=( (not A267)  and  a30209a );
 a30214a <=( (not A302)  and  A300 );
 a30215a <=( A299  and  a30214a );
 a30216a <=( a30215a  and  a30210a );
 a30220a <=( (not A167)  and  A168 );
 a30221a <=( A170  and  a30220a );
 a30225a <=( (not A203)  and  (not A201) );
 a30226a <=( A166  and  a30225a );
 a30227a <=( a30226a  and  a30221a );
 a30231a <=( A298  and  (not A269) );
 a30232a <=( (not A267)  and  a30231a );
 a30236a <=( A301  and  A300 );
 a30237a <=( (not A299)  and  a30236a );
 a30238a <=( a30237a  and  a30232a );
 a30242a <=( (not A167)  and  A168 );
 a30243a <=( A170  and  a30242a );
 a30247a <=( (not A203)  and  (not A201) );
 a30248a <=( A166  and  a30247a );
 a30249a <=( a30248a  and  a30243a );
 a30253a <=( A298  and  (not A269) );
 a30254a <=( (not A267)  and  a30253a );
 a30258a <=( (not A302)  and  A300 );
 a30259a <=( (not A299)  and  a30258a );
 a30260a <=( a30259a  and  a30254a );
 a30264a <=( (not A167)  and  A168 );
 a30265a <=( A170  and  a30264a );
 a30269a <=( (not A203)  and  (not A201) );
 a30270a <=( A166  and  a30269a );
 a30271a <=( a30270a  and  a30265a );
 a30275a <=( (not A298)  and  (not A269) );
 a30276a <=( (not A267)  and  a30275a );
 a30280a <=( A301  and  A300 );
 a30281a <=( A299  and  a30280a );
 a30282a <=( a30281a  and  a30276a );
 a30286a <=( (not A167)  and  A168 );
 a30287a <=( A170  and  a30286a );
 a30291a <=( (not A203)  and  (not A201) );
 a30292a <=( A166  and  a30291a );
 a30293a <=( a30292a  and  a30287a );
 a30297a <=( (not A298)  and  (not A269) );
 a30298a <=( (not A267)  and  a30297a );
 a30302a <=( (not A302)  and  A300 );
 a30303a <=( A299  and  a30302a );
 a30304a <=( a30303a  and  a30298a );
 a30308a <=( (not A167)  and  A168 );
 a30309a <=( A170  and  a30308a );
 a30313a <=( (not A203)  and  (not A201) );
 a30314a <=( A166  and  a30313a );
 a30315a <=( a30314a  and  a30309a );
 a30319a <=( A298  and  A266 );
 a30320a <=( A265  and  a30319a );
 a30324a <=( A301  and  A300 );
 a30325a <=( (not A299)  and  a30324a );
 a30326a <=( a30325a  and  a30320a );
 a30330a <=( (not A167)  and  A168 );
 a30331a <=( A170  and  a30330a );
 a30335a <=( (not A203)  and  (not A201) );
 a30336a <=( A166  and  a30335a );
 a30337a <=( a30336a  and  a30331a );
 a30341a <=( A298  and  A266 );
 a30342a <=( A265  and  a30341a );
 a30346a <=( (not A302)  and  A300 );
 a30347a <=( (not A299)  and  a30346a );
 a30348a <=( a30347a  and  a30342a );
 a30352a <=( (not A167)  and  A168 );
 a30353a <=( A170  and  a30352a );
 a30357a <=( (not A203)  and  (not A201) );
 a30358a <=( A166  and  a30357a );
 a30359a <=( a30358a  and  a30353a );
 a30363a <=( (not A298)  and  A266 );
 a30364a <=( A265  and  a30363a );
 a30368a <=( A301  and  A300 );
 a30369a <=( A299  and  a30368a );
 a30370a <=( a30369a  and  a30364a );
 a30374a <=( (not A167)  and  A168 );
 a30375a <=( A170  and  a30374a );
 a30379a <=( (not A203)  and  (not A201) );
 a30380a <=( A166  and  a30379a );
 a30381a <=( a30380a  and  a30375a );
 a30385a <=( (not A298)  and  A266 );
 a30386a <=( A265  and  a30385a );
 a30390a <=( (not A302)  and  A300 );
 a30391a <=( A299  and  a30390a );
 a30392a <=( a30391a  and  a30386a );
 a30396a <=( (not A167)  and  A168 );
 a30397a <=( A170  and  a30396a );
 a30401a <=( (not A203)  and  (not A201) );
 a30402a <=( A166  and  a30401a );
 a30403a <=( a30402a  and  a30397a );
 a30407a <=( A267  and  A266 );
 a30408a <=( (not A265)  and  a30407a );
 a30412a <=( A301  and  (not A300) );
 a30413a <=( A268  and  a30412a );
 a30414a <=( a30413a  and  a30408a );
 a30418a <=( (not A167)  and  A168 );
 a30419a <=( A170  and  a30418a );
 a30423a <=( (not A203)  and  (not A201) );
 a30424a <=( A166  and  a30423a );
 a30425a <=( a30424a  and  a30419a );
 a30429a <=( A267  and  A266 );
 a30430a <=( (not A265)  and  a30429a );
 a30434a <=( (not A302)  and  (not A300) );
 a30435a <=( A268  and  a30434a );
 a30436a <=( a30435a  and  a30430a );
 a30440a <=( (not A167)  and  A168 );
 a30441a <=( A170  and  a30440a );
 a30445a <=( (not A203)  and  (not A201) );
 a30446a <=( A166  and  a30445a );
 a30447a <=( a30446a  and  a30441a );
 a30451a <=( A267  and  A266 );
 a30452a <=( (not A265)  and  a30451a );
 a30456a <=( A299  and  A298 );
 a30457a <=( A268  and  a30456a );
 a30458a <=( a30457a  and  a30452a );
 a30462a <=( (not A167)  and  A168 );
 a30463a <=( A170  and  a30462a );
 a30467a <=( (not A203)  and  (not A201) );
 a30468a <=( A166  and  a30467a );
 a30469a <=( a30468a  and  a30463a );
 a30473a <=( A267  and  A266 );
 a30474a <=( (not A265)  and  a30473a );
 a30478a <=( (not A299)  and  (not A298) );
 a30479a <=( A268  and  a30478a );
 a30480a <=( a30479a  and  a30474a );
 a30484a <=( (not A167)  and  A168 );
 a30485a <=( A170  and  a30484a );
 a30489a <=( (not A203)  and  (not A201) );
 a30490a <=( A166  and  a30489a );
 a30491a <=( a30490a  and  a30485a );
 a30495a <=( A267  and  A266 );
 a30496a <=( (not A265)  and  a30495a );
 a30500a <=( A301  and  (not A300) );
 a30501a <=( (not A269)  and  a30500a );
 a30502a <=( a30501a  and  a30496a );
 a30506a <=( (not A167)  and  A168 );
 a30507a <=( A170  and  a30506a );
 a30511a <=( (not A203)  and  (not A201) );
 a30512a <=( A166  and  a30511a );
 a30513a <=( a30512a  and  a30507a );
 a30517a <=( A267  and  A266 );
 a30518a <=( (not A265)  and  a30517a );
 a30522a <=( (not A302)  and  (not A300) );
 a30523a <=( (not A269)  and  a30522a );
 a30524a <=( a30523a  and  a30518a );
 a30528a <=( (not A167)  and  A168 );
 a30529a <=( A170  and  a30528a );
 a30533a <=( (not A203)  and  (not A201) );
 a30534a <=( A166  and  a30533a );
 a30535a <=( a30534a  and  a30529a );
 a30539a <=( A267  and  A266 );
 a30540a <=( (not A265)  and  a30539a );
 a30544a <=( A299  and  A298 );
 a30545a <=( (not A269)  and  a30544a );
 a30546a <=( a30545a  and  a30540a );
 a30550a <=( (not A167)  and  A168 );
 a30551a <=( A170  and  a30550a );
 a30555a <=( (not A203)  and  (not A201) );
 a30556a <=( A166  and  a30555a );
 a30557a <=( a30556a  and  a30551a );
 a30561a <=( A267  and  A266 );
 a30562a <=( (not A265)  and  a30561a );
 a30566a <=( (not A299)  and  (not A298) );
 a30567a <=( (not A269)  and  a30566a );
 a30568a <=( a30567a  and  a30562a );
 a30572a <=( (not A167)  and  A168 );
 a30573a <=( A170  and  a30572a );
 a30577a <=( (not A203)  and  (not A201) );
 a30578a <=( A166  and  a30577a );
 a30579a <=( a30578a  and  a30573a );
 a30583a <=( A267  and  (not A266) );
 a30584a <=( A265  and  a30583a );
 a30588a <=( A301  and  (not A300) );
 a30589a <=( A268  and  a30588a );
 a30590a <=( a30589a  and  a30584a );
 a30594a <=( (not A167)  and  A168 );
 a30595a <=( A170  and  a30594a );
 a30599a <=( (not A203)  and  (not A201) );
 a30600a <=( A166  and  a30599a );
 a30601a <=( a30600a  and  a30595a );
 a30605a <=( A267  and  (not A266) );
 a30606a <=( A265  and  a30605a );
 a30610a <=( (not A302)  and  (not A300) );
 a30611a <=( A268  and  a30610a );
 a30612a <=( a30611a  and  a30606a );
 a30616a <=( (not A167)  and  A168 );
 a30617a <=( A170  and  a30616a );
 a30621a <=( (not A203)  and  (not A201) );
 a30622a <=( A166  and  a30621a );
 a30623a <=( a30622a  and  a30617a );
 a30627a <=( A267  and  (not A266) );
 a30628a <=( A265  and  a30627a );
 a30632a <=( A299  and  A298 );
 a30633a <=( A268  and  a30632a );
 a30634a <=( a30633a  and  a30628a );
 a30638a <=( (not A167)  and  A168 );
 a30639a <=( A170  and  a30638a );
 a30643a <=( (not A203)  and  (not A201) );
 a30644a <=( A166  and  a30643a );
 a30645a <=( a30644a  and  a30639a );
 a30649a <=( A267  and  (not A266) );
 a30650a <=( A265  and  a30649a );
 a30654a <=( (not A299)  and  (not A298) );
 a30655a <=( A268  and  a30654a );
 a30656a <=( a30655a  and  a30650a );
 a30660a <=( (not A167)  and  A168 );
 a30661a <=( A170  and  a30660a );
 a30665a <=( (not A203)  and  (not A201) );
 a30666a <=( A166  and  a30665a );
 a30667a <=( a30666a  and  a30661a );
 a30671a <=( A267  and  (not A266) );
 a30672a <=( A265  and  a30671a );
 a30676a <=( A301  and  (not A300) );
 a30677a <=( (not A269)  and  a30676a );
 a30678a <=( a30677a  and  a30672a );
 a30682a <=( (not A167)  and  A168 );
 a30683a <=( A170  and  a30682a );
 a30687a <=( (not A203)  and  (not A201) );
 a30688a <=( A166  and  a30687a );
 a30689a <=( a30688a  and  a30683a );
 a30693a <=( A267  and  (not A266) );
 a30694a <=( A265  and  a30693a );
 a30698a <=( (not A302)  and  (not A300) );
 a30699a <=( (not A269)  and  a30698a );
 a30700a <=( a30699a  and  a30694a );
 a30704a <=( (not A167)  and  A168 );
 a30705a <=( A170  and  a30704a );
 a30709a <=( (not A203)  and  (not A201) );
 a30710a <=( A166  and  a30709a );
 a30711a <=( a30710a  and  a30705a );
 a30715a <=( A267  and  (not A266) );
 a30716a <=( A265  and  a30715a );
 a30720a <=( A299  and  A298 );
 a30721a <=( (not A269)  and  a30720a );
 a30722a <=( a30721a  and  a30716a );
 a30726a <=( (not A167)  and  A168 );
 a30727a <=( A170  and  a30726a );
 a30731a <=( (not A203)  and  (not A201) );
 a30732a <=( A166  and  a30731a );
 a30733a <=( a30732a  and  a30727a );
 a30737a <=( A267  and  (not A266) );
 a30738a <=( A265  and  a30737a );
 a30742a <=( (not A299)  and  (not A298) );
 a30743a <=( (not A269)  and  a30742a );
 a30744a <=( a30743a  and  a30738a );
 a30748a <=( (not A167)  and  A168 );
 a30749a <=( A170  and  a30748a );
 a30753a <=( (not A203)  and  (not A201) );
 a30754a <=( A166  and  a30753a );
 a30755a <=( a30754a  and  a30749a );
 a30759a <=( A298  and  (not A266) );
 a30760a <=( (not A265)  and  a30759a );
 a30764a <=( A301  and  A300 );
 a30765a <=( (not A299)  and  a30764a );
 a30766a <=( a30765a  and  a30760a );
 a30770a <=( (not A167)  and  A168 );
 a30771a <=( A170  and  a30770a );
 a30775a <=( (not A203)  and  (not A201) );
 a30776a <=( A166  and  a30775a );
 a30777a <=( a30776a  and  a30771a );
 a30781a <=( A298  and  (not A266) );
 a30782a <=( (not A265)  and  a30781a );
 a30786a <=( (not A302)  and  A300 );
 a30787a <=( (not A299)  and  a30786a );
 a30788a <=( a30787a  and  a30782a );
 a30792a <=( (not A167)  and  A168 );
 a30793a <=( A170  and  a30792a );
 a30797a <=( (not A203)  and  (not A201) );
 a30798a <=( A166  and  a30797a );
 a30799a <=( a30798a  and  a30793a );
 a30803a <=( (not A298)  and  (not A266) );
 a30804a <=( (not A265)  and  a30803a );
 a30808a <=( A301  and  A300 );
 a30809a <=( A299  and  a30808a );
 a30810a <=( a30809a  and  a30804a );
 a30814a <=( (not A167)  and  A168 );
 a30815a <=( A170  and  a30814a );
 a30819a <=( (not A203)  and  (not A201) );
 a30820a <=( A166  and  a30819a );
 a30821a <=( a30820a  and  a30815a );
 a30825a <=( (not A298)  and  (not A266) );
 a30826a <=( (not A265)  and  a30825a );
 a30830a <=( (not A302)  and  A300 );
 a30831a <=( A299  and  a30830a );
 a30832a <=( a30831a  and  a30826a );
 a30836a <=( (not A167)  and  A168 );
 a30837a <=( A170  and  a30836a );
 a30841a <=( A200  and  A199 );
 a30842a <=( A166  and  a30841a );
 a30843a <=( a30842a  and  a30837a );
 a30847a <=( A298  and  A268 );
 a30848a <=( (not A267)  and  a30847a );
 a30852a <=( A301  and  A300 );
 a30853a <=( (not A299)  and  a30852a );
 a30854a <=( a30853a  and  a30848a );
 a30858a <=( (not A167)  and  A168 );
 a30859a <=( A170  and  a30858a );
 a30863a <=( A200  and  A199 );
 a30864a <=( A166  and  a30863a );
 a30865a <=( a30864a  and  a30859a );
 a30869a <=( A298  and  A268 );
 a30870a <=( (not A267)  and  a30869a );
 a30874a <=( (not A302)  and  A300 );
 a30875a <=( (not A299)  and  a30874a );
 a30876a <=( a30875a  and  a30870a );
 a30880a <=( (not A167)  and  A168 );
 a30881a <=( A170  and  a30880a );
 a30885a <=( A200  and  A199 );
 a30886a <=( A166  and  a30885a );
 a30887a <=( a30886a  and  a30881a );
 a30891a <=( (not A298)  and  A268 );
 a30892a <=( (not A267)  and  a30891a );
 a30896a <=( A301  and  A300 );
 a30897a <=( A299  and  a30896a );
 a30898a <=( a30897a  and  a30892a );
 a30902a <=( (not A167)  and  A168 );
 a30903a <=( A170  and  a30902a );
 a30907a <=( A200  and  A199 );
 a30908a <=( A166  and  a30907a );
 a30909a <=( a30908a  and  a30903a );
 a30913a <=( (not A298)  and  A268 );
 a30914a <=( (not A267)  and  a30913a );
 a30918a <=( (not A302)  and  A300 );
 a30919a <=( A299  and  a30918a );
 a30920a <=( a30919a  and  a30914a );
 a30924a <=( (not A167)  and  A168 );
 a30925a <=( A170  and  a30924a );
 a30929a <=( A200  and  A199 );
 a30930a <=( A166  and  a30929a );
 a30931a <=( a30930a  and  a30925a );
 a30935a <=( A298  and  (not A269) );
 a30936a <=( (not A267)  and  a30935a );
 a30940a <=( A301  and  A300 );
 a30941a <=( (not A299)  and  a30940a );
 a30942a <=( a30941a  and  a30936a );
 a30946a <=( (not A167)  and  A168 );
 a30947a <=( A170  and  a30946a );
 a30951a <=( A200  and  A199 );
 a30952a <=( A166  and  a30951a );
 a30953a <=( a30952a  and  a30947a );
 a30957a <=( A298  and  (not A269) );
 a30958a <=( (not A267)  and  a30957a );
 a30962a <=( (not A302)  and  A300 );
 a30963a <=( (not A299)  and  a30962a );
 a30964a <=( a30963a  and  a30958a );
 a30968a <=( (not A167)  and  A168 );
 a30969a <=( A170  and  a30968a );
 a30973a <=( A200  and  A199 );
 a30974a <=( A166  and  a30973a );
 a30975a <=( a30974a  and  a30969a );
 a30979a <=( (not A298)  and  (not A269) );
 a30980a <=( (not A267)  and  a30979a );
 a30984a <=( A301  and  A300 );
 a30985a <=( A299  and  a30984a );
 a30986a <=( a30985a  and  a30980a );
 a30990a <=( (not A167)  and  A168 );
 a30991a <=( A170  and  a30990a );
 a30995a <=( A200  and  A199 );
 a30996a <=( A166  and  a30995a );
 a30997a <=( a30996a  and  a30991a );
 a31001a <=( (not A298)  and  (not A269) );
 a31002a <=( (not A267)  and  a31001a );
 a31006a <=( (not A302)  and  A300 );
 a31007a <=( A299  and  a31006a );
 a31008a <=( a31007a  and  a31002a );
 a31012a <=( (not A167)  and  A168 );
 a31013a <=( A170  and  a31012a );
 a31017a <=( A200  and  A199 );
 a31018a <=( A166  and  a31017a );
 a31019a <=( a31018a  and  a31013a );
 a31023a <=( A298  and  A266 );
 a31024a <=( A265  and  a31023a );
 a31028a <=( A301  and  A300 );
 a31029a <=( (not A299)  and  a31028a );
 a31030a <=( a31029a  and  a31024a );
 a31034a <=( (not A167)  and  A168 );
 a31035a <=( A170  and  a31034a );
 a31039a <=( A200  and  A199 );
 a31040a <=( A166  and  a31039a );
 a31041a <=( a31040a  and  a31035a );
 a31045a <=( A298  and  A266 );
 a31046a <=( A265  and  a31045a );
 a31050a <=( (not A302)  and  A300 );
 a31051a <=( (not A299)  and  a31050a );
 a31052a <=( a31051a  and  a31046a );
 a31056a <=( (not A167)  and  A168 );
 a31057a <=( A170  and  a31056a );
 a31061a <=( A200  and  A199 );
 a31062a <=( A166  and  a31061a );
 a31063a <=( a31062a  and  a31057a );
 a31067a <=( (not A298)  and  A266 );
 a31068a <=( A265  and  a31067a );
 a31072a <=( A301  and  A300 );
 a31073a <=( A299  and  a31072a );
 a31074a <=( a31073a  and  a31068a );
 a31078a <=( (not A167)  and  A168 );
 a31079a <=( A170  and  a31078a );
 a31083a <=( A200  and  A199 );
 a31084a <=( A166  and  a31083a );
 a31085a <=( a31084a  and  a31079a );
 a31089a <=( (not A298)  and  A266 );
 a31090a <=( A265  and  a31089a );
 a31094a <=( (not A302)  and  A300 );
 a31095a <=( A299  and  a31094a );
 a31096a <=( a31095a  and  a31090a );
 a31100a <=( (not A167)  and  A168 );
 a31101a <=( A170  and  a31100a );
 a31105a <=( A200  and  A199 );
 a31106a <=( A166  and  a31105a );
 a31107a <=( a31106a  and  a31101a );
 a31111a <=( A267  and  A266 );
 a31112a <=( (not A265)  and  a31111a );
 a31116a <=( A301  and  (not A300) );
 a31117a <=( A268  and  a31116a );
 a31118a <=( a31117a  and  a31112a );
 a31122a <=( (not A167)  and  A168 );
 a31123a <=( A170  and  a31122a );
 a31127a <=( A200  and  A199 );
 a31128a <=( A166  and  a31127a );
 a31129a <=( a31128a  and  a31123a );
 a31133a <=( A267  and  A266 );
 a31134a <=( (not A265)  and  a31133a );
 a31138a <=( (not A302)  and  (not A300) );
 a31139a <=( A268  and  a31138a );
 a31140a <=( a31139a  and  a31134a );
 a31144a <=( (not A167)  and  A168 );
 a31145a <=( A170  and  a31144a );
 a31149a <=( A200  and  A199 );
 a31150a <=( A166  and  a31149a );
 a31151a <=( a31150a  and  a31145a );
 a31155a <=( A267  and  A266 );
 a31156a <=( (not A265)  and  a31155a );
 a31160a <=( A299  and  A298 );
 a31161a <=( A268  and  a31160a );
 a31162a <=( a31161a  and  a31156a );
 a31166a <=( (not A167)  and  A168 );
 a31167a <=( A170  and  a31166a );
 a31171a <=( A200  and  A199 );
 a31172a <=( A166  and  a31171a );
 a31173a <=( a31172a  and  a31167a );
 a31177a <=( A267  and  A266 );
 a31178a <=( (not A265)  and  a31177a );
 a31182a <=( (not A299)  and  (not A298) );
 a31183a <=( A268  and  a31182a );
 a31184a <=( a31183a  and  a31178a );
 a31188a <=( (not A167)  and  A168 );
 a31189a <=( A170  and  a31188a );
 a31193a <=( A200  and  A199 );
 a31194a <=( A166  and  a31193a );
 a31195a <=( a31194a  and  a31189a );
 a31199a <=( A267  and  A266 );
 a31200a <=( (not A265)  and  a31199a );
 a31204a <=( A301  and  (not A300) );
 a31205a <=( (not A269)  and  a31204a );
 a31206a <=( a31205a  and  a31200a );
 a31210a <=( (not A167)  and  A168 );
 a31211a <=( A170  and  a31210a );
 a31215a <=( A200  and  A199 );
 a31216a <=( A166  and  a31215a );
 a31217a <=( a31216a  and  a31211a );
 a31221a <=( A267  and  A266 );
 a31222a <=( (not A265)  and  a31221a );
 a31226a <=( (not A302)  and  (not A300) );
 a31227a <=( (not A269)  and  a31226a );
 a31228a <=( a31227a  and  a31222a );
 a31232a <=( (not A167)  and  A168 );
 a31233a <=( A170  and  a31232a );
 a31237a <=( A200  and  A199 );
 a31238a <=( A166  and  a31237a );
 a31239a <=( a31238a  and  a31233a );
 a31243a <=( A267  and  A266 );
 a31244a <=( (not A265)  and  a31243a );
 a31248a <=( A299  and  A298 );
 a31249a <=( (not A269)  and  a31248a );
 a31250a <=( a31249a  and  a31244a );
 a31254a <=( (not A167)  and  A168 );
 a31255a <=( A170  and  a31254a );
 a31259a <=( A200  and  A199 );
 a31260a <=( A166  and  a31259a );
 a31261a <=( a31260a  and  a31255a );
 a31265a <=( A267  and  A266 );
 a31266a <=( (not A265)  and  a31265a );
 a31270a <=( (not A299)  and  (not A298) );
 a31271a <=( (not A269)  and  a31270a );
 a31272a <=( a31271a  and  a31266a );
 a31276a <=( (not A167)  and  A168 );
 a31277a <=( A170  and  a31276a );
 a31281a <=( A200  and  A199 );
 a31282a <=( A166  and  a31281a );
 a31283a <=( a31282a  and  a31277a );
 a31287a <=( A267  and  (not A266) );
 a31288a <=( A265  and  a31287a );
 a31292a <=( A301  and  (not A300) );
 a31293a <=( A268  and  a31292a );
 a31294a <=( a31293a  and  a31288a );
 a31298a <=( (not A167)  and  A168 );
 a31299a <=( A170  and  a31298a );
 a31303a <=( A200  and  A199 );
 a31304a <=( A166  and  a31303a );
 a31305a <=( a31304a  and  a31299a );
 a31309a <=( A267  and  (not A266) );
 a31310a <=( A265  and  a31309a );
 a31314a <=( (not A302)  and  (not A300) );
 a31315a <=( A268  and  a31314a );
 a31316a <=( a31315a  and  a31310a );
 a31320a <=( (not A167)  and  A168 );
 a31321a <=( A170  and  a31320a );
 a31325a <=( A200  and  A199 );
 a31326a <=( A166  and  a31325a );
 a31327a <=( a31326a  and  a31321a );
 a31331a <=( A267  and  (not A266) );
 a31332a <=( A265  and  a31331a );
 a31336a <=( A299  and  A298 );
 a31337a <=( A268  and  a31336a );
 a31338a <=( a31337a  and  a31332a );
 a31342a <=( (not A167)  and  A168 );
 a31343a <=( A170  and  a31342a );
 a31347a <=( A200  and  A199 );
 a31348a <=( A166  and  a31347a );
 a31349a <=( a31348a  and  a31343a );
 a31353a <=( A267  and  (not A266) );
 a31354a <=( A265  and  a31353a );
 a31358a <=( (not A299)  and  (not A298) );
 a31359a <=( A268  and  a31358a );
 a31360a <=( a31359a  and  a31354a );
 a31364a <=( (not A167)  and  A168 );
 a31365a <=( A170  and  a31364a );
 a31369a <=( A200  and  A199 );
 a31370a <=( A166  and  a31369a );
 a31371a <=( a31370a  and  a31365a );
 a31375a <=( A267  and  (not A266) );
 a31376a <=( A265  and  a31375a );
 a31380a <=( A301  and  (not A300) );
 a31381a <=( (not A269)  and  a31380a );
 a31382a <=( a31381a  and  a31376a );
 a31386a <=( (not A167)  and  A168 );
 a31387a <=( A170  and  a31386a );
 a31391a <=( A200  and  A199 );
 a31392a <=( A166  and  a31391a );
 a31393a <=( a31392a  and  a31387a );
 a31397a <=( A267  and  (not A266) );
 a31398a <=( A265  and  a31397a );
 a31402a <=( (not A302)  and  (not A300) );
 a31403a <=( (not A269)  and  a31402a );
 a31404a <=( a31403a  and  a31398a );
 a31408a <=( (not A167)  and  A168 );
 a31409a <=( A170  and  a31408a );
 a31413a <=( A200  and  A199 );
 a31414a <=( A166  and  a31413a );
 a31415a <=( a31414a  and  a31409a );
 a31419a <=( A267  and  (not A266) );
 a31420a <=( A265  and  a31419a );
 a31424a <=( A299  and  A298 );
 a31425a <=( (not A269)  and  a31424a );
 a31426a <=( a31425a  and  a31420a );
 a31430a <=( (not A167)  and  A168 );
 a31431a <=( A170  and  a31430a );
 a31435a <=( A200  and  A199 );
 a31436a <=( A166  and  a31435a );
 a31437a <=( a31436a  and  a31431a );
 a31441a <=( A267  and  (not A266) );
 a31442a <=( A265  and  a31441a );
 a31446a <=( (not A299)  and  (not A298) );
 a31447a <=( (not A269)  and  a31446a );
 a31448a <=( a31447a  and  a31442a );
 a31452a <=( (not A167)  and  A168 );
 a31453a <=( A170  and  a31452a );
 a31457a <=( A200  and  A199 );
 a31458a <=( A166  and  a31457a );
 a31459a <=( a31458a  and  a31453a );
 a31463a <=( A298  and  (not A266) );
 a31464a <=( (not A265)  and  a31463a );
 a31468a <=( A301  and  A300 );
 a31469a <=( (not A299)  and  a31468a );
 a31470a <=( a31469a  and  a31464a );
 a31474a <=( (not A167)  and  A168 );
 a31475a <=( A170  and  a31474a );
 a31479a <=( A200  and  A199 );
 a31480a <=( A166  and  a31479a );
 a31481a <=( a31480a  and  a31475a );
 a31485a <=( A298  and  (not A266) );
 a31486a <=( (not A265)  and  a31485a );
 a31490a <=( (not A302)  and  A300 );
 a31491a <=( (not A299)  and  a31490a );
 a31492a <=( a31491a  and  a31486a );
 a31496a <=( (not A167)  and  A168 );
 a31497a <=( A170  and  a31496a );
 a31501a <=( A200  and  A199 );
 a31502a <=( A166  and  a31501a );
 a31503a <=( a31502a  and  a31497a );
 a31507a <=( (not A298)  and  (not A266) );
 a31508a <=( (not A265)  and  a31507a );
 a31512a <=( A301  and  A300 );
 a31513a <=( A299  and  a31512a );
 a31514a <=( a31513a  and  a31508a );
 a31518a <=( (not A167)  and  A168 );
 a31519a <=( A170  and  a31518a );
 a31523a <=( A200  and  A199 );
 a31524a <=( A166  and  a31523a );
 a31525a <=( a31524a  and  a31519a );
 a31529a <=( (not A298)  and  (not A266) );
 a31530a <=( (not A265)  and  a31529a );
 a31534a <=( (not A302)  and  A300 );
 a31535a <=( A299  and  a31534a );
 a31536a <=( a31535a  and  a31530a );
 a31540a <=( (not A167)  and  A168 );
 a31541a <=( A170  and  a31540a );
 a31545a <=( (not A200)  and  (not A199) );
 a31546a <=( A166  and  a31545a );
 a31547a <=( a31546a  and  a31541a );
 a31551a <=( A298  and  A268 );
 a31552a <=( (not A267)  and  a31551a );
 a31556a <=( A301  and  A300 );
 a31557a <=( (not A299)  and  a31556a );
 a31558a <=( a31557a  and  a31552a );
 a31562a <=( (not A167)  and  A168 );
 a31563a <=( A170  and  a31562a );
 a31567a <=( (not A200)  and  (not A199) );
 a31568a <=( A166  and  a31567a );
 a31569a <=( a31568a  and  a31563a );
 a31573a <=( A298  and  A268 );
 a31574a <=( (not A267)  and  a31573a );
 a31578a <=( (not A302)  and  A300 );
 a31579a <=( (not A299)  and  a31578a );
 a31580a <=( a31579a  and  a31574a );
 a31584a <=( (not A167)  and  A168 );
 a31585a <=( A170  and  a31584a );
 a31589a <=( (not A200)  and  (not A199) );
 a31590a <=( A166  and  a31589a );
 a31591a <=( a31590a  and  a31585a );
 a31595a <=( (not A298)  and  A268 );
 a31596a <=( (not A267)  and  a31595a );
 a31600a <=( A301  and  A300 );
 a31601a <=( A299  and  a31600a );
 a31602a <=( a31601a  and  a31596a );
 a31606a <=( (not A167)  and  A168 );
 a31607a <=( A170  and  a31606a );
 a31611a <=( (not A200)  and  (not A199) );
 a31612a <=( A166  and  a31611a );
 a31613a <=( a31612a  and  a31607a );
 a31617a <=( (not A298)  and  A268 );
 a31618a <=( (not A267)  and  a31617a );
 a31622a <=( (not A302)  and  A300 );
 a31623a <=( A299  and  a31622a );
 a31624a <=( a31623a  and  a31618a );
 a31628a <=( (not A167)  and  A168 );
 a31629a <=( A170  and  a31628a );
 a31633a <=( (not A200)  and  (not A199) );
 a31634a <=( A166  and  a31633a );
 a31635a <=( a31634a  and  a31629a );
 a31639a <=( A298  and  (not A269) );
 a31640a <=( (not A267)  and  a31639a );
 a31644a <=( A301  and  A300 );
 a31645a <=( (not A299)  and  a31644a );
 a31646a <=( a31645a  and  a31640a );
 a31650a <=( (not A167)  and  A168 );
 a31651a <=( A170  and  a31650a );
 a31655a <=( (not A200)  and  (not A199) );
 a31656a <=( A166  and  a31655a );
 a31657a <=( a31656a  and  a31651a );
 a31661a <=( A298  and  (not A269) );
 a31662a <=( (not A267)  and  a31661a );
 a31666a <=( (not A302)  and  A300 );
 a31667a <=( (not A299)  and  a31666a );
 a31668a <=( a31667a  and  a31662a );
 a31672a <=( (not A167)  and  A168 );
 a31673a <=( A170  and  a31672a );
 a31677a <=( (not A200)  and  (not A199) );
 a31678a <=( A166  and  a31677a );
 a31679a <=( a31678a  and  a31673a );
 a31683a <=( (not A298)  and  (not A269) );
 a31684a <=( (not A267)  and  a31683a );
 a31688a <=( A301  and  A300 );
 a31689a <=( A299  and  a31688a );
 a31690a <=( a31689a  and  a31684a );
 a31694a <=( (not A167)  and  A168 );
 a31695a <=( A170  and  a31694a );
 a31699a <=( (not A200)  and  (not A199) );
 a31700a <=( A166  and  a31699a );
 a31701a <=( a31700a  and  a31695a );
 a31705a <=( (not A298)  and  (not A269) );
 a31706a <=( (not A267)  and  a31705a );
 a31710a <=( (not A302)  and  A300 );
 a31711a <=( A299  and  a31710a );
 a31712a <=( a31711a  and  a31706a );
 a31716a <=( (not A167)  and  A168 );
 a31717a <=( A170  and  a31716a );
 a31721a <=( (not A200)  and  (not A199) );
 a31722a <=( A166  and  a31721a );
 a31723a <=( a31722a  and  a31717a );
 a31727a <=( A298  and  A266 );
 a31728a <=( A265  and  a31727a );
 a31732a <=( A301  and  A300 );
 a31733a <=( (not A299)  and  a31732a );
 a31734a <=( a31733a  and  a31728a );
 a31738a <=( (not A167)  and  A168 );
 a31739a <=( A170  and  a31738a );
 a31743a <=( (not A200)  and  (not A199) );
 a31744a <=( A166  and  a31743a );
 a31745a <=( a31744a  and  a31739a );
 a31749a <=( A298  and  A266 );
 a31750a <=( A265  and  a31749a );
 a31754a <=( (not A302)  and  A300 );
 a31755a <=( (not A299)  and  a31754a );
 a31756a <=( a31755a  and  a31750a );
 a31760a <=( (not A167)  and  A168 );
 a31761a <=( A170  and  a31760a );
 a31765a <=( (not A200)  and  (not A199) );
 a31766a <=( A166  and  a31765a );
 a31767a <=( a31766a  and  a31761a );
 a31771a <=( (not A298)  and  A266 );
 a31772a <=( A265  and  a31771a );
 a31776a <=( A301  and  A300 );
 a31777a <=( A299  and  a31776a );
 a31778a <=( a31777a  and  a31772a );
 a31782a <=( (not A167)  and  A168 );
 a31783a <=( A170  and  a31782a );
 a31787a <=( (not A200)  and  (not A199) );
 a31788a <=( A166  and  a31787a );
 a31789a <=( a31788a  and  a31783a );
 a31793a <=( (not A298)  and  A266 );
 a31794a <=( A265  and  a31793a );
 a31798a <=( (not A302)  and  A300 );
 a31799a <=( A299  and  a31798a );
 a31800a <=( a31799a  and  a31794a );
 a31804a <=( (not A167)  and  A168 );
 a31805a <=( A170  and  a31804a );
 a31809a <=( (not A200)  and  (not A199) );
 a31810a <=( A166  and  a31809a );
 a31811a <=( a31810a  and  a31805a );
 a31815a <=( A267  and  A266 );
 a31816a <=( (not A265)  and  a31815a );
 a31820a <=( A301  and  (not A300) );
 a31821a <=( A268  and  a31820a );
 a31822a <=( a31821a  and  a31816a );
 a31826a <=( (not A167)  and  A168 );
 a31827a <=( A170  and  a31826a );
 a31831a <=( (not A200)  and  (not A199) );
 a31832a <=( A166  and  a31831a );
 a31833a <=( a31832a  and  a31827a );
 a31837a <=( A267  and  A266 );
 a31838a <=( (not A265)  and  a31837a );
 a31842a <=( (not A302)  and  (not A300) );
 a31843a <=( A268  and  a31842a );
 a31844a <=( a31843a  and  a31838a );
 a31848a <=( (not A167)  and  A168 );
 a31849a <=( A170  and  a31848a );
 a31853a <=( (not A200)  and  (not A199) );
 a31854a <=( A166  and  a31853a );
 a31855a <=( a31854a  and  a31849a );
 a31859a <=( A267  and  A266 );
 a31860a <=( (not A265)  and  a31859a );
 a31864a <=( A299  and  A298 );
 a31865a <=( A268  and  a31864a );
 a31866a <=( a31865a  and  a31860a );
 a31870a <=( (not A167)  and  A168 );
 a31871a <=( A170  and  a31870a );
 a31875a <=( (not A200)  and  (not A199) );
 a31876a <=( A166  and  a31875a );
 a31877a <=( a31876a  and  a31871a );
 a31881a <=( A267  and  A266 );
 a31882a <=( (not A265)  and  a31881a );
 a31886a <=( (not A299)  and  (not A298) );
 a31887a <=( A268  and  a31886a );
 a31888a <=( a31887a  and  a31882a );
 a31892a <=( (not A167)  and  A168 );
 a31893a <=( A170  and  a31892a );
 a31897a <=( (not A200)  and  (not A199) );
 a31898a <=( A166  and  a31897a );
 a31899a <=( a31898a  and  a31893a );
 a31903a <=( A267  and  A266 );
 a31904a <=( (not A265)  and  a31903a );
 a31908a <=( A301  and  (not A300) );
 a31909a <=( (not A269)  and  a31908a );
 a31910a <=( a31909a  and  a31904a );
 a31914a <=( (not A167)  and  A168 );
 a31915a <=( A170  and  a31914a );
 a31919a <=( (not A200)  and  (not A199) );
 a31920a <=( A166  and  a31919a );
 a31921a <=( a31920a  and  a31915a );
 a31925a <=( A267  and  A266 );
 a31926a <=( (not A265)  and  a31925a );
 a31930a <=( (not A302)  and  (not A300) );
 a31931a <=( (not A269)  and  a31930a );
 a31932a <=( a31931a  and  a31926a );
 a31936a <=( (not A167)  and  A168 );
 a31937a <=( A170  and  a31936a );
 a31941a <=( (not A200)  and  (not A199) );
 a31942a <=( A166  and  a31941a );
 a31943a <=( a31942a  and  a31937a );
 a31947a <=( A267  and  A266 );
 a31948a <=( (not A265)  and  a31947a );
 a31952a <=( A299  and  A298 );
 a31953a <=( (not A269)  and  a31952a );
 a31954a <=( a31953a  and  a31948a );
 a31958a <=( (not A167)  and  A168 );
 a31959a <=( A170  and  a31958a );
 a31963a <=( (not A200)  and  (not A199) );
 a31964a <=( A166  and  a31963a );
 a31965a <=( a31964a  and  a31959a );
 a31969a <=( A267  and  A266 );
 a31970a <=( (not A265)  and  a31969a );
 a31974a <=( (not A299)  and  (not A298) );
 a31975a <=( (not A269)  and  a31974a );
 a31976a <=( a31975a  and  a31970a );
 a31980a <=( (not A167)  and  A168 );
 a31981a <=( A170  and  a31980a );
 a31985a <=( (not A200)  and  (not A199) );
 a31986a <=( A166  and  a31985a );
 a31987a <=( a31986a  and  a31981a );
 a31991a <=( A267  and  (not A266) );
 a31992a <=( A265  and  a31991a );
 a31996a <=( A301  and  (not A300) );
 a31997a <=( A268  and  a31996a );
 a31998a <=( a31997a  and  a31992a );
 a32002a <=( (not A167)  and  A168 );
 a32003a <=( A170  and  a32002a );
 a32007a <=( (not A200)  and  (not A199) );
 a32008a <=( A166  and  a32007a );
 a32009a <=( a32008a  and  a32003a );
 a32013a <=( A267  and  (not A266) );
 a32014a <=( A265  and  a32013a );
 a32018a <=( (not A302)  and  (not A300) );
 a32019a <=( A268  and  a32018a );
 a32020a <=( a32019a  and  a32014a );
 a32024a <=( (not A167)  and  A168 );
 a32025a <=( A170  and  a32024a );
 a32029a <=( (not A200)  and  (not A199) );
 a32030a <=( A166  and  a32029a );
 a32031a <=( a32030a  and  a32025a );
 a32035a <=( A267  and  (not A266) );
 a32036a <=( A265  and  a32035a );
 a32040a <=( A299  and  A298 );
 a32041a <=( A268  and  a32040a );
 a32042a <=( a32041a  and  a32036a );
 a32046a <=( (not A167)  and  A168 );
 a32047a <=( A170  and  a32046a );
 a32051a <=( (not A200)  and  (not A199) );
 a32052a <=( A166  and  a32051a );
 a32053a <=( a32052a  and  a32047a );
 a32057a <=( A267  and  (not A266) );
 a32058a <=( A265  and  a32057a );
 a32062a <=( (not A299)  and  (not A298) );
 a32063a <=( A268  and  a32062a );
 a32064a <=( a32063a  and  a32058a );
 a32068a <=( (not A167)  and  A168 );
 a32069a <=( A170  and  a32068a );
 a32073a <=( (not A200)  and  (not A199) );
 a32074a <=( A166  and  a32073a );
 a32075a <=( a32074a  and  a32069a );
 a32079a <=( A267  and  (not A266) );
 a32080a <=( A265  and  a32079a );
 a32084a <=( A301  and  (not A300) );
 a32085a <=( (not A269)  and  a32084a );
 a32086a <=( a32085a  and  a32080a );
 a32090a <=( (not A167)  and  A168 );
 a32091a <=( A170  and  a32090a );
 a32095a <=( (not A200)  and  (not A199) );
 a32096a <=( A166  and  a32095a );
 a32097a <=( a32096a  and  a32091a );
 a32101a <=( A267  and  (not A266) );
 a32102a <=( A265  and  a32101a );
 a32106a <=( (not A302)  and  (not A300) );
 a32107a <=( (not A269)  and  a32106a );
 a32108a <=( a32107a  and  a32102a );
 a32112a <=( (not A167)  and  A168 );
 a32113a <=( A170  and  a32112a );
 a32117a <=( (not A200)  and  (not A199) );
 a32118a <=( A166  and  a32117a );
 a32119a <=( a32118a  and  a32113a );
 a32123a <=( A267  and  (not A266) );
 a32124a <=( A265  and  a32123a );
 a32128a <=( A299  and  A298 );
 a32129a <=( (not A269)  and  a32128a );
 a32130a <=( a32129a  and  a32124a );
 a32134a <=( (not A167)  and  A168 );
 a32135a <=( A170  and  a32134a );
 a32139a <=( (not A200)  and  (not A199) );
 a32140a <=( A166  and  a32139a );
 a32141a <=( a32140a  and  a32135a );
 a32145a <=( A267  and  (not A266) );
 a32146a <=( A265  and  a32145a );
 a32150a <=( (not A299)  and  (not A298) );
 a32151a <=( (not A269)  and  a32150a );
 a32152a <=( a32151a  and  a32146a );
 a32156a <=( (not A167)  and  A168 );
 a32157a <=( A170  and  a32156a );
 a32161a <=( (not A200)  and  (not A199) );
 a32162a <=( A166  and  a32161a );
 a32163a <=( a32162a  and  a32157a );
 a32167a <=( A298  and  (not A266) );
 a32168a <=( (not A265)  and  a32167a );
 a32172a <=( A301  and  A300 );
 a32173a <=( (not A299)  and  a32172a );
 a32174a <=( a32173a  and  a32168a );
 a32178a <=( (not A167)  and  A168 );
 a32179a <=( A170  and  a32178a );
 a32183a <=( (not A200)  and  (not A199) );
 a32184a <=( A166  and  a32183a );
 a32185a <=( a32184a  and  a32179a );
 a32189a <=( A298  and  (not A266) );
 a32190a <=( (not A265)  and  a32189a );
 a32194a <=( (not A302)  and  A300 );
 a32195a <=( (not A299)  and  a32194a );
 a32196a <=( a32195a  and  a32190a );
 a32200a <=( (not A167)  and  A168 );
 a32201a <=( A170  and  a32200a );
 a32205a <=( (not A200)  and  (not A199) );
 a32206a <=( A166  and  a32205a );
 a32207a <=( a32206a  and  a32201a );
 a32211a <=( (not A298)  and  (not A266) );
 a32212a <=( (not A265)  and  a32211a );
 a32216a <=( A301  and  A300 );
 a32217a <=( A299  and  a32216a );
 a32218a <=( a32217a  and  a32212a );
 a32222a <=( (not A167)  and  A168 );
 a32223a <=( A170  and  a32222a );
 a32227a <=( (not A200)  and  (not A199) );
 a32228a <=( A166  and  a32227a );
 a32229a <=( a32228a  and  a32223a );
 a32233a <=( (not A298)  and  (not A266) );
 a32234a <=( (not A265)  and  a32233a );
 a32238a <=( (not A302)  and  A300 );
 a32239a <=( A299  and  a32238a );
 a32240a <=( a32239a  and  a32234a );
 a32244a <=( (not A232)  and  (not A168) );
 a32245a <=( A170  and  a32244a );
 a32249a <=( (not A235)  and  (not A234) );
 a32250a <=( A233  and  a32249a );
 a32251a <=( a32250a  and  a32245a );
 a32255a <=( A266  and  (not A265) );
 a32256a <=( A236  and  a32255a );
 a32260a <=( A269  and  (not A268) );
 a32261a <=( (not A267)  and  a32260a );
 a32262a <=( a32261a  and  a32256a );
 a32266a <=( (not A232)  and  (not A168) );
 a32267a <=( A170  and  a32266a );
 a32271a <=( (not A235)  and  (not A234) );
 a32272a <=( A233  and  a32271a );
 a32273a <=( a32272a  and  a32267a );
 a32277a <=( (not A266)  and  A265 );
 a32278a <=( A236  and  a32277a );
 a32282a <=( A269  and  (not A268) );
 a32283a <=( (not A267)  and  a32282a );
 a32284a <=( a32283a  and  a32278a );
 a32288a <=( A232  and  (not A168) );
 a32289a <=( A170  and  a32288a );
 a32293a <=( (not A235)  and  (not A234) );
 a32294a <=( (not A233)  and  a32293a );
 a32295a <=( a32294a  and  a32289a );
 a32299a <=( A266  and  (not A265) );
 a32300a <=( A236  and  a32299a );
 a32304a <=( A269  and  (not A268) );
 a32305a <=( (not A267)  and  a32304a );
 a32306a <=( a32305a  and  a32300a );
 a32310a <=( A232  and  (not A168) );
 a32311a <=( A170  and  a32310a );
 a32315a <=( (not A235)  and  (not A234) );
 a32316a <=( (not A233)  and  a32315a );
 a32317a <=( a32316a  and  a32311a );
 a32321a <=( (not A266)  and  A265 );
 a32322a <=( A236  and  a32321a );
 a32326a <=( A269  and  (not A268) );
 a32327a <=( (not A267)  and  a32326a );
 a32328a <=( a32327a  and  a32322a );
 a32332a <=( (not A199)  and  (not A168) );
 a32333a <=( A170  and  a32332a );
 a32337a <=( A202  and  A201 );
 a32338a <=( A200  and  a32337a );
 a32339a <=( a32338a  and  a32333a );
 a32343a <=( A269  and  (not A268) );
 a32344a <=( A267  and  a32343a );
 a32348a <=( A302  and  (not A301) );
 a32349a <=( A300  and  a32348a );
 a32350a <=( a32349a  and  a32344a );
 a32354a <=( (not A199)  and  (not A168) );
 a32355a <=( A170  and  a32354a );
 a32359a <=( (not A203)  and  A201 );
 a32360a <=( A200  and  a32359a );
 a32361a <=( a32360a  and  a32355a );
 a32365a <=( A269  and  (not A268) );
 a32366a <=( A267  and  a32365a );
 a32370a <=( A302  and  (not A301) );
 a32371a <=( A300  and  a32370a );
 a32372a <=( a32371a  and  a32366a );
 a32376a <=( (not A199)  and  (not A168) );
 a32377a <=( A170  and  a32376a );
 a32381a <=( (not A202)  and  (not A201) );
 a32382a <=( A200  and  a32381a );
 a32383a <=( a32382a  and  a32377a );
 a32387a <=( (not A268)  and  A267 );
 a32388a <=( A203  and  a32387a );
 a32392a <=( A301  and  (not A300) );
 a32393a <=( A269  and  a32392a );
 a32394a <=( a32393a  and  a32388a );
 a32398a <=( (not A199)  and  (not A168) );
 a32399a <=( A170  and  a32398a );
 a32403a <=( (not A202)  and  (not A201) );
 a32404a <=( A200  and  a32403a );
 a32405a <=( a32404a  and  a32399a );
 a32409a <=( (not A268)  and  A267 );
 a32410a <=( A203  and  a32409a );
 a32414a <=( (not A302)  and  (not A300) );
 a32415a <=( A269  and  a32414a );
 a32416a <=( a32415a  and  a32410a );
 a32420a <=( (not A199)  and  (not A168) );
 a32421a <=( A170  and  a32420a );
 a32425a <=( (not A202)  and  (not A201) );
 a32426a <=( A200  and  a32425a );
 a32427a <=( a32426a  and  a32421a );
 a32431a <=( (not A268)  and  A267 );
 a32432a <=( A203  and  a32431a );
 a32436a <=( A299  and  A298 );
 a32437a <=( A269  and  a32436a );
 a32438a <=( a32437a  and  a32432a );
 a32442a <=( (not A199)  and  (not A168) );
 a32443a <=( A170  and  a32442a );
 a32447a <=( (not A202)  and  (not A201) );
 a32448a <=( A200  and  a32447a );
 a32449a <=( a32448a  and  a32443a );
 a32453a <=( (not A268)  and  A267 );
 a32454a <=( A203  and  a32453a );
 a32458a <=( (not A299)  and  (not A298) );
 a32459a <=( A269  and  a32458a );
 a32460a <=( a32459a  and  a32454a );
 a32464a <=( (not A199)  and  (not A168) );
 a32465a <=( A170  and  a32464a );
 a32469a <=( (not A202)  and  (not A201) );
 a32470a <=( A200  and  a32469a );
 a32471a <=( a32470a  and  a32465a );
 a32475a <=( A268  and  (not A267) );
 a32476a <=( A203  and  a32475a );
 a32480a <=( A302  and  (not A301) );
 a32481a <=( A300  and  a32480a );
 a32482a <=( a32481a  and  a32476a );
 a32486a <=( (not A199)  and  (not A168) );
 a32487a <=( A170  and  a32486a );
 a32491a <=( (not A202)  and  (not A201) );
 a32492a <=( A200  and  a32491a );
 a32493a <=( a32492a  and  a32487a );
 a32497a <=( (not A269)  and  (not A267) );
 a32498a <=( A203  and  a32497a );
 a32502a <=( A302  and  (not A301) );
 a32503a <=( A300  and  a32502a );
 a32504a <=( a32503a  and  a32498a );
 a32508a <=( (not A199)  and  (not A168) );
 a32509a <=( A170  and  a32508a );
 a32513a <=( (not A202)  and  (not A201) );
 a32514a <=( A200  and  a32513a );
 a32515a <=( a32514a  and  a32509a );
 a32519a <=( A266  and  A265 );
 a32520a <=( A203  and  a32519a );
 a32524a <=( A302  and  (not A301) );
 a32525a <=( A300  and  a32524a );
 a32526a <=( a32525a  and  a32520a );
 a32530a <=( (not A199)  and  (not A168) );
 a32531a <=( A170  and  a32530a );
 a32535a <=( (not A202)  and  (not A201) );
 a32536a <=( A200  and  a32535a );
 a32537a <=( a32536a  and  a32531a );
 a32541a <=( (not A266)  and  (not A265) );
 a32542a <=( A203  and  a32541a );
 a32546a <=( A302  and  (not A301) );
 a32547a <=( A300  and  a32546a );
 a32548a <=( a32547a  and  a32542a );
 a32552a <=( A199  and  (not A168) );
 a32553a <=( A170  and  a32552a );
 a32557a <=( A202  and  A201 );
 a32558a <=( (not A200)  and  a32557a );
 a32559a <=( a32558a  and  a32553a );
 a32563a <=( A269  and  (not A268) );
 a32564a <=( A267  and  a32563a );
 a32568a <=( A302  and  (not A301) );
 a32569a <=( A300  and  a32568a );
 a32570a <=( a32569a  and  a32564a );
 a32574a <=( A199  and  (not A168) );
 a32575a <=( A170  and  a32574a );
 a32579a <=( (not A203)  and  A201 );
 a32580a <=( (not A200)  and  a32579a );
 a32581a <=( a32580a  and  a32575a );
 a32585a <=( A269  and  (not A268) );
 a32586a <=( A267  and  a32585a );
 a32590a <=( A302  and  (not A301) );
 a32591a <=( A300  and  a32590a );
 a32592a <=( a32591a  and  a32586a );
 a32596a <=( A199  and  (not A168) );
 a32597a <=( A170  and  a32596a );
 a32601a <=( (not A202)  and  (not A201) );
 a32602a <=( (not A200)  and  a32601a );
 a32603a <=( a32602a  and  a32597a );
 a32607a <=( (not A268)  and  A267 );
 a32608a <=( A203  and  a32607a );
 a32612a <=( A301  and  (not A300) );
 a32613a <=( A269  and  a32612a );
 a32614a <=( a32613a  and  a32608a );
 a32618a <=( A199  and  (not A168) );
 a32619a <=( A170  and  a32618a );
 a32623a <=( (not A202)  and  (not A201) );
 a32624a <=( (not A200)  and  a32623a );
 a32625a <=( a32624a  and  a32619a );
 a32629a <=( (not A268)  and  A267 );
 a32630a <=( A203  and  a32629a );
 a32634a <=( (not A302)  and  (not A300) );
 a32635a <=( A269  and  a32634a );
 a32636a <=( a32635a  and  a32630a );
 a32640a <=( A199  and  (not A168) );
 a32641a <=( A170  and  a32640a );
 a32645a <=( (not A202)  and  (not A201) );
 a32646a <=( (not A200)  and  a32645a );
 a32647a <=( a32646a  and  a32641a );
 a32651a <=( (not A268)  and  A267 );
 a32652a <=( A203  and  a32651a );
 a32656a <=( A299  and  A298 );
 a32657a <=( A269  and  a32656a );
 a32658a <=( a32657a  and  a32652a );
 a32662a <=( A199  and  (not A168) );
 a32663a <=( A170  and  a32662a );
 a32667a <=( (not A202)  and  (not A201) );
 a32668a <=( (not A200)  and  a32667a );
 a32669a <=( a32668a  and  a32663a );
 a32673a <=( (not A268)  and  A267 );
 a32674a <=( A203  and  a32673a );
 a32678a <=( (not A299)  and  (not A298) );
 a32679a <=( A269  and  a32678a );
 a32680a <=( a32679a  and  a32674a );
 a32684a <=( A199  and  (not A168) );
 a32685a <=( A170  and  a32684a );
 a32689a <=( (not A202)  and  (not A201) );
 a32690a <=( (not A200)  and  a32689a );
 a32691a <=( a32690a  and  a32685a );
 a32695a <=( A268  and  (not A267) );
 a32696a <=( A203  and  a32695a );
 a32700a <=( A302  and  (not A301) );
 a32701a <=( A300  and  a32700a );
 a32702a <=( a32701a  and  a32696a );
 a32706a <=( A199  and  (not A168) );
 a32707a <=( A170  and  a32706a );
 a32711a <=( (not A202)  and  (not A201) );
 a32712a <=( (not A200)  and  a32711a );
 a32713a <=( a32712a  and  a32707a );
 a32717a <=( (not A269)  and  (not A267) );
 a32718a <=( A203  and  a32717a );
 a32722a <=( A302  and  (not A301) );
 a32723a <=( A300  and  a32722a );
 a32724a <=( a32723a  and  a32718a );
 a32728a <=( A199  and  (not A168) );
 a32729a <=( A170  and  a32728a );
 a32733a <=( (not A202)  and  (not A201) );
 a32734a <=( (not A200)  and  a32733a );
 a32735a <=( a32734a  and  a32729a );
 a32739a <=( A266  and  A265 );
 a32740a <=( A203  and  a32739a );
 a32744a <=( A302  and  (not A301) );
 a32745a <=( A300  and  a32744a );
 a32746a <=( a32745a  and  a32740a );
 a32750a <=( A199  and  (not A168) );
 a32751a <=( A170  and  a32750a );
 a32755a <=( (not A202)  and  (not A201) );
 a32756a <=( (not A200)  and  a32755a );
 a32757a <=( a32756a  and  a32751a );
 a32761a <=( (not A266)  and  (not A265) );
 a32762a <=( A203  and  a32761a );
 a32766a <=( A302  and  (not A301) );
 a32767a <=( A300  and  a32766a );
 a32768a <=( a32767a  and  a32762a );
 a32772a <=( A167  and  A168 );
 a32773a <=( A169  and  a32772a );
 a32777a <=( A202  and  (not A201) );
 a32778a <=( (not A166)  and  a32777a );
 a32779a <=( a32778a  and  a32773a );
 a32783a <=( A298  and  A268 );
 a32784a <=( (not A267)  and  a32783a );
 a32788a <=( A301  and  A300 );
 a32789a <=( (not A299)  and  a32788a );
 a32790a <=( a32789a  and  a32784a );
 a32794a <=( A167  and  A168 );
 a32795a <=( A169  and  a32794a );
 a32799a <=( A202  and  (not A201) );
 a32800a <=( (not A166)  and  a32799a );
 a32801a <=( a32800a  and  a32795a );
 a32805a <=( A298  and  A268 );
 a32806a <=( (not A267)  and  a32805a );
 a32810a <=( (not A302)  and  A300 );
 a32811a <=( (not A299)  and  a32810a );
 a32812a <=( a32811a  and  a32806a );
 a32816a <=( A167  and  A168 );
 a32817a <=( A169  and  a32816a );
 a32821a <=( A202  and  (not A201) );
 a32822a <=( (not A166)  and  a32821a );
 a32823a <=( a32822a  and  a32817a );
 a32827a <=( (not A298)  and  A268 );
 a32828a <=( (not A267)  and  a32827a );
 a32832a <=( A301  and  A300 );
 a32833a <=( A299  and  a32832a );
 a32834a <=( a32833a  and  a32828a );
 a32838a <=( A167  and  A168 );
 a32839a <=( A169  and  a32838a );
 a32843a <=( A202  and  (not A201) );
 a32844a <=( (not A166)  and  a32843a );
 a32845a <=( a32844a  and  a32839a );
 a32849a <=( (not A298)  and  A268 );
 a32850a <=( (not A267)  and  a32849a );
 a32854a <=( (not A302)  and  A300 );
 a32855a <=( A299  and  a32854a );
 a32856a <=( a32855a  and  a32850a );
 a32860a <=( A167  and  A168 );
 a32861a <=( A169  and  a32860a );
 a32865a <=( A202  and  (not A201) );
 a32866a <=( (not A166)  and  a32865a );
 a32867a <=( a32866a  and  a32861a );
 a32871a <=( A298  and  (not A269) );
 a32872a <=( (not A267)  and  a32871a );
 a32876a <=( A301  and  A300 );
 a32877a <=( (not A299)  and  a32876a );
 a32878a <=( a32877a  and  a32872a );
 a32882a <=( A167  and  A168 );
 a32883a <=( A169  and  a32882a );
 a32887a <=( A202  and  (not A201) );
 a32888a <=( (not A166)  and  a32887a );
 a32889a <=( a32888a  and  a32883a );
 a32893a <=( A298  and  (not A269) );
 a32894a <=( (not A267)  and  a32893a );
 a32898a <=( (not A302)  and  A300 );
 a32899a <=( (not A299)  and  a32898a );
 a32900a <=( a32899a  and  a32894a );
 a32904a <=( A167  and  A168 );
 a32905a <=( A169  and  a32904a );
 a32909a <=( A202  and  (not A201) );
 a32910a <=( (not A166)  and  a32909a );
 a32911a <=( a32910a  and  a32905a );
 a32915a <=( (not A298)  and  (not A269) );
 a32916a <=( (not A267)  and  a32915a );
 a32920a <=( A301  and  A300 );
 a32921a <=( A299  and  a32920a );
 a32922a <=( a32921a  and  a32916a );
 a32926a <=( A167  and  A168 );
 a32927a <=( A169  and  a32926a );
 a32931a <=( A202  and  (not A201) );
 a32932a <=( (not A166)  and  a32931a );
 a32933a <=( a32932a  and  a32927a );
 a32937a <=( (not A298)  and  (not A269) );
 a32938a <=( (not A267)  and  a32937a );
 a32942a <=( (not A302)  and  A300 );
 a32943a <=( A299  and  a32942a );
 a32944a <=( a32943a  and  a32938a );
 a32948a <=( A167  and  A168 );
 a32949a <=( A169  and  a32948a );
 a32953a <=( A202  and  (not A201) );
 a32954a <=( (not A166)  and  a32953a );
 a32955a <=( a32954a  and  a32949a );
 a32959a <=( A298  and  A266 );
 a32960a <=( A265  and  a32959a );
 a32964a <=( A301  and  A300 );
 a32965a <=( (not A299)  and  a32964a );
 a32966a <=( a32965a  and  a32960a );
 a32970a <=( A167  and  A168 );
 a32971a <=( A169  and  a32970a );
 a32975a <=( A202  and  (not A201) );
 a32976a <=( (not A166)  and  a32975a );
 a32977a <=( a32976a  and  a32971a );
 a32981a <=( A298  and  A266 );
 a32982a <=( A265  and  a32981a );
 a32986a <=( (not A302)  and  A300 );
 a32987a <=( (not A299)  and  a32986a );
 a32988a <=( a32987a  and  a32982a );
 a32992a <=( A167  and  A168 );
 a32993a <=( A169  and  a32992a );
 a32997a <=( A202  and  (not A201) );
 a32998a <=( (not A166)  and  a32997a );
 a32999a <=( a32998a  and  a32993a );
 a33003a <=( (not A298)  and  A266 );
 a33004a <=( A265  and  a33003a );
 a33008a <=( A301  and  A300 );
 a33009a <=( A299  and  a33008a );
 a33010a <=( a33009a  and  a33004a );
 a33014a <=( A167  and  A168 );
 a33015a <=( A169  and  a33014a );
 a33019a <=( A202  and  (not A201) );
 a33020a <=( (not A166)  and  a33019a );
 a33021a <=( a33020a  and  a33015a );
 a33025a <=( (not A298)  and  A266 );
 a33026a <=( A265  and  a33025a );
 a33030a <=( (not A302)  and  A300 );
 a33031a <=( A299  and  a33030a );
 a33032a <=( a33031a  and  a33026a );
 a33036a <=( A167  and  A168 );
 a33037a <=( A169  and  a33036a );
 a33041a <=( A202  and  (not A201) );
 a33042a <=( (not A166)  and  a33041a );
 a33043a <=( a33042a  and  a33037a );
 a33047a <=( A267  and  A266 );
 a33048a <=( (not A265)  and  a33047a );
 a33052a <=( A301  and  (not A300) );
 a33053a <=( A268  and  a33052a );
 a33054a <=( a33053a  and  a33048a );
 a33058a <=( A167  and  A168 );
 a33059a <=( A169  and  a33058a );
 a33063a <=( A202  and  (not A201) );
 a33064a <=( (not A166)  and  a33063a );
 a33065a <=( a33064a  and  a33059a );
 a33069a <=( A267  and  A266 );
 a33070a <=( (not A265)  and  a33069a );
 a33074a <=( (not A302)  and  (not A300) );
 a33075a <=( A268  and  a33074a );
 a33076a <=( a33075a  and  a33070a );
 a33080a <=( A167  and  A168 );
 a33081a <=( A169  and  a33080a );
 a33085a <=( A202  and  (not A201) );
 a33086a <=( (not A166)  and  a33085a );
 a33087a <=( a33086a  and  a33081a );
 a33091a <=( A267  and  A266 );
 a33092a <=( (not A265)  and  a33091a );
 a33096a <=( A299  and  A298 );
 a33097a <=( A268  and  a33096a );
 a33098a <=( a33097a  and  a33092a );
 a33102a <=( A167  and  A168 );
 a33103a <=( A169  and  a33102a );
 a33107a <=( A202  and  (not A201) );
 a33108a <=( (not A166)  and  a33107a );
 a33109a <=( a33108a  and  a33103a );
 a33113a <=( A267  and  A266 );
 a33114a <=( (not A265)  and  a33113a );
 a33118a <=( (not A299)  and  (not A298) );
 a33119a <=( A268  and  a33118a );
 a33120a <=( a33119a  and  a33114a );
 a33124a <=( A167  and  A168 );
 a33125a <=( A169  and  a33124a );
 a33129a <=( A202  and  (not A201) );
 a33130a <=( (not A166)  and  a33129a );
 a33131a <=( a33130a  and  a33125a );
 a33135a <=( A267  and  A266 );
 a33136a <=( (not A265)  and  a33135a );
 a33140a <=( A301  and  (not A300) );
 a33141a <=( (not A269)  and  a33140a );
 a33142a <=( a33141a  and  a33136a );
 a33146a <=( A167  and  A168 );
 a33147a <=( A169  and  a33146a );
 a33151a <=( A202  and  (not A201) );
 a33152a <=( (not A166)  and  a33151a );
 a33153a <=( a33152a  and  a33147a );
 a33157a <=( A267  and  A266 );
 a33158a <=( (not A265)  and  a33157a );
 a33162a <=( (not A302)  and  (not A300) );
 a33163a <=( (not A269)  and  a33162a );
 a33164a <=( a33163a  and  a33158a );
 a33168a <=( A167  and  A168 );
 a33169a <=( A169  and  a33168a );
 a33173a <=( A202  and  (not A201) );
 a33174a <=( (not A166)  and  a33173a );
 a33175a <=( a33174a  and  a33169a );
 a33179a <=( A267  and  A266 );
 a33180a <=( (not A265)  and  a33179a );
 a33184a <=( A299  and  A298 );
 a33185a <=( (not A269)  and  a33184a );
 a33186a <=( a33185a  and  a33180a );
 a33190a <=( A167  and  A168 );
 a33191a <=( A169  and  a33190a );
 a33195a <=( A202  and  (not A201) );
 a33196a <=( (not A166)  and  a33195a );
 a33197a <=( a33196a  and  a33191a );
 a33201a <=( A267  and  A266 );
 a33202a <=( (not A265)  and  a33201a );
 a33206a <=( (not A299)  and  (not A298) );
 a33207a <=( (not A269)  and  a33206a );
 a33208a <=( a33207a  and  a33202a );
 a33212a <=( A167  and  A168 );
 a33213a <=( A169  and  a33212a );
 a33217a <=( A202  and  (not A201) );
 a33218a <=( (not A166)  and  a33217a );
 a33219a <=( a33218a  and  a33213a );
 a33223a <=( A267  and  (not A266) );
 a33224a <=( A265  and  a33223a );
 a33228a <=( A301  and  (not A300) );
 a33229a <=( A268  and  a33228a );
 a33230a <=( a33229a  and  a33224a );
 a33234a <=( A167  and  A168 );
 a33235a <=( A169  and  a33234a );
 a33239a <=( A202  and  (not A201) );
 a33240a <=( (not A166)  and  a33239a );
 a33241a <=( a33240a  and  a33235a );
 a33245a <=( A267  and  (not A266) );
 a33246a <=( A265  and  a33245a );
 a33250a <=( (not A302)  and  (not A300) );
 a33251a <=( A268  and  a33250a );
 a33252a <=( a33251a  and  a33246a );
 a33256a <=( A167  and  A168 );
 a33257a <=( A169  and  a33256a );
 a33261a <=( A202  and  (not A201) );
 a33262a <=( (not A166)  and  a33261a );
 a33263a <=( a33262a  and  a33257a );
 a33267a <=( A267  and  (not A266) );
 a33268a <=( A265  and  a33267a );
 a33272a <=( A299  and  A298 );
 a33273a <=( A268  and  a33272a );
 a33274a <=( a33273a  and  a33268a );
 a33278a <=( A167  and  A168 );
 a33279a <=( A169  and  a33278a );
 a33283a <=( A202  and  (not A201) );
 a33284a <=( (not A166)  and  a33283a );
 a33285a <=( a33284a  and  a33279a );
 a33289a <=( A267  and  (not A266) );
 a33290a <=( A265  and  a33289a );
 a33294a <=( (not A299)  and  (not A298) );
 a33295a <=( A268  and  a33294a );
 a33296a <=( a33295a  and  a33290a );
 a33300a <=( A167  and  A168 );
 a33301a <=( A169  and  a33300a );
 a33305a <=( A202  and  (not A201) );
 a33306a <=( (not A166)  and  a33305a );
 a33307a <=( a33306a  and  a33301a );
 a33311a <=( A267  and  (not A266) );
 a33312a <=( A265  and  a33311a );
 a33316a <=( A301  and  (not A300) );
 a33317a <=( (not A269)  and  a33316a );
 a33318a <=( a33317a  and  a33312a );
 a33322a <=( A167  and  A168 );
 a33323a <=( A169  and  a33322a );
 a33327a <=( A202  and  (not A201) );
 a33328a <=( (not A166)  and  a33327a );
 a33329a <=( a33328a  and  a33323a );
 a33333a <=( A267  and  (not A266) );
 a33334a <=( A265  and  a33333a );
 a33338a <=( (not A302)  and  (not A300) );
 a33339a <=( (not A269)  and  a33338a );
 a33340a <=( a33339a  and  a33334a );
 a33344a <=( A167  and  A168 );
 a33345a <=( A169  and  a33344a );
 a33349a <=( A202  and  (not A201) );
 a33350a <=( (not A166)  and  a33349a );
 a33351a <=( a33350a  and  a33345a );
 a33355a <=( A267  and  (not A266) );
 a33356a <=( A265  and  a33355a );
 a33360a <=( A299  and  A298 );
 a33361a <=( (not A269)  and  a33360a );
 a33362a <=( a33361a  and  a33356a );
 a33366a <=( A167  and  A168 );
 a33367a <=( A169  and  a33366a );
 a33371a <=( A202  and  (not A201) );
 a33372a <=( (not A166)  and  a33371a );
 a33373a <=( a33372a  and  a33367a );
 a33377a <=( A267  and  (not A266) );
 a33378a <=( A265  and  a33377a );
 a33382a <=( (not A299)  and  (not A298) );
 a33383a <=( (not A269)  and  a33382a );
 a33384a <=( a33383a  and  a33378a );
 a33388a <=( A167  and  A168 );
 a33389a <=( A169  and  a33388a );
 a33393a <=( A202  and  (not A201) );
 a33394a <=( (not A166)  and  a33393a );
 a33395a <=( a33394a  and  a33389a );
 a33399a <=( A298  and  (not A266) );
 a33400a <=( (not A265)  and  a33399a );
 a33404a <=( A301  and  A300 );
 a33405a <=( (not A299)  and  a33404a );
 a33406a <=( a33405a  and  a33400a );
 a33410a <=( A167  and  A168 );
 a33411a <=( A169  and  a33410a );
 a33415a <=( A202  and  (not A201) );
 a33416a <=( (not A166)  and  a33415a );
 a33417a <=( a33416a  and  a33411a );
 a33421a <=( A298  and  (not A266) );
 a33422a <=( (not A265)  and  a33421a );
 a33426a <=( (not A302)  and  A300 );
 a33427a <=( (not A299)  and  a33426a );
 a33428a <=( a33427a  and  a33422a );
 a33432a <=( A167  and  A168 );
 a33433a <=( A169  and  a33432a );
 a33437a <=( A202  and  (not A201) );
 a33438a <=( (not A166)  and  a33437a );
 a33439a <=( a33438a  and  a33433a );
 a33443a <=( (not A298)  and  (not A266) );
 a33444a <=( (not A265)  and  a33443a );
 a33448a <=( A301  and  A300 );
 a33449a <=( A299  and  a33448a );
 a33450a <=( a33449a  and  a33444a );
 a33454a <=( A167  and  A168 );
 a33455a <=( A169  and  a33454a );
 a33459a <=( A202  and  (not A201) );
 a33460a <=( (not A166)  and  a33459a );
 a33461a <=( a33460a  and  a33455a );
 a33465a <=( (not A298)  and  (not A266) );
 a33466a <=( (not A265)  and  a33465a );
 a33470a <=( (not A302)  and  A300 );
 a33471a <=( A299  and  a33470a );
 a33472a <=( a33471a  and  a33466a );
 a33476a <=( A167  and  A168 );
 a33477a <=( A169  and  a33476a );
 a33481a <=( (not A203)  and  (not A201) );
 a33482a <=( (not A166)  and  a33481a );
 a33483a <=( a33482a  and  a33477a );
 a33487a <=( A298  and  A268 );
 a33488a <=( (not A267)  and  a33487a );
 a33492a <=( A301  and  A300 );
 a33493a <=( (not A299)  and  a33492a );
 a33494a <=( a33493a  and  a33488a );
 a33498a <=( A167  and  A168 );
 a33499a <=( A169  and  a33498a );
 a33503a <=( (not A203)  and  (not A201) );
 a33504a <=( (not A166)  and  a33503a );
 a33505a <=( a33504a  and  a33499a );
 a33509a <=( A298  and  A268 );
 a33510a <=( (not A267)  and  a33509a );
 a33514a <=( (not A302)  and  A300 );
 a33515a <=( (not A299)  and  a33514a );
 a33516a <=( a33515a  and  a33510a );
 a33520a <=( A167  and  A168 );
 a33521a <=( A169  and  a33520a );
 a33525a <=( (not A203)  and  (not A201) );
 a33526a <=( (not A166)  and  a33525a );
 a33527a <=( a33526a  and  a33521a );
 a33531a <=( (not A298)  and  A268 );
 a33532a <=( (not A267)  and  a33531a );
 a33536a <=( A301  and  A300 );
 a33537a <=( A299  and  a33536a );
 a33538a <=( a33537a  and  a33532a );
 a33542a <=( A167  and  A168 );
 a33543a <=( A169  and  a33542a );
 a33547a <=( (not A203)  and  (not A201) );
 a33548a <=( (not A166)  and  a33547a );
 a33549a <=( a33548a  and  a33543a );
 a33553a <=( (not A298)  and  A268 );
 a33554a <=( (not A267)  and  a33553a );
 a33558a <=( (not A302)  and  A300 );
 a33559a <=( A299  and  a33558a );
 a33560a <=( a33559a  and  a33554a );
 a33564a <=( A167  and  A168 );
 a33565a <=( A169  and  a33564a );
 a33569a <=( (not A203)  and  (not A201) );
 a33570a <=( (not A166)  and  a33569a );
 a33571a <=( a33570a  and  a33565a );
 a33575a <=( A298  and  (not A269) );
 a33576a <=( (not A267)  and  a33575a );
 a33580a <=( A301  and  A300 );
 a33581a <=( (not A299)  and  a33580a );
 a33582a <=( a33581a  and  a33576a );
 a33586a <=( A167  and  A168 );
 a33587a <=( A169  and  a33586a );
 a33591a <=( (not A203)  and  (not A201) );
 a33592a <=( (not A166)  and  a33591a );
 a33593a <=( a33592a  and  a33587a );
 a33597a <=( A298  and  (not A269) );
 a33598a <=( (not A267)  and  a33597a );
 a33602a <=( (not A302)  and  A300 );
 a33603a <=( (not A299)  and  a33602a );
 a33604a <=( a33603a  and  a33598a );
 a33608a <=( A167  and  A168 );
 a33609a <=( A169  and  a33608a );
 a33613a <=( (not A203)  and  (not A201) );
 a33614a <=( (not A166)  and  a33613a );
 a33615a <=( a33614a  and  a33609a );
 a33619a <=( (not A298)  and  (not A269) );
 a33620a <=( (not A267)  and  a33619a );
 a33624a <=( A301  and  A300 );
 a33625a <=( A299  and  a33624a );
 a33626a <=( a33625a  and  a33620a );
 a33630a <=( A167  and  A168 );
 a33631a <=( A169  and  a33630a );
 a33635a <=( (not A203)  and  (not A201) );
 a33636a <=( (not A166)  and  a33635a );
 a33637a <=( a33636a  and  a33631a );
 a33641a <=( (not A298)  and  (not A269) );
 a33642a <=( (not A267)  and  a33641a );
 a33646a <=( (not A302)  and  A300 );
 a33647a <=( A299  and  a33646a );
 a33648a <=( a33647a  and  a33642a );
 a33652a <=( A167  and  A168 );
 a33653a <=( A169  and  a33652a );
 a33657a <=( (not A203)  and  (not A201) );
 a33658a <=( (not A166)  and  a33657a );
 a33659a <=( a33658a  and  a33653a );
 a33663a <=( A298  and  A266 );
 a33664a <=( A265  and  a33663a );
 a33668a <=( A301  and  A300 );
 a33669a <=( (not A299)  and  a33668a );
 a33670a <=( a33669a  and  a33664a );
 a33674a <=( A167  and  A168 );
 a33675a <=( A169  and  a33674a );
 a33679a <=( (not A203)  and  (not A201) );
 a33680a <=( (not A166)  and  a33679a );
 a33681a <=( a33680a  and  a33675a );
 a33685a <=( A298  and  A266 );
 a33686a <=( A265  and  a33685a );
 a33690a <=( (not A302)  and  A300 );
 a33691a <=( (not A299)  and  a33690a );
 a33692a <=( a33691a  and  a33686a );
 a33696a <=( A167  and  A168 );
 a33697a <=( A169  and  a33696a );
 a33701a <=( (not A203)  and  (not A201) );
 a33702a <=( (not A166)  and  a33701a );
 a33703a <=( a33702a  and  a33697a );
 a33707a <=( (not A298)  and  A266 );
 a33708a <=( A265  and  a33707a );
 a33712a <=( A301  and  A300 );
 a33713a <=( A299  and  a33712a );
 a33714a <=( a33713a  and  a33708a );
 a33718a <=( A167  and  A168 );
 a33719a <=( A169  and  a33718a );
 a33723a <=( (not A203)  and  (not A201) );
 a33724a <=( (not A166)  and  a33723a );
 a33725a <=( a33724a  and  a33719a );
 a33729a <=( (not A298)  and  A266 );
 a33730a <=( A265  and  a33729a );
 a33734a <=( (not A302)  and  A300 );
 a33735a <=( A299  and  a33734a );
 a33736a <=( a33735a  and  a33730a );
 a33740a <=( A167  and  A168 );
 a33741a <=( A169  and  a33740a );
 a33745a <=( (not A203)  and  (not A201) );
 a33746a <=( (not A166)  and  a33745a );
 a33747a <=( a33746a  and  a33741a );
 a33751a <=( A267  and  A266 );
 a33752a <=( (not A265)  and  a33751a );
 a33756a <=( A301  and  (not A300) );
 a33757a <=( A268  and  a33756a );
 a33758a <=( a33757a  and  a33752a );
 a33762a <=( A167  and  A168 );
 a33763a <=( A169  and  a33762a );
 a33767a <=( (not A203)  and  (not A201) );
 a33768a <=( (not A166)  and  a33767a );
 a33769a <=( a33768a  and  a33763a );
 a33773a <=( A267  and  A266 );
 a33774a <=( (not A265)  and  a33773a );
 a33778a <=( (not A302)  and  (not A300) );
 a33779a <=( A268  and  a33778a );
 a33780a <=( a33779a  and  a33774a );
 a33784a <=( A167  and  A168 );
 a33785a <=( A169  and  a33784a );
 a33789a <=( (not A203)  and  (not A201) );
 a33790a <=( (not A166)  and  a33789a );
 a33791a <=( a33790a  and  a33785a );
 a33795a <=( A267  and  A266 );
 a33796a <=( (not A265)  and  a33795a );
 a33800a <=( A299  and  A298 );
 a33801a <=( A268  and  a33800a );
 a33802a <=( a33801a  and  a33796a );
 a33806a <=( A167  and  A168 );
 a33807a <=( A169  and  a33806a );
 a33811a <=( (not A203)  and  (not A201) );
 a33812a <=( (not A166)  and  a33811a );
 a33813a <=( a33812a  and  a33807a );
 a33817a <=( A267  and  A266 );
 a33818a <=( (not A265)  and  a33817a );
 a33822a <=( (not A299)  and  (not A298) );
 a33823a <=( A268  and  a33822a );
 a33824a <=( a33823a  and  a33818a );
 a33828a <=( A167  and  A168 );
 a33829a <=( A169  and  a33828a );
 a33833a <=( (not A203)  and  (not A201) );
 a33834a <=( (not A166)  and  a33833a );
 a33835a <=( a33834a  and  a33829a );
 a33839a <=( A267  and  A266 );
 a33840a <=( (not A265)  and  a33839a );
 a33844a <=( A301  and  (not A300) );
 a33845a <=( (not A269)  and  a33844a );
 a33846a <=( a33845a  and  a33840a );
 a33850a <=( A167  and  A168 );
 a33851a <=( A169  and  a33850a );
 a33855a <=( (not A203)  and  (not A201) );
 a33856a <=( (not A166)  and  a33855a );
 a33857a <=( a33856a  and  a33851a );
 a33861a <=( A267  and  A266 );
 a33862a <=( (not A265)  and  a33861a );
 a33866a <=( (not A302)  and  (not A300) );
 a33867a <=( (not A269)  and  a33866a );
 a33868a <=( a33867a  and  a33862a );
 a33872a <=( A167  and  A168 );
 a33873a <=( A169  and  a33872a );
 a33877a <=( (not A203)  and  (not A201) );
 a33878a <=( (not A166)  and  a33877a );
 a33879a <=( a33878a  and  a33873a );
 a33883a <=( A267  and  A266 );
 a33884a <=( (not A265)  and  a33883a );
 a33888a <=( A299  and  A298 );
 a33889a <=( (not A269)  and  a33888a );
 a33890a <=( a33889a  and  a33884a );
 a33894a <=( A167  and  A168 );
 a33895a <=( A169  and  a33894a );
 a33899a <=( (not A203)  and  (not A201) );
 a33900a <=( (not A166)  and  a33899a );
 a33901a <=( a33900a  and  a33895a );
 a33905a <=( A267  and  A266 );
 a33906a <=( (not A265)  and  a33905a );
 a33910a <=( (not A299)  and  (not A298) );
 a33911a <=( (not A269)  and  a33910a );
 a33912a <=( a33911a  and  a33906a );
 a33916a <=( A167  and  A168 );
 a33917a <=( A169  and  a33916a );
 a33921a <=( (not A203)  and  (not A201) );
 a33922a <=( (not A166)  and  a33921a );
 a33923a <=( a33922a  and  a33917a );
 a33927a <=( A267  and  (not A266) );
 a33928a <=( A265  and  a33927a );
 a33932a <=( A301  and  (not A300) );
 a33933a <=( A268  and  a33932a );
 a33934a <=( a33933a  and  a33928a );
 a33938a <=( A167  and  A168 );
 a33939a <=( A169  and  a33938a );
 a33943a <=( (not A203)  and  (not A201) );
 a33944a <=( (not A166)  and  a33943a );
 a33945a <=( a33944a  and  a33939a );
 a33949a <=( A267  and  (not A266) );
 a33950a <=( A265  and  a33949a );
 a33954a <=( (not A302)  and  (not A300) );
 a33955a <=( A268  and  a33954a );
 a33956a <=( a33955a  and  a33950a );
 a33960a <=( A167  and  A168 );
 a33961a <=( A169  and  a33960a );
 a33965a <=( (not A203)  and  (not A201) );
 a33966a <=( (not A166)  and  a33965a );
 a33967a <=( a33966a  and  a33961a );
 a33971a <=( A267  and  (not A266) );
 a33972a <=( A265  and  a33971a );
 a33976a <=( A299  and  A298 );
 a33977a <=( A268  and  a33976a );
 a33978a <=( a33977a  and  a33972a );
 a33982a <=( A167  and  A168 );
 a33983a <=( A169  and  a33982a );
 a33987a <=( (not A203)  and  (not A201) );
 a33988a <=( (not A166)  and  a33987a );
 a33989a <=( a33988a  and  a33983a );
 a33993a <=( A267  and  (not A266) );
 a33994a <=( A265  and  a33993a );
 a33998a <=( (not A299)  and  (not A298) );
 a33999a <=( A268  and  a33998a );
 a34000a <=( a33999a  and  a33994a );
 a34004a <=( A167  and  A168 );
 a34005a <=( A169  and  a34004a );
 a34009a <=( (not A203)  and  (not A201) );
 a34010a <=( (not A166)  and  a34009a );
 a34011a <=( a34010a  and  a34005a );
 a34015a <=( A267  and  (not A266) );
 a34016a <=( A265  and  a34015a );
 a34020a <=( A301  and  (not A300) );
 a34021a <=( (not A269)  and  a34020a );
 a34022a <=( a34021a  and  a34016a );
 a34026a <=( A167  and  A168 );
 a34027a <=( A169  and  a34026a );
 a34031a <=( (not A203)  and  (not A201) );
 a34032a <=( (not A166)  and  a34031a );
 a34033a <=( a34032a  and  a34027a );
 a34037a <=( A267  and  (not A266) );
 a34038a <=( A265  and  a34037a );
 a34042a <=( (not A302)  and  (not A300) );
 a34043a <=( (not A269)  and  a34042a );
 a34044a <=( a34043a  and  a34038a );
 a34048a <=( A167  and  A168 );
 a34049a <=( A169  and  a34048a );
 a34053a <=( (not A203)  and  (not A201) );
 a34054a <=( (not A166)  and  a34053a );
 a34055a <=( a34054a  and  a34049a );
 a34059a <=( A267  and  (not A266) );
 a34060a <=( A265  and  a34059a );
 a34064a <=( A299  and  A298 );
 a34065a <=( (not A269)  and  a34064a );
 a34066a <=( a34065a  and  a34060a );
 a34070a <=( A167  and  A168 );
 a34071a <=( A169  and  a34070a );
 a34075a <=( (not A203)  and  (not A201) );
 a34076a <=( (not A166)  and  a34075a );
 a34077a <=( a34076a  and  a34071a );
 a34081a <=( A267  and  (not A266) );
 a34082a <=( A265  and  a34081a );
 a34086a <=( (not A299)  and  (not A298) );
 a34087a <=( (not A269)  and  a34086a );
 a34088a <=( a34087a  and  a34082a );
 a34092a <=( A167  and  A168 );
 a34093a <=( A169  and  a34092a );
 a34097a <=( (not A203)  and  (not A201) );
 a34098a <=( (not A166)  and  a34097a );
 a34099a <=( a34098a  and  a34093a );
 a34103a <=( A298  and  (not A266) );
 a34104a <=( (not A265)  and  a34103a );
 a34108a <=( A301  and  A300 );
 a34109a <=( (not A299)  and  a34108a );
 a34110a <=( a34109a  and  a34104a );
 a34114a <=( A167  and  A168 );
 a34115a <=( A169  and  a34114a );
 a34119a <=( (not A203)  and  (not A201) );
 a34120a <=( (not A166)  and  a34119a );
 a34121a <=( a34120a  and  a34115a );
 a34125a <=( A298  and  (not A266) );
 a34126a <=( (not A265)  and  a34125a );
 a34130a <=( (not A302)  and  A300 );
 a34131a <=( (not A299)  and  a34130a );
 a34132a <=( a34131a  and  a34126a );
 a34136a <=( A167  and  A168 );
 a34137a <=( A169  and  a34136a );
 a34141a <=( (not A203)  and  (not A201) );
 a34142a <=( (not A166)  and  a34141a );
 a34143a <=( a34142a  and  a34137a );
 a34147a <=( (not A298)  and  (not A266) );
 a34148a <=( (not A265)  and  a34147a );
 a34152a <=( A301  and  A300 );
 a34153a <=( A299  and  a34152a );
 a34154a <=( a34153a  and  a34148a );
 a34158a <=( A167  and  A168 );
 a34159a <=( A169  and  a34158a );
 a34163a <=( (not A203)  and  (not A201) );
 a34164a <=( (not A166)  and  a34163a );
 a34165a <=( a34164a  and  a34159a );
 a34169a <=( (not A298)  and  (not A266) );
 a34170a <=( (not A265)  and  a34169a );
 a34174a <=( (not A302)  and  A300 );
 a34175a <=( A299  and  a34174a );
 a34176a <=( a34175a  and  a34170a );
 a34180a <=( A167  and  A168 );
 a34181a <=( A169  and  a34180a );
 a34185a <=( A200  and  A199 );
 a34186a <=( (not A166)  and  a34185a );
 a34187a <=( a34186a  and  a34181a );
 a34191a <=( A298  and  A268 );
 a34192a <=( (not A267)  and  a34191a );
 a34196a <=( A301  and  A300 );
 a34197a <=( (not A299)  and  a34196a );
 a34198a <=( a34197a  and  a34192a );
 a34202a <=( A167  and  A168 );
 a34203a <=( A169  and  a34202a );
 a34207a <=( A200  and  A199 );
 a34208a <=( (not A166)  and  a34207a );
 a34209a <=( a34208a  and  a34203a );
 a34213a <=( A298  and  A268 );
 a34214a <=( (not A267)  and  a34213a );
 a34218a <=( (not A302)  and  A300 );
 a34219a <=( (not A299)  and  a34218a );
 a34220a <=( a34219a  and  a34214a );
 a34224a <=( A167  and  A168 );
 a34225a <=( A169  and  a34224a );
 a34229a <=( A200  and  A199 );
 a34230a <=( (not A166)  and  a34229a );
 a34231a <=( a34230a  and  a34225a );
 a34235a <=( (not A298)  and  A268 );
 a34236a <=( (not A267)  and  a34235a );
 a34240a <=( A301  and  A300 );
 a34241a <=( A299  and  a34240a );
 a34242a <=( a34241a  and  a34236a );
 a34246a <=( A167  and  A168 );
 a34247a <=( A169  and  a34246a );
 a34251a <=( A200  and  A199 );
 a34252a <=( (not A166)  and  a34251a );
 a34253a <=( a34252a  and  a34247a );
 a34257a <=( (not A298)  and  A268 );
 a34258a <=( (not A267)  and  a34257a );
 a34262a <=( (not A302)  and  A300 );
 a34263a <=( A299  and  a34262a );
 a34264a <=( a34263a  and  a34258a );
 a34268a <=( A167  and  A168 );
 a34269a <=( A169  and  a34268a );
 a34273a <=( A200  and  A199 );
 a34274a <=( (not A166)  and  a34273a );
 a34275a <=( a34274a  and  a34269a );
 a34279a <=( A298  and  (not A269) );
 a34280a <=( (not A267)  and  a34279a );
 a34284a <=( A301  and  A300 );
 a34285a <=( (not A299)  and  a34284a );
 a34286a <=( a34285a  and  a34280a );
 a34290a <=( A167  and  A168 );
 a34291a <=( A169  and  a34290a );
 a34295a <=( A200  and  A199 );
 a34296a <=( (not A166)  and  a34295a );
 a34297a <=( a34296a  and  a34291a );
 a34301a <=( A298  and  (not A269) );
 a34302a <=( (not A267)  and  a34301a );
 a34306a <=( (not A302)  and  A300 );
 a34307a <=( (not A299)  and  a34306a );
 a34308a <=( a34307a  and  a34302a );
 a34312a <=( A167  and  A168 );
 a34313a <=( A169  and  a34312a );
 a34317a <=( A200  and  A199 );
 a34318a <=( (not A166)  and  a34317a );
 a34319a <=( a34318a  and  a34313a );
 a34323a <=( (not A298)  and  (not A269) );
 a34324a <=( (not A267)  and  a34323a );
 a34328a <=( A301  and  A300 );
 a34329a <=( A299  and  a34328a );
 a34330a <=( a34329a  and  a34324a );
 a34334a <=( A167  and  A168 );
 a34335a <=( A169  and  a34334a );
 a34339a <=( A200  and  A199 );
 a34340a <=( (not A166)  and  a34339a );
 a34341a <=( a34340a  and  a34335a );
 a34345a <=( (not A298)  and  (not A269) );
 a34346a <=( (not A267)  and  a34345a );
 a34350a <=( (not A302)  and  A300 );
 a34351a <=( A299  and  a34350a );
 a34352a <=( a34351a  and  a34346a );
 a34356a <=( A167  and  A168 );
 a34357a <=( A169  and  a34356a );
 a34361a <=( A200  and  A199 );
 a34362a <=( (not A166)  and  a34361a );
 a34363a <=( a34362a  and  a34357a );
 a34367a <=( A298  and  A266 );
 a34368a <=( A265  and  a34367a );
 a34372a <=( A301  and  A300 );
 a34373a <=( (not A299)  and  a34372a );
 a34374a <=( a34373a  and  a34368a );
 a34378a <=( A167  and  A168 );
 a34379a <=( A169  and  a34378a );
 a34383a <=( A200  and  A199 );
 a34384a <=( (not A166)  and  a34383a );
 a34385a <=( a34384a  and  a34379a );
 a34389a <=( A298  and  A266 );
 a34390a <=( A265  and  a34389a );
 a34394a <=( (not A302)  and  A300 );
 a34395a <=( (not A299)  and  a34394a );
 a34396a <=( a34395a  and  a34390a );
 a34400a <=( A167  and  A168 );
 a34401a <=( A169  and  a34400a );
 a34405a <=( A200  and  A199 );
 a34406a <=( (not A166)  and  a34405a );
 a34407a <=( a34406a  and  a34401a );
 a34411a <=( (not A298)  and  A266 );
 a34412a <=( A265  and  a34411a );
 a34416a <=( A301  and  A300 );
 a34417a <=( A299  and  a34416a );
 a34418a <=( a34417a  and  a34412a );
 a34422a <=( A167  and  A168 );
 a34423a <=( A169  and  a34422a );
 a34427a <=( A200  and  A199 );
 a34428a <=( (not A166)  and  a34427a );
 a34429a <=( a34428a  and  a34423a );
 a34433a <=( (not A298)  and  A266 );
 a34434a <=( A265  and  a34433a );
 a34438a <=( (not A302)  and  A300 );
 a34439a <=( A299  and  a34438a );
 a34440a <=( a34439a  and  a34434a );
 a34444a <=( A167  and  A168 );
 a34445a <=( A169  and  a34444a );
 a34449a <=( A200  and  A199 );
 a34450a <=( (not A166)  and  a34449a );
 a34451a <=( a34450a  and  a34445a );
 a34455a <=( A267  and  A266 );
 a34456a <=( (not A265)  and  a34455a );
 a34460a <=( A301  and  (not A300) );
 a34461a <=( A268  and  a34460a );
 a34462a <=( a34461a  and  a34456a );
 a34466a <=( A167  and  A168 );
 a34467a <=( A169  and  a34466a );
 a34471a <=( A200  and  A199 );
 a34472a <=( (not A166)  and  a34471a );
 a34473a <=( a34472a  and  a34467a );
 a34477a <=( A267  and  A266 );
 a34478a <=( (not A265)  and  a34477a );
 a34482a <=( (not A302)  and  (not A300) );
 a34483a <=( A268  and  a34482a );
 a34484a <=( a34483a  and  a34478a );
 a34488a <=( A167  and  A168 );
 a34489a <=( A169  and  a34488a );
 a34493a <=( A200  and  A199 );
 a34494a <=( (not A166)  and  a34493a );
 a34495a <=( a34494a  and  a34489a );
 a34499a <=( A267  and  A266 );
 a34500a <=( (not A265)  and  a34499a );
 a34504a <=( A299  and  A298 );
 a34505a <=( A268  and  a34504a );
 a34506a <=( a34505a  and  a34500a );
 a34510a <=( A167  and  A168 );
 a34511a <=( A169  and  a34510a );
 a34515a <=( A200  and  A199 );
 a34516a <=( (not A166)  and  a34515a );
 a34517a <=( a34516a  and  a34511a );
 a34521a <=( A267  and  A266 );
 a34522a <=( (not A265)  and  a34521a );
 a34526a <=( (not A299)  and  (not A298) );
 a34527a <=( A268  and  a34526a );
 a34528a <=( a34527a  and  a34522a );
 a34532a <=( A167  and  A168 );
 a34533a <=( A169  and  a34532a );
 a34537a <=( A200  and  A199 );
 a34538a <=( (not A166)  and  a34537a );
 a34539a <=( a34538a  and  a34533a );
 a34543a <=( A267  and  A266 );
 a34544a <=( (not A265)  and  a34543a );
 a34548a <=( A301  and  (not A300) );
 a34549a <=( (not A269)  and  a34548a );
 a34550a <=( a34549a  and  a34544a );
 a34554a <=( A167  and  A168 );
 a34555a <=( A169  and  a34554a );
 a34559a <=( A200  and  A199 );
 a34560a <=( (not A166)  and  a34559a );
 a34561a <=( a34560a  and  a34555a );
 a34565a <=( A267  and  A266 );
 a34566a <=( (not A265)  and  a34565a );
 a34570a <=( (not A302)  and  (not A300) );
 a34571a <=( (not A269)  and  a34570a );
 a34572a <=( a34571a  and  a34566a );
 a34576a <=( A167  and  A168 );
 a34577a <=( A169  and  a34576a );
 a34581a <=( A200  and  A199 );
 a34582a <=( (not A166)  and  a34581a );
 a34583a <=( a34582a  and  a34577a );
 a34587a <=( A267  and  A266 );
 a34588a <=( (not A265)  and  a34587a );
 a34592a <=( A299  and  A298 );
 a34593a <=( (not A269)  and  a34592a );
 a34594a <=( a34593a  and  a34588a );
 a34598a <=( A167  and  A168 );
 a34599a <=( A169  and  a34598a );
 a34603a <=( A200  and  A199 );
 a34604a <=( (not A166)  and  a34603a );
 a34605a <=( a34604a  and  a34599a );
 a34609a <=( A267  and  A266 );
 a34610a <=( (not A265)  and  a34609a );
 a34614a <=( (not A299)  and  (not A298) );
 a34615a <=( (not A269)  and  a34614a );
 a34616a <=( a34615a  and  a34610a );
 a34620a <=( A167  and  A168 );
 a34621a <=( A169  and  a34620a );
 a34625a <=( A200  and  A199 );
 a34626a <=( (not A166)  and  a34625a );
 a34627a <=( a34626a  and  a34621a );
 a34631a <=( A267  and  (not A266) );
 a34632a <=( A265  and  a34631a );
 a34636a <=( A301  and  (not A300) );
 a34637a <=( A268  and  a34636a );
 a34638a <=( a34637a  and  a34632a );
 a34642a <=( A167  and  A168 );
 a34643a <=( A169  and  a34642a );
 a34647a <=( A200  and  A199 );
 a34648a <=( (not A166)  and  a34647a );
 a34649a <=( a34648a  and  a34643a );
 a34653a <=( A267  and  (not A266) );
 a34654a <=( A265  and  a34653a );
 a34658a <=( (not A302)  and  (not A300) );
 a34659a <=( A268  and  a34658a );
 a34660a <=( a34659a  and  a34654a );
 a34664a <=( A167  and  A168 );
 a34665a <=( A169  and  a34664a );
 a34669a <=( A200  and  A199 );
 a34670a <=( (not A166)  and  a34669a );
 a34671a <=( a34670a  and  a34665a );
 a34675a <=( A267  and  (not A266) );
 a34676a <=( A265  and  a34675a );
 a34680a <=( A299  and  A298 );
 a34681a <=( A268  and  a34680a );
 a34682a <=( a34681a  and  a34676a );
 a34686a <=( A167  and  A168 );
 a34687a <=( A169  and  a34686a );
 a34691a <=( A200  and  A199 );
 a34692a <=( (not A166)  and  a34691a );
 a34693a <=( a34692a  and  a34687a );
 a34697a <=( A267  and  (not A266) );
 a34698a <=( A265  and  a34697a );
 a34702a <=( (not A299)  and  (not A298) );
 a34703a <=( A268  and  a34702a );
 a34704a <=( a34703a  and  a34698a );
 a34708a <=( A167  and  A168 );
 a34709a <=( A169  and  a34708a );
 a34713a <=( A200  and  A199 );
 a34714a <=( (not A166)  and  a34713a );
 a34715a <=( a34714a  and  a34709a );
 a34719a <=( A267  and  (not A266) );
 a34720a <=( A265  and  a34719a );
 a34724a <=( A301  and  (not A300) );
 a34725a <=( (not A269)  and  a34724a );
 a34726a <=( a34725a  and  a34720a );
 a34730a <=( A167  and  A168 );
 a34731a <=( A169  and  a34730a );
 a34735a <=( A200  and  A199 );
 a34736a <=( (not A166)  and  a34735a );
 a34737a <=( a34736a  and  a34731a );
 a34741a <=( A267  and  (not A266) );
 a34742a <=( A265  and  a34741a );
 a34746a <=( (not A302)  and  (not A300) );
 a34747a <=( (not A269)  and  a34746a );
 a34748a <=( a34747a  and  a34742a );
 a34752a <=( A167  and  A168 );
 a34753a <=( A169  and  a34752a );
 a34757a <=( A200  and  A199 );
 a34758a <=( (not A166)  and  a34757a );
 a34759a <=( a34758a  and  a34753a );
 a34763a <=( A267  and  (not A266) );
 a34764a <=( A265  and  a34763a );
 a34768a <=( A299  and  A298 );
 a34769a <=( (not A269)  and  a34768a );
 a34770a <=( a34769a  and  a34764a );
 a34774a <=( A167  and  A168 );
 a34775a <=( A169  and  a34774a );
 a34779a <=( A200  and  A199 );
 a34780a <=( (not A166)  and  a34779a );
 a34781a <=( a34780a  and  a34775a );
 a34785a <=( A267  and  (not A266) );
 a34786a <=( A265  and  a34785a );
 a34790a <=( (not A299)  and  (not A298) );
 a34791a <=( (not A269)  and  a34790a );
 a34792a <=( a34791a  and  a34786a );
 a34796a <=( A167  and  A168 );
 a34797a <=( A169  and  a34796a );
 a34801a <=( A200  and  A199 );
 a34802a <=( (not A166)  and  a34801a );
 a34803a <=( a34802a  and  a34797a );
 a34807a <=( A298  and  (not A266) );
 a34808a <=( (not A265)  and  a34807a );
 a34812a <=( A301  and  A300 );
 a34813a <=( (not A299)  and  a34812a );
 a34814a <=( a34813a  and  a34808a );
 a34818a <=( A167  and  A168 );
 a34819a <=( A169  and  a34818a );
 a34823a <=( A200  and  A199 );
 a34824a <=( (not A166)  and  a34823a );
 a34825a <=( a34824a  and  a34819a );
 a34829a <=( A298  and  (not A266) );
 a34830a <=( (not A265)  and  a34829a );
 a34834a <=( (not A302)  and  A300 );
 a34835a <=( (not A299)  and  a34834a );
 a34836a <=( a34835a  and  a34830a );
 a34840a <=( A167  and  A168 );
 a34841a <=( A169  and  a34840a );
 a34845a <=( A200  and  A199 );
 a34846a <=( (not A166)  and  a34845a );
 a34847a <=( a34846a  and  a34841a );
 a34851a <=( (not A298)  and  (not A266) );
 a34852a <=( (not A265)  and  a34851a );
 a34856a <=( A301  and  A300 );
 a34857a <=( A299  and  a34856a );
 a34858a <=( a34857a  and  a34852a );
 a34862a <=( A167  and  A168 );
 a34863a <=( A169  and  a34862a );
 a34867a <=( A200  and  A199 );
 a34868a <=( (not A166)  and  a34867a );
 a34869a <=( a34868a  and  a34863a );
 a34873a <=( (not A298)  and  (not A266) );
 a34874a <=( (not A265)  and  a34873a );
 a34878a <=( (not A302)  and  A300 );
 a34879a <=( A299  and  a34878a );
 a34880a <=( a34879a  and  a34874a );
 a34884a <=( A167  and  A168 );
 a34885a <=( A169  and  a34884a );
 a34889a <=( (not A200)  and  (not A199) );
 a34890a <=( (not A166)  and  a34889a );
 a34891a <=( a34890a  and  a34885a );
 a34895a <=( A298  and  A268 );
 a34896a <=( (not A267)  and  a34895a );
 a34900a <=( A301  and  A300 );
 a34901a <=( (not A299)  and  a34900a );
 a34902a <=( a34901a  and  a34896a );
 a34906a <=( A167  and  A168 );
 a34907a <=( A169  and  a34906a );
 a34911a <=( (not A200)  and  (not A199) );
 a34912a <=( (not A166)  and  a34911a );
 a34913a <=( a34912a  and  a34907a );
 a34917a <=( A298  and  A268 );
 a34918a <=( (not A267)  and  a34917a );
 a34922a <=( (not A302)  and  A300 );
 a34923a <=( (not A299)  and  a34922a );
 a34924a <=( a34923a  and  a34918a );
 a34928a <=( A167  and  A168 );
 a34929a <=( A169  and  a34928a );
 a34933a <=( (not A200)  and  (not A199) );
 a34934a <=( (not A166)  and  a34933a );
 a34935a <=( a34934a  and  a34929a );
 a34939a <=( (not A298)  and  A268 );
 a34940a <=( (not A267)  and  a34939a );
 a34944a <=( A301  and  A300 );
 a34945a <=( A299  and  a34944a );
 a34946a <=( a34945a  and  a34940a );
 a34950a <=( A167  and  A168 );
 a34951a <=( A169  and  a34950a );
 a34955a <=( (not A200)  and  (not A199) );
 a34956a <=( (not A166)  and  a34955a );
 a34957a <=( a34956a  and  a34951a );
 a34961a <=( (not A298)  and  A268 );
 a34962a <=( (not A267)  and  a34961a );
 a34966a <=( (not A302)  and  A300 );
 a34967a <=( A299  and  a34966a );
 a34968a <=( a34967a  and  a34962a );
 a34972a <=( A167  and  A168 );
 a34973a <=( A169  and  a34972a );
 a34977a <=( (not A200)  and  (not A199) );
 a34978a <=( (not A166)  and  a34977a );
 a34979a <=( a34978a  and  a34973a );
 a34983a <=( A298  and  (not A269) );
 a34984a <=( (not A267)  and  a34983a );
 a34988a <=( A301  and  A300 );
 a34989a <=( (not A299)  and  a34988a );
 a34990a <=( a34989a  and  a34984a );
 a34994a <=( A167  and  A168 );
 a34995a <=( A169  and  a34994a );
 a34999a <=( (not A200)  and  (not A199) );
 a35000a <=( (not A166)  and  a34999a );
 a35001a <=( a35000a  and  a34995a );
 a35005a <=( A298  and  (not A269) );
 a35006a <=( (not A267)  and  a35005a );
 a35010a <=( (not A302)  and  A300 );
 a35011a <=( (not A299)  and  a35010a );
 a35012a <=( a35011a  and  a35006a );
 a35016a <=( A167  and  A168 );
 a35017a <=( A169  and  a35016a );
 a35021a <=( (not A200)  and  (not A199) );
 a35022a <=( (not A166)  and  a35021a );
 a35023a <=( a35022a  and  a35017a );
 a35027a <=( (not A298)  and  (not A269) );
 a35028a <=( (not A267)  and  a35027a );
 a35032a <=( A301  and  A300 );
 a35033a <=( A299  and  a35032a );
 a35034a <=( a35033a  and  a35028a );
 a35038a <=( A167  and  A168 );
 a35039a <=( A169  and  a35038a );
 a35043a <=( (not A200)  and  (not A199) );
 a35044a <=( (not A166)  and  a35043a );
 a35045a <=( a35044a  and  a35039a );
 a35049a <=( (not A298)  and  (not A269) );
 a35050a <=( (not A267)  and  a35049a );
 a35054a <=( (not A302)  and  A300 );
 a35055a <=( A299  and  a35054a );
 a35056a <=( a35055a  and  a35050a );
 a35060a <=( A167  and  A168 );
 a35061a <=( A169  and  a35060a );
 a35065a <=( (not A200)  and  (not A199) );
 a35066a <=( (not A166)  and  a35065a );
 a35067a <=( a35066a  and  a35061a );
 a35071a <=( A298  and  A266 );
 a35072a <=( A265  and  a35071a );
 a35076a <=( A301  and  A300 );
 a35077a <=( (not A299)  and  a35076a );
 a35078a <=( a35077a  and  a35072a );
 a35082a <=( A167  and  A168 );
 a35083a <=( A169  and  a35082a );
 a35087a <=( (not A200)  and  (not A199) );
 a35088a <=( (not A166)  and  a35087a );
 a35089a <=( a35088a  and  a35083a );
 a35093a <=( A298  and  A266 );
 a35094a <=( A265  and  a35093a );
 a35098a <=( (not A302)  and  A300 );
 a35099a <=( (not A299)  and  a35098a );
 a35100a <=( a35099a  and  a35094a );
 a35104a <=( A167  and  A168 );
 a35105a <=( A169  and  a35104a );
 a35109a <=( (not A200)  and  (not A199) );
 a35110a <=( (not A166)  and  a35109a );
 a35111a <=( a35110a  and  a35105a );
 a35115a <=( (not A298)  and  A266 );
 a35116a <=( A265  and  a35115a );
 a35120a <=( A301  and  A300 );
 a35121a <=( A299  and  a35120a );
 a35122a <=( a35121a  and  a35116a );
 a35126a <=( A167  and  A168 );
 a35127a <=( A169  and  a35126a );
 a35131a <=( (not A200)  and  (not A199) );
 a35132a <=( (not A166)  and  a35131a );
 a35133a <=( a35132a  and  a35127a );
 a35137a <=( (not A298)  and  A266 );
 a35138a <=( A265  and  a35137a );
 a35142a <=( (not A302)  and  A300 );
 a35143a <=( A299  and  a35142a );
 a35144a <=( a35143a  and  a35138a );
 a35148a <=( A167  and  A168 );
 a35149a <=( A169  and  a35148a );
 a35153a <=( (not A200)  and  (not A199) );
 a35154a <=( (not A166)  and  a35153a );
 a35155a <=( a35154a  and  a35149a );
 a35159a <=( A267  and  A266 );
 a35160a <=( (not A265)  and  a35159a );
 a35164a <=( A301  and  (not A300) );
 a35165a <=( A268  and  a35164a );
 a35166a <=( a35165a  and  a35160a );
 a35170a <=( A167  and  A168 );
 a35171a <=( A169  and  a35170a );
 a35175a <=( (not A200)  and  (not A199) );
 a35176a <=( (not A166)  and  a35175a );
 a35177a <=( a35176a  and  a35171a );
 a35181a <=( A267  and  A266 );
 a35182a <=( (not A265)  and  a35181a );
 a35186a <=( (not A302)  and  (not A300) );
 a35187a <=( A268  and  a35186a );
 a35188a <=( a35187a  and  a35182a );
 a35192a <=( A167  and  A168 );
 a35193a <=( A169  and  a35192a );
 a35197a <=( (not A200)  and  (not A199) );
 a35198a <=( (not A166)  and  a35197a );
 a35199a <=( a35198a  and  a35193a );
 a35203a <=( A267  and  A266 );
 a35204a <=( (not A265)  and  a35203a );
 a35208a <=( A299  and  A298 );
 a35209a <=( A268  and  a35208a );
 a35210a <=( a35209a  and  a35204a );
 a35214a <=( A167  and  A168 );
 a35215a <=( A169  and  a35214a );
 a35219a <=( (not A200)  and  (not A199) );
 a35220a <=( (not A166)  and  a35219a );
 a35221a <=( a35220a  and  a35215a );
 a35225a <=( A267  and  A266 );
 a35226a <=( (not A265)  and  a35225a );
 a35230a <=( (not A299)  and  (not A298) );
 a35231a <=( A268  and  a35230a );
 a35232a <=( a35231a  and  a35226a );
 a35236a <=( A167  and  A168 );
 a35237a <=( A169  and  a35236a );
 a35241a <=( (not A200)  and  (not A199) );
 a35242a <=( (not A166)  and  a35241a );
 a35243a <=( a35242a  and  a35237a );
 a35247a <=( A267  and  A266 );
 a35248a <=( (not A265)  and  a35247a );
 a35252a <=( A301  and  (not A300) );
 a35253a <=( (not A269)  and  a35252a );
 a35254a <=( a35253a  and  a35248a );
 a35258a <=( A167  and  A168 );
 a35259a <=( A169  and  a35258a );
 a35263a <=( (not A200)  and  (not A199) );
 a35264a <=( (not A166)  and  a35263a );
 a35265a <=( a35264a  and  a35259a );
 a35269a <=( A267  and  A266 );
 a35270a <=( (not A265)  and  a35269a );
 a35274a <=( (not A302)  and  (not A300) );
 a35275a <=( (not A269)  and  a35274a );
 a35276a <=( a35275a  and  a35270a );
 a35280a <=( A167  and  A168 );
 a35281a <=( A169  and  a35280a );
 a35285a <=( (not A200)  and  (not A199) );
 a35286a <=( (not A166)  and  a35285a );
 a35287a <=( a35286a  and  a35281a );
 a35291a <=( A267  and  A266 );
 a35292a <=( (not A265)  and  a35291a );
 a35296a <=( A299  and  A298 );
 a35297a <=( (not A269)  and  a35296a );
 a35298a <=( a35297a  and  a35292a );
 a35302a <=( A167  and  A168 );
 a35303a <=( A169  and  a35302a );
 a35307a <=( (not A200)  and  (not A199) );
 a35308a <=( (not A166)  and  a35307a );
 a35309a <=( a35308a  and  a35303a );
 a35313a <=( A267  and  A266 );
 a35314a <=( (not A265)  and  a35313a );
 a35318a <=( (not A299)  and  (not A298) );
 a35319a <=( (not A269)  and  a35318a );
 a35320a <=( a35319a  and  a35314a );
 a35324a <=( A167  and  A168 );
 a35325a <=( A169  and  a35324a );
 a35329a <=( (not A200)  and  (not A199) );
 a35330a <=( (not A166)  and  a35329a );
 a35331a <=( a35330a  and  a35325a );
 a35335a <=( A267  and  (not A266) );
 a35336a <=( A265  and  a35335a );
 a35340a <=( A301  and  (not A300) );
 a35341a <=( A268  and  a35340a );
 a35342a <=( a35341a  and  a35336a );
 a35346a <=( A167  and  A168 );
 a35347a <=( A169  and  a35346a );
 a35351a <=( (not A200)  and  (not A199) );
 a35352a <=( (not A166)  and  a35351a );
 a35353a <=( a35352a  and  a35347a );
 a35357a <=( A267  and  (not A266) );
 a35358a <=( A265  and  a35357a );
 a35362a <=( (not A302)  and  (not A300) );
 a35363a <=( A268  and  a35362a );
 a35364a <=( a35363a  and  a35358a );
 a35368a <=( A167  and  A168 );
 a35369a <=( A169  and  a35368a );
 a35373a <=( (not A200)  and  (not A199) );
 a35374a <=( (not A166)  and  a35373a );
 a35375a <=( a35374a  and  a35369a );
 a35379a <=( A267  and  (not A266) );
 a35380a <=( A265  and  a35379a );
 a35384a <=( A299  and  A298 );
 a35385a <=( A268  and  a35384a );
 a35386a <=( a35385a  and  a35380a );
 a35390a <=( A167  and  A168 );
 a35391a <=( A169  and  a35390a );
 a35395a <=( (not A200)  and  (not A199) );
 a35396a <=( (not A166)  and  a35395a );
 a35397a <=( a35396a  and  a35391a );
 a35401a <=( A267  and  (not A266) );
 a35402a <=( A265  and  a35401a );
 a35406a <=( (not A299)  and  (not A298) );
 a35407a <=( A268  and  a35406a );
 a35408a <=( a35407a  and  a35402a );
 a35412a <=( A167  and  A168 );
 a35413a <=( A169  and  a35412a );
 a35417a <=( (not A200)  and  (not A199) );
 a35418a <=( (not A166)  and  a35417a );
 a35419a <=( a35418a  and  a35413a );
 a35423a <=( A267  and  (not A266) );
 a35424a <=( A265  and  a35423a );
 a35428a <=( A301  and  (not A300) );
 a35429a <=( (not A269)  and  a35428a );
 a35430a <=( a35429a  and  a35424a );
 a35434a <=( A167  and  A168 );
 a35435a <=( A169  and  a35434a );
 a35439a <=( (not A200)  and  (not A199) );
 a35440a <=( (not A166)  and  a35439a );
 a35441a <=( a35440a  and  a35435a );
 a35445a <=( A267  and  (not A266) );
 a35446a <=( A265  and  a35445a );
 a35450a <=( (not A302)  and  (not A300) );
 a35451a <=( (not A269)  and  a35450a );
 a35452a <=( a35451a  and  a35446a );
 a35456a <=( A167  and  A168 );
 a35457a <=( A169  and  a35456a );
 a35461a <=( (not A200)  and  (not A199) );
 a35462a <=( (not A166)  and  a35461a );
 a35463a <=( a35462a  and  a35457a );
 a35467a <=( A267  and  (not A266) );
 a35468a <=( A265  and  a35467a );
 a35472a <=( A299  and  A298 );
 a35473a <=( (not A269)  and  a35472a );
 a35474a <=( a35473a  and  a35468a );
 a35478a <=( A167  and  A168 );
 a35479a <=( A169  and  a35478a );
 a35483a <=( (not A200)  and  (not A199) );
 a35484a <=( (not A166)  and  a35483a );
 a35485a <=( a35484a  and  a35479a );
 a35489a <=( A267  and  (not A266) );
 a35490a <=( A265  and  a35489a );
 a35494a <=( (not A299)  and  (not A298) );
 a35495a <=( (not A269)  and  a35494a );
 a35496a <=( a35495a  and  a35490a );
 a35500a <=( A167  and  A168 );
 a35501a <=( A169  and  a35500a );
 a35505a <=( (not A200)  and  (not A199) );
 a35506a <=( (not A166)  and  a35505a );
 a35507a <=( a35506a  and  a35501a );
 a35511a <=( A298  and  (not A266) );
 a35512a <=( (not A265)  and  a35511a );
 a35516a <=( A301  and  A300 );
 a35517a <=( (not A299)  and  a35516a );
 a35518a <=( a35517a  and  a35512a );
 a35522a <=( A167  and  A168 );
 a35523a <=( A169  and  a35522a );
 a35527a <=( (not A200)  and  (not A199) );
 a35528a <=( (not A166)  and  a35527a );
 a35529a <=( a35528a  and  a35523a );
 a35533a <=( A298  and  (not A266) );
 a35534a <=( (not A265)  and  a35533a );
 a35538a <=( (not A302)  and  A300 );
 a35539a <=( (not A299)  and  a35538a );
 a35540a <=( a35539a  and  a35534a );
 a35544a <=( A167  and  A168 );
 a35545a <=( A169  and  a35544a );
 a35549a <=( (not A200)  and  (not A199) );
 a35550a <=( (not A166)  and  a35549a );
 a35551a <=( a35550a  and  a35545a );
 a35555a <=( (not A298)  and  (not A266) );
 a35556a <=( (not A265)  and  a35555a );
 a35560a <=( A301  and  A300 );
 a35561a <=( A299  and  a35560a );
 a35562a <=( a35561a  and  a35556a );
 a35566a <=( A167  and  A168 );
 a35567a <=( A169  and  a35566a );
 a35571a <=( (not A200)  and  (not A199) );
 a35572a <=( (not A166)  and  a35571a );
 a35573a <=( a35572a  and  a35567a );
 a35577a <=( (not A298)  and  (not A266) );
 a35578a <=( (not A265)  and  a35577a );
 a35582a <=( (not A302)  and  A300 );
 a35583a <=( A299  and  a35582a );
 a35584a <=( a35583a  and  a35578a );
 a35588a <=( (not A167)  and  A168 );
 a35589a <=( A169  and  a35588a );
 a35593a <=( A202  and  (not A201) );
 a35594a <=( A166  and  a35593a );
 a35595a <=( a35594a  and  a35589a );
 a35599a <=( A298  and  A268 );
 a35600a <=( (not A267)  and  a35599a );
 a35604a <=( A301  and  A300 );
 a35605a <=( (not A299)  and  a35604a );
 a35606a <=( a35605a  and  a35600a );
 a35610a <=( (not A167)  and  A168 );
 a35611a <=( A169  and  a35610a );
 a35615a <=( A202  and  (not A201) );
 a35616a <=( A166  and  a35615a );
 a35617a <=( a35616a  and  a35611a );
 a35621a <=( A298  and  A268 );
 a35622a <=( (not A267)  and  a35621a );
 a35626a <=( (not A302)  and  A300 );
 a35627a <=( (not A299)  and  a35626a );
 a35628a <=( a35627a  and  a35622a );
 a35632a <=( (not A167)  and  A168 );
 a35633a <=( A169  and  a35632a );
 a35637a <=( A202  and  (not A201) );
 a35638a <=( A166  and  a35637a );
 a35639a <=( a35638a  and  a35633a );
 a35643a <=( (not A298)  and  A268 );
 a35644a <=( (not A267)  and  a35643a );
 a35648a <=( A301  and  A300 );
 a35649a <=( A299  and  a35648a );
 a35650a <=( a35649a  and  a35644a );
 a35654a <=( (not A167)  and  A168 );
 a35655a <=( A169  and  a35654a );
 a35659a <=( A202  and  (not A201) );
 a35660a <=( A166  and  a35659a );
 a35661a <=( a35660a  and  a35655a );
 a35665a <=( (not A298)  and  A268 );
 a35666a <=( (not A267)  and  a35665a );
 a35670a <=( (not A302)  and  A300 );
 a35671a <=( A299  and  a35670a );
 a35672a <=( a35671a  and  a35666a );
 a35676a <=( (not A167)  and  A168 );
 a35677a <=( A169  and  a35676a );
 a35681a <=( A202  and  (not A201) );
 a35682a <=( A166  and  a35681a );
 a35683a <=( a35682a  and  a35677a );
 a35687a <=( A298  and  (not A269) );
 a35688a <=( (not A267)  and  a35687a );
 a35692a <=( A301  and  A300 );
 a35693a <=( (not A299)  and  a35692a );
 a35694a <=( a35693a  and  a35688a );
 a35698a <=( (not A167)  and  A168 );
 a35699a <=( A169  and  a35698a );
 a35703a <=( A202  and  (not A201) );
 a35704a <=( A166  and  a35703a );
 a35705a <=( a35704a  and  a35699a );
 a35709a <=( A298  and  (not A269) );
 a35710a <=( (not A267)  and  a35709a );
 a35714a <=( (not A302)  and  A300 );
 a35715a <=( (not A299)  and  a35714a );
 a35716a <=( a35715a  and  a35710a );
 a35720a <=( (not A167)  and  A168 );
 a35721a <=( A169  and  a35720a );
 a35725a <=( A202  and  (not A201) );
 a35726a <=( A166  and  a35725a );
 a35727a <=( a35726a  and  a35721a );
 a35731a <=( (not A298)  and  (not A269) );
 a35732a <=( (not A267)  and  a35731a );
 a35736a <=( A301  and  A300 );
 a35737a <=( A299  and  a35736a );
 a35738a <=( a35737a  and  a35732a );
 a35742a <=( (not A167)  and  A168 );
 a35743a <=( A169  and  a35742a );
 a35747a <=( A202  and  (not A201) );
 a35748a <=( A166  and  a35747a );
 a35749a <=( a35748a  and  a35743a );
 a35753a <=( (not A298)  and  (not A269) );
 a35754a <=( (not A267)  and  a35753a );
 a35758a <=( (not A302)  and  A300 );
 a35759a <=( A299  and  a35758a );
 a35760a <=( a35759a  and  a35754a );
 a35764a <=( (not A167)  and  A168 );
 a35765a <=( A169  and  a35764a );
 a35769a <=( A202  and  (not A201) );
 a35770a <=( A166  and  a35769a );
 a35771a <=( a35770a  and  a35765a );
 a35775a <=( A298  and  A266 );
 a35776a <=( A265  and  a35775a );
 a35780a <=( A301  and  A300 );
 a35781a <=( (not A299)  and  a35780a );
 a35782a <=( a35781a  and  a35776a );
 a35786a <=( (not A167)  and  A168 );
 a35787a <=( A169  and  a35786a );
 a35791a <=( A202  and  (not A201) );
 a35792a <=( A166  and  a35791a );
 a35793a <=( a35792a  and  a35787a );
 a35797a <=( A298  and  A266 );
 a35798a <=( A265  and  a35797a );
 a35802a <=( (not A302)  and  A300 );
 a35803a <=( (not A299)  and  a35802a );
 a35804a <=( a35803a  and  a35798a );
 a35808a <=( (not A167)  and  A168 );
 a35809a <=( A169  and  a35808a );
 a35813a <=( A202  and  (not A201) );
 a35814a <=( A166  and  a35813a );
 a35815a <=( a35814a  and  a35809a );
 a35819a <=( (not A298)  and  A266 );
 a35820a <=( A265  and  a35819a );
 a35824a <=( A301  and  A300 );
 a35825a <=( A299  and  a35824a );
 a35826a <=( a35825a  and  a35820a );
 a35830a <=( (not A167)  and  A168 );
 a35831a <=( A169  and  a35830a );
 a35835a <=( A202  and  (not A201) );
 a35836a <=( A166  and  a35835a );
 a35837a <=( a35836a  and  a35831a );
 a35841a <=( (not A298)  and  A266 );
 a35842a <=( A265  and  a35841a );
 a35846a <=( (not A302)  and  A300 );
 a35847a <=( A299  and  a35846a );
 a35848a <=( a35847a  and  a35842a );
 a35852a <=( (not A167)  and  A168 );
 a35853a <=( A169  and  a35852a );
 a35857a <=( A202  and  (not A201) );
 a35858a <=( A166  and  a35857a );
 a35859a <=( a35858a  and  a35853a );
 a35863a <=( A267  and  A266 );
 a35864a <=( (not A265)  and  a35863a );
 a35868a <=( A301  and  (not A300) );
 a35869a <=( A268  and  a35868a );
 a35870a <=( a35869a  and  a35864a );
 a35874a <=( (not A167)  and  A168 );
 a35875a <=( A169  and  a35874a );
 a35879a <=( A202  and  (not A201) );
 a35880a <=( A166  and  a35879a );
 a35881a <=( a35880a  and  a35875a );
 a35885a <=( A267  and  A266 );
 a35886a <=( (not A265)  and  a35885a );
 a35890a <=( (not A302)  and  (not A300) );
 a35891a <=( A268  and  a35890a );
 a35892a <=( a35891a  and  a35886a );
 a35896a <=( (not A167)  and  A168 );
 a35897a <=( A169  and  a35896a );
 a35901a <=( A202  and  (not A201) );
 a35902a <=( A166  and  a35901a );
 a35903a <=( a35902a  and  a35897a );
 a35907a <=( A267  and  A266 );
 a35908a <=( (not A265)  and  a35907a );
 a35912a <=( A299  and  A298 );
 a35913a <=( A268  and  a35912a );
 a35914a <=( a35913a  and  a35908a );
 a35918a <=( (not A167)  and  A168 );
 a35919a <=( A169  and  a35918a );
 a35923a <=( A202  and  (not A201) );
 a35924a <=( A166  and  a35923a );
 a35925a <=( a35924a  and  a35919a );
 a35929a <=( A267  and  A266 );
 a35930a <=( (not A265)  and  a35929a );
 a35934a <=( (not A299)  and  (not A298) );
 a35935a <=( A268  and  a35934a );
 a35936a <=( a35935a  and  a35930a );
 a35940a <=( (not A167)  and  A168 );
 a35941a <=( A169  and  a35940a );
 a35945a <=( A202  and  (not A201) );
 a35946a <=( A166  and  a35945a );
 a35947a <=( a35946a  and  a35941a );
 a35951a <=( A267  and  A266 );
 a35952a <=( (not A265)  and  a35951a );
 a35956a <=( A301  and  (not A300) );
 a35957a <=( (not A269)  and  a35956a );
 a35958a <=( a35957a  and  a35952a );
 a35962a <=( (not A167)  and  A168 );
 a35963a <=( A169  and  a35962a );
 a35967a <=( A202  and  (not A201) );
 a35968a <=( A166  and  a35967a );
 a35969a <=( a35968a  and  a35963a );
 a35973a <=( A267  and  A266 );
 a35974a <=( (not A265)  and  a35973a );
 a35978a <=( (not A302)  and  (not A300) );
 a35979a <=( (not A269)  and  a35978a );
 a35980a <=( a35979a  and  a35974a );
 a35984a <=( (not A167)  and  A168 );
 a35985a <=( A169  and  a35984a );
 a35989a <=( A202  and  (not A201) );
 a35990a <=( A166  and  a35989a );
 a35991a <=( a35990a  and  a35985a );
 a35995a <=( A267  and  A266 );
 a35996a <=( (not A265)  and  a35995a );
 a36000a <=( A299  and  A298 );
 a36001a <=( (not A269)  and  a36000a );
 a36002a <=( a36001a  and  a35996a );
 a36006a <=( (not A167)  and  A168 );
 a36007a <=( A169  and  a36006a );
 a36011a <=( A202  and  (not A201) );
 a36012a <=( A166  and  a36011a );
 a36013a <=( a36012a  and  a36007a );
 a36017a <=( A267  and  A266 );
 a36018a <=( (not A265)  and  a36017a );
 a36022a <=( (not A299)  and  (not A298) );
 a36023a <=( (not A269)  and  a36022a );
 a36024a <=( a36023a  and  a36018a );
 a36028a <=( (not A167)  and  A168 );
 a36029a <=( A169  and  a36028a );
 a36033a <=( A202  and  (not A201) );
 a36034a <=( A166  and  a36033a );
 a36035a <=( a36034a  and  a36029a );
 a36039a <=( A267  and  (not A266) );
 a36040a <=( A265  and  a36039a );
 a36044a <=( A301  and  (not A300) );
 a36045a <=( A268  and  a36044a );
 a36046a <=( a36045a  and  a36040a );
 a36050a <=( (not A167)  and  A168 );
 a36051a <=( A169  and  a36050a );
 a36055a <=( A202  and  (not A201) );
 a36056a <=( A166  and  a36055a );
 a36057a <=( a36056a  and  a36051a );
 a36061a <=( A267  and  (not A266) );
 a36062a <=( A265  and  a36061a );
 a36066a <=( (not A302)  and  (not A300) );
 a36067a <=( A268  and  a36066a );
 a36068a <=( a36067a  and  a36062a );
 a36072a <=( (not A167)  and  A168 );
 a36073a <=( A169  and  a36072a );
 a36077a <=( A202  and  (not A201) );
 a36078a <=( A166  and  a36077a );
 a36079a <=( a36078a  and  a36073a );
 a36083a <=( A267  and  (not A266) );
 a36084a <=( A265  and  a36083a );
 a36088a <=( A299  and  A298 );
 a36089a <=( A268  and  a36088a );
 a36090a <=( a36089a  and  a36084a );
 a36094a <=( (not A167)  and  A168 );
 a36095a <=( A169  and  a36094a );
 a36099a <=( A202  and  (not A201) );
 a36100a <=( A166  and  a36099a );
 a36101a <=( a36100a  and  a36095a );
 a36105a <=( A267  and  (not A266) );
 a36106a <=( A265  and  a36105a );
 a36110a <=( (not A299)  and  (not A298) );
 a36111a <=( A268  and  a36110a );
 a36112a <=( a36111a  and  a36106a );
 a36116a <=( (not A167)  and  A168 );
 a36117a <=( A169  and  a36116a );
 a36121a <=( A202  and  (not A201) );
 a36122a <=( A166  and  a36121a );
 a36123a <=( a36122a  and  a36117a );
 a36127a <=( A267  and  (not A266) );
 a36128a <=( A265  and  a36127a );
 a36132a <=( A301  and  (not A300) );
 a36133a <=( (not A269)  and  a36132a );
 a36134a <=( a36133a  and  a36128a );
 a36138a <=( (not A167)  and  A168 );
 a36139a <=( A169  and  a36138a );
 a36143a <=( A202  and  (not A201) );
 a36144a <=( A166  and  a36143a );
 a36145a <=( a36144a  and  a36139a );
 a36149a <=( A267  and  (not A266) );
 a36150a <=( A265  and  a36149a );
 a36154a <=( (not A302)  and  (not A300) );
 a36155a <=( (not A269)  and  a36154a );
 a36156a <=( a36155a  and  a36150a );
 a36160a <=( (not A167)  and  A168 );
 a36161a <=( A169  and  a36160a );
 a36165a <=( A202  and  (not A201) );
 a36166a <=( A166  and  a36165a );
 a36167a <=( a36166a  and  a36161a );
 a36171a <=( A267  and  (not A266) );
 a36172a <=( A265  and  a36171a );
 a36176a <=( A299  and  A298 );
 a36177a <=( (not A269)  and  a36176a );
 a36178a <=( a36177a  and  a36172a );
 a36182a <=( (not A167)  and  A168 );
 a36183a <=( A169  and  a36182a );
 a36187a <=( A202  and  (not A201) );
 a36188a <=( A166  and  a36187a );
 a36189a <=( a36188a  and  a36183a );
 a36193a <=( A267  and  (not A266) );
 a36194a <=( A265  and  a36193a );
 a36198a <=( (not A299)  and  (not A298) );
 a36199a <=( (not A269)  and  a36198a );
 a36200a <=( a36199a  and  a36194a );
 a36204a <=( (not A167)  and  A168 );
 a36205a <=( A169  and  a36204a );
 a36209a <=( A202  and  (not A201) );
 a36210a <=( A166  and  a36209a );
 a36211a <=( a36210a  and  a36205a );
 a36215a <=( A298  and  (not A266) );
 a36216a <=( (not A265)  and  a36215a );
 a36220a <=( A301  and  A300 );
 a36221a <=( (not A299)  and  a36220a );
 a36222a <=( a36221a  and  a36216a );
 a36226a <=( (not A167)  and  A168 );
 a36227a <=( A169  and  a36226a );
 a36231a <=( A202  and  (not A201) );
 a36232a <=( A166  and  a36231a );
 a36233a <=( a36232a  and  a36227a );
 a36237a <=( A298  and  (not A266) );
 a36238a <=( (not A265)  and  a36237a );
 a36242a <=( (not A302)  and  A300 );
 a36243a <=( (not A299)  and  a36242a );
 a36244a <=( a36243a  and  a36238a );
 a36248a <=( (not A167)  and  A168 );
 a36249a <=( A169  and  a36248a );
 a36253a <=( A202  and  (not A201) );
 a36254a <=( A166  and  a36253a );
 a36255a <=( a36254a  and  a36249a );
 a36259a <=( (not A298)  and  (not A266) );
 a36260a <=( (not A265)  and  a36259a );
 a36264a <=( A301  and  A300 );
 a36265a <=( A299  and  a36264a );
 a36266a <=( a36265a  and  a36260a );
 a36270a <=( (not A167)  and  A168 );
 a36271a <=( A169  and  a36270a );
 a36275a <=( A202  and  (not A201) );
 a36276a <=( A166  and  a36275a );
 a36277a <=( a36276a  and  a36271a );
 a36281a <=( (not A298)  and  (not A266) );
 a36282a <=( (not A265)  and  a36281a );
 a36286a <=( (not A302)  and  A300 );
 a36287a <=( A299  and  a36286a );
 a36288a <=( a36287a  and  a36282a );
 a36292a <=( (not A167)  and  A168 );
 a36293a <=( A169  and  a36292a );
 a36297a <=( (not A203)  and  (not A201) );
 a36298a <=( A166  and  a36297a );
 a36299a <=( a36298a  and  a36293a );
 a36303a <=( A298  and  A268 );
 a36304a <=( (not A267)  and  a36303a );
 a36308a <=( A301  and  A300 );
 a36309a <=( (not A299)  and  a36308a );
 a36310a <=( a36309a  and  a36304a );
 a36314a <=( (not A167)  and  A168 );
 a36315a <=( A169  and  a36314a );
 a36319a <=( (not A203)  and  (not A201) );
 a36320a <=( A166  and  a36319a );
 a36321a <=( a36320a  and  a36315a );
 a36325a <=( A298  and  A268 );
 a36326a <=( (not A267)  and  a36325a );
 a36330a <=( (not A302)  and  A300 );
 a36331a <=( (not A299)  and  a36330a );
 a36332a <=( a36331a  and  a36326a );
 a36336a <=( (not A167)  and  A168 );
 a36337a <=( A169  and  a36336a );
 a36341a <=( (not A203)  and  (not A201) );
 a36342a <=( A166  and  a36341a );
 a36343a <=( a36342a  and  a36337a );
 a36347a <=( (not A298)  and  A268 );
 a36348a <=( (not A267)  and  a36347a );
 a36352a <=( A301  and  A300 );
 a36353a <=( A299  and  a36352a );
 a36354a <=( a36353a  and  a36348a );
 a36358a <=( (not A167)  and  A168 );
 a36359a <=( A169  and  a36358a );
 a36363a <=( (not A203)  and  (not A201) );
 a36364a <=( A166  and  a36363a );
 a36365a <=( a36364a  and  a36359a );
 a36369a <=( (not A298)  and  A268 );
 a36370a <=( (not A267)  and  a36369a );
 a36374a <=( (not A302)  and  A300 );
 a36375a <=( A299  and  a36374a );
 a36376a <=( a36375a  and  a36370a );
 a36380a <=( (not A167)  and  A168 );
 a36381a <=( A169  and  a36380a );
 a36385a <=( (not A203)  and  (not A201) );
 a36386a <=( A166  and  a36385a );
 a36387a <=( a36386a  and  a36381a );
 a36391a <=( A298  and  (not A269) );
 a36392a <=( (not A267)  and  a36391a );
 a36396a <=( A301  and  A300 );
 a36397a <=( (not A299)  and  a36396a );
 a36398a <=( a36397a  and  a36392a );
 a36402a <=( (not A167)  and  A168 );
 a36403a <=( A169  and  a36402a );
 a36407a <=( (not A203)  and  (not A201) );
 a36408a <=( A166  and  a36407a );
 a36409a <=( a36408a  and  a36403a );
 a36413a <=( A298  and  (not A269) );
 a36414a <=( (not A267)  and  a36413a );
 a36418a <=( (not A302)  and  A300 );
 a36419a <=( (not A299)  and  a36418a );
 a36420a <=( a36419a  and  a36414a );
 a36424a <=( (not A167)  and  A168 );
 a36425a <=( A169  and  a36424a );
 a36429a <=( (not A203)  and  (not A201) );
 a36430a <=( A166  and  a36429a );
 a36431a <=( a36430a  and  a36425a );
 a36435a <=( (not A298)  and  (not A269) );
 a36436a <=( (not A267)  and  a36435a );
 a36440a <=( A301  and  A300 );
 a36441a <=( A299  and  a36440a );
 a36442a <=( a36441a  and  a36436a );
 a36446a <=( (not A167)  and  A168 );
 a36447a <=( A169  and  a36446a );
 a36451a <=( (not A203)  and  (not A201) );
 a36452a <=( A166  and  a36451a );
 a36453a <=( a36452a  and  a36447a );
 a36457a <=( (not A298)  and  (not A269) );
 a36458a <=( (not A267)  and  a36457a );
 a36462a <=( (not A302)  and  A300 );
 a36463a <=( A299  and  a36462a );
 a36464a <=( a36463a  and  a36458a );
 a36468a <=( (not A167)  and  A168 );
 a36469a <=( A169  and  a36468a );
 a36473a <=( (not A203)  and  (not A201) );
 a36474a <=( A166  and  a36473a );
 a36475a <=( a36474a  and  a36469a );
 a36479a <=( A298  and  A266 );
 a36480a <=( A265  and  a36479a );
 a36484a <=( A301  and  A300 );
 a36485a <=( (not A299)  and  a36484a );
 a36486a <=( a36485a  and  a36480a );
 a36490a <=( (not A167)  and  A168 );
 a36491a <=( A169  and  a36490a );
 a36495a <=( (not A203)  and  (not A201) );
 a36496a <=( A166  and  a36495a );
 a36497a <=( a36496a  and  a36491a );
 a36501a <=( A298  and  A266 );
 a36502a <=( A265  and  a36501a );
 a36506a <=( (not A302)  and  A300 );
 a36507a <=( (not A299)  and  a36506a );
 a36508a <=( a36507a  and  a36502a );
 a36512a <=( (not A167)  and  A168 );
 a36513a <=( A169  and  a36512a );
 a36517a <=( (not A203)  and  (not A201) );
 a36518a <=( A166  and  a36517a );
 a36519a <=( a36518a  and  a36513a );
 a36523a <=( (not A298)  and  A266 );
 a36524a <=( A265  and  a36523a );
 a36528a <=( A301  and  A300 );
 a36529a <=( A299  and  a36528a );
 a36530a <=( a36529a  and  a36524a );
 a36534a <=( (not A167)  and  A168 );
 a36535a <=( A169  and  a36534a );
 a36539a <=( (not A203)  and  (not A201) );
 a36540a <=( A166  and  a36539a );
 a36541a <=( a36540a  and  a36535a );
 a36545a <=( (not A298)  and  A266 );
 a36546a <=( A265  and  a36545a );
 a36550a <=( (not A302)  and  A300 );
 a36551a <=( A299  and  a36550a );
 a36552a <=( a36551a  and  a36546a );
 a36556a <=( (not A167)  and  A168 );
 a36557a <=( A169  and  a36556a );
 a36561a <=( (not A203)  and  (not A201) );
 a36562a <=( A166  and  a36561a );
 a36563a <=( a36562a  and  a36557a );
 a36567a <=( A267  and  A266 );
 a36568a <=( (not A265)  and  a36567a );
 a36572a <=( A301  and  (not A300) );
 a36573a <=( A268  and  a36572a );
 a36574a <=( a36573a  and  a36568a );
 a36578a <=( (not A167)  and  A168 );
 a36579a <=( A169  and  a36578a );
 a36583a <=( (not A203)  and  (not A201) );
 a36584a <=( A166  and  a36583a );
 a36585a <=( a36584a  and  a36579a );
 a36589a <=( A267  and  A266 );
 a36590a <=( (not A265)  and  a36589a );
 a36594a <=( (not A302)  and  (not A300) );
 a36595a <=( A268  and  a36594a );
 a36596a <=( a36595a  and  a36590a );
 a36600a <=( (not A167)  and  A168 );
 a36601a <=( A169  and  a36600a );
 a36605a <=( (not A203)  and  (not A201) );
 a36606a <=( A166  and  a36605a );
 a36607a <=( a36606a  and  a36601a );
 a36611a <=( A267  and  A266 );
 a36612a <=( (not A265)  and  a36611a );
 a36616a <=( A299  and  A298 );
 a36617a <=( A268  and  a36616a );
 a36618a <=( a36617a  and  a36612a );
 a36622a <=( (not A167)  and  A168 );
 a36623a <=( A169  and  a36622a );
 a36627a <=( (not A203)  and  (not A201) );
 a36628a <=( A166  and  a36627a );
 a36629a <=( a36628a  and  a36623a );
 a36633a <=( A267  and  A266 );
 a36634a <=( (not A265)  and  a36633a );
 a36638a <=( (not A299)  and  (not A298) );
 a36639a <=( A268  and  a36638a );
 a36640a <=( a36639a  and  a36634a );
 a36644a <=( (not A167)  and  A168 );
 a36645a <=( A169  and  a36644a );
 a36649a <=( (not A203)  and  (not A201) );
 a36650a <=( A166  and  a36649a );
 a36651a <=( a36650a  and  a36645a );
 a36655a <=( A267  and  A266 );
 a36656a <=( (not A265)  and  a36655a );
 a36660a <=( A301  and  (not A300) );
 a36661a <=( (not A269)  and  a36660a );
 a36662a <=( a36661a  and  a36656a );
 a36666a <=( (not A167)  and  A168 );
 a36667a <=( A169  and  a36666a );
 a36671a <=( (not A203)  and  (not A201) );
 a36672a <=( A166  and  a36671a );
 a36673a <=( a36672a  and  a36667a );
 a36677a <=( A267  and  A266 );
 a36678a <=( (not A265)  and  a36677a );
 a36682a <=( (not A302)  and  (not A300) );
 a36683a <=( (not A269)  and  a36682a );
 a36684a <=( a36683a  and  a36678a );
 a36688a <=( (not A167)  and  A168 );
 a36689a <=( A169  and  a36688a );
 a36693a <=( (not A203)  and  (not A201) );
 a36694a <=( A166  and  a36693a );
 a36695a <=( a36694a  and  a36689a );
 a36699a <=( A267  and  A266 );
 a36700a <=( (not A265)  and  a36699a );
 a36704a <=( A299  and  A298 );
 a36705a <=( (not A269)  and  a36704a );
 a36706a <=( a36705a  and  a36700a );
 a36710a <=( (not A167)  and  A168 );
 a36711a <=( A169  and  a36710a );
 a36715a <=( (not A203)  and  (not A201) );
 a36716a <=( A166  and  a36715a );
 a36717a <=( a36716a  and  a36711a );
 a36721a <=( A267  and  A266 );
 a36722a <=( (not A265)  and  a36721a );
 a36726a <=( (not A299)  and  (not A298) );
 a36727a <=( (not A269)  and  a36726a );
 a36728a <=( a36727a  and  a36722a );
 a36732a <=( (not A167)  and  A168 );
 a36733a <=( A169  and  a36732a );
 a36737a <=( (not A203)  and  (not A201) );
 a36738a <=( A166  and  a36737a );
 a36739a <=( a36738a  and  a36733a );
 a36743a <=( A267  and  (not A266) );
 a36744a <=( A265  and  a36743a );
 a36748a <=( A301  and  (not A300) );
 a36749a <=( A268  and  a36748a );
 a36750a <=( a36749a  and  a36744a );
 a36754a <=( (not A167)  and  A168 );
 a36755a <=( A169  and  a36754a );
 a36759a <=( (not A203)  and  (not A201) );
 a36760a <=( A166  and  a36759a );
 a36761a <=( a36760a  and  a36755a );
 a36765a <=( A267  and  (not A266) );
 a36766a <=( A265  and  a36765a );
 a36770a <=( (not A302)  and  (not A300) );
 a36771a <=( A268  and  a36770a );
 a36772a <=( a36771a  and  a36766a );
 a36776a <=( (not A167)  and  A168 );
 a36777a <=( A169  and  a36776a );
 a36781a <=( (not A203)  and  (not A201) );
 a36782a <=( A166  and  a36781a );
 a36783a <=( a36782a  and  a36777a );
 a36787a <=( A267  and  (not A266) );
 a36788a <=( A265  and  a36787a );
 a36792a <=( A299  and  A298 );
 a36793a <=( A268  and  a36792a );
 a36794a <=( a36793a  and  a36788a );
 a36798a <=( (not A167)  and  A168 );
 a36799a <=( A169  and  a36798a );
 a36803a <=( (not A203)  and  (not A201) );
 a36804a <=( A166  and  a36803a );
 a36805a <=( a36804a  and  a36799a );
 a36809a <=( A267  and  (not A266) );
 a36810a <=( A265  and  a36809a );
 a36814a <=( (not A299)  and  (not A298) );
 a36815a <=( A268  and  a36814a );
 a36816a <=( a36815a  and  a36810a );
 a36820a <=( (not A167)  and  A168 );
 a36821a <=( A169  and  a36820a );
 a36825a <=( (not A203)  and  (not A201) );
 a36826a <=( A166  and  a36825a );
 a36827a <=( a36826a  and  a36821a );
 a36831a <=( A267  and  (not A266) );
 a36832a <=( A265  and  a36831a );
 a36836a <=( A301  and  (not A300) );
 a36837a <=( (not A269)  and  a36836a );
 a36838a <=( a36837a  and  a36832a );
 a36842a <=( (not A167)  and  A168 );
 a36843a <=( A169  and  a36842a );
 a36847a <=( (not A203)  and  (not A201) );
 a36848a <=( A166  and  a36847a );
 a36849a <=( a36848a  and  a36843a );
 a36853a <=( A267  and  (not A266) );
 a36854a <=( A265  and  a36853a );
 a36858a <=( (not A302)  and  (not A300) );
 a36859a <=( (not A269)  and  a36858a );
 a36860a <=( a36859a  and  a36854a );
 a36864a <=( (not A167)  and  A168 );
 a36865a <=( A169  and  a36864a );
 a36869a <=( (not A203)  and  (not A201) );
 a36870a <=( A166  and  a36869a );
 a36871a <=( a36870a  and  a36865a );
 a36875a <=( A267  and  (not A266) );
 a36876a <=( A265  and  a36875a );
 a36880a <=( A299  and  A298 );
 a36881a <=( (not A269)  and  a36880a );
 a36882a <=( a36881a  and  a36876a );
 a36886a <=( (not A167)  and  A168 );
 a36887a <=( A169  and  a36886a );
 a36891a <=( (not A203)  and  (not A201) );
 a36892a <=( A166  and  a36891a );
 a36893a <=( a36892a  and  a36887a );
 a36897a <=( A267  and  (not A266) );
 a36898a <=( A265  and  a36897a );
 a36902a <=( (not A299)  and  (not A298) );
 a36903a <=( (not A269)  and  a36902a );
 a36904a <=( a36903a  and  a36898a );
 a36908a <=( (not A167)  and  A168 );
 a36909a <=( A169  and  a36908a );
 a36913a <=( (not A203)  and  (not A201) );
 a36914a <=( A166  and  a36913a );
 a36915a <=( a36914a  and  a36909a );
 a36919a <=( A298  and  (not A266) );
 a36920a <=( (not A265)  and  a36919a );
 a36924a <=( A301  and  A300 );
 a36925a <=( (not A299)  and  a36924a );
 a36926a <=( a36925a  and  a36920a );
 a36930a <=( (not A167)  and  A168 );
 a36931a <=( A169  and  a36930a );
 a36935a <=( (not A203)  and  (not A201) );
 a36936a <=( A166  and  a36935a );
 a36937a <=( a36936a  and  a36931a );
 a36941a <=( A298  and  (not A266) );
 a36942a <=( (not A265)  and  a36941a );
 a36946a <=( (not A302)  and  A300 );
 a36947a <=( (not A299)  and  a36946a );
 a36948a <=( a36947a  and  a36942a );
 a36952a <=( (not A167)  and  A168 );
 a36953a <=( A169  and  a36952a );
 a36957a <=( (not A203)  and  (not A201) );
 a36958a <=( A166  and  a36957a );
 a36959a <=( a36958a  and  a36953a );
 a36963a <=( (not A298)  and  (not A266) );
 a36964a <=( (not A265)  and  a36963a );
 a36968a <=( A301  and  A300 );
 a36969a <=( A299  and  a36968a );
 a36970a <=( a36969a  and  a36964a );
 a36974a <=( (not A167)  and  A168 );
 a36975a <=( A169  and  a36974a );
 a36979a <=( (not A203)  and  (not A201) );
 a36980a <=( A166  and  a36979a );
 a36981a <=( a36980a  and  a36975a );
 a36985a <=( (not A298)  and  (not A266) );
 a36986a <=( (not A265)  and  a36985a );
 a36990a <=( (not A302)  and  A300 );
 a36991a <=( A299  and  a36990a );
 a36992a <=( a36991a  and  a36986a );
 a36996a <=( (not A167)  and  A168 );
 a36997a <=( A169  and  a36996a );
 a37001a <=( A200  and  A199 );
 a37002a <=( A166  and  a37001a );
 a37003a <=( a37002a  and  a36997a );
 a37007a <=( A298  and  A268 );
 a37008a <=( (not A267)  and  a37007a );
 a37012a <=( A301  and  A300 );
 a37013a <=( (not A299)  and  a37012a );
 a37014a <=( a37013a  and  a37008a );
 a37018a <=( (not A167)  and  A168 );
 a37019a <=( A169  and  a37018a );
 a37023a <=( A200  and  A199 );
 a37024a <=( A166  and  a37023a );
 a37025a <=( a37024a  and  a37019a );
 a37029a <=( A298  and  A268 );
 a37030a <=( (not A267)  and  a37029a );
 a37034a <=( (not A302)  and  A300 );
 a37035a <=( (not A299)  and  a37034a );
 a37036a <=( a37035a  and  a37030a );
 a37040a <=( (not A167)  and  A168 );
 a37041a <=( A169  and  a37040a );
 a37045a <=( A200  and  A199 );
 a37046a <=( A166  and  a37045a );
 a37047a <=( a37046a  and  a37041a );
 a37051a <=( (not A298)  and  A268 );
 a37052a <=( (not A267)  and  a37051a );
 a37056a <=( A301  and  A300 );
 a37057a <=( A299  and  a37056a );
 a37058a <=( a37057a  and  a37052a );
 a37062a <=( (not A167)  and  A168 );
 a37063a <=( A169  and  a37062a );
 a37067a <=( A200  and  A199 );
 a37068a <=( A166  and  a37067a );
 a37069a <=( a37068a  and  a37063a );
 a37073a <=( (not A298)  and  A268 );
 a37074a <=( (not A267)  and  a37073a );
 a37078a <=( (not A302)  and  A300 );
 a37079a <=( A299  and  a37078a );
 a37080a <=( a37079a  and  a37074a );
 a37084a <=( (not A167)  and  A168 );
 a37085a <=( A169  and  a37084a );
 a37089a <=( A200  and  A199 );
 a37090a <=( A166  and  a37089a );
 a37091a <=( a37090a  and  a37085a );
 a37095a <=( A298  and  (not A269) );
 a37096a <=( (not A267)  and  a37095a );
 a37100a <=( A301  and  A300 );
 a37101a <=( (not A299)  and  a37100a );
 a37102a <=( a37101a  and  a37096a );
 a37106a <=( (not A167)  and  A168 );
 a37107a <=( A169  and  a37106a );
 a37111a <=( A200  and  A199 );
 a37112a <=( A166  and  a37111a );
 a37113a <=( a37112a  and  a37107a );
 a37117a <=( A298  and  (not A269) );
 a37118a <=( (not A267)  and  a37117a );
 a37122a <=( (not A302)  and  A300 );
 a37123a <=( (not A299)  and  a37122a );
 a37124a <=( a37123a  and  a37118a );
 a37128a <=( (not A167)  and  A168 );
 a37129a <=( A169  and  a37128a );
 a37133a <=( A200  and  A199 );
 a37134a <=( A166  and  a37133a );
 a37135a <=( a37134a  and  a37129a );
 a37139a <=( (not A298)  and  (not A269) );
 a37140a <=( (not A267)  and  a37139a );
 a37144a <=( A301  and  A300 );
 a37145a <=( A299  and  a37144a );
 a37146a <=( a37145a  and  a37140a );
 a37150a <=( (not A167)  and  A168 );
 a37151a <=( A169  and  a37150a );
 a37155a <=( A200  and  A199 );
 a37156a <=( A166  and  a37155a );
 a37157a <=( a37156a  and  a37151a );
 a37161a <=( (not A298)  and  (not A269) );
 a37162a <=( (not A267)  and  a37161a );
 a37166a <=( (not A302)  and  A300 );
 a37167a <=( A299  and  a37166a );
 a37168a <=( a37167a  and  a37162a );
 a37172a <=( (not A167)  and  A168 );
 a37173a <=( A169  and  a37172a );
 a37177a <=( A200  and  A199 );
 a37178a <=( A166  and  a37177a );
 a37179a <=( a37178a  and  a37173a );
 a37183a <=( A298  and  A266 );
 a37184a <=( A265  and  a37183a );
 a37188a <=( A301  and  A300 );
 a37189a <=( (not A299)  and  a37188a );
 a37190a <=( a37189a  and  a37184a );
 a37194a <=( (not A167)  and  A168 );
 a37195a <=( A169  and  a37194a );
 a37199a <=( A200  and  A199 );
 a37200a <=( A166  and  a37199a );
 a37201a <=( a37200a  and  a37195a );
 a37205a <=( A298  and  A266 );
 a37206a <=( A265  and  a37205a );
 a37210a <=( (not A302)  and  A300 );
 a37211a <=( (not A299)  and  a37210a );
 a37212a <=( a37211a  and  a37206a );
 a37216a <=( (not A167)  and  A168 );
 a37217a <=( A169  and  a37216a );
 a37221a <=( A200  and  A199 );
 a37222a <=( A166  and  a37221a );
 a37223a <=( a37222a  and  a37217a );
 a37227a <=( (not A298)  and  A266 );
 a37228a <=( A265  and  a37227a );
 a37232a <=( A301  and  A300 );
 a37233a <=( A299  and  a37232a );
 a37234a <=( a37233a  and  a37228a );
 a37238a <=( (not A167)  and  A168 );
 a37239a <=( A169  and  a37238a );
 a37243a <=( A200  and  A199 );
 a37244a <=( A166  and  a37243a );
 a37245a <=( a37244a  and  a37239a );
 a37249a <=( (not A298)  and  A266 );
 a37250a <=( A265  and  a37249a );
 a37254a <=( (not A302)  and  A300 );
 a37255a <=( A299  and  a37254a );
 a37256a <=( a37255a  and  a37250a );
 a37260a <=( (not A167)  and  A168 );
 a37261a <=( A169  and  a37260a );
 a37265a <=( A200  and  A199 );
 a37266a <=( A166  and  a37265a );
 a37267a <=( a37266a  and  a37261a );
 a37271a <=( A267  and  A266 );
 a37272a <=( (not A265)  and  a37271a );
 a37276a <=( A301  and  (not A300) );
 a37277a <=( A268  and  a37276a );
 a37278a <=( a37277a  and  a37272a );
 a37282a <=( (not A167)  and  A168 );
 a37283a <=( A169  and  a37282a );
 a37287a <=( A200  and  A199 );
 a37288a <=( A166  and  a37287a );
 a37289a <=( a37288a  and  a37283a );
 a37293a <=( A267  and  A266 );
 a37294a <=( (not A265)  and  a37293a );
 a37298a <=( (not A302)  and  (not A300) );
 a37299a <=( A268  and  a37298a );
 a37300a <=( a37299a  and  a37294a );
 a37304a <=( (not A167)  and  A168 );
 a37305a <=( A169  and  a37304a );
 a37309a <=( A200  and  A199 );
 a37310a <=( A166  and  a37309a );
 a37311a <=( a37310a  and  a37305a );
 a37315a <=( A267  and  A266 );
 a37316a <=( (not A265)  and  a37315a );
 a37320a <=( A299  and  A298 );
 a37321a <=( A268  and  a37320a );
 a37322a <=( a37321a  and  a37316a );
 a37326a <=( (not A167)  and  A168 );
 a37327a <=( A169  and  a37326a );
 a37331a <=( A200  and  A199 );
 a37332a <=( A166  and  a37331a );
 a37333a <=( a37332a  and  a37327a );
 a37337a <=( A267  and  A266 );
 a37338a <=( (not A265)  and  a37337a );
 a37342a <=( (not A299)  and  (not A298) );
 a37343a <=( A268  and  a37342a );
 a37344a <=( a37343a  and  a37338a );
 a37348a <=( (not A167)  and  A168 );
 a37349a <=( A169  and  a37348a );
 a37353a <=( A200  and  A199 );
 a37354a <=( A166  and  a37353a );
 a37355a <=( a37354a  and  a37349a );
 a37359a <=( A267  and  A266 );
 a37360a <=( (not A265)  and  a37359a );
 a37364a <=( A301  and  (not A300) );
 a37365a <=( (not A269)  and  a37364a );
 a37366a <=( a37365a  and  a37360a );
 a37370a <=( (not A167)  and  A168 );
 a37371a <=( A169  and  a37370a );
 a37375a <=( A200  and  A199 );
 a37376a <=( A166  and  a37375a );
 a37377a <=( a37376a  and  a37371a );
 a37381a <=( A267  and  A266 );
 a37382a <=( (not A265)  and  a37381a );
 a37386a <=( (not A302)  and  (not A300) );
 a37387a <=( (not A269)  and  a37386a );
 a37388a <=( a37387a  and  a37382a );
 a37392a <=( (not A167)  and  A168 );
 a37393a <=( A169  and  a37392a );
 a37397a <=( A200  and  A199 );
 a37398a <=( A166  and  a37397a );
 a37399a <=( a37398a  and  a37393a );
 a37403a <=( A267  and  A266 );
 a37404a <=( (not A265)  and  a37403a );
 a37408a <=( A299  and  A298 );
 a37409a <=( (not A269)  and  a37408a );
 a37410a <=( a37409a  and  a37404a );
 a37414a <=( (not A167)  and  A168 );
 a37415a <=( A169  and  a37414a );
 a37419a <=( A200  and  A199 );
 a37420a <=( A166  and  a37419a );
 a37421a <=( a37420a  and  a37415a );
 a37425a <=( A267  and  A266 );
 a37426a <=( (not A265)  and  a37425a );
 a37430a <=( (not A299)  and  (not A298) );
 a37431a <=( (not A269)  and  a37430a );
 a37432a <=( a37431a  and  a37426a );
 a37436a <=( (not A167)  and  A168 );
 a37437a <=( A169  and  a37436a );
 a37441a <=( A200  and  A199 );
 a37442a <=( A166  and  a37441a );
 a37443a <=( a37442a  and  a37437a );
 a37447a <=( A267  and  (not A266) );
 a37448a <=( A265  and  a37447a );
 a37452a <=( A301  and  (not A300) );
 a37453a <=( A268  and  a37452a );
 a37454a <=( a37453a  and  a37448a );
 a37458a <=( (not A167)  and  A168 );
 a37459a <=( A169  and  a37458a );
 a37463a <=( A200  and  A199 );
 a37464a <=( A166  and  a37463a );
 a37465a <=( a37464a  and  a37459a );
 a37469a <=( A267  and  (not A266) );
 a37470a <=( A265  and  a37469a );
 a37474a <=( (not A302)  and  (not A300) );
 a37475a <=( A268  and  a37474a );
 a37476a <=( a37475a  and  a37470a );
 a37480a <=( (not A167)  and  A168 );
 a37481a <=( A169  and  a37480a );
 a37485a <=( A200  and  A199 );
 a37486a <=( A166  and  a37485a );
 a37487a <=( a37486a  and  a37481a );
 a37491a <=( A267  and  (not A266) );
 a37492a <=( A265  and  a37491a );
 a37496a <=( A299  and  A298 );
 a37497a <=( A268  and  a37496a );
 a37498a <=( a37497a  and  a37492a );
 a37502a <=( (not A167)  and  A168 );
 a37503a <=( A169  and  a37502a );
 a37507a <=( A200  and  A199 );
 a37508a <=( A166  and  a37507a );
 a37509a <=( a37508a  and  a37503a );
 a37513a <=( A267  and  (not A266) );
 a37514a <=( A265  and  a37513a );
 a37518a <=( (not A299)  and  (not A298) );
 a37519a <=( A268  and  a37518a );
 a37520a <=( a37519a  and  a37514a );
 a37524a <=( (not A167)  and  A168 );
 a37525a <=( A169  and  a37524a );
 a37529a <=( A200  and  A199 );
 a37530a <=( A166  and  a37529a );
 a37531a <=( a37530a  and  a37525a );
 a37535a <=( A267  and  (not A266) );
 a37536a <=( A265  and  a37535a );
 a37540a <=( A301  and  (not A300) );
 a37541a <=( (not A269)  and  a37540a );
 a37542a <=( a37541a  and  a37536a );
 a37546a <=( (not A167)  and  A168 );
 a37547a <=( A169  and  a37546a );
 a37551a <=( A200  and  A199 );
 a37552a <=( A166  and  a37551a );
 a37553a <=( a37552a  and  a37547a );
 a37557a <=( A267  and  (not A266) );
 a37558a <=( A265  and  a37557a );
 a37562a <=( (not A302)  and  (not A300) );
 a37563a <=( (not A269)  and  a37562a );
 a37564a <=( a37563a  and  a37558a );
 a37568a <=( (not A167)  and  A168 );
 a37569a <=( A169  and  a37568a );
 a37573a <=( A200  and  A199 );
 a37574a <=( A166  and  a37573a );
 a37575a <=( a37574a  and  a37569a );
 a37579a <=( A267  and  (not A266) );
 a37580a <=( A265  and  a37579a );
 a37584a <=( A299  and  A298 );
 a37585a <=( (not A269)  and  a37584a );
 a37586a <=( a37585a  and  a37580a );
 a37590a <=( (not A167)  and  A168 );
 a37591a <=( A169  and  a37590a );
 a37595a <=( A200  and  A199 );
 a37596a <=( A166  and  a37595a );
 a37597a <=( a37596a  and  a37591a );
 a37601a <=( A267  and  (not A266) );
 a37602a <=( A265  and  a37601a );
 a37606a <=( (not A299)  and  (not A298) );
 a37607a <=( (not A269)  and  a37606a );
 a37608a <=( a37607a  and  a37602a );
 a37612a <=( (not A167)  and  A168 );
 a37613a <=( A169  and  a37612a );
 a37617a <=( A200  and  A199 );
 a37618a <=( A166  and  a37617a );
 a37619a <=( a37618a  and  a37613a );
 a37623a <=( A298  and  (not A266) );
 a37624a <=( (not A265)  and  a37623a );
 a37628a <=( A301  and  A300 );
 a37629a <=( (not A299)  and  a37628a );
 a37630a <=( a37629a  and  a37624a );
 a37634a <=( (not A167)  and  A168 );
 a37635a <=( A169  and  a37634a );
 a37639a <=( A200  and  A199 );
 a37640a <=( A166  and  a37639a );
 a37641a <=( a37640a  and  a37635a );
 a37645a <=( A298  and  (not A266) );
 a37646a <=( (not A265)  and  a37645a );
 a37650a <=( (not A302)  and  A300 );
 a37651a <=( (not A299)  and  a37650a );
 a37652a <=( a37651a  and  a37646a );
 a37656a <=( (not A167)  and  A168 );
 a37657a <=( A169  and  a37656a );
 a37661a <=( A200  and  A199 );
 a37662a <=( A166  and  a37661a );
 a37663a <=( a37662a  and  a37657a );
 a37667a <=( (not A298)  and  (not A266) );
 a37668a <=( (not A265)  and  a37667a );
 a37672a <=( A301  and  A300 );
 a37673a <=( A299  and  a37672a );
 a37674a <=( a37673a  and  a37668a );
 a37678a <=( (not A167)  and  A168 );
 a37679a <=( A169  and  a37678a );
 a37683a <=( A200  and  A199 );
 a37684a <=( A166  and  a37683a );
 a37685a <=( a37684a  and  a37679a );
 a37689a <=( (not A298)  and  (not A266) );
 a37690a <=( (not A265)  and  a37689a );
 a37694a <=( (not A302)  and  A300 );
 a37695a <=( A299  and  a37694a );
 a37696a <=( a37695a  and  a37690a );
 a37700a <=( (not A167)  and  A168 );
 a37701a <=( A169  and  a37700a );
 a37705a <=( (not A200)  and  (not A199) );
 a37706a <=( A166  and  a37705a );
 a37707a <=( a37706a  and  a37701a );
 a37711a <=( A298  and  A268 );
 a37712a <=( (not A267)  and  a37711a );
 a37716a <=( A301  and  A300 );
 a37717a <=( (not A299)  and  a37716a );
 a37718a <=( a37717a  and  a37712a );
 a37722a <=( (not A167)  and  A168 );
 a37723a <=( A169  and  a37722a );
 a37727a <=( (not A200)  and  (not A199) );
 a37728a <=( A166  and  a37727a );
 a37729a <=( a37728a  and  a37723a );
 a37733a <=( A298  and  A268 );
 a37734a <=( (not A267)  and  a37733a );
 a37738a <=( (not A302)  and  A300 );
 a37739a <=( (not A299)  and  a37738a );
 a37740a <=( a37739a  and  a37734a );
 a37744a <=( (not A167)  and  A168 );
 a37745a <=( A169  and  a37744a );
 a37749a <=( (not A200)  and  (not A199) );
 a37750a <=( A166  and  a37749a );
 a37751a <=( a37750a  and  a37745a );
 a37755a <=( (not A298)  and  A268 );
 a37756a <=( (not A267)  and  a37755a );
 a37760a <=( A301  and  A300 );
 a37761a <=( A299  and  a37760a );
 a37762a <=( a37761a  and  a37756a );
 a37766a <=( (not A167)  and  A168 );
 a37767a <=( A169  and  a37766a );
 a37771a <=( (not A200)  and  (not A199) );
 a37772a <=( A166  and  a37771a );
 a37773a <=( a37772a  and  a37767a );
 a37777a <=( (not A298)  and  A268 );
 a37778a <=( (not A267)  and  a37777a );
 a37782a <=( (not A302)  and  A300 );
 a37783a <=( A299  and  a37782a );
 a37784a <=( a37783a  and  a37778a );
 a37788a <=( (not A167)  and  A168 );
 a37789a <=( A169  and  a37788a );
 a37793a <=( (not A200)  and  (not A199) );
 a37794a <=( A166  and  a37793a );
 a37795a <=( a37794a  and  a37789a );
 a37799a <=( A298  and  (not A269) );
 a37800a <=( (not A267)  and  a37799a );
 a37804a <=( A301  and  A300 );
 a37805a <=( (not A299)  and  a37804a );
 a37806a <=( a37805a  and  a37800a );
 a37810a <=( (not A167)  and  A168 );
 a37811a <=( A169  and  a37810a );
 a37815a <=( (not A200)  and  (not A199) );
 a37816a <=( A166  and  a37815a );
 a37817a <=( a37816a  and  a37811a );
 a37821a <=( A298  and  (not A269) );
 a37822a <=( (not A267)  and  a37821a );
 a37826a <=( (not A302)  and  A300 );
 a37827a <=( (not A299)  and  a37826a );
 a37828a <=( a37827a  and  a37822a );
 a37832a <=( (not A167)  and  A168 );
 a37833a <=( A169  and  a37832a );
 a37837a <=( (not A200)  and  (not A199) );
 a37838a <=( A166  and  a37837a );
 a37839a <=( a37838a  and  a37833a );
 a37843a <=( (not A298)  and  (not A269) );
 a37844a <=( (not A267)  and  a37843a );
 a37848a <=( A301  and  A300 );
 a37849a <=( A299  and  a37848a );
 a37850a <=( a37849a  and  a37844a );
 a37854a <=( (not A167)  and  A168 );
 a37855a <=( A169  and  a37854a );
 a37859a <=( (not A200)  and  (not A199) );
 a37860a <=( A166  and  a37859a );
 a37861a <=( a37860a  and  a37855a );
 a37865a <=( (not A298)  and  (not A269) );
 a37866a <=( (not A267)  and  a37865a );
 a37870a <=( (not A302)  and  A300 );
 a37871a <=( A299  and  a37870a );
 a37872a <=( a37871a  and  a37866a );
 a37876a <=( (not A167)  and  A168 );
 a37877a <=( A169  and  a37876a );
 a37881a <=( (not A200)  and  (not A199) );
 a37882a <=( A166  and  a37881a );
 a37883a <=( a37882a  and  a37877a );
 a37887a <=( A298  and  A266 );
 a37888a <=( A265  and  a37887a );
 a37892a <=( A301  and  A300 );
 a37893a <=( (not A299)  and  a37892a );
 a37894a <=( a37893a  and  a37888a );
 a37898a <=( (not A167)  and  A168 );
 a37899a <=( A169  and  a37898a );
 a37903a <=( (not A200)  and  (not A199) );
 a37904a <=( A166  and  a37903a );
 a37905a <=( a37904a  and  a37899a );
 a37909a <=( A298  and  A266 );
 a37910a <=( A265  and  a37909a );
 a37914a <=( (not A302)  and  A300 );
 a37915a <=( (not A299)  and  a37914a );
 a37916a <=( a37915a  and  a37910a );
 a37920a <=( (not A167)  and  A168 );
 a37921a <=( A169  and  a37920a );
 a37925a <=( (not A200)  and  (not A199) );
 a37926a <=( A166  and  a37925a );
 a37927a <=( a37926a  and  a37921a );
 a37931a <=( (not A298)  and  A266 );
 a37932a <=( A265  and  a37931a );
 a37936a <=( A301  and  A300 );
 a37937a <=( A299  and  a37936a );
 a37938a <=( a37937a  and  a37932a );
 a37942a <=( (not A167)  and  A168 );
 a37943a <=( A169  and  a37942a );
 a37947a <=( (not A200)  and  (not A199) );
 a37948a <=( A166  and  a37947a );
 a37949a <=( a37948a  and  a37943a );
 a37953a <=( (not A298)  and  A266 );
 a37954a <=( A265  and  a37953a );
 a37958a <=( (not A302)  and  A300 );
 a37959a <=( A299  and  a37958a );
 a37960a <=( a37959a  and  a37954a );
 a37964a <=( (not A167)  and  A168 );
 a37965a <=( A169  and  a37964a );
 a37969a <=( (not A200)  and  (not A199) );
 a37970a <=( A166  and  a37969a );
 a37971a <=( a37970a  and  a37965a );
 a37975a <=( A267  and  A266 );
 a37976a <=( (not A265)  and  a37975a );
 a37980a <=( A301  and  (not A300) );
 a37981a <=( A268  and  a37980a );
 a37982a <=( a37981a  and  a37976a );
 a37986a <=( (not A167)  and  A168 );
 a37987a <=( A169  and  a37986a );
 a37991a <=( (not A200)  and  (not A199) );
 a37992a <=( A166  and  a37991a );
 a37993a <=( a37992a  and  a37987a );
 a37997a <=( A267  and  A266 );
 a37998a <=( (not A265)  and  a37997a );
 a38002a <=( (not A302)  and  (not A300) );
 a38003a <=( A268  and  a38002a );
 a38004a <=( a38003a  and  a37998a );
 a38008a <=( (not A167)  and  A168 );
 a38009a <=( A169  and  a38008a );
 a38013a <=( (not A200)  and  (not A199) );
 a38014a <=( A166  and  a38013a );
 a38015a <=( a38014a  and  a38009a );
 a38019a <=( A267  and  A266 );
 a38020a <=( (not A265)  and  a38019a );
 a38024a <=( A299  and  A298 );
 a38025a <=( A268  and  a38024a );
 a38026a <=( a38025a  and  a38020a );
 a38030a <=( (not A167)  and  A168 );
 a38031a <=( A169  and  a38030a );
 a38035a <=( (not A200)  and  (not A199) );
 a38036a <=( A166  and  a38035a );
 a38037a <=( a38036a  and  a38031a );
 a38041a <=( A267  and  A266 );
 a38042a <=( (not A265)  and  a38041a );
 a38046a <=( (not A299)  and  (not A298) );
 a38047a <=( A268  and  a38046a );
 a38048a <=( a38047a  and  a38042a );
 a38052a <=( (not A167)  and  A168 );
 a38053a <=( A169  and  a38052a );
 a38057a <=( (not A200)  and  (not A199) );
 a38058a <=( A166  and  a38057a );
 a38059a <=( a38058a  and  a38053a );
 a38063a <=( A267  and  A266 );
 a38064a <=( (not A265)  and  a38063a );
 a38068a <=( A301  and  (not A300) );
 a38069a <=( (not A269)  and  a38068a );
 a38070a <=( a38069a  and  a38064a );
 a38074a <=( (not A167)  and  A168 );
 a38075a <=( A169  and  a38074a );
 a38079a <=( (not A200)  and  (not A199) );
 a38080a <=( A166  and  a38079a );
 a38081a <=( a38080a  and  a38075a );
 a38085a <=( A267  and  A266 );
 a38086a <=( (not A265)  and  a38085a );
 a38090a <=( (not A302)  and  (not A300) );
 a38091a <=( (not A269)  and  a38090a );
 a38092a <=( a38091a  and  a38086a );
 a38096a <=( (not A167)  and  A168 );
 a38097a <=( A169  and  a38096a );
 a38101a <=( (not A200)  and  (not A199) );
 a38102a <=( A166  and  a38101a );
 a38103a <=( a38102a  and  a38097a );
 a38107a <=( A267  and  A266 );
 a38108a <=( (not A265)  and  a38107a );
 a38112a <=( A299  and  A298 );
 a38113a <=( (not A269)  and  a38112a );
 a38114a <=( a38113a  and  a38108a );
 a38118a <=( (not A167)  and  A168 );
 a38119a <=( A169  and  a38118a );
 a38123a <=( (not A200)  and  (not A199) );
 a38124a <=( A166  and  a38123a );
 a38125a <=( a38124a  and  a38119a );
 a38129a <=( A267  and  A266 );
 a38130a <=( (not A265)  and  a38129a );
 a38134a <=( (not A299)  and  (not A298) );
 a38135a <=( (not A269)  and  a38134a );
 a38136a <=( a38135a  and  a38130a );
 a38140a <=( (not A167)  and  A168 );
 a38141a <=( A169  and  a38140a );
 a38145a <=( (not A200)  and  (not A199) );
 a38146a <=( A166  and  a38145a );
 a38147a <=( a38146a  and  a38141a );
 a38151a <=( A267  and  (not A266) );
 a38152a <=( A265  and  a38151a );
 a38156a <=( A301  and  (not A300) );
 a38157a <=( A268  and  a38156a );
 a38158a <=( a38157a  and  a38152a );
 a38162a <=( (not A167)  and  A168 );
 a38163a <=( A169  and  a38162a );
 a38167a <=( (not A200)  and  (not A199) );
 a38168a <=( A166  and  a38167a );
 a38169a <=( a38168a  and  a38163a );
 a38173a <=( A267  and  (not A266) );
 a38174a <=( A265  and  a38173a );
 a38178a <=( (not A302)  and  (not A300) );
 a38179a <=( A268  and  a38178a );
 a38180a <=( a38179a  and  a38174a );
 a38184a <=( (not A167)  and  A168 );
 a38185a <=( A169  and  a38184a );
 a38189a <=( (not A200)  and  (not A199) );
 a38190a <=( A166  and  a38189a );
 a38191a <=( a38190a  and  a38185a );
 a38195a <=( A267  and  (not A266) );
 a38196a <=( A265  and  a38195a );
 a38200a <=( A299  and  A298 );
 a38201a <=( A268  and  a38200a );
 a38202a <=( a38201a  and  a38196a );
 a38206a <=( (not A167)  and  A168 );
 a38207a <=( A169  and  a38206a );
 a38211a <=( (not A200)  and  (not A199) );
 a38212a <=( A166  and  a38211a );
 a38213a <=( a38212a  and  a38207a );
 a38217a <=( A267  and  (not A266) );
 a38218a <=( A265  and  a38217a );
 a38222a <=( (not A299)  and  (not A298) );
 a38223a <=( A268  and  a38222a );
 a38224a <=( a38223a  and  a38218a );
 a38228a <=( (not A167)  and  A168 );
 a38229a <=( A169  and  a38228a );
 a38233a <=( (not A200)  and  (not A199) );
 a38234a <=( A166  and  a38233a );
 a38235a <=( a38234a  and  a38229a );
 a38239a <=( A267  and  (not A266) );
 a38240a <=( A265  and  a38239a );
 a38244a <=( A301  and  (not A300) );
 a38245a <=( (not A269)  and  a38244a );
 a38246a <=( a38245a  and  a38240a );
 a38250a <=( (not A167)  and  A168 );
 a38251a <=( A169  and  a38250a );
 a38255a <=( (not A200)  and  (not A199) );
 a38256a <=( A166  and  a38255a );
 a38257a <=( a38256a  and  a38251a );
 a38261a <=( A267  and  (not A266) );
 a38262a <=( A265  and  a38261a );
 a38266a <=( (not A302)  and  (not A300) );
 a38267a <=( (not A269)  and  a38266a );
 a38268a <=( a38267a  and  a38262a );
 a38272a <=( (not A167)  and  A168 );
 a38273a <=( A169  and  a38272a );
 a38277a <=( (not A200)  and  (not A199) );
 a38278a <=( A166  and  a38277a );
 a38279a <=( a38278a  and  a38273a );
 a38283a <=( A267  and  (not A266) );
 a38284a <=( A265  and  a38283a );
 a38288a <=( A299  and  A298 );
 a38289a <=( (not A269)  and  a38288a );
 a38290a <=( a38289a  and  a38284a );
 a38294a <=( (not A167)  and  A168 );
 a38295a <=( A169  and  a38294a );
 a38299a <=( (not A200)  and  (not A199) );
 a38300a <=( A166  and  a38299a );
 a38301a <=( a38300a  and  a38295a );
 a38305a <=( A267  and  (not A266) );
 a38306a <=( A265  and  a38305a );
 a38310a <=( (not A299)  and  (not A298) );
 a38311a <=( (not A269)  and  a38310a );
 a38312a <=( a38311a  and  a38306a );
 a38316a <=( (not A167)  and  A168 );
 a38317a <=( A169  and  a38316a );
 a38321a <=( (not A200)  and  (not A199) );
 a38322a <=( A166  and  a38321a );
 a38323a <=( a38322a  and  a38317a );
 a38327a <=( A298  and  (not A266) );
 a38328a <=( (not A265)  and  a38327a );
 a38332a <=( A301  and  A300 );
 a38333a <=( (not A299)  and  a38332a );
 a38334a <=( a38333a  and  a38328a );
 a38338a <=( (not A167)  and  A168 );
 a38339a <=( A169  and  a38338a );
 a38343a <=( (not A200)  and  (not A199) );
 a38344a <=( A166  and  a38343a );
 a38345a <=( a38344a  and  a38339a );
 a38349a <=( A298  and  (not A266) );
 a38350a <=( (not A265)  and  a38349a );
 a38354a <=( (not A302)  and  A300 );
 a38355a <=( (not A299)  and  a38354a );
 a38356a <=( a38355a  and  a38350a );
 a38360a <=( (not A167)  and  A168 );
 a38361a <=( A169  and  a38360a );
 a38365a <=( (not A200)  and  (not A199) );
 a38366a <=( A166  and  a38365a );
 a38367a <=( a38366a  and  a38361a );
 a38371a <=( (not A298)  and  (not A266) );
 a38372a <=( (not A265)  and  a38371a );
 a38376a <=( A301  and  A300 );
 a38377a <=( A299  and  a38376a );
 a38378a <=( a38377a  and  a38372a );
 a38382a <=( (not A167)  and  A168 );
 a38383a <=( A169  and  a38382a );
 a38387a <=( (not A200)  and  (not A199) );
 a38388a <=( A166  and  a38387a );
 a38389a <=( a38388a  and  a38383a );
 a38393a <=( (not A298)  and  (not A266) );
 a38394a <=( (not A265)  and  a38393a );
 a38398a <=( (not A302)  and  A300 );
 a38399a <=( A299  and  a38398a );
 a38400a <=( a38399a  and  a38394a );
 a38404a <=( (not A232)  and  (not A168) );
 a38405a <=( A169  and  a38404a );
 a38409a <=( (not A235)  and  (not A234) );
 a38410a <=( A233  and  a38409a );
 a38411a <=( a38410a  and  a38405a );
 a38415a <=( A266  and  (not A265) );
 a38416a <=( A236  and  a38415a );
 a38420a <=( A269  and  (not A268) );
 a38421a <=( (not A267)  and  a38420a );
 a38422a <=( a38421a  and  a38416a );
 a38426a <=( (not A232)  and  (not A168) );
 a38427a <=( A169  and  a38426a );
 a38431a <=( (not A235)  and  (not A234) );
 a38432a <=( A233  and  a38431a );
 a38433a <=( a38432a  and  a38427a );
 a38437a <=( (not A266)  and  A265 );
 a38438a <=( A236  and  a38437a );
 a38442a <=( A269  and  (not A268) );
 a38443a <=( (not A267)  and  a38442a );
 a38444a <=( a38443a  and  a38438a );
 a38448a <=( A232  and  (not A168) );
 a38449a <=( A169  and  a38448a );
 a38453a <=( (not A235)  and  (not A234) );
 a38454a <=( (not A233)  and  a38453a );
 a38455a <=( a38454a  and  a38449a );
 a38459a <=( A266  and  (not A265) );
 a38460a <=( A236  and  a38459a );
 a38464a <=( A269  and  (not A268) );
 a38465a <=( (not A267)  and  a38464a );
 a38466a <=( a38465a  and  a38460a );
 a38470a <=( A232  and  (not A168) );
 a38471a <=( A169  and  a38470a );
 a38475a <=( (not A235)  and  (not A234) );
 a38476a <=( (not A233)  and  a38475a );
 a38477a <=( a38476a  and  a38471a );
 a38481a <=( (not A266)  and  A265 );
 a38482a <=( A236  and  a38481a );
 a38486a <=( A269  and  (not A268) );
 a38487a <=( (not A267)  and  a38486a );
 a38488a <=( a38487a  and  a38482a );
 a38492a <=( (not A199)  and  (not A168) );
 a38493a <=( A169  and  a38492a );
 a38497a <=( A202  and  A201 );
 a38498a <=( A200  and  a38497a );
 a38499a <=( a38498a  and  a38493a );
 a38503a <=( A269  and  (not A268) );
 a38504a <=( A267  and  a38503a );
 a38508a <=( A302  and  (not A301) );
 a38509a <=( A300  and  a38508a );
 a38510a <=( a38509a  and  a38504a );
 a38514a <=( (not A199)  and  (not A168) );
 a38515a <=( A169  and  a38514a );
 a38519a <=( (not A203)  and  A201 );
 a38520a <=( A200  and  a38519a );
 a38521a <=( a38520a  and  a38515a );
 a38525a <=( A269  and  (not A268) );
 a38526a <=( A267  and  a38525a );
 a38530a <=( A302  and  (not A301) );
 a38531a <=( A300  and  a38530a );
 a38532a <=( a38531a  and  a38526a );
 a38536a <=( (not A199)  and  (not A168) );
 a38537a <=( A169  and  a38536a );
 a38541a <=( (not A202)  and  (not A201) );
 a38542a <=( A200  and  a38541a );
 a38543a <=( a38542a  and  a38537a );
 a38547a <=( (not A268)  and  A267 );
 a38548a <=( A203  and  a38547a );
 a38552a <=( A301  and  (not A300) );
 a38553a <=( A269  and  a38552a );
 a38554a <=( a38553a  and  a38548a );
 a38558a <=( (not A199)  and  (not A168) );
 a38559a <=( A169  and  a38558a );
 a38563a <=( (not A202)  and  (not A201) );
 a38564a <=( A200  and  a38563a );
 a38565a <=( a38564a  and  a38559a );
 a38569a <=( (not A268)  and  A267 );
 a38570a <=( A203  and  a38569a );
 a38574a <=( (not A302)  and  (not A300) );
 a38575a <=( A269  and  a38574a );
 a38576a <=( a38575a  and  a38570a );
 a38580a <=( (not A199)  and  (not A168) );
 a38581a <=( A169  and  a38580a );
 a38585a <=( (not A202)  and  (not A201) );
 a38586a <=( A200  and  a38585a );
 a38587a <=( a38586a  and  a38581a );
 a38591a <=( (not A268)  and  A267 );
 a38592a <=( A203  and  a38591a );
 a38596a <=( A299  and  A298 );
 a38597a <=( A269  and  a38596a );
 a38598a <=( a38597a  and  a38592a );
 a38602a <=( (not A199)  and  (not A168) );
 a38603a <=( A169  and  a38602a );
 a38607a <=( (not A202)  and  (not A201) );
 a38608a <=( A200  and  a38607a );
 a38609a <=( a38608a  and  a38603a );
 a38613a <=( (not A268)  and  A267 );
 a38614a <=( A203  and  a38613a );
 a38618a <=( (not A299)  and  (not A298) );
 a38619a <=( A269  and  a38618a );
 a38620a <=( a38619a  and  a38614a );
 a38624a <=( (not A199)  and  (not A168) );
 a38625a <=( A169  and  a38624a );
 a38629a <=( (not A202)  and  (not A201) );
 a38630a <=( A200  and  a38629a );
 a38631a <=( a38630a  and  a38625a );
 a38635a <=( A268  and  (not A267) );
 a38636a <=( A203  and  a38635a );
 a38640a <=( A302  and  (not A301) );
 a38641a <=( A300  and  a38640a );
 a38642a <=( a38641a  and  a38636a );
 a38646a <=( (not A199)  and  (not A168) );
 a38647a <=( A169  and  a38646a );
 a38651a <=( (not A202)  and  (not A201) );
 a38652a <=( A200  and  a38651a );
 a38653a <=( a38652a  and  a38647a );
 a38657a <=( (not A269)  and  (not A267) );
 a38658a <=( A203  and  a38657a );
 a38662a <=( A302  and  (not A301) );
 a38663a <=( A300  and  a38662a );
 a38664a <=( a38663a  and  a38658a );
 a38668a <=( (not A199)  and  (not A168) );
 a38669a <=( A169  and  a38668a );
 a38673a <=( (not A202)  and  (not A201) );
 a38674a <=( A200  and  a38673a );
 a38675a <=( a38674a  and  a38669a );
 a38679a <=( A266  and  A265 );
 a38680a <=( A203  and  a38679a );
 a38684a <=( A302  and  (not A301) );
 a38685a <=( A300  and  a38684a );
 a38686a <=( a38685a  and  a38680a );
 a38690a <=( (not A199)  and  (not A168) );
 a38691a <=( A169  and  a38690a );
 a38695a <=( (not A202)  and  (not A201) );
 a38696a <=( A200  and  a38695a );
 a38697a <=( a38696a  and  a38691a );
 a38701a <=( (not A266)  and  (not A265) );
 a38702a <=( A203  and  a38701a );
 a38706a <=( A302  and  (not A301) );
 a38707a <=( A300  and  a38706a );
 a38708a <=( a38707a  and  a38702a );
 a38712a <=( A199  and  (not A168) );
 a38713a <=( A169  and  a38712a );
 a38717a <=( A202  and  A201 );
 a38718a <=( (not A200)  and  a38717a );
 a38719a <=( a38718a  and  a38713a );
 a38723a <=( A269  and  (not A268) );
 a38724a <=( A267  and  a38723a );
 a38728a <=( A302  and  (not A301) );
 a38729a <=( A300  and  a38728a );
 a38730a <=( a38729a  and  a38724a );
 a38734a <=( A199  and  (not A168) );
 a38735a <=( A169  and  a38734a );
 a38739a <=( (not A203)  and  A201 );
 a38740a <=( (not A200)  and  a38739a );
 a38741a <=( a38740a  and  a38735a );
 a38745a <=( A269  and  (not A268) );
 a38746a <=( A267  and  a38745a );
 a38750a <=( A302  and  (not A301) );
 a38751a <=( A300  and  a38750a );
 a38752a <=( a38751a  and  a38746a );
 a38756a <=( A199  and  (not A168) );
 a38757a <=( A169  and  a38756a );
 a38761a <=( (not A202)  and  (not A201) );
 a38762a <=( (not A200)  and  a38761a );
 a38763a <=( a38762a  and  a38757a );
 a38767a <=( (not A268)  and  A267 );
 a38768a <=( A203  and  a38767a );
 a38772a <=( A301  and  (not A300) );
 a38773a <=( A269  and  a38772a );
 a38774a <=( a38773a  and  a38768a );
 a38778a <=( A199  and  (not A168) );
 a38779a <=( A169  and  a38778a );
 a38783a <=( (not A202)  and  (not A201) );
 a38784a <=( (not A200)  and  a38783a );
 a38785a <=( a38784a  and  a38779a );
 a38789a <=( (not A268)  and  A267 );
 a38790a <=( A203  and  a38789a );
 a38794a <=( (not A302)  and  (not A300) );
 a38795a <=( A269  and  a38794a );
 a38796a <=( a38795a  and  a38790a );
 a38800a <=( A199  and  (not A168) );
 a38801a <=( A169  and  a38800a );
 a38805a <=( (not A202)  and  (not A201) );
 a38806a <=( (not A200)  and  a38805a );
 a38807a <=( a38806a  and  a38801a );
 a38811a <=( (not A268)  and  A267 );
 a38812a <=( A203  and  a38811a );
 a38816a <=( A299  and  A298 );
 a38817a <=( A269  and  a38816a );
 a38818a <=( a38817a  and  a38812a );
 a38822a <=( A199  and  (not A168) );
 a38823a <=( A169  and  a38822a );
 a38827a <=( (not A202)  and  (not A201) );
 a38828a <=( (not A200)  and  a38827a );
 a38829a <=( a38828a  and  a38823a );
 a38833a <=( (not A268)  and  A267 );
 a38834a <=( A203  and  a38833a );
 a38838a <=( (not A299)  and  (not A298) );
 a38839a <=( A269  and  a38838a );
 a38840a <=( a38839a  and  a38834a );
 a38844a <=( A199  and  (not A168) );
 a38845a <=( A169  and  a38844a );
 a38849a <=( (not A202)  and  (not A201) );
 a38850a <=( (not A200)  and  a38849a );
 a38851a <=( a38850a  and  a38845a );
 a38855a <=( A268  and  (not A267) );
 a38856a <=( A203  and  a38855a );
 a38860a <=( A302  and  (not A301) );
 a38861a <=( A300  and  a38860a );
 a38862a <=( a38861a  and  a38856a );
 a38866a <=( A199  and  (not A168) );
 a38867a <=( A169  and  a38866a );
 a38871a <=( (not A202)  and  (not A201) );
 a38872a <=( (not A200)  and  a38871a );
 a38873a <=( a38872a  and  a38867a );
 a38877a <=( (not A269)  and  (not A267) );
 a38878a <=( A203  and  a38877a );
 a38882a <=( A302  and  (not A301) );
 a38883a <=( A300  and  a38882a );
 a38884a <=( a38883a  and  a38878a );
 a38888a <=( A199  and  (not A168) );
 a38889a <=( A169  and  a38888a );
 a38893a <=( (not A202)  and  (not A201) );
 a38894a <=( (not A200)  and  a38893a );
 a38895a <=( a38894a  and  a38889a );
 a38899a <=( A266  and  A265 );
 a38900a <=( A203  and  a38899a );
 a38904a <=( A302  and  (not A301) );
 a38905a <=( A300  and  a38904a );
 a38906a <=( a38905a  and  a38900a );
 a38910a <=( A199  and  (not A168) );
 a38911a <=( A169  and  a38910a );
 a38915a <=( (not A202)  and  (not A201) );
 a38916a <=( (not A200)  and  a38915a );
 a38917a <=( a38916a  and  a38911a );
 a38921a <=( (not A266)  and  (not A265) );
 a38922a <=( A203  and  a38921a );
 a38926a <=( A302  and  (not A301) );
 a38927a <=( A300  and  a38926a );
 a38928a <=( a38927a  and  a38922a );
 a38932a <=( A168  and  (not A169) );
 a38933a <=( (not A170)  and  a38932a );
 a38937a <=( A201  and  A200 );
 a38938a <=( (not A199)  and  a38937a );
 a38939a <=( a38938a  and  a38933a );
 a38943a <=( (not A268)  and  A267 );
 a38944a <=( A202  and  a38943a );
 a38948a <=( A301  and  (not A300) );
 a38949a <=( A269  and  a38948a );
 a38950a <=( a38949a  and  a38944a );
 a38954a <=( A168  and  (not A169) );
 a38955a <=( (not A170)  and  a38954a );
 a38959a <=( A201  and  A200 );
 a38960a <=( (not A199)  and  a38959a );
 a38961a <=( a38960a  and  a38955a );
 a38965a <=( (not A268)  and  A267 );
 a38966a <=( A202  and  a38965a );
 a38970a <=( (not A302)  and  (not A300) );
 a38971a <=( A269  and  a38970a );
 a38972a <=( a38971a  and  a38966a );
 a38976a <=( A168  and  (not A169) );
 a38977a <=( (not A170)  and  a38976a );
 a38981a <=( A201  and  A200 );
 a38982a <=( (not A199)  and  a38981a );
 a38983a <=( a38982a  and  a38977a );
 a38987a <=( (not A268)  and  A267 );
 a38988a <=( A202  and  a38987a );
 a38992a <=( A299  and  A298 );
 a38993a <=( A269  and  a38992a );
 a38994a <=( a38993a  and  a38988a );
 a38998a <=( A168  and  (not A169) );
 a38999a <=( (not A170)  and  a38998a );
 a39003a <=( A201  and  A200 );
 a39004a <=( (not A199)  and  a39003a );
 a39005a <=( a39004a  and  a38999a );
 a39009a <=( (not A268)  and  A267 );
 a39010a <=( A202  and  a39009a );
 a39014a <=( (not A299)  and  (not A298) );
 a39015a <=( A269  and  a39014a );
 a39016a <=( a39015a  and  a39010a );
 a39020a <=( A168  and  (not A169) );
 a39021a <=( (not A170)  and  a39020a );
 a39025a <=( A201  and  A200 );
 a39026a <=( (not A199)  and  a39025a );
 a39027a <=( a39026a  and  a39021a );
 a39031a <=( A268  and  (not A267) );
 a39032a <=( A202  and  a39031a );
 a39036a <=( A302  and  (not A301) );
 a39037a <=( A300  and  a39036a );
 a39038a <=( a39037a  and  a39032a );
 a39042a <=( A168  and  (not A169) );
 a39043a <=( (not A170)  and  a39042a );
 a39047a <=( A201  and  A200 );
 a39048a <=( (not A199)  and  a39047a );
 a39049a <=( a39048a  and  a39043a );
 a39053a <=( (not A269)  and  (not A267) );
 a39054a <=( A202  and  a39053a );
 a39058a <=( A302  and  (not A301) );
 a39059a <=( A300  and  a39058a );
 a39060a <=( a39059a  and  a39054a );
 a39064a <=( A168  and  (not A169) );
 a39065a <=( (not A170)  and  a39064a );
 a39069a <=( A201  and  A200 );
 a39070a <=( (not A199)  and  a39069a );
 a39071a <=( a39070a  and  a39065a );
 a39075a <=( A266  and  A265 );
 a39076a <=( A202  and  a39075a );
 a39080a <=( A302  and  (not A301) );
 a39081a <=( A300  and  a39080a );
 a39082a <=( a39081a  and  a39076a );
 a39086a <=( A168  and  (not A169) );
 a39087a <=( (not A170)  and  a39086a );
 a39091a <=( A201  and  A200 );
 a39092a <=( (not A199)  and  a39091a );
 a39093a <=( a39092a  and  a39087a );
 a39097a <=( (not A266)  and  (not A265) );
 a39098a <=( A202  and  a39097a );
 a39102a <=( A302  and  (not A301) );
 a39103a <=( A300  and  a39102a );
 a39104a <=( a39103a  and  a39098a );
 a39108a <=( A168  and  (not A169) );
 a39109a <=( (not A170)  and  a39108a );
 a39113a <=( A201  and  A200 );
 a39114a <=( (not A199)  and  a39113a );
 a39115a <=( a39114a  and  a39109a );
 a39119a <=( (not A268)  and  A267 );
 a39120a <=( (not A203)  and  a39119a );
 a39124a <=( A301  and  (not A300) );
 a39125a <=( A269  and  a39124a );
 a39126a <=( a39125a  and  a39120a );
 a39130a <=( A168  and  (not A169) );
 a39131a <=( (not A170)  and  a39130a );
 a39135a <=( A201  and  A200 );
 a39136a <=( (not A199)  and  a39135a );
 a39137a <=( a39136a  and  a39131a );
 a39141a <=( (not A268)  and  A267 );
 a39142a <=( (not A203)  and  a39141a );
 a39146a <=( (not A302)  and  (not A300) );
 a39147a <=( A269  and  a39146a );
 a39148a <=( a39147a  and  a39142a );
 a39152a <=( A168  and  (not A169) );
 a39153a <=( (not A170)  and  a39152a );
 a39157a <=( A201  and  A200 );
 a39158a <=( (not A199)  and  a39157a );
 a39159a <=( a39158a  and  a39153a );
 a39163a <=( (not A268)  and  A267 );
 a39164a <=( (not A203)  and  a39163a );
 a39168a <=( A299  and  A298 );
 a39169a <=( A269  and  a39168a );
 a39170a <=( a39169a  and  a39164a );
 a39174a <=( A168  and  (not A169) );
 a39175a <=( (not A170)  and  a39174a );
 a39179a <=( A201  and  A200 );
 a39180a <=( (not A199)  and  a39179a );
 a39181a <=( a39180a  and  a39175a );
 a39185a <=( (not A268)  and  A267 );
 a39186a <=( (not A203)  and  a39185a );
 a39190a <=( (not A299)  and  (not A298) );
 a39191a <=( A269  and  a39190a );
 a39192a <=( a39191a  and  a39186a );
 a39196a <=( A168  and  (not A169) );
 a39197a <=( (not A170)  and  a39196a );
 a39201a <=( A201  and  A200 );
 a39202a <=( (not A199)  and  a39201a );
 a39203a <=( a39202a  and  a39197a );
 a39207a <=( A268  and  (not A267) );
 a39208a <=( (not A203)  and  a39207a );
 a39212a <=( A302  and  (not A301) );
 a39213a <=( A300  and  a39212a );
 a39214a <=( a39213a  and  a39208a );
 a39218a <=( A168  and  (not A169) );
 a39219a <=( (not A170)  and  a39218a );
 a39223a <=( A201  and  A200 );
 a39224a <=( (not A199)  and  a39223a );
 a39225a <=( a39224a  and  a39219a );
 a39229a <=( (not A269)  and  (not A267) );
 a39230a <=( (not A203)  and  a39229a );
 a39234a <=( A302  and  (not A301) );
 a39235a <=( A300  and  a39234a );
 a39236a <=( a39235a  and  a39230a );
 a39240a <=( A168  and  (not A169) );
 a39241a <=( (not A170)  and  a39240a );
 a39245a <=( A201  and  A200 );
 a39246a <=( (not A199)  and  a39245a );
 a39247a <=( a39246a  and  a39241a );
 a39251a <=( A266  and  A265 );
 a39252a <=( (not A203)  and  a39251a );
 a39256a <=( A302  and  (not A301) );
 a39257a <=( A300  and  a39256a );
 a39258a <=( a39257a  and  a39252a );
 a39262a <=( A168  and  (not A169) );
 a39263a <=( (not A170)  and  a39262a );
 a39267a <=( A201  and  A200 );
 a39268a <=( (not A199)  and  a39267a );
 a39269a <=( a39268a  and  a39263a );
 a39273a <=( (not A266)  and  (not A265) );
 a39274a <=( (not A203)  and  a39273a );
 a39278a <=( A302  and  (not A301) );
 a39279a <=( A300  and  a39278a );
 a39280a <=( a39279a  and  a39274a );
 a39284a <=( A168  and  (not A169) );
 a39285a <=( (not A170)  and  a39284a );
 a39289a <=( (not A201)  and  A200 );
 a39290a <=( (not A199)  and  a39289a );
 a39291a <=( a39290a  and  a39285a );
 a39295a <=( (not A267)  and  A203 );
 a39296a <=( (not A202)  and  a39295a );
 a39300a <=( A301  and  (not A300) );
 a39301a <=( A268  and  a39300a );
 a39302a <=( a39301a  and  a39296a );
 a39306a <=( A168  and  (not A169) );
 a39307a <=( (not A170)  and  a39306a );
 a39311a <=( (not A201)  and  A200 );
 a39312a <=( (not A199)  and  a39311a );
 a39313a <=( a39312a  and  a39307a );
 a39317a <=( (not A267)  and  A203 );
 a39318a <=( (not A202)  and  a39317a );
 a39322a <=( (not A302)  and  (not A300) );
 a39323a <=( A268  and  a39322a );
 a39324a <=( a39323a  and  a39318a );
 a39328a <=( A168  and  (not A169) );
 a39329a <=( (not A170)  and  a39328a );
 a39333a <=( (not A201)  and  A200 );
 a39334a <=( (not A199)  and  a39333a );
 a39335a <=( a39334a  and  a39329a );
 a39339a <=( (not A267)  and  A203 );
 a39340a <=( (not A202)  and  a39339a );
 a39344a <=( A299  and  A298 );
 a39345a <=( A268  and  a39344a );
 a39346a <=( a39345a  and  a39340a );
 a39350a <=( A168  and  (not A169) );
 a39351a <=( (not A170)  and  a39350a );
 a39355a <=( (not A201)  and  A200 );
 a39356a <=( (not A199)  and  a39355a );
 a39357a <=( a39356a  and  a39351a );
 a39361a <=( (not A267)  and  A203 );
 a39362a <=( (not A202)  and  a39361a );
 a39366a <=( (not A299)  and  (not A298) );
 a39367a <=( A268  and  a39366a );
 a39368a <=( a39367a  and  a39362a );
 a39372a <=( A168  and  (not A169) );
 a39373a <=( (not A170)  and  a39372a );
 a39377a <=( (not A201)  and  A200 );
 a39378a <=( (not A199)  and  a39377a );
 a39379a <=( a39378a  and  a39373a );
 a39383a <=( (not A267)  and  A203 );
 a39384a <=( (not A202)  and  a39383a );
 a39388a <=( A301  and  (not A300) );
 a39389a <=( (not A269)  and  a39388a );
 a39390a <=( a39389a  and  a39384a );
 a39394a <=( A168  and  (not A169) );
 a39395a <=( (not A170)  and  a39394a );
 a39399a <=( (not A201)  and  A200 );
 a39400a <=( (not A199)  and  a39399a );
 a39401a <=( a39400a  and  a39395a );
 a39405a <=( (not A267)  and  A203 );
 a39406a <=( (not A202)  and  a39405a );
 a39410a <=( (not A302)  and  (not A300) );
 a39411a <=( (not A269)  and  a39410a );
 a39412a <=( a39411a  and  a39406a );
 a39416a <=( A168  and  (not A169) );
 a39417a <=( (not A170)  and  a39416a );
 a39421a <=( (not A201)  and  A200 );
 a39422a <=( (not A199)  and  a39421a );
 a39423a <=( a39422a  and  a39417a );
 a39427a <=( (not A267)  and  A203 );
 a39428a <=( (not A202)  and  a39427a );
 a39432a <=( A299  and  A298 );
 a39433a <=( (not A269)  and  a39432a );
 a39434a <=( a39433a  and  a39428a );
 a39438a <=( A168  and  (not A169) );
 a39439a <=( (not A170)  and  a39438a );
 a39443a <=( (not A201)  and  A200 );
 a39444a <=( (not A199)  and  a39443a );
 a39445a <=( a39444a  and  a39439a );
 a39449a <=( (not A267)  and  A203 );
 a39450a <=( (not A202)  and  a39449a );
 a39454a <=( (not A299)  and  (not A298) );
 a39455a <=( (not A269)  and  a39454a );
 a39456a <=( a39455a  and  a39450a );
 a39460a <=( A168  and  (not A169) );
 a39461a <=( (not A170)  and  a39460a );
 a39465a <=( (not A201)  and  A200 );
 a39466a <=( (not A199)  and  a39465a );
 a39467a <=( a39466a  and  a39461a );
 a39471a <=( A265  and  A203 );
 a39472a <=( (not A202)  and  a39471a );
 a39476a <=( A301  and  (not A300) );
 a39477a <=( A266  and  a39476a );
 a39478a <=( a39477a  and  a39472a );
 a39482a <=( A168  and  (not A169) );
 a39483a <=( (not A170)  and  a39482a );
 a39487a <=( (not A201)  and  A200 );
 a39488a <=( (not A199)  and  a39487a );
 a39489a <=( a39488a  and  a39483a );
 a39493a <=( A265  and  A203 );
 a39494a <=( (not A202)  and  a39493a );
 a39498a <=( (not A302)  and  (not A300) );
 a39499a <=( A266  and  a39498a );
 a39500a <=( a39499a  and  a39494a );
 a39504a <=( A168  and  (not A169) );
 a39505a <=( (not A170)  and  a39504a );
 a39509a <=( (not A201)  and  A200 );
 a39510a <=( (not A199)  and  a39509a );
 a39511a <=( a39510a  and  a39505a );
 a39515a <=( A265  and  A203 );
 a39516a <=( (not A202)  and  a39515a );
 a39520a <=( A299  and  A298 );
 a39521a <=( A266  and  a39520a );
 a39522a <=( a39521a  and  a39516a );
 a39526a <=( A168  and  (not A169) );
 a39527a <=( (not A170)  and  a39526a );
 a39531a <=( (not A201)  and  A200 );
 a39532a <=( (not A199)  and  a39531a );
 a39533a <=( a39532a  and  a39527a );
 a39537a <=( A265  and  A203 );
 a39538a <=( (not A202)  and  a39537a );
 a39542a <=( (not A299)  and  (not A298) );
 a39543a <=( A266  and  a39542a );
 a39544a <=( a39543a  and  a39538a );
 a39548a <=( A168  and  (not A169) );
 a39549a <=( (not A170)  and  a39548a );
 a39553a <=( (not A201)  and  A200 );
 a39554a <=( (not A199)  and  a39553a );
 a39555a <=( a39554a  and  a39549a );
 a39559a <=( (not A265)  and  A203 );
 a39560a <=( (not A202)  and  a39559a );
 a39564a <=( A301  and  (not A300) );
 a39565a <=( (not A266)  and  a39564a );
 a39566a <=( a39565a  and  a39560a );
 a39570a <=( A168  and  (not A169) );
 a39571a <=( (not A170)  and  a39570a );
 a39575a <=( (not A201)  and  A200 );
 a39576a <=( (not A199)  and  a39575a );
 a39577a <=( a39576a  and  a39571a );
 a39581a <=( (not A265)  and  A203 );
 a39582a <=( (not A202)  and  a39581a );
 a39586a <=( (not A302)  and  (not A300) );
 a39587a <=( (not A266)  and  a39586a );
 a39588a <=( a39587a  and  a39582a );
 a39592a <=( A168  and  (not A169) );
 a39593a <=( (not A170)  and  a39592a );
 a39597a <=( (not A201)  and  A200 );
 a39598a <=( (not A199)  and  a39597a );
 a39599a <=( a39598a  and  a39593a );
 a39603a <=( (not A265)  and  A203 );
 a39604a <=( (not A202)  and  a39603a );
 a39608a <=( A299  and  A298 );
 a39609a <=( (not A266)  and  a39608a );
 a39610a <=( a39609a  and  a39604a );
 a39614a <=( A168  and  (not A169) );
 a39615a <=( (not A170)  and  a39614a );
 a39619a <=( (not A201)  and  A200 );
 a39620a <=( (not A199)  and  a39619a );
 a39621a <=( a39620a  and  a39615a );
 a39625a <=( (not A265)  and  A203 );
 a39626a <=( (not A202)  and  a39625a );
 a39630a <=( (not A299)  and  (not A298) );
 a39631a <=( (not A266)  and  a39630a );
 a39632a <=( a39631a  and  a39626a );
 a39636a <=( A168  and  (not A169) );
 a39637a <=( (not A170)  and  a39636a );
 a39641a <=( A201  and  (not A200) );
 a39642a <=( A199  and  a39641a );
 a39643a <=( a39642a  and  a39637a );
 a39647a <=( (not A268)  and  A267 );
 a39648a <=( A202  and  a39647a );
 a39652a <=( A301  and  (not A300) );
 a39653a <=( A269  and  a39652a );
 a39654a <=( a39653a  and  a39648a );
 a39658a <=( A168  and  (not A169) );
 a39659a <=( (not A170)  and  a39658a );
 a39663a <=( A201  and  (not A200) );
 a39664a <=( A199  and  a39663a );
 a39665a <=( a39664a  and  a39659a );
 a39669a <=( (not A268)  and  A267 );
 a39670a <=( A202  and  a39669a );
 a39674a <=( (not A302)  and  (not A300) );
 a39675a <=( A269  and  a39674a );
 a39676a <=( a39675a  and  a39670a );
 a39680a <=( A168  and  (not A169) );
 a39681a <=( (not A170)  and  a39680a );
 a39685a <=( A201  and  (not A200) );
 a39686a <=( A199  and  a39685a );
 a39687a <=( a39686a  and  a39681a );
 a39691a <=( (not A268)  and  A267 );
 a39692a <=( A202  and  a39691a );
 a39696a <=( A299  and  A298 );
 a39697a <=( A269  and  a39696a );
 a39698a <=( a39697a  and  a39692a );
 a39702a <=( A168  and  (not A169) );
 a39703a <=( (not A170)  and  a39702a );
 a39707a <=( A201  and  (not A200) );
 a39708a <=( A199  and  a39707a );
 a39709a <=( a39708a  and  a39703a );
 a39713a <=( (not A268)  and  A267 );
 a39714a <=( A202  and  a39713a );
 a39718a <=( (not A299)  and  (not A298) );
 a39719a <=( A269  and  a39718a );
 a39720a <=( a39719a  and  a39714a );
 a39724a <=( A168  and  (not A169) );
 a39725a <=( (not A170)  and  a39724a );
 a39729a <=( A201  and  (not A200) );
 a39730a <=( A199  and  a39729a );
 a39731a <=( a39730a  and  a39725a );
 a39735a <=( A268  and  (not A267) );
 a39736a <=( A202  and  a39735a );
 a39740a <=( A302  and  (not A301) );
 a39741a <=( A300  and  a39740a );
 a39742a <=( a39741a  and  a39736a );
 a39746a <=( A168  and  (not A169) );
 a39747a <=( (not A170)  and  a39746a );
 a39751a <=( A201  and  (not A200) );
 a39752a <=( A199  and  a39751a );
 a39753a <=( a39752a  and  a39747a );
 a39757a <=( (not A269)  and  (not A267) );
 a39758a <=( A202  and  a39757a );
 a39762a <=( A302  and  (not A301) );
 a39763a <=( A300  and  a39762a );
 a39764a <=( a39763a  and  a39758a );
 a39768a <=( A168  and  (not A169) );
 a39769a <=( (not A170)  and  a39768a );
 a39773a <=( A201  and  (not A200) );
 a39774a <=( A199  and  a39773a );
 a39775a <=( a39774a  and  a39769a );
 a39779a <=( A266  and  A265 );
 a39780a <=( A202  and  a39779a );
 a39784a <=( A302  and  (not A301) );
 a39785a <=( A300  and  a39784a );
 a39786a <=( a39785a  and  a39780a );
 a39790a <=( A168  and  (not A169) );
 a39791a <=( (not A170)  and  a39790a );
 a39795a <=( A201  and  (not A200) );
 a39796a <=( A199  and  a39795a );
 a39797a <=( a39796a  and  a39791a );
 a39801a <=( (not A266)  and  (not A265) );
 a39802a <=( A202  and  a39801a );
 a39806a <=( A302  and  (not A301) );
 a39807a <=( A300  and  a39806a );
 a39808a <=( a39807a  and  a39802a );
 a39812a <=( A168  and  (not A169) );
 a39813a <=( (not A170)  and  a39812a );
 a39817a <=( A201  and  (not A200) );
 a39818a <=( A199  and  a39817a );
 a39819a <=( a39818a  and  a39813a );
 a39823a <=( (not A268)  and  A267 );
 a39824a <=( (not A203)  and  a39823a );
 a39828a <=( A301  and  (not A300) );
 a39829a <=( A269  and  a39828a );
 a39830a <=( a39829a  and  a39824a );
 a39834a <=( A168  and  (not A169) );
 a39835a <=( (not A170)  and  a39834a );
 a39839a <=( A201  and  (not A200) );
 a39840a <=( A199  and  a39839a );
 a39841a <=( a39840a  and  a39835a );
 a39845a <=( (not A268)  and  A267 );
 a39846a <=( (not A203)  and  a39845a );
 a39850a <=( (not A302)  and  (not A300) );
 a39851a <=( A269  and  a39850a );
 a39852a <=( a39851a  and  a39846a );
 a39856a <=( A168  and  (not A169) );
 a39857a <=( (not A170)  and  a39856a );
 a39861a <=( A201  and  (not A200) );
 a39862a <=( A199  and  a39861a );
 a39863a <=( a39862a  and  a39857a );
 a39867a <=( (not A268)  and  A267 );
 a39868a <=( (not A203)  and  a39867a );
 a39872a <=( A299  and  A298 );
 a39873a <=( A269  and  a39872a );
 a39874a <=( a39873a  and  a39868a );
 a39878a <=( A168  and  (not A169) );
 a39879a <=( (not A170)  and  a39878a );
 a39883a <=( A201  and  (not A200) );
 a39884a <=( A199  and  a39883a );
 a39885a <=( a39884a  and  a39879a );
 a39889a <=( (not A268)  and  A267 );
 a39890a <=( (not A203)  and  a39889a );
 a39894a <=( (not A299)  and  (not A298) );
 a39895a <=( A269  and  a39894a );
 a39896a <=( a39895a  and  a39890a );
 a39900a <=( A168  and  (not A169) );
 a39901a <=( (not A170)  and  a39900a );
 a39905a <=( A201  and  (not A200) );
 a39906a <=( A199  and  a39905a );
 a39907a <=( a39906a  and  a39901a );
 a39911a <=( A268  and  (not A267) );
 a39912a <=( (not A203)  and  a39911a );
 a39916a <=( A302  and  (not A301) );
 a39917a <=( A300  and  a39916a );
 a39918a <=( a39917a  and  a39912a );
 a39922a <=( A168  and  (not A169) );
 a39923a <=( (not A170)  and  a39922a );
 a39927a <=( A201  and  (not A200) );
 a39928a <=( A199  and  a39927a );
 a39929a <=( a39928a  and  a39923a );
 a39933a <=( (not A269)  and  (not A267) );
 a39934a <=( (not A203)  and  a39933a );
 a39938a <=( A302  and  (not A301) );
 a39939a <=( A300  and  a39938a );
 a39940a <=( a39939a  and  a39934a );
 a39944a <=( A168  and  (not A169) );
 a39945a <=( (not A170)  and  a39944a );
 a39949a <=( A201  and  (not A200) );
 a39950a <=( A199  and  a39949a );
 a39951a <=( a39950a  and  a39945a );
 a39955a <=( A266  and  A265 );
 a39956a <=( (not A203)  and  a39955a );
 a39960a <=( A302  and  (not A301) );
 a39961a <=( A300  and  a39960a );
 a39962a <=( a39961a  and  a39956a );
 a39966a <=( A168  and  (not A169) );
 a39967a <=( (not A170)  and  a39966a );
 a39971a <=( A201  and  (not A200) );
 a39972a <=( A199  and  a39971a );
 a39973a <=( a39972a  and  a39967a );
 a39977a <=( (not A266)  and  (not A265) );
 a39978a <=( (not A203)  and  a39977a );
 a39982a <=( A302  and  (not A301) );
 a39983a <=( A300  and  a39982a );
 a39984a <=( a39983a  and  a39978a );
 a39988a <=( A168  and  (not A169) );
 a39989a <=( (not A170)  and  a39988a );
 a39993a <=( (not A201)  and  (not A200) );
 a39994a <=( A199  and  a39993a );
 a39995a <=( a39994a  and  a39989a );
 a39999a <=( (not A267)  and  A203 );
 a40000a <=( (not A202)  and  a39999a );
 a40004a <=( A301  and  (not A300) );
 a40005a <=( A268  and  a40004a );
 a40006a <=( a40005a  and  a40000a );
 a40010a <=( A168  and  (not A169) );
 a40011a <=( (not A170)  and  a40010a );
 a40015a <=( (not A201)  and  (not A200) );
 a40016a <=( A199  and  a40015a );
 a40017a <=( a40016a  and  a40011a );
 a40021a <=( (not A267)  and  A203 );
 a40022a <=( (not A202)  and  a40021a );
 a40026a <=( (not A302)  and  (not A300) );
 a40027a <=( A268  and  a40026a );
 a40028a <=( a40027a  and  a40022a );
 a40032a <=( A168  and  (not A169) );
 a40033a <=( (not A170)  and  a40032a );
 a40037a <=( (not A201)  and  (not A200) );
 a40038a <=( A199  and  a40037a );
 a40039a <=( a40038a  and  a40033a );
 a40043a <=( (not A267)  and  A203 );
 a40044a <=( (not A202)  and  a40043a );
 a40048a <=( A299  and  A298 );
 a40049a <=( A268  and  a40048a );
 a40050a <=( a40049a  and  a40044a );
 a40054a <=( A168  and  (not A169) );
 a40055a <=( (not A170)  and  a40054a );
 a40059a <=( (not A201)  and  (not A200) );
 a40060a <=( A199  and  a40059a );
 a40061a <=( a40060a  and  a40055a );
 a40065a <=( (not A267)  and  A203 );
 a40066a <=( (not A202)  and  a40065a );
 a40070a <=( (not A299)  and  (not A298) );
 a40071a <=( A268  and  a40070a );
 a40072a <=( a40071a  and  a40066a );
 a40076a <=( A168  and  (not A169) );
 a40077a <=( (not A170)  and  a40076a );
 a40081a <=( (not A201)  and  (not A200) );
 a40082a <=( A199  and  a40081a );
 a40083a <=( a40082a  and  a40077a );
 a40087a <=( (not A267)  and  A203 );
 a40088a <=( (not A202)  and  a40087a );
 a40092a <=( A301  and  (not A300) );
 a40093a <=( (not A269)  and  a40092a );
 a40094a <=( a40093a  and  a40088a );
 a40098a <=( A168  and  (not A169) );
 a40099a <=( (not A170)  and  a40098a );
 a40103a <=( (not A201)  and  (not A200) );
 a40104a <=( A199  and  a40103a );
 a40105a <=( a40104a  and  a40099a );
 a40109a <=( (not A267)  and  A203 );
 a40110a <=( (not A202)  and  a40109a );
 a40114a <=( (not A302)  and  (not A300) );
 a40115a <=( (not A269)  and  a40114a );
 a40116a <=( a40115a  and  a40110a );
 a40120a <=( A168  and  (not A169) );
 a40121a <=( (not A170)  and  a40120a );
 a40125a <=( (not A201)  and  (not A200) );
 a40126a <=( A199  and  a40125a );
 a40127a <=( a40126a  and  a40121a );
 a40131a <=( (not A267)  and  A203 );
 a40132a <=( (not A202)  and  a40131a );
 a40136a <=( A299  and  A298 );
 a40137a <=( (not A269)  and  a40136a );
 a40138a <=( a40137a  and  a40132a );
 a40142a <=( A168  and  (not A169) );
 a40143a <=( (not A170)  and  a40142a );
 a40147a <=( (not A201)  and  (not A200) );
 a40148a <=( A199  and  a40147a );
 a40149a <=( a40148a  and  a40143a );
 a40153a <=( (not A267)  and  A203 );
 a40154a <=( (not A202)  and  a40153a );
 a40158a <=( (not A299)  and  (not A298) );
 a40159a <=( (not A269)  and  a40158a );
 a40160a <=( a40159a  and  a40154a );
 a40164a <=( A168  and  (not A169) );
 a40165a <=( (not A170)  and  a40164a );
 a40169a <=( (not A201)  and  (not A200) );
 a40170a <=( A199  and  a40169a );
 a40171a <=( a40170a  and  a40165a );
 a40175a <=( A265  and  A203 );
 a40176a <=( (not A202)  and  a40175a );
 a40180a <=( A301  and  (not A300) );
 a40181a <=( A266  and  a40180a );
 a40182a <=( a40181a  and  a40176a );
 a40186a <=( A168  and  (not A169) );
 a40187a <=( (not A170)  and  a40186a );
 a40191a <=( (not A201)  and  (not A200) );
 a40192a <=( A199  and  a40191a );
 a40193a <=( a40192a  and  a40187a );
 a40197a <=( A265  and  A203 );
 a40198a <=( (not A202)  and  a40197a );
 a40202a <=( (not A302)  and  (not A300) );
 a40203a <=( A266  and  a40202a );
 a40204a <=( a40203a  and  a40198a );
 a40208a <=( A168  and  (not A169) );
 a40209a <=( (not A170)  and  a40208a );
 a40213a <=( (not A201)  and  (not A200) );
 a40214a <=( A199  and  a40213a );
 a40215a <=( a40214a  and  a40209a );
 a40219a <=( A265  and  A203 );
 a40220a <=( (not A202)  and  a40219a );
 a40224a <=( A299  and  A298 );
 a40225a <=( A266  and  a40224a );
 a40226a <=( a40225a  and  a40220a );
 a40230a <=( A168  and  (not A169) );
 a40231a <=( (not A170)  and  a40230a );
 a40235a <=( (not A201)  and  (not A200) );
 a40236a <=( A199  and  a40235a );
 a40237a <=( a40236a  and  a40231a );
 a40241a <=( A265  and  A203 );
 a40242a <=( (not A202)  and  a40241a );
 a40246a <=( (not A299)  and  (not A298) );
 a40247a <=( A266  and  a40246a );
 a40248a <=( a40247a  and  a40242a );
 a40252a <=( A168  and  (not A169) );
 a40253a <=( (not A170)  and  a40252a );
 a40257a <=( (not A201)  and  (not A200) );
 a40258a <=( A199  and  a40257a );
 a40259a <=( a40258a  and  a40253a );
 a40263a <=( (not A265)  and  A203 );
 a40264a <=( (not A202)  and  a40263a );
 a40268a <=( A301  and  (not A300) );
 a40269a <=( (not A266)  and  a40268a );
 a40270a <=( a40269a  and  a40264a );
 a40274a <=( A168  and  (not A169) );
 a40275a <=( (not A170)  and  a40274a );
 a40279a <=( (not A201)  and  (not A200) );
 a40280a <=( A199  and  a40279a );
 a40281a <=( a40280a  and  a40275a );
 a40285a <=( (not A265)  and  A203 );
 a40286a <=( (not A202)  and  a40285a );
 a40290a <=( (not A302)  and  (not A300) );
 a40291a <=( (not A266)  and  a40290a );
 a40292a <=( a40291a  and  a40286a );
 a40296a <=( A168  and  (not A169) );
 a40297a <=( (not A170)  and  a40296a );
 a40301a <=( (not A201)  and  (not A200) );
 a40302a <=( A199  and  a40301a );
 a40303a <=( a40302a  and  a40297a );
 a40307a <=( (not A265)  and  A203 );
 a40308a <=( (not A202)  and  a40307a );
 a40312a <=( A299  and  A298 );
 a40313a <=( (not A266)  and  a40312a );
 a40314a <=( a40313a  and  a40308a );
 a40318a <=( A168  and  (not A169) );
 a40319a <=( (not A170)  and  a40318a );
 a40323a <=( (not A201)  and  (not A200) );
 a40324a <=( A199  and  a40323a );
 a40325a <=( a40324a  and  a40319a );
 a40329a <=( (not A265)  and  A203 );
 a40330a <=( (not A202)  and  a40329a );
 a40334a <=( (not A299)  and  (not A298) );
 a40335a <=( (not A266)  and  a40334a );
 a40336a <=( a40335a  and  a40330a );
 a40340a <=( A202  and  A200 );
 a40341a <=( (not A199)  and  a40340a );
 a40345a <=( (not A234)  and  A233 );
 a40346a <=( (not A232)  and  a40345a );
 a40347a <=( a40346a  and  a40341a );
 a40351a <=( (not A265)  and  A236 );
 a40352a <=( (not A235)  and  a40351a );
 a40355a <=( (not A267)  and  A266 );
 a40358a <=( A269  and  (not A268) );
 a40359a <=( a40358a  and  a40355a );
 a40360a <=( a40359a  and  a40352a );
 a40364a <=( A202  and  A200 );
 a40365a <=( (not A199)  and  a40364a );
 a40369a <=( (not A234)  and  A233 );
 a40370a <=( (not A232)  and  a40369a );
 a40371a <=( a40370a  and  a40365a );
 a40375a <=( A265  and  A236 );
 a40376a <=( (not A235)  and  a40375a );
 a40379a <=( (not A267)  and  (not A266) );
 a40382a <=( A269  and  (not A268) );
 a40383a <=( a40382a  and  a40379a );
 a40384a <=( a40383a  and  a40376a );
 a40388a <=( A202  and  A200 );
 a40389a <=( (not A199)  and  a40388a );
 a40393a <=( (not A234)  and  (not A233) );
 a40394a <=( A232  and  a40393a );
 a40395a <=( a40394a  and  a40389a );
 a40399a <=( (not A265)  and  A236 );
 a40400a <=( (not A235)  and  a40399a );
 a40403a <=( (not A267)  and  A266 );
 a40406a <=( A269  and  (not A268) );
 a40407a <=( a40406a  and  a40403a );
 a40408a <=( a40407a  and  a40400a );
 a40412a <=( A202  and  A200 );
 a40413a <=( (not A199)  and  a40412a );
 a40417a <=( (not A234)  and  (not A233) );
 a40418a <=( A232  and  a40417a );
 a40419a <=( a40418a  and  a40413a );
 a40423a <=( A265  and  A236 );
 a40424a <=( (not A235)  and  a40423a );
 a40427a <=( (not A267)  and  (not A266) );
 a40430a <=( A269  and  (not A268) );
 a40431a <=( a40430a  and  a40427a );
 a40432a <=( a40431a  and  a40424a );
 a40436a <=( (not A203)  and  A200 );
 a40437a <=( (not A199)  and  a40436a );
 a40441a <=( (not A234)  and  A233 );
 a40442a <=( (not A232)  and  a40441a );
 a40443a <=( a40442a  and  a40437a );
 a40447a <=( (not A265)  and  A236 );
 a40448a <=( (not A235)  and  a40447a );
 a40451a <=( (not A267)  and  A266 );
 a40454a <=( A269  and  (not A268) );
 a40455a <=( a40454a  and  a40451a );
 a40456a <=( a40455a  and  a40448a );
 a40460a <=( (not A203)  and  A200 );
 a40461a <=( (not A199)  and  a40460a );
 a40465a <=( (not A234)  and  A233 );
 a40466a <=( (not A232)  and  a40465a );
 a40467a <=( a40466a  and  a40461a );
 a40471a <=( A265  and  A236 );
 a40472a <=( (not A235)  and  a40471a );
 a40475a <=( (not A267)  and  (not A266) );
 a40478a <=( A269  and  (not A268) );
 a40479a <=( a40478a  and  a40475a );
 a40480a <=( a40479a  and  a40472a );
 a40484a <=( (not A203)  and  A200 );
 a40485a <=( (not A199)  and  a40484a );
 a40489a <=( (not A234)  and  (not A233) );
 a40490a <=( A232  and  a40489a );
 a40491a <=( a40490a  and  a40485a );
 a40495a <=( (not A265)  and  A236 );
 a40496a <=( (not A235)  and  a40495a );
 a40499a <=( (not A267)  and  A266 );
 a40502a <=( A269  and  (not A268) );
 a40503a <=( a40502a  and  a40499a );
 a40504a <=( a40503a  and  a40496a );
 a40508a <=( (not A203)  and  A200 );
 a40509a <=( (not A199)  and  a40508a );
 a40513a <=( (not A234)  and  (not A233) );
 a40514a <=( A232  and  a40513a );
 a40515a <=( a40514a  and  a40509a );
 a40519a <=( A265  and  A236 );
 a40520a <=( (not A235)  and  a40519a );
 a40523a <=( (not A267)  and  (not A266) );
 a40526a <=( A269  and  (not A268) );
 a40527a <=( a40526a  and  a40523a );
 a40528a <=( a40527a  and  a40520a );
 a40532a <=( A202  and  (not A200) );
 a40533a <=( A199  and  a40532a );
 a40537a <=( (not A234)  and  A233 );
 a40538a <=( (not A232)  and  a40537a );
 a40539a <=( a40538a  and  a40533a );
 a40543a <=( (not A265)  and  A236 );
 a40544a <=( (not A235)  and  a40543a );
 a40547a <=( (not A267)  and  A266 );
 a40550a <=( A269  and  (not A268) );
 a40551a <=( a40550a  and  a40547a );
 a40552a <=( a40551a  and  a40544a );
 a40556a <=( A202  and  (not A200) );
 a40557a <=( A199  and  a40556a );
 a40561a <=( (not A234)  and  A233 );
 a40562a <=( (not A232)  and  a40561a );
 a40563a <=( a40562a  and  a40557a );
 a40567a <=( A265  and  A236 );
 a40568a <=( (not A235)  and  a40567a );
 a40571a <=( (not A267)  and  (not A266) );
 a40574a <=( A269  and  (not A268) );
 a40575a <=( a40574a  and  a40571a );
 a40576a <=( a40575a  and  a40568a );
 a40580a <=( A202  and  (not A200) );
 a40581a <=( A199  and  a40580a );
 a40585a <=( (not A234)  and  (not A233) );
 a40586a <=( A232  and  a40585a );
 a40587a <=( a40586a  and  a40581a );
 a40591a <=( (not A265)  and  A236 );
 a40592a <=( (not A235)  and  a40591a );
 a40595a <=( (not A267)  and  A266 );
 a40598a <=( A269  and  (not A268) );
 a40599a <=( a40598a  and  a40595a );
 a40600a <=( a40599a  and  a40592a );
 a40604a <=( A202  and  (not A200) );
 a40605a <=( A199  and  a40604a );
 a40609a <=( (not A234)  and  (not A233) );
 a40610a <=( A232  and  a40609a );
 a40611a <=( a40610a  and  a40605a );
 a40615a <=( A265  and  A236 );
 a40616a <=( (not A235)  and  a40615a );
 a40619a <=( (not A267)  and  (not A266) );
 a40622a <=( A269  and  (not A268) );
 a40623a <=( a40622a  and  a40619a );
 a40624a <=( a40623a  and  a40616a );
 a40628a <=( (not A203)  and  (not A200) );
 a40629a <=( A199  and  a40628a );
 a40633a <=( (not A234)  and  A233 );
 a40634a <=( (not A232)  and  a40633a );
 a40635a <=( a40634a  and  a40629a );
 a40639a <=( (not A265)  and  A236 );
 a40640a <=( (not A235)  and  a40639a );
 a40643a <=( (not A267)  and  A266 );
 a40646a <=( A269  and  (not A268) );
 a40647a <=( a40646a  and  a40643a );
 a40648a <=( a40647a  and  a40640a );
 a40652a <=( (not A203)  and  (not A200) );
 a40653a <=( A199  and  a40652a );
 a40657a <=( (not A234)  and  A233 );
 a40658a <=( (not A232)  and  a40657a );
 a40659a <=( a40658a  and  a40653a );
 a40663a <=( A265  and  A236 );
 a40664a <=( (not A235)  and  a40663a );
 a40667a <=( (not A267)  and  (not A266) );
 a40670a <=( A269  and  (not A268) );
 a40671a <=( a40670a  and  a40667a );
 a40672a <=( a40671a  and  a40664a );
 a40676a <=( (not A203)  and  (not A200) );
 a40677a <=( A199  and  a40676a );
 a40681a <=( (not A234)  and  (not A233) );
 a40682a <=( A232  and  a40681a );
 a40683a <=( a40682a  and  a40677a );
 a40687a <=( (not A265)  and  A236 );
 a40688a <=( (not A235)  and  a40687a );
 a40691a <=( (not A267)  and  A266 );
 a40694a <=( A269  and  (not A268) );
 a40695a <=( a40694a  and  a40691a );
 a40696a <=( a40695a  and  a40688a );
 a40700a <=( (not A203)  and  (not A200) );
 a40701a <=( A199  and  a40700a );
 a40705a <=( (not A234)  and  (not A233) );
 a40706a <=( A232  and  a40705a );
 a40707a <=( a40706a  and  a40701a );
 a40711a <=( A265  and  A236 );
 a40712a <=( (not A235)  and  a40711a );
 a40715a <=( (not A267)  and  (not A266) );
 a40718a <=( A269  and  (not A268) );
 a40719a <=( a40718a  and  a40715a );
 a40720a <=( a40719a  and  a40712a );
 a40724a <=( (not A199)  and  A166 );
 a40725a <=( A167  and  a40724a );
 a40729a <=( (not A202)  and  (not A201) );
 a40730a <=( A200  and  a40729a );
 a40731a <=( a40730a  and  a40725a );
 a40735a <=( (not A268)  and  A267 );
 a40736a <=( A203  and  a40735a );
 a40739a <=( A300  and  A269 );
 a40742a <=( A302  and  (not A301) );
 a40743a <=( a40742a  and  a40739a );
 a40744a <=( a40743a  and  a40736a );
 a40748a <=( A199  and  A166 );
 a40749a <=( A167  and  a40748a );
 a40753a <=( (not A202)  and  (not A201) );
 a40754a <=( (not A200)  and  a40753a );
 a40755a <=( a40754a  and  a40749a );
 a40759a <=( (not A268)  and  A267 );
 a40760a <=( A203  and  a40759a );
 a40763a <=( A300  and  A269 );
 a40766a <=( A302  and  (not A301) );
 a40767a <=( a40766a  and  a40763a );
 a40768a <=( a40767a  and  a40760a );
 a40772a <=( (not A199)  and  (not A166) );
 a40773a <=( (not A167)  and  a40772a );
 a40777a <=( (not A202)  and  (not A201) );
 a40778a <=( A200  and  a40777a );
 a40779a <=( a40778a  and  a40773a );
 a40783a <=( (not A268)  and  A267 );
 a40784a <=( A203  and  a40783a );
 a40787a <=( A300  and  A269 );
 a40790a <=( A302  and  (not A301) );
 a40791a <=( a40790a  and  a40787a );
 a40792a <=( a40791a  and  a40784a );
 a40796a <=( A199  and  (not A166) );
 a40797a <=( (not A167)  and  a40796a );
 a40801a <=( (not A202)  and  (not A201) );
 a40802a <=( (not A200)  and  a40801a );
 a40803a <=( a40802a  and  a40797a );
 a40807a <=( (not A268)  and  A267 );
 a40808a <=( A203  and  a40807a );
 a40811a <=( A300  and  A269 );
 a40814a <=( A302  and  (not A301) );
 a40815a <=( a40814a  and  a40811a );
 a40816a <=( a40815a  and  a40808a );
 a40820a <=( A200  and  (not A199) );
 a40821a <=( A170  and  a40820a );
 a40825a <=( (not A234)  and  A233 );
 a40826a <=( (not A232)  and  a40825a );
 a40827a <=( a40826a  and  a40821a );
 a40831a <=( (not A265)  and  A236 );
 a40832a <=( (not A235)  and  a40831a );
 a40835a <=( (not A267)  and  A266 );
 a40838a <=( A269  and  (not A268) );
 a40839a <=( a40838a  and  a40835a );
 a40840a <=( a40839a  and  a40832a );
 a40844a <=( A200  and  (not A199) );
 a40845a <=( A170  and  a40844a );
 a40849a <=( (not A234)  and  A233 );
 a40850a <=( (not A232)  and  a40849a );
 a40851a <=( a40850a  and  a40845a );
 a40855a <=( A265  and  A236 );
 a40856a <=( (not A235)  and  a40855a );
 a40859a <=( (not A267)  and  (not A266) );
 a40862a <=( A269  and  (not A268) );
 a40863a <=( a40862a  and  a40859a );
 a40864a <=( a40863a  and  a40856a );
 a40868a <=( A200  and  (not A199) );
 a40869a <=( A170  and  a40868a );
 a40873a <=( (not A234)  and  (not A233) );
 a40874a <=( A232  and  a40873a );
 a40875a <=( a40874a  and  a40869a );
 a40879a <=( (not A265)  and  A236 );
 a40880a <=( (not A235)  and  a40879a );
 a40883a <=( (not A267)  and  A266 );
 a40886a <=( A269  and  (not A268) );
 a40887a <=( a40886a  and  a40883a );
 a40888a <=( a40887a  and  a40880a );
 a40892a <=( A200  and  (not A199) );
 a40893a <=( A170  and  a40892a );
 a40897a <=( (not A234)  and  (not A233) );
 a40898a <=( A232  and  a40897a );
 a40899a <=( a40898a  and  a40893a );
 a40903a <=( A265  and  A236 );
 a40904a <=( (not A235)  and  a40903a );
 a40907a <=( (not A267)  and  (not A266) );
 a40910a <=( A269  and  (not A268) );
 a40911a <=( a40910a  and  a40907a );
 a40912a <=( a40911a  and  a40904a );
 a40916a <=( (not A200)  and  A199 );
 a40917a <=( A170  and  a40916a );
 a40921a <=( (not A234)  and  A233 );
 a40922a <=( (not A232)  and  a40921a );
 a40923a <=( a40922a  and  a40917a );
 a40927a <=( (not A265)  and  A236 );
 a40928a <=( (not A235)  and  a40927a );
 a40931a <=( (not A267)  and  A266 );
 a40934a <=( A269  and  (not A268) );
 a40935a <=( a40934a  and  a40931a );
 a40936a <=( a40935a  and  a40928a );
 a40940a <=( (not A200)  and  A199 );
 a40941a <=( A170  and  a40940a );
 a40945a <=( (not A234)  and  A233 );
 a40946a <=( (not A232)  and  a40945a );
 a40947a <=( a40946a  and  a40941a );
 a40951a <=( A265  and  A236 );
 a40952a <=( (not A235)  and  a40951a );
 a40955a <=( (not A267)  and  (not A266) );
 a40958a <=( A269  and  (not A268) );
 a40959a <=( a40958a  and  a40955a );
 a40960a <=( a40959a  and  a40952a );
 a40964a <=( (not A200)  and  A199 );
 a40965a <=( A170  and  a40964a );
 a40969a <=( (not A234)  and  (not A233) );
 a40970a <=( A232  and  a40969a );
 a40971a <=( a40970a  and  a40965a );
 a40975a <=( (not A265)  and  A236 );
 a40976a <=( (not A235)  and  a40975a );
 a40979a <=( (not A267)  and  A266 );
 a40982a <=( A269  and  (not A268) );
 a40983a <=( a40982a  and  a40979a );
 a40984a <=( a40983a  and  a40976a );
 a40988a <=( (not A200)  and  A199 );
 a40989a <=( A170  and  a40988a );
 a40993a <=( (not A234)  and  (not A233) );
 a40994a <=( A232  and  a40993a );
 a40995a <=( a40994a  and  a40989a );
 a40999a <=( A265  and  A236 );
 a41000a <=( (not A235)  and  a40999a );
 a41003a <=( (not A267)  and  (not A266) );
 a41006a <=( A269  and  (not A268) );
 a41007a <=( a41006a  and  a41003a );
 a41008a <=( a41007a  and  a41000a );
 a41012a <=( A167  and  A168 );
 a41013a <=( A170  and  a41012a );
 a41017a <=( (not A202)  and  A201 );
 a41018a <=( (not A166)  and  a41017a );
 a41019a <=( a41018a  and  a41013a );
 a41023a <=( A268  and  (not A267) );
 a41024a <=( A203  and  a41023a );
 a41027a <=( (not A299)  and  A298 );
 a41030a <=( A301  and  A300 );
 a41031a <=( a41030a  and  a41027a );
 a41032a <=( a41031a  and  a41024a );
 a41036a <=( A167  and  A168 );
 a41037a <=( A170  and  a41036a );
 a41041a <=( (not A202)  and  A201 );
 a41042a <=( (not A166)  and  a41041a );
 a41043a <=( a41042a  and  a41037a );
 a41047a <=( A268  and  (not A267) );
 a41048a <=( A203  and  a41047a );
 a41051a <=( (not A299)  and  A298 );
 a41054a <=( (not A302)  and  A300 );
 a41055a <=( a41054a  and  a41051a );
 a41056a <=( a41055a  and  a41048a );
 a41060a <=( A167  and  A168 );
 a41061a <=( A170  and  a41060a );
 a41065a <=( (not A202)  and  A201 );
 a41066a <=( (not A166)  and  a41065a );
 a41067a <=( a41066a  and  a41061a );
 a41071a <=( A268  and  (not A267) );
 a41072a <=( A203  and  a41071a );
 a41075a <=( A299  and  (not A298) );
 a41078a <=( A301  and  A300 );
 a41079a <=( a41078a  and  a41075a );
 a41080a <=( a41079a  and  a41072a );
 a41084a <=( A167  and  A168 );
 a41085a <=( A170  and  a41084a );
 a41089a <=( (not A202)  and  A201 );
 a41090a <=( (not A166)  and  a41089a );
 a41091a <=( a41090a  and  a41085a );
 a41095a <=( A268  and  (not A267) );
 a41096a <=( A203  and  a41095a );
 a41099a <=( A299  and  (not A298) );
 a41102a <=( (not A302)  and  A300 );
 a41103a <=( a41102a  and  a41099a );
 a41104a <=( a41103a  and  a41096a );
 a41108a <=( A167  and  A168 );
 a41109a <=( A170  and  a41108a );
 a41113a <=( (not A202)  and  A201 );
 a41114a <=( (not A166)  and  a41113a );
 a41115a <=( a41114a  and  a41109a );
 a41119a <=( (not A269)  and  (not A267) );
 a41120a <=( A203  and  a41119a );
 a41123a <=( (not A299)  and  A298 );
 a41126a <=( A301  and  A300 );
 a41127a <=( a41126a  and  a41123a );
 a41128a <=( a41127a  and  a41120a );
 a41132a <=( A167  and  A168 );
 a41133a <=( A170  and  a41132a );
 a41137a <=( (not A202)  and  A201 );
 a41138a <=( (not A166)  and  a41137a );
 a41139a <=( a41138a  and  a41133a );
 a41143a <=( (not A269)  and  (not A267) );
 a41144a <=( A203  and  a41143a );
 a41147a <=( (not A299)  and  A298 );
 a41150a <=( (not A302)  and  A300 );
 a41151a <=( a41150a  and  a41147a );
 a41152a <=( a41151a  and  a41144a );
 a41156a <=( A167  and  A168 );
 a41157a <=( A170  and  a41156a );
 a41161a <=( (not A202)  and  A201 );
 a41162a <=( (not A166)  and  a41161a );
 a41163a <=( a41162a  and  a41157a );
 a41167a <=( (not A269)  and  (not A267) );
 a41168a <=( A203  and  a41167a );
 a41171a <=( A299  and  (not A298) );
 a41174a <=( A301  and  A300 );
 a41175a <=( a41174a  and  a41171a );
 a41176a <=( a41175a  and  a41168a );
 a41180a <=( A167  and  A168 );
 a41181a <=( A170  and  a41180a );
 a41185a <=( (not A202)  and  A201 );
 a41186a <=( (not A166)  and  a41185a );
 a41187a <=( a41186a  and  a41181a );
 a41191a <=( (not A269)  and  (not A267) );
 a41192a <=( A203  and  a41191a );
 a41195a <=( A299  and  (not A298) );
 a41198a <=( (not A302)  and  A300 );
 a41199a <=( a41198a  and  a41195a );
 a41200a <=( a41199a  and  a41192a );
 a41204a <=( A167  and  A168 );
 a41205a <=( A170  and  a41204a );
 a41209a <=( (not A202)  and  A201 );
 a41210a <=( (not A166)  and  a41209a );
 a41211a <=( a41210a  and  a41205a );
 a41215a <=( A266  and  A265 );
 a41216a <=( A203  and  a41215a );
 a41219a <=( (not A299)  and  A298 );
 a41222a <=( A301  and  A300 );
 a41223a <=( a41222a  and  a41219a );
 a41224a <=( a41223a  and  a41216a );
 a41228a <=( A167  and  A168 );
 a41229a <=( A170  and  a41228a );
 a41233a <=( (not A202)  and  A201 );
 a41234a <=( (not A166)  and  a41233a );
 a41235a <=( a41234a  and  a41229a );
 a41239a <=( A266  and  A265 );
 a41240a <=( A203  and  a41239a );
 a41243a <=( (not A299)  and  A298 );
 a41246a <=( (not A302)  and  A300 );
 a41247a <=( a41246a  and  a41243a );
 a41248a <=( a41247a  and  a41240a );
 a41252a <=( A167  and  A168 );
 a41253a <=( A170  and  a41252a );
 a41257a <=( (not A202)  and  A201 );
 a41258a <=( (not A166)  and  a41257a );
 a41259a <=( a41258a  and  a41253a );
 a41263a <=( A266  and  A265 );
 a41264a <=( A203  and  a41263a );
 a41267a <=( A299  and  (not A298) );
 a41270a <=( A301  and  A300 );
 a41271a <=( a41270a  and  a41267a );
 a41272a <=( a41271a  and  a41264a );
 a41276a <=( A167  and  A168 );
 a41277a <=( A170  and  a41276a );
 a41281a <=( (not A202)  and  A201 );
 a41282a <=( (not A166)  and  a41281a );
 a41283a <=( a41282a  and  a41277a );
 a41287a <=( A266  and  A265 );
 a41288a <=( A203  and  a41287a );
 a41291a <=( A299  and  (not A298) );
 a41294a <=( (not A302)  and  A300 );
 a41295a <=( a41294a  and  a41291a );
 a41296a <=( a41295a  and  a41288a );
 a41300a <=( A167  and  A168 );
 a41301a <=( A170  and  a41300a );
 a41305a <=( (not A202)  and  A201 );
 a41306a <=( (not A166)  and  a41305a );
 a41307a <=( a41306a  and  a41301a );
 a41311a <=( A266  and  (not A265) );
 a41312a <=( A203  and  a41311a );
 a41315a <=( A268  and  A267 );
 a41318a <=( A301  and  (not A300) );
 a41319a <=( a41318a  and  a41315a );
 a41320a <=( a41319a  and  a41312a );
 a41324a <=( A167  and  A168 );
 a41325a <=( A170  and  a41324a );
 a41329a <=( (not A202)  and  A201 );
 a41330a <=( (not A166)  and  a41329a );
 a41331a <=( a41330a  and  a41325a );
 a41335a <=( A266  and  (not A265) );
 a41336a <=( A203  and  a41335a );
 a41339a <=( A268  and  A267 );
 a41342a <=( (not A302)  and  (not A300) );
 a41343a <=( a41342a  and  a41339a );
 a41344a <=( a41343a  and  a41336a );
 a41348a <=( A167  and  A168 );
 a41349a <=( A170  and  a41348a );
 a41353a <=( (not A202)  and  A201 );
 a41354a <=( (not A166)  and  a41353a );
 a41355a <=( a41354a  and  a41349a );
 a41359a <=( A266  and  (not A265) );
 a41360a <=( A203  and  a41359a );
 a41363a <=( A268  and  A267 );
 a41366a <=( A299  and  A298 );
 a41367a <=( a41366a  and  a41363a );
 a41368a <=( a41367a  and  a41360a );
 a41372a <=( A167  and  A168 );
 a41373a <=( A170  and  a41372a );
 a41377a <=( (not A202)  and  A201 );
 a41378a <=( (not A166)  and  a41377a );
 a41379a <=( a41378a  and  a41373a );
 a41383a <=( A266  and  (not A265) );
 a41384a <=( A203  and  a41383a );
 a41387a <=( A268  and  A267 );
 a41390a <=( (not A299)  and  (not A298) );
 a41391a <=( a41390a  and  a41387a );
 a41392a <=( a41391a  and  a41384a );
 a41396a <=( A167  and  A168 );
 a41397a <=( A170  and  a41396a );
 a41401a <=( (not A202)  and  A201 );
 a41402a <=( (not A166)  and  a41401a );
 a41403a <=( a41402a  and  a41397a );
 a41407a <=( A266  and  (not A265) );
 a41408a <=( A203  and  a41407a );
 a41411a <=( (not A269)  and  A267 );
 a41414a <=( A301  and  (not A300) );
 a41415a <=( a41414a  and  a41411a );
 a41416a <=( a41415a  and  a41408a );
 a41420a <=( A167  and  A168 );
 a41421a <=( A170  and  a41420a );
 a41425a <=( (not A202)  and  A201 );
 a41426a <=( (not A166)  and  a41425a );
 a41427a <=( a41426a  and  a41421a );
 a41431a <=( A266  and  (not A265) );
 a41432a <=( A203  and  a41431a );
 a41435a <=( (not A269)  and  A267 );
 a41438a <=( (not A302)  and  (not A300) );
 a41439a <=( a41438a  and  a41435a );
 a41440a <=( a41439a  and  a41432a );
 a41444a <=( A167  and  A168 );
 a41445a <=( A170  and  a41444a );
 a41449a <=( (not A202)  and  A201 );
 a41450a <=( (not A166)  and  a41449a );
 a41451a <=( a41450a  and  a41445a );
 a41455a <=( A266  and  (not A265) );
 a41456a <=( A203  and  a41455a );
 a41459a <=( (not A269)  and  A267 );
 a41462a <=( A299  and  A298 );
 a41463a <=( a41462a  and  a41459a );
 a41464a <=( a41463a  and  a41456a );
 a41468a <=( A167  and  A168 );
 a41469a <=( A170  and  a41468a );
 a41473a <=( (not A202)  and  A201 );
 a41474a <=( (not A166)  and  a41473a );
 a41475a <=( a41474a  and  a41469a );
 a41479a <=( A266  and  (not A265) );
 a41480a <=( A203  and  a41479a );
 a41483a <=( (not A269)  and  A267 );
 a41486a <=( (not A299)  and  (not A298) );
 a41487a <=( a41486a  and  a41483a );
 a41488a <=( a41487a  and  a41480a );
 a41492a <=( A167  and  A168 );
 a41493a <=( A170  and  a41492a );
 a41497a <=( (not A202)  and  A201 );
 a41498a <=( (not A166)  and  a41497a );
 a41499a <=( a41498a  and  a41493a );
 a41503a <=( (not A266)  and  A265 );
 a41504a <=( A203  and  a41503a );
 a41507a <=( A268  and  A267 );
 a41510a <=( A301  and  (not A300) );
 a41511a <=( a41510a  and  a41507a );
 a41512a <=( a41511a  and  a41504a );
 a41516a <=( A167  and  A168 );
 a41517a <=( A170  and  a41516a );
 a41521a <=( (not A202)  and  A201 );
 a41522a <=( (not A166)  and  a41521a );
 a41523a <=( a41522a  and  a41517a );
 a41527a <=( (not A266)  and  A265 );
 a41528a <=( A203  and  a41527a );
 a41531a <=( A268  and  A267 );
 a41534a <=( (not A302)  and  (not A300) );
 a41535a <=( a41534a  and  a41531a );
 a41536a <=( a41535a  and  a41528a );
 a41540a <=( A167  and  A168 );
 a41541a <=( A170  and  a41540a );
 a41545a <=( (not A202)  and  A201 );
 a41546a <=( (not A166)  and  a41545a );
 a41547a <=( a41546a  and  a41541a );
 a41551a <=( (not A266)  and  A265 );
 a41552a <=( A203  and  a41551a );
 a41555a <=( A268  and  A267 );
 a41558a <=( A299  and  A298 );
 a41559a <=( a41558a  and  a41555a );
 a41560a <=( a41559a  and  a41552a );
 a41564a <=( A167  and  A168 );
 a41565a <=( A170  and  a41564a );
 a41569a <=( (not A202)  and  A201 );
 a41570a <=( (not A166)  and  a41569a );
 a41571a <=( a41570a  and  a41565a );
 a41575a <=( (not A266)  and  A265 );
 a41576a <=( A203  and  a41575a );
 a41579a <=( A268  and  A267 );
 a41582a <=( (not A299)  and  (not A298) );
 a41583a <=( a41582a  and  a41579a );
 a41584a <=( a41583a  and  a41576a );
 a41588a <=( A167  and  A168 );
 a41589a <=( A170  and  a41588a );
 a41593a <=( (not A202)  and  A201 );
 a41594a <=( (not A166)  and  a41593a );
 a41595a <=( a41594a  and  a41589a );
 a41599a <=( (not A266)  and  A265 );
 a41600a <=( A203  and  a41599a );
 a41603a <=( (not A269)  and  A267 );
 a41606a <=( A301  and  (not A300) );
 a41607a <=( a41606a  and  a41603a );
 a41608a <=( a41607a  and  a41600a );
 a41612a <=( A167  and  A168 );
 a41613a <=( A170  and  a41612a );
 a41617a <=( (not A202)  and  A201 );
 a41618a <=( (not A166)  and  a41617a );
 a41619a <=( a41618a  and  a41613a );
 a41623a <=( (not A266)  and  A265 );
 a41624a <=( A203  and  a41623a );
 a41627a <=( (not A269)  and  A267 );
 a41630a <=( (not A302)  and  (not A300) );
 a41631a <=( a41630a  and  a41627a );
 a41632a <=( a41631a  and  a41624a );
 a41636a <=( A167  and  A168 );
 a41637a <=( A170  and  a41636a );
 a41641a <=( (not A202)  and  A201 );
 a41642a <=( (not A166)  and  a41641a );
 a41643a <=( a41642a  and  a41637a );
 a41647a <=( (not A266)  and  A265 );
 a41648a <=( A203  and  a41647a );
 a41651a <=( (not A269)  and  A267 );
 a41654a <=( A299  and  A298 );
 a41655a <=( a41654a  and  a41651a );
 a41656a <=( a41655a  and  a41648a );
 a41660a <=( A167  and  A168 );
 a41661a <=( A170  and  a41660a );
 a41665a <=( (not A202)  and  A201 );
 a41666a <=( (not A166)  and  a41665a );
 a41667a <=( a41666a  and  a41661a );
 a41671a <=( (not A266)  and  A265 );
 a41672a <=( A203  and  a41671a );
 a41675a <=( (not A269)  and  A267 );
 a41678a <=( (not A299)  and  (not A298) );
 a41679a <=( a41678a  and  a41675a );
 a41680a <=( a41679a  and  a41672a );
 a41684a <=( A167  and  A168 );
 a41685a <=( A170  and  a41684a );
 a41689a <=( (not A202)  and  A201 );
 a41690a <=( (not A166)  and  a41689a );
 a41691a <=( a41690a  and  a41685a );
 a41695a <=( (not A266)  and  (not A265) );
 a41696a <=( A203  and  a41695a );
 a41699a <=( (not A299)  and  A298 );
 a41702a <=( A301  and  A300 );
 a41703a <=( a41702a  and  a41699a );
 a41704a <=( a41703a  and  a41696a );
 a41708a <=( A167  and  A168 );
 a41709a <=( A170  and  a41708a );
 a41713a <=( (not A202)  and  A201 );
 a41714a <=( (not A166)  and  a41713a );
 a41715a <=( a41714a  and  a41709a );
 a41719a <=( (not A266)  and  (not A265) );
 a41720a <=( A203  and  a41719a );
 a41723a <=( (not A299)  and  A298 );
 a41726a <=( (not A302)  and  A300 );
 a41727a <=( a41726a  and  a41723a );
 a41728a <=( a41727a  and  a41720a );
 a41732a <=( A167  and  A168 );
 a41733a <=( A170  and  a41732a );
 a41737a <=( (not A202)  and  A201 );
 a41738a <=( (not A166)  and  a41737a );
 a41739a <=( a41738a  and  a41733a );
 a41743a <=( (not A266)  and  (not A265) );
 a41744a <=( A203  and  a41743a );
 a41747a <=( A299  and  (not A298) );
 a41750a <=( A301  and  A300 );
 a41751a <=( a41750a  and  a41747a );
 a41752a <=( a41751a  and  a41744a );
 a41756a <=( A167  and  A168 );
 a41757a <=( A170  and  a41756a );
 a41761a <=( (not A202)  and  A201 );
 a41762a <=( (not A166)  and  a41761a );
 a41763a <=( a41762a  and  a41757a );
 a41767a <=( (not A266)  and  (not A265) );
 a41768a <=( A203  and  a41767a );
 a41771a <=( A299  and  (not A298) );
 a41774a <=( (not A302)  and  A300 );
 a41775a <=( a41774a  and  a41771a );
 a41776a <=( a41775a  and  a41768a );
 a41780a <=( A167  and  A168 );
 a41781a <=( A170  and  a41780a );
 a41785a <=( A202  and  (not A201) );
 a41786a <=( (not A166)  and  a41785a );
 a41787a <=( a41786a  and  a41781a );
 a41791a <=( A269  and  (not A268) );
 a41792a <=( A267  and  a41791a );
 a41795a <=( (not A299)  and  A298 );
 a41798a <=( A301  and  A300 );
 a41799a <=( a41798a  and  a41795a );
 a41800a <=( a41799a  and  a41792a );
 a41804a <=( A167  and  A168 );
 a41805a <=( A170  and  a41804a );
 a41809a <=( A202  and  (not A201) );
 a41810a <=( (not A166)  and  a41809a );
 a41811a <=( a41810a  and  a41805a );
 a41815a <=( A269  and  (not A268) );
 a41816a <=( A267  and  a41815a );
 a41819a <=( (not A299)  and  A298 );
 a41822a <=( (not A302)  and  A300 );
 a41823a <=( a41822a  and  a41819a );
 a41824a <=( a41823a  and  a41816a );
 a41828a <=( A167  and  A168 );
 a41829a <=( A170  and  a41828a );
 a41833a <=( A202  and  (not A201) );
 a41834a <=( (not A166)  and  a41833a );
 a41835a <=( a41834a  and  a41829a );
 a41839a <=( A269  and  (not A268) );
 a41840a <=( A267  and  a41839a );
 a41843a <=( A299  and  (not A298) );
 a41846a <=( A301  and  A300 );
 a41847a <=( a41846a  and  a41843a );
 a41848a <=( a41847a  and  a41840a );
 a41852a <=( A167  and  A168 );
 a41853a <=( A170  and  a41852a );
 a41857a <=( A202  and  (not A201) );
 a41858a <=( (not A166)  and  a41857a );
 a41859a <=( a41858a  and  a41853a );
 a41863a <=( A269  and  (not A268) );
 a41864a <=( A267  and  a41863a );
 a41867a <=( A299  and  (not A298) );
 a41870a <=( (not A302)  and  A300 );
 a41871a <=( a41870a  and  a41867a );
 a41872a <=( a41871a  and  a41864a );
 a41876a <=( A167  and  A168 );
 a41877a <=( A170  and  a41876a );
 a41881a <=( A202  and  (not A201) );
 a41882a <=( (not A166)  and  a41881a );
 a41883a <=( a41882a  and  a41877a );
 a41887a <=( A298  and  A268 );
 a41888a <=( (not A267)  and  a41887a );
 a41891a <=( (not A300)  and  (not A299) );
 a41894a <=( A302  and  (not A301) );
 a41895a <=( a41894a  and  a41891a );
 a41896a <=( a41895a  and  a41888a );
 a41900a <=( A167  and  A168 );
 a41901a <=( A170  and  a41900a );
 a41905a <=( A202  and  (not A201) );
 a41906a <=( (not A166)  and  a41905a );
 a41907a <=( a41906a  and  a41901a );
 a41911a <=( (not A298)  and  A268 );
 a41912a <=( (not A267)  and  a41911a );
 a41915a <=( (not A300)  and  A299 );
 a41918a <=( A302  and  (not A301) );
 a41919a <=( a41918a  and  a41915a );
 a41920a <=( a41919a  and  a41912a );
 a41924a <=( A167  and  A168 );
 a41925a <=( A170  and  a41924a );
 a41929a <=( A202  and  (not A201) );
 a41930a <=( (not A166)  and  a41929a );
 a41931a <=( a41930a  and  a41925a );
 a41935a <=( A298  and  (not A269) );
 a41936a <=( (not A267)  and  a41935a );
 a41939a <=( (not A300)  and  (not A299) );
 a41942a <=( A302  and  (not A301) );
 a41943a <=( a41942a  and  a41939a );
 a41944a <=( a41943a  and  a41936a );
 a41948a <=( A167  and  A168 );
 a41949a <=( A170  and  a41948a );
 a41953a <=( A202  and  (not A201) );
 a41954a <=( (not A166)  and  a41953a );
 a41955a <=( a41954a  and  a41949a );
 a41959a <=( (not A298)  and  (not A269) );
 a41960a <=( (not A267)  and  a41959a );
 a41963a <=( (not A300)  and  A299 );
 a41966a <=( A302  and  (not A301) );
 a41967a <=( a41966a  and  a41963a );
 a41968a <=( a41967a  and  a41960a );
 a41972a <=( A167  and  A168 );
 a41973a <=( A170  and  a41972a );
 a41977a <=( A202  and  (not A201) );
 a41978a <=( (not A166)  and  a41977a );
 a41979a <=( a41978a  and  a41973a );
 a41983a <=( A298  and  A266 );
 a41984a <=( A265  and  a41983a );
 a41987a <=( (not A300)  and  (not A299) );
 a41990a <=( A302  and  (not A301) );
 a41991a <=( a41990a  and  a41987a );
 a41992a <=( a41991a  and  a41984a );
 a41996a <=( A167  and  A168 );
 a41997a <=( A170  and  a41996a );
 a42001a <=( A202  and  (not A201) );
 a42002a <=( (not A166)  and  a42001a );
 a42003a <=( a42002a  and  a41997a );
 a42007a <=( (not A298)  and  A266 );
 a42008a <=( A265  and  a42007a );
 a42011a <=( (not A300)  and  A299 );
 a42014a <=( A302  and  (not A301) );
 a42015a <=( a42014a  and  a42011a );
 a42016a <=( a42015a  and  a42008a );
 a42020a <=( A167  and  A168 );
 a42021a <=( A170  and  a42020a );
 a42025a <=( A202  and  (not A201) );
 a42026a <=( (not A166)  and  a42025a );
 a42027a <=( a42026a  and  a42021a );
 a42031a <=( A267  and  A266 );
 a42032a <=( (not A265)  and  a42031a );
 a42035a <=( A300  and  A268 );
 a42038a <=( A302  and  (not A301) );
 a42039a <=( a42038a  and  a42035a );
 a42040a <=( a42039a  and  a42032a );
 a42044a <=( A167  and  A168 );
 a42045a <=( A170  and  a42044a );
 a42049a <=( A202  and  (not A201) );
 a42050a <=( (not A166)  and  a42049a );
 a42051a <=( a42050a  and  a42045a );
 a42055a <=( A267  and  A266 );
 a42056a <=( (not A265)  and  a42055a );
 a42059a <=( A300  and  (not A269) );
 a42062a <=( A302  and  (not A301) );
 a42063a <=( a42062a  and  a42059a );
 a42064a <=( a42063a  and  a42056a );
 a42068a <=( A167  and  A168 );
 a42069a <=( A170  and  a42068a );
 a42073a <=( A202  and  (not A201) );
 a42074a <=( (not A166)  and  a42073a );
 a42075a <=( a42074a  and  a42069a );
 a42079a <=( (not A267)  and  A266 );
 a42080a <=( (not A265)  and  a42079a );
 a42083a <=( A269  and  (not A268) );
 a42086a <=( A301  and  (not A300) );
 a42087a <=( a42086a  and  a42083a );
 a42088a <=( a42087a  and  a42080a );
 a42092a <=( A167  and  A168 );
 a42093a <=( A170  and  a42092a );
 a42097a <=( A202  and  (not A201) );
 a42098a <=( (not A166)  and  a42097a );
 a42099a <=( a42098a  and  a42093a );
 a42103a <=( (not A267)  and  A266 );
 a42104a <=( (not A265)  and  a42103a );
 a42107a <=( A269  and  (not A268) );
 a42110a <=( (not A302)  and  (not A300) );
 a42111a <=( a42110a  and  a42107a );
 a42112a <=( a42111a  and  a42104a );
 a42116a <=( A167  and  A168 );
 a42117a <=( A170  and  a42116a );
 a42121a <=( A202  and  (not A201) );
 a42122a <=( (not A166)  and  a42121a );
 a42123a <=( a42122a  and  a42117a );
 a42127a <=( (not A267)  and  A266 );
 a42128a <=( (not A265)  and  a42127a );
 a42131a <=( A269  and  (not A268) );
 a42134a <=( A299  and  A298 );
 a42135a <=( a42134a  and  a42131a );
 a42136a <=( a42135a  and  a42128a );
 a42140a <=( A167  and  A168 );
 a42141a <=( A170  and  a42140a );
 a42145a <=( A202  and  (not A201) );
 a42146a <=( (not A166)  and  a42145a );
 a42147a <=( a42146a  and  a42141a );
 a42151a <=( (not A267)  and  A266 );
 a42152a <=( (not A265)  and  a42151a );
 a42155a <=( A269  and  (not A268) );
 a42158a <=( (not A299)  and  (not A298) );
 a42159a <=( a42158a  and  a42155a );
 a42160a <=( a42159a  and  a42152a );
 a42164a <=( A167  and  A168 );
 a42165a <=( A170  and  a42164a );
 a42169a <=( A202  and  (not A201) );
 a42170a <=( (not A166)  and  a42169a );
 a42171a <=( a42170a  and  a42165a );
 a42175a <=( A267  and  (not A266) );
 a42176a <=( A265  and  a42175a );
 a42179a <=( A300  and  A268 );
 a42182a <=( A302  and  (not A301) );
 a42183a <=( a42182a  and  a42179a );
 a42184a <=( a42183a  and  a42176a );
 a42188a <=( A167  and  A168 );
 a42189a <=( A170  and  a42188a );
 a42193a <=( A202  and  (not A201) );
 a42194a <=( (not A166)  and  a42193a );
 a42195a <=( a42194a  and  a42189a );
 a42199a <=( A267  and  (not A266) );
 a42200a <=( A265  and  a42199a );
 a42203a <=( A300  and  (not A269) );
 a42206a <=( A302  and  (not A301) );
 a42207a <=( a42206a  and  a42203a );
 a42208a <=( a42207a  and  a42200a );
 a42212a <=( A167  and  A168 );
 a42213a <=( A170  and  a42212a );
 a42217a <=( A202  and  (not A201) );
 a42218a <=( (not A166)  and  a42217a );
 a42219a <=( a42218a  and  a42213a );
 a42223a <=( (not A267)  and  (not A266) );
 a42224a <=( A265  and  a42223a );
 a42227a <=( A269  and  (not A268) );
 a42230a <=( A301  and  (not A300) );
 a42231a <=( a42230a  and  a42227a );
 a42232a <=( a42231a  and  a42224a );
 a42236a <=( A167  and  A168 );
 a42237a <=( A170  and  a42236a );
 a42241a <=( A202  and  (not A201) );
 a42242a <=( (not A166)  and  a42241a );
 a42243a <=( a42242a  and  a42237a );
 a42247a <=( (not A267)  and  (not A266) );
 a42248a <=( A265  and  a42247a );
 a42251a <=( A269  and  (not A268) );
 a42254a <=( (not A302)  and  (not A300) );
 a42255a <=( a42254a  and  a42251a );
 a42256a <=( a42255a  and  a42248a );
 a42260a <=( A167  and  A168 );
 a42261a <=( A170  and  a42260a );
 a42265a <=( A202  and  (not A201) );
 a42266a <=( (not A166)  and  a42265a );
 a42267a <=( a42266a  and  a42261a );
 a42271a <=( (not A267)  and  (not A266) );
 a42272a <=( A265  and  a42271a );
 a42275a <=( A269  and  (not A268) );
 a42278a <=( A299  and  A298 );
 a42279a <=( a42278a  and  a42275a );
 a42280a <=( a42279a  and  a42272a );
 a42284a <=( A167  and  A168 );
 a42285a <=( A170  and  a42284a );
 a42289a <=( A202  and  (not A201) );
 a42290a <=( (not A166)  and  a42289a );
 a42291a <=( a42290a  and  a42285a );
 a42295a <=( (not A267)  and  (not A266) );
 a42296a <=( A265  and  a42295a );
 a42299a <=( A269  and  (not A268) );
 a42302a <=( (not A299)  and  (not A298) );
 a42303a <=( a42302a  and  a42299a );
 a42304a <=( a42303a  and  a42296a );
 a42308a <=( A167  and  A168 );
 a42309a <=( A170  and  a42308a );
 a42313a <=( A202  and  (not A201) );
 a42314a <=( (not A166)  and  a42313a );
 a42315a <=( a42314a  and  a42309a );
 a42319a <=( A298  and  (not A266) );
 a42320a <=( (not A265)  and  a42319a );
 a42323a <=( (not A300)  and  (not A299) );
 a42326a <=( A302  and  (not A301) );
 a42327a <=( a42326a  and  a42323a );
 a42328a <=( a42327a  and  a42320a );
 a42332a <=( A167  and  A168 );
 a42333a <=( A170  and  a42332a );
 a42337a <=( A202  and  (not A201) );
 a42338a <=( (not A166)  and  a42337a );
 a42339a <=( a42338a  and  a42333a );
 a42343a <=( (not A298)  and  (not A266) );
 a42344a <=( (not A265)  and  a42343a );
 a42347a <=( (not A300)  and  A299 );
 a42350a <=( A302  and  (not A301) );
 a42351a <=( a42350a  and  a42347a );
 a42352a <=( a42351a  and  a42344a );
 a42356a <=( A167  and  A168 );
 a42357a <=( A170  and  a42356a );
 a42361a <=( (not A203)  and  (not A201) );
 a42362a <=( (not A166)  and  a42361a );
 a42363a <=( a42362a  and  a42357a );
 a42367a <=( A269  and  (not A268) );
 a42368a <=( A267  and  a42367a );
 a42371a <=( (not A299)  and  A298 );
 a42374a <=( A301  and  A300 );
 a42375a <=( a42374a  and  a42371a );
 a42376a <=( a42375a  and  a42368a );
 a42380a <=( A167  and  A168 );
 a42381a <=( A170  and  a42380a );
 a42385a <=( (not A203)  and  (not A201) );
 a42386a <=( (not A166)  and  a42385a );
 a42387a <=( a42386a  and  a42381a );
 a42391a <=( A269  and  (not A268) );
 a42392a <=( A267  and  a42391a );
 a42395a <=( (not A299)  and  A298 );
 a42398a <=( (not A302)  and  A300 );
 a42399a <=( a42398a  and  a42395a );
 a42400a <=( a42399a  and  a42392a );
 a42404a <=( A167  and  A168 );
 a42405a <=( A170  and  a42404a );
 a42409a <=( (not A203)  and  (not A201) );
 a42410a <=( (not A166)  and  a42409a );
 a42411a <=( a42410a  and  a42405a );
 a42415a <=( A269  and  (not A268) );
 a42416a <=( A267  and  a42415a );
 a42419a <=( A299  and  (not A298) );
 a42422a <=( A301  and  A300 );
 a42423a <=( a42422a  and  a42419a );
 a42424a <=( a42423a  and  a42416a );
 a42428a <=( A167  and  A168 );
 a42429a <=( A170  and  a42428a );
 a42433a <=( (not A203)  and  (not A201) );
 a42434a <=( (not A166)  and  a42433a );
 a42435a <=( a42434a  and  a42429a );
 a42439a <=( A269  and  (not A268) );
 a42440a <=( A267  and  a42439a );
 a42443a <=( A299  and  (not A298) );
 a42446a <=( (not A302)  and  A300 );
 a42447a <=( a42446a  and  a42443a );
 a42448a <=( a42447a  and  a42440a );
 a42452a <=( A167  and  A168 );
 a42453a <=( A170  and  a42452a );
 a42457a <=( (not A203)  and  (not A201) );
 a42458a <=( (not A166)  and  a42457a );
 a42459a <=( a42458a  and  a42453a );
 a42463a <=( A298  and  A268 );
 a42464a <=( (not A267)  and  a42463a );
 a42467a <=( (not A300)  and  (not A299) );
 a42470a <=( A302  and  (not A301) );
 a42471a <=( a42470a  and  a42467a );
 a42472a <=( a42471a  and  a42464a );
 a42476a <=( A167  and  A168 );
 a42477a <=( A170  and  a42476a );
 a42481a <=( (not A203)  and  (not A201) );
 a42482a <=( (not A166)  and  a42481a );
 a42483a <=( a42482a  and  a42477a );
 a42487a <=( (not A298)  and  A268 );
 a42488a <=( (not A267)  and  a42487a );
 a42491a <=( (not A300)  and  A299 );
 a42494a <=( A302  and  (not A301) );
 a42495a <=( a42494a  and  a42491a );
 a42496a <=( a42495a  and  a42488a );
 a42500a <=( A167  and  A168 );
 a42501a <=( A170  and  a42500a );
 a42505a <=( (not A203)  and  (not A201) );
 a42506a <=( (not A166)  and  a42505a );
 a42507a <=( a42506a  and  a42501a );
 a42511a <=( A298  and  (not A269) );
 a42512a <=( (not A267)  and  a42511a );
 a42515a <=( (not A300)  and  (not A299) );
 a42518a <=( A302  and  (not A301) );
 a42519a <=( a42518a  and  a42515a );
 a42520a <=( a42519a  and  a42512a );
 a42524a <=( A167  and  A168 );
 a42525a <=( A170  and  a42524a );
 a42529a <=( (not A203)  and  (not A201) );
 a42530a <=( (not A166)  and  a42529a );
 a42531a <=( a42530a  and  a42525a );
 a42535a <=( (not A298)  and  (not A269) );
 a42536a <=( (not A267)  and  a42535a );
 a42539a <=( (not A300)  and  A299 );
 a42542a <=( A302  and  (not A301) );
 a42543a <=( a42542a  and  a42539a );
 a42544a <=( a42543a  and  a42536a );
 a42548a <=( A167  and  A168 );
 a42549a <=( A170  and  a42548a );
 a42553a <=( (not A203)  and  (not A201) );
 a42554a <=( (not A166)  and  a42553a );
 a42555a <=( a42554a  and  a42549a );
 a42559a <=( A298  and  A266 );
 a42560a <=( A265  and  a42559a );
 a42563a <=( (not A300)  and  (not A299) );
 a42566a <=( A302  and  (not A301) );
 a42567a <=( a42566a  and  a42563a );
 a42568a <=( a42567a  and  a42560a );
 a42572a <=( A167  and  A168 );
 a42573a <=( A170  and  a42572a );
 a42577a <=( (not A203)  and  (not A201) );
 a42578a <=( (not A166)  and  a42577a );
 a42579a <=( a42578a  and  a42573a );
 a42583a <=( (not A298)  and  A266 );
 a42584a <=( A265  and  a42583a );
 a42587a <=( (not A300)  and  A299 );
 a42590a <=( A302  and  (not A301) );
 a42591a <=( a42590a  and  a42587a );
 a42592a <=( a42591a  and  a42584a );
 a42596a <=( A167  and  A168 );
 a42597a <=( A170  and  a42596a );
 a42601a <=( (not A203)  and  (not A201) );
 a42602a <=( (not A166)  and  a42601a );
 a42603a <=( a42602a  and  a42597a );
 a42607a <=( A267  and  A266 );
 a42608a <=( (not A265)  and  a42607a );
 a42611a <=( A300  and  A268 );
 a42614a <=( A302  and  (not A301) );
 a42615a <=( a42614a  and  a42611a );
 a42616a <=( a42615a  and  a42608a );
 a42620a <=( A167  and  A168 );
 a42621a <=( A170  and  a42620a );
 a42625a <=( (not A203)  and  (not A201) );
 a42626a <=( (not A166)  and  a42625a );
 a42627a <=( a42626a  and  a42621a );
 a42631a <=( A267  and  A266 );
 a42632a <=( (not A265)  and  a42631a );
 a42635a <=( A300  and  (not A269) );
 a42638a <=( A302  and  (not A301) );
 a42639a <=( a42638a  and  a42635a );
 a42640a <=( a42639a  and  a42632a );
 a42644a <=( A167  and  A168 );
 a42645a <=( A170  and  a42644a );
 a42649a <=( (not A203)  and  (not A201) );
 a42650a <=( (not A166)  and  a42649a );
 a42651a <=( a42650a  and  a42645a );
 a42655a <=( (not A267)  and  A266 );
 a42656a <=( (not A265)  and  a42655a );
 a42659a <=( A269  and  (not A268) );
 a42662a <=( A301  and  (not A300) );
 a42663a <=( a42662a  and  a42659a );
 a42664a <=( a42663a  and  a42656a );
 a42668a <=( A167  and  A168 );
 a42669a <=( A170  and  a42668a );
 a42673a <=( (not A203)  and  (not A201) );
 a42674a <=( (not A166)  and  a42673a );
 a42675a <=( a42674a  and  a42669a );
 a42679a <=( (not A267)  and  A266 );
 a42680a <=( (not A265)  and  a42679a );
 a42683a <=( A269  and  (not A268) );
 a42686a <=( (not A302)  and  (not A300) );
 a42687a <=( a42686a  and  a42683a );
 a42688a <=( a42687a  and  a42680a );
 a42692a <=( A167  and  A168 );
 a42693a <=( A170  and  a42692a );
 a42697a <=( (not A203)  and  (not A201) );
 a42698a <=( (not A166)  and  a42697a );
 a42699a <=( a42698a  and  a42693a );
 a42703a <=( (not A267)  and  A266 );
 a42704a <=( (not A265)  and  a42703a );
 a42707a <=( A269  and  (not A268) );
 a42710a <=( A299  and  A298 );
 a42711a <=( a42710a  and  a42707a );
 a42712a <=( a42711a  and  a42704a );
 a42716a <=( A167  and  A168 );
 a42717a <=( A170  and  a42716a );
 a42721a <=( (not A203)  and  (not A201) );
 a42722a <=( (not A166)  and  a42721a );
 a42723a <=( a42722a  and  a42717a );
 a42727a <=( (not A267)  and  A266 );
 a42728a <=( (not A265)  and  a42727a );
 a42731a <=( A269  and  (not A268) );
 a42734a <=( (not A299)  and  (not A298) );
 a42735a <=( a42734a  and  a42731a );
 a42736a <=( a42735a  and  a42728a );
 a42740a <=( A167  and  A168 );
 a42741a <=( A170  and  a42740a );
 a42745a <=( (not A203)  and  (not A201) );
 a42746a <=( (not A166)  and  a42745a );
 a42747a <=( a42746a  and  a42741a );
 a42751a <=( A267  and  (not A266) );
 a42752a <=( A265  and  a42751a );
 a42755a <=( A300  and  A268 );
 a42758a <=( A302  and  (not A301) );
 a42759a <=( a42758a  and  a42755a );
 a42760a <=( a42759a  and  a42752a );
 a42764a <=( A167  and  A168 );
 a42765a <=( A170  and  a42764a );
 a42769a <=( (not A203)  and  (not A201) );
 a42770a <=( (not A166)  and  a42769a );
 a42771a <=( a42770a  and  a42765a );
 a42775a <=( A267  and  (not A266) );
 a42776a <=( A265  and  a42775a );
 a42779a <=( A300  and  (not A269) );
 a42782a <=( A302  and  (not A301) );
 a42783a <=( a42782a  and  a42779a );
 a42784a <=( a42783a  and  a42776a );
 a42788a <=( A167  and  A168 );
 a42789a <=( A170  and  a42788a );
 a42793a <=( (not A203)  and  (not A201) );
 a42794a <=( (not A166)  and  a42793a );
 a42795a <=( a42794a  and  a42789a );
 a42799a <=( (not A267)  and  (not A266) );
 a42800a <=( A265  and  a42799a );
 a42803a <=( A269  and  (not A268) );
 a42806a <=( A301  and  (not A300) );
 a42807a <=( a42806a  and  a42803a );
 a42808a <=( a42807a  and  a42800a );
 a42812a <=( A167  and  A168 );
 a42813a <=( A170  and  a42812a );
 a42817a <=( (not A203)  and  (not A201) );
 a42818a <=( (not A166)  and  a42817a );
 a42819a <=( a42818a  and  a42813a );
 a42823a <=( (not A267)  and  (not A266) );
 a42824a <=( A265  and  a42823a );
 a42827a <=( A269  and  (not A268) );
 a42830a <=( (not A302)  and  (not A300) );
 a42831a <=( a42830a  and  a42827a );
 a42832a <=( a42831a  and  a42824a );
 a42836a <=( A167  and  A168 );
 a42837a <=( A170  and  a42836a );
 a42841a <=( (not A203)  and  (not A201) );
 a42842a <=( (not A166)  and  a42841a );
 a42843a <=( a42842a  and  a42837a );
 a42847a <=( (not A267)  and  (not A266) );
 a42848a <=( A265  and  a42847a );
 a42851a <=( A269  and  (not A268) );
 a42854a <=( A299  and  A298 );
 a42855a <=( a42854a  and  a42851a );
 a42856a <=( a42855a  and  a42848a );
 a42860a <=( A167  and  A168 );
 a42861a <=( A170  and  a42860a );
 a42865a <=( (not A203)  and  (not A201) );
 a42866a <=( (not A166)  and  a42865a );
 a42867a <=( a42866a  and  a42861a );
 a42871a <=( (not A267)  and  (not A266) );
 a42872a <=( A265  and  a42871a );
 a42875a <=( A269  and  (not A268) );
 a42878a <=( (not A299)  and  (not A298) );
 a42879a <=( a42878a  and  a42875a );
 a42880a <=( a42879a  and  a42872a );
 a42884a <=( A167  and  A168 );
 a42885a <=( A170  and  a42884a );
 a42889a <=( (not A203)  and  (not A201) );
 a42890a <=( (not A166)  and  a42889a );
 a42891a <=( a42890a  and  a42885a );
 a42895a <=( A298  and  (not A266) );
 a42896a <=( (not A265)  and  a42895a );
 a42899a <=( (not A300)  and  (not A299) );
 a42902a <=( A302  and  (not A301) );
 a42903a <=( a42902a  and  a42899a );
 a42904a <=( a42903a  and  a42896a );
 a42908a <=( A167  and  A168 );
 a42909a <=( A170  and  a42908a );
 a42913a <=( (not A203)  and  (not A201) );
 a42914a <=( (not A166)  and  a42913a );
 a42915a <=( a42914a  and  a42909a );
 a42919a <=( (not A298)  and  (not A266) );
 a42920a <=( (not A265)  and  a42919a );
 a42923a <=( (not A300)  and  A299 );
 a42926a <=( A302  and  (not A301) );
 a42927a <=( a42926a  and  a42923a );
 a42928a <=( a42927a  and  a42920a );
 a42932a <=( A167  and  A168 );
 a42933a <=( A170  and  a42932a );
 a42937a <=( A200  and  A199 );
 a42938a <=( (not A166)  and  a42937a );
 a42939a <=( a42938a  and  a42933a );
 a42943a <=( A269  and  (not A268) );
 a42944a <=( A267  and  a42943a );
 a42947a <=( (not A299)  and  A298 );
 a42950a <=( A301  and  A300 );
 a42951a <=( a42950a  and  a42947a );
 a42952a <=( a42951a  and  a42944a );
 a42956a <=( A167  and  A168 );
 a42957a <=( A170  and  a42956a );
 a42961a <=( A200  and  A199 );
 a42962a <=( (not A166)  and  a42961a );
 a42963a <=( a42962a  and  a42957a );
 a42967a <=( A269  and  (not A268) );
 a42968a <=( A267  and  a42967a );
 a42971a <=( (not A299)  and  A298 );
 a42974a <=( (not A302)  and  A300 );
 a42975a <=( a42974a  and  a42971a );
 a42976a <=( a42975a  and  a42968a );
 a42980a <=( A167  and  A168 );
 a42981a <=( A170  and  a42980a );
 a42985a <=( A200  and  A199 );
 a42986a <=( (not A166)  and  a42985a );
 a42987a <=( a42986a  and  a42981a );
 a42991a <=( A269  and  (not A268) );
 a42992a <=( A267  and  a42991a );
 a42995a <=( A299  and  (not A298) );
 a42998a <=( A301  and  A300 );
 a42999a <=( a42998a  and  a42995a );
 a43000a <=( a42999a  and  a42992a );
 a43004a <=( A167  and  A168 );
 a43005a <=( A170  and  a43004a );
 a43009a <=( A200  and  A199 );
 a43010a <=( (not A166)  and  a43009a );
 a43011a <=( a43010a  and  a43005a );
 a43015a <=( A269  and  (not A268) );
 a43016a <=( A267  and  a43015a );
 a43019a <=( A299  and  (not A298) );
 a43022a <=( (not A302)  and  A300 );
 a43023a <=( a43022a  and  a43019a );
 a43024a <=( a43023a  and  a43016a );
 a43028a <=( A167  and  A168 );
 a43029a <=( A170  and  a43028a );
 a43033a <=( A200  and  A199 );
 a43034a <=( (not A166)  and  a43033a );
 a43035a <=( a43034a  and  a43029a );
 a43039a <=( A298  and  A268 );
 a43040a <=( (not A267)  and  a43039a );
 a43043a <=( (not A300)  and  (not A299) );
 a43046a <=( A302  and  (not A301) );
 a43047a <=( a43046a  and  a43043a );
 a43048a <=( a43047a  and  a43040a );
 a43052a <=( A167  and  A168 );
 a43053a <=( A170  and  a43052a );
 a43057a <=( A200  and  A199 );
 a43058a <=( (not A166)  and  a43057a );
 a43059a <=( a43058a  and  a43053a );
 a43063a <=( (not A298)  and  A268 );
 a43064a <=( (not A267)  and  a43063a );
 a43067a <=( (not A300)  and  A299 );
 a43070a <=( A302  and  (not A301) );
 a43071a <=( a43070a  and  a43067a );
 a43072a <=( a43071a  and  a43064a );
 a43076a <=( A167  and  A168 );
 a43077a <=( A170  and  a43076a );
 a43081a <=( A200  and  A199 );
 a43082a <=( (not A166)  and  a43081a );
 a43083a <=( a43082a  and  a43077a );
 a43087a <=( A298  and  (not A269) );
 a43088a <=( (not A267)  and  a43087a );
 a43091a <=( (not A300)  and  (not A299) );
 a43094a <=( A302  and  (not A301) );
 a43095a <=( a43094a  and  a43091a );
 a43096a <=( a43095a  and  a43088a );
 a43100a <=( A167  and  A168 );
 a43101a <=( A170  and  a43100a );
 a43105a <=( A200  and  A199 );
 a43106a <=( (not A166)  and  a43105a );
 a43107a <=( a43106a  and  a43101a );
 a43111a <=( (not A298)  and  (not A269) );
 a43112a <=( (not A267)  and  a43111a );
 a43115a <=( (not A300)  and  A299 );
 a43118a <=( A302  and  (not A301) );
 a43119a <=( a43118a  and  a43115a );
 a43120a <=( a43119a  and  a43112a );
 a43124a <=( A167  and  A168 );
 a43125a <=( A170  and  a43124a );
 a43129a <=( A200  and  A199 );
 a43130a <=( (not A166)  and  a43129a );
 a43131a <=( a43130a  and  a43125a );
 a43135a <=( A298  and  A266 );
 a43136a <=( A265  and  a43135a );
 a43139a <=( (not A300)  and  (not A299) );
 a43142a <=( A302  and  (not A301) );
 a43143a <=( a43142a  and  a43139a );
 a43144a <=( a43143a  and  a43136a );
 a43148a <=( A167  and  A168 );
 a43149a <=( A170  and  a43148a );
 a43153a <=( A200  and  A199 );
 a43154a <=( (not A166)  and  a43153a );
 a43155a <=( a43154a  and  a43149a );
 a43159a <=( (not A298)  and  A266 );
 a43160a <=( A265  and  a43159a );
 a43163a <=( (not A300)  and  A299 );
 a43166a <=( A302  and  (not A301) );
 a43167a <=( a43166a  and  a43163a );
 a43168a <=( a43167a  and  a43160a );
 a43172a <=( A167  and  A168 );
 a43173a <=( A170  and  a43172a );
 a43177a <=( A200  and  A199 );
 a43178a <=( (not A166)  and  a43177a );
 a43179a <=( a43178a  and  a43173a );
 a43183a <=( A267  and  A266 );
 a43184a <=( (not A265)  and  a43183a );
 a43187a <=( A300  and  A268 );
 a43190a <=( A302  and  (not A301) );
 a43191a <=( a43190a  and  a43187a );
 a43192a <=( a43191a  and  a43184a );
 a43196a <=( A167  and  A168 );
 a43197a <=( A170  and  a43196a );
 a43201a <=( A200  and  A199 );
 a43202a <=( (not A166)  and  a43201a );
 a43203a <=( a43202a  and  a43197a );
 a43207a <=( A267  and  A266 );
 a43208a <=( (not A265)  and  a43207a );
 a43211a <=( A300  and  (not A269) );
 a43214a <=( A302  and  (not A301) );
 a43215a <=( a43214a  and  a43211a );
 a43216a <=( a43215a  and  a43208a );
 a43220a <=( A167  and  A168 );
 a43221a <=( A170  and  a43220a );
 a43225a <=( A200  and  A199 );
 a43226a <=( (not A166)  and  a43225a );
 a43227a <=( a43226a  and  a43221a );
 a43231a <=( (not A267)  and  A266 );
 a43232a <=( (not A265)  and  a43231a );
 a43235a <=( A269  and  (not A268) );
 a43238a <=( A301  and  (not A300) );
 a43239a <=( a43238a  and  a43235a );
 a43240a <=( a43239a  and  a43232a );
 a43244a <=( A167  and  A168 );
 a43245a <=( A170  and  a43244a );
 a43249a <=( A200  and  A199 );
 a43250a <=( (not A166)  and  a43249a );
 a43251a <=( a43250a  and  a43245a );
 a43255a <=( (not A267)  and  A266 );
 a43256a <=( (not A265)  and  a43255a );
 a43259a <=( A269  and  (not A268) );
 a43262a <=( (not A302)  and  (not A300) );
 a43263a <=( a43262a  and  a43259a );
 a43264a <=( a43263a  and  a43256a );
 a43268a <=( A167  and  A168 );
 a43269a <=( A170  and  a43268a );
 a43273a <=( A200  and  A199 );
 a43274a <=( (not A166)  and  a43273a );
 a43275a <=( a43274a  and  a43269a );
 a43279a <=( (not A267)  and  A266 );
 a43280a <=( (not A265)  and  a43279a );
 a43283a <=( A269  and  (not A268) );
 a43286a <=( A299  and  A298 );
 a43287a <=( a43286a  and  a43283a );
 a43288a <=( a43287a  and  a43280a );
 a43292a <=( A167  and  A168 );
 a43293a <=( A170  and  a43292a );
 a43297a <=( A200  and  A199 );
 a43298a <=( (not A166)  and  a43297a );
 a43299a <=( a43298a  and  a43293a );
 a43303a <=( (not A267)  and  A266 );
 a43304a <=( (not A265)  and  a43303a );
 a43307a <=( A269  and  (not A268) );
 a43310a <=( (not A299)  and  (not A298) );
 a43311a <=( a43310a  and  a43307a );
 a43312a <=( a43311a  and  a43304a );
 a43316a <=( A167  and  A168 );
 a43317a <=( A170  and  a43316a );
 a43321a <=( A200  and  A199 );
 a43322a <=( (not A166)  and  a43321a );
 a43323a <=( a43322a  and  a43317a );
 a43327a <=( A267  and  (not A266) );
 a43328a <=( A265  and  a43327a );
 a43331a <=( A300  and  A268 );
 a43334a <=( A302  and  (not A301) );
 a43335a <=( a43334a  and  a43331a );
 a43336a <=( a43335a  and  a43328a );
 a43340a <=( A167  and  A168 );
 a43341a <=( A170  and  a43340a );
 a43345a <=( A200  and  A199 );
 a43346a <=( (not A166)  and  a43345a );
 a43347a <=( a43346a  and  a43341a );
 a43351a <=( A267  and  (not A266) );
 a43352a <=( A265  and  a43351a );
 a43355a <=( A300  and  (not A269) );
 a43358a <=( A302  and  (not A301) );
 a43359a <=( a43358a  and  a43355a );
 a43360a <=( a43359a  and  a43352a );
 a43364a <=( A167  and  A168 );
 a43365a <=( A170  and  a43364a );
 a43369a <=( A200  and  A199 );
 a43370a <=( (not A166)  and  a43369a );
 a43371a <=( a43370a  and  a43365a );
 a43375a <=( (not A267)  and  (not A266) );
 a43376a <=( A265  and  a43375a );
 a43379a <=( A269  and  (not A268) );
 a43382a <=( A301  and  (not A300) );
 a43383a <=( a43382a  and  a43379a );
 a43384a <=( a43383a  and  a43376a );
 a43388a <=( A167  and  A168 );
 a43389a <=( A170  and  a43388a );
 a43393a <=( A200  and  A199 );
 a43394a <=( (not A166)  and  a43393a );
 a43395a <=( a43394a  and  a43389a );
 a43399a <=( (not A267)  and  (not A266) );
 a43400a <=( A265  and  a43399a );
 a43403a <=( A269  and  (not A268) );
 a43406a <=( (not A302)  and  (not A300) );
 a43407a <=( a43406a  and  a43403a );
 a43408a <=( a43407a  and  a43400a );
 a43412a <=( A167  and  A168 );
 a43413a <=( A170  and  a43412a );
 a43417a <=( A200  and  A199 );
 a43418a <=( (not A166)  and  a43417a );
 a43419a <=( a43418a  and  a43413a );
 a43423a <=( (not A267)  and  (not A266) );
 a43424a <=( A265  and  a43423a );
 a43427a <=( A269  and  (not A268) );
 a43430a <=( A299  and  A298 );
 a43431a <=( a43430a  and  a43427a );
 a43432a <=( a43431a  and  a43424a );
 a43436a <=( A167  and  A168 );
 a43437a <=( A170  and  a43436a );
 a43441a <=( A200  and  A199 );
 a43442a <=( (not A166)  and  a43441a );
 a43443a <=( a43442a  and  a43437a );
 a43447a <=( (not A267)  and  (not A266) );
 a43448a <=( A265  and  a43447a );
 a43451a <=( A269  and  (not A268) );
 a43454a <=( (not A299)  and  (not A298) );
 a43455a <=( a43454a  and  a43451a );
 a43456a <=( a43455a  and  a43448a );
 a43460a <=( A167  and  A168 );
 a43461a <=( A170  and  a43460a );
 a43465a <=( A200  and  A199 );
 a43466a <=( (not A166)  and  a43465a );
 a43467a <=( a43466a  and  a43461a );
 a43471a <=( A298  and  (not A266) );
 a43472a <=( (not A265)  and  a43471a );
 a43475a <=( (not A300)  and  (not A299) );
 a43478a <=( A302  and  (not A301) );
 a43479a <=( a43478a  and  a43475a );
 a43480a <=( a43479a  and  a43472a );
 a43484a <=( A167  and  A168 );
 a43485a <=( A170  and  a43484a );
 a43489a <=( A200  and  A199 );
 a43490a <=( (not A166)  and  a43489a );
 a43491a <=( a43490a  and  a43485a );
 a43495a <=( (not A298)  and  (not A266) );
 a43496a <=( (not A265)  and  a43495a );
 a43499a <=( (not A300)  and  A299 );
 a43502a <=( A302  and  (not A301) );
 a43503a <=( a43502a  and  a43499a );
 a43504a <=( a43503a  and  a43496a );
 a43508a <=( A167  and  A168 );
 a43509a <=( A170  and  a43508a );
 a43513a <=( (not A200)  and  (not A199) );
 a43514a <=( (not A166)  and  a43513a );
 a43515a <=( a43514a  and  a43509a );
 a43519a <=( A269  and  (not A268) );
 a43520a <=( A267  and  a43519a );
 a43523a <=( (not A299)  and  A298 );
 a43526a <=( A301  and  A300 );
 a43527a <=( a43526a  and  a43523a );
 a43528a <=( a43527a  and  a43520a );
 a43532a <=( A167  and  A168 );
 a43533a <=( A170  and  a43532a );
 a43537a <=( (not A200)  and  (not A199) );
 a43538a <=( (not A166)  and  a43537a );
 a43539a <=( a43538a  and  a43533a );
 a43543a <=( A269  and  (not A268) );
 a43544a <=( A267  and  a43543a );
 a43547a <=( (not A299)  and  A298 );
 a43550a <=( (not A302)  and  A300 );
 a43551a <=( a43550a  and  a43547a );
 a43552a <=( a43551a  and  a43544a );
 a43556a <=( A167  and  A168 );
 a43557a <=( A170  and  a43556a );
 a43561a <=( (not A200)  and  (not A199) );
 a43562a <=( (not A166)  and  a43561a );
 a43563a <=( a43562a  and  a43557a );
 a43567a <=( A269  and  (not A268) );
 a43568a <=( A267  and  a43567a );
 a43571a <=( A299  and  (not A298) );
 a43574a <=( A301  and  A300 );
 a43575a <=( a43574a  and  a43571a );
 a43576a <=( a43575a  and  a43568a );
 a43580a <=( A167  and  A168 );
 a43581a <=( A170  and  a43580a );
 a43585a <=( (not A200)  and  (not A199) );
 a43586a <=( (not A166)  and  a43585a );
 a43587a <=( a43586a  and  a43581a );
 a43591a <=( A269  and  (not A268) );
 a43592a <=( A267  and  a43591a );
 a43595a <=( A299  and  (not A298) );
 a43598a <=( (not A302)  and  A300 );
 a43599a <=( a43598a  and  a43595a );
 a43600a <=( a43599a  and  a43592a );
 a43604a <=( A167  and  A168 );
 a43605a <=( A170  and  a43604a );
 a43609a <=( (not A200)  and  (not A199) );
 a43610a <=( (not A166)  and  a43609a );
 a43611a <=( a43610a  and  a43605a );
 a43615a <=( A298  and  A268 );
 a43616a <=( (not A267)  and  a43615a );
 a43619a <=( (not A300)  and  (not A299) );
 a43622a <=( A302  and  (not A301) );
 a43623a <=( a43622a  and  a43619a );
 a43624a <=( a43623a  and  a43616a );
 a43628a <=( A167  and  A168 );
 a43629a <=( A170  and  a43628a );
 a43633a <=( (not A200)  and  (not A199) );
 a43634a <=( (not A166)  and  a43633a );
 a43635a <=( a43634a  and  a43629a );
 a43639a <=( (not A298)  and  A268 );
 a43640a <=( (not A267)  and  a43639a );
 a43643a <=( (not A300)  and  A299 );
 a43646a <=( A302  and  (not A301) );
 a43647a <=( a43646a  and  a43643a );
 a43648a <=( a43647a  and  a43640a );
 a43652a <=( A167  and  A168 );
 a43653a <=( A170  and  a43652a );
 a43657a <=( (not A200)  and  (not A199) );
 a43658a <=( (not A166)  and  a43657a );
 a43659a <=( a43658a  and  a43653a );
 a43663a <=( A298  and  (not A269) );
 a43664a <=( (not A267)  and  a43663a );
 a43667a <=( (not A300)  and  (not A299) );
 a43670a <=( A302  and  (not A301) );
 a43671a <=( a43670a  and  a43667a );
 a43672a <=( a43671a  and  a43664a );
 a43676a <=( A167  and  A168 );
 a43677a <=( A170  and  a43676a );
 a43681a <=( (not A200)  and  (not A199) );
 a43682a <=( (not A166)  and  a43681a );
 a43683a <=( a43682a  and  a43677a );
 a43687a <=( (not A298)  and  (not A269) );
 a43688a <=( (not A267)  and  a43687a );
 a43691a <=( (not A300)  and  A299 );
 a43694a <=( A302  and  (not A301) );
 a43695a <=( a43694a  and  a43691a );
 a43696a <=( a43695a  and  a43688a );
 a43700a <=( A167  and  A168 );
 a43701a <=( A170  and  a43700a );
 a43705a <=( (not A200)  and  (not A199) );
 a43706a <=( (not A166)  and  a43705a );
 a43707a <=( a43706a  and  a43701a );
 a43711a <=( A298  and  A266 );
 a43712a <=( A265  and  a43711a );
 a43715a <=( (not A300)  and  (not A299) );
 a43718a <=( A302  and  (not A301) );
 a43719a <=( a43718a  and  a43715a );
 a43720a <=( a43719a  and  a43712a );
 a43724a <=( A167  and  A168 );
 a43725a <=( A170  and  a43724a );
 a43729a <=( (not A200)  and  (not A199) );
 a43730a <=( (not A166)  and  a43729a );
 a43731a <=( a43730a  and  a43725a );
 a43735a <=( (not A298)  and  A266 );
 a43736a <=( A265  and  a43735a );
 a43739a <=( (not A300)  and  A299 );
 a43742a <=( A302  and  (not A301) );
 a43743a <=( a43742a  and  a43739a );
 a43744a <=( a43743a  and  a43736a );
 a43748a <=( A167  and  A168 );
 a43749a <=( A170  and  a43748a );
 a43753a <=( (not A200)  and  (not A199) );
 a43754a <=( (not A166)  and  a43753a );
 a43755a <=( a43754a  and  a43749a );
 a43759a <=( A267  and  A266 );
 a43760a <=( (not A265)  and  a43759a );
 a43763a <=( A300  and  A268 );
 a43766a <=( A302  and  (not A301) );
 a43767a <=( a43766a  and  a43763a );
 a43768a <=( a43767a  and  a43760a );
 a43772a <=( A167  and  A168 );
 a43773a <=( A170  and  a43772a );
 a43777a <=( (not A200)  and  (not A199) );
 a43778a <=( (not A166)  and  a43777a );
 a43779a <=( a43778a  and  a43773a );
 a43783a <=( A267  and  A266 );
 a43784a <=( (not A265)  and  a43783a );
 a43787a <=( A300  and  (not A269) );
 a43790a <=( A302  and  (not A301) );
 a43791a <=( a43790a  and  a43787a );
 a43792a <=( a43791a  and  a43784a );
 a43796a <=( A167  and  A168 );
 a43797a <=( A170  and  a43796a );
 a43801a <=( (not A200)  and  (not A199) );
 a43802a <=( (not A166)  and  a43801a );
 a43803a <=( a43802a  and  a43797a );
 a43807a <=( (not A267)  and  A266 );
 a43808a <=( (not A265)  and  a43807a );
 a43811a <=( A269  and  (not A268) );
 a43814a <=( A301  and  (not A300) );
 a43815a <=( a43814a  and  a43811a );
 a43816a <=( a43815a  and  a43808a );
 a43820a <=( A167  and  A168 );
 a43821a <=( A170  and  a43820a );
 a43825a <=( (not A200)  and  (not A199) );
 a43826a <=( (not A166)  and  a43825a );
 a43827a <=( a43826a  and  a43821a );
 a43831a <=( (not A267)  and  A266 );
 a43832a <=( (not A265)  and  a43831a );
 a43835a <=( A269  and  (not A268) );
 a43838a <=( (not A302)  and  (not A300) );
 a43839a <=( a43838a  and  a43835a );
 a43840a <=( a43839a  and  a43832a );
 a43844a <=( A167  and  A168 );
 a43845a <=( A170  and  a43844a );
 a43849a <=( (not A200)  and  (not A199) );
 a43850a <=( (not A166)  and  a43849a );
 a43851a <=( a43850a  and  a43845a );
 a43855a <=( (not A267)  and  A266 );
 a43856a <=( (not A265)  and  a43855a );
 a43859a <=( A269  and  (not A268) );
 a43862a <=( A299  and  A298 );
 a43863a <=( a43862a  and  a43859a );
 a43864a <=( a43863a  and  a43856a );
 a43868a <=( A167  and  A168 );
 a43869a <=( A170  and  a43868a );
 a43873a <=( (not A200)  and  (not A199) );
 a43874a <=( (not A166)  and  a43873a );
 a43875a <=( a43874a  and  a43869a );
 a43879a <=( (not A267)  and  A266 );
 a43880a <=( (not A265)  and  a43879a );
 a43883a <=( A269  and  (not A268) );
 a43886a <=( (not A299)  and  (not A298) );
 a43887a <=( a43886a  and  a43883a );
 a43888a <=( a43887a  and  a43880a );
 a43892a <=( A167  and  A168 );
 a43893a <=( A170  and  a43892a );
 a43897a <=( (not A200)  and  (not A199) );
 a43898a <=( (not A166)  and  a43897a );
 a43899a <=( a43898a  and  a43893a );
 a43903a <=( A267  and  (not A266) );
 a43904a <=( A265  and  a43903a );
 a43907a <=( A300  and  A268 );
 a43910a <=( A302  and  (not A301) );
 a43911a <=( a43910a  and  a43907a );
 a43912a <=( a43911a  and  a43904a );
 a43916a <=( A167  and  A168 );
 a43917a <=( A170  and  a43916a );
 a43921a <=( (not A200)  and  (not A199) );
 a43922a <=( (not A166)  and  a43921a );
 a43923a <=( a43922a  and  a43917a );
 a43927a <=( A267  and  (not A266) );
 a43928a <=( A265  and  a43927a );
 a43931a <=( A300  and  (not A269) );
 a43934a <=( A302  and  (not A301) );
 a43935a <=( a43934a  and  a43931a );
 a43936a <=( a43935a  and  a43928a );
 a43940a <=( A167  and  A168 );
 a43941a <=( A170  and  a43940a );
 a43945a <=( (not A200)  and  (not A199) );
 a43946a <=( (not A166)  and  a43945a );
 a43947a <=( a43946a  and  a43941a );
 a43951a <=( (not A267)  and  (not A266) );
 a43952a <=( A265  and  a43951a );
 a43955a <=( A269  and  (not A268) );
 a43958a <=( A301  and  (not A300) );
 a43959a <=( a43958a  and  a43955a );
 a43960a <=( a43959a  and  a43952a );
 a43964a <=( A167  and  A168 );
 a43965a <=( A170  and  a43964a );
 a43969a <=( (not A200)  and  (not A199) );
 a43970a <=( (not A166)  and  a43969a );
 a43971a <=( a43970a  and  a43965a );
 a43975a <=( (not A267)  and  (not A266) );
 a43976a <=( A265  and  a43975a );
 a43979a <=( A269  and  (not A268) );
 a43982a <=( (not A302)  and  (not A300) );
 a43983a <=( a43982a  and  a43979a );
 a43984a <=( a43983a  and  a43976a );
 a43988a <=( A167  and  A168 );
 a43989a <=( A170  and  a43988a );
 a43993a <=( (not A200)  and  (not A199) );
 a43994a <=( (not A166)  and  a43993a );
 a43995a <=( a43994a  and  a43989a );
 a43999a <=( (not A267)  and  (not A266) );
 a44000a <=( A265  and  a43999a );
 a44003a <=( A269  and  (not A268) );
 a44006a <=( A299  and  A298 );
 a44007a <=( a44006a  and  a44003a );
 a44008a <=( a44007a  and  a44000a );
 a44012a <=( A167  and  A168 );
 a44013a <=( A170  and  a44012a );
 a44017a <=( (not A200)  and  (not A199) );
 a44018a <=( (not A166)  and  a44017a );
 a44019a <=( a44018a  and  a44013a );
 a44023a <=( (not A267)  and  (not A266) );
 a44024a <=( A265  and  a44023a );
 a44027a <=( A269  and  (not A268) );
 a44030a <=( (not A299)  and  (not A298) );
 a44031a <=( a44030a  and  a44027a );
 a44032a <=( a44031a  and  a44024a );
 a44036a <=( A167  and  A168 );
 a44037a <=( A170  and  a44036a );
 a44041a <=( (not A200)  and  (not A199) );
 a44042a <=( (not A166)  and  a44041a );
 a44043a <=( a44042a  and  a44037a );
 a44047a <=( A298  and  (not A266) );
 a44048a <=( (not A265)  and  a44047a );
 a44051a <=( (not A300)  and  (not A299) );
 a44054a <=( A302  and  (not A301) );
 a44055a <=( a44054a  and  a44051a );
 a44056a <=( a44055a  and  a44048a );
 a44060a <=( A167  and  A168 );
 a44061a <=( A170  and  a44060a );
 a44065a <=( (not A200)  and  (not A199) );
 a44066a <=( (not A166)  and  a44065a );
 a44067a <=( a44066a  and  a44061a );
 a44071a <=( (not A298)  and  (not A266) );
 a44072a <=( (not A265)  and  a44071a );
 a44075a <=( (not A300)  and  A299 );
 a44078a <=( A302  and  (not A301) );
 a44079a <=( a44078a  and  a44075a );
 a44080a <=( a44079a  and  a44072a );
 a44084a <=( (not A167)  and  A168 );
 a44085a <=( A170  and  a44084a );
 a44089a <=( (not A202)  and  A201 );
 a44090a <=( A166  and  a44089a );
 a44091a <=( a44090a  and  a44085a );
 a44095a <=( A268  and  (not A267) );
 a44096a <=( A203  and  a44095a );
 a44099a <=( (not A299)  and  A298 );
 a44102a <=( A301  and  A300 );
 a44103a <=( a44102a  and  a44099a );
 a44104a <=( a44103a  and  a44096a );
 a44108a <=( (not A167)  and  A168 );
 a44109a <=( A170  and  a44108a );
 a44113a <=( (not A202)  and  A201 );
 a44114a <=( A166  and  a44113a );
 a44115a <=( a44114a  and  a44109a );
 a44119a <=( A268  and  (not A267) );
 a44120a <=( A203  and  a44119a );
 a44123a <=( (not A299)  and  A298 );
 a44126a <=( (not A302)  and  A300 );
 a44127a <=( a44126a  and  a44123a );
 a44128a <=( a44127a  and  a44120a );
 a44132a <=( (not A167)  and  A168 );
 a44133a <=( A170  and  a44132a );
 a44137a <=( (not A202)  and  A201 );
 a44138a <=( A166  and  a44137a );
 a44139a <=( a44138a  and  a44133a );
 a44143a <=( A268  and  (not A267) );
 a44144a <=( A203  and  a44143a );
 a44147a <=( A299  and  (not A298) );
 a44150a <=( A301  and  A300 );
 a44151a <=( a44150a  and  a44147a );
 a44152a <=( a44151a  and  a44144a );
 a44156a <=( (not A167)  and  A168 );
 a44157a <=( A170  and  a44156a );
 a44161a <=( (not A202)  and  A201 );
 a44162a <=( A166  and  a44161a );
 a44163a <=( a44162a  and  a44157a );
 a44167a <=( A268  and  (not A267) );
 a44168a <=( A203  and  a44167a );
 a44171a <=( A299  and  (not A298) );
 a44174a <=( (not A302)  and  A300 );
 a44175a <=( a44174a  and  a44171a );
 a44176a <=( a44175a  and  a44168a );
 a44180a <=( (not A167)  and  A168 );
 a44181a <=( A170  and  a44180a );
 a44185a <=( (not A202)  and  A201 );
 a44186a <=( A166  and  a44185a );
 a44187a <=( a44186a  and  a44181a );
 a44191a <=( (not A269)  and  (not A267) );
 a44192a <=( A203  and  a44191a );
 a44195a <=( (not A299)  and  A298 );
 a44198a <=( A301  and  A300 );
 a44199a <=( a44198a  and  a44195a );
 a44200a <=( a44199a  and  a44192a );
 a44204a <=( (not A167)  and  A168 );
 a44205a <=( A170  and  a44204a );
 a44209a <=( (not A202)  and  A201 );
 a44210a <=( A166  and  a44209a );
 a44211a <=( a44210a  and  a44205a );
 a44215a <=( (not A269)  and  (not A267) );
 a44216a <=( A203  and  a44215a );
 a44219a <=( (not A299)  and  A298 );
 a44222a <=( (not A302)  and  A300 );
 a44223a <=( a44222a  and  a44219a );
 a44224a <=( a44223a  and  a44216a );
 a44228a <=( (not A167)  and  A168 );
 a44229a <=( A170  and  a44228a );
 a44233a <=( (not A202)  and  A201 );
 a44234a <=( A166  and  a44233a );
 a44235a <=( a44234a  and  a44229a );
 a44239a <=( (not A269)  and  (not A267) );
 a44240a <=( A203  and  a44239a );
 a44243a <=( A299  and  (not A298) );
 a44246a <=( A301  and  A300 );
 a44247a <=( a44246a  and  a44243a );
 a44248a <=( a44247a  and  a44240a );
 a44252a <=( (not A167)  and  A168 );
 a44253a <=( A170  and  a44252a );
 a44257a <=( (not A202)  and  A201 );
 a44258a <=( A166  and  a44257a );
 a44259a <=( a44258a  and  a44253a );
 a44263a <=( (not A269)  and  (not A267) );
 a44264a <=( A203  and  a44263a );
 a44267a <=( A299  and  (not A298) );
 a44270a <=( (not A302)  and  A300 );
 a44271a <=( a44270a  and  a44267a );
 a44272a <=( a44271a  and  a44264a );
 a44276a <=( (not A167)  and  A168 );
 a44277a <=( A170  and  a44276a );
 a44281a <=( (not A202)  and  A201 );
 a44282a <=( A166  and  a44281a );
 a44283a <=( a44282a  and  a44277a );
 a44287a <=( A266  and  A265 );
 a44288a <=( A203  and  a44287a );
 a44291a <=( (not A299)  and  A298 );
 a44294a <=( A301  and  A300 );
 a44295a <=( a44294a  and  a44291a );
 a44296a <=( a44295a  and  a44288a );
 a44300a <=( (not A167)  and  A168 );
 a44301a <=( A170  and  a44300a );
 a44305a <=( (not A202)  and  A201 );
 a44306a <=( A166  and  a44305a );
 a44307a <=( a44306a  and  a44301a );
 a44311a <=( A266  and  A265 );
 a44312a <=( A203  and  a44311a );
 a44315a <=( (not A299)  and  A298 );
 a44318a <=( (not A302)  and  A300 );
 a44319a <=( a44318a  and  a44315a );
 a44320a <=( a44319a  and  a44312a );
 a44324a <=( (not A167)  and  A168 );
 a44325a <=( A170  and  a44324a );
 a44329a <=( (not A202)  and  A201 );
 a44330a <=( A166  and  a44329a );
 a44331a <=( a44330a  and  a44325a );
 a44335a <=( A266  and  A265 );
 a44336a <=( A203  and  a44335a );
 a44339a <=( A299  and  (not A298) );
 a44342a <=( A301  and  A300 );
 a44343a <=( a44342a  and  a44339a );
 a44344a <=( a44343a  and  a44336a );
 a44348a <=( (not A167)  and  A168 );
 a44349a <=( A170  and  a44348a );
 a44353a <=( (not A202)  and  A201 );
 a44354a <=( A166  and  a44353a );
 a44355a <=( a44354a  and  a44349a );
 a44359a <=( A266  and  A265 );
 a44360a <=( A203  and  a44359a );
 a44363a <=( A299  and  (not A298) );
 a44366a <=( (not A302)  and  A300 );
 a44367a <=( a44366a  and  a44363a );
 a44368a <=( a44367a  and  a44360a );
 a44372a <=( (not A167)  and  A168 );
 a44373a <=( A170  and  a44372a );
 a44377a <=( (not A202)  and  A201 );
 a44378a <=( A166  and  a44377a );
 a44379a <=( a44378a  and  a44373a );
 a44383a <=( A266  and  (not A265) );
 a44384a <=( A203  and  a44383a );
 a44387a <=( A268  and  A267 );
 a44390a <=( A301  and  (not A300) );
 a44391a <=( a44390a  and  a44387a );
 a44392a <=( a44391a  and  a44384a );
 a44396a <=( (not A167)  and  A168 );
 a44397a <=( A170  and  a44396a );
 a44401a <=( (not A202)  and  A201 );
 a44402a <=( A166  and  a44401a );
 a44403a <=( a44402a  and  a44397a );
 a44407a <=( A266  and  (not A265) );
 a44408a <=( A203  and  a44407a );
 a44411a <=( A268  and  A267 );
 a44414a <=( (not A302)  and  (not A300) );
 a44415a <=( a44414a  and  a44411a );
 a44416a <=( a44415a  and  a44408a );
 a44420a <=( (not A167)  and  A168 );
 a44421a <=( A170  and  a44420a );
 a44425a <=( (not A202)  and  A201 );
 a44426a <=( A166  and  a44425a );
 a44427a <=( a44426a  and  a44421a );
 a44431a <=( A266  and  (not A265) );
 a44432a <=( A203  and  a44431a );
 a44435a <=( A268  and  A267 );
 a44438a <=( A299  and  A298 );
 a44439a <=( a44438a  and  a44435a );
 a44440a <=( a44439a  and  a44432a );
 a44444a <=( (not A167)  and  A168 );
 a44445a <=( A170  and  a44444a );
 a44449a <=( (not A202)  and  A201 );
 a44450a <=( A166  and  a44449a );
 a44451a <=( a44450a  and  a44445a );
 a44455a <=( A266  and  (not A265) );
 a44456a <=( A203  and  a44455a );
 a44459a <=( A268  and  A267 );
 a44462a <=( (not A299)  and  (not A298) );
 a44463a <=( a44462a  and  a44459a );
 a44464a <=( a44463a  and  a44456a );
 a44468a <=( (not A167)  and  A168 );
 a44469a <=( A170  and  a44468a );
 a44473a <=( (not A202)  and  A201 );
 a44474a <=( A166  and  a44473a );
 a44475a <=( a44474a  and  a44469a );
 a44479a <=( A266  and  (not A265) );
 a44480a <=( A203  and  a44479a );
 a44483a <=( (not A269)  and  A267 );
 a44486a <=( A301  and  (not A300) );
 a44487a <=( a44486a  and  a44483a );
 a44488a <=( a44487a  and  a44480a );
 a44492a <=( (not A167)  and  A168 );
 a44493a <=( A170  and  a44492a );
 a44497a <=( (not A202)  and  A201 );
 a44498a <=( A166  and  a44497a );
 a44499a <=( a44498a  and  a44493a );
 a44503a <=( A266  and  (not A265) );
 a44504a <=( A203  and  a44503a );
 a44507a <=( (not A269)  and  A267 );
 a44510a <=( (not A302)  and  (not A300) );
 a44511a <=( a44510a  and  a44507a );
 a44512a <=( a44511a  and  a44504a );
 a44516a <=( (not A167)  and  A168 );
 a44517a <=( A170  and  a44516a );
 a44521a <=( (not A202)  and  A201 );
 a44522a <=( A166  and  a44521a );
 a44523a <=( a44522a  and  a44517a );
 a44527a <=( A266  and  (not A265) );
 a44528a <=( A203  and  a44527a );
 a44531a <=( (not A269)  and  A267 );
 a44534a <=( A299  and  A298 );
 a44535a <=( a44534a  and  a44531a );
 a44536a <=( a44535a  and  a44528a );
 a44540a <=( (not A167)  and  A168 );
 a44541a <=( A170  and  a44540a );
 a44545a <=( (not A202)  and  A201 );
 a44546a <=( A166  and  a44545a );
 a44547a <=( a44546a  and  a44541a );
 a44551a <=( A266  and  (not A265) );
 a44552a <=( A203  and  a44551a );
 a44555a <=( (not A269)  and  A267 );
 a44558a <=( (not A299)  and  (not A298) );
 a44559a <=( a44558a  and  a44555a );
 a44560a <=( a44559a  and  a44552a );
 a44564a <=( (not A167)  and  A168 );
 a44565a <=( A170  and  a44564a );
 a44569a <=( (not A202)  and  A201 );
 a44570a <=( A166  and  a44569a );
 a44571a <=( a44570a  and  a44565a );
 a44575a <=( (not A266)  and  A265 );
 a44576a <=( A203  and  a44575a );
 a44579a <=( A268  and  A267 );
 a44582a <=( A301  and  (not A300) );
 a44583a <=( a44582a  and  a44579a );
 a44584a <=( a44583a  and  a44576a );
 a44588a <=( (not A167)  and  A168 );
 a44589a <=( A170  and  a44588a );
 a44593a <=( (not A202)  and  A201 );
 a44594a <=( A166  and  a44593a );
 a44595a <=( a44594a  and  a44589a );
 a44599a <=( (not A266)  and  A265 );
 a44600a <=( A203  and  a44599a );
 a44603a <=( A268  and  A267 );
 a44606a <=( (not A302)  and  (not A300) );
 a44607a <=( a44606a  and  a44603a );
 a44608a <=( a44607a  and  a44600a );
 a44612a <=( (not A167)  and  A168 );
 a44613a <=( A170  and  a44612a );
 a44617a <=( (not A202)  and  A201 );
 a44618a <=( A166  and  a44617a );
 a44619a <=( a44618a  and  a44613a );
 a44623a <=( (not A266)  and  A265 );
 a44624a <=( A203  and  a44623a );
 a44627a <=( A268  and  A267 );
 a44630a <=( A299  and  A298 );
 a44631a <=( a44630a  and  a44627a );
 a44632a <=( a44631a  and  a44624a );
 a44636a <=( (not A167)  and  A168 );
 a44637a <=( A170  and  a44636a );
 a44641a <=( (not A202)  and  A201 );
 a44642a <=( A166  and  a44641a );
 a44643a <=( a44642a  and  a44637a );
 a44647a <=( (not A266)  and  A265 );
 a44648a <=( A203  and  a44647a );
 a44651a <=( A268  and  A267 );
 a44654a <=( (not A299)  and  (not A298) );
 a44655a <=( a44654a  and  a44651a );
 a44656a <=( a44655a  and  a44648a );
 a44660a <=( (not A167)  and  A168 );
 a44661a <=( A170  and  a44660a );
 a44665a <=( (not A202)  and  A201 );
 a44666a <=( A166  and  a44665a );
 a44667a <=( a44666a  and  a44661a );
 a44671a <=( (not A266)  and  A265 );
 a44672a <=( A203  and  a44671a );
 a44675a <=( (not A269)  and  A267 );
 a44678a <=( A301  and  (not A300) );
 a44679a <=( a44678a  and  a44675a );
 a44680a <=( a44679a  and  a44672a );
 a44684a <=( (not A167)  and  A168 );
 a44685a <=( A170  and  a44684a );
 a44689a <=( (not A202)  and  A201 );
 a44690a <=( A166  and  a44689a );
 a44691a <=( a44690a  and  a44685a );
 a44695a <=( (not A266)  and  A265 );
 a44696a <=( A203  and  a44695a );
 a44699a <=( (not A269)  and  A267 );
 a44702a <=( (not A302)  and  (not A300) );
 a44703a <=( a44702a  and  a44699a );
 a44704a <=( a44703a  and  a44696a );
 a44708a <=( (not A167)  and  A168 );
 a44709a <=( A170  and  a44708a );
 a44713a <=( (not A202)  and  A201 );
 a44714a <=( A166  and  a44713a );
 a44715a <=( a44714a  and  a44709a );
 a44719a <=( (not A266)  and  A265 );
 a44720a <=( A203  and  a44719a );
 a44723a <=( (not A269)  and  A267 );
 a44726a <=( A299  and  A298 );
 a44727a <=( a44726a  and  a44723a );
 a44728a <=( a44727a  and  a44720a );
 a44732a <=( (not A167)  and  A168 );
 a44733a <=( A170  and  a44732a );
 a44737a <=( (not A202)  and  A201 );
 a44738a <=( A166  and  a44737a );
 a44739a <=( a44738a  and  a44733a );
 a44743a <=( (not A266)  and  A265 );
 a44744a <=( A203  and  a44743a );
 a44747a <=( (not A269)  and  A267 );
 a44750a <=( (not A299)  and  (not A298) );
 a44751a <=( a44750a  and  a44747a );
 a44752a <=( a44751a  and  a44744a );
 a44756a <=( (not A167)  and  A168 );
 a44757a <=( A170  and  a44756a );
 a44761a <=( (not A202)  and  A201 );
 a44762a <=( A166  and  a44761a );
 a44763a <=( a44762a  and  a44757a );
 a44767a <=( (not A266)  and  (not A265) );
 a44768a <=( A203  and  a44767a );
 a44771a <=( (not A299)  and  A298 );
 a44774a <=( A301  and  A300 );
 a44775a <=( a44774a  and  a44771a );
 a44776a <=( a44775a  and  a44768a );
 a44780a <=( (not A167)  and  A168 );
 a44781a <=( A170  and  a44780a );
 a44785a <=( (not A202)  and  A201 );
 a44786a <=( A166  and  a44785a );
 a44787a <=( a44786a  and  a44781a );
 a44791a <=( (not A266)  and  (not A265) );
 a44792a <=( A203  and  a44791a );
 a44795a <=( (not A299)  and  A298 );
 a44798a <=( (not A302)  and  A300 );
 a44799a <=( a44798a  and  a44795a );
 a44800a <=( a44799a  and  a44792a );
 a44804a <=( (not A167)  and  A168 );
 a44805a <=( A170  and  a44804a );
 a44809a <=( (not A202)  and  A201 );
 a44810a <=( A166  and  a44809a );
 a44811a <=( a44810a  and  a44805a );
 a44815a <=( (not A266)  and  (not A265) );
 a44816a <=( A203  and  a44815a );
 a44819a <=( A299  and  (not A298) );
 a44822a <=( A301  and  A300 );
 a44823a <=( a44822a  and  a44819a );
 a44824a <=( a44823a  and  a44816a );
 a44828a <=( (not A167)  and  A168 );
 a44829a <=( A170  and  a44828a );
 a44833a <=( (not A202)  and  A201 );
 a44834a <=( A166  and  a44833a );
 a44835a <=( a44834a  and  a44829a );
 a44839a <=( (not A266)  and  (not A265) );
 a44840a <=( A203  and  a44839a );
 a44843a <=( A299  and  (not A298) );
 a44846a <=( (not A302)  and  A300 );
 a44847a <=( a44846a  and  a44843a );
 a44848a <=( a44847a  and  a44840a );
 a44852a <=( (not A167)  and  A168 );
 a44853a <=( A170  and  a44852a );
 a44857a <=( A202  and  (not A201) );
 a44858a <=( A166  and  a44857a );
 a44859a <=( a44858a  and  a44853a );
 a44863a <=( A269  and  (not A268) );
 a44864a <=( A267  and  a44863a );
 a44867a <=( (not A299)  and  A298 );
 a44870a <=( A301  and  A300 );
 a44871a <=( a44870a  and  a44867a );
 a44872a <=( a44871a  and  a44864a );
 a44876a <=( (not A167)  and  A168 );
 a44877a <=( A170  and  a44876a );
 a44881a <=( A202  and  (not A201) );
 a44882a <=( A166  and  a44881a );
 a44883a <=( a44882a  and  a44877a );
 a44887a <=( A269  and  (not A268) );
 a44888a <=( A267  and  a44887a );
 a44891a <=( (not A299)  and  A298 );
 a44894a <=( (not A302)  and  A300 );
 a44895a <=( a44894a  and  a44891a );
 a44896a <=( a44895a  and  a44888a );
 a44900a <=( (not A167)  and  A168 );
 a44901a <=( A170  and  a44900a );
 a44905a <=( A202  and  (not A201) );
 a44906a <=( A166  and  a44905a );
 a44907a <=( a44906a  and  a44901a );
 a44911a <=( A269  and  (not A268) );
 a44912a <=( A267  and  a44911a );
 a44915a <=( A299  and  (not A298) );
 a44918a <=( A301  and  A300 );
 a44919a <=( a44918a  and  a44915a );
 a44920a <=( a44919a  and  a44912a );
 a44924a <=( (not A167)  and  A168 );
 a44925a <=( A170  and  a44924a );
 a44929a <=( A202  and  (not A201) );
 a44930a <=( A166  and  a44929a );
 a44931a <=( a44930a  and  a44925a );
 a44935a <=( A269  and  (not A268) );
 a44936a <=( A267  and  a44935a );
 a44939a <=( A299  and  (not A298) );
 a44942a <=( (not A302)  and  A300 );
 a44943a <=( a44942a  and  a44939a );
 a44944a <=( a44943a  and  a44936a );
 a44948a <=( (not A167)  and  A168 );
 a44949a <=( A170  and  a44948a );
 a44953a <=( A202  and  (not A201) );
 a44954a <=( A166  and  a44953a );
 a44955a <=( a44954a  and  a44949a );
 a44959a <=( A298  and  A268 );
 a44960a <=( (not A267)  and  a44959a );
 a44963a <=( (not A300)  and  (not A299) );
 a44966a <=( A302  and  (not A301) );
 a44967a <=( a44966a  and  a44963a );
 a44968a <=( a44967a  and  a44960a );
 a44972a <=( (not A167)  and  A168 );
 a44973a <=( A170  and  a44972a );
 a44977a <=( A202  and  (not A201) );
 a44978a <=( A166  and  a44977a );
 a44979a <=( a44978a  and  a44973a );
 a44983a <=( (not A298)  and  A268 );
 a44984a <=( (not A267)  and  a44983a );
 a44987a <=( (not A300)  and  A299 );
 a44990a <=( A302  and  (not A301) );
 a44991a <=( a44990a  and  a44987a );
 a44992a <=( a44991a  and  a44984a );
 a44996a <=( (not A167)  and  A168 );
 a44997a <=( A170  and  a44996a );
 a45001a <=( A202  and  (not A201) );
 a45002a <=( A166  and  a45001a );
 a45003a <=( a45002a  and  a44997a );
 a45007a <=( A298  and  (not A269) );
 a45008a <=( (not A267)  and  a45007a );
 a45011a <=( (not A300)  and  (not A299) );
 a45014a <=( A302  and  (not A301) );
 a45015a <=( a45014a  and  a45011a );
 a45016a <=( a45015a  and  a45008a );
 a45020a <=( (not A167)  and  A168 );
 a45021a <=( A170  and  a45020a );
 a45025a <=( A202  and  (not A201) );
 a45026a <=( A166  and  a45025a );
 a45027a <=( a45026a  and  a45021a );
 a45031a <=( (not A298)  and  (not A269) );
 a45032a <=( (not A267)  and  a45031a );
 a45035a <=( (not A300)  and  A299 );
 a45038a <=( A302  and  (not A301) );
 a45039a <=( a45038a  and  a45035a );
 a45040a <=( a45039a  and  a45032a );
 a45044a <=( (not A167)  and  A168 );
 a45045a <=( A170  and  a45044a );
 a45049a <=( A202  and  (not A201) );
 a45050a <=( A166  and  a45049a );
 a45051a <=( a45050a  and  a45045a );
 a45055a <=( A298  and  A266 );
 a45056a <=( A265  and  a45055a );
 a45059a <=( (not A300)  and  (not A299) );
 a45062a <=( A302  and  (not A301) );
 a45063a <=( a45062a  and  a45059a );
 a45064a <=( a45063a  and  a45056a );
 a45068a <=( (not A167)  and  A168 );
 a45069a <=( A170  and  a45068a );
 a45073a <=( A202  and  (not A201) );
 a45074a <=( A166  and  a45073a );
 a45075a <=( a45074a  and  a45069a );
 a45079a <=( (not A298)  and  A266 );
 a45080a <=( A265  and  a45079a );
 a45083a <=( (not A300)  and  A299 );
 a45086a <=( A302  and  (not A301) );
 a45087a <=( a45086a  and  a45083a );
 a45088a <=( a45087a  and  a45080a );
 a45092a <=( (not A167)  and  A168 );
 a45093a <=( A170  and  a45092a );
 a45097a <=( A202  and  (not A201) );
 a45098a <=( A166  and  a45097a );
 a45099a <=( a45098a  and  a45093a );
 a45103a <=( A267  and  A266 );
 a45104a <=( (not A265)  and  a45103a );
 a45107a <=( A300  and  A268 );
 a45110a <=( A302  and  (not A301) );
 a45111a <=( a45110a  and  a45107a );
 a45112a <=( a45111a  and  a45104a );
 a45116a <=( (not A167)  and  A168 );
 a45117a <=( A170  and  a45116a );
 a45121a <=( A202  and  (not A201) );
 a45122a <=( A166  and  a45121a );
 a45123a <=( a45122a  and  a45117a );
 a45127a <=( A267  and  A266 );
 a45128a <=( (not A265)  and  a45127a );
 a45131a <=( A300  and  (not A269) );
 a45134a <=( A302  and  (not A301) );
 a45135a <=( a45134a  and  a45131a );
 a45136a <=( a45135a  and  a45128a );
 a45140a <=( (not A167)  and  A168 );
 a45141a <=( A170  and  a45140a );
 a45145a <=( A202  and  (not A201) );
 a45146a <=( A166  and  a45145a );
 a45147a <=( a45146a  and  a45141a );
 a45151a <=( (not A267)  and  A266 );
 a45152a <=( (not A265)  and  a45151a );
 a45155a <=( A269  and  (not A268) );
 a45158a <=( A301  and  (not A300) );
 a45159a <=( a45158a  and  a45155a );
 a45160a <=( a45159a  and  a45152a );
 a45164a <=( (not A167)  and  A168 );
 a45165a <=( A170  and  a45164a );
 a45169a <=( A202  and  (not A201) );
 a45170a <=( A166  and  a45169a );
 a45171a <=( a45170a  and  a45165a );
 a45175a <=( (not A267)  and  A266 );
 a45176a <=( (not A265)  and  a45175a );
 a45179a <=( A269  and  (not A268) );
 a45182a <=( (not A302)  and  (not A300) );
 a45183a <=( a45182a  and  a45179a );
 a45184a <=( a45183a  and  a45176a );
 a45188a <=( (not A167)  and  A168 );
 a45189a <=( A170  and  a45188a );
 a45193a <=( A202  and  (not A201) );
 a45194a <=( A166  and  a45193a );
 a45195a <=( a45194a  and  a45189a );
 a45199a <=( (not A267)  and  A266 );
 a45200a <=( (not A265)  and  a45199a );
 a45203a <=( A269  and  (not A268) );
 a45206a <=( A299  and  A298 );
 a45207a <=( a45206a  and  a45203a );
 a45208a <=( a45207a  and  a45200a );
 a45212a <=( (not A167)  and  A168 );
 a45213a <=( A170  and  a45212a );
 a45217a <=( A202  and  (not A201) );
 a45218a <=( A166  and  a45217a );
 a45219a <=( a45218a  and  a45213a );
 a45223a <=( (not A267)  and  A266 );
 a45224a <=( (not A265)  and  a45223a );
 a45227a <=( A269  and  (not A268) );
 a45230a <=( (not A299)  and  (not A298) );
 a45231a <=( a45230a  and  a45227a );
 a45232a <=( a45231a  and  a45224a );
 a45236a <=( (not A167)  and  A168 );
 a45237a <=( A170  and  a45236a );
 a45241a <=( A202  and  (not A201) );
 a45242a <=( A166  and  a45241a );
 a45243a <=( a45242a  and  a45237a );
 a45247a <=( A267  and  (not A266) );
 a45248a <=( A265  and  a45247a );
 a45251a <=( A300  and  A268 );
 a45254a <=( A302  and  (not A301) );
 a45255a <=( a45254a  and  a45251a );
 a45256a <=( a45255a  and  a45248a );
 a45260a <=( (not A167)  and  A168 );
 a45261a <=( A170  and  a45260a );
 a45265a <=( A202  and  (not A201) );
 a45266a <=( A166  and  a45265a );
 a45267a <=( a45266a  and  a45261a );
 a45271a <=( A267  and  (not A266) );
 a45272a <=( A265  and  a45271a );
 a45275a <=( A300  and  (not A269) );
 a45278a <=( A302  and  (not A301) );
 a45279a <=( a45278a  and  a45275a );
 a45280a <=( a45279a  and  a45272a );
 a45284a <=( (not A167)  and  A168 );
 a45285a <=( A170  and  a45284a );
 a45289a <=( A202  and  (not A201) );
 a45290a <=( A166  and  a45289a );
 a45291a <=( a45290a  and  a45285a );
 a45295a <=( (not A267)  and  (not A266) );
 a45296a <=( A265  and  a45295a );
 a45299a <=( A269  and  (not A268) );
 a45302a <=( A301  and  (not A300) );
 a45303a <=( a45302a  and  a45299a );
 a45304a <=( a45303a  and  a45296a );
 a45308a <=( (not A167)  and  A168 );
 a45309a <=( A170  and  a45308a );
 a45313a <=( A202  and  (not A201) );
 a45314a <=( A166  and  a45313a );
 a45315a <=( a45314a  and  a45309a );
 a45319a <=( (not A267)  and  (not A266) );
 a45320a <=( A265  and  a45319a );
 a45323a <=( A269  and  (not A268) );
 a45326a <=( (not A302)  and  (not A300) );
 a45327a <=( a45326a  and  a45323a );
 a45328a <=( a45327a  and  a45320a );
 a45332a <=( (not A167)  and  A168 );
 a45333a <=( A170  and  a45332a );
 a45337a <=( A202  and  (not A201) );
 a45338a <=( A166  and  a45337a );
 a45339a <=( a45338a  and  a45333a );
 a45343a <=( (not A267)  and  (not A266) );
 a45344a <=( A265  and  a45343a );
 a45347a <=( A269  and  (not A268) );
 a45350a <=( A299  and  A298 );
 a45351a <=( a45350a  and  a45347a );
 a45352a <=( a45351a  and  a45344a );
 a45356a <=( (not A167)  and  A168 );
 a45357a <=( A170  and  a45356a );
 a45361a <=( A202  and  (not A201) );
 a45362a <=( A166  and  a45361a );
 a45363a <=( a45362a  and  a45357a );
 a45367a <=( (not A267)  and  (not A266) );
 a45368a <=( A265  and  a45367a );
 a45371a <=( A269  and  (not A268) );
 a45374a <=( (not A299)  and  (not A298) );
 a45375a <=( a45374a  and  a45371a );
 a45376a <=( a45375a  and  a45368a );
 a45380a <=( (not A167)  and  A168 );
 a45381a <=( A170  and  a45380a );
 a45385a <=( A202  and  (not A201) );
 a45386a <=( A166  and  a45385a );
 a45387a <=( a45386a  and  a45381a );
 a45391a <=( A298  and  (not A266) );
 a45392a <=( (not A265)  and  a45391a );
 a45395a <=( (not A300)  and  (not A299) );
 a45398a <=( A302  and  (not A301) );
 a45399a <=( a45398a  and  a45395a );
 a45400a <=( a45399a  and  a45392a );
 a45404a <=( (not A167)  and  A168 );
 a45405a <=( A170  and  a45404a );
 a45409a <=( A202  and  (not A201) );
 a45410a <=( A166  and  a45409a );
 a45411a <=( a45410a  and  a45405a );
 a45415a <=( (not A298)  and  (not A266) );
 a45416a <=( (not A265)  and  a45415a );
 a45419a <=( (not A300)  and  A299 );
 a45422a <=( A302  and  (not A301) );
 a45423a <=( a45422a  and  a45419a );
 a45424a <=( a45423a  and  a45416a );
 a45428a <=( (not A167)  and  A168 );
 a45429a <=( A170  and  a45428a );
 a45433a <=( (not A203)  and  (not A201) );
 a45434a <=( A166  and  a45433a );
 a45435a <=( a45434a  and  a45429a );
 a45439a <=( A269  and  (not A268) );
 a45440a <=( A267  and  a45439a );
 a45443a <=( (not A299)  and  A298 );
 a45446a <=( A301  and  A300 );
 a45447a <=( a45446a  and  a45443a );
 a45448a <=( a45447a  and  a45440a );
 a45452a <=( (not A167)  and  A168 );
 a45453a <=( A170  and  a45452a );
 a45457a <=( (not A203)  and  (not A201) );
 a45458a <=( A166  and  a45457a );
 a45459a <=( a45458a  and  a45453a );
 a45463a <=( A269  and  (not A268) );
 a45464a <=( A267  and  a45463a );
 a45467a <=( (not A299)  and  A298 );
 a45470a <=( (not A302)  and  A300 );
 a45471a <=( a45470a  and  a45467a );
 a45472a <=( a45471a  and  a45464a );
 a45476a <=( (not A167)  and  A168 );
 a45477a <=( A170  and  a45476a );
 a45481a <=( (not A203)  and  (not A201) );
 a45482a <=( A166  and  a45481a );
 a45483a <=( a45482a  and  a45477a );
 a45487a <=( A269  and  (not A268) );
 a45488a <=( A267  and  a45487a );
 a45491a <=( A299  and  (not A298) );
 a45494a <=( A301  and  A300 );
 a45495a <=( a45494a  and  a45491a );
 a45496a <=( a45495a  and  a45488a );
 a45500a <=( (not A167)  and  A168 );
 a45501a <=( A170  and  a45500a );
 a45505a <=( (not A203)  and  (not A201) );
 a45506a <=( A166  and  a45505a );
 a45507a <=( a45506a  and  a45501a );
 a45511a <=( A269  and  (not A268) );
 a45512a <=( A267  and  a45511a );
 a45515a <=( A299  and  (not A298) );
 a45518a <=( (not A302)  and  A300 );
 a45519a <=( a45518a  and  a45515a );
 a45520a <=( a45519a  and  a45512a );
 a45524a <=( (not A167)  and  A168 );
 a45525a <=( A170  and  a45524a );
 a45529a <=( (not A203)  and  (not A201) );
 a45530a <=( A166  and  a45529a );
 a45531a <=( a45530a  and  a45525a );
 a45535a <=( A298  and  A268 );
 a45536a <=( (not A267)  and  a45535a );
 a45539a <=( (not A300)  and  (not A299) );
 a45542a <=( A302  and  (not A301) );
 a45543a <=( a45542a  and  a45539a );
 a45544a <=( a45543a  and  a45536a );
 a45548a <=( (not A167)  and  A168 );
 a45549a <=( A170  and  a45548a );
 a45553a <=( (not A203)  and  (not A201) );
 a45554a <=( A166  and  a45553a );
 a45555a <=( a45554a  and  a45549a );
 a45559a <=( (not A298)  and  A268 );
 a45560a <=( (not A267)  and  a45559a );
 a45563a <=( (not A300)  and  A299 );
 a45566a <=( A302  and  (not A301) );
 a45567a <=( a45566a  and  a45563a );
 a45568a <=( a45567a  and  a45560a );
 a45572a <=( (not A167)  and  A168 );
 a45573a <=( A170  and  a45572a );
 a45577a <=( (not A203)  and  (not A201) );
 a45578a <=( A166  and  a45577a );
 a45579a <=( a45578a  and  a45573a );
 a45583a <=( A298  and  (not A269) );
 a45584a <=( (not A267)  and  a45583a );
 a45587a <=( (not A300)  and  (not A299) );
 a45590a <=( A302  and  (not A301) );
 a45591a <=( a45590a  and  a45587a );
 a45592a <=( a45591a  and  a45584a );
 a45596a <=( (not A167)  and  A168 );
 a45597a <=( A170  and  a45596a );
 a45601a <=( (not A203)  and  (not A201) );
 a45602a <=( A166  and  a45601a );
 a45603a <=( a45602a  and  a45597a );
 a45607a <=( (not A298)  and  (not A269) );
 a45608a <=( (not A267)  and  a45607a );
 a45611a <=( (not A300)  and  A299 );
 a45614a <=( A302  and  (not A301) );
 a45615a <=( a45614a  and  a45611a );
 a45616a <=( a45615a  and  a45608a );
 a45620a <=( (not A167)  and  A168 );
 a45621a <=( A170  and  a45620a );
 a45625a <=( (not A203)  and  (not A201) );
 a45626a <=( A166  and  a45625a );
 a45627a <=( a45626a  and  a45621a );
 a45631a <=( A298  and  A266 );
 a45632a <=( A265  and  a45631a );
 a45635a <=( (not A300)  and  (not A299) );
 a45638a <=( A302  and  (not A301) );
 a45639a <=( a45638a  and  a45635a );
 a45640a <=( a45639a  and  a45632a );
 a45644a <=( (not A167)  and  A168 );
 a45645a <=( A170  and  a45644a );
 a45649a <=( (not A203)  and  (not A201) );
 a45650a <=( A166  and  a45649a );
 a45651a <=( a45650a  and  a45645a );
 a45655a <=( (not A298)  and  A266 );
 a45656a <=( A265  and  a45655a );
 a45659a <=( (not A300)  and  A299 );
 a45662a <=( A302  and  (not A301) );
 a45663a <=( a45662a  and  a45659a );
 a45664a <=( a45663a  and  a45656a );
 a45668a <=( (not A167)  and  A168 );
 a45669a <=( A170  and  a45668a );
 a45673a <=( (not A203)  and  (not A201) );
 a45674a <=( A166  and  a45673a );
 a45675a <=( a45674a  and  a45669a );
 a45679a <=( A267  and  A266 );
 a45680a <=( (not A265)  and  a45679a );
 a45683a <=( A300  and  A268 );
 a45686a <=( A302  and  (not A301) );
 a45687a <=( a45686a  and  a45683a );
 a45688a <=( a45687a  and  a45680a );
 a45692a <=( (not A167)  and  A168 );
 a45693a <=( A170  and  a45692a );
 a45697a <=( (not A203)  and  (not A201) );
 a45698a <=( A166  and  a45697a );
 a45699a <=( a45698a  and  a45693a );
 a45703a <=( A267  and  A266 );
 a45704a <=( (not A265)  and  a45703a );
 a45707a <=( A300  and  (not A269) );
 a45710a <=( A302  and  (not A301) );
 a45711a <=( a45710a  and  a45707a );
 a45712a <=( a45711a  and  a45704a );
 a45716a <=( (not A167)  and  A168 );
 a45717a <=( A170  and  a45716a );
 a45721a <=( (not A203)  and  (not A201) );
 a45722a <=( A166  and  a45721a );
 a45723a <=( a45722a  and  a45717a );
 a45727a <=( (not A267)  and  A266 );
 a45728a <=( (not A265)  and  a45727a );
 a45731a <=( A269  and  (not A268) );
 a45734a <=( A301  and  (not A300) );
 a45735a <=( a45734a  and  a45731a );
 a45736a <=( a45735a  and  a45728a );
 a45740a <=( (not A167)  and  A168 );
 a45741a <=( A170  and  a45740a );
 a45745a <=( (not A203)  and  (not A201) );
 a45746a <=( A166  and  a45745a );
 a45747a <=( a45746a  and  a45741a );
 a45751a <=( (not A267)  and  A266 );
 a45752a <=( (not A265)  and  a45751a );
 a45755a <=( A269  and  (not A268) );
 a45758a <=( (not A302)  and  (not A300) );
 a45759a <=( a45758a  and  a45755a );
 a45760a <=( a45759a  and  a45752a );
 a45764a <=( (not A167)  and  A168 );
 a45765a <=( A170  and  a45764a );
 a45769a <=( (not A203)  and  (not A201) );
 a45770a <=( A166  and  a45769a );
 a45771a <=( a45770a  and  a45765a );
 a45775a <=( (not A267)  and  A266 );
 a45776a <=( (not A265)  and  a45775a );
 a45779a <=( A269  and  (not A268) );
 a45782a <=( A299  and  A298 );
 a45783a <=( a45782a  and  a45779a );
 a45784a <=( a45783a  and  a45776a );
 a45788a <=( (not A167)  and  A168 );
 a45789a <=( A170  and  a45788a );
 a45793a <=( (not A203)  and  (not A201) );
 a45794a <=( A166  and  a45793a );
 a45795a <=( a45794a  and  a45789a );
 a45799a <=( (not A267)  and  A266 );
 a45800a <=( (not A265)  and  a45799a );
 a45803a <=( A269  and  (not A268) );
 a45806a <=( (not A299)  and  (not A298) );
 a45807a <=( a45806a  and  a45803a );
 a45808a <=( a45807a  and  a45800a );
 a45812a <=( (not A167)  and  A168 );
 a45813a <=( A170  and  a45812a );
 a45817a <=( (not A203)  and  (not A201) );
 a45818a <=( A166  and  a45817a );
 a45819a <=( a45818a  and  a45813a );
 a45823a <=( A267  and  (not A266) );
 a45824a <=( A265  and  a45823a );
 a45827a <=( A300  and  A268 );
 a45830a <=( A302  and  (not A301) );
 a45831a <=( a45830a  and  a45827a );
 a45832a <=( a45831a  and  a45824a );
 a45836a <=( (not A167)  and  A168 );
 a45837a <=( A170  and  a45836a );
 a45841a <=( (not A203)  and  (not A201) );
 a45842a <=( A166  and  a45841a );
 a45843a <=( a45842a  and  a45837a );
 a45847a <=( A267  and  (not A266) );
 a45848a <=( A265  and  a45847a );
 a45851a <=( A300  and  (not A269) );
 a45854a <=( A302  and  (not A301) );
 a45855a <=( a45854a  and  a45851a );
 a45856a <=( a45855a  and  a45848a );
 a45860a <=( (not A167)  and  A168 );
 a45861a <=( A170  and  a45860a );
 a45865a <=( (not A203)  and  (not A201) );
 a45866a <=( A166  and  a45865a );
 a45867a <=( a45866a  and  a45861a );
 a45871a <=( (not A267)  and  (not A266) );
 a45872a <=( A265  and  a45871a );
 a45875a <=( A269  and  (not A268) );
 a45878a <=( A301  and  (not A300) );
 a45879a <=( a45878a  and  a45875a );
 a45880a <=( a45879a  and  a45872a );
 a45884a <=( (not A167)  and  A168 );
 a45885a <=( A170  and  a45884a );
 a45889a <=( (not A203)  and  (not A201) );
 a45890a <=( A166  and  a45889a );
 a45891a <=( a45890a  and  a45885a );
 a45895a <=( (not A267)  and  (not A266) );
 a45896a <=( A265  and  a45895a );
 a45899a <=( A269  and  (not A268) );
 a45902a <=( (not A302)  and  (not A300) );
 a45903a <=( a45902a  and  a45899a );
 a45904a <=( a45903a  and  a45896a );
 a45908a <=( (not A167)  and  A168 );
 a45909a <=( A170  and  a45908a );
 a45913a <=( (not A203)  and  (not A201) );
 a45914a <=( A166  and  a45913a );
 a45915a <=( a45914a  and  a45909a );
 a45919a <=( (not A267)  and  (not A266) );
 a45920a <=( A265  and  a45919a );
 a45923a <=( A269  and  (not A268) );
 a45926a <=( A299  and  A298 );
 a45927a <=( a45926a  and  a45923a );
 a45928a <=( a45927a  and  a45920a );
 a45932a <=( (not A167)  and  A168 );
 a45933a <=( A170  and  a45932a );
 a45937a <=( (not A203)  and  (not A201) );
 a45938a <=( A166  and  a45937a );
 a45939a <=( a45938a  and  a45933a );
 a45943a <=( (not A267)  and  (not A266) );
 a45944a <=( A265  and  a45943a );
 a45947a <=( A269  and  (not A268) );
 a45950a <=( (not A299)  and  (not A298) );
 a45951a <=( a45950a  and  a45947a );
 a45952a <=( a45951a  and  a45944a );
 a45956a <=( (not A167)  and  A168 );
 a45957a <=( A170  and  a45956a );
 a45961a <=( (not A203)  and  (not A201) );
 a45962a <=( A166  and  a45961a );
 a45963a <=( a45962a  and  a45957a );
 a45967a <=( A298  and  (not A266) );
 a45968a <=( (not A265)  and  a45967a );
 a45971a <=( (not A300)  and  (not A299) );
 a45974a <=( A302  and  (not A301) );
 a45975a <=( a45974a  and  a45971a );
 a45976a <=( a45975a  and  a45968a );
 a45980a <=( (not A167)  and  A168 );
 a45981a <=( A170  and  a45980a );
 a45985a <=( (not A203)  and  (not A201) );
 a45986a <=( A166  and  a45985a );
 a45987a <=( a45986a  and  a45981a );
 a45991a <=( (not A298)  and  (not A266) );
 a45992a <=( (not A265)  and  a45991a );
 a45995a <=( (not A300)  and  A299 );
 a45998a <=( A302  and  (not A301) );
 a45999a <=( a45998a  and  a45995a );
 a46000a <=( a45999a  and  a45992a );
 a46004a <=( (not A167)  and  A168 );
 a46005a <=( A170  and  a46004a );
 a46009a <=( A200  and  A199 );
 a46010a <=( A166  and  a46009a );
 a46011a <=( a46010a  and  a46005a );
 a46015a <=( A269  and  (not A268) );
 a46016a <=( A267  and  a46015a );
 a46019a <=( (not A299)  and  A298 );
 a46022a <=( A301  and  A300 );
 a46023a <=( a46022a  and  a46019a );
 a46024a <=( a46023a  and  a46016a );
 a46028a <=( (not A167)  and  A168 );
 a46029a <=( A170  and  a46028a );
 a46033a <=( A200  and  A199 );
 a46034a <=( A166  and  a46033a );
 a46035a <=( a46034a  and  a46029a );
 a46039a <=( A269  and  (not A268) );
 a46040a <=( A267  and  a46039a );
 a46043a <=( (not A299)  and  A298 );
 a46046a <=( (not A302)  and  A300 );
 a46047a <=( a46046a  and  a46043a );
 a46048a <=( a46047a  and  a46040a );
 a46052a <=( (not A167)  and  A168 );
 a46053a <=( A170  and  a46052a );
 a46057a <=( A200  and  A199 );
 a46058a <=( A166  and  a46057a );
 a46059a <=( a46058a  and  a46053a );
 a46063a <=( A269  and  (not A268) );
 a46064a <=( A267  and  a46063a );
 a46067a <=( A299  and  (not A298) );
 a46070a <=( A301  and  A300 );
 a46071a <=( a46070a  and  a46067a );
 a46072a <=( a46071a  and  a46064a );
 a46076a <=( (not A167)  and  A168 );
 a46077a <=( A170  and  a46076a );
 a46081a <=( A200  and  A199 );
 a46082a <=( A166  and  a46081a );
 a46083a <=( a46082a  and  a46077a );
 a46087a <=( A269  and  (not A268) );
 a46088a <=( A267  and  a46087a );
 a46091a <=( A299  and  (not A298) );
 a46094a <=( (not A302)  and  A300 );
 a46095a <=( a46094a  and  a46091a );
 a46096a <=( a46095a  and  a46088a );
 a46100a <=( (not A167)  and  A168 );
 a46101a <=( A170  and  a46100a );
 a46105a <=( A200  and  A199 );
 a46106a <=( A166  and  a46105a );
 a46107a <=( a46106a  and  a46101a );
 a46111a <=( A298  and  A268 );
 a46112a <=( (not A267)  and  a46111a );
 a46115a <=( (not A300)  and  (not A299) );
 a46118a <=( A302  and  (not A301) );
 a46119a <=( a46118a  and  a46115a );
 a46120a <=( a46119a  and  a46112a );
 a46124a <=( (not A167)  and  A168 );
 a46125a <=( A170  and  a46124a );
 a46129a <=( A200  and  A199 );
 a46130a <=( A166  and  a46129a );
 a46131a <=( a46130a  and  a46125a );
 a46135a <=( (not A298)  and  A268 );
 a46136a <=( (not A267)  and  a46135a );
 a46139a <=( (not A300)  and  A299 );
 a46142a <=( A302  and  (not A301) );
 a46143a <=( a46142a  and  a46139a );
 a46144a <=( a46143a  and  a46136a );
 a46148a <=( (not A167)  and  A168 );
 a46149a <=( A170  and  a46148a );
 a46153a <=( A200  and  A199 );
 a46154a <=( A166  and  a46153a );
 a46155a <=( a46154a  and  a46149a );
 a46159a <=( A298  and  (not A269) );
 a46160a <=( (not A267)  and  a46159a );
 a46163a <=( (not A300)  and  (not A299) );
 a46166a <=( A302  and  (not A301) );
 a46167a <=( a46166a  and  a46163a );
 a46168a <=( a46167a  and  a46160a );
 a46172a <=( (not A167)  and  A168 );
 a46173a <=( A170  and  a46172a );
 a46177a <=( A200  and  A199 );
 a46178a <=( A166  and  a46177a );
 a46179a <=( a46178a  and  a46173a );
 a46183a <=( (not A298)  and  (not A269) );
 a46184a <=( (not A267)  and  a46183a );
 a46187a <=( (not A300)  and  A299 );
 a46190a <=( A302  and  (not A301) );
 a46191a <=( a46190a  and  a46187a );
 a46192a <=( a46191a  and  a46184a );
 a46196a <=( (not A167)  and  A168 );
 a46197a <=( A170  and  a46196a );
 a46201a <=( A200  and  A199 );
 a46202a <=( A166  and  a46201a );
 a46203a <=( a46202a  and  a46197a );
 a46207a <=( A298  and  A266 );
 a46208a <=( A265  and  a46207a );
 a46211a <=( (not A300)  and  (not A299) );
 a46214a <=( A302  and  (not A301) );
 a46215a <=( a46214a  and  a46211a );
 a46216a <=( a46215a  and  a46208a );
 a46220a <=( (not A167)  and  A168 );
 a46221a <=( A170  and  a46220a );
 a46225a <=( A200  and  A199 );
 a46226a <=( A166  and  a46225a );
 a46227a <=( a46226a  and  a46221a );
 a46231a <=( (not A298)  and  A266 );
 a46232a <=( A265  and  a46231a );
 a46235a <=( (not A300)  and  A299 );
 a46238a <=( A302  and  (not A301) );
 a46239a <=( a46238a  and  a46235a );
 a46240a <=( a46239a  and  a46232a );
 a46244a <=( (not A167)  and  A168 );
 a46245a <=( A170  and  a46244a );
 a46249a <=( A200  and  A199 );
 a46250a <=( A166  and  a46249a );
 a46251a <=( a46250a  and  a46245a );
 a46255a <=( A267  and  A266 );
 a46256a <=( (not A265)  and  a46255a );
 a46259a <=( A300  and  A268 );
 a46262a <=( A302  and  (not A301) );
 a46263a <=( a46262a  and  a46259a );
 a46264a <=( a46263a  and  a46256a );
 a46268a <=( (not A167)  and  A168 );
 a46269a <=( A170  and  a46268a );
 a46273a <=( A200  and  A199 );
 a46274a <=( A166  and  a46273a );
 a46275a <=( a46274a  and  a46269a );
 a46279a <=( A267  and  A266 );
 a46280a <=( (not A265)  and  a46279a );
 a46283a <=( A300  and  (not A269) );
 a46286a <=( A302  and  (not A301) );
 a46287a <=( a46286a  and  a46283a );
 a46288a <=( a46287a  and  a46280a );
 a46292a <=( (not A167)  and  A168 );
 a46293a <=( A170  and  a46292a );
 a46297a <=( A200  and  A199 );
 a46298a <=( A166  and  a46297a );
 a46299a <=( a46298a  and  a46293a );
 a46303a <=( (not A267)  and  A266 );
 a46304a <=( (not A265)  and  a46303a );
 a46307a <=( A269  and  (not A268) );
 a46310a <=( A301  and  (not A300) );
 a46311a <=( a46310a  and  a46307a );
 a46312a <=( a46311a  and  a46304a );
 a46316a <=( (not A167)  and  A168 );
 a46317a <=( A170  and  a46316a );
 a46321a <=( A200  and  A199 );
 a46322a <=( A166  and  a46321a );
 a46323a <=( a46322a  and  a46317a );
 a46327a <=( (not A267)  and  A266 );
 a46328a <=( (not A265)  and  a46327a );
 a46331a <=( A269  and  (not A268) );
 a46334a <=( (not A302)  and  (not A300) );
 a46335a <=( a46334a  and  a46331a );
 a46336a <=( a46335a  and  a46328a );
 a46340a <=( (not A167)  and  A168 );
 a46341a <=( A170  and  a46340a );
 a46345a <=( A200  and  A199 );
 a46346a <=( A166  and  a46345a );
 a46347a <=( a46346a  and  a46341a );
 a46351a <=( (not A267)  and  A266 );
 a46352a <=( (not A265)  and  a46351a );
 a46355a <=( A269  and  (not A268) );
 a46358a <=( A299  and  A298 );
 a46359a <=( a46358a  and  a46355a );
 a46360a <=( a46359a  and  a46352a );
 a46364a <=( (not A167)  and  A168 );
 a46365a <=( A170  and  a46364a );
 a46369a <=( A200  and  A199 );
 a46370a <=( A166  and  a46369a );
 a46371a <=( a46370a  and  a46365a );
 a46375a <=( (not A267)  and  A266 );
 a46376a <=( (not A265)  and  a46375a );
 a46379a <=( A269  and  (not A268) );
 a46382a <=( (not A299)  and  (not A298) );
 a46383a <=( a46382a  and  a46379a );
 a46384a <=( a46383a  and  a46376a );
 a46388a <=( (not A167)  and  A168 );
 a46389a <=( A170  and  a46388a );
 a46393a <=( A200  and  A199 );
 a46394a <=( A166  and  a46393a );
 a46395a <=( a46394a  and  a46389a );
 a46399a <=( A267  and  (not A266) );
 a46400a <=( A265  and  a46399a );
 a46403a <=( A300  and  A268 );
 a46406a <=( A302  and  (not A301) );
 a46407a <=( a46406a  and  a46403a );
 a46408a <=( a46407a  and  a46400a );
 a46412a <=( (not A167)  and  A168 );
 a46413a <=( A170  and  a46412a );
 a46417a <=( A200  and  A199 );
 a46418a <=( A166  and  a46417a );
 a46419a <=( a46418a  and  a46413a );
 a46423a <=( A267  and  (not A266) );
 a46424a <=( A265  and  a46423a );
 a46427a <=( A300  and  (not A269) );
 a46430a <=( A302  and  (not A301) );
 a46431a <=( a46430a  and  a46427a );
 a46432a <=( a46431a  and  a46424a );
 a46436a <=( (not A167)  and  A168 );
 a46437a <=( A170  and  a46436a );
 a46441a <=( A200  and  A199 );
 a46442a <=( A166  and  a46441a );
 a46443a <=( a46442a  and  a46437a );
 a46447a <=( (not A267)  and  (not A266) );
 a46448a <=( A265  and  a46447a );
 a46451a <=( A269  and  (not A268) );
 a46454a <=( A301  and  (not A300) );
 a46455a <=( a46454a  and  a46451a );
 a46456a <=( a46455a  and  a46448a );
 a46460a <=( (not A167)  and  A168 );
 a46461a <=( A170  and  a46460a );
 a46465a <=( A200  and  A199 );
 a46466a <=( A166  and  a46465a );
 a46467a <=( a46466a  and  a46461a );
 a46471a <=( (not A267)  and  (not A266) );
 a46472a <=( A265  and  a46471a );
 a46475a <=( A269  and  (not A268) );
 a46478a <=( (not A302)  and  (not A300) );
 a46479a <=( a46478a  and  a46475a );
 a46480a <=( a46479a  and  a46472a );
 a46484a <=( (not A167)  and  A168 );
 a46485a <=( A170  and  a46484a );
 a46489a <=( A200  and  A199 );
 a46490a <=( A166  and  a46489a );
 a46491a <=( a46490a  and  a46485a );
 a46495a <=( (not A267)  and  (not A266) );
 a46496a <=( A265  and  a46495a );
 a46499a <=( A269  and  (not A268) );
 a46502a <=( A299  and  A298 );
 a46503a <=( a46502a  and  a46499a );
 a46504a <=( a46503a  and  a46496a );
 a46508a <=( (not A167)  and  A168 );
 a46509a <=( A170  and  a46508a );
 a46513a <=( A200  and  A199 );
 a46514a <=( A166  and  a46513a );
 a46515a <=( a46514a  and  a46509a );
 a46519a <=( (not A267)  and  (not A266) );
 a46520a <=( A265  and  a46519a );
 a46523a <=( A269  and  (not A268) );
 a46526a <=( (not A299)  and  (not A298) );
 a46527a <=( a46526a  and  a46523a );
 a46528a <=( a46527a  and  a46520a );
 a46532a <=( (not A167)  and  A168 );
 a46533a <=( A170  and  a46532a );
 a46537a <=( A200  and  A199 );
 a46538a <=( A166  and  a46537a );
 a46539a <=( a46538a  and  a46533a );
 a46543a <=( A298  and  (not A266) );
 a46544a <=( (not A265)  and  a46543a );
 a46547a <=( (not A300)  and  (not A299) );
 a46550a <=( A302  and  (not A301) );
 a46551a <=( a46550a  and  a46547a );
 a46552a <=( a46551a  and  a46544a );
 a46556a <=( (not A167)  and  A168 );
 a46557a <=( A170  and  a46556a );
 a46561a <=( A200  and  A199 );
 a46562a <=( A166  and  a46561a );
 a46563a <=( a46562a  and  a46557a );
 a46567a <=( (not A298)  and  (not A266) );
 a46568a <=( (not A265)  and  a46567a );
 a46571a <=( (not A300)  and  A299 );
 a46574a <=( A302  and  (not A301) );
 a46575a <=( a46574a  and  a46571a );
 a46576a <=( a46575a  and  a46568a );
 a46580a <=( (not A167)  and  A168 );
 a46581a <=( A170  and  a46580a );
 a46585a <=( (not A200)  and  (not A199) );
 a46586a <=( A166  and  a46585a );
 a46587a <=( a46586a  and  a46581a );
 a46591a <=( A269  and  (not A268) );
 a46592a <=( A267  and  a46591a );
 a46595a <=( (not A299)  and  A298 );
 a46598a <=( A301  and  A300 );
 a46599a <=( a46598a  and  a46595a );
 a46600a <=( a46599a  and  a46592a );
 a46604a <=( (not A167)  and  A168 );
 a46605a <=( A170  and  a46604a );
 a46609a <=( (not A200)  and  (not A199) );
 a46610a <=( A166  and  a46609a );
 a46611a <=( a46610a  and  a46605a );
 a46615a <=( A269  and  (not A268) );
 a46616a <=( A267  and  a46615a );
 a46619a <=( (not A299)  and  A298 );
 a46622a <=( (not A302)  and  A300 );
 a46623a <=( a46622a  and  a46619a );
 a46624a <=( a46623a  and  a46616a );
 a46628a <=( (not A167)  and  A168 );
 a46629a <=( A170  and  a46628a );
 a46633a <=( (not A200)  and  (not A199) );
 a46634a <=( A166  and  a46633a );
 a46635a <=( a46634a  and  a46629a );
 a46639a <=( A269  and  (not A268) );
 a46640a <=( A267  and  a46639a );
 a46643a <=( A299  and  (not A298) );
 a46646a <=( A301  and  A300 );
 a46647a <=( a46646a  and  a46643a );
 a46648a <=( a46647a  and  a46640a );
 a46652a <=( (not A167)  and  A168 );
 a46653a <=( A170  and  a46652a );
 a46657a <=( (not A200)  and  (not A199) );
 a46658a <=( A166  and  a46657a );
 a46659a <=( a46658a  and  a46653a );
 a46663a <=( A269  and  (not A268) );
 a46664a <=( A267  and  a46663a );
 a46667a <=( A299  and  (not A298) );
 a46670a <=( (not A302)  and  A300 );
 a46671a <=( a46670a  and  a46667a );
 a46672a <=( a46671a  and  a46664a );
 a46676a <=( (not A167)  and  A168 );
 a46677a <=( A170  and  a46676a );
 a46681a <=( (not A200)  and  (not A199) );
 a46682a <=( A166  and  a46681a );
 a46683a <=( a46682a  and  a46677a );
 a46687a <=( A298  and  A268 );
 a46688a <=( (not A267)  and  a46687a );
 a46691a <=( (not A300)  and  (not A299) );
 a46694a <=( A302  and  (not A301) );
 a46695a <=( a46694a  and  a46691a );
 a46696a <=( a46695a  and  a46688a );
 a46700a <=( (not A167)  and  A168 );
 a46701a <=( A170  and  a46700a );
 a46705a <=( (not A200)  and  (not A199) );
 a46706a <=( A166  and  a46705a );
 a46707a <=( a46706a  and  a46701a );
 a46711a <=( (not A298)  and  A268 );
 a46712a <=( (not A267)  and  a46711a );
 a46715a <=( (not A300)  and  A299 );
 a46718a <=( A302  and  (not A301) );
 a46719a <=( a46718a  and  a46715a );
 a46720a <=( a46719a  and  a46712a );
 a46724a <=( (not A167)  and  A168 );
 a46725a <=( A170  and  a46724a );
 a46729a <=( (not A200)  and  (not A199) );
 a46730a <=( A166  and  a46729a );
 a46731a <=( a46730a  and  a46725a );
 a46735a <=( A298  and  (not A269) );
 a46736a <=( (not A267)  and  a46735a );
 a46739a <=( (not A300)  and  (not A299) );
 a46742a <=( A302  and  (not A301) );
 a46743a <=( a46742a  and  a46739a );
 a46744a <=( a46743a  and  a46736a );
 a46748a <=( (not A167)  and  A168 );
 a46749a <=( A170  and  a46748a );
 a46753a <=( (not A200)  and  (not A199) );
 a46754a <=( A166  and  a46753a );
 a46755a <=( a46754a  and  a46749a );
 a46759a <=( (not A298)  and  (not A269) );
 a46760a <=( (not A267)  and  a46759a );
 a46763a <=( (not A300)  and  A299 );
 a46766a <=( A302  and  (not A301) );
 a46767a <=( a46766a  and  a46763a );
 a46768a <=( a46767a  and  a46760a );
 a46772a <=( (not A167)  and  A168 );
 a46773a <=( A170  and  a46772a );
 a46777a <=( (not A200)  and  (not A199) );
 a46778a <=( A166  and  a46777a );
 a46779a <=( a46778a  and  a46773a );
 a46783a <=( A298  and  A266 );
 a46784a <=( A265  and  a46783a );
 a46787a <=( (not A300)  and  (not A299) );
 a46790a <=( A302  and  (not A301) );
 a46791a <=( a46790a  and  a46787a );
 a46792a <=( a46791a  and  a46784a );
 a46796a <=( (not A167)  and  A168 );
 a46797a <=( A170  and  a46796a );
 a46801a <=( (not A200)  and  (not A199) );
 a46802a <=( A166  and  a46801a );
 a46803a <=( a46802a  and  a46797a );
 a46807a <=( (not A298)  and  A266 );
 a46808a <=( A265  and  a46807a );
 a46811a <=( (not A300)  and  A299 );
 a46814a <=( A302  and  (not A301) );
 a46815a <=( a46814a  and  a46811a );
 a46816a <=( a46815a  and  a46808a );
 a46820a <=( (not A167)  and  A168 );
 a46821a <=( A170  and  a46820a );
 a46825a <=( (not A200)  and  (not A199) );
 a46826a <=( A166  and  a46825a );
 a46827a <=( a46826a  and  a46821a );
 a46831a <=( A267  and  A266 );
 a46832a <=( (not A265)  and  a46831a );
 a46835a <=( A300  and  A268 );
 a46838a <=( A302  and  (not A301) );
 a46839a <=( a46838a  and  a46835a );
 a46840a <=( a46839a  and  a46832a );
 a46844a <=( (not A167)  and  A168 );
 a46845a <=( A170  and  a46844a );
 a46849a <=( (not A200)  and  (not A199) );
 a46850a <=( A166  and  a46849a );
 a46851a <=( a46850a  and  a46845a );
 a46855a <=( A267  and  A266 );
 a46856a <=( (not A265)  and  a46855a );
 a46859a <=( A300  and  (not A269) );
 a46862a <=( A302  and  (not A301) );
 a46863a <=( a46862a  and  a46859a );
 a46864a <=( a46863a  and  a46856a );
 a46868a <=( (not A167)  and  A168 );
 a46869a <=( A170  and  a46868a );
 a46873a <=( (not A200)  and  (not A199) );
 a46874a <=( A166  and  a46873a );
 a46875a <=( a46874a  and  a46869a );
 a46879a <=( (not A267)  and  A266 );
 a46880a <=( (not A265)  and  a46879a );
 a46883a <=( A269  and  (not A268) );
 a46886a <=( A301  and  (not A300) );
 a46887a <=( a46886a  and  a46883a );
 a46888a <=( a46887a  and  a46880a );
 a46892a <=( (not A167)  and  A168 );
 a46893a <=( A170  and  a46892a );
 a46897a <=( (not A200)  and  (not A199) );
 a46898a <=( A166  and  a46897a );
 a46899a <=( a46898a  and  a46893a );
 a46903a <=( (not A267)  and  A266 );
 a46904a <=( (not A265)  and  a46903a );
 a46907a <=( A269  and  (not A268) );
 a46910a <=( (not A302)  and  (not A300) );
 a46911a <=( a46910a  and  a46907a );
 a46912a <=( a46911a  and  a46904a );
 a46916a <=( (not A167)  and  A168 );
 a46917a <=( A170  and  a46916a );
 a46921a <=( (not A200)  and  (not A199) );
 a46922a <=( A166  and  a46921a );
 a46923a <=( a46922a  and  a46917a );
 a46927a <=( (not A267)  and  A266 );
 a46928a <=( (not A265)  and  a46927a );
 a46931a <=( A269  and  (not A268) );
 a46934a <=( A299  and  A298 );
 a46935a <=( a46934a  and  a46931a );
 a46936a <=( a46935a  and  a46928a );
 a46940a <=( (not A167)  and  A168 );
 a46941a <=( A170  and  a46940a );
 a46945a <=( (not A200)  and  (not A199) );
 a46946a <=( A166  and  a46945a );
 a46947a <=( a46946a  and  a46941a );
 a46951a <=( (not A267)  and  A266 );
 a46952a <=( (not A265)  and  a46951a );
 a46955a <=( A269  and  (not A268) );
 a46958a <=( (not A299)  and  (not A298) );
 a46959a <=( a46958a  and  a46955a );
 a46960a <=( a46959a  and  a46952a );
 a46964a <=( (not A167)  and  A168 );
 a46965a <=( A170  and  a46964a );
 a46969a <=( (not A200)  and  (not A199) );
 a46970a <=( A166  and  a46969a );
 a46971a <=( a46970a  and  a46965a );
 a46975a <=( A267  and  (not A266) );
 a46976a <=( A265  and  a46975a );
 a46979a <=( A300  and  A268 );
 a46982a <=( A302  and  (not A301) );
 a46983a <=( a46982a  and  a46979a );
 a46984a <=( a46983a  and  a46976a );
 a46988a <=( (not A167)  and  A168 );
 a46989a <=( A170  and  a46988a );
 a46993a <=( (not A200)  and  (not A199) );
 a46994a <=( A166  and  a46993a );
 a46995a <=( a46994a  and  a46989a );
 a46999a <=( A267  and  (not A266) );
 a47000a <=( A265  and  a46999a );
 a47003a <=( A300  and  (not A269) );
 a47006a <=( A302  and  (not A301) );
 a47007a <=( a47006a  and  a47003a );
 a47008a <=( a47007a  and  a47000a );
 a47012a <=( (not A167)  and  A168 );
 a47013a <=( A170  and  a47012a );
 a47017a <=( (not A200)  and  (not A199) );
 a47018a <=( A166  and  a47017a );
 a47019a <=( a47018a  and  a47013a );
 a47023a <=( (not A267)  and  (not A266) );
 a47024a <=( A265  and  a47023a );
 a47027a <=( A269  and  (not A268) );
 a47030a <=( A301  and  (not A300) );
 a47031a <=( a47030a  and  a47027a );
 a47032a <=( a47031a  and  a47024a );
 a47036a <=( (not A167)  and  A168 );
 a47037a <=( A170  and  a47036a );
 a47041a <=( (not A200)  and  (not A199) );
 a47042a <=( A166  and  a47041a );
 a47043a <=( a47042a  and  a47037a );
 a47047a <=( (not A267)  and  (not A266) );
 a47048a <=( A265  and  a47047a );
 a47051a <=( A269  and  (not A268) );
 a47054a <=( (not A302)  and  (not A300) );
 a47055a <=( a47054a  and  a47051a );
 a47056a <=( a47055a  and  a47048a );
 a47060a <=( (not A167)  and  A168 );
 a47061a <=( A170  and  a47060a );
 a47065a <=( (not A200)  and  (not A199) );
 a47066a <=( A166  and  a47065a );
 a47067a <=( a47066a  and  a47061a );
 a47071a <=( (not A267)  and  (not A266) );
 a47072a <=( A265  and  a47071a );
 a47075a <=( A269  and  (not A268) );
 a47078a <=( A299  and  A298 );
 a47079a <=( a47078a  and  a47075a );
 a47080a <=( a47079a  and  a47072a );
 a47084a <=( (not A167)  and  A168 );
 a47085a <=( A170  and  a47084a );
 a47089a <=( (not A200)  and  (not A199) );
 a47090a <=( A166  and  a47089a );
 a47091a <=( a47090a  and  a47085a );
 a47095a <=( (not A267)  and  (not A266) );
 a47096a <=( A265  and  a47095a );
 a47099a <=( A269  and  (not A268) );
 a47102a <=( (not A299)  and  (not A298) );
 a47103a <=( a47102a  and  a47099a );
 a47104a <=( a47103a  and  a47096a );
 a47108a <=( (not A167)  and  A168 );
 a47109a <=( A170  and  a47108a );
 a47113a <=( (not A200)  and  (not A199) );
 a47114a <=( A166  and  a47113a );
 a47115a <=( a47114a  and  a47109a );
 a47119a <=( A298  and  (not A266) );
 a47120a <=( (not A265)  and  a47119a );
 a47123a <=( (not A300)  and  (not A299) );
 a47126a <=( A302  and  (not A301) );
 a47127a <=( a47126a  and  a47123a );
 a47128a <=( a47127a  and  a47120a );
 a47132a <=( (not A167)  and  A168 );
 a47133a <=( A170  and  a47132a );
 a47137a <=( (not A200)  and  (not A199) );
 a47138a <=( A166  and  a47137a );
 a47139a <=( a47138a  and  a47133a );
 a47143a <=( (not A298)  and  (not A266) );
 a47144a <=( (not A265)  and  a47143a );
 a47147a <=( (not A300)  and  A299 );
 a47150a <=( A302  and  (not A301) );
 a47151a <=( a47150a  and  a47147a );
 a47152a <=( a47151a  and  a47144a );
 a47156a <=( (not A199)  and  (not A168) );
 a47157a <=( A170  and  a47156a );
 a47161a <=( (not A202)  and  (not A201) );
 a47162a <=( A200  and  a47161a );
 a47163a <=( a47162a  and  a47157a );
 a47167a <=( (not A268)  and  A267 );
 a47168a <=( A203  and  a47167a );
 a47171a <=( A300  and  A269 );
 a47174a <=( A302  and  (not A301) );
 a47175a <=( a47174a  and  a47171a );
 a47176a <=( a47175a  and  a47168a );
 a47180a <=( A199  and  (not A168) );
 a47181a <=( A170  and  a47180a );
 a47185a <=( (not A202)  and  (not A201) );
 a47186a <=( (not A200)  and  a47185a );
 a47187a <=( a47186a  and  a47181a );
 a47191a <=( (not A268)  and  A267 );
 a47192a <=( A203  and  a47191a );
 a47195a <=( A300  and  A269 );
 a47198a <=( A302  and  (not A301) );
 a47199a <=( a47198a  and  a47195a );
 a47200a <=( a47199a  and  a47192a );
 a47204a <=( A167  and  A168 );
 a47205a <=( A169  and  a47204a );
 a47209a <=( (not A202)  and  A201 );
 a47210a <=( (not A166)  and  a47209a );
 a47211a <=( a47210a  and  a47205a );
 a47215a <=( A268  and  (not A267) );
 a47216a <=( A203  and  a47215a );
 a47219a <=( (not A299)  and  A298 );
 a47222a <=( A301  and  A300 );
 a47223a <=( a47222a  and  a47219a );
 a47224a <=( a47223a  and  a47216a );
 a47228a <=( A167  and  A168 );
 a47229a <=( A169  and  a47228a );
 a47233a <=( (not A202)  and  A201 );
 a47234a <=( (not A166)  and  a47233a );
 a47235a <=( a47234a  and  a47229a );
 a47239a <=( A268  and  (not A267) );
 a47240a <=( A203  and  a47239a );
 a47243a <=( (not A299)  and  A298 );
 a47246a <=( (not A302)  and  A300 );
 a47247a <=( a47246a  and  a47243a );
 a47248a <=( a47247a  and  a47240a );
 a47252a <=( A167  and  A168 );
 a47253a <=( A169  and  a47252a );
 a47257a <=( (not A202)  and  A201 );
 a47258a <=( (not A166)  and  a47257a );
 a47259a <=( a47258a  and  a47253a );
 a47263a <=( A268  and  (not A267) );
 a47264a <=( A203  and  a47263a );
 a47267a <=( A299  and  (not A298) );
 a47270a <=( A301  and  A300 );
 a47271a <=( a47270a  and  a47267a );
 a47272a <=( a47271a  and  a47264a );
 a47276a <=( A167  and  A168 );
 a47277a <=( A169  and  a47276a );
 a47281a <=( (not A202)  and  A201 );
 a47282a <=( (not A166)  and  a47281a );
 a47283a <=( a47282a  and  a47277a );
 a47287a <=( A268  and  (not A267) );
 a47288a <=( A203  and  a47287a );
 a47291a <=( A299  and  (not A298) );
 a47294a <=( (not A302)  and  A300 );
 a47295a <=( a47294a  and  a47291a );
 a47296a <=( a47295a  and  a47288a );
 a47300a <=( A167  and  A168 );
 a47301a <=( A169  and  a47300a );
 a47305a <=( (not A202)  and  A201 );
 a47306a <=( (not A166)  and  a47305a );
 a47307a <=( a47306a  and  a47301a );
 a47311a <=( (not A269)  and  (not A267) );
 a47312a <=( A203  and  a47311a );
 a47315a <=( (not A299)  and  A298 );
 a47318a <=( A301  and  A300 );
 a47319a <=( a47318a  and  a47315a );
 a47320a <=( a47319a  and  a47312a );
 a47324a <=( A167  and  A168 );
 a47325a <=( A169  and  a47324a );
 a47329a <=( (not A202)  and  A201 );
 a47330a <=( (not A166)  and  a47329a );
 a47331a <=( a47330a  and  a47325a );
 a47335a <=( (not A269)  and  (not A267) );
 a47336a <=( A203  and  a47335a );
 a47339a <=( (not A299)  and  A298 );
 a47342a <=( (not A302)  and  A300 );
 a47343a <=( a47342a  and  a47339a );
 a47344a <=( a47343a  and  a47336a );
 a47348a <=( A167  and  A168 );
 a47349a <=( A169  and  a47348a );
 a47353a <=( (not A202)  and  A201 );
 a47354a <=( (not A166)  and  a47353a );
 a47355a <=( a47354a  and  a47349a );
 a47359a <=( (not A269)  and  (not A267) );
 a47360a <=( A203  and  a47359a );
 a47363a <=( A299  and  (not A298) );
 a47366a <=( A301  and  A300 );
 a47367a <=( a47366a  and  a47363a );
 a47368a <=( a47367a  and  a47360a );
 a47372a <=( A167  and  A168 );
 a47373a <=( A169  and  a47372a );
 a47377a <=( (not A202)  and  A201 );
 a47378a <=( (not A166)  and  a47377a );
 a47379a <=( a47378a  and  a47373a );
 a47383a <=( (not A269)  and  (not A267) );
 a47384a <=( A203  and  a47383a );
 a47387a <=( A299  and  (not A298) );
 a47390a <=( (not A302)  and  A300 );
 a47391a <=( a47390a  and  a47387a );
 a47392a <=( a47391a  and  a47384a );
 a47396a <=( A167  and  A168 );
 a47397a <=( A169  and  a47396a );
 a47401a <=( (not A202)  and  A201 );
 a47402a <=( (not A166)  and  a47401a );
 a47403a <=( a47402a  and  a47397a );
 a47407a <=( A266  and  A265 );
 a47408a <=( A203  and  a47407a );
 a47411a <=( (not A299)  and  A298 );
 a47414a <=( A301  and  A300 );
 a47415a <=( a47414a  and  a47411a );
 a47416a <=( a47415a  and  a47408a );
 a47420a <=( A167  and  A168 );
 a47421a <=( A169  and  a47420a );
 a47425a <=( (not A202)  and  A201 );
 a47426a <=( (not A166)  and  a47425a );
 a47427a <=( a47426a  and  a47421a );
 a47431a <=( A266  and  A265 );
 a47432a <=( A203  and  a47431a );
 a47435a <=( (not A299)  and  A298 );
 a47438a <=( (not A302)  and  A300 );
 a47439a <=( a47438a  and  a47435a );
 a47440a <=( a47439a  and  a47432a );
 a47444a <=( A167  and  A168 );
 a47445a <=( A169  and  a47444a );
 a47449a <=( (not A202)  and  A201 );
 a47450a <=( (not A166)  and  a47449a );
 a47451a <=( a47450a  and  a47445a );
 a47455a <=( A266  and  A265 );
 a47456a <=( A203  and  a47455a );
 a47459a <=( A299  and  (not A298) );
 a47462a <=( A301  and  A300 );
 a47463a <=( a47462a  and  a47459a );
 a47464a <=( a47463a  and  a47456a );
 a47468a <=( A167  and  A168 );
 a47469a <=( A169  and  a47468a );
 a47473a <=( (not A202)  and  A201 );
 a47474a <=( (not A166)  and  a47473a );
 a47475a <=( a47474a  and  a47469a );
 a47479a <=( A266  and  A265 );
 a47480a <=( A203  and  a47479a );
 a47483a <=( A299  and  (not A298) );
 a47486a <=( (not A302)  and  A300 );
 a47487a <=( a47486a  and  a47483a );
 a47488a <=( a47487a  and  a47480a );
 a47492a <=( A167  and  A168 );
 a47493a <=( A169  and  a47492a );
 a47497a <=( (not A202)  and  A201 );
 a47498a <=( (not A166)  and  a47497a );
 a47499a <=( a47498a  and  a47493a );
 a47503a <=( A266  and  (not A265) );
 a47504a <=( A203  and  a47503a );
 a47507a <=( A268  and  A267 );
 a47510a <=( A301  and  (not A300) );
 a47511a <=( a47510a  and  a47507a );
 a47512a <=( a47511a  and  a47504a );
 a47516a <=( A167  and  A168 );
 a47517a <=( A169  and  a47516a );
 a47521a <=( (not A202)  and  A201 );
 a47522a <=( (not A166)  and  a47521a );
 a47523a <=( a47522a  and  a47517a );
 a47527a <=( A266  and  (not A265) );
 a47528a <=( A203  and  a47527a );
 a47531a <=( A268  and  A267 );
 a47534a <=( (not A302)  and  (not A300) );
 a47535a <=( a47534a  and  a47531a );
 a47536a <=( a47535a  and  a47528a );
 a47540a <=( A167  and  A168 );
 a47541a <=( A169  and  a47540a );
 a47545a <=( (not A202)  and  A201 );
 a47546a <=( (not A166)  and  a47545a );
 a47547a <=( a47546a  and  a47541a );
 a47551a <=( A266  and  (not A265) );
 a47552a <=( A203  and  a47551a );
 a47555a <=( A268  and  A267 );
 a47558a <=( A299  and  A298 );
 a47559a <=( a47558a  and  a47555a );
 a47560a <=( a47559a  and  a47552a );
 a47564a <=( A167  and  A168 );
 a47565a <=( A169  and  a47564a );
 a47569a <=( (not A202)  and  A201 );
 a47570a <=( (not A166)  and  a47569a );
 a47571a <=( a47570a  and  a47565a );
 a47575a <=( A266  and  (not A265) );
 a47576a <=( A203  and  a47575a );
 a47579a <=( A268  and  A267 );
 a47582a <=( (not A299)  and  (not A298) );
 a47583a <=( a47582a  and  a47579a );
 a47584a <=( a47583a  and  a47576a );
 a47588a <=( A167  and  A168 );
 a47589a <=( A169  and  a47588a );
 a47593a <=( (not A202)  and  A201 );
 a47594a <=( (not A166)  and  a47593a );
 a47595a <=( a47594a  and  a47589a );
 a47599a <=( A266  and  (not A265) );
 a47600a <=( A203  and  a47599a );
 a47603a <=( (not A269)  and  A267 );
 a47606a <=( A301  and  (not A300) );
 a47607a <=( a47606a  and  a47603a );
 a47608a <=( a47607a  and  a47600a );
 a47612a <=( A167  and  A168 );
 a47613a <=( A169  and  a47612a );
 a47617a <=( (not A202)  and  A201 );
 a47618a <=( (not A166)  and  a47617a );
 a47619a <=( a47618a  and  a47613a );
 a47623a <=( A266  and  (not A265) );
 a47624a <=( A203  and  a47623a );
 a47627a <=( (not A269)  and  A267 );
 a47630a <=( (not A302)  and  (not A300) );
 a47631a <=( a47630a  and  a47627a );
 a47632a <=( a47631a  and  a47624a );
 a47636a <=( A167  and  A168 );
 a47637a <=( A169  and  a47636a );
 a47641a <=( (not A202)  and  A201 );
 a47642a <=( (not A166)  and  a47641a );
 a47643a <=( a47642a  and  a47637a );
 a47647a <=( A266  and  (not A265) );
 a47648a <=( A203  and  a47647a );
 a47651a <=( (not A269)  and  A267 );
 a47654a <=( A299  and  A298 );
 a47655a <=( a47654a  and  a47651a );
 a47656a <=( a47655a  and  a47648a );
 a47660a <=( A167  and  A168 );
 a47661a <=( A169  and  a47660a );
 a47665a <=( (not A202)  and  A201 );
 a47666a <=( (not A166)  and  a47665a );
 a47667a <=( a47666a  and  a47661a );
 a47671a <=( A266  and  (not A265) );
 a47672a <=( A203  and  a47671a );
 a47675a <=( (not A269)  and  A267 );
 a47678a <=( (not A299)  and  (not A298) );
 a47679a <=( a47678a  and  a47675a );
 a47680a <=( a47679a  and  a47672a );
 a47684a <=( A167  and  A168 );
 a47685a <=( A169  and  a47684a );
 a47689a <=( (not A202)  and  A201 );
 a47690a <=( (not A166)  and  a47689a );
 a47691a <=( a47690a  and  a47685a );
 a47695a <=( (not A266)  and  A265 );
 a47696a <=( A203  and  a47695a );
 a47699a <=( A268  and  A267 );
 a47702a <=( A301  and  (not A300) );
 a47703a <=( a47702a  and  a47699a );
 a47704a <=( a47703a  and  a47696a );
 a47708a <=( A167  and  A168 );
 a47709a <=( A169  and  a47708a );
 a47713a <=( (not A202)  and  A201 );
 a47714a <=( (not A166)  and  a47713a );
 a47715a <=( a47714a  and  a47709a );
 a47719a <=( (not A266)  and  A265 );
 a47720a <=( A203  and  a47719a );
 a47723a <=( A268  and  A267 );
 a47726a <=( (not A302)  and  (not A300) );
 a47727a <=( a47726a  and  a47723a );
 a47728a <=( a47727a  and  a47720a );
 a47732a <=( A167  and  A168 );
 a47733a <=( A169  and  a47732a );
 a47737a <=( (not A202)  and  A201 );
 a47738a <=( (not A166)  and  a47737a );
 a47739a <=( a47738a  and  a47733a );
 a47743a <=( (not A266)  and  A265 );
 a47744a <=( A203  and  a47743a );
 a47747a <=( A268  and  A267 );
 a47750a <=( A299  and  A298 );
 a47751a <=( a47750a  and  a47747a );
 a47752a <=( a47751a  and  a47744a );
 a47756a <=( A167  and  A168 );
 a47757a <=( A169  and  a47756a );
 a47761a <=( (not A202)  and  A201 );
 a47762a <=( (not A166)  and  a47761a );
 a47763a <=( a47762a  and  a47757a );
 a47767a <=( (not A266)  and  A265 );
 a47768a <=( A203  and  a47767a );
 a47771a <=( A268  and  A267 );
 a47774a <=( (not A299)  and  (not A298) );
 a47775a <=( a47774a  and  a47771a );
 a47776a <=( a47775a  and  a47768a );
 a47780a <=( A167  and  A168 );
 a47781a <=( A169  and  a47780a );
 a47785a <=( (not A202)  and  A201 );
 a47786a <=( (not A166)  and  a47785a );
 a47787a <=( a47786a  and  a47781a );
 a47791a <=( (not A266)  and  A265 );
 a47792a <=( A203  and  a47791a );
 a47795a <=( (not A269)  and  A267 );
 a47798a <=( A301  and  (not A300) );
 a47799a <=( a47798a  and  a47795a );
 a47800a <=( a47799a  and  a47792a );
 a47804a <=( A167  and  A168 );
 a47805a <=( A169  and  a47804a );
 a47809a <=( (not A202)  and  A201 );
 a47810a <=( (not A166)  and  a47809a );
 a47811a <=( a47810a  and  a47805a );
 a47815a <=( (not A266)  and  A265 );
 a47816a <=( A203  and  a47815a );
 a47819a <=( (not A269)  and  A267 );
 a47822a <=( (not A302)  and  (not A300) );
 a47823a <=( a47822a  and  a47819a );
 a47824a <=( a47823a  and  a47816a );
 a47828a <=( A167  and  A168 );
 a47829a <=( A169  and  a47828a );
 a47833a <=( (not A202)  and  A201 );
 a47834a <=( (not A166)  and  a47833a );
 a47835a <=( a47834a  and  a47829a );
 a47839a <=( (not A266)  and  A265 );
 a47840a <=( A203  and  a47839a );
 a47843a <=( (not A269)  and  A267 );
 a47846a <=( A299  and  A298 );
 a47847a <=( a47846a  and  a47843a );
 a47848a <=( a47847a  and  a47840a );
 a47852a <=( A167  and  A168 );
 a47853a <=( A169  and  a47852a );
 a47857a <=( (not A202)  and  A201 );
 a47858a <=( (not A166)  and  a47857a );
 a47859a <=( a47858a  and  a47853a );
 a47863a <=( (not A266)  and  A265 );
 a47864a <=( A203  and  a47863a );
 a47867a <=( (not A269)  and  A267 );
 a47870a <=( (not A299)  and  (not A298) );
 a47871a <=( a47870a  and  a47867a );
 a47872a <=( a47871a  and  a47864a );
 a47876a <=( A167  and  A168 );
 a47877a <=( A169  and  a47876a );
 a47881a <=( (not A202)  and  A201 );
 a47882a <=( (not A166)  and  a47881a );
 a47883a <=( a47882a  and  a47877a );
 a47887a <=( (not A266)  and  (not A265) );
 a47888a <=( A203  and  a47887a );
 a47891a <=( (not A299)  and  A298 );
 a47894a <=( A301  and  A300 );
 a47895a <=( a47894a  and  a47891a );
 a47896a <=( a47895a  and  a47888a );
 a47900a <=( A167  and  A168 );
 a47901a <=( A169  and  a47900a );
 a47905a <=( (not A202)  and  A201 );
 a47906a <=( (not A166)  and  a47905a );
 a47907a <=( a47906a  and  a47901a );
 a47911a <=( (not A266)  and  (not A265) );
 a47912a <=( A203  and  a47911a );
 a47915a <=( (not A299)  and  A298 );
 a47918a <=( (not A302)  and  A300 );
 a47919a <=( a47918a  and  a47915a );
 a47920a <=( a47919a  and  a47912a );
 a47924a <=( A167  and  A168 );
 a47925a <=( A169  and  a47924a );
 a47929a <=( (not A202)  and  A201 );
 a47930a <=( (not A166)  and  a47929a );
 a47931a <=( a47930a  and  a47925a );
 a47935a <=( (not A266)  and  (not A265) );
 a47936a <=( A203  and  a47935a );
 a47939a <=( A299  and  (not A298) );
 a47942a <=( A301  and  A300 );
 a47943a <=( a47942a  and  a47939a );
 a47944a <=( a47943a  and  a47936a );
 a47948a <=( A167  and  A168 );
 a47949a <=( A169  and  a47948a );
 a47953a <=( (not A202)  and  A201 );
 a47954a <=( (not A166)  and  a47953a );
 a47955a <=( a47954a  and  a47949a );
 a47959a <=( (not A266)  and  (not A265) );
 a47960a <=( A203  and  a47959a );
 a47963a <=( A299  and  (not A298) );
 a47966a <=( (not A302)  and  A300 );
 a47967a <=( a47966a  and  a47963a );
 a47968a <=( a47967a  and  a47960a );
 a47972a <=( A167  and  A168 );
 a47973a <=( A169  and  a47972a );
 a47977a <=( A202  and  (not A201) );
 a47978a <=( (not A166)  and  a47977a );
 a47979a <=( a47978a  and  a47973a );
 a47983a <=( A269  and  (not A268) );
 a47984a <=( A267  and  a47983a );
 a47987a <=( (not A299)  and  A298 );
 a47990a <=( A301  and  A300 );
 a47991a <=( a47990a  and  a47987a );
 a47992a <=( a47991a  and  a47984a );
 a47996a <=( A167  and  A168 );
 a47997a <=( A169  and  a47996a );
 a48001a <=( A202  and  (not A201) );
 a48002a <=( (not A166)  and  a48001a );
 a48003a <=( a48002a  and  a47997a );
 a48007a <=( A269  and  (not A268) );
 a48008a <=( A267  and  a48007a );
 a48011a <=( (not A299)  and  A298 );
 a48014a <=( (not A302)  and  A300 );
 a48015a <=( a48014a  and  a48011a );
 a48016a <=( a48015a  and  a48008a );
 a48020a <=( A167  and  A168 );
 a48021a <=( A169  and  a48020a );
 a48025a <=( A202  and  (not A201) );
 a48026a <=( (not A166)  and  a48025a );
 a48027a <=( a48026a  and  a48021a );
 a48031a <=( A269  and  (not A268) );
 a48032a <=( A267  and  a48031a );
 a48035a <=( A299  and  (not A298) );
 a48038a <=( A301  and  A300 );
 a48039a <=( a48038a  and  a48035a );
 a48040a <=( a48039a  and  a48032a );
 a48044a <=( A167  and  A168 );
 a48045a <=( A169  and  a48044a );
 a48049a <=( A202  and  (not A201) );
 a48050a <=( (not A166)  and  a48049a );
 a48051a <=( a48050a  and  a48045a );
 a48055a <=( A269  and  (not A268) );
 a48056a <=( A267  and  a48055a );
 a48059a <=( A299  and  (not A298) );
 a48062a <=( (not A302)  and  A300 );
 a48063a <=( a48062a  and  a48059a );
 a48064a <=( a48063a  and  a48056a );
 a48068a <=( A167  and  A168 );
 a48069a <=( A169  and  a48068a );
 a48073a <=( A202  and  (not A201) );
 a48074a <=( (not A166)  and  a48073a );
 a48075a <=( a48074a  and  a48069a );
 a48079a <=( A298  and  A268 );
 a48080a <=( (not A267)  and  a48079a );
 a48083a <=( (not A300)  and  (not A299) );
 a48086a <=( A302  and  (not A301) );
 a48087a <=( a48086a  and  a48083a );
 a48088a <=( a48087a  and  a48080a );
 a48092a <=( A167  and  A168 );
 a48093a <=( A169  and  a48092a );
 a48097a <=( A202  and  (not A201) );
 a48098a <=( (not A166)  and  a48097a );
 a48099a <=( a48098a  and  a48093a );
 a48103a <=( (not A298)  and  A268 );
 a48104a <=( (not A267)  and  a48103a );
 a48107a <=( (not A300)  and  A299 );
 a48110a <=( A302  and  (not A301) );
 a48111a <=( a48110a  and  a48107a );
 a48112a <=( a48111a  and  a48104a );
 a48116a <=( A167  and  A168 );
 a48117a <=( A169  and  a48116a );
 a48121a <=( A202  and  (not A201) );
 a48122a <=( (not A166)  and  a48121a );
 a48123a <=( a48122a  and  a48117a );
 a48127a <=( A298  and  (not A269) );
 a48128a <=( (not A267)  and  a48127a );
 a48131a <=( (not A300)  and  (not A299) );
 a48134a <=( A302  and  (not A301) );
 a48135a <=( a48134a  and  a48131a );
 a48136a <=( a48135a  and  a48128a );
 a48140a <=( A167  and  A168 );
 a48141a <=( A169  and  a48140a );
 a48145a <=( A202  and  (not A201) );
 a48146a <=( (not A166)  and  a48145a );
 a48147a <=( a48146a  and  a48141a );
 a48151a <=( (not A298)  and  (not A269) );
 a48152a <=( (not A267)  and  a48151a );
 a48155a <=( (not A300)  and  A299 );
 a48158a <=( A302  and  (not A301) );
 a48159a <=( a48158a  and  a48155a );
 a48160a <=( a48159a  and  a48152a );
 a48164a <=( A167  and  A168 );
 a48165a <=( A169  and  a48164a );
 a48169a <=( A202  and  (not A201) );
 a48170a <=( (not A166)  and  a48169a );
 a48171a <=( a48170a  and  a48165a );
 a48175a <=( A298  and  A266 );
 a48176a <=( A265  and  a48175a );
 a48179a <=( (not A300)  and  (not A299) );
 a48182a <=( A302  and  (not A301) );
 a48183a <=( a48182a  and  a48179a );
 a48184a <=( a48183a  and  a48176a );
 a48188a <=( A167  and  A168 );
 a48189a <=( A169  and  a48188a );
 a48193a <=( A202  and  (not A201) );
 a48194a <=( (not A166)  and  a48193a );
 a48195a <=( a48194a  and  a48189a );
 a48199a <=( (not A298)  and  A266 );
 a48200a <=( A265  and  a48199a );
 a48203a <=( (not A300)  and  A299 );
 a48206a <=( A302  and  (not A301) );
 a48207a <=( a48206a  and  a48203a );
 a48208a <=( a48207a  and  a48200a );
 a48212a <=( A167  and  A168 );
 a48213a <=( A169  and  a48212a );
 a48217a <=( A202  and  (not A201) );
 a48218a <=( (not A166)  and  a48217a );
 a48219a <=( a48218a  and  a48213a );
 a48223a <=( A267  and  A266 );
 a48224a <=( (not A265)  and  a48223a );
 a48227a <=( A300  and  A268 );
 a48230a <=( A302  and  (not A301) );
 a48231a <=( a48230a  and  a48227a );
 a48232a <=( a48231a  and  a48224a );
 a48236a <=( A167  and  A168 );
 a48237a <=( A169  and  a48236a );
 a48241a <=( A202  and  (not A201) );
 a48242a <=( (not A166)  and  a48241a );
 a48243a <=( a48242a  and  a48237a );
 a48247a <=( A267  and  A266 );
 a48248a <=( (not A265)  and  a48247a );
 a48251a <=( A300  and  (not A269) );
 a48254a <=( A302  and  (not A301) );
 a48255a <=( a48254a  and  a48251a );
 a48256a <=( a48255a  and  a48248a );
 a48260a <=( A167  and  A168 );
 a48261a <=( A169  and  a48260a );
 a48265a <=( A202  and  (not A201) );
 a48266a <=( (not A166)  and  a48265a );
 a48267a <=( a48266a  and  a48261a );
 a48271a <=( (not A267)  and  A266 );
 a48272a <=( (not A265)  and  a48271a );
 a48275a <=( A269  and  (not A268) );
 a48278a <=( A301  and  (not A300) );
 a48279a <=( a48278a  and  a48275a );
 a48280a <=( a48279a  and  a48272a );
 a48284a <=( A167  and  A168 );
 a48285a <=( A169  and  a48284a );
 a48289a <=( A202  and  (not A201) );
 a48290a <=( (not A166)  and  a48289a );
 a48291a <=( a48290a  and  a48285a );
 a48295a <=( (not A267)  and  A266 );
 a48296a <=( (not A265)  and  a48295a );
 a48299a <=( A269  and  (not A268) );
 a48302a <=( (not A302)  and  (not A300) );
 a48303a <=( a48302a  and  a48299a );
 a48304a <=( a48303a  and  a48296a );
 a48308a <=( A167  and  A168 );
 a48309a <=( A169  and  a48308a );
 a48313a <=( A202  and  (not A201) );
 a48314a <=( (not A166)  and  a48313a );
 a48315a <=( a48314a  and  a48309a );
 a48319a <=( (not A267)  and  A266 );
 a48320a <=( (not A265)  and  a48319a );
 a48323a <=( A269  and  (not A268) );
 a48326a <=( A299  and  A298 );
 a48327a <=( a48326a  and  a48323a );
 a48328a <=( a48327a  and  a48320a );
 a48332a <=( A167  and  A168 );
 a48333a <=( A169  and  a48332a );
 a48337a <=( A202  and  (not A201) );
 a48338a <=( (not A166)  and  a48337a );
 a48339a <=( a48338a  and  a48333a );
 a48343a <=( (not A267)  and  A266 );
 a48344a <=( (not A265)  and  a48343a );
 a48347a <=( A269  and  (not A268) );
 a48350a <=( (not A299)  and  (not A298) );
 a48351a <=( a48350a  and  a48347a );
 a48352a <=( a48351a  and  a48344a );
 a48356a <=( A167  and  A168 );
 a48357a <=( A169  and  a48356a );
 a48361a <=( A202  and  (not A201) );
 a48362a <=( (not A166)  and  a48361a );
 a48363a <=( a48362a  and  a48357a );
 a48367a <=( A267  and  (not A266) );
 a48368a <=( A265  and  a48367a );
 a48371a <=( A300  and  A268 );
 a48374a <=( A302  and  (not A301) );
 a48375a <=( a48374a  and  a48371a );
 a48376a <=( a48375a  and  a48368a );
 a48380a <=( A167  and  A168 );
 a48381a <=( A169  and  a48380a );
 a48385a <=( A202  and  (not A201) );
 a48386a <=( (not A166)  and  a48385a );
 a48387a <=( a48386a  and  a48381a );
 a48391a <=( A267  and  (not A266) );
 a48392a <=( A265  and  a48391a );
 a48395a <=( A300  and  (not A269) );
 a48398a <=( A302  and  (not A301) );
 a48399a <=( a48398a  and  a48395a );
 a48400a <=( a48399a  and  a48392a );
 a48404a <=( A167  and  A168 );
 a48405a <=( A169  and  a48404a );
 a48409a <=( A202  and  (not A201) );
 a48410a <=( (not A166)  and  a48409a );
 a48411a <=( a48410a  and  a48405a );
 a48415a <=( (not A267)  and  (not A266) );
 a48416a <=( A265  and  a48415a );
 a48419a <=( A269  and  (not A268) );
 a48422a <=( A301  and  (not A300) );
 a48423a <=( a48422a  and  a48419a );
 a48424a <=( a48423a  and  a48416a );
 a48428a <=( A167  and  A168 );
 a48429a <=( A169  and  a48428a );
 a48433a <=( A202  and  (not A201) );
 a48434a <=( (not A166)  and  a48433a );
 a48435a <=( a48434a  and  a48429a );
 a48439a <=( (not A267)  and  (not A266) );
 a48440a <=( A265  and  a48439a );
 a48443a <=( A269  and  (not A268) );
 a48446a <=( (not A302)  and  (not A300) );
 a48447a <=( a48446a  and  a48443a );
 a48448a <=( a48447a  and  a48440a );
 a48452a <=( A167  and  A168 );
 a48453a <=( A169  and  a48452a );
 a48457a <=( A202  and  (not A201) );
 a48458a <=( (not A166)  and  a48457a );
 a48459a <=( a48458a  and  a48453a );
 a48463a <=( (not A267)  and  (not A266) );
 a48464a <=( A265  and  a48463a );
 a48467a <=( A269  and  (not A268) );
 a48470a <=( A299  and  A298 );
 a48471a <=( a48470a  and  a48467a );
 a48472a <=( a48471a  and  a48464a );
 a48476a <=( A167  and  A168 );
 a48477a <=( A169  and  a48476a );
 a48481a <=( A202  and  (not A201) );
 a48482a <=( (not A166)  and  a48481a );
 a48483a <=( a48482a  and  a48477a );
 a48487a <=( (not A267)  and  (not A266) );
 a48488a <=( A265  and  a48487a );
 a48491a <=( A269  and  (not A268) );
 a48494a <=( (not A299)  and  (not A298) );
 a48495a <=( a48494a  and  a48491a );
 a48496a <=( a48495a  and  a48488a );
 a48500a <=( A167  and  A168 );
 a48501a <=( A169  and  a48500a );
 a48505a <=( A202  and  (not A201) );
 a48506a <=( (not A166)  and  a48505a );
 a48507a <=( a48506a  and  a48501a );
 a48511a <=( A298  and  (not A266) );
 a48512a <=( (not A265)  and  a48511a );
 a48515a <=( (not A300)  and  (not A299) );
 a48518a <=( A302  and  (not A301) );
 a48519a <=( a48518a  and  a48515a );
 a48520a <=( a48519a  and  a48512a );
 a48524a <=( A167  and  A168 );
 a48525a <=( A169  and  a48524a );
 a48529a <=( A202  and  (not A201) );
 a48530a <=( (not A166)  and  a48529a );
 a48531a <=( a48530a  and  a48525a );
 a48535a <=( (not A298)  and  (not A266) );
 a48536a <=( (not A265)  and  a48535a );
 a48539a <=( (not A300)  and  A299 );
 a48542a <=( A302  and  (not A301) );
 a48543a <=( a48542a  and  a48539a );
 a48544a <=( a48543a  and  a48536a );
 a48548a <=( A167  and  A168 );
 a48549a <=( A169  and  a48548a );
 a48553a <=( (not A203)  and  (not A201) );
 a48554a <=( (not A166)  and  a48553a );
 a48555a <=( a48554a  and  a48549a );
 a48559a <=( A269  and  (not A268) );
 a48560a <=( A267  and  a48559a );
 a48563a <=( (not A299)  and  A298 );
 a48566a <=( A301  and  A300 );
 a48567a <=( a48566a  and  a48563a );
 a48568a <=( a48567a  and  a48560a );
 a48572a <=( A167  and  A168 );
 a48573a <=( A169  and  a48572a );
 a48577a <=( (not A203)  and  (not A201) );
 a48578a <=( (not A166)  and  a48577a );
 a48579a <=( a48578a  and  a48573a );
 a48583a <=( A269  and  (not A268) );
 a48584a <=( A267  and  a48583a );
 a48587a <=( (not A299)  and  A298 );
 a48590a <=( (not A302)  and  A300 );
 a48591a <=( a48590a  and  a48587a );
 a48592a <=( a48591a  and  a48584a );
 a48596a <=( A167  and  A168 );
 a48597a <=( A169  and  a48596a );
 a48601a <=( (not A203)  and  (not A201) );
 a48602a <=( (not A166)  and  a48601a );
 a48603a <=( a48602a  and  a48597a );
 a48607a <=( A269  and  (not A268) );
 a48608a <=( A267  and  a48607a );
 a48611a <=( A299  and  (not A298) );
 a48614a <=( A301  and  A300 );
 a48615a <=( a48614a  and  a48611a );
 a48616a <=( a48615a  and  a48608a );
 a48620a <=( A167  and  A168 );
 a48621a <=( A169  and  a48620a );
 a48625a <=( (not A203)  and  (not A201) );
 a48626a <=( (not A166)  and  a48625a );
 a48627a <=( a48626a  and  a48621a );
 a48631a <=( A269  and  (not A268) );
 a48632a <=( A267  and  a48631a );
 a48635a <=( A299  and  (not A298) );
 a48638a <=( (not A302)  and  A300 );
 a48639a <=( a48638a  and  a48635a );
 a48640a <=( a48639a  and  a48632a );
 a48644a <=( A167  and  A168 );
 a48645a <=( A169  and  a48644a );
 a48649a <=( (not A203)  and  (not A201) );
 a48650a <=( (not A166)  and  a48649a );
 a48651a <=( a48650a  and  a48645a );
 a48655a <=( A298  and  A268 );
 a48656a <=( (not A267)  and  a48655a );
 a48659a <=( (not A300)  and  (not A299) );
 a48662a <=( A302  and  (not A301) );
 a48663a <=( a48662a  and  a48659a );
 a48664a <=( a48663a  and  a48656a );
 a48668a <=( A167  and  A168 );
 a48669a <=( A169  and  a48668a );
 a48673a <=( (not A203)  and  (not A201) );
 a48674a <=( (not A166)  and  a48673a );
 a48675a <=( a48674a  and  a48669a );
 a48679a <=( (not A298)  and  A268 );
 a48680a <=( (not A267)  and  a48679a );
 a48683a <=( (not A300)  and  A299 );
 a48686a <=( A302  and  (not A301) );
 a48687a <=( a48686a  and  a48683a );
 a48688a <=( a48687a  and  a48680a );
 a48692a <=( A167  and  A168 );
 a48693a <=( A169  and  a48692a );
 a48697a <=( (not A203)  and  (not A201) );
 a48698a <=( (not A166)  and  a48697a );
 a48699a <=( a48698a  and  a48693a );
 a48703a <=( A298  and  (not A269) );
 a48704a <=( (not A267)  and  a48703a );
 a48707a <=( (not A300)  and  (not A299) );
 a48710a <=( A302  and  (not A301) );
 a48711a <=( a48710a  and  a48707a );
 a48712a <=( a48711a  and  a48704a );
 a48716a <=( A167  and  A168 );
 a48717a <=( A169  and  a48716a );
 a48721a <=( (not A203)  and  (not A201) );
 a48722a <=( (not A166)  and  a48721a );
 a48723a <=( a48722a  and  a48717a );
 a48727a <=( (not A298)  and  (not A269) );
 a48728a <=( (not A267)  and  a48727a );
 a48731a <=( (not A300)  and  A299 );
 a48734a <=( A302  and  (not A301) );
 a48735a <=( a48734a  and  a48731a );
 a48736a <=( a48735a  and  a48728a );
 a48740a <=( A167  and  A168 );
 a48741a <=( A169  and  a48740a );
 a48745a <=( (not A203)  and  (not A201) );
 a48746a <=( (not A166)  and  a48745a );
 a48747a <=( a48746a  and  a48741a );
 a48751a <=( A298  and  A266 );
 a48752a <=( A265  and  a48751a );
 a48755a <=( (not A300)  and  (not A299) );
 a48758a <=( A302  and  (not A301) );
 a48759a <=( a48758a  and  a48755a );
 a48760a <=( a48759a  and  a48752a );
 a48764a <=( A167  and  A168 );
 a48765a <=( A169  and  a48764a );
 a48769a <=( (not A203)  and  (not A201) );
 a48770a <=( (not A166)  and  a48769a );
 a48771a <=( a48770a  and  a48765a );
 a48775a <=( (not A298)  and  A266 );
 a48776a <=( A265  and  a48775a );
 a48779a <=( (not A300)  and  A299 );
 a48782a <=( A302  and  (not A301) );
 a48783a <=( a48782a  and  a48779a );
 a48784a <=( a48783a  and  a48776a );
 a48788a <=( A167  and  A168 );
 a48789a <=( A169  and  a48788a );
 a48793a <=( (not A203)  and  (not A201) );
 a48794a <=( (not A166)  and  a48793a );
 a48795a <=( a48794a  and  a48789a );
 a48799a <=( A267  and  A266 );
 a48800a <=( (not A265)  and  a48799a );
 a48803a <=( A300  and  A268 );
 a48806a <=( A302  and  (not A301) );
 a48807a <=( a48806a  and  a48803a );
 a48808a <=( a48807a  and  a48800a );
 a48812a <=( A167  and  A168 );
 a48813a <=( A169  and  a48812a );
 a48817a <=( (not A203)  and  (not A201) );
 a48818a <=( (not A166)  and  a48817a );
 a48819a <=( a48818a  and  a48813a );
 a48823a <=( A267  and  A266 );
 a48824a <=( (not A265)  and  a48823a );
 a48827a <=( A300  and  (not A269) );
 a48830a <=( A302  and  (not A301) );
 a48831a <=( a48830a  and  a48827a );
 a48832a <=( a48831a  and  a48824a );
 a48836a <=( A167  and  A168 );
 a48837a <=( A169  and  a48836a );
 a48841a <=( (not A203)  and  (not A201) );
 a48842a <=( (not A166)  and  a48841a );
 a48843a <=( a48842a  and  a48837a );
 a48847a <=( (not A267)  and  A266 );
 a48848a <=( (not A265)  and  a48847a );
 a48851a <=( A269  and  (not A268) );
 a48854a <=( A301  and  (not A300) );
 a48855a <=( a48854a  and  a48851a );
 a48856a <=( a48855a  and  a48848a );
 a48860a <=( A167  and  A168 );
 a48861a <=( A169  and  a48860a );
 a48865a <=( (not A203)  and  (not A201) );
 a48866a <=( (not A166)  and  a48865a );
 a48867a <=( a48866a  and  a48861a );
 a48871a <=( (not A267)  and  A266 );
 a48872a <=( (not A265)  and  a48871a );
 a48875a <=( A269  and  (not A268) );
 a48878a <=( (not A302)  and  (not A300) );
 a48879a <=( a48878a  and  a48875a );
 a48880a <=( a48879a  and  a48872a );
 a48884a <=( A167  and  A168 );
 a48885a <=( A169  and  a48884a );
 a48889a <=( (not A203)  and  (not A201) );
 a48890a <=( (not A166)  and  a48889a );
 a48891a <=( a48890a  and  a48885a );
 a48895a <=( (not A267)  and  A266 );
 a48896a <=( (not A265)  and  a48895a );
 a48899a <=( A269  and  (not A268) );
 a48902a <=( A299  and  A298 );
 a48903a <=( a48902a  and  a48899a );
 a48904a <=( a48903a  and  a48896a );
 a48908a <=( A167  and  A168 );
 a48909a <=( A169  and  a48908a );
 a48913a <=( (not A203)  and  (not A201) );
 a48914a <=( (not A166)  and  a48913a );
 a48915a <=( a48914a  and  a48909a );
 a48919a <=( (not A267)  and  A266 );
 a48920a <=( (not A265)  and  a48919a );
 a48923a <=( A269  and  (not A268) );
 a48926a <=( (not A299)  and  (not A298) );
 a48927a <=( a48926a  and  a48923a );
 a48928a <=( a48927a  and  a48920a );
 a48932a <=( A167  and  A168 );
 a48933a <=( A169  and  a48932a );
 a48937a <=( (not A203)  and  (not A201) );
 a48938a <=( (not A166)  and  a48937a );
 a48939a <=( a48938a  and  a48933a );
 a48943a <=( A267  and  (not A266) );
 a48944a <=( A265  and  a48943a );
 a48947a <=( A300  and  A268 );
 a48950a <=( A302  and  (not A301) );
 a48951a <=( a48950a  and  a48947a );
 a48952a <=( a48951a  and  a48944a );
 a48956a <=( A167  and  A168 );
 a48957a <=( A169  and  a48956a );
 a48961a <=( (not A203)  and  (not A201) );
 a48962a <=( (not A166)  and  a48961a );
 a48963a <=( a48962a  and  a48957a );
 a48967a <=( A267  and  (not A266) );
 a48968a <=( A265  and  a48967a );
 a48971a <=( A300  and  (not A269) );
 a48974a <=( A302  and  (not A301) );
 a48975a <=( a48974a  and  a48971a );
 a48976a <=( a48975a  and  a48968a );
 a48980a <=( A167  and  A168 );
 a48981a <=( A169  and  a48980a );
 a48985a <=( (not A203)  and  (not A201) );
 a48986a <=( (not A166)  and  a48985a );
 a48987a <=( a48986a  and  a48981a );
 a48991a <=( (not A267)  and  (not A266) );
 a48992a <=( A265  and  a48991a );
 a48995a <=( A269  and  (not A268) );
 a48998a <=( A301  and  (not A300) );
 a48999a <=( a48998a  and  a48995a );
 a49000a <=( a48999a  and  a48992a );
 a49004a <=( A167  and  A168 );
 a49005a <=( A169  and  a49004a );
 a49009a <=( (not A203)  and  (not A201) );
 a49010a <=( (not A166)  and  a49009a );
 a49011a <=( a49010a  and  a49005a );
 a49015a <=( (not A267)  and  (not A266) );
 a49016a <=( A265  and  a49015a );
 a49019a <=( A269  and  (not A268) );
 a49022a <=( (not A302)  and  (not A300) );
 a49023a <=( a49022a  and  a49019a );
 a49024a <=( a49023a  and  a49016a );
 a49028a <=( A167  and  A168 );
 a49029a <=( A169  and  a49028a );
 a49033a <=( (not A203)  and  (not A201) );
 a49034a <=( (not A166)  and  a49033a );
 a49035a <=( a49034a  and  a49029a );
 a49039a <=( (not A267)  and  (not A266) );
 a49040a <=( A265  and  a49039a );
 a49043a <=( A269  and  (not A268) );
 a49046a <=( A299  and  A298 );
 a49047a <=( a49046a  and  a49043a );
 a49048a <=( a49047a  and  a49040a );
 a49052a <=( A167  and  A168 );
 a49053a <=( A169  and  a49052a );
 a49057a <=( (not A203)  and  (not A201) );
 a49058a <=( (not A166)  and  a49057a );
 a49059a <=( a49058a  and  a49053a );
 a49063a <=( (not A267)  and  (not A266) );
 a49064a <=( A265  and  a49063a );
 a49067a <=( A269  and  (not A268) );
 a49070a <=( (not A299)  and  (not A298) );
 a49071a <=( a49070a  and  a49067a );
 a49072a <=( a49071a  and  a49064a );
 a49076a <=( A167  and  A168 );
 a49077a <=( A169  and  a49076a );
 a49081a <=( (not A203)  and  (not A201) );
 a49082a <=( (not A166)  and  a49081a );
 a49083a <=( a49082a  and  a49077a );
 a49087a <=( A298  and  (not A266) );
 a49088a <=( (not A265)  and  a49087a );
 a49091a <=( (not A300)  and  (not A299) );
 a49094a <=( A302  and  (not A301) );
 a49095a <=( a49094a  and  a49091a );
 a49096a <=( a49095a  and  a49088a );
 a49100a <=( A167  and  A168 );
 a49101a <=( A169  and  a49100a );
 a49105a <=( (not A203)  and  (not A201) );
 a49106a <=( (not A166)  and  a49105a );
 a49107a <=( a49106a  and  a49101a );
 a49111a <=( (not A298)  and  (not A266) );
 a49112a <=( (not A265)  and  a49111a );
 a49115a <=( (not A300)  and  A299 );
 a49118a <=( A302  and  (not A301) );
 a49119a <=( a49118a  and  a49115a );
 a49120a <=( a49119a  and  a49112a );
 a49124a <=( A167  and  A168 );
 a49125a <=( A169  and  a49124a );
 a49129a <=( A200  and  A199 );
 a49130a <=( (not A166)  and  a49129a );
 a49131a <=( a49130a  and  a49125a );
 a49135a <=( A269  and  (not A268) );
 a49136a <=( A267  and  a49135a );
 a49139a <=( (not A299)  and  A298 );
 a49142a <=( A301  and  A300 );
 a49143a <=( a49142a  and  a49139a );
 a49144a <=( a49143a  and  a49136a );
 a49148a <=( A167  and  A168 );
 a49149a <=( A169  and  a49148a );
 a49153a <=( A200  and  A199 );
 a49154a <=( (not A166)  and  a49153a );
 a49155a <=( a49154a  and  a49149a );
 a49159a <=( A269  and  (not A268) );
 a49160a <=( A267  and  a49159a );
 a49163a <=( (not A299)  and  A298 );
 a49166a <=( (not A302)  and  A300 );
 a49167a <=( a49166a  and  a49163a );
 a49168a <=( a49167a  and  a49160a );
 a49172a <=( A167  and  A168 );
 a49173a <=( A169  and  a49172a );
 a49177a <=( A200  and  A199 );
 a49178a <=( (not A166)  and  a49177a );
 a49179a <=( a49178a  and  a49173a );
 a49183a <=( A269  and  (not A268) );
 a49184a <=( A267  and  a49183a );
 a49187a <=( A299  and  (not A298) );
 a49190a <=( A301  and  A300 );
 a49191a <=( a49190a  and  a49187a );
 a49192a <=( a49191a  and  a49184a );
 a49196a <=( A167  and  A168 );
 a49197a <=( A169  and  a49196a );
 a49201a <=( A200  and  A199 );
 a49202a <=( (not A166)  and  a49201a );
 a49203a <=( a49202a  and  a49197a );
 a49207a <=( A269  and  (not A268) );
 a49208a <=( A267  and  a49207a );
 a49211a <=( A299  and  (not A298) );
 a49214a <=( (not A302)  and  A300 );
 a49215a <=( a49214a  and  a49211a );
 a49216a <=( a49215a  and  a49208a );
 a49220a <=( A167  and  A168 );
 a49221a <=( A169  and  a49220a );
 a49225a <=( A200  and  A199 );
 a49226a <=( (not A166)  and  a49225a );
 a49227a <=( a49226a  and  a49221a );
 a49231a <=( A298  and  A268 );
 a49232a <=( (not A267)  and  a49231a );
 a49235a <=( (not A300)  and  (not A299) );
 a49238a <=( A302  and  (not A301) );
 a49239a <=( a49238a  and  a49235a );
 a49240a <=( a49239a  and  a49232a );
 a49244a <=( A167  and  A168 );
 a49245a <=( A169  and  a49244a );
 a49249a <=( A200  and  A199 );
 a49250a <=( (not A166)  and  a49249a );
 a49251a <=( a49250a  and  a49245a );
 a49255a <=( (not A298)  and  A268 );
 a49256a <=( (not A267)  and  a49255a );
 a49259a <=( (not A300)  and  A299 );
 a49262a <=( A302  and  (not A301) );
 a49263a <=( a49262a  and  a49259a );
 a49264a <=( a49263a  and  a49256a );
 a49268a <=( A167  and  A168 );
 a49269a <=( A169  and  a49268a );
 a49273a <=( A200  and  A199 );
 a49274a <=( (not A166)  and  a49273a );
 a49275a <=( a49274a  and  a49269a );
 a49279a <=( A298  and  (not A269) );
 a49280a <=( (not A267)  and  a49279a );
 a49283a <=( (not A300)  and  (not A299) );
 a49286a <=( A302  and  (not A301) );
 a49287a <=( a49286a  and  a49283a );
 a49288a <=( a49287a  and  a49280a );
 a49292a <=( A167  and  A168 );
 a49293a <=( A169  and  a49292a );
 a49297a <=( A200  and  A199 );
 a49298a <=( (not A166)  and  a49297a );
 a49299a <=( a49298a  and  a49293a );
 a49303a <=( (not A298)  and  (not A269) );
 a49304a <=( (not A267)  and  a49303a );
 a49307a <=( (not A300)  and  A299 );
 a49310a <=( A302  and  (not A301) );
 a49311a <=( a49310a  and  a49307a );
 a49312a <=( a49311a  and  a49304a );
 a49316a <=( A167  and  A168 );
 a49317a <=( A169  and  a49316a );
 a49321a <=( A200  and  A199 );
 a49322a <=( (not A166)  and  a49321a );
 a49323a <=( a49322a  and  a49317a );
 a49327a <=( A298  and  A266 );
 a49328a <=( A265  and  a49327a );
 a49331a <=( (not A300)  and  (not A299) );
 a49334a <=( A302  and  (not A301) );
 a49335a <=( a49334a  and  a49331a );
 a49336a <=( a49335a  and  a49328a );
 a49340a <=( A167  and  A168 );
 a49341a <=( A169  and  a49340a );
 a49345a <=( A200  and  A199 );
 a49346a <=( (not A166)  and  a49345a );
 a49347a <=( a49346a  and  a49341a );
 a49351a <=( (not A298)  and  A266 );
 a49352a <=( A265  and  a49351a );
 a49355a <=( (not A300)  and  A299 );
 a49358a <=( A302  and  (not A301) );
 a49359a <=( a49358a  and  a49355a );
 a49360a <=( a49359a  and  a49352a );
 a49364a <=( A167  and  A168 );
 a49365a <=( A169  and  a49364a );
 a49369a <=( A200  and  A199 );
 a49370a <=( (not A166)  and  a49369a );
 a49371a <=( a49370a  and  a49365a );
 a49375a <=( A267  and  A266 );
 a49376a <=( (not A265)  and  a49375a );
 a49379a <=( A300  and  A268 );
 a49382a <=( A302  and  (not A301) );
 a49383a <=( a49382a  and  a49379a );
 a49384a <=( a49383a  and  a49376a );
 a49388a <=( A167  and  A168 );
 a49389a <=( A169  and  a49388a );
 a49393a <=( A200  and  A199 );
 a49394a <=( (not A166)  and  a49393a );
 a49395a <=( a49394a  and  a49389a );
 a49399a <=( A267  and  A266 );
 a49400a <=( (not A265)  and  a49399a );
 a49403a <=( A300  and  (not A269) );
 a49406a <=( A302  and  (not A301) );
 a49407a <=( a49406a  and  a49403a );
 a49408a <=( a49407a  and  a49400a );
 a49412a <=( A167  and  A168 );
 a49413a <=( A169  and  a49412a );
 a49417a <=( A200  and  A199 );
 a49418a <=( (not A166)  and  a49417a );
 a49419a <=( a49418a  and  a49413a );
 a49423a <=( (not A267)  and  A266 );
 a49424a <=( (not A265)  and  a49423a );
 a49427a <=( A269  and  (not A268) );
 a49430a <=( A301  and  (not A300) );
 a49431a <=( a49430a  and  a49427a );
 a49432a <=( a49431a  and  a49424a );
 a49436a <=( A167  and  A168 );
 a49437a <=( A169  and  a49436a );
 a49441a <=( A200  and  A199 );
 a49442a <=( (not A166)  and  a49441a );
 a49443a <=( a49442a  and  a49437a );
 a49447a <=( (not A267)  and  A266 );
 a49448a <=( (not A265)  and  a49447a );
 a49451a <=( A269  and  (not A268) );
 a49454a <=( (not A302)  and  (not A300) );
 a49455a <=( a49454a  and  a49451a );
 a49456a <=( a49455a  and  a49448a );
 a49460a <=( A167  and  A168 );
 a49461a <=( A169  and  a49460a );
 a49465a <=( A200  and  A199 );
 a49466a <=( (not A166)  and  a49465a );
 a49467a <=( a49466a  and  a49461a );
 a49471a <=( (not A267)  and  A266 );
 a49472a <=( (not A265)  and  a49471a );
 a49475a <=( A269  and  (not A268) );
 a49478a <=( A299  and  A298 );
 a49479a <=( a49478a  and  a49475a );
 a49480a <=( a49479a  and  a49472a );
 a49484a <=( A167  and  A168 );
 a49485a <=( A169  and  a49484a );
 a49489a <=( A200  and  A199 );
 a49490a <=( (not A166)  and  a49489a );
 a49491a <=( a49490a  and  a49485a );
 a49495a <=( (not A267)  and  A266 );
 a49496a <=( (not A265)  and  a49495a );
 a49499a <=( A269  and  (not A268) );
 a49502a <=( (not A299)  and  (not A298) );
 a49503a <=( a49502a  and  a49499a );
 a49504a <=( a49503a  and  a49496a );
 a49508a <=( A167  and  A168 );
 a49509a <=( A169  and  a49508a );
 a49513a <=( A200  and  A199 );
 a49514a <=( (not A166)  and  a49513a );
 a49515a <=( a49514a  and  a49509a );
 a49519a <=( A267  and  (not A266) );
 a49520a <=( A265  and  a49519a );
 a49523a <=( A300  and  A268 );
 a49526a <=( A302  and  (not A301) );
 a49527a <=( a49526a  and  a49523a );
 a49528a <=( a49527a  and  a49520a );
 a49532a <=( A167  and  A168 );
 a49533a <=( A169  and  a49532a );
 a49537a <=( A200  and  A199 );
 a49538a <=( (not A166)  and  a49537a );
 a49539a <=( a49538a  and  a49533a );
 a49543a <=( A267  and  (not A266) );
 a49544a <=( A265  and  a49543a );
 a49547a <=( A300  and  (not A269) );
 a49550a <=( A302  and  (not A301) );
 a49551a <=( a49550a  and  a49547a );
 a49552a <=( a49551a  and  a49544a );
 a49556a <=( A167  and  A168 );
 a49557a <=( A169  and  a49556a );
 a49561a <=( A200  and  A199 );
 a49562a <=( (not A166)  and  a49561a );
 a49563a <=( a49562a  and  a49557a );
 a49567a <=( (not A267)  and  (not A266) );
 a49568a <=( A265  and  a49567a );
 a49571a <=( A269  and  (not A268) );
 a49574a <=( A301  and  (not A300) );
 a49575a <=( a49574a  and  a49571a );
 a49576a <=( a49575a  and  a49568a );
 a49580a <=( A167  and  A168 );
 a49581a <=( A169  and  a49580a );
 a49585a <=( A200  and  A199 );
 a49586a <=( (not A166)  and  a49585a );
 a49587a <=( a49586a  and  a49581a );
 a49591a <=( (not A267)  and  (not A266) );
 a49592a <=( A265  and  a49591a );
 a49595a <=( A269  and  (not A268) );
 a49598a <=( (not A302)  and  (not A300) );
 a49599a <=( a49598a  and  a49595a );
 a49600a <=( a49599a  and  a49592a );
 a49604a <=( A167  and  A168 );
 a49605a <=( A169  and  a49604a );
 a49609a <=( A200  and  A199 );
 a49610a <=( (not A166)  and  a49609a );
 a49611a <=( a49610a  and  a49605a );
 a49615a <=( (not A267)  and  (not A266) );
 a49616a <=( A265  and  a49615a );
 a49619a <=( A269  and  (not A268) );
 a49622a <=( A299  and  A298 );
 a49623a <=( a49622a  and  a49619a );
 a49624a <=( a49623a  and  a49616a );
 a49628a <=( A167  and  A168 );
 a49629a <=( A169  and  a49628a );
 a49633a <=( A200  and  A199 );
 a49634a <=( (not A166)  and  a49633a );
 a49635a <=( a49634a  and  a49629a );
 a49639a <=( (not A267)  and  (not A266) );
 a49640a <=( A265  and  a49639a );
 a49643a <=( A269  and  (not A268) );
 a49646a <=( (not A299)  and  (not A298) );
 a49647a <=( a49646a  and  a49643a );
 a49648a <=( a49647a  and  a49640a );
 a49652a <=( A167  and  A168 );
 a49653a <=( A169  and  a49652a );
 a49657a <=( A200  and  A199 );
 a49658a <=( (not A166)  and  a49657a );
 a49659a <=( a49658a  and  a49653a );
 a49663a <=( A298  and  (not A266) );
 a49664a <=( (not A265)  and  a49663a );
 a49667a <=( (not A300)  and  (not A299) );
 a49670a <=( A302  and  (not A301) );
 a49671a <=( a49670a  and  a49667a );
 a49672a <=( a49671a  and  a49664a );
 a49676a <=( A167  and  A168 );
 a49677a <=( A169  and  a49676a );
 a49681a <=( A200  and  A199 );
 a49682a <=( (not A166)  and  a49681a );
 a49683a <=( a49682a  and  a49677a );
 a49687a <=( (not A298)  and  (not A266) );
 a49688a <=( (not A265)  and  a49687a );
 a49691a <=( (not A300)  and  A299 );
 a49694a <=( A302  and  (not A301) );
 a49695a <=( a49694a  and  a49691a );
 a49696a <=( a49695a  and  a49688a );
 a49700a <=( A167  and  A168 );
 a49701a <=( A169  and  a49700a );
 a49705a <=( (not A200)  and  (not A199) );
 a49706a <=( (not A166)  and  a49705a );
 a49707a <=( a49706a  and  a49701a );
 a49711a <=( A269  and  (not A268) );
 a49712a <=( A267  and  a49711a );
 a49715a <=( (not A299)  and  A298 );
 a49718a <=( A301  and  A300 );
 a49719a <=( a49718a  and  a49715a );
 a49720a <=( a49719a  and  a49712a );
 a49724a <=( A167  and  A168 );
 a49725a <=( A169  and  a49724a );
 a49729a <=( (not A200)  and  (not A199) );
 a49730a <=( (not A166)  and  a49729a );
 a49731a <=( a49730a  and  a49725a );
 a49735a <=( A269  and  (not A268) );
 a49736a <=( A267  and  a49735a );
 a49739a <=( (not A299)  and  A298 );
 a49742a <=( (not A302)  and  A300 );
 a49743a <=( a49742a  and  a49739a );
 a49744a <=( a49743a  and  a49736a );
 a49748a <=( A167  and  A168 );
 a49749a <=( A169  and  a49748a );
 a49753a <=( (not A200)  and  (not A199) );
 a49754a <=( (not A166)  and  a49753a );
 a49755a <=( a49754a  and  a49749a );
 a49759a <=( A269  and  (not A268) );
 a49760a <=( A267  and  a49759a );
 a49763a <=( A299  and  (not A298) );
 a49766a <=( A301  and  A300 );
 a49767a <=( a49766a  and  a49763a );
 a49768a <=( a49767a  and  a49760a );
 a49772a <=( A167  and  A168 );
 a49773a <=( A169  and  a49772a );
 a49777a <=( (not A200)  and  (not A199) );
 a49778a <=( (not A166)  and  a49777a );
 a49779a <=( a49778a  and  a49773a );
 a49783a <=( A269  and  (not A268) );
 a49784a <=( A267  and  a49783a );
 a49787a <=( A299  and  (not A298) );
 a49790a <=( (not A302)  and  A300 );
 a49791a <=( a49790a  and  a49787a );
 a49792a <=( a49791a  and  a49784a );
 a49796a <=( A167  and  A168 );
 a49797a <=( A169  and  a49796a );
 a49801a <=( (not A200)  and  (not A199) );
 a49802a <=( (not A166)  and  a49801a );
 a49803a <=( a49802a  and  a49797a );
 a49807a <=( A298  and  A268 );
 a49808a <=( (not A267)  and  a49807a );
 a49811a <=( (not A300)  and  (not A299) );
 a49814a <=( A302  and  (not A301) );
 a49815a <=( a49814a  and  a49811a );
 a49816a <=( a49815a  and  a49808a );
 a49820a <=( A167  and  A168 );
 a49821a <=( A169  and  a49820a );
 a49825a <=( (not A200)  and  (not A199) );
 a49826a <=( (not A166)  and  a49825a );
 a49827a <=( a49826a  and  a49821a );
 a49831a <=( (not A298)  and  A268 );
 a49832a <=( (not A267)  and  a49831a );
 a49835a <=( (not A300)  and  A299 );
 a49838a <=( A302  and  (not A301) );
 a49839a <=( a49838a  and  a49835a );
 a49840a <=( a49839a  and  a49832a );
 a49844a <=( A167  and  A168 );
 a49845a <=( A169  and  a49844a );
 a49849a <=( (not A200)  and  (not A199) );
 a49850a <=( (not A166)  and  a49849a );
 a49851a <=( a49850a  and  a49845a );
 a49855a <=( A298  and  (not A269) );
 a49856a <=( (not A267)  and  a49855a );
 a49859a <=( (not A300)  and  (not A299) );
 a49862a <=( A302  and  (not A301) );
 a49863a <=( a49862a  and  a49859a );
 a49864a <=( a49863a  and  a49856a );
 a49868a <=( A167  and  A168 );
 a49869a <=( A169  and  a49868a );
 a49873a <=( (not A200)  and  (not A199) );
 a49874a <=( (not A166)  and  a49873a );
 a49875a <=( a49874a  and  a49869a );
 a49879a <=( (not A298)  and  (not A269) );
 a49880a <=( (not A267)  and  a49879a );
 a49883a <=( (not A300)  and  A299 );
 a49886a <=( A302  and  (not A301) );
 a49887a <=( a49886a  and  a49883a );
 a49888a <=( a49887a  and  a49880a );
 a49892a <=( A167  and  A168 );
 a49893a <=( A169  and  a49892a );
 a49897a <=( (not A200)  and  (not A199) );
 a49898a <=( (not A166)  and  a49897a );
 a49899a <=( a49898a  and  a49893a );
 a49903a <=( A298  and  A266 );
 a49904a <=( A265  and  a49903a );
 a49907a <=( (not A300)  and  (not A299) );
 a49910a <=( A302  and  (not A301) );
 a49911a <=( a49910a  and  a49907a );
 a49912a <=( a49911a  and  a49904a );
 a49916a <=( A167  and  A168 );
 a49917a <=( A169  and  a49916a );
 a49921a <=( (not A200)  and  (not A199) );
 a49922a <=( (not A166)  and  a49921a );
 a49923a <=( a49922a  and  a49917a );
 a49927a <=( (not A298)  and  A266 );
 a49928a <=( A265  and  a49927a );
 a49931a <=( (not A300)  and  A299 );
 a49934a <=( A302  and  (not A301) );
 a49935a <=( a49934a  and  a49931a );
 a49936a <=( a49935a  and  a49928a );
 a49940a <=( A167  and  A168 );
 a49941a <=( A169  and  a49940a );
 a49945a <=( (not A200)  and  (not A199) );
 a49946a <=( (not A166)  and  a49945a );
 a49947a <=( a49946a  and  a49941a );
 a49951a <=( A267  and  A266 );
 a49952a <=( (not A265)  and  a49951a );
 a49955a <=( A300  and  A268 );
 a49958a <=( A302  and  (not A301) );
 a49959a <=( a49958a  and  a49955a );
 a49960a <=( a49959a  and  a49952a );
 a49964a <=( A167  and  A168 );
 a49965a <=( A169  and  a49964a );
 a49969a <=( (not A200)  and  (not A199) );
 a49970a <=( (not A166)  and  a49969a );
 a49971a <=( a49970a  and  a49965a );
 a49975a <=( A267  and  A266 );
 a49976a <=( (not A265)  and  a49975a );
 a49979a <=( A300  and  (not A269) );
 a49982a <=( A302  and  (not A301) );
 a49983a <=( a49982a  and  a49979a );
 a49984a <=( a49983a  and  a49976a );
 a49988a <=( A167  and  A168 );
 a49989a <=( A169  and  a49988a );
 a49993a <=( (not A200)  and  (not A199) );
 a49994a <=( (not A166)  and  a49993a );
 a49995a <=( a49994a  and  a49989a );
 a49999a <=( (not A267)  and  A266 );
 a50000a <=( (not A265)  and  a49999a );
 a50003a <=( A269  and  (not A268) );
 a50006a <=( A301  and  (not A300) );
 a50007a <=( a50006a  and  a50003a );
 a50008a <=( a50007a  and  a50000a );
 a50012a <=( A167  and  A168 );
 a50013a <=( A169  and  a50012a );
 a50017a <=( (not A200)  and  (not A199) );
 a50018a <=( (not A166)  and  a50017a );
 a50019a <=( a50018a  and  a50013a );
 a50023a <=( (not A267)  and  A266 );
 a50024a <=( (not A265)  and  a50023a );
 a50027a <=( A269  and  (not A268) );
 a50030a <=( (not A302)  and  (not A300) );
 a50031a <=( a50030a  and  a50027a );
 a50032a <=( a50031a  and  a50024a );
 a50036a <=( A167  and  A168 );
 a50037a <=( A169  and  a50036a );
 a50041a <=( (not A200)  and  (not A199) );
 a50042a <=( (not A166)  and  a50041a );
 a50043a <=( a50042a  and  a50037a );
 a50047a <=( (not A267)  and  A266 );
 a50048a <=( (not A265)  and  a50047a );
 a50051a <=( A269  and  (not A268) );
 a50054a <=( A299  and  A298 );
 a50055a <=( a50054a  and  a50051a );
 a50056a <=( a50055a  and  a50048a );
 a50060a <=( A167  and  A168 );
 a50061a <=( A169  and  a50060a );
 a50065a <=( (not A200)  and  (not A199) );
 a50066a <=( (not A166)  and  a50065a );
 a50067a <=( a50066a  and  a50061a );
 a50071a <=( (not A267)  and  A266 );
 a50072a <=( (not A265)  and  a50071a );
 a50075a <=( A269  and  (not A268) );
 a50078a <=( (not A299)  and  (not A298) );
 a50079a <=( a50078a  and  a50075a );
 a50080a <=( a50079a  and  a50072a );
 a50084a <=( A167  and  A168 );
 a50085a <=( A169  and  a50084a );
 a50089a <=( (not A200)  and  (not A199) );
 a50090a <=( (not A166)  and  a50089a );
 a50091a <=( a50090a  and  a50085a );
 a50095a <=( A267  and  (not A266) );
 a50096a <=( A265  and  a50095a );
 a50099a <=( A300  and  A268 );
 a50102a <=( A302  and  (not A301) );
 a50103a <=( a50102a  and  a50099a );
 a50104a <=( a50103a  and  a50096a );
 a50108a <=( A167  and  A168 );
 a50109a <=( A169  and  a50108a );
 a50113a <=( (not A200)  and  (not A199) );
 a50114a <=( (not A166)  and  a50113a );
 a50115a <=( a50114a  and  a50109a );
 a50119a <=( A267  and  (not A266) );
 a50120a <=( A265  and  a50119a );
 a50123a <=( A300  and  (not A269) );
 a50126a <=( A302  and  (not A301) );
 a50127a <=( a50126a  and  a50123a );
 a50128a <=( a50127a  and  a50120a );
 a50132a <=( A167  and  A168 );
 a50133a <=( A169  and  a50132a );
 a50137a <=( (not A200)  and  (not A199) );
 a50138a <=( (not A166)  and  a50137a );
 a50139a <=( a50138a  and  a50133a );
 a50143a <=( (not A267)  and  (not A266) );
 a50144a <=( A265  and  a50143a );
 a50147a <=( A269  and  (not A268) );
 a50150a <=( A301  and  (not A300) );
 a50151a <=( a50150a  and  a50147a );
 a50152a <=( a50151a  and  a50144a );
 a50156a <=( A167  and  A168 );
 a50157a <=( A169  and  a50156a );
 a50161a <=( (not A200)  and  (not A199) );
 a50162a <=( (not A166)  and  a50161a );
 a50163a <=( a50162a  and  a50157a );
 a50167a <=( (not A267)  and  (not A266) );
 a50168a <=( A265  and  a50167a );
 a50171a <=( A269  and  (not A268) );
 a50174a <=( (not A302)  and  (not A300) );
 a50175a <=( a50174a  and  a50171a );
 a50176a <=( a50175a  and  a50168a );
 a50180a <=( A167  and  A168 );
 a50181a <=( A169  and  a50180a );
 a50185a <=( (not A200)  and  (not A199) );
 a50186a <=( (not A166)  and  a50185a );
 a50187a <=( a50186a  and  a50181a );
 a50191a <=( (not A267)  and  (not A266) );
 a50192a <=( A265  and  a50191a );
 a50195a <=( A269  and  (not A268) );
 a50198a <=( A299  and  A298 );
 a50199a <=( a50198a  and  a50195a );
 a50200a <=( a50199a  and  a50192a );
 a50204a <=( A167  and  A168 );
 a50205a <=( A169  and  a50204a );
 a50209a <=( (not A200)  and  (not A199) );
 a50210a <=( (not A166)  and  a50209a );
 a50211a <=( a50210a  and  a50205a );
 a50215a <=( (not A267)  and  (not A266) );
 a50216a <=( A265  and  a50215a );
 a50219a <=( A269  and  (not A268) );
 a50222a <=( (not A299)  and  (not A298) );
 a50223a <=( a50222a  and  a50219a );
 a50224a <=( a50223a  and  a50216a );
 a50228a <=( A167  and  A168 );
 a50229a <=( A169  and  a50228a );
 a50233a <=( (not A200)  and  (not A199) );
 a50234a <=( (not A166)  and  a50233a );
 a50235a <=( a50234a  and  a50229a );
 a50239a <=( A298  and  (not A266) );
 a50240a <=( (not A265)  and  a50239a );
 a50243a <=( (not A300)  and  (not A299) );
 a50246a <=( A302  and  (not A301) );
 a50247a <=( a50246a  and  a50243a );
 a50248a <=( a50247a  and  a50240a );
 a50252a <=( A167  and  A168 );
 a50253a <=( A169  and  a50252a );
 a50257a <=( (not A200)  and  (not A199) );
 a50258a <=( (not A166)  and  a50257a );
 a50259a <=( a50258a  and  a50253a );
 a50263a <=( (not A298)  and  (not A266) );
 a50264a <=( (not A265)  and  a50263a );
 a50267a <=( (not A300)  and  A299 );
 a50270a <=( A302  and  (not A301) );
 a50271a <=( a50270a  and  a50267a );
 a50272a <=( a50271a  and  a50264a );
 a50276a <=( (not A167)  and  A168 );
 a50277a <=( A169  and  a50276a );
 a50281a <=( (not A202)  and  A201 );
 a50282a <=( A166  and  a50281a );
 a50283a <=( a50282a  and  a50277a );
 a50287a <=( A268  and  (not A267) );
 a50288a <=( A203  and  a50287a );
 a50291a <=( (not A299)  and  A298 );
 a50294a <=( A301  and  A300 );
 a50295a <=( a50294a  and  a50291a );
 a50296a <=( a50295a  and  a50288a );
 a50300a <=( (not A167)  and  A168 );
 a50301a <=( A169  and  a50300a );
 a50305a <=( (not A202)  and  A201 );
 a50306a <=( A166  and  a50305a );
 a50307a <=( a50306a  and  a50301a );
 a50311a <=( A268  and  (not A267) );
 a50312a <=( A203  and  a50311a );
 a50315a <=( (not A299)  and  A298 );
 a50318a <=( (not A302)  and  A300 );
 a50319a <=( a50318a  and  a50315a );
 a50320a <=( a50319a  and  a50312a );
 a50324a <=( (not A167)  and  A168 );
 a50325a <=( A169  and  a50324a );
 a50329a <=( (not A202)  and  A201 );
 a50330a <=( A166  and  a50329a );
 a50331a <=( a50330a  and  a50325a );
 a50335a <=( A268  and  (not A267) );
 a50336a <=( A203  and  a50335a );
 a50339a <=( A299  and  (not A298) );
 a50342a <=( A301  and  A300 );
 a50343a <=( a50342a  and  a50339a );
 a50344a <=( a50343a  and  a50336a );
 a50348a <=( (not A167)  and  A168 );
 a50349a <=( A169  and  a50348a );
 a50353a <=( (not A202)  and  A201 );
 a50354a <=( A166  and  a50353a );
 a50355a <=( a50354a  and  a50349a );
 a50359a <=( A268  and  (not A267) );
 a50360a <=( A203  and  a50359a );
 a50363a <=( A299  and  (not A298) );
 a50366a <=( (not A302)  and  A300 );
 a50367a <=( a50366a  and  a50363a );
 a50368a <=( a50367a  and  a50360a );
 a50372a <=( (not A167)  and  A168 );
 a50373a <=( A169  and  a50372a );
 a50377a <=( (not A202)  and  A201 );
 a50378a <=( A166  and  a50377a );
 a50379a <=( a50378a  and  a50373a );
 a50383a <=( (not A269)  and  (not A267) );
 a50384a <=( A203  and  a50383a );
 a50387a <=( (not A299)  and  A298 );
 a50390a <=( A301  and  A300 );
 a50391a <=( a50390a  and  a50387a );
 a50392a <=( a50391a  and  a50384a );
 a50396a <=( (not A167)  and  A168 );
 a50397a <=( A169  and  a50396a );
 a50401a <=( (not A202)  and  A201 );
 a50402a <=( A166  and  a50401a );
 a50403a <=( a50402a  and  a50397a );
 a50407a <=( (not A269)  and  (not A267) );
 a50408a <=( A203  and  a50407a );
 a50411a <=( (not A299)  and  A298 );
 a50414a <=( (not A302)  and  A300 );
 a50415a <=( a50414a  and  a50411a );
 a50416a <=( a50415a  and  a50408a );
 a50420a <=( (not A167)  and  A168 );
 a50421a <=( A169  and  a50420a );
 a50425a <=( (not A202)  and  A201 );
 a50426a <=( A166  and  a50425a );
 a50427a <=( a50426a  and  a50421a );
 a50431a <=( (not A269)  and  (not A267) );
 a50432a <=( A203  and  a50431a );
 a50435a <=( A299  and  (not A298) );
 a50438a <=( A301  and  A300 );
 a50439a <=( a50438a  and  a50435a );
 a50440a <=( a50439a  and  a50432a );
 a50444a <=( (not A167)  and  A168 );
 a50445a <=( A169  and  a50444a );
 a50449a <=( (not A202)  and  A201 );
 a50450a <=( A166  and  a50449a );
 a50451a <=( a50450a  and  a50445a );
 a50455a <=( (not A269)  and  (not A267) );
 a50456a <=( A203  and  a50455a );
 a50459a <=( A299  and  (not A298) );
 a50462a <=( (not A302)  and  A300 );
 a50463a <=( a50462a  and  a50459a );
 a50464a <=( a50463a  and  a50456a );
 a50468a <=( (not A167)  and  A168 );
 a50469a <=( A169  and  a50468a );
 a50473a <=( (not A202)  and  A201 );
 a50474a <=( A166  and  a50473a );
 a50475a <=( a50474a  and  a50469a );
 a50479a <=( A266  and  A265 );
 a50480a <=( A203  and  a50479a );
 a50483a <=( (not A299)  and  A298 );
 a50486a <=( A301  and  A300 );
 a50487a <=( a50486a  and  a50483a );
 a50488a <=( a50487a  and  a50480a );
 a50492a <=( (not A167)  and  A168 );
 a50493a <=( A169  and  a50492a );
 a50497a <=( (not A202)  and  A201 );
 a50498a <=( A166  and  a50497a );
 a50499a <=( a50498a  and  a50493a );
 a50503a <=( A266  and  A265 );
 a50504a <=( A203  and  a50503a );
 a50507a <=( (not A299)  and  A298 );
 a50510a <=( (not A302)  and  A300 );
 a50511a <=( a50510a  and  a50507a );
 a50512a <=( a50511a  and  a50504a );
 a50516a <=( (not A167)  and  A168 );
 a50517a <=( A169  and  a50516a );
 a50521a <=( (not A202)  and  A201 );
 a50522a <=( A166  and  a50521a );
 a50523a <=( a50522a  and  a50517a );
 a50527a <=( A266  and  A265 );
 a50528a <=( A203  and  a50527a );
 a50531a <=( A299  and  (not A298) );
 a50534a <=( A301  and  A300 );
 a50535a <=( a50534a  and  a50531a );
 a50536a <=( a50535a  and  a50528a );
 a50540a <=( (not A167)  and  A168 );
 a50541a <=( A169  and  a50540a );
 a50545a <=( (not A202)  and  A201 );
 a50546a <=( A166  and  a50545a );
 a50547a <=( a50546a  and  a50541a );
 a50551a <=( A266  and  A265 );
 a50552a <=( A203  and  a50551a );
 a50555a <=( A299  and  (not A298) );
 a50558a <=( (not A302)  and  A300 );
 a50559a <=( a50558a  and  a50555a );
 a50560a <=( a50559a  and  a50552a );
 a50564a <=( (not A167)  and  A168 );
 a50565a <=( A169  and  a50564a );
 a50569a <=( (not A202)  and  A201 );
 a50570a <=( A166  and  a50569a );
 a50571a <=( a50570a  and  a50565a );
 a50575a <=( A266  and  (not A265) );
 a50576a <=( A203  and  a50575a );
 a50579a <=( A268  and  A267 );
 a50582a <=( A301  and  (not A300) );
 a50583a <=( a50582a  and  a50579a );
 a50584a <=( a50583a  and  a50576a );
 a50588a <=( (not A167)  and  A168 );
 a50589a <=( A169  and  a50588a );
 a50593a <=( (not A202)  and  A201 );
 a50594a <=( A166  and  a50593a );
 a50595a <=( a50594a  and  a50589a );
 a50599a <=( A266  and  (not A265) );
 a50600a <=( A203  and  a50599a );
 a50603a <=( A268  and  A267 );
 a50606a <=( (not A302)  and  (not A300) );
 a50607a <=( a50606a  and  a50603a );
 a50608a <=( a50607a  and  a50600a );
 a50612a <=( (not A167)  and  A168 );
 a50613a <=( A169  and  a50612a );
 a50617a <=( (not A202)  and  A201 );
 a50618a <=( A166  and  a50617a );
 a50619a <=( a50618a  and  a50613a );
 a50623a <=( A266  and  (not A265) );
 a50624a <=( A203  and  a50623a );
 a50627a <=( A268  and  A267 );
 a50630a <=( A299  and  A298 );
 a50631a <=( a50630a  and  a50627a );
 a50632a <=( a50631a  and  a50624a );
 a50636a <=( (not A167)  and  A168 );
 a50637a <=( A169  and  a50636a );
 a50641a <=( (not A202)  and  A201 );
 a50642a <=( A166  and  a50641a );
 a50643a <=( a50642a  and  a50637a );
 a50647a <=( A266  and  (not A265) );
 a50648a <=( A203  and  a50647a );
 a50651a <=( A268  and  A267 );
 a50654a <=( (not A299)  and  (not A298) );
 a50655a <=( a50654a  and  a50651a );
 a50656a <=( a50655a  and  a50648a );
 a50660a <=( (not A167)  and  A168 );
 a50661a <=( A169  and  a50660a );
 a50665a <=( (not A202)  and  A201 );
 a50666a <=( A166  and  a50665a );
 a50667a <=( a50666a  and  a50661a );
 a50671a <=( A266  and  (not A265) );
 a50672a <=( A203  and  a50671a );
 a50675a <=( (not A269)  and  A267 );
 a50678a <=( A301  and  (not A300) );
 a50679a <=( a50678a  and  a50675a );
 a50680a <=( a50679a  and  a50672a );
 a50684a <=( (not A167)  and  A168 );
 a50685a <=( A169  and  a50684a );
 a50689a <=( (not A202)  and  A201 );
 a50690a <=( A166  and  a50689a );
 a50691a <=( a50690a  and  a50685a );
 a50695a <=( A266  and  (not A265) );
 a50696a <=( A203  and  a50695a );
 a50699a <=( (not A269)  and  A267 );
 a50702a <=( (not A302)  and  (not A300) );
 a50703a <=( a50702a  and  a50699a );
 a50704a <=( a50703a  and  a50696a );
 a50708a <=( (not A167)  and  A168 );
 a50709a <=( A169  and  a50708a );
 a50713a <=( (not A202)  and  A201 );
 a50714a <=( A166  and  a50713a );
 a50715a <=( a50714a  and  a50709a );
 a50719a <=( A266  and  (not A265) );
 a50720a <=( A203  and  a50719a );
 a50723a <=( (not A269)  and  A267 );
 a50726a <=( A299  and  A298 );
 a50727a <=( a50726a  and  a50723a );
 a50728a <=( a50727a  and  a50720a );
 a50732a <=( (not A167)  and  A168 );
 a50733a <=( A169  and  a50732a );
 a50737a <=( (not A202)  and  A201 );
 a50738a <=( A166  and  a50737a );
 a50739a <=( a50738a  and  a50733a );
 a50743a <=( A266  and  (not A265) );
 a50744a <=( A203  and  a50743a );
 a50747a <=( (not A269)  and  A267 );
 a50750a <=( (not A299)  and  (not A298) );
 a50751a <=( a50750a  and  a50747a );
 a50752a <=( a50751a  and  a50744a );
 a50756a <=( (not A167)  and  A168 );
 a50757a <=( A169  and  a50756a );
 a50761a <=( (not A202)  and  A201 );
 a50762a <=( A166  and  a50761a );
 a50763a <=( a50762a  and  a50757a );
 a50767a <=( (not A266)  and  A265 );
 a50768a <=( A203  and  a50767a );
 a50771a <=( A268  and  A267 );
 a50774a <=( A301  and  (not A300) );
 a50775a <=( a50774a  and  a50771a );
 a50776a <=( a50775a  and  a50768a );
 a50780a <=( (not A167)  and  A168 );
 a50781a <=( A169  and  a50780a );
 a50785a <=( (not A202)  and  A201 );
 a50786a <=( A166  and  a50785a );
 a50787a <=( a50786a  and  a50781a );
 a50791a <=( (not A266)  and  A265 );
 a50792a <=( A203  and  a50791a );
 a50795a <=( A268  and  A267 );
 a50798a <=( (not A302)  and  (not A300) );
 a50799a <=( a50798a  and  a50795a );
 a50800a <=( a50799a  and  a50792a );
 a50804a <=( (not A167)  and  A168 );
 a50805a <=( A169  and  a50804a );
 a50809a <=( (not A202)  and  A201 );
 a50810a <=( A166  and  a50809a );
 a50811a <=( a50810a  and  a50805a );
 a50815a <=( (not A266)  and  A265 );
 a50816a <=( A203  and  a50815a );
 a50819a <=( A268  and  A267 );
 a50822a <=( A299  and  A298 );
 a50823a <=( a50822a  and  a50819a );
 a50824a <=( a50823a  and  a50816a );
 a50828a <=( (not A167)  and  A168 );
 a50829a <=( A169  and  a50828a );
 a50833a <=( (not A202)  and  A201 );
 a50834a <=( A166  and  a50833a );
 a50835a <=( a50834a  and  a50829a );
 a50839a <=( (not A266)  and  A265 );
 a50840a <=( A203  and  a50839a );
 a50843a <=( A268  and  A267 );
 a50846a <=( (not A299)  and  (not A298) );
 a50847a <=( a50846a  and  a50843a );
 a50848a <=( a50847a  and  a50840a );
 a50852a <=( (not A167)  and  A168 );
 a50853a <=( A169  and  a50852a );
 a50857a <=( (not A202)  and  A201 );
 a50858a <=( A166  and  a50857a );
 a50859a <=( a50858a  and  a50853a );
 a50863a <=( (not A266)  and  A265 );
 a50864a <=( A203  and  a50863a );
 a50867a <=( (not A269)  and  A267 );
 a50870a <=( A301  and  (not A300) );
 a50871a <=( a50870a  and  a50867a );
 a50872a <=( a50871a  and  a50864a );
 a50876a <=( (not A167)  and  A168 );
 a50877a <=( A169  and  a50876a );
 a50881a <=( (not A202)  and  A201 );
 a50882a <=( A166  and  a50881a );
 a50883a <=( a50882a  and  a50877a );
 a50887a <=( (not A266)  and  A265 );
 a50888a <=( A203  and  a50887a );
 a50891a <=( (not A269)  and  A267 );
 a50894a <=( (not A302)  and  (not A300) );
 a50895a <=( a50894a  and  a50891a );
 a50896a <=( a50895a  and  a50888a );
 a50900a <=( (not A167)  and  A168 );
 a50901a <=( A169  and  a50900a );
 a50905a <=( (not A202)  and  A201 );
 a50906a <=( A166  and  a50905a );
 a50907a <=( a50906a  and  a50901a );
 a50911a <=( (not A266)  and  A265 );
 a50912a <=( A203  and  a50911a );
 a50915a <=( (not A269)  and  A267 );
 a50918a <=( A299  and  A298 );
 a50919a <=( a50918a  and  a50915a );
 a50920a <=( a50919a  and  a50912a );
 a50924a <=( (not A167)  and  A168 );
 a50925a <=( A169  and  a50924a );
 a50929a <=( (not A202)  and  A201 );
 a50930a <=( A166  and  a50929a );
 a50931a <=( a50930a  and  a50925a );
 a50935a <=( (not A266)  and  A265 );
 a50936a <=( A203  and  a50935a );
 a50939a <=( (not A269)  and  A267 );
 a50942a <=( (not A299)  and  (not A298) );
 a50943a <=( a50942a  and  a50939a );
 a50944a <=( a50943a  and  a50936a );
 a50948a <=( (not A167)  and  A168 );
 a50949a <=( A169  and  a50948a );
 a50953a <=( (not A202)  and  A201 );
 a50954a <=( A166  and  a50953a );
 a50955a <=( a50954a  and  a50949a );
 a50959a <=( (not A266)  and  (not A265) );
 a50960a <=( A203  and  a50959a );
 a50963a <=( (not A299)  and  A298 );
 a50966a <=( A301  and  A300 );
 a50967a <=( a50966a  and  a50963a );
 a50968a <=( a50967a  and  a50960a );
 a50972a <=( (not A167)  and  A168 );
 a50973a <=( A169  and  a50972a );
 a50977a <=( (not A202)  and  A201 );
 a50978a <=( A166  and  a50977a );
 a50979a <=( a50978a  and  a50973a );
 a50983a <=( (not A266)  and  (not A265) );
 a50984a <=( A203  and  a50983a );
 a50987a <=( (not A299)  and  A298 );
 a50990a <=( (not A302)  and  A300 );
 a50991a <=( a50990a  and  a50987a );
 a50992a <=( a50991a  and  a50984a );
 a50996a <=( (not A167)  and  A168 );
 a50997a <=( A169  and  a50996a );
 a51001a <=( (not A202)  and  A201 );
 a51002a <=( A166  and  a51001a );
 a51003a <=( a51002a  and  a50997a );
 a51007a <=( (not A266)  and  (not A265) );
 a51008a <=( A203  and  a51007a );
 a51011a <=( A299  and  (not A298) );
 a51014a <=( A301  and  A300 );
 a51015a <=( a51014a  and  a51011a );
 a51016a <=( a51015a  and  a51008a );
 a51020a <=( (not A167)  and  A168 );
 a51021a <=( A169  and  a51020a );
 a51025a <=( (not A202)  and  A201 );
 a51026a <=( A166  and  a51025a );
 a51027a <=( a51026a  and  a51021a );
 a51031a <=( (not A266)  and  (not A265) );
 a51032a <=( A203  and  a51031a );
 a51035a <=( A299  and  (not A298) );
 a51038a <=( (not A302)  and  A300 );
 a51039a <=( a51038a  and  a51035a );
 a51040a <=( a51039a  and  a51032a );
 a51044a <=( (not A167)  and  A168 );
 a51045a <=( A169  and  a51044a );
 a51049a <=( A202  and  (not A201) );
 a51050a <=( A166  and  a51049a );
 a51051a <=( a51050a  and  a51045a );
 a51055a <=( A269  and  (not A268) );
 a51056a <=( A267  and  a51055a );
 a51059a <=( (not A299)  and  A298 );
 a51062a <=( A301  and  A300 );
 a51063a <=( a51062a  and  a51059a );
 a51064a <=( a51063a  and  a51056a );
 a51068a <=( (not A167)  and  A168 );
 a51069a <=( A169  and  a51068a );
 a51073a <=( A202  and  (not A201) );
 a51074a <=( A166  and  a51073a );
 a51075a <=( a51074a  and  a51069a );
 a51079a <=( A269  and  (not A268) );
 a51080a <=( A267  and  a51079a );
 a51083a <=( (not A299)  and  A298 );
 a51086a <=( (not A302)  and  A300 );
 a51087a <=( a51086a  and  a51083a );
 a51088a <=( a51087a  and  a51080a );
 a51092a <=( (not A167)  and  A168 );
 a51093a <=( A169  and  a51092a );
 a51097a <=( A202  and  (not A201) );
 a51098a <=( A166  and  a51097a );
 a51099a <=( a51098a  and  a51093a );
 a51103a <=( A269  and  (not A268) );
 a51104a <=( A267  and  a51103a );
 a51107a <=( A299  and  (not A298) );
 a51110a <=( A301  and  A300 );
 a51111a <=( a51110a  and  a51107a );
 a51112a <=( a51111a  and  a51104a );
 a51116a <=( (not A167)  and  A168 );
 a51117a <=( A169  and  a51116a );
 a51121a <=( A202  and  (not A201) );
 a51122a <=( A166  and  a51121a );
 a51123a <=( a51122a  and  a51117a );
 a51127a <=( A269  and  (not A268) );
 a51128a <=( A267  and  a51127a );
 a51131a <=( A299  and  (not A298) );
 a51134a <=( (not A302)  and  A300 );
 a51135a <=( a51134a  and  a51131a );
 a51136a <=( a51135a  and  a51128a );
 a51140a <=( (not A167)  and  A168 );
 a51141a <=( A169  and  a51140a );
 a51145a <=( A202  and  (not A201) );
 a51146a <=( A166  and  a51145a );
 a51147a <=( a51146a  and  a51141a );
 a51151a <=( A298  and  A268 );
 a51152a <=( (not A267)  and  a51151a );
 a51155a <=( (not A300)  and  (not A299) );
 a51158a <=( A302  and  (not A301) );
 a51159a <=( a51158a  and  a51155a );
 a51160a <=( a51159a  and  a51152a );
 a51164a <=( (not A167)  and  A168 );
 a51165a <=( A169  and  a51164a );
 a51169a <=( A202  and  (not A201) );
 a51170a <=( A166  and  a51169a );
 a51171a <=( a51170a  and  a51165a );
 a51175a <=( (not A298)  and  A268 );
 a51176a <=( (not A267)  and  a51175a );
 a51179a <=( (not A300)  and  A299 );
 a51182a <=( A302  and  (not A301) );
 a51183a <=( a51182a  and  a51179a );
 a51184a <=( a51183a  and  a51176a );
 a51188a <=( (not A167)  and  A168 );
 a51189a <=( A169  and  a51188a );
 a51193a <=( A202  and  (not A201) );
 a51194a <=( A166  and  a51193a );
 a51195a <=( a51194a  and  a51189a );
 a51199a <=( A298  and  (not A269) );
 a51200a <=( (not A267)  and  a51199a );
 a51203a <=( (not A300)  and  (not A299) );
 a51206a <=( A302  and  (not A301) );
 a51207a <=( a51206a  and  a51203a );
 a51208a <=( a51207a  and  a51200a );
 a51212a <=( (not A167)  and  A168 );
 a51213a <=( A169  and  a51212a );
 a51217a <=( A202  and  (not A201) );
 a51218a <=( A166  and  a51217a );
 a51219a <=( a51218a  and  a51213a );
 a51223a <=( (not A298)  and  (not A269) );
 a51224a <=( (not A267)  and  a51223a );
 a51227a <=( (not A300)  and  A299 );
 a51230a <=( A302  and  (not A301) );
 a51231a <=( a51230a  and  a51227a );
 a51232a <=( a51231a  and  a51224a );
 a51236a <=( (not A167)  and  A168 );
 a51237a <=( A169  and  a51236a );
 a51241a <=( A202  and  (not A201) );
 a51242a <=( A166  and  a51241a );
 a51243a <=( a51242a  and  a51237a );
 a51247a <=( A298  and  A266 );
 a51248a <=( A265  and  a51247a );
 a51251a <=( (not A300)  and  (not A299) );
 a51254a <=( A302  and  (not A301) );
 a51255a <=( a51254a  and  a51251a );
 a51256a <=( a51255a  and  a51248a );
 a51260a <=( (not A167)  and  A168 );
 a51261a <=( A169  and  a51260a );
 a51265a <=( A202  and  (not A201) );
 a51266a <=( A166  and  a51265a );
 a51267a <=( a51266a  and  a51261a );
 a51271a <=( (not A298)  and  A266 );
 a51272a <=( A265  and  a51271a );
 a51275a <=( (not A300)  and  A299 );
 a51278a <=( A302  and  (not A301) );
 a51279a <=( a51278a  and  a51275a );
 a51280a <=( a51279a  and  a51272a );
 a51284a <=( (not A167)  and  A168 );
 a51285a <=( A169  and  a51284a );
 a51289a <=( A202  and  (not A201) );
 a51290a <=( A166  and  a51289a );
 a51291a <=( a51290a  and  a51285a );
 a51295a <=( A267  and  A266 );
 a51296a <=( (not A265)  and  a51295a );
 a51299a <=( A300  and  A268 );
 a51302a <=( A302  and  (not A301) );
 a51303a <=( a51302a  and  a51299a );
 a51304a <=( a51303a  and  a51296a );
 a51308a <=( (not A167)  and  A168 );
 a51309a <=( A169  and  a51308a );
 a51313a <=( A202  and  (not A201) );
 a51314a <=( A166  and  a51313a );
 a51315a <=( a51314a  and  a51309a );
 a51319a <=( A267  and  A266 );
 a51320a <=( (not A265)  and  a51319a );
 a51323a <=( A300  and  (not A269) );
 a51326a <=( A302  and  (not A301) );
 a51327a <=( a51326a  and  a51323a );
 a51328a <=( a51327a  and  a51320a );
 a51332a <=( (not A167)  and  A168 );
 a51333a <=( A169  and  a51332a );
 a51337a <=( A202  and  (not A201) );
 a51338a <=( A166  and  a51337a );
 a51339a <=( a51338a  and  a51333a );
 a51343a <=( (not A267)  and  A266 );
 a51344a <=( (not A265)  and  a51343a );
 a51347a <=( A269  and  (not A268) );
 a51350a <=( A301  and  (not A300) );
 a51351a <=( a51350a  and  a51347a );
 a51352a <=( a51351a  and  a51344a );
 a51356a <=( (not A167)  and  A168 );
 a51357a <=( A169  and  a51356a );
 a51361a <=( A202  and  (not A201) );
 a51362a <=( A166  and  a51361a );
 a51363a <=( a51362a  and  a51357a );
 a51367a <=( (not A267)  and  A266 );
 a51368a <=( (not A265)  and  a51367a );
 a51371a <=( A269  and  (not A268) );
 a51374a <=( (not A302)  and  (not A300) );
 a51375a <=( a51374a  and  a51371a );
 a51376a <=( a51375a  and  a51368a );
 a51380a <=( (not A167)  and  A168 );
 a51381a <=( A169  and  a51380a );
 a51385a <=( A202  and  (not A201) );
 a51386a <=( A166  and  a51385a );
 a51387a <=( a51386a  and  a51381a );
 a51391a <=( (not A267)  and  A266 );
 a51392a <=( (not A265)  and  a51391a );
 a51395a <=( A269  and  (not A268) );
 a51398a <=( A299  and  A298 );
 a51399a <=( a51398a  and  a51395a );
 a51400a <=( a51399a  and  a51392a );
 a51404a <=( (not A167)  and  A168 );
 a51405a <=( A169  and  a51404a );
 a51409a <=( A202  and  (not A201) );
 a51410a <=( A166  and  a51409a );
 a51411a <=( a51410a  and  a51405a );
 a51415a <=( (not A267)  and  A266 );
 a51416a <=( (not A265)  and  a51415a );
 a51419a <=( A269  and  (not A268) );
 a51422a <=( (not A299)  and  (not A298) );
 a51423a <=( a51422a  and  a51419a );
 a51424a <=( a51423a  and  a51416a );
 a51428a <=( (not A167)  and  A168 );
 a51429a <=( A169  and  a51428a );
 a51433a <=( A202  and  (not A201) );
 a51434a <=( A166  and  a51433a );
 a51435a <=( a51434a  and  a51429a );
 a51439a <=( A267  and  (not A266) );
 a51440a <=( A265  and  a51439a );
 a51443a <=( A300  and  A268 );
 a51446a <=( A302  and  (not A301) );
 a51447a <=( a51446a  and  a51443a );
 a51448a <=( a51447a  and  a51440a );
 a51452a <=( (not A167)  and  A168 );
 a51453a <=( A169  and  a51452a );
 a51457a <=( A202  and  (not A201) );
 a51458a <=( A166  and  a51457a );
 a51459a <=( a51458a  and  a51453a );
 a51463a <=( A267  and  (not A266) );
 a51464a <=( A265  and  a51463a );
 a51467a <=( A300  and  (not A269) );
 a51470a <=( A302  and  (not A301) );
 a51471a <=( a51470a  and  a51467a );
 a51472a <=( a51471a  and  a51464a );
 a51476a <=( (not A167)  and  A168 );
 a51477a <=( A169  and  a51476a );
 a51481a <=( A202  and  (not A201) );
 a51482a <=( A166  and  a51481a );
 a51483a <=( a51482a  and  a51477a );
 a51487a <=( (not A267)  and  (not A266) );
 a51488a <=( A265  and  a51487a );
 a51491a <=( A269  and  (not A268) );
 a51494a <=( A301  and  (not A300) );
 a51495a <=( a51494a  and  a51491a );
 a51496a <=( a51495a  and  a51488a );
 a51500a <=( (not A167)  and  A168 );
 a51501a <=( A169  and  a51500a );
 a51505a <=( A202  and  (not A201) );
 a51506a <=( A166  and  a51505a );
 a51507a <=( a51506a  and  a51501a );
 a51511a <=( (not A267)  and  (not A266) );
 a51512a <=( A265  and  a51511a );
 a51515a <=( A269  and  (not A268) );
 a51518a <=( (not A302)  and  (not A300) );
 a51519a <=( a51518a  and  a51515a );
 a51520a <=( a51519a  and  a51512a );
 a51524a <=( (not A167)  and  A168 );
 a51525a <=( A169  and  a51524a );
 a51529a <=( A202  and  (not A201) );
 a51530a <=( A166  and  a51529a );
 a51531a <=( a51530a  and  a51525a );
 a51535a <=( (not A267)  and  (not A266) );
 a51536a <=( A265  and  a51535a );
 a51539a <=( A269  and  (not A268) );
 a51542a <=( A299  and  A298 );
 a51543a <=( a51542a  and  a51539a );
 a51544a <=( a51543a  and  a51536a );
 a51548a <=( (not A167)  and  A168 );
 a51549a <=( A169  and  a51548a );
 a51553a <=( A202  and  (not A201) );
 a51554a <=( A166  and  a51553a );
 a51555a <=( a51554a  and  a51549a );
 a51559a <=( (not A267)  and  (not A266) );
 a51560a <=( A265  and  a51559a );
 a51563a <=( A269  and  (not A268) );
 a51566a <=( (not A299)  and  (not A298) );
 a51567a <=( a51566a  and  a51563a );
 a51568a <=( a51567a  and  a51560a );
 a51572a <=( (not A167)  and  A168 );
 a51573a <=( A169  and  a51572a );
 a51577a <=( A202  and  (not A201) );
 a51578a <=( A166  and  a51577a );
 a51579a <=( a51578a  and  a51573a );
 a51583a <=( A298  and  (not A266) );
 a51584a <=( (not A265)  and  a51583a );
 a51587a <=( (not A300)  and  (not A299) );
 a51590a <=( A302  and  (not A301) );
 a51591a <=( a51590a  and  a51587a );
 a51592a <=( a51591a  and  a51584a );
 a51596a <=( (not A167)  and  A168 );
 a51597a <=( A169  and  a51596a );
 a51601a <=( A202  and  (not A201) );
 a51602a <=( A166  and  a51601a );
 a51603a <=( a51602a  and  a51597a );
 a51607a <=( (not A298)  and  (not A266) );
 a51608a <=( (not A265)  and  a51607a );
 a51611a <=( (not A300)  and  A299 );
 a51614a <=( A302  and  (not A301) );
 a51615a <=( a51614a  and  a51611a );
 a51616a <=( a51615a  and  a51608a );
 a51620a <=( (not A167)  and  A168 );
 a51621a <=( A169  and  a51620a );
 a51625a <=( (not A203)  and  (not A201) );
 a51626a <=( A166  and  a51625a );
 a51627a <=( a51626a  and  a51621a );
 a51631a <=( A269  and  (not A268) );
 a51632a <=( A267  and  a51631a );
 a51635a <=( (not A299)  and  A298 );
 a51638a <=( A301  and  A300 );
 a51639a <=( a51638a  and  a51635a );
 a51640a <=( a51639a  and  a51632a );
 a51644a <=( (not A167)  and  A168 );
 a51645a <=( A169  and  a51644a );
 a51649a <=( (not A203)  and  (not A201) );
 a51650a <=( A166  and  a51649a );
 a51651a <=( a51650a  and  a51645a );
 a51655a <=( A269  and  (not A268) );
 a51656a <=( A267  and  a51655a );
 a51659a <=( (not A299)  and  A298 );
 a51662a <=( (not A302)  and  A300 );
 a51663a <=( a51662a  and  a51659a );
 a51664a <=( a51663a  and  a51656a );
 a51668a <=( (not A167)  and  A168 );
 a51669a <=( A169  and  a51668a );
 a51673a <=( (not A203)  and  (not A201) );
 a51674a <=( A166  and  a51673a );
 a51675a <=( a51674a  and  a51669a );
 a51679a <=( A269  and  (not A268) );
 a51680a <=( A267  and  a51679a );
 a51683a <=( A299  and  (not A298) );
 a51686a <=( A301  and  A300 );
 a51687a <=( a51686a  and  a51683a );
 a51688a <=( a51687a  and  a51680a );
 a51692a <=( (not A167)  and  A168 );
 a51693a <=( A169  and  a51692a );
 a51697a <=( (not A203)  and  (not A201) );
 a51698a <=( A166  and  a51697a );
 a51699a <=( a51698a  and  a51693a );
 a51703a <=( A269  and  (not A268) );
 a51704a <=( A267  and  a51703a );
 a51707a <=( A299  and  (not A298) );
 a51710a <=( (not A302)  and  A300 );
 a51711a <=( a51710a  and  a51707a );
 a51712a <=( a51711a  and  a51704a );
 a51716a <=( (not A167)  and  A168 );
 a51717a <=( A169  and  a51716a );
 a51721a <=( (not A203)  and  (not A201) );
 a51722a <=( A166  and  a51721a );
 a51723a <=( a51722a  and  a51717a );
 a51727a <=( A298  and  A268 );
 a51728a <=( (not A267)  and  a51727a );
 a51731a <=( (not A300)  and  (not A299) );
 a51734a <=( A302  and  (not A301) );
 a51735a <=( a51734a  and  a51731a );
 a51736a <=( a51735a  and  a51728a );
 a51740a <=( (not A167)  and  A168 );
 a51741a <=( A169  and  a51740a );
 a51745a <=( (not A203)  and  (not A201) );
 a51746a <=( A166  and  a51745a );
 a51747a <=( a51746a  and  a51741a );
 a51751a <=( (not A298)  and  A268 );
 a51752a <=( (not A267)  and  a51751a );
 a51755a <=( (not A300)  and  A299 );
 a51758a <=( A302  and  (not A301) );
 a51759a <=( a51758a  and  a51755a );
 a51760a <=( a51759a  and  a51752a );
 a51764a <=( (not A167)  and  A168 );
 a51765a <=( A169  and  a51764a );
 a51769a <=( (not A203)  and  (not A201) );
 a51770a <=( A166  and  a51769a );
 a51771a <=( a51770a  and  a51765a );
 a51775a <=( A298  and  (not A269) );
 a51776a <=( (not A267)  and  a51775a );
 a51779a <=( (not A300)  and  (not A299) );
 a51782a <=( A302  and  (not A301) );
 a51783a <=( a51782a  and  a51779a );
 a51784a <=( a51783a  and  a51776a );
 a51788a <=( (not A167)  and  A168 );
 a51789a <=( A169  and  a51788a );
 a51793a <=( (not A203)  and  (not A201) );
 a51794a <=( A166  and  a51793a );
 a51795a <=( a51794a  and  a51789a );
 a51799a <=( (not A298)  and  (not A269) );
 a51800a <=( (not A267)  and  a51799a );
 a51803a <=( (not A300)  and  A299 );
 a51806a <=( A302  and  (not A301) );
 a51807a <=( a51806a  and  a51803a );
 a51808a <=( a51807a  and  a51800a );
 a51812a <=( (not A167)  and  A168 );
 a51813a <=( A169  and  a51812a );
 a51817a <=( (not A203)  and  (not A201) );
 a51818a <=( A166  and  a51817a );
 a51819a <=( a51818a  and  a51813a );
 a51823a <=( A298  and  A266 );
 a51824a <=( A265  and  a51823a );
 a51827a <=( (not A300)  and  (not A299) );
 a51830a <=( A302  and  (not A301) );
 a51831a <=( a51830a  and  a51827a );
 a51832a <=( a51831a  and  a51824a );
 a51836a <=( (not A167)  and  A168 );
 a51837a <=( A169  and  a51836a );
 a51841a <=( (not A203)  and  (not A201) );
 a51842a <=( A166  and  a51841a );
 a51843a <=( a51842a  and  a51837a );
 a51847a <=( (not A298)  and  A266 );
 a51848a <=( A265  and  a51847a );
 a51851a <=( (not A300)  and  A299 );
 a51854a <=( A302  and  (not A301) );
 a51855a <=( a51854a  and  a51851a );
 a51856a <=( a51855a  and  a51848a );
 a51860a <=( (not A167)  and  A168 );
 a51861a <=( A169  and  a51860a );
 a51865a <=( (not A203)  and  (not A201) );
 a51866a <=( A166  and  a51865a );
 a51867a <=( a51866a  and  a51861a );
 a51871a <=( A267  and  A266 );
 a51872a <=( (not A265)  and  a51871a );
 a51875a <=( A300  and  A268 );
 a51878a <=( A302  and  (not A301) );
 a51879a <=( a51878a  and  a51875a );
 a51880a <=( a51879a  and  a51872a );
 a51884a <=( (not A167)  and  A168 );
 a51885a <=( A169  and  a51884a );
 a51889a <=( (not A203)  and  (not A201) );
 a51890a <=( A166  and  a51889a );
 a51891a <=( a51890a  and  a51885a );
 a51895a <=( A267  and  A266 );
 a51896a <=( (not A265)  and  a51895a );
 a51899a <=( A300  and  (not A269) );
 a51902a <=( A302  and  (not A301) );
 a51903a <=( a51902a  and  a51899a );
 a51904a <=( a51903a  and  a51896a );
 a51908a <=( (not A167)  and  A168 );
 a51909a <=( A169  and  a51908a );
 a51913a <=( (not A203)  and  (not A201) );
 a51914a <=( A166  and  a51913a );
 a51915a <=( a51914a  and  a51909a );
 a51919a <=( (not A267)  and  A266 );
 a51920a <=( (not A265)  and  a51919a );
 a51923a <=( A269  and  (not A268) );
 a51926a <=( A301  and  (not A300) );
 a51927a <=( a51926a  and  a51923a );
 a51928a <=( a51927a  and  a51920a );
 a51932a <=( (not A167)  and  A168 );
 a51933a <=( A169  and  a51932a );
 a51937a <=( (not A203)  and  (not A201) );
 a51938a <=( A166  and  a51937a );
 a51939a <=( a51938a  and  a51933a );
 a51943a <=( (not A267)  and  A266 );
 a51944a <=( (not A265)  and  a51943a );
 a51947a <=( A269  and  (not A268) );
 a51950a <=( (not A302)  and  (not A300) );
 a51951a <=( a51950a  and  a51947a );
 a51952a <=( a51951a  and  a51944a );
 a51956a <=( (not A167)  and  A168 );
 a51957a <=( A169  and  a51956a );
 a51961a <=( (not A203)  and  (not A201) );
 a51962a <=( A166  and  a51961a );
 a51963a <=( a51962a  and  a51957a );
 a51967a <=( (not A267)  and  A266 );
 a51968a <=( (not A265)  and  a51967a );
 a51971a <=( A269  and  (not A268) );
 a51974a <=( A299  and  A298 );
 a51975a <=( a51974a  and  a51971a );
 a51976a <=( a51975a  and  a51968a );
 a51980a <=( (not A167)  and  A168 );
 a51981a <=( A169  and  a51980a );
 a51985a <=( (not A203)  and  (not A201) );
 a51986a <=( A166  and  a51985a );
 a51987a <=( a51986a  and  a51981a );
 a51991a <=( (not A267)  and  A266 );
 a51992a <=( (not A265)  and  a51991a );
 a51995a <=( A269  and  (not A268) );
 a51998a <=( (not A299)  and  (not A298) );
 a51999a <=( a51998a  and  a51995a );
 a52000a <=( a51999a  and  a51992a );
 a52004a <=( (not A167)  and  A168 );
 a52005a <=( A169  and  a52004a );
 a52009a <=( (not A203)  and  (not A201) );
 a52010a <=( A166  and  a52009a );
 a52011a <=( a52010a  and  a52005a );
 a52015a <=( A267  and  (not A266) );
 a52016a <=( A265  and  a52015a );
 a52019a <=( A300  and  A268 );
 a52022a <=( A302  and  (not A301) );
 a52023a <=( a52022a  and  a52019a );
 a52024a <=( a52023a  and  a52016a );
 a52028a <=( (not A167)  and  A168 );
 a52029a <=( A169  and  a52028a );
 a52033a <=( (not A203)  and  (not A201) );
 a52034a <=( A166  and  a52033a );
 a52035a <=( a52034a  and  a52029a );
 a52039a <=( A267  and  (not A266) );
 a52040a <=( A265  and  a52039a );
 a52043a <=( A300  and  (not A269) );
 a52046a <=( A302  and  (not A301) );
 a52047a <=( a52046a  and  a52043a );
 a52048a <=( a52047a  and  a52040a );
 a52052a <=( (not A167)  and  A168 );
 a52053a <=( A169  and  a52052a );
 a52057a <=( (not A203)  and  (not A201) );
 a52058a <=( A166  and  a52057a );
 a52059a <=( a52058a  and  a52053a );
 a52063a <=( (not A267)  and  (not A266) );
 a52064a <=( A265  and  a52063a );
 a52067a <=( A269  and  (not A268) );
 a52070a <=( A301  and  (not A300) );
 a52071a <=( a52070a  and  a52067a );
 a52072a <=( a52071a  and  a52064a );
 a52076a <=( (not A167)  and  A168 );
 a52077a <=( A169  and  a52076a );
 a52081a <=( (not A203)  and  (not A201) );
 a52082a <=( A166  and  a52081a );
 a52083a <=( a52082a  and  a52077a );
 a52087a <=( (not A267)  and  (not A266) );
 a52088a <=( A265  and  a52087a );
 a52091a <=( A269  and  (not A268) );
 a52094a <=( (not A302)  and  (not A300) );
 a52095a <=( a52094a  and  a52091a );
 a52096a <=( a52095a  and  a52088a );
 a52100a <=( (not A167)  and  A168 );
 a52101a <=( A169  and  a52100a );
 a52105a <=( (not A203)  and  (not A201) );
 a52106a <=( A166  and  a52105a );
 a52107a <=( a52106a  and  a52101a );
 a52111a <=( (not A267)  and  (not A266) );
 a52112a <=( A265  and  a52111a );
 a52115a <=( A269  and  (not A268) );
 a52118a <=( A299  and  A298 );
 a52119a <=( a52118a  and  a52115a );
 a52120a <=( a52119a  and  a52112a );
 a52124a <=( (not A167)  and  A168 );
 a52125a <=( A169  and  a52124a );
 a52129a <=( (not A203)  and  (not A201) );
 a52130a <=( A166  and  a52129a );
 a52131a <=( a52130a  and  a52125a );
 a52135a <=( (not A267)  and  (not A266) );
 a52136a <=( A265  and  a52135a );
 a52139a <=( A269  and  (not A268) );
 a52142a <=( (not A299)  and  (not A298) );
 a52143a <=( a52142a  and  a52139a );
 a52144a <=( a52143a  and  a52136a );
 a52148a <=( (not A167)  and  A168 );
 a52149a <=( A169  and  a52148a );
 a52153a <=( (not A203)  and  (not A201) );
 a52154a <=( A166  and  a52153a );
 a52155a <=( a52154a  and  a52149a );
 a52159a <=( A298  and  (not A266) );
 a52160a <=( (not A265)  and  a52159a );
 a52163a <=( (not A300)  and  (not A299) );
 a52166a <=( A302  and  (not A301) );
 a52167a <=( a52166a  and  a52163a );
 a52168a <=( a52167a  and  a52160a );
 a52172a <=( (not A167)  and  A168 );
 a52173a <=( A169  and  a52172a );
 a52177a <=( (not A203)  and  (not A201) );
 a52178a <=( A166  and  a52177a );
 a52179a <=( a52178a  and  a52173a );
 a52183a <=( (not A298)  and  (not A266) );
 a52184a <=( (not A265)  and  a52183a );
 a52187a <=( (not A300)  and  A299 );
 a52190a <=( A302  and  (not A301) );
 a52191a <=( a52190a  and  a52187a );
 a52192a <=( a52191a  and  a52184a );
 a52196a <=( (not A167)  and  A168 );
 a52197a <=( A169  and  a52196a );
 a52201a <=( A200  and  A199 );
 a52202a <=( A166  and  a52201a );
 a52203a <=( a52202a  and  a52197a );
 a52207a <=( A269  and  (not A268) );
 a52208a <=( A267  and  a52207a );
 a52211a <=( (not A299)  and  A298 );
 a52214a <=( A301  and  A300 );
 a52215a <=( a52214a  and  a52211a );
 a52216a <=( a52215a  and  a52208a );
 a52220a <=( (not A167)  and  A168 );
 a52221a <=( A169  and  a52220a );
 a52225a <=( A200  and  A199 );
 a52226a <=( A166  and  a52225a );
 a52227a <=( a52226a  and  a52221a );
 a52231a <=( A269  and  (not A268) );
 a52232a <=( A267  and  a52231a );
 a52235a <=( (not A299)  and  A298 );
 a52238a <=( (not A302)  and  A300 );
 a52239a <=( a52238a  and  a52235a );
 a52240a <=( a52239a  and  a52232a );
 a52244a <=( (not A167)  and  A168 );
 a52245a <=( A169  and  a52244a );
 a52249a <=( A200  and  A199 );
 a52250a <=( A166  and  a52249a );
 a52251a <=( a52250a  and  a52245a );
 a52255a <=( A269  and  (not A268) );
 a52256a <=( A267  and  a52255a );
 a52259a <=( A299  and  (not A298) );
 a52262a <=( A301  and  A300 );
 a52263a <=( a52262a  and  a52259a );
 a52264a <=( a52263a  and  a52256a );
 a52268a <=( (not A167)  and  A168 );
 a52269a <=( A169  and  a52268a );
 a52273a <=( A200  and  A199 );
 a52274a <=( A166  and  a52273a );
 a52275a <=( a52274a  and  a52269a );
 a52279a <=( A269  and  (not A268) );
 a52280a <=( A267  and  a52279a );
 a52283a <=( A299  and  (not A298) );
 a52286a <=( (not A302)  and  A300 );
 a52287a <=( a52286a  and  a52283a );
 a52288a <=( a52287a  and  a52280a );
 a52292a <=( (not A167)  and  A168 );
 a52293a <=( A169  and  a52292a );
 a52297a <=( A200  and  A199 );
 a52298a <=( A166  and  a52297a );
 a52299a <=( a52298a  and  a52293a );
 a52303a <=( A298  and  A268 );
 a52304a <=( (not A267)  and  a52303a );
 a52307a <=( (not A300)  and  (not A299) );
 a52310a <=( A302  and  (not A301) );
 a52311a <=( a52310a  and  a52307a );
 a52312a <=( a52311a  and  a52304a );
 a52316a <=( (not A167)  and  A168 );
 a52317a <=( A169  and  a52316a );
 a52321a <=( A200  and  A199 );
 a52322a <=( A166  and  a52321a );
 a52323a <=( a52322a  and  a52317a );
 a52327a <=( (not A298)  and  A268 );
 a52328a <=( (not A267)  and  a52327a );
 a52331a <=( (not A300)  and  A299 );
 a52334a <=( A302  and  (not A301) );
 a52335a <=( a52334a  and  a52331a );
 a52336a <=( a52335a  and  a52328a );
 a52340a <=( (not A167)  and  A168 );
 a52341a <=( A169  and  a52340a );
 a52345a <=( A200  and  A199 );
 a52346a <=( A166  and  a52345a );
 a52347a <=( a52346a  and  a52341a );
 a52351a <=( A298  and  (not A269) );
 a52352a <=( (not A267)  and  a52351a );
 a52355a <=( (not A300)  and  (not A299) );
 a52358a <=( A302  and  (not A301) );
 a52359a <=( a52358a  and  a52355a );
 a52360a <=( a52359a  and  a52352a );
 a52364a <=( (not A167)  and  A168 );
 a52365a <=( A169  and  a52364a );
 a52369a <=( A200  and  A199 );
 a52370a <=( A166  and  a52369a );
 a52371a <=( a52370a  and  a52365a );
 a52375a <=( (not A298)  and  (not A269) );
 a52376a <=( (not A267)  and  a52375a );
 a52379a <=( (not A300)  and  A299 );
 a52382a <=( A302  and  (not A301) );
 a52383a <=( a52382a  and  a52379a );
 a52384a <=( a52383a  and  a52376a );
 a52388a <=( (not A167)  and  A168 );
 a52389a <=( A169  and  a52388a );
 a52393a <=( A200  and  A199 );
 a52394a <=( A166  and  a52393a );
 a52395a <=( a52394a  and  a52389a );
 a52399a <=( A298  and  A266 );
 a52400a <=( A265  and  a52399a );
 a52403a <=( (not A300)  and  (not A299) );
 a52406a <=( A302  and  (not A301) );
 a52407a <=( a52406a  and  a52403a );
 a52408a <=( a52407a  and  a52400a );
 a52412a <=( (not A167)  and  A168 );
 a52413a <=( A169  and  a52412a );
 a52417a <=( A200  and  A199 );
 a52418a <=( A166  and  a52417a );
 a52419a <=( a52418a  and  a52413a );
 a52423a <=( (not A298)  and  A266 );
 a52424a <=( A265  and  a52423a );
 a52427a <=( (not A300)  and  A299 );
 a52430a <=( A302  and  (not A301) );
 a52431a <=( a52430a  and  a52427a );
 a52432a <=( a52431a  and  a52424a );
 a52436a <=( (not A167)  and  A168 );
 a52437a <=( A169  and  a52436a );
 a52441a <=( A200  and  A199 );
 a52442a <=( A166  and  a52441a );
 a52443a <=( a52442a  and  a52437a );
 a52447a <=( A267  and  A266 );
 a52448a <=( (not A265)  and  a52447a );
 a52451a <=( A300  and  A268 );
 a52454a <=( A302  and  (not A301) );
 a52455a <=( a52454a  and  a52451a );
 a52456a <=( a52455a  and  a52448a );
 a52460a <=( (not A167)  and  A168 );
 a52461a <=( A169  and  a52460a );
 a52465a <=( A200  and  A199 );
 a52466a <=( A166  and  a52465a );
 a52467a <=( a52466a  and  a52461a );
 a52471a <=( A267  and  A266 );
 a52472a <=( (not A265)  and  a52471a );
 a52475a <=( A300  and  (not A269) );
 a52478a <=( A302  and  (not A301) );
 a52479a <=( a52478a  and  a52475a );
 a52480a <=( a52479a  and  a52472a );
 a52484a <=( (not A167)  and  A168 );
 a52485a <=( A169  and  a52484a );
 a52489a <=( A200  and  A199 );
 a52490a <=( A166  and  a52489a );
 a52491a <=( a52490a  and  a52485a );
 a52495a <=( (not A267)  and  A266 );
 a52496a <=( (not A265)  and  a52495a );
 a52499a <=( A269  and  (not A268) );
 a52502a <=( A301  and  (not A300) );
 a52503a <=( a52502a  and  a52499a );
 a52504a <=( a52503a  and  a52496a );
 a52508a <=( (not A167)  and  A168 );
 a52509a <=( A169  and  a52508a );
 a52513a <=( A200  and  A199 );
 a52514a <=( A166  and  a52513a );
 a52515a <=( a52514a  and  a52509a );
 a52519a <=( (not A267)  and  A266 );
 a52520a <=( (not A265)  and  a52519a );
 a52523a <=( A269  and  (not A268) );
 a52526a <=( (not A302)  and  (not A300) );
 a52527a <=( a52526a  and  a52523a );
 a52528a <=( a52527a  and  a52520a );
 a52532a <=( (not A167)  and  A168 );
 a52533a <=( A169  and  a52532a );
 a52537a <=( A200  and  A199 );
 a52538a <=( A166  and  a52537a );
 a52539a <=( a52538a  and  a52533a );
 a52543a <=( (not A267)  and  A266 );
 a52544a <=( (not A265)  and  a52543a );
 a52547a <=( A269  and  (not A268) );
 a52550a <=( A299  and  A298 );
 a52551a <=( a52550a  and  a52547a );
 a52552a <=( a52551a  and  a52544a );
 a52556a <=( (not A167)  and  A168 );
 a52557a <=( A169  and  a52556a );
 a52561a <=( A200  and  A199 );
 a52562a <=( A166  and  a52561a );
 a52563a <=( a52562a  and  a52557a );
 a52567a <=( (not A267)  and  A266 );
 a52568a <=( (not A265)  and  a52567a );
 a52571a <=( A269  and  (not A268) );
 a52574a <=( (not A299)  and  (not A298) );
 a52575a <=( a52574a  and  a52571a );
 a52576a <=( a52575a  and  a52568a );
 a52580a <=( (not A167)  and  A168 );
 a52581a <=( A169  and  a52580a );
 a52585a <=( A200  and  A199 );
 a52586a <=( A166  and  a52585a );
 a52587a <=( a52586a  and  a52581a );
 a52591a <=( A267  and  (not A266) );
 a52592a <=( A265  and  a52591a );
 a52595a <=( A300  and  A268 );
 a52598a <=( A302  and  (not A301) );
 a52599a <=( a52598a  and  a52595a );
 a52600a <=( a52599a  and  a52592a );
 a52604a <=( (not A167)  and  A168 );
 a52605a <=( A169  and  a52604a );
 a52609a <=( A200  and  A199 );
 a52610a <=( A166  and  a52609a );
 a52611a <=( a52610a  and  a52605a );
 a52615a <=( A267  and  (not A266) );
 a52616a <=( A265  and  a52615a );
 a52619a <=( A300  and  (not A269) );
 a52622a <=( A302  and  (not A301) );
 a52623a <=( a52622a  and  a52619a );
 a52624a <=( a52623a  and  a52616a );
 a52628a <=( (not A167)  and  A168 );
 a52629a <=( A169  and  a52628a );
 a52633a <=( A200  and  A199 );
 a52634a <=( A166  and  a52633a );
 a52635a <=( a52634a  and  a52629a );
 a52639a <=( (not A267)  and  (not A266) );
 a52640a <=( A265  and  a52639a );
 a52643a <=( A269  and  (not A268) );
 a52646a <=( A301  and  (not A300) );
 a52647a <=( a52646a  and  a52643a );
 a52648a <=( a52647a  and  a52640a );
 a52652a <=( (not A167)  and  A168 );
 a52653a <=( A169  and  a52652a );
 a52657a <=( A200  and  A199 );
 a52658a <=( A166  and  a52657a );
 a52659a <=( a52658a  and  a52653a );
 a52663a <=( (not A267)  and  (not A266) );
 a52664a <=( A265  and  a52663a );
 a52667a <=( A269  and  (not A268) );
 a52670a <=( (not A302)  and  (not A300) );
 a52671a <=( a52670a  and  a52667a );
 a52672a <=( a52671a  and  a52664a );
 a52676a <=( (not A167)  and  A168 );
 a52677a <=( A169  and  a52676a );
 a52681a <=( A200  and  A199 );
 a52682a <=( A166  and  a52681a );
 a52683a <=( a52682a  and  a52677a );
 a52687a <=( (not A267)  and  (not A266) );
 a52688a <=( A265  and  a52687a );
 a52691a <=( A269  and  (not A268) );
 a52694a <=( A299  and  A298 );
 a52695a <=( a52694a  and  a52691a );
 a52696a <=( a52695a  and  a52688a );
 a52700a <=( (not A167)  and  A168 );
 a52701a <=( A169  and  a52700a );
 a52705a <=( A200  and  A199 );
 a52706a <=( A166  and  a52705a );
 a52707a <=( a52706a  and  a52701a );
 a52711a <=( (not A267)  and  (not A266) );
 a52712a <=( A265  and  a52711a );
 a52715a <=( A269  and  (not A268) );
 a52718a <=( (not A299)  and  (not A298) );
 a52719a <=( a52718a  and  a52715a );
 a52720a <=( a52719a  and  a52712a );
 a52724a <=( (not A167)  and  A168 );
 a52725a <=( A169  and  a52724a );
 a52729a <=( A200  and  A199 );
 a52730a <=( A166  and  a52729a );
 a52731a <=( a52730a  and  a52725a );
 a52735a <=( A298  and  (not A266) );
 a52736a <=( (not A265)  and  a52735a );
 a52739a <=( (not A300)  and  (not A299) );
 a52742a <=( A302  and  (not A301) );
 a52743a <=( a52742a  and  a52739a );
 a52744a <=( a52743a  and  a52736a );
 a52748a <=( (not A167)  and  A168 );
 a52749a <=( A169  and  a52748a );
 a52753a <=( A200  and  A199 );
 a52754a <=( A166  and  a52753a );
 a52755a <=( a52754a  and  a52749a );
 a52759a <=( (not A298)  and  (not A266) );
 a52760a <=( (not A265)  and  a52759a );
 a52763a <=( (not A300)  and  A299 );
 a52766a <=( A302  and  (not A301) );
 a52767a <=( a52766a  and  a52763a );
 a52768a <=( a52767a  and  a52760a );
 a52772a <=( (not A167)  and  A168 );
 a52773a <=( A169  and  a52772a );
 a52777a <=( (not A200)  and  (not A199) );
 a52778a <=( A166  and  a52777a );
 a52779a <=( a52778a  and  a52773a );
 a52783a <=( A269  and  (not A268) );
 a52784a <=( A267  and  a52783a );
 a52787a <=( (not A299)  and  A298 );
 a52790a <=( A301  and  A300 );
 a52791a <=( a52790a  and  a52787a );
 a52792a <=( a52791a  and  a52784a );
 a52796a <=( (not A167)  and  A168 );
 a52797a <=( A169  and  a52796a );
 a52801a <=( (not A200)  and  (not A199) );
 a52802a <=( A166  and  a52801a );
 a52803a <=( a52802a  and  a52797a );
 a52807a <=( A269  and  (not A268) );
 a52808a <=( A267  and  a52807a );
 a52811a <=( (not A299)  and  A298 );
 a52814a <=( (not A302)  and  A300 );
 a52815a <=( a52814a  and  a52811a );
 a52816a <=( a52815a  and  a52808a );
 a52820a <=( (not A167)  and  A168 );
 a52821a <=( A169  and  a52820a );
 a52825a <=( (not A200)  and  (not A199) );
 a52826a <=( A166  and  a52825a );
 a52827a <=( a52826a  and  a52821a );
 a52831a <=( A269  and  (not A268) );
 a52832a <=( A267  and  a52831a );
 a52835a <=( A299  and  (not A298) );
 a52838a <=( A301  and  A300 );
 a52839a <=( a52838a  and  a52835a );
 a52840a <=( a52839a  and  a52832a );
 a52844a <=( (not A167)  and  A168 );
 a52845a <=( A169  and  a52844a );
 a52849a <=( (not A200)  and  (not A199) );
 a52850a <=( A166  and  a52849a );
 a52851a <=( a52850a  and  a52845a );
 a52855a <=( A269  and  (not A268) );
 a52856a <=( A267  and  a52855a );
 a52859a <=( A299  and  (not A298) );
 a52862a <=( (not A302)  and  A300 );
 a52863a <=( a52862a  and  a52859a );
 a52864a <=( a52863a  and  a52856a );
 a52868a <=( (not A167)  and  A168 );
 a52869a <=( A169  and  a52868a );
 a52873a <=( (not A200)  and  (not A199) );
 a52874a <=( A166  and  a52873a );
 a52875a <=( a52874a  and  a52869a );
 a52879a <=( A298  and  A268 );
 a52880a <=( (not A267)  and  a52879a );
 a52883a <=( (not A300)  and  (not A299) );
 a52886a <=( A302  and  (not A301) );
 a52887a <=( a52886a  and  a52883a );
 a52888a <=( a52887a  and  a52880a );
 a52892a <=( (not A167)  and  A168 );
 a52893a <=( A169  and  a52892a );
 a52897a <=( (not A200)  and  (not A199) );
 a52898a <=( A166  and  a52897a );
 a52899a <=( a52898a  and  a52893a );
 a52903a <=( (not A298)  and  A268 );
 a52904a <=( (not A267)  and  a52903a );
 a52907a <=( (not A300)  and  A299 );
 a52910a <=( A302  and  (not A301) );
 a52911a <=( a52910a  and  a52907a );
 a52912a <=( a52911a  and  a52904a );
 a52916a <=( (not A167)  and  A168 );
 a52917a <=( A169  and  a52916a );
 a52921a <=( (not A200)  and  (not A199) );
 a52922a <=( A166  and  a52921a );
 a52923a <=( a52922a  and  a52917a );
 a52927a <=( A298  and  (not A269) );
 a52928a <=( (not A267)  and  a52927a );
 a52931a <=( (not A300)  and  (not A299) );
 a52934a <=( A302  and  (not A301) );
 a52935a <=( a52934a  and  a52931a );
 a52936a <=( a52935a  and  a52928a );
 a52940a <=( (not A167)  and  A168 );
 a52941a <=( A169  and  a52940a );
 a52945a <=( (not A200)  and  (not A199) );
 a52946a <=( A166  and  a52945a );
 a52947a <=( a52946a  and  a52941a );
 a52951a <=( (not A298)  and  (not A269) );
 a52952a <=( (not A267)  and  a52951a );
 a52955a <=( (not A300)  and  A299 );
 a52958a <=( A302  and  (not A301) );
 a52959a <=( a52958a  and  a52955a );
 a52960a <=( a52959a  and  a52952a );
 a52964a <=( (not A167)  and  A168 );
 a52965a <=( A169  and  a52964a );
 a52969a <=( (not A200)  and  (not A199) );
 a52970a <=( A166  and  a52969a );
 a52971a <=( a52970a  and  a52965a );
 a52975a <=( A298  and  A266 );
 a52976a <=( A265  and  a52975a );
 a52979a <=( (not A300)  and  (not A299) );
 a52982a <=( A302  and  (not A301) );
 a52983a <=( a52982a  and  a52979a );
 a52984a <=( a52983a  and  a52976a );
 a52988a <=( (not A167)  and  A168 );
 a52989a <=( A169  and  a52988a );
 a52993a <=( (not A200)  and  (not A199) );
 a52994a <=( A166  and  a52993a );
 a52995a <=( a52994a  and  a52989a );
 a52999a <=( (not A298)  and  A266 );
 a53000a <=( A265  and  a52999a );
 a53003a <=( (not A300)  and  A299 );
 a53006a <=( A302  and  (not A301) );
 a53007a <=( a53006a  and  a53003a );
 a53008a <=( a53007a  and  a53000a );
 a53012a <=( (not A167)  and  A168 );
 a53013a <=( A169  and  a53012a );
 a53017a <=( (not A200)  and  (not A199) );
 a53018a <=( A166  and  a53017a );
 a53019a <=( a53018a  and  a53013a );
 a53023a <=( A267  and  A266 );
 a53024a <=( (not A265)  and  a53023a );
 a53027a <=( A300  and  A268 );
 a53030a <=( A302  and  (not A301) );
 a53031a <=( a53030a  and  a53027a );
 a53032a <=( a53031a  and  a53024a );
 a53036a <=( (not A167)  and  A168 );
 a53037a <=( A169  and  a53036a );
 a53041a <=( (not A200)  and  (not A199) );
 a53042a <=( A166  and  a53041a );
 a53043a <=( a53042a  and  a53037a );
 a53047a <=( A267  and  A266 );
 a53048a <=( (not A265)  and  a53047a );
 a53051a <=( A300  and  (not A269) );
 a53054a <=( A302  and  (not A301) );
 a53055a <=( a53054a  and  a53051a );
 a53056a <=( a53055a  and  a53048a );
 a53060a <=( (not A167)  and  A168 );
 a53061a <=( A169  and  a53060a );
 a53065a <=( (not A200)  and  (not A199) );
 a53066a <=( A166  and  a53065a );
 a53067a <=( a53066a  and  a53061a );
 a53071a <=( (not A267)  and  A266 );
 a53072a <=( (not A265)  and  a53071a );
 a53075a <=( A269  and  (not A268) );
 a53078a <=( A301  and  (not A300) );
 a53079a <=( a53078a  and  a53075a );
 a53080a <=( a53079a  and  a53072a );
 a53084a <=( (not A167)  and  A168 );
 a53085a <=( A169  and  a53084a );
 a53089a <=( (not A200)  and  (not A199) );
 a53090a <=( A166  and  a53089a );
 a53091a <=( a53090a  and  a53085a );
 a53095a <=( (not A267)  and  A266 );
 a53096a <=( (not A265)  and  a53095a );
 a53099a <=( A269  and  (not A268) );
 a53102a <=( (not A302)  and  (not A300) );
 a53103a <=( a53102a  and  a53099a );
 a53104a <=( a53103a  and  a53096a );
 a53108a <=( (not A167)  and  A168 );
 a53109a <=( A169  and  a53108a );
 a53113a <=( (not A200)  and  (not A199) );
 a53114a <=( A166  and  a53113a );
 a53115a <=( a53114a  and  a53109a );
 a53119a <=( (not A267)  and  A266 );
 a53120a <=( (not A265)  and  a53119a );
 a53123a <=( A269  and  (not A268) );
 a53126a <=( A299  and  A298 );
 a53127a <=( a53126a  and  a53123a );
 a53128a <=( a53127a  and  a53120a );
 a53132a <=( (not A167)  and  A168 );
 a53133a <=( A169  and  a53132a );
 a53137a <=( (not A200)  and  (not A199) );
 a53138a <=( A166  and  a53137a );
 a53139a <=( a53138a  and  a53133a );
 a53143a <=( (not A267)  and  A266 );
 a53144a <=( (not A265)  and  a53143a );
 a53147a <=( A269  and  (not A268) );
 a53150a <=( (not A299)  and  (not A298) );
 a53151a <=( a53150a  and  a53147a );
 a53152a <=( a53151a  and  a53144a );
 a53156a <=( (not A167)  and  A168 );
 a53157a <=( A169  and  a53156a );
 a53161a <=( (not A200)  and  (not A199) );
 a53162a <=( A166  and  a53161a );
 a53163a <=( a53162a  and  a53157a );
 a53167a <=( A267  and  (not A266) );
 a53168a <=( A265  and  a53167a );
 a53171a <=( A300  and  A268 );
 a53174a <=( A302  and  (not A301) );
 a53175a <=( a53174a  and  a53171a );
 a53176a <=( a53175a  and  a53168a );
 a53180a <=( (not A167)  and  A168 );
 a53181a <=( A169  and  a53180a );
 a53185a <=( (not A200)  and  (not A199) );
 a53186a <=( A166  and  a53185a );
 a53187a <=( a53186a  and  a53181a );
 a53191a <=( A267  and  (not A266) );
 a53192a <=( A265  and  a53191a );
 a53195a <=( A300  and  (not A269) );
 a53198a <=( A302  and  (not A301) );
 a53199a <=( a53198a  and  a53195a );
 a53200a <=( a53199a  and  a53192a );
 a53204a <=( (not A167)  and  A168 );
 a53205a <=( A169  and  a53204a );
 a53209a <=( (not A200)  and  (not A199) );
 a53210a <=( A166  and  a53209a );
 a53211a <=( a53210a  and  a53205a );
 a53215a <=( (not A267)  and  (not A266) );
 a53216a <=( A265  and  a53215a );
 a53219a <=( A269  and  (not A268) );
 a53222a <=( A301  and  (not A300) );
 a53223a <=( a53222a  and  a53219a );
 a53224a <=( a53223a  and  a53216a );
 a53228a <=( (not A167)  and  A168 );
 a53229a <=( A169  and  a53228a );
 a53233a <=( (not A200)  and  (not A199) );
 a53234a <=( A166  and  a53233a );
 a53235a <=( a53234a  and  a53229a );
 a53239a <=( (not A267)  and  (not A266) );
 a53240a <=( A265  and  a53239a );
 a53243a <=( A269  and  (not A268) );
 a53246a <=( (not A302)  and  (not A300) );
 a53247a <=( a53246a  and  a53243a );
 a53248a <=( a53247a  and  a53240a );
 a53252a <=( (not A167)  and  A168 );
 a53253a <=( A169  and  a53252a );
 a53257a <=( (not A200)  and  (not A199) );
 a53258a <=( A166  and  a53257a );
 a53259a <=( a53258a  and  a53253a );
 a53263a <=( (not A267)  and  (not A266) );
 a53264a <=( A265  and  a53263a );
 a53267a <=( A269  and  (not A268) );
 a53270a <=( A299  and  A298 );
 a53271a <=( a53270a  and  a53267a );
 a53272a <=( a53271a  and  a53264a );
 a53276a <=( (not A167)  and  A168 );
 a53277a <=( A169  and  a53276a );
 a53281a <=( (not A200)  and  (not A199) );
 a53282a <=( A166  and  a53281a );
 a53283a <=( a53282a  and  a53277a );
 a53287a <=( (not A267)  and  (not A266) );
 a53288a <=( A265  and  a53287a );
 a53291a <=( A269  and  (not A268) );
 a53294a <=( (not A299)  and  (not A298) );
 a53295a <=( a53294a  and  a53291a );
 a53296a <=( a53295a  and  a53288a );
 a53300a <=( (not A167)  and  A168 );
 a53301a <=( A169  and  a53300a );
 a53305a <=( (not A200)  and  (not A199) );
 a53306a <=( A166  and  a53305a );
 a53307a <=( a53306a  and  a53301a );
 a53311a <=( A298  and  (not A266) );
 a53312a <=( (not A265)  and  a53311a );
 a53315a <=( (not A300)  and  (not A299) );
 a53318a <=( A302  and  (not A301) );
 a53319a <=( a53318a  and  a53315a );
 a53320a <=( a53319a  and  a53312a );
 a53324a <=( (not A167)  and  A168 );
 a53325a <=( A169  and  a53324a );
 a53329a <=( (not A200)  and  (not A199) );
 a53330a <=( A166  and  a53329a );
 a53331a <=( a53330a  and  a53325a );
 a53335a <=( (not A298)  and  (not A266) );
 a53336a <=( (not A265)  and  a53335a );
 a53339a <=( (not A300)  and  A299 );
 a53342a <=( A302  and  (not A301) );
 a53343a <=( a53342a  and  a53339a );
 a53344a <=( a53343a  and  a53336a );
 a53348a <=( (not A199)  and  (not A168) );
 a53349a <=( A169  and  a53348a );
 a53353a <=( (not A202)  and  (not A201) );
 a53354a <=( A200  and  a53353a );
 a53355a <=( a53354a  and  a53349a );
 a53359a <=( (not A268)  and  A267 );
 a53360a <=( A203  and  a53359a );
 a53363a <=( A300  and  A269 );
 a53366a <=( A302  and  (not A301) );
 a53367a <=( a53366a  and  a53363a );
 a53368a <=( a53367a  and  a53360a );
 a53372a <=( A199  and  (not A168) );
 a53373a <=( A169  and  a53372a );
 a53377a <=( (not A202)  and  (not A201) );
 a53378a <=( (not A200)  and  a53377a );
 a53379a <=( a53378a  and  a53373a );
 a53383a <=( (not A268)  and  A267 );
 a53384a <=( A203  and  a53383a );
 a53387a <=( A300  and  A269 );
 a53390a <=( A302  and  (not A301) );
 a53391a <=( a53390a  and  a53387a );
 a53392a <=( a53391a  and  a53384a );
 a53396a <=( A168  and  (not A169) );
 a53397a <=( (not A170)  and  a53396a );
 a53401a <=( (not A234)  and  A233 );
 a53402a <=( (not A232)  and  a53401a );
 a53403a <=( a53402a  and  a53397a );
 a53407a <=( (not A265)  and  A236 );
 a53408a <=( (not A235)  and  a53407a );
 a53411a <=( (not A267)  and  A266 );
 a53414a <=( A269  and  (not A268) );
 a53415a <=( a53414a  and  a53411a );
 a53416a <=( a53415a  and  a53408a );
 a53420a <=( A168  and  (not A169) );
 a53421a <=( (not A170)  and  a53420a );
 a53425a <=( (not A234)  and  A233 );
 a53426a <=( (not A232)  and  a53425a );
 a53427a <=( a53426a  and  a53421a );
 a53431a <=( A265  and  A236 );
 a53432a <=( (not A235)  and  a53431a );
 a53435a <=( (not A267)  and  (not A266) );
 a53438a <=( A269  and  (not A268) );
 a53439a <=( a53438a  and  a53435a );
 a53440a <=( a53439a  and  a53432a );
 a53444a <=( A168  and  (not A169) );
 a53445a <=( (not A170)  and  a53444a );
 a53449a <=( (not A234)  and  (not A233) );
 a53450a <=( A232  and  a53449a );
 a53451a <=( a53450a  and  a53445a );
 a53455a <=( (not A265)  and  A236 );
 a53456a <=( (not A235)  and  a53455a );
 a53459a <=( (not A267)  and  A266 );
 a53462a <=( A269  and  (not A268) );
 a53463a <=( a53462a  and  a53459a );
 a53464a <=( a53463a  and  a53456a );
 a53468a <=( A168  and  (not A169) );
 a53469a <=( (not A170)  and  a53468a );
 a53473a <=( (not A234)  and  (not A233) );
 a53474a <=( A232  and  a53473a );
 a53475a <=( a53474a  and  a53469a );
 a53479a <=( A265  and  A236 );
 a53480a <=( (not A235)  and  a53479a );
 a53483a <=( (not A267)  and  (not A266) );
 a53486a <=( A269  and  (not A268) );
 a53487a <=( a53486a  and  a53483a );
 a53488a <=( a53487a  and  a53480a );
 a53492a <=( A168  and  (not A169) );
 a53493a <=( (not A170)  and  a53492a );
 a53497a <=( A201  and  A200 );
 a53498a <=( (not A199)  and  a53497a );
 a53499a <=( a53498a  and  a53493a );
 a53503a <=( (not A268)  and  A267 );
 a53504a <=( A202  and  a53503a );
 a53507a <=( A300  and  A269 );
 a53510a <=( A302  and  (not A301) );
 a53511a <=( a53510a  and  a53507a );
 a53512a <=( a53511a  and  a53504a );
 a53516a <=( A168  and  (not A169) );
 a53517a <=( (not A170)  and  a53516a );
 a53521a <=( A201  and  A200 );
 a53522a <=( (not A199)  and  a53521a );
 a53523a <=( a53522a  and  a53517a );
 a53527a <=( (not A268)  and  A267 );
 a53528a <=( (not A203)  and  a53527a );
 a53531a <=( A300  and  A269 );
 a53534a <=( A302  and  (not A301) );
 a53535a <=( a53534a  and  a53531a );
 a53536a <=( a53535a  and  a53528a );
 a53540a <=( A168  and  (not A169) );
 a53541a <=( (not A170)  and  a53540a );
 a53545a <=( (not A201)  and  A200 );
 a53546a <=( (not A199)  and  a53545a );
 a53547a <=( a53546a  and  a53541a );
 a53551a <=( A267  and  A203 );
 a53552a <=( (not A202)  and  a53551a );
 a53555a <=( A269  and  (not A268) );
 a53558a <=( A301  and  (not A300) );
 a53559a <=( a53558a  and  a53555a );
 a53560a <=( a53559a  and  a53552a );
 a53564a <=( A168  and  (not A169) );
 a53565a <=( (not A170)  and  a53564a );
 a53569a <=( (not A201)  and  A200 );
 a53570a <=( (not A199)  and  a53569a );
 a53571a <=( a53570a  and  a53565a );
 a53575a <=( A267  and  A203 );
 a53576a <=( (not A202)  and  a53575a );
 a53579a <=( A269  and  (not A268) );
 a53582a <=( (not A302)  and  (not A300) );
 a53583a <=( a53582a  and  a53579a );
 a53584a <=( a53583a  and  a53576a );
 a53588a <=( A168  and  (not A169) );
 a53589a <=( (not A170)  and  a53588a );
 a53593a <=( (not A201)  and  A200 );
 a53594a <=( (not A199)  and  a53593a );
 a53595a <=( a53594a  and  a53589a );
 a53599a <=( A267  and  A203 );
 a53600a <=( (not A202)  and  a53599a );
 a53603a <=( A269  and  (not A268) );
 a53606a <=( A299  and  A298 );
 a53607a <=( a53606a  and  a53603a );
 a53608a <=( a53607a  and  a53600a );
 a53612a <=( A168  and  (not A169) );
 a53613a <=( (not A170)  and  a53612a );
 a53617a <=( (not A201)  and  A200 );
 a53618a <=( (not A199)  and  a53617a );
 a53619a <=( a53618a  and  a53613a );
 a53623a <=( A267  and  A203 );
 a53624a <=( (not A202)  and  a53623a );
 a53627a <=( A269  and  (not A268) );
 a53630a <=( (not A299)  and  (not A298) );
 a53631a <=( a53630a  and  a53627a );
 a53632a <=( a53631a  and  a53624a );
 a53636a <=( A168  and  (not A169) );
 a53637a <=( (not A170)  and  a53636a );
 a53641a <=( (not A201)  and  A200 );
 a53642a <=( (not A199)  and  a53641a );
 a53643a <=( a53642a  and  a53637a );
 a53647a <=( (not A267)  and  A203 );
 a53648a <=( (not A202)  and  a53647a );
 a53651a <=( A300  and  A268 );
 a53654a <=( A302  and  (not A301) );
 a53655a <=( a53654a  and  a53651a );
 a53656a <=( a53655a  and  a53648a );
 a53660a <=( A168  and  (not A169) );
 a53661a <=( (not A170)  and  a53660a );
 a53665a <=( (not A201)  and  A200 );
 a53666a <=( (not A199)  and  a53665a );
 a53667a <=( a53666a  and  a53661a );
 a53671a <=( (not A267)  and  A203 );
 a53672a <=( (not A202)  and  a53671a );
 a53675a <=( A300  and  (not A269) );
 a53678a <=( A302  and  (not A301) );
 a53679a <=( a53678a  and  a53675a );
 a53680a <=( a53679a  and  a53672a );
 a53684a <=( A168  and  (not A169) );
 a53685a <=( (not A170)  and  a53684a );
 a53689a <=( (not A201)  and  A200 );
 a53690a <=( (not A199)  and  a53689a );
 a53691a <=( a53690a  and  a53685a );
 a53695a <=( A265  and  A203 );
 a53696a <=( (not A202)  and  a53695a );
 a53699a <=( A300  and  A266 );
 a53702a <=( A302  and  (not A301) );
 a53703a <=( a53702a  and  a53699a );
 a53704a <=( a53703a  and  a53696a );
 a53708a <=( A168  and  (not A169) );
 a53709a <=( (not A170)  and  a53708a );
 a53713a <=( (not A201)  and  A200 );
 a53714a <=( (not A199)  and  a53713a );
 a53715a <=( a53714a  and  a53709a );
 a53719a <=( (not A265)  and  A203 );
 a53720a <=( (not A202)  and  a53719a );
 a53723a <=( A300  and  (not A266) );
 a53726a <=( A302  and  (not A301) );
 a53727a <=( a53726a  and  a53723a );
 a53728a <=( a53727a  and  a53720a );
 a53732a <=( A168  and  (not A169) );
 a53733a <=( (not A170)  and  a53732a );
 a53737a <=( A201  and  (not A200) );
 a53738a <=( A199  and  a53737a );
 a53739a <=( a53738a  and  a53733a );
 a53743a <=( (not A268)  and  A267 );
 a53744a <=( A202  and  a53743a );
 a53747a <=( A300  and  A269 );
 a53750a <=( A302  and  (not A301) );
 a53751a <=( a53750a  and  a53747a );
 a53752a <=( a53751a  and  a53744a );
 a53756a <=( A168  and  (not A169) );
 a53757a <=( (not A170)  and  a53756a );
 a53761a <=( A201  and  (not A200) );
 a53762a <=( A199  and  a53761a );
 a53763a <=( a53762a  and  a53757a );
 a53767a <=( (not A268)  and  A267 );
 a53768a <=( (not A203)  and  a53767a );
 a53771a <=( A300  and  A269 );
 a53774a <=( A302  and  (not A301) );
 a53775a <=( a53774a  and  a53771a );
 a53776a <=( a53775a  and  a53768a );
 a53780a <=( A168  and  (not A169) );
 a53781a <=( (not A170)  and  a53780a );
 a53785a <=( (not A201)  and  (not A200) );
 a53786a <=( A199  and  a53785a );
 a53787a <=( a53786a  and  a53781a );
 a53791a <=( A267  and  A203 );
 a53792a <=( (not A202)  and  a53791a );
 a53795a <=( A269  and  (not A268) );
 a53798a <=( A301  and  (not A300) );
 a53799a <=( a53798a  and  a53795a );
 a53800a <=( a53799a  and  a53792a );
 a53804a <=( A168  and  (not A169) );
 a53805a <=( (not A170)  and  a53804a );
 a53809a <=( (not A201)  and  (not A200) );
 a53810a <=( A199  and  a53809a );
 a53811a <=( a53810a  and  a53805a );
 a53815a <=( A267  and  A203 );
 a53816a <=( (not A202)  and  a53815a );
 a53819a <=( A269  and  (not A268) );
 a53822a <=( (not A302)  and  (not A300) );
 a53823a <=( a53822a  and  a53819a );
 a53824a <=( a53823a  and  a53816a );
 a53828a <=( A168  and  (not A169) );
 a53829a <=( (not A170)  and  a53828a );
 a53833a <=( (not A201)  and  (not A200) );
 a53834a <=( A199  and  a53833a );
 a53835a <=( a53834a  and  a53829a );
 a53839a <=( A267  and  A203 );
 a53840a <=( (not A202)  and  a53839a );
 a53843a <=( A269  and  (not A268) );
 a53846a <=( A299  and  A298 );
 a53847a <=( a53846a  and  a53843a );
 a53848a <=( a53847a  and  a53840a );
 a53852a <=( A168  and  (not A169) );
 a53853a <=( (not A170)  and  a53852a );
 a53857a <=( (not A201)  and  (not A200) );
 a53858a <=( A199  and  a53857a );
 a53859a <=( a53858a  and  a53853a );
 a53863a <=( A267  and  A203 );
 a53864a <=( (not A202)  and  a53863a );
 a53867a <=( A269  and  (not A268) );
 a53870a <=( (not A299)  and  (not A298) );
 a53871a <=( a53870a  and  a53867a );
 a53872a <=( a53871a  and  a53864a );
 a53876a <=( A168  and  (not A169) );
 a53877a <=( (not A170)  and  a53876a );
 a53881a <=( (not A201)  and  (not A200) );
 a53882a <=( A199  and  a53881a );
 a53883a <=( a53882a  and  a53877a );
 a53887a <=( (not A267)  and  A203 );
 a53888a <=( (not A202)  and  a53887a );
 a53891a <=( A300  and  A268 );
 a53894a <=( A302  and  (not A301) );
 a53895a <=( a53894a  and  a53891a );
 a53896a <=( a53895a  and  a53888a );
 a53900a <=( A168  and  (not A169) );
 a53901a <=( (not A170)  and  a53900a );
 a53905a <=( (not A201)  and  (not A200) );
 a53906a <=( A199  and  a53905a );
 a53907a <=( a53906a  and  a53901a );
 a53911a <=( (not A267)  and  A203 );
 a53912a <=( (not A202)  and  a53911a );
 a53915a <=( A300  and  (not A269) );
 a53918a <=( A302  and  (not A301) );
 a53919a <=( a53918a  and  a53915a );
 a53920a <=( a53919a  and  a53912a );
 a53924a <=( A168  and  (not A169) );
 a53925a <=( (not A170)  and  a53924a );
 a53929a <=( (not A201)  and  (not A200) );
 a53930a <=( A199  and  a53929a );
 a53931a <=( a53930a  and  a53925a );
 a53935a <=( A265  and  A203 );
 a53936a <=( (not A202)  and  a53935a );
 a53939a <=( A300  and  A266 );
 a53942a <=( A302  and  (not A301) );
 a53943a <=( a53942a  and  a53939a );
 a53944a <=( a53943a  and  a53936a );
 a53948a <=( A168  and  (not A169) );
 a53949a <=( (not A170)  and  a53948a );
 a53953a <=( (not A201)  and  (not A200) );
 a53954a <=( A199  and  a53953a );
 a53955a <=( a53954a  and  a53949a );
 a53959a <=( (not A265)  and  A203 );
 a53960a <=( (not A202)  and  a53959a );
 a53963a <=( A300  and  (not A266) );
 a53966a <=( A302  and  (not A301) );
 a53967a <=( a53966a  and  a53963a );
 a53968a <=( a53967a  and  a53960a );
 a53972a <=( (not A168)  and  (not A169) );
 a53973a <=( (not A170)  and  a53972a );
 a53977a <=( (not A201)  and  (not A166) );
 a53978a <=( A167  and  a53977a );
 a53979a <=( a53978a  and  a53973a );
 a53983a <=( A268  and  (not A267) );
 a53984a <=( A202  and  a53983a );
 a53987a <=( (not A299)  and  A298 );
 a53990a <=( A301  and  A300 );
 a53991a <=( a53990a  and  a53987a );
 a53992a <=( a53991a  and  a53984a );
 a53996a <=( (not A168)  and  (not A169) );
 a53997a <=( (not A170)  and  a53996a );
 a54001a <=( (not A201)  and  (not A166) );
 a54002a <=( A167  and  a54001a );
 a54003a <=( a54002a  and  a53997a );
 a54007a <=( A268  and  (not A267) );
 a54008a <=( A202  and  a54007a );
 a54011a <=( (not A299)  and  A298 );
 a54014a <=( (not A302)  and  A300 );
 a54015a <=( a54014a  and  a54011a );
 a54016a <=( a54015a  and  a54008a );
 a54020a <=( (not A168)  and  (not A169) );
 a54021a <=( (not A170)  and  a54020a );
 a54025a <=( (not A201)  and  (not A166) );
 a54026a <=( A167  and  a54025a );
 a54027a <=( a54026a  and  a54021a );
 a54031a <=( A268  and  (not A267) );
 a54032a <=( A202  and  a54031a );
 a54035a <=( A299  and  (not A298) );
 a54038a <=( A301  and  A300 );
 a54039a <=( a54038a  and  a54035a );
 a54040a <=( a54039a  and  a54032a );
 a54044a <=( (not A168)  and  (not A169) );
 a54045a <=( (not A170)  and  a54044a );
 a54049a <=( (not A201)  and  (not A166) );
 a54050a <=( A167  and  a54049a );
 a54051a <=( a54050a  and  a54045a );
 a54055a <=( A268  and  (not A267) );
 a54056a <=( A202  and  a54055a );
 a54059a <=( A299  and  (not A298) );
 a54062a <=( (not A302)  and  A300 );
 a54063a <=( a54062a  and  a54059a );
 a54064a <=( a54063a  and  a54056a );
 a54068a <=( (not A168)  and  (not A169) );
 a54069a <=( (not A170)  and  a54068a );
 a54073a <=( (not A201)  and  (not A166) );
 a54074a <=( A167  and  a54073a );
 a54075a <=( a54074a  and  a54069a );
 a54079a <=( (not A269)  and  (not A267) );
 a54080a <=( A202  and  a54079a );
 a54083a <=( (not A299)  and  A298 );
 a54086a <=( A301  and  A300 );
 a54087a <=( a54086a  and  a54083a );
 a54088a <=( a54087a  and  a54080a );
 a54092a <=( (not A168)  and  (not A169) );
 a54093a <=( (not A170)  and  a54092a );
 a54097a <=( (not A201)  and  (not A166) );
 a54098a <=( A167  and  a54097a );
 a54099a <=( a54098a  and  a54093a );
 a54103a <=( (not A269)  and  (not A267) );
 a54104a <=( A202  and  a54103a );
 a54107a <=( (not A299)  and  A298 );
 a54110a <=( (not A302)  and  A300 );
 a54111a <=( a54110a  and  a54107a );
 a54112a <=( a54111a  and  a54104a );
 a54116a <=( (not A168)  and  (not A169) );
 a54117a <=( (not A170)  and  a54116a );
 a54121a <=( (not A201)  and  (not A166) );
 a54122a <=( A167  and  a54121a );
 a54123a <=( a54122a  and  a54117a );
 a54127a <=( (not A269)  and  (not A267) );
 a54128a <=( A202  and  a54127a );
 a54131a <=( A299  and  (not A298) );
 a54134a <=( A301  and  A300 );
 a54135a <=( a54134a  and  a54131a );
 a54136a <=( a54135a  and  a54128a );
 a54140a <=( (not A168)  and  (not A169) );
 a54141a <=( (not A170)  and  a54140a );
 a54145a <=( (not A201)  and  (not A166) );
 a54146a <=( A167  and  a54145a );
 a54147a <=( a54146a  and  a54141a );
 a54151a <=( (not A269)  and  (not A267) );
 a54152a <=( A202  and  a54151a );
 a54155a <=( A299  and  (not A298) );
 a54158a <=( (not A302)  and  A300 );
 a54159a <=( a54158a  and  a54155a );
 a54160a <=( a54159a  and  a54152a );
 a54164a <=( (not A168)  and  (not A169) );
 a54165a <=( (not A170)  and  a54164a );
 a54169a <=( (not A201)  and  (not A166) );
 a54170a <=( A167  and  a54169a );
 a54171a <=( a54170a  and  a54165a );
 a54175a <=( A266  and  A265 );
 a54176a <=( A202  and  a54175a );
 a54179a <=( (not A299)  and  A298 );
 a54182a <=( A301  and  A300 );
 a54183a <=( a54182a  and  a54179a );
 a54184a <=( a54183a  and  a54176a );
 a54188a <=( (not A168)  and  (not A169) );
 a54189a <=( (not A170)  and  a54188a );
 a54193a <=( (not A201)  and  (not A166) );
 a54194a <=( A167  and  a54193a );
 a54195a <=( a54194a  and  a54189a );
 a54199a <=( A266  and  A265 );
 a54200a <=( A202  and  a54199a );
 a54203a <=( (not A299)  and  A298 );
 a54206a <=( (not A302)  and  A300 );
 a54207a <=( a54206a  and  a54203a );
 a54208a <=( a54207a  and  a54200a );
 a54212a <=( (not A168)  and  (not A169) );
 a54213a <=( (not A170)  and  a54212a );
 a54217a <=( (not A201)  and  (not A166) );
 a54218a <=( A167  and  a54217a );
 a54219a <=( a54218a  and  a54213a );
 a54223a <=( A266  and  A265 );
 a54224a <=( A202  and  a54223a );
 a54227a <=( A299  and  (not A298) );
 a54230a <=( A301  and  A300 );
 a54231a <=( a54230a  and  a54227a );
 a54232a <=( a54231a  and  a54224a );
 a54236a <=( (not A168)  and  (not A169) );
 a54237a <=( (not A170)  and  a54236a );
 a54241a <=( (not A201)  and  (not A166) );
 a54242a <=( A167  and  a54241a );
 a54243a <=( a54242a  and  a54237a );
 a54247a <=( A266  and  A265 );
 a54248a <=( A202  and  a54247a );
 a54251a <=( A299  and  (not A298) );
 a54254a <=( (not A302)  and  A300 );
 a54255a <=( a54254a  and  a54251a );
 a54256a <=( a54255a  and  a54248a );
 a54260a <=( (not A168)  and  (not A169) );
 a54261a <=( (not A170)  and  a54260a );
 a54265a <=( (not A201)  and  (not A166) );
 a54266a <=( A167  and  a54265a );
 a54267a <=( a54266a  and  a54261a );
 a54271a <=( A266  and  (not A265) );
 a54272a <=( A202  and  a54271a );
 a54275a <=( A268  and  A267 );
 a54278a <=( A301  and  (not A300) );
 a54279a <=( a54278a  and  a54275a );
 a54280a <=( a54279a  and  a54272a );
 a54284a <=( (not A168)  and  (not A169) );
 a54285a <=( (not A170)  and  a54284a );
 a54289a <=( (not A201)  and  (not A166) );
 a54290a <=( A167  and  a54289a );
 a54291a <=( a54290a  and  a54285a );
 a54295a <=( A266  and  (not A265) );
 a54296a <=( A202  and  a54295a );
 a54299a <=( A268  and  A267 );
 a54302a <=( (not A302)  and  (not A300) );
 a54303a <=( a54302a  and  a54299a );
 a54304a <=( a54303a  and  a54296a );
 a54308a <=( (not A168)  and  (not A169) );
 a54309a <=( (not A170)  and  a54308a );
 a54313a <=( (not A201)  and  (not A166) );
 a54314a <=( A167  and  a54313a );
 a54315a <=( a54314a  and  a54309a );
 a54319a <=( A266  and  (not A265) );
 a54320a <=( A202  and  a54319a );
 a54323a <=( A268  and  A267 );
 a54326a <=( A299  and  A298 );
 a54327a <=( a54326a  and  a54323a );
 a54328a <=( a54327a  and  a54320a );
 a54332a <=( (not A168)  and  (not A169) );
 a54333a <=( (not A170)  and  a54332a );
 a54337a <=( (not A201)  and  (not A166) );
 a54338a <=( A167  and  a54337a );
 a54339a <=( a54338a  and  a54333a );
 a54343a <=( A266  and  (not A265) );
 a54344a <=( A202  and  a54343a );
 a54347a <=( A268  and  A267 );
 a54350a <=( (not A299)  and  (not A298) );
 a54351a <=( a54350a  and  a54347a );
 a54352a <=( a54351a  and  a54344a );
 a54356a <=( (not A168)  and  (not A169) );
 a54357a <=( (not A170)  and  a54356a );
 a54361a <=( (not A201)  and  (not A166) );
 a54362a <=( A167  and  a54361a );
 a54363a <=( a54362a  and  a54357a );
 a54367a <=( A266  and  (not A265) );
 a54368a <=( A202  and  a54367a );
 a54371a <=( (not A269)  and  A267 );
 a54374a <=( A301  and  (not A300) );
 a54375a <=( a54374a  and  a54371a );
 a54376a <=( a54375a  and  a54368a );
 a54380a <=( (not A168)  and  (not A169) );
 a54381a <=( (not A170)  and  a54380a );
 a54385a <=( (not A201)  and  (not A166) );
 a54386a <=( A167  and  a54385a );
 a54387a <=( a54386a  and  a54381a );
 a54391a <=( A266  and  (not A265) );
 a54392a <=( A202  and  a54391a );
 a54395a <=( (not A269)  and  A267 );
 a54398a <=( (not A302)  and  (not A300) );
 a54399a <=( a54398a  and  a54395a );
 a54400a <=( a54399a  and  a54392a );
 a54404a <=( (not A168)  and  (not A169) );
 a54405a <=( (not A170)  and  a54404a );
 a54409a <=( (not A201)  and  (not A166) );
 a54410a <=( A167  and  a54409a );
 a54411a <=( a54410a  and  a54405a );
 a54415a <=( A266  and  (not A265) );
 a54416a <=( A202  and  a54415a );
 a54419a <=( (not A269)  and  A267 );
 a54422a <=( A299  and  A298 );
 a54423a <=( a54422a  and  a54419a );
 a54424a <=( a54423a  and  a54416a );
 a54428a <=( (not A168)  and  (not A169) );
 a54429a <=( (not A170)  and  a54428a );
 a54433a <=( (not A201)  and  (not A166) );
 a54434a <=( A167  and  a54433a );
 a54435a <=( a54434a  and  a54429a );
 a54439a <=( A266  and  (not A265) );
 a54440a <=( A202  and  a54439a );
 a54443a <=( (not A269)  and  A267 );
 a54446a <=( (not A299)  and  (not A298) );
 a54447a <=( a54446a  and  a54443a );
 a54448a <=( a54447a  and  a54440a );
 a54452a <=( (not A168)  and  (not A169) );
 a54453a <=( (not A170)  and  a54452a );
 a54457a <=( (not A201)  and  (not A166) );
 a54458a <=( A167  and  a54457a );
 a54459a <=( a54458a  and  a54453a );
 a54463a <=( (not A266)  and  A265 );
 a54464a <=( A202  and  a54463a );
 a54467a <=( A268  and  A267 );
 a54470a <=( A301  and  (not A300) );
 a54471a <=( a54470a  and  a54467a );
 a54472a <=( a54471a  and  a54464a );
 a54476a <=( (not A168)  and  (not A169) );
 a54477a <=( (not A170)  and  a54476a );
 a54481a <=( (not A201)  and  (not A166) );
 a54482a <=( A167  and  a54481a );
 a54483a <=( a54482a  and  a54477a );
 a54487a <=( (not A266)  and  A265 );
 a54488a <=( A202  and  a54487a );
 a54491a <=( A268  and  A267 );
 a54494a <=( (not A302)  and  (not A300) );
 a54495a <=( a54494a  and  a54491a );
 a54496a <=( a54495a  and  a54488a );
 a54500a <=( (not A168)  and  (not A169) );
 a54501a <=( (not A170)  and  a54500a );
 a54505a <=( (not A201)  and  (not A166) );
 a54506a <=( A167  and  a54505a );
 a54507a <=( a54506a  and  a54501a );
 a54511a <=( (not A266)  and  A265 );
 a54512a <=( A202  and  a54511a );
 a54515a <=( A268  and  A267 );
 a54518a <=( A299  and  A298 );
 a54519a <=( a54518a  and  a54515a );
 a54520a <=( a54519a  and  a54512a );
 a54524a <=( (not A168)  and  (not A169) );
 a54525a <=( (not A170)  and  a54524a );
 a54529a <=( (not A201)  and  (not A166) );
 a54530a <=( A167  and  a54529a );
 a54531a <=( a54530a  and  a54525a );
 a54535a <=( (not A266)  and  A265 );
 a54536a <=( A202  and  a54535a );
 a54539a <=( A268  and  A267 );
 a54542a <=( (not A299)  and  (not A298) );
 a54543a <=( a54542a  and  a54539a );
 a54544a <=( a54543a  and  a54536a );
 a54548a <=( (not A168)  and  (not A169) );
 a54549a <=( (not A170)  and  a54548a );
 a54553a <=( (not A201)  and  (not A166) );
 a54554a <=( A167  and  a54553a );
 a54555a <=( a54554a  and  a54549a );
 a54559a <=( (not A266)  and  A265 );
 a54560a <=( A202  and  a54559a );
 a54563a <=( (not A269)  and  A267 );
 a54566a <=( A301  and  (not A300) );
 a54567a <=( a54566a  and  a54563a );
 a54568a <=( a54567a  and  a54560a );
 a54572a <=( (not A168)  and  (not A169) );
 a54573a <=( (not A170)  and  a54572a );
 a54577a <=( (not A201)  and  (not A166) );
 a54578a <=( A167  and  a54577a );
 a54579a <=( a54578a  and  a54573a );
 a54583a <=( (not A266)  and  A265 );
 a54584a <=( A202  and  a54583a );
 a54587a <=( (not A269)  and  A267 );
 a54590a <=( (not A302)  and  (not A300) );
 a54591a <=( a54590a  and  a54587a );
 a54592a <=( a54591a  and  a54584a );
 a54596a <=( (not A168)  and  (not A169) );
 a54597a <=( (not A170)  and  a54596a );
 a54601a <=( (not A201)  and  (not A166) );
 a54602a <=( A167  and  a54601a );
 a54603a <=( a54602a  and  a54597a );
 a54607a <=( (not A266)  and  A265 );
 a54608a <=( A202  and  a54607a );
 a54611a <=( (not A269)  and  A267 );
 a54614a <=( A299  and  A298 );
 a54615a <=( a54614a  and  a54611a );
 a54616a <=( a54615a  and  a54608a );
 a54620a <=( (not A168)  and  (not A169) );
 a54621a <=( (not A170)  and  a54620a );
 a54625a <=( (not A201)  and  (not A166) );
 a54626a <=( A167  and  a54625a );
 a54627a <=( a54626a  and  a54621a );
 a54631a <=( (not A266)  and  A265 );
 a54632a <=( A202  and  a54631a );
 a54635a <=( (not A269)  and  A267 );
 a54638a <=( (not A299)  and  (not A298) );
 a54639a <=( a54638a  and  a54635a );
 a54640a <=( a54639a  and  a54632a );
 a54644a <=( (not A168)  and  (not A169) );
 a54645a <=( (not A170)  and  a54644a );
 a54649a <=( (not A201)  and  (not A166) );
 a54650a <=( A167  and  a54649a );
 a54651a <=( a54650a  and  a54645a );
 a54655a <=( (not A266)  and  (not A265) );
 a54656a <=( A202  and  a54655a );
 a54659a <=( (not A299)  and  A298 );
 a54662a <=( A301  and  A300 );
 a54663a <=( a54662a  and  a54659a );
 a54664a <=( a54663a  and  a54656a );
 a54668a <=( (not A168)  and  (not A169) );
 a54669a <=( (not A170)  and  a54668a );
 a54673a <=( (not A201)  and  (not A166) );
 a54674a <=( A167  and  a54673a );
 a54675a <=( a54674a  and  a54669a );
 a54679a <=( (not A266)  and  (not A265) );
 a54680a <=( A202  and  a54679a );
 a54683a <=( (not A299)  and  A298 );
 a54686a <=( (not A302)  and  A300 );
 a54687a <=( a54686a  and  a54683a );
 a54688a <=( a54687a  and  a54680a );
 a54692a <=( (not A168)  and  (not A169) );
 a54693a <=( (not A170)  and  a54692a );
 a54697a <=( (not A201)  and  (not A166) );
 a54698a <=( A167  and  a54697a );
 a54699a <=( a54698a  and  a54693a );
 a54703a <=( (not A266)  and  (not A265) );
 a54704a <=( A202  and  a54703a );
 a54707a <=( A299  and  (not A298) );
 a54710a <=( A301  and  A300 );
 a54711a <=( a54710a  and  a54707a );
 a54712a <=( a54711a  and  a54704a );
 a54716a <=( (not A168)  and  (not A169) );
 a54717a <=( (not A170)  and  a54716a );
 a54721a <=( (not A201)  and  (not A166) );
 a54722a <=( A167  and  a54721a );
 a54723a <=( a54722a  and  a54717a );
 a54727a <=( (not A266)  and  (not A265) );
 a54728a <=( A202  and  a54727a );
 a54731a <=( A299  and  (not A298) );
 a54734a <=( (not A302)  and  A300 );
 a54735a <=( a54734a  and  a54731a );
 a54736a <=( a54735a  and  a54728a );
 a54740a <=( (not A168)  and  (not A169) );
 a54741a <=( (not A170)  and  a54740a );
 a54745a <=( (not A201)  and  (not A166) );
 a54746a <=( A167  and  a54745a );
 a54747a <=( a54746a  and  a54741a );
 a54751a <=( A268  and  (not A267) );
 a54752a <=( (not A203)  and  a54751a );
 a54755a <=( (not A299)  and  A298 );
 a54758a <=( A301  and  A300 );
 a54759a <=( a54758a  and  a54755a );
 a54760a <=( a54759a  and  a54752a );
 a54764a <=( (not A168)  and  (not A169) );
 a54765a <=( (not A170)  and  a54764a );
 a54769a <=( (not A201)  and  (not A166) );
 a54770a <=( A167  and  a54769a );
 a54771a <=( a54770a  and  a54765a );
 a54775a <=( A268  and  (not A267) );
 a54776a <=( (not A203)  and  a54775a );
 a54779a <=( (not A299)  and  A298 );
 a54782a <=( (not A302)  and  A300 );
 a54783a <=( a54782a  and  a54779a );
 a54784a <=( a54783a  and  a54776a );
 a54788a <=( (not A168)  and  (not A169) );
 a54789a <=( (not A170)  and  a54788a );
 a54793a <=( (not A201)  and  (not A166) );
 a54794a <=( A167  and  a54793a );
 a54795a <=( a54794a  and  a54789a );
 a54799a <=( A268  and  (not A267) );
 a54800a <=( (not A203)  and  a54799a );
 a54803a <=( A299  and  (not A298) );
 a54806a <=( A301  and  A300 );
 a54807a <=( a54806a  and  a54803a );
 a54808a <=( a54807a  and  a54800a );
 a54812a <=( (not A168)  and  (not A169) );
 a54813a <=( (not A170)  and  a54812a );
 a54817a <=( (not A201)  and  (not A166) );
 a54818a <=( A167  and  a54817a );
 a54819a <=( a54818a  and  a54813a );
 a54823a <=( A268  and  (not A267) );
 a54824a <=( (not A203)  and  a54823a );
 a54827a <=( A299  and  (not A298) );
 a54830a <=( (not A302)  and  A300 );
 a54831a <=( a54830a  and  a54827a );
 a54832a <=( a54831a  and  a54824a );
 a54836a <=( (not A168)  and  (not A169) );
 a54837a <=( (not A170)  and  a54836a );
 a54841a <=( (not A201)  and  (not A166) );
 a54842a <=( A167  and  a54841a );
 a54843a <=( a54842a  and  a54837a );
 a54847a <=( (not A269)  and  (not A267) );
 a54848a <=( (not A203)  and  a54847a );
 a54851a <=( (not A299)  and  A298 );
 a54854a <=( A301  and  A300 );
 a54855a <=( a54854a  and  a54851a );
 a54856a <=( a54855a  and  a54848a );
 a54860a <=( (not A168)  and  (not A169) );
 a54861a <=( (not A170)  and  a54860a );
 a54865a <=( (not A201)  and  (not A166) );
 a54866a <=( A167  and  a54865a );
 a54867a <=( a54866a  and  a54861a );
 a54871a <=( (not A269)  and  (not A267) );
 a54872a <=( (not A203)  and  a54871a );
 a54875a <=( (not A299)  and  A298 );
 a54878a <=( (not A302)  and  A300 );
 a54879a <=( a54878a  and  a54875a );
 a54880a <=( a54879a  and  a54872a );
 a54884a <=( (not A168)  and  (not A169) );
 a54885a <=( (not A170)  and  a54884a );
 a54889a <=( (not A201)  and  (not A166) );
 a54890a <=( A167  and  a54889a );
 a54891a <=( a54890a  and  a54885a );
 a54895a <=( (not A269)  and  (not A267) );
 a54896a <=( (not A203)  and  a54895a );
 a54899a <=( A299  and  (not A298) );
 a54902a <=( A301  and  A300 );
 a54903a <=( a54902a  and  a54899a );
 a54904a <=( a54903a  and  a54896a );
 a54908a <=( (not A168)  and  (not A169) );
 a54909a <=( (not A170)  and  a54908a );
 a54913a <=( (not A201)  and  (not A166) );
 a54914a <=( A167  and  a54913a );
 a54915a <=( a54914a  and  a54909a );
 a54919a <=( (not A269)  and  (not A267) );
 a54920a <=( (not A203)  and  a54919a );
 a54923a <=( A299  and  (not A298) );
 a54926a <=( (not A302)  and  A300 );
 a54927a <=( a54926a  and  a54923a );
 a54928a <=( a54927a  and  a54920a );
 a54932a <=( (not A168)  and  (not A169) );
 a54933a <=( (not A170)  and  a54932a );
 a54937a <=( (not A201)  and  (not A166) );
 a54938a <=( A167  and  a54937a );
 a54939a <=( a54938a  and  a54933a );
 a54943a <=( A266  and  A265 );
 a54944a <=( (not A203)  and  a54943a );
 a54947a <=( (not A299)  and  A298 );
 a54950a <=( A301  and  A300 );
 a54951a <=( a54950a  and  a54947a );
 a54952a <=( a54951a  and  a54944a );
 a54956a <=( (not A168)  and  (not A169) );
 a54957a <=( (not A170)  and  a54956a );
 a54961a <=( (not A201)  and  (not A166) );
 a54962a <=( A167  and  a54961a );
 a54963a <=( a54962a  and  a54957a );
 a54967a <=( A266  and  A265 );
 a54968a <=( (not A203)  and  a54967a );
 a54971a <=( (not A299)  and  A298 );
 a54974a <=( (not A302)  and  A300 );
 a54975a <=( a54974a  and  a54971a );
 a54976a <=( a54975a  and  a54968a );
 a54980a <=( (not A168)  and  (not A169) );
 a54981a <=( (not A170)  and  a54980a );
 a54985a <=( (not A201)  and  (not A166) );
 a54986a <=( A167  and  a54985a );
 a54987a <=( a54986a  and  a54981a );
 a54991a <=( A266  and  A265 );
 a54992a <=( (not A203)  and  a54991a );
 a54995a <=( A299  and  (not A298) );
 a54998a <=( A301  and  A300 );
 a54999a <=( a54998a  and  a54995a );
 a55000a <=( a54999a  and  a54992a );
 a55004a <=( (not A168)  and  (not A169) );
 a55005a <=( (not A170)  and  a55004a );
 a55009a <=( (not A201)  and  (not A166) );
 a55010a <=( A167  and  a55009a );
 a55011a <=( a55010a  and  a55005a );
 a55015a <=( A266  and  A265 );
 a55016a <=( (not A203)  and  a55015a );
 a55019a <=( A299  and  (not A298) );
 a55022a <=( (not A302)  and  A300 );
 a55023a <=( a55022a  and  a55019a );
 a55024a <=( a55023a  and  a55016a );
 a55028a <=( (not A168)  and  (not A169) );
 a55029a <=( (not A170)  and  a55028a );
 a55033a <=( (not A201)  and  (not A166) );
 a55034a <=( A167  and  a55033a );
 a55035a <=( a55034a  and  a55029a );
 a55039a <=( A266  and  (not A265) );
 a55040a <=( (not A203)  and  a55039a );
 a55043a <=( A268  and  A267 );
 a55046a <=( A301  and  (not A300) );
 a55047a <=( a55046a  and  a55043a );
 a55048a <=( a55047a  and  a55040a );
 a55052a <=( (not A168)  and  (not A169) );
 a55053a <=( (not A170)  and  a55052a );
 a55057a <=( (not A201)  and  (not A166) );
 a55058a <=( A167  and  a55057a );
 a55059a <=( a55058a  and  a55053a );
 a55063a <=( A266  and  (not A265) );
 a55064a <=( (not A203)  and  a55063a );
 a55067a <=( A268  and  A267 );
 a55070a <=( (not A302)  and  (not A300) );
 a55071a <=( a55070a  and  a55067a );
 a55072a <=( a55071a  and  a55064a );
 a55076a <=( (not A168)  and  (not A169) );
 a55077a <=( (not A170)  and  a55076a );
 a55081a <=( (not A201)  and  (not A166) );
 a55082a <=( A167  and  a55081a );
 a55083a <=( a55082a  and  a55077a );
 a55087a <=( A266  and  (not A265) );
 a55088a <=( (not A203)  and  a55087a );
 a55091a <=( A268  and  A267 );
 a55094a <=( A299  and  A298 );
 a55095a <=( a55094a  and  a55091a );
 a55096a <=( a55095a  and  a55088a );
 a55100a <=( (not A168)  and  (not A169) );
 a55101a <=( (not A170)  and  a55100a );
 a55105a <=( (not A201)  and  (not A166) );
 a55106a <=( A167  and  a55105a );
 a55107a <=( a55106a  and  a55101a );
 a55111a <=( A266  and  (not A265) );
 a55112a <=( (not A203)  and  a55111a );
 a55115a <=( A268  and  A267 );
 a55118a <=( (not A299)  and  (not A298) );
 a55119a <=( a55118a  and  a55115a );
 a55120a <=( a55119a  and  a55112a );
 a55124a <=( (not A168)  and  (not A169) );
 a55125a <=( (not A170)  and  a55124a );
 a55129a <=( (not A201)  and  (not A166) );
 a55130a <=( A167  and  a55129a );
 a55131a <=( a55130a  and  a55125a );
 a55135a <=( A266  and  (not A265) );
 a55136a <=( (not A203)  and  a55135a );
 a55139a <=( (not A269)  and  A267 );
 a55142a <=( A301  and  (not A300) );
 a55143a <=( a55142a  and  a55139a );
 a55144a <=( a55143a  and  a55136a );
 a55148a <=( (not A168)  and  (not A169) );
 a55149a <=( (not A170)  and  a55148a );
 a55153a <=( (not A201)  and  (not A166) );
 a55154a <=( A167  and  a55153a );
 a55155a <=( a55154a  and  a55149a );
 a55159a <=( A266  and  (not A265) );
 a55160a <=( (not A203)  and  a55159a );
 a55163a <=( (not A269)  and  A267 );
 a55166a <=( (not A302)  and  (not A300) );
 a55167a <=( a55166a  and  a55163a );
 a55168a <=( a55167a  and  a55160a );
 a55172a <=( (not A168)  and  (not A169) );
 a55173a <=( (not A170)  and  a55172a );
 a55177a <=( (not A201)  and  (not A166) );
 a55178a <=( A167  and  a55177a );
 a55179a <=( a55178a  and  a55173a );
 a55183a <=( A266  and  (not A265) );
 a55184a <=( (not A203)  and  a55183a );
 a55187a <=( (not A269)  and  A267 );
 a55190a <=( A299  and  A298 );
 a55191a <=( a55190a  and  a55187a );
 a55192a <=( a55191a  and  a55184a );
 a55196a <=( (not A168)  and  (not A169) );
 a55197a <=( (not A170)  and  a55196a );
 a55201a <=( (not A201)  and  (not A166) );
 a55202a <=( A167  and  a55201a );
 a55203a <=( a55202a  and  a55197a );
 a55207a <=( A266  and  (not A265) );
 a55208a <=( (not A203)  and  a55207a );
 a55211a <=( (not A269)  and  A267 );
 a55214a <=( (not A299)  and  (not A298) );
 a55215a <=( a55214a  and  a55211a );
 a55216a <=( a55215a  and  a55208a );
 a55220a <=( (not A168)  and  (not A169) );
 a55221a <=( (not A170)  and  a55220a );
 a55225a <=( (not A201)  and  (not A166) );
 a55226a <=( A167  and  a55225a );
 a55227a <=( a55226a  and  a55221a );
 a55231a <=( (not A266)  and  A265 );
 a55232a <=( (not A203)  and  a55231a );
 a55235a <=( A268  and  A267 );
 a55238a <=( A301  and  (not A300) );
 a55239a <=( a55238a  and  a55235a );
 a55240a <=( a55239a  and  a55232a );
 a55244a <=( (not A168)  and  (not A169) );
 a55245a <=( (not A170)  and  a55244a );
 a55249a <=( (not A201)  and  (not A166) );
 a55250a <=( A167  and  a55249a );
 a55251a <=( a55250a  and  a55245a );
 a55255a <=( (not A266)  and  A265 );
 a55256a <=( (not A203)  and  a55255a );
 a55259a <=( A268  and  A267 );
 a55262a <=( (not A302)  and  (not A300) );
 a55263a <=( a55262a  and  a55259a );
 a55264a <=( a55263a  and  a55256a );
 a55268a <=( (not A168)  and  (not A169) );
 a55269a <=( (not A170)  and  a55268a );
 a55273a <=( (not A201)  and  (not A166) );
 a55274a <=( A167  and  a55273a );
 a55275a <=( a55274a  and  a55269a );
 a55279a <=( (not A266)  and  A265 );
 a55280a <=( (not A203)  and  a55279a );
 a55283a <=( A268  and  A267 );
 a55286a <=( A299  and  A298 );
 a55287a <=( a55286a  and  a55283a );
 a55288a <=( a55287a  and  a55280a );
 a55292a <=( (not A168)  and  (not A169) );
 a55293a <=( (not A170)  and  a55292a );
 a55297a <=( (not A201)  and  (not A166) );
 a55298a <=( A167  and  a55297a );
 a55299a <=( a55298a  and  a55293a );
 a55303a <=( (not A266)  and  A265 );
 a55304a <=( (not A203)  and  a55303a );
 a55307a <=( A268  and  A267 );
 a55310a <=( (not A299)  and  (not A298) );
 a55311a <=( a55310a  and  a55307a );
 a55312a <=( a55311a  and  a55304a );
 a55316a <=( (not A168)  and  (not A169) );
 a55317a <=( (not A170)  and  a55316a );
 a55321a <=( (not A201)  and  (not A166) );
 a55322a <=( A167  and  a55321a );
 a55323a <=( a55322a  and  a55317a );
 a55327a <=( (not A266)  and  A265 );
 a55328a <=( (not A203)  and  a55327a );
 a55331a <=( (not A269)  and  A267 );
 a55334a <=( A301  and  (not A300) );
 a55335a <=( a55334a  and  a55331a );
 a55336a <=( a55335a  and  a55328a );
 a55340a <=( (not A168)  and  (not A169) );
 a55341a <=( (not A170)  and  a55340a );
 a55345a <=( (not A201)  and  (not A166) );
 a55346a <=( A167  and  a55345a );
 a55347a <=( a55346a  and  a55341a );
 a55351a <=( (not A266)  and  A265 );
 a55352a <=( (not A203)  and  a55351a );
 a55355a <=( (not A269)  and  A267 );
 a55358a <=( (not A302)  and  (not A300) );
 a55359a <=( a55358a  and  a55355a );
 a55360a <=( a55359a  and  a55352a );
 a55364a <=( (not A168)  and  (not A169) );
 a55365a <=( (not A170)  and  a55364a );
 a55369a <=( (not A201)  and  (not A166) );
 a55370a <=( A167  and  a55369a );
 a55371a <=( a55370a  and  a55365a );
 a55375a <=( (not A266)  and  A265 );
 a55376a <=( (not A203)  and  a55375a );
 a55379a <=( (not A269)  and  A267 );
 a55382a <=( A299  and  A298 );
 a55383a <=( a55382a  and  a55379a );
 a55384a <=( a55383a  and  a55376a );
 a55388a <=( (not A168)  and  (not A169) );
 a55389a <=( (not A170)  and  a55388a );
 a55393a <=( (not A201)  and  (not A166) );
 a55394a <=( A167  and  a55393a );
 a55395a <=( a55394a  and  a55389a );
 a55399a <=( (not A266)  and  A265 );
 a55400a <=( (not A203)  and  a55399a );
 a55403a <=( (not A269)  and  A267 );
 a55406a <=( (not A299)  and  (not A298) );
 a55407a <=( a55406a  and  a55403a );
 a55408a <=( a55407a  and  a55400a );
 a55412a <=( (not A168)  and  (not A169) );
 a55413a <=( (not A170)  and  a55412a );
 a55417a <=( (not A201)  and  (not A166) );
 a55418a <=( A167  and  a55417a );
 a55419a <=( a55418a  and  a55413a );
 a55423a <=( (not A266)  and  (not A265) );
 a55424a <=( (not A203)  and  a55423a );
 a55427a <=( (not A299)  and  A298 );
 a55430a <=( A301  and  A300 );
 a55431a <=( a55430a  and  a55427a );
 a55432a <=( a55431a  and  a55424a );
 a55436a <=( (not A168)  and  (not A169) );
 a55437a <=( (not A170)  and  a55436a );
 a55441a <=( (not A201)  and  (not A166) );
 a55442a <=( A167  and  a55441a );
 a55443a <=( a55442a  and  a55437a );
 a55447a <=( (not A266)  and  (not A265) );
 a55448a <=( (not A203)  and  a55447a );
 a55451a <=( (not A299)  and  A298 );
 a55454a <=( (not A302)  and  A300 );
 a55455a <=( a55454a  and  a55451a );
 a55456a <=( a55455a  and  a55448a );
 a55460a <=( (not A168)  and  (not A169) );
 a55461a <=( (not A170)  and  a55460a );
 a55465a <=( (not A201)  and  (not A166) );
 a55466a <=( A167  and  a55465a );
 a55467a <=( a55466a  and  a55461a );
 a55471a <=( (not A266)  and  (not A265) );
 a55472a <=( (not A203)  and  a55471a );
 a55475a <=( A299  and  (not A298) );
 a55478a <=( A301  and  A300 );
 a55479a <=( a55478a  and  a55475a );
 a55480a <=( a55479a  and  a55472a );
 a55484a <=( (not A168)  and  (not A169) );
 a55485a <=( (not A170)  and  a55484a );
 a55489a <=( (not A201)  and  (not A166) );
 a55490a <=( A167  and  a55489a );
 a55491a <=( a55490a  and  a55485a );
 a55495a <=( (not A266)  and  (not A265) );
 a55496a <=( (not A203)  and  a55495a );
 a55499a <=( A299  and  (not A298) );
 a55502a <=( (not A302)  and  A300 );
 a55503a <=( a55502a  and  a55499a );
 a55504a <=( a55503a  and  a55496a );
 a55508a <=( (not A168)  and  (not A169) );
 a55509a <=( (not A170)  and  a55508a );
 a55513a <=( A199  and  (not A166) );
 a55514a <=( A167  and  a55513a );
 a55515a <=( a55514a  and  a55509a );
 a55519a <=( A268  and  (not A267) );
 a55520a <=( A200  and  a55519a );
 a55523a <=( (not A299)  and  A298 );
 a55526a <=( A301  and  A300 );
 a55527a <=( a55526a  and  a55523a );
 a55528a <=( a55527a  and  a55520a );
 a55532a <=( (not A168)  and  (not A169) );
 a55533a <=( (not A170)  and  a55532a );
 a55537a <=( A199  and  (not A166) );
 a55538a <=( A167  and  a55537a );
 a55539a <=( a55538a  and  a55533a );
 a55543a <=( A268  and  (not A267) );
 a55544a <=( A200  and  a55543a );
 a55547a <=( (not A299)  and  A298 );
 a55550a <=( (not A302)  and  A300 );
 a55551a <=( a55550a  and  a55547a );
 a55552a <=( a55551a  and  a55544a );
 a55556a <=( (not A168)  and  (not A169) );
 a55557a <=( (not A170)  and  a55556a );
 a55561a <=( A199  and  (not A166) );
 a55562a <=( A167  and  a55561a );
 a55563a <=( a55562a  and  a55557a );
 a55567a <=( A268  and  (not A267) );
 a55568a <=( A200  and  a55567a );
 a55571a <=( A299  and  (not A298) );
 a55574a <=( A301  and  A300 );
 a55575a <=( a55574a  and  a55571a );
 a55576a <=( a55575a  and  a55568a );
 a55580a <=( (not A168)  and  (not A169) );
 a55581a <=( (not A170)  and  a55580a );
 a55585a <=( A199  and  (not A166) );
 a55586a <=( A167  and  a55585a );
 a55587a <=( a55586a  and  a55581a );
 a55591a <=( A268  and  (not A267) );
 a55592a <=( A200  and  a55591a );
 a55595a <=( A299  and  (not A298) );
 a55598a <=( (not A302)  and  A300 );
 a55599a <=( a55598a  and  a55595a );
 a55600a <=( a55599a  and  a55592a );
 a55604a <=( (not A168)  and  (not A169) );
 a55605a <=( (not A170)  and  a55604a );
 a55609a <=( A199  and  (not A166) );
 a55610a <=( A167  and  a55609a );
 a55611a <=( a55610a  and  a55605a );
 a55615a <=( (not A269)  and  (not A267) );
 a55616a <=( A200  and  a55615a );
 a55619a <=( (not A299)  and  A298 );
 a55622a <=( A301  and  A300 );
 a55623a <=( a55622a  and  a55619a );
 a55624a <=( a55623a  and  a55616a );
 a55628a <=( (not A168)  and  (not A169) );
 a55629a <=( (not A170)  and  a55628a );
 a55633a <=( A199  and  (not A166) );
 a55634a <=( A167  and  a55633a );
 a55635a <=( a55634a  and  a55629a );
 a55639a <=( (not A269)  and  (not A267) );
 a55640a <=( A200  and  a55639a );
 a55643a <=( (not A299)  and  A298 );
 a55646a <=( (not A302)  and  A300 );
 a55647a <=( a55646a  and  a55643a );
 a55648a <=( a55647a  and  a55640a );
 a55652a <=( (not A168)  and  (not A169) );
 a55653a <=( (not A170)  and  a55652a );
 a55657a <=( A199  and  (not A166) );
 a55658a <=( A167  and  a55657a );
 a55659a <=( a55658a  and  a55653a );
 a55663a <=( (not A269)  and  (not A267) );
 a55664a <=( A200  and  a55663a );
 a55667a <=( A299  and  (not A298) );
 a55670a <=( A301  and  A300 );
 a55671a <=( a55670a  and  a55667a );
 a55672a <=( a55671a  and  a55664a );
 a55676a <=( (not A168)  and  (not A169) );
 a55677a <=( (not A170)  and  a55676a );
 a55681a <=( A199  and  (not A166) );
 a55682a <=( A167  and  a55681a );
 a55683a <=( a55682a  and  a55677a );
 a55687a <=( (not A269)  and  (not A267) );
 a55688a <=( A200  and  a55687a );
 a55691a <=( A299  and  (not A298) );
 a55694a <=( (not A302)  and  A300 );
 a55695a <=( a55694a  and  a55691a );
 a55696a <=( a55695a  and  a55688a );
 a55700a <=( (not A168)  and  (not A169) );
 a55701a <=( (not A170)  and  a55700a );
 a55705a <=( A199  and  (not A166) );
 a55706a <=( A167  and  a55705a );
 a55707a <=( a55706a  and  a55701a );
 a55711a <=( A266  and  A265 );
 a55712a <=( A200  and  a55711a );
 a55715a <=( (not A299)  and  A298 );
 a55718a <=( A301  and  A300 );
 a55719a <=( a55718a  and  a55715a );
 a55720a <=( a55719a  and  a55712a );
 a55724a <=( (not A168)  and  (not A169) );
 a55725a <=( (not A170)  and  a55724a );
 a55729a <=( A199  and  (not A166) );
 a55730a <=( A167  and  a55729a );
 a55731a <=( a55730a  and  a55725a );
 a55735a <=( A266  and  A265 );
 a55736a <=( A200  and  a55735a );
 a55739a <=( (not A299)  and  A298 );
 a55742a <=( (not A302)  and  A300 );
 a55743a <=( a55742a  and  a55739a );
 a55744a <=( a55743a  and  a55736a );
 a55748a <=( (not A168)  and  (not A169) );
 a55749a <=( (not A170)  and  a55748a );
 a55753a <=( A199  and  (not A166) );
 a55754a <=( A167  and  a55753a );
 a55755a <=( a55754a  and  a55749a );
 a55759a <=( A266  and  A265 );
 a55760a <=( A200  and  a55759a );
 a55763a <=( A299  and  (not A298) );
 a55766a <=( A301  and  A300 );
 a55767a <=( a55766a  and  a55763a );
 a55768a <=( a55767a  and  a55760a );
 a55772a <=( (not A168)  and  (not A169) );
 a55773a <=( (not A170)  and  a55772a );
 a55777a <=( A199  and  (not A166) );
 a55778a <=( A167  and  a55777a );
 a55779a <=( a55778a  and  a55773a );
 a55783a <=( A266  and  A265 );
 a55784a <=( A200  and  a55783a );
 a55787a <=( A299  and  (not A298) );
 a55790a <=( (not A302)  and  A300 );
 a55791a <=( a55790a  and  a55787a );
 a55792a <=( a55791a  and  a55784a );
 a55796a <=( (not A168)  and  (not A169) );
 a55797a <=( (not A170)  and  a55796a );
 a55801a <=( A199  and  (not A166) );
 a55802a <=( A167  and  a55801a );
 a55803a <=( a55802a  and  a55797a );
 a55807a <=( A266  and  (not A265) );
 a55808a <=( A200  and  a55807a );
 a55811a <=( A268  and  A267 );
 a55814a <=( A301  and  (not A300) );
 a55815a <=( a55814a  and  a55811a );
 a55816a <=( a55815a  and  a55808a );
 a55820a <=( (not A168)  and  (not A169) );
 a55821a <=( (not A170)  and  a55820a );
 a55825a <=( A199  and  (not A166) );
 a55826a <=( A167  and  a55825a );
 a55827a <=( a55826a  and  a55821a );
 a55831a <=( A266  and  (not A265) );
 a55832a <=( A200  and  a55831a );
 a55835a <=( A268  and  A267 );
 a55838a <=( (not A302)  and  (not A300) );
 a55839a <=( a55838a  and  a55835a );
 a55840a <=( a55839a  and  a55832a );
 a55844a <=( (not A168)  and  (not A169) );
 a55845a <=( (not A170)  and  a55844a );
 a55849a <=( A199  and  (not A166) );
 a55850a <=( A167  and  a55849a );
 a55851a <=( a55850a  and  a55845a );
 a55855a <=( A266  and  (not A265) );
 a55856a <=( A200  and  a55855a );
 a55859a <=( A268  and  A267 );
 a55862a <=( A299  and  A298 );
 a55863a <=( a55862a  and  a55859a );
 a55864a <=( a55863a  and  a55856a );
 a55868a <=( (not A168)  and  (not A169) );
 a55869a <=( (not A170)  and  a55868a );
 a55873a <=( A199  and  (not A166) );
 a55874a <=( A167  and  a55873a );
 a55875a <=( a55874a  and  a55869a );
 a55879a <=( A266  and  (not A265) );
 a55880a <=( A200  and  a55879a );
 a55883a <=( A268  and  A267 );
 a55886a <=( (not A299)  and  (not A298) );
 a55887a <=( a55886a  and  a55883a );
 a55888a <=( a55887a  and  a55880a );
 a55892a <=( (not A168)  and  (not A169) );
 a55893a <=( (not A170)  and  a55892a );
 a55897a <=( A199  and  (not A166) );
 a55898a <=( A167  and  a55897a );
 a55899a <=( a55898a  and  a55893a );
 a55903a <=( A266  and  (not A265) );
 a55904a <=( A200  and  a55903a );
 a55907a <=( (not A269)  and  A267 );
 a55910a <=( A301  and  (not A300) );
 a55911a <=( a55910a  and  a55907a );
 a55912a <=( a55911a  and  a55904a );
 a55916a <=( (not A168)  and  (not A169) );
 a55917a <=( (not A170)  and  a55916a );
 a55921a <=( A199  and  (not A166) );
 a55922a <=( A167  and  a55921a );
 a55923a <=( a55922a  and  a55917a );
 a55927a <=( A266  and  (not A265) );
 a55928a <=( A200  and  a55927a );
 a55931a <=( (not A269)  and  A267 );
 a55934a <=( (not A302)  and  (not A300) );
 a55935a <=( a55934a  and  a55931a );
 a55936a <=( a55935a  and  a55928a );
 a55940a <=( (not A168)  and  (not A169) );
 a55941a <=( (not A170)  and  a55940a );
 a55945a <=( A199  and  (not A166) );
 a55946a <=( A167  and  a55945a );
 a55947a <=( a55946a  and  a55941a );
 a55951a <=( A266  and  (not A265) );
 a55952a <=( A200  and  a55951a );
 a55955a <=( (not A269)  and  A267 );
 a55958a <=( A299  and  A298 );
 a55959a <=( a55958a  and  a55955a );
 a55960a <=( a55959a  and  a55952a );
 a55964a <=( (not A168)  and  (not A169) );
 a55965a <=( (not A170)  and  a55964a );
 a55969a <=( A199  and  (not A166) );
 a55970a <=( A167  and  a55969a );
 a55971a <=( a55970a  and  a55965a );
 a55975a <=( A266  and  (not A265) );
 a55976a <=( A200  and  a55975a );
 a55979a <=( (not A269)  and  A267 );
 a55982a <=( (not A299)  and  (not A298) );
 a55983a <=( a55982a  and  a55979a );
 a55984a <=( a55983a  and  a55976a );
 a55988a <=( (not A168)  and  (not A169) );
 a55989a <=( (not A170)  and  a55988a );
 a55993a <=( A199  and  (not A166) );
 a55994a <=( A167  and  a55993a );
 a55995a <=( a55994a  and  a55989a );
 a55999a <=( (not A266)  and  A265 );
 a56000a <=( A200  and  a55999a );
 a56003a <=( A268  and  A267 );
 a56006a <=( A301  and  (not A300) );
 a56007a <=( a56006a  and  a56003a );
 a56008a <=( a56007a  and  a56000a );
 a56012a <=( (not A168)  and  (not A169) );
 a56013a <=( (not A170)  and  a56012a );
 a56017a <=( A199  and  (not A166) );
 a56018a <=( A167  and  a56017a );
 a56019a <=( a56018a  and  a56013a );
 a56023a <=( (not A266)  and  A265 );
 a56024a <=( A200  and  a56023a );
 a56027a <=( A268  and  A267 );
 a56030a <=( (not A302)  and  (not A300) );
 a56031a <=( a56030a  and  a56027a );
 a56032a <=( a56031a  and  a56024a );
 a56036a <=( (not A168)  and  (not A169) );
 a56037a <=( (not A170)  and  a56036a );
 a56041a <=( A199  and  (not A166) );
 a56042a <=( A167  and  a56041a );
 a56043a <=( a56042a  and  a56037a );
 a56047a <=( (not A266)  and  A265 );
 a56048a <=( A200  and  a56047a );
 a56051a <=( A268  and  A267 );
 a56054a <=( A299  and  A298 );
 a56055a <=( a56054a  and  a56051a );
 a56056a <=( a56055a  and  a56048a );
 a56060a <=( (not A168)  and  (not A169) );
 a56061a <=( (not A170)  and  a56060a );
 a56065a <=( A199  and  (not A166) );
 a56066a <=( A167  and  a56065a );
 a56067a <=( a56066a  and  a56061a );
 a56071a <=( (not A266)  and  A265 );
 a56072a <=( A200  and  a56071a );
 a56075a <=( A268  and  A267 );
 a56078a <=( (not A299)  and  (not A298) );
 a56079a <=( a56078a  and  a56075a );
 a56080a <=( a56079a  and  a56072a );
 a56084a <=( (not A168)  and  (not A169) );
 a56085a <=( (not A170)  and  a56084a );
 a56089a <=( A199  and  (not A166) );
 a56090a <=( A167  and  a56089a );
 a56091a <=( a56090a  and  a56085a );
 a56095a <=( (not A266)  and  A265 );
 a56096a <=( A200  and  a56095a );
 a56099a <=( (not A269)  and  A267 );
 a56102a <=( A301  and  (not A300) );
 a56103a <=( a56102a  and  a56099a );
 a56104a <=( a56103a  and  a56096a );
 a56108a <=( (not A168)  and  (not A169) );
 a56109a <=( (not A170)  and  a56108a );
 a56113a <=( A199  and  (not A166) );
 a56114a <=( A167  and  a56113a );
 a56115a <=( a56114a  and  a56109a );
 a56119a <=( (not A266)  and  A265 );
 a56120a <=( A200  and  a56119a );
 a56123a <=( (not A269)  and  A267 );
 a56126a <=( (not A302)  and  (not A300) );
 a56127a <=( a56126a  and  a56123a );
 a56128a <=( a56127a  and  a56120a );
 a56132a <=( (not A168)  and  (not A169) );
 a56133a <=( (not A170)  and  a56132a );
 a56137a <=( A199  and  (not A166) );
 a56138a <=( A167  and  a56137a );
 a56139a <=( a56138a  and  a56133a );
 a56143a <=( (not A266)  and  A265 );
 a56144a <=( A200  and  a56143a );
 a56147a <=( (not A269)  and  A267 );
 a56150a <=( A299  and  A298 );
 a56151a <=( a56150a  and  a56147a );
 a56152a <=( a56151a  and  a56144a );
 a56156a <=( (not A168)  and  (not A169) );
 a56157a <=( (not A170)  and  a56156a );
 a56161a <=( A199  and  (not A166) );
 a56162a <=( A167  and  a56161a );
 a56163a <=( a56162a  and  a56157a );
 a56167a <=( (not A266)  and  A265 );
 a56168a <=( A200  and  a56167a );
 a56171a <=( (not A269)  and  A267 );
 a56174a <=( (not A299)  and  (not A298) );
 a56175a <=( a56174a  and  a56171a );
 a56176a <=( a56175a  and  a56168a );
 a56180a <=( (not A168)  and  (not A169) );
 a56181a <=( (not A170)  and  a56180a );
 a56185a <=( A199  and  (not A166) );
 a56186a <=( A167  and  a56185a );
 a56187a <=( a56186a  and  a56181a );
 a56191a <=( (not A266)  and  (not A265) );
 a56192a <=( A200  and  a56191a );
 a56195a <=( (not A299)  and  A298 );
 a56198a <=( A301  and  A300 );
 a56199a <=( a56198a  and  a56195a );
 a56200a <=( a56199a  and  a56192a );
 a56204a <=( (not A168)  and  (not A169) );
 a56205a <=( (not A170)  and  a56204a );
 a56209a <=( A199  and  (not A166) );
 a56210a <=( A167  and  a56209a );
 a56211a <=( a56210a  and  a56205a );
 a56215a <=( (not A266)  and  (not A265) );
 a56216a <=( A200  and  a56215a );
 a56219a <=( (not A299)  and  A298 );
 a56222a <=( (not A302)  and  A300 );
 a56223a <=( a56222a  and  a56219a );
 a56224a <=( a56223a  and  a56216a );
 a56228a <=( (not A168)  and  (not A169) );
 a56229a <=( (not A170)  and  a56228a );
 a56233a <=( A199  and  (not A166) );
 a56234a <=( A167  and  a56233a );
 a56235a <=( a56234a  and  a56229a );
 a56239a <=( (not A266)  and  (not A265) );
 a56240a <=( A200  and  a56239a );
 a56243a <=( A299  and  (not A298) );
 a56246a <=( A301  and  A300 );
 a56247a <=( a56246a  and  a56243a );
 a56248a <=( a56247a  and  a56240a );
 a56252a <=( (not A168)  and  (not A169) );
 a56253a <=( (not A170)  and  a56252a );
 a56257a <=( A199  and  (not A166) );
 a56258a <=( A167  and  a56257a );
 a56259a <=( a56258a  and  a56253a );
 a56263a <=( (not A266)  and  (not A265) );
 a56264a <=( A200  and  a56263a );
 a56267a <=( A299  and  (not A298) );
 a56270a <=( (not A302)  and  A300 );
 a56271a <=( a56270a  and  a56267a );
 a56272a <=( a56271a  and  a56264a );
 a56276a <=( (not A168)  and  (not A169) );
 a56277a <=( (not A170)  and  a56276a );
 a56281a <=( (not A199)  and  (not A166) );
 a56282a <=( A167  and  a56281a );
 a56283a <=( a56282a  and  a56277a );
 a56287a <=( A268  and  (not A267) );
 a56288a <=( (not A200)  and  a56287a );
 a56291a <=( (not A299)  and  A298 );
 a56294a <=( A301  and  A300 );
 a56295a <=( a56294a  and  a56291a );
 a56296a <=( a56295a  and  a56288a );
 a56300a <=( (not A168)  and  (not A169) );
 a56301a <=( (not A170)  and  a56300a );
 a56305a <=( (not A199)  and  (not A166) );
 a56306a <=( A167  and  a56305a );
 a56307a <=( a56306a  and  a56301a );
 a56311a <=( A268  and  (not A267) );
 a56312a <=( (not A200)  and  a56311a );
 a56315a <=( (not A299)  and  A298 );
 a56318a <=( (not A302)  and  A300 );
 a56319a <=( a56318a  and  a56315a );
 a56320a <=( a56319a  and  a56312a );
 a56324a <=( (not A168)  and  (not A169) );
 a56325a <=( (not A170)  and  a56324a );
 a56329a <=( (not A199)  and  (not A166) );
 a56330a <=( A167  and  a56329a );
 a56331a <=( a56330a  and  a56325a );
 a56335a <=( A268  and  (not A267) );
 a56336a <=( (not A200)  and  a56335a );
 a56339a <=( A299  and  (not A298) );
 a56342a <=( A301  and  A300 );
 a56343a <=( a56342a  and  a56339a );
 a56344a <=( a56343a  and  a56336a );
 a56348a <=( (not A168)  and  (not A169) );
 a56349a <=( (not A170)  and  a56348a );
 a56353a <=( (not A199)  and  (not A166) );
 a56354a <=( A167  and  a56353a );
 a56355a <=( a56354a  and  a56349a );
 a56359a <=( A268  and  (not A267) );
 a56360a <=( (not A200)  and  a56359a );
 a56363a <=( A299  and  (not A298) );
 a56366a <=( (not A302)  and  A300 );
 a56367a <=( a56366a  and  a56363a );
 a56368a <=( a56367a  and  a56360a );
 a56372a <=( (not A168)  and  (not A169) );
 a56373a <=( (not A170)  and  a56372a );
 a56377a <=( (not A199)  and  (not A166) );
 a56378a <=( A167  and  a56377a );
 a56379a <=( a56378a  and  a56373a );
 a56383a <=( (not A269)  and  (not A267) );
 a56384a <=( (not A200)  and  a56383a );
 a56387a <=( (not A299)  and  A298 );
 a56390a <=( A301  and  A300 );
 a56391a <=( a56390a  and  a56387a );
 a56392a <=( a56391a  and  a56384a );
 a56396a <=( (not A168)  and  (not A169) );
 a56397a <=( (not A170)  and  a56396a );
 a56401a <=( (not A199)  and  (not A166) );
 a56402a <=( A167  and  a56401a );
 a56403a <=( a56402a  and  a56397a );
 a56407a <=( (not A269)  and  (not A267) );
 a56408a <=( (not A200)  and  a56407a );
 a56411a <=( (not A299)  and  A298 );
 a56414a <=( (not A302)  and  A300 );
 a56415a <=( a56414a  and  a56411a );
 a56416a <=( a56415a  and  a56408a );
 a56420a <=( (not A168)  and  (not A169) );
 a56421a <=( (not A170)  and  a56420a );
 a56425a <=( (not A199)  and  (not A166) );
 a56426a <=( A167  and  a56425a );
 a56427a <=( a56426a  and  a56421a );
 a56431a <=( (not A269)  and  (not A267) );
 a56432a <=( (not A200)  and  a56431a );
 a56435a <=( A299  and  (not A298) );
 a56438a <=( A301  and  A300 );
 a56439a <=( a56438a  and  a56435a );
 a56440a <=( a56439a  and  a56432a );
 a56444a <=( (not A168)  and  (not A169) );
 a56445a <=( (not A170)  and  a56444a );
 a56449a <=( (not A199)  and  (not A166) );
 a56450a <=( A167  and  a56449a );
 a56451a <=( a56450a  and  a56445a );
 a56455a <=( (not A269)  and  (not A267) );
 a56456a <=( (not A200)  and  a56455a );
 a56459a <=( A299  and  (not A298) );
 a56462a <=( (not A302)  and  A300 );
 a56463a <=( a56462a  and  a56459a );
 a56464a <=( a56463a  and  a56456a );
 a56468a <=( (not A168)  and  (not A169) );
 a56469a <=( (not A170)  and  a56468a );
 a56473a <=( (not A199)  and  (not A166) );
 a56474a <=( A167  and  a56473a );
 a56475a <=( a56474a  and  a56469a );
 a56479a <=( A266  and  A265 );
 a56480a <=( (not A200)  and  a56479a );
 a56483a <=( (not A299)  and  A298 );
 a56486a <=( A301  and  A300 );
 a56487a <=( a56486a  and  a56483a );
 a56488a <=( a56487a  and  a56480a );
 a56492a <=( (not A168)  and  (not A169) );
 a56493a <=( (not A170)  and  a56492a );
 a56497a <=( (not A199)  and  (not A166) );
 a56498a <=( A167  and  a56497a );
 a56499a <=( a56498a  and  a56493a );
 a56503a <=( A266  and  A265 );
 a56504a <=( (not A200)  and  a56503a );
 a56507a <=( (not A299)  and  A298 );
 a56510a <=( (not A302)  and  A300 );
 a56511a <=( a56510a  and  a56507a );
 a56512a <=( a56511a  and  a56504a );
 a56516a <=( (not A168)  and  (not A169) );
 a56517a <=( (not A170)  and  a56516a );
 a56521a <=( (not A199)  and  (not A166) );
 a56522a <=( A167  and  a56521a );
 a56523a <=( a56522a  and  a56517a );
 a56527a <=( A266  and  A265 );
 a56528a <=( (not A200)  and  a56527a );
 a56531a <=( A299  and  (not A298) );
 a56534a <=( A301  and  A300 );
 a56535a <=( a56534a  and  a56531a );
 a56536a <=( a56535a  and  a56528a );
 a56540a <=( (not A168)  and  (not A169) );
 a56541a <=( (not A170)  and  a56540a );
 a56545a <=( (not A199)  and  (not A166) );
 a56546a <=( A167  and  a56545a );
 a56547a <=( a56546a  and  a56541a );
 a56551a <=( A266  and  A265 );
 a56552a <=( (not A200)  and  a56551a );
 a56555a <=( A299  and  (not A298) );
 a56558a <=( (not A302)  and  A300 );
 a56559a <=( a56558a  and  a56555a );
 a56560a <=( a56559a  and  a56552a );
 a56564a <=( (not A168)  and  (not A169) );
 a56565a <=( (not A170)  and  a56564a );
 a56569a <=( (not A199)  and  (not A166) );
 a56570a <=( A167  and  a56569a );
 a56571a <=( a56570a  and  a56565a );
 a56575a <=( A266  and  (not A265) );
 a56576a <=( (not A200)  and  a56575a );
 a56579a <=( A268  and  A267 );
 a56582a <=( A301  and  (not A300) );
 a56583a <=( a56582a  and  a56579a );
 a56584a <=( a56583a  and  a56576a );
 a56588a <=( (not A168)  and  (not A169) );
 a56589a <=( (not A170)  and  a56588a );
 a56593a <=( (not A199)  and  (not A166) );
 a56594a <=( A167  and  a56593a );
 a56595a <=( a56594a  and  a56589a );
 a56599a <=( A266  and  (not A265) );
 a56600a <=( (not A200)  and  a56599a );
 a56603a <=( A268  and  A267 );
 a56606a <=( (not A302)  and  (not A300) );
 a56607a <=( a56606a  and  a56603a );
 a56608a <=( a56607a  and  a56600a );
 a56612a <=( (not A168)  and  (not A169) );
 a56613a <=( (not A170)  and  a56612a );
 a56617a <=( (not A199)  and  (not A166) );
 a56618a <=( A167  and  a56617a );
 a56619a <=( a56618a  and  a56613a );
 a56623a <=( A266  and  (not A265) );
 a56624a <=( (not A200)  and  a56623a );
 a56627a <=( A268  and  A267 );
 a56630a <=( A299  and  A298 );
 a56631a <=( a56630a  and  a56627a );
 a56632a <=( a56631a  and  a56624a );
 a56636a <=( (not A168)  and  (not A169) );
 a56637a <=( (not A170)  and  a56636a );
 a56641a <=( (not A199)  and  (not A166) );
 a56642a <=( A167  and  a56641a );
 a56643a <=( a56642a  and  a56637a );
 a56647a <=( A266  and  (not A265) );
 a56648a <=( (not A200)  and  a56647a );
 a56651a <=( A268  and  A267 );
 a56654a <=( (not A299)  and  (not A298) );
 a56655a <=( a56654a  and  a56651a );
 a56656a <=( a56655a  and  a56648a );
 a56660a <=( (not A168)  and  (not A169) );
 a56661a <=( (not A170)  and  a56660a );
 a56665a <=( (not A199)  and  (not A166) );
 a56666a <=( A167  and  a56665a );
 a56667a <=( a56666a  and  a56661a );
 a56671a <=( A266  and  (not A265) );
 a56672a <=( (not A200)  and  a56671a );
 a56675a <=( (not A269)  and  A267 );
 a56678a <=( A301  and  (not A300) );
 a56679a <=( a56678a  and  a56675a );
 a56680a <=( a56679a  and  a56672a );
 a56684a <=( (not A168)  and  (not A169) );
 a56685a <=( (not A170)  and  a56684a );
 a56689a <=( (not A199)  and  (not A166) );
 a56690a <=( A167  and  a56689a );
 a56691a <=( a56690a  and  a56685a );
 a56695a <=( A266  and  (not A265) );
 a56696a <=( (not A200)  and  a56695a );
 a56699a <=( (not A269)  and  A267 );
 a56702a <=( (not A302)  and  (not A300) );
 a56703a <=( a56702a  and  a56699a );
 a56704a <=( a56703a  and  a56696a );
 a56708a <=( (not A168)  and  (not A169) );
 a56709a <=( (not A170)  and  a56708a );
 a56713a <=( (not A199)  and  (not A166) );
 a56714a <=( A167  and  a56713a );
 a56715a <=( a56714a  and  a56709a );
 a56719a <=( A266  and  (not A265) );
 a56720a <=( (not A200)  and  a56719a );
 a56723a <=( (not A269)  and  A267 );
 a56726a <=( A299  and  A298 );
 a56727a <=( a56726a  and  a56723a );
 a56728a <=( a56727a  and  a56720a );
 a56732a <=( (not A168)  and  (not A169) );
 a56733a <=( (not A170)  and  a56732a );
 a56737a <=( (not A199)  and  (not A166) );
 a56738a <=( A167  and  a56737a );
 a56739a <=( a56738a  and  a56733a );
 a56743a <=( A266  and  (not A265) );
 a56744a <=( (not A200)  and  a56743a );
 a56747a <=( (not A269)  and  A267 );
 a56750a <=( (not A299)  and  (not A298) );
 a56751a <=( a56750a  and  a56747a );
 a56752a <=( a56751a  and  a56744a );
 a56756a <=( (not A168)  and  (not A169) );
 a56757a <=( (not A170)  and  a56756a );
 a56761a <=( (not A199)  and  (not A166) );
 a56762a <=( A167  and  a56761a );
 a56763a <=( a56762a  and  a56757a );
 a56767a <=( (not A266)  and  A265 );
 a56768a <=( (not A200)  and  a56767a );
 a56771a <=( A268  and  A267 );
 a56774a <=( A301  and  (not A300) );
 a56775a <=( a56774a  and  a56771a );
 a56776a <=( a56775a  and  a56768a );
 a56780a <=( (not A168)  and  (not A169) );
 a56781a <=( (not A170)  and  a56780a );
 a56785a <=( (not A199)  and  (not A166) );
 a56786a <=( A167  and  a56785a );
 a56787a <=( a56786a  and  a56781a );
 a56791a <=( (not A266)  and  A265 );
 a56792a <=( (not A200)  and  a56791a );
 a56795a <=( A268  and  A267 );
 a56798a <=( (not A302)  and  (not A300) );
 a56799a <=( a56798a  and  a56795a );
 a56800a <=( a56799a  and  a56792a );
 a56804a <=( (not A168)  and  (not A169) );
 a56805a <=( (not A170)  and  a56804a );
 a56809a <=( (not A199)  and  (not A166) );
 a56810a <=( A167  and  a56809a );
 a56811a <=( a56810a  and  a56805a );
 a56815a <=( (not A266)  and  A265 );
 a56816a <=( (not A200)  and  a56815a );
 a56819a <=( A268  and  A267 );
 a56822a <=( A299  and  A298 );
 a56823a <=( a56822a  and  a56819a );
 a56824a <=( a56823a  and  a56816a );
 a56828a <=( (not A168)  and  (not A169) );
 a56829a <=( (not A170)  and  a56828a );
 a56833a <=( (not A199)  and  (not A166) );
 a56834a <=( A167  and  a56833a );
 a56835a <=( a56834a  and  a56829a );
 a56839a <=( (not A266)  and  A265 );
 a56840a <=( (not A200)  and  a56839a );
 a56843a <=( A268  and  A267 );
 a56846a <=( (not A299)  and  (not A298) );
 a56847a <=( a56846a  and  a56843a );
 a56848a <=( a56847a  and  a56840a );
 a56852a <=( (not A168)  and  (not A169) );
 a56853a <=( (not A170)  and  a56852a );
 a56857a <=( (not A199)  and  (not A166) );
 a56858a <=( A167  and  a56857a );
 a56859a <=( a56858a  and  a56853a );
 a56863a <=( (not A266)  and  A265 );
 a56864a <=( (not A200)  and  a56863a );
 a56867a <=( (not A269)  and  A267 );
 a56870a <=( A301  and  (not A300) );
 a56871a <=( a56870a  and  a56867a );
 a56872a <=( a56871a  and  a56864a );
 a56876a <=( (not A168)  and  (not A169) );
 a56877a <=( (not A170)  and  a56876a );
 a56881a <=( (not A199)  and  (not A166) );
 a56882a <=( A167  and  a56881a );
 a56883a <=( a56882a  and  a56877a );
 a56887a <=( (not A266)  and  A265 );
 a56888a <=( (not A200)  and  a56887a );
 a56891a <=( (not A269)  and  A267 );
 a56894a <=( (not A302)  and  (not A300) );
 a56895a <=( a56894a  and  a56891a );
 a56896a <=( a56895a  and  a56888a );
 a56900a <=( (not A168)  and  (not A169) );
 a56901a <=( (not A170)  and  a56900a );
 a56905a <=( (not A199)  and  (not A166) );
 a56906a <=( A167  and  a56905a );
 a56907a <=( a56906a  and  a56901a );
 a56911a <=( (not A266)  and  A265 );
 a56912a <=( (not A200)  and  a56911a );
 a56915a <=( (not A269)  and  A267 );
 a56918a <=( A299  and  A298 );
 a56919a <=( a56918a  and  a56915a );
 a56920a <=( a56919a  and  a56912a );
 a56924a <=( (not A168)  and  (not A169) );
 a56925a <=( (not A170)  and  a56924a );
 a56929a <=( (not A199)  and  (not A166) );
 a56930a <=( A167  and  a56929a );
 a56931a <=( a56930a  and  a56925a );
 a56935a <=( (not A266)  and  A265 );
 a56936a <=( (not A200)  and  a56935a );
 a56939a <=( (not A269)  and  A267 );
 a56942a <=( (not A299)  and  (not A298) );
 a56943a <=( a56942a  and  a56939a );
 a56944a <=( a56943a  and  a56936a );
 a56948a <=( (not A168)  and  (not A169) );
 a56949a <=( (not A170)  and  a56948a );
 a56953a <=( (not A199)  and  (not A166) );
 a56954a <=( A167  and  a56953a );
 a56955a <=( a56954a  and  a56949a );
 a56959a <=( (not A266)  and  (not A265) );
 a56960a <=( (not A200)  and  a56959a );
 a56963a <=( (not A299)  and  A298 );
 a56966a <=( A301  and  A300 );
 a56967a <=( a56966a  and  a56963a );
 a56968a <=( a56967a  and  a56960a );
 a56972a <=( (not A168)  and  (not A169) );
 a56973a <=( (not A170)  and  a56972a );
 a56977a <=( (not A199)  and  (not A166) );
 a56978a <=( A167  and  a56977a );
 a56979a <=( a56978a  and  a56973a );
 a56983a <=( (not A266)  and  (not A265) );
 a56984a <=( (not A200)  and  a56983a );
 a56987a <=( (not A299)  and  A298 );
 a56990a <=( (not A302)  and  A300 );
 a56991a <=( a56990a  and  a56987a );
 a56992a <=( a56991a  and  a56984a );
 a56996a <=( (not A168)  and  (not A169) );
 a56997a <=( (not A170)  and  a56996a );
 a57001a <=( (not A199)  and  (not A166) );
 a57002a <=( A167  and  a57001a );
 a57003a <=( a57002a  and  a56997a );
 a57007a <=( (not A266)  and  (not A265) );
 a57008a <=( (not A200)  and  a57007a );
 a57011a <=( A299  and  (not A298) );
 a57014a <=( A301  and  A300 );
 a57015a <=( a57014a  and  a57011a );
 a57016a <=( a57015a  and  a57008a );
 a57020a <=( (not A168)  and  (not A169) );
 a57021a <=( (not A170)  and  a57020a );
 a57025a <=( (not A199)  and  (not A166) );
 a57026a <=( A167  and  a57025a );
 a57027a <=( a57026a  and  a57021a );
 a57031a <=( (not A266)  and  (not A265) );
 a57032a <=( (not A200)  and  a57031a );
 a57035a <=( A299  and  (not A298) );
 a57038a <=( (not A302)  and  A300 );
 a57039a <=( a57038a  and  a57035a );
 a57040a <=( a57039a  and  a57032a );
 a57044a <=( (not A168)  and  (not A169) );
 a57045a <=( (not A170)  and  a57044a );
 a57049a <=( (not A201)  and  A166 );
 a57050a <=( (not A167)  and  a57049a );
 a57051a <=( a57050a  and  a57045a );
 a57055a <=( A268  and  (not A267) );
 a57056a <=( A202  and  a57055a );
 a57059a <=( (not A299)  and  A298 );
 a57062a <=( A301  and  A300 );
 a57063a <=( a57062a  and  a57059a );
 a57064a <=( a57063a  and  a57056a );
 a57068a <=( (not A168)  and  (not A169) );
 a57069a <=( (not A170)  and  a57068a );
 a57073a <=( (not A201)  and  A166 );
 a57074a <=( (not A167)  and  a57073a );
 a57075a <=( a57074a  and  a57069a );
 a57079a <=( A268  and  (not A267) );
 a57080a <=( A202  and  a57079a );
 a57083a <=( (not A299)  and  A298 );
 a57086a <=( (not A302)  and  A300 );
 a57087a <=( a57086a  and  a57083a );
 a57088a <=( a57087a  and  a57080a );
 a57092a <=( (not A168)  and  (not A169) );
 a57093a <=( (not A170)  and  a57092a );
 a57097a <=( (not A201)  and  A166 );
 a57098a <=( (not A167)  and  a57097a );
 a57099a <=( a57098a  and  a57093a );
 a57103a <=( A268  and  (not A267) );
 a57104a <=( A202  and  a57103a );
 a57107a <=( A299  and  (not A298) );
 a57110a <=( A301  and  A300 );
 a57111a <=( a57110a  and  a57107a );
 a57112a <=( a57111a  and  a57104a );
 a57116a <=( (not A168)  and  (not A169) );
 a57117a <=( (not A170)  and  a57116a );
 a57121a <=( (not A201)  and  A166 );
 a57122a <=( (not A167)  and  a57121a );
 a57123a <=( a57122a  and  a57117a );
 a57127a <=( A268  and  (not A267) );
 a57128a <=( A202  and  a57127a );
 a57131a <=( A299  and  (not A298) );
 a57134a <=( (not A302)  and  A300 );
 a57135a <=( a57134a  and  a57131a );
 a57136a <=( a57135a  and  a57128a );
 a57140a <=( (not A168)  and  (not A169) );
 a57141a <=( (not A170)  and  a57140a );
 a57145a <=( (not A201)  and  A166 );
 a57146a <=( (not A167)  and  a57145a );
 a57147a <=( a57146a  and  a57141a );
 a57151a <=( (not A269)  and  (not A267) );
 a57152a <=( A202  and  a57151a );
 a57155a <=( (not A299)  and  A298 );
 a57158a <=( A301  and  A300 );
 a57159a <=( a57158a  and  a57155a );
 a57160a <=( a57159a  and  a57152a );
 a57164a <=( (not A168)  and  (not A169) );
 a57165a <=( (not A170)  and  a57164a );
 a57169a <=( (not A201)  and  A166 );
 a57170a <=( (not A167)  and  a57169a );
 a57171a <=( a57170a  and  a57165a );
 a57175a <=( (not A269)  and  (not A267) );
 a57176a <=( A202  and  a57175a );
 a57179a <=( (not A299)  and  A298 );
 a57182a <=( (not A302)  and  A300 );
 a57183a <=( a57182a  and  a57179a );
 a57184a <=( a57183a  and  a57176a );
 a57188a <=( (not A168)  and  (not A169) );
 a57189a <=( (not A170)  and  a57188a );
 a57193a <=( (not A201)  and  A166 );
 a57194a <=( (not A167)  and  a57193a );
 a57195a <=( a57194a  and  a57189a );
 a57199a <=( (not A269)  and  (not A267) );
 a57200a <=( A202  and  a57199a );
 a57203a <=( A299  and  (not A298) );
 a57206a <=( A301  and  A300 );
 a57207a <=( a57206a  and  a57203a );
 a57208a <=( a57207a  and  a57200a );
 a57212a <=( (not A168)  and  (not A169) );
 a57213a <=( (not A170)  and  a57212a );
 a57217a <=( (not A201)  and  A166 );
 a57218a <=( (not A167)  and  a57217a );
 a57219a <=( a57218a  and  a57213a );
 a57223a <=( (not A269)  and  (not A267) );
 a57224a <=( A202  and  a57223a );
 a57227a <=( A299  and  (not A298) );
 a57230a <=( (not A302)  and  A300 );
 a57231a <=( a57230a  and  a57227a );
 a57232a <=( a57231a  and  a57224a );
 a57236a <=( (not A168)  and  (not A169) );
 a57237a <=( (not A170)  and  a57236a );
 a57241a <=( (not A201)  and  A166 );
 a57242a <=( (not A167)  and  a57241a );
 a57243a <=( a57242a  and  a57237a );
 a57247a <=( A266  and  A265 );
 a57248a <=( A202  and  a57247a );
 a57251a <=( (not A299)  and  A298 );
 a57254a <=( A301  and  A300 );
 a57255a <=( a57254a  and  a57251a );
 a57256a <=( a57255a  and  a57248a );
 a57260a <=( (not A168)  and  (not A169) );
 a57261a <=( (not A170)  and  a57260a );
 a57265a <=( (not A201)  and  A166 );
 a57266a <=( (not A167)  and  a57265a );
 a57267a <=( a57266a  and  a57261a );
 a57271a <=( A266  and  A265 );
 a57272a <=( A202  and  a57271a );
 a57275a <=( (not A299)  and  A298 );
 a57278a <=( (not A302)  and  A300 );
 a57279a <=( a57278a  and  a57275a );
 a57280a <=( a57279a  and  a57272a );
 a57284a <=( (not A168)  and  (not A169) );
 a57285a <=( (not A170)  and  a57284a );
 a57289a <=( (not A201)  and  A166 );
 a57290a <=( (not A167)  and  a57289a );
 a57291a <=( a57290a  and  a57285a );
 a57295a <=( A266  and  A265 );
 a57296a <=( A202  and  a57295a );
 a57299a <=( A299  and  (not A298) );
 a57302a <=( A301  and  A300 );
 a57303a <=( a57302a  and  a57299a );
 a57304a <=( a57303a  and  a57296a );
 a57308a <=( (not A168)  and  (not A169) );
 a57309a <=( (not A170)  and  a57308a );
 a57313a <=( (not A201)  and  A166 );
 a57314a <=( (not A167)  and  a57313a );
 a57315a <=( a57314a  and  a57309a );
 a57319a <=( A266  and  A265 );
 a57320a <=( A202  and  a57319a );
 a57323a <=( A299  and  (not A298) );
 a57326a <=( (not A302)  and  A300 );
 a57327a <=( a57326a  and  a57323a );
 a57328a <=( a57327a  and  a57320a );
 a57332a <=( (not A168)  and  (not A169) );
 a57333a <=( (not A170)  and  a57332a );
 a57337a <=( (not A201)  and  A166 );
 a57338a <=( (not A167)  and  a57337a );
 a57339a <=( a57338a  and  a57333a );
 a57343a <=( A266  and  (not A265) );
 a57344a <=( A202  and  a57343a );
 a57347a <=( A268  and  A267 );
 a57350a <=( A301  and  (not A300) );
 a57351a <=( a57350a  and  a57347a );
 a57352a <=( a57351a  and  a57344a );
 a57356a <=( (not A168)  and  (not A169) );
 a57357a <=( (not A170)  and  a57356a );
 a57361a <=( (not A201)  and  A166 );
 a57362a <=( (not A167)  and  a57361a );
 a57363a <=( a57362a  and  a57357a );
 a57367a <=( A266  and  (not A265) );
 a57368a <=( A202  and  a57367a );
 a57371a <=( A268  and  A267 );
 a57374a <=( (not A302)  and  (not A300) );
 a57375a <=( a57374a  and  a57371a );
 a57376a <=( a57375a  and  a57368a );
 a57380a <=( (not A168)  and  (not A169) );
 a57381a <=( (not A170)  and  a57380a );
 a57385a <=( (not A201)  and  A166 );
 a57386a <=( (not A167)  and  a57385a );
 a57387a <=( a57386a  and  a57381a );
 a57391a <=( A266  and  (not A265) );
 a57392a <=( A202  and  a57391a );
 a57395a <=( A268  and  A267 );
 a57398a <=( A299  and  A298 );
 a57399a <=( a57398a  and  a57395a );
 a57400a <=( a57399a  and  a57392a );
 a57404a <=( (not A168)  and  (not A169) );
 a57405a <=( (not A170)  and  a57404a );
 a57409a <=( (not A201)  and  A166 );
 a57410a <=( (not A167)  and  a57409a );
 a57411a <=( a57410a  and  a57405a );
 a57415a <=( A266  and  (not A265) );
 a57416a <=( A202  and  a57415a );
 a57419a <=( A268  and  A267 );
 a57422a <=( (not A299)  and  (not A298) );
 a57423a <=( a57422a  and  a57419a );
 a57424a <=( a57423a  and  a57416a );
 a57428a <=( (not A168)  and  (not A169) );
 a57429a <=( (not A170)  and  a57428a );
 a57433a <=( (not A201)  and  A166 );
 a57434a <=( (not A167)  and  a57433a );
 a57435a <=( a57434a  and  a57429a );
 a57439a <=( A266  and  (not A265) );
 a57440a <=( A202  and  a57439a );
 a57443a <=( (not A269)  and  A267 );
 a57446a <=( A301  and  (not A300) );
 a57447a <=( a57446a  and  a57443a );
 a57448a <=( a57447a  and  a57440a );
 a57452a <=( (not A168)  and  (not A169) );
 a57453a <=( (not A170)  and  a57452a );
 a57457a <=( (not A201)  and  A166 );
 a57458a <=( (not A167)  and  a57457a );
 a57459a <=( a57458a  and  a57453a );
 a57463a <=( A266  and  (not A265) );
 a57464a <=( A202  and  a57463a );
 a57467a <=( (not A269)  and  A267 );
 a57470a <=( (not A302)  and  (not A300) );
 a57471a <=( a57470a  and  a57467a );
 a57472a <=( a57471a  and  a57464a );
 a57476a <=( (not A168)  and  (not A169) );
 a57477a <=( (not A170)  and  a57476a );
 a57481a <=( (not A201)  and  A166 );
 a57482a <=( (not A167)  and  a57481a );
 a57483a <=( a57482a  and  a57477a );
 a57487a <=( A266  and  (not A265) );
 a57488a <=( A202  and  a57487a );
 a57491a <=( (not A269)  and  A267 );
 a57494a <=( A299  and  A298 );
 a57495a <=( a57494a  and  a57491a );
 a57496a <=( a57495a  and  a57488a );
 a57500a <=( (not A168)  and  (not A169) );
 a57501a <=( (not A170)  and  a57500a );
 a57505a <=( (not A201)  and  A166 );
 a57506a <=( (not A167)  and  a57505a );
 a57507a <=( a57506a  and  a57501a );
 a57511a <=( A266  and  (not A265) );
 a57512a <=( A202  and  a57511a );
 a57515a <=( (not A269)  and  A267 );
 a57518a <=( (not A299)  and  (not A298) );
 a57519a <=( a57518a  and  a57515a );
 a57520a <=( a57519a  and  a57512a );
 a57524a <=( (not A168)  and  (not A169) );
 a57525a <=( (not A170)  and  a57524a );
 a57529a <=( (not A201)  and  A166 );
 a57530a <=( (not A167)  and  a57529a );
 a57531a <=( a57530a  and  a57525a );
 a57535a <=( (not A266)  and  A265 );
 a57536a <=( A202  and  a57535a );
 a57539a <=( A268  and  A267 );
 a57542a <=( A301  and  (not A300) );
 a57543a <=( a57542a  and  a57539a );
 a57544a <=( a57543a  and  a57536a );
 a57548a <=( (not A168)  and  (not A169) );
 a57549a <=( (not A170)  and  a57548a );
 a57553a <=( (not A201)  and  A166 );
 a57554a <=( (not A167)  and  a57553a );
 a57555a <=( a57554a  and  a57549a );
 a57559a <=( (not A266)  and  A265 );
 a57560a <=( A202  and  a57559a );
 a57563a <=( A268  and  A267 );
 a57566a <=( (not A302)  and  (not A300) );
 a57567a <=( a57566a  and  a57563a );
 a57568a <=( a57567a  and  a57560a );
 a57572a <=( (not A168)  and  (not A169) );
 a57573a <=( (not A170)  and  a57572a );
 a57577a <=( (not A201)  and  A166 );
 a57578a <=( (not A167)  and  a57577a );
 a57579a <=( a57578a  and  a57573a );
 a57583a <=( (not A266)  and  A265 );
 a57584a <=( A202  and  a57583a );
 a57587a <=( A268  and  A267 );
 a57590a <=( A299  and  A298 );
 a57591a <=( a57590a  and  a57587a );
 a57592a <=( a57591a  and  a57584a );
 a57596a <=( (not A168)  and  (not A169) );
 a57597a <=( (not A170)  and  a57596a );
 a57601a <=( (not A201)  and  A166 );
 a57602a <=( (not A167)  and  a57601a );
 a57603a <=( a57602a  and  a57597a );
 a57607a <=( (not A266)  and  A265 );
 a57608a <=( A202  and  a57607a );
 a57611a <=( A268  and  A267 );
 a57614a <=( (not A299)  and  (not A298) );
 a57615a <=( a57614a  and  a57611a );
 a57616a <=( a57615a  and  a57608a );
 a57620a <=( (not A168)  and  (not A169) );
 a57621a <=( (not A170)  and  a57620a );
 a57625a <=( (not A201)  and  A166 );
 a57626a <=( (not A167)  and  a57625a );
 a57627a <=( a57626a  and  a57621a );
 a57631a <=( (not A266)  and  A265 );
 a57632a <=( A202  and  a57631a );
 a57635a <=( (not A269)  and  A267 );
 a57638a <=( A301  and  (not A300) );
 a57639a <=( a57638a  and  a57635a );
 a57640a <=( a57639a  and  a57632a );
 a57644a <=( (not A168)  and  (not A169) );
 a57645a <=( (not A170)  and  a57644a );
 a57649a <=( (not A201)  and  A166 );
 a57650a <=( (not A167)  and  a57649a );
 a57651a <=( a57650a  and  a57645a );
 a57655a <=( (not A266)  and  A265 );
 a57656a <=( A202  and  a57655a );
 a57659a <=( (not A269)  and  A267 );
 a57662a <=( (not A302)  and  (not A300) );
 a57663a <=( a57662a  and  a57659a );
 a57664a <=( a57663a  and  a57656a );
 a57668a <=( (not A168)  and  (not A169) );
 a57669a <=( (not A170)  and  a57668a );
 a57673a <=( (not A201)  and  A166 );
 a57674a <=( (not A167)  and  a57673a );
 a57675a <=( a57674a  and  a57669a );
 a57679a <=( (not A266)  and  A265 );
 a57680a <=( A202  and  a57679a );
 a57683a <=( (not A269)  and  A267 );
 a57686a <=( A299  and  A298 );
 a57687a <=( a57686a  and  a57683a );
 a57688a <=( a57687a  and  a57680a );
 a57692a <=( (not A168)  and  (not A169) );
 a57693a <=( (not A170)  and  a57692a );
 a57697a <=( (not A201)  and  A166 );
 a57698a <=( (not A167)  and  a57697a );
 a57699a <=( a57698a  and  a57693a );
 a57703a <=( (not A266)  and  A265 );
 a57704a <=( A202  and  a57703a );
 a57707a <=( (not A269)  and  A267 );
 a57710a <=( (not A299)  and  (not A298) );
 a57711a <=( a57710a  and  a57707a );
 a57712a <=( a57711a  and  a57704a );
 a57716a <=( (not A168)  and  (not A169) );
 a57717a <=( (not A170)  and  a57716a );
 a57721a <=( (not A201)  and  A166 );
 a57722a <=( (not A167)  and  a57721a );
 a57723a <=( a57722a  and  a57717a );
 a57727a <=( (not A266)  and  (not A265) );
 a57728a <=( A202  and  a57727a );
 a57731a <=( (not A299)  and  A298 );
 a57734a <=( A301  and  A300 );
 a57735a <=( a57734a  and  a57731a );
 a57736a <=( a57735a  and  a57728a );
 a57740a <=( (not A168)  and  (not A169) );
 a57741a <=( (not A170)  and  a57740a );
 a57745a <=( (not A201)  and  A166 );
 a57746a <=( (not A167)  and  a57745a );
 a57747a <=( a57746a  and  a57741a );
 a57751a <=( (not A266)  and  (not A265) );
 a57752a <=( A202  and  a57751a );
 a57755a <=( (not A299)  and  A298 );
 a57758a <=( (not A302)  and  A300 );
 a57759a <=( a57758a  and  a57755a );
 a57760a <=( a57759a  and  a57752a );
 a57764a <=( (not A168)  and  (not A169) );
 a57765a <=( (not A170)  and  a57764a );
 a57769a <=( (not A201)  and  A166 );
 a57770a <=( (not A167)  and  a57769a );
 a57771a <=( a57770a  and  a57765a );
 a57775a <=( (not A266)  and  (not A265) );
 a57776a <=( A202  and  a57775a );
 a57779a <=( A299  and  (not A298) );
 a57782a <=( A301  and  A300 );
 a57783a <=( a57782a  and  a57779a );
 a57784a <=( a57783a  and  a57776a );
 a57788a <=( (not A168)  and  (not A169) );
 a57789a <=( (not A170)  and  a57788a );
 a57793a <=( (not A201)  and  A166 );
 a57794a <=( (not A167)  and  a57793a );
 a57795a <=( a57794a  and  a57789a );
 a57799a <=( (not A266)  and  (not A265) );
 a57800a <=( A202  and  a57799a );
 a57803a <=( A299  and  (not A298) );
 a57806a <=( (not A302)  and  A300 );
 a57807a <=( a57806a  and  a57803a );
 a57808a <=( a57807a  and  a57800a );
 a57812a <=( (not A168)  and  (not A169) );
 a57813a <=( (not A170)  and  a57812a );
 a57817a <=( (not A201)  and  A166 );
 a57818a <=( (not A167)  and  a57817a );
 a57819a <=( a57818a  and  a57813a );
 a57823a <=( A268  and  (not A267) );
 a57824a <=( (not A203)  and  a57823a );
 a57827a <=( (not A299)  and  A298 );
 a57830a <=( A301  and  A300 );
 a57831a <=( a57830a  and  a57827a );
 a57832a <=( a57831a  and  a57824a );
 a57836a <=( (not A168)  and  (not A169) );
 a57837a <=( (not A170)  and  a57836a );
 a57841a <=( (not A201)  and  A166 );
 a57842a <=( (not A167)  and  a57841a );
 a57843a <=( a57842a  and  a57837a );
 a57847a <=( A268  and  (not A267) );
 a57848a <=( (not A203)  and  a57847a );
 a57851a <=( (not A299)  and  A298 );
 a57854a <=( (not A302)  and  A300 );
 a57855a <=( a57854a  and  a57851a );
 a57856a <=( a57855a  and  a57848a );
 a57860a <=( (not A168)  and  (not A169) );
 a57861a <=( (not A170)  and  a57860a );
 a57865a <=( (not A201)  and  A166 );
 a57866a <=( (not A167)  and  a57865a );
 a57867a <=( a57866a  and  a57861a );
 a57871a <=( A268  and  (not A267) );
 a57872a <=( (not A203)  and  a57871a );
 a57875a <=( A299  and  (not A298) );
 a57878a <=( A301  and  A300 );
 a57879a <=( a57878a  and  a57875a );
 a57880a <=( a57879a  and  a57872a );
 a57884a <=( (not A168)  and  (not A169) );
 a57885a <=( (not A170)  and  a57884a );
 a57889a <=( (not A201)  and  A166 );
 a57890a <=( (not A167)  and  a57889a );
 a57891a <=( a57890a  and  a57885a );
 a57895a <=( A268  and  (not A267) );
 a57896a <=( (not A203)  and  a57895a );
 a57899a <=( A299  and  (not A298) );
 a57902a <=( (not A302)  and  A300 );
 a57903a <=( a57902a  and  a57899a );
 a57904a <=( a57903a  and  a57896a );
 a57908a <=( (not A168)  and  (not A169) );
 a57909a <=( (not A170)  and  a57908a );
 a57913a <=( (not A201)  and  A166 );
 a57914a <=( (not A167)  and  a57913a );
 a57915a <=( a57914a  and  a57909a );
 a57919a <=( (not A269)  and  (not A267) );
 a57920a <=( (not A203)  and  a57919a );
 a57923a <=( (not A299)  and  A298 );
 a57926a <=( A301  and  A300 );
 a57927a <=( a57926a  and  a57923a );
 a57928a <=( a57927a  and  a57920a );
 a57932a <=( (not A168)  and  (not A169) );
 a57933a <=( (not A170)  and  a57932a );
 a57937a <=( (not A201)  and  A166 );
 a57938a <=( (not A167)  and  a57937a );
 a57939a <=( a57938a  and  a57933a );
 a57943a <=( (not A269)  and  (not A267) );
 a57944a <=( (not A203)  and  a57943a );
 a57947a <=( (not A299)  and  A298 );
 a57950a <=( (not A302)  and  A300 );
 a57951a <=( a57950a  and  a57947a );
 a57952a <=( a57951a  and  a57944a );
 a57956a <=( (not A168)  and  (not A169) );
 a57957a <=( (not A170)  and  a57956a );
 a57961a <=( (not A201)  and  A166 );
 a57962a <=( (not A167)  and  a57961a );
 a57963a <=( a57962a  and  a57957a );
 a57967a <=( (not A269)  and  (not A267) );
 a57968a <=( (not A203)  and  a57967a );
 a57971a <=( A299  and  (not A298) );
 a57974a <=( A301  and  A300 );
 a57975a <=( a57974a  and  a57971a );
 a57976a <=( a57975a  and  a57968a );
 a57980a <=( (not A168)  and  (not A169) );
 a57981a <=( (not A170)  and  a57980a );
 a57985a <=( (not A201)  and  A166 );
 a57986a <=( (not A167)  and  a57985a );
 a57987a <=( a57986a  and  a57981a );
 a57991a <=( (not A269)  and  (not A267) );
 a57992a <=( (not A203)  and  a57991a );
 a57995a <=( A299  and  (not A298) );
 a57998a <=( (not A302)  and  A300 );
 a57999a <=( a57998a  and  a57995a );
 a58000a <=( a57999a  and  a57992a );
 a58004a <=( (not A168)  and  (not A169) );
 a58005a <=( (not A170)  and  a58004a );
 a58009a <=( (not A201)  and  A166 );
 a58010a <=( (not A167)  and  a58009a );
 a58011a <=( a58010a  and  a58005a );
 a58015a <=( A266  and  A265 );
 a58016a <=( (not A203)  and  a58015a );
 a58019a <=( (not A299)  and  A298 );
 a58022a <=( A301  and  A300 );
 a58023a <=( a58022a  and  a58019a );
 a58024a <=( a58023a  and  a58016a );
 a58028a <=( (not A168)  and  (not A169) );
 a58029a <=( (not A170)  and  a58028a );
 a58033a <=( (not A201)  and  A166 );
 a58034a <=( (not A167)  and  a58033a );
 a58035a <=( a58034a  and  a58029a );
 a58039a <=( A266  and  A265 );
 a58040a <=( (not A203)  and  a58039a );
 a58043a <=( (not A299)  and  A298 );
 a58046a <=( (not A302)  and  A300 );
 a58047a <=( a58046a  and  a58043a );
 a58048a <=( a58047a  and  a58040a );
 a58052a <=( (not A168)  and  (not A169) );
 a58053a <=( (not A170)  and  a58052a );
 a58057a <=( (not A201)  and  A166 );
 a58058a <=( (not A167)  and  a58057a );
 a58059a <=( a58058a  and  a58053a );
 a58063a <=( A266  and  A265 );
 a58064a <=( (not A203)  and  a58063a );
 a58067a <=( A299  and  (not A298) );
 a58070a <=( A301  and  A300 );
 a58071a <=( a58070a  and  a58067a );
 a58072a <=( a58071a  and  a58064a );
 a58076a <=( (not A168)  and  (not A169) );
 a58077a <=( (not A170)  and  a58076a );
 a58081a <=( (not A201)  and  A166 );
 a58082a <=( (not A167)  and  a58081a );
 a58083a <=( a58082a  and  a58077a );
 a58087a <=( A266  and  A265 );
 a58088a <=( (not A203)  and  a58087a );
 a58091a <=( A299  and  (not A298) );
 a58094a <=( (not A302)  and  A300 );
 a58095a <=( a58094a  and  a58091a );
 a58096a <=( a58095a  and  a58088a );
 a58100a <=( (not A168)  and  (not A169) );
 a58101a <=( (not A170)  and  a58100a );
 a58105a <=( (not A201)  and  A166 );
 a58106a <=( (not A167)  and  a58105a );
 a58107a <=( a58106a  and  a58101a );
 a58111a <=( A266  and  (not A265) );
 a58112a <=( (not A203)  and  a58111a );
 a58115a <=( A268  and  A267 );
 a58118a <=( A301  and  (not A300) );
 a58119a <=( a58118a  and  a58115a );
 a58120a <=( a58119a  and  a58112a );
 a58124a <=( (not A168)  and  (not A169) );
 a58125a <=( (not A170)  and  a58124a );
 a58129a <=( (not A201)  and  A166 );
 a58130a <=( (not A167)  and  a58129a );
 a58131a <=( a58130a  and  a58125a );
 a58135a <=( A266  and  (not A265) );
 a58136a <=( (not A203)  and  a58135a );
 a58139a <=( A268  and  A267 );
 a58142a <=( (not A302)  and  (not A300) );
 a58143a <=( a58142a  and  a58139a );
 a58144a <=( a58143a  and  a58136a );
 a58148a <=( (not A168)  and  (not A169) );
 a58149a <=( (not A170)  and  a58148a );
 a58153a <=( (not A201)  and  A166 );
 a58154a <=( (not A167)  and  a58153a );
 a58155a <=( a58154a  and  a58149a );
 a58159a <=( A266  and  (not A265) );
 a58160a <=( (not A203)  and  a58159a );
 a58163a <=( A268  and  A267 );
 a58166a <=( A299  and  A298 );
 a58167a <=( a58166a  and  a58163a );
 a58168a <=( a58167a  and  a58160a );
 a58172a <=( (not A168)  and  (not A169) );
 a58173a <=( (not A170)  and  a58172a );
 a58177a <=( (not A201)  and  A166 );
 a58178a <=( (not A167)  and  a58177a );
 a58179a <=( a58178a  and  a58173a );
 a58183a <=( A266  and  (not A265) );
 a58184a <=( (not A203)  and  a58183a );
 a58187a <=( A268  and  A267 );
 a58190a <=( (not A299)  and  (not A298) );
 a58191a <=( a58190a  and  a58187a );
 a58192a <=( a58191a  and  a58184a );
 a58196a <=( (not A168)  and  (not A169) );
 a58197a <=( (not A170)  and  a58196a );
 a58201a <=( (not A201)  and  A166 );
 a58202a <=( (not A167)  and  a58201a );
 a58203a <=( a58202a  and  a58197a );
 a58207a <=( A266  and  (not A265) );
 a58208a <=( (not A203)  and  a58207a );
 a58211a <=( (not A269)  and  A267 );
 a58214a <=( A301  and  (not A300) );
 a58215a <=( a58214a  and  a58211a );
 a58216a <=( a58215a  and  a58208a );
 a58220a <=( (not A168)  and  (not A169) );
 a58221a <=( (not A170)  and  a58220a );
 a58225a <=( (not A201)  and  A166 );
 a58226a <=( (not A167)  and  a58225a );
 a58227a <=( a58226a  and  a58221a );
 a58231a <=( A266  and  (not A265) );
 a58232a <=( (not A203)  and  a58231a );
 a58235a <=( (not A269)  and  A267 );
 a58238a <=( (not A302)  and  (not A300) );
 a58239a <=( a58238a  and  a58235a );
 a58240a <=( a58239a  and  a58232a );
 a58244a <=( (not A168)  and  (not A169) );
 a58245a <=( (not A170)  and  a58244a );
 a58249a <=( (not A201)  and  A166 );
 a58250a <=( (not A167)  and  a58249a );
 a58251a <=( a58250a  and  a58245a );
 a58255a <=( A266  and  (not A265) );
 a58256a <=( (not A203)  and  a58255a );
 a58259a <=( (not A269)  and  A267 );
 a58262a <=( A299  and  A298 );
 a58263a <=( a58262a  and  a58259a );
 a58264a <=( a58263a  and  a58256a );
 a58268a <=( (not A168)  and  (not A169) );
 a58269a <=( (not A170)  and  a58268a );
 a58273a <=( (not A201)  and  A166 );
 a58274a <=( (not A167)  and  a58273a );
 a58275a <=( a58274a  and  a58269a );
 a58279a <=( A266  and  (not A265) );
 a58280a <=( (not A203)  and  a58279a );
 a58283a <=( (not A269)  and  A267 );
 a58286a <=( (not A299)  and  (not A298) );
 a58287a <=( a58286a  and  a58283a );
 a58288a <=( a58287a  and  a58280a );
 a58292a <=( (not A168)  and  (not A169) );
 a58293a <=( (not A170)  and  a58292a );
 a58297a <=( (not A201)  and  A166 );
 a58298a <=( (not A167)  and  a58297a );
 a58299a <=( a58298a  and  a58293a );
 a58303a <=( (not A266)  and  A265 );
 a58304a <=( (not A203)  and  a58303a );
 a58307a <=( A268  and  A267 );
 a58310a <=( A301  and  (not A300) );
 a58311a <=( a58310a  and  a58307a );
 a58312a <=( a58311a  and  a58304a );
 a58316a <=( (not A168)  and  (not A169) );
 a58317a <=( (not A170)  and  a58316a );
 a58321a <=( (not A201)  and  A166 );
 a58322a <=( (not A167)  and  a58321a );
 a58323a <=( a58322a  and  a58317a );
 a58327a <=( (not A266)  and  A265 );
 a58328a <=( (not A203)  and  a58327a );
 a58331a <=( A268  and  A267 );
 a58334a <=( (not A302)  and  (not A300) );
 a58335a <=( a58334a  and  a58331a );
 a58336a <=( a58335a  and  a58328a );
 a58340a <=( (not A168)  and  (not A169) );
 a58341a <=( (not A170)  and  a58340a );
 a58345a <=( (not A201)  and  A166 );
 a58346a <=( (not A167)  and  a58345a );
 a58347a <=( a58346a  and  a58341a );
 a58351a <=( (not A266)  and  A265 );
 a58352a <=( (not A203)  and  a58351a );
 a58355a <=( A268  and  A267 );
 a58358a <=( A299  and  A298 );
 a58359a <=( a58358a  and  a58355a );
 a58360a <=( a58359a  and  a58352a );
 a58364a <=( (not A168)  and  (not A169) );
 a58365a <=( (not A170)  and  a58364a );
 a58369a <=( (not A201)  and  A166 );
 a58370a <=( (not A167)  and  a58369a );
 a58371a <=( a58370a  and  a58365a );
 a58375a <=( (not A266)  and  A265 );
 a58376a <=( (not A203)  and  a58375a );
 a58379a <=( A268  and  A267 );
 a58382a <=( (not A299)  and  (not A298) );
 a58383a <=( a58382a  and  a58379a );
 a58384a <=( a58383a  and  a58376a );
 a58388a <=( (not A168)  and  (not A169) );
 a58389a <=( (not A170)  and  a58388a );
 a58393a <=( (not A201)  and  A166 );
 a58394a <=( (not A167)  and  a58393a );
 a58395a <=( a58394a  and  a58389a );
 a58399a <=( (not A266)  and  A265 );
 a58400a <=( (not A203)  and  a58399a );
 a58403a <=( (not A269)  and  A267 );
 a58406a <=( A301  and  (not A300) );
 a58407a <=( a58406a  and  a58403a );
 a58408a <=( a58407a  and  a58400a );
 a58412a <=( (not A168)  and  (not A169) );
 a58413a <=( (not A170)  and  a58412a );
 a58417a <=( (not A201)  and  A166 );
 a58418a <=( (not A167)  and  a58417a );
 a58419a <=( a58418a  and  a58413a );
 a58423a <=( (not A266)  and  A265 );
 a58424a <=( (not A203)  and  a58423a );
 a58427a <=( (not A269)  and  A267 );
 a58430a <=( (not A302)  and  (not A300) );
 a58431a <=( a58430a  and  a58427a );
 a58432a <=( a58431a  and  a58424a );
 a58436a <=( (not A168)  and  (not A169) );
 a58437a <=( (not A170)  and  a58436a );
 a58441a <=( (not A201)  and  A166 );
 a58442a <=( (not A167)  and  a58441a );
 a58443a <=( a58442a  and  a58437a );
 a58447a <=( (not A266)  and  A265 );
 a58448a <=( (not A203)  and  a58447a );
 a58451a <=( (not A269)  and  A267 );
 a58454a <=( A299  and  A298 );
 a58455a <=( a58454a  and  a58451a );
 a58456a <=( a58455a  and  a58448a );
 a58460a <=( (not A168)  and  (not A169) );
 a58461a <=( (not A170)  and  a58460a );
 a58465a <=( (not A201)  and  A166 );
 a58466a <=( (not A167)  and  a58465a );
 a58467a <=( a58466a  and  a58461a );
 a58471a <=( (not A266)  and  A265 );
 a58472a <=( (not A203)  and  a58471a );
 a58475a <=( (not A269)  and  A267 );
 a58478a <=( (not A299)  and  (not A298) );
 a58479a <=( a58478a  and  a58475a );
 a58480a <=( a58479a  and  a58472a );
 a58484a <=( (not A168)  and  (not A169) );
 a58485a <=( (not A170)  and  a58484a );
 a58489a <=( (not A201)  and  A166 );
 a58490a <=( (not A167)  and  a58489a );
 a58491a <=( a58490a  and  a58485a );
 a58495a <=( (not A266)  and  (not A265) );
 a58496a <=( (not A203)  and  a58495a );
 a58499a <=( (not A299)  and  A298 );
 a58502a <=( A301  and  A300 );
 a58503a <=( a58502a  and  a58499a );
 a58504a <=( a58503a  and  a58496a );
 a58508a <=( (not A168)  and  (not A169) );
 a58509a <=( (not A170)  and  a58508a );
 a58513a <=( (not A201)  and  A166 );
 a58514a <=( (not A167)  and  a58513a );
 a58515a <=( a58514a  and  a58509a );
 a58519a <=( (not A266)  and  (not A265) );
 a58520a <=( (not A203)  and  a58519a );
 a58523a <=( (not A299)  and  A298 );
 a58526a <=( (not A302)  and  A300 );
 a58527a <=( a58526a  and  a58523a );
 a58528a <=( a58527a  and  a58520a );
 a58532a <=( (not A168)  and  (not A169) );
 a58533a <=( (not A170)  and  a58532a );
 a58537a <=( (not A201)  and  A166 );
 a58538a <=( (not A167)  and  a58537a );
 a58539a <=( a58538a  and  a58533a );
 a58543a <=( (not A266)  and  (not A265) );
 a58544a <=( (not A203)  and  a58543a );
 a58547a <=( A299  and  (not A298) );
 a58550a <=( A301  and  A300 );
 a58551a <=( a58550a  and  a58547a );
 a58552a <=( a58551a  and  a58544a );
 a58556a <=( (not A168)  and  (not A169) );
 a58557a <=( (not A170)  and  a58556a );
 a58561a <=( (not A201)  and  A166 );
 a58562a <=( (not A167)  and  a58561a );
 a58563a <=( a58562a  and  a58557a );
 a58567a <=( (not A266)  and  (not A265) );
 a58568a <=( (not A203)  and  a58567a );
 a58571a <=( A299  and  (not A298) );
 a58574a <=( (not A302)  and  A300 );
 a58575a <=( a58574a  and  a58571a );
 a58576a <=( a58575a  and  a58568a );
 a58580a <=( (not A168)  and  (not A169) );
 a58581a <=( (not A170)  and  a58580a );
 a58585a <=( A199  and  A166 );
 a58586a <=( (not A167)  and  a58585a );
 a58587a <=( a58586a  and  a58581a );
 a58591a <=( A268  and  (not A267) );
 a58592a <=( A200  and  a58591a );
 a58595a <=( (not A299)  and  A298 );
 a58598a <=( A301  and  A300 );
 a58599a <=( a58598a  and  a58595a );
 a58600a <=( a58599a  and  a58592a );
 a58604a <=( (not A168)  and  (not A169) );
 a58605a <=( (not A170)  and  a58604a );
 a58609a <=( A199  and  A166 );
 a58610a <=( (not A167)  and  a58609a );
 a58611a <=( a58610a  and  a58605a );
 a58615a <=( A268  and  (not A267) );
 a58616a <=( A200  and  a58615a );
 a58619a <=( (not A299)  and  A298 );
 a58622a <=( (not A302)  and  A300 );
 a58623a <=( a58622a  and  a58619a );
 a58624a <=( a58623a  and  a58616a );
 a58628a <=( (not A168)  and  (not A169) );
 a58629a <=( (not A170)  and  a58628a );
 a58633a <=( A199  and  A166 );
 a58634a <=( (not A167)  and  a58633a );
 a58635a <=( a58634a  and  a58629a );
 a58639a <=( A268  and  (not A267) );
 a58640a <=( A200  and  a58639a );
 a58643a <=( A299  and  (not A298) );
 a58646a <=( A301  and  A300 );
 a58647a <=( a58646a  and  a58643a );
 a58648a <=( a58647a  and  a58640a );
 a58652a <=( (not A168)  and  (not A169) );
 a58653a <=( (not A170)  and  a58652a );
 a58657a <=( A199  and  A166 );
 a58658a <=( (not A167)  and  a58657a );
 a58659a <=( a58658a  and  a58653a );
 a58663a <=( A268  and  (not A267) );
 a58664a <=( A200  and  a58663a );
 a58667a <=( A299  and  (not A298) );
 a58670a <=( (not A302)  and  A300 );
 a58671a <=( a58670a  and  a58667a );
 a58672a <=( a58671a  and  a58664a );
 a58676a <=( (not A168)  and  (not A169) );
 a58677a <=( (not A170)  and  a58676a );
 a58681a <=( A199  and  A166 );
 a58682a <=( (not A167)  and  a58681a );
 a58683a <=( a58682a  and  a58677a );
 a58687a <=( (not A269)  and  (not A267) );
 a58688a <=( A200  and  a58687a );
 a58691a <=( (not A299)  and  A298 );
 a58694a <=( A301  and  A300 );
 a58695a <=( a58694a  and  a58691a );
 a58696a <=( a58695a  and  a58688a );
 a58700a <=( (not A168)  and  (not A169) );
 a58701a <=( (not A170)  and  a58700a );
 a58705a <=( A199  and  A166 );
 a58706a <=( (not A167)  and  a58705a );
 a58707a <=( a58706a  and  a58701a );
 a58711a <=( (not A269)  and  (not A267) );
 a58712a <=( A200  and  a58711a );
 a58715a <=( (not A299)  and  A298 );
 a58718a <=( (not A302)  and  A300 );
 a58719a <=( a58718a  and  a58715a );
 a58720a <=( a58719a  and  a58712a );
 a58724a <=( (not A168)  and  (not A169) );
 a58725a <=( (not A170)  and  a58724a );
 a58729a <=( A199  and  A166 );
 a58730a <=( (not A167)  and  a58729a );
 a58731a <=( a58730a  and  a58725a );
 a58735a <=( (not A269)  and  (not A267) );
 a58736a <=( A200  and  a58735a );
 a58739a <=( A299  and  (not A298) );
 a58742a <=( A301  and  A300 );
 a58743a <=( a58742a  and  a58739a );
 a58744a <=( a58743a  and  a58736a );
 a58748a <=( (not A168)  and  (not A169) );
 a58749a <=( (not A170)  and  a58748a );
 a58753a <=( A199  and  A166 );
 a58754a <=( (not A167)  and  a58753a );
 a58755a <=( a58754a  and  a58749a );
 a58759a <=( (not A269)  and  (not A267) );
 a58760a <=( A200  and  a58759a );
 a58763a <=( A299  and  (not A298) );
 a58766a <=( (not A302)  and  A300 );
 a58767a <=( a58766a  and  a58763a );
 a58768a <=( a58767a  and  a58760a );
 a58772a <=( (not A168)  and  (not A169) );
 a58773a <=( (not A170)  and  a58772a );
 a58777a <=( A199  and  A166 );
 a58778a <=( (not A167)  and  a58777a );
 a58779a <=( a58778a  and  a58773a );
 a58783a <=( A266  and  A265 );
 a58784a <=( A200  and  a58783a );
 a58787a <=( (not A299)  and  A298 );
 a58790a <=( A301  and  A300 );
 a58791a <=( a58790a  and  a58787a );
 a58792a <=( a58791a  and  a58784a );
 a58796a <=( (not A168)  and  (not A169) );
 a58797a <=( (not A170)  and  a58796a );
 a58801a <=( A199  and  A166 );
 a58802a <=( (not A167)  and  a58801a );
 a58803a <=( a58802a  and  a58797a );
 a58807a <=( A266  and  A265 );
 a58808a <=( A200  and  a58807a );
 a58811a <=( (not A299)  and  A298 );
 a58814a <=( (not A302)  and  A300 );
 a58815a <=( a58814a  and  a58811a );
 a58816a <=( a58815a  and  a58808a );
 a58820a <=( (not A168)  and  (not A169) );
 a58821a <=( (not A170)  and  a58820a );
 a58825a <=( A199  and  A166 );
 a58826a <=( (not A167)  and  a58825a );
 a58827a <=( a58826a  and  a58821a );
 a58831a <=( A266  and  A265 );
 a58832a <=( A200  and  a58831a );
 a58835a <=( A299  and  (not A298) );
 a58838a <=( A301  and  A300 );
 a58839a <=( a58838a  and  a58835a );
 a58840a <=( a58839a  and  a58832a );
 a58844a <=( (not A168)  and  (not A169) );
 a58845a <=( (not A170)  and  a58844a );
 a58849a <=( A199  and  A166 );
 a58850a <=( (not A167)  and  a58849a );
 a58851a <=( a58850a  and  a58845a );
 a58855a <=( A266  and  A265 );
 a58856a <=( A200  and  a58855a );
 a58859a <=( A299  and  (not A298) );
 a58862a <=( (not A302)  and  A300 );
 a58863a <=( a58862a  and  a58859a );
 a58864a <=( a58863a  and  a58856a );
 a58868a <=( (not A168)  and  (not A169) );
 a58869a <=( (not A170)  and  a58868a );
 a58873a <=( A199  and  A166 );
 a58874a <=( (not A167)  and  a58873a );
 a58875a <=( a58874a  and  a58869a );
 a58879a <=( A266  and  (not A265) );
 a58880a <=( A200  and  a58879a );
 a58883a <=( A268  and  A267 );
 a58886a <=( A301  and  (not A300) );
 a58887a <=( a58886a  and  a58883a );
 a58888a <=( a58887a  and  a58880a );
 a58892a <=( (not A168)  and  (not A169) );
 a58893a <=( (not A170)  and  a58892a );
 a58897a <=( A199  and  A166 );
 a58898a <=( (not A167)  and  a58897a );
 a58899a <=( a58898a  and  a58893a );
 a58903a <=( A266  and  (not A265) );
 a58904a <=( A200  and  a58903a );
 a58907a <=( A268  and  A267 );
 a58910a <=( (not A302)  and  (not A300) );
 a58911a <=( a58910a  and  a58907a );
 a58912a <=( a58911a  and  a58904a );
 a58916a <=( (not A168)  and  (not A169) );
 a58917a <=( (not A170)  and  a58916a );
 a58921a <=( A199  and  A166 );
 a58922a <=( (not A167)  and  a58921a );
 a58923a <=( a58922a  and  a58917a );
 a58927a <=( A266  and  (not A265) );
 a58928a <=( A200  and  a58927a );
 a58931a <=( A268  and  A267 );
 a58934a <=( A299  and  A298 );
 a58935a <=( a58934a  and  a58931a );
 a58936a <=( a58935a  and  a58928a );
 a58940a <=( (not A168)  and  (not A169) );
 a58941a <=( (not A170)  and  a58940a );
 a58945a <=( A199  and  A166 );
 a58946a <=( (not A167)  and  a58945a );
 a58947a <=( a58946a  and  a58941a );
 a58951a <=( A266  and  (not A265) );
 a58952a <=( A200  and  a58951a );
 a58955a <=( A268  and  A267 );
 a58958a <=( (not A299)  and  (not A298) );
 a58959a <=( a58958a  and  a58955a );
 a58960a <=( a58959a  and  a58952a );
 a58964a <=( (not A168)  and  (not A169) );
 a58965a <=( (not A170)  and  a58964a );
 a58969a <=( A199  and  A166 );
 a58970a <=( (not A167)  and  a58969a );
 a58971a <=( a58970a  and  a58965a );
 a58975a <=( A266  and  (not A265) );
 a58976a <=( A200  and  a58975a );
 a58979a <=( (not A269)  and  A267 );
 a58982a <=( A301  and  (not A300) );
 a58983a <=( a58982a  and  a58979a );
 a58984a <=( a58983a  and  a58976a );
 a58988a <=( (not A168)  and  (not A169) );
 a58989a <=( (not A170)  and  a58988a );
 a58993a <=( A199  and  A166 );
 a58994a <=( (not A167)  and  a58993a );
 a58995a <=( a58994a  and  a58989a );
 a58999a <=( A266  and  (not A265) );
 a59000a <=( A200  and  a58999a );
 a59003a <=( (not A269)  and  A267 );
 a59006a <=( (not A302)  and  (not A300) );
 a59007a <=( a59006a  and  a59003a );
 a59008a <=( a59007a  and  a59000a );
 a59012a <=( (not A168)  and  (not A169) );
 a59013a <=( (not A170)  and  a59012a );
 a59017a <=( A199  and  A166 );
 a59018a <=( (not A167)  and  a59017a );
 a59019a <=( a59018a  and  a59013a );
 a59023a <=( A266  and  (not A265) );
 a59024a <=( A200  and  a59023a );
 a59027a <=( (not A269)  and  A267 );
 a59030a <=( A299  and  A298 );
 a59031a <=( a59030a  and  a59027a );
 a59032a <=( a59031a  and  a59024a );
 a59036a <=( (not A168)  and  (not A169) );
 a59037a <=( (not A170)  and  a59036a );
 a59041a <=( A199  and  A166 );
 a59042a <=( (not A167)  and  a59041a );
 a59043a <=( a59042a  and  a59037a );
 a59047a <=( A266  and  (not A265) );
 a59048a <=( A200  and  a59047a );
 a59051a <=( (not A269)  and  A267 );
 a59054a <=( (not A299)  and  (not A298) );
 a59055a <=( a59054a  and  a59051a );
 a59056a <=( a59055a  and  a59048a );
 a59060a <=( (not A168)  and  (not A169) );
 a59061a <=( (not A170)  and  a59060a );
 a59065a <=( A199  and  A166 );
 a59066a <=( (not A167)  and  a59065a );
 a59067a <=( a59066a  and  a59061a );
 a59071a <=( (not A266)  and  A265 );
 a59072a <=( A200  and  a59071a );
 a59075a <=( A268  and  A267 );
 a59078a <=( A301  and  (not A300) );
 a59079a <=( a59078a  and  a59075a );
 a59080a <=( a59079a  and  a59072a );
 a59084a <=( (not A168)  and  (not A169) );
 a59085a <=( (not A170)  and  a59084a );
 a59089a <=( A199  and  A166 );
 a59090a <=( (not A167)  and  a59089a );
 a59091a <=( a59090a  and  a59085a );
 a59095a <=( (not A266)  and  A265 );
 a59096a <=( A200  and  a59095a );
 a59099a <=( A268  and  A267 );
 a59102a <=( (not A302)  and  (not A300) );
 a59103a <=( a59102a  and  a59099a );
 a59104a <=( a59103a  and  a59096a );
 a59108a <=( (not A168)  and  (not A169) );
 a59109a <=( (not A170)  and  a59108a );
 a59113a <=( A199  and  A166 );
 a59114a <=( (not A167)  and  a59113a );
 a59115a <=( a59114a  and  a59109a );
 a59119a <=( (not A266)  and  A265 );
 a59120a <=( A200  and  a59119a );
 a59123a <=( A268  and  A267 );
 a59126a <=( A299  and  A298 );
 a59127a <=( a59126a  and  a59123a );
 a59128a <=( a59127a  and  a59120a );
 a59132a <=( (not A168)  and  (not A169) );
 a59133a <=( (not A170)  and  a59132a );
 a59137a <=( A199  and  A166 );
 a59138a <=( (not A167)  and  a59137a );
 a59139a <=( a59138a  and  a59133a );
 a59143a <=( (not A266)  and  A265 );
 a59144a <=( A200  and  a59143a );
 a59147a <=( A268  and  A267 );
 a59150a <=( (not A299)  and  (not A298) );
 a59151a <=( a59150a  and  a59147a );
 a59152a <=( a59151a  and  a59144a );
 a59156a <=( (not A168)  and  (not A169) );
 a59157a <=( (not A170)  and  a59156a );
 a59161a <=( A199  and  A166 );
 a59162a <=( (not A167)  and  a59161a );
 a59163a <=( a59162a  and  a59157a );
 a59167a <=( (not A266)  and  A265 );
 a59168a <=( A200  and  a59167a );
 a59171a <=( (not A269)  and  A267 );
 a59174a <=( A301  and  (not A300) );
 a59175a <=( a59174a  and  a59171a );
 a59176a <=( a59175a  and  a59168a );
 a59180a <=( (not A168)  and  (not A169) );
 a59181a <=( (not A170)  and  a59180a );
 a59185a <=( A199  and  A166 );
 a59186a <=( (not A167)  and  a59185a );
 a59187a <=( a59186a  and  a59181a );
 a59191a <=( (not A266)  and  A265 );
 a59192a <=( A200  and  a59191a );
 a59195a <=( (not A269)  and  A267 );
 a59198a <=( (not A302)  and  (not A300) );
 a59199a <=( a59198a  and  a59195a );
 a59200a <=( a59199a  and  a59192a );
 a59204a <=( (not A168)  and  (not A169) );
 a59205a <=( (not A170)  and  a59204a );
 a59209a <=( A199  and  A166 );
 a59210a <=( (not A167)  and  a59209a );
 a59211a <=( a59210a  and  a59205a );
 a59215a <=( (not A266)  and  A265 );
 a59216a <=( A200  and  a59215a );
 a59219a <=( (not A269)  and  A267 );
 a59222a <=( A299  and  A298 );
 a59223a <=( a59222a  and  a59219a );
 a59224a <=( a59223a  and  a59216a );
 a59228a <=( (not A168)  and  (not A169) );
 a59229a <=( (not A170)  and  a59228a );
 a59233a <=( A199  and  A166 );
 a59234a <=( (not A167)  and  a59233a );
 a59235a <=( a59234a  and  a59229a );
 a59239a <=( (not A266)  and  A265 );
 a59240a <=( A200  and  a59239a );
 a59243a <=( (not A269)  and  A267 );
 a59246a <=( (not A299)  and  (not A298) );
 a59247a <=( a59246a  and  a59243a );
 a59248a <=( a59247a  and  a59240a );
 a59252a <=( (not A168)  and  (not A169) );
 a59253a <=( (not A170)  and  a59252a );
 a59257a <=( A199  and  A166 );
 a59258a <=( (not A167)  and  a59257a );
 a59259a <=( a59258a  and  a59253a );
 a59263a <=( (not A266)  and  (not A265) );
 a59264a <=( A200  and  a59263a );
 a59267a <=( (not A299)  and  A298 );
 a59270a <=( A301  and  A300 );
 a59271a <=( a59270a  and  a59267a );
 a59272a <=( a59271a  and  a59264a );
 a59276a <=( (not A168)  and  (not A169) );
 a59277a <=( (not A170)  and  a59276a );
 a59281a <=( A199  and  A166 );
 a59282a <=( (not A167)  and  a59281a );
 a59283a <=( a59282a  and  a59277a );
 a59287a <=( (not A266)  and  (not A265) );
 a59288a <=( A200  and  a59287a );
 a59291a <=( (not A299)  and  A298 );
 a59294a <=( (not A302)  and  A300 );
 a59295a <=( a59294a  and  a59291a );
 a59296a <=( a59295a  and  a59288a );
 a59300a <=( (not A168)  and  (not A169) );
 a59301a <=( (not A170)  and  a59300a );
 a59305a <=( A199  and  A166 );
 a59306a <=( (not A167)  and  a59305a );
 a59307a <=( a59306a  and  a59301a );
 a59311a <=( (not A266)  and  (not A265) );
 a59312a <=( A200  and  a59311a );
 a59315a <=( A299  and  (not A298) );
 a59318a <=( A301  and  A300 );
 a59319a <=( a59318a  and  a59315a );
 a59320a <=( a59319a  and  a59312a );
 a59324a <=( (not A168)  and  (not A169) );
 a59325a <=( (not A170)  and  a59324a );
 a59329a <=( A199  and  A166 );
 a59330a <=( (not A167)  and  a59329a );
 a59331a <=( a59330a  and  a59325a );
 a59335a <=( (not A266)  and  (not A265) );
 a59336a <=( A200  and  a59335a );
 a59339a <=( A299  and  (not A298) );
 a59342a <=( (not A302)  and  A300 );
 a59343a <=( a59342a  and  a59339a );
 a59344a <=( a59343a  and  a59336a );
 a59348a <=( (not A168)  and  (not A169) );
 a59349a <=( (not A170)  and  a59348a );
 a59353a <=( (not A199)  and  A166 );
 a59354a <=( (not A167)  and  a59353a );
 a59355a <=( a59354a  and  a59349a );
 a59359a <=( A268  and  (not A267) );
 a59360a <=( (not A200)  and  a59359a );
 a59363a <=( (not A299)  and  A298 );
 a59366a <=( A301  and  A300 );
 a59367a <=( a59366a  and  a59363a );
 a59368a <=( a59367a  and  a59360a );
 a59372a <=( (not A168)  and  (not A169) );
 a59373a <=( (not A170)  and  a59372a );
 a59377a <=( (not A199)  and  A166 );
 a59378a <=( (not A167)  and  a59377a );
 a59379a <=( a59378a  and  a59373a );
 a59383a <=( A268  and  (not A267) );
 a59384a <=( (not A200)  and  a59383a );
 a59387a <=( (not A299)  and  A298 );
 a59390a <=( (not A302)  and  A300 );
 a59391a <=( a59390a  and  a59387a );
 a59392a <=( a59391a  and  a59384a );
 a59396a <=( (not A168)  and  (not A169) );
 a59397a <=( (not A170)  and  a59396a );
 a59401a <=( (not A199)  and  A166 );
 a59402a <=( (not A167)  and  a59401a );
 a59403a <=( a59402a  and  a59397a );
 a59407a <=( A268  and  (not A267) );
 a59408a <=( (not A200)  and  a59407a );
 a59411a <=( A299  and  (not A298) );
 a59414a <=( A301  and  A300 );
 a59415a <=( a59414a  and  a59411a );
 a59416a <=( a59415a  and  a59408a );
 a59420a <=( (not A168)  and  (not A169) );
 a59421a <=( (not A170)  and  a59420a );
 a59425a <=( (not A199)  and  A166 );
 a59426a <=( (not A167)  and  a59425a );
 a59427a <=( a59426a  and  a59421a );
 a59431a <=( A268  and  (not A267) );
 a59432a <=( (not A200)  and  a59431a );
 a59435a <=( A299  and  (not A298) );
 a59438a <=( (not A302)  and  A300 );
 a59439a <=( a59438a  and  a59435a );
 a59440a <=( a59439a  and  a59432a );
 a59444a <=( (not A168)  and  (not A169) );
 a59445a <=( (not A170)  and  a59444a );
 a59449a <=( (not A199)  and  A166 );
 a59450a <=( (not A167)  and  a59449a );
 a59451a <=( a59450a  and  a59445a );
 a59455a <=( (not A269)  and  (not A267) );
 a59456a <=( (not A200)  and  a59455a );
 a59459a <=( (not A299)  and  A298 );
 a59462a <=( A301  and  A300 );
 a59463a <=( a59462a  and  a59459a );
 a59464a <=( a59463a  and  a59456a );
 a59468a <=( (not A168)  and  (not A169) );
 a59469a <=( (not A170)  and  a59468a );
 a59473a <=( (not A199)  and  A166 );
 a59474a <=( (not A167)  and  a59473a );
 a59475a <=( a59474a  and  a59469a );
 a59479a <=( (not A269)  and  (not A267) );
 a59480a <=( (not A200)  and  a59479a );
 a59483a <=( (not A299)  and  A298 );
 a59486a <=( (not A302)  and  A300 );
 a59487a <=( a59486a  and  a59483a );
 a59488a <=( a59487a  and  a59480a );
 a59492a <=( (not A168)  and  (not A169) );
 a59493a <=( (not A170)  and  a59492a );
 a59497a <=( (not A199)  and  A166 );
 a59498a <=( (not A167)  and  a59497a );
 a59499a <=( a59498a  and  a59493a );
 a59503a <=( (not A269)  and  (not A267) );
 a59504a <=( (not A200)  and  a59503a );
 a59507a <=( A299  and  (not A298) );
 a59510a <=( A301  and  A300 );
 a59511a <=( a59510a  and  a59507a );
 a59512a <=( a59511a  and  a59504a );
 a59516a <=( (not A168)  and  (not A169) );
 a59517a <=( (not A170)  and  a59516a );
 a59521a <=( (not A199)  and  A166 );
 a59522a <=( (not A167)  and  a59521a );
 a59523a <=( a59522a  and  a59517a );
 a59527a <=( (not A269)  and  (not A267) );
 a59528a <=( (not A200)  and  a59527a );
 a59531a <=( A299  and  (not A298) );
 a59534a <=( (not A302)  and  A300 );
 a59535a <=( a59534a  and  a59531a );
 a59536a <=( a59535a  and  a59528a );
 a59540a <=( (not A168)  and  (not A169) );
 a59541a <=( (not A170)  and  a59540a );
 a59545a <=( (not A199)  and  A166 );
 a59546a <=( (not A167)  and  a59545a );
 a59547a <=( a59546a  and  a59541a );
 a59551a <=( A266  and  A265 );
 a59552a <=( (not A200)  and  a59551a );
 a59555a <=( (not A299)  and  A298 );
 a59558a <=( A301  and  A300 );
 a59559a <=( a59558a  and  a59555a );
 a59560a <=( a59559a  and  a59552a );
 a59564a <=( (not A168)  and  (not A169) );
 a59565a <=( (not A170)  and  a59564a );
 a59569a <=( (not A199)  and  A166 );
 a59570a <=( (not A167)  and  a59569a );
 a59571a <=( a59570a  and  a59565a );
 a59575a <=( A266  and  A265 );
 a59576a <=( (not A200)  and  a59575a );
 a59579a <=( (not A299)  and  A298 );
 a59582a <=( (not A302)  and  A300 );
 a59583a <=( a59582a  and  a59579a );
 a59584a <=( a59583a  and  a59576a );
 a59588a <=( (not A168)  and  (not A169) );
 a59589a <=( (not A170)  and  a59588a );
 a59593a <=( (not A199)  and  A166 );
 a59594a <=( (not A167)  and  a59593a );
 a59595a <=( a59594a  and  a59589a );
 a59599a <=( A266  and  A265 );
 a59600a <=( (not A200)  and  a59599a );
 a59603a <=( A299  and  (not A298) );
 a59606a <=( A301  and  A300 );
 a59607a <=( a59606a  and  a59603a );
 a59608a <=( a59607a  and  a59600a );
 a59612a <=( (not A168)  and  (not A169) );
 a59613a <=( (not A170)  and  a59612a );
 a59617a <=( (not A199)  and  A166 );
 a59618a <=( (not A167)  and  a59617a );
 a59619a <=( a59618a  and  a59613a );
 a59623a <=( A266  and  A265 );
 a59624a <=( (not A200)  and  a59623a );
 a59627a <=( A299  and  (not A298) );
 a59630a <=( (not A302)  and  A300 );
 a59631a <=( a59630a  and  a59627a );
 a59632a <=( a59631a  and  a59624a );
 a59636a <=( (not A168)  and  (not A169) );
 a59637a <=( (not A170)  and  a59636a );
 a59641a <=( (not A199)  and  A166 );
 a59642a <=( (not A167)  and  a59641a );
 a59643a <=( a59642a  and  a59637a );
 a59647a <=( A266  and  (not A265) );
 a59648a <=( (not A200)  and  a59647a );
 a59651a <=( A268  and  A267 );
 a59654a <=( A301  and  (not A300) );
 a59655a <=( a59654a  and  a59651a );
 a59656a <=( a59655a  and  a59648a );
 a59660a <=( (not A168)  and  (not A169) );
 a59661a <=( (not A170)  and  a59660a );
 a59665a <=( (not A199)  and  A166 );
 a59666a <=( (not A167)  and  a59665a );
 a59667a <=( a59666a  and  a59661a );
 a59671a <=( A266  and  (not A265) );
 a59672a <=( (not A200)  and  a59671a );
 a59675a <=( A268  and  A267 );
 a59678a <=( (not A302)  and  (not A300) );
 a59679a <=( a59678a  and  a59675a );
 a59680a <=( a59679a  and  a59672a );
 a59684a <=( (not A168)  and  (not A169) );
 a59685a <=( (not A170)  and  a59684a );
 a59689a <=( (not A199)  and  A166 );
 a59690a <=( (not A167)  and  a59689a );
 a59691a <=( a59690a  and  a59685a );
 a59695a <=( A266  and  (not A265) );
 a59696a <=( (not A200)  and  a59695a );
 a59699a <=( A268  and  A267 );
 a59702a <=( A299  and  A298 );
 a59703a <=( a59702a  and  a59699a );
 a59704a <=( a59703a  and  a59696a );
 a59708a <=( (not A168)  and  (not A169) );
 a59709a <=( (not A170)  and  a59708a );
 a59713a <=( (not A199)  and  A166 );
 a59714a <=( (not A167)  and  a59713a );
 a59715a <=( a59714a  and  a59709a );
 a59719a <=( A266  and  (not A265) );
 a59720a <=( (not A200)  and  a59719a );
 a59723a <=( A268  and  A267 );
 a59726a <=( (not A299)  and  (not A298) );
 a59727a <=( a59726a  and  a59723a );
 a59728a <=( a59727a  and  a59720a );
 a59732a <=( (not A168)  and  (not A169) );
 a59733a <=( (not A170)  and  a59732a );
 a59737a <=( (not A199)  and  A166 );
 a59738a <=( (not A167)  and  a59737a );
 a59739a <=( a59738a  and  a59733a );
 a59743a <=( A266  and  (not A265) );
 a59744a <=( (not A200)  and  a59743a );
 a59747a <=( (not A269)  and  A267 );
 a59750a <=( A301  and  (not A300) );
 a59751a <=( a59750a  and  a59747a );
 a59752a <=( a59751a  and  a59744a );
 a59756a <=( (not A168)  and  (not A169) );
 a59757a <=( (not A170)  and  a59756a );
 a59761a <=( (not A199)  and  A166 );
 a59762a <=( (not A167)  and  a59761a );
 a59763a <=( a59762a  and  a59757a );
 a59767a <=( A266  and  (not A265) );
 a59768a <=( (not A200)  and  a59767a );
 a59771a <=( (not A269)  and  A267 );
 a59774a <=( (not A302)  and  (not A300) );
 a59775a <=( a59774a  and  a59771a );
 a59776a <=( a59775a  and  a59768a );
 a59780a <=( (not A168)  and  (not A169) );
 a59781a <=( (not A170)  and  a59780a );
 a59785a <=( (not A199)  and  A166 );
 a59786a <=( (not A167)  and  a59785a );
 a59787a <=( a59786a  and  a59781a );
 a59791a <=( A266  and  (not A265) );
 a59792a <=( (not A200)  and  a59791a );
 a59795a <=( (not A269)  and  A267 );
 a59798a <=( A299  and  A298 );
 a59799a <=( a59798a  and  a59795a );
 a59800a <=( a59799a  and  a59792a );
 a59804a <=( (not A168)  and  (not A169) );
 a59805a <=( (not A170)  and  a59804a );
 a59809a <=( (not A199)  and  A166 );
 a59810a <=( (not A167)  and  a59809a );
 a59811a <=( a59810a  and  a59805a );
 a59815a <=( A266  and  (not A265) );
 a59816a <=( (not A200)  and  a59815a );
 a59819a <=( (not A269)  and  A267 );
 a59822a <=( (not A299)  and  (not A298) );
 a59823a <=( a59822a  and  a59819a );
 a59824a <=( a59823a  and  a59816a );
 a59828a <=( (not A168)  and  (not A169) );
 a59829a <=( (not A170)  and  a59828a );
 a59833a <=( (not A199)  and  A166 );
 a59834a <=( (not A167)  and  a59833a );
 a59835a <=( a59834a  and  a59829a );
 a59839a <=( (not A266)  and  A265 );
 a59840a <=( (not A200)  and  a59839a );
 a59843a <=( A268  and  A267 );
 a59846a <=( A301  and  (not A300) );
 a59847a <=( a59846a  and  a59843a );
 a59848a <=( a59847a  and  a59840a );
 a59852a <=( (not A168)  and  (not A169) );
 a59853a <=( (not A170)  and  a59852a );
 a59857a <=( (not A199)  and  A166 );
 a59858a <=( (not A167)  and  a59857a );
 a59859a <=( a59858a  and  a59853a );
 a59863a <=( (not A266)  and  A265 );
 a59864a <=( (not A200)  and  a59863a );
 a59867a <=( A268  and  A267 );
 a59870a <=( (not A302)  and  (not A300) );
 a59871a <=( a59870a  and  a59867a );
 a59872a <=( a59871a  and  a59864a );
 a59876a <=( (not A168)  and  (not A169) );
 a59877a <=( (not A170)  and  a59876a );
 a59881a <=( (not A199)  and  A166 );
 a59882a <=( (not A167)  and  a59881a );
 a59883a <=( a59882a  and  a59877a );
 a59887a <=( (not A266)  and  A265 );
 a59888a <=( (not A200)  and  a59887a );
 a59891a <=( A268  and  A267 );
 a59894a <=( A299  and  A298 );
 a59895a <=( a59894a  and  a59891a );
 a59896a <=( a59895a  and  a59888a );
 a59900a <=( (not A168)  and  (not A169) );
 a59901a <=( (not A170)  and  a59900a );
 a59905a <=( (not A199)  and  A166 );
 a59906a <=( (not A167)  and  a59905a );
 a59907a <=( a59906a  and  a59901a );
 a59911a <=( (not A266)  and  A265 );
 a59912a <=( (not A200)  and  a59911a );
 a59915a <=( A268  and  A267 );
 a59918a <=( (not A299)  and  (not A298) );
 a59919a <=( a59918a  and  a59915a );
 a59920a <=( a59919a  and  a59912a );
 a59924a <=( (not A168)  and  (not A169) );
 a59925a <=( (not A170)  and  a59924a );
 a59929a <=( (not A199)  and  A166 );
 a59930a <=( (not A167)  and  a59929a );
 a59931a <=( a59930a  and  a59925a );
 a59935a <=( (not A266)  and  A265 );
 a59936a <=( (not A200)  and  a59935a );
 a59939a <=( (not A269)  and  A267 );
 a59942a <=( A301  and  (not A300) );
 a59943a <=( a59942a  and  a59939a );
 a59944a <=( a59943a  and  a59936a );
 a59948a <=( (not A168)  and  (not A169) );
 a59949a <=( (not A170)  and  a59948a );
 a59953a <=( (not A199)  and  A166 );
 a59954a <=( (not A167)  and  a59953a );
 a59955a <=( a59954a  and  a59949a );
 a59959a <=( (not A266)  and  A265 );
 a59960a <=( (not A200)  and  a59959a );
 a59963a <=( (not A269)  and  A267 );
 a59966a <=( (not A302)  and  (not A300) );
 a59967a <=( a59966a  and  a59963a );
 a59968a <=( a59967a  and  a59960a );
 a59972a <=( (not A168)  and  (not A169) );
 a59973a <=( (not A170)  and  a59972a );
 a59977a <=( (not A199)  and  A166 );
 a59978a <=( (not A167)  and  a59977a );
 a59979a <=( a59978a  and  a59973a );
 a59983a <=( (not A266)  and  A265 );
 a59984a <=( (not A200)  and  a59983a );
 a59987a <=( (not A269)  and  A267 );
 a59990a <=( A299  and  A298 );
 a59991a <=( a59990a  and  a59987a );
 a59992a <=( a59991a  and  a59984a );
 a59996a <=( (not A168)  and  (not A169) );
 a59997a <=( (not A170)  and  a59996a );
 a60001a <=( (not A199)  and  A166 );
 a60002a <=( (not A167)  and  a60001a );
 a60003a <=( a60002a  and  a59997a );
 a60007a <=( (not A266)  and  A265 );
 a60008a <=( (not A200)  and  a60007a );
 a60011a <=( (not A269)  and  A267 );
 a60014a <=( (not A299)  and  (not A298) );
 a60015a <=( a60014a  and  a60011a );
 a60016a <=( a60015a  and  a60008a );
 a60020a <=( (not A168)  and  (not A169) );
 a60021a <=( (not A170)  and  a60020a );
 a60025a <=( (not A199)  and  A166 );
 a60026a <=( (not A167)  and  a60025a );
 a60027a <=( a60026a  and  a60021a );
 a60031a <=( (not A266)  and  (not A265) );
 a60032a <=( (not A200)  and  a60031a );
 a60035a <=( (not A299)  and  A298 );
 a60038a <=( A301  and  A300 );
 a60039a <=( a60038a  and  a60035a );
 a60040a <=( a60039a  and  a60032a );
 a60044a <=( (not A168)  and  (not A169) );
 a60045a <=( (not A170)  and  a60044a );
 a60049a <=( (not A199)  and  A166 );
 a60050a <=( (not A167)  and  a60049a );
 a60051a <=( a60050a  and  a60045a );
 a60055a <=( (not A266)  and  (not A265) );
 a60056a <=( (not A200)  and  a60055a );
 a60059a <=( (not A299)  and  A298 );
 a60062a <=( (not A302)  and  A300 );
 a60063a <=( a60062a  and  a60059a );
 a60064a <=( a60063a  and  a60056a );
 a60068a <=( (not A168)  and  (not A169) );
 a60069a <=( (not A170)  and  a60068a );
 a60073a <=( (not A199)  and  A166 );
 a60074a <=( (not A167)  and  a60073a );
 a60075a <=( a60074a  and  a60069a );
 a60079a <=( (not A266)  and  (not A265) );
 a60080a <=( (not A200)  and  a60079a );
 a60083a <=( A299  and  (not A298) );
 a60086a <=( A301  and  A300 );
 a60087a <=( a60086a  and  a60083a );
 a60088a <=( a60087a  and  a60080a );
 a60092a <=( (not A168)  and  (not A169) );
 a60093a <=( (not A170)  and  a60092a );
 a60097a <=( (not A199)  and  A166 );
 a60098a <=( (not A167)  and  a60097a );
 a60099a <=( a60098a  and  a60093a );
 a60103a <=( (not A266)  and  (not A265) );
 a60104a <=( (not A200)  and  a60103a );
 a60107a <=( A299  and  (not A298) );
 a60110a <=( (not A302)  and  A300 );
 a60111a <=( a60110a  and  a60107a );
 a60112a <=( a60111a  and  a60104a );
 a60116a <=( (not A199)  and  A166 );
 a60117a <=( A167  and  a60116a );
 a60120a <=( A201  and  A200 );
 a60123a <=( (not A265)  and  A202 );
 a60124a <=( a60123a  and  a60120a );
 a60125a <=( a60124a  and  a60117a );
 a60129a <=( A268  and  A267 );
 a60130a <=( A266  and  a60129a );
 a60133a <=( (not A299)  and  A298 );
 a60136a <=( A301  and  A300 );
 a60137a <=( a60136a  and  a60133a );
 a60138a <=( a60137a  and  a60130a );
 a60142a <=( (not A199)  and  A166 );
 a60143a <=( A167  and  a60142a );
 a60146a <=( A201  and  A200 );
 a60149a <=( (not A265)  and  A202 );
 a60150a <=( a60149a  and  a60146a );
 a60151a <=( a60150a  and  a60143a );
 a60155a <=( A268  and  A267 );
 a60156a <=( A266  and  a60155a );
 a60159a <=( (not A299)  and  A298 );
 a60162a <=( (not A302)  and  A300 );
 a60163a <=( a60162a  and  a60159a );
 a60164a <=( a60163a  and  a60156a );
 a60168a <=( (not A199)  and  A166 );
 a60169a <=( A167  and  a60168a );
 a60172a <=( A201  and  A200 );
 a60175a <=( (not A265)  and  A202 );
 a60176a <=( a60175a  and  a60172a );
 a60177a <=( a60176a  and  a60169a );
 a60181a <=( A268  and  A267 );
 a60182a <=( A266  and  a60181a );
 a60185a <=( A299  and  (not A298) );
 a60188a <=( A301  and  A300 );
 a60189a <=( a60188a  and  a60185a );
 a60190a <=( a60189a  and  a60182a );
 a60194a <=( (not A199)  and  A166 );
 a60195a <=( A167  and  a60194a );
 a60198a <=( A201  and  A200 );
 a60201a <=( (not A265)  and  A202 );
 a60202a <=( a60201a  and  a60198a );
 a60203a <=( a60202a  and  a60195a );
 a60207a <=( A268  and  A267 );
 a60208a <=( A266  and  a60207a );
 a60211a <=( A299  and  (not A298) );
 a60214a <=( (not A302)  and  A300 );
 a60215a <=( a60214a  and  a60211a );
 a60216a <=( a60215a  and  a60208a );
 a60220a <=( (not A199)  and  A166 );
 a60221a <=( A167  and  a60220a );
 a60224a <=( A201  and  A200 );
 a60227a <=( (not A265)  and  A202 );
 a60228a <=( a60227a  and  a60224a );
 a60229a <=( a60228a  and  a60221a );
 a60233a <=( (not A269)  and  A267 );
 a60234a <=( A266  and  a60233a );
 a60237a <=( (not A299)  and  A298 );
 a60240a <=( A301  and  A300 );
 a60241a <=( a60240a  and  a60237a );
 a60242a <=( a60241a  and  a60234a );
 a60246a <=( (not A199)  and  A166 );
 a60247a <=( A167  and  a60246a );
 a60250a <=( A201  and  A200 );
 a60253a <=( (not A265)  and  A202 );
 a60254a <=( a60253a  and  a60250a );
 a60255a <=( a60254a  and  a60247a );
 a60259a <=( (not A269)  and  A267 );
 a60260a <=( A266  and  a60259a );
 a60263a <=( (not A299)  and  A298 );
 a60266a <=( (not A302)  and  A300 );
 a60267a <=( a60266a  and  a60263a );
 a60268a <=( a60267a  and  a60260a );
 a60272a <=( (not A199)  and  A166 );
 a60273a <=( A167  and  a60272a );
 a60276a <=( A201  and  A200 );
 a60279a <=( (not A265)  and  A202 );
 a60280a <=( a60279a  and  a60276a );
 a60281a <=( a60280a  and  a60273a );
 a60285a <=( (not A269)  and  A267 );
 a60286a <=( A266  and  a60285a );
 a60289a <=( A299  and  (not A298) );
 a60292a <=( A301  and  A300 );
 a60293a <=( a60292a  and  a60289a );
 a60294a <=( a60293a  and  a60286a );
 a60298a <=( (not A199)  and  A166 );
 a60299a <=( A167  and  a60298a );
 a60302a <=( A201  and  A200 );
 a60305a <=( (not A265)  and  A202 );
 a60306a <=( a60305a  and  a60302a );
 a60307a <=( a60306a  and  a60299a );
 a60311a <=( (not A269)  and  A267 );
 a60312a <=( A266  and  a60311a );
 a60315a <=( A299  and  (not A298) );
 a60318a <=( (not A302)  and  A300 );
 a60319a <=( a60318a  and  a60315a );
 a60320a <=( a60319a  and  a60312a );
 a60324a <=( (not A199)  and  A166 );
 a60325a <=( A167  and  a60324a );
 a60328a <=( A201  and  A200 );
 a60331a <=( A265  and  A202 );
 a60332a <=( a60331a  and  a60328a );
 a60333a <=( a60332a  and  a60325a );
 a60337a <=( A268  and  A267 );
 a60338a <=( (not A266)  and  a60337a );
 a60341a <=( (not A299)  and  A298 );
 a60344a <=( A301  and  A300 );
 a60345a <=( a60344a  and  a60341a );
 a60346a <=( a60345a  and  a60338a );
 a60350a <=( (not A199)  and  A166 );
 a60351a <=( A167  and  a60350a );
 a60354a <=( A201  and  A200 );
 a60357a <=( A265  and  A202 );
 a60358a <=( a60357a  and  a60354a );
 a60359a <=( a60358a  and  a60351a );
 a60363a <=( A268  and  A267 );
 a60364a <=( (not A266)  and  a60363a );
 a60367a <=( (not A299)  and  A298 );
 a60370a <=( (not A302)  and  A300 );
 a60371a <=( a60370a  and  a60367a );
 a60372a <=( a60371a  and  a60364a );
 a60376a <=( (not A199)  and  A166 );
 a60377a <=( A167  and  a60376a );
 a60380a <=( A201  and  A200 );
 a60383a <=( A265  and  A202 );
 a60384a <=( a60383a  and  a60380a );
 a60385a <=( a60384a  and  a60377a );
 a60389a <=( A268  and  A267 );
 a60390a <=( (not A266)  and  a60389a );
 a60393a <=( A299  and  (not A298) );
 a60396a <=( A301  and  A300 );
 a60397a <=( a60396a  and  a60393a );
 a60398a <=( a60397a  and  a60390a );
 a60402a <=( (not A199)  and  A166 );
 a60403a <=( A167  and  a60402a );
 a60406a <=( A201  and  A200 );
 a60409a <=( A265  and  A202 );
 a60410a <=( a60409a  and  a60406a );
 a60411a <=( a60410a  and  a60403a );
 a60415a <=( A268  and  A267 );
 a60416a <=( (not A266)  and  a60415a );
 a60419a <=( A299  and  (not A298) );
 a60422a <=( (not A302)  and  A300 );
 a60423a <=( a60422a  and  a60419a );
 a60424a <=( a60423a  and  a60416a );
 a60428a <=( (not A199)  and  A166 );
 a60429a <=( A167  and  a60428a );
 a60432a <=( A201  and  A200 );
 a60435a <=( A265  and  A202 );
 a60436a <=( a60435a  and  a60432a );
 a60437a <=( a60436a  and  a60429a );
 a60441a <=( (not A269)  and  A267 );
 a60442a <=( (not A266)  and  a60441a );
 a60445a <=( (not A299)  and  A298 );
 a60448a <=( A301  and  A300 );
 a60449a <=( a60448a  and  a60445a );
 a60450a <=( a60449a  and  a60442a );
 a60454a <=( (not A199)  and  A166 );
 a60455a <=( A167  and  a60454a );
 a60458a <=( A201  and  A200 );
 a60461a <=( A265  and  A202 );
 a60462a <=( a60461a  and  a60458a );
 a60463a <=( a60462a  and  a60455a );
 a60467a <=( (not A269)  and  A267 );
 a60468a <=( (not A266)  and  a60467a );
 a60471a <=( (not A299)  and  A298 );
 a60474a <=( (not A302)  and  A300 );
 a60475a <=( a60474a  and  a60471a );
 a60476a <=( a60475a  and  a60468a );
 a60480a <=( (not A199)  and  A166 );
 a60481a <=( A167  and  a60480a );
 a60484a <=( A201  and  A200 );
 a60487a <=( A265  and  A202 );
 a60488a <=( a60487a  and  a60484a );
 a60489a <=( a60488a  and  a60481a );
 a60493a <=( (not A269)  and  A267 );
 a60494a <=( (not A266)  and  a60493a );
 a60497a <=( A299  and  (not A298) );
 a60500a <=( A301  and  A300 );
 a60501a <=( a60500a  and  a60497a );
 a60502a <=( a60501a  and  a60494a );
 a60506a <=( (not A199)  and  A166 );
 a60507a <=( A167  and  a60506a );
 a60510a <=( A201  and  A200 );
 a60513a <=( A265  and  A202 );
 a60514a <=( a60513a  and  a60510a );
 a60515a <=( a60514a  and  a60507a );
 a60519a <=( (not A269)  and  A267 );
 a60520a <=( (not A266)  and  a60519a );
 a60523a <=( A299  and  (not A298) );
 a60526a <=( (not A302)  and  A300 );
 a60527a <=( a60526a  and  a60523a );
 a60528a <=( a60527a  and  a60520a );
 a60532a <=( (not A199)  and  A166 );
 a60533a <=( A167  and  a60532a );
 a60536a <=( A201  and  A200 );
 a60539a <=( (not A265)  and  (not A203) );
 a60540a <=( a60539a  and  a60536a );
 a60541a <=( a60540a  and  a60533a );
 a60545a <=( A268  and  A267 );
 a60546a <=( A266  and  a60545a );
 a60549a <=( (not A299)  and  A298 );
 a60552a <=( A301  and  A300 );
 a60553a <=( a60552a  and  a60549a );
 a60554a <=( a60553a  and  a60546a );
 a60558a <=( (not A199)  and  A166 );
 a60559a <=( A167  and  a60558a );
 a60562a <=( A201  and  A200 );
 a60565a <=( (not A265)  and  (not A203) );
 a60566a <=( a60565a  and  a60562a );
 a60567a <=( a60566a  and  a60559a );
 a60571a <=( A268  and  A267 );
 a60572a <=( A266  and  a60571a );
 a60575a <=( (not A299)  and  A298 );
 a60578a <=( (not A302)  and  A300 );
 a60579a <=( a60578a  and  a60575a );
 a60580a <=( a60579a  and  a60572a );
 a60584a <=( (not A199)  and  A166 );
 a60585a <=( A167  and  a60584a );
 a60588a <=( A201  and  A200 );
 a60591a <=( (not A265)  and  (not A203) );
 a60592a <=( a60591a  and  a60588a );
 a60593a <=( a60592a  and  a60585a );
 a60597a <=( A268  and  A267 );
 a60598a <=( A266  and  a60597a );
 a60601a <=( A299  and  (not A298) );
 a60604a <=( A301  and  A300 );
 a60605a <=( a60604a  and  a60601a );
 a60606a <=( a60605a  and  a60598a );
 a60610a <=( (not A199)  and  A166 );
 a60611a <=( A167  and  a60610a );
 a60614a <=( A201  and  A200 );
 a60617a <=( (not A265)  and  (not A203) );
 a60618a <=( a60617a  and  a60614a );
 a60619a <=( a60618a  and  a60611a );
 a60623a <=( A268  and  A267 );
 a60624a <=( A266  and  a60623a );
 a60627a <=( A299  and  (not A298) );
 a60630a <=( (not A302)  and  A300 );
 a60631a <=( a60630a  and  a60627a );
 a60632a <=( a60631a  and  a60624a );
 a60636a <=( (not A199)  and  A166 );
 a60637a <=( A167  and  a60636a );
 a60640a <=( A201  and  A200 );
 a60643a <=( (not A265)  and  (not A203) );
 a60644a <=( a60643a  and  a60640a );
 a60645a <=( a60644a  and  a60637a );
 a60649a <=( (not A269)  and  A267 );
 a60650a <=( A266  and  a60649a );
 a60653a <=( (not A299)  and  A298 );
 a60656a <=( A301  and  A300 );
 a60657a <=( a60656a  and  a60653a );
 a60658a <=( a60657a  and  a60650a );
 a60662a <=( (not A199)  and  A166 );
 a60663a <=( A167  and  a60662a );
 a60666a <=( A201  and  A200 );
 a60669a <=( (not A265)  and  (not A203) );
 a60670a <=( a60669a  and  a60666a );
 a60671a <=( a60670a  and  a60663a );
 a60675a <=( (not A269)  and  A267 );
 a60676a <=( A266  and  a60675a );
 a60679a <=( (not A299)  and  A298 );
 a60682a <=( (not A302)  and  A300 );
 a60683a <=( a60682a  and  a60679a );
 a60684a <=( a60683a  and  a60676a );
 a60688a <=( (not A199)  and  A166 );
 a60689a <=( A167  and  a60688a );
 a60692a <=( A201  and  A200 );
 a60695a <=( (not A265)  and  (not A203) );
 a60696a <=( a60695a  and  a60692a );
 a60697a <=( a60696a  and  a60689a );
 a60701a <=( (not A269)  and  A267 );
 a60702a <=( A266  and  a60701a );
 a60705a <=( A299  and  (not A298) );
 a60708a <=( A301  and  A300 );
 a60709a <=( a60708a  and  a60705a );
 a60710a <=( a60709a  and  a60702a );
 a60714a <=( (not A199)  and  A166 );
 a60715a <=( A167  and  a60714a );
 a60718a <=( A201  and  A200 );
 a60721a <=( (not A265)  and  (not A203) );
 a60722a <=( a60721a  and  a60718a );
 a60723a <=( a60722a  and  a60715a );
 a60727a <=( (not A269)  and  A267 );
 a60728a <=( A266  and  a60727a );
 a60731a <=( A299  and  (not A298) );
 a60734a <=( (not A302)  and  A300 );
 a60735a <=( a60734a  and  a60731a );
 a60736a <=( a60735a  and  a60728a );
 a60740a <=( (not A199)  and  A166 );
 a60741a <=( A167  and  a60740a );
 a60744a <=( A201  and  A200 );
 a60747a <=( A265  and  (not A203) );
 a60748a <=( a60747a  and  a60744a );
 a60749a <=( a60748a  and  a60741a );
 a60753a <=( A268  and  A267 );
 a60754a <=( (not A266)  and  a60753a );
 a60757a <=( (not A299)  and  A298 );
 a60760a <=( A301  and  A300 );
 a60761a <=( a60760a  and  a60757a );
 a60762a <=( a60761a  and  a60754a );
 a60766a <=( (not A199)  and  A166 );
 a60767a <=( A167  and  a60766a );
 a60770a <=( A201  and  A200 );
 a60773a <=( A265  and  (not A203) );
 a60774a <=( a60773a  and  a60770a );
 a60775a <=( a60774a  and  a60767a );
 a60779a <=( A268  and  A267 );
 a60780a <=( (not A266)  and  a60779a );
 a60783a <=( (not A299)  and  A298 );
 a60786a <=( (not A302)  and  A300 );
 a60787a <=( a60786a  and  a60783a );
 a60788a <=( a60787a  and  a60780a );
 a60792a <=( (not A199)  and  A166 );
 a60793a <=( A167  and  a60792a );
 a60796a <=( A201  and  A200 );
 a60799a <=( A265  and  (not A203) );
 a60800a <=( a60799a  and  a60796a );
 a60801a <=( a60800a  and  a60793a );
 a60805a <=( A268  and  A267 );
 a60806a <=( (not A266)  and  a60805a );
 a60809a <=( A299  and  (not A298) );
 a60812a <=( A301  and  A300 );
 a60813a <=( a60812a  and  a60809a );
 a60814a <=( a60813a  and  a60806a );
 a60818a <=( (not A199)  and  A166 );
 a60819a <=( A167  and  a60818a );
 a60822a <=( A201  and  A200 );
 a60825a <=( A265  and  (not A203) );
 a60826a <=( a60825a  and  a60822a );
 a60827a <=( a60826a  and  a60819a );
 a60831a <=( A268  and  A267 );
 a60832a <=( (not A266)  and  a60831a );
 a60835a <=( A299  and  (not A298) );
 a60838a <=( (not A302)  and  A300 );
 a60839a <=( a60838a  and  a60835a );
 a60840a <=( a60839a  and  a60832a );
 a60844a <=( (not A199)  and  A166 );
 a60845a <=( A167  and  a60844a );
 a60848a <=( A201  and  A200 );
 a60851a <=( A265  and  (not A203) );
 a60852a <=( a60851a  and  a60848a );
 a60853a <=( a60852a  and  a60845a );
 a60857a <=( (not A269)  and  A267 );
 a60858a <=( (not A266)  and  a60857a );
 a60861a <=( (not A299)  and  A298 );
 a60864a <=( A301  and  A300 );
 a60865a <=( a60864a  and  a60861a );
 a60866a <=( a60865a  and  a60858a );
 a60870a <=( (not A199)  and  A166 );
 a60871a <=( A167  and  a60870a );
 a60874a <=( A201  and  A200 );
 a60877a <=( A265  and  (not A203) );
 a60878a <=( a60877a  and  a60874a );
 a60879a <=( a60878a  and  a60871a );
 a60883a <=( (not A269)  and  A267 );
 a60884a <=( (not A266)  and  a60883a );
 a60887a <=( (not A299)  and  A298 );
 a60890a <=( (not A302)  and  A300 );
 a60891a <=( a60890a  and  a60887a );
 a60892a <=( a60891a  and  a60884a );
 a60896a <=( (not A199)  and  A166 );
 a60897a <=( A167  and  a60896a );
 a60900a <=( A201  and  A200 );
 a60903a <=( A265  and  (not A203) );
 a60904a <=( a60903a  and  a60900a );
 a60905a <=( a60904a  and  a60897a );
 a60909a <=( (not A269)  and  A267 );
 a60910a <=( (not A266)  and  a60909a );
 a60913a <=( A299  and  (not A298) );
 a60916a <=( A301  and  A300 );
 a60917a <=( a60916a  and  a60913a );
 a60918a <=( a60917a  and  a60910a );
 a60922a <=( (not A199)  and  A166 );
 a60923a <=( A167  and  a60922a );
 a60926a <=( A201  and  A200 );
 a60929a <=( A265  and  (not A203) );
 a60930a <=( a60929a  and  a60926a );
 a60931a <=( a60930a  and  a60923a );
 a60935a <=( (not A269)  and  A267 );
 a60936a <=( (not A266)  and  a60935a );
 a60939a <=( A299  and  (not A298) );
 a60942a <=( (not A302)  and  A300 );
 a60943a <=( a60942a  and  a60939a );
 a60944a <=( a60943a  and  a60936a );
 a60948a <=( A199  and  A166 );
 a60949a <=( A167  and  a60948a );
 a60952a <=( A201  and  (not A200) );
 a60955a <=( (not A265)  and  A202 );
 a60956a <=( a60955a  and  a60952a );
 a60957a <=( a60956a  and  a60949a );
 a60961a <=( A268  and  A267 );
 a60962a <=( A266  and  a60961a );
 a60965a <=( (not A299)  and  A298 );
 a60968a <=( A301  and  A300 );
 a60969a <=( a60968a  and  a60965a );
 a60970a <=( a60969a  and  a60962a );
 a60974a <=( A199  and  A166 );
 a60975a <=( A167  and  a60974a );
 a60978a <=( A201  and  (not A200) );
 a60981a <=( (not A265)  and  A202 );
 a60982a <=( a60981a  and  a60978a );
 a60983a <=( a60982a  and  a60975a );
 a60987a <=( A268  and  A267 );
 a60988a <=( A266  and  a60987a );
 a60991a <=( (not A299)  and  A298 );
 a60994a <=( (not A302)  and  A300 );
 a60995a <=( a60994a  and  a60991a );
 a60996a <=( a60995a  and  a60988a );
 a61000a <=( A199  and  A166 );
 a61001a <=( A167  and  a61000a );
 a61004a <=( A201  and  (not A200) );
 a61007a <=( (not A265)  and  A202 );
 a61008a <=( a61007a  and  a61004a );
 a61009a <=( a61008a  and  a61001a );
 a61013a <=( A268  and  A267 );
 a61014a <=( A266  and  a61013a );
 a61017a <=( A299  and  (not A298) );
 a61020a <=( A301  and  A300 );
 a61021a <=( a61020a  and  a61017a );
 a61022a <=( a61021a  and  a61014a );
 a61026a <=( A199  and  A166 );
 a61027a <=( A167  and  a61026a );
 a61030a <=( A201  and  (not A200) );
 a61033a <=( (not A265)  and  A202 );
 a61034a <=( a61033a  and  a61030a );
 a61035a <=( a61034a  and  a61027a );
 a61039a <=( A268  and  A267 );
 a61040a <=( A266  and  a61039a );
 a61043a <=( A299  and  (not A298) );
 a61046a <=( (not A302)  and  A300 );
 a61047a <=( a61046a  and  a61043a );
 a61048a <=( a61047a  and  a61040a );
 a61052a <=( A199  and  A166 );
 a61053a <=( A167  and  a61052a );
 a61056a <=( A201  and  (not A200) );
 a61059a <=( (not A265)  and  A202 );
 a61060a <=( a61059a  and  a61056a );
 a61061a <=( a61060a  and  a61053a );
 a61065a <=( (not A269)  and  A267 );
 a61066a <=( A266  and  a61065a );
 a61069a <=( (not A299)  and  A298 );
 a61072a <=( A301  and  A300 );
 a61073a <=( a61072a  and  a61069a );
 a61074a <=( a61073a  and  a61066a );
 a61078a <=( A199  and  A166 );
 a61079a <=( A167  and  a61078a );
 a61082a <=( A201  and  (not A200) );
 a61085a <=( (not A265)  and  A202 );
 a61086a <=( a61085a  and  a61082a );
 a61087a <=( a61086a  and  a61079a );
 a61091a <=( (not A269)  and  A267 );
 a61092a <=( A266  and  a61091a );
 a61095a <=( (not A299)  and  A298 );
 a61098a <=( (not A302)  and  A300 );
 a61099a <=( a61098a  and  a61095a );
 a61100a <=( a61099a  and  a61092a );
 a61104a <=( A199  and  A166 );
 a61105a <=( A167  and  a61104a );
 a61108a <=( A201  and  (not A200) );
 a61111a <=( (not A265)  and  A202 );
 a61112a <=( a61111a  and  a61108a );
 a61113a <=( a61112a  and  a61105a );
 a61117a <=( (not A269)  and  A267 );
 a61118a <=( A266  and  a61117a );
 a61121a <=( A299  and  (not A298) );
 a61124a <=( A301  and  A300 );
 a61125a <=( a61124a  and  a61121a );
 a61126a <=( a61125a  and  a61118a );
 a61130a <=( A199  and  A166 );
 a61131a <=( A167  and  a61130a );
 a61134a <=( A201  and  (not A200) );
 a61137a <=( (not A265)  and  A202 );
 a61138a <=( a61137a  and  a61134a );
 a61139a <=( a61138a  and  a61131a );
 a61143a <=( (not A269)  and  A267 );
 a61144a <=( A266  and  a61143a );
 a61147a <=( A299  and  (not A298) );
 a61150a <=( (not A302)  and  A300 );
 a61151a <=( a61150a  and  a61147a );
 a61152a <=( a61151a  and  a61144a );
 a61156a <=( A199  and  A166 );
 a61157a <=( A167  and  a61156a );
 a61160a <=( A201  and  (not A200) );
 a61163a <=( A265  and  A202 );
 a61164a <=( a61163a  and  a61160a );
 a61165a <=( a61164a  and  a61157a );
 a61169a <=( A268  and  A267 );
 a61170a <=( (not A266)  and  a61169a );
 a61173a <=( (not A299)  and  A298 );
 a61176a <=( A301  and  A300 );
 a61177a <=( a61176a  and  a61173a );
 a61178a <=( a61177a  and  a61170a );
 a61182a <=( A199  and  A166 );
 a61183a <=( A167  and  a61182a );
 a61186a <=( A201  and  (not A200) );
 a61189a <=( A265  and  A202 );
 a61190a <=( a61189a  and  a61186a );
 a61191a <=( a61190a  and  a61183a );
 a61195a <=( A268  and  A267 );
 a61196a <=( (not A266)  and  a61195a );
 a61199a <=( (not A299)  and  A298 );
 a61202a <=( (not A302)  and  A300 );
 a61203a <=( a61202a  and  a61199a );
 a61204a <=( a61203a  and  a61196a );
 a61208a <=( A199  and  A166 );
 a61209a <=( A167  and  a61208a );
 a61212a <=( A201  and  (not A200) );
 a61215a <=( A265  and  A202 );
 a61216a <=( a61215a  and  a61212a );
 a61217a <=( a61216a  and  a61209a );
 a61221a <=( A268  and  A267 );
 a61222a <=( (not A266)  and  a61221a );
 a61225a <=( A299  and  (not A298) );
 a61228a <=( A301  and  A300 );
 a61229a <=( a61228a  and  a61225a );
 a61230a <=( a61229a  and  a61222a );
 a61234a <=( A199  and  A166 );
 a61235a <=( A167  and  a61234a );
 a61238a <=( A201  and  (not A200) );
 a61241a <=( A265  and  A202 );
 a61242a <=( a61241a  and  a61238a );
 a61243a <=( a61242a  and  a61235a );
 a61247a <=( A268  and  A267 );
 a61248a <=( (not A266)  and  a61247a );
 a61251a <=( A299  and  (not A298) );
 a61254a <=( (not A302)  and  A300 );
 a61255a <=( a61254a  and  a61251a );
 a61256a <=( a61255a  and  a61248a );
 a61260a <=( A199  and  A166 );
 a61261a <=( A167  and  a61260a );
 a61264a <=( A201  and  (not A200) );
 a61267a <=( A265  and  A202 );
 a61268a <=( a61267a  and  a61264a );
 a61269a <=( a61268a  and  a61261a );
 a61273a <=( (not A269)  and  A267 );
 a61274a <=( (not A266)  and  a61273a );
 a61277a <=( (not A299)  and  A298 );
 a61280a <=( A301  and  A300 );
 a61281a <=( a61280a  and  a61277a );
 a61282a <=( a61281a  and  a61274a );
 a61286a <=( A199  and  A166 );
 a61287a <=( A167  and  a61286a );
 a61290a <=( A201  and  (not A200) );
 a61293a <=( A265  and  A202 );
 a61294a <=( a61293a  and  a61290a );
 a61295a <=( a61294a  and  a61287a );
 a61299a <=( (not A269)  and  A267 );
 a61300a <=( (not A266)  and  a61299a );
 a61303a <=( (not A299)  and  A298 );
 a61306a <=( (not A302)  and  A300 );
 a61307a <=( a61306a  and  a61303a );
 a61308a <=( a61307a  and  a61300a );
 a61312a <=( A199  and  A166 );
 a61313a <=( A167  and  a61312a );
 a61316a <=( A201  and  (not A200) );
 a61319a <=( A265  and  A202 );
 a61320a <=( a61319a  and  a61316a );
 a61321a <=( a61320a  and  a61313a );
 a61325a <=( (not A269)  and  A267 );
 a61326a <=( (not A266)  and  a61325a );
 a61329a <=( A299  and  (not A298) );
 a61332a <=( A301  and  A300 );
 a61333a <=( a61332a  and  a61329a );
 a61334a <=( a61333a  and  a61326a );
 a61338a <=( A199  and  A166 );
 a61339a <=( A167  and  a61338a );
 a61342a <=( A201  and  (not A200) );
 a61345a <=( A265  and  A202 );
 a61346a <=( a61345a  and  a61342a );
 a61347a <=( a61346a  and  a61339a );
 a61351a <=( (not A269)  and  A267 );
 a61352a <=( (not A266)  and  a61351a );
 a61355a <=( A299  and  (not A298) );
 a61358a <=( (not A302)  and  A300 );
 a61359a <=( a61358a  and  a61355a );
 a61360a <=( a61359a  and  a61352a );
 a61364a <=( A199  and  A166 );
 a61365a <=( A167  and  a61364a );
 a61368a <=( A201  and  (not A200) );
 a61371a <=( (not A265)  and  (not A203) );
 a61372a <=( a61371a  and  a61368a );
 a61373a <=( a61372a  and  a61365a );
 a61377a <=( A268  and  A267 );
 a61378a <=( A266  and  a61377a );
 a61381a <=( (not A299)  and  A298 );
 a61384a <=( A301  and  A300 );
 a61385a <=( a61384a  and  a61381a );
 a61386a <=( a61385a  and  a61378a );
 a61390a <=( A199  and  A166 );
 a61391a <=( A167  and  a61390a );
 a61394a <=( A201  and  (not A200) );
 a61397a <=( (not A265)  and  (not A203) );
 a61398a <=( a61397a  and  a61394a );
 a61399a <=( a61398a  and  a61391a );
 a61403a <=( A268  and  A267 );
 a61404a <=( A266  and  a61403a );
 a61407a <=( (not A299)  and  A298 );
 a61410a <=( (not A302)  and  A300 );
 a61411a <=( a61410a  and  a61407a );
 a61412a <=( a61411a  and  a61404a );
 a61416a <=( A199  and  A166 );
 a61417a <=( A167  and  a61416a );
 a61420a <=( A201  and  (not A200) );
 a61423a <=( (not A265)  and  (not A203) );
 a61424a <=( a61423a  and  a61420a );
 a61425a <=( a61424a  and  a61417a );
 a61429a <=( A268  and  A267 );
 a61430a <=( A266  and  a61429a );
 a61433a <=( A299  and  (not A298) );
 a61436a <=( A301  and  A300 );
 a61437a <=( a61436a  and  a61433a );
 a61438a <=( a61437a  and  a61430a );
 a61442a <=( A199  and  A166 );
 a61443a <=( A167  and  a61442a );
 a61446a <=( A201  and  (not A200) );
 a61449a <=( (not A265)  and  (not A203) );
 a61450a <=( a61449a  and  a61446a );
 a61451a <=( a61450a  and  a61443a );
 a61455a <=( A268  and  A267 );
 a61456a <=( A266  and  a61455a );
 a61459a <=( A299  and  (not A298) );
 a61462a <=( (not A302)  and  A300 );
 a61463a <=( a61462a  and  a61459a );
 a61464a <=( a61463a  and  a61456a );
 a61468a <=( A199  and  A166 );
 a61469a <=( A167  and  a61468a );
 a61472a <=( A201  and  (not A200) );
 a61475a <=( (not A265)  and  (not A203) );
 a61476a <=( a61475a  and  a61472a );
 a61477a <=( a61476a  and  a61469a );
 a61481a <=( (not A269)  and  A267 );
 a61482a <=( A266  and  a61481a );
 a61485a <=( (not A299)  and  A298 );
 a61488a <=( A301  and  A300 );
 a61489a <=( a61488a  and  a61485a );
 a61490a <=( a61489a  and  a61482a );
 a61494a <=( A199  and  A166 );
 a61495a <=( A167  and  a61494a );
 a61498a <=( A201  and  (not A200) );
 a61501a <=( (not A265)  and  (not A203) );
 a61502a <=( a61501a  and  a61498a );
 a61503a <=( a61502a  and  a61495a );
 a61507a <=( (not A269)  and  A267 );
 a61508a <=( A266  and  a61507a );
 a61511a <=( (not A299)  and  A298 );
 a61514a <=( (not A302)  and  A300 );
 a61515a <=( a61514a  and  a61511a );
 a61516a <=( a61515a  and  a61508a );
 a61520a <=( A199  and  A166 );
 a61521a <=( A167  and  a61520a );
 a61524a <=( A201  and  (not A200) );
 a61527a <=( (not A265)  and  (not A203) );
 a61528a <=( a61527a  and  a61524a );
 a61529a <=( a61528a  and  a61521a );
 a61533a <=( (not A269)  and  A267 );
 a61534a <=( A266  and  a61533a );
 a61537a <=( A299  and  (not A298) );
 a61540a <=( A301  and  A300 );
 a61541a <=( a61540a  and  a61537a );
 a61542a <=( a61541a  and  a61534a );
 a61546a <=( A199  and  A166 );
 a61547a <=( A167  and  a61546a );
 a61550a <=( A201  and  (not A200) );
 a61553a <=( (not A265)  and  (not A203) );
 a61554a <=( a61553a  and  a61550a );
 a61555a <=( a61554a  and  a61547a );
 a61559a <=( (not A269)  and  A267 );
 a61560a <=( A266  and  a61559a );
 a61563a <=( A299  and  (not A298) );
 a61566a <=( (not A302)  and  A300 );
 a61567a <=( a61566a  and  a61563a );
 a61568a <=( a61567a  and  a61560a );
 a61572a <=( A199  and  A166 );
 a61573a <=( A167  and  a61572a );
 a61576a <=( A201  and  (not A200) );
 a61579a <=( A265  and  (not A203) );
 a61580a <=( a61579a  and  a61576a );
 a61581a <=( a61580a  and  a61573a );
 a61585a <=( A268  and  A267 );
 a61586a <=( (not A266)  and  a61585a );
 a61589a <=( (not A299)  and  A298 );
 a61592a <=( A301  and  A300 );
 a61593a <=( a61592a  and  a61589a );
 a61594a <=( a61593a  and  a61586a );
 a61598a <=( A199  and  A166 );
 a61599a <=( A167  and  a61598a );
 a61602a <=( A201  and  (not A200) );
 a61605a <=( A265  and  (not A203) );
 a61606a <=( a61605a  and  a61602a );
 a61607a <=( a61606a  and  a61599a );
 a61611a <=( A268  and  A267 );
 a61612a <=( (not A266)  and  a61611a );
 a61615a <=( (not A299)  and  A298 );
 a61618a <=( (not A302)  and  A300 );
 a61619a <=( a61618a  and  a61615a );
 a61620a <=( a61619a  and  a61612a );
 a61624a <=( A199  and  A166 );
 a61625a <=( A167  and  a61624a );
 a61628a <=( A201  and  (not A200) );
 a61631a <=( A265  and  (not A203) );
 a61632a <=( a61631a  and  a61628a );
 a61633a <=( a61632a  and  a61625a );
 a61637a <=( A268  and  A267 );
 a61638a <=( (not A266)  and  a61637a );
 a61641a <=( A299  and  (not A298) );
 a61644a <=( A301  and  A300 );
 a61645a <=( a61644a  and  a61641a );
 a61646a <=( a61645a  and  a61638a );
 a61650a <=( A199  and  A166 );
 a61651a <=( A167  and  a61650a );
 a61654a <=( A201  and  (not A200) );
 a61657a <=( A265  and  (not A203) );
 a61658a <=( a61657a  and  a61654a );
 a61659a <=( a61658a  and  a61651a );
 a61663a <=( A268  and  A267 );
 a61664a <=( (not A266)  and  a61663a );
 a61667a <=( A299  and  (not A298) );
 a61670a <=( (not A302)  and  A300 );
 a61671a <=( a61670a  and  a61667a );
 a61672a <=( a61671a  and  a61664a );
 a61676a <=( A199  and  A166 );
 a61677a <=( A167  and  a61676a );
 a61680a <=( A201  and  (not A200) );
 a61683a <=( A265  and  (not A203) );
 a61684a <=( a61683a  and  a61680a );
 a61685a <=( a61684a  and  a61677a );
 a61689a <=( (not A269)  and  A267 );
 a61690a <=( (not A266)  and  a61689a );
 a61693a <=( (not A299)  and  A298 );
 a61696a <=( A301  and  A300 );
 a61697a <=( a61696a  and  a61693a );
 a61698a <=( a61697a  and  a61690a );
 a61702a <=( A199  and  A166 );
 a61703a <=( A167  and  a61702a );
 a61706a <=( A201  and  (not A200) );
 a61709a <=( A265  and  (not A203) );
 a61710a <=( a61709a  and  a61706a );
 a61711a <=( a61710a  and  a61703a );
 a61715a <=( (not A269)  and  A267 );
 a61716a <=( (not A266)  and  a61715a );
 a61719a <=( (not A299)  and  A298 );
 a61722a <=( (not A302)  and  A300 );
 a61723a <=( a61722a  and  a61719a );
 a61724a <=( a61723a  and  a61716a );
 a61728a <=( A199  and  A166 );
 a61729a <=( A167  and  a61728a );
 a61732a <=( A201  and  (not A200) );
 a61735a <=( A265  and  (not A203) );
 a61736a <=( a61735a  and  a61732a );
 a61737a <=( a61736a  and  a61729a );
 a61741a <=( (not A269)  and  A267 );
 a61742a <=( (not A266)  and  a61741a );
 a61745a <=( A299  and  (not A298) );
 a61748a <=( A301  and  A300 );
 a61749a <=( a61748a  and  a61745a );
 a61750a <=( a61749a  and  a61742a );
 a61754a <=( A199  and  A166 );
 a61755a <=( A167  and  a61754a );
 a61758a <=( A201  and  (not A200) );
 a61761a <=( A265  and  (not A203) );
 a61762a <=( a61761a  and  a61758a );
 a61763a <=( a61762a  and  a61755a );
 a61767a <=( (not A269)  and  A267 );
 a61768a <=( (not A266)  and  a61767a );
 a61771a <=( A299  and  (not A298) );
 a61774a <=( (not A302)  and  A300 );
 a61775a <=( a61774a  and  a61771a );
 a61776a <=( a61775a  and  a61768a );
 a61780a <=( (not A199)  and  (not A166) );
 a61781a <=( (not A167)  and  a61780a );
 a61784a <=( A201  and  A200 );
 a61787a <=( (not A265)  and  A202 );
 a61788a <=( a61787a  and  a61784a );
 a61789a <=( a61788a  and  a61781a );
 a61793a <=( A268  and  A267 );
 a61794a <=( A266  and  a61793a );
 a61797a <=( (not A299)  and  A298 );
 a61800a <=( A301  and  A300 );
 a61801a <=( a61800a  and  a61797a );
 a61802a <=( a61801a  and  a61794a );
 a61806a <=( (not A199)  and  (not A166) );
 a61807a <=( (not A167)  and  a61806a );
 a61810a <=( A201  and  A200 );
 a61813a <=( (not A265)  and  A202 );
 a61814a <=( a61813a  and  a61810a );
 a61815a <=( a61814a  and  a61807a );
 a61819a <=( A268  and  A267 );
 a61820a <=( A266  and  a61819a );
 a61823a <=( (not A299)  and  A298 );
 a61826a <=( (not A302)  and  A300 );
 a61827a <=( a61826a  and  a61823a );
 a61828a <=( a61827a  and  a61820a );
 a61832a <=( (not A199)  and  (not A166) );
 a61833a <=( (not A167)  and  a61832a );
 a61836a <=( A201  and  A200 );
 a61839a <=( (not A265)  and  A202 );
 a61840a <=( a61839a  and  a61836a );
 a61841a <=( a61840a  and  a61833a );
 a61845a <=( A268  and  A267 );
 a61846a <=( A266  and  a61845a );
 a61849a <=( A299  and  (not A298) );
 a61852a <=( A301  and  A300 );
 a61853a <=( a61852a  and  a61849a );
 a61854a <=( a61853a  and  a61846a );
 a61858a <=( (not A199)  and  (not A166) );
 a61859a <=( (not A167)  and  a61858a );
 a61862a <=( A201  and  A200 );
 a61865a <=( (not A265)  and  A202 );
 a61866a <=( a61865a  and  a61862a );
 a61867a <=( a61866a  and  a61859a );
 a61871a <=( A268  and  A267 );
 a61872a <=( A266  and  a61871a );
 a61875a <=( A299  and  (not A298) );
 a61878a <=( (not A302)  and  A300 );
 a61879a <=( a61878a  and  a61875a );
 a61880a <=( a61879a  and  a61872a );
 a61884a <=( (not A199)  and  (not A166) );
 a61885a <=( (not A167)  and  a61884a );
 a61888a <=( A201  and  A200 );
 a61891a <=( (not A265)  and  A202 );
 a61892a <=( a61891a  and  a61888a );
 a61893a <=( a61892a  and  a61885a );
 a61897a <=( (not A269)  and  A267 );
 a61898a <=( A266  and  a61897a );
 a61901a <=( (not A299)  and  A298 );
 a61904a <=( A301  and  A300 );
 a61905a <=( a61904a  and  a61901a );
 a61906a <=( a61905a  and  a61898a );
 a61910a <=( (not A199)  and  (not A166) );
 a61911a <=( (not A167)  and  a61910a );
 a61914a <=( A201  and  A200 );
 a61917a <=( (not A265)  and  A202 );
 a61918a <=( a61917a  and  a61914a );
 a61919a <=( a61918a  and  a61911a );
 a61923a <=( (not A269)  and  A267 );
 a61924a <=( A266  and  a61923a );
 a61927a <=( (not A299)  and  A298 );
 a61930a <=( (not A302)  and  A300 );
 a61931a <=( a61930a  and  a61927a );
 a61932a <=( a61931a  and  a61924a );
 a61936a <=( (not A199)  and  (not A166) );
 a61937a <=( (not A167)  and  a61936a );
 a61940a <=( A201  and  A200 );
 a61943a <=( (not A265)  and  A202 );
 a61944a <=( a61943a  and  a61940a );
 a61945a <=( a61944a  and  a61937a );
 a61949a <=( (not A269)  and  A267 );
 a61950a <=( A266  and  a61949a );
 a61953a <=( A299  and  (not A298) );
 a61956a <=( A301  and  A300 );
 a61957a <=( a61956a  and  a61953a );
 a61958a <=( a61957a  and  a61950a );
 a61962a <=( (not A199)  and  (not A166) );
 a61963a <=( (not A167)  and  a61962a );
 a61966a <=( A201  and  A200 );
 a61969a <=( (not A265)  and  A202 );
 a61970a <=( a61969a  and  a61966a );
 a61971a <=( a61970a  and  a61963a );
 a61975a <=( (not A269)  and  A267 );
 a61976a <=( A266  and  a61975a );
 a61979a <=( A299  and  (not A298) );
 a61982a <=( (not A302)  and  A300 );
 a61983a <=( a61982a  and  a61979a );
 a61984a <=( a61983a  and  a61976a );
 a61988a <=( (not A199)  and  (not A166) );
 a61989a <=( (not A167)  and  a61988a );
 a61992a <=( A201  and  A200 );
 a61995a <=( A265  and  A202 );
 a61996a <=( a61995a  and  a61992a );
 a61997a <=( a61996a  and  a61989a );
 a62001a <=( A268  and  A267 );
 a62002a <=( (not A266)  and  a62001a );
 a62005a <=( (not A299)  and  A298 );
 a62008a <=( A301  and  A300 );
 a62009a <=( a62008a  and  a62005a );
 a62010a <=( a62009a  and  a62002a );
 a62014a <=( (not A199)  and  (not A166) );
 a62015a <=( (not A167)  and  a62014a );
 a62018a <=( A201  and  A200 );
 a62021a <=( A265  and  A202 );
 a62022a <=( a62021a  and  a62018a );
 a62023a <=( a62022a  and  a62015a );
 a62027a <=( A268  and  A267 );
 a62028a <=( (not A266)  and  a62027a );
 a62031a <=( (not A299)  and  A298 );
 a62034a <=( (not A302)  and  A300 );
 a62035a <=( a62034a  and  a62031a );
 a62036a <=( a62035a  and  a62028a );
 a62040a <=( (not A199)  and  (not A166) );
 a62041a <=( (not A167)  and  a62040a );
 a62044a <=( A201  and  A200 );
 a62047a <=( A265  and  A202 );
 a62048a <=( a62047a  and  a62044a );
 a62049a <=( a62048a  and  a62041a );
 a62053a <=( A268  and  A267 );
 a62054a <=( (not A266)  and  a62053a );
 a62057a <=( A299  and  (not A298) );
 a62060a <=( A301  and  A300 );
 a62061a <=( a62060a  and  a62057a );
 a62062a <=( a62061a  and  a62054a );
 a62066a <=( (not A199)  and  (not A166) );
 a62067a <=( (not A167)  and  a62066a );
 a62070a <=( A201  and  A200 );
 a62073a <=( A265  and  A202 );
 a62074a <=( a62073a  and  a62070a );
 a62075a <=( a62074a  and  a62067a );
 a62079a <=( A268  and  A267 );
 a62080a <=( (not A266)  and  a62079a );
 a62083a <=( A299  and  (not A298) );
 a62086a <=( (not A302)  and  A300 );
 a62087a <=( a62086a  and  a62083a );
 a62088a <=( a62087a  and  a62080a );
 a62092a <=( (not A199)  and  (not A166) );
 a62093a <=( (not A167)  and  a62092a );
 a62096a <=( A201  and  A200 );
 a62099a <=( A265  and  A202 );
 a62100a <=( a62099a  and  a62096a );
 a62101a <=( a62100a  and  a62093a );
 a62105a <=( (not A269)  and  A267 );
 a62106a <=( (not A266)  and  a62105a );
 a62109a <=( (not A299)  and  A298 );
 a62112a <=( A301  and  A300 );
 a62113a <=( a62112a  and  a62109a );
 a62114a <=( a62113a  and  a62106a );
 a62118a <=( (not A199)  and  (not A166) );
 a62119a <=( (not A167)  and  a62118a );
 a62122a <=( A201  and  A200 );
 a62125a <=( A265  and  A202 );
 a62126a <=( a62125a  and  a62122a );
 a62127a <=( a62126a  and  a62119a );
 a62131a <=( (not A269)  and  A267 );
 a62132a <=( (not A266)  and  a62131a );
 a62135a <=( (not A299)  and  A298 );
 a62138a <=( (not A302)  and  A300 );
 a62139a <=( a62138a  and  a62135a );
 a62140a <=( a62139a  and  a62132a );
 a62144a <=( (not A199)  and  (not A166) );
 a62145a <=( (not A167)  and  a62144a );
 a62148a <=( A201  and  A200 );
 a62151a <=( A265  and  A202 );
 a62152a <=( a62151a  and  a62148a );
 a62153a <=( a62152a  and  a62145a );
 a62157a <=( (not A269)  and  A267 );
 a62158a <=( (not A266)  and  a62157a );
 a62161a <=( A299  and  (not A298) );
 a62164a <=( A301  and  A300 );
 a62165a <=( a62164a  and  a62161a );
 a62166a <=( a62165a  and  a62158a );
 a62170a <=( (not A199)  and  (not A166) );
 a62171a <=( (not A167)  and  a62170a );
 a62174a <=( A201  and  A200 );
 a62177a <=( A265  and  A202 );
 a62178a <=( a62177a  and  a62174a );
 a62179a <=( a62178a  and  a62171a );
 a62183a <=( (not A269)  and  A267 );
 a62184a <=( (not A266)  and  a62183a );
 a62187a <=( A299  and  (not A298) );
 a62190a <=( (not A302)  and  A300 );
 a62191a <=( a62190a  and  a62187a );
 a62192a <=( a62191a  and  a62184a );
 a62196a <=( (not A199)  and  (not A166) );
 a62197a <=( (not A167)  and  a62196a );
 a62200a <=( A201  and  A200 );
 a62203a <=( (not A265)  and  (not A203) );
 a62204a <=( a62203a  and  a62200a );
 a62205a <=( a62204a  and  a62197a );
 a62209a <=( A268  and  A267 );
 a62210a <=( A266  and  a62209a );
 a62213a <=( (not A299)  and  A298 );
 a62216a <=( A301  and  A300 );
 a62217a <=( a62216a  and  a62213a );
 a62218a <=( a62217a  and  a62210a );
 a62222a <=( (not A199)  and  (not A166) );
 a62223a <=( (not A167)  and  a62222a );
 a62226a <=( A201  and  A200 );
 a62229a <=( (not A265)  and  (not A203) );
 a62230a <=( a62229a  and  a62226a );
 a62231a <=( a62230a  and  a62223a );
 a62235a <=( A268  and  A267 );
 a62236a <=( A266  and  a62235a );
 a62239a <=( (not A299)  and  A298 );
 a62242a <=( (not A302)  and  A300 );
 a62243a <=( a62242a  and  a62239a );
 a62244a <=( a62243a  and  a62236a );
 a62248a <=( (not A199)  and  (not A166) );
 a62249a <=( (not A167)  and  a62248a );
 a62252a <=( A201  and  A200 );
 a62255a <=( (not A265)  and  (not A203) );
 a62256a <=( a62255a  and  a62252a );
 a62257a <=( a62256a  and  a62249a );
 a62261a <=( A268  and  A267 );
 a62262a <=( A266  and  a62261a );
 a62265a <=( A299  and  (not A298) );
 a62268a <=( A301  and  A300 );
 a62269a <=( a62268a  and  a62265a );
 a62270a <=( a62269a  and  a62262a );
 a62274a <=( (not A199)  and  (not A166) );
 a62275a <=( (not A167)  and  a62274a );
 a62278a <=( A201  and  A200 );
 a62281a <=( (not A265)  and  (not A203) );
 a62282a <=( a62281a  and  a62278a );
 a62283a <=( a62282a  and  a62275a );
 a62287a <=( A268  and  A267 );
 a62288a <=( A266  and  a62287a );
 a62291a <=( A299  and  (not A298) );
 a62294a <=( (not A302)  and  A300 );
 a62295a <=( a62294a  and  a62291a );
 a62296a <=( a62295a  and  a62288a );
 a62300a <=( (not A199)  and  (not A166) );
 a62301a <=( (not A167)  and  a62300a );
 a62304a <=( A201  and  A200 );
 a62307a <=( (not A265)  and  (not A203) );
 a62308a <=( a62307a  and  a62304a );
 a62309a <=( a62308a  and  a62301a );
 a62313a <=( (not A269)  and  A267 );
 a62314a <=( A266  and  a62313a );
 a62317a <=( (not A299)  and  A298 );
 a62320a <=( A301  and  A300 );
 a62321a <=( a62320a  and  a62317a );
 a62322a <=( a62321a  and  a62314a );
 a62326a <=( (not A199)  and  (not A166) );
 a62327a <=( (not A167)  and  a62326a );
 a62330a <=( A201  and  A200 );
 a62333a <=( (not A265)  and  (not A203) );
 a62334a <=( a62333a  and  a62330a );
 a62335a <=( a62334a  and  a62327a );
 a62339a <=( (not A269)  and  A267 );
 a62340a <=( A266  and  a62339a );
 a62343a <=( (not A299)  and  A298 );
 a62346a <=( (not A302)  and  A300 );
 a62347a <=( a62346a  and  a62343a );
 a62348a <=( a62347a  and  a62340a );
 a62352a <=( (not A199)  and  (not A166) );
 a62353a <=( (not A167)  and  a62352a );
 a62356a <=( A201  and  A200 );
 a62359a <=( (not A265)  and  (not A203) );
 a62360a <=( a62359a  and  a62356a );
 a62361a <=( a62360a  and  a62353a );
 a62365a <=( (not A269)  and  A267 );
 a62366a <=( A266  and  a62365a );
 a62369a <=( A299  and  (not A298) );
 a62372a <=( A301  and  A300 );
 a62373a <=( a62372a  and  a62369a );
 a62374a <=( a62373a  and  a62366a );
 a62378a <=( (not A199)  and  (not A166) );
 a62379a <=( (not A167)  and  a62378a );
 a62382a <=( A201  and  A200 );
 a62385a <=( (not A265)  and  (not A203) );
 a62386a <=( a62385a  and  a62382a );
 a62387a <=( a62386a  and  a62379a );
 a62391a <=( (not A269)  and  A267 );
 a62392a <=( A266  and  a62391a );
 a62395a <=( A299  and  (not A298) );
 a62398a <=( (not A302)  and  A300 );
 a62399a <=( a62398a  and  a62395a );
 a62400a <=( a62399a  and  a62392a );
 a62404a <=( (not A199)  and  (not A166) );
 a62405a <=( (not A167)  and  a62404a );
 a62408a <=( A201  and  A200 );
 a62411a <=( A265  and  (not A203) );
 a62412a <=( a62411a  and  a62408a );
 a62413a <=( a62412a  and  a62405a );
 a62417a <=( A268  and  A267 );
 a62418a <=( (not A266)  and  a62417a );
 a62421a <=( (not A299)  and  A298 );
 a62424a <=( A301  and  A300 );
 a62425a <=( a62424a  and  a62421a );
 a62426a <=( a62425a  and  a62418a );
 a62430a <=( (not A199)  and  (not A166) );
 a62431a <=( (not A167)  and  a62430a );
 a62434a <=( A201  and  A200 );
 a62437a <=( A265  and  (not A203) );
 a62438a <=( a62437a  and  a62434a );
 a62439a <=( a62438a  and  a62431a );
 a62443a <=( A268  and  A267 );
 a62444a <=( (not A266)  and  a62443a );
 a62447a <=( (not A299)  and  A298 );
 a62450a <=( (not A302)  and  A300 );
 a62451a <=( a62450a  and  a62447a );
 a62452a <=( a62451a  and  a62444a );
 a62456a <=( (not A199)  and  (not A166) );
 a62457a <=( (not A167)  and  a62456a );
 a62460a <=( A201  and  A200 );
 a62463a <=( A265  and  (not A203) );
 a62464a <=( a62463a  and  a62460a );
 a62465a <=( a62464a  and  a62457a );
 a62469a <=( A268  and  A267 );
 a62470a <=( (not A266)  and  a62469a );
 a62473a <=( A299  and  (not A298) );
 a62476a <=( A301  and  A300 );
 a62477a <=( a62476a  and  a62473a );
 a62478a <=( a62477a  and  a62470a );
 a62482a <=( (not A199)  and  (not A166) );
 a62483a <=( (not A167)  and  a62482a );
 a62486a <=( A201  and  A200 );
 a62489a <=( A265  and  (not A203) );
 a62490a <=( a62489a  and  a62486a );
 a62491a <=( a62490a  and  a62483a );
 a62495a <=( A268  and  A267 );
 a62496a <=( (not A266)  and  a62495a );
 a62499a <=( A299  and  (not A298) );
 a62502a <=( (not A302)  and  A300 );
 a62503a <=( a62502a  and  a62499a );
 a62504a <=( a62503a  and  a62496a );
 a62508a <=( (not A199)  and  (not A166) );
 a62509a <=( (not A167)  and  a62508a );
 a62512a <=( A201  and  A200 );
 a62515a <=( A265  and  (not A203) );
 a62516a <=( a62515a  and  a62512a );
 a62517a <=( a62516a  and  a62509a );
 a62521a <=( (not A269)  and  A267 );
 a62522a <=( (not A266)  and  a62521a );
 a62525a <=( (not A299)  and  A298 );
 a62528a <=( A301  and  A300 );
 a62529a <=( a62528a  and  a62525a );
 a62530a <=( a62529a  and  a62522a );
 a62534a <=( (not A199)  and  (not A166) );
 a62535a <=( (not A167)  and  a62534a );
 a62538a <=( A201  and  A200 );
 a62541a <=( A265  and  (not A203) );
 a62542a <=( a62541a  and  a62538a );
 a62543a <=( a62542a  and  a62535a );
 a62547a <=( (not A269)  and  A267 );
 a62548a <=( (not A266)  and  a62547a );
 a62551a <=( (not A299)  and  A298 );
 a62554a <=( (not A302)  and  A300 );
 a62555a <=( a62554a  and  a62551a );
 a62556a <=( a62555a  and  a62548a );
 a62560a <=( (not A199)  and  (not A166) );
 a62561a <=( (not A167)  and  a62560a );
 a62564a <=( A201  and  A200 );
 a62567a <=( A265  and  (not A203) );
 a62568a <=( a62567a  and  a62564a );
 a62569a <=( a62568a  and  a62561a );
 a62573a <=( (not A269)  and  A267 );
 a62574a <=( (not A266)  and  a62573a );
 a62577a <=( A299  and  (not A298) );
 a62580a <=( A301  and  A300 );
 a62581a <=( a62580a  and  a62577a );
 a62582a <=( a62581a  and  a62574a );
 a62586a <=( (not A199)  and  (not A166) );
 a62587a <=( (not A167)  and  a62586a );
 a62590a <=( A201  and  A200 );
 a62593a <=( A265  and  (not A203) );
 a62594a <=( a62593a  and  a62590a );
 a62595a <=( a62594a  and  a62587a );
 a62599a <=( (not A269)  and  A267 );
 a62600a <=( (not A266)  and  a62599a );
 a62603a <=( A299  and  (not A298) );
 a62606a <=( (not A302)  and  A300 );
 a62607a <=( a62606a  and  a62603a );
 a62608a <=( a62607a  and  a62600a );
 a62612a <=( A199  and  (not A166) );
 a62613a <=( (not A167)  and  a62612a );
 a62616a <=( A201  and  (not A200) );
 a62619a <=( (not A265)  and  A202 );
 a62620a <=( a62619a  and  a62616a );
 a62621a <=( a62620a  and  a62613a );
 a62625a <=( A268  and  A267 );
 a62626a <=( A266  and  a62625a );
 a62629a <=( (not A299)  and  A298 );
 a62632a <=( A301  and  A300 );
 a62633a <=( a62632a  and  a62629a );
 a62634a <=( a62633a  and  a62626a );
 a62638a <=( A199  and  (not A166) );
 a62639a <=( (not A167)  and  a62638a );
 a62642a <=( A201  and  (not A200) );
 a62645a <=( (not A265)  and  A202 );
 a62646a <=( a62645a  and  a62642a );
 a62647a <=( a62646a  and  a62639a );
 a62651a <=( A268  and  A267 );
 a62652a <=( A266  and  a62651a );
 a62655a <=( (not A299)  and  A298 );
 a62658a <=( (not A302)  and  A300 );
 a62659a <=( a62658a  and  a62655a );
 a62660a <=( a62659a  and  a62652a );
 a62664a <=( A199  and  (not A166) );
 a62665a <=( (not A167)  and  a62664a );
 a62668a <=( A201  and  (not A200) );
 a62671a <=( (not A265)  and  A202 );
 a62672a <=( a62671a  and  a62668a );
 a62673a <=( a62672a  and  a62665a );
 a62677a <=( A268  and  A267 );
 a62678a <=( A266  and  a62677a );
 a62681a <=( A299  and  (not A298) );
 a62684a <=( A301  and  A300 );
 a62685a <=( a62684a  and  a62681a );
 a62686a <=( a62685a  and  a62678a );
 a62690a <=( A199  and  (not A166) );
 a62691a <=( (not A167)  and  a62690a );
 a62694a <=( A201  and  (not A200) );
 a62697a <=( (not A265)  and  A202 );
 a62698a <=( a62697a  and  a62694a );
 a62699a <=( a62698a  and  a62691a );
 a62703a <=( A268  and  A267 );
 a62704a <=( A266  and  a62703a );
 a62707a <=( A299  and  (not A298) );
 a62710a <=( (not A302)  and  A300 );
 a62711a <=( a62710a  and  a62707a );
 a62712a <=( a62711a  and  a62704a );
 a62716a <=( A199  and  (not A166) );
 a62717a <=( (not A167)  and  a62716a );
 a62720a <=( A201  and  (not A200) );
 a62723a <=( (not A265)  and  A202 );
 a62724a <=( a62723a  and  a62720a );
 a62725a <=( a62724a  and  a62717a );
 a62729a <=( (not A269)  and  A267 );
 a62730a <=( A266  and  a62729a );
 a62733a <=( (not A299)  and  A298 );
 a62736a <=( A301  and  A300 );
 a62737a <=( a62736a  and  a62733a );
 a62738a <=( a62737a  and  a62730a );
 a62742a <=( A199  and  (not A166) );
 a62743a <=( (not A167)  and  a62742a );
 a62746a <=( A201  and  (not A200) );
 a62749a <=( (not A265)  and  A202 );
 a62750a <=( a62749a  and  a62746a );
 a62751a <=( a62750a  and  a62743a );
 a62755a <=( (not A269)  and  A267 );
 a62756a <=( A266  and  a62755a );
 a62759a <=( (not A299)  and  A298 );
 a62762a <=( (not A302)  and  A300 );
 a62763a <=( a62762a  and  a62759a );
 a62764a <=( a62763a  and  a62756a );
 a62768a <=( A199  and  (not A166) );
 a62769a <=( (not A167)  and  a62768a );
 a62772a <=( A201  and  (not A200) );
 a62775a <=( (not A265)  and  A202 );
 a62776a <=( a62775a  and  a62772a );
 a62777a <=( a62776a  and  a62769a );
 a62781a <=( (not A269)  and  A267 );
 a62782a <=( A266  and  a62781a );
 a62785a <=( A299  and  (not A298) );
 a62788a <=( A301  and  A300 );
 a62789a <=( a62788a  and  a62785a );
 a62790a <=( a62789a  and  a62782a );
 a62794a <=( A199  and  (not A166) );
 a62795a <=( (not A167)  and  a62794a );
 a62798a <=( A201  and  (not A200) );
 a62801a <=( (not A265)  and  A202 );
 a62802a <=( a62801a  and  a62798a );
 a62803a <=( a62802a  and  a62795a );
 a62807a <=( (not A269)  and  A267 );
 a62808a <=( A266  and  a62807a );
 a62811a <=( A299  and  (not A298) );
 a62814a <=( (not A302)  and  A300 );
 a62815a <=( a62814a  and  a62811a );
 a62816a <=( a62815a  and  a62808a );
 a62820a <=( A199  and  (not A166) );
 a62821a <=( (not A167)  and  a62820a );
 a62824a <=( A201  and  (not A200) );
 a62827a <=( A265  and  A202 );
 a62828a <=( a62827a  and  a62824a );
 a62829a <=( a62828a  and  a62821a );
 a62833a <=( A268  and  A267 );
 a62834a <=( (not A266)  and  a62833a );
 a62837a <=( (not A299)  and  A298 );
 a62840a <=( A301  and  A300 );
 a62841a <=( a62840a  and  a62837a );
 a62842a <=( a62841a  and  a62834a );
 a62846a <=( A199  and  (not A166) );
 a62847a <=( (not A167)  and  a62846a );
 a62850a <=( A201  and  (not A200) );
 a62853a <=( A265  and  A202 );
 a62854a <=( a62853a  and  a62850a );
 a62855a <=( a62854a  and  a62847a );
 a62859a <=( A268  and  A267 );
 a62860a <=( (not A266)  and  a62859a );
 a62863a <=( (not A299)  and  A298 );
 a62866a <=( (not A302)  and  A300 );
 a62867a <=( a62866a  and  a62863a );
 a62868a <=( a62867a  and  a62860a );
 a62872a <=( A199  and  (not A166) );
 a62873a <=( (not A167)  and  a62872a );
 a62876a <=( A201  and  (not A200) );
 a62879a <=( A265  and  A202 );
 a62880a <=( a62879a  and  a62876a );
 a62881a <=( a62880a  and  a62873a );
 a62885a <=( A268  and  A267 );
 a62886a <=( (not A266)  and  a62885a );
 a62889a <=( A299  and  (not A298) );
 a62892a <=( A301  and  A300 );
 a62893a <=( a62892a  and  a62889a );
 a62894a <=( a62893a  and  a62886a );
 a62898a <=( A199  and  (not A166) );
 a62899a <=( (not A167)  and  a62898a );
 a62902a <=( A201  and  (not A200) );
 a62905a <=( A265  and  A202 );
 a62906a <=( a62905a  and  a62902a );
 a62907a <=( a62906a  and  a62899a );
 a62911a <=( A268  and  A267 );
 a62912a <=( (not A266)  and  a62911a );
 a62915a <=( A299  and  (not A298) );
 a62918a <=( (not A302)  and  A300 );
 a62919a <=( a62918a  and  a62915a );
 a62920a <=( a62919a  and  a62912a );
 a62924a <=( A199  and  (not A166) );
 a62925a <=( (not A167)  and  a62924a );
 a62928a <=( A201  and  (not A200) );
 a62931a <=( A265  and  A202 );
 a62932a <=( a62931a  and  a62928a );
 a62933a <=( a62932a  and  a62925a );
 a62937a <=( (not A269)  and  A267 );
 a62938a <=( (not A266)  and  a62937a );
 a62941a <=( (not A299)  and  A298 );
 a62944a <=( A301  and  A300 );
 a62945a <=( a62944a  and  a62941a );
 a62946a <=( a62945a  and  a62938a );
 a62950a <=( A199  and  (not A166) );
 a62951a <=( (not A167)  and  a62950a );
 a62954a <=( A201  and  (not A200) );
 a62957a <=( A265  and  A202 );
 a62958a <=( a62957a  and  a62954a );
 a62959a <=( a62958a  and  a62951a );
 a62963a <=( (not A269)  and  A267 );
 a62964a <=( (not A266)  and  a62963a );
 a62967a <=( (not A299)  and  A298 );
 a62970a <=( (not A302)  and  A300 );
 a62971a <=( a62970a  and  a62967a );
 a62972a <=( a62971a  and  a62964a );
 a62976a <=( A199  and  (not A166) );
 a62977a <=( (not A167)  and  a62976a );
 a62980a <=( A201  and  (not A200) );
 a62983a <=( A265  and  A202 );
 a62984a <=( a62983a  and  a62980a );
 a62985a <=( a62984a  and  a62977a );
 a62989a <=( (not A269)  and  A267 );
 a62990a <=( (not A266)  and  a62989a );
 a62993a <=( A299  and  (not A298) );
 a62996a <=( A301  and  A300 );
 a62997a <=( a62996a  and  a62993a );
 a62998a <=( a62997a  and  a62990a );
 a63002a <=( A199  and  (not A166) );
 a63003a <=( (not A167)  and  a63002a );
 a63006a <=( A201  and  (not A200) );
 a63009a <=( A265  and  A202 );
 a63010a <=( a63009a  and  a63006a );
 a63011a <=( a63010a  and  a63003a );
 a63015a <=( (not A269)  and  A267 );
 a63016a <=( (not A266)  and  a63015a );
 a63019a <=( A299  and  (not A298) );
 a63022a <=( (not A302)  and  A300 );
 a63023a <=( a63022a  and  a63019a );
 a63024a <=( a63023a  and  a63016a );
 a63028a <=( A199  and  (not A166) );
 a63029a <=( (not A167)  and  a63028a );
 a63032a <=( A201  and  (not A200) );
 a63035a <=( (not A265)  and  (not A203) );
 a63036a <=( a63035a  and  a63032a );
 a63037a <=( a63036a  and  a63029a );
 a63041a <=( A268  and  A267 );
 a63042a <=( A266  and  a63041a );
 a63045a <=( (not A299)  and  A298 );
 a63048a <=( A301  and  A300 );
 a63049a <=( a63048a  and  a63045a );
 a63050a <=( a63049a  and  a63042a );
 a63054a <=( A199  and  (not A166) );
 a63055a <=( (not A167)  and  a63054a );
 a63058a <=( A201  and  (not A200) );
 a63061a <=( (not A265)  and  (not A203) );
 a63062a <=( a63061a  and  a63058a );
 a63063a <=( a63062a  and  a63055a );
 a63067a <=( A268  and  A267 );
 a63068a <=( A266  and  a63067a );
 a63071a <=( (not A299)  and  A298 );
 a63074a <=( (not A302)  and  A300 );
 a63075a <=( a63074a  and  a63071a );
 a63076a <=( a63075a  and  a63068a );
 a63080a <=( A199  and  (not A166) );
 a63081a <=( (not A167)  and  a63080a );
 a63084a <=( A201  and  (not A200) );
 a63087a <=( (not A265)  and  (not A203) );
 a63088a <=( a63087a  and  a63084a );
 a63089a <=( a63088a  and  a63081a );
 a63093a <=( A268  and  A267 );
 a63094a <=( A266  and  a63093a );
 a63097a <=( A299  and  (not A298) );
 a63100a <=( A301  and  A300 );
 a63101a <=( a63100a  and  a63097a );
 a63102a <=( a63101a  and  a63094a );
 a63106a <=( A199  and  (not A166) );
 a63107a <=( (not A167)  and  a63106a );
 a63110a <=( A201  and  (not A200) );
 a63113a <=( (not A265)  and  (not A203) );
 a63114a <=( a63113a  and  a63110a );
 a63115a <=( a63114a  and  a63107a );
 a63119a <=( A268  and  A267 );
 a63120a <=( A266  and  a63119a );
 a63123a <=( A299  and  (not A298) );
 a63126a <=( (not A302)  and  A300 );
 a63127a <=( a63126a  and  a63123a );
 a63128a <=( a63127a  and  a63120a );
 a63132a <=( A199  and  (not A166) );
 a63133a <=( (not A167)  and  a63132a );
 a63136a <=( A201  and  (not A200) );
 a63139a <=( (not A265)  and  (not A203) );
 a63140a <=( a63139a  and  a63136a );
 a63141a <=( a63140a  and  a63133a );
 a63145a <=( (not A269)  and  A267 );
 a63146a <=( A266  and  a63145a );
 a63149a <=( (not A299)  and  A298 );
 a63152a <=( A301  and  A300 );
 a63153a <=( a63152a  and  a63149a );
 a63154a <=( a63153a  and  a63146a );
 a63158a <=( A199  and  (not A166) );
 a63159a <=( (not A167)  and  a63158a );
 a63162a <=( A201  and  (not A200) );
 a63165a <=( (not A265)  and  (not A203) );
 a63166a <=( a63165a  and  a63162a );
 a63167a <=( a63166a  and  a63159a );
 a63171a <=( (not A269)  and  A267 );
 a63172a <=( A266  and  a63171a );
 a63175a <=( (not A299)  and  A298 );
 a63178a <=( (not A302)  and  A300 );
 a63179a <=( a63178a  and  a63175a );
 a63180a <=( a63179a  and  a63172a );
 a63184a <=( A199  and  (not A166) );
 a63185a <=( (not A167)  and  a63184a );
 a63188a <=( A201  and  (not A200) );
 a63191a <=( (not A265)  and  (not A203) );
 a63192a <=( a63191a  and  a63188a );
 a63193a <=( a63192a  and  a63185a );
 a63197a <=( (not A269)  and  A267 );
 a63198a <=( A266  and  a63197a );
 a63201a <=( A299  and  (not A298) );
 a63204a <=( A301  and  A300 );
 a63205a <=( a63204a  and  a63201a );
 a63206a <=( a63205a  and  a63198a );
 a63210a <=( A199  and  (not A166) );
 a63211a <=( (not A167)  and  a63210a );
 a63214a <=( A201  and  (not A200) );
 a63217a <=( (not A265)  and  (not A203) );
 a63218a <=( a63217a  and  a63214a );
 a63219a <=( a63218a  and  a63211a );
 a63223a <=( (not A269)  and  A267 );
 a63224a <=( A266  and  a63223a );
 a63227a <=( A299  and  (not A298) );
 a63230a <=( (not A302)  and  A300 );
 a63231a <=( a63230a  and  a63227a );
 a63232a <=( a63231a  and  a63224a );
 a63236a <=( A199  and  (not A166) );
 a63237a <=( (not A167)  and  a63236a );
 a63240a <=( A201  and  (not A200) );
 a63243a <=( A265  and  (not A203) );
 a63244a <=( a63243a  and  a63240a );
 a63245a <=( a63244a  and  a63237a );
 a63249a <=( A268  and  A267 );
 a63250a <=( (not A266)  and  a63249a );
 a63253a <=( (not A299)  and  A298 );
 a63256a <=( A301  and  A300 );
 a63257a <=( a63256a  and  a63253a );
 a63258a <=( a63257a  and  a63250a );
 a63262a <=( A199  and  (not A166) );
 a63263a <=( (not A167)  and  a63262a );
 a63266a <=( A201  and  (not A200) );
 a63269a <=( A265  and  (not A203) );
 a63270a <=( a63269a  and  a63266a );
 a63271a <=( a63270a  and  a63263a );
 a63275a <=( A268  and  A267 );
 a63276a <=( (not A266)  and  a63275a );
 a63279a <=( (not A299)  and  A298 );
 a63282a <=( (not A302)  and  A300 );
 a63283a <=( a63282a  and  a63279a );
 a63284a <=( a63283a  and  a63276a );
 a63288a <=( A199  and  (not A166) );
 a63289a <=( (not A167)  and  a63288a );
 a63292a <=( A201  and  (not A200) );
 a63295a <=( A265  and  (not A203) );
 a63296a <=( a63295a  and  a63292a );
 a63297a <=( a63296a  and  a63289a );
 a63301a <=( A268  and  A267 );
 a63302a <=( (not A266)  and  a63301a );
 a63305a <=( A299  and  (not A298) );
 a63308a <=( A301  and  A300 );
 a63309a <=( a63308a  and  a63305a );
 a63310a <=( a63309a  and  a63302a );
 a63314a <=( A199  and  (not A166) );
 a63315a <=( (not A167)  and  a63314a );
 a63318a <=( A201  and  (not A200) );
 a63321a <=( A265  and  (not A203) );
 a63322a <=( a63321a  and  a63318a );
 a63323a <=( a63322a  and  a63315a );
 a63327a <=( A268  and  A267 );
 a63328a <=( (not A266)  and  a63327a );
 a63331a <=( A299  and  (not A298) );
 a63334a <=( (not A302)  and  A300 );
 a63335a <=( a63334a  and  a63331a );
 a63336a <=( a63335a  and  a63328a );
 a63340a <=( A199  and  (not A166) );
 a63341a <=( (not A167)  and  a63340a );
 a63344a <=( A201  and  (not A200) );
 a63347a <=( A265  and  (not A203) );
 a63348a <=( a63347a  and  a63344a );
 a63349a <=( a63348a  and  a63341a );
 a63353a <=( (not A269)  and  A267 );
 a63354a <=( (not A266)  and  a63353a );
 a63357a <=( (not A299)  and  A298 );
 a63360a <=( A301  and  A300 );
 a63361a <=( a63360a  and  a63357a );
 a63362a <=( a63361a  and  a63354a );
 a63366a <=( A199  and  (not A166) );
 a63367a <=( (not A167)  and  a63366a );
 a63370a <=( A201  and  (not A200) );
 a63373a <=( A265  and  (not A203) );
 a63374a <=( a63373a  and  a63370a );
 a63375a <=( a63374a  and  a63367a );
 a63379a <=( (not A269)  and  A267 );
 a63380a <=( (not A266)  and  a63379a );
 a63383a <=( (not A299)  and  A298 );
 a63386a <=( (not A302)  and  A300 );
 a63387a <=( a63386a  and  a63383a );
 a63388a <=( a63387a  and  a63380a );
 a63392a <=( A199  and  (not A166) );
 a63393a <=( (not A167)  and  a63392a );
 a63396a <=( A201  and  (not A200) );
 a63399a <=( A265  and  (not A203) );
 a63400a <=( a63399a  and  a63396a );
 a63401a <=( a63400a  and  a63393a );
 a63405a <=( (not A269)  and  A267 );
 a63406a <=( (not A266)  and  a63405a );
 a63409a <=( A299  and  (not A298) );
 a63412a <=( A301  and  A300 );
 a63413a <=( a63412a  and  a63409a );
 a63414a <=( a63413a  and  a63406a );
 a63418a <=( A199  and  (not A166) );
 a63419a <=( (not A167)  and  a63418a );
 a63422a <=( A201  and  (not A200) );
 a63425a <=( A265  and  (not A203) );
 a63426a <=( a63425a  and  a63422a );
 a63427a <=( a63426a  and  a63419a );
 a63431a <=( (not A269)  and  A267 );
 a63432a <=( (not A266)  and  a63431a );
 a63435a <=( A299  and  (not A298) );
 a63438a <=( (not A302)  and  A300 );
 a63439a <=( a63438a  and  a63435a );
 a63440a <=( a63439a  and  a63432a );
 a63444a <=( A167  and  A168 );
 a63445a <=( A170  and  a63444a );
 a63448a <=( A201  and  (not A166) );
 a63451a <=( A203  and  (not A202) );
 a63452a <=( a63451a  and  a63448a );
 a63453a <=( a63452a  and  a63445a );
 a63457a <=( A269  and  (not A268) );
 a63458a <=( A267  and  a63457a );
 a63461a <=( (not A299)  and  A298 );
 a63464a <=( A301  and  A300 );
 a63465a <=( a63464a  and  a63461a );
 a63466a <=( a63465a  and  a63458a );
 a63470a <=( A167  and  A168 );
 a63471a <=( A170  and  a63470a );
 a63474a <=( A201  and  (not A166) );
 a63477a <=( A203  and  (not A202) );
 a63478a <=( a63477a  and  a63474a );
 a63479a <=( a63478a  and  a63471a );
 a63483a <=( A269  and  (not A268) );
 a63484a <=( A267  and  a63483a );
 a63487a <=( (not A299)  and  A298 );
 a63490a <=( (not A302)  and  A300 );
 a63491a <=( a63490a  and  a63487a );
 a63492a <=( a63491a  and  a63484a );
 a63496a <=( A167  and  A168 );
 a63497a <=( A170  and  a63496a );
 a63500a <=( A201  and  (not A166) );
 a63503a <=( A203  and  (not A202) );
 a63504a <=( a63503a  and  a63500a );
 a63505a <=( a63504a  and  a63497a );
 a63509a <=( A269  and  (not A268) );
 a63510a <=( A267  and  a63509a );
 a63513a <=( A299  and  (not A298) );
 a63516a <=( A301  and  A300 );
 a63517a <=( a63516a  and  a63513a );
 a63518a <=( a63517a  and  a63510a );
 a63522a <=( A167  and  A168 );
 a63523a <=( A170  and  a63522a );
 a63526a <=( A201  and  (not A166) );
 a63529a <=( A203  and  (not A202) );
 a63530a <=( a63529a  and  a63526a );
 a63531a <=( a63530a  and  a63523a );
 a63535a <=( A269  and  (not A268) );
 a63536a <=( A267  and  a63535a );
 a63539a <=( A299  and  (not A298) );
 a63542a <=( (not A302)  and  A300 );
 a63543a <=( a63542a  and  a63539a );
 a63544a <=( a63543a  and  a63536a );
 a63548a <=( A167  and  A168 );
 a63549a <=( A170  and  a63548a );
 a63552a <=( A201  and  (not A166) );
 a63555a <=( A203  and  (not A202) );
 a63556a <=( a63555a  and  a63552a );
 a63557a <=( a63556a  and  a63549a );
 a63561a <=( A298  and  A268 );
 a63562a <=( (not A267)  and  a63561a );
 a63565a <=( (not A300)  and  (not A299) );
 a63568a <=( A302  and  (not A301) );
 a63569a <=( a63568a  and  a63565a );
 a63570a <=( a63569a  and  a63562a );
 a63574a <=( A167  and  A168 );
 a63575a <=( A170  and  a63574a );
 a63578a <=( A201  and  (not A166) );
 a63581a <=( A203  and  (not A202) );
 a63582a <=( a63581a  and  a63578a );
 a63583a <=( a63582a  and  a63575a );
 a63587a <=( (not A298)  and  A268 );
 a63588a <=( (not A267)  and  a63587a );
 a63591a <=( (not A300)  and  A299 );
 a63594a <=( A302  and  (not A301) );
 a63595a <=( a63594a  and  a63591a );
 a63596a <=( a63595a  and  a63588a );
 a63600a <=( A167  and  A168 );
 a63601a <=( A170  and  a63600a );
 a63604a <=( A201  and  (not A166) );
 a63607a <=( A203  and  (not A202) );
 a63608a <=( a63607a  and  a63604a );
 a63609a <=( a63608a  and  a63601a );
 a63613a <=( A298  and  (not A269) );
 a63614a <=( (not A267)  and  a63613a );
 a63617a <=( (not A300)  and  (not A299) );
 a63620a <=( A302  and  (not A301) );
 a63621a <=( a63620a  and  a63617a );
 a63622a <=( a63621a  and  a63614a );
 a63626a <=( A167  and  A168 );
 a63627a <=( A170  and  a63626a );
 a63630a <=( A201  and  (not A166) );
 a63633a <=( A203  and  (not A202) );
 a63634a <=( a63633a  and  a63630a );
 a63635a <=( a63634a  and  a63627a );
 a63639a <=( (not A298)  and  (not A269) );
 a63640a <=( (not A267)  and  a63639a );
 a63643a <=( (not A300)  and  A299 );
 a63646a <=( A302  and  (not A301) );
 a63647a <=( a63646a  and  a63643a );
 a63648a <=( a63647a  and  a63640a );
 a63652a <=( A167  and  A168 );
 a63653a <=( A170  and  a63652a );
 a63656a <=( A201  and  (not A166) );
 a63659a <=( A203  and  (not A202) );
 a63660a <=( a63659a  and  a63656a );
 a63661a <=( a63660a  and  a63653a );
 a63665a <=( A298  and  A266 );
 a63666a <=( A265  and  a63665a );
 a63669a <=( (not A300)  and  (not A299) );
 a63672a <=( A302  and  (not A301) );
 a63673a <=( a63672a  and  a63669a );
 a63674a <=( a63673a  and  a63666a );
 a63678a <=( A167  and  A168 );
 a63679a <=( A170  and  a63678a );
 a63682a <=( A201  and  (not A166) );
 a63685a <=( A203  and  (not A202) );
 a63686a <=( a63685a  and  a63682a );
 a63687a <=( a63686a  and  a63679a );
 a63691a <=( (not A298)  and  A266 );
 a63692a <=( A265  and  a63691a );
 a63695a <=( (not A300)  and  A299 );
 a63698a <=( A302  and  (not A301) );
 a63699a <=( a63698a  and  a63695a );
 a63700a <=( a63699a  and  a63692a );
 a63704a <=( A167  and  A168 );
 a63705a <=( A170  and  a63704a );
 a63708a <=( A201  and  (not A166) );
 a63711a <=( A203  and  (not A202) );
 a63712a <=( a63711a  and  a63708a );
 a63713a <=( a63712a  and  a63705a );
 a63717a <=( A267  and  A266 );
 a63718a <=( (not A265)  and  a63717a );
 a63721a <=( A300  and  A268 );
 a63724a <=( A302  and  (not A301) );
 a63725a <=( a63724a  and  a63721a );
 a63726a <=( a63725a  and  a63718a );
 a63730a <=( A167  and  A168 );
 a63731a <=( A170  and  a63730a );
 a63734a <=( A201  and  (not A166) );
 a63737a <=( A203  and  (not A202) );
 a63738a <=( a63737a  and  a63734a );
 a63739a <=( a63738a  and  a63731a );
 a63743a <=( A267  and  A266 );
 a63744a <=( (not A265)  and  a63743a );
 a63747a <=( A300  and  (not A269) );
 a63750a <=( A302  and  (not A301) );
 a63751a <=( a63750a  and  a63747a );
 a63752a <=( a63751a  and  a63744a );
 a63756a <=( A167  and  A168 );
 a63757a <=( A170  and  a63756a );
 a63760a <=( A201  and  (not A166) );
 a63763a <=( A203  and  (not A202) );
 a63764a <=( a63763a  and  a63760a );
 a63765a <=( a63764a  and  a63757a );
 a63769a <=( (not A267)  and  A266 );
 a63770a <=( (not A265)  and  a63769a );
 a63773a <=( A269  and  (not A268) );
 a63776a <=( A301  and  (not A300) );
 a63777a <=( a63776a  and  a63773a );
 a63778a <=( a63777a  and  a63770a );
 a63782a <=( A167  and  A168 );
 a63783a <=( A170  and  a63782a );
 a63786a <=( A201  and  (not A166) );
 a63789a <=( A203  and  (not A202) );
 a63790a <=( a63789a  and  a63786a );
 a63791a <=( a63790a  and  a63783a );
 a63795a <=( (not A267)  and  A266 );
 a63796a <=( (not A265)  and  a63795a );
 a63799a <=( A269  and  (not A268) );
 a63802a <=( (not A302)  and  (not A300) );
 a63803a <=( a63802a  and  a63799a );
 a63804a <=( a63803a  and  a63796a );
 a63808a <=( A167  and  A168 );
 a63809a <=( A170  and  a63808a );
 a63812a <=( A201  and  (not A166) );
 a63815a <=( A203  and  (not A202) );
 a63816a <=( a63815a  and  a63812a );
 a63817a <=( a63816a  and  a63809a );
 a63821a <=( (not A267)  and  A266 );
 a63822a <=( (not A265)  and  a63821a );
 a63825a <=( A269  and  (not A268) );
 a63828a <=( A299  and  A298 );
 a63829a <=( a63828a  and  a63825a );
 a63830a <=( a63829a  and  a63822a );
 a63834a <=( A167  and  A168 );
 a63835a <=( A170  and  a63834a );
 a63838a <=( A201  and  (not A166) );
 a63841a <=( A203  and  (not A202) );
 a63842a <=( a63841a  and  a63838a );
 a63843a <=( a63842a  and  a63835a );
 a63847a <=( (not A267)  and  A266 );
 a63848a <=( (not A265)  and  a63847a );
 a63851a <=( A269  and  (not A268) );
 a63854a <=( (not A299)  and  (not A298) );
 a63855a <=( a63854a  and  a63851a );
 a63856a <=( a63855a  and  a63848a );
 a63860a <=( A167  and  A168 );
 a63861a <=( A170  and  a63860a );
 a63864a <=( A201  and  (not A166) );
 a63867a <=( A203  and  (not A202) );
 a63868a <=( a63867a  and  a63864a );
 a63869a <=( a63868a  and  a63861a );
 a63873a <=( A267  and  (not A266) );
 a63874a <=( A265  and  a63873a );
 a63877a <=( A300  and  A268 );
 a63880a <=( A302  and  (not A301) );
 a63881a <=( a63880a  and  a63877a );
 a63882a <=( a63881a  and  a63874a );
 a63886a <=( A167  and  A168 );
 a63887a <=( A170  and  a63886a );
 a63890a <=( A201  and  (not A166) );
 a63893a <=( A203  and  (not A202) );
 a63894a <=( a63893a  and  a63890a );
 a63895a <=( a63894a  and  a63887a );
 a63899a <=( A267  and  (not A266) );
 a63900a <=( A265  and  a63899a );
 a63903a <=( A300  and  (not A269) );
 a63906a <=( A302  and  (not A301) );
 a63907a <=( a63906a  and  a63903a );
 a63908a <=( a63907a  and  a63900a );
 a63912a <=( A167  and  A168 );
 a63913a <=( A170  and  a63912a );
 a63916a <=( A201  and  (not A166) );
 a63919a <=( A203  and  (not A202) );
 a63920a <=( a63919a  and  a63916a );
 a63921a <=( a63920a  and  a63913a );
 a63925a <=( (not A267)  and  (not A266) );
 a63926a <=( A265  and  a63925a );
 a63929a <=( A269  and  (not A268) );
 a63932a <=( A301  and  (not A300) );
 a63933a <=( a63932a  and  a63929a );
 a63934a <=( a63933a  and  a63926a );
 a63938a <=( A167  and  A168 );
 a63939a <=( A170  and  a63938a );
 a63942a <=( A201  and  (not A166) );
 a63945a <=( A203  and  (not A202) );
 a63946a <=( a63945a  and  a63942a );
 a63947a <=( a63946a  and  a63939a );
 a63951a <=( (not A267)  and  (not A266) );
 a63952a <=( A265  and  a63951a );
 a63955a <=( A269  and  (not A268) );
 a63958a <=( (not A302)  and  (not A300) );
 a63959a <=( a63958a  and  a63955a );
 a63960a <=( a63959a  and  a63952a );
 a63964a <=( A167  and  A168 );
 a63965a <=( A170  and  a63964a );
 a63968a <=( A201  and  (not A166) );
 a63971a <=( A203  and  (not A202) );
 a63972a <=( a63971a  and  a63968a );
 a63973a <=( a63972a  and  a63965a );
 a63977a <=( (not A267)  and  (not A266) );
 a63978a <=( A265  and  a63977a );
 a63981a <=( A269  and  (not A268) );
 a63984a <=( A299  and  A298 );
 a63985a <=( a63984a  and  a63981a );
 a63986a <=( a63985a  and  a63978a );
 a63990a <=( A167  and  A168 );
 a63991a <=( A170  and  a63990a );
 a63994a <=( A201  and  (not A166) );
 a63997a <=( A203  and  (not A202) );
 a63998a <=( a63997a  and  a63994a );
 a63999a <=( a63998a  and  a63991a );
 a64003a <=( (not A267)  and  (not A266) );
 a64004a <=( A265  and  a64003a );
 a64007a <=( A269  and  (not A268) );
 a64010a <=( (not A299)  and  (not A298) );
 a64011a <=( a64010a  and  a64007a );
 a64012a <=( a64011a  and  a64004a );
 a64016a <=( A167  and  A168 );
 a64017a <=( A170  and  a64016a );
 a64020a <=( A201  and  (not A166) );
 a64023a <=( A203  and  (not A202) );
 a64024a <=( a64023a  and  a64020a );
 a64025a <=( a64024a  and  a64017a );
 a64029a <=( A298  and  (not A266) );
 a64030a <=( (not A265)  and  a64029a );
 a64033a <=( (not A300)  and  (not A299) );
 a64036a <=( A302  and  (not A301) );
 a64037a <=( a64036a  and  a64033a );
 a64038a <=( a64037a  and  a64030a );
 a64042a <=( A167  and  A168 );
 a64043a <=( A170  and  a64042a );
 a64046a <=( A201  and  (not A166) );
 a64049a <=( A203  and  (not A202) );
 a64050a <=( a64049a  and  a64046a );
 a64051a <=( a64050a  and  a64043a );
 a64055a <=( (not A298)  and  (not A266) );
 a64056a <=( (not A265)  and  a64055a );
 a64059a <=( (not A300)  and  A299 );
 a64062a <=( A302  and  (not A301) );
 a64063a <=( a64062a  and  a64059a );
 a64064a <=( a64063a  and  a64056a );
 a64068a <=( A167  and  A168 );
 a64069a <=( A170  and  a64068a );
 a64072a <=( (not A201)  and  (not A166) );
 a64075a <=( A267  and  A202 );
 a64076a <=( a64075a  and  a64072a );
 a64077a <=( a64076a  and  a64069a );
 a64081a <=( A298  and  A269 );
 a64082a <=( (not A268)  and  a64081a );
 a64085a <=( (not A300)  and  (not A299) );
 a64088a <=( A302  and  (not A301) );
 a64089a <=( a64088a  and  a64085a );
 a64090a <=( a64089a  and  a64082a );
 a64094a <=( A167  and  A168 );
 a64095a <=( A170  and  a64094a );
 a64098a <=( (not A201)  and  (not A166) );
 a64101a <=( A267  and  A202 );
 a64102a <=( a64101a  and  a64098a );
 a64103a <=( a64102a  and  a64095a );
 a64107a <=( (not A298)  and  A269 );
 a64108a <=( (not A268)  and  a64107a );
 a64111a <=( (not A300)  and  A299 );
 a64114a <=( A302  and  (not A301) );
 a64115a <=( a64114a  and  a64111a );
 a64116a <=( a64115a  and  a64108a );
 a64120a <=( A167  and  A168 );
 a64121a <=( A170  and  a64120a );
 a64124a <=( (not A201)  and  (not A166) );
 a64127a <=( (not A265)  and  A202 );
 a64128a <=( a64127a  and  a64124a );
 a64129a <=( a64128a  and  a64121a );
 a64133a <=( (not A268)  and  (not A267) );
 a64134a <=( A266  and  a64133a );
 a64137a <=( A300  and  A269 );
 a64140a <=( A302  and  (not A301) );
 a64141a <=( a64140a  and  a64137a );
 a64142a <=( a64141a  and  a64134a );
 a64146a <=( A167  and  A168 );
 a64147a <=( A170  and  a64146a );
 a64150a <=( (not A201)  and  (not A166) );
 a64153a <=( A265  and  A202 );
 a64154a <=( a64153a  and  a64150a );
 a64155a <=( a64154a  and  a64147a );
 a64159a <=( (not A268)  and  (not A267) );
 a64160a <=( (not A266)  and  a64159a );
 a64163a <=( A300  and  A269 );
 a64166a <=( A302  and  (not A301) );
 a64167a <=( a64166a  and  a64163a );
 a64168a <=( a64167a  and  a64160a );
 a64172a <=( A167  and  A168 );
 a64173a <=( A170  and  a64172a );
 a64176a <=( (not A201)  and  (not A166) );
 a64179a <=( A267  and  (not A203) );
 a64180a <=( a64179a  and  a64176a );
 a64181a <=( a64180a  and  a64173a );
 a64185a <=( A298  and  A269 );
 a64186a <=( (not A268)  and  a64185a );
 a64189a <=( (not A300)  and  (not A299) );
 a64192a <=( A302  and  (not A301) );
 a64193a <=( a64192a  and  a64189a );
 a64194a <=( a64193a  and  a64186a );
 a64198a <=( A167  and  A168 );
 a64199a <=( A170  and  a64198a );
 a64202a <=( (not A201)  and  (not A166) );
 a64205a <=( A267  and  (not A203) );
 a64206a <=( a64205a  and  a64202a );
 a64207a <=( a64206a  and  a64199a );
 a64211a <=( (not A298)  and  A269 );
 a64212a <=( (not A268)  and  a64211a );
 a64215a <=( (not A300)  and  A299 );
 a64218a <=( A302  and  (not A301) );
 a64219a <=( a64218a  and  a64215a );
 a64220a <=( a64219a  and  a64212a );
 a64224a <=( A167  and  A168 );
 a64225a <=( A170  and  a64224a );
 a64228a <=( (not A201)  and  (not A166) );
 a64231a <=( (not A265)  and  (not A203) );
 a64232a <=( a64231a  and  a64228a );
 a64233a <=( a64232a  and  a64225a );
 a64237a <=( (not A268)  and  (not A267) );
 a64238a <=( A266  and  a64237a );
 a64241a <=( A300  and  A269 );
 a64244a <=( A302  and  (not A301) );
 a64245a <=( a64244a  and  a64241a );
 a64246a <=( a64245a  and  a64238a );
 a64250a <=( A167  and  A168 );
 a64251a <=( A170  and  a64250a );
 a64254a <=( (not A201)  and  (not A166) );
 a64257a <=( A265  and  (not A203) );
 a64258a <=( a64257a  and  a64254a );
 a64259a <=( a64258a  and  a64251a );
 a64263a <=( (not A268)  and  (not A267) );
 a64264a <=( (not A266)  and  a64263a );
 a64267a <=( A300  and  A269 );
 a64270a <=( A302  and  (not A301) );
 a64271a <=( a64270a  and  a64267a );
 a64272a <=( a64271a  and  a64264a );
 a64276a <=( A167  and  A168 );
 a64277a <=( A170  and  a64276a );
 a64280a <=( A199  and  (not A166) );
 a64283a <=( A267  and  A200 );
 a64284a <=( a64283a  and  a64280a );
 a64285a <=( a64284a  and  a64277a );
 a64289a <=( A298  and  A269 );
 a64290a <=( (not A268)  and  a64289a );
 a64293a <=( (not A300)  and  (not A299) );
 a64296a <=( A302  and  (not A301) );
 a64297a <=( a64296a  and  a64293a );
 a64298a <=( a64297a  and  a64290a );
 a64302a <=( A167  and  A168 );
 a64303a <=( A170  and  a64302a );
 a64306a <=( A199  and  (not A166) );
 a64309a <=( A267  and  A200 );
 a64310a <=( a64309a  and  a64306a );
 a64311a <=( a64310a  and  a64303a );
 a64315a <=( (not A298)  and  A269 );
 a64316a <=( (not A268)  and  a64315a );
 a64319a <=( (not A300)  and  A299 );
 a64322a <=( A302  and  (not A301) );
 a64323a <=( a64322a  and  a64319a );
 a64324a <=( a64323a  and  a64316a );
 a64328a <=( A167  and  A168 );
 a64329a <=( A170  and  a64328a );
 a64332a <=( A199  and  (not A166) );
 a64335a <=( (not A265)  and  A200 );
 a64336a <=( a64335a  and  a64332a );
 a64337a <=( a64336a  and  a64329a );
 a64341a <=( (not A268)  and  (not A267) );
 a64342a <=( A266  and  a64341a );
 a64345a <=( A300  and  A269 );
 a64348a <=( A302  and  (not A301) );
 a64349a <=( a64348a  and  a64345a );
 a64350a <=( a64349a  and  a64342a );
 a64354a <=( A167  and  A168 );
 a64355a <=( A170  and  a64354a );
 a64358a <=( A199  and  (not A166) );
 a64361a <=( A265  and  A200 );
 a64362a <=( a64361a  and  a64358a );
 a64363a <=( a64362a  and  a64355a );
 a64367a <=( (not A268)  and  (not A267) );
 a64368a <=( (not A266)  and  a64367a );
 a64371a <=( A300  and  A269 );
 a64374a <=( A302  and  (not A301) );
 a64375a <=( a64374a  and  a64371a );
 a64376a <=( a64375a  and  a64368a );
 a64380a <=( A167  and  A168 );
 a64381a <=( A170  and  a64380a );
 a64384a <=( (not A199)  and  (not A166) );
 a64387a <=( A267  and  (not A200) );
 a64388a <=( a64387a  and  a64384a );
 a64389a <=( a64388a  and  a64381a );
 a64393a <=( A298  and  A269 );
 a64394a <=( (not A268)  and  a64393a );
 a64397a <=( (not A300)  and  (not A299) );
 a64400a <=( A302  and  (not A301) );
 a64401a <=( a64400a  and  a64397a );
 a64402a <=( a64401a  and  a64394a );
 a64406a <=( A167  and  A168 );
 a64407a <=( A170  and  a64406a );
 a64410a <=( (not A199)  and  (not A166) );
 a64413a <=( A267  and  (not A200) );
 a64414a <=( a64413a  and  a64410a );
 a64415a <=( a64414a  and  a64407a );
 a64419a <=( (not A298)  and  A269 );
 a64420a <=( (not A268)  and  a64419a );
 a64423a <=( (not A300)  and  A299 );
 a64426a <=( A302  and  (not A301) );
 a64427a <=( a64426a  and  a64423a );
 a64428a <=( a64427a  and  a64420a );
 a64432a <=( A167  and  A168 );
 a64433a <=( A170  and  a64432a );
 a64436a <=( (not A199)  and  (not A166) );
 a64439a <=( (not A265)  and  (not A200) );
 a64440a <=( a64439a  and  a64436a );
 a64441a <=( a64440a  and  a64433a );
 a64445a <=( (not A268)  and  (not A267) );
 a64446a <=( A266  and  a64445a );
 a64449a <=( A300  and  A269 );
 a64452a <=( A302  and  (not A301) );
 a64453a <=( a64452a  and  a64449a );
 a64454a <=( a64453a  and  a64446a );
 a64458a <=( A167  and  A168 );
 a64459a <=( A170  and  a64458a );
 a64462a <=( (not A199)  and  (not A166) );
 a64465a <=( A265  and  (not A200) );
 a64466a <=( a64465a  and  a64462a );
 a64467a <=( a64466a  and  a64459a );
 a64471a <=( (not A268)  and  (not A267) );
 a64472a <=( (not A266)  and  a64471a );
 a64475a <=( A300  and  A269 );
 a64478a <=( A302  and  (not A301) );
 a64479a <=( a64478a  and  a64475a );
 a64480a <=( a64479a  and  a64472a );
 a64484a <=( (not A167)  and  A168 );
 a64485a <=( A170  and  a64484a );
 a64488a <=( A201  and  A166 );
 a64491a <=( A203  and  (not A202) );
 a64492a <=( a64491a  and  a64488a );
 a64493a <=( a64492a  and  a64485a );
 a64497a <=( A269  and  (not A268) );
 a64498a <=( A267  and  a64497a );
 a64501a <=( (not A299)  and  A298 );
 a64504a <=( A301  and  A300 );
 a64505a <=( a64504a  and  a64501a );
 a64506a <=( a64505a  and  a64498a );
 a64510a <=( (not A167)  and  A168 );
 a64511a <=( A170  and  a64510a );
 a64514a <=( A201  and  A166 );
 a64517a <=( A203  and  (not A202) );
 a64518a <=( a64517a  and  a64514a );
 a64519a <=( a64518a  and  a64511a );
 a64523a <=( A269  and  (not A268) );
 a64524a <=( A267  and  a64523a );
 a64527a <=( (not A299)  and  A298 );
 a64530a <=( (not A302)  and  A300 );
 a64531a <=( a64530a  and  a64527a );
 a64532a <=( a64531a  and  a64524a );
 a64536a <=( (not A167)  and  A168 );
 a64537a <=( A170  and  a64536a );
 a64540a <=( A201  and  A166 );
 a64543a <=( A203  and  (not A202) );
 a64544a <=( a64543a  and  a64540a );
 a64545a <=( a64544a  and  a64537a );
 a64549a <=( A269  and  (not A268) );
 a64550a <=( A267  and  a64549a );
 a64553a <=( A299  and  (not A298) );
 a64556a <=( A301  and  A300 );
 a64557a <=( a64556a  and  a64553a );
 a64558a <=( a64557a  and  a64550a );
 a64562a <=( (not A167)  and  A168 );
 a64563a <=( A170  and  a64562a );
 a64566a <=( A201  and  A166 );
 a64569a <=( A203  and  (not A202) );
 a64570a <=( a64569a  and  a64566a );
 a64571a <=( a64570a  and  a64563a );
 a64575a <=( A269  and  (not A268) );
 a64576a <=( A267  and  a64575a );
 a64579a <=( A299  and  (not A298) );
 a64582a <=( (not A302)  and  A300 );
 a64583a <=( a64582a  and  a64579a );
 a64584a <=( a64583a  and  a64576a );
 a64588a <=( (not A167)  and  A168 );
 a64589a <=( A170  and  a64588a );
 a64592a <=( A201  and  A166 );
 a64595a <=( A203  and  (not A202) );
 a64596a <=( a64595a  and  a64592a );
 a64597a <=( a64596a  and  a64589a );
 a64601a <=( A298  and  A268 );
 a64602a <=( (not A267)  and  a64601a );
 a64605a <=( (not A300)  and  (not A299) );
 a64608a <=( A302  and  (not A301) );
 a64609a <=( a64608a  and  a64605a );
 a64610a <=( a64609a  and  a64602a );
 a64614a <=( (not A167)  and  A168 );
 a64615a <=( A170  and  a64614a );
 a64618a <=( A201  and  A166 );
 a64621a <=( A203  and  (not A202) );
 a64622a <=( a64621a  and  a64618a );
 a64623a <=( a64622a  and  a64615a );
 a64627a <=( (not A298)  and  A268 );
 a64628a <=( (not A267)  and  a64627a );
 a64631a <=( (not A300)  and  A299 );
 a64634a <=( A302  and  (not A301) );
 a64635a <=( a64634a  and  a64631a );
 a64636a <=( a64635a  and  a64628a );
 a64640a <=( (not A167)  and  A168 );
 a64641a <=( A170  and  a64640a );
 a64644a <=( A201  and  A166 );
 a64647a <=( A203  and  (not A202) );
 a64648a <=( a64647a  and  a64644a );
 a64649a <=( a64648a  and  a64641a );
 a64653a <=( A298  and  (not A269) );
 a64654a <=( (not A267)  and  a64653a );
 a64657a <=( (not A300)  and  (not A299) );
 a64660a <=( A302  and  (not A301) );
 a64661a <=( a64660a  and  a64657a );
 a64662a <=( a64661a  and  a64654a );
 a64666a <=( (not A167)  and  A168 );
 a64667a <=( A170  and  a64666a );
 a64670a <=( A201  and  A166 );
 a64673a <=( A203  and  (not A202) );
 a64674a <=( a64673a  and  a64670a );
 a64675a <=( a64674a  and  a64667a );
 a64679a <=( (not A298)  and  (not A269) );
 a64680a <=( (not A267)  and  a64679a );
 a64683a <=( (not A300)  and  A299 );
 a64686a <=( A302  and  (not A301) );
 a64687a <=( a64686a  and  a64683a );
 a64688a <=( a64687a  and  a64680a );
 a64692a <=( (not A167)  and  A168 );
 a64693a <=( A170  and  a64692a );
 a64696a <=( A201  and  A166 );
 a64699a <=( A203  and  (not A202) );
 a64700a <=( a64699a  and  a64696a );
 a64701a <=( a64700a  and  a64693a );
 a64705a <=( A298  and  A266 );
 a64706a <=( A265  and  a64705a );
 a64709a <=( (not A300)  and  (not A299) );
 a64712a <=( A302  and  (not A301) );
 a64713a <=( a64712a  and  a64709a );
 a64714a <=( a64713a  and  a64706a );
 a64718a <=( (not A167)  and  A168 );
 a64719a <=( A170  and  a64718a );
 a64722a <=( A201  and  A166 );
 a64725a <=( A203  and  (not A202) );
 a64726a <=( a64725a  and  a64722a );
 a64727a <=( a64726a  and  a64719a );
 a64731a <=( (not A298)  and  A266 );
 a64732a <=( A265  and  a64731a );
 a64735a <=( (not A300)  and  A299 );
 a64738a <=( A302  and  (not A301) );
 a64739a <=( a64738a  and  a64735a );
 a64740a <=( a64739a  and  a64732a );
 a64744a <=( (not A167)  and  A168 );
 a64745a <=( A170  and  a64744a );
 a64748a <=( A201  and  A166 );
 a64751a <=( A203  and  (not A202) );
 a64752a <=( a64751a  and  a64748a );
 a64753a <=( a64752a  and  a64745a );
 a64757a <=( A267  and  A266 );
 a64758a <=( (not A265)  and  a64757a );
 a64761a <=( A300  and  A268 );
 a64764a <=( A302  and  (not A301) );
 a64765a <=( a64764a  and  a64761a );
 a64766a <=( a64765a  and  a64758a );
 a64770a <=( (not A167)  and  A168 );
 a64771a <=( A170  and  a64770a );
 a64774a <=( A201  and  A166 );
 a64777a <=( A203  and  (not A202) );
 a64778a <=( a64777a  and  a64774a );
 a64779a <=( a64778a  and  a64771a );
 a64783a <=( A267  and  A266 );
 a64784a <=( (not A265)  and  a64783a );
 a64787a <=( A300  and  (not A269) );
 a64790a <=( A302  and  (not A301) );
 a64791a <=( a64790a  and  a64787a );
 a64792a <=( a64791a  and  a64784a );
 a64796a <=( (not A167)  and  A168 );
 a64797a <=( A170  and  a64796a );
 a64800a <=( A201  and  A166 );
 a64803a <=( A203  and  (not A202) );
 a64804a <=( a64803a  and  a64800a );
 a64805a <=( a64804a  and  a64797a );
 a64809a <=( (not A267)  and  A266 );
 a64810a <=( (not A265)  and  a64809a );
 a64813a <=( A269  and  (not A268) );
 a64816a <=( A301  and  (not A300) );
 a64817a <=( a64816a  and  a64813a );
 a64818a <=( a64817a  and  a64810a );
 a64822a <=( (not A167)  and  A168 );
 a64823a <=( A170  and  a64822a );
 a64826a <=( A201  and  A166 );
 a64829a <=( A203  and  (not A202) );
 a64830a <=( a64829a  and  a64826a );
 a64831a <=( a64830a  and  a64823a );
 a64835a <=( (not A267)  and  A266 );
 a64836a <=( (not A265)  and  a64835a );
 a64839a <=( A269  and  (not A268) );
 a64842a <=( (not A302)  and  (not A300) );
 a64843a <=( a64842a  and  a64839a );
 a64844a <=( a64843a  and  a64836a );
 a64848a <=( (not A167)  and  A168 );
 a64849a <=( A170  and  a64848a );
 a64852a <=( A201  and  A166 );
 a64855a <=( A203  and  (not A202) );
 a64856a <=( a64855a  and  a64852a );
 a64857a <=( a64856a  and  a64849a );
 a64861a <=( (not A267)  and  A266 );
 a64862a <=( (not A265)  and  a64861a );
 a64865a <=( A269  and  (not A268) );
 a64868a <=( A299  and  A298 );
 a64869a <=( a64868a  and  a64865a );
 a64870a <=( a64869a  and  a64862a );
 a64874a <=( (not A167)  and  A168 );
 a64875a <=( A170  and  a64874a );
 a64878a <=( A201  and  A166 );
 a64881a <=( A203  and  (not A202) );
 a64882a <=( a64881a  and  a64878a );
 a64883a <=( a64882a  and  a64875a );
 a64887a <=( (not A267)  and  A266 );
 a64888a <=( (not A265)  and  a64887a );
 a64891a <=( A269  and  (not A268) );
 a64894a <=( (not A299)  and  (not A298) );
 a64895a <=( a64894a  and  a64891a );
 a64896a <=( a64895a  and  a64888a );
 a64900a <=( (not A167)  and  A168 );
 a64901a <=( A170  and  a64900a );
 a64904a <=( A201  and  A166 );
 a64907a <=( A203  and  (not A202) );
 a64908a <=( a64907a  and  a64904a );
 a64909a <=( a64908a  and  a64901a );
 a64913a <=( A267  and  (not A266) );
 a64914a <=( A265  and  a64913a );
 a64917a <=( A300  and  A268 );
 a64920a <=( A302  and  (not A301) );
 a64921a <=( a64920a  and  a64917a );
 a64922a <=( a64921a  and  a64914a );
 a64926a <=( (not A167)  and  A168 );
 a64927a <=( A170  and  a64926a );
 a64930a <=( A201  and  A166 );
 a64933a <=( A203  and  (not A202) );
 a64934a <=( a64933a  and  a64930a );
 a64935a <=( a64934a  and  a64927a );
 a64939a <=( A267  and  (not A266) );
 a64940a <=( A265  and  a64939a );
 a64943a <=( A300  and  (not A269) );
 a64946a <=( A302  and  (not A301) );
 a64947a <=( a64946a  and  a64943a );
 a64948a <=( a64947a  and  a64940a );
 a64952a <=( (not A167)  and  A168 );
 a64953a <=( A170  and  a64952a );
 a64956a <=( A201  and  A166 );
 a64959a <=( A203  and  (not A202) );
 a64960a <=( a64959a  and  a64956a );
 a64961a <=( a64960a  and  a64953a );
 a64965a <=( (not A267)  and  (not A266) );
 a64966a <=( A265  and  a64965a );
 a64969a <=( A269  and  (not A268) );
 a64972a <=( A301  and  (not A300) );
 a64973a <=( a64972a  and  a64969a );
 a64974a <=( a64973a  and  a64966a );
 a64978a <=( (not A167)  and  A168 );
 a64979a <=( A170  and  a64978a );
 a64982a <=( A201  and  A166 );
 a64985a <=( A203  and  (not A202) );
 a64986a <=( a64985a  and  a64982a );
 a64987a <=( a64986a  and  a64979a );
 a64991a <=( (not A267)  and  (not A266) );
 a64992a <=( A265  and  a64991a );
 a64995a <=( A269  and  (not A268) );
 a64998a <=( (not A302)  and  (not A300) );
 a64999a <=( a64998a  and  a64995a );
 a65000a <=( a64999a  and  a64992a );
 a65004a <=( (not A167)  and  A168 );
 a65005a <=( A170  and  a65004a );
 a65008a <=( A201  and  A166 );
 a65011a <=( A203  and  (not A202) );
 a65012a <=( a65011a  and  a65008a );
 a65013a <=( a65012a  and  a65005a );
 a65017a <=( (not A267)  and  (not A266) );
 a65018a <=( A265  and  a65017a );
 a65021a <=( A269  and  (not A268) );
 a65024a <=( A299  and  A298 );
 a65025a <=( a65024a  and  a65021a );
 a65026a <=( a65025a  and  a65018a );
 a65030a <=( (not A167)  and  A168 );
 a65031a <=( A170  and  a65030a );
 a65034a <=( A201  and  A166 );
 a65037a <=( A203  and  (not A202) );
 a65038a <=( a65037a  and  a65034a );
 a65039a <=( a65038a  and  a65031a );
 a65043a <=( (not A267)  and  (not A266) );
 a65044a <=( A265  and  a65043a );
 a65047a <=( A269  and  (not A268) );
 a65050a <=( (not A299)  and  (not A298) );
 a65051a <=( a65050a  and  a65047a );
 a65052a <=( a65051a  and  a65044a );
 a65056a <=( (not A167)  and  A168 );
 a65057a <=( A170  and  a65056a );
 a65060a <=( A201  and  A166 );
 a65063a <=( A203  and  (not A202) );
 a65064a <=( a65063a  and  a65060a );
 a65065a <=( a65064a  and  a65057a );
 a65069a <=( A298  and  (not A266) );
 a65070a <=( (not A265)  and  a65069a );
 a65073a <=( (not A300)  and  (not A299) );
 a65076a <=( A302  and  (not A301) );
 a65077a <=( a65076a  and  a65073a );
 a65078a <=( a65077a  and  a65070a );
 a65082a <=( (not A167)  and  A168 );
 a65083a <=( A170  and  a65082a );
 a65086a <=( A201  and  A166 );
 a65089a <=( A203  and  (not A202) );
 a65090a <=( a65089a  and  a65086a );
 a65091a <=( a65090a  and  a65083a );
 a65095a <=( (not A298)  and  (not A266) );
 a65096a <=( (not A265)  and  a65095a );
 a65099a <=( (not A300)  and  A299 );
 a65102a <=( A302  and  (not A301) );
 a65103a <=( a65102a  and  a65099a );
 a65104a <=( a65103a  and  a65096a );
 a65108a <=( (not A167)  and  A168 );
 a65109a <=( A170  and  a65108a );
 a65112a <=( (not A201)  and  A166 );
 a65115a <=( A267  and  A202 );
 a65116a <=( a65115a  and  a65112a );
 a65117a <=( a65116a  and  a65109a );
 a65121a <=( A298  and  A269 );
 a65122a <=( (not A268)  and  a65121a );
 a65125a <=( (not A300)  and  (not A299) );
 a65128a <=( A302  and  (not A301) );
 a65129a <=( a65128a  and  a65125a );
 a65130a <=( a65129a  and  a65122a );
 a65134a <=( (not A167)  and  A168 );
 a65135a <=( A170  and  a65134a );
 a65138a <=( (not A201)  and  A166 );
 a65141a <=( A267  and  A202 );
 a65142a <=( a65141a  and  a65138a );
 a65143a <=( a65142a  and  a65135a );
 a65147a <=( (not A298)  and  A269 );
 a65148a <=( (not A268)  and  a65147a );
 a65151a <=( (not A300)  and  A299 );
 a65154a <=( A302  and  (not A301) );
 a65155a <=( a65154a  and  a65151a );
 a65156a <=( a65155a  and  a65148a );
 a65160a <=( (not A167)  and  A168 );
 a65161a <=( A170  and  a65160a );
 a65164a <=( (not A201)  and  A166 );
 a65167a <=( (not A265)  and  A202 );
 a65168a <=( a65167a  and  a65164a );
 a65169a <=( a65168a  and  a65161a );
 a65173a <=( (not A268)  and  (not A267) );
 a65174a <=( A266  and  a65173a );
 a65177a <=( A300  and  A269 );
 a65180a <=( A302  and  (not A301) );
 a65181a <=( a65180a  and  a65177a );
 a65182a <=( a65181a  and  a65174a );
 a65186a <=( (not A167)  and  A168 );
 a65187a <=( A170  and  a65186a );
 a65190a <=( (not A201)  and  A166 );
 a65193a <=( A265  and  A202 );
 a65194a <=( a65193a  and  a65190a );
 a65195a <=( a65194a  and  a65187a );
 a65199a <=( (not A268)  and  (not A267) );
 a65200a <=( (not A266)  and  a65199a );
 a65203a <=( A300  and  A269 );
 a65206a <=( A302  and  (not A301) );
 a65207a <=( a65206a  and  a65203a );
 a65208a <=( a65207a  and  a65200a );
 a65212a <=( (not A167)  and  A168 );
 a65213a <=( A170  and  a65212a );
 a65216a <=( (not A201)  and  A166 );
 a65219a <=( A267  and  (not A203) );
 a65220a <=( a65219a  and  a65216a );
 a65221a <=( a65220a  and  a65213a );
 a65225a <=( A298  and  A269 );
 a65226a <=( (not A268)  and  a65225a );
 a65229a <=( (not A300)  and  (not A299) );
 a65232a <=( A302  and  (not A301) );
 a65233a <=( a65232a  and  a65229a );
 a65234a <=( a65233a  and  a65226a );
 a65238a <=( (not A167)  and  A168 );
 a65239a <=( A170  and  a65238a );
 a65242a <=( (not A201)  and  A166 );
 a65245a <=( A267  and  (not A203) );
 a65246a <=( a65245a  and  a65242a );
 a65247a <=( a65246a  and  a65239a );
 a65251a <=( (not A298)  and  A269 );
 a65252a <=( (not A268)  and  a65251a );
 a65255a <=( (not A300)  and  A299 );
 a65258a <=( A302  and  (not A301) );
 a65259a <=( a65258a  and  a65255a );
 a65260a <=( a65259a  and  a65252a );
 a65264a <=( (not A167)  and  A168 );
 a65265a <=( A170  and  a65264a );
 a65268a <=( (not A201)  and  A166 );
 a65271a <=( (not A265)  and  (not A203) );
 a65272a <=( a65271a  and  a65268a );
 a65273a <=( a65272a  and  a65265a );
 a65277a <=( (not A268)  and  (not A267) );
 a65278a <=( A266  and  a65277a );
 a65281a <=( A300  and  A269 );
 a65284a <=( A302  and  (not A301) );
 a65285a <=( a65284a  and  a65281a );
 a65286a <=( a65285a  and  a65278a );
 a65290a <=( (not A167)  and  A168 );
 a65291a <=( A170  and  a65290a );
 a65294a <=( (not A201)  and  A166 );
 a65297a <=( A265  and  (not A203) );
 a65298a <=( a65297a  and  a65294a );
 a65299a <=( a65298a  and  a65291a );
 a65303a <=( (not A268)  and  (not A267) );
 a65304a <=( (not A266)  and  a65303a );
 a65307a <=( A300  and  A269 );
 a65310a <=( A302  and  (not A301) );
 a65311a <=( a65310a  and  a65307a );
 a65312a <=( a65311a  and  a65304a );
 a65316a <=( (not A167)  and  A168 );
 a65317a <=( A170  and  a65316a );
 a65320a <=( A199  and  A166 );
 a65323a <=( A267  and  A200 );
 a65324a <=( a65323a  and  a65320a );
 a65325a <=( a65324a  and  a65317a );
 a65329a <=( A298  and  A269 );
 a65330a <=( (not A268)  and  a65329a );
 a65333a <=( (not A300)  and  (not A299) );
 a65336a <=( A302  and  (not A301) );
 a65337a <=( a65336a  and  a65333a );
 a65338a <=( a65337a  and  a65330a );
 a65342a <=( (not A167)  and  A168 );
 a65343a <=( A170  and  a65342a );
 a65346a <=( A199  and  A166 );
 a65349a <=( A267  and  A200 );
 a65350a <=( a65349a  and  a65346a );
 a65351a <=( a65350a  and  a65343a );
 a65355a <=( (not A298)  and  A269 );
 a65356a <=( (not A268)  and  a65355a );
 a65359a <=( (not A300)  and  A299 );
 a65362a <=( A302  and  (not A301) );
 a65363a <=( a65362a  and  a65359a );
 a65364a <=( a65363a  and  a65356a );
 a65368a <=( (not A167)  and  A168 );
 a65369a <=( A170  and  a65368a );
 a65372a <=( A199  and  A166 );
 a65375a <=( (not A265)  and  A200 );
 a65376a <=( a65375a  and  a65372a );
 a65377a <=( a65376a  and  a65369a );
 a65381a <=( (not A268)  and  (not A267) );
 a65382a <=( A266  and  a65381a );
 a65385a <=( A300  and  A269 );
 a65388a <=( A302  and  (not A301) );
 a65389a <=( a65388a  and  a65385a );
 a65390a <=( a65389a  and  a65382a );
 a65394a <=( (not A167)  and  A168 );
 a65395a <=( A170  and  a65394a );
 a65398a <=( A199  and  A166 );
 a65401a <=( A265  and  A200 );
 a65402a <=( a65401a  and  a65398a );
 a65403a <=( a65402a  and  a65395a );
 a65407a <=( (not A268)  and  (not A267) );
 a65408a <=( (not A266)  and  a65407a );
 a65411a <=( A300  and  A269 );
 a65414a <=( A302  and  (not A301) );
 a65415a <=( a65414a  and  a65411a );
 a65416a <=( a65415a  and  a65408a );
 a65420a <=( (not A167)  and  A168 );
 a65421a <=( A170  and  a65420a );
 a65424a <=( (not A199)  and  A166 );
 a65427a <=( A267  and  (not A200) );
 a65428a <=( a65427a  and  a65424a );
 a65429a <=( a65428a  and  a65421a );
 a65433a <=( A298  and  A269 );
 a65434a <=( (not A268)  and  a65433a );
 a65437a <=( (not A300)  and  (not A299) );
 a65440a <=( A302  and  (not A301) );
 a65441a <=( a65440a  and  a65437a );
 a65442a <=( a65441a  and  a65434a );
 a65446a <=( (not A167)  and  A168 );
 a65447a <=( A170  and  a65446a );
 a65450a <=( (not A199)  and  A166 );
 a65453a <=( A267  and  (not A200) );
 a65454a <=( a65453a  and  a65450a );
 a65455a <=( a65454a  and  a65447a );
 a65459a <=( (not A298)  and  A269 );
 a65460a <=( (not A268)  and  a65459a );
 a65463a <=( (not A300)  and  A299 );
 a65466a <=( A302  and  (not A301) );
 a65467a <=( a65466a  and  a65463a );
 a65468a <=( a65467a  and  a65460a );
 a65472a <=( (not A167)  and  A168 );
 a65473a <=( A170  and  a65472a );
 a65476a <=( (not A199)  and  A166 );
 a65479a <=( (not A265)  and  (not A200) );
 a65480a <=( a65479a  and  a65476a );
 a65481a <=( a65480a  and  a65473a );
 a65485a <=( (not A268)  and  (not A267) );
 a65486a <=( A266  and  a65485a );
 a65489a <=( A300  and  A269 );
 a65492a <=( A302  and  (not A301) );
 a65493a <=( a65492a  and  a65489a );
 a65494a <=( a65493a  and  a65486a );
 a65498a <=( (not A167)  and  A168 );
 a65499a <=( A170  and  a65498a );
 a65502a <=( (not A199)  and  A166 );
 a65505a <=( A265  and  (not A200) );
 a65506a <=( a65505a  and  a65502a );
 a65507a <=( a65506a  and  a65499a );
 a65511a <=( (not A268)  and  (not A267) );
 a65512a <=( (not A266)  and  a65511a );
 a65515a <=( A300  and  A269 );
 a65518a <=( A302  and  (not A301) );
 a65519a <=( a65518a  and  a65515a );
 a65520a <=( a65519a  and  a65512a );
 a65524a <=( (not A199)  and  (not A168) );
 a65525a <=( A170  and  a65524a );
 a65528a <=( A201  and  A200 );
 a65531a <=( (not A265)  and  A202 );
 a65532a <=( a65531a  and  a65528a );
 a65533a <=( a65532a  and  a65525a );
 a65537a <=( A268  and  A267 );
 a65538a <=( A266  and  a65537a );
 a65541a <=( (not A299)  and  A298 );
 a65544a <=( A301  and  A300 );
 a65545a <=( a65544a  and  a65541a );
 a65546a <=( a65545a  and  a65538a );
 a65550a <=( (not A199)  and  (not A168) );
 a65551a <=( A170  and  a65550a );
 a65554a <=( A201  and  A200 );
 a65557a <=( (not A265)  and  A202 );
 a65558a <=( a65557a  and  a65554a );
 a65559a <=( a65558a  and  a65551a );
 a65563a <=( A268  and  A267 );
 a65564a <=( A266  and  a65563a );
 a65567a <=( (not A299)  and  A298 );
 a65570a <=( (not A302)  and  A300 );
 a65571a <=( a65570a  and  a65567a );
 a65572a <=( a65571a  and  a65564a );
 a65576a <=( (not A199)  and  (not A168) );
 a65577a <=( A170  and  a65576a );
 a65580a <=( A201  and  A200 );
 a65583a <=( (not A265)  and  A202 );
 a65584a <=( a65583a  and  a65580a );
 a65585a <=( a65584a  and  a65577a );
 a65589a <=( A268  and  A267 );
 a65590a <=( A266  and  a65589a );
 a65593a <=( A299  and  (not A298) );
 a65596a <=( A301  and  A300 );
 a65597a <=( a65596a  and  a65593a );
 a65598a <=( a65597a  and  a65590a );
 a65602a <=( (not A199)  and  (not A168) );
 a65603a <=( A170  and  a65602a );
 a65606a <=( A201  and  A200 );
 a65609a <=( (not A265)  and  A202 );
 a65610a <=( a65609a  and  a65606a );
 a65611a <=( a65610a  and  a65603a );
 a65615a <=( A268  and  A267 );
 a65616a <=( A266  and  a65615a );
 a65619a <=( A299  and  (not A298) );
 a65622a <=( (not A302)  and  A300 );
 a65623a <=( a65622a  and  a65619a );
 a65624a <=( a65623a  and  a65616a );
 a65628a <=( (not A199)  and  (not A168) );
 a65629a <=( A170  and  a65628a );
 a65632a <=( A201  and  A200 );
 a65635a <=( (not A265)  and  A202 );
 a65636a <=( a65635a  and  a65632a );
 a65637a <=( a65636a  and  a65629a );
 a65641a <=( (not A269)  and  A267 );
 a65642a <=( A266  and  a65641a );
 a65645a <=( (not A299)  and  A298 );
 a65648a <=( A301  and  A300 );
 a65649a <=( a65648a  and  a65645a );
 a65650a <=( a65649a  and  a65642a );
 a65654a <=( (not A199)  and  (not A168) );
 a65655a <=( A170  and  a65654a );
 a65658a <=( A201  and  A200 );
 a65661a <=( (not A265)  and  A202 );
 a65662a <=( a65661a  and  a65658a );
 a65663a <=( a65662a  and  a65655a );
 a65667a <=( (not A269)  and  A267 );
 a65668a <=( A266  and  a65667a );
 a65671a <=( (not A299)  and  A298 );
 a65674a <=( (not A302)  and  A300 );
 a65675a <=( a65674a  and  a65671a );
 a65676a <=( a65675a  and  a65668a );
 a65680a <=( (not A199)  and  (not A168) );
 a65681a <=( A170  and  a65680a );
 a65684a <=( A201  and  A200 );
 a65687a <=( (not A265)  and  A202 );
 a65688a <=( a65687a  and  a65684a );
 a65689a <=( a65688a  and  a65681a );
 a65693a <=( (not A269)  and  A267 );
 a65694a <=( A266  and  a65693a );
 a65697a <=( A299  and  (not A298) );
 a65700a <=( A301  and  A300 );
 a65701a <=( a65700a  and  a65697a );
 a65702a <=( a65701a  and  a65694a );
 a65706a <=( (not A199)  and  (not A168) );
 a65707a <=( A170  and  a65706a );
 a65710a <=( A201  and  A200 );
 a65713a <=( (not A265)  and  A202 );
 a65714a <=( a65713a  and  a65710a );
 a65715a <=( a65714a  and  a65707a );
 a65719a <=( (not A269)  and  A267 );
 a65720a <=( A266  and  a65719a );
 a65723a <=( A299  and  (not A298) );
 a65726a <=( (not A302)  and  A300 );
 a65727a <=( a65726a  and  a65723a );
 a65728a <=( a65727a  and  a65720a );
 a65732a <=( (not A199)  and  (not A168) );
 a65733a <=( A170  and  a65732a );
 a65736a <=( A201  and  A200 );
 a65739a <=( A265  and  A202 );
 a65740a <=( a65739a  and  a65736a );
 a65741a <=( a65740a  and  a65733a );
 a65745a <=( A268  and  A267 );
 a65746a <=( (not A266)  and  a65745a );
 a65749a <=( (not A299)  and  A298 );
 a65752a <=( A301  and  A300 );
 a65753a <=( a65752a  and  a65749a );
 a65754a <=( a65753a  and  a65746a );
 a65758a <=( (not A199)  and  (not A168) );
 a65759a <=( A170  and  a65758a );
 a65762a <=( A201  and  A200 );
 a65765a <=( A265  and  A202 );
 a65766a <=( a65765a  and  a65762a );
 a65767a <=( a65766a  and  a65759a );
 a65771a <=( A268  and  A267 );
 a65772a <=( (not A266)  and  a65771a );
 a65775a <=( (not A299)  and  A298 );
 a65778a <=( (not A302)  and  A300 );
 a65779a <=( a65778a  and  a65775a );
 a65780a <=( a65779a  and  a65772a );
 a65784a <=( (not A199)  and  (not A168) );
 a65785a <=( A170  and  a65784a );
 a65788a <=( A201  and  A200 );
 a65791a <=( A265  and  A202 );
 a65792a <=( a65791a  and  a65788a );
 a65793a <=( a65792a  and  a65785a );
 a65797a <=( A268  and  A267 );
 a65798a <=( (not A266)  and  a65797a );
 a65801a <=( A299  and  (not A298) );
 a65804a <=( A301  and  A300 );
 a65805a <=( a65804a  and  a65801a );
 a65806a <=( a65805a  and  a65798a );
 a65810a <=( (not A199)  and  (not A168) );
 a65811a <=( A170  and  a65810a );
 a65814a <=( A201  and  A200 );
 a65817a <=( A265  and  A202 );
 a65818a <=( a65817a  and  a65814a );
 a65819a <=( a65818a  and  a65811a );
 a65823a <=( A268  and  A267 );
 a65824a <=( (not A266)  and  a65823a );
 a65827a <=( A299  and  (not A298) );
 a65830a <=( (not A302)  and  A300 );
 a65831a <=( a65830a  and  a65827a );
 a65832a <=( a65831a  and  a65824a );
 a65836a <=( (not A199)  and  (not A168) );
 a65837a <=( A170  and  a65836a );
 a65840a <=( A201  and  A200 );
 a65843a <=( A265  and  A202 );
 a65844a <=( a65843a  and  a65840a );
 a65845a <=( a65844a  and  a65837a );
 a65849a <=( (not A269)  and  A267 );
 a65850a <=( (not A266)  and  a65849a );
 a65853a <=( (not A299)  and  A298 );
 a65856a <=( A301  and  A300 );
 a65857a <=( a65856a  and  a65853a );
 a65858a <=( a65857a  and  a65850a );
 a65862a <=( (not A199)  and  (not A168) );
 a65863a <=( A170  and  a65862a );
 a65866a <=( A201  and  A200 );
 a65869a <=( A265  and  A202 );
 a65870a <=( a65869a  and  a65866a );
 a65871a <=( a65870a  and  a65863a );
 a65875a <=( (not A269)  and  A267 );
 a65876a <=( (not A266)  and  a65875a );
 a65879a <=( (not A299)  and  A298 );
 a65882a <=( (not A302)  and  A300 );
 a65883a <=( a65882a  and  a65879a );
 a65884a <=( a65883a  and  a65876a );
 a65888a <=( (not A199)  and  (not A168) );
 a65889a <=( A170  and  a65888a );
 a65892a <=( A201  and  A200 );
 a65895a <=( A265  and  A202 );
 a65896a <=( a65895a  and  a65892a );
 a65897a <=( a65896a  and  a65889a );
 a65901a <=( (not A269)  and  A267 );
 a65902a <=( (not A266)  and  a65901a );
 a65905a <=( A299  and  (not A298) );
 a65908a <=( A301  and  A300 );
 a65909a <=( a65908a  and  a65905a );
 a65910a <=( a65909a  and  a65902a );
 a65914a <=( (not A199)  and  (not A168) );
 a65915a <=( A170  and  a65914a );
 a65918a <=( A201  and  A200 );
 a65921a <=( A265  and  A202 );
 a65922a <=( a65921a  and  a65918a );
 a65923a <=( a65922a  and  a65915a );
 a65927a <=( (not A269)  and  A267 );
 a65928a <=( (not A266)  and  a65927a );
 a65931a <=( A299  and  (not A298) );
 a65934a <=( (not A302)  and  A300 );
 a65935a <=( a65934a  and  a65931a );
 a65936a <=( a65935a  and  a65928a );
 a65940a <=( (not A199)  and  (not A168) );
 a65941a <=( A170  and  a65940a );
 a65944a <=( A201  and  A200 );
 a65947a <=( (not A265)  and  (not A203) );
 a65948a <=( a65947a  and  a65944a );
 a65949a <=( a65948a  and  a65941a );
 a65953a <=( A268  and  A267 );
 a65954a <=( A266  and  a65953a );
 a65957a <=( (not A299)  and  A298 );
 a65960a <=( A301  and  A300 );
 a65961a <=( a65960a  and  a65957a );
 a65962a <=( a65961a  and  a65954a );
 a65966a <=( (not A199)  and  (not A168) );
 a65967a <=( A170  and  a65966a );
 a65970a <=( A201  and  A200 );
 a65973a <=( (not A265)  and  (not A203) );
 a65974a <=( a65973a  and  a65970a );
 a65975a <=( a65974a  and  a65967a );
 a65979a <=( A268  and  A267 );
 a65980a <=( A266  and  a65979a );
 a65983a <=( (not A299)  and  A298 );
 a65986a <=( (not A302)  and  A300 );
 a65987a <=( a65986a  and  a65983a );
 a65988a <=( a65987a  and  a65980a );
 a65992a <=( (not A199)  and  (not A168) );
 a65993a <=( A170  and  a65992a );
 a65996a <=( A201  and  A200 );
 a65999a <=( (not A265)  and  (not A203) );
 a66000a <=( a65999a  and  a65996a );
 a66001a <=( a66000a  and  a65993a );
 a66005a <=( A268  and  A267 );
 a66006a <=( A266  and  a66005a );
 a66009a <=( A299  and  (not A298) );
 a66012a <=( A301  and  A300 );
 a66013a <=( a66012a  and  a66009a );
 a66014a <=( a66013a  and  a66006a );
 a66018a <=( (not A199)  and  (not A168) );
 a66019a <=( A170  and  a66018a );
 a66022a <=( A201  and  A200 );
 a66025a <=( (not A265)  and  (not A203) );
 a66026a <=( a66025a  and  a66022a );
 a66027a <=( a66026a  and  a66019a );
 a66031a <=( A268  and  A267 );
 a66032a <=( A266  and  a66031a );
 a66035a <=( A299  and  (not A298) );
 a66038a <=( (not A302)  and  A300 );
 a66039a <=( a66038a  and  a66035a );
 a66040a <=( a66039a  and  a66032a );
 a66044a <=( (not A199)  and  (not A168) );
 a66045a <=( A170  and  a66044a );
 a66048a <=( A201  and  A200 );
 a66051a <=( (not A265)  and  (not A203) );
 a66052a <=( a66051a  and  a66048a );
 a66053a <=( a66052a  and  a66045a );
 a66057a <=( (not A269)  and  A267 );
 a66058a <=( A266  and  a66057a );
 a66061a <=( (not A299)  and  A298 );
 a66064a <=( A301  and  A300 );
 a66065a <=( a66064a  and  a66061a );
 a66066a <=( a66065a  and  a66058a );
 a66070a <=( (not A199)  and  (not A168) );
 a66071a <=( A170  and  a66070a );
 a66074a <=( A201  and  A200 );
 a66077a <=( (not A265)  and  (not A203) );
 a66078a <=( a66077a  and  a66074a );
 a66079a <=( a66078a  and  a66071a );
 a66083a <=( (not A269)  and  A267 );
 a66084a <=( A266  and  a66083a );
 a66087a <=( (not A299)  and  A298 );
 a66090a <=( (not A302)  and  A300 );
 a66091a <=( a66090a  and  a66087a );
 a66092a <=( a66091a  and  a66084a );
 a66096a <=( (not A199)  and  (not A168) );
 a66097a <=( A170  and  a66096a );
 a66100a <=( A201  and  A200 );
 a66103a <=( (not A265)  and  (not A203) );
 a66104a <=( a66103a  and  a66100a );
 a66105a <=( a66104a  and  a66097a );
 a66109a <=( (not A269)  and  A267 );
 a66110a <=( A266  and  a66109a );
 a66113a <=( A299  and  (not A298) );
 a66116a <=( A301  and  A300 );
 a66117a <=( a66116a  and  a66113a );
 a66118a <=( a66117a  and  a66110a );
 a66122a <=( (not A199)  and  (not A168) );
 a66123a <=( A170  and  a66122a );
 a66126a <=( A201  and  A200 );
 a66129a <=( (not A265)  and  (not A203) );
 a66130a <=( a66129a  and  a66126a );
 a66131a <=( a66130a  and  a66123a );
 a66135a <=( (not A269)  and  A267 );
 a66136a <=( A266  and  a66135a );
 a66139a <=( A299  and  (not A298) );
 a66142a <=( (not A302)  and  A300 );
 a66143a <=( a66142a  and  a66139a );
 a66144a <=( a66143a  and  a66136a );
 a66148a <=( (not A199)  and  (not A168) );
 a66149a <=( A170  and  a66148a );
 a66152a <=( A201  and  A200 );
 a66155a <=( A265  and  (not A203) );
 a66156a <=( a66155a  and  a66152a );
 a66157a <=( a66156a  and  a66149a );
 a66161a <=( A268  and  A267 );
 a66162a <=( (not A266)  and  a66161a );
 a66165a <=( (not A299)  and  A298 );
 a66168a <=( A301  and  A300 );
 a66169a <=( a66168a  and  a66165a );
 a66170a <=( a66169a  and  a66162a );
 a66174a <=( (not A199)  and  (not A168) );
 a66175a <=( A170  and  a66174a );
 a66178a <=( A201  and  A200 );
 a66181a <=( A265  and  (not A203) );
 a66182a <=( a66181a  and  a66178a );
 a66183a <=( a66182a  and  a66175a );
 a66187a <=( A268  and  A267 );
 a66188a <=( (not A266)  and  a66187a );
 a66191a <=( (not A299)  and  A298 );
 a66194a <=( (not A302)  and  A300 );
 a66195a <=( a66194a  and  a66191a );
 a66196a <=( a66195a  and  a66188a );
 a66200a <=( (not A199)  and  (not A168) );
 a66201a <=( A170  and  a66200a );
 a66204a <=( A201  and  A200 );
 a66207a <=( A265  and  (not A203) );
 a66208a <=( a66207a  and  a66204a );
 a66209a <=( a66208a  and  a66201a );
 a66213a <=( A268  and  A267 );
 a66214a <=( (not A266)  and  a66213a );
 a66217a <=( A299  and  (not A298) );
 a66220a <=( A301  and  A300 );
 a66221a <=( a66220a  and  a66217a );
 a66222a <=( a66221a  and  a66214a );
 a66226a <=( (not A199)  and  (not A168) );
 a66227a <=( A170  and  a66226a );
 a66230a <=( A201  and  A200 );
 a66233a <=( A265  and  (not A203) );
 a66234a <=( a66233a  and  a66230a );
 a66235a <=( a66234a  and  a66227a );
 a66239a <=( A268  and  A267 );
 a66240a <=( (not A266)  and  a66239a );
 a66243a <=( A299  and  (not A298) );
 a66246a <=( (not A302)  and  A300 );
 a66247a <=( a66246a  and  a66243a );
 a66248a <=( a66247a  and  a66240a );
 a66252a <=( (not A199)  and  (not A168) );
 a66253a <=( A170  and  a66252a );
 a66256a <=( A201  and  A200 );
 a66259a <=( A265  and  (not A203) );
 a66260a <=( a66259a  and  a66256a );
 a66261a <=( a66260a  and  a66253a );
 a66265a <=( (not A269)  and  A267 );
 a66266a <=( (not A266)  and  a66265a );
 a66269a <=( (not A299)  and  A298 );
 a66272a <=( A301  and  A300 );
 a66273a <=( a66272a  and  a66269a );
 a66274a <=( a66273a  and  a66266a );
 a66278a <=( (not A199)  and  (not A168) );
 a66279a <=( A170  and  a66278a );
 a66282a <=( A201  and  A200 );
 a66285a <=( A265  and  (not A203) );
 a66286a <=( a66285a  and  a66282a );
 a66287a <=( a66286a  and  a66279a );
 a66291a <=( (not A269)  and  A267 );
 a66292a <=( (not A266)  and  a66291a );
 a66295a <=( (not A299)  and  A298 );
 a66298a <=( (not A302)  and  A300 );
 a66299a <=( a66298a  and  a66295a );
 a66300a <=( a66299a  and  a66292a );
 a66304a <=( (not A199)  and  (not A168) );
 a66305a <=( A170  and  a66304a );
 a66308a <=( A201  and  A200 );
 a66311a <=( A265  and  (not A203) );
 a66312a <=( a66311a  and  a66308a );
 a66313a <=( a66312a  and  a66305a );
 a66317a <=( (not A269)  and  A267 );
 a66318a <=( (not A266)  and  a66317a );
 a66321a <=( A299  and  (not A298) );
 a66324a <=( A301  and  A300 );
 a66325a <=( a66324a  and  a66321a );
 a66326a <=( a66325a  and  a66318a );
 a66330a <=( (not A199)  and  (not A168) );
 a66331a <=( A170  and  a66330a );
 a66334a <=( A201  and  A200 );
 a66337a <=( A265  and  (not A203) );
 a66338a <=( a66337a  and  a66334a );
 a66339a <=( a66338a  and  a66331a );
 a66343a <=( (not A269)  and  A267 );
 a66344a <=( (not A266)  and  a66343a );
 a66347a <=( A299  and  (not A298) );
 a66350a <=( (not A302)  and  A300 );
 a66351a <=( a66350a  and  a66347a );
 a66352a <=( a66351a  and  a66344a );
 a66356a <=( A199  and  (not A168) );
 a66357a <=( A170  and  a66356a );
 a66360a <=( A201  and  (not A200) );
 a66363a <=( (not A265)  and  A202 );
 a66364a <=( a66363a  and  a66360a );
 a66365a <=( a66364a  and  a66357a );
 a66369a <=( A268  and  A267 );
 a66370a <=( A266  and  a66369a );
 a66373a <=( (not A299)  and  A298 );
 a66376a <=( A301  and  A300 );
 a66377a <=( a66376a  and  a66373a );
 a66378a <=( a66377a  and  a66370a );
 a66382a <=( A199  and  (not A168) );
 a66383a <=( A170  and  a66382a );
 a66386a <=( A201  and  (not A200) );
 a66389a <=( (not A265)  and  A202 );
 a66390a <=( a66389a  and  a66386a );
 a66391a <=( a66390a  and  a66383a );
 a66395a <=( A268  and  A267 );
 a66396a <=( A266  and  a66395a );
 a66399a <=( (not A299)  and  A298 );
 a66402a <=( (not A302)  and  A300 );
 a66403a <=( a66402a  and  a66399a );
 a66404a <=( a66403a  and  a66396a );
 a66408a <=( A199  and  (not A168) );
 a66409a <=( A170  and  a66408a );
 a66412a <=( A201  and  (not A200) );
 a66415a <=( (not A265)  and  A202 );
 a66416a <=( a66415a  and  a66412a );
 a66417a <=( a66416a  and  a66409a );
 a66421a <=( A268  and  A267 );
 a66422a <=( A266  and  a66421a );
 a66425a <=( A299  and  (not A298) );
 a66428a <=( A301  and  A300 );
 a66429a <=( a66428a  and  a66425a );
 a66430a <=( a66429a  and  a66422a );
 a66434a <=( A199  and  (not A168) );
 a66435a <=( A170  and  a66434a );
 a66438a <=( A201  and  (not A200) );
 a66441a <=( (not A265)  and  A202 );
 a66442a <=( a66441a  and  a66438a );
 a66443a <=( a66442a  and  a66435a );
 a66447a <=( A268  and  A267 );
 a66448a <=( A266  and  a66447a );
 a66451a <=( A299  and  (not A298) );
 a66454a <=( (not A302)  and  A300 );
 a66455a <=( a66454a  and  a66451a );
 a66456a <=( a66455a  and  a66448a );
 a66460a <=( A199  and  (not A168) );
 a66461a <=( A170  and  a66460a );
 a66464a <=( A201  and  (not A200) );
 a66467a <=( (not A265)  and  A202 );
 a66468a <=( a66467a  and  a66464a );
 a66469a <=( a66468a  and  a66461a );
 a66473a <=( (not A269)  and  A267 );
 a66474a <=( A266  and  a66473a );
 a66477a <=( (not A299)  and  A298 );
 a66480a <=( A301  and  A300 );
 a66481a <=( a66480a  and  a66477a );
 a66482a <=( a66481a  and  a66474a );
 a66486a <=( A199  and  (not A168) );
 a66487a <=( A170  and  a66486a );
 a66490a <=( A201  and  (not A200) );
 a66493a <=( (not A265)  and  A202 );
 a66494a <=( a66493a  and  a66490a );
 a66495a <=( a66494a  and  a66487a );
 a66499a <=( (not A269)  and  A267 );
 a66500a <=( A266  and  a66499a );
 a66503a <=( (not A299)  and  A298 );
 a66506a <=( (not A302)  and  A300 );
 a66507a <=( a66506a  and  a66503a );
 a66508a <=( a66507a  and  a66500a );
 a66512a <=( A199  and  (not A168) );
 a66513a <=( A170  and  a66512a );
 a66516a <=( A201  and  (not A200) );
 a66519a <=( (not A265)  and  A202 );
 a66520a <=( a66519a  and  a66516a );
 a66521a <=( a66520a  and  a66513a );
 a66525a <=( (not A269)  and  A267 );
 a66526a <=( A266  and  a66525a );
 a66529a <=( A299  and  (not A298) );
 a66532a <=( A301  and  A300 );
 a66533a <=( a66532a  and  a66529a );
 a66534a <=( a66533a  and  a66526a );
 a66538a <=( A199  and  (not A168) );
 a66539a <=( A170  and  a66538a );
 a66542a <=( A201  and  (not A200) );
 a66545a <=( (not A265)  and  A202 );
 a66546a <=( a66545a  and  a66542a );
 a66547a <=( a66546a  and  a66539a );
 a66551a <=( (not A269)  and  A267 );
 a66552a <=( A266  and  a66551a );
 a66555a <=( A299  and  (not A298) );
 a66558a <=( (not A302)  and  A300 );
 a66559a <=( a66558a  and  a66555a );
 a66560a <=( a66559a  and  a66552a );
 a66564a <=( A199  and  (not A168) );
 a66565a <=( A170  and  a66564a );
 a66568a <=( A201  and  (not A200) );
 a66571a <=( A265  and  A202 );
 a66572a <=( a66571a  and  a66568a );
 a66573a <=( a66572a  and  a66565a );
 a66577a <=( A268  and  A267 );
 a66578a <=( (not A266)  and  a66577a );
 a66581a <=( (not A299)  and  A298 );
 a66584a <=( A301  and  A300 );
 a66585a <=( a66584a  and  a66581a );
 a66586a <=( a66585a  and  a66578a );
 a66590a <=( A199  and  (not A168) );
 a66591a <=( A170  and  a66590a );
 a66594a <=( A201  and  (not A200) );
 a66597a <=( A265  and  A202 );
 a66598a <=( a66597a  and  a66594a );
 a66599a <=( a66598a  and  a66591a );
 a66603a <=( A268  and  A267 );
 a66604a <=( (not A266)  and  a66603a );
 a66607a <=( (not A299)  and  A298 );
 a66610a <=( (not A302)  and  A300 );
 a66611a <=( a66610a  and  a66607a );
 a66612a <=( a66611a  and  a66604a );
 a66616a <=( A199  and  (not A168) );
 a66617a <=( A170  and  a66616a );
 a66620a <=( A201  and  (not A200) );
 a66623a <=( A265  and  A202 );
 a66624a <=( a66623a  and  a66620a );
 a66625a <=( a66624a  and  a66617a );
 a66629a <=( A268  and  A267 );
 a66630a <=( (not A266)  and  a66629a );
 a66633a <=( A299  and  (not A298) );
 a66636a <=( A301  and  A300 );
 a66637a <=( a66636a  and  a66633a );
 a66638a <=( a66637a  and  a66630a );
 a66642a <=( A199  and  (not A168) );
 a66643a <=( A170  and  a66642a );
 a66646a <=( A201  and  (not A200) );
 a66649a <=( A265  and  A202 );
 a66650a <=( a66649a  and  a66646a );
 a66651a <=( a66650a  and  a66643a );
 a66655a <=( A268  and  A267 );
 a66656a <=( (not A266)  and  a66655a );
 a66659a <=( A299  and  (not A298) );
 a66662a <=( (not A302)  and  A300 );
 a66663a <=( a66662a  and  a66659a );
 a66664a <=( a66663a  and  a66656a );
 a66668a <=( A199  and  (not A168) );
 a66669a <=( A170  and  a66668a );
 a66672a <=( A201  and  (not A200) );
 a66675a <=( A265  and  A202 );
 a66676a <=( a66675a  and  a66672a );
 a66677a <=( a66676a  and  a66669a );
 a66681a <=( (not A269)  and  A267 );
 a66682a <=( (not A266)  and  a66681a );
 a66685a <=( (not A299)  and  A298 );
 a66688a <=( A301  and  A300 );
 a66689a <=( a66688a  and  a66685a );
 a66690a <=( a66689a  and  a66682a );
 a66694a <=( A199  and  (not A168) );
 a66695a <=( A170  and  a66694a );
 a66698a <=( A201  and  (not A200) );
 a66701a <=( A265  and  A202 );
 a66702a <=( a66701a  and  a66698a );
 a66703a <=( a66702a  and  a66695a );
 a66707a <=( (not A269)  and  A267 );
 a66708a <=( (not A266)  and  a66707a );
 a66711a <=( (not A299)  and  A298 );
 a66714a <=( (not A302)  and  A300 );
 a66715a <=( a66714a  and  a66711a );
 a66716a <=( a66715a  and  a66708a );
 a66720a <=( A199  and  (not A168) );
 a66721a <=( A170  and  a66720a );
 a66724a <=( A201  and  (not A200) );
 a66727a <=( A265  and  A202 );
 a66728a <=( a66727a  and  a66724a );
 a66729a <=( a66728a  and  a66721a );
 a66733a <=( (not A269)  and  A267 );
 a66734a <=( (not A266)  and  a66733a );
 a66737a <=( A299  and  (not A298) );
 a66740a <=( A301  and  A300 );
 a66741a <=( a66740a  and  a66737a );
 a66742a <=( a66741a  and  a66734a );
 a66746a <=( A199  and  (not A168) );
 a66747a <=( A170  and  a66746a );
 a66750a <=( A201  and  (not A200) );
 a66753a <=( A265  and  A202 );
 a66754a <=( a66753a  and  a66750a );
 a66755a <=( a66754a  and  a66747a );
 a66759a <=( (not A269)  and  A267 );
 a66760a <=( (not A266)  and  a66759a );
 a66763a <=( A299  and  (not A298) );
 a66766a <=( (not A302)  and  A300 );
 a66767a <=( a66766a  and  a66763a );
 a66768a <=( a66767a  and  a66760a );
 a66772a <=( A199  and  (not A168) );
 a66773a <=( A170  and  a66772a );
 a66776a <=( A201  and  (not A200) );
 a66779a <=( (not A265)  and  (not A203) );
 a66780a <=( a66779a  and  a66776a );
 a66781a <=( a66780a  and  a66773a );
 a66785a <=( A268  and  A267 );
 a66786a <=( A266  and  a66785a );
 a66789a <=( (not A299)  and  A298 );
 a66792a <=( A301  and  A300 );
 a66793a <=( a66792a  and  a66789a );
 a66794a <=( a66793a  and  a66786a );
 a66798a <=( A199  and  (not A168) );
 a66799a <=( A170  and  a66798a );
 a66802a <=( A201  and  (not A200) );
 a66805a <=( (not A265)  and  (not A203) );
 a66806a <=( a66805a  and  a66802a );
 a66807a <=( a66806a  and  a66799a );
 a66811a <=( A268  and  A267 );
 a66812a <=( A266  and  a66811a );
 a66815a <=( (not A299)  and  A298 );
 a66818a <=( (not A302)  and  A300 );
 a66819a <=( a66818a  and  a66815a );
 a66820a <=( a66819a  and  a66812a );
 a66824a <=( A199  and  (not A168) );
 a66825a <=( A170  and  a66824a );
 a66828a <=( A201  and  (not A200) );
 a66831a <=( (not A265)  and  (not A203) );
 a66832a <=( a66831a  and  a66828a );
 a66833a <=( a66832a  and  a66825a );
 a66837a <=( A268  and  A267 );
 a66838a <=( A266  and  a66837a );
 a66841a <=( A299  and  (not A298) );
 a66844a <=( A301  and  A300 );
 a66845a <=( a66844a  and  a66841a );
 a66846a <=( a66845a  and  a66838a );
 a66850a <=( A199  and  (not A168) );
 a66851a <=( A170  and  a66850a );
 a66854a <=( A201  and  (not A200) );
 a66857a <=( (not A265)  and  (not A203) );
 a66858a <=( a66857a  and  a66854a );
 a66859a <=( a66858a  and  a66851a );
 a66863a <=( A268  and  A267 );
 a66864a <=( A266  and  a66863a );
 a66867a <=( A299  and  (not A298) );
 a66870a <=( (not A302)  and  A300 );
 a66871a <=( a66870a  and  a66867a );
 a66872a <=( a66871a  and  a66864a );
 a66876a <=( A199  and  (not A168) );
 a66877a <=( A170  and  a66876a );
 a66880a <=( A201  and  (not A200) );
 a66883a <=( (not A265)  and  (not A203) );
 a66884a <=( a66883a  and  a66880a );
 a66885a <=( a66884a  and  a66877a );
 a66889a <=( (not A269)  and  A267 );
 a66890a <=( A266  and  a66889a );
 a66893a <=( (not A299)  and  A298 );
 a66896a <=( A301  and  A300 );
 a66897a <=( a66896a  and  a66893a );
 a66898a <=( a66897a  and  a66890a );
 a66902a <=( A199  and  (not A168) );
 a66903a <=( A170  and  a66902a );
 a66906a <=( A201  and  (not A200) );
 a66909a <=( (not A265)  and  (not A203) );
 a66910a <=( a66909a  and  a66906a );
 a66911a <=( a66910a  and  a66903a );
 a66915a <=( (not A269)  and  A267 );
 a66916a <=( A266  and  a66915a );
 a66919a <=( (not A299)  and  A298 );
 a66922a <=( (not A302)  and  A300 );
 a66923a <=( a66922a  and  a66919a );
 a66924a <=( a66923a  and  a66916a );
 a66928a <=( A199  and  (not A168) );
 a66929a <=( A170  and  a66928a );
 a66932a <=( A201  and  (not A200) );
 a66935a <=( (not A265)  and  (not A203) );
 a66936a <=( a66935a  and  a66932a );
 a66937a <=( a66936a  and  a66929a );
 a66941a <=( (not A269)  and  A267 );
 a66942a <=( A266  and  a66941a );
 a66945a <=( A299  and  (not A298) );
 a66948a <=( A301  and  A300 );
 a66949a <=( a66948a  and  a66945a );
 a66950a <=( a66949a  and  a66942a );
 a66954a <=( A199  and  (not A168) );
 a66955a <=( A170  and  a66954a );
 a66958a <=( A201  and  (not A200) );
 a66961a <=( (not A265)  and  (not A203) );
 a66962a <=( a66961a  and  a66958a );
 a66963a <=( a66962a  and  a66955a );
 a66967a <=( (not A269)  and  A267 );
 a66968a <=( A266  and  a66967a );
 a66971a <=( A299  and  (not A298) );
 a66974a <=( (not A302)  and  A300 );
 a66975a <=( a66974a  and  a66971a );
 a66976a <=( a66975a  and  a66968a );
 a66980a <=( A199  and  (not A168) );
 a66981a <=( A170  and  a66980a );
 a66984a <=( A201  and  (not A200) );
 a66987a <=( A265  and  (not A203) );
 a66988a <=( a66987a  and  a66984a );
 a66989a <=( a66988a  and  a66981a );
 a66993a <=( A268  and  A267 );
 a66994a <=( (not A266)  and  a66993a );
 a66997a <=( (not A299)  and  A298 );
 a67000a <=( A301  and  A300 );
 a67001a <=( a67000a  and  a66997a );
 a67002a <=( a67001a  and  a66994a );
 a67006a <=( A199  and  (not A168) );
 a67007a <=( A170  and  a67006a );
 a67010a <=( A201  and  (not A200) );
 a67013a <=( A265  and  (not A203) );
 a67014a <=( a67013a  and  a67010a );
 a67015a <=( a67014a  and  a67007a );
 a67019a <=( A268  and  A267 );
 a67020a <=( (not A266)  and  a67019a );
 a67023a <=( (not A299)  and  A298 );
 a67026a <=( (not A302)  and  A300 );
 a67027a <=( a67026a  and  a67023a );
 a67028a <=( a67027a  and  a67020a );
 a67032a <=( A199  and  (not A168) );
 a67033a <=( A170  and  a67032a );
 a67036a <=( A201  and  (not A200) );
 a67039a <=( A265  and  (not A203) );
 a67040a <=( a67039a  and  a67036a );
 a67041a <=( a67040a  and  a67033a );
 a67045a <=( A268  and  A267 );
 a67046a <=( (not A266)  and  a67045a );
 a67049a <=( A299  and  (not A298) );
 a67052a <=( A301  and  A300 );
 a67053a <=( a67052a  and  a67049a );
 a67054a <=( a67053a  and  a67046a );
 a67058a <=( A199  and  (not A168) );
 a67059a <=( A170  and  a67058a );
 a67062a <=( A201  and  (not A200) );
 a67065a <=( A265  and  (not A203) );
 a67066a <=( a67065a  and  a67062a );
 a67067a <=( a67066a  and  a67059a );
 a67071a <=( A268  and  A267 );
 a67072a <=( (not A266)  and  a67071a );
 a67075a <=( A299  and  (not A298) );
 a67078a <=( (not A302)  and  A300 );
 a67079a <=( a67078a  and  a67075a );
 a67080a <=( a67079a  and  a67072a );
 a67084a <=( A199  and  (not A168) );
 a67085a <=( A170  and  a67084a );
 a67088a <=( A201  and  (not A200) );
 a67091a <=( A265  and  (not A203) );
 a67092a <=( a67091a  and  a67088a );
 a67093a <=( a67092a  and  a67085a );
 a67097a <=( (not A269)  and  A267 );
 a67098a <=( (not A266)  and  a67097a );
 a67101a <=( (not A299)  and  A298 );
 a67104a <=( A301  and  A300 );
 a67105a <=( a67104a  and  a67101a );
 a67106a <=( a67105a  and  a67098a );
 a67110a <=( A199  and  (not A168) );
 a67111a <=( A170  and  a67110a );
 a67114a <=( A201  and  (not A200) );
 a67117a <=( A265  and  (not A203) );
 a67118a <=( a67117a  and  a67114a );
 a67119a <=( a67118a  and  a67111a );
 a67123a <=( (not A269)  and  A267 );
 a67124a <=( (not A266)  and  a67123a );
 a67127a <=( (not A299)  and  A298 );
 a67130a <=( (not A302)  and  A300 );
 a67131a <=( a67130a  and  a67127a );
 a67132a <=( a67131a  and  a67124a );
 a67136a <=( A199  and  (not A168) );
 a67137a <=( A170  and  a67136a );
 a67140a <=( A201  and  (not A200) );
 a67143a <=( A265  and  (not A203) );
 a67144a <=( a67143a  and  a67140a );
 a67145a <=( a67144a  and  a67137a );
 a67149a <=( (not A269)  and  A267 );
 a67150a <=( (not A266)  and  a67149a );
 a67153a <=( A299  and  (not A298) );
 a67156a <=( A301  and  A300 );
 a67157a <=( a67156a  and  a67153a );
 a67158a <=( a67157a  and  a67150a );
 a67162a <=( A199  and  (not A168) );
 a67163a <=( A170  and  a67162a );
 a67166a <=( A201  and  (not A200) );
 a67169a <=( A265  and  (not A203) );
 a67170a <=( a67169a  and  a67166a );
 a67171a <=( a67170a  and  a67163a );
 a67175a <=( (not A269)  and  A267 );
 a67176a <=( (not A266)  and  a67175a );
 a67179a <=( A299  and  (not A298) );
 a67182a <=( (not A302)  and  A300 );
 a67183a <=( a67182a  and  a67179a );
 a67184a <=( a67183a  and  a67176a );
 a67188a <=( A167  and  A168 );
 a67189a <=( A169  and  a67188a );
 a67192a <=( A201  and  (not A166) );
 a67195a <=( A203  and  (not A202) );
 a67196a <=( a67195a  and  a67192a );
 a67197a <=( a67196a  and  a67189a );
 a67201a <=( A269  and  (not A268) );
 a67202a <=( A267  and  a67201a );
 a67205a <=( (not A299)  and  A298 );
 a67208a <=( A301  and  A300 );
 a67209a <=( a67208a  and  a67205a );
 a67210a <=( a67209a  and  a67202a );
 a67214a <=( A167  and  A168 );
 a67215a <=( A169  and  a67214a );
 a67218a <=( A201  and  (not A166) );
 a67221a <=( A203  and  (not A202) );
 a67222a <=( a67221a  and  a67218a );
 a67223a <=( a67222a  and  a67215a );
 a67227a <=( A269  and  (not A268) );
 a67228a <=( A267  and  a67227a );
 a67231a <=( (not A299)  and  A298 );
 a67234a <=( (not A302)  and  A300 );
 a67235a <=( a67234a  and  a67231a );
 a67236a <=( a67235a  and  a67228a );
 a67240a <=( A167  and  A168 );
 a67241a <=( A169  and  a67240a );
 a67244a <=( A201  and  (not A166) );
 a67247a <=( A203  and  (not A202) );
 a67248a <=( a67247a  and  a67244a );
 a67249a <=( a67248a  and  a67241a );
 a67253a <=( A269  and  (not A268) );
 a67254a <=( A267  and  a67253a );
 a67257a <=( A299  and  (not A298) );
 a67260a <=( A301  and  A300 );
 a67261a <=( a67260a  and  a67257a );
 a67262a <=( a67261a  and  a67254a );
 a67266a <=( A167  and  A168 );
 a67267a <=( A169  and  a67266a );
 a67270a <=( A201  and  (not A166) );
 a67273a <=( A203  and  (not A202) );
 a67274a <=( a67273a  and  a67270a );
 a67275a <=( a67274a  and  a67267a );
 a67279a <=( A269  and  (not A268) );
 a67280a <=( A267  and  a67279a );
 a67283a <=( A299  and  (not A298) );
 a67286a <=( (not A302)  and  A300 );
 a67287a <=( a67286a  and  a67283a );
 a67288a <=( a67287a  and  a67280a );
 a67292a <=( A167  and  A168 );
 a67293a <=( A169  and  a67292a );
 a67296a <=( A201  and  (not A166) );
 a67299a <=( A203  and  (not A202) );
 a67300a <=( a67299a  and  a67296a );
 a67301a <=( a67300a  and  a67293a );
 a67305a <=( A298  and  A268 );
 a67306a <=( (not A267)  and  a67305a );
 a67309a <=( (not A300)  and  (not A299) );
 a67312a <=( A302  and  (not A301) );
 a67313a <=( a67312a  and  a67309a );
 a67314a <=( a67313a  and  a67306a );
 a67318a <=( A167  and  A168 );
 a67319a <=( A169  and  a67318a );
 a67322a <=( A201  and  (not A166) );
 a67325a <=( A203  and  (not A202) );
 a67326a <=( a67325a  and  a67322a );
 a67327a <=( a67326a  and  a67319a );
 a67331a <=( (not A298)  and  A268 );
 a67332a <=( (not A267)  and  a67331a );
 a67335a <=( (not A300)  and  A299 );
 a67338a <=( A302  and  (not A301) );
 a67339a <=( a67338a  and  a67335a );
 a67340a <=( a67339a  and  a67332a );
 a67344a <=( A167  and  A168 );
 a67345a <=( A169  and  a67344a );
 a67348a <=( A201  and  (not A166) );
 a67351a <=( A203  and  (not A202) );
 a67352a <=( a67351a  and  a67348a );
 a67353a <=( a67352a  and  a67345a );
 a67357a <=( A298  and  (not A269) );
 a67358a <=( (not A267)  and  a67357a );
 a67361a <=( (not A300)  and  (not A299) );
 a67364a <=( A302  and  (not A301) );
 a67365a <=( a67364a  and  a67361a );
 a67366a <=( a67365a  and  a67358a );
 a67370a <=( A167  and  A168 );
 a67371a <=( A169  and  a67370a );
 a67374a <=( A201  and  (not A166) );
 a67377a <=( A203  and  (not A202) );
 a67378a <=( a67377a  and  a67374a );
 a67379a <=( a67378a  and  a67371a );
 a67383a <=( (not A298)  and  (not A269) );
 a67384a <=( (not A267)  and  a67383a );
 a67387a <=( (not A300)  and  A299 );
 a67390a <=( A302  and  (not A301) );
 a67391a <=( a67390a  and  a67387a );
 a67392a <=( a67391a  and  a67384a );
 a67396a <=( A167  and  A168 );
 a67397a <=( A169  and  a67396a );
 a67400a <=( A201  and  (not A166) );
 a67403a <=( A203  and  (not A202) );
 a67404a <=( a67403a  and  a67400a );
 a67405a <=( a67404a  and  a67397a );
 a67409a <=( A298  and  A266 );
 a67410a <=( A265  and  a67409a );
 a67413a <=( (not A300)  and  (not A299) );
 a67416a <=( A302  and  (not A301) );
 a67417a <=( a67416a  and  a67413a );
 a67418a <=( a67417a  and  a67410a );
 a67422a <=( A167  and  A168 );
 a67423a <=( A169  and  a67422a );
 a67426a <=( A201  and  (not A166) );
 a67429a <=( A203  and  (not A202) );
 a67430a <=( a67429a  and  a67426a );
 a67431a <=( a67430a  and  a67423a );
 a67435a <=( (not A298)  and  A266 );
 a67436a <=( A265  and  a67435a );
 a67439a <=( (not A300)  and  A299 );
 a67442a <=( A302  and  (not A301) );
 a67443a <=( a67442a  and  a67439a );
 a67444a <=( a67443a  and  a67436a );
 a67448a <=( A167  and  A168 );
 a67449a <=( A169  and  a67448a );
 a67452a <=( A201  and  (not A166) );
 a67455a <=( A203  and  (not A202) );
 a67456a <=( a67455a  and  a67452a );
 a67457a <=( a67456a  and  a67449a );
 a67461a <=( A267  and  A266 );
 a67462a <=( (not A265)  and  a67461a );
 a67465a <=( A300  and  A268 );
 a67468a <=( A302  and  (not A301) );
 a67469a <=( a67468a  and  a67465a );
 a67470a <=( a67469a  and  a67462a );
 a67474a <=( A167  and  A168 );
 a67475a <=( A169  and  a67474a );
 a67478a <=( A201  and  (not A166) );
 a67481a <=( A203  and  (not A202) );
 a67482a <=( a67481a  and  a67478a );
 a67483a <=( a67482a  and  a67475a );
 a67487a <=( A267  and  A266 );
 a67488a <=( (not A265)  and  a67487a );
 a67491a <=( A300  and  (not A269) );
 a67494a <=( A302  and  (not A301) );
 a67495a <=( a67494a  and  a67491a );
 a67496a <=( a67495a  and  a67488a );
 a67500a <=( A167  and  A168 );
 a67501a <=( A169  and  a67500a );
 a67504a <=( A201  and  (not A166) );
 a67507a <=( A203  and  (not A202) );
 a67508a <=( a67507a  and  a67504a );
 a67509a <=( a67508a  and  a67501a );
 a67513a <=( (not A267)  and  A266 );
 a67514a <=( (not A265)  and  a67513a );
 a67517a <=( A269  and  (not A268) );
 a67520a <=( A301  and  (not A300) );
 a67521a <=( a67520a  and  a67517a );
 a67522a <=( a67521a  and  a67514a );
 a67526a <=( A167  and  A168 );
 a67527a <=( A169  and  a67526a );
 a67530a <=( A201  and  (not A166) );
 a67533a <=( A203  and  (not A202) );
 a67534a <=( a67533a  and  a67530a );
 a67535a <=( a67534a  and  a67527a );
 a67539a <=( (not A267)  and  A266 );
 a67540a <=( (not A265)  and  a67539a );
 a67543a <=( A269  and  (not A268) );
 a67546a <=( (not A302)  and  (not A300) );
 a67547a <=( a67546a  and  a67543a );
 a67548a <=( a67547a  and  a67540a );
 a67552a <=( A167  and  A168 );
 a67553a <=( A169  and  a67552a );
 a67556a <=( A201  and  (not A166) );
 a67559a <=( A203  and  (not A202) );
 a67560a <=( a67559a  and  a67556a );
 a67561a <=( a67560a  and  a67553a );
 a67565a <=( (not A267)  and  A266 );
 a67566a <=( (not A265)  and  a67565a );
 a67569a <=( A269  and  (not A268) );
 a67572a <=( A299  and  A298 );
 a67573a <=( a67572a  and  a67569a );
 a67574a <=( a67573a  and  a67566a );
 a67578a <=( A167  and  A168 );
 a67579a <=( A169  and  a67578a );
 a67582a <=( A201  and  (not A166) );
 a67585a <=( A203  and  (not A202) );
 a67586a <=( a67585a  and  a67582a );
 a67587a <=( a67586a  and  a67579a );
 a67591a <=( (not A267)  and  A266 );
 a67592a <=( (not A265)  and  a67591a );
 a67595a <=( A269  and  (not A268) );
 a67598a <=( (not A299)  and  (not A298) );
 a67599a <=( a67598a  and  a67595a );
 a67600a <=( a67599a  and  a67592a );
 a67604a <=( A167  and  A168 );
 a67605a <=( A169  and  a67604a );
 a67608a <=( A201  and  (not A166) );
 a67611a <=( A203  and  (not A202) );
 a67612a <=( a67611a  and  a67608a );
 a67613a <=( a67612a  and  a67605a );
 a67617a <=( A267  and  (not A266) );
 a67618a <=( A265  and  a67617a );
 a67621a <=( A300  and  A268 );
 a67624a <=( A302  and  (not A301) );
 a67625a <=( a67624a  and  a67621a );
 a67626a <=( a67625a  and  a67618a );
 a67630a <=( A167  and  A168 );
 a67631a <=( A169  and  a67630a );
 a67634a <=( A201  and  (not A166) );
 a67637a <=( A203  and  (not A202) );
 a67638a <=( a67637a  and  a67634a );
 a67639a <=( a67638a  and  a67631a );
 a67643a <=( A267  and  (not A266) );
 a67644a <=( A265  and  a67643a );
 a67647a <=( A300  and  (not A269) );
 a67650a <=( A302  and  (not A301) );
 a67651a <=( a67650a  and  a67647a );
 a67652a <=( a67651a  and  a67644a );
 a67656a <=( A167  and  A168 );
 a67657a <=( A169  and  a67656a );
 a67660a <=( A201  and  (not A166) );
 a67663a <=( A203  and  (not A202) );
 a67664a <=( a67663a  and  a67660a );
 a67665a <=( a67664a  and  a67657a );
 a67669a <=( (not A267)  and  (not A266) );
 a67670a <=( A265  and  a67669a );
 a67673a <=( A269  and  (not A268) );
 a67676a <=( A301  and  (not A300) );
 a67677a <=( a67676a  and  a67673a );
 a67678a <=( a67677a  and  a67670a );
 a67682a <=( A167  and  A168 );
 a67683a <=( A169  and  a67682a );
 a67686a <=( A201  and  (not A166) );
 a67689a <=( A203  and  (not A202) );
 a67690a <=( a67689a  and  a67686a );
 a67691a <=( a67690a  and  a67683a );
 a67695a <=( (not A267)  and  (not A266) );
 a67696a <=( A265  and  a67695a );
 a67699a <=( A269  and  (not A268) );
 a67702a <=( (not A302)  and  (not A300) );
 a67703a <=( a67702a  and  a67699a );
 a67704a <=( a67703a  and  a67696a );
 a67708a <=( A167  and  A168 );
 a67709a <=( A169  and  a67708a );
 a67712a <=( A201  and  (not A166) );
 a67715a <=( A203  and  (not A202) );
 a67716a <=( a67715a  and  a67712a );
 a67717a <=( a67716a  and  a67709a );
 a67721a <=( (not A267)  and  (not A266) );
 a67722a <=( A265  and  a67721a );
 a67725a <=( A269  and  (not A268) );
 a67728a <=( A299  and  A298 );
 a67729a <=( a67728a  and  a67725a );
 a67730a <=( a67729a  and  a67722a );
 a67734a <=( A167  and  A168 );
 a67735a <=( A169  and  a67734a );
 a67738a <=( A201  and  (not A166) );
 a67741a <=( A203  and  (not A202) );
 a67742a <=( a67741a  and  a67738a );
 a67743a <=( a67742a  and  a67735a );
 a67747a <=( (not A267)  and  (not A266) );
 a67748a <=( A265  and  a67747a );
 a67751a <=( A269  and  (not A268) );
 a67754a <=( (not A299)  and  (not A298) );
 a67755a <=( a67754a  and  a67751a );
 a67756a <=( a67755a  and  a67748a );
 a67760a <=( A167  and  A168 );
 a67761a <=( A169  and  a67760a );
 a67764a <=( A201  and  (not A166) );
 a67767a <=( A203  and  (not A202) );
 a67768a <=( a67767a  and  a67764a );
 a67769a <=( a67768a  and  a67761a );
 a67773a <=( A298  and  (not A266) );
 a67774a <=( (not A265)  and  a67773a );
 a67777a <=( (not A300)  and  (not A299) );
 a67780a <=( A302  and  (not A301) );
 a67781a <=( a67780a  and  a67777a );
 a67782a <=( a67781a  and  a67774a );
 a67786a <=( A167  and  A168 );
 a67787a <=( A169  and  a67786a );
 a67790a <=( A201  and  (not A166) );
 a67793a <=( A203  and  (not A202) );
 a67794a <=( a67793a  and  a67790a );
 a67795a <=( a67794a  and  a67787a );
 a67799a <=( (not A298)  and  (not A266) );
 a67800a <=( (not A265)  and  a67799a );
 a67803a <=( (not A300)  and  A299 );
 a67806a <=( A302  and  (not A301) );
 a67807a <=( a67806a  and  a67803a );
 a67808a <=( a67807a  and  a67800a );
 a67812a <=( A167  and  A168 );
 a67813a <=( A169  and  a67812a );
 a67816a <=( (not A201)  and  (not A166) );
 a67819a <=( A267  and  A202 );
 a67820a <=( a67819a  and  a67816a );
 a67821a <=( a67820a  and  a67813a );
 a67825a <=( A298  and  A269 );
 a67826a <=( (not A268)  and  a67825a );
 a67829a <=( (not A300)  and  (not A299) );
 a67832a <=( A302  and  (not A301) );
 a67833a <=( a67832a  and  a67829a );
 a67834a <=( a67833a  and  a67826a );
 a67838a <=( A167  and  A168 );
 a67839a <=( A169  and  a67838a );
 a67842a <=( (not A201)  and  (not A166) );
 a67845a <=( A267  and  A202 );
 a67846a <=( a67845a  and  a67842a );
 a67847a <=( a67846a  and  a67839a );
 a67851a <=( (not A298)  and  A269 );
 a67852a <=( (not A268)  and  a67851a );
 a67855a <=( (not A300)  and  A299 );
 a67858a <=( A302  and  (not A301) );
 a67859a <=( a67858a  and  a67855a );
 a67860a <=( a67859a  and  a67852a );
 a67864a <=( A167  and  A168 );
 a67865a <=( A169  and  a67864a );
 a67868a <=( (not A201)  and  (not A166) );
 a67871a <=( (not A265)  and  A202 );
 a67872a <=( a67871a  and  a67868a );
 a67873a <=( a67872a  and  a67865a );
 a67877a <=( (not A268)  and  (not A267) );
 a67878a <=( A266  and  a67877a );
 a67881a <=( A300  and  A269 );
 a67884a <=( A302  and  (not A301) );
 a67885a <=( a67884a  and  a67881a );
 a67886a <=( a67885a  and  a67878a );
 a67890a <=( A167  and  A168 );
 a67891a <=( A169  and  a67890a );
 a67894a <=( (not A201)  and  (not A166) );
 a67897a <=( A265  and  A202 );
 a67898a <=( a67897a  and  a67894a );
 a67899a <=( a67898a  and  a67891a );
 a67903a <=( (not A268)  and  (not A267) );
 a67904a <=( (not A266)  and  a67903a );
 a67907a <=( A300  and  A269 );
 a67910a <=( A302  and  (not A301) );
 a67911a <=( a67910a  and  a67907a );
 a67912a <=( a67911a  and  a67904a );
 a67916a <=( A167  and  A168 );
 a67917a <=( A169  and  a67916a );
 a67920a <=( (not A201)  and  (not A166) );
 a67923a <=( A267  and  (not A203) );
 a67924a <=( a67923a  and  a67920a );
 a67925a <=( a67924a  and  a67917a );
 a67929a <=( A298  and  A269 );
 a67930a <=( (not A268)  and  a67929a );
 a67933a <=( (not A300)  and  (not A299) );
 a67936a <=( A302  and  (not A301) );
 a67937a <=( a67936a  and  a67933a );
 a67938a <=( a67937a  and  a67930a );
 a67942a <=( A167  and  A168 );
 a67943a <=( A169  and  a67942a );
 a67946a <=( (not A201)  and  (not A166) );
 a67949a <=( A267  and  (not A203) );
 a67950a <=( a67949a  and  a67946a );
 a67951a <=( a67950a  and  a67943a );
 a67955a <=( (not A298)  and  A269 );
 a67956a <=( (not A268)  and  a67955a );
 a67959a <=( (not A300)  and  A299 );
 a67962a <=( A302  and  (not A301) );
 a67963a <=( a67962a  and  a67959a );
 a67964a <=( a67963a  and  a67956a );
 a67968a <=( A167  and  A168 );
 a67969a <=( A169  and  a67968a );
 a67972a <=( (not A201)  and  (not A166) );
 a67975a <=( (not A265)  and  (not A203) );
 a67976a <=( a67975a  and  a67972a );
 a67977a <=( a67976a  and  a67969a );
 a67981a <=( (not A268)  and  (not A267) );
 a67982a <=( A266  and  a67981a );
 a67985a <=( A300  and  A269 );
 a67988a <=( A302  and  (not A301) );
 a67989a <=( a67988a  and  a67985a );
 a67990a <=( a67989a  and  a67982a );
 a67994a <=( A167  and  A168 );
 a67995a <=( A169  and  a67994a );
 a67998a <=( (not A201)  and  (not A166) );
 a68001a <=( A265  and  (not A203) );
 a68002a <=( a68001a  and  a67998a );
 a68003a <=( a68002a  and  a67995a );
 a68007a <=( (not A268)  and  (not A267) );
 a68008a <=( (not A266)  and  a68007a );
 a68011a <=( A300  and  A269 );
 a68014a <=( A302  and  (not A301) );
 a68015a <=( a68014a  and  a68011a );
 a68016a <=( a68015a  and  a68008a );
 a68020a <=( A167  and  A168 );
 a68021a <=( A169  and  a68020a );
 a68024a <=( A199  and  (not A166) );
 a68027a <=( A267  and  A200 );
 a68028a <=( a68027a  and  a68024a );
 a68029a <=( a68028a  and  a68021a );
 a68033a <=( A298  and  A269 );
 a68034a <=( (not A268)  and  a68033a );
 a68037a <=( (not A300)  and  (not A299) );
 a68040a <=( A302  and  (not A301) );
 a68041a <=( a68040a  and  a68037a );
 a68042a <=( a68041a  and  a68034a );
 a68046a <=( A167  and  A168 );
 a68047a <=( A169  and  a68046a );
 a68050a <=( A199  and  (not A166) );
 a68053a <=( A267  and  A200 );
 a68054a <=( a68053a  and  a68050a );
 a68055a <=( a68054a  and  a68047a );
 a68059a <=( (not A298)  and  A269 );
 a68060a <=( (not A268)  and  a68059a );
 a68063a <=( (not A300)  and  A299 );
 a68066a <=( A302  and  (not A301) );
 a68067a <=( a68066a  and  a68063a );
 a68068a <=( a68067a  and  a68060a );
 a68072a <=( A167  and  A168 );
 a68073a <=( A169  and  a68072a );
 a68076a <=( A199  and  (not A166) );
 a68079a <=( (not A265)  and  A200 );
 a68080a <=( a68079a  and  a68076a );
 a68081a <=( a68080a  and  a68073a );
 a68085a <=( (not A268)  and  (not A267) );
 a68086a <=( A266  and  a68085a );
 a68089a <=( A300  and  A269 );
 a68092a <=( A302  and  (not A301) );
 a68093a <=( a68092a  and  a68089a );
 a68094a <=( a68093a  and  a68086a );
 a68098a <=( A167  and  A168 );
 a68099a <=( A169  and  a68098a );
 a68102a <=( A199  and  (not A166) );
 a68105a <=( A265  and  A200 );
 a68106a <=( a68105a  and  a68102a );
 a68107a <=( a68106a  and  a68099a );
 a68111a <=( (not A268)  and  (not A267) );
 a68112a <=( (not A266)  and  a68111a );
 a68115a <=( A300  and  A269 );
 a68118a <=( A302  and  (not A301) );
 a68119a <=( a68118a  and  a68115a );
 a68120a <=( a68119a  and  a68112a );
 a68124a <=( A167  and  A168 );
 a68125a <=( A169  and  a68124a );
 a68128a <=( (not A199)  and  (not A166) );
 a68131a <=( A267  and  (not A200) );
 a68132a <=( a68131a  and  a68128a );
 a68133a <=( a68132a  and  a68125a );
 a68137a <=( A298  and  A269 );
 a68138a <=( (not A268)  and  a68137a );
 a68141a <=( (not A300)  and  (not A299) );
 a68144a <=( A302  and  (not A301) );
 a68145a <=( a68144a  and  a68141a );
 a68146a <=( a68145a  and  a68138a );
 a68150a <=( A167  and  A168 );
 a68151a <=( A169  and  a68150a );
 a68154a <=( (not A199)  and  (not A166) );
 a68157a <=( A267  and  (not A200) );
 a68158a <=( a68157a  and  a68154a );
 a68159a <=( a68158a  and  a68151a );
 a68163a <=( (not A298)  and  A269 );
 a68164a <=( (not A268)  and  a68163a );
 a68167a <=( (not A300)  and  A299 );
 a68170a <=( A302  and  (not A301) );
 a68171a <=( a68170a  and  a68167a );
 a68172a <=( a68171a  and  a68164a );
 a68176a <=( A167  and  A168 );
 a68177a <=( A169  and  a68176a );
 a68180a <=( (not A199)  and  (not A166) );
 a68183a <=( (not A265)  and  (not A200) );
 a68184a <=( a68183a  and  a68180a );
 a68185a <=( a68184a  and  a68177a );
 a68189a <=( (not A268)  and  (not A267) );
 a68190a <=( A266  and  a68189a );
 a68193a <=( A300  and  A269 );
 a68196a <=( A302  and  (not A301) );
 a68197a <=( a68196a  and  a68193a );
 a68198a <=( a68197a  and  a68190a );
 a68202a <=( A167  and  A168 );
 a68203a <=( A169  and  a68202a );
 a68206a <=( (not A199)  and  (not A166) );
 a68209a <=( A265  and  (not A200) );
 a68210a <=( a68209a  and  a68206a );
 a68211a <=( a68210a  and  a68203a );
 a68215a <=( (not A268)  and  (not A267) );
 a68216a <=( (not A266)  and  a68215a );
 a68219a <=( A300  and  A269 );
 a68222a <=( A302  and  (not A301) );
 a68223a <=( a68222a  and  a68219a );
 a68224a <=( a68223a  and  a68216a );
 a68228a <=( (not A167)  and  A168 );
 a68229a <=( A169  and  a68228a );
 a68232a <=( A201  and  A166 );
 a68235a <=( A203  and  (not A202) );
 a68236a <=( a68235a  and  a68232a );
 a68237a <=( a68236a  and  a68229a );
 a68241a <=( A269  and  (not A268) );
 a68242a <=( A267  and  a68241a );
 a68245a <=( (not A299)  and  A298 );
 a68248a <=( A301  and  A300 );
 a68249a <=( a68248a  and  a68245a );
 a68250a <=( a68249a  and  a68242a );
 a68254a <=( (not A167)  and  A168 );
 a68255a <=( A169  and  a68254a );
 a68258a <=( A201  and  A166 );
 a68261a <=( A203  and  (not A202) );
 a68262a <=( a68261a  and  a68258a );
 a68263a <=( a68262a  and  a68255a );
 a68267a <=( A269  and  (not A268) );
 a68268a <=( A267  and  a68267a );
 a68271a <=( (not A299)  and  A298 );
 a68274a <=( (not A302)  and  A300 );
 a68275a <=( a68274a  and  a68271a );
 a68276a <=( a68275a  and  a68268a );
 a68280a <=( (not A167)  and  A168 );
 a68281a <=( A169  and  a68280a );
 a68284a <=( A201  and  A166 );
 a68287a <=( A203  and  (not A202) );
 a68288a <=( a68287a  and  a68284a );
 a68289a <=( a68288a  and  a68281a );
 a68293a <=( A269  and  (not A268) );
 a68294a <=( A267  and  a68293a );
 a68297a <=( A299  and  (not A298) );
 a68300a <=( A301  and  A300 );
 a68301a <=( a68300a  and  a68297a );
 a68302a <=( a68301a  and  a68294a );
 a68306a <=( (not A167)  and  A168 );
 a68307a <=( A169  and  a68306a );
 a68310a <=( A201  and  A166 );
 a68313a <=( A203  and  (not A202) );
 a68314a <=( a68313a  and  a68310a );
 a68315a <=( a68314a  and  a68307a );
 a68319a <=( A269  and  (not A268) );
 a68320a <=( A267  and  a68319a );
 a68323a <=( A299  and  (not A298) );
 a68326a <=( (not A302)  and  A300 );
 a68327a <=( a68326a  and  a68323a );
 a68328a <=( a68327a  and  a68320a );
 a68332a <=( (not A167)  and  A168 );
 a68333a <=( A169  and  a68332a );
 a68336a <=( A201  and  A166 );
 a68339a <=( A203  and  (not A202) );
 a68340a <=( a68339a  and  a68336a );
 a68341a <=( a68340a  and  a68333a );
 a68345a <=( A298  and  A268 );
 a68346a <=( (not A267)  and  a68345a );
 a68349a <=( (not A300)  and  (not A299) );
 a68352a <=( A302  and  (not A301) );
 a68353a <=( a68352a  and  a68349a );
 a68354a <=( a68353a  and  a68346a );
 a68358a <=( (not A167)  and  A168 );
 a68359a <=( A169  and  a68358a );
 a68362a <=( A201  and  A166 );
 a68365a <=( A203  and  (not A202) );
 a68366a <=( a68365a  and  a68362a );
 a68367a <=( a68366a  and  a68359a );
 a68371a <=( (not A298)  and  A268 );
 a68372a <=( (not A267)  and  a68371a );
 a68375a <=( (not A300)  and  A299 );
 a68378a <=( A302  and  (not A301) );
 a68379a <=( a68378a  and  a68375a );
 a68380a <=( a68379a  and  a68372a );
 a68384a <=( (not A167)  and  A168 );
 a68385a <=( A169  and  a68384a );
 a68388a <=( A201  and  A166 );
 a68391a <=( A203  and  (not A202) );
 a68392a <=( a68391a  and  a68388a );
 a68393a <=( a68392a  and  a68385a );
 a68397a <=( A298  and  (not A269) );
 a68398a <=( (not A267)  and  a68397a );
 a68401a <=( (not A300)  and  (not A299) );
 a68404a <=( A302  and  (not A301) );
 a68405a <=( a68404a  and  a68401a );
 a68406a <=( a68405a  and  a68398a );
 a68410a <=( (not A167)  and  A168 );
 a68411a <=( A169  and  a68410a );
 a68414a <=( A201  and  A166 );
 a68417a <=( A203  and  (not A202) );
 a68418a <=( a68417a  and  a68414a );
 a68419a <=( a68418a  and  a68411a );
 a68423a <=( (not A298)  and  (not A269) );
 a68424a <=( (not A267)  and  a68423a );
 a68427a <=( (not A300)  and  A299 );
 a68430a <=( A302  and  (not A301) );
 a68431a <=( a68430a  and  a68427a );
 a68432a <=( a68431a  and  a68424a );
 a68436a <=( (not A167)  and  A168 );
 a68437a <=( A169  and  a68436a );
 a68440a <=( A201  and  A166 );
 a68443a <=( A203  and  (not A202) );
 a68444a <=( a68443a  and  a68440a );
 a68445a <=( a68444a  and  a68437a );
 a68449a <=( A298  and  A266 );
 a68450a <=( A265  and  a68449a );
 a68453a <=( (not A300)  and  (not A299) );
 a68456a <=( A302  and  (not A301) );
 a68457a <=( a68456a  and  a68453a );
 a68458a <=( a68457a  and  a68450a );
 a68462a <=( (not A167)  and  A168 );
 a68463a <=( A169  and  a68462a );
 a68466a <=( A201  and  A166 );
 a68469a <=( A203  and  (not A202) );
 a68470a <=( a68469a  and  a68466a );
 a68471a <=( a68470a  and  a68463a );
 a68475a <=( (not A298)  and  A266 );
 a68476a <=( A265  and  a68475a );
 a68479a <=( (not A300)  and  A299 );
 a68482a <=( A302  and  (not A301) );
 a68483a <=( a68482a  and  a68479a );
 a68484a <=( a68483a  and  a68476a );
 a68488a <=( (not A167)  and  A168 );
 a68489a <=( A169  and  a68488a );
 a68492a <=( A201  and  A166 );
 a68495a <=( A203  and  (not A202) );
 a68496a <=( a68495a  and  a68492a );
 a68497a <=( a68496a  and  a68489a );
 a68501a <=( A267  and  A266 );
 a68502a <=( (not A265)  and  a68501a );
 a68505a <=( A300  and  A268 );
 a68508a <=( A302  and  (not A301) );
 a68509a <=( a68508a  and  a68505a );
 a68510a <=( a68509a  and  a68502a );
 a68514a <=( (not A167)  and  A168 );
 a68515a <=( A169  and  a68514a );
 a68518a <=( A201  and  A166 );
 a68521a <=( A203  and  (not A202) );
 a68522a <=( a68521a  and  a68518a );
 a68523a <=( a68522a  and  a68515a );
 a68527a <=( A267  and  A266 );
 a68528a <=( (not A265)  and  a68527a );
 a68531a <=( A300  and  (not A269) );
 a68534a <=( A302  and  (not A301) );
 a68535a <=( a68534a  and  a68531a );
 a68536a <=( a68535a  and  a68528a );
 a68540a <=( (not A167)  and  A168 );
 a68541a <=( A169  and  a68540a );
 a68544a <=( A201  and  A166 );
 a68547a <=( A203  and  (not A202) );
 a68548a <=( a68547a  and  a68544a );
 a68549a <=( a68548a  and  a68541a );
 a68553a <=( (not A267)  and  A266 );
 a68554a <=( (not A265)  and  a68553a );
 a68557a <=( A269  and  (not A268) );
 a68560a <=( A301  and  (not A300) );
 a68561a <=( a68560a  and  a68557a );
 a68562a <=( a68561a  and  a68554a );
 a68566a <=( (not A167)  and  A168 );
 a68567a <=( A169  and  a68566a );
 a68570a <=( A201  and  A166 );
 a68573a <=( A203  and  (not A202) );
 a68574a <=( a68573a  and  a68570a );
 a68575a <=( a68574a  and  a68567a );
 a68579a <=( (not A267)  and  A266 );
 a68580a <=( (not A265)  and  a68579a );
 a68583a <=( A269  and  (not A268) );
 a68586a <=( (not A302)  and  (not A300) );
 a68587a <=( a68586a  and  a68583a );
 a68588a <=( a68587a  and  a68580a );
 a68592a <=( (not A167)  and  A168 );
 a68593a <=( A169  and  a68592a );
 a68596a <=( A201  and  A166 );
 a68599a <=( A203  and  (not A202) );
 a68600a <=( a68599a  and  a68596a );
 a68601a <=( a68600a  and  a68593a );
 a68605a <=( (not A267)  and  A266 );
 a68606a <=( (not A265)  and  a68605a );
 a68609a <=( A269  and  (not A268) );
 a68612a <=( A299  and  A298 );
 a68613a <=( a68612a  and  a68609a );
 a68614a <=( a68613a  and  a68606a );
 a68618a <=( (not A167)  and  A168 );
 a68619a <=( A169  and  a68618a );
 a68622a <=( A201  and  A166 );
 a68625a <=( A203  and  (not A202) );
 a68626a <=( a68625a  and  a68622a );
 a68627a <=( a68626a  and  a68619a );
 a68631a <=( (not A267)  and  A266 );
 a68632a <=( (not A265)  and  a68631a );
 a68635a <=( A269  and  (not A268) );
 a68638a <=( (not A299)  and  (not A298) );
 a68639a <=( a68638a  and  a68635a );
 a68640a <=( a68639a  and  a68632a );
 a68644a <=( (not A167)  and  A168 );
 a68645a <=( A169  and  a68644a );
 a68648a <=( A201  and  A166 );
 a68651a <=( A203  and  (not A202) );
 a68652a <=( a68651a  and  a68648a );
 a68653a <=( a68652a  and  a68645a );
 a68657a <=( A267  and  (not A266) );
 a68658a <=( A265  and  a68657a );
 a68661a <=( A300  and  A268 );
 a68664a <=( A302  and  (not A301) );
 a68665a <=( a68664a  and  a68661a );
 a68666a <=( a68665a  and  a68658a );
 a68670a <=( (not A167)  and  A168 );
 a68671a <=( A169  and  a68670a );
 a68674a <=( A201  and  A166 );
 a68677a <=( A203  and  (not A202) );
 a68678a <=( a68677a  and  a68674a );
 a68679a <=( a68678a  and  a68671a );
 a68683a <=( A267  and  (not A266) );
 a68684a <=( A265  and  a68683a );
 a68687a <=( A300  and  (not A269) );
 a68690a <=( A302  and  (not A301) );
 a68691a <=( a68690a  and  a68687a );
 a68692a <=( a68691a  and  a68684a );
 a68696a <=( (not A167)  and  A168 );
 a68697a <=( A169  and  a68696a );
 a68700a <=( A201  and  A166 );
 a68703a <=( A203  and  (not A202) );
 a68704a <=( a68703a  and  a68700a );
 a68705a <=( a68704a  and  a68697a );
 a68709a <=( (not A267)  and  (not A266) );
 a68710a <=( A265  and  a68709a );
 a68713a <=( A269  and  (not A268) );
 a68716a <=( A301  and  (not A300) );
 a68717a <=( a68716a  and  a68713a );
 a68718a <=( a68717a  and  a68710a );
 a68722a <=( (not A167)  and  A168 );
 a68723a <=( A169  and  a68722a );
 a68726a <=( A201  and  A166 );
 a68729a <=( A203  and  (not A202) );
 a68730a <=( a68729a  and  a68726a );
 a68731a <=( a68730a  and  a68723a );
 a68735a <=( (not A267)  and  (not A266) );
 a68736a <=( A265  and  a68735a );
 a68739a <=( A269  and  (not A268) );
 a68742a <=( (not A302)  and  (not A300) );
 a68743a <=( a68742a  and  a68739a );
 a68744a <=( a68743a  and  a68736a );
 a68748a <=( (not A167)  and  A168 );
 a68749a <=( A169  and  a68748a );
 a68752a <=( A201  and  A166 );
 a68755a <=( A203  and  (not A202) );
 a68756a <=( a68755a  and  a68752a );
 a68757a <=( a68756a  and  a68749a );
 a68761a <=( (not A267)  and  (not A266) );
 a68762a <=( A265  and  a68761a );
 a68765a <=( A269  and  (not A268) );
 a68768a <=( A299  and  A298 );
 a68769a <=( a68768a  and  a68765a );
 a68770a <=( a68769a  and  a68762a );
 a68774a <=( (not A167)  and  A168 );
 a68775a <=( A169  and  a68774a );
 a68778a <=( A201  and  A166 );
 a68781a <=( A203  and  (not A202) );
 a68782a <=( a68781a  and  a68778a );
 a68783a <=( a68782a  and  a68775a );
 a68787a <=( (not A267)  and  (not A266) );
 a68788a <=( A265  and  a68787a );
 a68791a <=( A269  and  (not A268) );
 a68794a <=( (not A299)  and  (not A298) );
 a68795a <=( a68794a  and  a68791a );
 a68796a <=( a68795a  and  a68788a );
 a68800a <=( (not A167)  and  A168 );
 a68801a <=( A169  and  a68800a );
 a68804a <=( A201  and  A166 );
 a68807a <=( A203  and  (not A202) );
 a68808a <=( a68807a  and  a68804a );
 a68809a <=( a68808a  and  a68801a );
 a68813a <=( A298  and  (not A266) );
 a68814a <=( (not A265)  and  a68813a );
 a68817a <=( (not A300)  and  (not A299) );
 a68820a <=( A302  and  (not A301) );
 a68821a <=( a68820a  and  a68817a );
 a68822a <=( a68821a  and  a68814a );
 a68826a <=( (not A167)  and  A168 );
 a68827a <=( A169  and  a68826a );
 a68830a <=( A201  and  A166 );
 a68833a <=( A203  and  (not A202) );
 a68834a <=( a68833a  and  a68830a );
 a68835a <=( a68834a  and  a68827a );
 a68839a <=( (not A298)  and  (not A266) );
 a68840a <=( (not A265)  and  a68839a );
 a68843a <=( (not A300)  and  A299 );
 a68846a <=( A302  and  (not A301) );
 a68847a <=( a68846a  and  a68843a );
 a68848a <=( a68847a  and  a68840a );
 a68852a <=( (not A167)  and  A168 );
 a68853a <=( A169  and  a68852a );
 a68856a <=( (not A201)  and  A166 );
 a68859a <=( A267  and  A202 );
 a68860a <=( a68859a  and  a68856a );
 a68861a <=( a68860a  and  a68853a );
 a68865a <=( A298  and  A269 );
 a68866a <=( (not A268)  and  a68865a );
 a68869a <=( (not A300)  and  (not A299) );
 a68872a <=( A302  and  (not A301) );
 a68873a <=( a68872a  and  a68869a );
 a68874a <=( a68873a  and  a68866a );
 a68878a <=( (not A167)  and  A168 );
 a68879a <=( A169  and  a68878a );
 a68882a <=( (not A201)  and  A166 );
 a68885a <=( A267  and  A202 );
 a68886a <=( a68885a  and  a68882a );
 a68887a <=( a68886a  and  a68879a );
 a68891a <=( (not A298)  and  A269 );
 a68892a <=( (not A268)  and  a68891a );
 a68895a <=( (not A300)  and  A299 );
 a68898a <=( A302  and  (not A301) );
 a68899a <=( a68898a  and  a68895a );
 a68900a <=( a68899a  and  a68892a );
 a68904a <=( (not A167)  and  A168 );
 a68905a <=( A169  and  a68904a );
 a68908a <=( (not A201)  and  A166 );
 a68911a <=( (not A265)  and  A202 );
 a68912a <=( a68911a  and  a68908a );
 a68913a <=( a68912a  and  a68905a );
 a68917a <=( (not A268)  and  (not A267) );
 a68918a <=( A266  and  a68917a );
 a68921a <=( A300  and  A269 );
 a68924a <=( A302  and  (not A301) );
 a68925a <=( a68924a  and  a68921a );
 a68926a <=( a68925a  and  a68918a );
 a68930a <=( (not A167)  and  A168 );
 a68931a <=( A169  and  a68930a );
 a68934a <=( (not A201)  and  A166 );
 a68937a <=( A265  and  A202 );
 a68938a <=( a68937a  and  a68934a );
 a68939a <=( a68938a  and  a68931a );
 a68943a <=( (not A268)  and  (not A267) );
 a68944a <=( (not A266)  and  a68943a );
 a68947a <=( A300  and  A269 );
 a68950a <=( A302  and  (not A301) );
 a68951a <=( a68950a  and  a68947a );
 a68952a <=( a68951a  and  a68944a );
 a68956a <=( (not A167)  and  A168 );
 a68957a <=( A169  and  a68956a );
 a68960a <=( (not A201)  and  A166 );
 a68963a <=( A267  and  (not A203) );
 a68964a <=( a68963a  and  a68960a );
 a68965a <=( a68964a  and  a68957a );
 a68969a <=( A298  and  A269 );
 a68970a <=( (not A268)  and  a68969a );
 a68973a <=( (not A300)  and  (not A299) );
 a68976a <=( A302  and  (not A301) );
 a68977a <=( a68976a  and  a68973a );
 a68978a <=( a68977a  and  a68970a );
 a68982a <=( (not A167)  and  A168 );
 a68983a <=( A169  and  a68982a );
 a68986a <=( (not A201)  and  A166 );
 a68989a <=( A267  and  (not A203) );
 a68990a <=( a68989a  and  a68986a );
 a68991a <=( a68990a  and  a68983a );
 a68995a <=( (not A298)  and  A269 );
 a68996a <=( (not A268)  and  a68995a );
 a68999a <=( (not A300)  and  A299 );
 a69002a <=( A302  and  (not A301) );
 a69003a <=( a69002a  and  a68999a );
 a69004a <=( a69003a  and  a68996a );
 a69008a <=( (not A167)  and  A168 );
 a69009a <=( A169  and  a69008a );
 a69012a <=( (not A201)  and  A166 );
 a69015a <=( (not A265)  and  (not A203) );
 a69016a <=( a69015a  and  a69012a );
 a69017a <=( a69016a  and  a69009a );
 a69021a <=( (not A268)  and  (not A267) );
 a69022a <=( A266  and  a69021a );
 a69025a <=( A300  and  A269 );
 a69028a <=( A302  and  (not A301) );
 a69029a <=( a69028a  and  a69025a );
 a69030a <=( a69029a  and  a69022a );
 a69034a <=( (not A167)  and  A168 );
 a69035a <=( A169  and  a69034a );
 a69038a <=( (not A201)  and  A166 );
 a69041a <=( A265  and  (not A203) );
 a69042a <=( a69041a  and  a69038a );
 a69043a <=( a69042a  and  a69035a );
 a69047a <=( (not A268)  and  (not A267) );
 a69048a <=( (not A266)  and  a69047a );
 a69051a <=( A300  and  A269 );
 a69054a <=( A302  and  (not A301) );
 a69055a <=( a69054a  and  a69051a );
 a69056a <=( a69055a  and  a69048a );
 a69060a <=( (not A167)  and  A168 );
 a69061a <=( A169  and  a69060a );
 a69064a <=( A199  and  A166 );
 a69067a <=( A267  and  A200 );
 a69068a <=( a69067a  and  a69064a );
 a69069a <=( a69068a  and  a69061a );
 a69073a <=( A298  and  A269 );
 a69074a <=( (not A268)  and  a69073a );
 a69077a <=( (not A300)  and  (not A299) );
 a69080a <=( A302  and  (not A301) );
 a69081a <=( a69080a  and  a69077a );
 a69082a <=( a69081a  and  a69074a );
 a69086a <=( (not A167)  and  A168 );
 a69087a <=( A169  and  a69086a );
 a69090a <=( A199  and  A166 );
 a69093a <=( A267  and  A200 );
 a69094a <=( a69093a  and  a69090a );
 a69095a <=( a69094a  and  a69087a );
 a69099a <=( (not A298)  and  A269 );
 a69100a <=( (not A268)  and  a69099a );
 a69103a <=( (not A300)  and  A299 );
 a69106a <=( A302  and  (not A301) );
 a69107a <=( a69106a  and  a69103a );
 a69108a <=( a69107a  and  a69100a );
 a69112a <=( (not A167)  and  A168 );
 a69113a <=( A169  and  a69112a );
 a69116a <=( A199  and  A166 );
 a69119a <=( (not A265)  and  A200 );
 a69120a <=( a69119a  and  a69116a );
 a69121a <=( a69120a  and  a69113a );
 a69125a <=( (not A268)  and  (not A267) );
 a69126a <=( A266  and  a69125a );
 a69129a <=( A300  and  A269 );
 a69132a <=( A302  and  (not A301) );
 a69133a <=( a69132a  and  a69129a );
 a69134a <=( a69133a  and  a69126a );
 a69138a <=( (not A167)  and  A168 );
 a69139a <=( A169  and  a69138a );
 a69142a <=( A199  and  A166 );
 a69145a <=( A265  and  A200 );
 a69146a <=( a69145a  and  a69142a );
 a69147a <=( a69146a  and  a69139a );
 a69151a <=( (not A268)  and  (not A267) );
 a69152a <=( (not A266)  and  a69151a );
 a69155a <=( A300  and  A269 );
 a69158a <=( A302  and  (not A301) );
 a69159a <=( a69158a  and  a69155a );
 a69160a <=( a69159a  and  a69152a );
 a69164a <=( (not A167)  and  A168 );
 a69165a <=( A169  and  a69164a );
 a69168a <=( (not A199)  and  A166 );
 a69171a <=( A267  and  (not A200) );
 a69172a <=( a69171a  and  a69168a );
 a69173a <=( a69172a  and  a69165a );
 a69177a <=( A298  and  A269 );
 a69178a <=( (not A268)  and  a69177a );
 a69181a <=( (not A300)  and  (not A299) );
 a69184a <=( A302  and  (not A301) );
 a69185a <=( a69184a  and  a69181a );
 a69186a <=( a69185a  and  a69178a );
 a69190a <=( (not A167)  and  A168 );
 a69191a <=( A169  and  a69190a );
 a69194a <=( (not A199)  and  A166 );
 a69197a <=( A267  and  (not A200) );
 a69198a <=( a69197a  and  a69194a );
 a69199a <=( a69198a  and  a69191a );
 a69203a <=( (not A298)  and  A269 );
 a69204a <=( (not A268)  and  a69203a );
 a69207a <=( (not A300)  and  A299 );
 a69210a <=( A302  and  (not A301) );
 a69211a <=( a69210a  and  a69207a );
 a69212a <=( a69211a  and  a69204a );
 a69216a <=( (not A167)  and  A168 );
 a69217a <=( A169  and  a69216a );
 a69220a <=( (not A199)  and  A166 );
 a69223a <=( (not A265)  and  (not A200) );
 a69224a <=( a69223a  and  a69220a );
 a69225a <=( a69224a  and  a69217a );
 a69229a <=( (not A268)  and  (not A267) );
 a69230a <=( A266  and  a69229a );
 a69233a <=( A300  and  A269 );
 a69236a <=( A302  and  (not A301) );
 a69237a <=( a69236a  and  a69233a );
 a69238a <=( a69237a  and  a69230a );
 a69242a <=( (not A167)  and  A168 );
 a69243a <=( A169  and  a69242a );
 a69246a <=( (not A199)  and  A166 );
 a69249a <=( A265  and  (not A200) );
 a69250a <=( a69249a  and  a69246a );
 a69251a <=( a69250a  and  a69243a );
 a69255a <=( (not A268)  and  (not A267) );
 a69256a <=( (not A266)  and  a69255a );
 a69259a <=( A300  and  A269 );
 a69262a <=( A302  and  (not A301) );
 a69263a <=( a69262a  and  a69259a );
 a69264a <=( a69263a  and  a69256a );
 a69268a <=( (not A199)  and  (not A168) );
 a69269a <=( A169  and  a69268a );
 a69272a <=( A201  and  A200 );
 a69275a <=( (not A265)  and  A202 );
 a69276a <=( a69275a  and  a69272a );
 a69277a <=( a69276a  and  a69269a );
 a69281a <=( A268  and  A267 );
 a69282a <=( A266  and  a69281a );
 a69285a <=( (not A299)  and  A298 );
 a69288a <=( A301  and  A300 );
 a69289a <=( a69288a  and  a69285a );
 a69290a <=( a69289a  and  a69282a );
 a69294a <=( (not A199)  and  (not A168) );
 a69295a <=( A169  and  a69294a );
 a69298a <=( A201  and  A200 );
 a69301a <=( (not A265)  and  A202 );
 a69302a <=( a69301a  and  a69298a );
 a69303a <=( a69302a  and  a69295a );
 a69307a <=( A268  and  A267 );
 a69308a <=( A266  and  a69307a );
 a69311a <=( (not A299)  and  A298 );
 a69314a <=( (not A302)  and  A300 );
 a69315a <=( a69314a  and  a69311a );
 a69316a <=( a69315a  and  a69308a );
 a69320a <=( (not A199)  and  (not A168) );
 a69321a <=( A169  and  a69320a );
 a69324a <=( A201  and  A200 );
 a69327a <=( (not A265)  and  A202 );
 a69328a <=( a69327a  and  a69324a );
 a69329a <=( a69328a  and  a69321a );
 a69333a <=( A268  and  A267 );
 a69334a <=( A266  and  a69333a );
 a69337a <=( A299  and  (not A298) );
 a69340a <=( A301  and  A300 );
 a69341a <=( a69340a  and  a69337a );
 a69342a <=( a69341a  and  a69334a );
 a69346a <=( (not A199)  and  (not A168) );
 a69347a <=( A169  and  a69346a );
 a69350a <=( A201  and  A200 );
 a69353a <=( (not A265)  and  A202 );
 a69354a <=( a69353a  and  a69350a );
 a69355a <=( a69354a  and  a69347a );
 a69359a <=( A268  and  A267 );
 a69360a <=( A266  and  a69359a );
 a69363a <=( A299  and  (not A298) );
 a69366a <=( (not A302)  and  A300 );
 a69367a <=( a69366a  and  a69363a );
 a69368a <=( a69367a  and  a69360a );
 a69372a <=( (not A199)  and  (not A168) );
 a69373a <=( A169  and  a69372a );
 a69376a <=( A201  and  A200 );
 a69379a <=( (not A265)  and  A202 );
 a69380a <=( a69379a  and  a69376a );
 a69381a <=( a69380a  and  a69373a );
 a69385a <=( (not A269)  and  A267 );
 a69386a <=( A266  and  a69385a );
 a69389a <=( (not A299)  and  A298 );
 a69392a <=( A301  and  A300 );
 a69393a <=( a69392a  and  a69389a );
 a69394a <=( a69393a  and  a69386a );
 a69398a <=( (not A199)  and  (not A168) );
 a69399a <=( A169  and  a69398a );
 a69402a <=( A201  and  A200 );
 a69405a <=( (not A265)  and  A202 );
 a69406a <=( a69405a  and  a69402a );
 a69407a <=( a69406a  and  a69399a );
 a69411a <=( (not A269)  and  A267 );
 a69412a <=( A266  and  a69411a );
 a69415a <=( (not A299)  and  A298 );
 a69418a <=( (not A302)  and  A300 );
 a69419a <=( a69418a  and  a69415a );
 a69420a <=( a69419a  and  a69412a );
 a69424a <=( (not A199)  and  (not A168) );
 a69425a <=( A169  and  a69424a );
 a69428a <=( A201  and  A200 );
 a69431a <=( (not A265)  and  A202 );
 a69432a <=( a69431a  and  a69428a );
 a69433a <=( a69432a  and  a69425a );
 a69437a <=( (not A269)  and  A267 );
 a69438a <=( A266  and  a69437a );
 a69441a <=( A299  and  (not A298) );
 a69444a <=( A301  and  A300 );
 a69445a <=( a69444a  and  a69441a );
 a69446a <=( a69445a  and  a69438a );
 a69450a <=( (not A199)  and  (not A168) );
 a69451a <=( A169  and  a69450a );
 a69454a <=( A201  and  A200 );
 a69457a <=( (not A265)  and  A202 );
 a69458a <=( a69457a  and  a69454a );
 a69459a <=( a69458a  and  a69451a );
 a69463a <=( (not A269)  and  A267 );
 a69464a <=( A266  and  a69463a );
 a69467a <=( A299  and  (not A298) );
 a69470a <=( (not A302)  and  A300 );
 a69471a <=( a69470a  and  a69467a );
 a69472a <=( a69471a  and  a69464a );
 a69476a <=( (not A199)  and  (not A168) );
 a69477a <=( A169  and  a69476a );
 a69480a <=( A201  and  A200 );
 a69483a <=( A265  and  A202 );
 a69484a <=( a69483a  and  a69480a );
 a69485a <=( a69484a  and  a69477a );
 a69489a <=( A268  and  A267 );
 a69490a <=( (not A266)  and  a69489a );
 a69493a <=( (not A299)  and  A298 );
 a69496a <=( A301  and  A300 );
 a69497a <=( a69496a  and  a69493a );
 a69498a <=( a69497a  and  a69490a );
 a69502a <=( (not A199)  and  (not A168) );
 a69503a <=( A169  and  a69502a );
 a69506a <=( A201  and  A200 );
 a69509a <=( A265  and  A202 );
 a69510a <=( a69509a  and  a69506a );
 a69511a <=( a69510a  and  a69503a );
 a69515a <=( A268  and  A267 );
 a69516a <=( (not A266)  and  a69515a );
 a69519a <=( (not A299)  and  A298 );
 a69522a <=( (not A302)  and  A300 );
 a69523a <=( a69522a  and  a69519a );
 a69524a <=( a69523a  and  a69516a );
 a69528a <=( (not A199)  and  (not A168) );
 a69529a <=( A169  and  a69528a );
 a69532a <=( A201  and  A200 );
 a69535a <=( A265  and  A202 );
 a69536a <=( a69535a  and  a69532a );
 a69537a <=( a69536a  and  a69529a );
 a69541a <=( A268  and  A267 );
 a69542a <=( (not A266)  and  a69541a );
 a69545a <=( A299  and  (not A298) );
 a69548a <=( A301  and  A300 );
 a69549a <=( a69548a  and  a69545a );
 a69550a <=( a69549a  and  a69542a );
 a69554a <=( (not A199)  and  (not A168) );
 a69555a <=( A169  and  a69554a );
 a69558a <=( A201  and  A200 );
 a69561a <=( A265  and  A202 );
 a69562a <=( a69561a  and  a69558a );
 a69563a <=( a69562a  and  a69555a );
 a69567a <=( A268  and  A267 );
 a69568a <=( (not A266)  and  a69567a );
 a69571a <=( A299  and  (not A298) );
 a69574a <=( (not A302)  and  A300 );
 a69575a <=( a69574a  and  a69571a );
 a69576a <=( a69575a  and  a69568a );
 a69580a <=( (not A199)  and  (not A168) );
 a69581a <=( A169  and  a69580a );
 a69584a <=( A201  and  A200 );
 a69587a <=( A265  and  A202 );
 a69588a <=( a69587a  and  a69584a );
 a69589a <=( a69588a  and  a69581a );
 a69593a <=( (not A269)  and  A267 );
 a69594a <=( (not A266)  and  a69593a );
 a69597a <=( (not A299)  and  A298 );
 a69600a <=( A301  and  A300 );
 a69601a <=( a69600a  and  a69597a );
 a69602a <=( a69601a  and  a69594a );
 a69606a <=( (not A199)  and  (not A168) );
 a69607a <=( A169  and  a69606a );
 a69610a <=( A201  and  A200 );
 a69613a <=( A265  and  A202 );
 a69614a <=( a69613a  and  a69610a );
 a69615a <=( a69614a  and  a69607a );
 a69619a <=( (not A269)  and  A267 );
 a69620a <=( (not A266)  and  a69619a );
 a69623a <=( (not A299)  and  A298 );
 a69626a <=( (not A302)  and  A300 );
 a69627a <=( a69626a  and  a69623a );
 a69628a <=( a69627a  and  a69620a );
 a69632a <=( (not A199)  and  (not A168) );
 a69633a <=( A169  and  a69632a );
 a69636a <=( A201  and  A200 );
 a69639a <=( A265  and  A202 );
 a69640a <=( a69639a  and  a69636a );
 a69641a <=( a69640a  and  a69633a );
 a69645a <=( (not A269)  and  A267 );
 a69646a <=( (not A266)  and  a69645a );
 a69649a <=( A299  and  (not A298) );
 a69652a <=( A301  and  A300 );
 a69653a <=( a69652a  and  a69649a );
 a69654a <=( a69653a  and  a69646a );
 a69658a <=( (not A199)  and  (not A168) );
 a69659a <=( A169  and  a69658a );
 a69662a <=( A201  and  A200 );
 a69665a <=( A265  and  A202 );
 a69666a <=( a69665a  and  a69662a );
 a69667a <=( a69666a  and  a69659a );
 a69671a <=( (not A269)  and  A267 );
 a69672a <=( (not A266)  and  a69671a );
 a69675a <=( A299  and  (not A298) );
 a69678a <=( (not A302)  and  A300 );
 a69679a <=( a69678a  and  a69675a );
 a69680a <=( a69679a  and  a69672a );
 a69684a <=( (not A199)  and  (not A168) );
 a69685a <=( A169  and  a69684a );
 a69688a <=( A201  and  A200 );
 a69691a <=( (not A265)  and  (not A203) );
 a69692a <=( a69691a  and  a69688a );
 a69693a <=( a69692a  and  a69685a );
 a69697a <=( A268  and  A267 );
 a69698a <=( A266  and  a69697a );
 a69701a <=( (not A299)  and  A298 );
 a69704a <=( A301  and  A300 );
 a69705a <=( a69704a  and  a69701a );
 a69706a <=( a69705a  and  a69698a );
 a69710a <=( (not A199)  and  (not A168) );
 a69711a <=( A169  and  a69710a );
 a69714a <=( A201  and  A200 );
 a69717a <=( (not A265)  and  (not A203) );
 a69718a <=( a69717a  and  a69714a );
 a69719a <=( a69718a  and  a69711a );
 a69723a <=( A268  and  A267 );
 a69724a <=( A266  and  a69723a );
 a69727a <=( (not A299)  and  A298 );
 a69730a <=( (not A302)  and  A300 );
 a69731a <=( a69730a  and  a69727a );
 a69732a <=( a69731a  and  a69724a );
 a69736a <=( (not A199)  and  (not A168) );
 a69737a <=( A169  and  a69736a );
 a69740a <=( A201  and  A200 );
 a69743a <=( (not A265)  and  (not A203) );
 a69744a <=( a69743a  and  a69740a );
 a69745a <=( a69744a  and  a69737a );
 a69749a <=( A268  and  A267 );
 a69750a <=( A266  and  a69749a );
 a69753a <=( A299  and  (not A298) );
 a69756a <=( A301  and  A300 );
 a69757a <=( a69756a  and  a69753a );
 a69758a <=( a69757a  and  a69750a );
 a69762a <=( (not A199)  and  (not A168) );
 a69763a <=( A169  and  a69762a );
 a69766a <=( A201  and  A200 );
 a69769a <=( (not A265)  and  (not A203) );
 a69770a <=( a69769a  and  a69766a );
 a69771a <=( a69770a  and  a69763a );
 a69775a <=( A268  and  A267 );
 a69776a <=( A266  and  a69775a );
 a69779a <=( A299  and  (not A298) );
 a69782a <=( (not A302)  and  A300 );
 a69783a <=( a69782a  and  a69779a );
 a69784a <=( a69783a  and  a69776a );
 a69788a <=( (not A199)  and  (not A168) );
 a69789a <=( A169  and  a69788a );
 a69792a <=( A201  and  A200 );
 a69795a <=( (not A265)  and  (not A203) );
 a69796a <=( a69795a  and  a69792a );
 a69797a <=( a69796a  and  a69789a );
 a69801a <=( (not A269)  and  A267 );
 a69802a <=( A266  and  a69801a );
 a69805a <=( (not A299)  and  A298 );
 a69808a <=( A301  and  A300 );
 a69809a <=( a69808a  and  a69805a );
 a69810a <=( a69809a  and  a69802a );
 a69814a <=( (not A199)  and  (not A168) );
 a69815a <=( A169  and  a69814a );
 a69818a <=( A201  and  A200 );
 a69821a <=( (not A265)  and  (not A203) );
 a69822a <=( a69821a  and  a69818a );
 a69823a <=( a69822a  and  a69815a );
 a69827a <=( (not A269)  and  A267 );
 a69828a <=( A266  and  a69827a );
 a69831a <=( (not A299)  and  A298 );
 a69834a <=( (not A302)  and  A300 );
 a69835a <=( a69834a  and  a69831a );
 a69836a <=( a69835a  and  a69828a );
 a69840a <=( (not A199)  and  (not A168) );
 a69841a <=( A169  and  a69840a );
 a69844a <=( A201  and  A200 );
 a69847a <=( (not A265)  and  (not A203) );
 a69848a <=( a69847a  and  a69844a );
 a69849a <=( a69848a  and  a69841a );
 a69853a <=( (not A269)  and  A267 );
 a69854a <=( A266  and  a69853a );
 a69857a <=( A299  and  (not A298) );
 a69860a <=( A301  and  A300 );
 a69861a <=( a69860a  and  a69857a );
 a69862a <=( a69861a  and  a69854a );
 a69866a <=( (not A199)  and  (not A168) );
 a69867a <=( A169  and  a69866a );
 a69870a <=( A201  and  A200 );
 a69873a <=( (not A265)  and  (not A203) );
 a69874a <=( a69873a  and  a69870a );
 a69875a <=( a69874a  and  a69867a );
 a69879a <=( (not A269)  and  A267 );
 a69880a <=( A266  and  a69879a );
 a69883a <=( A299  and  (not A298) );
 a69886a <=( (not A302)  and  A300 );
 a69887a <=( a69886a  and  a69883a );
 a69888a <=( a69887a  and  a69880a );
 a69892a <=( (not A199)  and  (not A168) );
 a69893a <=( A169  and  a69892a );
 a69896a <=( A201  and  A200 );
 a69899a <=( A265  and  (not A203) );
 a69900a <=( a69899a  and  a69896a );
 a69901a <=( a69900a  and  a69893a );
 a69905a <=( A268  and  A267 );
 a69906a <=( (not A266)  and  a69905a );
 a69909a <=( (not A299)  and  A298 );
 a69912a <=( A301  and  A300 );
 a69913a <=( a69912a  and  a69909a );
 a69914a <=( a69913a  and  a69906a );
 a69918a <=( (not A199)  and  (not A168) );
 a69919a <=( A169  and  a69918a );
 a69922a <=( A201  and  A200 );
 a69925a <=( A265  and  (not A203) );
 a69926a <=( a69925a  and  a69922a );
 a69927a <=( a69926a  and  a69919a );
 a69931a <=( A268  and  A267 );
 a69932a <=( (not A266)  and  a69931a );
 a69935a <=( (not A299)  and  A298 );
 a69938a <=( (not A302)  and  A300 );
 a69939a <=( a69938a  and  a69935a );
 a69940a <=( a69939a  and  a69932a );
 a69944a <=( (not A199)  and  (not A168) );
 a69945a <=( A169  and  a69944a );
 a69948a <=( A201  and  A200 );
 a69951a <=( A265  and  (not A203) );
 a69952a <=( a69951a  and  a69948a );
 a69953a <=( a69952a  and  a69945a );
 a69957a <=( A268  and  A267 );
 a69958a <=( (not A266)  and  a69957a );
 a69961a <=( A299  and  (not A298) );
 a69964a <=( A301  and  A300 );
 a69965a <=( a69964a  and  a69961a );
 a69966a <=( a69965a  and  a69958a );
 a69970a <=( (not A199)  and  (not A168) );
 a69971a <=( A169  and  a69970a );
 a69974a <=( A201  and  A200 );
 a69977a <=( A265  and  (not A203) );
 a69978a <=( a69977a  and  a69974a );
 a69979a <=( a69978a  and  a69971a );
 a69983a <=( A268  and  A267 );
 a69984a <=( (not A266)  and  a69983a );
 a69987a <=( A299  and  (not A298) );
 a69990a <=( (not A302)  and  A300 );
 a69991a <=( a69990a  and  a69987a );
 a69992a <=( a69991a  and  a69984a );
 a69996a <=( (not A199)  and  (not A168) );
 a69997a <=( A169  and  a69996a );
 a70000a <=( A201  and  A200 );
 a70003a <=( A265  and  (not A203) );
 a70004a <=( a70003a  and  a70000a );
 a70005a <=( a70004a  and  a69997a );
 a70009a <=( (not A269)  and  A267 );
 a70010a <=( (not A266)  and  a70009a );
 a70013a <=( (not A299)  and  A298 );
 a70016a <=( A301  and  A300 );
 a70017a <=( a70016a  and  a70013a );
 a70018a <=( a70017a  and  a70010a );
 a70022a <=( (not A199)  and  (not A168) );
 a70023a <=( A169  and  a70022a );
 a70026a <=( A201  and  A200 );
 a70029a <=( A265  and  (not A203) );
 a70030a <=( a70029a  and  a70026a );
 a70031a <=( a70030a  and  a70023a );
 a70035a <=( (not A269)  and  A267 );
 a70036a <=( (not A266)  and  a70035a );
 a70039a <=( (not A299)  and  A298 );
 a70042a <=( (not A302)  and  A300 );
 a70043a <=( a70042a  and  a70039a );
 a70044a <=( a70043a  and  a70036a );
 a70048a <=( (not A199)  and  (not A168) );
 a70049a <=( A169  and  a70048a );
 a70052a <=( A201  and  A200 );
 a70055a <=( A265  and  (not A203) );
 a70056a <=( a70055a  and  a70052a );
 a70057a <=( a70056a  and  a70049a );
 a70061a <=( (not A269)  and  A267 );
 a70062a <=( (not A266)  and  a70061a );
 a70065a <=( A299  and  (not A298) );
 a70068a <=( A301  and  A300 );
 a70069a <=( a70068a  and  a70065a );
 a70070a <=( a70069a  and  a70062a );
 a70074a <=( (not A199)  and  (not A168) );
 a70075a <=( A169  and  a70074a );
 a70078a <=( A201  and  A200 );
 a70081a <=( A265  and  (not A203) );
 a70082a <=( a70081a  and  a70078a );
 a70083a <=( a70082a  and  a70075a );
 a70087a <=( (not A269)  and  A267 );
 a70088a <=( (not A266)  and  a70087a );
 a70091a <=( A299  and  (not A298) );
 a70094a <=( (not A302)  and  A300 );
 a70095a <=( a70094a  and  a70091a );
 a70096a <=( a70095a  and  a70088a );
 a70100a <=( A199  and  (not A168) );
 a70101a <=( A169  and  a70100a );
 a70104a <=( A201  and  (not A200) );
 a70107a <=( (not A265)  and  A202 );
 a70108a <=( a70107a  and  a70104a );
 a70109a <=( a70108a  and  a70101a );
 a70113a <=( A268  and  A267 );
 a70114a <=( A266  and  a70113a );
 a70117a <=( (not A299)  and  A298 );
 a70120a <=( A301  and  A300 );
 a70121a <=( a70120a  and  a70117a );
 a70122a <=( a70121a  and  a70114a );
 a70126a <=( A199  and  (not A168) );
 a70127a <=( A169  and  a70126a );
 a70130a <=( A201  and  (not A200) );
 a70133a <=( (not A265)  and  A202 );
 a70134a <=( a70133a  and  a70130a );
 a70135a <=( a70134a  and  a70127a );
 a70139a <=( A268  and  A267 );
 a70140a <=( A266  and  a70139a );
 a70143a <=( (not A299)  and  A298 );
 a70146a <=( (not A302)  and  A300 );
 a70147a <=( a70146a  and  a70143a );
 a70148a <=( a70147a  and  a70140a );
 a70152a <=( A199  and  (not A168) );
 a70153a <=( A169  and  a70152a );
 a70156a <=( A201  and  (not A200) );
 a70159a <=( (not A265)  and  A202 );
 a70160a <=( a70159a  and  a70156a );
 a70161a <=( a70160a  and  a70153a );
 a70165a <=( A268  and  A267 );
 a70166a <=( A266  and  a70165a );
 a70169a <=( A299  and  (not A298) );
 a70172a <=( A301  and  A300 );
 a70173a <=( a70172a  and  a70169a );
 a70174a <=( a70173a  and  a70166a );
 a70178a <=( A199  and  (not A168) );
 a70179a <=( A169  and  a70178a );
 a70182a <=( A201  and  (not A200) );
 a70185a <=( (not A265)  and  A202 );
 a70186a <=( a70185a  and  a70182a );
 a70187a <=( a70186a  and  a70179a );
 a70191a <=( A268  and  A267 );
 a70192a <=( A266  and  a70191a );
 a70195a <=( A299  and  (not A298) );
 a70198a <=( (not A302)  and  A300 );
 a70199a <=( a70198a  and  a70195a );
 a70200a <=( a70199a  and  a70192a );
 a70204a <=( A199  and  (not A168) );
 a70205a <=( A169  and  a70204a );
 a70208a <=( A201  and  (not A200) );
 a70211a <=( (not A265)  and  A202 );
 a70212a <=( a70211a  and  a70208a );
 a70213a <=( a70212a  and  a70205a );
 a70217a <=( (not A269)  and  A267 );
 a70218a <=( A266  and  a70217a );
 a70221a <=( (not A299)  and  A298 );
 a70224a <=( A301  and  A300 );
 a70225a <=( a70224a  and  a70221a );
 a70226a <=( a70225a  and  a70218a );
 a70230a <=( A199  and  (not A168) );
 a70231a <=( A169  and  a70230a );
 a70234a <=( A201  and  (not A200) );
 a70237a <=( (not A265)  and  A202 );
 a70238a <=( a70237a  and  a70234a );
 a70239a <=( a70238a  and  a70231a );
 a70243a <=( (not A269)  and  A267 );
 a70244a <=( A266  and  a70243a );
 a70247a <=( (not A299)  and  A298 );
 a70250a <=( (not A302)  and  A300 );
 a70251a <=( a70250a  and  a70247a );
 a70252a <=( a70251a  and  a70244a );
 a70256a <=( A199  and  (not A168) );
 a70257a <=( A169  and  a70256a );
 a70260a <=( A201  and  (not A200) );
 a70263a <=( (not A265)  and  A202 );
 a70264a <=( a70263a  and  a70260a );
 a70265a <=( a70264a  and  a70257a );
 a70269a <=( (not A269)  and  A267 );
 a70270a <=( A266  and  a70269a );
 a70273a <=( A299  and  (not A298) );
 a70276a <=( A301  and  A300 );
 a70277a <=( a70276a  and  a70273a );
 a70278a <=( a70277a  and  a70270a );
 a70282a <=( A199  and  (not A168) );
 a70283a <=( A169  and  a70282a );
 a70286a <=( A201  and  (not A200) );
 a70289a <=( (not A265)  and  A202 );
 a70290a <=( a70289a  and  a70286a );
 a70291a <=( a70290a  and  a70283a );
 a70295a <=( (not A269)  and  A267 );
 a70296a <=( A266  and  a70295a );
 a70299a <=( A299  and  (not A298) );
 a70302a <=( (not A302)  and  A300 );
 a70303a <=( a70302a  and  a70299a );
 a70304a <=( a70303a  and  a70296a );
 a70308a <=( A199  and  (not A168) );
 a70309a <=( A169  and  a70308a );
 a70312a <=( A201  and  (not A200) );
 a70315a <=( A265  and  A202 );
 a70316a <=( a70315a  and  a70312a );
 a70317a <=( a70316a  and  a70309a );
 a70321a <=( A268  and  A267 );
 a70322a <=( (not A266)  and  a70321a );
 a70325a <=( (not A299)  and  A298 );
 a70328a <=( A301  and  A300 );
 a70329a <=( a70328a  and  a70325a );
 a70330a <=( a70329a  and  a70322a );
 a70334a <=( A199  and  (not A168) );
 a70335a <=( A169  and  a70334a );
 a70338a <=( A201  and  (not A200) );
 a70341a <=( A265  and  A202 );
 a70342a <=( a70341a  and  a70338a );
 a70343a <=( a70342a  and  a70335a );
 a70347a <=( A268  and  A267 );
 a70348a <=( (not A266)  and  a70347a );
 a70351a <=( (not A299)  and  A298 );
 a70354a <=( (not A302)  and  A300 );
 a70355a <=( a70354a  and  a70351a );
 a70356a <=( a70355a  and  a70348a );
 a70360a <=( A199  and  (not A168) );
 a70361a <=( A169  and  a70360a );
 a70364a <=( A201  and  (not A200) );
 a70367a <=( A265  and  A202 );
 a70368a <=( a70367a  and  a70364a );
 a70369a <=( a70368a  and  a70361a );
 a70373a <=( A268  and  A267 );
 a70374a <=( (not A266)  and  a70373a );
 a70377a <=( A299  and  (not A298) );
 a70380a <=( A301  and  A300 );
 a70381a <=( a70380a  and  a70377a );
 a70382a <=( a70381a  and  a70374a );
 a70386a <=( A199  and  (not A168) );
 a70387a <=( A169  and  a70386a );
 a70390a <=( A201  and  (not A200) );
 a70393a <=( A265  and  A202 );
 a70394a <=( a70393a  and  a70390a );
 a70395a <=( a70394a  and  a70387a );
 a70399a <=( A268  and  A267 );
 a70400a <=( (not A266)  and  a70399a );
 a70403a <=( A299  and  (not A298) );
 a70406a <=( (not A302)  and  A300 );
 a70407a <=( a70406a  and  a70403a );
 a70408a <=( a70407a  and  a70400a );
 a70412a <=( A199  and  (not A168) );
 a70413a <=( A169  and  a70412a );
 a70416a <=( A201  and  (not A200) );
 a70419a <=( A265  and  A202 );
 a70420a <=( a70419a  and  a70416a );
 a70421a <=( a70420a  and  a70413a );
 a70425a <=( (not A269)  and  A267 );
 a70426a <=( (not A266)  and  a70425a );
 a70429a <=( (not A299)  and  A298 );
 a70432a <=( A301  and  A300 );
 a70433a <=( a70432a  and  a70429a );
 a70434a <=( a70433a  and  a70426a );
 a70438a <=( A199  and  (not A168) );
 a70439a <=( A169  and  a70438a );
 a70442a <=( A201  and  (not A200) );
 a70445a <=( A265  and  A202 );
 a70446a <=( a70445a  and  a70442a );
 a70447a <=( a70446a  and  a70439a );
 a70451a <=( (not A269)  and  A267 );
 a70452a <=( (not A266)  and  a70451a );
 a70455a <=( (not A299)  and  A298 );
 a70458a <=( (not A302)  and  A300 );
 a70459a <=( a70458a  and  a70455a );
 a70460a <=( a70459a  and  a70452a );
 a70464a <=( A199  and  (not A168) );
 a70465a <=( A169  and  a70464a );
 a70468a <=( A201  and  (not A200) );
 a70471a <=( A265  and  A202 );
 a70472a <=( a70471a  and  a70468a );
 a70473a <=( a70472a  and  a70465a );
 a70477a <=( (not A269)  and  A267 );
 a70478a <=( (not A266)  and  a70477a );
 a70481a <=( A299  and  (not A298) );
 a70484a <=( A301  and  A300 );
 a70485a <=( a70484a  and  a70481a );
 a70486a <=( a70485a  and  a70478a );
 a70490a <=( A199  and  (not A168) );
 a70491a <=( A169  and  a70490a );
 a70494a <=( A201  and  (not A200) );
 a70497a <=( A265  and  A202 );
 a70498a <=( a70497a  and  a70494a );
 a70499a <=( a70498a  and  a70491a );
 a70503a <=( (not A269)  and  A267 );
 a70504a <=( (not A266)  and  a70503a );
 a70507a <=( A299  and  (not A298) );
 a70510a <=( (not A302)  and  A300 );
 a70511a <=( a70510a  and  a70507a );
 a70512a <=( a70511a  and  a70504a );
 a70516a <=( A199  and  (not A168) );
 a70517a <=( A169  and  a70516a );
 a70520a <=( A201  and  (not A200) );
 a70523a <=( (not A265)  and  (not A203) );
 a70524a <=( a70523a  and  a70520a );
 a70525a <=( a70524a  and  a70517a );
 a70529a <=( A268  and  A267 );
 a70530a <=( A266  and  a70529a );
 a70533a <=( (not A299)  and  A298 );
 a70536a <=( A301  and  A300 );
 a70537a <=( a70536a  and  a70533a );
 a70538a <=( a70537a  and  a70530a );
 a70542a <=( A199  and  (not A168) );
 a70543a <=( A169  and  a70542a );
 a70546a <=( A201  and  (not A200) );
 a70549a <=( (not A265)  and  (not A203) );
 a70550a <=( a70549a  and  a70546a );
 a70551a <=( a70550a  and  a70543a );
 a70555a <=( A268  and  A267 );
 a70556a <=( A266  and  a70555a );
 a70559a <=( (not A299)  and  A298 );
 a70562a <=( (not A302)  and  A300 );
 a70563a <=( a70562a  and  a70559a );
 a70564a <=( a70563a  and  a70556a );
 a70568a <=( A199  and  (not A168) );
 a70569a <=( A169  and  a70568a );
 a70572a <=( A201  and  (not A200) );
 a70575a <=( (not A265)  and  (not A203) );
 a70576a <=( a70575a  and  a70572a );
 a70577a <=( a70576a  and  a70569a );
 a70581a <=( A268  and  A267 );
 a70582a <=( A266  and  a70581a );
 a70585a <=( A299  and  (not A298) );
 a70588a <=( A301  and  A300 );
 a70589a <=( a70588a  and  a70585a );
 a70590a <=( a70589a  and  a70582a );
 a70594a <=( A199  and  (not A168) );
 a70595a <=( A169  and  a70594a );
 a70598a <=( A201  and  (not A200) );
 a70601a <=( (not A265)  and  (not A203) );
 a70602a <=( a70601a  and  a70598a );
 a70603a <=( a70602a  and  a70595a );
 a70607a <=( A268  and  A267 );
 a70608a <=( A266  and  a70607a );
 a70611a <=( A299  and  (not A298) );
 a70614a <=( (not A302)  and  A300 );
 a70615a <=( a70614a  and  a70611a );
 a70616a <=( a70615a  and  a70608a );
 a70620a <=( A199  and  (not A168) );
 a70621a <=( A169  and  a70620a );
 a70624a <=( A201  and  (not A200) );
 a70627a <=( (not A265)  and  (not A203) );
 a70628a <=( a70627a  and  a70624a );
 a70629a <=( a70628a  and  a70621a );
 a70633a <=( (not A269)  and  A267 );
 a70634a <=( A266  and  a70633a );
 a70637a <=( (not A299)  and  A298 );
 a70640a <=( A301  and  A300 );
 a70641a <=( a70640a  and  a70637a );
 a70642a <=( a70641a  and  a70634a );
 a70646a <=( A199  and  (not A168) );
 a70647a <=( A169  and  a70646a );
 a70650a <=( A201  and  (not A200) );
 a70653a <=( (not A265)  and  (not A203) );
 a70654a <=( a70653a  and  a70650a );
 a70655a <=( a70654a  and  a70647a );
 a70659a <=( (not A269)  and  A267 );
 a70660a <=( A266  and  a70659a );
 a70663a <=( (not A299)  and  A298 );
 a70666a <=( (not A302)  and  A300 );
 a70667a <=( a70666a  and  a70663a );
 a70668a <=( a70667a  and  a70660a );
 a70672a <=( A199  and  (not A168) );
 a70673a <=( A169  and  a70672a );
 a70676a <=( A201  and  (not A200) );
 a70679a <=( (not A265)  and  (not A203) );
 a70680a <=( a70679a  and  a70676a );
 a70681a <=( a70680a  and  a70673a );
 a70685a <=( (not A269)  and  A267 );
 a70686a <=( A266  and  a70685a );
 a70689a <=( A299  and  (not A298) );
 a70692a <=( A301  and  A300 );
 a70693a <=( a70692a  and  a70689a );
 a70694a <=( a70693a  and  a70686a );
 a70698a <=( A199  and  (not A168) );
 a70699a <=( A169  and  a70698a );
 a70702a <=( A201  and  (not A200) );
 a70705a <=( (not A265)  and  (not A203) );
 a70706a <=( a70705a  and  a70702a );
 a70707a <=( a70706a  and  a70699a );
 a70711a <=( (not A269)  and  A267 );
 a70712a <=( A266  and  a70711a );
 a70715a <=( A299  and  (not A298) );
 a70718a <=( (not A302)  and  A300 );
 a70719a <=( a70718a  and  a70715a );
 a70720a <=( a70719a  and  a70712a );
 a70724a <=( A199  and  (not A168) );
 a70725a <=( A169  and  a70724a );
 a70728a <=( A201  and  (not A200) );
 a70731a <=( A265  and  (not A203) );
 a70732a <=( a70731a  and  a70728a );
 a70733a <=( a70732a  and  a70725a );
 a70737a <=( A268  and  A267 );
 a70738a <=( (not A266)  and  a70737a );
 a70741a <=( (not A299)  and  A298 );
 a70744a <=( A301  and  A300 );
 a70745a <=( a70744a  and  a70741a );
 a70746a <=( a70745a  and  a70738a );
 a70750a <=( A199  and  (not A168) );
 a70751a <=( A169  and  a70750a );
 a70754a <=( A201  and  (not A200) );
 a70757a <=( A265  and  (not A203) );
 a70758a <=( a70757a  and  a70754a );
 a70759a <=( a70758a  and  a70751a );
 a70763a <=( A268  and  A267 );
 a70764a <=( (not A266)  and  a70763a );
 a70767a <=( (not A299)  and  A298 );
 a70770a <=( (not A302)  and  A300 );
 a70771a <=( a70770a  and  a70767a );
 a70772a <=( a70771a  and  a70764a );
 a70776a <=( A199  and  (not A168) );
 a70777a <=( A169  and  a70776a );
 a70780a <=( A201  and  (not A200) );
 a70783a <=( A265  and  (not A203) );
 a70784a <=( a70783a  and  a70780a );
 a70785a <=( a70784a  and  a70777a );
 a70789a <=( A268  and  A267 );
 a70790a <=( (not A266)  and  a70789a );
 a70793a <=( A299  and  (not A298) );
 a70796a <=( A301  and  A300 );
 a70797a <=( a70796a  and  a70793a );
 a70798a <=( a70797a  and  a70790a );
 a70802a <=( A199  and  (not A168) );
 a70803a <=( A169  and  a70802a );
 a70806a <=( A201  and  (not A200) );
 a70809a <=( A265  and  (not A203) );
 a70810a <=( a70809a  and  a70806a );
 a70811a <=( a70810a  and  a70803a );
 a70815a <=( A268  and  A267 );
 a70816a <=( (not A266)  and  a70815a );
 a70819a <=( A299  and  (not A298) );
 a70822a <=( (not A302)  and  A300 );
 a70823a <=( a70822a  and  a70819a );
 a70824a <=( a70823a  and  a70816a );
 a70828a <=( A199  and  (not A168) );
 a70829a <=( A169  and  a70828a );
 a70832a <=( A201  and  (not A200) );
 a70835a <=( A265  and  (not A203) );
 a70836a <=( a70835a  and  a70832a );
 a70837a <=( a70836a  and  a70829a );
 a70841a <=( (not A269)  and  A267 );
 a70842a <=( (not A266)  and  a70841a );
 a70845a <=( (not A299)  and  A298 );
 a70848a <=( A301  and  A300 );
 a70849a <=( a70848a  and  a70845a );
 a70850a <=( a70849a  and  a70842a );
 a70854a <=( A199  and  (not A168) );
 a70855a <=( A169  and  a70854a );
 a70858a <=( A201  and  (not A200) );
 a70861a <=( A265  and  (not A203) );
 a70862a <=( a70861a  and  a70858a );
 a70863a <=( a70862a  and  a70855a );
 a70867a <=( (not A269)  and  A267 );
 a70868a <=( (not A266)  and  a70867a );
 a70871a <=( (not A299)  and  A298 );
 a70874a <=( (not A302)  and  A300 );
 a70875a <=( a70874a  and  a70871a );
 a70876a <=( a70875a  and  a70868a );
 a70880a <=( A199  and  (not A168) );
 a70881a <=( A169  and  a70880a );
 a70884a <=( A201  and  (not A200) );
 a70887a <=( A265  and  (not A203) );
 a70888a <=( a70887a  and  a70884a );
 a70889a <=( a70888a  and  a70881a );
 a70893a <=( (not A269)  and  A267 );
 a70894a <=( (not A266)  and  a70893a );
 a70897a <=( A299  and  (not A298) );
 a70900a <=( A301  and  A300 );
 a70901a <=( a70900a  and  a70897a );
 a70902a <=( a70901a  and  a70894a );
 a70906a <=( A199  and  (not A168) );
 a70907a <=( A169  and  a70906a );
 a70910a <=( A201  and  (not A200) );
 a70913a <=( A265  and  (not A203) );
 a70914a <=( a70913a  and  a70910a );
 a70915a <=( a70914a  and  a70907a );
 a70919a <=( (not A269)  and  A267 );
 a70920a <=( (not A266)  and  a70919a );
 a70923a <=( A299  and  (not A298) );
 a70926a <=( (not A302)  and  A300 );
 a70927a <=( a70926a  and  a70923a );
 a70928a <=( a70927a  and  a70920a );
 a70932a <=( A168  and  (not A169) );
 a70933a <=( (not A170)  and  a70932a );
 a70936a <=( A200  and  (not A199) );
 a70939a <=( (not A202)  and  (not A201) );
 a70940a <=( a70939a  and  a70936a );
 a70941a <=( a70940a  and  a70933a );
 a70945a <=( (not A268)  and  A267 );
 a70946a <=( A203  and  a70945a );
 a70949a <=( A300  and  A269 );
 a70952a <=( A302  and  (not A301) );
 a70953a <=( a70952a  and  a70949a );
 a70954a <=( a70953a  and  a70946a );
 a70958a <=( A168  and  (not A169) );
 a70959a <=( (not A170)  and  a70958a );
 a70962a <=( (not A200)  and  A199 );
 a70965a <=( (not A202)  and  (not A201) );
 a70966a <=( a70965a  and  a70962a );
 a70967a <=( a70966a  and  a70959a );
 a70971a <=( (not A268)  and  A267 );
 a70972a <=( A203  and  a70971a );
 a70975a <=( A300  and  A269 );
 a70978a <=( A302  and  (not A301) );
 a70979a <=( a70978a  and  a70975a );
 a70980a <=( a70979a  and  a70972a );
 a70984a <=( (not A168)  and  (not A169) );
 a70985a <=( (not A170)  and  a70984a );
 a70988a <=( (not A166)  and  A167 );
 a70991a <=( (not A202)  and  A201 );
 a70992a <=( a70991a  and  a70988a );
 a70993a <=( a70992a  and  a70985a );
 a70997a <=( A268  and  (not A267) );
 a70998a <=( A203  and  a70997a );
 a71001a <=( (not A299)  and  A298 );
 a71004a <=( A301  and  A300 );
 a71005a <=( a71004a  and  a71001a );
 a71006a <=( a71005a  and  a70998a );
 a71010a <=( (not A168)  and  (not A169) );
 a71011a <=( (not A170)  and  a71010a );
 a71014a <=( (not A166)  and  A167 );
 a71017a <=( (not A202)  and  A201 );
 a71018a <=( a71017a  and  a71014a );
 a71019a <=( a71018a  and  a71011a );
 a71023a <=( A268  and  (not A267) );
 a71024a <=( A203  and  a71023a );
 a71027a <=( (not A299)  and  A298 );
 a71030a <=( (not A302)  and  A300 );
 a71031a <=( a71030a  and  a71027a );
 a71032a <=( a71031a  and  a71024a );
 a71036a <=( (not A168)  and  (not A169) );
 a71037a <=( (not A170)  and  a71036a );
 a71040a <=( (not A166)  and  A167 );
 a71043a <=( (not A202)  and  A201 );
 a71044a <=( a71043a  and  a71040a );
 a71045a <=( a71044a  and  a71037a );
 a71049a <=( A268  and  (not A267) );
 a71050a <=( A203  and  a71049a );
 a71053a <=( A299  and  (not A298) );
 a71056a <=( A301  and  A300 );
 a71057a <=( a71056a  and  a71053a );
 a71058a <=( a71057a  and  a71050a );
 a71062a <=( (not A168)  and  (not A169) );
 a71063a <=( (not A170)  and  a71062a );
 a71066a <=( (not A166)  and  A167 );
 a71069a <=( (not A202)  and  A201 );
 a71070a <=( a71069a  and  a71066a );
 a71071a <=( a71070a  and  a71063a );
 a71075a <=( A268  and  (not A267) );
 a71076a <=( A203  and  a71075a );
 a71079a <=( A299  and  (not A298) );
 a71082a <=( (not A302)  and  A300 );
 a71083a <=( a71082a  and  a71079a );
 a71084a <=( a71083a  and  a71076a );
 a71088a <=( (not A168)  and  (not A169) );
 a71089a <=( (not A170)  and  a71088a );
 a71092a <=( (not A166)  and  A167 );
 a71095a <=( (not A202)  and  A201 );
 a71096a <=( a71095a  and  a71092a );
 a71097a <=( a71096a  and  a71089a );
 a71101a <=( (not A269)  and  (not A267) );
 a71102a <=( A203  and  a71101a );
 a71105a <=( (not A299)  and  A298 );
 a71108a <=( A301  and  A300 );
 a71109a <=( a71108a  and  a71105a );
 a71110a <=( a71109a  and  a71102a );
 a71114a <=( (not A168)  and  (not A169) );
 a71115a <=( (not A170)  and  a71114a );
 a71118a <=( (not A166)  and  A167 );
 a71121a <=( (not A202)  and  A201 );
 a71122a <=( a71121a  and  a71118a );
 a71123a <=( a71122a  and  a71115a );
 a71127a <=( (not A269)  and  (not A267) );
 a71128a <=( A203  and  a71127a );
 a71131a <=( (not A299)  and  A298 );
 a71134a <=( (not A302)  and  A300 );
 a71135a <=( a71134a  and  a71131a );
 a71136a <=( a71135a  and  a71128a );
 a71140a <=( (not A168)  and  (not A169) );
 a71141a <=( (not A170)  and  a71140a );
 a71144a <=( (not A166)  and  A167 );
 a71147a <=( (not A202)  and  A201 );
 a71148a <=( a71147a  and  a71144a );
 a71149a <=( a71148a  and  a71141a );
 a71153a <=( (not A269)  and  (not A267) );
 a71154a <=( A203  and  a71153a );
 a71157a <=( A299  and  (not A298) );
 a71160a <=( A301  and  A300 );
 a71161a <=( a71160a  and  a71157a );
 a71162a <=( a71161a  and  a71154a );
 a71166a <=( (not A168)  and  (not A169) );
 a71167a <=( (not A170)  and  a71166a );
 a71170a <=( (not A166)  and  A167 );
 a71173a <=( (not A202)  and  A201 );
 a71174a <=( a71173a  and  a71170a );
 a71175a <=( a71174a  and  a71167a );
 a71179a <=( (not A269)  and  (not A267) );
 a71180a <=( A203  and  a71179a );
 a71183a <=( A299  and  (not A298) );
 a71186a <=( (not A302)  and  A300 );
 a71187a <=( a71186a  and  a71183a );
 a71188a <=( a71187a  and  a71180a );
 a71192a <=( (not A168)  and  (not A169) );
 a71193a <=( (not A170)  and  a71192a );
 a71196a <=( (not A166)  and  A167 );
 a71199a <=( (not A202)  and  A201 );
 a71200a <=( a71199a  and  a71196a );
 a71201a <=( a71200a  and  a71193a );
 a71205a <=( A266  and  A265 );
 a71206a <=( A203  and  a71205a );
 a71209a <=( (not A299)  and  A298 );
 a71212a <=( A301  and  A300 );
 a71213a <=( a71212a  and  a71209a );
 a71214a <=( a71213a  and  a71206a );
 a71218a <=( (not A168)  and  (not A169) );
 a71219a <=( (not A170)  and  a71218a );
 a71222a <=( (not A166)  and  A167 );
 a71225a <=( (not A202)  and  A201 );
 a71226a <=( a71225a  and  a71222a );
 a71227a <=( a71226a  and  a71219a );
 a71231a <=( A266  and  A265 );
 a71232a <=( A203  and  a71231a );
 a71235a <=( (not A299)  and  A298 );
 a71238a <=( (not A302)  and  A300 );
 a71239a <=( a71238a  and  a71235a );
 a71240a <=( a71239a  and  a71232a );
 a71244a <=( (not A168)  and  (not A169) );
 a71245a <=( (not A170)  and  a71244a );
 a71248a <=( (not A166)  and  A167 );
 a71251a <=( (not A202)  and  A201 );
 a71252a <=( a71251a  and  a71248a );
 a71253a <=( a71252a  and  a71245a );
 a71257a <=( A266  and  A265 );
 a71258a <=( A203  and  a71257a );
 a71261a <=( A299  and  (not A298) );
 a71264a <=( A301  and  A300 );
 a71265a <=( a71264a  and  a71261a );
 a71266a <=( a71265a  and  a71258a );
 a71270a <=( (not A168)  and  (not A169) );
 a71271a <=( (not A170)  and  a71270a );
 a71274a <=( (not A166)  and  A167 );
 a71277a <=( (not A202)  and  A201 );
 a71278a <=( a71277a  and  a71274a );
 a71279a <=( a71278a  and  a71271a );
 a71283a <=( A266  and  A265 );
 a71284a <=( A203  and  a71283a );
 a71287a <=( A299  and  (not A298) );
 a71290a <=( (not A302)  and  A300 );
 a71291a <=( a71290a  and  a71287a );
 a71292a <=( a71291a  and  a71284a );
 a71296a <=( (not A168)  and  (not A169) );
 a71297a <=( (not A170)  and  a71296a );
 a71300a <=( (not A166)  and  A167 );
 a71303a <=( (not A202)  and  A201 );
 a71304a <=( a71303a  and  a71300a );
 a71305a <=( a71304a  and  a71297a );
 a71309a <=( A266  and  (not A265) );
 a71310a <=( A203  and  a71309a );
 a71313a <=( A268  and  A267 );
 a71316a <=( A301  and  (not A300) );
 a71317a <=( a71316a  and  a71313a );
 a71318a <=( a71317a  and  a71310a );
 a71322a <=( (not A168)  and  (not A169) );
 a71323a <=( (not A170)  and  a71322a );
 a71326a <=( (not A166)  and  A167 );
 a71329a <=( (not A202)  and  A201 );
 a71330a <=( a71329a  and  a71326a );
 a71331a <=( a71330a  and  a71323a );
 a71335a <=( A266  and  (not A265) );
 a71336a <=( A203  and  a71335a );
 a71339a <=( A268  and  A267 );
 a71342a <=( (not A302)  and  (not A300) );
 a71343a <=( a71342a  and  a71339a );
 a71344a <=( a71343a  and  a71336a );
 a71348a <=( (not A168)  and  (not A169) );
 a71349a <=( (not A170)  and  a71348a );
 a71352a <=( (not A166)  and  A167 );
 a71355a <=( (not A202)  and  A201 );
 a71356a <=( a71355a  and  a71352a );
 a71357a <=( a71356a  and  a71349a );
 a71361a <=( A266  and  (not A265) );
 a71362a <=( A203  and  a71361a );
 a71365a <=( A268  and  A267 );
 a71368a <=( A299  and  A298 );
 a71369a <=( a71368a  and  a71365a );
 a71370a <=( a71369a  and  a71362a );
 a71374a <=( (not A168)  and  (not A169) );
 a71375a <=( (not A170)  and  a71374a );
 a71378a <=( (not A166)  and  A167 );
 a71381a <=( (not A202)  and  A201 );
 a71382a <=( a71381a  and  a71378a );
 a71383a <=( a71382a  and  a71375a );
 a71387a <=( A266  and  (not A265) );
 a71388a <=( A203  and  a71387a );
 a71391a <=( A268  and  A267 );
 a71394a <=( (not A299)  and  (not A298) );
 a71395a <=( a71394a  and  a71391a );
 a71396a <=( a71395a  and  a71388a );
 a71400a <=( (not A168)  and  (not A169) );
 a71401a <=( (not A170)  and  a71400a );
 a71404a <=( (not A166)  and  A167 );
 a71407a <=( (not A202)  and  A201 );
 a71408a <=( a71407a  and  a71404a );
 a71409a <=( a71408a  and  a71401a );
 a71413a <=( A266  and  (not A265) );
 a71414a <=( A203  and  a71413a );
 a71417a <=( (not A269)  and  A267 );
 a71420a <=( A301  and  (not A300) );
 a71421a <=( a71420a  and  a71417a );
 a71422a <=( a71421a  and  a71414a );
 a71426a <=( (not A168)  and  (not A169) );
 a71427a <=( (not A170)  and  a71426a );
 a71430a <=( (not A166)  and  A167 );
 a71433a <=( (not A202)  and  A201 );
 a71434a <=( a71433a  and  a71430a );
 a71435a <=( a71434a  and  a71427a );
 a71439a <=( A266  and  (not A265) );
 a71440a <=( A203  and  a71439a );
 a71443a <=( (not A269)  and  A267 );
 a71446a <=( (not A302)  and  (not A300) );
 a71447a <=( a71446a  and  a71443a );
 a71448a <=( a71447a  and  a71440a );
 a71452a <=( (not A168)  and  (not A169) );
 a71453a <=( (not A170)  and  a71452a );
 a71456a <=( (not A166)  and  A167 );
 a71459a <=( (not A202)  and  A201 );
 a71460a <=( a71459a  and  a71456a );
 a71461a <=( a71460a  and  a71453a );
 a71465a <=( A266  and  (not A265) );
 a71466a <=( A203  and  a71465a );
 a71469a <=( (not A269)  and  A267 );
 a71472a <=( A299  and  A298 );
 a71473a <=( a71472a  and  a71469a );
 a71474a <=( a71473a  and  a71466a );
 a71478a <=( (not A168)  and  (not A169) );
 a71479a <=( (not A170)  and  a71478a );
 a71482a <=( (not A166)  and  A167 );
 a71485a <=( (not A202)  and  A201 );
 a71486a <=( a71485a  and  a71482a );
 a71487a <=( a71486a  and  a71479a );
 a71491a <=( A266  and  (not A265) );
 a71492a <=( A203  and  a71491a );
 a71495a <=( (not A269)  and  A267 );
 a71498a <=( (not A299)  and  (not A298) );
 a71499a <=( a71498a  and  a71495a );
 a71500a <=( a71499a  and  a71492a );
 a71504a <=( (not A168)  and  (not A169) );
 a71505a <=( (not A170)  and  a71504a );
 a71508a <=( (not A166)  and  A167 );
 a71511a <=( (not A202)  and  A201 );
 a71512a <=( a71511a  and  a71508a );
 a71513a <=( a71512a  and  a71505a );
 a71517a <=( (not A266)  and  A265 );
 a71518a <=( A203  and  a71517a );
 a71521a <=( A268  and  A267 );
 a71524a <=( A301  and  (not A300) );
 a71525a <=( a71524a  and  a71521a );
 a71526a <=( a71525a  and  a71518a );
 a71530a <=( (not A168)  and  (not A169) );
 a71531a <=( (not A170)  and  a71530a );
 a71534a <=( (not A166)  and  A167 );
 a71537a <=( (not A202)  and  A201 );
 a71538a <=( a71537a  and  a71534a );
 a71539a <=( a71538a  and  a71531a );
 a71543a <=( (not A266)  and  A265 );
 a71544a <=( A203  and  a71543a );
 a71547a <=( A268  and  A267 );
 a71550a <=( (not A302)  and  (not A300) );
 a71551a <=( a71550a  and  a71547a );
 a71552a <=( a71551a  and  a71544a );
 a71556a <=( (not A168)  and  (not A169) );
 a71557a <=( (not A170)  and  a71556a );
 a71560a <=( (not A166)  and  A167 );
 a71563a <=( (not A202)  and  A201 );
 a71564a <=( a71563a  and  a71560a );
 a71565a <=( a71564a  and  a71557a );
 a71569a <=( (not A266)  and  A265 );
 a71570a <=( A203  and  a71569a );
 a71573a <=( A268  and  A267 );
 a71576a <=( A299  and  A298 );
 a71577a <=( a71576a  and  a71573a );
 a71578a <=( a71577a  and  a71570a );
 a71582a <=( (not A168)  and  (not A169) );
 a71583a <=( (not A170)  and  a71582a );
 a71586a <=( (not A166)  and  A167 );
 a71589a <=( (not A202)  and  A201 );
 a71590a <=( a71589a  and  a71586a );
 a71591a <=( a71590a  and  a71583a );
 a71595a <=( (not A266)  and  A265 );
 a71596a <=( A203  and  a71595a );
 a71599a <=( A268  and  A267 );
 a71602a <=( (not A299)  and  (not A298) );
 a71603a <=( a71602a  and  a71599a );
 a71604a <=( a71603a  and  a71596a );
 a71608a <=( (not A168)  and  (not A169) );
 a71609a <=( (not A170)  and  a71608a );
 a71612a <=( (not A166)  and  A167 );
 a71615a <=( (not A202)  and  A201 );
 a71616a <=( a71615a  and  a71612a );
 a71617a <=( a71616a  and  a71609a );
 a71621a <=( (not A266)  and  A265 );
 a71622a <=( A203  and  a71621a );
 a71625a <=( (not A269)  and  A267 );
 a71628a <=( A301  and  (not A300) );
 a71629a <=( a71628a  and  a71625a );
 a71630a <=( a71629a  and  a71622a );
 a71634a <=( (not A168)  and  (not A169) );
 a71635a <=( (not A170)  and  a71634a );
 a71638a <=( (not A166)  and  A167 );
 a71641a <=( (not A202)  and  A201 );
 a71642a <=( a71641a  and  a71638a );
 a71643a <=( a71642a  and  a71635a );
 a71647a <=( (not A266)  and  A265 );
 a71648a <=( A203  and  a71647a );
 a71651a <=( (not A269)  and  A267 );
 a71654a <=( (not A302)  and  (not A300) );
 a71655a <=( a71654a  and  a71651a );
 a71656a <=( a71655a  and  a71648a );
 a71660a <=( (not A168)  and  (not A169) );
 a71661a <=( (not A170)  and  a71660a );
 a71664a <=( (not A166)  and  A167 );
 a71667a <=( (not A202)  and  A201 );
 a71668a <=( a71667a  and  a71664a );
 a71669a <=( a71668a  and  a71661a );
 a71673a <=( (not A266)  and  A265 );
 a71674a <=( A203  and  a71673a );
 a71677a <=( (not A269)  and  A267 );
 a71680a <=( A299  and  A298 );
 a71681a <=( a71680a  and  a71677a );
 a71682a <=( a71681a  and  a71674a );
 a71686a <=( (not A168)  and  (not A169) );
 a71687a <=( (not A170)  and  a71686a );
 a71690a <=( (not A166)  and  A167 );
 a71693a <=( (not A202)  and  A201 );
 a71694a <=( a71693a  and  a71690a );
 a71695a <=( a71694a  and  a71687a );
 a71699a <=( (not A266)  and  A265 );
 a71700a <=( A203  and  a71699a );
 a71703a <=( (not A269)  and  A267 );
 a71706a <=( (not A299)  and  (not A298) );
 a71707a <=( a71706a  and  a71703a );
 a71708a <=( a71707a  and  a71700a );
 a71712a <=( (not A168)  and  (not A169) );
 a71713a <=( (not A170)  and  a71712a );
 a71716a <=( (not A166)  and  A167 );
 a71719a <=( (not A202)  and  A201 );
 a71720a <=( a71719a  and  a71716a );
 a71721a <=( a71720a  and  a71713a );
 a71725a <=( (not A266)  and  (not A265) );
 a71726a <=( A203  and  a71725a );
 a71729a <=( (not A299)  and  A298 );
 a71732a <=( A301  and  A300 );
 a71733a <=( a71732a  and  a71729a );
 a71734a <=( a71733a  and  a71726a );
 a71738a <=( (not A168)  and  (not A169) );
 a71739a <=( (not A170)  and  a71738a );
 a71742a <=( (not A166)  and  A167 );
 a71745a <=( (not A202)  and  A201 );
 a71746a <=( a71745a  and  a71742a );
 a71747a <=( a71746a  and  a71739a );
 a71751a <=( (not A266)  and  (not A265) );
 a71752a <=( A203  and  a71751a );
 a71755a <=( (not A299)  and  A298 );
 a71758a <=( (not A302)  and  A300 );
 a71759a <=( a71758a  and  a71755a );
 a71760a <=( a71759a  and  a71752a );
 a71764a <=( (not A168)  and  (not A169) );
 a71765a <=( (not A170)  and  a71764a );
 a71768a <=( (not A166)  and  A167 );
 a71771a <=( (not A202)  and  A201 );
 a71772a <=( a71771a  and  a71768a );
 a71773a <=( a71772a  and  a71765a );
 a71777a <=( (not A266)  and  (not A265) );
 a71778a <=( A203  and  a71777a );
 a71781a <=( A299  and  (not A298) );
 a71784a <=( A301  and  A300 );
 a71785a <=( a71784a  and  a71781a );
 a71786a <=( a71785a  and  a71778a );
 a71790a <=( (not A168)  and  (not A169) );
 a71791a <=( (not A170)  and  a71790a );
 a71794a <=( (not A166)  and  A167 );
 a71797a <=( (not A202)  and  A201 );
 a71798a <=( a71797a  and  a71794a );
 a71799a <=( a71798a  and  a71791a );
 a71803a <=( (not A266)  and  (not A265) );
 a71804a <=( A203  and  a71803a );
 a71807a <=( A299  and  (not A298) );
 a71810a <=( (not A302)  and  A300 );
 a71811a <=( a71810a  and  a71807a );
 a71812a <=( a71811a  and  a71804a );
 a71816a <=( (not A168)  and  (not A169) );
 a71817a <=( (not A170)  and  a71816a );
 a71820a <=( (not A166)  and  A167 );
 a71823a <=( A202  and  (not A201) );
 a71824a <=( a71823a  and  a71820a );
 a71825a <=( a71824a  and  a71817a );
 a71829a <=( A269  and  (not A268) );
 a71830a <=( A267  and  a71829a );
 a71833a <=( (not A299)  and  A298 );
 a71836a <=( A301  and  A300 );
 a71837a <=( a71836a  and  a71833a );
 a71838a <=( a71837a  and  a71830a );
 a71842a <=( (not A168)  and  (not A169) );
 a71843a <=( (not A170)  and  a71842a );
 a71846a <=( (not A166)  and  A167 );
 a71849a <=( A202  and  (not A201) );
 a71850a <=( a71849a  and  a71846a );
 a71851a <=( a71850a  and  a71843a );
 a71855a <=( A269  and  (not A268) );
 a71856a <=( A267  and  a71855a );
 a71859a <=( (not A299)  and  A298 );
 a71862a <=( (not A302)  and  A300 );
 a71863a <=( a71862a  and  a71859a );
 a71864a <=( a71863a  and  a71856a );
 a71868a <=( (not A168)  and  (not A169) );
 a71869a <=( (not A170)  and  a71868a );
 a71872a <=( (not A166)  and  A167 );
 a71875a <=( A202  and  (not A201) );
 a71876a <=( a71875a  and  a71872a );
 a71877a <=( a71876a  and  a71869a );
 a71881a <=( A269  and  (not A268) );
 a71882a <=( A267  and  a71881a );
 a71885a <=( A299  and  (not A298) );
 a71888a <=( A301  and  A300 );
 a71889a <=( a71888a  and  a71885a );
 a71890a <=( a71889a  and  a71882a );
 a71894a <=( (not A168)  and  (not A169) );
 a71895a <=( (not A170)  and  a71894a );
 a71898a <=( (not A166)  and  A167 );
 a71901a <=( A202  and  (not A201) );
 a71902a <=( a71901a  and  a71898a );
 a71903a <=( a71902a  and  a71895a );
 a71907a <=( A269  and  (not A268) );
 a71908a <=( A267  and  a71907a );
 a71911a <=( A299  and  (not A298) );
 a71914a <=( (not A302)  and  A300 );
 a71915a <=( a71914a  and  a71911a );
 a71916a <=( a71915a  and  a71908a );
 a71920a <=( (not A168)  and  (not A169) );
 a71921a <=( (not A170)  and  a71920a );
 a71924a <=( (not A166)  and  A167 );
 a71927a <=( A202  and  (not A201) );
 a71928a <=( a71927a  and  a71924a );
 a71929a <=( a71928a  and  a71921a );
 a71933a <=( A298  and  A268 );
 a71934a <=( (not A267)  and  a71933a );
 a71937a <=( (not A300)  and  (not A299) );
 a71940a <=( A302  and  (not A301) );
 a71941a <=( a71940a  and  a71937a );
 a71942a <=( a71941a  and  a71934a );
 a71946a <=( (not A168)  and  (not A169) );
 a71947a <=( (not A170)  and  a71946a );
 a71950a <=( (not A166)  and  A167 );
 a71953a <=( A202  and  (not A201) );
 a71954a <=( a71953a  and  a71950a );
 a71955a <=( a71954a  and  a71947a );
 a71959a <=( (not A298)  and  A268 );
 a71960a <=( (not A267)  and  a71959a );
 a71963a <=( (not A300)  and  A299 );
 a71966a <=( A302  and  (not A301) );
 a71967a <=( a71966a  and  a71963a );
 a71968a <=( a71967a  and  a71960a );
 a71972a <=( (not A168)  and  (not A169) );
 a71973a <=( (not A170)  and  a71972a );
 a71976a <=( (not A166)  and  A167 );
 a71979a <=( A202  and  (not A201) );
 a71980a <=( a71979a  and  a71976a );
 a71981a <=( a71980a  and  a71973a );
 a71985a <=( A298  and  (not A269) );
 a71986a <=( (not A267)  and  a71985a );
 a71989a <=( (not A300)  and  (not A299) );
 a71992a <=( A302  and  (not A301) );
 a71993a <=( a71992a  and  a71989a );
 a71994a <=( a71993a  and  a71986a );
 a71998a <=( (not A168)  and  (not A169) );
 a71999a <=( (not A170)  and  a71998a );
 a72002a <=( (not A166)  and  A167 );
 a72005a <=( A202  and  (not A201) );
 a72006a <=( a72005a  and  a72002a );
 a72007a <=( a72006a  and  a71999a );
 a72011a <=( (not A298)  and  (not A269) );
 a72012a <=( (not A267)  and  a72011a );
 a72015a <=( (not A300)  and  A299 );
 a72018a <=( A302  and  (not A301) );
 a72019a <=( a72018a  and  a72015a );
 a72020a <=( a72019a  and  a72012a );
 a72024a <=( (not A168)  and  (not A169) );
 a72025a <=( (not A170)  and  a72024a );
 a72028a <=( (not A166)  and  A167 );
 a72031a <=( A202  and  (not A201) );
 a72032a <=( a72031a  and  a72028a );
 a72033a <=( a72032a  and  a72025a );
 a72037a <=( A298  and  A266 );
 a72038a <=( A265  and  a72037a );
 a72041a <=( (not A300)  and  (not A299) );
 a72044a <=( A302  and  (not A301) );
 a72045a <=( a72044a  and  a72041a );
 a72046a <=( a72045a  and  a72038a );
 a72050a <=( (not A168)  and  (not A169) );
 a72051a <=( (not A170)  and  a72050a );
 a72054a <=( (not A166)  and  A167 );
 a72057a <=( A202  and  (not A201) );
 a72058a <=( a72057a  and  a72054a );
 a72059a <=( a72058a  and  a72051a );
 a72063a <=( (not A298)  and  A266 );
 a72064a <=( A265  and  a72063a );
 a72067a <=( (not A300)  and  A299 );
 a72070a <=( A302  and  (not A301) );
 a72071a <=( a72070a  and  a72067a );
 a72072a <=( a72071a  and  a72064a );
 a72076a <=( (not A168)  and  (not A169) );
 a72077a <=( (not A170)  and  a72076a );
 a72080a <=( (not A166)  and  A167 );
 a72083a <=( A202  and  (not A201) );
 a72084a <=( a72083a  and  a72080a );
 a72085a <=( a72084a  and  a72077a );
 a72089a <=( A267  and  A266 );
 a72090a <=( (not A265)  and  a72089a );
 a72093a <=( A300  and  A268 );
 a72096a <=( A302  and  (not A301) );
 a72097a <=( a72096a  and  a72093a );
 a72098a <=( a72097a  and  a72090a );
 a72102a <=( (not A168)  and  (not A169) );
 a72103a <=( (not A170)  and  a72102a );
 a72106a <=( (not A166)  and  A167 );
 a72109a <=( A202  and  (not A201) );
 a72110a <=( a72109a  and  a72106a );
 a72111a <=( a72110a  and  a72103a );
 a72115a <=( A267  and  A266 );
 a72116a <=( (not A265)  and  a72115a );
 a72119a <=( A300  and  (not A269) );
 a72122a <=( A302  and  (not A301) );
 a72123a <=( a72122a  and  a72119a );
 a72124a <=( a72123a  and  a72116a );
 a72128a <=( (not A168)  and  (not A169) );
 a72129a <=( (not A170)  and  a72128a );
 a72132a <=( (not A166)  and  A167 );
 a72135a <=( A202  and  (not A201) );
 a72136a <=( a72135a  and  a72132a );
 a72137a <=( a72136a  and  a72129a );
 a72141a <=( (not A267)  and  A266 );
 a72142a <=( (not A265)  and  a72141a );
 a72145a <=( A269  and  (not A268) );
 a72148a <=( A301  and  (not A300) );
 a72149a <=( a72148a  and  a72145a );
 a72150a <=( a72149a  and  a72142a );
 a72154a <=( (not A168)  and  (not A169) );
 a72155a <=( (not A170)  and  a72154a );
 a72158a <=( (not A166)  and  A167 );
 a72161a <=( A202  and  (not A201) );
 a72162a <=( a72161a  and  a72158a );
 a72163a <=( a72162a  and  a72155a );
 a72167a <=( (not A267)  and  A266 );
 a72168a <=( (not A265)  and  a72167a );
 a72171a <=( A269  and  (not A268) );
 a72174a <=( (not A302)  and  (not A300) );
 a72175a <=( a72174a  and  a72171a );
 a72176a <=( a72175a  and  a72168a );
 a72180a <=( (not A168)  and  (not A169) );
 a72181a <=( (not A170)  and  a72180a );
 a72184a <=( (not A166)  and  A167 );
 a72187a <=( A202  and  (not A201) );
 a72188a <=( a72187a  and  a72184a );
 a72189a <=( a72188a  and  a72181a );
 a72193a <=( (not A267)  and  A266 );
 a72194a <=( (not A265)  and  a72193a );
 a72197a <=( A269  and  (not A268) );
 a72200a <=( A299  and  A298 );
 a72201a <=( a72200a  and  a72197a );
 a72202a <=( a72201a  and  a72194a );
 a72206a <=( (not A168)  and  (not A169) );
 a72207a <=( (not A170)  and  a72206a );
 a72210a <=( (not A166)  and  A167 );
 a72213a <=( A202  and  (not A201) );
 a72214a <=( a72213a  and  a72210a );
 a72215a <=( a72214a  and  a72207a );
 a72219a <=( (not A267)  and  A266 );
 a72220a <=( (not A265)  and  a72219a );
 a72223a <=( A269  and  (not A268) );
 a72226a <=( (not A299)  and  (not A298) );
 a72227a <=( a72226a  and  a72223a );
 a72228a <=( a72227a  and  a72220a );
 a72232a <=( (not A168)  and  (not A169) );
 a72233a <=( (not A170)  and  a72232a );
 a72236a <=( (not A166)  and  A167 );
 a72239a <=( A202  and  (not A201) );
 a72240a <=( a72239a  and  a72236a );
 a72241a <=( a72240a  and  a72233a );
 a72245a <=( A267  and  (not A266) );
 a72246a <=( A265  and  a72245a );
 a72249a <=( A300  and  A268 );
 a72252a <=( A302  and  (not A301) );
 a72253a <=( a72252a  and  a72249a );
 a72254a <=( a72253a  and  a72246a );
 a72258a <=( (not A168)  and  (not A169) );
 a72259a <=( (not A170)  and  a72258a );
 a72262a <=( (not A166)  and  A167 );
 a72265a <=( A202  and  (not A201) );
 a72266a <=( a72265a  and  a72262a );
 a72267a <=( a72266a  and  a72259a );
 a72271a <=( A267  and  (not A266) );
 a72272a <=( A265  and  a72271a );
 a72275a <=( A300  and  (not A269) );
 a72278a <=( A302  and  (not A301) );
 a72279a <=( a72278a  and  a72275a );
 a72280a <=( a72279a  and  a72272a );
 a72284a <=( (not A168)  and  (not A169) );
 a72285a <=( (not A170)  and  a72284a );
 a72288a <=( (not A166)  and  A167 );
 a72291a <=( A202  and  (not A201) );
 a72292a <=( a72291a  and  a72288a );
 a72293a <=( a72292a  and  a72285a );
 a72297a <=( (not A267)  and  (not A266) );
 a72298a <=( A265  and  a72297a );
 a72301a <=( A269  and  (not A268) );
 a72304a <=( A301  and  (not A300) );
 a72305a <=( a72304a  and  a72301a );
 a72306a <=( a72305a  and  a72298a );
 a72310a <=( (not A168)  and  (not A169) );
 a72311a <=( (not A170)  and  a72310a );
 a72314a <=( (not A166)  and  A167 );
 a72317a <=( A202  and  (not A201) );
 a72318a <=( a72317a  and  a72314a );
 a72319a <=( a72318a  and  a72311a );
 a72323a <=( (not A267)  and  (not A266) );
 a72324a <=( A265  and  a72323a );
 a72327a <=( A269  and  (not A268) );
 a72330a <=( (not A302)  and  (not A300) );
 a72331a <=( a72330a  and  a72327a );
 a72332a <=( a72331a  and  a72324a );
 a72336a <=( (not A168)  and  (not A169) );
 a72337a <=( (not A170)  and  a72336a );
 a72340a <=( (not A166)  and  A167 );
 a72343a <=( A202  and  (not A201) );
 a72344a <=( a72343a  and  a72340a );
 a72345a <=( a72344a  and  a72337a );
 a72349a <=( (not A267)  and  (not A266) );
 a72350a <=( A265  and  a72349a );
 a72353a <=( A269  and  (not A268) );
 a72356a <=( A299  and  A298 );
 a72357a <=( a72356a  and  a72353a );
 a72358a <=( a72357a  and  a72350a );
 a72362a <=( (not A168)  and  (not A169) );
 a72363a <=( (not A170)  and  a72362a );
 a72366a <=( (not A166)  and  A167 );
 a72369a <=( A202  and  (not A201) );
 a72370a <=( a72369a  and  a72366a );
 a72371a <=( a72370a  and  a72363a );
 a72375a <=( (not A267)  and  (not A266) );
 a72376a <=( A265  and  a72375a );
 a72379a <=( A269  and  (not A268) );
 a72382a <=( (not A299)  and  (not A298) );
 a72383a <=( a72382a  and  a72379a );
 a72384a <=( a72383a  and  a72376a );
 a72388a <=( (not A168)  and  (not A169) );
 a72389a <=( (not A170)  and  a72388a );
 a72392a <=( (not A166)  and  A167 );
 a72395a <=( A202  and  (not A201) );
 a72396a <=( a72395a  and  a72392a );
 a72397a <=( a72396a  and  a72389a );
 a72401a <=( A298  and  (not A266) );
 a72402a <=( (not A265)  and  a72401a );
 a72405a <=( (not A300)  and  (not A299) );
 a72408a <=( A302  and  (not A301) );
 a72409a <=( a72408a  and  a72405a );
 a72410a <=( a72409a  and  a72402a );
 a72414a <=( (not A168)  and  (not A169) );
 a72415a <=( (not A170)  and  a72414a );
 a72418a <=( (not A166)  and  A167 );
 a72421a <=( A202  and  (not A201) );
 a72422a <=( a72421a  and  a72418a );
 a72423a <=( a72422a  and  a72415a );
 a72427a <=( (not A298)  and  (not A266) );
 a72428a <=( (not A265)  and  a72427a );
 a72431a <=( (not A300)  and  A299 );
 a72434a <=( A302  and  (not A301) );
 a72435a <=( a72434a  and  a72431a );
 a72436a <=( a72435a  and  a72428a );
 a72440a <=( (not A168)  and  (not A169) );
 a72441a <=( (not A170)  and  a72440a );
 a72444a <=( (not A166)  and  A167 );
 a72447a <=( (not A203)  and  (not A201) );
 a72448a <=( a72447a  and  a72444a );
 a72449a <=( a72448a  and  a72441a );
 a72453a <=( A269  and  (not A268) );
 a72454a <=( A267  and  a72453a );
 a72457a <=( (not A299)  and  A298 );
 a72460a <=( A301  and  A300 );
 a72461a <=( a72460a  and  a72457a );
 a72462a <=( a72461a  and  a72454a );
 a72466a <=( (not A168)  and  (not A169) );
 a72467a <=( (not A170)  and  a72466a );
 a72470a <=( (not A166)  and  A167 );
 a72473a <=( (not A203)  and  (not A201) );
 a72474a <=( a72473a  and  a72470a );
 a72475a <=( a72474a  and  a72467a );
 a72479a <=( A269  and  (not A268) );
 a72480a <=( A267  and  a72479a );
 a72483a <=( (not A299)  and  A298 );
 a72486a <=( (not A302)  and  A300 );
 a72487a <=( a72486a  and  a72483a );
 a72488a <=( a72487a  and  a72480a );
 a72492a <=( (not A168)  and  (not A169) );
 a72493a <=( (not A170)  and  a72492a );
 a72496a <=( (not A166)  and  A167 );
 a72499a <=( (not A203)  and  (not A201) );
 a72500a <=( a72499a  and  a72496a );
 a72501a <=( a72500a  and  a72493a );
 a72505a <=( A269  and  (not A268) );
 a72506a <=( A267  and  a72505a );
 a72509a <=( A299  and  (not A298) );
 a72512a <=( A301  and  A300 );
 a72513a <=( a72512a  and  a72509a );
 a72514a <=( a72513a  and  a72506a );
 a72518a <=( (not A168)  and  (not A169) );
 a72519a <=( (not A170)  and  a72518a );
 a72522a <=( (not A166)  and  A167 );
 a72525a <=( (not A203)  and  (not A201) );
 a72526a <=( a72525a  and  a72522a );
 a72527a <=( a72526a  and  a72519a );
 a72531a <=( A269  and  (not A268) );
 a72532a <=( A267  and  a72531a );
 a72535a <=( A299  and  (not A298) );
 a72538a <=( (not A302)  and  A300 );
 a72539a <=( a72538a  and  a72535a );
 a72540a <=( a72539a  and  a72532a );
 a72544a <=( (not A168)  and  (not A169) );
 a72545a <=( (not A170)  and  a72544a );
 a72548a <=( (not A166)  and  A167 );
 a72551a <=( (not A203)  and  (not A201) );
 a72552a <=( a72551a  and  a72548a );
 a72553a <=( a72552a  and  a72545a );
 a72557a <=( A298  and  A268 );
 a72558a <=( (not A267)  and  a72557a );
 a72561a <=( (not A300)  and  (not A299) );
 a72564a <=( A302  and  (not A301) );
 a72565a <=( a72564a  and  a72561a );
 a72566a <=( a72565a  and  a72558a );
 a72570a <=( (not A168)  and  (not A169) );
 a72571a <=( (not A170)  and  a72570a );
 a72574a <=( (not A166)  and  A167 );
 a72577a <=( (not A203)  and  (not A201) );
 a72578a <=( a72577a  and  a72574a );
 a72579a <=( a72578a  and  a72571a );
 a72583a <=( (not A298)  and  A268 );
 a72584a <=( (not A267)  and  a72583a );
 a72587a <=( (not A300)  and  A299 );
 a72590a <=( A302  and  (not A301) );
 a72591a <=( a72590a  and  a72587a );
 a72592a <=( a72591a  and  a72584a );
 a72596a <=( (not A168)  and  (not A169) );
 a72597a <=( (not A170)  and  a72596a );
 a72600a <=( (not A166)  and  A167 );
 a72603a <=( (not A203)  and  (not A201) );
 a72604a <=( a72603a  and  a72600a );
 a72605a <=( a72604a  and  a72597a );
 a72609a <=( A298  and  (not A269) );
 a72610a <=( (not A267)  and  a72609a );
 a72613a <=( (not A300)  and  (not A299) );
 a72616a <=( A302  and  (not A301) );
 a72617a <=( a72616a  and  a72613a );
 a72618a <=( a72617a  and  a72610a );
 a72622a <=( (not A168)  and  (not A169) );
 a72623a <=( (not A170)  and  a72622a );
 a72626a <=( (not A166)  and  A167 );
 a72629a <=( (not A203)  and  (not A201) );
 a72630a <=( a72629a  and  a72626a );
 a72631a <=( a72630a  and  a72623a );
 a72635a <=( (not A298)  and  (not A269) );
 a72636a <=( (not A267)  and  a72635a );
 a72639a <=( (not A300)  and  A299 );
 a72642a <=( A302  and  (not A301) );
 a72643a <=( a72642a  and  a72639a );
 a72644a <=( a72643a  and  a72636a );
 a72648a <=( (not A168)  and  (not A169) );
 a72649a <=( (not A170)  and  a72648a );
 a72652a <=( (not A166)  and  A167 );
 a72655a <=( (not A203)  and  (not A201) );
 a72656a <=( a72655a  and  a72652a );
 a72657a <=( a72656a  and  a72649a );
 a72661a <=( A298  and  A266 );
 a72662a <=( A265  and  a72661a );
 a72665a <=( (not A300)  and  (not A299) );
 a72668a <=( A302  and  (not A301) );
 a72669a <=( a72668a  and  a72665a );
 a72670a <=( a72669a  and  a72662a );
 a72674a <=( (not A168)  and  (not A169) );
 a72675a <=( (not A170)  and  a72674a );
 a72678a <=( (not A166)  and  A167 );
 a72681a <=( (not A203)  and  (not A201) );
 a72682a <=( a72681a  and  a72678a );
 a72683a <=( a72682a  and  a72675a );
 a72687a <=( (not A298)  and  A266 );
 a72688a <=( A265  and  a72687a );
 a72691a <=( (not A300)  and  A299 );
 a72694a <=( A302  and  (not A301) );
 a72695a <=( a72694a  and  a72691a );
 a72696a <=( a72695a  and  a72688a );
 a72700a <=( (not A168)  and  (not A169) );
 a72701a <=( (not A170)  and  a72700a );
 a72704a <=( (not A166)  and  A167 );
 a72707a <=( (not A203)  and  (not A201) );
 a72708a <=( a72707a  and  a72704a );
 a72709a <=( a72708a  and  a72701a );
 a72713a <=( A267  and  A266 );
 a72714a <=( (not A265)  and  a72713a );
 a72717a <=( A300  and  A268 );
 a72720a <=( A302  and  (not A301) );
 a72721a <=( a72720a  and  a72717a );
 a72722a <=( a72721a  and  a72714a );
 a72726a <=( (not A168)  and  (not A169) );
 a72727a <=( (not A170)  and  a72726a );
 a72730a <=( (not A166)  and  A167 );
 a72733a <=( (not A203)  and  (not A201) );
 a72734a <=( a72733a  and  a72730a );
 a72735a <=( a72734a  and  a72727a );
 a72739a <=( A267  and  A266 );
 a72740a <=( (not A265)  and  a72739a );
 a72743a <=( A300  and  (not A269) );
 a72746a <=( A302  and  (not A301) );
 a72747a <=( a72746a  and  a72743a );
 a72748a <=( a72747a  and  a72740a );
 a72752a <=( (not A168)  and  (not A169) );
 a72753a <=( (not A170)  and  a72752a );
 a72756a <=( (not A166)  and  A167 );
 a72759a <=( (not A203)  and  (not A201) );
 a72760a <=( a72759a  and  a72756a );
 a72761a <=( a72760a  and  a72753a );
 a72765a <=( (not A267)  and  A266 );
 a72766a <=( (not A265)  and  a72765a );
 a72769a <=( A269  and  (not A268) );
 a72772a <=( A301  and  (not A300) );
 a72773a <=( a72772a  and  a72769a );
 a72774a <=( a72773a  and  a72766a );
 a72778a <=( (not A168)  and  (not A169) );
 a72779a <=( (not A170)  and  a72778a );
 a72782a <=( (not A166)  and  A167 );
 a72785a <=( (not A203)  and  (not A201) );
 a72786a <=( a72785a  and  a72782a );
 a72787a <=( a72786a  and  a72779a );
 a72791a <=( (not A267)  and  A266 );
 a72792a <=( (not A265)  and  a72791a );
 a72795a <=( A269  and  (not A268) );
 a72798a <=( (not A302)  and  (not A300) );
 a72799a <=( a72798a  and  a72795a );
 a72800a <=( a72799a  and  a72792a );
 a72804a <=( (not A168)  and  (not A169) );
 a72805a <=( (not A170)  and  a72804a );
 a72808a <=( (not A166)  and  A167 );
 a72811a <=( (not A203)  and  (not A201) );
 a72812a <=( a72811a  and  a72808a );
 a72813a <=( a72812a  and  a72805a );
 a72817a <=( (not A267)  and  A266 );
 a72818a <=( (not A265)  and  a72817a );
 a72821a <=( A269  and  (not A268) );
 a72824a <=( A299  and  A298 );
 a72825a <=( a72824a  and  a72821a );
 a72826a <=( a72825a  and  a72818a );
 a72830a <=( (not A168)  and  (not A169) );
 a72831a <=( (not A170)  and  a72830a );
 a72834a <=( (not A166)  and  A167 );
 a72837a <=( (not A203)  and  (not A201) );
 a72838a <=( a72837a  and  a72834a );
 a72839a <=( a72838a  and  a72831a );
 a72843a <=( (not A267)  and  A266 );
 a72844a <=( (not A265)  and  a72843a );
 a72847a <=( A269  and  (not A268) );
 a72850a <=( (not A299)  and  (not A298) );
 a72851a <=( a72850a  and  a72847a );
 a72852a <=( a72851a  and  a72844a );
 a72856a <=( (not A168)  and  (not A169) );
 a72857a <=( (not A170)  and  a72856a );
 a72860a <=( (not A166)  and  A167 );
 a72863a <=( (not A203)  and  (not A201) );
 a72864a <=( a72863a  and  a72860a );
 a72865a <=( a72864a  and  a72857a );
 a72869a <=( A267  and  (not A266) );
 a72870a <=( A265  and  a72869a );
 a72873a <=( A300  and  A268 );
 a72876a <=( A302  and  (not A301) );
 a72877a <=( a72876a  and  a72873a );
 a72878a <=( a72877a  and  a72870a );
 a72882a <=( (not A168)  and  (not A169) );
 a72883a <=( (not A170)  and  a72882a );
 a72886a <=( (not A166)  and  A167 );
 a72889a <=( (not A203)  and  (not A201) );
 a72890a <=( a72889a  and  a72886a );
 a72891a <=( a72890a  and  a72883a );
 a72895a <=( A267  and  (not A266) );
 a72896a <=( A265  and  a72895a );
 a72899a <=( A300  and  (not A269) );
 a72902a <=( A302  and  (not A301) );
 a72903a <=( a72902a  and  a72899a );
 a72904a <=( a72903a  and  a72896a );
 a72908a <=( (not A168)  and  (not A169) );
 a72909a <=( (not A170)  and  a72908a );
 a72912a <=( (not A166)  and  A167 );
 a72915a <=( (not A203)  and  (not A201) );
 a72916a <=( a72915a  and  a72912a );
 a72917a <=( a72916a  and  a72909a );
 a72921a <=( (not A267)  and  (not A266) );
 a72922a <=( A265  and  a72921a );
 a72925a <=( A269  and  (not A268) );
 a72928a <=( A301  and  (not A300) );
 a72929a <=( a72928a  and  a72925a );
 a72930a <=( a72929a  and  a72922a );
 a72934a <=( (not A168)  and  (not A169) );
 a72935a <=( (not A170)  and  a72934a );
 a72938a <=( (not A166)  and  A167 );
 a72941a <=( (not A203)  and  (not A201) );
 a72942a <=( a72941a  and  a72938a );
 a72943a <=( a72942a  and  a72935a );
 a72947a <=( (not A267)  and  (not A266) );
 a72948a <=( A265  and  a72947a );
 a72951a <=( A269  and  (not A268) );
 a72954a <=( (not A302)  and  (not A300) );
 a72955a <=( a72954a  and  a72951a );
 a72956a <=( a72955a  and  a72948a );
 a72960a <=( (not A168)  and  (not A169) );
 a72961a <=( (not A170)  and  a72960a );
 a72964a <=( (not A166)  and  A167 );
 a72967a <=( (not A203)  and  (not A201) );
 a72968a <=( a72967a  and  a72964a );
 a72969a <=( a72968a  and  a72961a );
 a72973a <=( (not A267)  and  (not A266) );
 a72974a <=( A265  and  a72973a );
 a72977a <=( A269  and  (not A268) );
 a72980a <=( A299  and  A298 );
 a72981a <=( a72980a  and  a72977a );
 a72982a <=( a72981a  and  a72974a );
 a72986a <=( (not A168)  and  (not A169) );
 a72987a <=( (not A170)  and  a72986a );
 a72990a <=( (not A166)  and  A167 );
 a72993a <=( (not A203)  and  (not A201) );
 a72994a <=( a72993a  and  a72990a );
 a72995a <=( a72994a  and  a72987a );
 a72999a <=( (not A267)  and  (not A266) );
 a73000a <=( A265  and  a72999a );
 a73003a <=( A269  and  (not A268) );
 a73006a <=( (not A299)  and  (not A298) );
 a73007a <=( a73006a  and  a73003a );
 a73008a <=( a73007a  and  a73000a );
 a73012a <=( (not A168)  and  (not A169) );
 a73013a <=( (not A170)  and  a73012a );
 a73016a <=( (not A166)  and  A167 );
 a73019a <=( (not A203)  and  (not A201) );
 a73020a <=( a73019a  and  a73016a );
 a73021a <=( a73020a  and  a73013a );
 a73025a <=( A298  and  (not A266) );
 a73026a <=( (not A265)  and  a73025a );
 a73029a <=( (not A300)  and  (not A299) );
 a73032a <=( A302  and  (not A301) );
 a73033a <=( a73032a  and  a73029a );
 a73034a <=( a73033a  and  a73026a );
 a73038a <=( (not A168)  and  (not A169) );
 a73039a <=( (not A170)  and  a73038a );
 a73042a <=( (not A166)  and  A167 );
 a73045a <=( (not A203)  and  (not A201) );
 a73046a <=( a73045a  and  a73042a );
 a73047a <=( a73046a  and  a73039a );
 a73051a <=( (not A298)  and  (not A266) );
 a73052a <=( (not A265)  and  a73051a );
 a73055a <=( (not A300)  and  A299 );
 a73058a <=( A302  and  (not A301) );
 a73059a <=( a73058a  and  a73055a );
 a73060a <=( a73059a  and  a73052a );
 a73064a <=( (not A168)  and  (not A169) );
 a73065a <=( (not A170)  and  a73064a );
 a73068a <=( (not A166)  and  A167 );
 a73071a <=( A200  and  A199 );
 a73072a <=( a73071a  and  a73068a );
 a73073a <=( a73072a  and  a73065a );
 a73077a <=( A269  and  (not A268) );
 a73078a <=( A267  and  a73077a );
 a73081a <=( (not A299)  and  A298 );
 a73084a <=( A301  and  A300 );
 a73085a <=( a73084a  and  a73081a );
 a73086a <=( a73085a  and  a73078a );
 a73090a <=( (not A168)  and  (not A169) );
 a73091a <=( (not A170)  and  a73090a );
 a73094a <=( (not A166)  and  A167 );
 a73097a <=( A200  and  A199 );
 a73098a <=( a73097a  and  a73094a );
 a73099a <=( a73098a  and  a73091a );
 a73103a <=( A269  and  (not A268) );
 a73104a <=( A267  and  a73103a );
 a73107a <=( (not A299)  and  A298 );
 a73110a <=( (not A302)  and  A300 );
 a73111a <=( a73110a  and  a73107a );
 a73112a <=( a73111a  and  a73104a );
 a73116a <=( (not A168)  and  (not A169) );
 a73117a <=( (not A170)  and  a73116a );
 a73120a <=( (not A166)  and  A167 );
 a73123a <=( A200  and  A199 );
 a73124a <=( a73123a  and  a73120a );
 a73125a <=( a73124a  and  a73117a );
 a73129a <=( A269  and  (not A268) );
 a73130a <=( A267  and  a73129a );
 a73133a <=( A299  and  (not A298) );
 a73136a <=( A301  and  A300 );
 a73137a <=( a73136a  and  a73133a );
 a73138a <=( a73137a  and  a73130a );
 a73142a <=( (not A168)  and  (not A169) );
 a73143a <=( (not A170)  and  a73142a );
 a73146a <=( (not A166)  and  A167 );
 a73149a <=( A200  and  A199 );
 a73150a <=( a73149a  and  a73146a );
 a73151a <=( a73150a  and  a73143a );
 a73155a <=( A269  and  (not A268) );
 a73156a <=( A267  and  a73155a );
 a73159a <=( A299  and  (not A298) );
 a73162a <=( (not A302)  and  A300 );
 a73163a <=( a73162a  and  a73159a );
 a73164a <=( a73163a  and  a73156a );
 a73168a <=( (not A168)  and  (not A169) );
 a73169a <=( (not A170)  and  a73168a );
 a73172a <=( (not A166)  and  A167 );
 a73175a <=( A200  and  A199 );
 a73176a <=( a73175a  and  a73172a );
 a73177a <=( a73176a  and  a73169a );
 a73181a <=( A298  and  A268 );
 a73182a <=( (not A267)  and  a73181a );
 a73185a <=( (not A300)  and  (not A299) );
 a73188a <=( A302  and  (not A301) );
 a73189a <=( a73188a  and  a73185a );
 a73190a <=( a73189a  and  a73182a );
 a73194a <=( (not A168)  and  (not A169) );
 a73195a <=( (not A170)  and  a73194a );
 a73198a <=( (not A166)  and  A167 );
 a73201a <=( A200  and  A199 );
 a73202a <=( a73201a  and  a73198a );
 a73203a <=( a73202a  and  a73195a );
 a73207a <=( (not A298)  and  A268 );
 a73208a <=( (not A267)  and  a73207a );
 a73211a <=( (not A300)  and  A299 );
 a73214a <=( A302  and  (not A301) );
 a73215a <=( a73214a  and  a73211a );
 a73216a <=( a73215a  and  a73208a );
 a73220a <=( (not A168)  and  (not A169) );
 a73221a <=( (not A170)  and  a73220a );
 a73224a <=( (not A166)  and  A167 );
 a73227a <=( A200  and  A199 );
 a73228a <=( a73227a  and  a73224a );
 a73229a <=( a73228a  and  a73221a );
 a73233a <=( A298  and  (not A269) );
 a73234a <=( (not A267)  and  a73233a );
 a73237a <=( (not A300)  and  (not A299) );
 a73240a <=( A302  and  (not A301) );
 a73241a <=( a73240a  and  a73237a );
 a73242a <=( a73241a  and  a73234a );
 a73246a <=( (not A168)  and  (not A169) );
 a73247a <=( (not A170)  and  a73246a );
 a73250a <=( (not A166)  and  A167 );
 a73253a <=( A200  and  A199 );
 a73254a <=( a73253a  and  a73250a );
 a73255a <=( a73254a  and  a73247a );
 a73259a <=( (not A298)  and  (not A269) );
 a73260a <=( (not A267)  and  a73259a );
 a73263a <=( (not A300)  and  A299 );
 a73266a <=( A302  and  (not A301) );
 a73267a <=( a73266a  and  a73263a );
 a73268a <=( a73267a  and  a73260a );
 a73272a <=( (not A168)  and  (not A169) );
 a73273a <=( (not A170)  and  a73272a );
 a73276a <=( (not A166)  and  A167 );
 a73279a <=( A200  and  A199 );
 a73280a <=( a73279a  and  a73276a );
 a73281a <=( a73280a  and  a73273a );
 a73285a <=( A298  and  A266 );
 a73286a <=( A265  and  a73285a );
 a73289a <=( (not A300)  and  (not A299) );
 a73292a <=( A302  and  (not A301) );
 a73293a <=( a73292a  and  a73289a );
 a73294a <=( a73293a  and  a73286a );
 a73298a <=( (not A168)  and  (not A169) );
 a73299a <=( (not A170)  and  a73298a );
 a73302a <=( (not A166)  and  A167 );
 a73305a <=( A200  and  A199 );
 a73306a <=( a73305a  and  a73302a );
 a73307a <=( a73306a  and  a73299a );
 a73311a <=( (not A298)  and  A266 );
 a73312a <=( A265  and  a73311a );
 a73315a <=( (not A300)  and  A299 );
 a73318a <=( A302  and  (not A301) );
 a73319a <=( a73318a  and  a73315a );
 a73320a <=( a73319a  and  a73312a );
 a73324a <=( (not A168)  and  (not A169) );
 a73325a <=( (not A170)  and  a73324a );
 a73328a <=( (not A166)  and  A167 );
 a73331a <=( A200  and  A199 );
 a73332a <=( a73331a  and  a73328a );
 a73333a <=( a73332a  and  a73325a );
 a73337a <=( A267  and  A266 );
 a73338a <=( (not A265)  and  a73337a );
 a73341a <=( A300  and  A268 );
 a73344a <=( A302  and  (not A301) );
 a73345a <=( a73344a  and  a73341a );
 a73346a <=( a73345a  and  a73338a );
 a73350a <=( (not A168)  and  (not A169) );
 a73351a <=( (not A170)  and  a73350a );
 a73354a <=( (not A166)  and  A167 );
 a73357a <=( A200  and  A199 );
 a73358a <=( a73357a  and  a73354a );
 a73359a <=( a73358a  and  a73351a );
 a73363a <=( A267  and  A266 );
 a73364a <=( (not A265)  and  a73363a );
 a73367a <=( A300  and  (not A269) );
 a73370a <=( A302  and  (not A301) );
 a73371a <=( a73370a  and  a73367a );
 a73372a <=( a73371a  and  a73364a );
 a73376a <=( (not A168)  and  (not A169) );
 a73377a <=( (not A170)  and  a73376a );
 a73380a <=( (not A166)  and  A167 );
 a73383a <=( A200  and  A199 );
 a73384a <=( a73383a  and  a73380a );
 a73385a <=( a73384a  and  a73377a );
 a73389a <=( (not A267)  and  A266 );
 a73390a <=( (not A265)  and  a73389a );
 a73393a <=( A269  and  (not A268) );
 a73396a <=( A301  and  (not A300) );
 a73397a <=( a73396a  and  a73393a );
 a73398a <=( a73397a  and  a73390a );
 a73402a <=( (not A168)  and  (not A169) );
 a73403a <=( (not A170)  and  a73402a );
 a73406a <=( (not A166)  and  A167 );
 a73409a <=( A200  and  A199 );
 a73410a <=( a73409a  and  a73406a );
 a73411a <=( a73410a  and  a73403a );
 a73415a <=( (not A267)  and  A266 );
 a73416a <=( (not A265)  and  a73415a );
 a73419a <=( A269  and  (not A268) );
 a73422a <=( (not A302)  and  (not A300) );
 a73423a <=( a73422a  and  a73419a );
 a73424a <=( a73423a  and  a73416a );
 a73428a <=( (not A168)  and  (not A169) );
 a73429a <=( (not A170)  and  a73428a );
 a73432a <=( (not A166)  and  A167 );
 a73435a <=( A200  and  A199 );
 a73436a <=( a73435a  and  a73432a );
 a73437a <=( a73436a  and  a73429a );
 a73441a <=( (not A267)  and  A266 );
 a73442a <=( (not A265)  and  a73441a );
 a73445a <=( A269  and  (not A268) );
 a73448a <=( A299  and  A298 );
 a73449a <=( a73448a  and  a73445a );
 a73450a <=( a73449a  and  a73442a );
 a73454a <=( (not A168)  and  (not A169) );
 a73455a <=( (not A170)  and  a73454a );
 a73458a <=( (not A166)  and  A167 );
 a73461a <=( A200  and  A199 );
 a73462a <=( a73461a  and  a73458a );
 a73463a <=( a73462a  and  a73455a );
 a73467a <=( (not A267)  and  A266 );
 a73468a <=( (not A265)  and  a73467a );
 a73471a <=( A269  and  (not A268) );
 a73474a <=( (not A299)  and  (not A298) );
 a73475a <=( a73474a  and  a73471a );
 a73476a <=( a73475a  and  a73468a );
 a73480a <=( (not A168)  and  (not A169) );
 a73481a <=( (not A170)  and  a73480a );
 a73484a <=( (not A166)  and  A167 );
 a73487a <=( A200  and  A199 );
 a73488a <=( a73487a  and  a73484a );
 a73489a <=( a73488a  and  a73481a );
 a73493a <=( A267  and  (not A266) );
 a73494a <=( A265  and  a73493a );
 a73497a <=( A300  and  A268 );
 a73500a <=( A302  and  (not A301) );
 a73501a <=( a73500a  and  a73497a );
 a73502a <=( a73501a  and  a73494a );
 a73506a <=( (not A168)  and  (not A169) );
 a73507a <=( (not A170)  and  a73506a );
 a73510a <=( (not A166)  and  A167 );
 a73513a <=( A200  and  A199 );
 a73514a <=( a73513a  and  a73510a );
 a73515a <=( a73514a  and  a73507a );
 a73519a <=( A267  and  (not A266) );
 a73520a <=( A265  and  a73519a );
 a73523a <=( A300  and  (not A269) );
 a73526a <=( A302  and  (not A301) );
 a73527a <=( a73526a  and  a73523a );
 a73528a <=( a73527a  and  a73520a );
 a73532a <=( (not A168)  and  (not A169) );
 a73533a <=( (not A170)  and  a73532a );
 a73536a <=( (not A166)  and  A167 );
 a73539a <=( A200  and  A199 );
 a73540a <=( a73539a  and  a73536a );
 a73541a <=( a73540a  and  a73533a );
 a73545a <=( (not A267)  and  (not A266) );
 a73546a <=( A265  and  a73545a );
 a73549a <=( A269  and  (not A268) );
 a73552a <=( A301  and  (not A300) );
 a73553a <=( a73552a  and  a73549a );
 a73554a <=( a73553a  and  a73546a );
 a73558a <=( (not A168)  and  (not A169) );
 a73559a <=( (not A170)  and  a73558a );
 a73562a <=( (not A166)  and  A167 );
 a73565a <=( A200  and  A199 );
 a73566a <=( a73565a  and  a73562a );
 a73567a <=( a73566a  and  a73559a );
 a73571a <=( (not A267)  and  (not A266) );
 a73572a <=( A265  and  a73571a );
 a73575a <=( A269  and  (not A268) );
 a73578a <=( (not A302)  and  (not A300) );
 a73579a <=( a73578a  and  a73575a );
 a73580a <=( a73579a  and  a73572a );
 a73584a <=( (not A168)  and  (not A169) );
 a73585a <=( (not A170)  and  a73584a );
 a73588a <=( (not A166)  and  A167 );
 a73591a <=( A200  and  A199 );
 a73592a <=( a73591a  and  a73588a );
 a73593a <=( a73592a  and  a73585a );
 a73597a <=( (not A267)  and  (not A266) );
 a73598a <=( A265  and  a73597a );
 a73601a <=( A269  and  (not A268) );
 a73604a <=( A299  and  A298 );
 a73605a <=( a73604a  and  a73601a );
 a73606a <=( a73605a  and  a73598a );
 a73610a <=( (not A168)  and  (not A169) );
 a73611a <=( (not A170)  and  a73610a );
 a73614a <=( (not A166)  and  A167 );
 a73617a <=( A200  and  A199 );
 a73618a <=( a73617a  and  a73614a );
 a73619a <=( a73618a  and  a73611a );
 a73623a <=( (not A267)  and  (not A266) );
 a73624a <=( A265  and  a73623a );
 a73627a <=( A269  and  (not A268) );
 a73630a <=( (not A299)  and  (not A298) );
 a73631a <=( a73630a  and  a73627a );
 a73632a <=( a73631a  and  a73624a );
 a73636a <=( (not A168)  and  (not A169) );
 a73637a <=( (not A170)  and  a73636a );
 a73640a <=( (not A166)  and  A167 );
 a73643a <=( A200  and  A199 );
 a73644a <=( a73643a  and  a73640a );
 a73645a <=( a73644a  and  a73637a );
 a73649a <=( A298  and  (not A266) );
 a73650a <=( (not A265)  and  a73649a );
 a73653a <=( (not A300)  and  (not A299) );
 a73656a <=( A302  and  (not A301) );
 a73657a <=( a73656a  and  a73653a );
 a73658a <=( a73657a  and  a73650a );
 a73662a <=( (not A168)  and  (not A169) );
 a73663a <=( (not A170)  and  a73662a );
 a73666a <=( (not A166)  and  A167 );
 a73669a <=( A200  and  A199 );
 a73670a <=( a73669a  and  a73666a );
 a73671a <=( a73670a  and  a73663a );
 a73675a <=( (not A298)  and  (not A266) );
 a73676a <=( (not A265)  and  a73675a );
 a73679a <=( (not A300)  and  A299 );
 a73682a <=( A302  and  (not A301) );
 a73683a <=( a73682a  and  a73679a );
 a73684a <=( a73683a  and  a73676a );
 a73688a <=( (not A168)  and  (not A169) );
 a73689a <=( (not A170)  and  a73688a );
 a73692a <=( (not A166)  and  A167 );
 a73695a <=( (not A200)  and  (not A199) );
 a73696a <=( a73695a  and  a73692a );
 a73697a <=( a73696a  and  a73689a );
 a73701a <=( A269  and  (not A268) );
 a73702a <=( A267  and  a73701a );
 a73705a <=( (not A299)  and  A298 );
 a73708a <=( A301  and  A300 );
 a73709a <=( a73708a  and  a73705a );
 a73710a <=( a73709a  and  a73702a );
 a73714a <=( (not A168)  and  (not A169) );
 a73715a <=( (not A170)  and  a73714a );
 a73718a <=( (not A166)  and  A167 );
 a73721a <=( (not A200)  and  (not A199) );
 a73722a <=( a73721a  and  a73718a );
 a73723a <=( a73722a  and  a73715a );
 a73727a <=( A269  and  (not A268) );
 a73728a <=( A267  and  a73727a );
 a73731a <=( (not A299)  and  A298 );
 a73734a <=( (not A302)  and  A300 );
 a73735a <=( a73734a  and  a73731a );
 a73736a <=( a73735a  and  a73728a );
 a73740a <=( (not A168)  and  (not A169) );
 a73741a <=( (not A170)  and  a73740a );
 a73744a <=( (not A166)  and  A167 );
 a73747a <=( (not A200)  and  (not A199) );
 a73748a <=( a73747a  and  a73744a );
 a73749a <=( a73748a  and  a73741a );
 a73753a <=( A269  and  (not A268) );
 a73754a <=( A267  and  a73753a );
 a73757a <=( A299  and  (not A298) );
 a73760a <=( A301  and  A300 );
 a73761a <=( a73760a  and  a73757a );
 a73762a <=( a73761a  and  a73754a );
 a73766a <=( (not A168)  and  (not A169) );
 a73767a <=( (not A170)  and  a73766a );
 a73770a <=( (not A166)  and  A167 );
 a73773a <=( (not A200)  and  (not A199) );
 a73774a <=( a73773a  and  a73770a );
 a73775a <=( a73774a  and  a73767a );
 a73779a <=( A269  and  (not A268) );
 a73780a <=( A267  and  a73779a );
 a73783a <=( A299  and  (not A298) );
 a73786a <=( (not A302)  and  A300 );
 a73787a <=( a73786a  and  a73783a );
 a73788a <=( a73787a  and  a73780a );
 a73792a <=( (not A168)  and  (not A169) );
 a73793a <=( (not A170)  and  a73792a );
 a73796a <=( (not A166)  and  A167 );
 a73799a <=( (not A200)  and  (not A199) );
 a73800a <=( a73799a  and  a73796a );
 a73801a <=( a73800a  and  a73793a );
 a73805a <=( A298  and  A268 );
 a73806a <=( (not A267)  and  a73805a );
 a73809a <=( (not A300)  and  (not A299) );
 a73812a <=( A302  and  (not A301) );
 a73813a <=( a73812a  and  a73809a );
 a73814a <=( a73813a  and  a73806a );
 a73818a <=( (not A168)  and  (not A169) );
 a73819a <=( (not A170)  and  a73818a );
 a73822a <=( (not A166)  and  A167 );
 a73825a <=( (not A200)  and  (not A199) );
 a73826a <=( a73825a  and  a73822a );
 a73827a <=( a73826a  and  a73819a );
 a73831a <=( (not A298)  and  A268 );
 a73832a <=( (not A267)  and  a73831a );
 a73835a <=( (not A300)  and  A299 );
 a73838a <=( A302  and  (not A301) );
 a73839a <=( a73838a  and  a73835a );
 a73840a <=( a73839a  and  a73832a );
 a73844a <=( (not A168)  and  (not A169) );
 a73845a <=( (not A170)  and  a73844a );
 a73848a <=( (not A166)  and  A167 );
 a73851a <=( (not A200)  and  (not A199) );
 a73852a <=( a73851a  and  a73848a );
 a73853a <=( a73852a  and  a73845a );
 a73857a <=( A298  and  (not A269) );
 a73858a <=( (not A267)  and  a73857a );
 a73861a <=( (not A300)  and  (not A299) );
 a73864a <=( A302  and  (not A301) );
 a73865a <=( a73864a  and  a73861a );
 a73866a <=( a73865a  and  a73858a );
 a73870a <=( (not A168)  and  (not A169) );
 a73871a <=( (not A170)  and  a73870a );
 a73874a <=( (not A166)  and  A167 );
 a73877a <=( (not A200)  and  (not A199) );
 a73878a <=( a73877a  and  a73874a );
 a73879a <=( a73878a  and  a73871a );
 a73883a <=( (not A298)  and  (not A269) );
 a73884a <=( (not A267)  and  a73883a );
 a73887a <=( (not A300)  and  A299 );
 a73890a <=( A302  and  (not A301) );
 a73891a <=( a73890a  and  a73887a );
 a73892a <=( a73891a  and  a73884a );
 a73896a <=( (not A168)  and  (not A169) );
 a73897a <=( (not A170)  and  a73896a );
 a73900a <=( (not A166)  and  A167 );
 a73903a <=( (not A200)  and  (not A199) );
 a73904a <=( a73903a  and  a73900a );
 a73905a <=( a73904a  and  a73897a );
 a73909a <=( A298  and  A266 );
 a73910a <=( A265  and  a73909a );
 a73913a <=( (not A300)  and  (not A299) );
 a73916a <=( A302  and  (not A301) );
 a73917a <=( a73916a  and  a73913a );
 a73918a <=( a73917a  and  a73910a );
 a73922a <=( (not A168)  and  (not A169) );
 a73923a <=( (not A170)  and  a73922a );
 a73926a <=( (not A166)  and  A167 );
 a73929a <=( (not A200)  and  (not A199) );
 a73930a <=( a73929a  and  a73926a );
 a73931a <=( a73930a  and  a73923a );
 a73935a <=( (not A298)  and  A266 );
 a73936a <=( A265  and  a73935a );
 a73939a <=( (not A300)  and  A299 );
 a73942a <=( A302  and  (not A301) );
 a73943a <=( a73942a  and  a73939a );
 a73944a <=( a73943a  and  a73936a );
 a73948a <=( (not A168)  and  (not A169) );
 a73949a <=( (not A170)  and  a73948a );
 a73952a <=( (not A166)  and  A167 );
 a73955a <=( (not A200)  and  (not A199) );
 a73956a <=( a73955a  and  a73952a );
 a73957a <=( a73956a  and  a73949a );
 a73961a <=( A267  and  A266 );
 a73962a <=( (not A265)  and  a73961a );
 a73965a <=( A300  and  A268 );
 a73968a <=( A302  and  (not A301) );
 a73969a <=( a73968a  and  a73965a );
 a73970a <=( a73969a  and  a73962a );
 a73974a <=( (not A168)  and  (not A169) );
 a73975a <=( (not A170)  and  a73974a );
 a73978a <=( (not A166)  and  A167 );
 a73981a <=( (not A200)  and  (not A199) );
 a73982a <=( a73981a  and  a73978a );
 a73983a <=( a73982a  and  a73975a );
 a73987a <=( A267  and  A266 );
 a73988a <=( (not A265)  and  a73987a );
 a73991a <=( A300  and  (not A269) );
 a73994a <=( A302  and  (not A301) );
 a73995a <=( a73994a  and  a73991a );
 a73996a <=( a73995a  and  a73988a );
 a74000a <=( (not A168)  and  (not A169) );
 a74001a <=( (not A170)  and  a74000a );
 a74004a <=( (not A166)  and  A167 );
 a74007a <=( (not A200)  and  (not A199) );
 a74008a <=( a74007a  and  a74004a );
 a74009a <=( a74008a  and  a74001a );
 a74013a <=( (not A267)  and  A266 );
 a74014a <=( (not A265)  and  a74013a );
 a74017a <=( A269  and  (not A268) );
 a74020a <=( A301  and  (not A300) );
 a74021a <=( a74020a  and  a74017a );
 a74022a <=( a74021a  and  a74014a );
 a74026a <=( (not A168)  and  (not A169) );
 a74027a <=( (not A170)  and  a74026a );
 a74030a <=( (not A166)  and  A167 );
 a74033a <=( (not A200)  and  (not A199) );
 a74034a <=( a74033a  and  a74030a );
 a74035a <=( a74034a  and  a74027a );
 a74039a <=( (not A267)  and  A266 );
 a74040a <=( (not A265)  and  a74039a );
 a74043a <=( A269  and  (not A268) );
 a74046a <=( (not A302)  and  (not A300) );
 a74047a <=( a74046a  and  a74043a );
 a74048a <=( a74047a  and  a74040a );
 a74052a <=( (not A168)  and  (not A169) );
 a74053a <=( (not A170)  and  a74052a );
 a74056a <=( (not A166)  and  A167 );
 a74059a <=( (not A200)  and  (not A199) );
 a74060a <=( a74059a  and  a74056a );
 a74061a <=( a74060a  and  a74053a );
 a74065a <=( (not A267)  and  A266 );
 a74066a <=( (not A265)  and  a74065a );
 a74069a <=( A269  and  (not A268) );
 a74072a <=( A299  and  A298 );
 a74073a <=( a74072a  and  a74069a );
 a74074a <=( a74073a  and  a74066a );
 a74078a <=( (not A168)  and  (not A169) );
 a74079a <=( (not A170)  and  a74078a );
 a74082a <=( (not A166)  and  A167 );
 a74085a <=( (not A200)  and  (not A199) );
 a74086a <=( a74085a  and  a74082a );
 a74087a <=( a74086a  and  a74079a );
 a74091a <=( (not A267)  and  A266 );
 a74092a <=( (not A265)  and  a74091a );
 a74095a <=( A269  and  (not A268) );
 a74098a <=( (not A299)  and  (not A298) );
 a74099a <=( a74098a  and  a74095a );
 a74100a <=( a74099a  and  a74092a );
 a74104a <=( (not A168)  and  (not A169) );
 a74105a <=( (not A170)  and  a74104a );
 a74108a <=( (not A166)  and  A167 );
 a74111a <=( (not A200)  and  (not A199) );
 a74112a <=( a74111a  and  a74108a );
 a74113a <=( a74112a  and  a74105a );
 a74117a <=( A267  and  (not A266) );
 a74118a <=( A265  and  a74117a );
 a74121a <=( A300  and  A268 );
 a74124a <=( A302  and  (not A301) );
 a74125a <=( a74124a  and  a74121a );
 a74126a <=( a74125a  and  a74118a );
 a74130a <=( (not A168)  and  (not A169) );
 a74131a <=( (not A170)  and  a74130a );
 a74134a <=( (not A166)  and  A167 );
 a74137a <=( (not A200)  and  (not A199) );
 a74138a <=( a74137a  and  a74134a );
 a74139a <=( a74138a  and  a74131a );
 a74143a <=( A267  and  (not A266) );
 a74144a <=( A265  and  a74143a );
 a74147a <=( A300  and  (not A269) );
 a74150a <=( A302  and  (not A301) );
 a74151a <=( a74150a  and  a74147a );
 a74152a <=( a74151a  and  a74144a );
 a74156a <=( (not A168)  and  (not A169) );
 a74157a <=( (not A170)  and  a74156a );
 a74160a <=( (not A166)  and  A167 );
 a74163a <=( (not A200)  and  (not A199) );
 a74164a <=( a74163a  and  a74160a );
 a74165a <=( a74164a  and  a74157a );
 a74169a <=( (not A267)  and  (not A266) );
 a74170a <=( A265  and  a74169a );
 a74173a <=( A269  and  (not A268) );
 a74176a <=( A301  and  (not A300) );
 a74177a <=( a74176a  and  a74173a );
 a74178a <=( a74177a  and  a74170a );
 a74182a <=( (not A168)  and  (not A169) );
 a74183a <=( (not A170)  and  a74182a );
 a74186a <=( (not A166)  and  A167 );
 a74189a <=( (not A200)  and  (not A199) );
 a74190a <=( a74189a  and  a74186a );
 a74191a <=( a74190a  and  a74183a );
 a74195a <=( (not A267)  and  (not A266) );
 a74196a <=( A265  and  a74195a );
 a74199a <=( A269  and  (not A268) );
 a74202a <=( (not A302)  and  (not A300) );
 a74203a <=( a74202a  and  a74199a );
 a74204a <=( a74203a  and  a74196a );
 a74208a <=( (not A168)  and  (not A169) );
 a74209a <=( (not A170)  and  a74208a );
 a74212a <=( (not A166)  and  A167 );
 a74215a <=( (not A200)  and  (not A199) );
 a74216a <=( a74215a  and  a74212a );
 a74217a <=( a74216a  and  a74209a );
 a74221a <=( (not A267)  and  (not A266) );
 a74222a <=( A265  and  a74221a );
 a74225a <=( A269  and  (not A268) );
 a74228a <=( A299  and  A298 );
 a74229a <=( a74228a  and  a74225a );
 a74230a <=( a74229a  and  a74222a );
 a74234a <=( (not A168)  and  (not A169) );
 a74235a <=( (not A170)  and  a74234a );
 a74238a <=( (not A166)  and  A167 );
 a74241a <=( (not A200)  and  (not A199) );
 a74242a <=( a74241a  and  a74238a );
 a74243a <=( a74242a  and  a74235a );
 a74247a <=( (not A267)  and  (not A266) );
 a74248a <=( A265  and  a74247a );
 a74251a <=( A269  and  (not A268) );
 a74254a <=( (not A299)  and  (not A298) );
 a74255a <=( a74254a  and  a74251a );
 a74256a <=( a74255a  and  a74248a );
 a74260a <=( (not A168)  and  (not A169) );
 a74261a <=( (not A170)  and  a74260a );
 a74264a <=( (not A166)  and  A167 );
 a74267a <=( (not A200)  and  (not A199) );
 a74268a <=( a74267a  and  a74264a );
 a74269a <=( a74268a  and  a74261a );
 a74273a <=( A298  and  (not A266) );
 a74274a <=( (not A265)  and  a74273a );
 a74277a <=( (not A300)  and  (not A299) );
 a74280a <=( A302  and  (not A301) );
 a74281a <=( a74280a  and  a74277a );
 a74282a <=( a74281a  and  a74274a );
 a74286a <=( (not A168)  and  (not A169) );
 a74287a <=( (not A170)  and  a74286a );
 a74290a <=( (not A166)  and  A167 );
 a74293a <=( (not A200)  and  (not A199) );
 a74294a <=( a74293a  and  a74290a );
 a74295a <=( a74294a  and  a74287a );
 a74299a <=( (not A298)  and  (not A266) );
 a74300a <=( (not A265)  and  a74299a );
 a74303a <=( (not A300)  and  A299 );
 a74306a <=( A302  and  (not A301) );
 a74307a <=( a74306a  and  a74303a );
 a74308a <=( a74307a  and  a74300a );
 a74312a <=( (not A168)  and  (not A169) );
 a74313a <=( (not A170)  and  a74312a );
 a74316a <=( A166  and  (not A167) );
 a74319a <=( (not A202)  and  A201 );
 a74320a <=( a74319a  and  a74316a );
 a74321a <=( a74320a  and  a74313a );
 a74325a <=( A268  and  (not A267) );
 a74326a <=( A203  and  a74325a );
 a74329a <=( (not A299)  and  A298 );
 a74332a <=( A301  and  A300 );
 a74333a <=( a74332a  and  a74329a );
 a74334a <=( a74333a  and  a74326a );
 a74338a <=( (not A168)  and  (not A169) );
 a74339a <=( (not A170)  and  a74338a );
 a74342a <=( A166  and  (not A167) );
 a74345a <=( (not A202)  and  A201 );
 a74346a <=( a74345a  and  a74342a );
 a74347a <=( a74346a  and  a74339a );
 a74351a <=( A268  and  (not A267) );
 a74352a <=( A203  and  a74351a );
 a74355a <=( (not A299)  and  A298 );
 a74358a <=( (not A302)  and  A300 );
 a74359a <=( a74358a  and  a74355a );
 a74360a <=( a74359a  and  a74352a );
 a74364a <=( (not A168)  and  (not A169) );
 a74365a <=( (not A170)  and  a74364a );
 a74368a <=( A166  and  (not A167) );
 a74371a <=( (not A202)  and  A201 );
 a74372a <=( a74371a  and  a74368a );
 a74373a <=( a74372a  and  a74365a );
 a74377a <=( A268  and  (not A267) );
 a74378a <=( A203  and  a74377a );
 a74381a <=( A299  and  (not A298) );
 a74384a <=( A301  and  A300 );
 a74385a <=( a74384a  and  a74381a );
 a74386a <=( a74385a  and  a74378a );
 a74390a <=( (not A168)  and  (not A169) );
 a74391a <=( (not A170)  and  a74390a );
 a74394a <=( A166  and  (not A167) );
 a74397a <=( (not A202)  and  A201 );
 a74398a <=( a74397a  and  a74394a );
 a74399a <=( a74398a  and  a74391a );
 a74403a <=( A268  and  (not A267) );
 a74404a <=( A203  and  a74403a );
 a74407a <=( A299  and  (not A298) );
 a74410a <=( (not A302)  and  A300 );
 a74411a <=( a74410a  and  a74407a );
 a74412a <=( a74411a  and  a74404a );
 a74416a <=( (not A168)  and  (not A169) );
 a74417a <=( (not A170)  and  a74416a );
 a74420a <=( A166  and  (not A167) );
 a74423a <=( (not A202)  and  A201 );
 a74424a <=( a74423a  and  a74420a );
 a74425a <=( a74424a  and  a74417a );
 a74429a <=( (not A269)  and  (not A267) );
 a74430a <=( A203  and  a74429a );
 a74433a <=( (not A299)  and  A298 );
 a74436a <=( A301  and  A300 );
 a74437a <=( a74436a  and  a74433a );
 a74438a <=( a74437a  and  a74430a );
 a74442a <=( (not A168)  and  (not A169) );
 a74443a <=( (not A170)  and  a74442a );
 a74446a <=( A166  and  (not A167) );
 a74449a <=( (not A202)  and  A201 );
 a74450a <=( a74449a  and  a74446a );
 a74451a <=( a74450a  and  a74443a );
 a74455a <=( (not A269)  and  (not A267) );
 a74456a <=( A203  and  a74455a );
 a74459a <=( (not A299)  and  A298 );
 a74462a <=( (not A302)  and  A300 );
 a74463a <=( a74462a  and  a74459a );
 a74464a <=( a74463a  and  a74456a );
 a74468a <=( (not A168)  and  (not A169) );
 a74469a <=( (not A170)  and  a74468a );
 a74472a <=( A166  and  (not A167) );
 a74475a <=( (not A202)  and  A201 );
 a74476a <=( a74475a  and  a74472a );
 a74477a <=( a74476a  and  a74469a );
 a74481a <=( (not A269)  and  (not A267) );
 a74482a <=( A203  and  a74481a );
 a74485a <=( A299  and  (not A298) );
 a74488a <=( A301  and  A300 );
 a74489a <=( a74488a  and  a74485a );
 a74490a <=( a74489a  and  a74482a );
 a74494a <=( (not A168)  and  (not A169) );
 a74495a <=( (not A170)  and  a74494a );
 a74498a <=( A166  and  (not A167) );
 a74501a <=( (not A202)  and  A201 );
 a74502a <=( a74501a  and  a74498a );
 a74503a <=( a74502a  and  a74495a );
 a74507a <=( (not A269)  and  (not A267) );
 a74508a <=( A203  and  a74507a );
 a74511a <=( A299  and  (not A298) );
 a74514a <=( (not A302)  and  A300 );
 a74515a <=( a74514a  and  a74511a );
 a74516a <=( a74515a  and  a74508a );
 a74520a <=( (not A168)  and  (not A169) );
 a74521a <=( (not A170)  and  a74520a );
 a74524a <=( A166  and  (not A167) );
 a74527a <=( (not A202)  and  A201 );
 a74528a <=( a74527a  and  a74524a );
 a74529a <=( a74528a  and  a74521a );
 a74533a <=( A266  and  A265 );
 a74534a <=( A203  and  a74533a );
 a74537a <=( (not A299)  and  A298 );
 a74540a <=( A301  and  A300 );
 a74541a <=( a74540a  and  a74537a );
 a74542a <=( a74541a  and  a74534a );
 a74546a <=( (not A168)  and  (not A169) );
 a74547a <=( (not A170)  and  a74546a );
 a74550a <=( A166  and  (not A167) );
 a74553a <=( (not A202)  and  A201 );
 a74554a <=( a74553a  and  a74550a );
 a74555a <=( a74554a  and  a74547a );
 a74559a <=( A266  and  A265 );
 a74560a <=( A203  and  a74559a );
 a74563a <=( (not A299)  and  A298 );
 a74566a <=( (not A302)  and  A300 );
 a74567a <=( a74566a  and  a74563a );
 a74568a <=( a74567a  and  a74560a );
 a74572a <=( (not A168)  and  (not A169) );
 a74573a <=( (not A170)  and  a74572a );
 a74576a <=( A166  and  (not A167) );
 a74579a <=( (not A202)  and  A201 );
 a74580a <=( a74579a  and  a74576a );
 a74581a <=( a74580a  and  a74573a );
 a74585a <=( A266  and  A265 );
 a74586a <=( A203  and  a74585a );
 a74589a <=( A299  and  (not A298) );
 a74592a <=( A301  and  A300 );
 a74593a <=( a74592a  and  a74589a );
 a74594a <=( a74593a  and  a74586a );
 a74598a <=( (not A168)  and  (not A169) );
 a74599a <=( (not A170)  and  a74598a );
 a74602a <=( A166  and  (not A167) );
 a74605a <=( (not A202)  and  A201 );
 a74606a <=( a74605a  and  a74602a );
 a74607a <=( a74606a  and  a74599a );
 a74611a <=( A266  and  A265 );
 a74612a <=( A203  and  a74611a );
 a74615a <=( A299  and  (not A298) );
 a74618a <=( (not A302)  and  A300 );
 a74619a <=( a74618a  and  a74615a );
 a74620a <=( a74619a  and  a74612a );
 a74624a <=( (not A168)  and  (not A169) );
 a74625a <=( (not A170)  and  a74624a );
 a74628a <=( A166  and  (not A167) );
 a74631a <=( (not A202)  and  A201 );
 a74632a <=( a74631a  and  a74628a );
 a74633a <=( a74632a  and  a74625a );
 a74637a <=( A266  and  (not A265) );
 a74638a <=( A203  and  a74637a );
 a74641a <=( A268  and  A267 );
 a74644a <=( A301  and  (not A300) );
 a74645a <=( a74644a  and  a74641a );
 a74646a <=( a74645a  and  a74638a );
 a74650a <=( (not A168)  and  (not A169) );
 a74651a <=( (not A170)  and  a74650a );
 a74654a <=( A166  and  (not A167) );
 a74657a <=( (not A202)  and  A201 );
 a74658a <=( a74657a  and  a74654a );
 a74659a <=( a74658a  and  a74651a );
 a74663a <=( A266  and  (not A265) );
 a74664a <=( A203  and  a74663a );
 a74667a <=( A268  and  A267 );
 a74670a <=( (not A302)  and  (not A300) );
 a74671a <=( a74670a  and  a74667a );
 a74672a <=( a74671a  and  a74664a );
 a74676a <=( (not A168)  and  (not A169) );
 a74677a <=( (not A170)  and  a74676a );
 a74680a <=( A166  and  (not A167) );
 a74683a <=( (not A202)  and  A201 );
 a74684a <=( a74683a  and  a74680a );
 a74685a <=( a74684a  and  a74677a );
 a74689a <=( A266  and  (not A265) );
 a74690a <=( A203  and  a74689a );
 a74693a <=( A268  and  A267 );
 a74696a <=( A299  and  A298 );
 a74697a <=( a74696a  and  a74693a );
 a74698a <=( a74697a  and  a74690a );
 a74702a <=( (not A168)  and  (not A169) );
 a74703a <=( (not A170)  and  a74702a );
 a74706a <=( A166  and  (not A167) );
 a74709a <=( (not A202)  and  A201 );
 a74710a <=( a74709a  and  a74706a );
 a74711a <=( a74710a  and  a74703a );
 a74715a <=( A266  and  (not A265) );
 a74716a <=( A203  and  a74715a );
 a74719a <=( A268  and  A267 );
 a74722a <=( (not A299)  and  (not A298) );
 a74723a <=( a74722a  and  a74719a );
 a74724a <=( a74723a  and  a74716a );
 a74728a <=( (not A168)  and  (not A169) );
 a74729a <=( (not A170)  and  a74728a );
 a74732a <=( A166  and  (not A167) );
 a74735a <=( (not A202)  and  A201 );
 a74736a <=( a74735a  and  a74732a );
 a74737a <=( a74736a  and  a74729a );
 a74741a <=( A266  and  (not A265) );
 a74742a <=( A203  and  a74741a );
 a74745a <=( (not A269)  and  A267 );
 a74748a <=( A301  and  (not A300) );
 a74749a <=( a74748a  and  a74745a );
 a74750a <=( a74749a  and  a74742a );
 a74754a <=( (not A168)  and  (not A169) );
 a74755a <=( (not A170)  and  a74754a );
 a74758a <=( A166  and  (not A167) );
 a74761a <=( (not A202)  and  A201 );
 a74762a <=( a74761a  and  a74758a );
 a74763a <=( a74762a  and  a74755a );
 a74767a <=( A266  and  (not A265) );
 a74768a <=( A203  and  a74767a );
 a74771a <=( (not A269)  and  A267 );
 a74774a <=( (not A302)  and  (not A300) );
 a74775a <=( a74774a  and  a74771a );
 a74776a <=( a74775a  and  a74768a );
 a74780a <=( (not A168)  and  (not A169) );
 a74781a <=( (not A170)  and  a74780a );
 a74784a <=( A166  and  (not A167) );
 a74787a <=( (not A202)  and  A201 );
 a74788a <=( a74787a  and  a74784a );
 a74789a <=( a74788a  and  a74781a );
 a74793a <=( A266  and  (not A265) );
 a74794a <=( A203  and  a74793a );
 a74797a <=( (not A269)  and  A267 );
 a74800a <=( A299  and  A298 );
 a74801a <=( a74800a  and  a74797a );
 a74802a <=( a74801a  and  a74794a );
 a74806a <=( (not A168)  and  (not A169) );
 a74807a <=( (not A170)  and  a74806a );
 a74810a <=( A166  and  (not A167) );
 a74813a <=( (not A202)  and  A201 );
 a74814a <=( a74813a  and  a74810a );
 a74815a <=( a74814a  and  a74807a );
 a74819a <=( A266  and  (not A265) );
 a74820a <=( A203  and  a74819a );
 a74823a <=( (not A269)  and  A267 );
 a74826a <=( (not A299)  and  (not A298) );
 a74827a <=( a74826a  and  a74823a );
 a74828a <=( a74827a  and  a74820a );
 a74832a <=( (not A168)  and  (not A169) );
 a74833a <=( (not A170)  and  a74832a );
 a74836a <=( A166  and  (not A167) );
 a74839a <=( (not A202)  and  A201 );
 a74840a <=( a74839a  and  a74836a );
 a74841a <=( a74840a  and  a74833a );
 a74845a <=( (not A266)  and  A265 );
 a74846a <=( A203  and  a74845a );
 a74849a <=( A268  and  A267 );
 a74852a <=( A301  and  (not A300) );
 a74853a <=( a74852a  and  a74849a );
 a74854a <=( a74853a  and  a74846a );
 a74858a <=( (not A168)  and  (not A169) );
 a74859a <=( (not A170)  and  a74858a );
 a74862a <=( A166  and  (not A167) );
 a74865a <=( (not A202)  and  A201 );
 a74866a <=( a74865a  and  a74862a );
 a74867a <=( a74866a  and  a74859a );
 a74871a <=( (not A266)  and  A265 );
 a74872a <=( A203  and  a74871a );
 a74875a <=( A268  and  A267 );
 a74878a <=( (not A302)  and  (not A300) );
 a74879a <=( a74878a  and  a74875a );
 a74880a <=( a74879a  and  a74872a );
 a74884a <=( (not A168)  and  (not A169) );
 a74885a <=( (not A170)  and  a74884a );
 a74888a <=( A166  and  (not A167) );
 a74891a <=( (not A202)  and  A201 );
 a74892a <=( a74891a  and  a74888a );
 a74893a <=( a74892a  and  a74885a );
 a74897a <=( (not A266)  and  A265 );
 a74898a <=( A203  and  a74897a );
 a74901a <=( A268  and  A267 );
 a74904a <=( A299  and  A298 );
 a74905a <=( a74904a  and  a74901a );
 a74906a <=( a74905a  and  a74898a );
 a74910a <=( (not A168)  and  (not A169) );
 a74911a <=( (not A170)  and  a74910a );
 a74914a <=( A166  and  (not A167) );
 a74917a <=( (not A202)  and  A201 );
 a74918a <=( a74917a  and  a74914a );
 a74919a <=( a74918a  and  a74911a );
 a74923a <=( (not A266)  and  A265 );
 a74924a <=( A203  and  a74923a );
 a74927a <=( A268  and  A267 );
 a74930a <=( (not A299)  and  (not A298) );
 a74931a <=( a74930a  and  a74927a );
 a74932a <=( a74931a  and  a74924a );
 a74936a <=( (not A168)  and  (not A169) );
 a74937a <=( (not A170)  and  a74936a );
 a74940a <=( A166  and  (not A167) );
 a74943a <=( (not A202)  and  A201 );
 a74944a <=( a74943a  and  a74940a );
 a74945a <=( a74944a  and  a74937a );
 a74949a <=( (not A266)  and  A265 );
 a74950a <=( A203  and  a74949a );
 a74953a <=( (not A269)  and  A267 );
 a74956a <=( A301  and  (not A300) );
 a74957a <=( a74956a  and  a74953a );
 a74958a <=( a74957a  and  a74950a );
 a74962a <=( (not A168)  and  (not A169) );
 a74963a <=( (not A170)  and  a74962a );
 a74966a <=( A166  and  (not A167) );
 a74969a <=( (not A202)  and  A201 );
 a74970a <=( a74969a  and  a74966a );
 a74971a <=( a74970a  and  a74963a );
 a74975a <=( (not A266)  and  A265 );
 a74976a <=( A203  and  a74975a );
 a74979a <=( (not A269)  and  A267 );
 a74982a <=( (not A302)  and  (not A300) );
 a74983a <=( a74982a  and  a74979a );
 a74984a <=( a74983a  and  a74976a );
 a74988a <=( (not A168)  and  (not A169) );
 a74989a <=( (not A170)  and  a74988a );
 a74992a <=( A166  and  (not A167) );
 a74995a <=( (not A202)  and  A201 );
 a74996a <=( a74995a  and  a74992a );
 a74997a <=( a74996a  and  a74989a );
 a75001a <=( (not A266)  and  A265 );
 a75002a <=( A203  and  a75001a );
 a75005a <=( (not A269)  and  A267 );
 a75008a <=( A299  and  A298 );
 a75009a <=( a75008a  and  a75005a );
 a75010a <=( a75009a  and  a75002a );
 a75014a <=( (not A168)  and  (not A169) );
 a75015a <=( (not A170)  and  a75014a );
 a75018a <=( A166  and  (not A167) );
 a75021a <=( (not A202)  and  A201 );
 a75022a <=( a75021a  and  a75018a );
 a75023a <=( a75022a  and  a75015a );
 a75027a <=( (not A266)  and  A265 );
 a75028a <=( A203  and  a75027a );
 a75031a <=( (not A269)  and  A267 );
 a75034a <=( (not A299)  and  (not A298) );
 a75035a <=( a75034a  and  a75031a );
 a75036a <=( a75035a  and  a75028a );
 a75040a <=( (not A168)  and  (not A169) );
 a75041a <=( (not A170)  and  a75040a );
 a75044a <=( A166  and  (not A167) );
 a75047a <=( (not A202)  and  A201 );
 a75048a <=( a75047a  and  a75044a );
 a75049a <=( a75048a  and  a75041a );
 a75053a <=( (not A266)  and  (not A265) );
 a75054a <=( A203  and  a75053a );
 a75057a <=( (not A299)  and  A298 );
 a75060a <=( A301  and  A300 );
 a75061a <=( a75060a  and  a75057a );
 a75062a <=( a75061a  and  a75054a );
 a75066a <=( (not A168)  and  (not A169) );
 a75067a <=( (not A170)  and  a75066a );
 a75070a <=( A166  and  (not A167) );
 a75073a <=( (not A202)  and  A201 );
 a75074a <=( a75073a  and  a75070a );
 a75075a <=( a75074a  and  a75067a );
 a75079a <=( (not A266)  and  (not A265) );
 a75080a <=( A203  and  a75079a );
 a75083a <=( (not A299)  and  A298 );
 a75086a <=( (not A302)  and  A300 );
 a75087a <=( a75086a  and  a75083a );
 a75088a <=( a75087a  and  a75080a );
 a75092a <=( (not A168)  and  (not A169) );
 a75093a <=( (not A170)  and  a75092a );
 a75096a <=( A166  and  (not A167) );
 a75099a <=( (not A202)  and  A201 );
 a75100a <=( a75099a  and  a75096a );
 a75101a <=( a75100a  and  a75093a );
 a75105a <=( (not A266)  and  (not A265) );
 a75106a <=( A203  and  a75105a );
 a75109a <=( A299  and  (not A298) );
 a75112a <=( A301  and  A300 );
 a75113a <=( a75112a  and  a75109a );
 a75114a <=( a75113a  and  a75106a );
 a75118a <=( (not A168)  and  (not A169) );
 a75119a <=( (not A170)  and  a75118a );
 a75122a <=( A166  and  (not A167) );
 a75125a <=( (not A202)  and  A201 );
 a75126a <=( a75125a  and  a75122a );
 a75127a <=( a75126a  and  a75119a );
 a75131a <=( (not A266)  and  (not A265) );
 a75132a <=( A203  and  a75131a );
 a75135a <=( A299  and  (not A298) );
 a75138a <=( (not A302)  and  A300 );
 a75139a <=( a75138a  and  a75135a );
 a75140a <=( a75139a  and  a75132a );
 a75144a <=( (not A168)  and  (not A169) );
 a75145a <=( (not A170)  and  a75144a );
 a75148a <=( A166  and  (not A167) );
 a75151a <=( A202  and  (not A201) );
 a75152a <=( a75151a  and  a75148a );
 a75153a <=( a75152a  and  a75145a );
 a75157a <=( A269  and  (not A268) );
 a75158a <=( A267  and  a75157a );
 a75161a <=( (not A299)  and  A298 );
 a75164a <=( A301  and  A300 );
 a75165a <=( a75164a  and  a75161a );
 a75166a <=( a75165a  and  a75158a );
 a75170a <=( (not A168)  and  (not A169) );
 a75171a <=( (not A170)  and  a75170a );
 a75174a <=( A166  and  (not A167) );
 a75177a <=( A202  and  (not A201) );
 a75178a <=( a75177a  and  a75174a );
 a75179a <=( a75178a  and  a75171a );
 a75183a <=( A269  and  (not A268) );
 a75184a <=( A267  and  a75183a );
 a75187a <=( (not A299)  and  A298 );
 a75190a <=( (not A302)  and  A300 );
 a75191a <=( a75190a  and  a75187a );
 a75192a <=( a75191a  and  a75184a );
 a75196a <=( (not A168)  and  (not A169) );
 a75197a <=( (not A170)  and  a75196a );
 a75200a <=( A166  and  (not A167) );
 a75203a <=( A202  and  (not A201) );
 a75204a <=( a75203a  and  a75200a );
 a75205a <=( a75204a  and  a75197a );
 a75209a <=( A269  and  (not A268) );
 a75210a <=( A267  and  a75209a );
 a75213a <=( A299  and  (not A298) );
 a75216a <=( A301  and  A300 );
 a75217a <=( a75216a  and  a75213a );
 a75218a <=( a75217a  and  a75210a );
 a75222a <=( (not A168)  and  (not A169) );
 a75223a <=( (not A170)  and  a75222a );
 a75226a <=( A166  and  (not A167) );
 a75229a <=( A202  and  (not A201) );
 a75230a <=( a75229a  and  a75226a );
 a75231a <=( a75230a  and  a75223a );
 a75235a <=( A269  and  (not A268) );
 a75236a <=( A267  and  a75235a );
 a75239a <=( A299  and  (not A298) );
 a75242a <=( (not A302)  and  A300 );
 a75243a <=( a75242a  and  a75239a );
 a75244a <=( a75243a  and  a75236a );
 a75248a <=( (not A168)  and  (not A169) );
 a75249a <=( (not A170)  and  a75248a );
 a75252a <=( A166  and  (not A167) );
 a75255a <=( A202  and  (not A201) );
 a75256a <=( a75255a  and  a75252a );
 a75257a <=( a75256a  and  a75249a );
 a75261a <=( A298  and  A268 );
 a75262a <=( (not A267)  and  a75261a );
 a75265a <=( (not A300)  and  (not A299) );
 a75268a <=( A302  and  (not A301) );
 a75269a <=( a75268a  and  a75265a );
 a75270a <=( a75269a  and  a75262a );
 a75274a <=( (not A168)  and  (not A169) );
 a75275a <=( (not A170)  and  a75274a );
 a75278a <=( A166  and  (not A167) );
 a75281a <=( A202  and  (not A201) );
 a75282a <=( a75281a  and  a75278a );
 a75283a <=( a75282a  and  a75275a );
 a75287a <=( (not A298)  and  A268 );
 a75288a <=( (not A267)  and  a75287a );
 a75291a <=( (not A300)  and  A299 );
 a75294a <=( A302  and  (not A301) );
 a75295a <=( a75294a  and  a75291a );
 a75296a <=( a75295a  and  a75288a );
 a75300a <=( (not A168)  and  (not A169) );
 a75301a <=( (not A170)  and  a75300a );
 a75304a <=( A166  and  (not A167) );
 a75307a <=( A202  and  (not A201) );
 a75308a <=( a75307a  and  a75304a );
 a75309a <=( a75308a  and  a75301a );
 a75313a <=( A298  and  (not A269) );
 a75314a <=( (not A267)  and  a75313a );
 a75317a <=( (not A300)  and  (not A299) );
 a75320a <=( A302  and  (not A301) );
 a75321a <=( a75320a  and  a75317a );
 a75322a <=( a75321a  and  a75314a );
 a75326a <=( (not A168)  and  (not A169) );
 a75327a <=( (not A170)  and  a75326a );
 a75330a <=( A166  and  (not A167) );
 a75333a <=( A202  and  (not A201) );
 a75334a <=( a75333a  and  a75330a );
 a75335a <=( a75334a  and  a75327a );
 a75339a <=( (not A298)  and  (not A269) );
 a75340a <=( (not A267)  and  a75339a );
 a75343a <=( (not A300)  and  A299 );
 a75346a <=( A302  and  (not A301) );
 a75347a <=( a75346a  and  a75343a );
 a75348a <=( a75347a  and  a75340a );
 a75352a <=( (not A168)  and  (not A169) );
 a75353a <=( (not A170)  and  a75352a );
 a75356a <=( A166  and  (not A167) );
 a75359a <=( A202  and  (not A201) );
 a75360a <=( a75359a  and  a75356a );
 a75361a <=( a75360a  and  a75353a );
 a75365a <=( A298  and  A266 );
 a75366a <=( A265  and  a75365a );
 a75369a <=( (not A300)  and  (not A299) );
 a75372a <=( A302  and  (not A301) );
 a75373a <=( a75372a  and  a75369a );
 a75374a <=( a75373a  and  a75366a );
 a75378a <=( (not A168)  and  (not A169) );
 a75379a <=( (not A170)  and  a75378a );
 a75382a <=( A166  and  (not A167) );
 a75385a <=( A202  and  (not A201) );
 a75386a <=( a75385a  and  a75382a );
 a75387a <=( a75386a  and  a75379a );
 a75391a <=( (not A298)  and  A266 );
 a75392a <=( A265  and  a75391a );
 a75395a <=( (not A300)  and  A299 );
 a75398a <=( A302  and  (not A301) );
 a75399a <=( a75398a  and  a75395a );
 a75400a <=( a75399a  and  a75392a );
 a75404a <=( (not A168)  and  (not A169) );
 a75405a <=( (not A170)  and  a75404a );
 a75408a <=( A166  and  (not A167) );
 a75411a <=( A202  and  (not A201) );
 a75412a <=( a75411a  and  a75408a );
 a75413a <=( a75412a  and  a75405a );
 a75417a <=( A267  and  A266 );
 a75418a <=( (not A265)  and  a75417a );
 a75421a <=( A300  and  A268 );
 a75424a <=( A302  and  (not A301) );
 a75425a <=( a75424a  and  a75421a );
 a75426a <=( a75425a  and  a75418a );
 a75430a <=( (not A168)  and  (not A169) );
 a75431a <=( (not A170)  and  a75430a );
 a75434a <=( A166  and  (not A167) );
 a75437a <=( A202  and  (not A201) );
 a75438a <=( a75437a  and  a75434a );
 a75439a <=( a75438a  and  a75431a );
 a75443a <=( A267  and  A266 );
 a75444a <=( (not A265)  and  a75443a );
 a75447a <=( A300  and  (not A269) );
 a75450a <=( A302  and  (not A301) );
 a75451a <=( a75450a  and  a75447a );
 a75452a <=( a75451a  and  a75444a );
 a75456a <=( (not A168)  and  (not A169) );
 a75457a <=( (not A170)  and  a75456a );
 a75460a <=( A166  and  (not A167) );
 a75463a <=( A202  and  (not A201) );
 a75464a <=( a75463a  and  a75460a );
 a75465a <=( a75464a  and  a75457a );
 a75469a <=( (not A267)  and  A266 );
 a75470a <=( (not A265)  and  a75469a );
 a75473a <=( A269  and  (not A268) );
 a75476a <=( A301  and  (not A300) );
 a75477a <=( a75476a  and  a75473a );
 a75478a <=( a75477a  and  a75470a );
 a75482a <=( (not A168)  and  (not A169) );
 a75483a <=( (not A170)  and  a75482a );
 a75486a <=( A166  and  (not A167) );
 a75489a <=( A202  and  (not A201) );
 a75490a <=( a75489a  and  a75486a );
 a75491a <=( a75490a  and  a75483a );
 a75495a <=( (not A267)  and  A266 );
 a75496a <=( (not A265)  and  a75495a );
 a75499a <=( A269  and  (not A268) );
 a75502a <=( (not A302)  and  (not A300) );
 a75503a <=( a75502a  and  a75499a );
 a75504a <=( a75503a  and  a75496a );
 a75508a <=( (not A168)  and  (not A169) );
 a75509a <=( (not A170)  and  a75508a );
 a75512a <=( A166  and  (not A167) );
 a75515a <=( A202  and  (not A201) );
 a75516a <=( a75515a  and  a75512a );
 a75517a <=( a75516a  and  a75509a );
 a75521a <=( (not A267)  and  A266 );
 a75522a <=( (not A265)  and  a75521a );
 a75525a <=( A269  and  (not A268) );
 a75528a <=( A299  and  A298 );
 a75529a <=( a75528a  and  a75525a );
 a75530a <=( a75529a  and  a75522a );
 a75534a <=( (not A168)  and  (not A169) );
 a75535a <=( (not A170)  and  a75534a );
 a75538a <=( A166  and  (not A167) );
 a75541a <=( A202  and  (not A201) );
 a75542a <=( a75541a  and  a75538a );
 a75543a <=( a75542a  and  a75535a );
 a75547a <=( (not A267)  and  A266 );
 a75548a <=( (not A265)  and  a75547a );
 a75551a <=( A269  and  (not A268) );
 a75554a <=( (not A299)  and  (not A298) );
 a75555a <=( a75554a  and  a75551a );
 a75556a <=( a75555a  and  a75548a );
 a75560a <=( (not A168)  and  (not A169) );
 a75561a <=( (not A170)  and  a75560a );
 a75564a <=( A166  and  (not A167) );
 a75567a <=( A202  and  (not A201) );
 a75568a <=( a75567a  and  a75564a );
 a75569a <=( a75568a  and  a75561a );
 a75573a <=( A267  and  (not A266) );
 a75574a <=( A265  and  a75573a );
 a75577a <=( A300  and  A268 );
 a75580a <=( A302  and  (not A301) );
 a75581a <=( a75580a  and  a75577a );
 a75582a <=( a75581a  and  a75574a );
 a75586a <=( (not A168)  and  (not A169) );
 a75587a <=( (not A170)  and  a75586a );
 a75590a <=( A166  and  (not A167) );
 a75593a <=( A202  and  (not A201) );
 a75594a <=( a75593a  and  a75590a );
 a75595a <=( a75594a  and  a75587a );
 a75599a <=( A267  and  (not A266) );
 a75600a <=( A265  and  a75599a );
 a75603a <=( A300  and  (not A269) );
 a75606a <=( A302  and  (not A301) );
 a75607a <=( a75606a  and  a75603a );
 a75608a <=( a75607a  and  a75600a );
 a75612a <=( (not A168)  and  (not A169) );
 a75613a <=( (not A170)  and  a75612a );
 a75616a <=( A166  and  (not A167) );
 a75619a <=( A202  and  (not A201) );
 a75620a <=( a75619a  and  a75616a );
 a75621a <=( a75620a  and  a75613a );
 a75625a <=( (not A267)  and  (not A266) );
 a75626a <=( A265  and  a75625a );
 a75629a <=( A269  and  (not A268) );
 a75632a <=( A301  and  (not A300) );
 a75633a <=( a75632a  and  a75629a );
 a75634a <=( a75633a  and  a75626a );
 a75638a <=( (not A168)  and  (not A169) );
 a75639a <=( (not A170)  and  a75638a );
 a75642a <=( A166  and  (not A167) );
 a75645a <=( A202  and  (not A201) );
 a75646a <=( a75645a  and  a75642a );
 a75647a <=( a75646a  and  a75639a );
 a75651a <=( (not A267)  and  (not A266) );
 a75652a <=( A265  and  a75651a );
 a75655a <=( A269  and  (not A268) );
 a75658a <=( (not A302)  and  (not A300) );
 a75659a <=( a75658a  and  a75655a );
 a75660a <=( a75659a  and  a75652a );
 a75664a <=( (not A168)  and  (not A169) );
 a75665a <=( (not A170)  and  a75664a );
 a75668a <=( A166  and  (not A167) );
 a75671a <=( A202  and  (not A201) );
 a75672a <=( a75671a  and  a75668a );
 a75673a <=( a75672a  and  a75665a );
 a75677a <=( (not A267)  and  (not A266) );
 a75678a <=( A265  and  a75677a );
 a75681a <=( A269  and  (not A268) );
 a75684a <=( A299  and  A298 );
 a75685a <=( a75684a  and  a75681a );
 a75686a <=( a75685a  and  a75678a );
 a75690a <=( (not A168)  and  (not A169) );
 a75691a <=( (not A170)  and  a75690a );
 a75694a <=( A166  and  (not A167) );
 a75697a <=( A202  and  (not A201) );
 a75698a <=( a75697a  and  a75694a );
 a75699a <=( a75698a  and  a75691a );
 a75703a <=( (not A267)  and  (not A266) );
 a75704a <=( A265  and  a75703a );
 a75707a <=( A269  and  (not A268) );
 a75710a <=( (not A299)  and  (not A298) );
 a75711a <=( a75710a  and  a75707a );
 a75712a <=( a75711a  and  a75704a );
 a75716a <=( (not A168)  and  (not A169) );
 a75717a <=( (not A170)  and  a75716a );
 a75720a <=( A166  and  (not A167) );
 a75723a <=( A202  and  (not A201) );
 a75724a <=( a75723a  and  a75720a );
 a75725a <=( a75724a  and  a75717a );
 a75729a <=( A298  and  (not A266) );
 a75730a <=( (not A265)  and  a75729a );
 a75733a <=( (not A300)  and  (not A299) );
 a75736a <=( A302  and  (not A301) );
 a75737a <=( a75736a  and  a75733a );
 a75738a <=( a75737a  and  a75730a );
 a75742a <=( (not A168)  and  (not A169) );
 a75743a <=( (not A170)  and  a75742a );
 a75746a <=( A166  and  (not A167) );
 a75749a <=( A202  and  (not A201) );
 a75750a <=( a75749a  and  a75746a );
 a75751a <=( a75750a  and  a75743a );
 a75755a <=( (not A298)  and  (not A266) );
 a75756a <=( (not A265)  and  a75755a );
 a75759a <=( (not A300)  and  A299 );
 a75762a <=( A302  and  (not A301) );
 a75763a <=( a75762a  and  a75759a );
 a75764a <=( a75763a  and  a75756a );
 a75768a <=( (not A168)  and  (not A169) );
 a75769a <=( (not A170)  and  a75768a );
 a75772a <=( A166  and  (not A167) );
 a75775a <=( (not A203)  and  (not A201) );
 a75776a <=( a75775a  and  a75772a );
 a75777a <=( a75776a  and  a75769a );
 a75781a <=( A269  and  (not A268) );
 a75782a <=( A267  and  a75781a );
 a75785a <=( (not A299)  and  A298 );
 a75788a <=( A301  and  A300 );
 a75789a <=( a75788a  and  a75785a );
 a75790a <=( a75789a  and  a75782a );
 a75794a <=( (not A168)  and  (not A169) );
 a75795a <=( (not A170)  and  a75794a );
 a75798a <=( A166  and  (not A167) );
 a75801a <=( (not A203)  and  (not A201) );
 a75802a <=( a75801a  and  a75798a );
 a75803a <=( a75802a  and  a75795a );
 a75807a <=( A269  and  (not A268) );
 a75808a <=( A267  and  a75807a );
 a75811a <=( (not A299)  and  A298 );
 a75814a <=( (not A302)  and  A300 );
 a75815a <=( a75814a  and  a75811a );
 a75816a <=( a75815a  and  a75808a );
 a75820a <=( (not A168)  and  (not A169) );
 a75821a <=( (not A170)  and  a75820a );
 a75824a <=( A166  and  (not A167) );
 a75827a <=( (not A203)  and  (not A201) );
 a75828a <=( a75827a  and  a75824a );
 a75829a <=( a75828a  and  a75821a );
 a75833a <=( A269  and  (not A268) );
 a75834a <=( A267  and  a75833a );
 a75837a <=( A299  and  (not A298) );
 a75840a <=( A301  and  A300 );
 a75841a <=( a75840a  and  a75837a );
 a75842a <=( a75841a  and  a75834a );
 a75846a <=( (not A168)  and  (not A169) );
 a75847a <=( (not A170)  and  a75846a );
 a75850a <=( A166  and  (not A167) );
 a75853a <=( (not A203)  and  (not A201) );
 a75854a <=( a75853a  and  a75850a );
 a75855a <=( a75854a  and  a75847a );
 a75859a <=( A269  and  (not A268) );
 a75860a <=( A267  and  a75859a );
 a75863a <=( A299  and  (not A298) );
 a75866a <=( (not A302)  and  A300 );
 a75867a <=( a75866a  and  a75863a );
 a75868a <=( a75867a  and  a75860a );
 a75872a <=( (not A168)  and  (not A169) );
 a75873a <=( (not A170)  and  a75872a );
 a75876a <=( A166  and  (not A167) );
 a75879a <=( (not A203)  and  (not A201) );
 a75880a <=( a75879a  and  a75876a );
 a75881a <=( a75880a  and  a75873a );
 a75885a <=( A298  and  A268 );
 a75886a <=( (not A267)  and  a75885a );
 a75889a <=( (not A300)  and  (not A299) );
 a75892a <=( A302  and  (not A301) );
 a75893a <=( a75892a  and  a75889a );
 a75894a <=( a75893a  and  a75886a );
 a75898a <=( (not A168)  and  (not A169) );
 a75899a <=( (not A170)  and  a75898a );
 a75902a <=( A166  and  (not A167) );
 a75905a <=( (not A203)  and  (not A201) );
 a75906a <=( a75905a  and  a75902a );
 a75907a <=( a75906a  and  a75899a );
 a75911a <=( (not A298)  and  A268 );
 a75912a <=( (not A267)  and  a75911a );
 a75915a <=( (not A300)  and  A299 );
 a75918a <=( A302  and  (not A301) );
 a75919a <=( a75918a  and  a75915a );
 a75920a <=( a75919a  and  a75912a );
 a75924a <=( (not A168)  and  (not A169) );
 a75925a <=( (not A170)  and  a75924a );
 a75928a <=( A166  and  (not A167) );
 a75931a <=( (not A203)  and  (not A201) );
 a75932a <=( a75931a  and  a75928a );
 a75933a <=( a75932a  and  a75925a );
 a75937a <=( A298  and  (not A269) );
 a75938a <=( (not A267)  and  a75937a );
 a75941a <=( (not A300)  and  (not A299) );
 a75944a <=( A302  and  (not A301) );
 a75945a <=( a75944a  and  a75941a );
 a75946a <=( a75945a  and  a75938a );
 a75950a <=( (not A168)  and  (not A169) );
 a75951a <=( (not A170)  and  a75950a );
 a75954a <=( A166  and  (not A167) );
 a75957a <=( (not A203)  and  (not A201) );
 a75958a <=( a75957a  and  a75954a );
 a75959a <=( a75958a  and  a75951a );
 a75963a <=( (not A298)  and  (not A269) );
 a75964a <=( (not A267)  and  a75963a );
 a75967a <=( (not A300)  and  A299 );
 a75970a <=( A302  and  (not A301) );
 a75971a <=( a75970a  and  a75967a );
 a75972a <=( a75971a  and  a75964a );
 a75976a <=( (not A168)  and  (not A169) );
 a75977a <=( (not A170)  and  a75976a );
 a75980a <=( A166  and  (not A167) );
 a75983a <=( (not A203)  and  (not A201) );
 a75984a <=( a75983a  and  a75980a );
 a75985a <=( a75984a  and  a75977a );
 a75989a <=( A298  and  A266 );
 a75990a <=( A265  and  a75989a );
 a75993a <=( (not A300)  and  (not A299) );
 a75996a <=( A302  and  (not A301) );
 a75997a <=( a75996a  and  a75993a );
 a75998a <=( a75997a  and  a75990a );
 a76002a <=( (not A168)  and  (not A169) );
 a76003a <=( (not A170)  and  a76002a );
 a76006a <=( A166  and  (not A167) );
 a76009a <=( (not A203)  and  (not A201) );
 a76010a <=( a76009a  and  a76006a );
 a76011a <=( a76010a  and  a76003a );
 a76015a <=( (not A298)  and  A266 );
 a76016a <=( A265  and  a76015a );
 a76019a <=( (not A300)  and  A299 );
 a76022a <=( A302  and  (not A301) );
 a76023a <=( a76022a  and  a76019a );
 a76024a <=( a76023a  and  a76016a );
 a76028a <=( (not A168)  and  (not A169) );
 a76029a <=( (not A170)  and  a76028a );
 a76032a <=( A166  and  (not A167) );
 a76035a <=( (not A203)  and  (not A201) );
 a76036a <=( a76035a  and  a76032a );
 a76037a <=( a76036a  and  a76029a );
 a76041a <=( A267  and  A266 );
 a76042a <=( (not A265)  and  a76041a );
 a76045a <=( A300  and  A268 );
 a76048a <=( A302  and  (not A301) );
 a76049a <=( a76048a  and  a76045a );
 a76050a <=( a76049a  and  a76042a );
 a76054a <=( (not A168)  and  (not A169) );
 a76055a <=( (not A170)  and  a76054a );
 a76058a <=( A166  and  (not A167) );
 a76061a <=( (not A203)  and  (not A201) );
 a76062a <=( a76061a  and  a76058a );
 a76063a <=( a76062a  and  a76055a );
 a76067a <=( A267  and  A266 );
 a76068a <=( (not A265)  and  a76067a );
 a76071a <=( A300  and  (not A269) );
 a76074a <=( A302  and  (not A301) );
 a76075a <=( a76074a  and  a76071a );
 a76076a <=( a76075a  and  a76068a );
 a76080a <=( (not A168)  and  (not A169) );
 a76081a <=( (not A170)  and  a76080a );
 a76084a <=( A166  and  (not A167) );
 a76087a <=( (not A203)  and  (not A201) );
 a76088a <=( a76087a  and  a76084a );
 a76089a <=( a76088a  and  a76081a );
 a76093a <=( (not A267)  and  A266 );
 a76094a <=( (not A265)  and  a76093a );
 a76097a <=( A269  and  (not A268) );
 a76100a <=( A301  and  (not A300) );
 a76101a <=( a76100a  and  a76097a );
 a76102a <=( a76101a  and  a76094a );
 a76106a <=( (not A168)  and  (not A169) );
 a76107a <=( (not A170)  and  a76106a );
 a76110a <=( A166  and  (not A167) );
 a76113a <=( (not A203)  and  (not A201) );
 a76114a <=( a76113a  and  a76110a );
 a76115a <=( a76114a  and  a76107a );
 a76119a <=( (not A267)  and  A266 );
 a76120a <=( (not A265)  and  a76119a );
 a76123a <=( A269  and  (not A268) );
 a76126a <=( (not A302)  and  (not A300) );
 a76127a <=( a76126a  and  a76123a );
 a76128a <=( a76127a  and  a76120a );
 a76132a <=( (not A168)  and  (not A169) );
 a76133a <=( (not A170)  and  a76132a );
 a76136a <=( A166  and  (not A167) );
 a76139a <=( (not A203)  and  (not A201) );
 a76140a <=( a76139a  and  a76136a );
 a76141a <=( a76140a  and  a76133a );
 a76145a <=( (not A267)  and  A266 );
 a76146a <=( (not A265)  and  a76145a );
 a76149a <=( A269  and  (not A268) );
 a76152a <=( A299  and  A298 );
 a76153a <=( a76152a  and  a76149a );
 a76154a <=( a76153a  and  a76146a );
 a76158a <=( (not A168)  and  (not A169) );
 a76159a <=( (not A170)  and  a76158a );
 a76162a <=( A166  and  (not A167) );
 a76165a <=( (not A203)  and  (not A201) );
 a76166a <=( a76165a  and  a76162a );
 a76167a <=( a76166a  and  a76159a );
 a76171a <=( (not A267)  and  A266 );
 a76172a <=( (not A265)  and  a76171a );
 a76175a <=( A269  and  (not A268) );
 a76178a <=( (not A299)  and  (not A298) );
 a76179a <=( a76178a  and  a76175a );
 a76180a <=( a76179a  and  a76172a );
 a76184a <=( (not A168)  and  (not A169) );
 a76185a <=( (not A170)  and  a76184a );
 a76188a <=( A166  and  (not A167) );
 a76191a <=( (not A203)  and  (not A201) );
 a76192a <=( a76191a  and  a76188a );
 a76193a <=( a76192a  and  a76185a );
 a76197a <=( A267  and  (not A266) );
 a76198a <=( A265  and  a76197a );
 a76201a <=( A300  and  A268 );
 a76204a <=( A302  and  (not A301) );
 a76205a <=( a76204a  and  a76201a );
 a76206a <=( a76205a  and  a76198a );
 a76210a <=( (not A168)  and  (not A169) );
 a76211a <=( (not A170)  and  a76210a );
 a76214a <=( A166  and  (not A167) );
 a76217a <=( (not A203)  and  (not A201) );
 a76218a <=( a76217a  and  a76214a );
 a76219a <=( a76218a  and  a76211a );
 a76223a <=( A267  and  (not A266) );
 a76224a <=( A265  and  a76223a );
 a76227a <=( A300  and  (not A269) );
 a76230a <=( A302  and  (not A301) );
 a76231a <=( a76230a  and  a76227a );
 a76232a <=( a76231a  and  a76224a );
 a76236a <=( (not A168)  and  (not A169) );
 a76237a <=( (not A170)  and  a76236a );
 a76240a <=( A166  and  (not A167) );
 a76243a <=( (not A203)  and  (not A201) );
 a76244a <=( a76243a  and  a76240a );
 a76245a <=( a76244a  and  a76237a );
 a76249a <=( (not A267)  and  (not A266) );
 a76250a <=( A265  and  a76249a );
 a76253a <=( A269  and  (not A268) );
 a76256a <=( A301  and  (not A300) );
 a76257a <=( a76256a  and  a76253a );
 a76258a <=( a76257a  and  a76250a );
 a76262a <=( (not A168)  and  (not A169) );
 a76263a <=( (not A170)  and  a76262a );
 a76266a <=( A166  and  (not A167) );
 a76269a <=( (not A203)  and  (not A201) );
 a76270a <=( a76269a  and  a76266a );
 a76271a <=( a76270a  and  a76263a );
 a76275a <=( (not A267)  and  (not A266) );
 a76276a <=( A265  and  a76275a );
 a76279a <=( A269  and  (not A268) );
 a76282a <=( (not A302)  and  (not A300) );
 a76283a <=( a76282a  and  a76279a );
 a76284a <=( a76283a  and  a76276a );
 a76288a <=( (not A168)  and  (not A169) );
 a76289a <=( (not A170)  and  a76288a );
 a76292a <=( A166  and  (not A167) );
 a76295a <=( (not A203)  and  (not A201) );
 a76296a <=( a76295a  and  a76292a );
 a76297a <=( a76296a  and  a76289a );
 a76301a <=( (not A267)  and  (not A266) );
 a76302a <=( A265  and  a76301a );
 a76305a <=( A269  and  (not A268) );
 a76308a <=( A299  and  A298 );
 a76309a <=( a76308a  and  a76305a );
 a76310a <=( a76309a  and  a76302a );
 a76314a <=( (not A168)  and  (not A169) );
 a76315a <=( (not A170)  and  a76314a );
 a76318a <=( A166  and  (not A167) );
 a76321a <=( (not A203)  and  (not A201) );
 a76322a <=( a76321a  and  a76318a );
 a76323a <=( a76322a  and  a76315a );
 a76327a <=( (not A267)  and  (not A266) );
 a76328a <=( A265  and  a76327a );
 a76331a <=( A269  and  (not A268) );
 a76334a <=( (not A299)  and  (not A298) );
 a76335a <=( a76334a  and  a76331a );
 a76336a <=( a76335a  and  a76328a );
 a76340a <=( (not A168)  and  (not A169) );
 a76341a <=( (not A170)  and  a76340a );
 a76344a <=( A166  and  (not A167) );
 a76347a <=( (not A203)  and  (not A201) );
 a76348a <=( a76347a  and  a76344a );
 a76349a <=( a76348a  and  a76341a );
 a76353a <=( A298  and  (not A266) );
 a76354a <=( (not A265)  and  a76353a );
 a76357a <=( (not A300)  and  (not A299) );
 a76360a <=( A302  and  (not A301) );
 a76361a <=( a76360a  and  a76357a );
 a76362a <=( a76361a  and  a76354a );
 a76366a <=( (not A168)  and  (not A169) );
 a76367a <=( (not A170)  and  a76366a );
 a76370a <=( A166  and  (not A167) );
 a76373a <=( (not A203)  and  (not A201) );
 a76374a <=( a76373a  and  a76370a );
 a76375a <=( a76374a  and  a76367a );
 a76379a <=( (not A298)  and  (not A266) );
 a76380a <=( (not A265)  and  a76379a );
 a76383a <=( (not A300)  and  A299 );
 a76386a <=( A302  and  (not A301) );
 a76387a <=( a76386a  and  a76383a );
 a76388a <=( a76387a  and  a76380a );
 a76392a <=( (not A168)  and  (not A169) );
 a76393a <=( (not A170)  and  a76392a );
 a76396a <=( A166  and  (not A167) );
 a76399a <=( A200  and  A199 );
 a76400a <=( a76399a  and  a76396a );
 a76401a <=( a76400a  and  a76393a );
 a76405a <=( A269  and  (not A268) );
 a76406a <=( A267  and  a76405a );
 a76409a <=( (not A299)  and  A298 );
 a76412a <=( A301  and  A300 );
 a76413a <=( a76412a  and  a76409a );
 a76414a <=( a76413a  and  a76406a );
 a76418a <=( (not A168)  and  (not A169) );
 a76419a <=( (not A170)  and  a76418a );
 a76422a <=( A166  and  (not A167) );
 a76425a <=( A200  and  A199 );
 a76426a <=( a76425a  and  a76422a );
 a76427a <=( a76426a  and  a76419a );
 a76431a <=( A269  and  (not A268) );
 a76432a <=( A267  and  a76431a );
 a76435a <=( (not A299)  and  A298 );
 a76438a <=( (not A302)  and  A300 );
 a76439a <=( a76438a  and  a76435a );
 a76440a <=( a76439a  and  a76432a );
 a76444a <=( (not A168)  and  (not A169) );
 a76445a <=( (not A170)  and  a76444a );
 a76448a <=( A166  and  (not A167) );
 a76451a <=( A200  and  A199 );
 a76452a <=( a76451a  and  a76448a );
 a76453a <=( a76452a  and  a76445a );
 a76457a <=( A269  and  (not A268) );
 a76458a <=( A267  and  a76457a );
 a76461a <=( A299  and  (not A298) );
 a76464a <=( A301  and  A300 );
 a76465a <=( a76464a  and  a76461a );
 a76466a <=( a76465a  and  a76458a );
 a76470a <=( (not A168)  and  (not A169) );
 a76471a <=( (not A170)  and  a76470a );
 a76474a <=( A166  and  (not A167) );
 a76477a <=( A200  and  A199 );
 a76478a <=( a76477a  and  a76474a );
 a76479a <=( a76478a  and  a76471a );
 a76483a <=( A269  and  (not A268) );
 a76484a <=( A267  and  a76483a );
 a76487a <=( A299  and  (not A298) );
 a76490a <=( (not A302)  and  A300 );
 a76491a <=( a76490a  and  a76487a );
 a76492a <=( a76491a  and  a76484a );
 a76496a <=( (not A168)  and  (not A169) );
 a76497a <=( (not A170)  and  a76496a );
 a76500a <=( A166  and  (not A167) );
 a76503a <=( A200  and  A199 );
 a76504a <=( a76503a  and  a76500a );
 a76505a <=( a76504a  and  a76497a );
 a76509a <=( A298  and  A268 );
 a76510a <=( (not A267)  and  a76509a );
 a76513a <=( (not A300)  and  (not A299) );
 a76516a <=( A302  and  (not A301) );
 a76517a <=( a76516a  and  a76513a );
 a76518a <=( a76517a  and  a76510a );
 a76522a <=( (not A168)  and  (not A169) );
 a76523a <=( (not A170)  and  a76522a );
 a76526a <=( A166  and  (not A167) );
 a76529a <=( A200  and  A199 );
 a76530a <=( a76529a  and  a76526a );
 a76531a <=( a76530a  and  a76523a );
 a76535a <=( (not A298)  and  A268 );
 a76536a <=( (not A267)  and  a76535a );
 a76539a <=( (not A300)  and  A299 );
 a76542a <=( A302  and  (not A301) );
 a76543a <=( a76542a  and  a76539a );
 a76544a <=( a76543a  and  a76536a );
 a76548a <=( (not A168)  and  (not A169) );
 a76549a <=( (not A170)  and  a76548a );
 a76552a <=( A166  and  (not A167) );
 a76555a <=( A200  and  A199 );
 a76556a <=( a76555a  and  a76552a );
 a76557a <=( a76556a  and  a76549a );
 a76561a <=( A298  and  (not A269) );
 a76562a <=( (not A267)  and  a76561a );
 a76565a <=( (not A300)  and  (not A299) );
 a76568a <=( A302  and  (not A301) );
 a76569a <=( a76568a  and  a76565a );
 a76570a <=( a76569a  and  a76562a );
 a76574a <=( (not A168)  and  (not A169) );
 a76575a <=( (not A170)  and  a76574a );
 a76578a <=( A166  and  (not A167) );
 a76581a <=( A200  and  A199 );
 a76582a <=( a76581a  and  a76578a );
 a76583a <=( a76582a  and  a76575a );
 a76587a <=( (not A298)  and  (not A269) );
 a76588a <=( (not A267)  and  a76587a );
 a76591a <=( (not A300)  and  A299 );
 a76594a <=( A302  and  (not A301) );
 a76595a <=( a76594a  and  a76591a );
 a76596a <=( a76595a  and  a76588a );
 a76600a <=( (not A168)  and  (not A169) );
 a76601a <=( (not A170)  and  a76600a );
 a76604a <=( A166  and  (not A167) );
 a76607a <=( A200  and  A199 );
 a76608a <=( a76607a  and  a76604a );
 a76609a <=( a76608a  and  a76601a );
 a76613a <=( A298  and  A266 );
 a76614a <=( A265  and  a76613a );
 a76617a <=( (not A300)  and  (not A299) );
 a76620a <=( A302  and  (not A301) );
 a76621a <=( a76620a  and  a76617a );
 a76622a <=( a76621a  and  a76614a );
 a76626a <=( (not A168)  and  (not A169) );
 a76627a <=( (not A170)  and  a76626a );
 a76630a <=( A166  and  (not A167) );
 a76633a <=( A200  and  A199 );
 a76634a <=( a76633a  and  a76630a );
 a76635a <=( a76634a  and  a76627a );
 a76639a <=( (not A298)  and  A266 );
 a76640a <=( A265  and  a76639a );
 a76643a <=( (not A300)  and  A299 );
 a76646a <=( A302  and  (not A301) );
 a76647a <=( a76646a  and  a76643a );
 a76648a <=( a76647a  and  a76640a );
 a76652a <=( (not A168)  and  (not A169) );
 a76653a <=( (not A170)  and  a76652a );
 a76656a <=( A166  and  (not A167) );
 a76659a <=( A200  and  A199 );
 a76660a <=( a76659a  and  a76656a );
 a76661a <=( a76660a  and  a76653a );
 a76665a <=( A267  and  A266 );
 a76666a <=( (not A265)  and  a76665a );
 a76669a <=( A300  and  A268 );
 a76672a <=( A302  and  (not A301) );
 a76673a <=( a76672a  and  a76669a );
 a76674a <=( a76673a  and  a76666a );
 a76678a <=( (not A168)  and  (not A169) );
 a76679a <=( (not A170)  and  a76678a );
 a76682a <=( A166  and  (not A167) );
 a76685a <=( A200  and  A199 );
 a76686a <=( a76685a  and  a76682a );
 a76687a <=( a76686a  and  a76679a );
 a76691a <=( A267  and  A266 );
 a76692a <=( (not A265)  and  a76691a );
 a76695a <=( A300  and  (not A269) );
 a76698a <=( A302  and  (not A301) );
 a76699a <=( a76698a  and  a76695a );
 a76700a <=( a76699a  and  a76692a );
 a76704a <=( (not A168)  and  (not A169) );
 a76705a <=( (not A170)  and  a76704a );
 a76708a <=( A166  and  (not A167) );
 a76711a <=( A200  and  A199 );
 a76712a <=( a76711a  and  a76708a );
 a76713a <=( a76712a  and  a76705a );
 a76717a <=( (not A267)  and  A266 );
 a76718a <=( (not A265)  and  a76717a );
 a76721a <=( A269  and  (not A268) );
 a76724a <=( A301  and  (not A300) );
 a76725a <=( a76724a  and  a76721a );
 a76726a <=( a76725a  and  a76718a );
 a76730a <=( (not A168)  and  (not A169) );
 a76731a <=( (not A170)  and  a76730a );
 a76734a <=( A166  and  (not A167) );
 a76737a <=( A200  and  A199 );
 a76738a <=( a76737a  and  a76734a );
 a76739a <=( a76738a  and  a76731a );
 a76743a <=( (not A267)  and  A266 );
 a76744a <=( (not A265)  and  a76743a );
 a76747a <=( A269  and  (not A268) );
 a76750a <=( (not A302)  and  (not A300) );
 a76751a <=( a76750a  and  a76747a );
 a76752a <=( a76751a  and  a76744a );
 a76756a <=( (not A168)  and  (not A169) );
 a76757a <=( (not A170)  and  a76756a );
 a76760a <=( A166  and  (not A167) );
 a76763a <=( A200  and  A199 );
 a76764a <=( a76763a  and  a76760a );
 a76765a <=( a76764a  and  a76757a );
 a76769a <=( (not A267)  and  A266 );
 a76770a <=( (not A265)  and  a76769a );
 a76773a <=( A269  and  (not A268) );
 a76776a <=( A299  and  A298 );
 a76777a <=( a76776a  and  a76773a );
 a76778a <=( a76777a  and  a76770a );
 a76782a <=( (not A168)  and  (not A169) );
 a76783a <=( (not A170)  and  a76782a );
 a76786a <=( A166  and  (not A167) );
 a76789a <=( A200  and  A199 );
 a76790a <=( a76789a  and  a76786a );
 a76791a <=( a76790a  and  a76783a );
 a76795a <=( (not A267)  and  A266 );
 a76796a <=( (not A265)  and  a76795a );
 a76799a <=( A269  and  (not A268) );
 a76802a <=( (not A299)  and  (not A298) );
 a76803a <=( a76802a  and  a76799a );
 a76804a <=( a76803a  and  a76796a );
 a76808a <=( (not A168)  and  (not A169) );
 a76809a <=( (not A170)  and  a76808a );
 a76812a <=( A166  and  (not A167) );
 a76815a <=( A200  and  A199 );
 a76816a <=( a76815a  and  a76812a );
 a76817a <=( a76816a  and  a76809a );
 a76821a <=( A267  and  (not A266) );
 a76822a <=( A265  and  a76821a );
 a76825a <=( A300  and  A268 );
 a76828a <=( A302  and  (not A301) );
 a76829a <=( a76828a  and  a76825a );
 a76830a <=( a76829a  and  a76822a );
 a76834a <=( (not A168)  and  (not A169) );
 a76835a <=( (not A170)  and  a76834a );
 a76838a <=( A166  and  (not A167) );
 a76841a <=( A200  and  A199 );
 a76842a <=( a76841a  and  a76838a );
 a76843a <=( a76842a  and  a76835a );
 a76847a <=( A267  and  (not A266) );
 a76848a <=( A265  and  a76847a );
 a76851a <=( A300  and  (not A269) );
 a76854a <=( A302  and  (not A301) );
 a76855a <=( a76854a  and  a76851a );
 a76856a <=( a76855a  and  a76848a );
 a76860a <=( (not A168)  and  (not A169) );
 a76861a <=( (not A170)  and  a76860a );
 a76864a <=( A166  and  (not A167) );
 a76867a <=( A200  and  A199 );
 a76868a <=( a76867a  and  a76864a );
 a76869a <=( a76868a  and  a76861a );
 a76873a <=( (not A267)  and  (not A266) );
 a76874a <=( A265  and  a76873a );
 a76877a <=( A269  and  (not A268) );
 a76880a <=( A301  and  (not A300) );
 a76881a <=( a76880a  and  a76877a );
 a76882a <=( a76881a  and  a76874a );
 a76886a <=( (not A168)  and  (not A169) );
 a76887a <=( (not A170)  and  a76886a );
 a76890a <=( A166  and  (not A167) );
 a76893a <=( A200  and  A199 );
 a76894a <=( a76893a  and  a76890a );
 a76895a <=( a76894a  and  a76887a );
 a76899a <=( (not A267)  and  (not A266) );
 a76900a <=( A265  and  a76899a );
 a76903a <=( A269  and  (not A268) );
 a76906a <=( (not A302)  and  (not A300) );
 a76907a <=( a76906a  and  a76903a );
 a76908a <=( a76907a  and  a76900a );
 a76912a <=( (not A168)  and  (not A169) );
 a76913a <=( (not A170)  and  a76912a );
 a76916a <=( A166  and  (not A167) );
 a76919a <=( A200  and  A199 );
 a76920a <=( a76919a  and  a76916a );
 a76921a <=( a76920a  and  a76913a );
 a76925a <=( (not A267)  and  (not A266) );
 a76926a <=( A265  and  a76925a );
 a76929a <=( A269  and  (not A268) );
 a76932a <=( A299  and  A298 );
 a76933a <=( a76932a  and  a76929a );
 a76934a <=( a76933a  and  a76926a );
 a76938a <=( (not A168)  and  (not A169) );
 a76939a <=( (not A170)  and  a76938a );
 a76942a <=( A166  and  (not A167) );
 a76945a <=( A200  and  A199 );
 a76946a <=( a76945a  and  a76942a );
 a76947a <=( a76946a  and  a76939a );
 a76951a <=( (not A267)  and  (not A266) );
 a76952a <=( A265  and  a76951a );
 a76955a <=( A269  and  (not A268) );
 a76958a <=( (not A299)  and  (not A298) );
 a76959a <=( a76958a  and  a76955a );
 a76960a <=( a76959a  and  a76952a );
 a76964a <=( (not A168)  and  (not A169) );
 a76965a <=( (not A170)  and  a76964a );
 a76968a <=( A166  and  (not A167) );
 a76971a <=( A200  and  A199 );
 a76972a <=( a76971a  and  a76968a );
 a76973a <=( a76972a  and  a76965a );
 a76977a <=( A298  and  (not A266) );
 a76978a <=( (not A265)  and  a76977a );
 a76981a <=( (not A300)  and  (not A299) );
 a76984a <=( A302  and  (not A301) );
 a76985a <=( a76984a  and  a76981a );
 a76986a <=( a76985a  and  a76978a );
 a76990a <=( (not A168)  and  (not A169) );
 a76991a <=( (not A170)  and  a76990a );
 a76994a <=( A166  and  (not A167) );
 a76997a <=( A200  and  A199 );
 a76998a <=( a76997a  and  a76994a );
 a76999a <=( a76998a  and  a76991a );
 a77003a <=( (not A298)  and  (not A266) );
 a77004a <=( (not A265)  and  a77003a );
 a77007a <=( (not A300)  and  A299 );
 a77010a <=( A302  and  (not A301) );
 a77011a <=( a77010a  and  a77007a );
 a77012a <=( a77011a  and  a77004a );
 a77016a <=( (not A168)  and  (not A169) );
 a77017a <=( (not A170)  and  a77016a );
 a77020a <=( A166  and  (not A167) );
 a77023a <=( (not A200)  and  (not A199) );
 a77024a <=( a77023a  and  a77020a );
 a77025a <=( a77024a  and  a77017a );
 a77029a <=( A269  and  (not A268) );
 a77030a <=( A267  and  a77029a );
 a77033a <=( (not A299)  and  A298 );
 a77036a <=( A301  and  A300 );
 a77037a <=( a77036a  and  a77033a );
 a77038a <=( a77037a  and  a77030a );
 a77042a <=( (not A168)  and  (not A169) );
 a77043a <=( (not A170)  and  a77042a );
 a77046a <=( A166  and  (not A167) );
 a77049a <=( (not A200)  and  (not A199) );
 a77050a <=( a77049a  and  a77046a );
 a77051a <=( a77050a  and  a77043a );
 a77055a <=( A269  and  (not A268) );
 a77056a <=( A267  and  a77055a );
 a77059a <=( (not A299)  and  A298 );
 a77062a <=( (not A302)  and  A300 );
 a77063a <=( a77062a  and  a77059a );
 a77064a <=( a77063a  and  a77056a );
 a77068a <=( (not A168)  and  (not A169) );
 a77069a <=( (not A170)  and  a77068a );
 a77072a <=( A166  and  (not A167) );
 a77075a <=( (not A200)  and  (not A199) );
 a77076a <=( a77075a  and  a77072a );
 a77077a <=( a77076a  and  a77069a );
 a77081a <=( A269  and  (not A268) );
 a77082a <=( A267  and  a77081a );
 a77085a <=( A299  and  (not A298) );
 a77088a <=( A301  and  A300 );
 a77089a <=( a77088a  and  a77085a );
 a77090a <=( a77089a  and  a77082a );
 a77094a <=( (not A168)  and  (not A169) );
 a77095a <=( (not A170)  and  a77094a );
 a77098a <=( A166  and  (not A167) );
 a77101a <=( (not A200)  and  (not A199) );
 a77102a <=( a77101a  and  a77098a );
 a77103a <=( a77102a  and  a77095a );
 a77107a <=( A269  and  (not A268) );
 a77108a <=( A267  and  a77107a );
 a77111a <=( A299  and  (not A298) );
 a77114a <=( (not A302)  and  A300 );
 a77115a <=( a77114a  and  a77111a );
 a77116a <=( a77115a  and  a77108a );
 a77120a <=( (not A168)  and  (not A169) );
 a77121a <=( (not A170)  and  a77120a );
 a77124a <=( A166  and  (not A167) );
 a77127a <=( (not A200)  and  (not A199) );
 a77128a <=( a77127a  and  a77124a );
 a77129a <=( a77128a  and  a77121a );
 a77133a <=( A298  and  A268 );
 a77134a <=( (not A267)  and  a77133a );
 a77137a <=( (not A300)  and  (not A299) );
 a77140a <=( A302  and  (not A301) );
 a77141a <=( a77140a  and  a77137a );
 a77142a <=( a77141a  and  a77134a );
 a77146a <=( (not A168)  and  (not A169) );
 a77147a <=( (not A170)  and  a77146a );
 a77150a <=( A166  and  (not A167) );
 a77153a <=( (not A200)  and  (not A199) );
 a77154a <=( a77153a  and  a77150a );
 a77155a <=( a77154a  and  a77147a );
 a77159a <=( (not A298)  and  A268 );
 a77160a <=( (not A267)  and  a77159a );
 a77163a <=( (not A300)  and  A299 );
 a77166a <=( A302  and  (not A301) );
 a77167a <=( a77166a  and  a77163a );
 a77168a <=( a77167a  and  a77160a );
 a77172a <=( (not A168)  and  (not A169) );
 a77173a <=( (not A170)  and  a77172a );
 a77176a <=( A166  and  (not A167) );
 a77179a <=( (not A200)  and  (not A199) );
 a77180a <=( a77179a  and  a77176a );
 a77181a <=( a77180a  and  a77173a );
 a77185a <=( A298  and  (not A269) );
 a77186a <=( (not A267)  and  a77185a );
 a77189a <=( (not A300)  and  (not A299) );
 a77192a <=( A302  and  (not A301) );
 a77193a <=( a77192a  and  a77189a );
 a77194a <=( a77193a  and  a77186a );
 a77198a <=( (not A168)  and  (not A169) );
 a77199a <=( (not A170)  and  a77198a );
 a77202a <=( A166  and  (not A167) );
 a77205a <=( (not A200)  and  (not A199) );
 a77206a <=( a77205a  and  a77202a );
 a77207a <=( a77206a  and  a77199a );
 a77211a <=( (not A298)  and  (not A269) );
 a77212a <=( (not A267)  and  a77211a );
 a77215a <=( (not A300)  and  A299 );
 a77218a <=( A302  and  (not A301) );
 a77219a <=( a77218a  and  a77215a );
 a77220a <=( a77219a  and  a77212a );
 a77224a <=( (not A168)  and  (not A169) );
 a77225a <=( (not A170)  and  a77224a );
 a77228a <=( A166  and  (not A167) );
 a77231a <=( (not A200)  and  (not A199) );
 a77232a <=( a77231a  and  a77228a );
 a77233a <=( a77232a  and  a77225a );
 a77237a <=( A298  and  A266 );
 a77238a <=( A265  and  a77237a );
 a77241a <=( (not A300)  and  (not A299) );
 a77244a <=( A302  and  (not A301) );
 a77245a <=( a77244a  and  a77241a );
 a77246a <=( a77245a  and  a77238a );
 a77250a <=( (not A168)  and  (not A169) );
 a77251a <=( (not A170)  and  a77250a );
 a77254a <=( A166  and  (not A167) );
 a77257a <=( (not A200)  and  (not A199) );
 a77258a <=( a77257a  and  a77254a );
 a77259a <=( a77258a  and  a77251a );
 a77263a <=( (not A298)  and  A266 );
 a77264a <=( A265  and  a77263a );
 a77267a <=( (not A300)  and  A299 );
 a77270a <=( A302  and  (not A301) );
 a77271a <=( a77270a  and  a77267a );
 a77272a <=( a77271a  and  a77264a );
 a77276a <=( (not A168)  and  (not A169) );
 a77277a <=( (not A170)  and  a77276a );
 a77280a <=( A166  and  (not A167) );
 a77283a <=( (not A200)  and  (not A199) );
 a77284a <=( a77283a  and  a77280a );
 a77285a <=( a77284a  and  a77277a );
 a77289a <=( A267  and  A266 );
 a77290a <=( (not A265)  and  a77289a );
 a77293a <=( A300  and  A268 );
 a77296a <=( A302  and  (not A301) );
 a77297a <=( a77296a  and  a77293a );
 a77298a <=( a77297a  and  a77290a );
 a77302a <=( (not A168)  and  (not A169) );
 a77303a <=( (not A170)  and  a77302a );
 a77306a <=( A166  and  (not A167) );
 a77309a <=( (not A200)  and  (not A199) );
 a77310a <=( a77309a  and  a77306a );
 a77311a <=( a77310a  and  a77303a );
 a77315a <=( A267  and  A266 );
 a77316a <=( (not A265)  and  a77315a );
 a77319a <=( A300  and  (not A269) );
 a77322a <=( A302  and  (not A301) );
 a77323a <=( a77322a  and  a77319a );
 a77324a <=( a77323a  and  a77316a );
 a77328a <=( (not A168)  and  (not A169) );
 a77329a <=( (not A170)  and  a77328a );
 a77332a <=( A166  and  (not A167) );
 a77335a <=( (not A200)  and  (not A199) );
 a77336a <=( a77335a  and  a77332a );
 a77337a <=( a77336a  and  a77329a );
 a77341a <=( (not A267)  and  A266 );
 a77342a <=( (not A265)  and  a77341a );
 a77345a <=( A269  and  (not A268) );
 a77348a <=( A301  and  (not A300) );
 a77349a <=( a77348a  and  a77345a );
 a77350a <=( a77349a  and  a77342a );
 a77354a <=( (not A168)  and  (not A169) );
 a77355a <=( (not A170)  and  a77354a );
 a77358a <=( A166  and  (not A167) );
 a77361a <=( (not A200)  and  (not A199) );
 a77362a <=( a77361a  and  a77358a );
 a77363a <=( a77362a  and  a77355a );
 a77367a <=( (not A267)  and  A266 );
 a77368a <=( (not A265)  and  a77367a );
 a77371a <=( A269  and  (not A268) );
 a77374a <=( (not A302)  and  (not A300) );
 a77375a <=( a77374a  and  a77371a );
 a77376a <=( a77375a  and  a77368a );
 a77380a <=( (not A168)  and  (not A169) );
 a77381a <=( (not A170)  and  a77380a );
 a77384a <=( A166  and  (not A167) );
 a77387a <=( (not A200)  and  (not A199) );
 a77388a <=( a77387a  and  a77384a );
 a77389a <=( a77388a  and  a77381a );
 a77393a <=( (not A267)  and  A266 );
 a77394a <=( (not A265)  and  a77393a );
 a77397a <=( A269  and  (not A268) );
 a77400a <=( A299  and  A298 );
 a77401a <=( a77400a  and  a77397a );
 a77402a <=( a77401a  and  a77394a );
 a77406a <=( (not A168)  and  (not A169) );
 a77407a <=( (not A170)  and  a77406a );
 a77410a <=( A166  and  (not A167) );
 a77413a <=( (not A200)  and  (not A199) );
 a77414a <=( a77413a  and  a77410a );
 a77415a <=( a77414a  and  a77407a );
 a77419a <=( (not A267)  and  A266 );
 a77420a <=( (not A265)  and  a77419a );
 a77423a <=( A269  and  (not A268) );
 a77426a <=( (not A299)  and  (not A298) );
 a77427a <=( a77426a  and  a77423a );
 a77428a <=( a77427a  and  a77420a );
 a77432a <=( (not A168)  and  (not A169) );
 a77433a <=( (not A170)  and  a77432a );
 a77436a <=( A166  and  (not A167) );
 a77439a <=( (not A200)  and  (not A199) );
 a77440a <=( a77439a  and  a77436a );
 a77441a <=( a77440a  and  a77433a );
 a77445a <=( A267  and  (not A266) );
 a77446a <=( A265  and  a77445a );
 a77449a <=( A300  and  A268 );
 a77452a <=( A302  and  (not A301) );
 a77453a <=( a77452a  and  a77449a );
 a77454a <=( a77453a  and  a77446a );
 a77458a <=( (not A168)  and  (not A169) );
 a77459a <=( (not A170)  and  a77458a );
 a77462a <=( A166  and  (not A167) );
 a77465a <=( (not A200)  and  (not A199) );
 a77466a <=( a77465a  and  a77462a );
 a77467a <=( a77466a  and  a77459a );
 a77471a <=( A267  and  (not A266) );
 a77472a <=( A265  and  a77471a );
 a77475a <=( A300  and  (not A269) );
 a77478a <=( A302  and  (not A301) );
 a77479a <=( a77478a  and  a77475a );
 a77480a <=( a77479a  and  a77472a );
 a77484a <=( (not A168)  and  (not A169) );
 a77485a <=( (not A170)  and  a77484a );
 a77488a <=( A166  and  (not A167) );
 a77491a <=( (not A200)  and  (not A199) );
 a77492a <=( a77491a  and  a77488a );
 a77493a <=( a77492a  and  a77485a );
 a77497a <=( (not A267)  and  (not A266) );
 a77498a <=( A265  and  a77497a );
 a77501a <=( A269  and  (not A268) );
 a77504a <=( A301  and  (not A300) );
 a77505a <=( a77504a  and  a77501a );
 a77506a <=( a77505a  and  a77498a );
 a77510a <=( (not A168)  and  (not A169) );
 a77511a <=( (not A170)  and  a77510a );
 a77514a <=( A166  and  (not A167) );
 a77517a <=( (not A200)  and  (not A199) );
 a77518a <=( a77517a  and  a77514a );
 a77519a <=( a77518a  and  a77511a );
 a77523a <=( (not A267)  and  (not A266) );
 a77524a <=( A265  and  a77523a );
 a77527a <=( A269  and  (not A268) );
 a77530a <=( (not A302)  and  (not A300) );
 a77531a <=( a77530a  and  a77527a );
 a77532a <=( a77531a  and  a77524a );
 a77536a <=( (not A168)  and  (not A169) );
 a77537a <=( (not A170)  and  a77536a );
 a77540a <=( A166  and  (not A167) );
 a77543a <=( (not A200)  and  (not A199) );
 a77544a <=( a77543a  and  a77540a );
 a77545a <=( a77544a  and  a77537a );
 a77549a <=( (not A267)  and  (not A266) );
 a77550a <=( A265  and  a77549a );
 a77553a <=( A269  and  (not A268) );
 a77556a <=( A299  and  A298 );
 a77557a <=( a77556a  and  a77553a );
 a77558a <=( a77557a  and  a77550a );
 a77562a <=( (not A168)  and  (not A169) );
 a77563a <=( (not A170)  and  a77562a );
 a77566a <=( A166  and  (not A167) );
 a77569a <=( (not A200)  and  (not A199) );
 a77570a <=( a77569a  and  a77566a );
 a77571a <=( a77570a  and  a77563a );
 a77575a <=( (not A267)  and  (not A266) );
 a77576a <=( A265  and  a77575a );
 a77579a <=( A269  and  (not A268) );
 a77582a <=( (not A299)  and  (not A298) );
 a77583a <=( a77582a  and  a77579a );
 a77584a <=( a77583a  and  a77576a );
 a77588a <=( (not A168)  and  (not A169) );
 a77589a <=( (not A170)  and  a77588a );
 a77592a <=( A166  and  (not A167) );
 a77595a <=( (not A200)  and  (not A199) );
 a77596a <=( a77595a  and  a77592a );
 a77597a <=( a77596a  and  a77589a );
 a77601a <=( A298  and  (not A266) );
 a77602a <=( (not A265)  and  a77601a );
 a77605a <=( (not A300)  and  (not A299) );
 a77608a <=( A302  and  (not A301) );
 a77609a <=( a77608a  and  a77605a );
 a77610a <=( a77609a  and  a77602a );
 a77614a <=( (not A168)  and  (not A169) );
 a77615a <=( (not A170)  and  a77614a );
 a77618a <=( A166  and  (not A167) );
 a77621a <=( (not A200)  and  (not A199) );
 a77622a <=( a77621a  and  a77618a );
 a77623a <=( a77622a  and  a77615a );
 a77627a <=( (not A298)  and  (not A266) );
 a77628a <=( (not A265)  and  a77627a );
 a77631a <=( (not A300)  and  A299 );
 a77634a <=( A302  and  (not A301) );
 a77635a <=( a77634a  and  a77631a );
 a77636a <=( a77635a  and  a77628a );
 a77640a <=( (not A199)  and  A166 );
 a77641a <=( A167  and  a77640a );
 a77644a <=( A201  and  A200 );
 a77647a <=( (not A265)  and  A202 );
 a77648a <=( a77647a  and  a77644a );
 a77649a <=( a77648a  and  a77641a );
 a77652a <=( A267  and  A266 );
 a77655a <=( A298  and  A268 );
 a77656a <=( a77655a  and  a77652a );
 a77659a <=( (not A300)  and  (not A299) );
 a77662a <=( A302  and  (not A301) );
 a77663a <=( a77662a  and  a77659a );
 a77664a <=( a77663a  and  a77656a );
 a77668a <=( (not A199)  and  A166 );
 a77669a <=( A167  and  a77668a );
 a77672a <=( A201  and  A200 );
 a77675a <=( (not A265)  and  A202 );
 a77676a <=( a77675a  and  a77672a );
 a77677a <=( a77676a  and  a77669a );
 a77680a <=( A267  and  A266 );
 a77683a <=( (not A298)  and  A268 );
 a77684a <=( a77683a  and  a77680a );
 a77687a <=( (not A300)  and  A299 );
 a77690a <=( A302  and  (not A301) );
 a77691a <=( a77690a  and  a77687a );
 a77692a <=( a77691a  and  a77684a );
 a77696a <=( (not A199)  and  A166 );
 a77697a <=( A167  and  a77696a );
 a77700a <=( A201  and  A200 );
 a77703a <=( (not A265)  and  A202 );
 a77704a <=( a77703a  and  a77700a );
 a77705a <=( a77704a  and  a77697a );
 a77708a <=( A267  and  A266 );
 a77711a <=( A298  and  (not A269) );
 a77712a <=( a77711a  and  a77708a );
 a77715a <=( (not A300)  and  (not A299) );
 a77718a <=( A302  and  (not A301) );
 a77719a <=( a77718a  and  a77715a );
 a77720a <=( a77719a  and  a77712a );
 a77724a <=( (not A199)  and  A166 );
 a77725a <=( A167  and  a77724a );
 a77728a <=( A201  and  A200 );
 a77731a <=( (not A265)  and  A202 );
 a77732a <=( a77731a  and  a77728a );
 a77733a <=( a77732a  and  a77725a );
 a77736a <=( A267  and  A266 );
 a77739a <=( (not A298)  and  (not A269) );
 a77740a <=( a77739a  and  a77736a );
 a77743a <=( (not A300)  and  A299 );
 a77746a <=( A302  and  (not A301) );
 a77747a <=( a77746a  and  a77743a );
 a77748a <=( a77747a  and  a77740a );
 a77752a <=( (not A199)  and  A166 );
 a77753a <=( A167  and  a77752a );
 a77756a <=( A201  and  A200 );
 a77759a <=( (not A265)  and  A202 );
 a77760a <=( a77759a  and  a77756a );
 a77761a <=( a77760a  and  a77753a );
 a77764a <=( (not A267)  and  A266 );
 a77767a <=( A269  and  (not A268) );
 a77768a <=( a77767a  and  a77764a );
 a77771a <=( (not A299)  and  A298 );
 a77774a <=( A301  and  A300 );
 a77775a <=( a77774a  and  a77771a );
 a77776a <=( a77775a  and  a77768a );
 a77780a <=( (not A199)  and  A166 );
 a77781a <=( A167  and  a77780a );
 a77784a <=( A201  and  A200 );
 a77787a <=( (not A265)  and  A202 );
 a77788a <=( a77787a  and  a77784a );
 a77789a <=( a77788a  and  a77781a );
 a77792a <=( (not A267)  and  A266 );
 a77795a <=( A269  and  (not A268) );
 a77796a <=( a77795a  and  a77792a );
 a77799a <=( (not A299)  and  A298 );
 a77802a <=( (not A302)  and  A300 );
 a77803a <=( a77802a  and  a77799a );
 a77804a <=( a77803a  and  a77796a );
 a77808a <=( (not A199)  and  A166 );
 a77809a <=( A167  and  a77808a );
 a77812a <=( A201  and  A200 );
 a77815a <=( (not A265)  and  A202 );
 a77816a <=( a77815a  and  a77812a );
 a77817a <=( a77816a  and  a77809a );
 a77820a <=( (not A267)  and  A266 );
 a77823a <=( A269  and  (not A268) );
 a77824a <=( a77823a  and  a77820a );
 a77827a <=( A299  and  (not A298) );
 a77830a <=( A301  and  A300 );
 a77831a <=( a77830a  and  a77827a );
 a77832a <=( a77831a  and  a77824a );
 a77836a <=( (not A199)  and  A166 );
 a77837a <=( A167  and  a77836a );
 a77840a <=( A201  and  A200 );
 a77843a <=( (not A265)  and  A202 );
 a77844a <=( a77843a  and  a77840a );
 a77845a <=( a77844a  and  a77837a );
 a77848a <=( (not A267)  and  A266 );
 a77851a <=( A269  and  (not A268) );
 a77852a <=( a77851a  and  a77848a );
 a77855a <=( A299  and  (not A298) );
 a77858a <=( (not A302)  and  A300 );
 a77859a <=( a77858a  and  a77855a );
 a77860a <=( a77859a  and  a77852a );
 a77864a <=( (not A199)  and  A166 );
 a77865a <=( A167  and  a77864a );
 a77868a <=( A201  and  A200 );
 a77871a <=( A265  and  A202 );
 a77872a <=( a77871a  and  a77868a );
 a77873a <=( a77872a  and  a77865a );
 a77876a <=( A267  and  (not A266) );
 a77879a <=( A298  and  A268 );
 a77880a <=( a77879a  and  a77876a );
 a77883a <=( (not A300)  and  (not A299) );
 a77886a <=( A302  and  (not A301) );
 a77887a <=( a77886a  and  a77883a );
 a77888a <=( a77887a  and  a77880a );
 a77892a <=( (not A199)  and  A166 );
 a77893a <=( A167  and  a77892a );
 a77896a <=( A201  and  A200 );
 a77899a <=( A265  and  A202 );
 a77900a <=( a77899a  and  a77896a );
 a77901a <=( a77900a  and  a77893a );
 a77904a <=( A267  and  (not A266) );
 a77907a <=( (not A298)  and  A268 );
 a77908a <=( a77907a  and  a77904a );
 a77911a <=( (not A300)  and  A299 );
 a77914a <=( A302  and  (not A301) );
 a77915a <=( a77914a  and  a77911a );
 a77916a <=( a77915a  and  a77908a );
 a77920a <=( (not A199)  and  A166 );
 a77921a <=( A167  and  a77920a );
 a77924a <=( A201  and  A200 );
 a77927a <=( A265  and  A202 );
 a77928a <=( a77927a  and  a77924a );
 a77929a <=( a77928a  and  a77921a );
 a77932a <=( A267  and  (not A266) );
 a77935a <=( A298  and  (not A269) );
 a77936a <=( a77935a  and  a77932a );
 a77939a <=( (not A300)  and  (not A299) );
 a77942a <=( A302  and  (not A301) );
 a77943a <=( a77942a  and  a77939a );
 a77944a <=( a77943a  and  a77936a );
 a77948a <=( (not A199)  and  A166 );
 a77949a <=( A167  and  a77948a );
 a77952a <=( A201  and  A200 );
 a77955a <=( A265  and  A202 );
 a77956a <=( a77955a  and  a77952a );
 a77957a <=( a77956a  and  a77949a );
 a77960a <=( A267  and  (not A266) );
 a77963a <=( (not A298)  and  (not A269) );
 a77964a <=( a77963a  and  a77960a );
 a77967a <=( (not A300)  and  A299 );
 a77970a <=( A302  and  (not A301) );
 a77971a <=( a77970a  and  a77967a );
 a77972a <=( a77971a  and  a77964a );
 a77976a <=( (not A199)  and  A166 );
 a77977a <=( A167  and  a77976a );
 a77980a <=( A201  and  A200 );
 a77983a <=( A265  and  A202 );
 a77984a <=( a77983a  and  a77980a );
 a77985a <=( a77984a  and  a77977a );
 a77988a <=( (not A267)  and  (not A266) );
 a77991a <=( A269  and  (not A268) );
 a77992a <=( a77991a  and  a77988a );
 a77995a <=( (not A299)  and  A298 );
 a77998a <=( A301  and  A300 );
 a77999a <=( a77998a  and  a77995a );
 a78000a <=( a77999a  and  a77992a );
 a78004a <=( (not A199)  and  A166 );
 a78005a <=( A167  and  a78004a );
 a78008a <=( A201  and  A200 );
 a78011a <=( A265  and  A202 );
 a78012a <=( a78011a  and  a78008a );
 a78013a <=( a78012a  and  a78005a );
 a78016a <=( (not A267)  and  (not A266) );
 a78019a <=( A269  and  (not A268) );
 a78020a <=( a78019a  and  a78016a );
 a78023a <=( (not A299)  and  A298 );
 a78026a <=( (not A302)  and  A300 );
 a78027a <=( a78026a  and  a78023a );
 a78028a <=( a78027a  and  a78020a );
 a78032a <=( (not A199)  and  A166 );
 a78033a <=( A167  and  a78032a );
 a78036a <=( A201  and  A200 );
 a78039a <=( A265  and  A202 );
 a78040a <=( a78039a  and  a78036a );
 a78041a <=( a78040a  and  a78033a );
 a78044a <=( (not A267)  and  (not A266) );
 a78047a <=( A269  and  (not A268) );
 a78048a <=( a78047a  and  a78044a );
 a78051a <=( A299  and  (not A298) );
 a78054a <=( A301  and  A300 );
 a78055a <=( a78054a  and  a78051a );
 a78056a <=( a78055a  and  a78048a );
 a78060a <=( (not A199)  and  A166 );
 a78061a <=( A167  and  a78060a );
 a78064a <=( A201  and  A200 );
 a78067a <=( A265  and  A202 );
 a78068a <=( a78067a  and  a78064a );
 a78069a <=( a78068a  and  a78061a );
 a78072a <=( (not A267)  and  (not A266) );
 a78075a <=( A269  and  (not A268) );
 a78076a <=( a78075a  and  a78072a );
 a78079a <=( A299  and  (not A298) );
 a78082a <=( (not A302)  and  A300 );
 a78083a <=( a78082a  and  a78079a );
 a78084a <=( a78083a  and  a78076a );
 a78088a <=( (not A199)  and  A166 );
 a78089a <=( A167  and  a78088a );
 a78092a <=( A201  and  A200 );
 a78095a <=( (not A265)  and  (not A203) );
 a78096a <=( a78095a  and  a78092a );
 a78097a <=( a78096a  and  a78089a );
 a78100a <=( A267  and  A266 );
 a78103a <=( A298  and  A268 );
 a78104a <=( a78103a  and  a78100a );
 a78107a <=( (not A300)  and  (not A299) );
 a78110a <=( A302  and  (not A301) );
 a78111a <=( a78110a  and  a78107a );
 a78112a <=( a78111a  and  a78104a );
 a78116a <=( (not A199)  and  A166 );
 a78117a <=( A167  and  a78116a );
 a78120a <=( A201  and  A200 );
 a78123a <=( (not A265)  and  (not A203) );
 a78124a <=( a78123a  and  a78120a );
 a78125a <=( a78124a  and  a78117a );
 a78128a <=( A267  and  A266 );
 a78131a <=( (not A298)  and  A268 );
 a78132a <=( a78131a  and  a78128a );
 a78135a <=( (not A300)  and  A299 );
 a78138a <=( A302  and  (not A301) );
 a78139a <=( a78138a  and  a78135a );
 a78140a <=( a78139a  and  a78132a );
 a78144a <=( (not A199)  and  A166 );
 a78145a <=( A167  and  a78144a );
 a78148a <=( A201  and  A200 );
 a78151a <=( (not A265)  and  (not A203) );
 a78152a <=( a78151a  and  a78148a );
 a78153a <=( a78152a  and  a78145a );
 a78156a <=( A267  and  A266 );
 a78159a <=( A298  and  (not A269) );
 a78160a <=( a78159a  and  a78156a );
 a78163a <=( (not A300)  and  (not A299) );
 a78166a <=( A302  and  (not A301) );
 a78167a <=( a78166a  and  a78163a );
 a78168a <=( a78167a  and  a78160a );
 a78172a <=( (not A199)  and  A166 );
 a78173a <=( A167  and  a78172a );
 a78176a <=( A201  and  A200 );
 a78179a <=( (not A265)  and  (not A203) );
 a78180a <=( a78179a  and  a78176a );
 a78181a <=( a78180a  and  a78173a );
 a78184a <=( A267  and  A266 );
 a78187a <=( (not A298)  and  (not A269) );
 a78188a <=( a78187a  and  a78184a );
 a78191a <=( (not A300)  and  A299 );
 a78194a <=( A302  and  (not A301) );
 a78195a <=( a78194a  and  a78191a );
 a78196a <=( a78195a  and  a78188a );
 a78200a <=( (not A199)  and  A166 );
 a78201a <=( A167  and  a78200a );
 a78204a <=( A201  and  A200 );
 a78207a <=( (not A265)  and  (not A203) );
 a78208a <=( a78207a  and  a78204a );
 a78209a <=( a78208a  and  a78201a );
 a78212a <=( (not A267)  and  A266 );
 a78215a <=( A269  and  (not A268) );
 a78216a <=( a78215a  and  a78212a );
 a78219a <=( (not A299)  and  A298 );
 a78222a <=( A301  and  A300 );
 a78223a <=( a78222a  and  a78219a );
 a78224a <=( a78223a  and  a78216a );
 a78228a <=( (not A199)  and  A166 );
 a78229a <=( A167  and  a78228a );
 a78232a <=( A201  and  A200 );
 a78235a <=( (not A265)  and  (not A203) );
 a78236a <=( a78235a  and  a78232a );
 a78237a <=( a78236a  and  a78229a );
 a78240a <=( (not A267)  and  A266 );
 a78243a <=( A269  and  (not A268) );
 a78244a <=( a78243a  and  a78240a );
 a78247a <=( (not A299)  and  A298 );
 a78250a <=( (not A302)  and  A300 );
 a78251a <=( a78250a  and  a78247a );
 a78252a <=( a78251a  and  a78244a );
 a78256a <=( (not A199)  and  A166 );
 a78257a <=( A167  and  a78256a );
 a78260a <=( A201  and  A200 );
 a78263a <=( (not A265)  and  (not A203) );
 a78264a <=( a78263a  and  a78260a );
 a78265a <=( a78264a  and  a78257a );
 a78268a <=( (not A267)  and  A266 );
 a78271a <=( A269  and  (not A268) );
 a78272a <=( a78271a  and  a78268a );
 a78275a <=( A299  and  (not A298) );
 a78278a <=( A301  and  A300 );
 a78279a <=( a78278a  and  a78275a );
 a78280a <=( a78279a  and  a78272a );
 a78284a <=( (not A199)  and  A166 );
 a78285a <=( A167  and  a78284a );
 a78288a <=( A201  and  A200 );
 a78291a <=( (not A265)  and  (not A203) );
 a78292a <=( a78291a  and  a78288a );
 a78293a <=( a78292a  and  a78285a );
 a78296a <=( (not A267)  and  A266 );
 a78299a <=( A269  and  (not A268) );
 a78300a <=( a78299a  and  a78296a );
 a78303a <=( A299  and  (not A298) );
 a78306a <=( (not A302)  and  A300 );
 a78307a <=( a78306a  and  a78303a );
 a78308a <=( a78307a  and  a78300a );
 a78312a <=( (not A199)  and  A166 );
 a78313a <=( A167  and  a78312a );
 a78316a <=( A201  and  A200 );
 a78319a <=( A265  and  (not A203) );
 a78320a <=( a78319a  and  a78316a );
 a78321a <=( a78320a  and  a78313a );
 a78324a <=( A267  and  (not A266) );
 a78327a <=( A298  and  A268 );
 a78328a <=( a78327a  and  a78324a );
 a78331a <=( (not A300)  and  (not A299) );
 a78334a <=( A302  and  (not A301) );
 a78335a <=( a78334a  and  a78331a );
 a78336a <=( a78335a  and  a78328a );
 a78340a <=( (not A199)  and  A166 );
 a78341a <=( A167  and  a78340a );
 a78344a <=( A201  and  A200 );
 a78347a <=( A265  and  (not A203) );
 a78348a <=( a78347a  and  a78344a );
 a78349a <=( a78348a  and  a78341a );
 a78352a <=( A267  and  (not A266) );
 a78355a <=( (not A298)  and  A268 );
 a78356a <=( a78355a  and  a78352a );
 a78359a <=( (not A300)  and  A299 );
 a78362a <=( A302  and  (not A301) );
 a78363a <=( a78362a  and  a78359a );
 a78364a <=( a78363a  and  a78356a );
 a78368a <=( (not A199)  and  A166 );
 a78369a <=( A167  and  a78368a );
 a78372a <=( A201  and  A200 );
 a78375a <=( A265  and  (not A203) );
 a78376a <=( a78375a  and  a78372a );
 a78377a <=( a78376a  and  a78369a );
 a78380a <=( A267  and  (not A266) );
 a78383a <=( A298  and  (not A269) );
 a78384a <=( a78383a  and  a78380a );
 a78387a <=( (not A300)  and  (not A299) );
 a78390a <=( A302  and  (not A301) );
 a78391a <=( a78390a  and  a78387a );
 a78392a <=( a78391a  and  a78384a );
 a78396a <=( (not A199)  and  A166 );
 a78397a <=( A167  and  a78396a );
 a78400a <=( A201  and  A200 );
 a78403a <=( A265  and  (not A203) );
 a78404a <=( a78403a  and  a78400a );
 a78405a <=( a78404a  and  a78397a );
 a78408a <=( A267  and  (not A266) );
 a78411a <=( (not A298)  and  (not A269) );
 a78412a <=( a78411a  and  a78408a );
 a78415a <=( (not A300)  and  A299 );
 a78418a <=( A302  and  (not A301) );
 a78419a <=( a78418a  and  a78415a );
 a78420a <=( a78419a  and  a78412a );
 a78424a <=( (not A199)  and  A166 );
 a78425a <=( A167  and  a78424a );
 a78428a <=( A201  and  A200 );
 a78431a <=( A265  and  (not A203) );
 a78432a <=( a78431a  and  a78428a );
 a78433a <=( a78432a  and  a78425a );
 a78436a <=( (not A267)  and  (not A266) );
 a78439a <=( A269  and  (not A268) );
 a78440a <=( a78439a  and  a78436a );
 a78443a <=( (not A299)  and  A298 );
 a78446a <=( A301  and  A300 );
 a78447a <=( a78446a  and  a78443a );
 a78448a <=( a78447a  and  a78440a );
 a78452a <=( (not A199)  and  A166 );
 a78453a <=( A167  and  a78452a );
 a78456a <=( A201  and  A200 );
 a78459a <=( A265  and  (not A203) );
 a78460a <=( a78459a  and  a78456a );
 a78461a <=( a78460a  and  a78453a );
 a78464a <=( (not A267)  and  (not A266) );
 a78467a <=( A269  and  (not A268) );
 a78468a <=( a78467a  and  a78464a );
 a78471a <=( (not A299)  and  A298 );
 a78474a <=( (not A302)  and  A300 );
 a78475a <=( a78474a  and  a78471a );
 a78476a <=( a78475a  and  a78468a );
 a78480a <=( (not A199)  and  A166 );
 a78481a <=( A167  and  a78480a );
 a78484a <=( A201  and  A200 );
 a78487a <=( A265  and  (not A203) );
 a78488a <=( a78487a  and  a78484a );
 a78489a <=( a78488a  and  a78481a );
 a78492a <=( (not A267)  and  (not A266) );
 a78495a <=( A269  and  (not A268) );
 a78496a <=( a78495a  and  a78492a );
 a78499a <=( A299  and  (not A298) );
 a78502a <=( A301  and  A300 );
 a78503a <=( a78502a  and  a78499a );
 a78504a <=( a78503a  and  a78496a );
 a78508a <=( (not A199)  and  A166 );
 a78509a <=( A167  and  a78508a );
 a78512a <=( A201  and  A200 );
 a78515a <=( A265  and  (not A203) );
 a78516a <=( a78515a  and  a78512a );
 a78517a <=( a78516a  and  a78509a );
 a78520a <=( (not A267)  and  (not A266) );
 a78523a <=( A269  and  (not A268) );
 a78524a <=( a78523a  and  a78520a );
 a78527a <=( A299  and  (not A298) );
 a78530a <=( (not A302)  and  A300 );
 a78531a <=( a78530a  and  a78527a );
 a78532a <=( a78531a  and  a78524a );
 a78536a <=( (not A199)  and  A166 );
 a78537a <=( A167  and  a78536a );
 a78540a <=( (not A201)  and  A200 );
 a78543a <=( A203  and  (not A202) );
 a78544a <=( a78543a  and  a78540a );
 a78545a <=( a78544a  and  a78537a );
 a78548a <=( A266  and  (not A265) );
 a78551a <=( A268  and  A267 );
 a78552a <=( a78551a  and  a78548a );
 a78555a <=( (not A299)  and  A298 );
 a78558a <=( A301  and  A300 );
 a78559a <=( a78558a  and  a78555a );
 a78560a <=( a78559a  and  a78552a );
 a78564a <=( (not A199)  and  A166 );
 a78565a <=( A167  and  a78564a );
 a78568a <=( (not A201)  and  A200 );
 a78571a <=( A203  and  (not A202) );
 a78572a <=( a78571a  and  a78568a );
 a78573a <=( a78572a  and  a78565a );
 a78576a <=( A266  and  (not A265) );
 a78579a <=( A268  and  A267 );
 a78580a <=( a78579a  and  a78576a );
 a78583a <=( (not A299)  and  A298 );
 a78586a <=( (not A302)  and  A300 );
 a78587a <=( a78586a  and  a78583a );
 a78588a <=( a78587a  and  a78580a );
 a78592a <=( (not A199)  and  A166 );
 a78593a <=( A167  and  a78592a );
 a78596a <=( (not A201)  and  A200 );
 a78599a <=( A203  and  (not A202) );
 a78600a <=( a78599a  and  a78596a );
 a78601a <=( a78600a  and  a78593a );
 a78604a <=( A266  and  (not A265) );
 a78607a <=( A268  and  A267 );
 a78608a <=( a78607a  and  a78604a );
 a78611a <=( A299  and  (not A298) );
 a78614a <=( A301  and  A300 );
 a78615a <=( a78614a  and  a78611a );
 a78616a <=( a78615a  and  a78608a );
 a78620a <=( (not A199)  and  A166 );
 a78621a <=( A167  and  a78620a );
 a78624a <=( (not A201)  and  A200 );
 a78627a <=( A203  and  (not A202) );
 a78628a <=( a78627a  and  a78624a );
 a78629a <=( a78628a  and  a78621a );
 a78632a <=( A266  and  (not A265) );
 a78635a <=( A268  and  A267 );
 a78636a <=( a78635a  and  a78632a );
 a78639a <=( A299  and  (not A298) );
 a78642a <=( (not A302)  and  A300 );
 a78643a <=( a78642a  and  a78639a );
 a78644a <=( a78643a  and  a78636a );
 a78648a <=( (not A199)  and  A166 );
 a78649a <=( A167  and  a78648a );
 a78652a <=( (not A201)  and  A200 );
 a78655a <=( A203  and  (not A202) );
 a78656a <=( a78655a  and  a78652a );
 a78657a <=( a78656a  and  a78649a );
 a78660a <=( A266  and  (not A265) );
 a78663a <=( (not A269)  and  A267 );
 a78664a <=( a78663a  and  a78660a );
 a78667a <=( (not A299)  and  A298 );
 a78670a <=( A301  and  A300 );
 a78671a <=( a78670a  and  a78667a );
 a78672a <=( a78671a  and  a78664a );
 a78676a <=( (not A199)  and  A166 );
 a78677a <=( A167  and  a78676a );
 a78680a <=( (not A201)  and  A200 );
 a78683a <=( A203  and  (not A202) );
 a78684a <=( a78683a  and  a78680a );
 a78685a <=( a78684a  and  a78677a );
 a78688a <=( A266  and  (not A265) );
 a78691a <=( (not A269)  and  A267 );
 a78692a <=( a78691a  and  a78688a );
 a78695a <=( (not A299)  and  A298 );
 a78698a <=( (not A302)  and  A300 );
 a78699a <=( a78698a  and  a78695a );
 a78700a <=( a78699a  and  a78692a );
 a78704a <=( (not A199)  and  A166 );
 a78705a <=( A167  and  a78704a );
 a78708a <=( (not A201)  and  A200 );
 a78711a <=( A203  and  (not A202) );
 a78712a <=( a78711a  and  a78708a );
 a78713a <=( a78712a  and  a78705a );
 a78716a <=( A266  and  (not A265) );
 a78719a <=( (not A269)  and  A267 );
 a78720a <=( a78719a  and  a78716a );
 a78723a <=( A299  and  (not A298) );
 a78726a <=( A301  and  A300 );
 a78727a <=( a78726a  and  a78723a );
 a78728a <=( a78727a  and  a78720a );
 a78732a <=( (not A199)  and  A166 );
 a78733a <=( A167  and  a78732a );
 a78736a <=( (not A201)  and  A200 );
 a78739a <=( A203  and  (not A202) );
 a78740a <=( a78739a  and  a78736a );
 a78741a <=( a78740a  and  a78733a );
 a78744a <=( A266  and  (not A265) );
 a78747a <=( (not A269)  and  A267 );
 a78748a <=( a78747a  and  a78744a );
 a78751a <=( A299  and  (not A298) );
 a78754a <=( (not A302)  and  A300 );
 a78755a <=( a78754a  and  a78751a );
 a78756a <=( a78755a  and  a78748a );
 a78760a <=( (not A199)  and  A166 );
 a78761a <=( A167  and  a78760a );
 a78764a <=( (not A201)  and  A200 );
 a78767a <=( A203  and  (not A202) );
 a78768a <=( a78767a  and  a78764a );
 a78769a <=( a78768a  and  a78761a );
 a78772a <=( (not A266)  and  A265 );
 a78775a <=( A268  and  A267 );
 a78776a <=( a78775a  and  a78772a );
 a78779a <=( (not A299)  and  A298 );
 a78782a <=( A301  and  A300 );
 a78783a <=( a78782a  and  a78779a );
 a78784a <=( a78783a  and  a78776a );
 a78788a <=( (not A199)  and  A166 );
 a78789a <=( A167  and  a78788a );
 a78792a <=( (not A201)  and  A200 );
 a78795a <=( A203  and  (not A202) );
 a78796a <=( a78795a  and  a78792a );
 a78797a <=( a78796a  and  a78789a );
 a78800a <=( (not A266)  and  A265 );
 a78803a <=( A268  and  A267 );
 a78804a <=( a78803a  and  a78800a );
 a78807a <=( (not A299)  and  A298 );
 a78810a <=( (not A302)  and  A300 );
 a78811a <=( a78810a  and  a78807a );
 a78812a <=( a78811a  and  a78804a );
 a78816a <=( (not A199)  and  A166 );
 a78817a <=( A167  and  a78816a );
 a78820a <=( (not A201)  and  A200 );
 a78823a <=( A203  and  (not A202) );
 a78824a <=( a78823a  and  a78820a );
 a78825a <=( a78824a  and  a78817a );
 a78828a <=( (not A266)  and  A265 );
 a78831a <=( A268  and  A267 );
 a78832a <=( a78831a  and  a78828a );
 a78835a <=( A299  and  (not A298) );
 a78838a <=( A301  and  A300 );
 a78839a <=( a78838a  and  a78835a );
 a78840a <=( a78839a  and  a78832a );
 a78844a <=( (not A199)  and  A166 );
 a78845a <=( A167  and  a78844a );
 a78848a <=( (not A201)  and  A200 );
 a78851a <=( A203  and  (not A202) );
 a78852a <=( a78851a  and  a78848a );
 a78853a <=( a78852a  and  a78845a );
 a78856a <=( (not A266)  and  A265 );
 a78859a <=( A268  and  A267 );
 a78860a <=( a78859a  and  a78856a );
 a78863a <=( A299  and  (not A298) );
 a78866a <=( (not A302)  and  A300 );
 a78867a <=( a78866a  and  a78863a );
 a78868a <=( a78867a  and  a78860a );
 a78872a <=( (not A199)  and  A166 );
 a78873a <=( A167  and  a78872a );
 a78876a <=( (not A201)  and  A200 );
 a78879a <=( A203  and  (not A202) );
 a78880a <=( a78879a  and  a78876a );
 a78881a <=( a78880a  and  a78873a );
 a78884a <=( (not A266)  and  A265 );
 a78887a <=( (not A269)  and  A267 );
 a78888a <=( a78887a  and  a78884a );
 a78891a <=( (not A299)  and  A298 );
 a78894a <=( A301  and  A300 );
 a78895a <=( a78894a  and  a78891a );
 a78896a <=( a78895a  and  a78888a );
 a78900a <=( (not A199)  and  A166 );
 a78901a <=( A167  and  a78900a );
 a78904a <=( (not A201)  and  A200 );
 a78907a <=( A203  and  (not A202) );
 a78908a <=( a78907a  and  a78904a );
 a78909a <=( a78908a  and  a78901a );
 a78912a <=( (not A266)  and  A265 );
 a78915a <=( (not A269)  and  A267 );
 a78916a <=( a78915a  and  a78912a );
 a78919a <=( (not A299)  and  A298 );
 a78922a <=( (not A302)  and  A300 );
 a78923a <=( a78922a  and  a78919a );
 a78924a <=( a78923a  and  a78916a );
 a78928a <=( (not A199)  and  A166 );
 a78929a <=( A167  and  a78928a );
 a78932a <=( (not A201)  and  A200 );
 a78935a <=( A203  and  (not A202) );
 a78936a <=( a78935a  and  a78932a );
 a78937a <=( a78936a  and  a78929a );
 a78940a <=( (not A266)  and  A265 );
 a78943a <=( (not A269)  and  A267 );
 a78944a <=( a78943a  and  a78940a );
 a78947a <=( A299  and  (not A298) );
 a78950a <=( A301  and  A300 );
 a78951a <=( a78950a  and  a78947a );
 a78952a <=( a78951a  and  a78944a );
 a78956a <=( (not A199)  and  A166 );
 a78957a <=( A167  and  a78956a );
 a78960a <=( (not A201)  and  A200 );
 a78963a <=( A203  and  (not A202) );
 a78964a <=( a78963a  and  a78960a );
 a78965a <=( a78964a  and  a78957a );
 a78968a <=( (not A266)  and  A265 );
 a78971a <=( (not A269)  and  A267 );
 a78972a <=( a78971a  and  a78968a );
 a78975a <=( A299  and  (not A298) );
 a78978a <=( (not A302)  and  A300 );
 a78979a <=( a78978a  and  a78975a );
 a78980a <=( a78979a  and  a78972a );
 a78984a <=( A199  and  A166 );
 a78985a <=( A167  and  a78984a );
 a78988a <=( A201  and  (not A200) );
 a78991a <=( (not A265)  and  A202 );
 a78992a <=( a78991a  and  a78988a );
 a78993a <=( a78992a  and  a78985a );
 a78996a <=( A267  and  A266 );
 a78999a <=( A298  and  A268 );
 a79000a <=( a78999a  and  a78996a );
 a79003a <=( (not A300)  and  (not A299) );
 a79006a <=( A302  and  (not A301) );
 a79007a <=( a79006a  and  a79003a );
 a79008a <=( a79007a  and  a79000a );
 a79012a <=( A199  and  A166 );
 a79013a <=( A167  and  a79012a );
 a79016a <=( A201  and  (not A200) );
 a79019a <=( (not A265)  and  A202 );
 a79020a <=( a79019a  and  a79016a );
 a79021a <=( a79020a  and  a79013a );
 a79024a <=( A267  and  A266 );
 a79027a <=( (not A298)  and  A268 );
 a79028a <=( a79027a  and  a79024a );
 a79031a <=( (not A300)  and  A299 );
 a79034a <=( A302  and  (not A301) );
 a79035a <=( a79034a  and  a79031a );
 a79036a <=( a79035a  and  a79028a );
 a79040a <=( A199  and  A166 );
 a79041a <=( A167  and  a79040a );
 a79044a <=( A201  and  (not A200) );
 a79047a <=( (not A265)  and  A202 );
 a79048a <=( a79047a  and  a79044a );
 a79049a <=( a79048a  and  a79041a );
 a79052a <=( A267  and  A266 );
 a79055a <=( A298  and  (not A269) );
 a79056a <=( a79055a  and  a79052a );
 a79059a <=( (not A300)  and  (not A299) );
 a79062a <=( A302  and  (not A301) );
 a79063a <=( a79062a  and  a79059a );
 a79064a <=( a79063a  and  a79056a );
 a79068a <=( A199  and  A166 );
 a79069a <=( A167  and  a79068a );
 a79072a <=( A201  and  (not A200) );
 a79075a <=( (not A265)  and  A202 );
 a79076a <=( a79075a  and  a79072a );
 a79077a <=( a79076a  and  a79069a );
 a79080a <=( A267  and  A266 );
 a79083a <=( (not A298)  and  (not A269) );
 a79084a <=( a79083a  and  a79080a );
 a79087a <=( (not A300)  and  A299 );
 a79090a <=( A302  and  (not A301) );
 a79091a <=( a79090a  and  a79087a );
 a79092a <=( a79091a  and  a79084a );
 a79096a <=( A199  and  A166 );
 a79097a <=( A167  and  a79096a );
 a79100a <=( A201  and  (not A200) );
 a79103a <=( (not A265)  and  A202 );
 a79104a <=( a79103a  and  a79100a );
 a79105a <=( a79104a  and  a79097a );
 a79108a <=( (not A267)  and  A266 );
 a79111a <=( A269  and  (not A268) );
 a79112a <=( a79111a  and  a79108a );
 a79115a <=( (not A299)  and  A298 );
 a79118a <=( A301  and  A300 );
 a79119a <=( a79118a  and  a79115a );
 a79120a <=( a79119a  and  a79112a );
 a79124a <=( A199  and  A166 );
 a79125a <=( A167  and  a79124a );
 a79128a <=( A201  and  (not A200) );
 a79131a <=( (not A265)  and  A202 );
 a79132a <=( a79131a  and  a79128a );
 a79133a <=( a79132a  and  a79125a );
 a79136a <=( (not A267)  and  A266 );
 a79139a <=( A269  and  (not A268) );
 a79140a <=( a79139a  and  a79136a );
 a79143a <=( (not A299)  and  A298 );
 a79146a <=( (not A302)  and  A300 );
 a79147a <=( a79146a  and  a79143a );
 a79148a <=( a79147a  and  a79140a );
 a79152a <=( A199  and  A166 );
 a79153a <=( A167  and  a79152a );
 a79156a <=( A201  and  (not A200) );
 a79159a <=( (not A265)  and  A202 );
 a79160a <=( a79159a  and  a79156a );
 a79161a <=( a79160a  and  a79153a );
 a79164a <=( (not A267)  and  A266 );
 a79167a <=( A269  and  (not A268) );
 a79168a <=( a79167a  and  a79164a );
 a79171a <=( A299  and  (not A298) );
 a79174a <=( A301  and  A300 );
 a79175a <=( a79174a  and  a79171a );
 a79176a <=( a79175a  and  a79168a );
 a79180a <=( A199  and  A166 );
 a79181a <=( A167  and  a79180a );
 a79184a <=( A201  and  (not A200) );
 a79187a <=( (not A265)  and  A202 );
 a79188a <=( a79187a  and  a79184a );
 a79189a <=( a79188a  and  a79181a );
 a79192a <=( (not A267)  and  A266 );
 a79195a <=( A269  and  (not A268) );
 a79196a <=( a79195a  and  a79192a );
 a79199a <=( A299  and  (not A298) );
 a79202a <=( (not A302)  and  A300 );
 a79203a <=( a79202a  and  a79199a );
 a79204a <=( a79203a  and  a79196a );
 a79208a <=( A199  and  A166 );
 a79209a <=( A167  and  a79208a );
 a79212a <=( A201  and  (not A200) );
 a79215a <=( A265  and  A202 );
 a79216a <=( a79215a  and  a79212a );
 a79217a <=( a79216a  and  a79209a );
 a79220a <=( A267  and  (not A266) );
 a79223a <=( A298  and  A268 );
 a79224a <=( a79223a  and  a79220a );
 a79227a <=( (not A300)  and  (not A299) );
 a79230a <=( A302  and  (not A301) );
 a79231a <=( a79230a  and  a79227a );
 a79232a <=( a79231a  and  a79224a );
 a79236a <=( A199  and  A166 );
 a79237a <=( A167  and  a79236a );
 a79240a <=( A201  and  (not A200) );
 a79243a <=( A265  and  A202 );
 a79244a <=( a79243a  and  a79240a );
 a79245a <=( a79244a  and  a79237a );
 a79248a <=( A267  and  (not A266) );
 a79251a <=( (not A298)  and  A268 );
 a79252a <=( a79251a  and  a79248a );
 a79255a <=( (not A300)  and  A299 );
 a79258a <=( A302  and  (not A301) );
 a79259a <=( a79258a  and  a79255a );
 a79260a <=( a79259a  and  a79252a );
 a79264a <=( A199  and  A166 );
 a79265a <=( A167  and  a79264a );
 a79268a <=( A201  and  (not A200) );
 a79271a <=( A265  and  A202 );
 a79272a <=( a79271a  and  a79268a );
 a79273a <=( a79272a  and  a79265a );
 a79276a <=( A267  and  (not A266) );
 a79279a <=( A298  and  (not A269) );
 a79280a <=( a79279a  and  a79276a );
 a79283a <=( (not A300)  and  (not A299) );
 a79286a <=( A302  and  (not A301) );
 a79287a <=( a79286a  and  a79283a );
 a79288a <=( a79287a  and  a79280a );
 a79292a <=( A199  and  A166 );
 a79293a <=( A167  and  a79292a );
 a79296a <=( A201  and  (not A200) );
 a79299a <=( A265  and  A202 );
 a79300a <=( a79299a  and  a79296a );
 a79301a <=( a79300a  and  a79293a );
 a79304a <=( A267  and  (not A266) );
 a79307a <=( (not A298)  and  (not A269) );
 a79308a <=( a79307a  and  a79304a );
 a79311a <=( (not A300)  and  A299 );
 a79314a <=( A302  and  (not A301) );
 a79315a <=( a79314a  and  a79311a );
 a79316a <=( a79315a  and  a79308a );
 a79320a <=( A199  and  A166 );
 a79321a <=( A167  and  a79320a );
 a79324a <=( A201  and  (not A200) );
 a79327a <=( A265  and  A202 );
 a79328a <=( a79327a  and  a79324a );
 a79329a <=( a79328a  and  a79321a );
 a79332a <=( (not A267)  and  (not A266) );
 a79335a <=( A269  and  (not A268) );
 a79336a <=( a79335a  and  a79332a );
 a79339a <=( (not A299)  and  A298 );
 a79342a <=( A301  and  A300 );
 a79343a <=( a79342a  and  a79339a );
 a79344a <=( a79343a  and  a79336a );
 a79348a <=( A199  and  A166 );
 a79349a <=( A167  and  a79348a );
 a79352a <=( A201  and  (not A200) );
 a79355a <=( A265  and  A202 );
 a79356a <=( a79355a  and  a79352a );
 a79357a <=( a79356a  and  a79349a );
 a79360a <=( (not A267)  and  (not A266) );
 a79363a <=( A269  and  (not A268) );
 a79364a <=( a79363a  and  a79360a );
 a79367a <=( (not A299)  and  A298 );
 a79370a <=( (not A302)  and  A300 );
 a79371a <=( a79370a  and  a79367a );
 a79372a <=( a79371a  and  a79364a );
 a79376a <=( A199  and  A166 );
 a79377a <=( A167  and  a79376a );
 a79380a <=( A201  and  (not A200) );
 a79383a <=( A265  and  A202 );
 a79384a <=( a79383a  and  a79380a );
 a79385a <=( a79384a  and  a79377a );
 a79388a <=( (not A267)  and  (not A266) );
 a79391a <=( A269  and  (not A268) );
 a79392a <=( a79391a  and  a79388a );
 a79395a <=( A299  and  (not A298) );
 a79398a <=( A301  and  A300 );
 a79399a <=( a79398a  and  a79395a );
 a79400a <=( a79399a  and  a79392a );
 a79404a <=( A199  and  A166 );
 a79405a <=( A167  and  a79404a );
 a79408a <=( A201  and  (not A200) );
 a79411a <=( A265  and  A202 );
 a79412a <=( a79411a  and  a79408a );
 a79413a <=( a79412a  and  a79405a );
 a79416a <=( (not A267)  and  (not A266) );
 a79419a <=( A269  and  (not A268) );
 a79420a <=( a79419a  and  a79416a );
 a79423a <=( A299  and  (not A298) );
 a79426a <=( (not A302)  and  A300 );
 a79427a <=( a79426a  and  a79423a );
 a79428a <=( a79427a  and  a79420a );
 a79432a <=( A199  and  A166 );
 a79433a <=( A167  and  a79432a );
 a79436a <=( A201  and  (not A200) );
 a79439a <=( (not A265)  and  (not A203) );
 a79440a <=( a79439a  and  a79436a );
 a79441a <=( a79440a  and  a79433a );
 a79444a <=( A267  and  A266 );
 a79447a <=( A298  and  A268 );
 a79448a <=( a79447a  and  a79444a );
 a79451a <=( (not A300)  and  (not A299) );
 a79454a <=( A302  and  (not A301) );
 a79455a <=( a79454a  and  a79451a );
 a79456a <=( a79455a  and  a79448a );
 a79460a <=( A199  and  A166 );
 a79461a <=( A167  and  a79460a );
 a79464a <=( A201  and  (not A200) );
 a79467a <=( (not A265)  and  (not A203) );
 a79468a <=( a79467a  and  a79464a );
 a79469a <=( a79468a  and  a79461a );
 a79472a <=( A267  and  A266 );
 a79475a <=( (not A298)  and  A268 );
 a79476a <=( a79475a  and  a79472a );
 a79479a <=( (not A300)  and  A299 );
 a79482a <=( A302  and  (not A301) );
 a79483a <=( a79482a  and  a79479a );
 a79484a <=( a79483a  and  a79476a );
 a79488a <=( A199  and  A166 );
 a79489a <=( A167  and  a79488a );
 a79492a <=( A201  and  (not A200) );
 a79495a <=( (not A265)  and  (not A203) );
 a79496a <=( a79495a  and  a79492a );
 a79497a <=( a79496a  and  a79489a );
 a79500a <=( A267  and  A266 );
 a79503a <=( A298  and  (not A269) );
 a79504a <=( a79503a  and  a79500a );
 a79507a <=( (not A300)  and  (not A299) );
 a79510a <=( A302  and  (not A301) );
 a79511a <=( a79510a  and  a79507a );
 a79512a <=( a79511a  and  a79504a );
 a79516a <=( A199  and  A166 );
 a79517a <=( A167  and  a79516a );
 a79520a <=( A201  and  (not A200) );
 a79523a <=( (not A265)  and  (not A203) );
 a79524a <=( a79523a  and  a79520a );
 a79525a <=( a79524a  and  a79517a );
 a79528a <=( A267  and  A266 );
 a79531a <=( (not A298)  and  (not A269) );
 a79532a <=( a79531a  and  a79528a );
 a79535a <=( (not A300)  and  A299 );
 a79538a <=( A302  and  (not A301) );
 a79539a <=( a79538a  and  a79535a );
 a79540a <=( a79539a  and  a79532a );
 a79544a <=( A199  and  A166 );
 a79545a <=( A167  and  a79544a );
 a79548a <=( A201  and  (not A200) );
 a79551a <=( (not A265)  and  (not A203) );
 a79552a <=( a79551a  and  a79548a );
 a79553a <=( a79552a  and  a79545a );
 a79556a <=( (not A267)  and  A266 );
 a79559a <=( A269  and  (not A268) );
 a79560a <=( a79559a  and  a79556a );
 a79563a <=( (not A299)  and  A298 );
 a79566a <=( A301  and  A300 );
 a79567a <=( a79566a  and  a79563a );
 a79568a <=( a79567a  and  a79560a );
 a79572a <=( A199  and  A166 );
 a79573a <=( A167  and  a79572a );
 a79576a <=( A201  and  (not A200) );
 a79579a <=( (not A265)  and  (not A203) );
 a79580a <=( a79579a  and  a79576a );
 a79581a <=( a79580a  and  a79573a );
 a79584a <=( (not A267)  and  A266 );
 a79587a <=( A269  and  (not A268) );
 a79588a <=( a79587a  and  a79584a );
 a79591a <=( (not A299)  and  A298 );
 a79594a <=( (not A302)  and  A300 );
 a79595a <=( a79594a  and  a79591a );
 a79596a <=( a79595a  and  a79588a );
 a79600a <=( A199  and  A166 );
 a79601a <=( A167  and  a79600a );
 a79604a <=( A201  and  (not A200) );
 a79607a <=( (not A265)  and  (not A203) );
 a79608a <=( a79607a  and  a79604a );
 a79609a <=( a79608a  and  a79601a );
 a79612a <=( (not A267)  and  A266 );
 a79615a <=( A269  and  (not A268) );
 a79616a <=( a79615a  and  a79612a );
 a79619a <=( A299  and  (not A298) );
 a79622a <=( A301  and  A300 );
 a79623a <=( a79622a  and  a79619a );
 a79624a <=( a79623a  and  a79616a );
 a79628a <=( A199  and  A166 );
 a79629a <=( A167  and  a79628a );
 a79632a <=( A201  and  (not A200) );
 a79635a <=( (not A265)  and  (not A203) );
 a79636a <=( a79635a  and  a79632a );
 a79637a <=( a79636a  and  a79629a );
 a79640a <=( (not A267)  and  A266 );
 a79643a <=( A269  and  (not A268) );
 a79644a <=( a79643a  and  a79640a );
 a79647a <=( A299  and  (not A298) );
 a79650a <=( (not A302)  and  A300 );
 a79651a <=( a79650a  and  a79647a );
 a79652a <=( a79651a  and  a79644a );
 a79656a <=( A199  and  A166 );
 a79657a <=( A167  and  a79656a );
 a79660a <=( A201  and  (not A200) );
 a79663a <=( A265  and  (not A203) );
 a79664a <=( a79663a  and  a79660a );
 a79665a <=( a79664a  and  a79657a );
 a79668a <=( A267  and  (not A266) );
 a79671a <=( A298  and  A268 );
 a79672a <=( a79671a  and  a79668a );
 a79675a <=( (not A300)  and  (not A299) );
 a79678a <=( A302  and  (not A301) );
 a79679a <=( a79678a  and  a79675a );
 a79680a <=( a79679a  and  a79672a );
 a79684a <=( A199  and  A166 );
 a79685a <=( A167  and  a79684a );
 a79688a <=( A201  and  (not A200) );
 a79691a <=( A265  and  (not A203) );
 a79692a <=( a79691a  and  a79688a );
 a79693a <=( a79692a  and  a79685a );
 a79696a <=( A267  and  (not A266) );
 a79699a <=( (not A298)  and  A268 );
 a79700a <=( a79699a  and  a79696a );
 a79703a <=( (not A300)  and  A299 );
 a79706a <=( A302  and  (not A301) );
 a79707a <=( a79706a  and  a79703a );
 a79708a <=( a79707a  and  a79700a );
 a79712a <=( A199  and  A166 );
 a79713a <=( A167  and  a79712a );
 a79716a <=( A201  and  (not A200) );
 a79719a <=( A265  and  (not A203) );
 a79720a <=( a79719a  and  a79716a );
 a79721a <=( a79720a  and  a79713a );
 a79724a <=( A267  and  (not A266) );
 a79727a <=( A298  and  (not A269) );
 a79728a <=( a79727a  and  a79724a );
 a79731a <=( (not A300)  and  (not A299) );
 a79734a <=( A302  and  (not A301) );
 a79735a <=( a79734a  and  a79731a );
 a79736a <=( a79735a  and  a79728a );
 a79740a <=( A199  and  A166 );
 a79741a <=( A167  and  a79740a );
 a79744a <=( A201  and  (not A200) );
 a79747a <=( A265  and  (not A203) );
 a79748a <=( a79747a  and  a79744a );
 a79749a <=( a79748a  and  a79741a );
 a79752a <=( A267  and  (not A266) );
 a79755a <=( (not A298)  and  (not A269) );
 a79756a <=( a79755a  and  a79752a );
 a79759a <=( (not A300)  and  A299 );
 a79762a <=( A302  and  (not A301) );
 a79763a <=( a79762a  and  a79759a );
 a79764a <=( a79763a  and  a79756a );
 a79768a <=( A199  and  A166 );
 a79769a <=( A167  and  a79768a );
 a79772a <=( A201  and  (not A200) );
 a79775a <=( A265  and  (not A203) );
 a79776a <=( a79775a  and  a79772a );
 a79777a <=( a79776a  and  a79769a );
 a79780a <=( (not A267)  and  (not A266) );
 a79783a <=( A269  and  (not A268) );
 a79784a <=( a79783a  and  a79780a );
 a79787a <=( (not A299)  and  A298 );
 a79790a <=( A301  and  A300 );
 a79791a <=( a79790a  and  a79787a );
 a79792a <=( a79791a  and  a79784a );
 a79796a <=( A199  and  A166 );
 a79797a <=( A167  and  a79796a );
 a79800a <=( A201  and  (not A200) );
 a79803a <=( A265  and  (not A203) );
 a79804a <=( a79803a  and  a79800a );
 a79805a <=( a79804a  and  a79797a );
 a79808a <=( (not A267)  and  (not A266) );
 a79811a <=( A269  and  (not A268) );
 a79812a <=( a79811a  and  a79808a );
 a79815a <=( (not A299)  and  A298 );
 a79818a <=( (not A302)  and  A300 );
 a79819a <=( a79818a  and  a79815a );
 a79820a <=( a79819a  and  a79812a );
 a79824a <=( A199  and  A166 );
 a79825a <=( A167  and  a79824a );
 a79828a <=( A201  and  (not A200) );
 a79831a <=( A265  and  (not A203) );
 a79832a <=( a79831a  and  a79828a );
 a79833a <=( a79832a  and  a79825a );
 a79836a <=( (not A267)  and  (not A266) );
 a79839a <=( A269  and  (not A268) );
 a79840a <=( a79839a  and  a79836a );
 a79843a <=( A299  and  (not A298) );
 a79846a <=( A301  and  A300 );
 a79847a <=( a79846a  and  a79843a );
 a79848a <=( a79847a  and  a79840a );
 a79852a <=( A199  and  A166 );
 a79853a <=( A167  and  a79852a );
 a79856a <=( A201  and  (not A200) );
 a79859a <=( A265  and  (not A203) );
 a79860a <=( a79859a  and  a79856a );
 a79861a <=( a79860a  and  a79853a );
 a79864a <=( (not A267)  and  (not A266) );
 a79867a <=( A269  and  (not A268) );
 a79868a <=( a79867a  and  a79864a );
 a79871a <=( A299  and  (not A298) );
 a79874a <=( (not A302)  and  A300 );
 a79875a <=( a79874a  and  a79871a );
 a79876a <=( a79875a  and  a79868a );
 a79880a <=( A199  and  A166 );
 a79881a <=( A167  and  a79880a );
 a79884a <=( (not A201)  and  (not A200) );
 a79887a <=( A203  and  (not A202) );
 a79888a <=( a79887a  and  a79884a );
 a79889a <=( a79888a  and  a79881a );
 a79892a <=( A266  and  (not A265) );
 a79895a <=( A268  and  A267 );
 a79896a <=( a79895a  and  a79892a );
 a79899a <=( (not A299)  and  A298 );
 a79902a <=( A301  and  A300 );
 a79903a <=( a79902a  and  a79899a );
 a79904a <=( a79903a  and  a79896a );
 a79908a <=( A199  and  A166 );
 a79909a <=( A167  and  a79908a );
 a79912a <=( (not A201)  and  (not A200) );
 a79915a <=( A203  and  (not A202) );
 a79916a <=( a79915a  and  a79912a );
 a79917a <=( a79916a  and  a79909a );
 a79920a <=( A266  and  (not A265) );
 a79923a <=( A268  and  A267 );
 a79924a <=( a79923a  and  a79920a );
 a79927a <=( (not A299)  and  A298 );
 a79930a <=( (not A302)  and  A300 );
 a79931a <=( a79930a  and  a79927a );
 a79932a <=( a79931a  and  a79924a );
 a79936a <=( A199  and  A166 );
 a79937a <=( A167  and  a79936a );
 a79940a <=( (not A201)  and  (not A200) );
 a79943a <=( A203  and  (not A202) );
 a79944a <=( a79943a  and  a79940a );
 a79945a <=( a79944a  and  a79937a );
 a79948a <=( A266  and  (not A265) );
 a79951a <=( A268  and  A267 );
 a79952a <=( a79951a  and  a79948a );
 a79955a <=( A299  and  (not A298) );
 a79958a <=( A301  and  A300 );
 a79959a <=( a79958a  and  a79955a );
 a79960a <=( a79959a  and  a79952a );
 a79964a <=( A199  and  A166 );
 a79965a <=( A167  and  a79964a );
 a79968a <=( (not A201)  and  (not A200) );
 a79971a <=( A203  and  (not A202) );
 a79972a <=( a79971a  and  a79968a );
 a79973a <=( a79972a  and  a79965a );
 a79976a <=( A266  and  (not A265) );
 a79979a <=( A268  and  A267 );
 a79980a <=( a79979a  and  a79976a );
 a79983a <=( A299  and  (not A298) );
 a79986a <=( (not A302)  and  A300 );
 a79987a <=( a79986a  and  a79983a );
 a79988a <=( a79987a  and  a79980a );
 a79992a <=( A199  and  A166 );
 a79993a <=( A167  and  a79992a );
 a79996a <=( (not A201)  and  (not A200) );
 a79999a <=( A203  and  (not A202) );
 a80000a <=( a79999a  and  a79996a );
 a80001a <=( a80000a  and  a79993a );
 a80004a <=( A266  and  (not A265) );
 a80007a <=( (not A269)  and  A267 );
 a80008a <=( a80007a  and  a80004a );
 a80011a <=( (not A299)  and  A298 );
 a80014a <=( A301  and  A300 );
 a80015a <=( a80014a  and  a80011a );
 a80016a <=( a80015a  and  a80008a );
 a80020a <=( A199  and  A166 );
 a80021a <=( A167  and  a80020a );
 a80024a <=( (not A201)  and  (not A200) );
 a80027a <=( A203  and  (not A202) );
 a80028a <=( a80027a  and  a80024a );
 a80029a <=( a80028a  and  a80021a );
 a80032a <=( A266  and  (not A265) );
 a80035a <=( (not A269)  and  A267 );
 a80036a <=( a80035a  and  a80032a );
 a80039a <=( (not A299)  and  A298 );
 a80042a <=( (not A302)  and  A300 );
 a80043a <=( a80042a  and  a80039a );
 a80044a <=( a80043a  and  a80036a );
 a80048a <=( A199  and  A166 );
 a80049a <=( A167  and  a80048a );
 a80052a <=( (not A201)  and  (not A200) );
 a80055a <=( A203  and  (not A202) );
 a80056a <=( a80055a  and  a80052a );
 a80057a <=( a80056a  and  a80049a );
 a80060a <=( A266  and  (not A265) );
 a80063a <=( (not A269)  and  A267 );
 a80064a <=( a80063a  and  a80060a );
 a80067a <=( A299  and  (not A298) );
 a80070a <=( A301  and  A300 );
 a80071a <=( a80070a  and  a80067a );
 a80072a <=( a80071a  and  a80064a );
 a80076a <=( A199  and  A166 );
 a80077a <=( A167  and  a80076a );
 a80080a <=( (not A201)  and  (not A200) );
 a80083a <=( A203  and  (not A202) );
 a80084a <=( a80083a  and  a80080a );
 a80085a <=( a80084a  and  a80077a );
 a80088a <=( A266  and  (not A265) );
 a80091a <=( (not A269)  and  A267 );
 a80092a <=( a80091a  and  a80088a );
 a80095a <=( A299  and  (not A298) );
 a80098a <=( (not A302)  and  A300 );
 a80099a <=( a80098a  and  a80095a );
 a80100a <=( a80099a  and  a80092a );
 a80104a <=( A199  and  A166 );
 a80105a <=( A167  and  a80104a );
 a80108a <=( (not A201)  and  (not A200) );
 a80111a <=( A203  and  (not A202) );
 a80112a <=( a80111a  and  a80108a );
 a80113a <=( a80112a  and  a80105a );
 a80116a <=( (not A266)  and  A265 );
 a80119a <=( A268  and  A267 );
 a80120a <=( a80119a  and  a80116a );
 a80123a <=( (not A299)  and  A298 );
 a80126a <=( A301  and  A300 );
 a80127a <=( a80126a  and  a80123a );
 a80128a <=( a80127a  and  a80120a );
 a80132a <=( A199  and  A166 );
 a80133a <=( A167  and  a80132a );
 a80136a <=( (not A201)  and  (not A200) );
 a80139a <=( A203  and  (not A202) );
 a80140a <=( a80139a  and  a80136a );
 a80141a <=( a80140a  and  a80133a );
 a80144a <=( (not A266)  and  A265 );
 a80147a <=( A268  and  A267 );
 a80148a <=( a80147a  and  a80144a );
 a80151a <=( (not A299)  and  A298 );
 a80154a <=( (not A302)  and  A300 );
 a80155a <=( a80154a  and  a80151a );
 a80156a <=( a80155a  and  a80148a );
 a80160a <=( A199  and  A166 );
 a80161a <=( A167  and  a80160a );
 a80164a <=( (not A201)  and  (not A200) );
 a80167a <=( A203  and  (not A202) );
 a80168a <=( a80167a  and  a80164a );
 a80169a <=( a80168a  and  a80161a );
 a80172a <=( (not A266)  and  A265 );
 a80175a <=( A268  and  A267 );
 a80176a <=( a80175a  and  a80172a );
 a80179a <=( A299  and  (not A298) );
 a80182a <=( A301  and  A300 );
 a80183a <=( a80182a  and  a80179a );
 a80184a <=( a80183a  and  a80176a );
 a80188a <=( A199  and  A166 );
 a80189a <=( A167  and  a80188a );
 a80192a <=( (not A201)  and  (not A200) );
 a80195a <=( A203  and  (not A202) );
 a80196a <=( a80195a  and  a80192a );
 a80197a <=( a80196a  and  a80189a );
 a80200a <=( (not A266)  and  A265 );
 a80203a <=( A268  and  A267 );
 a80204a <=( a80203a  and  a80200a );
 a80207a <=( A299  and  (not A298) );
 a80210a <=( (not A302)  and  A300 );
 a80211a <=( a80210a  and  a80207a );
 a80212a <=( a80211a  and  a80204a );
 a80216a <=( A199  and  A166 );
 a80217a <=( A167  and  a80216a );
 a80220a <=( (not A201)  and  (not A200) );
 a80223a <=( A203  and  (not A202) );
 a80224a <=( a80223a  and  a80220a );
 a80225a <=( a80224a  and  a80217a );
 a80228a <=( (not A266)  and  A265 );
 a80231a <=( (not A269)  and  A267 );
 a80232a <=( a80231a  and  a80228a );
 a80235a <=( (not A299)  and  A298 );
 a80238a <=( A301  and  A300 );
 a80239a <=( a80238a  and  a80235a );
 a80240a <=( a80239a  and  a80232a );
 a80244a <=( A199  and  A166 );
 a80245a <=( A167  and  a80244a );
 a80248a <=( (not A201)  and  (not A200) );
 a80251a <=( A203  and  (not A202) );
 a80252a <=( a80251a  and  a80248a );
 a80253a <=( a80252a  and  a80245a );
 a80256a <=( (not A266)  and  A265 );
 a80259a <=( (not A269)  and  A267 );
 a80260a <=( a80259a  and  a80256a );
 a80263a <=( (not A299)  and  A298 );
 a80266a <=( (not A302)  and  A300 );
 a80267a <=( a80266a  and  a80263a );
 a80268a <=( a80267a  and  a80260a );
 a80272a <=( A199  and  A166 );
 a80273a <=( A167  and  a80272a );
 a80276a <=( (not A201)  and  (not A200) );
 a80279a <=( A203  and  (not A202) );
 a80280a <=( a80279a  and  a80276a );
 a80281a <=( a80280a  and  a80273a );
 a80284a <=( (not A266)  and  A265 );
 a80287a <=( (not A269)  and  A267 );
 a80288a <=( a80287a  and  a80284a );
 a80291a <=( A299  and  (not A298) );
 a80294a <=( A301  and  A300 );
 a80295a <=( a80294a  and  a80291a );
 a80296a <=( a80295a  and  a80288a );
 a80300a <=( A199  and  A166 );
 a80301a <=( A167  and  a80300a );
 a80304a <=( (not A201)  and  (not A200) );
 a80307a <=( A203  and  (not A202) );
 a80308a <=( a80307a  and  a80304a );
 a80309a <=( a80308a  and  a80301a );
 a80312a <=( (not A266)  and  A265 );
 a80315a <=( (not A269)  and  A267 );
 a80316a <=( a80315a  and  a80312a );
 a80319a <=( A299  and  (not A298) );
 a80322a <=( (not A302)  and  A300 );
 a80323a <=( a80322a  and  a80319a );
 a80324a <=( a80323a  and  a80316a );
 a80328a <=( (not A199)  and  (not A166) );
 a80329a <=( (not A167)  and  a80328a );
 a80332a <=( A201  and  A200 );
 a80335a <=( (not A265)  and  A202 );
 a80336a <=( a80335a  and  a80332a );
 a80337a <=( a80336a  and  a80329a );
 a80340a <=( A267  and  A266 );
 a80343a <=( A298  and  A268 );
 a80344a <=( a80343a  and  a80340a );
 a80347a <=( (not A300)  and  (not A299) );
 a80350a <=( A302  and  (not A301) );
 a80351a <=( a80350a  and  a80347a );
 a80352a <=( a80351a  and  a80344a );
 a80356a <=( (not A199)  and  (not A166) );
 a80357a <=( (not A167)  and  a80356a );
 a80360a <=( A201  and  A200 );
 a80363a <=( (not A265)  and  A202 );
 a80364a <=( a80363a  and  a80360a );
 a80365a <=( a80364a  and  a80357a );
 a80368a <=( A267  and  A266 );
 a80371a <=( (not A298)  and  A268 );
 a80372a <=( a80371a  and  a80368a );
 a80375a <=( (not A300)  and  A299 );
 a80378a <=( A302  and  (not A301) );
 a80379a <=( a80378a  and  a80375a );
 a80380a <=( a80379a  and  a80372a );
 a80384a <=( (not A199)  and  (not A166) );
 a80385a <=( (not A167)  and  a80384a );
 a80388a <=( A201  and  A200 );
 a80391a <=( (not A265)  and  A202 );
 a80392a <=( a80391a  and  a80388a );
 a80393a <=( a80392a  and  a80385a );
 a80396a <=( A267  and  A266 );
 a80399a <=( A298  and  (not A269) );
 a80400a <=( a80399a  and  a80396a );
 a80403a <=( (not A300)  and  (not A299) );
 a80406a <=( A302  and  (not A301) );
 a80407a <=( a80406a  and  a80403a );
 a80408a <=( a80407a  and  a80400a );
 a80412a <=( (not A199)  and  (not A166) );
 a80413a <=( (not A167)  and  a80412a );
 a80416a <=( A201  and  A200 );
 a80419a <=( (not A265)  and  A202 );
 a80420a <=( a80419a  and  a80416a );
 a80421a <=( a80420a  and  a80413a );
 a80424a <=( A267  and  A266 );
 a80427a <=( (not A298)  and  (not A269) );
 a80428a <=( a80427a  and  a80424a );
 a80431a <=( (not A300)  and  A299 );
 a80434a <=( A302  and  (not A301) );
 a80435a <=( a80434a  and  a80431a );
 a80436a <=( a80435a  and  a80428a );
 a80440a <=( (not A199)  and  (not A166) );
 a80441a <=( (not A167)  and  a80440a );
 a80444a <=( A201  and  A200 );
 a80447a <=( (not A265)  and  A202 );
 a80448a <=( a80447a  and  a80444a );
 a80449a <=( a80448a  and  a80441a );
 a80452a <=( (not A267)  and  A266 );
 a80455a <=( A269  and  (not A268) );
 a80456a <=( a80455a  and  a80452a );
 a80459a <=( (not A299)  and  A298 );
 a80462a <=( A301  and  A300 );
 a80463a <=( a80462a  and  a80459a );
 a80464a <=( a80463a  and  a80456a );
 a80468a <=( (not A199)  and  (not A166) );
 a80469a <=( (not A167)  and  a80468a );
 a80472a <=( A201  and  A200 );
 a80475a <=( (not A265)  and  A202 );
 a80476a <=( a80475a  and  a80472a );
 a80477a <=( a80476a  and  a80469a );
 a80480a <=( (not A267)  and  A266 );
 a80483a <=( A269  and  (not A268) );
 a80484a <=( a80483a  and  a80480a );
 a80487a <=( (not A299)  and  A298 );
 a80490a <=( (not A302)  and  A300 );
 a80491a <=( a80490a  and  a80487a );
 a80492a <=( a80491a  and  a80484a );
 a80496a <=( (not A199)  and  (not A166) );
 a80497a <=( (not A167)  and  a80496a );
 a80500a <=( A201  and  A200 );
 a80503a <=( (not A265)  and  A202 );
 a80504a <=( a80503a  and  a80500a );
 a80505a <=( a80504a  and  a80497a );
 a80508a <=( (not A267)  and  A266 );
 a80511a <=( A269  and  (not A268) );
 a80512a <=( a80511a  and  a80508a );
 a80515a <=( A299  and  (not A298) );
 a80518a <=( A301  and  A300 );
 a80519a <=( a80518a  and  a80515a );
 a80520a <=( a80519a  and  a80512a );
 a80524a <=( (not A199)  and  (not A166) );
 a80525a <=( (not A167)  and  a80524a );
 a80528a <=( A201  and  A200 );
 a80531a <=( (not A265)  and  A202 );
 a80532a <=( a80531a  and  a80528a );
 a80533a <=( a80532a  and  a80525a );
 a80536a <=( (not A267)  and  A266 );
 a80539a <=( A269  and  (not A268) );
 a80540a <=( a80539a  and  a80536a );
 a80543a <=( A299  and  (not A298) );
 a80546a <=( (not A302)  and  A300 );
 a80547a <=( a80546a  and  a80543a );
 a80548a <=( a80547a  and  a80540a );
 a80552a <=( (not A199)  and  (not A166) );
 a80553a <=( (not A167)  and  a80552a );
 a80556a <=( A201  and  A200 );
 a80559a <=( A265  and  A202 );
 a80560a <=( a80559a  and  a80556a );
 a80561a <=( a80560a  and  a80553a );
 a80564a <=( A267  and  (not A266) );
 a80567a <=( A298  and  A268 );
 a80568a <=( a80567a  and  a80564a );
 a80571a <=( (not A300)  and  (not A299) );
 a80574a <=( A302  and  (not A301) );
 a80575a <=( a80574a  and  a80571a );
 a80576a <=( a80575a  and  a80568a );
 a80580a <=( (not A199)  and  (not A166) );
 a80581a <=( (not A167)  and  a80580a );
 a80584a <=( A201  and  A200 );
 a80587a <=( A265  and  A202 );
 a80588a <=( a80587a  and  a80584a );
 a80589a <=( a80588a  and  a80581a );
 a80592a <=( A267  and  (not A266) );
 a80595a <=( (not A298)  and  A268 );
 a80596a <=( a80595a  and  a80592a );
 a80599a <=( (not A300)  and  A299 );
 a80602a <=( A302  and  (not A301) );
 a80603a <=( a80602a  and  a80599a );
 a80604a <=( a80603a  and  a80596a );
 a80608a <=( (not A199)  and  (not A166) );
 a80609a <=( (not A167)  and  a80608a );
 a80612a <=( A201  and  A200 );
 a80615a <=( A265  and  A202 );
 a80616a <=( a80615a  and  a80612a );
 a80617a <=( a80616a  and  a80609a );
 a80620a <=( A267  and  (not A266) );
 a80623a <=( A298  and  (not A269) );
 a80624a <=( a80623a  and  a80620a );
 a80627a <=( (not A300)  and  (not A299) );
 a80630a <=( A302  and  (not A301) );
 a80631a <=( a80630a  and  a80627a );
 a80632a <=( a80631a  and  a80624a );
 a80636a <=( (not A199)  and  (not A166) );
 a80637a <=( (not A167)  and  a80636a );
 a80640a <=( A201  and  A200 );
 a80643a <=( A265  and  A202 );
 a80644a <=( a80643a  and  a80640a );
 a80645a <=( a80644a  and  a80637a );
 a80648a <=( A267  and  (not A266) );
 a80651a <=( (not A298)  and  (not A269) );
 a80652a <=( a80651a  and  a80648a );
 a80655a <=( (not A300)  and  A299 );
 a80658a <=( A302  and  (not A301) );
 a80659a <=( a80658a  and  a80655a );
 a80660a <=( a80659a  and  a80652a );
 a80664a <=( (not A199)  and  (not A166) );
 a80665a <=( (not A167)  and  a80664a );
 a80668a <=( A201  and  A200 );
 a80671a <=( A265  and  A202 );
 a80672a <=( a80671a  and  a80668a );
 a80673a <=( a80672a  and  a80665a );
 a80676a <=( (not A267)  and  (not A266) );
 a80679a <=( A269  and  (not A268) );
 a80680a <=( a80679a  and  a80676a );
 a80683a <=( (not A299)  and  A298 );
 a80686a <=( A301  and  A300 );
 a80687a <=( a80686a  and  a80683a );
 a80688a <=( a80687a  and  a80680a );
 a80692a <=( (not A199)  and  (not A166) );
 a80693a <=( (not A167)  and  a80692a );
 a80696a <=( A201  and  A200 );
 a80699a <=( A265  and  A202 );
 a80700a <=( a80699a  and  a80696a );
 a80701a <=( a80700a  and  a80693a );
 a80704a <=( (not A267)  and  (not A266) );
 a80707a <=( A269  and  (not A268) );
 a80708a <=( a80707a  and  a80704a );
 a80711a <=( (not A299)  and  A298 );
 a80714a <=( (not A302)  and  A300 );
 a80715a <=( a80714a  and  a80711a );
 a80716a <=( a80715a  and  a80708a );
 a80720a <=( (not A199)  and  (not A166) );
 a80721a <=( (not A167)  and  a80720a );
 a80724a <=( A201  and  A200 );
 a80727a <=( A265  and  A202 );
 a80728a <=( a80727a  and  a80724a );
 a80729a <=( a80728a  and  a80721a );
 a80732a <=( (not A267)  and  (not A266) );
 a80735a <=( A269  and  (not A268) );
 a80736a <=( a80735a  and  a80732a );
 a80739a <=( A299  and  (not A298) );
 a80742a <=( A301  and  A300 );
 a80743a <=( a80742a  and  a80739a );
 a80744a <=( a80743a  and  a80736a );
 a80748a <=( (not A199)  and  (not A166) );
 a80749a <=( (not A167)  and  a80748a );
 a80752a <=( A201  and  A200 );
 a80755a <=( A265  and  A202 );
 a80756a <=( a80755a  and  a80752a );
 a80757a <=( a80756a  and  a80749a );
 a80760a <=( (not A267)  and  (not A266) );
 a80763a <=( A269  and  (not A268) );
 a80764a <=( a80763a  and  a80760a );
 a80767a <=( A299  and  (not A298) );
 a80770a <=( (not A302)  and  A300 );
 a80771a <=( a80770a  and  a80767a );
 a80772a <=( a80771a  and  a80764a );
 a80776a <=( (not A199)  and  (not A166) );
 a80777a <=( (not A167)  and  a80776a );
 a80780a <=( A201  and  A200 );
 a80783a <=( (not A265)  and  (not A203) );
 a80784a <=( a80783a  and  a80780a );
 a80785a <=( a80784a  and  a80777a );
 a80788a <=( A267  and  A266 );
 a80791a <=( A298  and  A268 );
 a80792a <=( a80791a  and  a80788a );
 a80795a <=( (not A300)  and  (not A299) );
 a80798a <=( A302  and  (not A301) );
 a80799a <=( a80798a  and  a80795a );
 a80800a <=( a80799a  and  a80792a );
 a80804a <=( (not A199)  and  (not A166) );
 a80805a <=( (not A167)  and  a80804a );
 a80808a <=( A201  and  A200 );
 a80811a <=( (not A265)  and  (not A203) );
 a80812a <=( a80811a  and  a80808a );
 a80813a <=( a80812a  and  a80805a );
 a80816a <=( A267  and  A266 );
 a80819a <=( (not A298)  and  A268 );
 a80820a <=( a80819a  and  a80816a );
 a80823a <=( (not A300)  and  A299 );
 a80826a <=( A302  and  (not A301) );
 a80827a <=( a80826a  and  a80823a );
 a80828a <=( a80827a  and  a80820a );
 a80832a <=( (not A199)  and  (not A166) );
 a80833a <=( (not A167)  and  a80832a );
 a80836a <=( A201  and  A200 );
 a80839a <=( (not A265)  and  (not A203) );
 a80840a <=( a80839a  and  a80836a );
 a80841a <=( a80840a  and  a80833a );
 a80844a <=( A267  and  A266 );
 a80847a <=( A298  and  (not A269) );
 a80848a <=( a80847a  and  a80844a );
 a80851a <=( (not A300)  and  (not A299) );
 a80854a <=( A302  and  (not A301) );
 a80855a <=( a80854a  and  a80851a );
 a80856a <=( a80855a  and  a80848a );
 a80860a <=( (not A199)  and  (not A166) );
 a80861a <=( (not A167)  and  a80860a );
 a80864a <=( A201  and  A200 );
 a80867a <=( (not A265)  and  (not A203) );
 a80868a <=( a80867a  and  a80864a );
 a80869a <=( a80868a  and  a80861a );
 a80872a <=( A267  and  A266 );
 a80875a <=( (not A298)  and  (not A269) );
 a80876a <=( a80875a  and  a80872a );
 a80879a <=( (not A300)  and  A299 );
 a80882a <=( A302  and  (not A301) );
 a80883a <=( a80882a  and  a80879a );
 a80884a <=( a80883a  and  a80876a );
 a80888a <=( (not A199)  and  (not A166) );
 a80889a <=( (not A167)  and  a80888a );
 a80892a <=( A201  and  A200 );
 a80895a <=( (not A265)  and  (not A203) );
 a80896a <=( a80895a  and  a80892a );
 a80897a <=( a80896a  and  a80889a );
 a80900a <=( (not A267)  and  A266 );
 a80903a <=( A269  and  (not A268) );
 a80904a <=( a80903a  and  a80900a );
 a80907a <=( (not A299)  and  A298 );
 a80910a <=( A301  and  A300 );
 a80911a <=( a80910a  and  a80907a );
 a80912a <=( a80911a  and  a80904a );
 a80916a <=( (not A199)  and  (not A166) );
 a80917a <=( (not A167)  and  a80916a );
 a80920a <=( A201  and  A200 );
 a80923a <=( (not A265)  and  (not A203) );
 a80924a <=( a80923a  and  a80920a );
 a80925a <=( a80924a  and  a80917a );
 a80928a <=( (not A267)  and  A266 );
 a80931a <=( A269  and  (not A268) );
 a80932a <=( a80931a  and  a80928a );
 a80935a <=( (not A299)  and  A298 );
 a80938a <=( (not A302)  and  A300 );
 a80939a <=( a80938a  and  a80935a );
 a80940a <=( a80939a  and  a80932a );
 a80944a <=( (not A199)  and  (not A166) );
 a80945a <=( (not A167)  and  a80944a );
 a80948a <=( A201  and  A200 );
 a80951a <=( (not A265)  and  (not A203) );
 a80952a <=( a80951a  and  a80948a );
 a80953a <=( a80952a  and  a80945a );
 a80956a <=( (not A267)  and  A266 );
 a80959a <=( A269  and  (not A268) );
 a80960a <=( a80959a  and  a80956a );
 a80963a <=( A299  and  (not A298) );
 a80966a <=( A301  and  A300 );
 a80967a <=( a80966a  and  a80963a );
 a80968a <=( a80967a  and  a80960a );
 a80972a <=( (not A199)  and  (not A166) );
 a80973a <=( (not A167)  and  a80972a );
 a80976a <=( A201  and  A200 );
 a80979a <=( (not A265)  and  (not A203) );
 a80980a <=( a80979a  and  a80976a );
 a80981a <=( a80980a  and  a80973a );
 a80984a <=( (not A267)  and  A266 );
 a80987a <=( A269  and  (not A268) );
 a80988a <=( a80987a  and  a80984a );
 a80991a <=( A299  and  (not A298) );
 a80994a <=( (not A302)  and  A300 );
 a80995a <=( a80994a  and  a80991a );
 a80996a <=( a80995a  and  a80988a );
 a81000a <=( (not A199)  and  (not A166) );
 a81001a <=( (not A167)  and  a81000a );
 a81004a <=( A201  and  A200 );
 a81007a <=( A265  and  (not A203) );
 a81008a <=( a81007a  and  a81004a );
 a81009a <=( a81008a  and  a81001a );
 a81012a <=( A267  and  (not A266) );
 a81015a <=( A298  and  A268 );
 a81016a <=( a81015a  and  a81012a );
 a81019a <=( (not A300)  and  (not A299) );
 a81022a <=( A302  and  (not A301) );
 a81023a <=( a81022a  and  a81019a );
 a81024a <=( a81023a  and  a81016a );
 a81028a <=( (not A199)  and  (not A166) );
 a81029a <=( (not A167)  and  a81028a );
 a81032a <=( A201  and  A200 );
 a81035a <=( A265  and  (not A203) );
 a81036a <=( a81035a  and  a81032a );
 a81037a <=( a81036a  and  a81029a );
 a81040a <=( A267  and  (not A266) );
 a81043a <=( (not A298)  and  A268 );
 a81044a <=( a81043a  and  a81040a );
 a81047a <=( (not A300)  and  A299 );
 a81050a <=( A302  and  (not A301) );
 a81051a <=( a81050a  and  a81047a );
 a81052a <=( a81051a  and  a81044a );
 a81056a <=( (not A199)  and  (not A166) );
 a81057a <=( (not A167)  and  a81056a );
 a81060a <=( A201  and  A200 );
 a81063a <=( A265  and  (not A203) );
 a81064a <=( a81063a  and  a81060a );
 a81065a <=( a81064a  and  a81057a );
 a81068a <=( A267  and  (not A266) );
 a81071a <=( A298  and  (not A269) );
 a81072a <=( a81071a  and  a81068a );
 a81075a <=( (not A300)  and  (not A299) );
 a81078a <=( A302  and  (not A301) );
 a81079a <=( a81078a  and  a81075a );
 a81080a <=( a81079a  and  a81072a );
 a81084a <=( (not A199)  and  (not A166) );
 a81085a <=( (not A167)  and  a81084a );
 a81088a <=( A201  and  A200 );
 a81091a <=( A265  and  (not A203) );
 a81092a <=( a81091a  and  a81088a );
 a81093a <=( a81092a  and  a81085a );
 a81096a <=( A267  and  (not A266) );
 a81099a <=( (not A298)  and  (not A269) );
 a81100a <=( a81099a  and  a81096a );
 a81103a <=( (not A300)  and  A299 );
 a81106a <=( A302  and  (not A301) );
 a81107a <=( a81106a  and  a81103a );
 a81108a <=( a81107a  and  a81100a );
 a81112a <=( (not A199)  and  (not A166) );
 a81113a <=( (not A167)  and  a81112a );
 a81116a <=( A201  and  A200 );
 a81119a <=( A265  and  (not A203) );
 a81120a <=( a81119a  and  a81116a );
 a81121a <=( a81120a  and  a81113a );
 a81124a <=( (not A267)  and  (not A266) );
 a81127a <=( A269  and  (not A268) );
 a81128a <=( a81127a  and  a81124a );
 a81131a <=( (not A299)  and  A298 );
 a81134a <=( A301  and  A300 );
 a81135a <=( a81134a  and  a81131a );
 a81136a <=( a81135a  and  a81128a );
 a81140a <=( (not A199)  and  (not A166) );
 a81141a <=( (not A167)  and  a81140a );
 a81144a <=( A201  and  A200 );
 a81147a <=( A265  and  (not A203) );
 a81148a <=( a81147a  and  a81144a );
 a81149a <=( a81148a  and  a81141a );
 a81152a <=( (not A267)  and  (not A266) );
 a81155a <=( A269  and  (not A268) );
 a81156a <=( a81155a  and  a81152a );
 a81159a <=( (not A299)  and  A298 );
 a81162a <=( (not A302)  and  A300 );
 a81163a <=( a81162a  and  a81159a );
 a81164a <=( a81163a  and  a81156a );
 a81168a <=( (not A199)  and  (not A166) );
 a81169a <=( (not A167)  and  a81168a );
 a81172a <=( A201  and  A200 );
 a81175a <=( A265  and  (not A203) );
 a81176a <=( a81175a  and  a81172a );
 a81177a <=( a81176a  and  a81169a );
 a81180a <=( (not A267)  and  (not A266) );
 a81183a <=( A269  and  (not A268) );
 a81184a <=( a81183a  and  a81180a );
 a81187a <=( A299  and  (not A298) );
 a81190a <=( A301  and  A300 );
 a81191a <=( a81190a  and  a81187a );
 a81192a <=( a81191a  and  a81184a );
 a81196a <=( (not A199)  and  (not A166) );
 a81197a <=( (not A167)  and  a81196a );
 a81200a <=( A201  and  A200 );
 a81203a <=( A265  and  (not A203) );
 a81204a <=( a81203a  and  a81200a );
 a81205a <=( a81204a  and  a81197a );
 a81208a <=( (not A267)  and  (not A266) );
 a81211a <=( A269  and  (not A268) );
 a81212a <=( a81211a  and  a81208a );
 a81215a <=( A299  and  (not A298) );
 a81218a <=( (not A302)  and  A300 );
 a81219a <=( a81218a  and  a81215a );
 a81220a <=( a81219a  and  a81212a );
 a81224a <=( (not A199)  and  (not A166) );
 a81225a <=( (not A167)  and  a81224a );
 a81228a <=( (not A201)  and  A200 );
 a81231a <=( A203  and  (not A202) );
 a81232a <=( a81231a  and  a81228a );
 a81233a <=( a81232a  and  a81225a );
 a81236a <=( A266  and  (not A265) );
 a81239a <=( A268  and  A267 );
 a81240a <=( a81239a  and  a81236a );
 a81243a <=( (not A299)  and  A298 );
 a81246a <=( A301  and  A300 );
 a81247a <=( a81246a  and  a81243a );
 a81248a <=( a81247a  and  a81240a );
 a81252a <=( (not A199)  and  (not A166) );
 a81253a <=( (not A167)  and  a81252a );
 a81256a <=( (not A201)  and  A200 );
 a81259a <=( A203  and  (not A202) );
 a81260a <=( a81259a  and  a81256a );
 a81261a <=( a81260a  and  a81253a );
 a81264a <=( A266  and  (not A265) );
 a81267a <=( A268  and  A267 );
 a81268a <=( a81267a  and  a81264a );
 a81271a <=( (not A299)  and  A298 );
 a81274a <=( (not A302)  and  A300 );
 a81275a <=( a81274a  and  a81271a );
 a81276a <=( a81275a  and  a81268a );
 a81280a <=( (not A199)  and  (not A166) );
 a81281a <=( (not A167)  and  a81280a );
 a81284a <=( (not A201)  and  A200 );
 a81287a <=( A203  and  (not A202) );
 a81288a <=( a81287a  and  a81284a );
 a81289a <=( a81288a  and  a81281a );
 a81292a <=( A266  and  (not A265) );
 a81295a <=( A268  and  A267 );
 a81296a <=( a81295a  and  a81292a );
 a81299a <=( A299  and  (not A298) );
 a81302a <=( A301  and  A300 );
 a81303a <=( a81302a  and  a81299a );
 a81304a <=( a81303a  and  a81296a );
 a81308a <=( (not A199)  and  (not A166) );
 a81309a <=( (not A167)  and  a81308a );
 a81312a <=( (not A201)  and  A200 );
 a81315a <=( A203  and  (not A202) );
 a81316a <=( a81315a  and  a81312a );
 a81317a <=( a81316a  and  a81309a );
 a81320a <=( A266  and  (not A265) );
 a81323a <=( A268  and  A267 );
 a81324a <=( a81323a  and  a81320a );
 a81327a <=( A299  and  (not A298) );
 a81330a <=( (not A302)  and  A300 );
 a81331a <=( a81330a  and  a81327a );
 a81332a <=( a81331a  and  a81324a );
 a81336a <=( (not A199)  and  (not A166) );
 a81337a <=( (not A167)  and  a81336a );
 a81340a <=( (not A201)  and  A200 );
 a81343a <=( A203  and  (not A202) );
 a81344a <=( a81343a  and  a81340a );
 a81345a <=( a81344a  and  a81337a );
 a81348a <=( A266  and  (not A265) );
 a81351a <=( (not A269)  and  A267 );
 a81352a <=( a81351a  and  a81348a );
 a81355a <=( (not A299)  and  A298 );
 a81358a <=( A301  and  A300 );
 a81359a <=( a81358a  and  a81355a );
 a81360a <=( a81359a  and  a81352a );
 a81364a <=( (not A199)  and  (not A166) );
 a81365a <=( (not A167)  and  a81364a );
 a81368a <=( (not A201)  and  A200 );
 a81371a <=( A203  and  (not A202) );
 a81372a <=( a81371a  and  a81368a );
 a81373a <=( a81372a  and  a81365a );
 a81376a <=( A266  and  (not A265) );
 a81379a <=( (not A269)  and  A267 );
 a81380a <=( a81379a  and  a81376a );
 a81383a <=( (not A299)  and  A298 );
 a81386a <=( (not A302)  and  A300 );
 a81387a <=( a81386a  and  a81383a );
 a81388a <=( a81387a  and  a81380a );
 a81392a <=( (not A199)  and  (not A166) );
 a81393a <=( (not A167)  and  a81392a );
 a81396a <=( (not A201)  and  A200 );
 a81399a <=( A203  and  (not A202) );
 a81400a <=( a81399a  and  a81396a );
 a81401a <=( a81400a  and  a81393a );
 a81404a <=( A266  and  (not A265) );
 a81407a <=( (not A269)  and  A267 );
 a81408a <=( a81407a  and  a81404a );
 a81411a <=( A299  and  (not A298) );
 a81414a <=( A301  and  A300 );
 a81415a <=( a81414a  and  a81411a );
 a81416a <=( a81415a  and  a81408a );
 a81420a <=( (not A199)  and  (not A166) );
 a81421a <=( (not A167)  and  a81420a );
 a81424a <=( (not A201)  and  A200 );
 a81427a <=( A203  and  (not A202) );
 a81428a <=( a81427a  and  a81424a );
 a81429a <=( a81428a  and  a81421a );
 a81432a <=( A266  and  (not A265) );
 a81435a <=( (not A269)  and  A267 );
 a81436a <=( a81435a  and  a81432a );
 a81439a <=( A299  and  (not A298) );
 a81442a <=( (not A302)  and  A300 );
 a81443a <=( a81442a  and  a81439a );
 a81444a <=( a81443a  and  a81436a );
 a81448a <=( (not A199)  and  (not A166) );
 a81449a <=( (not A167)  and  a81448a );
 a81452a <=( (not A201)  and  A200 );
 a81455a <=( A203  and  (not A202) );
 a81456a <=( a81455a  and  a81452a );
 a81457a <=( a81456a  and  a81449a );
 a81460a <=( (not A266)  and  A265 );
 a81463a <=( A268  and  A267 );
 a81464a <=( a81463a  and  a81460a );
 a81467a <=( (not A299)  and  A298 );
 a81470a <=( A301  and  A300 );
 a81471a <=( a81470a  and  a81467a );
 a81472a <=( a81471a  and  a81464a );
 a81476a <=( (not A199)  and  (not A166) );
 a81477a <=( (not A167)  and  a81476a );
 a81480a <=( (not A201)  and  A200 );
 a81483a <=( A203  and  (not A202) );
 a81484a <=( a81483a  and  a81480a );
 a81485a <=( a81484a  and  a81477a );
 a81488a <=( (not A266)  and  A265 );
 a81491a <=( A268  and  A267 );
 a81492a <=( a81491a  and  a81488a );
 a81495a <=( (not A299)  and  A298 );
 a81498a <=( (not A302)  and  A300 );
 a81499a <=( a81498a  and  a81495a );
 a81500a <=( a81499a  and  a81492a );
 a81504a <=( (not A199)  and  (not A166) );
 a81505a <=( (not A167)  and  a81504a );
 a81508a <=( (not A201)  and  A200 );
 a81511a <=( A203  and  (not A202) );
 a81512a <=( a81511a  and  a81508a );
 a81513a <=( a81512a  and  a81505a );
 a81516a <=( (not A266)  and  A265 );
 a81519a <=( A268  and  A267 );
 a81520a <=( a81519a  and  a81516a );
 a81523a <=( A299  and  (not A298) );
 a81526a <=( A301  and  A300 );
 a81527a <=( a81526a  and  a81523a );
 a81528a <=( a81527a  and  a81520a );
 a81532a <=( (not A199)  and  (not A166) );
 a81533a <=( (not A167)  and  a81532a );
 a81536a <=( (not A201)  and  A200 );
 a81539a <=( A203  and  (not A202) );
 a81540a <=( a81539a  and  a81536a );
 a81541a <=( a81540a  and  a81533a );
 a81544a <=( (not A266)  and  A265 );
 a81547a <=( A268  and  A267 );
 a81548a <=( a81547a  and  a81544a );
 a81551a <=( A299  and  (not A298) );
 a81554a <=( (not A302)  and  A300 );
 a81555a <=( a81554a  and  a81551a );
 a81556a <=( a81555a  and  a81548a );
 a81560a <=( (not A199)  and  (not A166) );
 a81561a <=( (not A167)  and  a81560a );
 a81564a <=( (not A201)  and  A200 );
 a81567a <=( A203  and  (not A202) );
 a81568a <=( a81567a  and  a81564a );
 a81569a <=( a81568a  and  a81561a );
 a81572a <=( (not A266)  and  A265 );
 a81575a <=( (not A269)  and  A267 );
 a81576a <=( a81575a  and  a81572a );
 a81579a <=( (not A299)  and  A298 );
 a81582a <=( A301  and  A300 );
 a81583a <=( a81582a  and  a81579a );
 a81584a <=( a81583a  and  a81576a );
 a81588a <=( (not A199)  and  (not A166) );
 a81589a <=( (not A167)  and  a81588a );
 a81592a <=( (not A201)  and  A200 );
 a81595a <=( A203  and  (not A202) );
 a81596a <=( a81595a  and  a81592a );
 a81597a <=( a81596a  and  a81589a );
 a81600a <=( (not A266)  and  A265 );
 a81603a <=( (not A269)  and  A267 );
 a81604a <=( a81603a  and  a81600a );
 a81607a <=( (not A299)  and  A298 );
 a81610a <=( (not A302)  and  A300 );
 a81611a <=( a81610a  and  a81607a );
 a81612a <=( a81611a  and  a81604a );
 a81616a <=( (not A199)  and  (not A166) );
 a81617a <=( (not A167)  and  a81616a );
 a81620a <=( (not A201)  and  A200 );
 a81623a <=( A203  and  (not A202) );
 a81624a <=( a81623a  and  a81620a );
 a81625a <=( a81624a  and  a81617a );
 a81628a <=( (not A266)  and  A265 );
 a81631a <=( (not A269)  and  A267 );
 a81632a <=( a81631a  and  a81628a );
 a81635a <=( A299  and  (not A298) );
 a81638a <=( A301  and  A300 );
 a81639a <=( a81638a  and  a81635a );
 a81640a <=( a81639a  and  a81632a );
 a81644a <=( (not A199)  and  (not A166) );
 a81645a <=( (not A167)  and  a81644a );
 a81648a <=( (not A201)  and  A200 );
 a81651a <=( A203  and  (not A202) );
 a81652a <=( a81651a  and  a81648a );
 a81653a <=( a81652a  and  a81645a );
 a81656a <=( (not A266)  and  A265 );
 a81659a <=( (not A269)  and  A267 );
 a81660a <=( a81659a  and  a81656a );
 a81663a <=( A299  and  (not A298) );
 a81666a <=( (not A302)  and  A300 );
 a81667a <=( a81666a  and  a81663a );
 a81668a <=( a81667a  and  a81660a );
 a81672a <=( A199  and  (not A166) );
 a81673a <=( (not A167)  and  a81672a );
 a81676a <=( A201  and  (not A200) );
 a81679a <=( (not A265)  and  A202 );
 a81680a <=( a81679a  and  a81676a );
 a81681a <=( a81680a  and  a81673a );
 a81684a <=( A267  and  A266 );
 a81687a <=( A298  and  A268 );
 a81688a <=( a81687a  and  a81684a );
 a81691a <=( (not A300)  and  (not A299) );
 a81694a <=( A302  and  (not A301) );
 a81695a <=( a81694a  and  a81691a );
 a81696a <=( a81695a  and  a81688a );
 a81700a <=( A199  and  (not A166) );
 a81701a <=( (not A167)  and  a81700a );
 a81704a <=( A201  and  (not A200) );
 a81707a <=( (not A265)  and  A202 );
 a81708a <=( a81707a  and  a81704a );
 a81709a <=( a81708a  and  a81701a );
 a81712a <=( A267  and  A266 );
 a81715a <=( (not A298)  and  A268 );
 a81716a <=( a81715a  and  a81712a );
 a81719a <=( (not A300)  and  A299 );
 a81722a <=( A302  and  (not A301) );
 a81723a <=( a81722a  and  a81719a );
 a81724a <=( a81723a  and  a81716a );
 a81728a <=( A199  and  (not A166) );
 a81729a <=( (not A167)  and  a81728a );
 a81732a <=( A201  and  (not A200) );
 a81735a <=( (not A265)  and  A202 );
 a81736a <=( a81735a  and  a81732a );
 a81737a <=( a81736a  and  a81729a );
 a81740a <=( A267  and  A266 );
 a81743a <=( A298  and  (not A269) );
 a81744a <=( a81743a  and  a81740a );
 a81747a <=( (not A300)  and  (not A299) );
 a81750a <=( A302  and  (not A301) );
 a81751a <=( a81750a  and  a81747a );
 a81752a <=( a81751a  and  a81744a );
 a81756a <=( A199  and  (not A166) );
 a81757a <=( (not A167)  and  a81756a );
 a81760a <=( A201  and  (not A200) );
 a81763a <=( (not A265)  and  A202 );
 a81764a <=( a81763a  and  a81760a );
 a81765a <=( a81764a  and  a81757a );
 a81768a <=( A267  and  A266 );
 a81771a <=( (not A298)  and  (not A269) );
 a81772a <=( a81771a  and  a81768a );
 a81775a <=( (not A300)  and  A299 );
 a81778a <=( A302  and  (not A301) );
 a81779a <=( a81778a  and  a81775a );
 a81780a <=( a81779a  and  a81772a );
 a81784a <=( A199  and  (not A166) );
 a81785a <=( (not A167)  and  a81784a );
 a81788a <=( A201  and  (not A200) );
 a81791a <=( (not A265)  and  A202 );
 a81792a <=( a81791a  and  a81788a );
 a81793a <=( a81792a  and  a81785a );
 a81796a <=( (not A267)  and  A266 );
 a81799a <=( A269  and  (not A268) );
 a81800a <=( a81799a  and  a81796a );
 a81803a <=( (not A299)  and  A298 );
 a81806a <=( A301  and  A300 );
 a81807a <=( a81806a  and  a81803a );
 a81808a <=( a81807a  and  a81800a );
 a81812a <=( A199  and  (not A166) );
 a81813a <=( (not A167)  and  a81812a );
 a81816a <=( A201  and  (not A200) );
 a81819a <=( (not A265)  and  A202 );
 a81820a <=( a81819a  and  a81816a );
 a81821a <=( a81820a  and  a81813a );
 a81824a <=( (not A267)  and  A266 );
 a81827a <=( A269  and  (not A268) );
 a81828a <=( a81827a  and  a81824a );
 a81831a <=( (not A299)  and  A298 );
 a81834a <=( (not A302)  and  A300 );
 a81835a <=( a81834a  and  a81831a );
 a81836a <=( a81835a  and  a81828a );
 a81840a <=( A199  and  (not A166) );
 a81841a <=( (not A167)  and  a81840a );
 a81844a <=( A201  and  (not A200) );
 a81847a <=( (not A265)  and  A202 );
 a81848a <=( a81847a  and  a81844a );
 a81849a <=( a81848a  and  a81841a );
 a81852a <=( (not A267)  and  A266 );
 a81855a <=( A269  and  (not A268) );
 a81856a <=( a81855a  and  a81852a );
 a81859a <=( A299  and  (not A298) );
 a81862a <=( A301  and  A300 );
 a81863a <=( a81862a  and  a81859a );
 a81864a <=( a81863a  and  a81856a );
 a81868a <=( A199  and  (not A166) );
 a81869a <=( (not A167)  and  a81868a );
 a81872a <=( A201  and  (not A200) );
 a81875a <=( (not A265)  and  A202 );
 a81876a <=( a81875a  and  a81872a );
 a81877a <=( a81876a  and  a81869a );
 a81880a <=( (not A267)  and  A266 );
 a81883a <=( A269  and  (not A268) );
 a81884a <=( a81883a  and  a81880a );
 a81887a <=( A299  and  (not A298) );
 a81890a <=( (not A302)  and  A300 );
 a81891a <=( a81890a  and  a81887a );
 a81892a <=( a81891a  and  a81884a );
 a81896a <=( A199  and  (not A166) );
 a81897a <=( (not A167)  and  a81896a );
 a81900a <=( A201  and  (not A200) );
 a81903a <=( A265  and  A202 );
 a81904a <=( a81903a  and  a81900a );
 a81905a <=( a81904a  and  a81897a );
 a81908a <=( A267  and  (not A266) );
 a81911a <=( A298  and  A268 );
 a81912a <=( a81911a  and  a81908a );
 a81915a <=( (not A300)  and  (not A299) );
 a81918a <=( A302  and  (not A301) );
 a81919a <=( a81918a  and  a81915a );
 a81920a <=( a81919a  and  a81912a );
 a81924a <=( A199  and  (not A166) );
 a81925a <=( (not A167)  and  a81924a );
 a81928a <=( A201  and  (not A200) );
 a81931a <=( A265  and  A202 );
 a81932a <=( a81931a  and  a81928a );
 a81933a <=( a81932a  and  a81925a );
 a81936a <=( A267  and  (not A266) );
 a81939a <=( (not A298)  and  A268 );
 a81940a <=( a81939a  and  a81936a );
 a81943a <=( (not A300)  and  A299 );
 a81946a <=( A302  and  (not A301) );
 a81947a <=( a81946a  and  a81943a );
 a81948a <=( a81947a  and  a81940a );
 a81952a <=( A199  and  (not A166) );
 a81953a <=( (not A167)  and  a81952a );
 a81956a <=( A201  and  (not A200) );
 a81959a <=( A265  and  A202 );
 a81960a <=( a81959a  and  a81956a );
 a81961a <=( a81960a  and  a81953a );
 a81964a <=( A267  and  (not A266) );
 a81967a <=( A298  and  (not A269) );
 a81968a <=( a81967a  and  a81964a );
 a81971a <=( (not A300)  and  (not A299) );
 a81974a <=( A302  and  (not A301) );
 a81975a <=( a81974a  and  a81971a );
 a81976a <=( a81975a  and  a81968a );
 a81980a <=( A199  and  (not A166) );
 a81981a <=( (not A167)  and  a81980a );
 a81984a <=( A201  and  (not A200) );
 a81987a <=( A265  and  A202 );
 a81988a <=( a81987a  and  a81984a );
 a81989a <=( a81988a  and  a81981a );
 a81992a <=( A267  and  (not A266) );
 a81995a <=( (not A298)  and  (not A269) );
 a81996a <=( a81995a  and  a81992a );
 a81999a <=( (not A300)  and  A299 );
 a82002a <=( A302  and  (not A301) );
 a82003a <=( a82002a  and  a81999a );
 a82004a <=( a82003a  and  a81996a );
 a82008a <=( A199  and  (not A166) );
 a82009a <=( (not A167)  and  a82008a );
 a82012a <=( A201  and  (not A200) );
 a82015a <=( A265  and  A202 );
 a82016a <=( a82015a  and  a82012a );
 a82017a <=( a82016a  and  a82009a );
 a82020a <=( (not A267)  and  (not A266) );
 a82023a <=( A269  and  (not A268) );
 a82024a <=( a82023a  and  a82020a );
 a82027a <=( (not A299)  and  A298 );
 a82030a <=( A301  and  A300 );
 a82031a <=( a82030a  and  a82027a );
 a82032a <=( a82031a  and  a82024a );
 a82036a <=( A199  and  (not A166) );
 a82037a <=( (not A167)  and  a82036a );
 a82040a <=( A201  and  (not A200) );
 a82043a <=( A265  and  A202 );
 a82044a <=( a82043a  and  a82040a );
 a82045a <=( a82044a  and  a82037a );
 a82048a <=( (not A267)  and  (not A266) );
 a82051a <=( A269  and  (not A268) );
 a82052a <=( a82051a  and  a82048a );
 a82055a <=( (not A299)  and  A298 );
 a82058a <=( (not A302)  and  A300 );
 a82059a <=( a82058a  and  a82055a );
 a82060a <=( a82059a  and  a82052a );
 a82064a <=( A199  and  (not A166) );
 a82065a <=( (not A167)  and  a82064a );
 a82068a <=( A201  and  (not A200) );
 a82071a <=( A265  and  A202 );
 a82072a <=( a82071a  and  a82068a );
 a82073a <=( a82072a  and  a82065a );
 a82076a <=( (not A267)  and  (not A266) );
 a82079a <=( A269  and  (not A268) );
 a82080a <=( a82079a  and  a82076a );
 a82083a <=( A299  and  (not A298) );
 a82086a <=( A301  and  A300 );
 a82087a <=( a82086a  and  a82083a );
 a82088a <=( a82087a  and  a82080a );
 a82092a <=( A199  and  (not A166) );
 a82093a <=( (not A167)  and  a82092a );
 a82096a <=( A201  and  (not A200) );
 a82099a <=( A265  and  A202 );
 a82100a <=( a82099a  and  a82096a );
 a82101a <=( a82100a  and  a82093a );
 a82104a <=( (not A267)  and  (not A266) );
 a82107a <=( A269  and  (not A268) );
 a82108a <=( a82107a  and  a82104a );
 a82111a <=( A299  and  (not A298) );
 a82114a <=( (not A302)  and  A300 );
 a82115a <=( a82114a  and  a82111a );
 a82116a <=( a82115a  and  a82108a );
 a82120a <=( A199  and  (not A166) );
 a82121a <=( (not A167)  and  a82120a );
 a82124a <=( A201  and  (not A200) );
 a82127a <=( (not A265)  and  (not A203) );
 a82128a <=( a82127a  and  a82124a );
 a82129a <=( a82128a  and  a82121a );
 a82132a <=( A267  and  A266 );
 a82135a <=( A298  and  A268 );
 a82136a <=( a82135a  and  a82132a );
 a82139a <=( (not A300)  and  (not A299) );
 a82142a <=( A302  and  (not A301) );
 a82143a <=( a82142a  and  a82139a );
 a82144a <=( a82143a  and  a82136a );
 a82148a <=( A199  and  (not A166) );
 a82149a <=( (not A167)  and  a82148a );
 a82152a <=( A201  and  (not A200) );
 a82155a <=( (not A265)  and  (not A203) );
 a82156a <=( a82155a  and  a82152a );
 a82157a <=( a82156a  and  a82149a );
 a82160a <=( A267  and  A266 );
 a82163a <=( (not A298)  and  A268 );
 a82164a <=( a82163a  and  a82160a );
 a82167a <=( (not A300)  and  A299 );
 a82170a <=( A302  and  (not A301) );
 a82171a <=( a82170a  and  a82167a );
 a82172a <=( a82171a  and  a82164a );
 a82176a <=( A199  and  (not A166) );
 a82177a <=( (not A167)  and  a82176a );
 a82180a <=( A201  and  (not A200) );
 a82183a <=( (not A265)  and  (not A203) );
 a82184a <=( a82183a  and  a82180a );
 a82185a <=( a82184a  and  a82177a );
 a82188a <=( A267  and  A266 );
 a82191a <=( A298  and  (not A269) );
 a82192a <=( a82191a  and  a82188a );
 a82195a <=( (not A300)  and  (not A299) );
 a82198a <=( A302  and  (not A301) );
 a82199a <=( a82198a  and  a82195a );
 a82200a <=( a82199a  and  a82192a );
 a82204a <=( A199  and  (not A166) );
 a82205a <=( (not A167)  and  a82204a );
 a82208a <=( A201  and  (not A200) );
 a82211a <=( (not A265)  and  (not A203) );
 a82212a <=( a82211a  and  a82208a );
 a82213a <=( a82212a  and  a82205a );
 a82216a <=( A267  and  A266 );
 a82219a <=( (not A298)  and  (not A269) );
 a82220a <=( a82219a  and  a82216a );
 a82223a <=( (not A300)  and  A299 );
 a82226a <=( A302  and  (not A301) );
 a82227a <=( a82226a  and  a82223a );
 a82228a <=( a82227a  and  a82220a );
 a82232a <=( A199  and  (not A166) );
 a82233a <=( (not A167)  and  a82232a );
 a82236a <=( A201  and  (not A200) );
 a82239a <=( (not A265)  and  (not A203) );
 a82240a <=( a82239a  and  a82236a );
 a82241a <=( a82240a  and  a82233a );
 a82244a <=( (not A267)  and  A266 );
 a82247a <=( A269  and  (not A268) );
 a82248a <=( a82247a  and  a82244a );
 a82251a <=( (not A299)  and  A298 );
 a82254a <=( A301  and  A300 );
 a82255a <=( a82254a  and  a82251a );
 a82256a <=( a82255a  and  a82248a );
 a82260a <=( A199  and  (not A166) );
 a82261a <=( (not A167)  and  a82260a );
 a82264a <=( A201  and  (not A200) );
 a82267a <=( (not A265)  and  (not A203) );
 a82268a <=( a82267a  and  a82264a );
 a82269a <=( a82268a  and  a82261a );
 a82272a <=( (not A267)  and  A266 );
 a82275a <=( A269  and  (not A268) );
 a82276a <=( a82275a  and  a82272a );
 a82279a <=( (not A299)  and  A298 );
 a82282a <=( (not A302)  and  A300 );
 a82283a <=( a82282a  and  a82279a );
 a82284a <=( a82283a  and  a82276a );
 a82288a <=( A199  and  (not A166) );
 a82289a <=( (not A167)  and  a82288a );
 a82292a <=( A201  and  (not A200) );
 a82295a <=( (not A265)  and  (not A203) );
 a82296a <=( a82295a  and  a82292a );
 a82297a <=( a82296a  and  a82289a );
 a82300a <=( (not A267)  and  A266 );
 a82303a <=( A269  and  (not A268) );
 a82304a <=( a82303a  and  a82300a );
 a82307a <=( A299  and  (not A298) );
 a82310a <=( A301  and  A300 );
 a82311a <=( a82310a  and  a82307a );
 a82312a <=( a82311a  and  a82304a );
 a82316a <=( A199  and  (not A166) );
 a82317a <=( (not A167)  and  a82316a );
 a82320a <=( A201  and  (not A200) );
 a82323a <=( (not A265)  and  (not A203) );
 a82324a <=( a82323a  and  a82320a );
 a82325a <=( a82324a  and  a82317a );
 a82328a <=( (not A267)  and  A266 );
 a82331a <=( A269  and  (not A268) );
 a82332a <=( a82331a  and  a82328a );
 a82335a <=( A299  and  (not A298) );
 a82338a <=( (not A302)  and  A300 );
 a82339a <=( a82338a  and  a82335a );
 a82340a <=( a82339a  and  a82332a );
 a82344a <=( A199  and  (not A166) );
 a82345a <=( (not A167)  and  a82344a );
 a82348a <=( A201  and  (not A200) );
 a82351a <=( A265  and  (not A203) );
 a82352a <=( a82351a  and  a82348a );
 a82353a <=( a82352a  and  a82345a );
 a82356a <=( A267  and  (not A266) );
 a82359a <=( A298  and  A268 );
 a82360a <=( a82359a  and  a82356a );
 a82363a <=( (not A300)  and  (not A299) );
 a82366a <=( A302  and  (not A301) );
 a82367a <=( a82366a  and  a82363a );
 a82368a <=( a82367a  and  a82360a );
 a82372a <=( A199  and  (not A166) );
 a82373a <=( (not A167)  and  a82372a );
 a82376a <=( A201  and  (not A200) );
 a82379a <=( A265  and  (not A203) );
 a82380a <=( a82379a  and  a82376a );
 a82381a <=( a82380a  and  a82373a );
 a82384a <=( A267  and  (not A266) );
 a82387a <=( (not A298)  and  A268 );
 a82388a <=( a82387a  and  a82384a );
 a82391a <=( (not A300)  and  A299 );
 a82394a <=( A302  and  (not A301) );
 a82395a <=( a82394a  and  a82391a );
 a82396a <=( a82395a  and  a82388a );
 a82400a <=( A199  and  (not A166) );
 a82401a <=( (not A167)  and  a82400a );
 a82404a <=( A201  and  (not A200) );
 a82407a <=( A265  and  (not A203) );
 a82408a <=( a82407a  and  a82404a );
 a82409a <=( a82408a  and  a82401a );
 a82412a <=( A267  and  (not A266) );
 a82415a <=( A298  and  (not A269) );
 a82416a <=( a82415a  and  a82412a );
 a82419a <=( (not A300)  and  (not A299) );
 a82422a <=( A302  and  (not A301) );
 a82423a <=( a82422a  and  a82419a );
 a82424a <=( a82423a  and  a82416a );
 a82428a <=( A199  and  (not A166) );
 a82429a <=( (not A167)  and  a82428a );
 a82432a <=( A201  and  (not A200) );
 a82435a <=( A265  and  (not A203) );
 a82436a <=( a82435a  and  a82432a );
 a82437a <=( a82436a  and  a82429a );
 a82440a <=( A267  and  (not A266) );
 a82443a <=( (not A298)  and  (not A269) );
 a82444a <=( a82443a  and  a82440a );
 a82447a <=( (not A300)  and  A299 );
 a82450a <=( A302  and  (not A301) );
 a82451a <=( a82450a  and  a82447a );
 a82452a <=( a82451a  and  a82444a );
 a82456a <=( A199  and  (not A166) );
 a82457a <=( (not A167)  and  a82456a );
 a82460a <=( A201  and  (not A200) );
 a82463a <=( A265  and  (not A203) );
 a82464a <=( a82463a  and  a82460a );
 a82465a <=( a82464a  and  a82457a );
 a82468a <=( (not A267)  and  (not A266) );
 a82471a <=( A269  and  (not A268) );
 a82472a <=( a82471a  and  a82468a );
 a82475a <=( (not A299)  and  A298 );
 a82478a <=( A301  and  A300 );
 a82479a <=( a82478a  and  a82475a );
 a82480a <=( a82479a  and  a82472a );
 a82484a <=( A199  and  (not A166) );
 a82485a <=( (not A167)  and  a82484a );
 a82488a <=( A201  and  (not A200) );
 a82491a <=( A265  and  (not A203) );
 a82492a <=( a82491a  and  a82488a );
 a82493a <=( a82492a  and  a82485a );
 a82496a <=( (not A267)  and  (not A266) );
 a82499a <=( A269  and  (not A268) );
 a82500a <=( a82499a  and  a82496a );
 a82503a <=( (not A299)  and  A298 );
 a82506a <=( (not A302)  and  A300 );
 a82507a <=( a82506a  and  a82503a );
 a82508a <=( a82507a  and  a82500a );
 a82512a <=( A199  and  (not A166) );
 a82513a <=( (not A167)  and  a82512a );
 a82516a <=( A201  and  (not A200) );
 a82519a <=( A265  and  (not A203) );
 a82520a <=( a82519a  and  a82516a );
 a82521a <=( a82520a  and  a82513a );
 a82524a <=( (not A267)  and  (not A266) );
 a82527a <=( A269  and  (not A268) );
 a82528a <=( a82527a  and  a82524a );
 a82531a <=( A299  and  (not A298) );
 a82534a <=( A301  and  A300 );
 a82535a <=( a82534a  and  a82531a );
 a82536a <=( a82535a  and  a82528a );
 a82540a <=( A199  and  (not A166) );
 a82541a <=( (not A167)  and  a82540a );
 a82544a <=( A201  and  (not A200) );
 a82547a <=( A265  and  (not A203) );
 a82548a <=( a82547a  and  a82544a );
 a82549a <=( a82548a  and  a82541a );
 a82552a <=( (not A267)  and  (not A266) );
 a82555a <=( A269  and  (not A268) );
 a82556a <=( a82555a  and  a82552a );
 a82559a <=( A299  and  (not A298) );
 a82562a <=( (not A302)  and  A300 );
 a82563a <=( a82562a  and  a82559a );
 a82564a <=( a82563a  and  a82556a );
 a82568a <=( A199  and  (not A166) );
 a82569a <=( (not A167)  and  a82568a );
 a82572a <=( (not A201)  and  (not A200) );
 a82575a <=( A203  and  (not A202) );
 a82576a <=( a82575a  and  a82572a );
 a82577a <=( a82576a  and  a82569a );
 a82580a <=( A266  and  (not A265) );
 a82583a <=( A268  and  A267 );
 a82584a <=( a82583a  and  a82580a );
 a82587a <=( (not A299)  and  A298 );
 a82590a <=( A301  and  A300 );
 a82591a <=( a82590a  and  a82587a );
 a82592a <=( a82591a  and  a82584a );
 a82596a <=( A199  and  (not A166) );
 a82597a <=( (not A167)  and  a82596a );
 a82600a <=( (not A201)  and  (not A200) );
 a82603a <=( A203  and  (not A202) );
 a82604a <=( a82603a  and  a82600a );
 a82605a <=( a82604a  and  a82597a );
 a82608a <=( A266  and  (not A265) );
 a82611a <=( A268  and  A267 );
 a82612a <=( a82611a  and  a82608a );
 a82615a <=( (not A299)  and  A298 );
 a82618a <=( (not A302)  and  A300 );
 a82619a <=( a82618a  and  a82615a );
 a82620a <=( a82619a  and  a82612a );
 a82624a <=( A199  and  (not A166) );
 a82625a <=( (not A167)  and  a82624a );
 a82628a <=( (not A201)  and  (not A200) );
 a82631a <=( A203  and  (not A202) );
 a82632a <=( a82631a  and  a82628a );
 a82633a <=( a82632a  and  a82625a );
 a82636a <=( A266  and  (not A265) );
 a82639a <=( A268  and  A267 );
 a82640a <=( a82639a  and  a82636a );
 a82643a <=( A299  and  (not A298) );
 a82646a <=( A301  and  A300 );
 a82647a <=( a82646a  and  a82643a );
 a82648a <=( a82647a  and  a82640a );
 a82652a <=( A199  and  (not A166) );
 a82653a <=( (not A167)  and  a82652a );
 a82656a <=( (not A201)  and  (not A200) );
 a82659a <=( A203  and  (not A202) );
 a82660a <=( a82659a  and  a82656a );
 a82661a <=( a82660a  and  a82653a );
 a82664a <=( A266  and  (not A265) );
 a82667a <=( A268  and  A267 );
 a82668a <=( a82667a  and  a82664a );
 a82671a <=( A299  and  (not A298) );
 a82674a <=( (not A302)  and  A300 );
 a82675a <=( a82674a  and  a82671a );
 a82676a <=( a82675a  and  a82668a );
 a82680a <=( A199  and  (not A166) );
 a82681a <=( (not A167)  and  a82680a );
 a82684a <=( (not A201)  and  (not A200) );
 a82687a <=( A203  and  (not A202) );
 a82688a <=( a82687a  and  a82684a );
 a82689a <=( a82688a  and  a82681a );
 a82692a <=( A266  and  (not A265) );
 a82695a <=( (not A269)  and  A267 );
 a82696a <=( a82695a  and  a82692a );
 a82699a <=( (not A299)  and  A298 );
 a82702a <=( A301  and  A300 );
 a82703a <=( a82702a  and  a82699a );
 a82704a <=( a82703a  and  a82696a );
 a82708a <=( A199  and  (not A166) );
 a82709a <=( (not A167)  and  a82708a );
 a82712a <=( (not A201)  and  (not A200) );
 a82715a <=( A203  and  (not A202) );
 a82716a <=( a82715a  and  a82712a );
 a82717a <=( a82716a  and  a82709a );
 a82720a <=( A266  and  (not A265) );
 a82723a <=( (not A269)  and  A267 );
 a82724a <=( a82723a  and  a82720a );
 a82727a <=( (not A299)  and  A298 );
 a82730a <=( (not A302)  and  A300 );
 a82731a <=( a82730a  and  a82727a );
 a82732a <=( a82731a  and  a82724a );
 a82736a <=( A199  and  (not A166) );
 a82737a <=( (not A167)  and  a82736a );
 a82740a <=( (not A201)  and  (not A200) );
 a82743a <=( A203  and  (not A202) );
 a82744a <=( a82743a  and  a82740a );
 a82745a <=( a82744a  and  a82737a );
 a82748a <=( A266  and  (not A265) );
 a82751a <=( (not A269)  and  A267 );
 a82752a <=( a82751a  and  a82748a );
 a82755a <=( A299  and  (not A298) );
 a82758a <=( A301  and  A300 );
 a82759a <=( a82758a  and  a82755a );
 a82760a <=( a82759a  and  a82752a );
 a82764a <=( A199  and  (not A166) );
 a82765a <=( (not A167)  and  a82764a );
 a82768a <=( (not A201)  and  (not A200) );
 a82771a <=( A203  and  (not A202) );
 a82772a <=( a82771a  and  a82768a );
 a82773a <=( a82772a  and  a82765a );
 a82776a <=( A266  and  (not A265) );
 a82779a <=( (not A269)  and  A267 );
 a82780a <=( a82779a  and  a82776a );
 a82783a <=( A299  and  (not A298) );
 a82786a <=( (not A302)  and  A300 );
 a82787a <=( a82786a  and  a82783a );
 a82788a <=( a82787a  and  a82780a );
 a82792a <=( A199  and  (not A166) );
 a82793a <=( (not A167)  and  a82792a );
 a82796a <=( (not A201)  and  (not A200) );
 a82799a <=( A203  and  (not A202) );
 a82800a <=( a82799a  and  a82796a );
 a82801a <=( a82800a  and  a82793a );
 a82804a <=( (not A266)  and  A265 );
 a82807a <=( A268  and  A267 );
 a82808a <=( a82807a  and  a82804a );
 a82811a <=( (not A299)  and  A298 );
 a82814a <=( A301  and  A300 );
 a82815a <=( a82814a  and  a82811a );
 a82816a <=( a82815a  and  a82808a );
 a82820a <=( A199  and  (not A166) );
 a82821a <=( (not A167)  and  a82820a );
 a82824a <=( (not A201)  and  (not A200) );
 a82827a <=( A203  and  (not A202) );
 a82828a <=( a82827a  and  a82824a );
 a82829a <=( a82828a  and  a82821a );
 a82832a <=( (not A266)  and  A265 );
 a82835a <=( A268  and  A267 );
 a82836a <=( a82835a  and  a82832a );
 a82839a <=( (not A299)  and  A298 );
 a82842a <=( (not A302)  and  A300 );
 a82843a <=( a82842a  and  a82839a );
 a82844a <=( a82843a  and  a82836a );
 a82848a <=( A199  and  (not A166) );
 a82849a <=( (not A167)  and  a82848a );
 a82852a <=( (not A201)  and  (not A200) );
 a82855a <=( A203  and  (not A202) );
 a82856a <=( a82855a  and  a82852a );
 a82857a <=( a82856a  and  a82849a );
 a82860a <=( (not A266)  and  A265 );
 a82863a <=( A268  and  A267 );
 a82864a <=( a82863a  and  a82860a );
 a82867a <=( A299  and  (not A298) );
 a82870a <=( A301  and  A300 );
 a82871a <=( a82870a  and  a82867a );
 a82872a <=( a82871a  and  a82864a );
 a82876a <=( A199  and  (not A166) );
 a82877a <=( (not A167)  and  a82876a );
 a82880a <=( (not A201)  and  (not A200) );
 a82883a <=( A203  and  (not A202) );
 a82884a <=( a82883a  and  a82880a );
 a82885a <=( a82884a  and  a82877a );
 a82888a <=( (not A266)  and  A265 );
 a82891a <=( A268  and  A267 );
 a82892a <=( a82891a  and  a82888a );
 a82895a <=( A299  and  (not A298) );
 a82898a <=( (not A302)  and  A300 );
 a82899a <=( a82898a  and  a82895a );
 a82900a <=( a82899a  and  a82892a );
 a82904a <=( A199  and  (not A166) );
 a82905a <=( (not A167)  and  a82904a );
 a82908a <=( (not A201)  and  (not A200) );
 a82911a <=( A203  and  (not A202) );
 a82912a <=( a82911a  and  a82908a );
 a82913a <=( a82912a  and  a82905a );
 a82916a <=( (not A266)  and  A265 );
 a82919a <=( (not A269)  and  A267 );
 a82920a <=( a82919a  and  a82916a );
 a82923a <=( (not A299)  and  A298 );
 a82926a <=( A301  and  A300 );
 a82927a <=( a82926a  and  a82923a );
 a82928a <=( a82927a  and  a82920a );
 a82932a <=( A199  and  (not A166) );
 a82933a <=( (not A167)  and  a82932a );
 a82936a <=( (not A201)  and  (not A200) );
 a82939a <=( A203  and  (not A202) );
 a82940a <=( a82939a  and  a82936a );
 a82941a <=( a82940a  and  a82933a );
 a82944a <=( (not A266)  and  A265 );
 a82947a <=( (not A269)  and  A267 );
 a82948a <=( a82947a  and  a82944a );
 a82951a <=( (not A299)  and  A298 );
 a82954a <=( (not A302)  and  A300 );
 a82955a <=( a82954a  and  a82951a );
 a82956a <=( a82955a  and  a82948a );
 a82960a <=( A199  and  (not A166) );
 a82961a <=( (not A167)  and  a82960a );
 a82964a <=( (not A201)  and  (not A200) );
 a82967a <=( A203  and  (not A202) );
 a82968a <=( a82967a  and  a82964a );
 a82969a <=( a82968a  and  a82961a );
 a82972a <=( (not A266)  and  A265 );
 a82975a <=( (not A269)  and  A267 );
 a82976a <=( a82975a  and  a82972a );
 a82979a <=( A299  and  (not A298) );
 a82982a <=( A301  and  A300 );
 a82983a <=( a82982a  and  a82979a );
 a82984a <=( a82983a  and  a82976a );
 a82988a <=( A199  and  (not A166) );
 a82989a <=( (not A167)  and  a82988a );
 a82992a <=( (not A201)  and  (not A200) );
 a82995a <=( A203  and  (not A202) );
 a82996a <=( a82995a  and  a82992a );
 a82997a <=( a82996a  and  a82989a );
 a83000a <=( (not A266)  and  A265 );
 a83003a <=( (not A269)  and  A267 );
 a83004a <=( a83003a  and  a83000a );
 a83007a <=( A299  and  (not A298) );
 a83010a <=( (not A302)  and  A300 );
 a83011a <=( a83010a  and  a83007a );
 a83012a <=( a83011a  and  a83004a );
 a83016a <=( A167  and  A168 );
 a83017a <=( A170  and  a83016a );
 a83020a <=( A201  and  (not A166) );
 a83023a <=( A203  and  (not A202) );
 a83024a <=( a83023a  and  a83020a );
 a83025a <=( a83024a  and  a83017a );
 a83028a <=( (not A268)  and  A267 );
 a83031a <=( A298  and  A269 );
 a83032a <=( a83031a  and  a83028a );
 a83035a <=( (not A300)  and  (not A299) );
 a83038a <=( A302  and  (not A301) );
 a83039a <=( a83038a  and  a83035a );
 a83040a <=( a83039a  and  a83032a );
 a83044a <=( A167  and  A168 );
 a83045a <=( A170  and  a83044a );
 a83048a <=( A201  and  (not A166) );
 a83051a <=( A203  and  (not A202) );
 a83052a <=( a83051a  and  a83048a );
 a83053a <=( a83052a  and  a83045a );
 a83056a <=( (not A268)  and  A267 );
 a83059a <=( (not A298)  and  A269 );
 a83060a <=( a83059a  and  a83056a );
 a83063a <=( (not A300)  and  A299 );
 a83066a <=( A302  and  (not A301) );
 a83067a <=( a83066a  and  a83063a );
 a83068a <=( a83067a  and  a83060a );
 a83072a <=( A167  and  A168 );
 a83073a <=( A170  and  a83072a );
 a83076a <=( A201  and  (not A166) );
 a83079a <=( A203  and  (not A202) );
 a83080a <=( a83079a  and  a83076a );
 a83081a <=( a83080a  and  a83073a );
 a83084a <=( A266  and  (not A265) );
 a83087a <=( (not A268)  and  (not A267) );
 a83088a <=( a83087a  and  a83084a );
 a83091a <=( A300  and  A269 );
 a83094a <=( A302  and  (not A301) );
 a83095a <=( a83094a  and  a83091a );
 a83096a <=( a83095a  and  a83088a );
 a83100a <=( A167  and  A168 );
 a83101a <=( A170  and  a83100a );
 a83104a <=( A201  and  (not A166) );
 a83107a <=( A203  and  (not A202) );
 a83108a <=( a83107a  and  a83104a );
 a83109a <=( a83108a  and  a83101a );
 a83112a <=( (not A266)  and  A265 );
 a83115a <=( (not A268)  and  (not A267) );
 a83116a <=( a83115a  and  a83112a );
 a83119a <=( A300  and  A269 );
 a83122a <=( A302  and  (not A301) );
 a83123a <=( a83122a  and  a83119a );
 a83124a <=( a83123a  and  a83116a );
 a83128a <=( (not A167)  and  A168 );
 a83129a <=( A170  and  a83128a );
 a83132a <=( A201  and  A166 );
 a83135a <=( A203  and  (not A202) );
 a83136a <=( a83135a  and  a83132a );
 a83137a <=( a83136a  and  a83129a );
 a83140a <=( (not A268)  and  A267 );
 a83143a <=( A298  and  A269 );
 a83144a <=( a83143a  and  a83140a );
 a83147a <=( (not A300)  and  (not A299) );
 a83150a <=( A302  and  (not A301) );
 a83151a <=( a83150a  and  a83147a );
 a83152a <=( a83151a  and  a83144a );
 a83156a <=( (not A167)  and  A168 );
 a83157a <=( A170  and  a83156a );
 a83160a <=( A201  and  A166 );
 a83163a <=( A203  and  (not A202) );
 a83164a <=( a83163a  and  a83160a );
 a83165a <=( a83164a  and  a83157a );
 a83168a <=( (not A268)  and  A267 );
 a83171a <=( (not A298)  and  A269 );
 a83172a <=( a83171a  and  a83168a );
 a83175a <=( (not A300)  and  A299 );
 a83178a <=( A302  and  (not A301) );
 a83179a <=( a83178a  and  a83175a );
 a83180a <=( a83179a  and  a83172a );
 a83184a <=( (not A167)  and  A168 );
 a83185a <=( A170  and  a83184a );
 a83188a <=( A201  and  A166 );
 a83191a <=( A203  and  (not A202) );
 a83192a <=( a83191a  and  a83188a );
 a83193a <=( a83192a  and  a83185a );
 a83196a <=( A266  and  (not A265) );
 a83199a <=( (not A268)  and  (not A267) );
 a83200a <=( a83199a  and  a83196a );
 a83203a <=( A300  and  A269 );
 a83206a <=( A302  and  (not A301) );
 a83207a <=( a83206a  and  a83203a );
 a83208a <=( a83207a  and  a83200a );
 a83212a <=( (not A167)  and  A168 );
 a83213a <=( A170  and  a83212a );
 a83216a <=( A201  and  A166 );
 a83219a <=( A203  and  (not A202) );
 a83220a <=( a83219a  and  a83216a );
 a83221a <=( a83220a  and  a83213a );
 a83224a <=( (not A266)  and  A265 );
 a83227a <=( (not A268)  and  (not A267) );
 a83228a <=( a83227a  and  a83224a );
 a83231a <=( A300  and  A269 );
 a83234a <=( A302  and  (not A301) );
 a83235a <=( a83234a  and  a83231a );
 a83236a <=( a83235a  and  a83228a );
 a83240a <=( (not A199)  and  (not A168) );
 a83241a <=( A170  and  a83240a );
 a83244a <=( A201  and  A200 );
 a83247a <=( (not A265)  and  A202 );
 a83248a <=( a83247a  and  a83244a );
 a83249a <=( a83248a  and  a83241a );
 a83252a <=( A267  and  A266 );
 a83255a <=( A298  and  A268 );
 a83256a <=( a83255a  and  a83252a );
 a83259a <=( (not A300)  and  (not A299) );
 a83262a <=( A302  and  (not A301) );
 a83263a <=( a83262a  and  a83259a );
 a83264a <=( a83263a  and  a83256a );
 a83268a <=( (not A199)  and  (not A168) );
 a83269a <=( A170  and  a83268a );
 a83272a <=( A201  and  A200 );
 a83275a <=( (not A265)  and  A202 );
 a83276a <=( a83275a  and  a83272a );
 a83277a <=( a83276a  and  a83269a );
 a83280a <=( A267  and  A266 );
 a83283a <=( (not A298)  and  A268 );
 a83284a <=( a83283a  and  a83280a );
 a83287a <=( (not A300)  and  A299 );
 a83290a <=( A302  and  (not A301) );
 a83291a <=( a83290a  and  a83287a );
 a83292a <=( a83291a  and  a83284a );
 a83296a <=( (not A199)  and  (not A168) );
 a83297a <=( A170  and  a83296a );
 a83300a <=( A201  and  A200 );
 a83303a <=( (not A265)  and  A202 );
 a83304a <=( a83303a  and  a83300a );
 a83305a <=( a83304a  and  a83297a );
 a83308a <=( A267  and  A266 );
 a83311a <=( A298  and  (not A269) );
 a83312a <=( a83311a  and  a83308a );
 a83315a <=( (not A300)  and  (not A299) );
 a83318a <=( A302  and  (not A301) );
 a83319a <=( a83318a  and  a83315a );
 a83320a <=( a83319a  and  a83312a );
 a83324a <=( (not A199)  and  (not A168) );
 a83325a <=( A170  and  a83324a );
 a83328a <=( A201  and  A200 );
 a83331a <=( (not A265)  and  A202 );
 a83332a <=( a83331a  and  a83328a );
 a83333a <=( a83332a  and  a83325a );
 a83336a <=( A267  and  A266 );
 a83339a <=( (not A298)  and  (not A269) );
 a83340a <=( a83339a  and  a83336a );
 a83343a <=( (not A300)  and  A299 );
 a83346a <=( A302  and  (not A301) );
 a83347a <=( a83346a  and  a83343a );
 a83348a <=( a83347a  and  a83340a );
 a83352a <=( (not A199)  and  (not A168) );
 a83353a <=( A170  and  a83352a );
 a83356a <=( A201  and  A200 );
 a83359a <=( (not A265)  and  A202 );
 a83360a <=( a83359a  and  a83356a );
 a83361a <=( a83360a  and  a83353a );
 a83364a <=( (not A267)  and  A266 );
 a83367a <=( A269  and  (not A268) );
 a83368a <=( a83367a  and  a83364a );
 a83371a <=( (not A299)  and  A298 );
 a83374a <=( A301  and  A300 );
 a83375a <=( a83374a  and  a83371a );
 a83376a <=( a83375a  and  a83368a );
 a83380a <=( (not A199)  and  (not A168) );
 a83381a <=( A170  and  a83380a );
 a83384a <=( A201  and  A200 );
 a83387a <=( (not A265)  and  A202 );
 a83388a <=( a83387a  and  a83384a );
 a83389a <=( a83388a  and  a83381a );
 a83392a <=( (not A267)  and  A266 );
 a83395a <=( A269  and  (not A268) );
 a83396a <=( a83395a  and  a83392a );
 a83399a <=( (not A299)  and  A298 );
 a83402a <=( (not A302)  and  A300 );
 a83403a <=( a83402a  and  a83399a );
 a83404a <=( a83403a  and  a83396a );
 a83408a <=( (not A199)  and  (not A168) );
 a83409a <=( A170  and  a83408a );
 a83412a <=( A201  and  A200 );
 a83415a <=( (not A265)  and  A202 );
 a83416a <=( a83415a  and  a83412a );
 a83417a <=( a83416a  and  a83409a );
 a83420a <=( (not A267)  and  A266 );
 a83423a <=( A269  and  (not A268) );
 a83424a <=( a83423a  and  a83420a );
 a83427a <=( A299  and  (not A298) );
 a83430a <=( A301  and  A300 );
 a83431a <=( a83430a  and  a83427a );
 a83432a <=( a83431a  and  a83424a );
 a83436a <=( (not A199)  and  (not A168) );
 a83437a <=( A170  and  a83436a );
 a83440a <=( A201  and  A200 );
 a83443a <=( (not A265)  and  A202 );
 a83444a <=( a83443a  and  a83440a );
 a83445a <=( a83444a  and  a83437a );
 a83448a <=( (not A267)  and  A266 );
 a83451a <=( A269  and  (not A268) );
 a83452a <=( a83451a  and  a83448a );
 a83455a <=( A299  and  (not A298) );
 a83458a <=( (not A302)  and  A300 );
 a83459a <=( a83458a  and  a83455a );
 a83460a <=( a83459a  and  a83452a );
 a83464a <=( (not A199)  and  (not A168) );
 a83465a <=( A170  and  a83464a );
 a83468a <=( A201  and  A200 );
 a83471a <=( A265  and  A202 );
 a83472a <=( a83471a  and  a83468a );
 a83473a <=( a83472a  and  a83465a );
 a83476a <=( A267  and  (not A266) );
 a83479a <=( A298  and  A268 );
 a83480a <=( a83479a  and  a83476a );
 a83483a <=( (not A300)  and  (not A299) );
 a83486a <=( A302  and  (not A301) );
 a83487a <=( a83486a  and  a83483a );
 a83488a <=( a83487a  and  a83480a );
 a83492a <=( (not A199)  and  (not A168) );
 a83493a <=( A170  and  a83492a );
 a83496a <=( A201  and  A200 );
 a83499a <=( A265  and  A202 );
 a83500a <=( a83499a  and  a83496a );
 a83501a <=( a83500a  and  a83493a );
 a83504a <=( A267  and  (not A266) );
 a83507a <=( (not A298)  and  A268 );
 a83508a <=( a83507a  and  a83504a );
 a83511a <=( (not A300)  and  A299 );
 a83514a <=( A302  and  (not A301) );
 a83515a <=( a83514a  and  a83511a );
 a83516a <=( a83515a  and  a83508a );
 a83520a <=( (not A199)  and  (not A168) );
 a83521a <=( A170  and  a83520a );
 a83524a <=( A201  and  A200 );
 a83527a <=( A265  and  A202 );
 a83528a <=( a83527a  and  a83524a );
 a83529a <=( a83528a  and  a83521a );
 a83532a <=( A267  and  (not A266) );
 a83535a <=( A298  and  (not A269) );
 a83536a <=( a83535a  and  a83532a );
 a83539a <=( (not A300)  and  (not A299) );
 a83542a <=( A302  and  (not A301) );
 a83543a <=( a83542a  and  a83539a );
 a83544a <=( a83543a  and  a83536a );
 a83548a <=( (not A199)  and  (not A168) );
 a83549a <=( A170  and  a83548a );
 a83552a <=( A201  and  A200 );
 a83555a <=( A265  and  A202 );
 a83556a <=( a83555a  and  a83552a );
 a83557a <=( a83556a  and  a83549a );
 a83560a <=( A267  and  (not A266) );
 a83563a <=( (not A298)  and  (not A269) );
 a83564a <=( a83563a  and  a83560a );
 a83567a <=( (not A300)  and  A299 );
 a83570a <=( A302  and  (not A301) );
 a83571a <=( a83570a  and  a83567a );
 a83572a <=( a83571a  and  a83564a );
 a83576a <=( (not A199)  and  (not A168) );
 a83577a <=( A170  and  a83576a );
 a83580a <=( A201  and  A200 );
 a83583a <=( A265  and  A202 );
 a83584a <=( a83583a  and  a83580a );
 a83585a <=( a83584a  and  a83577a );
 a83588a <=( (not A267)  and  (not A266) );
 a83591a <=( A269  and  (not A268) );
 a83592a <=( a83591a  and  a83588a );
 a83595a <=( (not A299)  and  A298 );
 a83598a <=( A301  and  A300 );
 a83599a <=( a83598a  and  a83595a );
 a83600a <=( a83599a  and  a83592a );
 a83604a <=( (not A199)  and  (not A168) );
 a83605a <=( A170  and  a83604a );
 a83608a <=( A201  and  A200 );
 a83611a <=( A265  and  A202 );
 a83612a <=( a83611a  and  a83608a );
 a83613a <=( a83612a  and  a83605a );
 a83616a <=( (not A267)  and  (not A266) );
 a83619a <=( A269  and  (not A268) );
 a83620a <=( a83619a  and  a83616a );
 a83623a <=( (not A299)  and  A298 );
 a83626a <=( (not A302)  and  A300 );
 a83627a <=( a83626a  and  a83623a );
 a83628a <=( a83627a  and  a83620a );
 a83632a <=( (not A199)  and  (not A168) );
 a83633a <=( A170  and  a83632a );
 a83636a <=( A201  and  A200 );
 a83639a <=( A265  and  A202 );
 a83640a <=( a83639a  and  a83636a );
 a83641a <=( a83640a  and  a83633a );
 a83644a <=( (not A267)  and  (not A266) );
 a83647a <=( A269  and  (not A268) );
 a83648a <=( a83647a  and  a83644a );
 a83651a <=( A299  and  (not A298) );
 a83654a <=( A301  and  A300 );
 a83655a <=( a83654a  and  a83651a );
 a83656a <=( a83655a  and  a83648a );
 a83660a <=( (not A199)  and  (not A168) );
 a83661a <=( A170  and  a83660a );
 a83664a <=( A201  and  A200 );
 a83667a <=( A265  and  A202 );
 a83668a <=( a83667a  and  a83664a );
 a83669a <=( a83668a  and  a83661a );
 a83672a <=( (not A267)  and  (not A266) );
 a83675a <=( A269  and  (not A268) );
 a83676a <=( a83675a  and  a83672a );
 a83679a <=( A299  and  (not A298) );
 a83682a <=( (not A302)  and  A300 );
 a83683a <=( a83682a  and  a83679a );
 a83684a <=( a83683a  and  a83676a );
 a83688a <=( (not A199)  and  (not A168) );
 a83689a <=( A170  and  a83688a );
 a83692a <=( A201  and  A200 );
 a83695a <=( (not A265)  and  (not A203) );
 a83696a <=( a83695a  and  a83692a );
 a83697a <=( a83696a  and  a83689a );
 a83700a <=( A267  and  A266 );
 a83703a <=( A298  and  A268 );
 a83704a <=( a83703a  and  a83700a );
 a83707a <=( (not A300)  and  (not A299) );
 a83710a <=( A302  and  (not A301) );
 a83711a <=( a83710a  and  a83707a );
 a83712a <=( a83711a  and  a83704a );
 a83716a <=( (not A199)  and  (not A168) );
 a83717a <=( A170  and  a83716a );
 a83720a <=( A201  and  A200 );
 a83723a <=( (not A265)  and  (not A203) );
 a83724a <=( a83723a  and  a83720a );
 a83725a <=( a83724a  and  a83717a );
 a83728a <=( A267  and  A266 );
 a83731a <=( (not A298)  and  A268 );
 a83732a <=( a83731a  and  a83728a );
 a83735a <=( (not A300)  and  A299 );
 a83738a <=( A302  and  (not A301) );
 a83739a <=( a83738a  and  a83735a );
 a83740a <=( a83739a  and  a83732a );
 a83744a <=( (not A199)  and  (not A168) );
 a83745a <=( A170  and  a83744a );
 a83748a <=( A201  and  A200 );
 a83751a <=( (not A265)  and  (not A203) );
 a83752a <=( a83751a  and  a83748a );
 a83753a <=( a83752a  and  a83745a );
 a83756a <=( A267  and  A266 );
 a83759a <=( A298  and  (not A269) );
 a83760a <=( a83759a  and  a83756a );
 a83763a <=( (not A300)  and  (not A299) );
 a83766a <=( A302  and  (not A301) );
 a83767a <=( a83766a  and  a83763a );
 a83768a <=( a83767a  and  a83760a );
 a83772a <=( (not A199)  and  (not A168) );
 a83773a <=( A170  and  a83772a );
 a83776a <=( A201  and  A200 );
 a83779a <=( (not A265)  and  (not A203) );
 a83780a <=( a83779a  and  a83776a );
 a83781a <=( a83780a  and  a83773a );
 a83784a <=( A267  and  A266 );
 a83787a <=( (not A298)  and  (not A269) );
 a83788a <=( a83787a  and  a83784a );
 a83791a <=( (not A300)  and  A299 );
 a83794a <=( A302  and  (not A301) );
 a83795a <=( a83794a  and  a83791a );
 a83796a <=( a83795a  and  a83788a );
 a83800a <=( (not A199)  and  (not A168) );
 a83801a <=( A170  and  a83800a );
 a83804a <=( A201  and  A200 );
 a83807a <=( (not A265)  and  (not A203) );
 a83808a <=( a83807a  and  a83804a );
 a83809a <=( a83808a  and  a83801a );
 a83812a <=( (not A267)  and  A266 );
 a83815a <=( A269  and  (not A268) );
 a83816a <=( a83815a  and  a83812a );
 a83819a <=( (not A299)  and  A298 );
 a83822a <=( A301  and  A300 );
 a83823a <=( a83822a  and  a83819a );
 a83824a <=( a83823a  and  a83816a );
 a83828a <=( (not A199)  and  (not A168) );
 a83829a <=( A170  and  a83828a );
 a83832a <=( A201  and  A200 );
 a83835a <=( (not A265)  and  (not A203) );
 a83836a <=( a83835a  and  a83832a );
 a83837a <=( a83836a  and  a83829a );
 a83840a <=( (not A267)  and  A266 );
 a83843a <=( A269  and  (not A268) );
 a83844a <=( a83843a  and  a83840a );
 a83847a <=( (not A299)  and  A298 );
 a83850a <=( (not A302)  and  A300 );
 a83851a <=( a83850a  and  a83847a );
 a83852a <=( a83851a  and  a83844a );
 a83856a <=( (not A199)  and  (not A168) );
 a83857a <=( A170  and  a83856a );
 a83860a <=( A201  and  A200 );
 a83863a <=( (not A265)  and  (not A203) );
 a83864a <=( a83863a  and  a83860a );
 a83865a <=( a83864a  and  a83857a );
 a83868a <=( (not A267)  and  A266 );
 a83871a <=( A269  and  (not A268) );
 a83872a <=( a83871a  and  a83868a );
 a83875a <=( A299  and  (not A298) );
 a83878a <=( A301  and  A300 );
 a83879a <=( a83878a  and  a83875a );
 a83880a <=( a83879a  and  a83872a );
 a83884a <=( (not A199)  and  (not A168) );
 a83885a <=( A170  and  a83884a );
 a83888a <=( A201  and  A200 );
 a83891a <=( (not A265)  and  (not A203) );
 a83892a <=( a83891a  and  a83888a );
 a83893a <=( a83892a  and  a83885a );
 a83896a <=( (not A267)  and  A266 );
 a83899a <=( A269  and  (not A268) );
 a83900a <=( a83899a  and  a83896a );
 a83903a <=( A299  and  (not A298) );
 a83906a <=( (not A302)  and  A300 );
 a83907a <=( a83906a  and  a83903a );
 a83908a <=( a83907a  and  a83900a );
 a83912a <=( (not A199)  and  (not A168) );
 a83913a <=( A170  and  a83912a );
 a83916a <=( A201  and  A200 );
 a83919a <=( A265  and  (not A203) );
 a83920a <=( a83919a  and  a83916a );
 a83921a <=( a83920a  and  a83913a );
 a83924a <=( A267  and  (not A266) );
 a83927a <=( A298  and  A268 );
 a83928a <=( a83927a  and  a83924a );
 a83931a <=( (not A300)  and  (not A299) );
 a83934a <=( A302  and  (not A301) );
 a83935a <=( a83934a  and  a83931a );
 a83936a <=( a83935a  and  a83928a );
 a83940a <=( (not A199)  and  (not A168) );
 a83941a <=( A170  and  a83940a );
 a83944a <=( A201  and  A200 );
 a83947a <=( A265  and  (not A203) );
 a83948a <=( a83947a  and  a83944a );
 a83949a <=( a83948a  and  a83941a );
 a83952a <=( A267  and  (not A266) );
 a83955a <=( (not A298)  and  A268 );
 a83956a <=( a83955a  and  a83952a );
 a83959a <=( (not A300)  and  A299 );
 a83962a <=( A302  and  (not A301) );
 a83963a <=( a83962a  and  a83959a );
 a83964a <=( a83963a  and  a83956a );
 a83968a <=( (not A199)  and  (not A168) );
 a83969a <=( A170  and  a83968a );
 a83972a <=( A201  and  A200 );
 a83975a <=( A265  and  (not A203) );
 a83976a <=( a83975a  and  a83972a );
 a83977a <=( a83976a  and  a83969a );
 a83980a <=( A267  and  (not A266) );
 a83983a <=( A298  and  (not A269) );
 a83984a <=( a83983a  and  a83980a );
 a83987a <=( (not A300)  and  (not A299) );
 a83990a <=( A302  and  (not A301) );
 a83991a <=( a83990a  and  a83987a );
 a83992a <=( a83991a  and  a83984a );
 a83996a <=( (not A199)  and  (not A168) );
 a83997a <=( A170  and  a83996a );
 a84000a <=( A201  and  A200 );
 a84003a <=( A265  and  (not A203) );
 a84004a <=( a84003a  and  a84000a );
 a84005a <=( a84004a  and  a83997a );
 a84008a <=( A267  and  (not A266) );
 a84011a <=( (not A298)  and  (not A269) );
 a84012a <=( a84011a  and  a84008a );
 a84015a <=( (not A300)  and  A299 );
 a84018a <=( A302  and  (not A301) );
 a84019a <=( a84018a  and  a84015a );
 a84020a <=( a84019a  and  a84012a );
 a84024a <=( (not A199)  and  (not A168) );
 a84025a <=( A170  and  a84024a );
 a84028a <=( A201  and  A200 );
 a84031a <=( A265  and  (not A203) );
 a84032a <=( a84031a  and  a84028a );
 a84033a <=( a84032a  and  a84025a );
 a84036a <=( (not A267)  and  (not A266) );
 a84039a <=( A269  and  (not A268) );
 a84040a <=( a84039a  and  a84036a );
 a84043a <=( (not A299)  and  A298 );
 a84046a <=( A301  and  A300 );
 a84047a <=( a84046a  and  a84043a );
 a84048a <=( a84047a  and  a84040a );
 a84052a <=( (not A199)  and  (not A168) );
 a84053a <=( A170  and  a84052a );
 a84056a <=( A201  and  A200 );
 a84059a <=( A265  and  (not A203) );
 a84060a <=( a84059a  and  a84056a );
 a84061a <=( a84060a  and  a84053a );
 a84064a <=( (not A267)  and  (not A266) );
 a84067a <=( A269  and  (not A268) );
 a84068a <=( a84067a  and  a84064a );
 a84071a <=( (not A299)  and  A298 );
 a84074a <=( (not A302)  and  A300 );
 a84075a <=( a84074a  and  a84071a );
 a84076a <=( a84075a  and  a84068a );
 a84080a <=( (not A199)  and  (not A168) );
 a84081a <=( A170  and  a84080a );
 a84084a <=( A201  and  A200 );
 a84087a <=( A265  and  (not A203) );
 a84088a <=( a84087a  and  a84084a );
 a84089a <=( a84088a  and  a84081a );
 a84092a <=( (not A267)  and  (not A266) );
 a84095a <=( A269  and  (not A268) );
 a84096a <=( a84095a  and  a84092a );
 a84099a <=( A299  and  (not A298) );
 a84102a <=( A301  and  A300 );
 a84103a <=( a84102a  and  a84099a );
 a84104a <=( a84103a  and  a84096a );
 a84108a <=( (not A199)  and  (not A168) );
 a84109a <=( A170  and  a84108a );
 a84112a <=( A201  and  A200 );
 a84115a <=( A265  and  (not A203) );
 a84116a <=( a84115a  and  a84112a );
 a84117a <=( a84116a  and  a84109a );
 a84120a <=( (not A267)  and  (not A266) );
 a84123a <=( A269  and  (not A268) );
 a84124a <=( a84123a  and  a84120a );
 a84127a <=( A299  and  (not A298) );
 a84130a <=( (not A302)  and  A300 );
 a84131a <=( a84130a  and  a84127a );
 a84132a <=( a84131a  and  a84124a );
 a84136a <=( (not A199)  and  (not A168) );
 a84137a <=( A170  and  a84136a );
 a84140a <=( (not A201)  and  A200 );
 a84143a <=( A203  and  (not A202) );
 a84144a <=( a84143a  and  a84140a );
 a84145a <=( a84144a  and  a84137a );
 a84148a <=( A266  and  (not A265) );
 a84151a <=( A268  and  A267 );
 a84152a <=( a84151a  and  a84148a );
 a84155a <=( (not A299)  and  A298 );
 a84158a <=( A301  and  A300 );
 a84159a <=( a84158a  and  a84155a );
 a84160a <=( a84159a  and  a84152a );
 a84164a <=( (not A199)  and  (not A168) );
 a84165a <=( A170  and  a84164a );
 a84168a <=( (not A201)  and  A200 );
 a84171a <=( A203  and  (not A202) );
 a84172a <=( a84171a  and  a84168a );
 a84173a <=( a84172a  and  a84165a );
 a84176a <=( A266  and  (not A265) );
 a84179a <=( A268  and  A267 );
 a84180a <=( a84179a  and  a84176a );
 a84183a <=( (not A299)  and  A298 );
 a84186a <=( (not A302)  and  A300 );
 a84187a <=( a84186a  and  a84183a );
 a84188a <=( a84187a  and  a84180a );
 a84192a <=( (not A199)  and  (not A168) );
 a84193a <=( A170  and  a84192a );
 a84196a <=( (not A201)  and  A200 );
 a84199a <=( A203  and  (not A202) );
 a84200a <=( a84199a  and  a84196a );
 a84201a <=( a84200a  and  a84193a );
 a84204a <=( A266  and  (not A265) );
 a84207a <=( A268  and  A267 );
 a84208a <=( a84207a  and  a84204a );
 a84211a <=( A299  and  (not A298) );
 a84214a <=( A301  and  A300 );
 a84215a <=( a84214a  and  a84211a );
 a84216a <=( a84215a  and  a84208a );
 a84220a <=( (not A199)  and  (not A168) );
 a84221a <=( A170  and  a84220a );
 a84224a <=( (not A201)  and  A200 );
 a84227a <=( A203  and  (not A202) );
 a84228a <=( a84227a  and  a84224a );
 a84229a <=( a84228a  and  a84221a );
 a84232a <=( A266  and  (not A265) );
 a84235a <=( A268  and  A267 );
 a84236a <=( a84235a  and  a84232a );
 a84239a <=( A299  and  (not A298) );
 a84242a <=( (not A302)  and  A300 );
 a84243a <=( a84242a  and  a84239a );
 a84244a <=( a84243a  and  a84236a );
 a84248a <=( (not A199)  and  (not A168) );
 a84249a <=( A170  and  a84248a );
 a84252a <=( (not A201)  and  A200 );
 a84255a <=( A203  and  (not A202) );
 a84256a <=( a84255a  and  a84252a );
 a84257a <=( a84256a  and  a84249a );
 a84260a <=( A266  and  (not A265) );
 a84263a <=( (not A269)  and  A267 );
 a84264a <=( a84263a  and  a84260a );
 a84267a <=( (not A299)  and  A298 );
 a84270a <=( A301  and  A300 );
 a84271a <=( a84270a  and  a84267a );
 a84272a <=( a84271a  and  a84264a );
 a84276a <=( (not A199)  and  (not A168) );
 a84277a <=( A170  and  a84276a );
 a84280a <=( (not A201)  and  A200 );
 a84283a <=( A203  and  (not A202) );
 a84284a <=( a84283a  and  a84280a );
 a84285a <=( a84284a  and  a84277a );
 a84288a <=( A266  and  (not A265) );
 a84291a <=( (not A269)  and  A267 );
 a84292a <=( a84291a  and  a84288a );
 a84295a <=( (not A299)  and  A298 );
 a84298a <=( (not A302)  and  A300 );
 a84299a <=( a84298a  and  a84295a );
 a84300a <=( a84299a  and  a84292a );
 a84304a <=( (not A199)  and  (not A168) );
 a84305a <=( A170  and  a84304a );
 a84308a <=( (not A201)  and  A200 );
 a84311a <=( A203  and  (not A202) );
 a84312a <=( a84311a  and  a84308a );
 a84313a <=( a84312a  and  a84305a );
 a84316a <=( A266  and  (not A265) );
 a84319a <=( (not A269)  and  A267 );
 a84320a <=( a84319a  and  a84316a );
 a84323a <=( A299  and  (not A298) );
 a84326a <=( A301  and  A300 );
 a84327a <=( a84326a  and  a84323a );
 a84328a <=( a84327a  and  a84320a );
 a84332a <=( (not A199)  and  (not A168) );
 a84333a <=( A170  and  a84332a );
 a84336a <=( (not A201)  and  A200 );
 a84339a <=( A203  and  (not A202) );
 a84340a <=( a84339a  and  a84336a );
 a84341a <=( a84340a  and  a84333a );
 a84344a <=( A266  and  (not A265) );
 a84347a <=( (not A269)  and  A267 );
 a84348a <=( a84347a  and  a84344a );
 a84351a <=( A299  and  (not A298) );
 a84354a <=( (not A302)  and  A300 );
 a84355a <=( a84354a  and  a84351a );
 a84356a <=( a84355a  and  a84348a );
 a84360a <=( (not A199)  and  (not A168) );
 a84361a <=( A170  and  a84360a );
 a84364a <=( (not A201)  and  A200 );
 a84367a <=( A203  and  (not A202) );
 a84368a <=( a84367a  and  a84364a );
 a84369a <=( a84368a  and  a84361a );
 a84372a <=( (not A266)  and  A265 );
 a84375a <=( A268  and  A267 );
 a84376a <=( a84375a  and  a84372a );
 a84379a <=( (not A299)  and  A298 );
 a84382a <=( A301  and  A300 );
 a84383a <=( a84382a  and  a84379a );
 a84384a <=( a84383a  and  a84376a );
 a84388a <=( (not A199)  and  (not A168) );
 a84389a <=( A170  and  a84388a );
 a84392a <=( (not A201)  and  A200 );
 a84395a <=( A203  and  (not A202) );
 a84396a <=( a84395a  and  a84392a );
 a84397a <=( a84396a  and  a84389a );
 a84400a <=( (not A266)  and  A265 );
 a84403a <=( A268  and  A267 );
 a84404a <=( a84403a  and  a84400a );
 a84407a <=( (not A299)  and  A298 );
 a84410a <=( (not A302)  and  A300 );
 a84411a <=( a84410a  and  a84407a );
 a84412a <=( a84411a  and  a84404a );
 a84416a <=( (not A199)  and  (not A168) );
 a84417a <=( A170  and  a84416a );
 a84420a <=( (not A201)  and  A200 );
 a84423a <=( A203  and  (not A202) );
 a84424a <=( a84423a  and  a84420a );
 a84425a <=( a84424a  and  a84417a );
 a84428a <=( (not A266)  and  A265 );
 a84431a <=( A268  and  A267 );
 a84432a <=( a84431a  and  a84428a );
 a84435a <=( A299  and  (not A298) );
 a84438a <=( A301  and  A300 );
 a84439a <=( a84438a  and  a84435a );
 a84440a <=( a84439a  and  a84432a );
 a84444a <=( (not A199)  and  (not A168) );
 a84445a <=( A170  and  a84444a );
 a84448a <=( (not A201)  and  A200 );
 a84451a <=( A203  and  (not A202) );
 a84452a <=( a84451a  and  a84448a );
 a84453a <=( a84452a  and  a84445a );
 a84456a <=( (not A266)  and  A265 );
 a84459a <=( A268  and  A267 );
 a84460a <=( a84459a  and  a84456a );
 a84463a <=( A299  and  (not A298) );
 a84466a <=( (not A302)  and  A300 );
 a84467a <=( a84466a  and  a84463a );
 a84468a <=( a84467a  and  a84460a );
 a84472a <=( (not A199)  and  (not A168) );
 a84473a <=( A170  and  a84472a );
 a84476a <=( (not A201)  and  A200 );
 a84479a <=( A203  and  (not A202) );
 a84480a <=( a84479a  and  a84476a );
 a84481a <=( a84480a  and  a84473a );
 a84484a <=( (not A266)  and  A265 );
 a84487a <=( (not A269)  and  A267 );
 a84488a <=( a84487a  and  a84484a );
 a84491a <=( (not A299)  and  A298 );
 a84494a <=( A301  and  A300 );
 a84495a <=( a84494a  and  a84491a );
 a84496a <=( a84495a  and  a84488a );
 a84500a <=( (not A199)  and  (not A168) );
 a84501a <=( A170  and  a84500a );
 a84504a <=( (not A201)  and  A200 );
 a84507a <=( A203  and  (not A202) );
 a84508a <=( a84507a  and  a84504a );
 a84509a <=( a84508a  and  a84501a );
 a84512a <=( (not A266)  and  A265 );
 a84515a <=( (not A269)  and  A267 );
 a84516a <=( a84515a  and  a84512a );
 a84519a <=( (not A299)  and  A298 );
 a84522a <=( (not A302)  and  A300 );
 a84523a <=( a84522a  and  a84519a );
 a84524a <=( a84523a  and  a84516a );
 a84528a <=( (not A199)  and  (not A168) );
 a84529a <=( A170  and  a84528a );
 a84532a <=( (not A201)  and  A200 );
 a84535a <=( A203  and  (not A202) );
 a84536a <=( a84535a  and  a84532a );
 a84537a <=( a84536a  and  a84529a );
 a84540a <=( (not A266)  and  A265 );
 a84543a <=( (not A269)  and  A267 );
 a84544a <=( a84543a  and  a84540a );
 a84547a <=( A299  and  (not A298) );
 a84550a <=( A301  and  A300 );
 a84551a <=( a84550a  and  a84547a );
 a84552a <=( a84551a  and  a84544a );
 a84556a <=( (not A199)  and  (not A168) );
 a84557a <=( A170  and  a84556a );
 a84560a <=( (not A201)  and  A200 );
 a84563a <=( A203  and  (not A202) );
 a84564a <=( a84563a  and  a84560a );
 a84565a <=( a84564a  and  a84557a );
 a84568a <=( (not A266)  and  A265 );
 a84571a <=( (not A269)  and  A267 );
 a84572a <=( a84571a  and  a84568a );
 a84575a <=( A299  and  (not A298) );
 a84578a <=( (not A302)  and  A300 );
 a84579a <=( a84578a  and  a84575a );
 a84580a <=( a84579a  and  a84572a );
 a84584a <=( A199  and  (not A168) );
 a84585a <=( A170  and  a84584a );
 a84588a <=( A201  and  (not A200) );
 a84591a <=( (not A265)  and  A202 );
 a84592a <=( a84591a  and  a84588a );
 a84593a <=( a84592a  and  a84585a );
 a84596a <=( A267  and  A266 );
 a84599a <=( A298  and  A268 );
 a84600a <=( a84599a  and  a84596a );
 a84603a <=( (not A300)  and  (not A299) );
 a84606a <=( A302  and  (not A301) );
 a84607a <=( a84606a  and  a84603a );
 a84608a <=( a84607a  and  a84600a );
 a84612a <=( A199  and  (not A168) );
 a84613a <=( A170  and  a84612a );
 a84616a <=( A201  and  (not A200) );
 a84619a <=( (not A265)  and  A202 );
 a84620a <=( a84619a  and  a84616a );
 a84621a <=( a84620a  and  a84613a );
 a84624a <=( A267  and  A266 );
 a84627a <=( (not A298)  and  A268 );
 a84628a <=( a84627a  and  a84624a );
 a84631a <=( (not A300)  and  A299 );
 a84634a <=( A302  and  (not A301) );
 a84635a <=( a84634a  and  a84631a );
 a84636a <=( a84635a  and  a84628a );
 a84640a <=( A199  and  (not A168) );
 a84641a <=( A170  and  a84640a );
 a84644a <=( A201  and  (not A200) );
 a84647a <=( (not A265)  and  A202 );
 a84648a <=( a84647a  and  a84644a );
 a84649a <=( a84648a  and  a84641a );
 a84652a <=( A267  and  A266 );
 a84655a <=( A298  and  (not A269) );
 a84656a <=( a84655a  and  a84652a );
 a84659a <=( (not A300)  and  (not A299) );
 a84662a <=( A302  and  (not A301) );
 a84663a <=( a84662a  and  a84659a );
 a84664a <=( a84663a  and  a84656a );
 a84668a <=( A199  and  (not A168) );
 a84669a <=( A170  and  a84668a );
 a84672a <=( A201  and  (not A200) );
 a84675a <=( (not A265)  and  A202 );
 a84676a <=( a84675a  and  a84672a );
 a84677a <=( a84676a  and  a84669a );
 a84680a <=( A267  and  A266 );
 a84683a <=( (not A298)  and  (not A269) );
 a84684a <=( a84683a  and  a84680a );
 a84687a <=( (not A300)  and  A299 );
 a84690a <=( A302  and  (not A301) );
 a84691a <=( a84690a  and  a84687a );
 a84692a <=( a84691a  and  a84684a );
 a84696a <=( A199  and  (not A168) );
 a84697a <=( A170  and  a84696a );
 a84700a <=( A201  and  (not A200) );
 a84703a <=( (not A265)  and  A202 );
 a84704a <=( a84703a  and  a84700a );
 a84705a <=( a84704a  and  a84697a );
 a84708a <=( (not A267)  and  A266 );
 a84711a <=( A269  and  (not A268) );
 a84712a <=( a84711a  and  a84708a );
 a84715a <=( (not A299)  and  A298 );
 a84718a <=( A301  and  A300 );
 a84719a <=( a84718a  and  a84715a );
 a84720a <=( a84719a  and  a84712a );
 a84724a <=( A199  and  (not A168) );
 a84725a <=( A170  and  a84724a );
 a84728a <=( A201  and  (not A200) );
 a84731a <=( (not A265)  and  A202 );
 a84732a <=( a84731a  and  a84728a );
 a84733a <=( a84732a  and  a84725a );
 a84736a <=( (not A267)  and  A266 );
 a84739a <=( A269  and  (not A268) );
 a84740a <=( a84739a  and  a84736a );
 a84743a <=( (not A299)  and  A298 );
 a84746a <=( (not A302)  and  A300 );
 a84747a <=( a84746a  and  a84743a );
 a84748a <=( a84747a  and  a84740a );
 a84752a <=( A199  and  (not A168) );
 a84753a <=( A170  and  a84752a );
 a84756a <=( A201  and  (not A200) );
 a84759a <=( (not A265)  and  A202 );
 a84760a <=( a84759a  and  a84756a );
 a84761a <=( a84760a  and  a84753a );
 a84764a <=( (not A267)  and  A266 );
 a84767a <=( A269  and  (not A268) );
 a84768a <=( a84767a  and  a84764a );
 a84771a <=( A299  and  (not A298) );
 a84774a <=( A301  and  A300 );
 a84775a <=( a84774a  and  a84771a );
 a84776a <=( a84775a  and  a84768a );
 a84780a <=( A199  and  (not A168) );
 a84781a <=( A170  and  a84780a );
 a84784a <=( A201  and  (not A200) );
 a84787a <=( (not A265)  and  A202 );
 a84788a <=( a84787a  and  a84784a );
 a84789a <=( a84788a  and  a84781a );
 a84792a <=( (not A267)  and  A266 );
 a84795a <=( A269  and  (not A268) );
 a84796a <=( a84795a  and  a84792a );
 a84799a <=( A299  and  (not A298) );
 a84802a <=( (not A302)  and  A300 );
 a84803a <=( a84802a  and  a84799a );
 a84804a <=( a84803a  and  a84796a );
 a84808a <=( A199  and  (not A168) );
 a84809a <=( A170  and  a84808a );
 a84812a <=( A201  and  (not A200) );
 a84815a <=( A265  and  A202 );
 a84816a <=( a84815a  and  a84812a );
 a84817a <=( a84816a  and  a84809a );
 a84820a <=( A267  and  (not A266) );
 a84823a <=( A298  and  A268 );
 a84824a <=( a84823a  and  a84820a );
 a84827a <=( (not A300)  and  (not A299) );
 a84830a <=( A302  and  (not A301) );
 a84831a <=( a84830a  and  a84827a );
 a84832a <=( a84831a  and  a84824a );
 a84836a <=( A199  and  (not A168) );
 a84837a <=( A170  and  a84836a );
 a84840a <=( A201  and  (not A200) );
 a84843a <=( A265  and  A202 );
 a84844a <=( a84843a  and  a84840a );
 a84845a <=( a84844a  and  a84837a );
 a84848a <=( A267  and  (not A266) );
 a84851a <=( (not A298)  and  A268 );
 a84852a <=( a84851a  and  a84848a );
 a84855a <=( (not A300)  and  A299 );
 a84858a <=( A302  and  (not A301) );
 a84859a <=( a84858a  and  a84855a );
 a84860a <=( a84859a  and  a84852a );
 a84864a <=( A199  and  (not A168) );
 a84865a <=( A170  and  a84864a );
 a84868a <=( A201  and  (not A200) );
 a84871a <=( A265  and  A202 );
 a84872a <=( a84871a  and  a84868a );
 a84873a <=( a84872a  and  a84865a );
 a84876a <=( A267  and  (not A266) );
 a84879a <=( A298  and  (not A269) );
 a84880a <=( a84879a  and  a84876a );
 a84883a <=( (not A300)  and  (not A299) );
 a84886a <=( A302  and  (not A301) );
 a84887a <=( a84886a  and  a84883a );
 a84888a <=( a84887a  and  a84880a );
 a84892a <=( A199  and  (not A168) );
 a84893a <=( A170  and  a84892a );
 a84896a <=( A201  and  (not A200) );
 a84899a <=( A265  and  A202 );
 a84900a <=( a84899a  and  a84896a );
 a84901a <=( a84900a  and  a84893a );
 a84904a <=( A267  and  (not A266) );
 a84907a <=( (not A298)  and  (not A269) );
 a84908a <=( a84907a  and  a84904a );
 a84911a <=( (not A300)  and  A299 );
 a84914a <=( A302  and  (not A301) );
 a84915a <=( a84914a  and  a84911a );
 a84916a <=( a84915a  and  a84908a );
 a84920a <=( A199  and  (not A168) );
 a84921a <=( A170  and  a84920a );
 a84924a <=( A201  and  (not A200) );
 a84927a <=( A265  and  A202 );
 a84928a <=( a84927a  and  a84924a );
 a84929a <=( a84928a  and  a84921a );
 a84932a <=( (not A267)  and  (not A266) );
 a84935a <=( A269  and  (not A268) );
 a84936a <=( a84935a  and  a84932a );
 a84939a <=( (not A299)  and  A298 );
 a84942a <=( A301  and  A300 );
 a84943a <=( a84942a  and  a84939a );
 a84944a <=( a84943a  and  a84936a );
 a84948a <=( A199  and  (not A168) );
 a84949a <=( A170  and  a84948a );
 a84952a <=( A201  and  (not A200) );
 a84955a <=( A265  and  A202 );
 a84956a <=( a84955a  and  a84952a );
 a84957a <=( a84956a  and  a84949a );
 a84960a <=( (not A267)  and  (not A266) );
 a84963a <=( A269  and  (not A268) );
 a84964a <=( a84963a  and  a84960a );
 a84967a <=( (not A299)  and  A298 );
 a84970a <=( (not A302)  and  A300 );
 a84971a <=( a84970a  and  a84967a );
 a84972a <=( a84971a  and  a84964a );
 a84976a <=( A199  and  (not A168) );
 a84977a <=( A170  and  a84976a );
 a84980a <=( A201  and  (not A200) );
 a84983a <=( A265  and  A202 );
 a84984a <=( a84983a  and  a84980a );
 a84985a <=( a84984a  and  a84977a );
 a84988a <=( (not A267)  and  (not A266) );
 a84991a <=( A269  and  (not A268) );
 a84992a <=( a84991a  and  a84988a );
 a84995a <=( A299  and  (not A298) );
 a84998a <=( A301  and  A300 );
 a84999a <=( a84998a  and  a84995a );
 a85000a <=( a84999a  and  a84992a );
 a85004a <=( A199  and  (not A168) );
 a85005a <=( A170  and  a85004a );
 a85008a <=( A201  and  (not A200) );
 a85011a <=( A265  and  A202 );
 a85012a <=( a85011a  and  a85008a );
 a85013a <=( a85012a  and  a85005a );
 a85016a <=( (not A267)  and  (not A266) );
 a85019a <=( A269  and  (not A268) );
 a85020a <=( a85019a  and  a85016a );
 a85023a <=( A299  and  (not A298) );
 a85026a <=( (not A302)  and  A300 );
 a85027a <=( a85026a  and  a85023a );
 a85028a <=( a85027a  and  a85020a );
 a85032a <=( A199  and  (not A168) );
 a85033a <=( A170  and  a85032a );
 a85036a <=( A201  and  (not A200) );
 a85039a <=( (not A265)  and  (not A203) );
 a85040a <=( a85039a  and  a85036a );
 a85041a <=( a85040a  and  a85033a );
 a85044a <=( A267  and  A266 );
 a85047a <=( A298  and  A268 );
 a85048a <=( a85047a  and  a85044a );
 a85051a <=( (not A300)  and  (not A299) );
 a85054a <=( A302  and  (not A301) );
 a85055a <=( a85054a  and  a85051a );
 a85056a <=( a85055a  and  a85048a );
 a85060a <=( A199  and  (not A168) );
 a85061a <=( A170  and  a85060a );
 a85064a <=( A201  and  (not A200) );
 a85067a <=( (not A265)  and  (not A203) );
 a85068a <=( a85067a  and  a85064a );
 a85069a <=( a85068a  and  a85061a );
 a85072a <=( A267  and  A266 );
 a85075a <=( (not A298)  and  A268 );
 a85076a <=( a85075a  and  a85072a );
 a85079a <=( (not A300)  and  A299 );
 a85082a <=( A302  and  (not A301) );
 a85083a <=( a85082a  and  a85079a );
 a85084a <=( a85083a  and  a85076a );
 a85088a <=( A199  and  (not A168) );
 a85089a <=( A170  and  a85088a );
 a85092a <=( A201  and  (not A200) );
 a85095a <=( (not A265)  and  (not A203) );
 a85096a <=( a85095a  and  a85092a );
 a85097a <=( a85096a  and  a85089a );
 a85100a <=( A267  and  A266 );
 a85103a <=( A298  and  (not A269) );
 a85104a <=( a85103a  and  a85100a );
 a85107a <=( (not A300)  and  (not A299) );
 a85110a <=( A302  and  (not A301) );
 a85111a <=( a85110a  and  a85107a );
 a85112a <=( a85111a  and  a85104a );
 a85116a <=( A199  and  (not A168) );
 a85117a <=( A170  and  a85116a );
 a85120a <=( A201  and  (not A200) );
 a85123a <=( (not A265)  and  (not A203) );
 a85124a <=( a85123a  and  a85120a );
 a85125a <=( a85124a  and  a85117a );
 a85128a <=( A267  and  A266 );
 a85131a <=( (not A298)  and  (not A269) );
 a85132a <=( a85131a  and  a85128a );
 a85135a <=( (not A300)  and  A299 );
 a85138a <=( A302  and  (not A301) );
 a85139a <=( a85138a  and  a85135a );
 a85140a <=( a85139a  and  a85132a );
 a85144a <=( A199  and  (not A168) );
 a85145a <=( A170  and  a85144a );
 a85148a <=( A201  and  (not A200) );
 a85151a <=( (not A265)  and  (not A203) );
 a85152a <=( a85151a  and  a85148a );
 a85153a <=( a85152a  and  a85145a );
 a85156a <=( (not A267)  and  A266 );
 a85159a <=( A269  and  (not A268) );
 a85160a <=( a85159a  and  a85156a );
 a85163a <=( (not A299)  and  A298 );
 a85166a <=( A301  and  A300 );
 a85167a <=( a85166a  and  a85163a );
 a85168a <=( a85167a  and  a85160a );
 a85172a <=( A199  and  (not A168) );
 a85173a <=( A170  and  a85172a );
 a85176a <=( A201  and  (not A200) );
 a85179a <=( (not A265)  and  (not A203) );
 a85180a <=( a85179a  and  a85176a );
 a85181a <=( a85180a  and  a85173a );
 a85184a <=( (not A267)  and  A266 );
 a85187a <=( A269  and  (not A268) );
 a85188a <=( a85187a  and  a85184a );
 a85191a <=( (not A299)  and  A298 );
 a85194a <=( (not A302)  and  A300 );
 a85195a <=( a85194a  and  a85191a );
 a85196a <=( a85195a  and  a85188a );
 a85200a <=( A199  and  (not A168) );
 a85201a <=( A170  and  a85200a );
 a85204a <=( A201  and  (not A200) );
 a85207a <=( (not A265)  and  (not A203) );
 a85208a <=( a85207a  and  a85204a );
 a85209a <=( a85208a  and  a85201a );
 a85212a <=( (not A267)  and  A266 );
 a85215a <=( A269  and  (not A268) );
 a85216a <=( a85215a  and  a85212a );
 a85219a <=( A299  and  (not A298) );
 a85222a <=( A301  and  A300 );
 a85223a <=( a85222a  and  a85219a );
 a85224a <=( a85223a  and  a85216a );
 a85228a <=( A199  and  (not A168) );
 a85229a <=( A170  and  a85228a );
 a85232a <=( A201  and  (not A200) );
 a85235a <=( (not A265)  and  (not A203) );
 a85236a <=( a85235a  and  a85232a );
 a85237a <=( a85236a  and  a85229a );
 a85240a <=( (not A267)  and  A266 );
 a85243a <=( A269  and  (not A268) );
 a85244a <=( a85243a  and  a85240a );
 a85247a <=( A299  and  (not A298) );
 a85250a <=( (not A302)  and  A300 );
 a85251a <=( a85250a  and  a85247a );
 a85252a <=( a85251a  and  a85244a );
 a85256a <=( A199  and  (not A168) );
 a85257a <=( A170  and  a85256a );
 a85260a <=( A201  and  (not A200) );
 a85263a <=( A265  and  (not A203) );
 a85264a <=( a85263a  and  a85260a );
 a85265a <=( a85264a  and  a85257a );
 a85268a <=( A267  and  (not A266) );
 a85271a <=( A298  and  A268 );
 a85272a <=( a85271a  and  a85268a );
 a85275a <=( (not A300)  and  (not A299) );
 a85278a <=( A302  and  (not A301) );
 a85279a <=( a85278a  and  a85275a );
 a85280a <=( a85279a  and  a85272a );
 a85284a <=( A199  and  (not A168) );
 a85285a <=( A170  and  a85284a );
 a85288a <=( A201  and  (not A200) );
 a85291a <=( A265  and  (not A203) );
 a85292a <=( a85291a  and  a85288a );
 a85293a <=( a85292a  and  a85285a );
 a85296a <=( A267  and  (not A266) );
 a85299a <=( (not A298)  and  A268 );
 a85300a <=( a85299a  and  a85296a );
 a85303a <=( (not A300)  and  A299 );
 a85306a <=( A302  and  (not A301) );
 a85307a <=( a85306a  and  a85303a );
 a85308a <=( a85307a  and  a85300a );
 a85312a <=( A199  and  (not A168) );
 a85313a <=( A170  and  a85312a );
 a85316a <=( A201  and  (not A200) );
 a85319a <=( A265  and  (not A203) );
 a85320a <=( a85319a  and  a85316a );
 a85321a <=( a85320a  and  a85313a );
 a85324a <=( A267  and  (not A266) );
 a85327a <=( A298  and  (not A269) );
 a85328a <=( a85327a  and  a85324a );
 a85331a <=( (not A300)  and  (not A299) );
 a85334a <=( A302  and  (not A301) );
 a85335a <=( a85334a  and  a85331a );
 a85336a <=( a85335a  and  a85328a );
 a85340a <=( A199  and  (not A168) );
 a85341a <=( A170  and  a85340a );
 a85344a <=( A201  and  (not A200) );
 a85347a <=( A265  and  (not A203) );
 a85348a <=( a85347a  and  a85344a );
 a85349a <=( a85348a  and  a85341a );
 a85352a <=( A267  and  (not A266) );
 a85355a <=( (not A298)  and  (not A269) );
 a85356a <=( a85355a  and  a85352a );
 a85359a <=( (not A300)  and  A299 );
 a85362a <=( A302  and  (not A301) );
 a85363a <=( a85362a  and  a85359a );
 a85364a <=( a85363a  and  a85356a );
 a85368a <=( A199  and  (not A168) );
 a85369a <=( A170  and  a85368a );
 a85372a <=( A201  and  (not A200) );
 a85375a <=( A265  and  (not A203) );
 a85376a <=( a85375a  and  a85372a );
 a85377a <=( a85376a  and  a85369a );
 a85380a <=( (not A267)  and  (not A266) );
 a85383a <=( A269  and  (not A268) );
 a85384a <=( a85383a  and  a85380a );
 a85387a <=( (not A299)  and  A298 );
 a85390a <=( A301  and  A300 );
 a85391a <=( a85390a  and  a85387a );
 a85392a <=( a85391a  and  a85384a );
 a85396a <=( A199  and  (not A168) );
 a85397a <=( A170  and  a85396a );
 a85400a <=( A201  and  (not A200) );
 a85403a <=( A265  and  (not A203) );
 a85404a <=( a85403a  and  a85400a );
 a85405a <=( a85404a  and  a85397a );
 a85408a <=( (not A267)  and  (not A266) );
 a85411a <=( A269  and  (not A268) );
 a85412a <=( a85411a  and  a85408a );
 a85415a <=( (not A299)  and  A298 );
 a85418a <=( (not A302)  and  A300 );
 a85419a <=( a85418a  and  a85415a );
 a85420a <=( a85419a  and  a85412a );
 a85424a <=( A199  and  (not A168) );
 a85425a <=( A170  and  a85424a );
 a85428a <=( A201  and  (not A200) );
 a85431a <=( A265  and  (not A203) );
 a85432a <=( a85431a  and  a85428a );
 a85433a <=( a85432a  and  a85425a );
 a85436a <=( (not A267)  and  (not A266) );
 a85439a <=( A269  and  (not A268) );
 a85440a <=( a85439a  and  a85436a );
 a85443a <=( A299  and  (not A298) );
 a85446a <=( A301  and  A300 );
 a85447a <=( a85446a  and  a85443a );
 a85448a <=( a85447a  and  a85440a );
 a85452a <=( A199  and  (not A168) );
 a85453a <=( A170  and  a85452a );
 a85456a <=( A201  and  (not A200) );
 a85459a <=( A265  and  (not A203) );
 a85460a <=( a85459a  and  a85456a );
 a85461a <=( a85460a  and  a85453a );
 a85464a <=( (not A267)  and  (not A266) );
 a85467a <=( A269  and  (not A268) );
 a85468a <=( a85467a  and  a85464a );
 a85471a <=( A299  and  (not A298) );
 a85474a <=( (not A302)  and  A300 );
 a85475a <=( a85474a  and  a85471a );
 a85476a <=( a85475a  and  a85468a );
 a85480a <=( A199  and  (not A168) );
 a85481a <=( A170  and  a85480a );
 a85484a <=( (not A201)  and  (not A200) );
 a85487a <=( A203  and  (not A202) );
 a85488a <=( a85487a  and  a85484a );
 a85489a <=( a85488a  and  a85481a );
 a85492a <=( A266  and  (not A265) );
 a85495a <=( A268  and  A267 );
 a85496a <=( a85495a  and  a85492a );
 a85499a <=( (not A299)  and  A298 );
 a85502a <=( A301  and  A300 );
 a85503a <=( a85502a  and  a85499a );
 a85504a <=( a85503a  and  a85496a );
 a85508a <=( A199  and  (not A168) );
 a85509a <=( A170  and  a85508a );
 a85512a <=( (not A201)  and  (not A200) );
 a85515a <=( A203  and  (not A202) );
 a85516a <=( a85515a  and  a85512a );
 a85517a <=( a85516a  and  a85509a );
 a85520a <=( A266  and  (not A265) );
 a85523a <=( A268  and  A267 );
 a85524a <=( a85523a  and  a85520a );
 a85527a <=( (not A299)  and  A298 );
 a85530a <=( (not A302)  and  A300 );
 a85531a <=( a85530a  and  a85527a );
 a85532a <=( a85531a  and  a85524a );
 a85536a <=( A199  and  (not A168) );
 a85537a <=( A170  and  a85536a );
 a85540a <=( (not A201)  and  (not A200) );
 a85543a <=( A203  and  (not A202) );
 a85544a <=( a85543a  and  a85540a );
 a85545a <=( a85544a  and  a85537a );
 a85548a <=( A266  and  (not A265) );
 a85551a <=( A268  and  A267 );
 a85552a <=( a85551a  and  a85548a );
 a85555a <=( A299  and  (not A298) );
 a85558a <=( A301  and  A300 );
 a85559a <=( a85558a  and  a85555a );
 a85560a <=( a85559a  and  a85552a );
 a85564a <=( A199  and  (not A168) );
 a85565a <=( A170  and  a85564a );
 a85568a <=( (not A201)  and  (not A200) );
 a85571a <=( A203  and  (not A202) );
 a85572a <=( a85571a  and  a85568a );
 a85573a <=( a85572a  and  a85565a );
 a85576a <=( A266  and  (not A265) );
 a85579a <=( A268  and  A267 );
 a85580a <=( a85579a  and  a85576a );
 a85583a <=( A299  and  (not A298) );
 a85586a <=( (not A302)  and  A300 );
 a85587a <=( a85586a  and  a85583a );
 a85588a <=( a85587a  and  a85580a );
 a85592a <=( A199  and  (not A168) );
 a85593a <=( A170  and  a85592a );
 a85596a <=( (not A201)  and  (not A200) );
 a85599a <=( A203  and  (not A202) );
 a85600a <=( a85599a  and  a85596a );
 a85601a <=( a85600a  and  a85593a );
 a85604a <=( A266  and  (not A265) );
 a85607a <=( (not A269)  and  A267 );
 a85608a <=( a85607a  and  a85604a );
 a85611a <=( (not A299)  and  A298 );
 a85614a <=( A301  and  A300 );
 a85615a <=( a85614a  and  a85611a );
 a85616a <=( a85615a  and  a85608a );
 a85620a <=( A199  and  (not A168) );
 a85621a <=( A170  and  a85620a );
 a85624a <=( (not A201)  and  (not A200) );
 a85627a <=( A203  and  (not A202) );
 a85628a <=( a85627a  and  a85624a );
 a85629a <=( a85628a  and  a85621a );
 a85632a <=( A266  and  (not A265) );
 a85635a <=( (not A269)  and  A267 );
 a85636a <=( a85635a  and  a85632a );
 a85639a <=( (not A299)  and  A298 );
 a85642a <=( (not A302)  and  A300 );
 a85643a <=( a85642a  and  a85639a );
 a85644a <=( a85643a  and  a85636a );
 a85648a <=( A199  and  (not A168) );
 a85649a <=( A170  and  a85648a );
 a85652a <=( (not A201)  and  (not A200) );
 a85655a <=( A203  and  (not A202) );
 a85656a <=( a85655a  and  a85652a );
 a85657a <=( a85656a  and  a85649a );
 a85660a <=( A266  and  (not A265) );
 a85663a <=( (not A269)  and  A267 );
 a85664a <=( a85663a  and  a85660a );
 a85667a <=( A299  and  (not A298) );
 a85670a <=( A301  and  A300 );
 a85671a <=( a85670a  and  a85667a );
 a85672a <=( a85671a  and  a85664a );
 a85676a <=( A199  and  (not A168) );
 a85677a <=( A170  and  a85676a );
 a85680a <=( (not A201)  and  (not A200) );
 a85683a <=( A203  and  (not A202) );
 a85684a <=( a85683a  and  a85680a );
 a85685a <=( a85684a  and  a85677a );
 a85688a <=( A266  and  (not A265) );
 a85691a <=( (not A269)  and  A267 );
 a85692a <=( a85691a  and  a85688a );
 a85695a <=( A299  and  (not A298) );
 a85698a <=( (not A302)  and  A300 );
 a85699a <=( a85698a  and  a85695a );
 a85700a <=( a85699a  and  a85692a );
 a85704a <=( A199  and  (not A168) );
 a85705a <=( A170  and  a85704a );
 a85708a <=( (not A201)  and  (not A200) );
 a85711a <=( A203  and  (not A202) );
 a85712a <=( a85711a  and  a85708a );
 a85713a <=( a85712a  and  a85705a );
 a85716a <=( (not A266)  and  A265 );
 a85719a <=( A268  and  A267 );
 a85720a <=( a85719a  and  a85716a );
 a85723a <=( (not A299)  and  A298 );
 a85726a <=( A301  and  A300 );
 a85727a <=( a85726a  and  a85723a );
 a85728a <=( a85727a  and  a85720a );
 a85732a <=( A199  and  (not A168) );
 a85733a <=( A170  and  a85732a );
 a85736a <=( (not A201)  and  (not A200) );
 a85739a <=( A203  and  (not A202) );
 a85740a <=( a85739a  and  a85736a );
 a85741a <=( a85740a  and  a85733a );
 a85744a <=( (not A266)  and  A265 );
 a85747a <=( A268  and  A267 );
 a85748a <=( a85747a  and  a85744a );
 a85751a <=( (not A299)  and  A298 );
 a85754a <=( (not A302)  and  A300 );
 a85755a <=( a85754a  and  a85751a );
 a85756a <=( a85755a  and  a85748a );
 a85760a <=( A199  and  (not A168) );
 a85761a <=( A170  and  a85760a );
 a85764a <=( (not A201)  and  (not A200) );
 a85767a <=( A203  and  (not A202) );
 a85768a <=( a85767a  and  a85764a );
 a85769a <=( a85768a  and  a85761a );
 a85772a <=( (not A266)  and  A265 );
 a85775a <=( A268  and  A267 );
 a85776a <=( a85775a  and  a85772a );
 a85779a <=( A299  and  (not A298) );
 a85782a <=( A301  and  A300 );
 a85783a <=( a85782a  and  a85779a );
 a85784a <=( a85783a  and  a85776a );
 a85788a <=( A199  and  (not A168) );
 a85789a <=( A170  and  a85788a );
 a85792a <=( (not A201)  and  (not A200) );
 a85795a <=( A203  and  (not A202) );
 a85796a <=( a85795a  and  a85792a );
 a85797a <=( a85796a  and  a85789a );
 a85800a <=( (not A266)  and  A265 );
 a85803a <=( A268  and  A267 );
 a85804a <=( a85803a  and  a85800a );
 a85807a <=( A299  and  (not A298) );
 a85810a <=( (not A302)  and  A300 );
 a85811a <=( a85810a  and  a85807a );
 a85812a <=( a85811a  and  a85804a );
 a85816a <=( A199  and  (not A168) );
 a85817a <=( A170  and  a85816a );
 a85820a <=( (not A201)  and  (not A200) );
 a85823a <=( A203  and  (not A202) );
 a85824a <=( a85823a  and  a85820a );
 a85825a <=( a85824a  and  a85817a );
 a85828a <=( (not A266)  and  A265 );
 a85831a <=( (not A269)  and  A267 );
 a85832a <=( a85831a  and  a85828a );
 a85835a <=( (not A299)  and  A298 );
 a85838a <=( A301  and  A300 );
 a85839a <=( a85838a  and  a85835a );
 a85840a <=( a85839a  and  a85832a );
 a85844a <=( A199  and  (not A168) );
 a85845a <=( A170  and  a85844a );
 a85848a <=( (not A201)  and  (not A200) );
 a85851a <=( A203  and  (not A202) );
 a85852a <=( a85851a  and  a85848a );
 a85853a <=( a85852a  and  a85845a );
 a85856a <=( (not A266)  and  A265 );
 a85859a <=( (not A269)  and  A267 );
 a85860a <=( a85859a  and  a85856a );
 a85863a <=( (not A299)  and  A298 );
 a85866a <=( (not A302)  and  A300 );
 a85867a <=( a85866a  and  a85863a );
 a85868a <=( a85867a  and  a85860a );
 a85872a <=( A199  and  (not A168) );
 a85873a <=( A170  and  a85872a );
 a85876a <=( (not A201)  and  (not A200) );
 a85879a <=( A203  and  (not A202) );
 a85880a <=( a85879a  and  a85876a );
 a85881a <=( a85880a  and  a85873a );
 a85884a <=( (not A266)  and  A265 );
 a85887a <=( (not A269)  and  A267 );
 a85888a <=( a85887a  and  a85884a );
 a85891a <=( A299  and  (not A298) );
 a85894a <=( A301  and  A300 );
 a85895a <=( a85894a  and  a85891a );
 a85896a <=( a85895a  and  a85888a );
 a85900a <=( A199  and  (not A168) );
 a85901a <=( A170  and  a85900a );
 a85904a <=( (not A201)  and  (not A200) );
 a85907a <=( A203  and  (not A202) );
 a85908a <=( a85907a  and  a85904a );
 a85909a <=( a85908a  and  a85901a );
 a85912a <=( (not A266)  and  A265 );
 a85915a <=( (not A269)  and  A267 );
 a85916a <=( a85915a  and  a85912a );
 a85919a <=( A299  and  (not A298) );
 a85922a <=( (not A302)  and  A300 );
 a85923a <=( a85922a  and  a85919a );
 a85924a <=( a85923a  and  a85916a );
 a85928a <=( A167  and  A168 );
 a85929a <=( A169  and  a85928a );
 a85932a <=( A201  and  (not A166) );
 a85935a <=( A203  and  (not A202) );
 a85936a <=( a85935a  and  a85932a );
 a85937a <=( a85936a  and  a85929a );
 a85940a <=( (not A268)  and  A267 );
 a85943a <=( A298  and  A269 );
 a85944a <=( a85943a  and  a85940a );
 a85947a <=( (not A300)  and  (not A299) );
 a85950a <=( A302  and  (not A301) );
 a85951a <=( a85950a  and  a85947a );
 a85952a <=( a85951a  and  a85944a );
 a85956a <=( A167  and  A168 );
 a85957a <=( A169  and  a85956a );
 a85960a <=( A201  and  (not A166) );
 a85963a <=( A203  and  (not A202) );
 a85964a <=( a85963a  and  a85960a );
 a85965a <=( a85964a  and  a85957a );
 a85968a <=( (not A268)  and  A267 );
 a85971a <=( (not A298)  and  A269 );
 a85972a <=( a85971a  and  a85968a );
 a85975a <=( (not A300)  and  A299 );
 a85978a <=( A302  and  (not A301) );
 a85979a <=( a85978a  and  a85975a );
 a85980a <=( a85979a  and  a85972a );
 a85984a <=( A167  and  A168 );
 a85985a <=( A169  and  a85984a );
 a85988a <=( A201  and  (not A166) );
 a85991a <=( A203  and  (not A202) );
 a85992a <=( a85991a  and  a85988a );
 a85993a <=( a85992a  and  a85985a );
 a85996a <=( A266  and  (not A265) );
 a85999a <=( (not A268)  and  (not A267) );
 a86000a <=( a85999a  and  a85996a );
 a86003a <=( A300  and  A269 );
 a86006a <=( A302  and  (not A301) );
 a86007a <=( a86006a  and  a86003a );
 a86008a <=( a86007a  and  a86000a );
 a86012a <=( A167  and  A168 );
 a86013a <=( A169  and  a86012a );
 a86016a <=( A201  and  (not A166) );
 a86019a <=( A203  and  (not A202) );
 a86020a <=( a86019a  and  a86016a );
 a86021a <=( a86020a  and  a86013a );
 a86024a <=( (not A266)  and  A265 );
 a86027a <=( (not A268)  and  (not A267) );
 a86028a <=( a86027a  and  a86024a );
 a86031a <=( A300  and  A269 );
 a86034a <=( A302  and  (not A301) );
 a86035a <=( a86034a  and  a86031a );
 a86036a <=( a86035a  and  a86028a );
 a86040a <=( (not A167)  and  A168 );
 a86041a <=( A169  and  a86040a );
 a86044a <=( A201  and  A166 );
 a86047a <=( A203  and  (not A202) );
 a86048a <=( a86047a  and  a86044a );
 a86049a <=( a86048a  and  a86041a );
 a86052a <=( (not A268)  and  A267 );
 a86055a <=( A298  and  A269 );
 a86056a <=( a86055a  and  a86052a );
 a86059a <=( (not A300)  and  (not A299) );
 a86062a <=( A302  and  (not A301) );
 a86063a <=( a86062a  and  a86059a );
 a86064a <=( a86063a  and  a86056a );
 a86068a <=( (not A167)  and  A168 );
 a86069a <=( A169  and  a86068a );
 a86072a <=( A201  and  A166 );
 a86075a <=( A203  and  (not A202) );
 a86076a <=( a86075a  and  a86072a );
 a86077a <=( a86076a  and  a86069a );
 a86080a <=( (not A268)  and  A267 );
 a86083a <=( (not A298)  and  A269 );
 a86084a <=( a86083a  and  a86080a );
 a86087a <=( (not A300)  and  A299 );
 a86090a <=( A302  and  (not A301) );
 a86091a <=( a86090a  and  a86087a );
 a86092a <=( a86091a  and  a86084a );
 a86096a <=( (not A167)  and  A168 );
 a86097a <=( A169  and  a86096a );
 a86100a <=( A201  and  A166 );
 a86103a <=( A203  and  (not A202) );
 a86104a <=( a86103a  and  a86100a );
 a86105a <=( a86104a  and  a86097a );
 a86108a <=( A266  and  (not A265) );
 a86111a <=( (not A268)  and  (not A267) );
 a86112a <=( a86111a  and  a86108a );
 a86115a <=( A300  and  A269 );
 a86118a <=( A302  and  (not A301) );
 a86119a <=( a86118a  and  a86115a );
 a86120a <=( a86119a  and  a86112a );
 a86124a <=( (not A167)  and  A168 );
 a86125a <=( A169  and  a86124a );
 a86128a <=( A201  and  A166 );
 a86131a <=( A203  and  (not A202) );
 a86132a <=( a86131a  and  a86128a );
 a86133a <=( a86132a  and  a86125a );
 a86136a <=( (not A266)  and  A265 );
 a86139a <=( (not A268)  and  (not A267) );
 a86140a <=( a86139a  and  a86136a );
 a86143a <=( A300  and  A269 );
 a86146a <=( A302  and  (not A301) );
 a86147a <=( a86146a  and  a86143a );
 a86148a <=( a86147a  and  a86140a );
 a86152a <=( (not A199)  and  (not A168) );
 a86153a <=( A169  and  a86152a );
 a86156a <=( A201  and  A200 );
 a86159a <=( (not A265)  and  A202 );
 a86160a <=( a86159a  and  a86156a );
 a86161a <=( a86160a  and  a86153a );
 a86164a <=( A267  and  A266 );
 a86167a <=( A298  and  A268 );
 a86168a <=( a86167a  and  a86164a );
 a86171a <=( (not A300)  and  (not A299) );
 a86174a <=( A302  and  (not A301) );
 a86175a <=( a86174a  and  a86171a );
 a86176a <=( a86175a  and  a86168a );
 a86180a <=( (not A199)  and  (not A168) );
 a86181a <=( A169  and  a86180a );
 a86184a <=( A201  and  A200 );
 a86187a <=( (not A265)  and  A202 );
 a86188a <=( a86187a  and  a86184a );
 a86189a <=( a86188a  and  a86181a );
 a86192a <=( A267  and  A266 );
 a86195a <=( (not A298)  and  A268 );
 a86196a <=( a86195a  and  a86192a );
 a86199a <=( (not A300)  and  A299 );
 a86202a <=( A302  and  (not A301) );
 a86203a <=( a86202a  and  a86199a );
 a86204a <=( a86203a  and  a86196a );
 a86208a <=( (not A199)  and  (not A168) );
 a86209a <=( A169  and  a86208a );
 a86212a <=( A201  and  A200 );
 a86215a <=( (not A265)  and  A202 );
 a86216a <=( a86215a  and  a86212a );
 a86217a <=( a86216a  and  a86209a );
 a86220a <=( A267  and  A266 );
 a86223a <=( A298  and  (not A269) );
 a86224a <=( a86223a  and  a86220a );
 a86227a <=( (not A300)  and  (not A299) );
 a86230a <=( A302  and  (not A301) );
 a86231a <=( a86230a  and  a86227a );
 a86232a <=( a86231a  and  a86224a );
 a86236a <=( (not A199)  and  (not A168) );
 a86237a <=( A169  and  a86236a );
 a86240a <=( A201  and  A200 );
 a86243a <=( (not A265)  and  A202 );
 a86244a <=( a86243a  and  a86240a );
 a86245a <=( a86244a  and  a86237a );
 a86248a <=( A267  and  A266 );
 a86251a <=( (not A298)  and  (not A269) );
 a86252a <=( a86251a  and  a86248a );
 a86255a <=( (not A300)  and  A299 );
 a86258a <=( A302  and  (not A301) );
 a86259a <=( a86258a  and  a86255a );
 a86260a <=( a86259a  and  a86252a );
 a86264a <=( (not A199)  and  (not A168) );
 a86265a <=( A169  and  a86264a );
 a86268a <=( A201  and  A200 );
 a86271a <=( (not A265)  and  A202 );
 a86272a <=( a86271a  and  a86268a );
 a86273a <=( a86272a  and  a86265a );
 a86276a <=( (not A267)  and  A266 );
 a86279a <=( A269  and  (not A268) );
 a86280a <=( a86279a  and  a86276a );
 a86283a <=( (not A299)  and  A298 );
 a86286a <=( A301  and  A300 );
 a86287a <=( a86286a  and  a86283a );
 a86288a <=( a86287a  and  a86280a );
 a86292a <=( (not A199)  and  (not A168) );
 a86293a <=( A169  and  a86292a );
 a86296a <=( A201  and  A200 );
 a86299a <=( (not A265)  and  A202 );
 a86300a <=( a86299a  and  a86296a );
 a86301a <=( a86300a  and  a86293a );
 a86304a <=( (not A267)  and  A266 );
 a86307a <=( A269  and  (not A268) );
 a86308a <=( a86307a  and  a86304a );
 a86311a <=( (not A299)  and  A298 );
 a86314a <=( (not A302)  and  A300 );
 a86315a <=( a86314a  and  a86311a );
 a86316a <=( a86315a  and  a86308a );
 a86320a <=( (not A199)  and  (not A168) );
 a86321a <=( A169  and  a86320a );
 a86324a <=( A201  and  A200 );
 a86327a <=( (not A265)  and  A202 );
 a86328a <=( a86327a  and  a86324a );
 a86329a <=( a86328a  and  a86321a );
 a86332a <=( (not A267)  and  A266 );
 a86335a <=( A269  and  (not A268) );
 a86336a <=( a86335a  and  a86332a );
 a86339a <=( A299  and  (not A298) );
 a86342a <=( A301  and  A300 );
 a86343a <=( a86342a  and  a86339a );
 a86344a <=( a86343a  and  a86336a );
 a86348a <=( (not A199)  and  (not A168) );
 a86349a <=( A169  and  a86348a );
 a86352a <=( A201  and  A200 );
 a86355a <=( (not A265)  and  A202 );
 a86356a <=( a86355a  and  a86352a );
 a86357a <=( a86356a  and  a86349a );
 a86360a <=( (not A267)  and  A266 );
 a86363a <=( A269  and  (not A268) );
 a86364a <=( a86363a  and  a86360a );
 a86367a <=( A299  and  (not A298) );
 a86370a <=( (not A302)  and  A300 );
 a86371a <=( a86370a  and  a86367a );
 a86372a <=( a86371a  and  a86364a );
 a86376a <=( (not A199)  and  (not A168) );
 a86377a <=( A169  and  a86376a );
 a86380a <=( A201  and  A200 );
 a86383a <=( A265  and  A202 );
 a86384a <=( a86383a  and  a86380a );
 a86385a <=( a86384a  and  a86377a );
 a86388a <=( A267  and  (not A266) );
 a86391a <=( A298  and  A268 );
 a86392a <=( a86391a  and  a86388a );
 a86395a <=( (not A300)  and  (not A299) );
 a86398a <=( A302  and  (not A301) );
 a86399a <=( a86398a  and  a86395a );
 a86400a <=( a86399a  and  a86392a );
 a86404a <=( (not A199)  and  (not A168) );
 a86405a <=( A169  and  a86404a );
 a86408a <=( A201  and  A200 );
 a86411a <=( A265  and  A202 );
 a86412a <=( a86411a  and  a86408a );
 a86413a <=( a86412a  and  a86405a );
 a86416a <=( A267  and  (not A266) );
 a86419a <=( (not A298)  and  A268 );
 a86420a <=( a86419a  and  a86416a );
 a86423a <=( (not A300)  and  A299 );
 a86426a <=( A302  and  (not A301) );
 a86427a <=( a86426a  and  a86423a );
 a86428a <=( a86427a  and  a86420a );
 a86432a <=( (not A199)  and  (not A168) );
 a86433a <=( A169  and  a86432a );
 a86436a <=( A201  and  A200 );
 a86439a <=( A265  and  A202 );
 a86440a <=( a86439a  and  a86436a );
 a86441a <=( a86440a  and  a86433a );
 a86444a <=( A267  and  (not A266) );
 a86447a <=( A298  and  (not A269) );
 a86448a <=( a86447a  and  a86444a );
 a86451a <=( (not A300)  and  (not A299) );
 a86454a <=( A302  and  (not A301) );
 a86455a <=( a86454a  and  a86451a );
 a86456a <=( a86455a  and  a86448a );
 a86460a <=( (not A199)  and  (not A168) );
 a86461a <=( A169  and  a86460a );
 a86464a <=( A201  and  A200 );
 a86467a <=( A265  and  A202 );
 a86468a <=( a86467a  and  a86464a );
 a86469a <=( a86468a  and  a86461a );
 a86472a <=( A267  and  (not A266) );
 a86475a <=( (not A298)  and  (not A269) );
 a86476a <=( a86475a  and  a86472a );
 a86479a <=( (not A300)  and  A299 );
 a86482a <=( A302  and  (not A301) );
 a86483a <=( a86482a  and  a86479a );
 a86484a <=( a86483a  and  a86476a );
 a86488a <=( (not A199)  and  (not A168) );
 a86489a <=( A169  and  a86488a );
 a86492a <=( A201  and  A200 );
 a86495a <=( A265  and  A202 );
 a86496a <=( a86495a  and  a86492a );
 a86497a <=( a86496a  and  a86489a );
 a86500a <=( (not A267)  and  (not A266) );
 a86503a <=( A269  and  (not A268) );
 a86504a <=( a86503a  and  a86500a );
 a86507a <=( (not A299)  and  A298 );
 a86510a <=( A301  and  A300 );
 a86511a <=( a86510a  and  a86507a );
 a86512a <=( a86511a  and  a86504a );
 a86516a <=( (not A199)  and  (not A168) );
 a86517a <=( A169  and  a86516a );
 a86520a <=( A201  and  A200 );
 a86523a <=( A265  and  A202 );
 a86524a <=( a86523a  and  a86520a );
 a86525a <=( a86524a  and  a86517a );
 a86528a <=( (not A267)  and  (not A266) );
 a86531a <=( A269  and  (not A268) );
 a86532a <=( a86531a  and  a86528a );
 a86535a <=( (not A299)  and  A298 );
 a86538a <=( (not A302)  and  A300 );
 a86539a <=( a86538a  and  a86535a );
 a86540a <=( a86539a  and  a86532a );
 a86544a <=( (not A199)  and  (not A168) );
 a86545a <=( A169  and  a86544a );
 a86548a <=( A201  and  A200 );
 a86551a <=( A265  and  A202 );
 a86552a <=( a86551a  and  a86548a );
 a86553a <=( a86552a  and  a86545a );
 a86556a <=( (not A267)  and  (not A266) );
 a86559a <=( A269  and  (not A268) );
 a86560a <=( a86559a  and  a86556a );
 a86563a <=( A299  and  (not A298) );
 a86566a <=( A301  and  A300 );
 a86567a <=( a86566a  and  a86563a );
 a86568a <=( a86567a  and  a86560a );
 a86572a <=( (not A199)  and  (not A168) );
 a86573a <=( A169  and  a86572a );
 a86576a <=( A201  and  A200 );
 a86579a <=( A265  and  A202 );
 a86580a <=( a86579a  and  a86576a );
 a86581a <=( a86580a  and  a86573a );
 a86584a <=( (not A267)  and  (not A266) );
 a86587a <=( A269  and  (not A268) );
 a86588a <=( a86587a  and  a86584a );
 a86591a <=( A299  and  (not A298) );
 a86594a <=( (not A302)  and  A300 );
 a86595a <=( a86594a  and  a86591a );
 a86596a <=( a86595a  and  a86588a );
 a86600a <=( (not A199)  and  (not A168) );
 a86601a <=( A169  and  a86600a );
 a86604a <=( A201  and  A200 );
 a86607a <=( (not A265)  and  (not A203) );
 a86608a <=( a86607a  and  a86604a );
 a86609a <=( a86608a  and  a86601a );
 a86612a <=( A267  and  A266 );
 a86615a <=( A298  and  A268 );
 a86616a <=( a86615a  and  a86612a );
 a86619a <=( (not A300)  and  (not A299) );
 a86622a <=( A302  and  (not A301) );
 a86623a <=( a86622a  and  a86619a );
 a86624a <=( a86623a  and  a86616a );
 a86628a <=( (not A199)  and  (not A168) );
 a86629a <=( A169  and  a86628a );
 a86632a <=( A201  and  A200 );
 a86635a <=( (not A265)  and  (not A203) );
 a86636a <=( a86635a  and  a86632a );
 a86637a <=( a86636a  and  a86629a );
 a86640a <=( A267  and  A266 );
 a86643a <=( (not A298)  and  A268 );
 a86644a <=( a86643a  and  a86640a );
 a86647a <=( (not A300)  and  A299 );
 a86650a <=( A302  and  (not A301) );
 a86651a <=( a86650a  and  a86647a );
 a86652a <=( a86651a  and  a86644a );
 a86656a <=( (not A199)  and  (not A168) );
 a86657a <=( A169  and  a86656a );
 a86660a <=( A201  and  A200 );
 a86663a <=( (not A265)  and  (not A203) );
 a86664a <=( a86663a  and  a86660a );
 a86665a <=( a86664a  and  a86657a );
 a86668a <=( A267  and  A266 );
 a86671a <=( A298  and  (not A269) );
 a86672a <=( a86671a  and  a86668a );
 a86675a <=( (not A300)  and  (not A299) );
 a86678a <=( A302  and  (not A301) );
 a86679a <=( a86678a  and  a86675a );
 a86680a <=( a86679a  and  a86672a );
 a86684a <=( (not A199)  and  (not A168) );
 a86685a <=( A169  and  a86684a );
 a86688a <=( A201  and  A200 );
 a86691a <=( (not A265)  and  (not A203) );
 a86692a <=( a86691a  and  a86688a );
 a86693a <=( a86692a  and  a86685a );
 a86696a <=( A267  and  A266 );
 a86699a <=( (not A298)  and  (not A269) );
 a86700a <=( a86699a  and  a86696a );
 a86703a <=( (not A300)  and  A299 );
 a86706a <=( A302  and  (not A301) );
 a86707a <=( a86706a  and  a86703a );
 a86708a <=( a86707a  and  a86700a );
 a86712a <=( (not A199)  and  (not A168) );
 a86713a <=( A169  and  a86712a );
 a86716a <=( A201  and  A200 );
 a86719a <=( (not A265)  and  (not A203) );
 a86720a <=( a86719a  and  a86716a );
 a86721a <=( a86720a  and  a86713a );
 a86724a <=( (not A267)  and  A266 );
 a86727a <=( A269  and  (not A268) );
 a86728a <=( a86727a  and  a86724a );
 a86731a <=( (not A299)  and  A298 );
 a86734a <=( A301  and  A300 );
 a86735a <=( a86734a  and  a86731a );
 a86736a <=( a86735a  and  a86728a );
 a86740a <=( (not A199)  and  (not A168) );
 a86741a <=( A169  and  a86740a );
 a86744a <=( A201  and  A200 );
 a86747a <=( (not A265)  and  (not A203) );
 a86748a <=( a86747a  and  a86744a );
 a86749a <=( a86748a  and  a86741a );
 a86752a <=( (not A267)  and  A266 );
 a86755a <=( A269  and  (not A268) );
 a86756a <=( a86755a  and  a86752a );
 a86759a <=( (not A299)  and  A298 );
 a86762a <=( (not A302)  and  A300 );
 a86763a <=( a86762a  and  a86759a );
 a86764a <=( a86763a  and  a86756a );
 a86768a <=( (not A199)  and  (not A168) );
 a86769a <=( A169  and  a86768a );
 a86772a <=( A201  and  A200 );
 a86775a <=( (not A265)  and  (not A203) );
 a86776a <=( a86775a  and  a86772a );
 a86777a <=( a86776a  and  a86769a );
 a86780a <=( (not A267)  and  A266 );
 a86783a <=( A269  and  (not A268) );
 a86784a <=( a86783a  and  a86780a );
 a86787a <=( A299  and  (not A298) );
 a86790a <=( A301  and  A300 );
 a86791a <=( a86790a  and  a86787a );
 a86792a <=( a86791a  and  a86784a );
 a86796a <=( (not A199)  and  (not A168) );
 a86797a <=( A169  and  a86796a );
 a86800a <=( A201  and  A200 );
 a86803a <=( (not A265)  and  (not A203) );
 a86804a <=( a86803a  and  a86800a );
 a86805a <=( a86804a  and  a86797a );
 a86808a <=( (not A267)  and  A266 );
 a86811a <=( A269  and  (not A268) );
 a86812a <=( a86811a  and  a86808a );
 a86815a <=( A299  and  (not A298) );
 a86818a <=( (not A302)  and  A300 );
 a86819a <=( a86818a  and  a86815a );
 a86820a <=( a86819a  and  a86812a );
 a86824a <=( (not A199)  and  (not A168) );
 a86825a <=( A169  and  a86824a );
 a86828a <=( A201  and  A200 );
 a86831a <=( A265  and  (not A203) );
 a86832a <=( a86831a  and  a86828a );
 a86833a <=( a86832a  and  a86825a );
 a86836a <=( A267  and  (not A266) );
 a86839a <=( A298  and  A268 );
 a86840a <=( a86839a  and  a86836a );
 a86843a <=( (not A300)  and  (not A299) );
 a86846a <=( A302  and  (not A301) );
 a86847a <=( a86846a  and  a86843a );
 a86848a <=( a86847a  and  a86840a );
 a86852a <=( (not A199)  and  (not A168) );
 a86853a <=( A169  and  a86852a );
 a86856a <=( A201  and  A200 );
 a86859a <=( A265  and  (not A203) );
 a86860a <=( a86859a  and  a86856a );
 a86861a <=( a86860a  and  a86853a );
 a86864a <=( A267  and  (not A266) );
 a86867a <=( (not A298)  and  A268 );
 a86868a <=( a86867a  and  a86864a );
 a86871a <=( (not A300)  and  A299 );
 a86874a <=( A302  and  (not A301) );
 a86875a <=( a86874a  and  a86871a );
 a86876a <=( a86875a  and  a86868a );
 a86880a <=( (not A199)  and  (not A168) );
 a86881a <=( A169  and  a86880a );
 a86884a <=( A201  and  A200 );
 a86887a <=( A265  and  (not A203) );
 a86888a <=( a86887a  and  a86884a );
 a86889a <=( a86888a  and  a86881a );
 a86892a <=( A267  and  (not A266) );
 a86895a <=( A298  and  (not A269) );
 a86896a <=( a86895a  and  a86892a );
 a86899a <=( (not A300)  and  (not A299) );
 a86902a <=( A302  and  (not A301) );
 a86903a <=( a86902a  and  a86899a );
 a86904a <=( a86903a  and  a86896a );
 a86908a <=( (not A199)  and  (not A168) );
 a86909a <=( A169  and  a86908a );
 a86912a <=( A201  and  A200 );
 a86915a <=( A265  and  (not A203) );
 a86916a <=( a86915a  and  a86912a );
 a86917a <=( a86916a  and  a86909a );
 a86920a <=( A267  and  (not A266) );
 a86923a <=( (not A298)  and  (not A269) );
 a86924a <=( a86923a  and  a86920a );
 a86927a <=( (not A300)  and  A299 );
 a86930a <=( A302  and  (not A301) );
 a86931a <=( a86930a  and  a86927a );
 a86932a <=( a86931a  and  a86924a );
 a86936a <=( (not A199)  and  (not A168) );
 a86937a <=( A169  and  a86936a );
 a86940a <=( A201  and  A200 );
 a86943a <=( A265  and  (not A203) );
 a86944a <=( a86943a  and  a86940a );
 a86945a <=( a86944a  and  a86937a );
 a86948a <=( (not A267)  and  (not A266) );
 a86951a <=( A269  and  (not A268) );
 a86952a <=( a86951a  and  a86948a );
 a86955a <=( (not A299)  and  A298 );
 a86958a <=( A301  and  A300 );
 a86959a <=( a86958a  and  a86955a );
 a86960a <=( a86959a  and  a86952a );
 a86964a <=( (not A199)  and  (not A168) );
 a86965a <=( A169  and  a86964a );
 a86968a <=( A201  and  A200 );
 a86971a <=( A265  and  (not A203) );
 a86972a <=( a86971a  and  a86968a );
 a86973a <=( a86972a  and  a86965a );
 a86976a <=( (not A267)  and  (not A266) );
 a86979a <=( A269  and  (not A268) );
 a86980a <=( a86979a  and  a86976a );
 a86983a <=( (not A299)  and  A298 );
 a86986a <=( (not A302)  and  A300 );
 a86987a <=( a86986a  and  a86983a );
 a86988a <=( a86987a  and  a86980a );
 a86992a <=( (not A199)  and  (not A168) );
 a86993a <=( A169  and  a86992a );
 a86996a <=( A201  and  A200 );
 a86999a <=( A265  and  (not A203) );
 a87000a <=( a86999a  and  a86996a );
 a87001a <=( a87000a  and  a86993a );
 a87004a <=( (not A267)  and  (not A266) );
 a87007a <=( A269  and  (not A268) );
 a87008a <=( a87007a  and  a87004a );
 a87011a <=( A299  and  (not A298) );
 a87014a <=( A301  and  A300 );
 a87015a <=( a87014a  and  a87011a );
 a87016a <=( a87015a  and  a87008a );
 a87020a <=( (not A199)  and  (not A168) );
 a87021a <=( A169  and  a87020a );
 a87024a <=( A201  and  A200 );
 a87027a <=( A265  and  (not A203) );
 a87028a <=( a87027a  and  a87024a );
 a87029a <=( a87028a  and  a87021a );
 a87032a <=( (not A267)  and  (not A266) );
 a87035a <=( A269  and  (not A268) );
 a87036a <=( a87035a  and  a87032a );
 a87039a <=( A299  and  (not A298) );
 a87042a <=( (not A302)  and  A300 );
 a87043a <=( a87042a  and  a87039a );
 a87044a <=( a87043a  and  a87036a );
 a87048a <=( (not A199)  and  (not A168) );
 a87049a <=( A169  and  a87048a );
 a87052a <=( (not A201)  and  A200 );
 a87055a <=( A203  and  (not A202) );
 a87056a <=( a87055a  and  a87052a );
 a87057a <=( a87056a  and  a87049a );
 a87060a <=( A266  and  (not A265) );
 a87063a <=( A268  and  A267 );
 a87064a <=( a87063a  and  a87060a );
 a87067a <=( (not A299)  and  A298 );
 a87070a <=( A301  and  A300 );
 a87071a <=( a87070a  and  a87067a );
 a87072a <=( a87071a  and  a87064a );
 a87076a <=( (not A199)  and  (not A168) );
 a87077a <=( A169  and  a87076a );
 a87080a <=( (not A201)  and  A200 );
 a87083a <=( A203  and  (not A202) );
 a87084a <=( a87083a  and  a87080a );
 a87085a <=( a87084a  and  a87077a );
 a87088a <=( A266  and  (not A265) );
 a87091a <=( A268  and  A267 );
 a87092a <=( a87091a  and  a87088a );
 a87095a <=( (not A299)  and  A298 );
 a87098a <=( (not A302)  and  A300 );
 a87099a <=( a87098a  and  a87095a );
 a87100a <=( a87099a  and  a87092a );
 a87104a <=( (not A199)  and  (not A168) );
 a87105a <=( A169  and  a87104a );
 a87108a <=( (not A201)  and  A200 );
 a87111a <=( A203  and  (not A202) );
 a87112a <=( a87111a  and  a87108a );
 a87113a <=( a87112a  and  a87105a );
 a87116a <=( A266  and  (not A265) );
 a87119a <=( A268  and  A267 );
 a87120a <=( a87119a  and  a87116a );
 a87123a <=( A299  and  (not A298) );
 a87126a <=( A301  and  A300 );
 a87127a <=( a87126a  and  a87123a );
 a87128a <=( a87127a  and  a87120a );
 a87132a <=( (not A199)  and  (not A168) );
 a87133a <=( A169  and  a87132a );
 a87136a <=( (not A201)  and  A200 );
 a87139a <=( A203  and  (not A202) );
 a87140a <=( a87139a  and  a87136a );
 a87141a <=( a87140a  and  a87133a );
 a87144a <=( A266  and  (not A265) );
 a87147a <=( A268  and  A267 );
 a87148a <=( a87147a  and  a87144a );
 a87151a <=( A299  and  (not A298) );
 a87154a <=( (not A302)  and  A300 );
 a87155a <=( a87154a  and  a87151a );
 a87156a <=( a87155a  and  a87148a );
 a87160a <=( (not A199)  and  (not A168) );
 a87161a <=( A169  and  a87160a );
 a87164a <=( (not A201)  and  A200 );
 a87167a <=( A203  and  (not A202) );
 a87168a <=( a87167a  and  a87164a );
 a87169a <=( a87168a  and  a87161a );
 a87172a <=( A266  and  (not A265) );
 a87175a <=( (not A269)  and  A267 );
 a87176a <=( a87175a  and  a87172a );
 a87179a <=( (not A299)  and  A298 );
 a87182a <=( A301  and  A300 );
 a87183a <=( a87182a  and  a87179a );
 a87184a <=( a87183a  and  a87176a );
 a87188a <=( (not A199)  and  (not A168) );
 a87189a <=( A169  and  a87188a );
 a87192a <=( (not A201)  and  A200 );
 a87195a <=( A203  and  (not A202) );
 a87196a <=( a87195a  and  a87192a );
 a87197a <=( a87196a  and  a87189a );
 a87200a <=( A266  and  (not A265) );
 a87203a <=( (not A269)  and  A267 );
 a87204a <=( a87203a  and  a87200a );
 a87207a <=( (not A299)  and  A298 );
 a87210a <=( (not A302)  and  A300 );
 a87211a <=( a87210a  and  a87207a );
 a87212a <=( a87211a  and  a87204a );
 a87216a <=( (not A199)  and  (not A168) );
 a87217a <=( A169  and  a87216a );
 a87220a <=( (not A201)  and  A200 );
 a87223a <=( A203  and  (not A202) );
 a87224a <=( a87223a  and  a87220a );
 a87225a <=( a87224a  and  a87217a );
 a87228a <=( A266  and  (not A265) );
 a87231a <=( (not A269)  and  A267 );
 a87232a <=( a87231a  and  a87228a );
 a87235a <=( A299  and  (not A298) );
 a87238a <=( A301  and  A300 );
 a87239a <=( a87238a  and  a87235a );
 a87240a <=( a87239a  and  a87232a );
 a87244a <=( (not A199)  and  (not A168) );
 a87245a <=( A169  and  a87244a );
 a87248a <=( (not A201)  and  A200 );
 a87251a <=( A203  and  (not A202) );
 a87252a <=( a87251a  and  a87248a );
 a87253a <=( a87252a  and  a87245a );
 a87256a <=( A266  and  (not A265) );
 a87259a <=( (not A269)  and  A267 );
 a87260a <=( a87259a  and  a87256a );
 a87263a <=( A299  and  (not A298) );
 a87266a <=( (not A302)  and  A300 );
 a87267a <=( a87266a  and  a87263a );
 a87268a <=( a87267a  and  a87260a );
 a87272a <=( (not A199)  and  (not A168) );
 a87273a <=( A169  and  a87272a );
 a87276a <=( (not A201)  and  A200 );
 a87279a <=( A203  and  (not A202) );
 a87280a <=( a87279a  and  a87276a );
 a87281a <=( a87280a  and  a87273a );
 a87284a <=( (not A266)  and  A265 );
 a87287a <=( A268  and  A267 );
 a87288a <=( a87287a  and  a87284a );
 a87291a <=( (not A299)  and  A298 );
 a87294a <=( A301  and  A300 );
 a87295a <=( a87294a  and  a87291a );
 a87296a <=( a87295a  and  a87288a );
 a87300a <=( (not A199)  and  (not A168) );
 a87301a <=( A169  and  a87300a );
 a87304a <=( (not A201)  and  A200 );
 a87307a <=( A203  and  (not A202) );
 a87308a <=( a87307a  and  a87304a );
 a87309a <=( a87308a  and  a87301a );
 a87312a <=( (not A266)  and  A265 );
 a87315a <=( A268  and  A267 );
 a87316a <=( a87315a  and  a87312a );
 a87319a <=( (not A299)  and  A298 );
 a87322a <=( (not A302)  and  A300 );
 a87323a <=( a87322a  and  a87319a );
 a87324a <=( a87323a  and  a87316a );
 a87328a <=( (not A199)  and  (not A168) );
 a87329a <=( A169  and  a87328a );
 a87332a <=( (not A201)  and  A200 );
 a87335a <=( A203  and  (not A202) );
 a87336a <=( a87335a  and  a87332a );
 a87337a <=( a87336a  and  a87329a );
 a87340a <=( (not A266)  and  A265 );
 a87343a <=( A268  and  A267 );
 a87344a <=( a87343a  and  a87340a );
 a87347a <=( A299  and  (not A298) );
 a87350a <=( A301  and  A300 );
 a87351a <=( a87350a  and  a87347a );
 a87352a <=( a87351a  and  a87344a );
 a87356a <=( (not A199)  and  (not A168) );
 a87357a <=( A169  and  a87356a );
 a87360a <=( (not A201)  and  A200 );
 a87363a <=( A203  and  (not A202) );
 a87364a <=( a87363a  and  a87360a );
 a87365a <=( a87364a  and  a87357a );
 a87368a <=( (not A266)  and  A265 );
 a87371a <=( A268  and  A267 );
 a87372a <=( a87371a  and  a87368a );
 a87375a <=( A299  and  (not A298) );
 a87378a <=( (not A302)  and  A300 );
 a87379a <=( a87378a  and  a87375a );
 a87380a <=( a87379a  and  a87372a );
 a87384a <=( (not A199)  and  (not A168) );
 a87385a <=( A169  and  a87384a );
 a87388a <=( (not A201)  and  A200 );
 a87391a <=( A203  and  (not A202) );
 a87392a <=( a87391a  and  a87388a );
 a87393a <=( a87392a  and  a87385a );
 a87396a <=( (not A266)  and  A265 );
 a87399a <=( (not A269)  and  A267 );
 a87400a <=( a87399a  and  a87396a );
 a87403a <=( (not A299)  and  A298 );
 a87406a <=( A301  and  A300 );
 a87407a <=( a87406a  and  a87403a );
 a87408a <=( a87407a  and  a87400a );
 a87412a <=( (not A199)  and  (not A168) );
 a87413a <=( A169  and  a87412a );
 a87416a <=( (not A201)  and  A200 );
 a87419a <=( A203  and  (not A202) );
 a87420a <=( a87419a  and  a87416a );
 a87421a <=( a87420a  and  a87413a );
 a87424a <=( (not A266)  and  A265 );
 a87427a <=( (not A269)  and  A267 );
 a87428a <=( a87427a  and  a87424a );
 a87431a <=( (not A299)  and  A298 );
 a87434a <=( (not A302)  and  A300 );
 a87435a <=( a87434a  and  a87431a );
 a87436a <=( a87435a  and  a87428a );
 a87440a <=( (not A199)  and  (not A168) );
 a87441a <=( A169  and  a87440a );
 a87444a <=( (not A201)  and  A200 );
 a87447a <=( A203  and  (not A202) );
 a87448a <=( a87447a  and  a87444a );
 a87449a <=( a87448a  and  a87441a );
 a87452a <=( (not A266)  and  A265 );
 a87455a <=( (not A269)  and  A267 );
 a87456a <=( a87455a  and  a87452a );
 a87459a <=( A299  and  (not A298) );
 a87462a <=( A301  and  A300 );
 a87463a <=( a87462a  and  a87459a );
 a87464a <=( a87463a  and  a87456a );
 a87468a <=( (not A199)  and  (not A168) );
 a87469a <=( A169  and  a87468a );
 a87472a <=( (not A201)  and  A200 );
 a87475a <=( A203  and  (not A202) );
 a87476a <=( a87475a  and  a87472a );
 a87477a <=( a87476a  and  a87469a );
 a87480a <=( (not A266)  and  A265 );
 a87483a <=( (not A269)  and  A267 );
 a87484a <=( a87483a  and  a87480a );
 a87487a <=( A299  and  (not A298) );
 a87490a <=( (not A302)  and  A300 );
 a87491a <=( a87490a  and  a87487a );
 a87492a <=( a87491a  and  a87484a );
 a87496a <=( A199  and  (not A168) );
 a87497a <=( A169  and  a87496a );
 a87500a <=( A201  and  (not A200) );
 a87503a <=( (not A265)  and  A202 );
 a87504a <=( a87503a  and  a87500a );
 a87505a <=( a87504a  and  a87497a );
 a87508a <=( A267  and  A266 );
 a87511a <=( A298  and  A268 );
 a87512a <=( a87511a  and  a87508a );
 a87515a <=( (not A300)  and  (not A299) );
 a87518a <=( A302  and  (not A301) );
 a87519a <=( a87518a  and  a87515a );
 a87520a <=( a87519a  and  a87512a );
 a87524a <=( A199  and  (not A168) );
 a87525a <=( A169  and  a87524a );
 a87528a <=( A201  and  (not A200) );
 a87531a <=( (not A265)  and  A202 );
 a87532a <=( a87531a  and  a87528a );
 a87533a <=( a87532a  and  a87525a );
 a87536a <=( A267  and  A266 );
 a87539a <=( (not A298)  and  A268 );
 a87540a <=( a87539a  and  a87536a );
 a87543a <=( (not A300)  and  A299 );
 a87546a <=( A302  and  (not A301) );
 a87547a <=( a87546a  and  a87543a );
 a87548a <=( a87547a  and  a87540a );
 a87552a <=( A199  and  (not A168) );
 a87553a <=( A169  and  a87552a );
 a87556a <=( A201  and  (not A200) );
 a87559a <=( (not A265)  and  A202 );
 a87560a <=( a87559a  and  a87556a );
 a87561a <=( a87560a  and  a87553a );
 a87564a <=( A267  and  A266 );
 a87567a <=( A298  and  (not A269) );
 a87568a <=( a87567a  and  a87564a );
 a87571a <=( (not A300)  and  (not A299) );
 a87574a <=( A302  and  (not A301) );
 a87575a <=( a87574a  and  a87571a );
 a87576a <=( a87575a  and  a87568a );
 a87580a <=( A199  and  (not A168) );
 a87581a <=( A169  and  a87580a );
 a87584a <=( A201  and  (not A200) );
 a87587a <=( (not A265)  and  A202 );
 a87588a <=( a87587a  and  a87584a );
 a87589a <=( a87588a  and  a87581a );
 a87592a <=( A267  and  A266 );
 a87595a <=( (not A298)  and  (not A269) );
 a87596a <=( a87595a  and  a87592a );
 a87599a <=( (not A300)  and  A299 );
 a87602a <=( A302  and  (not A301) );
 a87603a <=( a87602a  and  a87599a );
 a87604a <=( a87603a  and  a87596a );
 a87608a <=( A199  and  (not A168) );
 a87609a <=( A169  and  a87608a );
 a87612a <=( A201  and  (not A200) );
 a87615a <=( (not A265)  and  A202 );
 a87616a <=( a87615a  and  a87612a );
 a87617a <=( a87616a  and  a87609a );
 a87620a <=( (not A267)  and  A266 );
 a87623a <=( A269  and  (not A268) );
 a87624a <=( a87623a  and  a87620a );
 a87627a <=( (not A299)  and  A298 );
 a87630a <=( A301  and  A300 );
 a87631a <=( a87630a  and  a87627a );
 a87632a <=( a87631a  and  a87624a );
 a87636a <=( A199  and  (not A168) );
 a87637a <=( A169  and  a87636a );
 a87640a <=( A201  and  (not A200) );
 a87643a <=( (not A265)  and  A202 );
 a87644a <=( a87643a  and  a87640a );
 a87645a <=( a87644a  and  a87637a );
 a87648a <=( (not A267)  and  A266 );
 a87651a <=( A269  and  (not A268) );
 a87652a <=( a87651a  and  a87648a );
 a87655a <=( (not A299)  and  A298 );
 a87658a <=( (not A302)  and  A300 );
 a87659a <=( a87658a  and  a87655a );
 a87660a <=( a87659a  and  a87652a );
 a87664a <=( A199  and  (not A168) );
 a87665a <=( A169  and  a87664a );
 a87668a <=( A201  and  (not A200) );
 a87671a <=( (not A265)  and  A202 );
 a87672a <=( a87671a  and  a87668a );
 a87673a <=( a87672a  and  a87665a );
 a87676a <=( (not A267)  and  A266 );
 a87679a <=( A269  and  (not A268) );
 a87680a <=( a87679a  and  a87676a );
 a87683a <=( A299  and  (not A298) );
 a87686a <=( A301  and  A300 );
 a87687a <=( a87686a  and  a87683a );
 a87688a <=( a87687a  and  a87680a );
 a87692a <=( A199  and  (not A168) );
 a87693a <=( A169  and  a87692a );
 a87696a <=( A201  and  (not A200) );
 a87699a <=( (not A265)  and  A202 );
 a87700a <=( a87699a  and  a87696a );
 a87701a <=( a87700a  and  a87693a );
 a87704a <=( (not A267)  and  A266 );
 a87707a <=( A269  and  (not A268) );
 a87708a <=( a87707a  and  a87704a );
 a87711a <=( A299  and  (not A298) );
 a87714a <=( (not A302)  and  A300 );
 a87715a <=( a87714a  and  a87711a );
 a87716a <=( a87715a  and  a87708a );
 a87720a <=( A199  and  (not A168) );
 a87721a <=( A169  and  a87720a );
 a87724a <=( A201  and  (not A200) );
 a87727a <=( A265  and  A202 );
 a87728a <=( a87727a  and  a87724a );
 a87729a <=( a87728a  and  a87721a );
 a87732a <=( A267  and  (not A266) );
 a87735a <=( A298  and  A268 );
 a87736a <=( a87735a  and  a87732a );
 a87739a <=( (not A300)  and  (not A299) );
 a87742a <=( A302  and  (not A301) );
 a87743a <=( a87742a  and  a87739a );
 a87744a <=( a87743a  and  a87736a );
 a87748a <=( A199  and  (not A168) );
 a87749a <=( A169  and  a87748a );
 a87752a <=( A201  and  (not A200) );
 a87755a <=( A265  and  A202 );
 a87756a <=( a87755a  and  a87752a );
 a87757a <=( a87756a  and  a87749a );
 a87760a <=( A267  and  (not A266) );
 a87763a <=( (not A298)  and  A268 );
 a87764a <=( a87763a  and  a87760a );
 a87767a <=( (not A300)  and  A299 );
 a87770a <=( A302  and  (not A301) );
 a87771a <=( a87770a  and  a87767a );
 a87772a <=( a87771a  and  a87764a );
 a87776a <=( A199  and  (not A168) );
 a87777a <=( A169  and  a87776a );
 a87780a <=( A201  and  (not A200) );
 a87783a <=( A265  and  A202 );
 a87784a <=( a87783a  and  a87780a );
 a87785a <=( a87784a  and  a87777a );
 a87788a <=( A267  and  (not A266) );
 a87791a <=( A298  and  (not A269) );
 a87792a <=( a87791a  and  a87788a );
 a87795a <=( (not A300)  and  (not A299) );
 a87798a <=( A302  and  (not A301) );
 a87799a <=( a87798a  and  a87795a );
 a87800a <=( a87799a  and  a87792a );
 a87804a <=( A199  and  (not A168) );
 a87805a <=( A169  and  a87804a );
 a87808a <=( A201  and  (not A200) );
 a87811a <=( A265  and  A202 );
 a87812a <=( a87811a  and  a87808a );
 a87813a <=( a87812a  and  a87805a );
 a87816a <=( A267  and  (not A266) );
 a87819a <=( (not A298)  and  (not A269) );
 a87820a <=( a87819a  and  a87816a );
 a87823a <=( (not A300)  and  A299 );
 a87826a <=( A302  and  (not A301) );
 a87827a <=( a87826a  and  a87823a );
 a87828a <=( a87827a  and  a87820a );
 a87832a <=( A199  and  (not A168) );
 a87833a <=( A169  and  a87832a );
 a87836a <=( A201  and  (not A200) );
 a87839a <=( A265  and  A202 );
 a87840a <=( a87839a  and  a87836a );
 a87841a <=( a87840a  and  a87833a );
 a87844a <=( (not A267)  and  (not A266) );
 a87847a <=( A269  and  (not A268) );
 a87848a <=( a87847a  and  a87844a );
 a87851a <=( (not A299)  and  A298 );
 a87854a <=( A301  and  A300 );
 a87855a <=( a87854a  and  a87851a );
 a87856a <=( a87855a  and  a87848a );
 a87860a <=( A199  and  (not A168) );
 a87861a <=( A169  and  a87860a );
 a87864a <=( A201  and  (not A200) );
 a87867a <=( A265  and  A202 );
 a87868a <=( a87867a  and  a87864a );
 a87869a <=( a87868a  and  a87861a );
 a87872a <=( (not A267)  and  (not A266) );
 a87875a <=( A269  and  (not A268) );
 a87876a <=( a87875a  and  a87872a );
 a87879a <=( (not A299)  and  A298 );
 a87882a <=( (not A302)  and  A300 );
 a87883a <=( a87882a  and  a87879a );
 a87884a <=( a87883a  and  a87876a );
 a87888a <=( A199  and  (not A168) );
 a87889a <=( A169  and  a87888a );
 a87892a <=( A201  and  (not A200) );
 a87895a <=( A265  and  A202 );
 a87896a <=( a87895a  and  a87892a );
 a87897a <=( a87896a  and  a87889a );
 a87900a <=( (not A267)  and  (not A266) );
 a87903a <=( A269  and  (not A268) );
 a87904a <=( a87903a  and  a87900a );
 a87907a <=( A299  and  (not A298) );
 a87910a <=( A301  and  A300 );
 a87911a <=( a87910a  and  a87907a );
 a87912a <=( a87911a  and  a87904a );
 a87916a <=( A199  and  (not A168) );
 a87917a <=( A169  and  a87916a );
 a87920a <=( A201  and  (not A200) );
 a87923a <=( A265  and  A202 );
 a87924a <=( a87923a  and  a87920a );
 a87925a <=( a87924a  and  a87917a );
 a87928a <=( (not A267)  and  (not A266) );
 a87931a <=( A269  and  (not A268) );
 a87932a <=( a87931a  and  a87928a );
 a87935a <=( A299  and  (not A298) );
 a87938a <=( (not A302)  and  A300 );
 a87939a <=( a87938a  and  a87935a );
 a87940a <=( a87939a  and  a87932a );
 a87944a <=( A199  and  (not A168) );
 a87945a <=( A169  and  a87944a );
 a87948a <=( A201  and  (not A200) );
 a87951a <=( (not A265)  and  (not A203) );
 a87952a <=( a87951a  and  a87948a );
 a87953a <=( a87952a  and  a87945a );
 a87956a <=( A267  and  A266 );
 a87959a <=( A298  and  A268 );
 a87960a <=( a87959a  and  a87956a );
 a87963a <=( (not A300)  and  (not A299) );
 a87966a <=( A302  and  (not A301) );
 a87967a <=( a87966a  and  a87963a );
 a87968a <=( a87967a  and  a87960a );
 a87972a <=( A199  and  (not A168) );
 a87973a <=( A169  and  a87972a );
 a87976a <=( A201  and  (not A200) );
 a87979a <=( (not A265)  and  (not A203) );
 a87980a <=( a87979a  and  a87976a );
 a87981a <=( a87980a  and  a87973a );
 a87984a <=( A267  and  A266 );
 a87987a <=( (not A298)  and  A268 );
 a87988a <=( a87987a  and  a87984a );
 a87991a <=( (not A300)  and  A299 );
 a87994a <=( A302  and  (not A301) );
 a87995a <=( a87994a  and  a87991a );
 a87996a <=( a87995a  and  a87988a );
 a88000a <=( A199  and  (not A168) );
 a88001a <=( A169  and  a88000a );
 a88004a <=( A201  and  (not A200) );
 a88007a <=( (not A265)  and  (not A203) );
 a88008a <=( a88007a  and  a88004a );
 a88009a <=( a88008a  and  a88001a );
 a88012a <=( A267  and  A266 );
 a88015a <=( A298  and  (not A269) );
 a88016a <=( a88015a  and  a88012a );
 a88019a <=( (not A300)  and  (not A299) );
 a88022a <=( A302  and  (not A301) );
 a88023a <=( a88022a  and  a88019a );
 a88024a <=( a88023a  and  a88016a );
 a88028a <=( A199  and  (not A168) );
 a88029a <=( A169  and  a88028a );
 a88032a <=( A201  and  (not A200) );
 a88035a <=( (not A265)  and  (not A203) );
 a88036a <=( a88035a  and  a88032a );
 a88037a <=( a88036a  and  a88029a );
 a88040a <=( A267  and  A266 );
 a88043a <=( (not A298)  and  (not A269) );
 a88044a <=( a88043a  and  a88040a );
 a88047a <=( (not A300)  and  A299 );
 a88050a <=( A302  and  (not A301) );
 a88051a <=( a88050a  and  a88047a );
 a88052a <=( a88051a  and  a88044a );
 a88056a <=( A199  and  (not A168) );
 a88057a <=( A169  and  a88056a );
 a88060a <=( A201  and  (not A200) );
 a88063a <=( (not A265)  and  (not A203) );
 a88064a <=( a88063a  and  a88060a );
 a88065a <=( a88064a  and  a88057a );
 a88068a <=( (not A267)  and  A266 );
 a88071a <=( A269  and  (not A268) );
 a88072a <=( a88071a  and  a88068a );
 a88075a <=( (not A299)  and  A298 );
 a88078a <=( A301  and  A300 );
 a88079a <=( a88078a  and  a88075a );
 a88080a <=( a88079a  and  a88072a );
 a88084a <=( A199  and  (not A168) );
 a88085a <=( A169  and  a88084a );
 a88088a <=( A201  and  (not A200) );
 a88091a <=( (not A265)  and  (not A203) );
 a88092a <=( a88091a  and  a88088a );
 a88093a <=( a88092a  and  a88085a );
 a88096a <=( (not A267)  and  A266 );
 a88099a <=( A269  and  (not A268) );
 a88100a <=( a88099a  and  a88096a );
 a88103a <=( (not A299)  and  A298 );
 a88106a <=( (not A302)  and  A300 );
 a88107a <=( a88106a  and  a88103a );
 a88108a <=( a88107a  and  a88100a );
 a88112a <=( A199  and  (not A168) );
 a88113a <=( A169  and  a88112a );
 a88116a <=( A201  and  (not A200) );
 a88119a <=( (not A265)  and  (not A203) );
 a88120a <=( a88119a  and  a88116a );
 a88121a <=( a88120a  and  a88113a );
 a88124a <=( (not A267)  and  A266 );
 a88127a <=( A269  and  (not A268) );
 a88128a <=( a88127a  and  a88124a );
 a88131a <=( A299  and  (not A298) );
 a88134a <=( A301  and  A300 );
 a88135a <=( a88134a  and  a88131a );
 a88136a <=( a88135a  and  a88128a );
 a88140a <=( A199  and  (not A168) );
 a88141a <=( A169  and  a88140a );
 a88144a <=( A201  and  (not A200) );
 a88147a <=( (not A265)  and  (not A203) );
 a88148a <=( a88147a  and  a88144a );
 a88149a <=( a88148a  and  a88141a );
 a88152a <=( (not A267)  and  A266 );
 a88155a <=( A269  and  (not A268) );
 a88156a <=( a88155a  and  a88152a );
 a88159a <=( A299  and  (not A298) );
 a88162a <=( (not A302)  and  A300 );
 a88163a <=( a88162a  and  a88159a );
 a88164a <=( a88163a  and  a88156a );
 a88168a <=( A199  and  (not A168) );
 a88169a <=( A169  and  a88168a );
 a88172a <=( A201  and  (not A200) );
 a88175a <=( A265  and  (not A203) );
 a88176a <=( a88175a  and  a88172a );
 a88177a <=( a88176a  and  a88169a );
 a88180a <=( A267  and  (not A266) );
 a88183a <=( A298  and  A268 );
 a88184a <=( a88183a  and  a88180a );
 a88187a <=( (not A300)  and  (not A299) );
 a88190a <=( A302  and  (not A301) );
 a88191a <=( a88190a  and  a88187a );
 a88192a <=( a88191a  and  a88184a );
 a88196a <=( A199  and  (not A168) );
 a88197a <=( A169  and  a88196a );
 a88200a <=( A201  and  (not A200) );
 a88203a <=( A265  and  (not A203) );
 a88204a <=( a88203a  and  a88200a );
 a88205a <=( a88204a  and  a88197a );
 a88208a <=( A267  and  (not A266) );
 a88211a <=( (not A298)  and  A268 );
 a88212a <=( a88211a  and  a88208a );
 a88215a <=( (not A300)  and  A299 );
 a88218a <=( A302  and  (not A301) );
 a88219a <=( a88218a  and  a88215a );
 a88220a <=( a88219a  and  a88212a );
 a88224a <=( A199  and  (not A168) );
 a88225a <=( A169  and  a88224a );
 a88228a <=( A201  and  (not A200) );
 a88231a <=( A265  and  (not A203) );
 a88232a <=( a88231a  and  a88228a );
 a88233a <=( a88232a  and  a88225a );
 a88236a <=( A267  and  (not A266) );
 a88239a <=( A298  and  (not A269) );
 a88240a <=( a88239a  and  a88236a );
 a88243a <=( (not A300)  and  (not A299) );
 a88246a <=( A302  and  (not A301) );
 a88247a <=( a88246a  and  a88243a );
 a88248a <=( a88247a  and  a88240a );
 a88252a <=( A199  and  (not A168) );
 a88253a <=( A169  and  a88252a );
 a88256a <=( A201  and  (not A200) );
 a88259a <=( A265  and  (not A203) );
 a88260a <=( a88259a  and  a88256a );
 a88261a <=( a88260a  and  a88253a );
 a88264a <=( A267  and  (not A266) );
 a88267a <=( (not A298)  and  (not A269) );
 a88268a <=( a88267a  and  a88264a );
 a88271a <=( (not A300)  and  A299 );
 a88274a <=( A302  and  (not A301) );
 a88275a <=( a88274a  and  a88271a );
 a88276a <=( a88275a  and  a88268a );
 a88280a <=( A199  and  (not A168) );
 a88281a <=( A169  and  a88280a );
 a88284a <=( A201  and  (not A200) );
 a88287a <=( A265  and  (not A203) );
 a88288a <=( a88287a  and  a88284a );
 a88289a <=( a88288a  and  a88281a );
 a88292a <=( (not A267)  and  (not A266) );
 a88295a <=( A269  and  (not A268) );
 a88296a <=( a88295a  and  a88292a );
 a88299a <=( (not A299)  and  A298 );
 a88302a <=( A301  and  A300 );
 a88303a <=( a88302a  and  a88299a );
 a88304a <=( a88303a  and  a88296a );
 a88308a <=( A199  and  (not A168) );
 a88309a <=( A169  and  a88308a );
 a88312a <=( A201  and  (not A200) );
 a88315a <=( A265  and  (not A203) );
 a88316a <=( a88315a  and  a88312a );
 a88317a <=( a88316a  and  a88309a );
 a88320a <=( (not A267)  and  (not A266) );
 a88323a <=( A269  and  (not A268) );
 a88324a <=( a88323a  and  a88320a );
 a88327a <=( (not A299)  and  A298 );
 a88330a <=( (not A302)  and  A300 );
 a88331a <=( a88330a  and  a88327a );
 a88332a <=( a88331a  and  a88324a );
 a88336a <=( A199  and  (not A168) );
 a88337a <=( A169  and  a88336a );
 a88340a <=( A201  and  (not A200) );
 a88343a <=( A265  and  (not A203) );
 a88344a <=( a88343a  and  a88340a );
 a88345a <=( a88344a  and  a88337a );
 a88348a <=( (not A267)  and  (not A266) );
 a88351a <=( A269  and  (not A268) );
 a88352a <=( a88351a  and  a88348a );
 a88355a <=( A299  and  (not A298) );
 a88358a <=( A301  and  A300 );
 a88359a <=( a88358a  and  a88355a );
 a88360a <=( a88359a  and  a88352a );
 a88364a <=( A199  and  (not A168) );
 a88365a <=( A169  and  a88364a );
 a88368a <=( A201  and  (not A200) );
 a88371a <=( A265  and  (not A203) );
 a88372a <=( a88371a  and  a88368a );
 a88373a <=( a88372a  and  a88365a );
 a88376a <=( (not A267)  and  (not A266) );
 a88379a <=( A269  and  (not A268) );
 a88380a <=( a88379a  and  a88376a );
 a88383a <=( A299  and  (not A298) );
 a88386a <=( (not A302)  and  A300 );
 a88387a <=( a88386a  and  a88383a );
 a88388a <=( a88387a  and  a88380a );
 a88392a <=( A199  and  (not A168) );
 a88393a <=( A169  and  a88392a );
 a88396a <=( (not A201)  and  (not A200) );
 a88399a <=( A203  and  (not A202) );
 a88400a <=( a88399a  and  a88396a );
 a88401a <=( a88400a  and  a88393a );
 a88404a <=( A266  and  (not A265) );
 a88407a <=( A268  and  A267 );
 a88408a <=( a88407a  and  a88404a );
 a88411a <=( (not A299)  and  A298 );
 a88414a <=( A301  and  A300 );
 a88415a <=( a88414a  and  a88411a );
 a88416a <=( a88415a  and  a88408a );
 a88420a <=( A199  and  (not A168) );
 a88421a <=( A169  and  a88420a );
 a88424a <=( (not A201)  and  (not A200) );
 a88427a <=( A203  and  (not A202) );
 a88428a <=( a88427a  and  a88424a );
 a88429a <=( a88428a  and  a88421a );
 a88432a <=( A266  and  (not A265) );
 a88435a <=( A268  and  A267 );
 a88436a <=( a88435a  and  a88432a );
 a88439a <=( (not A299)  and  A298 );
 a88442a <=( (not A302)  and  A300 );
 a88443a <=( a88442a  and  a88439a );
 a88444a <=( a88443a  and  a88436a );
 a88448a <=( A199  and  (not A168) );
 a88449a <=( A169  and  a88448a );
 a88452a <=( (not A201)  and  (not A200) );
 a88455a <=( A203  and  (not A202) );
 a88456a <=( a88455a  and  a88452a );
 a88457a <=( a88456a  and  a88449a );
 a88460a <=( A266  and  (not A265) );
 a88463a <=( A268  and  A267 );
 a88464a <=( a88463a  and  a88460a );
 a88467a <=( A299  and  (not A298) );
 a88470a <=( A301  and  A300 );
 a88471a <=( a88470a  and  a88467a );
 a88472a <=( a88471a  and  a88464a );
 a88476a <=( A199  and  (not A168) );
 a88477a <=( A169  and  a88476a );
 a88480a <=( (not A201)  and  (not A200) );
 a88483a <=( A203  and  (not A202) );
 a88484a <=( a88483a  and  a88480a );
 a88485a <=( a88484a  and  a88477a );
 a88488a <=( A266  and  (not A265) );
 a88491a <=( A268  and  A267 );
 a88492a <=( a88491a  and  a88488a );
 a88495a <=( A299  and  (not A298) );
 a88498a <=( (not A302)  and  A300 );
 a88499a <=( a88498a  and  a88495a );
 a88500a <=( a88499a  and  a88492a );
 a88504a <=( A199  and  (not A168) );
 a88505a <=( A169  and  a88504a );
 a88508a <=( (not A201)  and  (not A200) );
 a88511a <=( A203  and  (not A202) );
 a88512a <=( a88511a  and  a88508a );
 a88513a <=( a88512a  and  a88505a );
 a88516a <=( A266  and  (not A265) );
 a88519a <=( (not A269)  and  A267 );
 a88520a <=( a88519a  and  a88516a );
 a88523a <=( (not A299)  and  A298 );
 a88526a <=( A301  and  A300 );
 a88527a <=( a88526a  and  a88523a );
 a88528a <=( a88527a  and  a88520a );
 a88532a <=( A199  and  (not A168) );
 a88533a <=( A169  and  a88532a );
 a88536a <=( (not A201)  and  (not A200) );
 a88539a <=( A203  and  (not A202) );
 a88540a <=( a88539a  and  a88536a );
 a88541a <=( a88540a  and  a88533a );
 a88544a <=( A266  and  (not A265) );
 a88547a <=( (not A269)  and  A267 );
 a88548a <=( a88547a  and  a88544a );
 a88551a <=( (not A299)  and  A298 );
 a88554a <=( (not A302)  and  A300 );
 a88555a <=( a88554a  and  a88551a );
 a88556a <=( a88555a  and  a88548a );
 a88560a <=( A199  and  (not A168) );
 a88561a <=( A169  and  a88560a );
 a88564a <=( (not A201)  and  (not A200) );
 a88567a <=( A203  and  (not A202) );
 a88568a <=( a88567a  and  a88564a );
 a88569a <=( a88568a  and  a88561a );
 a88572a <=( A266  and  (not A265) );
 a88575a <=( (not A269)  and  A267 );
 a88576a <=( a88575a  and  a88572a );
 a88579a <=( A299  and  (not A298) );
 a88582a <=( A301  and  A300 );
 a88583a <=( a88582a  and  a88579a );
 a88584a <=( a88583a  and  a88576a );
 a88588a <=( A199  and  (not A168) );
 a88589a <=( A169  and  a88588a );
 a88592a <=( (not A201)  and  (not A200) );
 a88595a <=( A203  and  (not A202) );
 a88596a <=( a88595a  and  a88592a );
 a88597a <=( a88596a  and  a88589a );
 a88600a <=( A266  and  (not A265) );
 a88603a <=( (not A269)  and  A267 );
 a88604a <=( a88603a  and  a88600a );
 a88607a <=( A299  and  (not A298) );
 a88610a <=( (not A302)  and  A300 );
 a88611a <=( a88610a  and  a88607a );
 a88612a <=( a88611a  and  a88604a );
 a88616a <=( A199  and  (not A168) );
 a88617a <=( A169  and  a88616a );
 a88620a <=( (not A201)  and  (not A200) );
 a88623a <=( A203  and  (not A202) );
 a88624a <=( a88623a  and  a88620a );
 a88625a <=( a88624a  and  a88617a );
 a88628a <=( (not A266)  and  A265 );
 a88631a <=( A268  and  A267 );
 a88632a <=( a88631a  and  a88628a );
 a88635a <=( (not A299)  and  A298 );
 a88638a <=( A301  and  A300 );
 a88639a <=( a88638a  and  a88635a );
 a88640a <=( a88639a  and  a88632a );
 a88644a <=( A199  and  (not A168) );
 a88645a <=( A169  and  a88644a );
 a88648a <=( (not A201)  and  (not A200) );
 a88651a <=( A203  and  (not A202) );
 a88652a <=( a88651a  and  a88648a );
 a88653a <=( a88652a  and  a88645a );
 a88656a <=( (not A266)  and  A265 );
 a88659a <=( A268  and  A267 );
 a88660a <=( a88659a  and  a88656a );
 a88663a <=( (not A299)  and  A298 );
 a88666a <=( (not A302)  and  A300 );
 a88667a <=( a88666a  and  a88663a );
 a88668a <=( a88667a  and  a88660a );
 a88672a <=( A199  and  (not A168) );
 a88673a <=( A169  and  a88672a );
 a88676a <=( (not A201)  and  (not A200) );
 a88679a <=( A203  and  (not A202) );
 a88680a <=( a88679a  and  a88676a );
 a88681a <=( a88680a  and  a88673a );
 a88684a <=( (not A266)  and  A265 );
 a88687a <=( A268  and  A267 );
 a88688a <=( a88687a  and  a88684a );
 a88691a <=( A299  and  (not A298) );
 a88694a <=( A301  and  A300 );
 a88695a <=( a88694a  and  a88691a );
 a88696a <=( a88695a  and  a88688a );
 a88700a <=( A199  and  (not A168) );
 a88701a <=( A169  and  a88700a );
 a88704a <=( (not A201)  and  (not A200) );
 a88707a <=( A203  and  (not A202) );
 a88708a <=( a88707a  and  a88704a );
 a88709a <=( a88708a  and  a88701a );
 a88712a <=( (not A266)  and  A265 );
 a88715a <=( A268  and  A267 );
 a88716a <=( a88715a  and  a88712a );
 a88719a <=( A299  and  (not A298) );
 a88722a <=( (not A302)  and  A300 );
 a88723a <=( a88722a  and  a88719a );
 a88724a <=( a88723a  and  a88716a );
 a88728a <=( A199  and  (not A168) );
 a88729a <=( A169  and  a88728a );
 a88732a <=( (not A201)  and  (not A200) );
 a88735a <=( A203  and  (not A202) );
 a88736a <=( a88735a  and  a88732a );
 a88737a <=( a88736a  and  a88729a );
 a88740a <=( (not A266)  and  A265 );
 a88743a <=( (not A269)  and  A267 );
 a88744a <=( a88743a  and  a88740a );
 a88747a <=( (not A299)  and  A298 );
 a88750a <=( A301  and  A300 );
 a88751a <=( a88750a  and  a88747a );
 a88752a <=( a88751a  and  a88744a );
 a88756a <=( A199  and  (not A168) );
 a88757a <=( A169  and  a88756a );
 a88760a <=( (not A201)  and  (not A200) );
 a88763a <=( A203  and  (not A202) );
 a88764a <=( a88763a  and  a88760a );
 a88765a <=( a88764a  and  a88757a );
 a88768a <=( (not A266)  and  A265 );
 a88771a <=( (not A269)  and  A267 );
 a88772a <=( a88771a  and  a88768a );
 a88775a <=( (not A299)  and  A298 );
 a88778a <=( (not A302)  and  A300 );
 a88779a <=( a88778a  and  a88775a );
 a88780a <=( a88779a  and  a88772a );
 a88784a <=( A199  and  (not A168) );
 a88785a <=( A169  and  a88784a );
 a88788a <=( (not A201)  and  (not A200) );
 a88791a <=( A203  and  (not A202) );
 a88792a <=( a88791a  and  a88788a );
 a88793a <=( a88792a  and  a88785a );
 a88796a <=( (not A266)  and  A265 );
 a88799a <=( (not A269)  and  A267 );
 a88800a <=( a88799a  and  a88796a );
 a88803a <=( A299  and  (not A298) );
 a88806a <=( A301  and  A300 );
 a88807a <=( a88806a  and  a88803a );
 a88808a <=( a88807a  and  a88800a );
 a88812a <=( A199  and  (not A168) );
 a88813a <=( A169  and  a88812a );
 a88816a <=( (not A201)  and  (not A200) );
 a88819a <=( A203  and  (not A202) );
 a88820a <=( a88819a  and  a88816a );
 a88821a <=( a88820a  and  a88813a );
 a88824a <=( (not A266)  and  A265 );
 a88827a <=( (not A269)  and  A267 );
 a88828a <=( a88827a  and  a88824a );
 a88831a <=( A299  and  (not A298) );
 a88834a <=( (not A302)  and  A300 );
 a88835a <=( a88834a  and  a88831a );
 a88836a <=( a88835a  and  a88828a );
 a88840a <=( A168  and  (not A169) );
 a88841a <=( (not A170)  and  a88840a );
 a88844a <=( A200  and  (not A199) );
 a88847a <=( A202  and  A201 );
 a88848a <=( a88847a  and  a88844a );
 a88849a <=( a88848a  and  a88841a );
 a88852a <=( A266  and  (not A265) );
 a88855a <=( A268  and  A267 );
 a88856a <=( a88855a  and  a88852a );
 a88859a <=( (not A299)  and  A298 );
 a88862a <=( A301  and  A300 );
 a88863a <=( a88862a  and  a88859a );
 a88864a <=( a88863a  and  a88856a );
 a88868a <=( A168  and  (not A169) );
 a88869a <=( (not A170)  and  a88868a );
 a88872a <=( A200  and  (not A199) );
 a88875a <=( A202  and  A201 );
 a88876a <=( a88875a  and  a88872a );
 a88877a <=( a88876a  and  a88869a );
 a88880a <=( A266  and  (not A265) );
 a88883a <=( A268  and  A267 );
 a88884a <=( a88883a  and  a88880a );
 a88887a <=( (not A299)  and  A298 );
 a88890a <=( (not A302)  and  A300 );
 a88891a <=( a88890a  and  a88887a );
 a88892a <=( a88891a  and  a88884a );
 a88896a <=( A168  and  (not A169) );
 a88897a <=( (not A170)  and  a88896a );
 a88900a <=( A200  and  (not A199) );
 a88903a <=( A202  and  A201 );
 a88904a <=( a88903a  and  a88900a );
 a88905a <=( a88904a  and  a88897a );
 a88908a <=( A266  and  (not A265) );
 a88911a <=( A268  and  A267 );
 a88912a <=( a88911a  and  a88908a );
 a88915a <=( A299  and  (not A298) );
 a88918a <=( A301  and  A300 );
 a88919a <=( a88918a  and  a88915a );
 a88920a <=( a88919a  and  a88912a );
 a88924a <=( A168  and  (not A169) );
 a88925a <=( (not A170)  and  a88924a );
 a88928a <=( A200  and  (not A199) );
 a88931a <=( A202  and  A201 );
 a88932a <=( a88931a  and  a88928a );
 a88933a <=( a88932a  and  a88925a );
 a88936a <=( A266  and  (not A265) );
 a88939a <=( A268  and  A267 );
 a88940a <=( a88939a  and  a88936a );
 a88943a <=( A299  and  (not A298) );
 a88946a <=( (not A302)  and  A300 );
 a88947a <=( a88946a  and  a88943a );
 a88948a <=( a88947a  and  a88940a );
 a88952a <=( A168  and  (not A169) );
 a88953a <=( (not A170)  and  a88952a );
 a88956a <=( A200  and  (not A199) );
 a88959a <=( A202  and  A201 );
 a88960a <=( a88959a  and  a88956a );
 a88961a <=( a88960a  and  a88953a );
 a88964a <=( A266  and  (not A265) );
 a88967a <=( (not A269)  and  A267 );
 a88968a <=( a88967a  and  a88964a );
 a88971a <=( (not A299)  and  A298 );
 a88974a <=( A301  and  A300 );
 a88975a <=( a88974a  and  a88971a );
 a88976a <=( a88975a  and  a88968a );
 a88980a <=( A168  and  (not A169) );
 a88981a <=( (not A170)  and  a88980a );
 a88984a <=( A200  and  (not A199) );
 a88987a <=( A202  and  A201 );
 a88988a <=( a88987a  and  a88984a );
 a88989a <=( a88988a  and  a88981a );
 a88992a <=( A266  and  (not A265) );
 a88995a <=( (not A269)  and  A267 );
 a88996a <=( a88995a  and  a88992a );
 a88999a <=( (not A299)  and  A298 );
 a89002a <=( (not A302)  and  A300 );
 a89003a <=( a89002a  and  a88999a );
 a89004a <=( a89003a  and  a88996a );
 a89008a <=( A168  and  (not A169) );
 a89009a <=( (not A170)  and  a89008a );
 a89012a <=( A200  and  (not A199) );
 a89015a <=( A202  and  A201 );
 a89016a <=( a89015a  and  a89012a );
 a89017a <=( a89016a  and  a89009a );
 a89020a <=( A266  and  (not A265) );
 a89023a <=( (not A269)  and  A267 );
 a89024a <=( a89023a  and  a89020a );
 a89027a <=( A299  and  (not A298) );
 a89030a <=( A301  and  A300 );
 a89031a <=( a89030a  and  a89027a );
 a89032a <=( a89031a  and  a89024a );
 a89036a <=( A168  and  (not A169) );
 a89037a <=( (not A170)  and  a89036a );
 a89040a <=( A200  and  (not A199) );
 a89043a <=( A202  and  A201 );
 a89044a <=( a89043a  and  a89040a );
 a89045a <=( a89044a  and  a89037a );
 a89048a <=( A266  and  (not A265) );
 a89051a <=( (not A269)  and  A267 );
 a89052a <=( a89051a  and  a89048a );
 a89055a <=( A299  and  (not A298) );
 a89058a <=( (not A302)  and  A300 );
 a89059a <=( a89058a  and  a89055a );
 a89060a <=( a89059a  and  a89052a );
 a89064a <=( A168  and  (not A169) );
 a89065a <=( (not A170)  and  a89064a );
 a89068a <=( A200  and  (not A199) );
 a89071a <=( A202  and  A201 );
 a89072a <=( a89071a  and  a89068a );
 a89073a <=( a89072a  and  a89065a );
 a89076a <=( (not A266)  and  A265 );
 a89079a <=( A268  and  A267 );
 a89080a <=( a89079a  and  a89076a );
 a89083a <=( (not A299)  and  A298 );
 a89086a <=( A301  and  A300 );
 a89087a <=( a89086a  and  a89083a );
 a89088a <=( a89087a  and  a89080a );
 a89092a <=( A168  and  (not A169) );
 a89093a <=( (not A170)  and  a89092a );
 a89096a <=( A200  and  (not A199) );
 a89099a <=( A202  and  A201 );
 a89100a <=( a89099a  and  a89096a );
 a89101a <=( a89100a  and  a89093a );
 a89104a <=( (not A266)  and  A265 );
 a89107a <=( A268  and  A267 );
 a89108a <=( a89107a  and  a89104a );
 a89111a <=( (not A299)  and  A298 );
 a89114a <=( (not A302)  and  A300 );
 a89115a <=( a89114a  and  a89111a );
 a89116a <=( a89115a  and  a89108a );
 a89120a <=( A168  and  (not A169) );
 a89121a <=( (not A170)  and  a89120a );
 a89124a <=( A200  and  (not A199) );
 a89127a <=( A202  and  A201 );
 a89128a <=( a89127a  and  a89124a );
 a89129a <=( a89128a  and  a89121a );
 a89132a <=( (not A266)  and  A265 );
 a89135a <=( A268  and  A267 );
 a89136a <=( a89135a  and  a89132a );
 a89139a <=( A299  and  (not A298) );
 a89142a <=( A301  and  A300 );
 a89143a <=( a89142a  and  a89139a );
 a89144a <=( a89143a  and  a89136a );
 a89148a <=( A168  and  (not A169) );
 a89149a <=( (not A170)  and  a89148a );
 a89152a <=( A200  and  (not A199) );
 a89155a <=( A202  and  A201 );
 a89156a <=( a89155a  and  a89152a );
 a89157a <=( a89156a  and  a89149a );
 a89160a <=( (not A266)  and  A265 );
 a89163a <=( A268  and  A267 );
 a89164a <=( a89163a  and  a89160a );
 a89167a <=( A299  and  (not A298) );
 a89170a <=( (not A302)  and  A300 );
 a89171a <=( a89170a  and  a89167a );
 a89172a <=( a89171a  and  a89164a );
 a89176a <=( A168  and  (not A169) );
 a89177a <=( (not A170)  and  a89176a );
 a89180a <=( A200  and  (not A199) );
 a89183a <=( A202  and  A201 );
 a89184a <=( a89183a  and  a89180a );
 a89185a <=( a89184a  and  a89177a );
 a89188a <=( (not A266)  and  A265 );
 a89191a <=( (not A269)  and  A267 );
 a89192a <=( a89191a  and  a89188a );
 a89195a <=( (not A299)  and  A298 );
 a89198a <=( A301  and  A300 );
 a89199a <=( a89198a  and  a89195a );
 a89200a <=( a89199a  and  a89192a );
 a89204a <=( A168  and  (not A169) );
 a89205a <=( (not A170)  and  a89204a );
 a89208a <=( A200  and  (not A199) );
 a89211a <=( A202  and  A201 );
 a89212a <=( a89211a  and  a89208a );
 a89213a <=( a89212a  and  a89205a );
 a89216a <=( (not A266)  and  A265 );
 a89219a <=( (not A269)  and  A267 );
 a89220a <=( a89219a  and  a89216a );
 a89223a <=( (not A299)  and  A298 );
 a89226a <=( (not A302)  and  A300 );
 a89227a <=( a89226a  and  a89223a );
 a89228a <=( a89227a  and  a89220a );
 a89232a <=( A168  and  (not A169) );
 a89233a <=( (not A170)  and  a89232a );
 a89236a <=( A200  and  (not A199) );
 a89239a <=( A202  and  A201 );
 a89240a <=( a89239a  and  a89236a );
 a89241a <=( a89240a  and  a89233a );
 a89244a <=( (not A266)  and  A265 );
 a89247a <=( (not A269)  and  A267 );
 a89248a <=( a89247a  and  a89244a );
 a89251a <=( A299  and  (not A298) );
 a89254a <=( A301  and  A300 );
 a89255a <=( a89254a  and  a89251a );
 a89256a <=( a89255a  and  a89248a );
 a89260a <=( A168  and  (not A169) );
 a89261a <=( (not A170)  and  a89260a );
 a89264a <=( A200  and  (not A199) );
 a89267a <=( A202  and  A201 );
 a89268a <=( a89267a  and  a89264a );
 a89269a <=( a89268a  and  a89261a );
 a89272a <=( (not A266)  and  A265 );
 a89275a <=( (not A269)  and  A267 );
 a89276a <=( a89275a  and  a89272a );
 a89279a <=( A299  and  (not A298) );
 a89282a <=( (not A302)  and  A300 );
 a89283a <=( a89282a  and  a89279a );
 a89284a <=( a89283a  and  a89276a );
 a89288a <=( A168  and  (not A169) );
 a89289a <=( (not A170)  and  a89288a );
 a89292a <=( A200  and  (not A199) );
 a89295a <=( (not A203)  and  A201 );
 a89296a <=( a89295a  and  a89292a );
 a89297a <=( a89296a  and  a89289a );
 a89300a <=( A266  and  (not A265) );
 a89303a <=( A268  and  A267 );
 a89304a <=( a89303a  and  a89300a );
 a89307a <=( (not A299)  and  A298 );
 a89310a <=( A301  and  A300 );
 a89311a <=( a89310a  and  a89307a );
 a89312a <=( a89311a  and  a89304a );
 a89316a <=( A168  and  (not A169) );
 a89317a <=( (not A170)  and  a89316a );
 a89320a <=( A200  and  (not A199) );
 a89323a <=( (not A203)  and  A201 );
 a89324a <=( a89323a  and  a89320a );
 a89325a <=( a89324a  and  a89317a );
 a89328a <=( A266  and  (not A265) );
 a89331a <=( A268  and  A267 );
 a89332a <=( a89331a  and  a89328a );
 a89335a <=( (not A299)  and  A298 );
 a89338a <=( (not A302)  and  A300 );
 a89339a <=( a89338a  and  a89335a );
 a89340a <=( a89339a  and  a89332a );
 a89344a <=( A168  and  (not A169) );
 a89345a <=( (not A170)  and  a89344a );
 a89348a <=( A200  and  (not A199) );
 a89351a <=( (not A203)  and  A201 );
 a89352a <=( a89351a  and  a89348a );
 a89353a <=( a89352a  and  a89345a );
 a89356a <=( A266  and  (not A265) );
 a89359a <=( A268  and  A267 );
 a89360a <=( a89359a  and  a89356a );
 a89363a <=( A299  and  (not A298) );
 a89366a <=( A301  and  A300 );
 a89367a <=( a89366a  and  a89363a );
 a89368a <=( a89367a  and  a89360a );
 a89372a <=( A168  and  (not A169) );
 a89373a <=( (not A170)  and  a89372a );
 a89376a <=( A200  and  (not A199) );
 a89379a <=( (not A203)  and  A201 );
 a89380a <=( a89379a  and  a89376a );
 a89381a <=( a89380a  and  a89373a );
 a89384a <=( A266  and  (not A265) );
 a89387a <=( A268  and  A267 );
 a89388a <=( a89387a  and  a89384a );
 a89391a <=( A299  and  (not A298) );
 a89394a <=( (not A302)  and  A300 );
 a89395a <=( a89394a  and  a89391a );
 a89396a <=( a89395a  and  a89388a );
 a89400a <=( A168  and  (not A169) );
 a89401a <=( (not A170)  and  a89400a );
 a89404a <=( A200  and  (not A199) );
 a89407a <=( (not A203)  and  A201 );
 a89408a <=( a89407a  and  a89404a );
 a89409a <=( a89408a  and  a89401a );
 a89412a <=( A266  and  (not A265) );
 a89415a <=( (not A269)  and  A267 );
 a89416a <=( a89415a  and  a89412a );
 a89419a <=( (not A299)  and  A298 );
 a89422a <=( A301  and  A300 );
 a89423a <=( a89422a  and  a89419a );
 a89424a <=( a89423a  and  a89416a );
 a89428a <=( A168  and  (not A169) );
 a89429a <=( (not A170)  and  a89428a );
 a89432a <=( A200  and  (not A199) );
 a89435a <=( (not A203)  and  A201 );
 a89436a <=( a89435a  and  a89432a );
 a89437a <=( a89436a  and  a89429a );
 a89440a <=( A266  and  (not A265) );
 a89443a <=( (not A269)  and  A267 );
 a89444a <=( a89443a  and  a89440a );
 a89447a <=( (not A299)  and  A298 );
 a89450a <=( (not A302)  and  A300 );
 a89451a <=( a89450a  and  a89447a );
 a89452a <=( a89451a  and  a89444a );
 a89456a <=( A168  and  (not A169) );
 a89457a <=( (not A170)  and  a89456a );
 a89460a <=( A200  and  (not A199) );
 a89463a <=( (not A203)  and  A201 );
 a89464a <=( a89463a  and  a89460a );
 a89465a <=( a89464a  and  a89457a );
 a89468a <=( A266  and  (not A265) );
 a89471a <=( (not A269)  and  A267 );
 a89472a <=( a89471a  and  a89468a );
 a89475a <=( A299  and  (not A298) );
 a89478a <=( A301  and  A300 );
 a89479a <=( a89478a  and  a89475a );
 a89480a <=( a89479a  and  a89472a );
 a89484a <=( A168  and  (not A169) );
 a89485a <=( (not A170)  and  a89484a );
 a89488a <=( A200  and  (not A199) );
 a89491a <=( (not A203)  and  A201 );
 a89492a <=( a89491a  and  a89488a );
 a89493a <=( a89492a  and  a89485a );
 a89496a <=( A266  and  (not A265) );
 a89499a <=( (not A269)  and  A267 );
 a89500a <=( a89499a  and  a89496a );
 a89503a <=( A299  and  (not A298) );
 a89506a <=( (not A302)  and  A300 );
 a89507a <=( a89506a  and  a89503a );
 a89508a <=( a89507a  and  a89500a );
 a89512a <=( A168  and  (not A169) );
 a89513a <=( (not A170)  and  a89512a );
 a89516a <=( A200  and  (not A199) );
 a89519a <=( (not A203)  and  A201 );
 a89520a <=( a89519a  and  a89516a );
 a89521a <=( a89520a  and  a89513a );
 a89524a <=( (not A266)  and  A265 );
 a89527a <=( A268  and  A267 );
 a89528a <=( a89527a  and  a89524a );
 a89531a <=( (not A299)  and  A298 );
 a89534a <=( A301  and  A300 );
 a89535a <=( a89534a  and  a89531a );
 a89536a <=( a89535a  and  a89528a );
 a89540a <=( A168  and  (not A169) );
 a89541a <=( (not A170)  and  a89540a );
 a89544a <=( A200  and  (not A199) );
 a89547a <=( (not A203)  and  A201 );
 a89548a <=( a89547a  and  a89544a );
 a89549a <=( a89548a  and  a89541a );
 a89552a <=( (not A266)  and  A265 );
 a89555a <=( A268  and  A267 );
 a89556a <=( a89555a  and  a89552a );
 a89559a <=( (not A299)  and  A298 );
 a89562a <=( (not A302)  and  A300 );
 a89563a <=( a89562a  and  a89559a );
 a89564a <=( a89563a  and  a89556a );
 a89568a <=( A168  and  (not A169) );
 a89569a <=( (not A170)  and  a89568a );
 a89572a <=( A200  and  (not A199) );
 a89575a <=( (not A203)  and  A201 );
 a89576a <=( a89575a  and  a89572a );
 a89577a <=( a89576a  and  a89569a );
 a89580a <=( (not A266)  and  A265 );
 a89583a <=( A268  and  A267 );
 a89584a <=( a89583a  and  a89580a );
 a89587a <=( A299  and  (not A298) );
 a89590a <=( A301  and  A300 );
 a89591a <=( a89590a  and  a89587a );
 a89592a <=( a89591a  and  a89584a );
 a89596a <=( A168  and  (not A169) );
 a89597a <=( (not A170)  and  a89596a );
 a89600a <=( A200  and  (not A199) );
 a89603a <=( (not A203)  and  A201 );
 a89604a <=( a89603a  and  a89600a );
 a89605a <=( a89604a  and  a89597a );
 a89608a <=( (not A266)  and  A265 );
 a89611a <=( A268  and  A267 );
 a89612a <=( a89611a  and  a89608a );
 a89615a <=( A299  and  (not A298) );
 a89618a <=( (not A302)  and  A300 );
 a89619a <=( a89618a  and  a89615a );
 a89620a <=( a89619a  and  a89612a );
 a89624a <=( A168  and  (not A169) );
 a89625a <=( (not A170)  and  a89624a );
 a89628a <=( A200  and  (not A199) );
 a89631a <=( (not A203)  and  A201 );
 a89632a <=( a89631a  and  a89628a );
 a89633a <=( a89632a  and  a89625a );
 a89636a <=( (not A266)  and  A265 );
 a89639a <=( (not A269)  and  A267 );
 a89640a <=( a89639a  and  a89636a );
 a89643a <=( (not A299)  and  A298 );
 a89646a <=( A301  and  A300 );
 a89647a <=( a89646a  and  a89643a );
 a89648a <=( a89647a  and  a89640a );
 a89652a <=( A168  and  (not A169) );
 a89653a <=( (not A170)  and  a89652a );
 a89656a <=( A200  and  (not A199) );
 a89659a <=( (not A203)  and  A201 );
 a89660a <=( a89659a  and  a89656a );
 a89661a <=( a89660a  and  a89653a );
 a89664a <=( (not A266)  and  A265 );
 a89667a <=( (not A269)  and  A267 );
 a89668a <=( a89667a  and  a89664a );
 a89671a <=( (not A299)  and  A298 );
 a89674a <=( (not A302)  and  A300 );
 a89675a <=( a89674a  and  a89671a );
 a89676a <=( a89675a  and  a89668a );
 a89680a <=( A168  and  (not A169) );
 a89681a <=( (not A170)  and  a89680a );
 a89684a <=( A200  and  (not A199) );
 a89687a <=( (not A203)  and  A201 );
 a89688a <=( a89687a  and  a89684a );
 a89689a <=( a89688a  and  a89681a );
 a89692a <=( (not A266)  and  A265 );
 a89695a <=( (not A269)  and  A267 );
 a89696a <=( a89695a  and  a89692a );
 a89699a <=( A299  and  (not A298) );
 a89702a <=( A301  and  A300 );
 a89703a <=( a89702a  and  a89699a );
 a89704a <=( a89703a  and  a89696a );
 a89708a <=( A168  and  (not A169) );
 a89709a <=( (not A170)  and  a89708a );
 a89712a <=( A200  and  (not A199) );
 a89715a <=( (not A203)  and  A201 );
 a89716a <=( a89715a  and  a89712a );
 a89717a <=( a89716a  and  a89709a );
 a89720a <=( (not A266)  and  A265 );
 a89723a <=( (not A269)  and  A267 );
 a89724a <=( a89723a  and  a89720a );
 a89727a <=( A299  and  (not A298) );
 a89730a <=( (not A302)  and  A300 );
 a89731a <=( a89730a  and  a89727a );
 a89732a <=( a89731a  and  a89724a );
 a89736a <=( A168  and  (not A169) );
 a89737a <=( (not A170)  and  a89736a );
 a89740a <=( (not A200)  and  A199 );
 a89743a <=( A202  and  A201 );
 a89744a <=( a89743a  and  a89740a );
 a89745a <=( a89744a  and  a89737a );
 a89748a <=( A266  and  (not A265) );
 a89751a <=( A268  and  A267 );
 a89752a <=( a89751a  and  a89748a );
 a89755a <=( (not A299)  and  A298 );
 a89758a <=( A301  and  A300 );
 a89759a <=( a89758a  and  a89755a );
 a89760a <=( a89759a  and  a89752a );
 a89764a <=( A168  and  (not A169) );
 a89765a <=( (not A170)  and  a89764a );
 a89768a <=( (not A200)  and  A199 );
 a89771a <=( A202  and  A201 );
 a89772a <=( a89771a  and  a89768a );
 a89773a <=( a89772a  and  a89765a );
 a89776a <=( A266  and  (not A265) );
 a89779a <=( A268  and  A267 );
 a89780a <=( a89779a  and  a89776a );
 a89783a <=( (not A299)  and  A298 );
 a89786a <=( (not A302)  and  A300 );
 a89787a <=( a89786a  and  a89783a );
 a89788a <=( a89787a  and  a89780a );
 a89792a <=( A168  and  (not A169) );
 a89793a <=( (not A170)  and  a89792a );
 a89796a <=( (not A200)  and  A199 );
 a89799a <=( A202  and  A201 );
 a89800a <=( a89799a  and  a89796a );
 a89801a <=( a89800a  and  a89793a );
 a89804a <=( A266  and  (not A265) );
 a89807a <=( A268  and  A267 );
 a89808a <=( a89807a  and  a89804a );
 a89811a <=( A299  and  (not A298) );
 a89814a <=( A301  and  A300 );
 a89815a <=( a89814a  and  a89811a );
 a89816a <=( a89815a  and  a89808a );
 a89820a <=( A168  and  (not A169) );
 a89821a <=( (not A170)  and  a89820a );
 a89824a <=( (not A200)  and  A199 );
 a89827a <=( A202  and  A201 );
 a89828a <=( a89827a  and  a89824a );
 a89829a <=( a89828a  and  a89821a );
 a89832a <=( A266  and  (not A265) );
 a89835a <=( A268  and  A267 );
 a89836a <=( a89835a  and  a89832a );
 a89839a <=( A299  and  (not A298) );
 a89842a <=( (not A302)  and  A300 );
 a89843a <=( a89842a  and  a89839a );
 a89844a <=( a89843a  and  a89836a );
 a89848a <=( A168  and  (not A169) );
 a89849a <=( (not A170)  and  a89848a );
 a89852a <=( (not A200)  and  A199 );
 a89855a <=( A202  and  A201 );
 a89856a <=( a89855a  and  a89852a );
 a89857a <=( a89856a  and  a89849a );
 a89860a <=( A266  and  (not A265) );
 a89863a <=( (not A269)  and  A267 );
 a89864a <=( a89863a  and  a89860a );
 a89867a <=( (not A299)  and  A298 );
 a89870a <=( A301  and  A300 );
 a89871a <=( a89870a  and  a89867a );
 a89872a <=( a89871a  and  a89864a );
 a89876a <=( A168  and  (not A169) );
 a89877a <=( (not A170)  and  a89876a );
 a89880a <=( (not A200)  and  A199 );
 a89883a <=( A202  and  A201 );
 a89884a <=( a89883a  and  a89880a );
 a89885a <=( a89884a  and  a89877a );
 a89888a <=( A266  and  (not A265) );
 a89891a <=( (not A269)  and  A267 );
 a89892a <=( a89891a  and  a89888a );
 a89895a <=( (not A299)  and  A298 );
 a89898a <=( (not A302)  and  A300 );
 a89899a <=( a89898a  and  a89895a );
 a89900a <=( a89899a  and  a89892a );
 a89904a <=( A168  and  (not A169) );
 a89905a <=( (not A170)  and  a89904a );
 a89908a <=( (not A200)  and  A199 );
 a89911a <=( A202  and  A201 );
 a89912a <=( a89911a  and  a89908a );
 a89913a <=( a89912a  and  a89905a );
 a89916a <=( A266  and  (not A265) );
 a89919a <=( (not A269)  and  A267 );
 a89920a <=( a89919a  and  a89916a );
 a89923a <=( A299  and  (not A298) );
 a89926a <=( A301  and  A300 );
 a89927a <=( a89926a  and  a89923a );
 a89928a <=( a89927a  and  a89920a );
 a89932a <=( A168  and  (not A169) );
 a89933a <=( (not A170)  and  a89932a );
 a89936a <=( (not A200)  and  A199 );
 a89939a <=( A202  and  A201 );
 a89940a <=( a89939a  and  a89936a );
 a89941a <=( a89940a  and  a89933a );
 a89944a <=( A266  and  (not A265) );
 a89947a <=( (not A269)  and  A267 );
 a89948a <=( a89947a  and  a89944a );
 a89951a <=( A299  and  (not A298) );
 a89954a <=( (not A302)  and  A300 );
 a89955a <=( a89954a  and  a89951a );
 a89956a <=( a89955a  and  a89948a );
 a89960a <=( A168  and  (not A169) );
 a89961a <=( (not A170)  and  a89960a );
 a89964a <=( (not A200)  and  A199 );
 a89967a <=( A202  and  A201 );
 a89968a <=( a89967a  and  a89964a );
 a89969a <=( a89968a  and  a89961a );
 a89972a <=( (not A266)  and  A265 );
 a89975a <=( A268  and  A267 );
 a89976a <=( a89975a  and  a89972a );
 a89979a <=( (not A299)  and  A298 );
 a89982a <=( A301  and  A300 );
 a89983a <=( a89982a  and  a89979a );
 a89984a <=( a89983a  and  a89976a );
 a89988a <=( A168  and  (not A169) );
 a89989a <=( (not A170)  and  a89988a );
 a89992a <=( (not A200)  and  A199 );
 a89995a <=( A202  and  A201 );
 a89996a <=( a89995a  and  a89992a );
 a89997a <=( a89996a  and  a89989a );
 a90000a <=( (not A266)  and  A265 );
 a90003a <=( A268  and  A267 );
 a90004a <=( a90003a  and  a90000a );
 a90007a <=( (not A299)  and  A298 );
 a90010a <=( (not A302)  and  A300 );
 a90011a <=( a90010a  and  a90007a );
 a90012a <=( a90011a  and  a90004a );
 a90016a <=( A168  and  (not A169) );
 a90017a <=( (not A170)  and  a90016a );
 a90020a <=( (not A200)  and  A199 );
 a90023a <=( A202  and  A201 );
 a90024a <=( a90023a  and  a90020a );
 a90025a <=( a90024a  and  a90017a );
 a90028a <=( (not A266)  and  A265 );
 a90031a <=( A268  and  A267 );
 a90032a <=( a90031a  and  a90028a );
 a90035a <=( A299  and  (not A298) );
 a90038a <=( A301  and  A300 );
 a90039a <=( a90038a  and  a90035a );
 a90040a <=( a90039a  and  a90032a );
 a90044a <=( A168  and  (not A169) );
 a90045a <=( (not A170)  and  a90044a );
 a90048a <=( (not A200)  and  A199 );
 a90051a <=( A202  and  A201 );
 a90052a <=( a90051a  and  a90048a );
 a90053a <=( a90052a  and  a90045a );
 a90056a <=( (not A266)  and  A265 );
 a90059a <=( A268  and  A267 );
 a90060a <=( a90059a  and  a90056a );
 a90063a <=( A299  and  (not A298) );
 a90066a <=( (not A302)  and  A300 );
 a90067a <=( a90066a  and  a90063a );
 a90068a <=( a90067a  and  a90060a );
 a90072a <=( A168  and  (not A169) );
 a90073a <=( (not A170)  and  a90072a );
 a90076a <=( (not A200)  and  A199 );
 a90079a <=( A202  and  A201 );
 a90080a <=( a90079a  and  a90076a );
 a90081a <=( a90080a  and  a90073a );
 a90084a <=( (not A266)  and  A265 );
 a90087a <=( (not A269)  and  A267 );
 a90088a <=( a90087a  and  a90084a );
 a90091a <=( (not A299)  and  A298 );
 a90094a <=( A301  and  A300 );
 a90095a <=( a90094a  and  a90091a );
 a90096a <=( a90095a  and  a90088a );
 a90100a <=( A168  and  (not A169) );
 a90101a <=( (not A170)  and  a90100a );
 a90104a <=( (not A200)  and  A199 );
 a90107a <=( A202  and  A201 );
 a90108a <=( a90107a  and  a90104a );
 a90109a <=( a90108a  and  a90101a );
 a90112a <=( (not A266)  and  A265 );
 a90115a <=( (not A269)  and  A267 );
 a90116a <=( a90115a  and  a90112a );
 a90119a <=( (not A299)  and  A298 );
 a90122a <=( (not A302)  and  A300 );
 a90123a <=( a90122a  and  a90119a );
 a90124a <=( a90123a  and  a90116a );
 a90128a <=( A168  and  (not A169) );
 a90129a <=( (not A170)  and  a90128a );
 a90132a <=( (not A200)  and  A199 );
 a90135a <=( A202  and  A201 );
 a90136a <=( a90135a  and  a90132a );
 a90137a <=( a90136a  and  a90129a );
 a90140a <=( (not A266)  and  A265 );
 a90143a <=( (not A269)  and  A267 );
 a90144a <=( a90143a  and  a90140a );
 a90147a <=( A299  and  (not A298) );
 a90150a <=( A301  and  A300 );
 a90151a <=( a90150a  and  a90147a );
 a90152a <=( a90151a  and  a90144a );
 a90156a <=( A168  and  (not A169) );
 a90157a <=( (not A170)  and  a90156a );
 a90160a <=( (not A200)  and  A199 );
 a90163a <=( A202  and  A201 );
 a90164a <=( a90163a  and  a90160a );
 a90165a <=( a90164a  and  a90157a );
 a90168a <=( (not A266)  and  A265 );
 a90171a <=( (not A269)  and  A267 );
 a90172a <=( a90171a  and  a90168a );
 a90175a <=( A299  and  (not A298) );
 a90178a <=( (not A302)  and  A300 );
 a90179a <=( a90178a  and  a90175a );
 a90180a <=( a90179a  and  a90172a );
 a90184a <=( A168  and  (not A169) );
 a90185a <=( (not A170)  and  a90184a );
 a90188a <=( (not A200)  and  A199 );
 a90191a <=( (not A203)  and  A201 );
 a90192a <=( a90191a  and  a90188a );
 a90193a <=( a90192a  and  a90185a );
 a90196a <=( A266  and  (not A265) );
 a90199a <=( A268  and  A267 );
 a90200a <=( a90199a  and  a90196a );
 a90203a <=( (not A299)  and  A298 );
 a90206a <=( A301  and  A300 );
 a90207a <=( a90206a  and  a90203a );
 a90208a <=( a90207a  and  a90200a );
 a90212a <=( A168  and  (not A169) );
 a90213a <=( (not A170)  and  a90212a );
 a90216a <=( (not A200)  and  A199 );
 a90219a <=( (not A203)  and  A201 );
 a90220a <=( a90219a  and  a90216a );
 a90221a <=( a90220a  and  a90213a );
 a90224a <=( A266  and  (not A265) );
 a90227a <=( A268  and  A267 );
 a90228a <=( a90227a  and  a90224a );
 a90231a <=( (not A299)  and  A298 );
 a90234a <=( (not A302)  and  A300 );
 a90235a <=( a90234a  and  a90231a );
 a90236a <=( a90235a  and  a90228a );
 a90240a <=( A168  and  (not A169) );
 a90241a <=( (not A170)  and  a90240a );
 a90244a <=( (not A200)  and  A199 );
 a90247a <=( (not A203)  and  A201 );
 a90248a <=( a90247a  and  a90244a );
 a90249a <=( a90248a  and  a90241a );
 a90252a <=( A266  and  (not A265) );
 a90255a <=( A268  and  A267 );
 a90256a <=( a90255a  and  a90252a );
 a90259a <=( A299  and  (not A298) );
 a90262a <=( A301  and  A300 );
 a90263a <=( a90262a  and  a90259a );
 a90264a <=( a90263a  and  a90256a );
 a90268a <=( A168  and  (not A169) );
 a90269a <=( (not A170)  and  a90268a );
 a90272a <=( (not A200)  and  A199 );
 a90275a <=( (not A203)  and  A201 );
 a90276a <=( a90275a  and  a90272a );
 a90277a <=( a90276a  and  a90269a );
 a90280a <=( A266  and  (not A265) );
 a90283a <=( A268  and  A267 );
 a90284a <=( a90283a  and  a90280a );
 a90287a <=( A299  and  (not A298) );
 a90290a <=( (not A302)  and  A300 );
 a90291a <=( a90290a  and  a90287a );
 a90292a <=( a90291a  and  a90284a );
 a90296a <=( A168  and  (not A169) );
 a90297a <=( (not A170)  and  a90296a );
 a90300a <=( (not A200)  and  A199 );
 a90303a <=( (not A203)  and  A201 );
 a90304a <=( a90303a  and  a90300a );
 a90305a <=( a90304a  and  a90297a );
 a90308a <=( A266  and  (not A265) );
 a90311a <=( (not A269)  and  A267 );
 a90312a <=( a90311a  and  a90308a );
 a90315a <=( (not A299)  and  A298 );
 a90318a <=( A301  and  A300 );
 a90319a <=( a90318a  and  a90315a );
 a90320a <=( a90319a  and  a90312a );
 a90324a <=( A168  and  (not A169) );
 a90325a <=( (not A170)  and  a90324a );
 a90328a <=( (not A200)  and  A199 );
 a90331a <=( (not A203)  and  A201 );
 a90332a <=( a90331a  and  a90328a );
 a90333a <=( a90332a  and  a90325a );
 a90336a <=( A266  and  (not A265) );
 a90339a <=( (not A269)  and  A267 );
 a90340a <=( a90339a  and  a90336a );
 a90343a <=( (not A299)  and  A298 );
 a90346a <=( (not A302)  and  A300 );
 a90347a <=( a90346a  and  a90343a );
 a90348a <=( a90347a  and  a90340a );
 a90352a <=( A168  and  (not A169) );
 a90353a <=( (not A170)  and  a90352a );
 a90356a <=( (not A200)  and  A199 );
 a90359a <=( (not A203)  and  A201 );
 a90360a <=( a90359a  and  a90356a );
 a90361a <=( a90360a  and  a90353a );
 a90364a <=( A266  and  (not A265) );
 a90367a <=( (not A269)  and  A267 );
 a90368a <=( a90367a  and  a90364a );
 a90371a <=( A299  and  (not A298) );
 a90374a <=( A301  and  A300 );
 a90375a <=( a90374a  and  a90371a );
 a90376a <=( a90375a  and  a90368a );
 a90380a <=( A168  and  (not A169) );
 a90381a <=( (not A170)  and  a90380a );
 a90384a <=( (not A200)  and  A199 );
 a90387a <=( (not A203)  and  A201 );
 a90388a <=( a90387a  and  a90384a );
 a90389a <=( a90388a  and  a90381a );
 a90392a <=( A266  and  (not A265) );
 a90395a <=( (not A269)  and  A267 );
 a90396a <=( a90395a  and  a90392a );
 a90399a <=( A299  and  (not A298) );
 a90402a <=( (not A302)  and  A300 );
 a90403a <=( a90402a  and  a90399a );
 a90404a <=( a90403a  and  a90396a );
 a90408a <=( A168  and  (not A169) );
 a90409a <=( (not A170)  and  a90408a );
 a90412a <=( (not A200)  and  A199 );
 a90415a <=( (not A203)  and  A201 );
 a90416a <=( a90415a  and  a90412a );
 a90417a <=( a90416a  and  a90409a );
 a90420a <=( (not A266)  and  A265 );
 a90423a <=( A268  and  A267 );
 a90424a <=( a90423a  and  a90420a );
 a90427a <=( (not A299)  and  A298 );
 a90430a <=( A301  and  A300 );
 a90431a <=( a90430a  and  a90427a );
 a90432a <=( a90431a  and  a90424a );
 a90436a <=( A168  and  (not A169) );
 a90437a <=( (not A170)  and  a90436a );
 a90440a <=( (not A200)  and  A199 );
 a90443a <=( (not A203)  and  A201 );
 a90444a <=( a90443a  and  a90440a );
 a90445a <=( a90444a  and  a90437a );
 a90448a <=( (not A266)  and  A265 );
 a90451a <=( A268  and  A267 );
 a90452a <=( a90451a  and  a90448a );
 a90455a <=( (not A299)  and  A298 );
 a90458a <=( (not A302)  and  A300 );
 a90459a <=( a90458a  and  a90455a );
 a90460a <=( a90459a  and  a90452a );
 a90464a <=( A168  and  (not A169) );
 a90465a <=( (not A170)  and  a90464a );
 a90468a <=( (not A200)  and  A199 );
 a90471a <=( (not A203)  and  A201 );
 a90472a <=( a90471a  and  a90468a );
 a90473a <=( a90472a  and  a90465a );
 a90476a <=( (not A266)  and  A265 );
 a90479a <=( A268  and  A267 );
 a90480a <=( a90479a  and  a90476a );
 a90483a <=( A299  and  (not A298) );
 a90486a <=( A301  and  A300 );
 a90487a <=( a90486a  and  a90483a );
 a90488a <=( a90487a  and  a90480a );
 a90492a <=( A168  and  (not A169) );
 a90493a <=( (not A170)  and  a90492a );
 a90496a <=( (not A200)  and  A199 );
 a90499a <=( (not A203)  and  A201 );
 a90500a <=( a90499a  and  a90496a );
 a90501a <=( a90500a  and  a90493a );
 a90504a <=( (not A266)  and  A265 );
 a90507a <=( A268  and  A267 );
 a90508a <=( a90507a  and  a90504a );
 a90511a <=( A299  and  (not A298) );
 a90514a <=( (not A302)  and  A300 );
 a90515a <=( a90514a  and  a90511a );
 a90516a <=( a90515a  and  a90508a );
 a90520a <=( A168  and  (not A169) );
 a90521a <=( (not A170)  and  a90520a );
 a90524a <=( (not A200)  and  A199 );
 a90527a <=( (not A203)  and  A201 );
 a90528a <=( a90527a  and  a90524a );
 a90529a <=( a90528a  and  a90521a );
 a90532a <=( (not A266)  and  A265 );
 a90535a <=( (not A269)  and  A267 );
 a90536a <=( a90535a  and  a90532a );
 a90539a <=( (not A299)  and  A298 );
 a90542a <=( A301  and  A300 );
 a90543a <=( a90542a  and  a90539a );
 a90544a <=( a90543a  and  a90536a );
 a90548a <=( A168  and  (not A169) );
 a90549a <=( (not A170)  and  a90548a );
 a90552a <=( (not A200)  and  A199 );
 a90555a <=( (not A203)  and  A201 );
 a90556a <=( a90555a  and  a90552a );
 a90557a <=( a90556a  and  a90549a );
 a90560a <=( (not A266)  and  A265 );
 a90563a <=( (not A269)  and  A267 );
 a90564a <=( a90563a  and  a90560a );
 a90567a <=( (not A299)  and  A298 );
 a90570a <=( (not A302)  and  A300 );
 a90571a <=( a90570a  and  a90567a );
 a90572a <=( a90571a  and  a90564a );
 a90576a <=( A168  and  (not A169) );
 a90577a <=( (not A170)  and  a90576a );
 a90580a <=( (not A200)  and  A199 );
 a90583a <=( (not A203)  and  A201 );
 a90584a <=( a90583a  and  a90580a );
 a90585a <=( a90584a  and  a90577a );
 a90588a <=( (not A266)  and  A265 );
 a90591a <=( (not A269)  and  A267 );
 a90592a <=( a90591a  and  a90588a );
 a90595a <=( A299  and  (not A298) );
 a90598a <=( A301  and  A300 );
 a90599a <=( a90598a  and  a90595a );
 a90600a <=( a90599a  and  a90592a );
 a90604a <=( A168  and  (not A169) );
 a90605a <=( (not A170)  and  a90604a );
 a90608a <=( (not A200)  and  A199 );
 a90611a <=( (not A203)  and  A201 );
 a90612a <=( a90611a  and  a90608a );
 a90613a <=( a90612a  and  a90605a );
 a90616a <=( (not A266)  and  A265 );
 a90619a <=( (not A269)  and  A267 );
 a90620a <=( a90619a  and  a90616a );
 a90623a <=( A299  and  (not A298) );
 a90626a <=( (not A302)  and  A300 );
 a90627a <=( a90626a  and  a90623a );
 a90628a <=( a90627a  and  a90620a );
 a90632a <=( (not A168)  and  (not A169) );
 a90633a <=( (not A170)  and  a90632a );
 a90636a <=( (not A166)  and  A167 );
 a90639a <=( (not A202)  and  A201 );
 a90640a <=( a90639a  and  a90636a );
 a90641a <=( a90640a  and  a90633a );
 a90644a <=( A267  and  A203 );
 a90647a <=( A269  and  (not A268) );
 a90648a <=( a90647a  and  a90644a );
 a90651a <=( (not A299)  and  A298 );
 a90654a <=( A301  and  A300 );
 a90655a <=( a90654a  and  a90651a );
 a90656a <=( a90655a  and  a90648a );
 a90660a <=( (not A168)  and  (not A169) );
 a90661a <=( (not A170)  and  a90660a );
 a90664a <=( (not A166)  and  A167 );
 a90667a <=( (not A202)  and  A201 );
 a90668a <=( a90667a  and  a90664a );
 a90669a <=( a90668a  and  a90661a );
 a90672a <=( A267  and  A203 );
 a90675a <=( A269  and  (not A268) );
 a90676a <=( a90675a  and  a90672a );
 a90679a <=( (not A299)  and  A298 );
 a90682a <=( (not A302)  and  A300 );
 a90683a <=( a90682a  and  a90679a );
 a90684a <=( a90683a  and  a90676a );
 a90688a <=( (not A168)  and  (not A169) );
 a90689a <=( (not A170)  and  a90688a );
 a90692a <=( (not A166)  and  A167 );
 a90695a <=( (not A202)  and  A201 );
 a90696a <=( a90695a  and  a90692a );
 a90697a <=( a90696a  and  a90689a );
 a90700a <=( A267  and  A203 );
 a90703a <=( A269  and  (not A268) );
 a90704a <=( a90703a  and  a90700a );
 a90707a <=( A299  and  (not A298) );
 a90710a <=( A301  and  A300 );
 a90711a <=( a90710a  and  a90707a );
 a90712a <=( a90711a  and  a90704a );
 a90716a <=( (not A168)  and  (not A169) );
 a90717a <=( (not A170)  and  a90716a );
 a90720a <=( (not A166)  and  A167 );
 a90723a <=( (not A202)  and  A201 );
 a90724a <=( a90723a  and  a90720a );
 a90725a <=( a90724a  and  a90717a );
 a90728a <=( A267  and  A203 );
 a90731a <=( A269  and  (not A268) );
 a90732a <=( a90731a  and  a90728a );
 a90735a <=( A299  and  (not A298) );
 a90738a <=( (not A302)  and  A300 );
 a90739a <=( a90738a  and  a90735a );
 a90740a <=( a90739a  and  a90732a );
 a90744a <=( (not A168)  and  (not A169) );
 a90745a <=( (not A170)  and  a90744a );
 a90748a <=( (not A166)  and  A167 );
 a90751a <=( (not A202)  and  A201 );
 a90752a <=( a90751a  and  a90748a );
 a90753a <=( a90752a  and  a90745a );
 a90756a <=( (not A267)  and  A203 );
 a90759a <=( A298  and  A268 );
 a90760a <=( a90759a  and  a90756a );
 a90763a <=( (not A300)  and  (not A299) );
 a90766a <=( A302  and  (not A301) );
 a90767a <=( a90766a  and  a90763a );
 a90768a <=( a90767a  and  a90760a );
 a90772a <=( (not A168)  and  (not A169) );
 a90773a <=( (not A170)  and  a90772a );
 a90776a <=( (not A166)  and  A167 );
 a90779a <=( (not A202)  and  A201 );
 a90780a <=( a90779a  and  a90776a );
 a90781a <=( a90780a  and  a90773a );
 a90784a <=( (not A267)  and  A203 );
 a90787a <=( (not A298)  and  A268 );
 a90788a <=( a90787a  and  a90784a );
 a90791a <=( (not A300)  and  A299 );
 a90794a <=( A302  and  (not A301) );
 a90795a <=( a90794a  and  a90791a );
 a90796a <=( a90795a  and  a90788a );
 a90800a <=( (not A168)  and  (not A169) );
 a90801a <=( (not A170)  and  a90800a );
 a90804a <=( (not A166)  and  A167 );
 a90807a <=( (not A202)  and  A201 );
 a90808a <=( a90807a  and  a90804a );
 a90809a <=( a90808a  and  a90801a );
 a90812a <=( (not A267)  and  A203 );
 a90815a <=( A298  and  (not A269) );
 a90816a <=( a90815a  and  a90812a );
 a90819a <=( (not A300)  and  (not A299) );
 a90822a <=( A302  and  (not A301) );
 a90823a <=( a90822a  and  a90819a );
 a90824a <=( a90823a  and  a90816a );
 a90828a <=( (not A168)  and  (not A169) );
 a90829a <=( (not A170)  and  a90828a );
 a90832a <=( (not A166)  and  A167 );
 a90835a <=( (not A202)  and  A201 );
 a90836a <=( a90835a  and  a90832a );
 a90837a <=( a90836a  and  a90829a );
 a90840a <=( (not A267)  and  A203 );
 a90843a <=( (not A298)  and  (not A269) );
 a90844a <=( a90843a  and  a90840a );
 a90847a <=( (not A300)  and  A299 );
 a90850a <=( A302  and  (not A301) );
 a90851a <=( a90850a  and  a90847a );
 a90852a <=( a90851a  and  a90844a );
 a90856a <=( (not A168)  and  (not A169) );
 a90857a <=( (not A170)  and  a90856a );
 a90860a <=( (not A166)  and  A167 );
 a90863a <=( (not A202)  and  A201 );
 a90864a <=( a90863a  and  a90860a );
 a90865a <=( a90864a  and  a90857a );
 a90868a <=( A265  and  A203 );
 a90871a <=( A298  and  A266 );
 a90872a <=( a90871a  and  a90868a );
 a90875a <=( (not A300)  and  (not A299) );
 a90878a <=( A302  and  (not A301) );
 a90879a <=( a90878a  and  a90875a );
 a90880a <=( a90879a  and  a90872a );
 a90884a <=( (not A168)  and  (not A169) );
 a90885a <=( (not A170)  and  a90884a );
 a90888a <=( (not A166)  and  A167 );
 a90891a <=( (not A202)  and  A201 );
 a90892a <=( a90891a  and  a90888a );
 a90893a <=( a90892a  and  a90885a );
 a90896a <=( A265  and  A203 );
 a90899a <=( (not A298)  and  A266 );
 a90900a <=( a90899a  and  a90896a );
 a90903a <=( (not A300)  and  A299 );
 a90906a <=( A302  and  (not A301) );
 a90907a <=( a90906a  and  a90903a );
 a90908a <=( a90907a  and  a90900a );
 a90912a <=( (not A168)  and  (not A169) );
 a90913a <=( (not A170)  and  a90912a );
 a90916a <=( (not A166)  and  A167 );
 a90919a <=( (not A202)  and  A201 );
 a90920a <=( a90919a  and  a90916a );
 a90921a <=( a90920a  and  a90913a );
 a90924a <=( (not A265)  and  A203 );
 a90927a <=( A267  and  A266 );
 a90928a <=( a90927a  and  a90924a );
 a90931a <=( A300  and  A268 );
 a90934a <=( A302  and  (not A301) );
 a90935a <=( a90934a  and  a90931a );
 a90936a <=( a90935a  and  a90928a );
 a90940a <=( (not A168)  and  (not A169) );
 a90941a <=( (not A170)  and  a90940a );
 a90944a <=( (not A166)  and  A167 );
 a90947a <=( (not A202)  and  A201 );
 a90948a <=( a90947a  and  a90944a );
 a90949a <=( a90948a  and  a90941a );
 a90952a <=( (not A265)  and  A203 );
 a90955a <=( A267  and  A266 );
 a90956a <=( a90955a  and  a90952a );
 a90959a <=( A300  and  (not A269) );
 a90962a <=( A302  and  (not A301) );
 a90963a <=( a90962a  and  a90959a );
 a90964a <=( a90963a  and  a90956a );
 a90968a <=( (not A168)  and  (not A169) );
 a90969a <=( (not A170)  and  a90968a );
 a90972a <=( (not A166)  and  A167 );
 a90975a <=( (not A202)  and  A201 );
 a90976a <=( a90975a  and  a90972a );
 a90977a <=( a90976a  and  a90969a );
 a90980a <=( (not A265)  and  A203 );
 a90983a <=( (not A267)  and  A266 );
 a90984a <=( a90983a  and  a90980a );
 a90987a <=( A269  and  (not A268) );
 a90990a <=( A301  and  (not A300) );
 a90991a <=( a90990a  and  a90987a );
 a90992a <=( a90991a  and  a90984a );
 a90996a <=( (not A168)  and  (not A169) );
 a90997a <=( (not A170)  and  a90996a );
 a91000a <=( (not A166)  and  A167 );
 a91003a <=( (not A202)  and  A201 );
 a91004a <=( a91003a  and  a91000a );
 a91005a <=( a91004a  and  a90997a );
 a91008a <=( (not A265)  and  A203 );
 a91011a <=( (not A267)  and  A266 );
 a91012a <=( a91011a  and  a91008a );
 a91015a <=( A269  and  (not A268) );
 a91018a <=( (not A302)  and  (not A300) );
 a91019a <=( a91018a  and  a91015a );
 a91020a <=( a91019a  and  a91012a );
 a91024a <=( (not A168)  and  (not A169) );
 a91025a <=( (not A170)  and  a91024a );
 a91028a <=( (not A166)  and  A167 );
 a91031a <=( (not A202)  and  A201 );
 a91032a <=( a91031a  and  a91028a );
 a91033a <=( a91032a  and  a91025a );
 a91036a <=( (not A265)  and  A203 );
 a91039a <=( (not A267)  and  A266 );
 a91040a <=( a91039a  and  a91036a );
 a91043a <=( A269  and  (not A268) );
 a91046a <=( A299  and  A298 );
 a91047a <=( a91046a  and  a91043a );
 a91048a <=( a91047a  and  a91040a );
 a91052a <=( (not A168)  and  (not A169) );
 a91053a <=( (not A170)  and  a91052a );
 a91056a <=( (not A166)  and  A167 );
 a91059a <=( (not A202)  and  A201 );
 a91060a <=( a91059a  and  a91056a );
 a91061a <=( a91060a  and  a91053a );
 a91064a <=( (not A265)  and  A203 );
 a91067a <=( (not A267)  and  A266 );
 a91068a <=( a91067a  and  a91064a );
 a91071a <=( A269  and  (not A268) );
 a91074a <=( (not A299)  and  (not A298) );
 a91075a <=( a91074a  and  a91071a );
 a91076a <=( a91075a  and  a91068a );
 a91080a <=( (not A168)  and  (not A169) );
 a91081a <=( (not A170)  and  a91080a );
 a91084a <=( (not A166)  and  A167 );
 a91087a <=( (not A202)  and  A201 );
 a91088a <=( a91087a  and  a91084a );
 a91089a <=( a91088a  and  a91081a );
 a91092a <=( A265  and  A203 );
 a91095a <=( A267  and  (not A266) );
 a91096a <=( a91095a  and  a91092a );
 a91099a <=( A300  and  A268 );
 a91102a <=( A302  and  (not A301) );
 a91103a <=( a91102a  and  a91099a );
 a91104a <=( a91103a  and  a91096a );
 a91108a <=( (not A168)  and  (not A169) );
 a91109a <=( (not A170)  and  a91108a );
 a91112a <=( (not A166)  and  A167 );
 a91115a <=( (not A202)  and  A201 );
 a91116a <=( a91115a  and  a91112a );
 a91117a <=( a91116a  and  a91109a );
 a91120a <=( A265  and  A203 );
 a91123a <=( A267  and  (not A266) );
 a91124a <=( a91123a  and  a91120a );
 a91127a <=( A300  and  (not A269) );
 a91130a <=( A302  and  (not A301) );
 a91131a <=( a91130a  and  a91127a );
 a91132a <=( a91131a  and  a91124a );
 a91136a <=( (not A168)  and  (not A169) );
 a91137a <=( (not A170)  and  a91136a );
 a91140a <=( (not A166)  and  A167 );
 a91143a <=( (not A202)  and  A201 );
 a91144a <=( a91143a  and  a91140a );
 a91145a <=( a91144a  and  a91137a );
 a91148a <=( A265  and  A203 );
 a91151a <=( (not A267)  and  (not A266) );
 a91152a <=( a91151a  and  a91148a );
 a91155a <=( A269  and  (not A268) );
 a91158a <=( A301  and  (not A300) );
 a91159a <=( a91158a  and  a91155a );
 a91160a <=( a91159a  and  a91152a );
 a91164a <=( (not A168)  and  (not A169) );
 a91165a <=( (not A170)  and  a91164a );
 a91168a <=( (not A166)  and  A167 );
 a91171a <=( (not A202)  and  A201 );
 a91172a <=( a91171a  and  a91168a );
 a91173a <=( a91172a  and  a91165a );
 a91176a <=( A265  and  A203 );
 a91179a <=( (not A267)  and  (not A266) );
 a91180a <=( a91179a  and  a91176a );
 a91183a <=( A269  and  (not A268) );
 a91186a <=( (not A302)  and  (not A300) );
 a91187a <=( a91186a  and  a91183a );
 a91188a <=( a91187a  and  a91180a );
 a91192a <=( (not A168)  and  (not A169) );
 a91193a <=( (not A170)  and  a91192a );
 a91196a <=( (not A166)  and  A167 );
 a91199a <=( (not A202)  and  A201 );
 a91200a <=( a91199a  and  a91196a );
 a91201a <=( a91200a  and  a91193a );
 a91204a <=( A265  and  A203 );
 a91207a <=( (not A267)  and  (not A266) );
 a91208a <=( a91207a  and  a91204a );
 a91211a <=( A269  and  (not A268) );
 a91214a <=( A299  and  A298 );
 a91215a <=( a91214a  and  a91211a );
 a91216a <=( a91215a  and  a91208a );
 a91220a <=( (not A168)  and  (not A169) );
 a91221a <=( (not A170)  and  a91220a );
 a91224a <=( (not A166)  and  A167 );
 a91227a <=( (not A202)  and  A201 );
 a91228a <=( a91227a  and  a91224a );
 a91229a <=( a91228a  and  a91221a );
 a91232a <=( A265  and  A203 );
 a91235a <=( (not A267)  and  (not A266) );
 a91236a <=( a91235a  and  a91232a );
 a91239a <=( A269  and  (not A268) );
 a91242a <=( (not A299)  and  (not A298) );
 a91243a <=( a91242a  and  a91239a );
 a91244a <=( a91243a  and  a91236a );
 a91248a <=( (not A168)  and  (not A169) );
 a91249a <=( (not A170)  and  a91248a );
 a91252a <=( (not A166)  and  A167 );
 a91255a <=( (not A202)  and  A201 );
 a91256a <=( a91255a  and  a91252a );
 a91257a <=( a91256a  and  a91249a );
 a91260a <=( (not A265)  and  A203 );
 a91263a <=( A298  and  (not A266) );
 a91264a <=( a91263a  and  a91260a );
 a91267a <=( (not A300)  and  (not A299) );
 a91270a <=( A302  and  (not A301) );
 a91271a <=( a91270a  and  a91267a );
 a91272a <=( a91271a  and  a91264a );
 a91276a <=( (not A168)  and  (not A169) );
 a91277a <=( (not A170)  and  a91276a );
 a91280a <=( (not A166)  and  A167 );
 a91283a <=( (not A202)  and  A201 );
 a91284a <=( a91283a  and  a91280a );
 a91285a <=( a91284a  and  a91277a );
 a91288a <=( (not A265)  and  A203 );
 a91291a <=( (not A298)  and  (not A266) );
 a91292a <=( a91291a  and  a91288a );
 a91295a <=( (not A300)  and  A299 );
 a91298a <=( A302  and  (not A301) );
 a91299a <=( a91298a  and  a91295a );
 a91300a <=( a91299a  and  a91292a );
 a91304a <=( (not A168)  and  (not A169) );
 a91305a <=( (not A170)  and  a91304a );
 a91308a <=( (not A166)  and  A167 );
 a91311a <=( A202  and  (not A201) );
 a91312a <=( a91311a  and  a91308a );
 a91313a <=( a91312a  and  a91305a );
 a91316a <=( (not A268)  and  A267 );
 a91319a <=( A298  and  A269 );
 a91320a <=( a91319a  and  a91316a );
 a91323a <=( (not A300)  and  (not A299) );
 a91326a <=( A302  and  (not A301) );
 a91327a <=( a91326a  and  a91323a );
 a91328a <=( a91327a  and  a91320a );
 a91332a <=( (not A168)  and  (not A169) );
 a91333a <=( (not A170)  and  a91332a );
 a91336a <=( (not A166)  and  A167 );
 a91339a <=( A202  and  (not A201) );
 a91340a <=( a91339a  and  a91336a );
 a91341a <=( a91340a  and  a91333a );
 a91344a <=( (not A268)  and  A267 );
 a91347a <=( (not A298)  and  A269 );
 a91348a <=( a91347a  and  a91344a );
 a91351a <=( (not A300)  and  A299 );
 a91354a <=( A302  and  (not A301) );
 a91355a <=( a91354a  and  a91351a );
 a91356a <=( a91355a  and  a91348a );
 a91360a <=( (not A168)  and  (not A169) );
 a91361a <=( (not A170)  and  a91360a );
 a91364a <=( (not A166)  and  A167 );
 a91367a <=( A202  and  (not A201) );
 a91368a <=( a91367a  and  a91364a );
 a91369a <=( a91368a  and  a91361a );
 a91372a <=( A266  and  (not A265) );
 a91375a <=( (not A268)  and  (not A267) );
 a91376a <=( a91375a  and  a91372a );
 a91379a <=( A300  and  A269 );
 a91382a <=( A302  and  (not A301) );
 a91383a <=( a91382a  and  a91379a );
 a91384a <=( a91383a  and  a91376a );
 a91388a <=( (not A168)  and  (not A169) );
 a91389a <=( (not A170)  and  a91388a );
 a91392a <=( (not A166)  and  A167 );
 a91395a <=( A202  and  (not A201) );
 a91396a <=( a91395a  and  a91392a );
 a91397a <=( a91396a  and  a91389a );
 a91400a <=( (not A266)  and  A265 );
 a91403a <=( (not A268)  and  (not A267) );
 a91404a <=( a91403a  and  a91400a );
 a91407a <=( A300  and  A269 );
 a91410a <=( A302  and  (not A301) );
 a91411a <=( a91410a  and  a91407a );
 a91412a <=( a91411a  and  a91404a );
 a91416a <=( (not A168)  and  (not A169) );
 a91417a <=( (not A170)  and  a91416a );
 a91420a <=( (not A166)  and  A167 );
 a91423a <=( (not A203)  and  (not A201) );
 a91424a <=( a91423a  and  a91420a );
 a91425a <=( a91424a  and  a91417a );
 a91428a <=( (not A268)  and  A267 );
 a91431a <=( A298  and  A269 );
 a91432a <=( a91431a  and  a91428a );
 a91435a <=( (not A300)  and  (not A299) );
 a91438a <=( A302  and  (not A301) );
 a91439a <=( a91438a  and  a91435a );
 a91440a <=( a91439a  and  a91432a );
 a91444a <=( (not A168)  and  (not A169) );
 a91445a <=( (not A170)  and  a91444a );
 a91448a <=( (not A166)  and  A167 );
 a91451a <=( (not A203)  and  (not A201) );
 a91452a <=( a91451a  and  a91448a );
 a91453a <=( a91452a  and  a91445a );
 a91456a <=( (not A268)  and  A267 );
 a91459a <=( (not A298)  and  A269 );
 a91460a <=( a91459a  and  a91456a );
 a91463a <=( (not A300)  and  A299 );
 a91466a <=( A302  and  (not A301) );
 a91467a <=( a91466a  and  a91463a );
 a91468a <=( a91467a  and  a91460a );
 a91472a <=( (not A168)  and  (not A169) );
 a91473a <=( (not A170)  and  a91472a );
 a91476a <=( (not A166)  and  A167 );
 a91479a <=( (not A203)  and  (not A201) );
 a91480a <=( a91479a  and  a91476a );
 a91481a <=( a91480a  and  a91473a );
 a91484a <=( A266  and  (not A265) );
 a91487a <=( (not A268)  and  (not A267) );
 a91488a <=( a91487a  and  a91484a );
 a91491a <=( A300  and  A269 );
 a91494a <=( A302  and  (not A301) );
 a91495a <=( a91494a  and  a91491a );
 a91496a <=( a91495a  and  a91488a );
 a91500a <=( (not A168)  and  (not A169) );
 a91501a <=( (not A170)  and  a91500a );
 a91504a <=( (not A166)  and  A167 );
 a91507a <=( (not A203)  and  (not A201) );
 a91508a <=( a91507a  and  a91504a );
 a91509a <=( a91508a  and  a91501a );
 a91512a <=( (not A266)  and  A265 );
 a91515a <=( (not A268)  and  (not A267) );
 a91516a <=( a91515a  and  a91512a );
 a91519a <=( A300  and  A269 );
 a91522a <=( A302  and  (not A301) );
 a91523a <=( a91522a  and  a91519a );
 a91524a <=( a91523a  and  a91516a );
 a91528a <=( (not A168)  and  (not A169) );
 a91529a <=( (not A170)  and  a91528a );
 a91532a <=( (not A166)  and  A167 );
 a91535a <=( A200  and  A199 );
 a91536a <=( a91535a  and  a91532a );
 a91537a <=( a91536a  and  a91529a );
 a91540a <=( (not A268)  and  A267 );
 a91543a <=( A298  and  A269 );
 a91544a <=( a91543a  and  a91540a );
 a91547a <=( (not A300)  and  (not A299) );
 a91550a <=( A302  and  (not A301) );
 a91551a <=( a91550a  and  a91547a );
 a91552a <=( a91551a  and  a91544a );
 a91556a <=( (not A168)  and  (not A169) );
 a91557a <=( (not A170)  and  a91556a );
 a91560a <=( (not A166)  and  A167 );
 a91563a <=( A200  and  A199 );
 a91564a <=( a91563a  and  a91560a );
 a91565a <=( a91564a  and  a91557a );
 a91568a <=( (not A268)  and  A267 );
 a91571a <=( (not A298)  and  A269 );
 a91572a <=( a91571a  and  a91568a );
 a91575a <=( (not A300)  and  A299 );
 a91578a <=( A302  and  (not A301) );
 a91579a <=( a91578a  and  a91575a );
 a91580a <=( a91579a  and  a91572a );
 a91584a <=( (not A168)  and  (not A169) );
 a91585a <=( (not A170)  and  a91584a );
 a91588a <=( (not A166)  and  A167 );
 a91591a <=( A200  and  A199 );
 a91592a <=( a91591a  and  a91588a );
 a91593a <=( a91592a  and  a91585a );
 a91596a <=( A266  and  (not A265) );
 a91599a <=( (not A268)  and  (not A267) );
 a91600a <=( a91599a  and  a91596a );
 a91603a <=( A300  and  A269 );
 a91606a <=( A302  and  (not A301) );
 a91607a <=( a91606a  and  a91603a );
 a91608a <=( a91607a  and  a91600a );
 a91612a <=( (not A168)  and  (not A169) );
 a91613a <=( (not A170)  and  a91612a );
 a91616a <=( (not A166)  and  A167 );
 a91619a <=( A200  and  A199 );
 a91620a <=( a91619a  and  a91616a );
 a91621a <=( a91620a  and  a91613a );
 a91624a <=( (not A266)  and  A265 );
 a91627a <=( (not A268)  and  (not A267) );
 a91628a <=( a91627a  and  a91624a );
 a91631a <=( A300  and  A269 );
 a91634a <=( A302  and  (not A301) );
 a91635a <=( a91634a  and  a91631a );
 a91636a <=( a91635a  and  a91628a );
 a91640a <=( (not A168)  and  (not A169) );
 a91641a <=( (not A170)  and  a91640a );
 a91644a <=( (not A166)  and  A167 );
 a91647a <=( (not A200)  and  (not A199) );
 a91648a <=( a91647a  and  a91644a );
 a91649a <=( a91648a  and  a91641a );
 a91652a <=( (not A268)  and  A267 );
 a91655a <=( A298  and  A269 );
 a91656a <=( a91655a  and  a91652a );
 a91659a <=( (not A300)  and  (not A299) );
 a91662a <=( A302  and  (not A301) );
 a91663a <=( a91662a  and  a91659a );
 a91664a <=( a91663a  and  a91656a );
 a91668a <=( (not A168)  and  (not A169) );
 a91669a <=( (not A170)  and  a91668a );
 a91672a <=( (not A166)  and  A167 );
 a91675a <=( (not A200)  and  (not A199) );
 a91676a <=( a91675a  and  a91672a );
 a91677a <=( a91676a  and  a91669a );
 a91680a <=( (not A268)  and  A267 );
 a91683a <=( (not A298)  and  A269 );
 a91684a <=( a91683a  and  a91680a );
 a91687a <=( (not A300)  and  A299 );
 a91690a <=( A302  and  (not A301) );
 a91691a <=( a91690a  and  a91687a );
 a91692a <=( a91691a  and  a91684a );
 a91696a <=( (not A168)  and  (not A169) );
 a91697a <=( (not A170)  and  a91696a );
 a91700a <=( (not A166)  and  A167 );
 a91703a <=( (not A200)  and  (not A199) );
 a91704a <=( a91703a  and  a91700a );
 a91705a <=( a91704a  and  a91697a );
 a91708a <=( A266  and  (not A265) );
 a91711a <=( (not A268)  and  (not A267) );
 a91712a <=( a91711a  and  a91708a );
 a91715a <=( A300  and  A269 );
 a91718a <=( A302  and  (not A301) );
 a91719a <=( a91718a  and  a91715a );
 a91720a <=( a91719a  and  a91712a );
 a91724a <=( (not A168)  and  (not A169) );
 a91725a <=( (not A170)  and  a91724a );
 a91728a <=( (not A166)  and  A167 );
 a91731a <=( (not A200)  and  (not A199) );
 a91732a <=( a91731a  and  a91728a );
 a91733a <=( a91732a  and  a91725a );
 a91736a <=( (not A266)  and  A265 );
 a91739a <=( (not A268)  and  (not A267) );
 a91740a <=( a91739a  and  a91736a );
 a91743a <=( A300  and  A269 );
 a91746a <=( A302  and  (not A301) );
 a91747a <=( a91746a  and  a91743a );
 a91748a <=( a91747a  and  a91740a );
 a91752a <=( (not A168)  and  (not A169) );
 a91753a <=( (not A170)  and  a91752a );
 a91756a <=( A166  and  (not A167) );
 a91759a <=( (not A202)  and  A201 );
 a91760a <=( a91759a  and  a91756a );
 a91761a <=( a91760a  and  a91753a );
 a91764a <=( A267  and  A203 );
 a91767a <=( A269  and  (not A268) );
 a91768a <=( a91767a  and  a91764a );
 a91771a <=( (not A299)  and  A298 );
 a91774a <=( A301  and  A300 );
 a91775a <=( a91774a  and  a91771a );
 a91776a <=( a91775a  and  a91768a );
 a91780a <=( (not A168)  and  (not A169) );
 a91781a <=( (not A170)  and  a91780a );
 a91784a <=( A166  and  (not A167) );
 a91787a <=( (not A202)  and  A201 );
 a91788a <=( a91787a  and  a91784a );
 a91789a <=( a91788a  and  a91781a );
 a91792a <=( A267  and  A203 );
 a91795a <=( A269  and  (not A268) );
 a91796a <=( a91795a  and  a91792a );
 a91799a <=( (not A299)  and  A298 );
 a91802a <=( (not A302)  and  A300 );
 a91803a <=( a91802a  and  a91799a );
 a91804a <=( a91803a  and  a91796a );
 a91808a <=( (not A168)  and  (not A169) );
 a91809a <=( (not A170)  and  a91808a );
 a91812a <=( A166  and  (not A167) );
 a91815a <=( (not A202)  and  A201 );
 a91816a <=( a91815a  and  a91812a );
 a91817a <=( a91816a  and  a91809a );
 a91820a <=( A267  and  A203 );
 a91823a <=( A269  and  (not A268) );
 a91824a <=( a91823a  and  a91820a );
 a91827a <=( A299  and  (not A298) );
 a91830a <=( A301  and  A300 );
 a91831a <=( a91830a  and  a91827a );
 a91832a <=( a91831a  and  a91824a );
 a91836a <=( (not A168)  and  (not A169) );
 a91837a <=( (not A170)  and  a91836a );
 a91840a <=( A166  and  (not A167) );
 a91843a <=( (not A202)  and  A201 );
 a91844a <=( a91843a  and  a91840a );
 a91845a <=( a91844a  and  a91837a );
 a91848a <=( A267  and  A203 );
 a91851a <=( A269  and  (not A268) );
 a91852a <=( a91851a  and  a91848a );
 a91855a <=( A299  and  (not A298) );
 a91858a <=( (not A302)  and  A300 );
 a91859a <=( a91858a  and  a91855a );
 a91860a <=( a91859a  and  a91852a );
 a91864a <=( (not A168)  and  (not A169) );
 a91865a <=( (not A170)  and  a91864a );
 a91868a <=( A166  and  (not A167) );
 a91871a <=( (not A202)  and  A201 );
 a91872a <=( a91871a  and  a91868a );
 a91873a <=( a91872a  and  a91865a );
 a91876a <=( (not A267)  and  A203 );
 a91879a <=( A298  and  A268 );
 a91880a <=( a91879a  and  a91876a );
 a91883a <=( (not A300)  and  (not A299) );
 a91886a <=( A302  and  (not A301) );
 a91887a <=( a91886a  and  a91883a );
 a91888a <=( a91887a  and  a91880a );
 a91892a <=( (not A168)  and  (not A169) );
 a91893a <=( (not A170)  and  a91892a );
 a91896a <=( A166  and  (not A167) );
 a91899a <=( (not A202)  and  A201 );
 a91900a <=( a91899a  and  a91896a );
 a91901a <=( a91900a  and  a91893a );
 a91904a <=( (not A267)  and  A203 );
 a91907a <=( (not A298)  and  A268 );
 a91908a <=( a91907a  and  a91904a );
 a91911a <=( (not A300)  and  A299 );
 a91914a <=( A302  and  (not A301) );
 a91915a <=( a91914a  and  a91911a );
 a91916a <=( a91915a  and  a91908a );
 a91920a <=( (not A168)  and  (not A169) );
 a91921a <=( (not A170)  and  a91920a );
 a91924a <=( A166  and  (not A167) );
 a91927a <=( (not A202)  and  A201 );
 a91928a <=( a91927a  and  a91924a );
 a91929a <=( a91928a  and  a91921a );
 a91932a <=( (not A267)  and  A203 );
 a91935a <=( A298  and  (not A269) );
 a91936a <=( a91935a  and  a91932a );
 a91939a <=( (not A300)  and  (not A299) );
 a91942a <=( A302  and  (not A301) );
 a91943a <=( a91942a  and  a91939a );
 a91944a <=( a91943a  and  a91936a );
 a91948a <=( (not A168)  and  (not A169) );
 a91949a <=( (not A170)  and  a91948a );
 a91952a <=( A166  and  (not A167) );
 a91955a <=( (not A202)  and  A201 );
 a91956a <=( a91955a  and  a91952a );
 a91957a <=( a91956a  and  a91949a );
 a91960a <=( (not A267)  and  A203 );
 a91963a <=( (not A298)  and  (not A269) );
 a91964a <=( a91963a  and  a91960a );
 a91967a <=( (not A300)  and  A299 );
 a91970a <=( A302  and  (not A301) );
 a91971a <=( a91970a  and  a91967a );
 a91972a <=( a91971a  and  a91964a );
 a91976a <=( (not A168)  and  (not A169) );
 a91977a <=( (not A170)  and  a91976a );
 a91980a <=( A166  and  (not A167) );
 a91983a <=( (not A202)  and  A201 );
 a91984a <=( a91983a  and  a91980a );
 a91985a <=( a91984a  and  a91977a );
 a91988a <=( A265  and  A203 );
 a91991a <=( A298  and  A266 );
 a91992a <=( a91991a  and  a91988a );
 a91995a <=( (not A300)  and  (not A299) );
 a91998a <=( A302  and  (not A301) );
 a91999a <=( a91998a  and  a91995a );
 a92000a <=( a91999a  and  a91992a );
 a92004a <=( (not A168)  and  (not A169) );
 a92005a <=( (not A170)  and  a92004a );
 a92008a <=( A166  and  (not A167) );
 a92011a <=( (not A202)  and  A201 );
 a92012a <=( a92011a  and  a92008a );
 a92013a <=( a92012a  and  a92005a );
 a92016a <=( A265  and  A203 );
 a92019a <=( (not A298)  and  A266 );
 a92020a <=( a92019a  and  a92016a );
 a92023a <=( (not A300)  and  A299 );
 a92026a <=( A302  and  (not A301) );
 a92027a <=( a92026a  and  a92023a );
 a92028a <=( a92027a  and  a92020a );
 a92032a <=( (not A168)  and  (not A169) );
 a92033a <=( (not A170)  and  a92032a );
 a92036a <=( A166  and  (not A167) );
 a92039a <=( (not A202)  and  A201 );
 a92040a <=( a92039a  and  a92036a );
 a92041a <=( a92040a  and  a92033a );
 a92044a <=( (not A265)  and  A203 );
 a92047a <=( A267  and  A266 );
 a92048a <=( a92047a  and  a92044a );
 a92051a <=( A300  and  A268 );
 a92054a <=( A302  and  (not A301) );
 a92055a <=( a92054a  and  a92051a );
 a92056a <=( a92055a  and  a92048a );
 a92060a <=( (not A168)  and  (not A169) );
 a92061a <=( (not A170)  and  a92060a );
 a92064a <=( A166  and  (not A167) );
 a92067a <=( (not A202)  and  A201 );
 a92068a <=( a92067a  and  a92064a );
 a92069a <=( a92068a  and  a92061a );
 a92072a <=( (not A265)  and  A203 );
 a92075a <=( A267  and  A266 );
 a92076a <=( a92075a  and  a92072a );
 a92079a <=( A300  and  (not A269) );
 a92082a <=( A302  and  (not A301) );
 a92083a <=( a92082a  and  a92079a );
 a92084a <=( a92083a  and  a92076a );
 a92088a <=( (not A168)  and  (not A169) );
 a92089a <=( (not A170)  and  a92088a );
 a92092a <=( A166  and  (not A167) );
 a92095a <=( (not A202)  and  A201 );
 a92096a <=( a92095a  and  a92092a );
 a92097a <=( a92096a  and  a92089a );
 a92100a <=( (not A265)  and  A203 );
 a92103a <=( (not A267)  and  A266 );
 a92104a <=( a92103a  and  a92100a );
 a92107a <=( A269  and  (not A268) );
 a92110a <=( A301  and  (not A300) );
 a92111a <=( a92110a  and  a92107a );
 a92112a <=( a92111a  and  a92104a );
 a92116a <=( (not A168)  and  (not A169) );
 a92117a <=( (not A170)  and  a92116a );
 a92120a <=( A166  and  (not A167) );
 a92123a <=( (not A202)  and  A201 );
 a92124a <=( a92123a  and  a92120a );
 a92125a <=( a92124a  and  a92117a );
 a92128a <=( (not A265)  and  A203 );
 a92131a <=( (not A267)  and  A266 );
 a92132a <=( a92131a  and  a92128a );
 a92135a <=( A269  and  (not A268) );
 a92138a <=( (not A302)  and  (not A300) );
 a92139a <=( a92138a  and  a92135a );
 a92140a <=( a92139a  and  a92132a );
 a92144a <=( (not A168)  and  (not A169) );
 a92145a <=( (not A170)  and  a92144a );
 a92148a <=( A166  and  (not A167) );
 a92151a <=( (not A202)  and  A201 );
 a92152a <=( a92151a  and  a92148a );
 a92153a <=( a92152a  and  a92145a );
 a92156a <=( (not A265)  and  A203 );
 a92159a <=( (not A267)  and  A266 );
 a92160a <=( a92159a  and  a92156a );
 a92163a <=( A269  and  (not A268) );
 a92166a <=( A299  and  A298 );
 a92167a <=( a92166a  and  a92163a );
 a92168a <=( a92167a  and  a92160a );
 a92172a <=( (not A168)  and  (not A169) );
 a92173a <=( (not A170)  and  a92172a );
 a92176a <=( A166  and  (not A167) );
 a92179a <=( (not A202)  and  A201 );
 a92180a <=( a92179a  and  a92176a );
 a92181a <=( a92180a  and  a92173a );
 a92184a <=( (not A265)  and  A203 );
 a92187a <=( (not A267)  and  A266 );
 a92188a <=( a92187a  and  a92184a );
 a92191a <=( A269  and  (not A268) );
 a92194a <=( (not A299)  and  (not A298) );
 a92195a <=( a92194a  and  a92191a );
 a92196a <=( a92195a  and  a92188a );
 a92200a <=( (not A168)  and  (not A169) );
 a92201a <=( (not A170)  and  a92200a );
 a92204a <=( A166  and  (not A167) );
 a92207a <=( (not A202)  and  A201 );
 a92208a <=( a92207a  and  a92204a );
 a92209a <=( a92208a  and  a92201a );
 a92212a <=( A265  and  A203 );
 a92215a <=( A267  and  (not A266) );
 a92216a <=( a92215a  and  a92212a );
 a92219a <=( A300  and  A268 );
 a92222a <=( A302  and  (not A301) );
 a92223a <=( a92222a  and  a92219a );
 a92224a <=( a92223a  and  a92216a );
 a92228a <=( (not A168)  and  (not A169) );
 a92229a <=( (not A170)  and  a92228a );
 a92232a <=( A166  and  (not A167) );
 a92235a <=( (not A202)  and  A201 );
 a92236a <=( a92235a  and  a92232a );
 a92237a <=( a92236a  and  a92229a );
 a92240a <=( A265  and  A203 );
 a92243a <=( A267  and  (not A266) );
 a92244a <=( a92243a  and  a92240a );
 a92247a <=( A300  and  (not A269) );
 a92250a <=( A302  and  (not A301) );
 a92251a <=( a92250a  and  a92247a );
 a92252a <=( a92251a  and  a92244a );
 a92256a <=( (not A168)  and  (not A169) );
 a92257a <=( (not A170)  and  a92256a );
 a92260a <=( A166  and  (not A167) );
 a92263a <=( (not A202)  and  A201 );
 a92264a <=( a92263a  and  a92260a );
 a92265a <=( a92264a  and  a92257a );
 a92268a <=( A265  and  A203 );
 a92271a <=( (not A267)  and  (not A266) );
 a92272a <=( a92271a  and  a92268a );
 a92275a <=( A269  and  (not A268) );
 a92278a <=( A301  and  (not A300) );
 a92279a <=( a92278a  and  a92275a );
 a92280a <=( a92279a  and  a92272a );
 a92284a <=( (not A168)  and  (not A169) );
 a92285a <=( (not A170)  and  a92284a );
 a92288a <=( A166  and  (not A167) );
 a92291a <=( (not A202)  and  A201 );
 a92292a <=( a92291a  and  a92288a );
 a92293a <=( a92292a  and  a92285a );
 a92296a <=( A265  and  A203 );
 a92299a <=( (not A267)  and  (not A266) );
 a92300a <=( a92299a  and  a92296a );
 a92303a <=( A269  and  (not A268) );
 a92306a <=( (not A302)  and  (not A300) );
 a92307a <=( a92306a  and  a92303a );
 a92308a <=( a92307a  and  a92300a );
 a92312a <=( (not A168)  and  (not A169) );
 a92313a <=( (not A170)  and  a92312a );
 a92316a <=( A166  and  (not A167) );
 a92319a <=( (not A202)  and  A201 );
 a92320a <=( a92319a  and  a92316a );
 a92321a <=( a92320a  and  a92313a );
 a92324a <=( A265  and  A203 );
 a92327a <=( (not A267)  and  (not A266) );
 a92328a <=( a92327a  and  a92324a );
 a92331a <=( A269  and  (not A268) );
 a92334a <=( A299  and  A298 );
 a92335a <=( a92334a  and  a92331a );
 a92336a <=( a92335a  and  a92328a );
 a92340a <=( (not A168)  and  (not A169) );
 a92341a <=( (not A170)  and  a92340a );
 a92344a <=( A166  and  (not A167) );
 a92347a <=( (not A202)  and  A201 );
 a92348a <=( a92347a  and  a92344a );
 a92349a <=( a92348a  and  a92341a );
 a92352a <=( A265  and  A203 );
 a92355a <=( (not A267)  and  (not A266) );
 a92356a <=( a92355a  and  a92352a );
 a92359a <=( A269  and  (not A268) );
 a92362a <=( (not A299)  and  (not A298) );
 a92363a <=( a92362a  and  a92359a );
 a92364a <=( a92363a  and  a92356a );
 a92368a <=( (not A168)  and  (not A169) );
 a92369a <=( (not A170)  and  a92368a );
 a92372a <=( A166  and  (not A167) );
 a92375a <=( (not A202)  and  A201 );
 a92376a <=( a92375a  and  a92372a );
 a92377a <=( a92376a  and  a92369a );
 a92380a <=( (not A265)  and  A203 );
 a92383a <=( A298  and  (not A266) );
 a92384a <=( a92383a  and  a92380a );
 a92387a <=( (not A300)  and  (not A299) );
 a92390a <=( A302  and  (not A301) );
 a92391a <=( a92390a  and  a92387a );
 a92392a <=( a92391a  and  a92384a );
 a92396a <=( (not A168)  and  (not A169) );
 a92397a <=( (not A170)  and  a92396a );
 a92400a <=( A166  and  (not A167) );
 a92403a <=( (not A202)  and  A201 );
 a92404a <=( a92403a  and  a92400a );
 a92405a <=( a92404a  and  a92397a );
 a92408a <=( (not A265)  and  A203 );
 a92411a <=( (not A298)  and  (not A266) );
 a92412a <=( a92411a  and  a92408a );
 a92415a <=( (not A300)  and  A299 );
 a92418a <=( A302  and  (not A301) );
 a92419a <=( a92418a  and  a92415a );
 a92420a <=( a92419a  and  a92412a );
 a92424a <=( (not A168)  and  (not A169) );
 a92425a <=( (not A170)  and  a92424a );
 a92428a <=( A166  and  (not A167) );
 a92431a <=( A202  and  (not A201) );
 a92432a <=( a92431a  and  a92428a );
 a92433a <=( a92432a  and  a92425a );
 a92436a <=( (not A268)  and  A267 );
 a92439a <=( A298  and  A269 );
 a92440a <=( a92439a  and  a92436a );
 a92443a <=( (not A300)  and  (not A299) );
 a92446a <=( A302  and  (not A301) );
 a92447a <=( a92446a  and  a92443a );
 a92448a <=( a92447a  and  a92440a );
 a92452a <=( (not A168)  and  (not A169) );
 a92453a <=( (not A170)  and  a92452a );
 a92456a <=( A166  and  (not A167) );
 a92459a <=( A202  and  (not A201) );
 a92460a <=( a92459a  and  a92456a );
 a92461a <=( a92460a  and  a92453a );
 a92464a <=( (not A268)  and  A267 );
 a92467a <=( (not A298)  and  A269 );
 a92468a <=( a92467a  and  a92464a );
 a92471a <=( (not A300)  and  A299 );
 a92474a <=( A302  and  (not A301) );
 a92475a <=( a92474a  and  a92471a );
 a92476a <=( a92475a  and  a92468a );
 a92480a <=( (not A168)  and  (not A169) );
 a92481a <=( (not A170)  and  a92480a );
 a92484a <=( A166  and  (not A167) );
 a92487a <=( A202  and  (not A201) );
 a92488a <=( a92487a  and  a92484a );
 a92489a <=( a92488a  and  a92481a );
 a92492a <=( A266  and  (not A265) );
 a92495a <=( (not A268)  and  (not A267) );
 a92496a <=( a92495a  and  a92492a );
 a92499a <=( A300  and  A269 );
 a92502a <=( A302  and  (not A301) );
 a92503a <=( a92502a  and  a92499a );
 a92504a <=( a92503a  and  a92496a );
 a92508a <=( (not A168)  and  (not A169) );
 a92509a <=( (not A170)  and  a92508a );
 a92512a <=( A166  and  (not A167) );
 a92515a <=( A202  and  (not A201) );
 a92516a <=( a92515a  and  a92512a );
 a92517a <=( a92516a  and  a92509a );
 a92520a <=( (not A266)  and  A265 );
 a92523a <=( (not A268)  and  (not A267) );
 a92524a <=( a92523a  and  a92520a );
 a92527a <=( A300  and  A269 );
 a92530a <=( A302  and  (not A301) );
 a92531a <=( a92530a  and  a92527a );
 a92532a <=( a92531a  and  a92524a );
 a92536a <=( (not A168)  and  (not A169) );
 a92537a <=( (not A170)  and  a92536a );
 a92540a <=( A166  and  (not A167) );
 a92543a <=( (not A203)  and  (not A201) );
 a92544a <=( a92543a  and  a92540a );
 a92545a <=( a92544a  and  a92537a );
 a92548a <=( (not A268)  and  A267 );
 a92551a <=( A298  and  A269 );
 a92552a <=( a92551a  and  a92548a );
 a92555a <=( (not A300)  and  (not A299) );
 a92558a <=( A302  and  (not A301) );
 a92559a <=( a92558a  and  a92555a );
 a92560a <=( a92559a  and  a92552a );
 a92564a <=( (not A168)  and  (not A169) );
 a92565a <=( (not A170)  and  a92564a );
 a92568a <=( A166  and  (not A167) );
 a92571a <=( (not A203)  and  (not A201) );
 a92572a <=( a92571a  and  a92568a );
 a92573a <=( a92572a  and  a92565a );
 a92576a <=( (not A268)  and  A267 );
 a92579a <=( (not A298)  and  A269 );
 a92580a <=( a92579a  and  a92576a );
 a92583a <=( (not A300)  and  A299 );
 a92586a <=( A302  and  (not A301) );
 a92587a <=( a92586a  and  a92583a );
 a92588a <=( a92587a  and  a92580a );
 a92592a <=( (not A168)  and  (not A169) );
 a92593a <=( (not A170)  and  a92592a );
 a92596a <=( A166  and  (not A167) );
 a92599a <=( (not A203)  and  (not A201) );
 a92600a <=( a92599a  and  a92596a );
 a92601a <=( a92600a  and  a92593a );
 a92604a <=( A266  and  (not A265) );
 a92607a <=( (not A268)  and  (not A267) );
 a92608a <=( a92607a  and  a92604a );
 a92611a <=( A300  and  A269 );
 a92614a <=( A302  and  (not A301) );
 a92615a <=( a92614a  and  a92611a );
 a92616a <=( a92615a  and  a92608a );
 a92620a <=( (not A168)  and  (not A169) );
 a92621a <=( (not A170)  and  a92620a );
 a92624a <=( A166  and  (not A167) );
 a92627a <=( (not A203)  and  (not A201) );
 a92628a <=( a92627a  and  a92624a );
 a92629a <=( a92628a  and  a92621a );
 a92632a <=( (not A266)  and  A265 );
 a92635a <=( (not A268)  and  (not A267) );
 a92636a <=( a92635a  and  a92632a );
 a92639a <=( A300  and  A269 );
 a92642a <=( A302  and  (not A301) );
 a92643a <=( a92642a  and  a92639a );
 a92644a <=( a92643a  and  a92636a );
 a92648a <=( (not A168)  and  (not A169) );
 a92649a <=( (not A170)  and  a92648a );
 a92652a <=( A166  and  (not A167) );
 a92655a <=( A200  and  A199 );
 a92656a <=( a92655a  and  a92652a );
 a92657a <=( a92656a  and  a92649a );
 a92660a <=( (not A268)  and  A267 );
 a92663a <=( A298  and  A269 );
 a92664a <=( a92663a  and  a92660a );
 a92667a <=( (not A300)  and  (not A299) );
 a92670a <=( A302  and  (not A301) );
 a92671a <=( a92670a  and  a92667a );
 a92672a <=( a92671a  and  a92664a );
 a92676a <=( (not A168)  and  (not A169) );
 a92677a <=( (not A170)  and  a92676a );
 a92680a <=( A166  and  (not A167) );
 a92683a <=( A200  and  A199 );
 a92684a <=( a92683a  and  a92680a );
 a92685a <=( a92684a  and  a92677a );
 a92688a <=( (not A268)  and  A267 );
 a92691a <=( (not A298)  and  A269 );
 a92692a <=( a92691a  and  a92688a );
 a92695a <=( (not A300)  and  A299 );
 a92698a <=( A302  and  (not A301) );
 a92699a <=( a92698a  and  a92695a );
 a92700a <=( a92699a  and  a92692a );
 a92704a <=( (not A168)  and  (not A169) );
 a92705a <=( (not A170)  and  a92704a );
 a92708a <=( A166  and  (not A167) );
 a92711a <=( A200  and  A199 );
 a92712a <=( a92711a  and  a92708a );
 a92713a <=( a92712a  and  a92705a );
 a92716a <=( A266  and  (not A265) );
 a92719a <=( (not A268)  and  (not A267) );
 a92720a <=( a92719a  and  a92716a );
 a92723a <=( A300  and  A269 );
 a92726a <=( A302  and  (not A301) );
 a92727a <=( a92726a  and  a92723a );
 a92728a <=( a92727a  and  a92720a );
 a92732a <=( (not A168)  and  (not A169) );
 a92733a <=( (not A170)  and  a92732a );
 a92736a <=( A166  and  (not A167) );
 a92739a <=( A200  and  A199 );
 a92740a <=( a92739a  and  a92736a );
 a92741a <=( a92740a  and  a92733a );
 a92744a <=( (not A266)  and  A265 );
 a92747a <=( (not A268)  and  (not A267) );
 a92748a <=( a92747a  and  a92744a );
 a92751a <=( A300  and  A269 );
 a92754a <=( A302  and  (not A301) );
 a92755a <=( a92754a  and  a92751a );
 a92756a <=( a92755a  and  a92748a );
 a92760a <=( (not A168)  and  (not A169) );
 a92761a <=( (not A170)  and  a92760a );
 a92764a <=( A166  and  (not A167) );
 a92767a <=( (not A200)  and  (not A199) );
 a92768a <=( a92767a  and  a92764a );
 a92769a <=( a92768a  and  a92761a );
 a92772a <=( (not A268)  and  A267 );
 a92775a <=( A298  and  A269 );
 a92776a <=( a92775a  and  a92772a );
 a92779a <=( (not A300)  and  (not A299) );
 a92782a <=( A302  and  (not A301) );
 a92783a <=( a92782a  and  a92779a );
 a92784a <=( a92783a  and  a92776a );
 a92788a <=( (not A168)  and  (not A169) );
 a92789a <=( (not A170)  and  a92788a );
 a92792a <=( A166  and  (not A167) );
 a92795a <=( (not A200)  and  (not A199) );
 a92796a <=( a92795a  and  a92792a );
 a92797a <=( a92796a  and  a92789a );
 a92800a <=( (not A268)  and  A267 );
 a92803a <=( (not A298)  and  A269 );
 a92804a <=( a92803a  and  a92800a );
 a92807a <=( (not A300)  and  A299 );
 a92810a <=( A302  and  (not A301) );
 a92811a <=( a92810a  and  a92807a );
 a92812a <=( a92811a  and  a92804a );
 a92816a <=( (not A168)  and  (not A169) );
 a92817a <=( (not A170)  and  a92816a );
 a92820a <=( A166  and  (not A167) );
 a92823a <=( (not A200)  and  (not A199) );
 a92824a <=( a92823a  and  a92820a );
 a92825a <=( a92824a  and  a92817a );
 a92828a <=( A266  and  (not A265) );
 a92831a <=( (not A268)  and  (not A267) );
 a92832a <=( a92831a  and  a92828a );
 a92835a <=( A300  and  A269 );
 a92838a <=( A302  and  (not A301) );
 a92839a <=( a92838a  and  a92835a );
 a92840a <=( a92839a  and  a92832a );
 a92844a <=( (not A168)  and  (not A169) );
 a92845a <=( (not A170)  and  a92844a );
 a92848a <=( A166  and  (not A167) );
 a92851a <=( (not A200)  and  (not A199) );
 a92852a <=( a92851a  and  a92848a );
 a92853a <=( a92852a  and  a92845a );
 a92856a <=( (not A266)  and  A265 );
 a92859a <=( (not A268)  and  (not A267) );
 a92860a <=( a92859a  and  a92856a );
 a92863a <=( A300  and  A269 );
 a92866a <=( A302  and  (not A301) );
 a92867a <=( a92866a  and  a92863a );
 a92868a <=( a92867a  and  a92860a );
 a92871a <=( A166  and  A167 );
 a92874a <=( A200  and  (not A199) );
 a92875a <=( a92874a  and  a92871a );
 a92878a <=( A202  and  A201 );
 a92881a <=( A266  and  (not A265) );
 a92882a <=( a92881a  and  a92878a );
 a92883a <=( a92882a  and  a92875a );
 a92886a <=( (not A268)  and  (not A267) );
 a92889a <=( A298  and  A269 );
 a92890a <=( a92889a  and  a92886a );
 a92893a <=( (not A300)  and  (not A299) );
 a92896a <=( A302  and  (not A301) );
 a92897a <=( a92896a  and  a92893a );
 a92898a <=( a92897a  and  a92890a );
 a92901a <=( A166  and  A167 );
 a92904a <=( A200  and  (not A199) );
 a92905a <=( a92904a  and  a92901a );
 a92908a <=( A202  and  A201 );
 a92911a <=( A266  and  (not A265) );
 a92912a <=( a92911a  and  a92908a );
 a92913a <=( a92912a  and  a92905a );
 a92916a <=( (not A268)  and  (not A267) );
 a92919a <=( (not A298)  and  A269 );
 a92920a <=( a92919a  and  a92916a );
 a92923a <=( (not A300)  and  A299 );
 a92926a <=( A302  and  (not A301) );
 a92927a <=( a92926a  and  a92923a );
 a92928a <=( a92927a  and  a92920a );
 a92931a <=( A166  and  A167 );
 a92934a <=( A200  and  (not A199) );
 a92935a <=( a92934a  and  a92931a );
 a92938a <=( A202  and  A201 );
 a92941a <=( (not A266)  and  A265 );
 a92942a <=( a92941a  and  a92938a );
 a92943a <=( a92942a  and  a92935a );
 a92946a <=( (not A268)  and  (not A267) );
 a92949a <=( A298  and  A269 );
 a92950a <=( a92949a  and  a92946a );
 a92953a <=( (not A300)  and  (not A299) );
 a92956a <=( A302  and  (not A301) );
 a92957a <=( a92956a  and  a92953a );
 a92958a <=( a92957a  and  a92950a );
 a92961a <=( A166  and  A167 );
 a92964a <=( A200  and  (not A199) );
 a92965a <=( a92964a  and  a92961a );
 a92968a <=( A202  and  A201 );
 a92971a <=( (not A266)  and  A265 );
 a92972a <=( a92971a  and  a92968a );
 a92973a <=( a92972a  and  a92965a );
 a92976a <=( (not A268)  and  (not A267) );
 a92979a <=( (not A298)  and  A269 );
 a92980a <=( a92979a  and  a92976a );
 a92983a <=( (not A300)  and  A299 );
 a92986a <=( A302  and  (not A301) );
 a92987a <=( a92986a  and  a92983a );
 a92988a <=( a92987a  and  a92980a );
 a92991a <=( A166  and  A167 );
 a92994a <=( A200  and  (not A199) );
 a92995a <=( a92994a  and  a92991a );
 a92998a <=( (not A203)  and  A201 );
 a93001a <=( A266  and  (not A265) );
 a93002a <=( a93001a  and  a92998a );
 a93003a <=( a93002a  and  a92995a );
 a93006a <=( (not A268)  and  (not A267) );
 a93009a <=( A298  and  A269 );
 a93010a <=( a93009a  and  a93006a );
 a93013a <=( (not A300)  and  (not A299) );
 a93016a <=( A302  and  (not A301) );
 a93017a <=( a93016a  and  a93013a );
 a93018a <=( a93017a  and  a93010a );
 a93021a <=( A166  and  A167 );
 a93024a <=( A200  and  (not A199) );
 a93025a <=( a93024a  and  a93021a );
 a93028a <=( (not A203)  and  A201 );
 a93031a <=( A266  and  (not A265) );
 a93032a <=( a93031a  and  a93028a );
 a93033a <=( a93032a  and  a93025a );
 a93036a <=( (not A268)  and  (not A267) );
 a93039a <=( (not A298)  and  A269 );
 a93040a <=( a93039a  and  a93036a );
 a93043a <=( (not A300)  and  A299 );
 a93046a <=( A302  and  (not A301) );
 a93047a <=( a93046a  and  a93043a );
 a93048a <=( a93047a  and  a93040a );
 a93051a <=( A166  and  A167 );
 a93054a <=( A200  and  (not A199) );
 a93055a <=( a93054a  and  a93051a );
 a93058a <=( (not A203)  and  A201 );
 a93061a <=( (not A266)  and  A265 );
 a93062a <=( a93061a  and  a93058a );
 a93063a <=( a93062a  and  a93055a );
 a93066a <=( (not A268)  and  (not A267) );
 a93069a <=( A298  and  A269 );
 a93070a <=( a93069a  and  a93066a );
 a93073a <=( (not A300)  and  (not A299) );
 a93076a <=( A302  and  (not A301) );
 a93077a <=( a93076a  and  a93073a );
 a93078a <=( a93077a  and  a93070a );
 a93081a <=( A166  and  A167 );
 a93084a <=( A200  and  (not A199) );
 a93085a <=( a93084a  and  a93081a );
 a93088a <=( (not A203)  and  A201 );
 a93091a <=( (not A266)  and  A265 );
 a93092a <=( a93091a  and  a93088a );
 a93093a <=( a93092a  and  a93085a );
 a93096a <=( (not A268)  and  (not A267) );
 a93099a <=( (not A298)  and  A269 );
 a93100a <=( a93099a  and  a93096a );
 a93103a <=( (not A300)  and  A299 );
 a93106a <=( A302  and  (not A301) );
 a93107a <=( a93106a  and  a93103a );
 a93108a <=( a93107a  and  a93100a );
 a93111a <=( A166  and  A167 );
 a93114a <=( A200  and  (not A199) );
 a93115a <=( a93114a  and  a93111a );
 a93118a <=( (not A202)  and  (not A201) );
 a93121a <=( (not A265)  and  A203 );
 a93122a <=( a93121a  and  a93118a );
 a93123a <=( a93122a  and  a93115a );
 a93126a <=( A267  and  A266 );
 a93129a <=( A298  and  A268 );
 a93130a <=( a93129a  and  a93126a );
 a93133a <=( (not A300)  and  (not A299) );
 a93136a <=( A302  and  (not A301) );
 a93137a <=( a93136a  and  a93133a );
 a93138a <=( a93137a  and  a93130a );
 a93141a <=( A166  and  A167 );
 a93144a <=( A200  and  (not A199) );
 a93145a <=( a93144a  and  a93141a );
 a93148a <=( (not A202)  and  (not A201) );
 a93151a <=( (not A265)  and  A203 );
 a93152a <=( a93151a  and  a93148a );
 a93153a <=( a93152a  and  a93145a );
 a93156a <=( A267  and  A266 );
 a93159a <=( (not A298)  and  A268 );
 a93160a <=( a93159a  and  a93156a );
 a93163a <=( (not A300)  and  A299 );
 a93166a <=( A302  and  (not A301) );
 a93167a <=( a93166a  and  a93163a );
 a93168a <=( a93167a  and  a93160a );
 a93171a <=( A166  and  A167 );
 a93174a <=( A200  and  (not A199) );
 a93175a <=( a93174a  and  a93171a );
 a93178a <=( (not A202)  and  (not A201) );
 a93181a <=( (not A265)  and  A203 );
 a93182a <=( a93181a  and  a93178a );
 a93183a <=( a93182a  and  a93175a );
 a93186a <=( A267  and  A266 );
 a93189a <=( A298  and  (not A269) );
 a93190a <=( a93189a  and  a93186a );
 a93193a <=( (not A300)  and  (not A299) );
 a93196a <=( A302  and  (not A301) );
 a93197a <=( a93196a  and  a93193a );
 a93198a <=( a93197a  and  a93190a );
 a93201a <=( A166  and  A167 );
 a93204a <=( A200  and  (not A199) );
 a93205a <=( a93204a  and  a93201a );
 a93208a <=( (not A202)  and  (not A201) );
 a93211a <=( (not A265)  and  A203 );
 a93212a <=( a93211a  and  a93208a );
 a93213a <=( a93212a  and  a93205a );
 a93216a <=( A267  and  A266 );
 a93219a <=( (not A298)  and  (not A269) );
 a93220a <=( a93219a  and  a93216a );
 a93223a <=( (not A300)  and  A299 );
 a93226a <=( A302  and  (not A301) );
 a93227a <=( a93226a  and  a93223a );
 a93228a <=( a93227a  and  a93220a );
 a93231a <=( A166  and  A167 );
 a93234a <=( A200  and  (not A199) );
 a93235a <=( a93234a  and  a93231a );
 a93238a <=( (not A202)  and  (not A201) );
 a93241a <=( (not A265)  and  A203 );
 a93242a <=( a93241a  and  a93238a );
 a93243a <=( a93242a  and  a93235a );
 a93246a <=( (not A267)  and  A266 );
 a93249a <=( A269  and  (not A268) );
 a93250a <=( a93249a  and  a93246a );
 a93253a <=( (not A299)  and  A298 );
 a93256a <=( A301  and  A300 );
 a93257a <=( a93256a  and  a93253a );
 a93258a <=( a93257a  and  a93250a );
 a93261a <=( A166  and  A167 );
 a93264a <=( A200  and  (not A199) );
 a93265a <=( a93264a  and  a93261a );
 a93268a <=( (not A202)  and  (not A201) );
 a93271a <=( (not A265)  and  A203 );
 a93272a <=( a93271a  and  a93268a );
 a93273a <=( a93272a  and  a93265a );
 a93276a <=( (not A267)  and  A266 );
 a93279a <=( A269  and  (not A268) );
 a93280a <=( a93279a  and  a93276a );
 a93283a <=( (not A299)  and  A298 );
 a93286a <=( (not A302)  and  A300 );
 a93287a <=( a93286a  and  a93283a );
 a93288a <=( a93287a  and  a93280a );
 a93291a <=( A166  and  A167 );
 a93294a <=( A200  and  (not A199) );
 a93295a <=( a93294a  and  a93291a );
 a93298a <=( (not A202)  and  (not A201) );
 a93301a <=( (not A265)  and  A203 );
 a93302a <=( a93301a  and  a93298a );
 a93303a <=( a93302a  and  a93295a );
 a93306a <=( (not A267)  and  A266 );
 a93309a <=( A269  and  (not A268) );
 a93310a <=( a93309a  and  a93306a );
 a93313a <=( A299  and  (not A298) );
 a93316a <=( A301  and  A300 );
 a93317a <=( a93316a  and  a93313a );
 a93318a <=( a93317a  and  a93310a );
 a93321a <=( A166  and  A167 );
 a93324a <=( A200  and  (not A199) );
 a93325a <=( a93324a  and  a93321a );
 a93328a <=( (not A202)  and  (not A201) );
 a93331a <=( (not A265)  and  A203 );
 a93332a <=( a93331a  and  a93328a );
 a93333a <=( a93332a  and  a93325a );
 a93336a <=( (not A267)  and  A266 );
 a93339a <=( A269  and  (not A268) );
 a93340a <=( a93339a  and  a93336a );
 a93343a <=( A299  and  (not A298) );
 a93346a <=( (not A302)  and  A300 );
 a93347a <=( a93346a  and  a93343a );
 a93348a <=( a93347a  and  a93340a );
 a93351a <=( A166  and  A167 );
 a93354a <=( A200  and  (not A199) );
 a93355a <=( a93354a  and  a93351a );
 a93358a <=( (not A202)  and  (not A201) );
 a93361a <=( A265  and  A203 );
 a93362a <=( a93361a  and  a93358a );
 a93363a <=( a93362a  and  a93355a );
 a93366a <=( A267  and  (not A266) );
 a93369a <=( A298  and  A268 );
 a93370a <=( a93369a  and  a93366a );
 a93373a <=( (not A300)  and  (not A299) );
 a93376a <=( A302  and  (not A301) );
 a93377a <=( a93376a  and  a93373a );
 a93378a <=( a93377a  and  a93370a );
 a93381a <=( A166  and  A167 );
 a93384a <=( A200  and  (not A199) );
 a93385a <=( a93384a  and  a93381a );
 a93388a <=( (not A202)  and  (not A201) );
 a93391a <=( A265  and  A203 );
 a93392a <=( a93391a  and  a93388a );
 a93393a <=( a93392a  and  a93385a );
 a93396a <=( A267  and  (not A266) );
 a93399a <=( (not A298)  and  A268 );
 a93400a <=( a93399a  and  a93396a );
 a93403a <=( (not A300)  and  A299 );
 a93406a <=( A302  and  (not A301) );
 a93407a <=( a93406a  and  a93403a );
 a93408a <=( a93407a  and  a93400a );
 a93411a <=( A166  and  A167 );
 a93414a <=( A200  and  (not A199) );
 a93415a <=( a93414a  and  a93411a );
 a93418a <=( (not A202)  and  (not A201) );
 a93421a <=( A265  and  A203 );
 a93422a <=( a93421a  and  a93418a );
 a93423a <=( a93422a  and  a93415a );
 a93426a <=( A267  and  (not A266) );
 a93429a <=( A298  and  (not A269) );
 a93430a <=( a93429a  and  a93426a );
 a93433a <=( (not A300)  and  (not A299) );
 a93436a <=( A302  and  (not A301) );
 a93437a <=( a93436a  and  a93433a );
 a93438a <=( a93437a  and  a93430a );
 a93441a <=( A166  and  A167 );
 a93444a <=( A200  and  (not A199) );
 a93445a <=( a93444a  and  a93441a );
 a93448a <=( (not A202)  and  (not A201) );
 a93451a <=( A265  and  A203 );
 a93452a <=( a93451a  and  a93448a );
 a93453a <=( a93452a  and  a93445a );
 a93456a <=( A267  and  (not A266) );
 a93459a <=( (not A298)  and  (not A269) );
 a93460a <=( a93459a  and  a93456a );
 a93463a <=( (not A300)  and  A299 );
 a93466a <=( A302  and  (not A301) );
 a93467a <=( a93466a  and  a93463a );
 a93468a <=( a93467a  and  a93460a );
 a93471a <=( A166  and  A167 );
 a93474a <=( A200  and  (not A199) );
 a93475a <=( a93474a  and  a93471a );
 a93478a <=( (not A202)  and  (not A201) );
 a93481a <=( A265  and  A203 );
 a93482a <=( a93481a  and  a93478a );
 a93483a <=( a93482a  and  a93475a );
 a93486a <=( (not A267)  and  (not A266) );
 a93489a <=( A269  and  (not A268) );
 a93490a <=( a93489a  and  a93486a );
 a93493a <=( (not A299)  and  A298 );
 a93496a <=( A301  and  A300 );
 a93497a <=( a93496a  and  a93493a );
 a93498a <=( a93497a  and  a93490a );
 a93501a <=( A166  and  A167 );
 a93504a <=( A200  and  (not A199) );
 a93505a <=( a93504a  and  a93501a );
 a93508a <=( (not A202)  and  (not A201) );
 a93511a <=( A265  and  A203 );
 a93512a <=( a93511a  and  a93508a );
 a93513a <=( a93512a  and  a93505a );
 a93516a <=( (not A267)  and  (not A266) );
 a93519a <=( A269  and  (not A268) );
 a93520a <=( a93519a  and  a93516a );
 a93523a <=( (not A299)  and  A298 );
 a93526a <=( (not A302)  and  A300 );
 a93527a <=( a93526a  and  a93523a );
 a93528a <=( a93527a  and  a93520a );
 a93531a <=( A166  and  A167 );
 a93534a <=( A200  and  (not A199) );
 a93535a <=( a93534a  and  a93531a );
 a93538a <=( (not A202)  and  (not A201) );
 a93541a <=( A265  and  A203 );
 a93542a <=( a93541a  and  a93538a );
 a93543a <=( a93542a  and  a93535a );
 a93546a <=( (not A267)  and  (not A266) );
 a93549a <=( A269  and  (not A268) );
 a93550a <=( a93549a  and  a93546a );
 a93553a <=( A299  and  (not A298) );
 a93556a <=( A301  and  A300 );
 a93557a <=( a93556a  and  a93553a );
 a93558a <=( a93557a  and  a93550a );
 a93561a <=( A166  and  A167 );
 a93564a <=( A200  and  (not A199) );
 a93565a <=( a93564a  and  a93561a );
 a93568a <=( (not A202)  and  (not A201) );
 a93571a <=( A265  and  A203 );
 a93572a <=( a93571a  and  a93568a );
 a93573a <=( a93572a  and  a93565a );
 a93576a <=( (not A267)  and  (not A266) );
 a93579a <=( A269  and  (not A268) );
 a93580a <=( a93579a  and  a93576a );
 a93583a <=( A299  and  (not A298) );
 a93586a <=( (not A302)  and  A300 );
 a93587a <=( a93586a  and  a93583a );
 a93588a <=( a93587a  and  a93580a );
 a93591a <=( A166  and  A167 );
 a93594a <=( (not A200)  and  A199 );
 a93595a <=( a93594a  and  a93591a );
 a93598a <=( A202  and  A201 );
 a93601a <=( A266  and  (not A265) );
 a93602a <=( a93601a  and  a93598a );
 a93603a <=( a93602a  and  a93595a );
 a93606a <=( (not A268)  and  (not A267) );
 a93609a <=( A298  and  A269 );
 a93610a <=( a93609a  and  a93606a );
 a93613a <=( (not A300)  and  (not A299) );
 a93616a <=( A302  and  (not A301) );
 a93617a <=( a93616a  and  a93613a );
 a93618a <=( a93617a  and  a93610a );
 a93621a <=( A166  and  A167 );
 a93624a <=( (not A200)  and  A199 );
 a93625a <=( a93624a  and  a93621a );
 a93628a <=( A202  and  A201 );
 a93631a <=( A266  and  (not A265) );
 a93632a <=( a93631a  and  a93628a );
 a93633a <=( a93632a  and  a93625a );
 a93636a <=( (not A268)  and  (not A267) );
 a93639a <=( (not A298)  and  A269 );
 a93640a <=( a93639a  and  a93636a );
 a93643a <=( (not A300)  and  A299 );
 a93646a <=( A302  and  (not A301) );
 a93647a <=( a93646a  and  a93643a );
 a93648a <=( a93647a  and  a93640a );
 a93651a <=( A166  and  A167 );
 a93654a <=( (not A200)  and  A199 );
 a93655a <=( a93654a  and  a93651a );
 a93658a <=( A202  and  A201 );
 a93661a <=( (not A266)  and  A265 );
 a93662a <=( a93661a  and  a93658a );
 a93663a <=( a93662a  and  a93655a );
 a93666a <=( (not A268)  and  (not A267) );
 a93669a <=( A298  and  A269 );
 a93670a <=( a93669a  and  a93666a );
 a93673a <=( (not A300)  and  (not A299) );
 a93676a <=( A302  and  (not A301) );
 a93677a <=( a93676a  and  a93673a );
 a93678a <=( a93677a  and  a93670a );
 a93681a <=( A166  and  A167 );
 a93684a <=( (not A200)  and  A199 );
 a93685a <=( a93684a  and  a93681a );
 a93688a <=( A202  and  A201 );
 a93691a <=( (not A266)  and  A265 );
 a93692a <=( a93691a  and  a93688a );
 a93693a <=( a93692a  and  a93685a );
 a93696a <=( (not A268)  and  (not A267) );
 a93699a <=( (not A298)  and  A269 );
 a93700a <=( a93699a  and  a93696a );
 a93703a <=( (not A300)  and  A299 );
 a93706a <=( A302  and  (not A301) );
 a93707a <=( a93706a  and  a93703a );
 a93708a <=( a93707a  and  a93700a );
 a93711a <=( A166  and  A167 );
 a93714a <=( (not A200)  and  A199 );
 a93715a <=( a93714a  and  a93711a );
 a93718a <=( (not A203)  and  A201 );
 a93721a <=( A266  and  (not A265) );
 a93722a <=( a93721a  and  a93718a );
 a93723a <=( a93722a  and  a93715a );
 a93726a <=( (not A268)  and  (not A267) );
 a93729a <=( A298  and  A269 );
 a93730a <=( a93729a  and  a93726a );
 a93733a <=( (not A300)  and  (not A299) );
 a93736a <=( A302  and  (not A301) );
 a93737a <=( a93736a  and  a93733a );
 a93738a <=( a93737a  and  a93730a );
 a93741a <=( A166  and  A167 );
 a93744a <=( (not A200)  and  A199 );
 a93745a <=( a93744a  and  a93741a );
 a93748a <=( (not A203)  and  A201 );
 a93751a <=( A266  and  (not A265) );
 a93752a <=( a93751a  and  a93748a );
 a93753a <=( a93752a  and  a93745a );
 a93756a <=( (not A268)  and  (not A267) );
 a93759a <=( (not A298)  and  A269 );
 a93760a <=( a93759a  and  a93756a );
 a93763a <=( (not A300)  and  A299 );
 a93766a <=( A302  and  (not A301) );
 a93767a <=( a93766a  and  a93763a );
 a93768a <=( a93767a  and  a93760a );
 a93771a <=( A166  and  A167 );
 a93774a <=( (not A200)  and  A199 );
 a93775a <=( a93774a  and  a93771a );
 a93778a <=( (not A203)  and  A201 );
 a93781a <=( (not A266)  and  A265 );
 a93782a <=( a93781a  and  a93778a );
 a93783a <=( a93782a  and  a93775a );
 a93786a <=( (not A268)  and  (not A267) );
 a93789a <=( A298  and  A269 );
 a93790a <=( a93789a  and  a93786a );
 a93793a <=( (not A300)  and  (not A299) );
 a93796a <=( A302  and  (not A301) );
 a93797a <=( a93796a  and  a93793a );
 a93798a <=( a93797a  and  a93790a );
 a93801a <=( A166  and  A167 );
 a93804a <=( (not A200)  and  A199 );
 a93805a <=( a93804a  and  a93801a );
 a93808a <=( (not A203)  and  A201 );
 a93811a <=( (not A266)  and  A265 );
 a93812a <=( a93811a  and  a93808a );
 a93813a <=( a93812a  and  a93805a );
 a93816a <=( (not A268)  and  (not A267) );
 a93819a <=( (not A298)  and  A269 );
 a93820a <=( a93819a  and  a93816a );
 a93823a <=( (not A300)  and  A299 );
 a93826a <=( A302  and  (not A301) );
 a93827a <=( a93826a  and  a93823a );
 a93828a <=( a93827a  and  a93820a );
 a93831a <=( A166  and  A167 );
 a93834a <=( (not A200)  and  A199 );
 a93835a <=( a93834a  and  a93831a );
 a93838a <=( (not A202)  and  (not A201) );
 a93841a <=( (not A265)  and  A203 );
 a93842a <=( a93841a  and  a93838a );
 a93843a <=( a93842a  and  a93835a );
 a93846a <=( A267  and  A266 );
 a93849a <=( A298  and  A268 );
 a93850a <=( a93849a  and  a93846a );
 a93853a <=( (not A300)  and  (not A299) );
 a93856a <=( A302  and  (not A301) );
 a93857a <=( a93856a  and  a93853a );
 a93858a <=( a93857a  and  a93850a );
 a93861a <=( A166  and  A167 );
 a93864a <=( (not A200)  and  A199 );
 a93865a <=( a93864a  and  a93861a );
 a93868a <=( (not A202)  and  (not A201) );
 a93871a <=( (not A265)  and  A203 );
 a93872a <=( a93871a  and  a93868a );
 a93873a <=( a93872a  and  a93865a );
 a93876a <=( A267  and  A266 );
 a93879a <=( (not A298)  and  A268 );
 a93880a <=( a93879a  and  a93876a );
 a93883a <=( (not A300)  and  A299 );
 a93886a <=( A302  and  (not A301) );
 a93887a <=( a93886a  and  a93883a );
 a93888a <=( a93887a  and  a93880a );
 a93891a <=( A166  and  A167 );
 a93894a <=( (not A200)  and  A199 );
 a93895a <=( a93894a  and  a93891a );
 a93898a <=( (not A202)  and  (not A201) );
 a93901a <=( (not A265)  and  A203 );
 a93902a <=( a93901a  and  a93898a );
 a93903a <=( a93902a  and  a93895a );
 a93906a <=( A267  and  A266 );
 a93909a <=( A298  and  (not A269) );
 a93910a <=( a93909a  and  a93906a );
 a93913a <=( (not A300)  and  (not A299) );
 a93916a <=( A302  and  (not A301) );
 a93917a <=( a93916a  and  a93913a );
 a93918a <=( a93917a  and  a93910a );
 a93921a <=( A166  and  A167 );
 a93924a <=( (not A200)  and  A199 );
 a93925a <=( a93924a  and  a93921a );
 a93928a <=( (not A202)  and  (not A201) );
 a93931a <=( (not A265)  and  A203 );
 a93932a <=( a93931a  and  a93928a );
 a93933a <=( a93932a  and  a93925a );
 a93936a <=( A267  and  A266 );
 a93939a <=( (not A298)  and  (not A269) );
 a93940a <=( a93939a  and  a93936a );
 a93943a <=( (not A300)  and  A299 );
 a93946a <=( A302  and  (not A301) );
 a93947a <=( a93946a  and  a93943a );
 a93948a <=( a93947a  and  a93940a );
 a93951a <=( A166  and  A167 );
 a93954a <=( (not A200)  and  A199 );
 a93955a <=( a93954a  and  a93951a );
 a93958a <=( (not A202)  and  (not A201) );
 a93961a <=( (not A265)  and  A203 );
 a93962a <=( a93961a  and  a93958a );
 a93963a <=( a93962a  and  a93955a );
 a93966a <=( (not A267)  and  A266 );
 a93969a <=( A269  and  (not A268) );
 a93970a <=( a93969a  and  a93966a );
 a93973a <=( (not A299)  and  A298 );
 a93976a <=( A301  and  A300 );
 a93977a <=( a93976a  and  a93973a );
 a93978a <=( a93977a  and  a93970a );
 a93981a <=( A166  and  A167 );
 a93984a <=( (not A200)  and  A199 );
 a93985a <=( a93984a  and  a93981a );
 a93988a <=( (not A202)  and  (not A201) );
 a93991a <=( (not A265)  and  A203 );
 a93992a <=( a93991a  and  a93988a );
 a93993a <=( a93992a  and  a93985a );
 a93996a <=( (not A267)  and  A266 );
 a93999a <=( A269  and  (not A268) );
 a94000a <=( a93999a  and  a93996a );
 a94003a <=( (not A299)  and  A298 );
 a94006a <=( (not A302)  and  A300 );
 a94007a <=( a94006a  and  a94003a );
 a94008a <=( a94007a  and  a94000a );
 a94011a <=( A166  and  A167 );
 a94014a <=( (not A200)  and  A199 );
 a94015a <=( a94014a  and  a94011a );
 a94018a <=( (not A202)  and  (not A201) );
 a94021a <=( (not A265)  and  A203 );
 a94022a <=( a94021a  and  a94018a );
 a94023a <=( a94022a  and  a94015a );
 a94026a <=( (not A267)  and  A266 );
 a94029a <=( A269  and  (not A268) );
 a94030a <=( a94029a  and  a94026a );
 a94033a <=( A299  and  (not A298) );
 a94036a <=( A301  and  A300 );
 a94037a <=( a94036a  and  a94033a );
 a94038a <=( a94037a  and  a94030a );
 a94041a <=( A166  and  A167 );
 a94044a <=( (not A200)  and  A199 );
 a94045a <=( a94044a  and  a94041a );
 a94048a <=( (not A202)  and  (not A201) );
 a94051a <=( (not A265)  and  A203 );
 a94052a <=( a94051a  and  a94048a );
 a94053a <=( a94052a  and  a94045a );
 a94056a <=( (not A267)  and  A266 );
 a94059a <=( A269  and  (not A268) );
 a94060a <=( a94059a  and  a94056a );
 a94063a <=( A299  and  (not A298) );
 a94066a <=( (not A302)  and  A300 );
 a94067a <=( a94066a  and  a94063a );
 a94068a <=( a94067a  and  a94060a );
 a94071a <=( A166  and  A167 );
 a94074a <=( (not A200)  and  A199 );
 a94075a <=( a94074a  and  a94071a );
 a94078a <=( (not A202)  and  (not A201) );
 a94081a <=( A265  and  A203 );
 a94082a <=( a94081a  and  a94078a );
 a94083a <=( a94082a  and  a94075a );
 a94086a <=( A267  and  (not A266) );
 a94089a <=( A298  and  A268 );
 a94090a <=( a94089a  and  a94086a );
 a94093a <=( (not A300)  and  (not A299) );
 a94096a <=( A302  and  (not A301) );
 a94097a <=( a94096a  and  a94093a );
 a94098a <=( a94097a  and  a94090a );
 a94101a <=( A166  and  A167 );
 a94104a <=( (not A200)  and  A199 );
 a94105a <=( a94104a  and  a94101a );
 a94108a <=( (not A202)  and  (not A201) );
 a94111a <=( A265  and  A203 );
 a94112a <=( a94111a  and  a94108a );
 a94113a <=( a94112a  and  a94105a );
 a94116a <=( A267  and  (not A266) );
 a94119a <=( (not A298)  and  A268 );
 a94120a <=( a94119a  and  a94116a );
 a94123a <=( (not A300)  and  A299 );
 a94126a <=( A302  and  (not A301) );
 a94127a <=( a94126a  and  a94123a );
 a94128a <=( a94127a  and  a94120a );
 a94131a <=( A166  and  A167 );
 a94134a <=( (not A200)  and  A199 );
 a94135a <=( a94134a  and  a94131a );
 a94138a <=( (not A202)  and  (not A201) );
 a94141a <=( A265  and  A203 );
 a94142a <=( a94141a  and  a94138a );
 a94143a <=( a94142a  and  a94135a );
 a94146a <=( A267  and  (not A266) );
 a94149a <=( A298  and  (not A269) );
 a94150a <=( a94149a  and  a94146a );
 a94153a <=( (not A300)  and  (not A299) );
 a94156a <=( A302  and  (not A301) );
 a94157a <=( a94156a  and  a94153a );
 a94158a <=( a94157a  and  a94150a );
 a94161a <=( A166  and  A167 );
 a94164a <=( (not A200)  and  A199 );
 a94165a <=( a94164a  and  a94161a );
 a94168a <=( (not A202)  and  (not A201) );
 a94171a <=( A265  and  A203 );
 a94172a <=( a94171a  and  a94168a );
 a94173a <=( a94172a  and  a94165a );
 a94176a <=( A267  and  (not A266) );
 a94179a <=( (not A298)  and  (not A269) );
 a94180a <=( a94179a  and  a94176a );
 a94183a <=( (not A300)  and  A299 );
 a94186a <=( A302  and  (not A301) );
 a94187a <=( a94186a  and  a94183a );
 a94188a <=( a94187a  and  a94180a );
 a94191a <=( A166  and  A167 );
 a94194a <=( (not A200)  and  A199 );
 a94195a <=( a94194a  and  a94191a );
 a94198a <=( (not A202)  and  (not A201) );
 a94201a <=( A265  and  A203 );
 a94202a <=( a94201a  and  a94198a );
 a94203a <=( a94202a  and  a94195a );
 a94206a <=( (not A267)  and  (not A266) );
 a94209a <=( A269  and  (not A268) );
 a94210a <=( a94209a  and  a94206a );
 a94213a <=( (not A299)  and  A298 );
 a94216a <=( A301  and  A300 );
 a94217a <=( a94216a  and  a94213a );
 a94218a <=( a94217a  and  a94210a );
 a94221a <=( A166  and  A167 );
 a94224a <=( (not A200)  and  A199 );
 a94225a <=( a94224a  and  a94221a );
 a94228a <=( (not A202)  and  (not A201) );
 a94231a <=( A265  and  A203 );
 a94232a <=( a94231a  and  a94228a );
 a94233a <=( a94232a  and  a94225a );
 a94236a <=( (not A267)  and  (not A266) );
 a94239a <=( A269  and  (not A268) );
 a94240a <=( a94239a  and  a94236a );
 a94243a <=( (not A299)  and  A298 );
 a94246a <=( (not A302)  and  A300 );
 a94247a <=( a94246a  and  a94243a );
 a94248a <=( a94247a  and  a94240a );
 a94251a <=( A166  and  A167 );
 a94254a <=( (not A200)  and  A199 );
 a94255a <=( a94254a  and  a94251a );
 a94258a <=( (not A202)  and  (not A201) );
 a94261a <=( A265  and  A203 );
 a94262a <=( a94261a  and  a94258a );
 a94263a <=( a94262a  and  a94255a );
 a94266a <=( (not A267)  and  (not A266) );
 a94269a <=( A269  and  (not A268) );
 a94270a <=( a94269a  and  a94266a );
 a94273a <=( A299  and  (not A298) );
 a94276a <=( A301  and  A300 );
 a94277a <=( a94276a  and  a94273a );
 a94278a <=( a94277a  and  a94270a );
 a94281a <=( A166  and  A167 );
 a94284a <=( (not A200)  and  A199 );
 a94285a <=( a94284a  and  a94281a );
 a94288a <=( (not A202)  and  (not A201) );
 a94291a <=( A265  and  A203 );
 a94292a <=( a94291a  and  a94288a );
 a94293a <=( a94292a  and  a94285a );
 a94296a <=( (not A267)  and  (not A266) );
 a94299a <=( A269  and  (not A268) );
 a94300a <=( a94299a  and  a94296a );
 a94303a <=( A299  and  (not A298) );
 a94306a <=( (not A302)  and  A300 );
 a94307a <=( a94306a  and  a94303a );
 a94308a <=( a94307a  and  a94300a );
 a94311a <=( (not A166)  and  (not A167) );
 a94314a <=( A200  and  (not A199) );
 a94315a <=( a94314a  and  a94311a );
 a94318a <=( A202  and  A201 );
 a94321a <=( A266  and  (not A265) );
 a94322a <=( a94321a  and  a94318a );
 a94323a <=( a94322a  and  a94315a );
 a94326a <=( (not A268)  and  (not A267) );
 a94329a <=( A298  and  A269 );
 a94330a <=( a94329a  and  a94326a );
 a94333a <=( (not A300)  and  (not A299) );
 a94336a <=( A302  and  (not A301) );
 a94337a <=( a94336a  and  a94333a );
 a94338a <=( a94337a  and  a94330a );
 a94341a <=( (not A166)  and  (not A167) );
 a94344a <=( A200  and  (not A199) );
 a94345a <=( a94344a  and  a94341a );
 a94348a <=( A202  and  A201 );
 a94351a <=( A266  and  (not A265) );
 a94352a <=( a94351a  and  a94348a );
 a94353a <=( a94352a  and  a94345a );
 a94356a <=( (not A268)  and  (not A267) );
 a94359a <=( (not A298)  and  A269 );
 a94360a <=( a94359a  and  a94356a );
 a94363a <=( (not A300)  and  A299 );
 a94366a <=( A302  and  (not A301) );
 a94367a <=( a94366a  and  a94363a );
 a94368a <=( a94367a  and  a94360a );
 a94371a <=( (not A166)  and  (not A167) );
 a94374a <=( A200  and  (not A199) );
 a94375a <=( a94374a  and  a94371a );
 a94378a <=( A202  and  A201 );
 a94381a <=( (not A266)  and  A265 );
 a94382a <=( a94381a  and  a94378a );
 a94383a <=( a94382a  and  a94375a );
 a94386a <=( (not A268)  and  (not A267) );
 a94389a <=( A298  and  A269 );
 a94390a <=( a94389a  and  a94386a );
 a94393a <=( (not A300)  and  (not A299) );
 a94396a <=( A302  and  (not A301) );
 a94397a <=( a94396a  and  a94393a );
 a94398a <=( a94397a  and  a94390a );
 a94401a <=( (not A166)  and  (not A167) );
 a94404a <=( A200  and  (not A199) );
 a94405a <=( a94404a  and  a94401a );
 a94408a <=( A202  and  A201 );
 a94411a <=( (not A266)  and  A265 );
 a94412a <=( a94411a  and  a94408a );
 a94413a <=( a94412a  and  a94405a );
 a94416a <=( (not A268)  and  (not A267) );
 a94419a <=( (not A298)  and  A269 );
 a94420a <=( a94419a  and  a94416a );
 a94423a <=( (not A300)  and  A299 );
 a94426a <=( A302  and  (not A301) );
 a94427a <=( a94426a  and  a94423a );
 a94428a <=( a94427a  and  a94420a );
 a94431a <=( (not A166)  and  (not A167) );
 a94434a <=( A200  and  (not A199) );
 a94435a <=( a94434a  and  a94431a );
 a94438a <=( (not A203)  and  A201 );
 a94441a <=( A266  and  (not A265) );
 a94442a <=( a94441a  and  a94438a );
 a94443a <=( a94442a  and  a94435a );
 a94446a <=( (not A268)  and  (not A267) );
 a94449a <=( A298  and  A269 );
 a94450a <=( a94449a  and  a94446a );
 a94453a <=( (not A300)  and  (not A299) );
 a94456a <=( A302  and  (not A301) );
 a94457a <=( a94456a  and  a94453a );
 a94458a <=( a94457a  and  a94450a );
 a94461a <=( (not A166)  and  (not A167) );
 a94464a <=( A200  and  (not A199) );
 a94465a <=( a94464a  and  a94461a );
 a94468a <=( (not A203)  and  A201 );
 a94471a <=( A266  and  (not A265) );
 a94472a <=( a94471a  and  a94468a );
 a94473a <=( a94472a  and  a94465a );
 a94476a <=( (not A268)  and  (not A267) );
 a94479a <=( (not A298)  and  A269 );
 a94480a <=( a94479a  and  a94476a );
 a94483a <=( (not A300)  and  A299 );
 a94486a <=( A302  and  (not A301) );
 a94487a <=( a94486a  and  a94483a );
 a94488a <=( a94487a  and  a94480a );
 a94491a <=( (not A166)  and  (not A167) );
 a94494a <=( A200  and  (not A199) );
 a94495a <=( a94494a  and  a94491a );
 a94498a <=( (not A203)  and  A201 );
 a94501a <=( (not A266)  and  A265 );
 a94502a <=( a94501a  and  a94498a );
 a94503a <=( a94502a  and  a94495a );
 a94506a <=( (not A268)  and  (not A267) );
 a94509a <=( A298  and  A269 );
 a94510a <=( a94509a  and  a94506a );
 a94513a <=( (not A300)  and  (not A299) );
 a94516a <=( A302  and  (not A301) );
 a94517a <=( a94516a  and  a94513a );
 a94518a <=( a94517a  and  a94510a );
 a94521a <=( (not A166)  and  (not A167) );
 a94524a <=( A200  and  (not A199) );
 a94525a <=( a94524a  and  a94521a );
 a94528a <=( (not A203)  and  A201 );
 a94531a <=( (not A266)  and  A265 );
 a94532a <=( a94531a  and  a94528a );
 a94533a <=( a94532a  and  a94525a );
 a94536a <=( (not A268)  and  (not A267) );
 a94539a <=( (not A298)  and  A269 );
 a94540a <=( a94539a  and  a94536a );
 a94543a <=( (not A300)  and  A299 );
 a94546a <=( A302  and  (not A301) );
 a94547a <=( a94546a  and  a94543a );
 a94548a <=( a94547a  and  a94540a );
 a94551a <=( (not A166)  and  (not A167) );
 a94554a <=( A200  and  (not A199) );
 a94555a <=( a94554a  and  a94551a );
 a94558a <=( (not A202)  and  (not A201) );
 a94561a <=( (not A265)  and  A203 );
 a94562a <=( a94561a  and  a94558a );
 a94563a <=( a94562a  and  a94555a );
 a94566a <=( A267  and  A266 );
 a94569a <=( A298  and  A268 );
 a94570a <=( a94569a  and  a94566a );
 a94573a <=( (not A300)  and  (not A299) );
 a94576a <=( A302  and  (not A301) );
 a94577a <=( a94576a  and  a94573a );
 a94578a <=( a94577a  and  a94570a );
 a94581a <=( (not A166)  and  (not A167) );
 a94584a <=( A200  and  (not A199) );
 a94585a <=( a94584a  and  a94581a );
 a94588a <=( (not A202)  and  (not A201) );
 a94591a <=( (not A265)  and  A203 );
 a94592a <=( a94591a  and  a94588a );
 a94593a <=( a94592a  and  a94585a );
 a94596a <=( A267  and  A266 );
 a94599a <=( (not A298)  and  A268 );
 a94600a <=( a94599a  and  a94596a );
 a94603a <=( (not A300)  and  A299 );
 a94606a <=( A302  and  (not A301) );
 a94607a <=( a94606a  and  a94603a );
 a94608a <=( a94607a  and  a94600a );
 a94611a <=( (not A166)  and  (not A167) );
 a94614a <=( A200  and  (not A199) );
 a94615a <=( a94614a  and  a94611a );
 a94618a <=( (not A202)  and  (not A201) );
 a94621a <=( (not A265)  and  A203 );
 a94622a <=( a94621a  and  a94618a );
 a94623a <=( a94622a  and  a94615a );
 a94626a <=( A267  and  A266 );
 a94629a <=( A298  and  (not A269) );
 a94630a <=( a94629a  and  a94626a );
 a94633a <=( (not A300)  and  (not A299) );
 a94636a <=( A302  and  (not A301) );
 a94637a <=( a94636a  and  a94633a );
 a94638a <=( a94637a  and  a94630a );
 a94641a <=( (not A166)  and  (not A167) );
 a94644a <=( A200  and  (not A199) );
 a94645a <=( a94644a  and  a94641a );
 a94648a <=( (not A202)  and  (not A201) );
 a94651a <=( (not A265)  and  A203 );
 a94652a <=( a94651a  and  a94648a );
 a94653a <=( a94652a  and  a94645a );
 a94656a <=( A267  and  A266 );
 a94659a <=( (not A298)  and  (not A269) );
 a94660a <=( a94659a  and  a94656a );
 a94663a <=( (not A300)  and  A299 );
 a94666a <=( A302  and  (not A301) );
 a94667a <=( a94666a  and  a94663a );
 a94668a <=( a94667a  and  a94660a );
 a94671a <=( (not A166)  and  (not A167) );
 a94674a <=( A200  and  (not A199) );
 a94675a <=( a94674a  and  a94671a );
 a94678a <=( (not A202)  and  (not A201) );
 a94681a <=( (not A265)  and  A203 );
 a94682a <=( a94681a  and  a94678a );
 a94683a <=( a94682a  and  a94675a );
 a94686a <=( (not A267)  and  A266 );
 a94689a <=( A269  and  (not A268) );
 a94690a <=( a94689a  and  a94686a );
 a94693a <=( (not A299)  and  A298 );
 a94696a <=( A301  and  A300 );
 a94697a <=( a94696a  and  a94693a );
 a94698a <=( a94697a  and  a94690a );
 a94701a <=( (not A166)  and  (not A167) );
 a94704a <=( A200  and  (not A199) );
 a94705a <=( a94704a  and  a94701a );
 a94708a <=( (not A202)  and  (not A201) );
 a94711a <=( (not A265)  and  A203 );
 a94712a <=( a94711a  and  a94708a );
 a94713a <=( a94712a  and  a94705a );
 a94716a <=( (not A267)  and  A266 );
 a94719a <=( A269  and  (not A268) );
 a94720a <=( a94719a  and  a94716a );
 a94723a <=( (not A299)  and  A298 );
 a94726a <=( (not A302)  and  A300 );
 a94727a <=( a94726a  and  a94723a );
 a94728a <=( a94727a  and  a94720a );
 a94731a <=( (not A166)  and  (not A167) );
 a94734a <=( A200  and  (not A199) );
 a94735a <=( a94734a  and  a94731a );
 a94738a <=( (not A202)  and  (not A201) );
 a94741a <=( (not A265)  and  A203 );
 a94742a <=( a94741a  and  a94738a );
 a94743a <=( a94742a  and  a94735a );
 a94746a <=( (not A267)  and  A266 );
 a94749a <=( A269  and  (not A268) );
 a94750a <=( a94749a  and  a94746a );
 a94753a <=( A299  and  (not A298) );
 a94756a <=( A301  and  A300 );
 a94757a <=( a94756a  and  a94753a );
 a94758a <=( a94757a  and  a94750a );
 a94761a <=( (not A166)  and  (not A167) );
 a94764a <=( A200  and  (not A199) );
 a94765a <=( a94764a  and  a94761a );
 a94768a <=( (not A202)  and  (not A201) );
 a94771a <=( (not A265)  and  A203 );
 a94772a <=( a94771a  and  a94768a );
 a94773a <=( a94772a  and  a94765a );
 a94776a <=( (not A267)  and  A266 );
 a94779a <=( A269  and  (not A268) );
 a94780a <=( a94779a  and  a94776a );
 a94783a <=( A299  and  (not A298) );
 a94786a <=( (not A302)  and  A300 );
 a94787a <=( a94786a  and  a94783a );
 a94788a <=( a94787a  and  a94780a );
 a94791a <=( (not A166)  and  (not A167) );
 a94794a <=( A200  and  (not A199) );
 a94795a <=( a94794a  and  a94791a );
 a94798a <=( (not A202)  and  (not A201) );
 a94801a <=( A265  and  A203 );
 a94802a <=( a94801a  and  a94798a );
 a94803a <=( a94802a  and  a94795a );
 a94806a <=( A267  and  (not A266) );
 a94809a <=( A298  and  A268 );
 a94810a <=( a94809a  and  a94806a );
 a94813a <=( (not A300)  and  (not A299) );
 a94816a <=( A302  and  (not A301) );
 a94817a <=( a94816a  and  a94813a );
 a94818a <=( a94817a  and  a94810a );
 a94821a <=( (not A166)  and  (not A167) );
 a94824a <=( A200  and  (not A199) );
 a94825a <=( a94824a  and  a94821a );
 a94828a <=( (not A202)  and  (not A201) );
 a94831a <=( A265  and  A203 );
 a94832a <=( a94831a  and  a94828a );
 a94833a <=( a94832a  and  a94825a );
 a94836a <=( A267  and  (not A266) );
 a94839a <=( (not A298)  and  A268 );
 a94840a <=( a94839a  and  a94836a );
 a94843a <=( (not A300)  and  A299 );
 a94846a <=( A302  and  (not A301) );
 a94847a <=( a94846a  and  a94843a );
 a94848a <=( a94847a  and  a94840a );
 a94851a <=( (not A166)  and  (not A167) );
 a94854a <=( A200  and  (not A199) );
 a94855a <=( a94854a  and  a94851a );
 a94858a <=( (not A202)  and  (not A201) );
 a94861a <=( A265  and  A203 );
 a94862a <=( a94861a  and  a94858a );
 a94863a <=( a94862a  and  a94855a );
 a94866a <=( A267  and  (not A266) );
 a94869a <=( A298  and  (not A269) );
 a94870a <=( a94869a  and  a94866a );
 a94873a <=( (not A300)  and  (not A299) );
 a94876a <=( A302  and  (not A301) );
 a94877a <=( a94876a  and  a94873a );
 a94878a <=( a94877a  and  a94870a );
 a94881a <=( (not A166)  and  (not A167) );
 a94884a <=( A200  and  (not A199) );
 a94885a <=( a94884a  and  a94881a );
 a94888a <=( (not A202)  and  (not A201) );
 a94891a <=( A265  and  A203 );
 a94892a <=( a94891a  and  a94888a );
 a94893a <=( a94892a  and  a94885a );
 a94896a <=( A267  and  (not A266) );
 a94899a <=( (not A298)  and  (not A269) );
 a94900a <=( a94899a  and  a94896a );
 a94903a <=( (not A300)  and  A299 );
 a94906a <=( A302  and  (not A301) );
 a94907a <=( a94906a  and  a94903a );
 a94908a <=( a94907a  and  a94900a );
 a94911a <=( (not A166)  and  (not A167) );
 a94914a <=( A200  and  (not A199) );
 a94915a <=( a94914a  and  a94911a );
 a94918a <=( (not A202)  and  (not A201) );
 a94921a <=( A265  and  A203 );
 a94922a <=( a94921a  and  a94918a );
 a94923a <=( a94922a  and  a94915a );
 a94926a <=( (not A267)  and  (not A266) );
 a94929a <=( A269  and  (not A268) );
 a94930a <=( a94929a  and  a94926a );
 a94933a <=( (not A299)  and  A298 );
 a94936a <=( A301  and  A300 );
 a94937a <=( a94936a  and  a94933a );
 a94938a <=( a94937a  and  a94930a );
 a94941a <=( (not A166)  and  (not A167) );
 a94944a <=( A200  and  (not A199) );
 a94945a <=( a94944a  and  a94941a );
 a94948a <=( (not A202)  and  (not A201) );
 a94951a <=( A265  and  A203 );
 a94952a <=( a94951a  and  a94948a );
 a94953a <=( a94952a  and  a94945a );
 a94956a <=( (not A267)  and  (not A266) );
 a94959a <=( A269  and  (not A268) );
 a94960a <=( a94959a  and  a94956a );
 a94963a <=( (not A299)  and  A298 );
 a94966a <=( (not A302)  and  A300 );
 a94967a <=( a94966a  and  a94963a );
 a94968a <=( a94967a  and  a94960a );
 a94971a <=( (not A166)  and  (not A167) );
 a94974a <=( A200  and  (not A199) );
 a94975a <=( a94974a  and  a94971a );
 a94978a <=( (not A202)  and  (not A201) );
 a94981a <=( A265  and  A203 );
 a94982a <=( a94981a  and  a94978a );
 a94983a <=( a94982a  and  a94975a );
 a94986a <=( (not A267)  and  (not A266) );
 a94989a <=( A269  and  (not A268) );
 a94990a <=( a94989a  and  a94986a );
 a94993a <=( A299  and  (not A298) );
 a94996a <=( A301  and  A300 );
 a94997a <=( a94996a  and  a94993a );
 a94998a <=( a94997a  and  a94990a );
 a95001a <=( (not A166)  and  (not A167) );
 a95004a <=( A200  and  (not A199) );
 a95005a <=( a95004a  and  a95001a );
 a95008a <=( (not A202)  and  (not A201) );
 a95011a <=( A265  and  A203 );
 a95012a <=( a95011a  and  a95008a );
 a95013a <=( a95012a  and  a95005a );
 a95016a <=( (not A267)  and  (not A266) );
 a95019a <=( A269  and  (not A268) );
 a95020a <=( a95019a  and  a95016a );
 a95023a <=( A299  and  (not A298) );
 a95026a <=( (not A302)  and  A300 );
 a95027a <=( a95026a  and  a95023a );
 a95028a <=( a95027a  and  a95020a );
 a95031a <=( (not A166)  and  (not A167) );
 a95034a <=( (not A200)  and  A199 );
 a95035a <=( a95034a  and  a95031a );
 a95038a <=( A202  and  A201 );
 a95041a <=( A266  and  (not A265) );
 a95042a <=( a95041a  and  a95038a );
 a95043a <=( a95042a  and  a95035a );
 a95046a <=( (not A268)  and  (not A267) );
 a95049a <=( A298  and  A269 );
 a95050a <=( a95049a  and  a95046a );
 a95053a <=( (not A300)  and  (not A299) );
 a95056a <=( A302  and  (not A301) );
 a95057a <=( a95056a  and  a95053a );
 a95058a <=( a95057a  and  a95050a );
 a95061a <=( (not A166)  and  (not A167) );
 a95064a <=( (not A200)  and  A199 );
 a95065a <=( a95064a  and  a95061a );
 a95068a <=( A202  and  A201 );
 a95071a <=( A266  and  (not A265) );
 a95072a <=( a95071a  and  a95068a );
 a95073a <=( a95072a  and  a95065a );
 a95076a <=( (not A268)  and  (not A267) );
 a95079a <=( (not A298)  and  A269 );
 a95080a <=( a95079a  and  a95076a );
 a95083a <=( (not A300)  and  A299 );
 a95086a <=( A302  and  (not A301) );
 a95087a <=( a95086a  and  a95083a );
 a95088a <=( a95087a  and  a95080a );
 a95091a <=( (not A166)  and  (not A167) );
 a95094a <=( (not A200)  and  A199 );
 a95095a <=( a95094a  and  a95091a );
 a95098a <=( A202  and  A201 );
 a95101a <=( (not A266)  and  A265 );
 a95102a <=( a95101a  and  a95098a );
 a95103a <=( a95102a  and  a95095a );
 a95106a <=( (not A268)  and  (not A267) );
 a95109a <=( A298  and  A269 );
 a95110a <=( a95109a  and  a95106a );
 a95113a <=( (not A300)  and  (not A299) );
 a95116a <=( A302  and  (not A301) );
 a95117a <=( a95116a  and  a95113a );
 a95118a <=( a95117a  and  a95110a );
 a95121a <=( (not A166)  and  (not A167) );
 a95124a <=( (not A200)  and  A199 );
 a95125a <=( a95124a  and  a95121a );
 a95128a <=( A202  and  A201 );
 a95131a <=( (not A266)  and  A265 );
 a95132a <=( a95131a  and  a95128a );
 a95133a <=( a95132a  and  a95125a );
 a95136a <=( (not A268)  and  (not A267) );
 a95139a <=( (not A298)  and  A269 );
 a95140a <=( a95139a  and  a95136a );
 a95143a <=( (not A300)  and  A299 );
 a95146a <=( A302  and  (not A301) );
 a95147a <=( a95146a  and  a95143a );
 a95148a <=( a95147a  and  a95140a );
 a95151a <=( (not A166)  and  (not A167) );
 a95154a <=( (not A200)  and  A199 );
 a95155a <=( a95154a  and  a95151a );
 a95158a <=( (not A203)  and  A201 );
 a95161a <=( A266  and  (not A265) );
 a95162a <=( a95161a  and  a95158a );
 a95163a <=( a95162a  and  a95155a );
 a95166a <=( (not A268)  and  (not A267) );
 a95169a <=( A298  and  A269 );
 a95170a <=( a95169a  and  a95166a );
 a95173a <=( (not A300)  and  (not A299) );
 a95176a <=( A302  and  (not A301) );
 a95177a <=( a95176a  and  a95173a );
 a95178a <=( a95177a  and  a95170a );
 a95181a <=( (not A166)  and  (not A167) );
 a95184a <=( (not A200)  and  A199 );
 a95185a <=( a95184a  and  a95181a );
 a95188a <=( (not A203)  and  A201 );
 a95191a <=( A266  and  (not A265) );
 a95192a <=( a95191a  and  a95188a );
 a95193a <=( a95192a  and  a95185a );
 a95196a <=( (not A268)  and  (not A267) );
 a95199a <=( (not A298)  and  A269 );
 a95200a <=( a95199a  and  a95196a );
 a95203a <=( (not A300)  and  A299 );
 a95206a <=( A302  and  (not A301) );
 a95207a <=( a95206a  and  a95203a );
 a95208a <=( a95207a  and  a95200a );
 a95211a <=( (not A166)  and  (not A167) );
 a95214a <=( (not A200)  and  A199 );
 a95215a <=( a95214a  and  a95211a );
 a95218a <=( (not A203)  and  A201 );
 a95221a <=( (not A266)  and  A265 );
 a95222a <=( a95221a  and  a95218a );
 a95223a <=( a95222a  and  a95215a );
 a95226a <=( (not A268)  and  (not A267) );
 a95229a <=( A298  and  A269 );
 a95230a <=( a95229a  and  a95226a );
 a95233a <=( (not A300)  and  (not A299) );
 a95236a <=( A302  and  (not A301) );
 a95237a <=( a95236a  and  a95233a );
 a95238a <=( a95237a  and  a95230a );
 a95241a <=( (not A166)  and  (not A167) );
 a95244a <=( (not A200)  and  A199 );
 a95245a <=( a95244a  and  a95241a );
 a95248a <=( (not A203)  and  A201 );
 a95251a <=( (not A266)  and  A265 );
 a95252a <=( a95251a  and  a95248a );
 a95253a <=( a95252a  and  a95245a );
 a95256a <=( (not A268)  and  (not A267) );
 a95259a <=( (not A298)  and  A269 );
 a95260a <=( a95259a  and  a95256a );
 a95263a <=( (not A300)  and  A299 );
 a95266a <=( A302  and  (not A301) );
 a95267a <=( a95266a  and  a95263a );
 a95268a <=( a95267a  and  a95260a );
 a95271a <=( (not A166)  and  (not A167) );
 a95274a <=( (not A200)  and  A199 );
 a95275a <=( a95274a  and  a95271a );
 a95278a <=( (not A202)  and  (not A201) );
 a95281a <=( (not A265)  and  A203 );
 a95282a <=( a95281a  and  a95278a );
 a95283a <=( a95282a  and  a95275a );
 a95286a <=( A267  and  A266 );
 a95289a <=( A298  and  A268 );
 a95290a <=( a95289a  and  a95286a );
 a95293a <=( (not A300)  and  (not A299) );
 a95296a <=( A302  and  (not A301) );
 a95297a <=( a95296a  and  a95293a );
 a95298a <=( a95297a  and  a95290a );
 a95301a <=( (not A166)  and  (not A167) );
 a95304a <=( (not A200)  and  A199 );
 a95305a <=( a95304a  and  a95301a );
 a95308a <=( (not A202)  and  (not A201) );
 a95311a <=( (not A265)  and  A203 );
 a95312a <=( a95311a  and  a95308a );
 a95313a <=( a95312a  and  a95305a );
 a95316a <=( A267  and  A266 );
 a95319a <=( (not A298)  and  A268 );
 a95320a <=( a95319a  and  a95316a );
 a95323a <=( (not A300)  and  A299 );
 a95326a <=( A302  and  (not A301) );
 a95327a <=( a95326a  and  a95323a );
 a95328a <=( a95327a  and  a95320a );
 a95331a <=( (not A166)  and  (not A167) );
 a95334a <=( (not A200)  and  A199 );
 a95335a <=( a95334a  and  a95331a );
 a95338a <=( (not A202)  and  (not A201) );
 a95341a <=( (not A265)  and  A203 );
 a95342a <=( a95341a  and  a95338a );
 a95343a <=( a95342a  and  a95335a );
 a95346a <=( A267  and  A266 );
 a95349a <=( A298  and  (not A269) );
 a95350a <=( a95349a  and  a95346a );
 a95353a <=( (not A300)  and  (not A299) );
 a95356a <=( A302  and  (not A301) );
 a95357a <=( a95356a  and  a95353a );
 a95358a <=( a95357a  and  a95350a );
 a95361a <=( (not A166)  and  (not A167) );
 a95364a <=( (not A200)  and  A199 );
 a95365a <=( a95364a  and  a95361a );
 a95368a <=( (not A202)  and  (not A201) );
 a95371a <=( (not A265)  and  A203 );
 a95372a <=( a95371a  and  a95368a );
 a95373a <=( a95372a  and  a95365a );
 a95376a <=( A267  and  A266 );
 a95379a <=( (not A298)  and  (not A269) );
 a95380a <=( a95379a  and  a95376a );
 a95383a <=( (not A300)  and  A299 );
 a95386a <=( A302  and  (not A301) );
 a95387a <=( a95386a  and  a95383a );
 a95388a <=( a95387a  and  a95380a );
 a95391a <=( (not A166)  and  (not A167) );
 a95394a <=( (not A200)  and  A199 );
 a95395a <=( a95394a  and  a95391a );
 a95398a <=( (not A202)  and  (not A201) );
 a95401a <=( (not A265)  and  A203 );
 a95402a <=( a95401a  and  a95398a );
 a95403a <=( a95402a  and  a95395a );
 a95406a <=( (not A267)  and  A266 );
 a95409a <=( A269  and  (not A268) );
 a95410a <=( a95409a  and  a95406a );
 a95413a <=( (not A299)  and  A298 );
 a95416a <=( A301  and  A300 );
 a95417a <=( a95416a  and  a95413a );
 a95418a <=( a95417a  and  a95410a );
 a95421a <=( (not A166)  and  (not A167) );
 a95424a <=( (not A200)  and  A199 );
 a95425a <=( a95424a  and  a95421a );
 a95428a <=( (not A202)  and  (not A201) );
 a95431a <=( (not A265)  and  A203 );
 a95432a <=( a95431a  and  a95428a );
 a95433a <=( a95432a  and  a95425a );
 a95436a <=( (not A267)  and  A266 );
 a95439a <=( A269  and  (not A268) );
 a95440a <=( a95439a  and  a95436a );
 a95443a <=( (not A299)  and  A298 );
 a95446a <=( (not A302)  and  A300 );
 a95447a <=( a95446a  and  a95443a );
 a95448a <=( a95447a  and  a95440a );
 a95451a <=( (not A166)  and  (not A167) );
 a95454a <=( (not A200)  and  A199 );
 a95455a <=( a95454a  and  a95451a );
 a95458a <=( (not A202)  and  (not A201) );
 a95461a <=( (not A265)  and  A203 );
 a95462a <=( a95461a  and  a95458a );
 a95463a <=( a95462a  and  a95455a );
 a95466a <=( (not A267)  and  A266 );
 a95469a <=( A269  and  (not A268) );
 a95470a <=( a95469a  and  a95466a );
 a95473a <=( A299  and  (not A298) );
 a95476a <=( A301  and  A300 );
 a95477a <=( a95476a  and  a95473a );
 a95478a <=( a95477a  and  a95470a );
 a95481a <=( (not A166)  and  (not A167) );
 a95484a <=( (not A200)  and  A199 );
 a95485a <=( a95484a  and  a95481a );
 a95488a <=( (not A202)  and  (not A201) );
 a95491a <=( (not A265)  and  A203 );
 a95492a <=( a95491a  and  a95488a );
 a95493a <=( a95492a  and  a95485a );
 a95496a <=( (not A267)  and  A266 );
 a95499a <=( A269  and  (not A268) );
 a95500a <=( a95499a  and  a95496a );
 a95503a <=( A299  and  (not A298) );
 a95506a <=( (not A302)  and  A300 );
 a95507a <=( a95506a  and  a95503a );
 a95508a <=( a95507a  and  a95500a );
 a95511a <=( (not A166)  and  (not A167) );
 a95514a <=( (not A200)  and  A199 );
 a95515a <=( a95514a  and  a95511a );
 a95518a <=( (not A202)  and  (not A201) );
 a95521a <=( A265  and  A203 );
 a95522a <=( a95521a  and  a95518a );
 a95523a <=( a95522a  and  a95515a );
 a95526a <=( A267  and  (not A266) );
 a95529a <=( A298  and  A268 );
 a95530a <=( a95529a  and  a95526a );
 a95533a <=( (not A300)  and  (not A299) );
 a95536a <=( A302  and  (not A301) );
 a95537a <=( a95536a  and  a95533a );
 a95538a <=( a95537a  and  a95530a );
 a95541a <=( (not A166)  and  (not A167) );
 a95544a <=( (not A200)  and  A199 );
 a95545a <=( a95544a  and  a95541a );
 a95548a <=( (not A202)  and  (not A201) );
 a95551a <=( A265  and  A203 );
 a95552a <=( a95551a  and  a95548a );
 a95553a <=( a95552a  and  a95545a );
 a95556a <=( A267  and  (not A266) );
 a95559a <=( (not A298)  and  A268 );
 a95560a <=( a95559a  and  a95556a );
 a95563a <=( (not A300)  and  A299 );
 a95566a <=( A302  and  (not A301) );
 a95567a <=( a95566a  and  a95563a );
 a95568a <=( a95567a  and  a95560a );
 a95571a <=( (not A166)  and  (not A167) );
 a95574a <=( (not A200)  and  A199 );
 a95575a <=( a95574a  and  a95571a );
 a95578a <=( (not A202)  and  (not A201) );
 a95581a <=( A265  and  A203 );
 a95582a <=( a95581a  and  a95578a );
 a95583a <=( a95582a  and  a95575a );
 a95586a <=( A267  and  (not A266) );
 a95589a <=( A298  and  (not A269) );
 a95590a <=( a95589a  and  a95586a );
 a95593a <=( (not A300)  and  (not A299) );
 a95596a <=( A302  and  (not A301) );
 a95597a <=( a95596a  and  a95593a );
 a95598a <=( a95597a  and  a95590a );
 a95601a <=( (not A166)  and  (not A167) );
 a95604a <=( (not A200)  and  A199 );
 a95605a <=( a95604a  and  a95601a );
 a95608a <=( (not A202)  and  (not A201) );
 a95611a <=( A265  and  A203 );
 a95612a <=( a95611a  and  a95608a );
 a95613a <=( a95612a  and  a95605a );
 a95616a <=( A267  and  (not A266) );
 a95619a <=( (not A298)  and  (not A269) );
 a95620a <=( a95619a  and  a95616a );
 a95623a <=( (not A300)  and  A299 );
 a95626a <=( A302  and  (not A301) );
 a95627a <=( a95626a  and  a95623a );
 a95628a <=( a95627a  and  a95620a );
 a95631a <=( (not A166)  and  (not A167) );
 a95634a <=( (not A200)  and  A199 );
 a95635a <=( a95634a  and  a95631a );
 a95638a <=( (not A202)  and  (not A201) );
 a95641a <=( A265  and  A203 );
 a95642a <=( a95641a  and  a95638a );
 a95643a <=( a95642a  and  a95635a );
 a95646a <=( (not A267)  and  (not A266) );
 a95649a <=( A269  and  (not A268) );
 a95650a <=( a95649a  and  a95646a );
 a95653a <=( (not A299)  and  A298 );
 a95656a <=( A301  and  A300 );
 a95657a <=( a95656a  and  a95653a );
 a95658a <=( a95657a  and  a95650a );
 a95661a <=( (not A166)  and  (not A167) );
 a95664a <=( (not A200)  and  A199 );
 a95665a <=( a95664a  and  a95661a );
 a95668a <=( (not A202)  and  (not A201) );
 a95671a <=( A265  and  A203 );
 a95672a <=( a95671a  and  a95668a );
 a95673a <=( a95672a  and  a95665a );
 a95676a <=( (not A267)  and  (not A266) );
 a95679a <=( A269  and  (not A268) );
 a95680a <=( a95679a  and  a95676a );
 a95683a <=( (not A299)  and  A298 );
 a95686a <=( (not A302)  and  A300 );
 a95687a <=( a95686a  and  a95683a );
 a95688a <=( a95687a  and  a95680a );
 a95691a <=( (not A166)  and  (not A167) );
 a95694a <=( (not A200)  and  A199 );
 a95695a <=( a95694a  and  a95691a );
 a95698a <=( (not A202)  and  (not A201) );
 a95701a <=( A265  and  A203 );
 a95702a <=( a95701a  and  a95698a );
 a95703a <=( a95702a  and  a95695a );
 a95706a <=( (not A267)  and  (not A266) );
 a95709a <=( A269  and  (not A268) );
 a95710a <=( a95709a  and  a95706a );
 a95713a <=( A299  and  (not A298) );
 a95716a <=( A301  and  A300 );
 a95717a <=( a95716a  and  a95713a );
 a95718a <=( a95717a  and  a95710a );
 a95721a <=( (not A166)  and  (not A167) );
 a95724a <=( (not A200)  and  A199 );
 a95725a <=( a95724a  and  a95721a );
 a95728a <=( (not A202)  and  (not A201) );
 a95731a <=( A265  and  A203 );
 a95732a <=( a95731a  and  a95728a );
 a95733a <=( a95732a  and  a95725a );
 a95736a <=( (not A267)  and  (not A266) );
 a95739a <=( A269  and  (not A268) );
 a95740a <=( a95739a  and  a95736a );
 a95743a <=( A299  and  (not A298) );
 a95746a <=( (not A302)  and  A300 );
 a95747a <=( a95746a  and  a95743a );
 a95748a <=( a95747a  and  a95740a );
 a95751a <=( (not A168)  and  A170 );
 a95754a <=( A200  and  (not A199) );
 a95755a <=( a95754a  and  a95751a );
 a95758a <=( A202  and  A201 );
 a95761a <=( A266  and  (not A265) );
 a95762a <=( a95761a  and  a95758a );
 a95763a <=( a95762a  and  a95755a );
 a95766a <=( (not A268)  and  (not A267) );
 a95769a <=( A298  and  A269 );
 a95770a <=( a95769a  and  a95766a );
 a95773a <=( (not A300)  and  (not A299) );
 a95776a <=( A302  and  (not A301) );
 a95777a <=( a95776a  and  a95773a );
 a95778a <=( a95777a  and  a95770a );
 a95781a <=( (not A168)  and  A170 );
 a95784a <=( A200  and  (not A199) );
 a95785a <=( a95784a  and  a95781a );
 a95788a <=( A202  and  A201 );
 a95791a <=( A266  and  (not A265) );
 a95792a <=( a95791a  and  a95788a );
 a95793a <=( a95792a  and  a95785a );
 a95796a <=( (not A268)  and  (not A267) );
 a95799a <=( (not A298)  and  A269 );
 a95800a <=( a95799a  and  a95796a );
 a95803a <=( (not A300)  and  A299 );
 a95806a <=( A302  and  (not A301) );
 a95807a <=( a95806a  and  a95803a );
 a95808a <=( a95807a  and  a95800a );
 a95811a <=( (not A168)  and  A170 );
 a95814a <=( A200  and  (not A199) );
 a95815a <=( a95814a  and  a95811a );
 a95818a <=( A202  and  A201 );
 a95821a <=( (not A266)  and  A265 );
 a95822a <=( a95821a  and  a95818a );
 a95823a <=( a95822a  and  a95815a );
 a95826a <=( (not A268)  and  (not A267) );
 a95829a <=( A298  and  A269 );
 a95830a <=( a95829a  and  a95826a );
 a95833a <=( (not A300)  and  (not A299) );
 a95836a <=( A302  and  (not A301) );
 a95837a <=( a95836a  and  a95833a );
 a95838a <=( a95837a  and  a95830a );
 a95841a <=( (not A168)  and  A170 );
 a95844a <=( A200  and  (not A199) );
 a95845a <=( a95844a  and  a95841a );
 a95848a <=( A202  and  A201 );
 a95851a <=( (not A266)  and  A265 );
 a95852a <=( a95851a  and  a95848a );
 a95853a <=( a95852a  and  a95845a );
 a95856a <=( (not A268)  and  (not A267) );
 a95859a <=( (not A298)  and  A269 );
 a95860a <=( a95859a  and  a95856a );
 a95863a <=( (not A300)  and  A299 );
 a95866a <=( A302  and  (not A301) );
 a95867a <=( a95866a  and  a95863a );
 a95868a <=( a95867a  and  a95860a );
 a95871a <=( (not A168)  and  A170 );
 a95874a <=( A200  and  (not A199) );
 a95875a <=( a95874a  and  a95871a );
 a95878a <=( (not A203)  and  A201 );
 a95881a <=( A266  and  (not A265) );
 a95882a <=( a95881a  and  a95878a );
 a95883a <=( a95882a  and  a95875a );
 a95886a <=( (not A268)  and  (not A267) );
 a95889a <=( A298  and  A269 );
 a95890a <=( a95889a  and  a95886a );
 a95893a <=( (not A300)  and  (not A299) );
 a95896a <=( A302  and  (not A301) );
 a95897a <=( a95896a  and  a95893a );
 a95898a <=( a95897a  and  a95890a );
 a95901a <=( (not A168)  and  A170 );
 a95904a <=( A200  and  (not A199) );
 a95905a <=( a95904a  and  a95901a );
 a95908a <=( (not A203)  and  A201 );
 a95911a <=( A266  and  (not A265) );
 a95912a <=( a95911a  and  a95908a );
 a95913a <=( a95912a  and  a95905a );
 a95916a <=( (not A268)  and  (not A267) );
 a95919a <=( (not A298)  and  A269 );
 a95920a <=( a95919a  and  a95916a );
 a95923a <=( (not A300)  and  A299 );
 a95926a <=( A302  and  (not A301) );
 a95927a <=( a95926a  and  a95923a );
 a95928a <=( a95927a  and  a95920a );
 a95931a <=( (not A168)  and  A170 );
 a95934a <=( A200  and  (not A199) );
 a95935a <=( a95934a  and  a95931a );
 a95938a <=( (not A203)  and  A201 );
 a95941a <=( (not A266)  and  A265 );
 a95942a <=( a95941a  and  a95938a );
 a95943a <=( a95942a  and  a95935a );
 a95946a <=( (not A268)  and  (not A267) );
 a95949a <=( A298  and  A269 );
 a95950a <=( a95949a  and  a95946a );
 a95953a <=( (not A300)  and  (not A299) );
 a95956a <=( A302  and  (not A301) );
 a95957a <=( a95956a  and  a95953a );
 a95958a <=( a95957a  and  a95950a );
 a95961a <=( (not A168)  and  A170 );
 a95964a <=( A200  and  (not A199) );
 a95965a <=( a95964a  and  a95961a );
 a95968a <=( (not A203)  and  A201 );
 a95971a <=( (not A266)  and  A265 );
 a95972a <=( a95971a  and  a95968a );
 a95973a <=( a95972a  and  a95965a );
 a95976a <=( (not A268)  and  (not A267) );
 a95979a <=( (not A298)  and  A269 );
 a95980a <=( a95979a  and  a95976a );
 a95983a <=( (not A300)  and  A299 );
 a95986a <=( A302  and  (not A301) );
 a95987a <=( a95986a  and  a95983a );
 a95988a <=( a95987a  and  a95980a );
 a95991a <=( (not A168)  and  A170 );
 a95994a <=( A200  and  (not A199) );
 a95995a <=( a95994a  and  a95991a );
 a95998a <=( (not A202)  and  (not A201) );
 a96001a <=( (not A265)  and  A203 );
 a96002a <=( a96001a  and  a95998a );
 a96003a <=( a96002a  and  a95995a );
 a96006a <=( A267  and  A266 );
 a96009a <=( A298  and  A268 );
 a96010a <=( a96009a  and  a96006a );
 a96013a <=( (not A300)  and  (not A299) );
 a96016a <=( A302  and  (not A301) );
 a96017a <=( a96016a  and  a96013a );
 a96018a <=( a96017a  and  a96010a );
 a96021a <=( (not A168)  and  A170 );
 a96024a <=( A200  and  (not A199) );
 a96025a <=( a96024a  and  a96021a );
 a96028a <=( (not A202)  and  (not A201) );
 a96031a <=( (not A265)  and  A203 );
 a96032a <=( a96031a  and  a96028a );
 a96033a <=( a96032a  and  a96025a );
 a96036a <=( A267  and  A266 );
 a96039a <=( (not A298)  and  A268 );
 a96040a <=( a96039a  and  a96036a );
 a96043a <=( (not A300)  and  A299 );
 a96046a <=( A302  and  (not A301) );
 a96047a <=( a96046a  and  a96043a );
 a96048a <=( a96047a  and  a96040a );
 a96051a <=( (not A168)  and  A170 );
 a96054a <=( A200  and  (not A199) );
 a96055a <=( a96054a  and  a96051a );
 a96058a <=( (not A202)  and  (not A201) );
 a96061a <=( (not A265)  and  A203 );
 a96062a <=( a96061a  and  a96058a );
 a96063a <=( a96062a  and  a96055a );
 a96066a <=( A267  and  A266 );
 a96069a <=( A298  and  (not A269) );
 a96070a <=( a96069a  and  a96066a );
 a96073a <=( (not A300)  and  (not A299) );
 a96076a <=( A302  and  (not A301) );
 a96077a <=( a96076a  and  a96073a );
 a96078a <=( a96077a  and  a96070a );
 a96081a <=( (not A168)  and  A170 );
 a96084a <=( A200  and  (not A199) );
 a96085a <=( a96084a  and  a96081a );
 a96088a <=( (not A202)  and  (not A201) );
 a96091a <=( (not A265)  and  A203 );
 a96092a <=( a96091a  and  a96088a );
 a96093a <=( a96092a  and  a96085a );
 a96096a <=( A267  and  A266 );
 a96099a <=( (not A298)  and  (not A269) );
 a96100a <=( a96099a  and  a96096a );
 a96103a <=( (not A300)  and  A299 );
 a96106a <=( A302  and  (not A301) );
 a96107a <=( a96106a  and  a96103a );
 a96108a <=( a96107a  and  a96100a );
 a96111a <=( (not A168)  and  A170 );
 a96114a <=( A200  and  (not A199) );
 a96115a <=( a96114a  and  a96111a );
 a96118a <=( (not A202)  and  (not A201) );
 a96121a <=( (not A265)  and  A203 );
 a96122a <=( a96121a  and  a96118a );
 a96123a <=( a96122a  and  a96115a );
 a96126a <=( (not A267)  and  A266 );
 a96129a <=( A269  and  (not A268) );
 a96130a <=( a96129a  and  a96126a );
 a96133a <=( (not A299)  and  A298 );
 a96136a <=( A301  and  A300 );
 a96137a <=( a96136a  and  a96133a );
 a96138a <=( a96137a  and  a96130a );
 a96141a <=( (not A168)  and  A170 );
 a96144a <=( A200  and  (not A199) );
 a96145a <=( a96144a  and  a96141a );
 a96148a <=( (not A202)  and  (not A201) );
 a96151a <=( (not A265)  and  A203 );
 a96152a <=( a96151a  and  a96148a );
 a96153a <=( a96152a  and  a96145a );
 a96156a <=( (not A267)  and  A266 );
 a96159a <=( A269  and  (not A268) );
 a96160a <=( a96159a  and  a96156a );
 a96163a <=( (not A299)  and  A298 );
 a96166a <=( (not A302)  and  A300 );
 a96167a <=( a96166a  and  a96163a );
 a96168a <=( a96167a  and  a96160a );
 a96171a <=( (not A168)  and  A170 );
 a96174a <=( A200  and  (not A199) );
 a96175a <=( a96174a  and  a96171a );
 a96178a <=( (not A202)  and  (not A201) );
 a96181a <=( (not A265)  and  A203 );
 a96182a <=( a96181a  and  a96178a );
 a96183a <=( a96182a  and  a96175a );
 a96186a <=( (not A267)  and  A266 );
 a96189a <=( A269  and  (not A268) );
 a96190a <=( a96189a  and  a96186a );
 a96193a <=( A299  and  (not A298) );
 a96196a <=( A301  and  A300 );
 a96197a <=( a96196a  and  a96193a );
 a96198a <=( a96197a  and  a96190a );
 a96201a <=( (not A168)  and  A170 );
 a96204a <=( A200  and  (not A199) );
 a96205a <=( a96204a  and  a96201a );
 a96208a <=( (not A202)  and  (not A201) );
 a96211a <=( (not A265)  and  A203 );
 a96212a <=( a96211a  and  a96208a );
 a96213a <=( a96212a  and  a96205a );
 a96216a <=( (not A267)  and  A266 );
 a96219a <=( A269  and  (not A268) );
 a96220a <=( a96219a  and  a96216a );
 a96223a <=( A299  and  (not A298) );
 a96226a <=( (not A302)  and  A300 );
 a96227a <=( a96226a  and  a96223a );
 a96228a <=( a96227a  and  a96220a );
 a96231a <=( (not A168)  and  A170 );
 a96234a <=( A200  and  (not A199) );
 a96235a <=( a96234a  and  a96231a );
 a96238a <=( (not A202)  and  (not A201) );
 a96241a <=( A265  and  A203 );
 a96242a <=( a96241a  and  a96238a );
 a96243a <=( a96242a  and  a96235a );
 a96246a <=( A267  and  (not A266) );
 a96249a <=( A298  and  A268 );
 a96250a <=( a96249a  and  a96246a );
 a96253a <=( (not A300)  and  (not A299) );
 a96256a <=( A302  and  (not A301) );
 a96257a <=( a96256a  and  a96253a );
 a96258a <=( a96257a  and  a96250a );
 a96261a <=( (not A168)  and  A170 );
 a96264a <=( A200  and  (not A199) );
 a96265a <=( a96264a  and  a96261a );
 a96268a <=( (not A202)  and  (not A201) );
 a96271a <=( A265  and  A203 );
 a96272a <=( a96271a  and  a96268a );
 a96273a <=( a96272a  and  a96265a );
 a96276a <=( A267  and  (not A266) );
 a96279a <=( (not A298)  and  A268 );
 a96280a <=( a96279a  and  a96276a );
 a96283a <=( (not A300)  and  A299 );
 a96286a <=( A302  and  (not A301) );
 a96287a <=( a96286a  and  a96283a );
 a96288a <=( a96287a  and  a96280a );
 a96291a <=( (not A168)  and  A170 );
 a96294a <=( A200  and  (not A199) );
 a96295a <=( a96294a  and  a96291a );
 a96298a <=( (not A202)  and  (not A201) );
 a96301a <=( A265  and  A203 );
 a96302a <=( a96301a  and  a96298a );
 a96303a <=( a96302a  and  a96295a );
 a96306a <=( A267  and  (not A266) );
 a96309a <=( A298  and  (not A269) );
 a96310a <=( a96309a  and  a96306a );
 a96313a <=( (not A300)  and  (not A299) );
 a96316a <=( A302  and  (not A301) );
 a96317a <=( a96316a  and  a96313a );
 a96318a <=( a96317a  and  a96310a );
 a96321a <=( (not A168)  and  A170 );
 a96324a <=( A200  and  (not A199) );
 a96325a <=( a96324a  and  a96321a );
 a96328a <=( (not A202)  and  (not A201) );
 a96331a <=( A265  and  A203 );
 a96332a <=( a96331a  and  a96328a );
 a96333a <=( a96332a  and  a96325a );
 a96336a <=( A267  and  (not A266) );
 a96339a <=( (not A298)  and  (not A269) );
 a96340a <=( a96339a  and  a96336a );
 a96343a <=( (not A300)  and  A299 );
 a96346a <=( A302  and  (not A301) );
 a96347a <=( a96346a  and  a96343a );
 a96348a <=( a96347a  and  a96340a );
 a96351a <=( (not A168)  and  A170 );
 a96354a <=( A200  and  (not A199) );
 a96355a <=( a96354a  and  a96351a );
 a96358a <=( (not A202)  and  (not A201) );
 a96361a <=( A265  and  A203 );
 a96362a <=( a96361a  and  a96358a );
 a96363a <=( a96362a  and  a96355a );
 a96366a <=( (not A267)  and  (not A266) );
 a96369a <=( A269  and  (not A268) );
 a96370a <=( a96369a  and  a96366a );
 a96373a <=( (not A299)  and  A298 );
 a96376a <=( A301  and  A300 );
 a96377a <=( a96376a  and  a96373a );
 a96378a <=( a96377a  and  a96370a );
 a96381a <=( (not A168)  and  A170 );
 a96384a <=( A200  and  (not A199) );
 a96385a <=( a96384a  and  a96381a );
 a96388a <=( (not A202)  and  (not A201) );
 a96391a <=( A265  and  A203 );
 a96392a <=( a96391a  and  a96388a );
 a96393a <=( a96392a  and  a96385a );
 a96396a <=( (not A267)  and  (not A266) );
 a96399a <=( A269  and  (not A268) );
 a96400a <=( a96399a  and  a96396a );
 a96403a <=( (not A299)  and  A298 );
 a96406a <=( (not A302)  and  A300 );
 a96407a <=( a96406a  and  a96403a );
 a96408a <=( a96407a  and  a96400a );
 a96411a <=( (not A168)  and  A170 );
 a96414a <=( A200  and  (not A199) );
 a96415a <=( a96414a  and  a96411a );
 a96418a <=( (not A202)  and  (not A201) );
 a96421a <=( A265  and  A203 );
 a96422a <=( a96421a  and  a96418a );
 a96423a <=( a96422a  and  a96415a );
 a96426a <=( (not A267)  and  (not A266) );
 a96429a <=( A269  and  (not A268) );
 a96430a <=( a96429a  and  a96426a );
 a96433a <=( A299  and  (not A298) );
 a96436a <=( A301  and  A300 );
 a96437a <=( a96436a  and  a96433a );
 a96438a <=( a96437a  and  a96430a );
 a96441a <=( (not A168)  and  A170 );
 a96444a <=( A200  and  (not A199) );
 a96445a <=( a96444a  and  a96441a );
 a96448a <=( (not A202)  and  (not A201) );
 a96451a <=( A265  and  A203 );
 a96452a <=( a96451a  and  a96448a );
 a96453a <=( a96452a  and  a96445a );
 a96456a <=( (not A267)  and  (not A266) );
 a96459a <=( A269  and  (not A268) );
 a96460a <=( a96459a  and  a96456a );
 a96463a <=( A299  and  (not A298) );
 a96466a <=( (not A302)  and  A300 );
 a96467a <=( a96466a  and  a96463a );
 a96468a <=( a96467a  and  a96460a );
 a96471a <=( (not A168)  and  A170 );
 a96474a <=( (not A200)  and  A199 );
 a96475a <=( a96474a  and  a96471a );
 a96478a <=( A202  and  A201 );
 a96481a <=( A266  and  (not A265) );
 a96482a <=( a96481a  and  a96478a );
 a96483a <=( a96482a  and  a96475a );
 a96486a <=( (not A268)  and  (not A267) );
 a96489a <=( A298  and  A269 );
 a96490a <=( a96489a  and  a96486a );
 a96493a <=( (not A300)  and  (not A299) );
 a96496a <=( A302  and  (not A301) );
 a96497a <=( a96496a  and  a96493a );
 a96498a <=( a96497a  and  a96490a );
 a96501a <=( (not A168)  and  A170 );
 a96504a <=( (not A200)  and  A199 );
 a96505a <=( a96504a  and  a96501a );
 a96508a <=( A202  and  A201 );
 a96511a <=( A266  and  (not A265) );
 a96512a <=( a96511a  and  a96508a );
 a96513a <=( a96512a  and  a96505a );
 a96516a <=( (not A268)  and  (not A267) );
 a96519a <=( (not A298)  and  A269 );
 a96520a <=( a96519a  and  a96516a );
 a96523a <=( (not A300)  and  A299 );
 a96526a <=( A302  and  (not A301) );
 a96527a <=( a96526a  and  a96523a );
 a96528a <=( a96527a  and  a96520a );
 a96531a <=( (not A168)  and  A170 );
 a96534a <=( (not A200)  and  A199 );
 a96535a <=( a96534a  and  a96531a );
 a96538a <=( A202  and  A201 );
 a96541a <=( (not A266)  and  A265 );
 a96542a <=( a96541a  and  a96538a );
 a96543a <=( a96542a  and  a96535a );
 a96546a <=( (not A268)  and  (not A267) );
 a96549a <=( A298  and  A269 );
 a96550a <=( a96549a  and  a96546a );
 a96553a <=( (not A300)  and  (not A299) );
 a96556a <=( A302  and  (not A301) );
 a96557a <=( a96556a  and  a96553a );
 a96558a <=( a96557a  and  a96550a );
 a96561a <=( (not A168)  and  A170 );
 a96564a <=( (not A200)  and  A199 );
 a96565a <=( a96564a  and  a96561a );
 a96568a <=( A202  and  A201 );
 a96571a <=( (not A266)  and  A265 );
 a96572a <=( a96571a  and  a96568a );
 a96573a <=( a96572a  and  a96565a );
 a96576a <=( (not A268)  and  (not A267) );
 a96579a <=( (not A298)  and  A269 );
 a96580a <=( a96579a  and  a96576a );
 a96583a <=( (not A300)  and  A299 );
 a96586a <=( A302  and  (not A301) );
 a96587a <=( a96586a  and  a96583a );
 a96588a <=( a96587a  and  a96580a );
 a96591a <=( (not A168)  and  A170 );
 a96594a <=( (not A200)  and  A199 );
 a96595a <=( a96594a  and  a96591a );
 a96598a <=( (not A203)  and  A201 );
 a96601a <=( A266  and  (not A265) );
 a96602a <=( a96601a  and  a96598a );
 a96603a <=( a96602a  and  a96595a );
 a96606a <=( (not A268)  and  (not A267) );
 a96609a <=( A298  and  A269 );
 a96610a <=( a96609a  and  a96606a );
 a96613a <=( (not A300)  and  (not A299) );
 a96616a <=( A302  and  (not A301) );
 a96617a <=( a96616a  and  a96613a );
 a96618a <=( a96617a  and  a96610a );
 a96621a <=( (not A168)  and  A170 );
 a96624a <=( (not A200)  and  A199 );
 a96625a <=( a96624a  and  a96621a );
 a96628a <=( (not A203)  and  A201 );
 a96631a <=( A266  and  (not A265) );
 a96632a <=( a96631a  and  a96628a );
 a96633a <=( a96632a  and  a96625a );
 a96636a <=( (not A268)  and  (not A267) );
 a96639a <=( (not A298)  and  A269 );
 a96640a <=( a96639a  and  a96636a );
 a96643a <=( (not A300)  and  A299 );
 a96646a <=( A302  and  (not A301) );
 a96647a <=( a96646a  and  a96643a );
 a96648a <=( a96647a  and  a96640a );
 a96651a <=( (not A168)  and  A170 );
 a96654a <=( (not A200)  and  A199 );
 a96655a <=( a96654a  and  a96651a );
 a96658a <=( (not A203)  and  A201 );
 a96661a <=( (not A266)  and  A265 );
 a96662a <=( a96661a  and  a96658a );
 a96663a <=( a96662a  and  a96655a );
 a96666a <=( (not A268)  and  (not A267) );
 a96669a <=( A298  and  A269 );
 a96670a <=( a96669a  and  a96666a );
 a96673a <=( (not A300)  and  (not A299) );
 a96676a <=( A302  and  (not A301) );
 a96677a <=( a96676a  and  a96673a );
 a96678a <=( a96677a  and  a96670a );
 a96681a <=( (not A168)  and  A170 );
 a96684a <=( (not A200)  and  A199 );
 a96685a <=( a96684a  and  a96681a );
 a96688a <=( (not A203)  and  A201 );
 a96691a <=( (not A266)  and  A265 );
 a96692a <=( a96691a  and  a96688a );
 a96693a <=( a96692a  and  a96685a );
 a96696a <=( (not A268)  and  (not A267) );
 a96699a <=( (not A298)  and  A269 );
 a96700a <=( a96699a  and  a96696a );
 a96703a <=( (not A300)  and  A299 );
 a96706a <=( A302  and  (not A301) );
 a96707a <=( a96706a  and  a96703a );
 a96708a <=( a96707a  and  a96700a );
 a96711a <=( (not A168)  and  A170 );
 a96714a <=( (not A200)  and  A199 );
 a96715a <=( a96714a  and  a96711a );
 a96718a <=( (not A202)  and  (not A201) );
 a96721a <=( (not A265)  and  A203 );
 a96722a <=( a96721a  and  a96718a );
 a96723a <=( a96722a  and  a96715a );
 a96726a <=( A267  and  A266 );
 a96729a <=( A298  and  A268 );
 a96730a <=( a96729a  and  a96726a );
 a96733a <=( (not A300)  and  (not A299) );
 a96736a <=( A302  and  (not A301) );
 a96737a <=( a96736a  and  a96733a );
 a96738a <=( a96737a  and  a96730a );
 a96741a <=( (not A168)  and  A170 );
 a96744a <=( (not A200)  and  A199 );
 a96745a <=( a96744a  and  a96741a );
 a96748a <=( (not A202)  and  (not A201) );
 a96751a <=( (not A265)  and  A203 );
 a96752a <=( a96751a  and  a96748a );
 a96753a <=( a96752a  and  a96745a );
 a96756a <=( A267  and  A266 );
 a96759a <=( (not A298)  and  A268 );
 a96760a <=( a96759a  and  a96756a );
 a96763a <=( (not A300)  and  A299 );
 a96766a <=( A302  and  (not A301) );
 a96767a <=( a96766a  and  a96763a );
 a96768a <=( a96767a  and  a96760a );
 a96771a <=( (not A168)  and  A170 );
 a96774a <=( (not A200)  and  A199 );
 a96775a <=( a96774a  and  a96771a );
 a96778a <=( (not A202)  and  (not A201) );
 a96781a <=( (not A265)  and  A203 );
 a96782a <=( a96781a  and  a96778a );
 a96783a <=( a96782a  and  a96775a );
 a96786a <=( A267  and  A266 );
 a96789a <=( A298  and  (not A269) );
 a96790a <=( a96789a  and  a96786a );
 a96793a <=( (not A300)  and  (not A299) );
 a96796a <=( A302  and  (not A301) );
 a96797a <=( a96796a  and  a96793a );
 a96798a <=( a96797a  and  a96790a );
 a96801a <=( (not A168)  and  A170 );
 a96804a <=( (not A200)  and  A199 );
 a96805a <=( a96804a  and  a96801a );
 a96808a <=( (not A202)  and  (not A201) );
 a96811a <=( (not A265)  and  A203 );
 a96812a <=( a96811a  and  a96808a );
 a96813a <=( a96812a  and  a96805a );
 a96816a <=( A267  and  A266 );
 a96819a <=( (not A298)  and  (not A269) );
 a96820a <=( a96819a  and  a96816a );
 a96823a <=( (not A300)  and  A299 );
 a96826a <=( A302  and  (not A301) );
 a96827a <=( a96826a  and  a96823a );
 a96828a <=( a96827a  and  a96820a );
 a96831a <=( (not A168)  and  A170 );
 a96834a <=( (not A200)  and  A199 );
 a96835a <=( a96834a  and  a96831a );
 a96838a <=( (not A202)  and  (not A201) );
 a96841a <=( (not A265)  and  A203 );
 a96842a <=( a96841a  and  a96838a );
 a96843a <=( a96842a  and  a96835a );
 a96846a <=( (not A267)  and  A266 );
 a96849a <=( A269  and  (not A268) );
 a96850a <=( a96849a  and  a96846a );
 a96853a <=( (not A299)  and  A298 );
 a96856a <=( A301  and  A300 );
 a96857a <=( a96856a  and  a96853a );
 a96858a <=( a96857a  and  a96850a );
 a96861a <=( (not A168)  and  A170 );
 a96864a <=( (not A200)  and  A199 );
 a96865a <=( a96864a  and  a96861a );
 a96868a <=( (not A202)  and  (not A201) );
 a96871a <=( (not A265)  and  A203 );
 a96872a <=( a96871a  and  a96868a );
 a96873a <=( a96872a  and  a96865a );
 a96876a <=( (not A267)  and  A266 );
 a96879a <=( A269  and  (not A268) );
 a96880a <=( a96879a  and  a96876a );
 a96883a <=( (not A299)  and  A298 );
 a96886a <=( (not A302)  and  A300 );
 a96887a <=( a96886a  and  a96883a );
 a96888a <=( a96887a  and  a96880a );
 a96891a <=( (not A168)  and  A170 );
 a96894a <=( (not A200)  and  A199 );
 a96895a <=( a96894a  and  a96891a );
 a96898a <=( (not A202)  and  (not A201) );
 a96901a <=( (not A265)  and  A203 );
 a96902a <=( a96901a  and  a96898a );
 a96903a <=( a96902a  and  a96895a );
 a96906a <=( (not A267)  and  A266 );
 a96909a <=( A269  and  (not A268) );
 a96910a <=( a96909a  and  a96906a );
 a96913a <=( A299  and  (not A298) );
 a96916a <=( A301  and  A300 );
 a96917a <=( a96916a  and  a96913a );
 a96918a <=( a96917a  and  a96910a );
 a96921a <=( (not A168)  and  A170 );
 a96924a <=( (not A200)  and  A199 );
 a96925a <=( a96924a  and  a96921a );
 a96928a <=( (not A202)  and  (not A201) );
 a96931a <=( (not A265)  and  A203 );
 a96932a <=( a96931a  and  a96928a );
 a96933a <=( a96932a  and  a96925a );
 a96936a <=( (not A267)  and  A266 );
 a96939a <=( A269  and  (not A268) );
 a96940a <=( a96939a  and  a96936a );
 a96943a <=( A299  and  (not A298) );
 a96946a <=( (not A302)  and  A300 );
 a96947a <=( a96946a  and  a96943a );
 a96948a <=( a96947a  and  a96940a );
 a96951a <=( (not A168)  and  A170 );
 a96954a <=( (not A200)  and  A199 );
 a96955a <=( a96954a  and  a96951a );
 a96958a <=( (not A202)  and  (not A201) );
 a96961a <=( A265  and  A203 );
 a96962a <=( a96961a  and  a96958a );
 a96963a <=( a96962a  and  a96955a );
 a96966a <=( A267  and  (not A266) );
 a96969a <=( A298  and  A268 );
 a96970a <=( a96969a  and  a96966a );
 a96973a <=( (not A300)  and  (not A299) );
 a96976a <=( A302  and  (not A301) );
 a96977a <=( a96976a  and  a96973a );
 a96978a <=( a96977a  and  a96970a );
 a96981a <=( (not A168)  and  A170 );
 a96984a <=( (not A200)  and  A199 );
 a96985a <=( a96984a  and  a96981a );
 a96988a <=( (not A202)  and  (not A201) );
 a96991a <=( A265  and  A203 );
 a96992a <=( a96991a  and  a96988a );
 a96993a <=( a96992a  and  a96985a );
 a96996a <=( A267  and  (not A266) );
 a96999a <=( (not A298)  and  A268 );
 a97000a <=( a96999a  and  a96996a );
 a97003a <=( (not A300)  and  A299 );
 a97006a <=( A302  and  (not A301) );
 a97007a <=( a97006a  and  a97003a );
 a97008a <=( a97007a  and  a97000a );
 a97011a <=( (not A168)  and  A170 );
 a97014a <=( (not A200)  and  A199 );
 a97015a <=( a97014a  and  a97011a );
 a97018a <=( (not A202)  and  (not A201) );
 a97021a <=( A265  and  A203 );
 a97022a <=( a97021a  and  a97018a );
 a97023a <=( a97022a  and  a97015a );
 a97026a <=( A267  and  (not A266) );
 a97029a <=( A298  and  (not A269) );
 a97030a <=( a97029a  and  a97026a );
 a97033a <=( (not A300)  and  (not A299) );
 a97036a <=( A302  and  (not A301) );
 a97037a <=( a97036a  and  a97033a );
 a97038a <=( a97037a  and  a97030a );
 a97041a <=( (not A168)  and  A170 );
 a97044a <=( (not A200)  and  A199 );
 a97045a <=( a97044a  and  a97041a );
 a97048a <=( (not A202)  and  (not A201) );
 a97051a <=( A265  and  A203 );
 a97052a <=( a97051a  and  a97048a );
 a97053a <=( a97052a  and  a97045a );
 a97056a <=( A267  and  (not A266) );
 a97059a <=( (not A298)  and  (not A269) );
 a97060a <=( a97059a  and  a97056a );
 a97063a <=( (not A300)  and  A299 );
 a97066a <=( A302  and  (not A301) );
 a97067a <=( a97066a  and  a97063a );
 a97068a <=( a97067a  and  a97060a );
 a97071a <=( (not A168)  and  A170 );
 a97074a <=( (not A200)  and  A199 );
 a97075a <=( a97074a  and  a97071a );
 a97078a <=( (not A202)  and  (not A201) );
 a97081a <=( A265  and  A203 );
 a97082a <=( a97081a  and  a97078a );
 a97083a <=( a97082a  and  a97075a );
 a97086a <=( (not A267)  and  (not A266) );
 a97089a <=( A269  and  (not A268) );
 a97090a <=( a97089a  and  a97086a );
 a97093a <=( (not A299)  and  A298 );
 a97096a <=( A301  and  A300 );
 a97097a <=( a97096a  and  a97093a );
 a97098a <=( a97097a  and  a97090a );
 a97101a <=( (not A168)  and  A170 );
 a97104a <=( (not A200)  and  A199 );
 a97105a <=( a97104a  and  a97101a );
 a97108a <=( (not A202)  and  (not A201) );
 a97111a <=( A265  and  A203 );
 a97112a <=( a97111a  and  a97108a );
 a97113a <=( a97112a  and  a97105a );
 a97116a <=( (not A267)  and  (not A266) );
 a97119a <=( A269  and  (not A268) );
 a97120a <=( a97119a  and  a97116a );
 a97123a <=( (not A299)  and  A298 );
 a97126a <=( (not A302)  and  A300 );
 a97127a <=( a97126a  and  a97123a );
 a97128a <=( a97127a  and  a97120a );
 a97131a <=( (not A168)  and  A170 );
 a97134a <=( (not A200)  and  A199 );
 a97135a <=( a97134a  and  a97131a );
 a97138a <=( (not A202)  and  (not A201) );
 a97141a <=( A265  and  A203 );
 a97142a <=( a97141a  and  a97138a );
 a97143a <=( a97142a  and  a97135a );
 a97146a <=( (not A267)  and  (not A266) );
 a97149a <=( A269  and  (not A268) );
 a97150a <=( a97149a  and  a97146a );
 a97153a <=( A299  and  (not A298) );
 a97156a <=( A301  and  A300 );
 a97157a <=( a97156a  and  a97153a );
 a97158a <=( a97157a  and  a97150a );
 a97161a <=( (not A168)  and  A170 );
 a97164a <=( (not A200)  and  A199 );
 a97165a <=( a97164a  and  a97161a );
 a97168a <=( (not A202)  and  (not A201) );
 a97171a <=( A265  and  A203 );
 a97172a <=( a97171a  and  a97168a );
 a97173a <=( a97172a  and  a97165a );
 a97176a <=( (not A267)  and  (not A266) );
 a97179a <=( A269  and  (not A268) );
 a97180a <=( a97179a  and  a97176a );
 a97183a <=( A299  and  (not A298) );
 a97186a <=( (not A302)  and  A300 );
 a97187a <=( a97186a  and  a97183a );
 a97188a <=( a97187a  and  a97180a );
 a97191a <=( (not A168)  and  A169 );
 a97194a <=( A200  and  (not A199) );
 a97195a <=( a97194a  and  a97191a );
 a97198a <=( A202  and  A201 );
 a97201a <=( A266  and  (not A265) );
 a97202a <=( a97201a  and  a97198a );
 a97203a <=( a97202a  and  a97195a );
 a97206a <=( (not A268)  and  (not A267) );
 a97209a <=( A298  and  A269 );
 a97210a <=( a97209a  and  a97206a );
 a97213a <=( (not A300)  and  (not A299) );
 a97216a <=( A302  and  (not A301) );
 a97217a <=( a97216a  and  a97213a );
 a97218a <=( a97217a  and  a97210a );
 a97221a <=( (not A168)  and  A169 );
 a97224a <=( A200  and  (not A199) );
 a97225a <=( a97224a  and  a97221a );
 a97228a <=( A202  and  A201 );
 a97231a <=( A266  and  (not A265) );
 a97232a <=( a97231a  and  a97228a );
 a97233a <=( a97232a  and  a97225a );
 a97236a <=( (not A268)  and  (not A267) );
 a97239a <=( (not A298)  and  A269 );
 a97240a <=( a97239a  and  a97236a );
 a97243a <=( (not A300)  and  A299 );
 a97246a <=( A302  and  (not A301) );
 a97247a <=( a97246a  and  a97243a );
 a97248a <=( a97247a  and  a97240a );
 a97251a <=( (not A168)  and  A169 );
 a97254a <=( A200  and  (not A199) );
 a97255a <=( a97254a  and  a97251a );
 a97258a <=( A202  and  A201 );
 a97261a <=( (not A266)  and  A265 );
 a97262a <=( a97261a  and  a97258a );
 a97263a <=( a97262a  and  a97255a );
 a97266a <=( (not A268)  and  (not A267) );
 a97269a <=( A298  and  A269 );
 a97270a <=( a97269a  and  a97266a );
 a97273a <=( (not A300)  and  (not A299) );
 a97276a <=( A302  and  (not A301) );
 a97277a <=( a97276a  and  a97273a );
 a97278a <=( a97277a  and  a97270a );
 a97281a <=( (not A168)  and  A169 );
 a97284a <=( A200  and  (not A199) );
 a97285a <=( a97284a  and  a97281a );
 a97288a <=( A202  and  A201 );
 a97291a <=( (not A266)  and  A265 );
 a97292a <=( a97291a  and  a97288a );
 a97293a <=( a97292a  and  a97285a );
 a97296a <=( (not A268)  and  (not A267) );
 a97299a <=( (not A298)  and  A269 );
 a97300a <=( a97299a  and  a97296a );
 a97303a <=( (not A300)  and  A299 );
 a97306a <=( A302  and  (not A301) );
 a97307a <=( a97306a  and  a97303a );
 a97308a <=( a97307a  and  a97300a );
 a97311a <=( (not A168)  and  A169 );
 a97314a <=( A200  and  (not A199) );
 a97315a <=( a97314a  and  a97311a );
 a97318a <=( (not A203)  and  A201 );
 a97321a <=( A266  and  (not A265) );
 a97322a <=( a97321a  and  a97318a );
 a97323a <=( a97322a  and  a97315a );
 a97326a <=( (not A268)  and  (not A267) );
 a97329a <=( A298  and  A269 );
 a97330a <=( a97329a  and  a97326a );
 a97333a <=( (not A300)  and  (not A299) );
 a97336a <=( A302  and  (not A301) );
 a97337a <=( a97336a  and  a97333a );
 a97338a <=( a97337a  and  a97330a );
 a97341a <=( (not A168)  and  A169 );
 a97344a <=( A200  and  (not A199) );
 a97345a <=( a97344a  and  a97341a );
 a97348a <=( (not A203)  and  A201 );
 a97351a <=( A266  and  (not A265) );
 a97352a <=( a97351a  and  a97348a );
 a97353a <=( a97352a  and  a97345a );
 a97356a <=( (not A268)  and  (not A267) );
 a97359a <=( (not A298)  and  A269 );
 a97360a <=( a97359a  and  a97356a );
 a97363a <=( (not A300)  and  A299 );
 a97366a <=( A302  and  (not A301) );
 a97367a <=( a97366a  and  a97363a );
 a97368a <=( a97367a  and  a97360a );
 a97371a <=( (not A168)  and  A169 );
 a97374a <=( A200  and  (not A199) );
 a97375a <=( a97374a  and  a97371a );
 a97378a <=( (not A203)  and  A201 );
 a97381a <=( (not A266)  and  A265 );
 a97382a <=( a97381a  and  a97378a );
 a97383a <=( a97382a  and  a97375a );
 a97386a <=( (not A268)  and  (not A267) );
 a97389a <=( A298  and  A269 );
 a97390a <=( a97389a  and  a97386a );
 a97393a <=( (not A300)  and  (not A299) );
 a97396a <=( A302  and  (not A301) );
 a97397a <=( a97396a  and  a97393a );
 a97398a <=( a97397a  and  a97390a );
 a97401a <=( (not A168)  and  A169 );
 a97404a <=( A200  and  (not A199) );
 a97405a <=( a97404a  and  a97401a );
 a97408a <=( (not A203)  and  A201 );
 a97411a <=( (not A266)  and  A265 );
 a97412a <=( a97411a  and  a97408a );
 a97413a <=( a97412a  and  a97405a );
 a97416a <=( (not A268)  and  (not A267) );
 a97419a <=( (not A298)  and  A269 );
 a97420a <=( a97419a  and  a97416a );
 a97423a <=( (not A300)  and  A299 );
 a97426a <=( A302  and  (not A301) );
 a97427a <=( a97426a  and  a97423a );
 a97428a <=( a97427a  and  a97420a );
 a97431a <=( (not A168)  and  A169 );
 a97434a <=( A200  and  (not A199) );
 a97435a <=( a97434a  and  a97431a );
 a97438a <=( (not A202)  and  (not A201) );
 a97441a <=( (not A265)  and  A203 );
 a97442a <=( a97441a  and  a97438a );
 a97443a <=( a97442a  and  a97435a );
 a97446a <=( A267  and  A266 );
 a97449a <=( A298  and  A268 );
 a97450a <=( a97449a  and  a97446a );
 a97453a <=( (not A300)  and  (not A299) );
 a97456a <=( A302  and  (not A301) );
 a97457a <=( a97456a  and  a97453a );
 a97458a <=( a97457a  and  a97450a );
 a97461a <=( (not A168)  and  A169 );
 a97464a <=( A200  and  (not A199) );
 a97465a <=( a97464a  and  a97461a );
 a97468a <=( (not A202)  and  (not A201) );
 a97471a <=( (not A265)  and  A203 );
 a97472a <=( a97471a  and  a97468a );
 a97473a <=( a97472a  and  a97465a );
 a97476a <=( A267  and  A266 );
 a97479a <=( (not A298)  and  A268 );
 a97480a <=( a97479a  and  a97476a );
 a97483a <=( (not A300)  and  A299 );
 a97486a <=( A302  and  (not A301) );
 a97487a <=( a97486a  and  a97483a );
 a97488a <=( a97487a  and  a97480a );
 a97491a <=( (not A168)  and  A169 );
 a97494a <=( A200  and  (not A199) );
 a97495a <=( a97494a  and  a97491a );
 a97498a <=( (not A202)  and  (not A201) );
 a97501a <=( (not A265)  and  A203 );
 a97502a <=( a97501a  and  a97498a );
 a97503a <=( a97502a  and  a97495a );
 a97506a <=( A267  and  A266 );
 a97509a <=( A298  and  (not A269) );
 a97510a <=( a97509a  and  a97506a );
 a97513a <=( (not A300)  and  (not A299) );
 a97516a <=( A302  and  (not A301) );
 a97517a <=( a97516a  and  a97513a );
 a97518a <=( a97517a  and  a97510a );
 a97521a <=( (not A168)  and  A169 );
 a97524a <=( A200  and  (not A199) );
 a97525a <=( a97524a  and  a97521a );
 a97528a <=( (not A202)  and  (not A201) );
 a97531a <=( (not A265)  and  A203 );
 a97532a <=( a97531a  and  a97528a );
 a97533a <=( a97532a  and  a97525a );
 a97536a <=( A267  and  A266 );
 a97539a <=( (not A298)  and  (not A269) );
 a97540a <=( a97539a  and  a97536a );
 a97543a <=( (not A300)  and  A299 );
 a97546a <=( A302  and  (not A301) );
 a97547a <=( a97546a  and  a97543a );
 a97548a <=( a97547a  and  a97540a );
 a97551a <=( (not A168)  and  A169 );
 a97554a <=( A200  and  (not A199) );
 a97555a <=( a97554a  and  a97551a );
 a97558a <=( (not A202)  and  (not A201) );
 a97561a <=( (not A265)  and  A203 );
 a97562a <=( a97561a  and  a97558a );
 a97563a <=( a97562a  and  a97555a );
 a97566a <=( (not A267)  and  A266 );
 a97569a <=( A269  and  (not A268) );
 a97570a <=( a97569a  and  a97566a );
 a97573a <=( (not A299)  and  A298 );
 a97576a <=( A301  and  A300 );
 a97577a <=( a97576a  and  a97573a );
 a97578a <=( a97577a  and  a97570a );
 a97581a <=( (not A168)  and  A169 );
 a97584a <=( A200  and  (not A199) );
 a97585a <=( a97584a  and  a97581a );
 a97588a <=( (not A202)  and  (not A201) );
 a97591a <=( (not A265)  and  A203 );
 a97592a <=( a97591a  and  a97588a );
 a97593a <=( a97592a  and  a97585a );
 a97596a <=( (not A267)  and  A266 );
 a97599a <=( A269  and  (not A268) );
 a97600a <=( a97599a  and  a97596a );
 a97603a <=( (not A299)  and  A298 );
 a97606a <=( (not A302)  and  A300 );
 a97607a <=( a97606a  and  a97603a );
 a97608a <=( a97607a  and  a97600a );
 a97611a <=( (not A168)  and  A169 );
 a97614a <=( A200  and  (not A199) );
 a97615a <=( a97614a  and  a97611a );
 a97618a <=( (not A202)  and  (not A201) );
 a97621a <=( (not A265)  and  A203 );
 a97622a <=( a97621a  and  a97618a );
 a97623a <=( a97622a  and  a97615a );
 a97626a <=( (not A267)  and  A266 );
 a97629a <=( A269  and  (not A268) );
 a97630a <=( a97629a  and  a97626a );
 a97633a <=( A299  and  (not A298) );
 a97636a <=( A301  and  A300 );
 a97637a <=( a97636a  and  a97633a );
 a97638a <=( a97637a  and  a97630a );
 a97641a <=( (not A168)  and  A169 );
 a97644a <=( A200  and  (not A199) );
 a97645a <=( a97644a  and  a97641a );
 a97648a <=( (not A202)  and  (not A201) );
 a97651a <=( (not A265)  and  A203 );
 a97652a <=( a97651a  and  a97648a );
 a97653a <=( a97652a  and  a97645a );
 a97656a <=( (not A267)  and  A266 );
 a97659a <=( A269  and  (not A268) );
 a97660a <=( a97659a  and  a97656a );
 a97663a <=( A299  and  (not A298) );
 a97666a <=( (not A302)  and  A300 );
 a97667a <=( a97666a  and  a97663a );
 a97668a <=( a97667a  and  a97660a );
 a97671a <=( (not A168)  and  A169 );
 a97674a <=( A200  and  (not A199) );
 a97675a <=( a97674a  and  a97671a );
 a97678a <=( (not A202)  and  (not A201) );
 a97681a <=( A265  and  A203 );
 a97682a <=( a97681a  and  a97678a );
 a97683a <=( a97682a  and  a97675a );
 a97686a <=( A267  and  (not A266) );
 a97689a <=( A298  and  A268 );
 a97690a <=( a97689a  and  a97686a );
 a97693a <=( (not A300)  and  (not A299) );
 a97696a <=( A302  and  (not A301) );
 a97697a <=( a97696a  and  a97693a );
 a97698a <=( a97697a  and  a97690a );
 a97701a <=( (not A168)  and  A169 );
 a97704a <=( A200  and  (not A199) );
 a97705a <=( a97704a  and  a97701a );
 a97708a <=( (not A202)  and  (not A201) );
 a97711a <=( A265  and  A203 );
 a97712a <=( a97711a  and  a97708a );
 a97713a <=( a97712a  and  a97705a );
 a97716a <=( A267  and  (not A266) );
 a97719a <=( (not A298)  and  A268 );
 a97720a <=( a97719a  and  a97716a );
 a97723a <=( (not A300)  and  A299 );
 a97726a <=( A302  and  (not A301) );
 a97727a <=( a97726a  and  a97723a );
 a97728a <=( a97727a  and  a97720a );
 a97731a <=( (not A168)  and  A169 );
 a97734a <=( A200  and  (not A199) );
 a97735a <=( a97734a  and  a97731a );
 a97738a <=( (not A202)  and  (not A201) );
 a97741a <=( A265  and  A203 );
 a97742a <=( a97741a  and  a97738a );
 a97743a <=( a97742a  and  a97735a );
 a97746a <=( A267  and  (not A266) );
 a97749a <=( A298  and  (not A269) );
 a97750a <=( a97749a  and  a97746a );
 a97753a <=( (not A300)  and  (not A299) );
 a97756a <=( A302  and  (not A301) );
 a97757a <=( a97756a  and  a97753a );
 a97758a <=( a97757a  and  a97750a );
 a97761a <=( (not A168)  and  A169 );
 a97764a <=( A200  and  (not A199) );
 a97765a <=( a97764a  and  a97761a );
 a97768a <=( (not A202)  and  (not A201) );
 a97771a <=( A265  and  A203 );
 a97772a <=( a97771a  and  a97768a );
 a97773a <=( a97772a  and  a97765a );
 a97776a <=( A267  and  (not A266) );
 a97779a <=( (not A298)  and  (not A269) );
 a97780a <=( a97779a  and  a97776a );
 a97783a <=( (not A300)  and  A299 );
 a97786a <=( A302  and  (not A301) );
 a97787a <=( a97786a  and  a97783a );
 a97788a <=( a97787a  and  a97780a );
 a97791a <=( (not A168)  and  A169 );
 a97794a <=( A200  and  (not A199) );
 a97795a <=( a97794a  and  a97791a );
 a97798a <=( (not A202)  and  (not A201) );
 a97801a <=( A265  and  A203 );
 a97802a <=( a97801a  and  a97798a );
 a97803a <=( a97802a  and  a97795a );
 a97806a <=( (not A267)  and  (not A266) );
 a97809a <=( A269  and  (not A268) );
 a97810a <=( a97809a  and  a97806a );
 a97813a <=( (not A299)  and  A298 );
 a97816a <=( A301  and  A300 );
 a97817a <=( a97816a  and  a97813a );
 a97818a <=( a97817a  and  a97810a );
 a97821a <=( (not A168)  and  A169 );
 a97824a <=( A200  and  (not A199) );
 a97825a <=( a97824a  and  a97821a );
 a97828a <=( (not A202)  and  (not A201) );
 a97831a <=( A265  and  A203 );
 a97832a <=( a97831a  and  a97828a );
 a97833a <=( a97832a  and  a97825a );
 a97836a <=( (not A267)  and  (not A266) );
 a97839a <=( A269  and  (not A268) );
 a97840a <=( a97839a  and  a97836a );
 a97843a <=( (not A299)  and  A298 );
 a97846a <=( (not A302)  and  A300 );
 a97847a <=( a97846a  and  a97843a );
 a97848a <=( a97847a  and  a97840a );
 a97851a <=( (not A168)  and  A169 );
 a97854a <=( A200  and  (not A199) );
 a97855a <=( a97854a  and  a97851a );
 a97858a <=( (not A202)  and  (not A201) );
 a97861a <=( A265  and  A203 );
 a97862a <=( a97861a  and  a97858a );
 a97863a <=( a97862a  and  a97855a );
 a97866a <=( (not A267)  and  (not A266) );
 a97869a <=( A269  and  (not A268) );
 a97870a <=( a97869a  and  a97866a );
 a97873a <=( A299  and  (not A298) );
 a97876a <=( A301  and  A300 );
 a97877a <=( a97876a  and  a97873a );
 a97878a <=( a97877a  and  a97870a );
 a97881a <=( (not A168)  and  A169 );
 a97884a <=( A200  and  (not A199) );
 a97885a <=( a97884a  and  a97881a );
 a97888a <=( (not A202)  and  (not A201) );
 a97891a <=( A265  and  A203 );
 a97892a <=( a97891a  and  a97888a );
 a97893a <=( a97892a  and  a97885a );
 a97896a <=( (not A267)  and  (not A266) );
 a97899a <=( A269  and  (not A268) );
 a97900a <=( a97899a  and  a97896a );
 a97903a <=( A299  and  (not A298) );
 a97906a <=( (not A302)  and  A300 );
 a97907a <=( a97906a  and  a97903a );
 a97908a <=( a97907a  and  a97900a );
 a97911a <=( (not A168)  and  A169 );
 a97914a <=( (not A200)  and  A199 );
 a97915a <=( a97914a  and  a97911a );
 a97918a <=( A202  and  A201 );
 a97921a <=( A266  and  (not A265) );
 a97922a <=( a97921a  and  a97918a );
 a97923a <=( a97922a  and  a97915a );
 a97926a <=( (not A268)  and  (not A267) );
 a97929a <=( A298  and  A269 );
 a97930a <=( a97929a  and  a97926a );
 a97933a <=( (not A300)  and  (not A299) );
 a97936a <=( A302  and  (not A301) );
 a97937a <=( a97936a  and  a97933a );
 a97938a <=( a97937a  and  a97930a );
 a97941a <=( (not A168)  and  A169 );
 a97944a <=( (not A200)  and  A199 );
 a97945a <=( a97944a  and  a97941a );
 a97948a <=( A202  and  A201 );
 a97951a <=( A266  and  (not A265) );
 a97952a <=( a97951a  and  a97948a );
 a97953a <=( a97952a  and  a97945a );
 a97956a <=( (not A268)  and  (not A267) );
 a97959a <=( (not A298)  and  A269 );
 a97960a <=( a97959a  and  a97956a );
 a97963a <=( (not A300)  and  A299 );
 a97966a <=( A302  and  (not A301) );
 a97967a <=( a97966a  and  a97963a );
 a97968a <=( a97967a  and  a97960a );
 a97971a <=( (not A168)  and  A169 );
 a97974a <=( (not A200)  and  A199 );
 a97975a <=( a97974a  and  a97971a );
 a97978a <=( A202  and  A201 );
 a97981a <=( (not A266)  and  A265 );
 a97982a <=( a97981a  and  a97978a );
 a97983a <=( a97982a  and  a97975a );
 a97986a <=( (not A268)  and  (not A267) );
 a97989a <=( A298  and  A269 );
 a97990a <=( a97989a  and  a97986a );
 a97993a <=( (not A300)  and  (not A299) );
 a97996a <=( A302  and  (not A301) );
 a97997a <=( a97996a  and  a97993a );
 a97998a <=( a97997a  and  a97990a );
 a98001a <=( (not A168)  and  A169 );
 a98004a <=( (not A200)  and  A199 );
 a98005a <=( a98004a  and  a98001a );
 a98008a <=( A202  and  A201 );
 a98011a <=( (not A266)  and  A265 );
 a98012a <=( a98011a  and  a98008a );
 a98013a <=( a98012a  and  a98005a );
 a98016a <=( (not A268)  and  (not A267) );
 a98019a <=( (not A298)  and  A269 );
 a98020a <=( a98019a  and  a98016a );
 a98023a <=( (not A300)  and  A299 );
 a98026a <=( A302  and  (not A301) );
 a98027a <=( a98026a  and  a98023a );
 a98028a <=( a98027a  and  a98020a );
 a98031a <=( (not A168)  and  A169 );
 a98034a <=( (not A200)  and  A199 );
 a98035a <=( a98034a  and  a98031a );
 a98038a <=( (not A203)  and  A201 );
 a98041a <=( A266  and  (not A265) );
 a98042a <=( a98041a  and  a98038a );
 a98043a <=( a98042a  and  a98035a );
 a98046a <=( (not A268)  and  (not A267) );
 a98049a <=( A298  and  A269 );
 a98050a <=( a98049a  and  a98046a );
 a98053a <=( (not A300)  and  (not A299) );
 a98056a <=( A302  and  (not A301) );
 a98057a <=( a98056a  and  a98053a );
 a98058a <=( a98057a  and  a98050a );
 a98061a <=( (not A168)  and  A169 );
 a98064a <=( (not A200)  and  A199 );
 a98065a <=( a98064a  and  a98061a );
 a98068a <=( (not A203)  and  A201 );
 a98071a <=( A266  and  (not A265) );
 a98072a <=( a98071a  and  a98068a );
 a98073a <=( a98072a  and  a98065a );
 a98076a <=( (not A268)  and  (not A267) );
 a98079a <=( (not A298)  and  A269 );
 a98080a <=( a98079a  and  a98076a );
 a98083a <=( (not A300)  and  A299 );
 a98086a <=( A302  and  (not A301) );
 a98087a <=( a98086a  and  a98083a );
 a98088a <=( a98087a  and  a98080a );
 a98091a <=( (not A168)  and  A169 );
 a98094a <=( (not A200)  and  A199 );
 a98095a <=( a98094a  and  a98091a );
 a98098a <=( (not A203)  and  A201 );
 a98101a <=( (not A266)  and  A265 );
 a98102a <=( a98101a  and  a98098a );
 a98103a <=( a98102a  and  a98095a );
 a98106a <=( (not A268)  and  (not A267) );
 a98109a <=( A298  and  A269 );
 a98110a <=( a98109a  and  a98106a );
 a98113a <=( (not A300)  and  (not A299) );
 a98116a <=( A302  and  (not A301) );
 a98117a <=( a98116a  and  a98113a );
 a98118a <=( a98117a  and  a98110a );
 a98121a <=( (not A168)  and  A169 );
 a98124a <=( (not A200)  and  A199 );
 a98125a <=( a98124a  and  a98121a );
 a98128a <=( (not A203)  and  A201 );
 a98131a <=( (not A266)  and  A265 );
 a98132a <=( a98131a  and  a98128a );
 a98133a <=( a98132a  and  a98125a );
 a98136a <=( (not A268)  and  (not A267) );
 a98139a <=( (not A298)  and  A269 );
 a98140a <=( a98139a  and  a98136a );
 a98143a <=( (not A300)  and  A299 );
 a98146a <=( A302  and  (not A301) );
 a98147a <=( a98146a  and  a98143a );
 a98148a <=( a98147a  and  a98140a );
 a98151a <=( (not A168)  and  A169 );
 a98154a <=( (not A200)  and  A199 );
 a98155a <=( a98154a  and  a98151a );
 a98158a <=( (not A202)  and  (not A201) );
 a98161a <=( (not A265)  and  A203 );
 a98162a <=( a98161a  and  a98158a );
 a98163a <=( a98162a  and  a98155a );
 a98166a <=( A267  and  A266 );
 a98169a <=( A298  and  A268 );
 a98170a <=( a98169a  and  a98166a );
 a98173a <=( (not A300)  and  (not A299) );
 a98176a <=( A302  and  (not A301) );
 a98177a <=( a98176a  and  a98173a );
 a98178a <=( a98177a  and  a98170a );
 a98181a <=( (not A168)  and  A169 );
 a98184a <=( (not A200)  and  A199 );
 a98185a <=( a98184a  and  a98181a );
 a98188a <=( (not A202)  and  (not A201) );
 a98191a <=( (not A265)  and  A203 );
 a98192a <=( a98191a  and  a98188a );
 a98193a <=( a98192a  and  a98185a );
 a98196a <=( A267  and  A266 );
 a98199a <=( (not A298)  and  A268 );
 a98200a <=( a98199a  and  a98196a );
 a98203a <=( (not A300)  and  A299 );
 a98206a <=( A302  and  (not A301) );
 a98207a <=( a98206a  and  a98203a );
 a98208a <=( a98207a  and  a98200a );
 a98211a <=( (not A168)  and  A169 );
 a98214a <=( (not A200)  and  A199 );
 a98215a <=( a98214a  and  a98211a );
 a98218a <=( (not A202)  and  (not A201) );
 a98221a <=( (not A265)  and  A203 );
 a98222a <=( a98221a  and  a98218a );
 a98223a <=( a98222a  and  a98215a );
 a98226a <=( A267  and  A266 );
 a98229a <=( A298  and  (not A269) );
 a98230a <=( a98229a  and  a98226a );
 a98233a <=( (not A300)  and  (not A299) );
 a98236a <=( A302  and  (not A301) );
 a98237a <=( a98236a  and  a98233a );
 a98238a <=( a98237a  and  a98230a );
 a98241a <=( (not A168)  and  A169 );
 a98244a <=( (not A200)  and  A199 );
 a98245a <=( a98244a  and  a98241a );
 a98248a <=( (not A202)  and  (not A201) );
 a98251a <=( (not A265)  and  A203 );
 a98252a <=( a98251a  and  a98248a );
 a98253a <=( a98252a  and  a98245a );
 a98256a <=( A267  and  A266 );
 a98259a <=( (not A298)  and  (not A269) );
 a98260a <=( a98259a  and  a98256a );
 a98263a <=( (not A300)  and  A299 );
 a98266a <=( A302  and  (not A301) );
 a98267a <=( a98266a  and  a98263a );
 a98268a <=( a98267a  and  a98260a );
 a98271a <=( (not A168)  and  A169 );
 a98274a <=( (not A200)  and  A199 );
 a98275a <=( a98274a  and  a98271a );
 a98278a <=( (not A202)  and  (not A201) );
 a98281a <=( (not A265)  and  A203 );
 a98282a <=( a98281a  and  a98278a );
 a98283a <=( a98282a  and  a98275a );
 a98286a <=( (not A267)  and  A266 );
 a98289a <=( A269  and  (not A268) );
 a98290a <=( a98289a  and  a98286a );
 a98293a <=( (not A299)  and  A298 );
 a98296a <=( A301  and  A300 );
 a98297a <=( a98296a  and  a98293a );
 a98298a <=( a98297a  and  a98290a );
 a98301a <=( (not A168)  and  A169 );
 a98304a <=( (not A200)  and  A199 );
 a98305a <=( a98304a  and  a98301a );
 a98308a <=( (not A202)  and  (not A201) );
 a98311a <=( (not A265)  and  A203 );
 a98312a <=( a98311a  and  a98308a );
 a98313a <=( a98312a  and  a98305a );
 a98316a <=( (not A267)  and  A266 );
 a98319a <=( A269  and  (not A268) );
 a98320a <=( a98319a  and  a98316a );
 a98323a <=( (not A299)  and  A298 );
 a98326a <=( (not A302)  and  A300 );
 a98327a <=( a98326a  and  a98323a );
 a98328a <=( a98327a  and  a98320a );
 a98331a <=( (not A168)  and  A169 );
 a98334a <=( (not A200)  and  A199 );
 a98335a <=( a98334a  and  a98331a );
 a98338a <=( (not A202)  and  (not A201) );
 a98341a <=( (not A265)  and  A203 );
 a98342a <=( a98341a  and  a98338a );
 a98343a <=( a98342a  and  a98335a );
 a98346a <=( (not A267)  and  A266 );
 a98349a <=( A269  and  (not A268) );
 a98350a <=( a98349a  and  a98346a );
 a98353a <=( A299  and  (not A298) );
 a98356a <=( A301  and  A300 );
 a98357a <=( a98356a  and  a98353a );
 a98358a <=( a98357a  and  a98350a );
 a98361a <=( (not A168)  and  A169 );
 a98364a <=( (not A200)  and  A199 );
 a98365a <=( a98364a  and  a98361a );
 a98368a <=( (not A202)  and  (not A201) );
 a98371a <=( (not A265)  and  A203 );
 a98372a <=( a98371a  and  a98368a );
 a98373a <=( a98372a  and  a98365a );
 a98376a <=( (not A267)  and  A266 );
 a98379a <=( A269  and  (not A268) );
 a98380a <=( a98379a  and  a98376a );
 a98383a <=( A299  and  (not A298) );
 a98386a <=( (not A302)  and  A300 );
 a98387a <=( a98386a  and  a98383a );
 a98388a <=( a98387a  and  a98380a );
 a98391a <=( (not A168)  and  A169 );
 a98394a <=( (not A200)  and  A199 );
 a98395a <=( a98394a  and  a98391a );
 a98398a <=( (not A202)  and  (not A201) );
 a98401a <=( A265  and  A203 );
 a98402a <=( a98401a  and  a98398a );
 a98403a <=( a98402a  and  a98395a );
 a98406a <=( A267  and  (not A266) );
 a98409a <=( A298  and  A268 );
 a98410a <=( a98409a  and  a98406a );
 a98413a <=( (not A300)  and  (not A299) );
 a98416a <=( A302  and  (not A301) );
 a98417a <=( a98416a  and  a98413a );
 a98418a <=( a98417a  and  a98410a );
 a98421a <=( (not A168)  and  A169 );
 a98424a <=( (not A200)  and  A199 );
 a98425a <=( a98424a  and  a98421a );
 a98428a <=( (not A202)  and  (not A201) );
 a98431a <=( A265  and  A203 );
 a98432a <=( a98431a  and  a98428a );
 a98433a <=( a98432a  and  a98425a );
 a98436a <=( A267  and  (not A266) );
 a98439a <=( (not A298)  and  A268 );
 a98440a <=( a98439a  and  a98436a );
 a98443a <=( (not A300)  and  A299 );
 a98446a <=( A302  and  (not A301) );
 a98447a <=( a98446a  and  a98443a );
 a98448a <=( a98447a  and  a98440a );
 a98451a <=( (not A168)  and  A169 );
 a98454a <=( (not A200)  and  A199 );
 a98455a <=( a98454a  and  a98451a );
 a98458a <=( (not A202)  and  (not A201) );
 a98461a <=( A265  and  A203 );
 a98462a <=( a98461a  and  a98458a );
 a98463a <=( a98462a  and  a98455a );
 a98466a <=( A267  and  (not A266) );
 a98469a <=( A298  and  (not A269) );
 a98470a <=( a98469a  and  a98466a );
 a98473a <=( (not A300)  and  (not A299) );
 a98476a <=( A302  and  (not A301) );
 a98477a <=( a98476a  and  a98473a );
 a98478a <=( a98477a  and  a98470a );
 a98481a <=( (not A168)  and  A169 );
 a98484a <=( (not A200)  and  A199 );
 a98485a <=( a98484a  and  a98481a );
 a98488a <=( (not A202)  and  (not A201) );
 a98491a <=( A265  and  A203 );
 a98492a <=( a98491a  and  a98488a );
 a98493a <=( a98492a  and  a98485a );
 a98496a <=( A267  and  (not A266) );
 a98499a <=( (not A298)  and  (not A269) );
 a98500a <=( a98499a  and  a98496a );
 a98503a <=( (not A300)  and  A299 );
 a98506a <=( A302  and  (not A301) );
 a98507a <=( a98506a  and  a98503a );
 a98508a <=( a98507a  and  a98500a );
 a98511a <=( (not A168)  and  A169 );
 a98514a <=( (not A200)  and  A199 );
 a98515a <=( a98514a  and  a98511a );
 a98518a <=( (not A202)  and  (not A201) );
 a98521a <=( A265  and  A203 );
 a98522a <=( a98521a  and  a98518a );
 a98523a <=( a98522a  and  a98515a );
 a98526a <=( (not A267)  and  (not A266) );
 a98529a <=( A269  and  (not A268) );
 a98530a <=( a98529a  and  a98526a );
 a98533a <=( (not A299)  and  A298 );
 a98536a <=( A301  and  A300 );
 a98537a <=( a98536a  and  a98533a );
 a98538a <=( a98537a  and  a98530a );
 a98541a <=( (not A168)  and  A169 );
 a98544a <=( (not A200)  and  A199 );
 a98545a <=( a98544a  and  a98541a );
 a98548a <=( (not A202)  and  (not A201) );
 a98551a <=( A265  and  A203 );
 a98552a <=( a98551a  and  a98548a );
 a98553a <=( a98552a  and  a98545a );
 a98556a <=( (not A267)  and  (not A266) );
 a98559a <=( A269  and  (not A268) );
 a98560a <=( a98559a  and  a98556a );
 a98563a <=( (not A299)  and  A298 );
 a98566a <=( (not A302)  and  A300 );
 a98567a <=( a98566a  and  a98563a );
 a98568a <=( a98567a  and  a98560a );
 a98571a <=( (not A168)  and  A169 );
 a98574a <=( (not A200)  and  A199 );
 a98575a <=( a98574a  and  a98571a );
 a98578a <=( (not A202)  and  (not A201) );
 a98581a <=( A265  and  A203 );
 a98582a <=( a98581a  and  a98578a );
 a98583a <=( a98582a  and  a98575a );
 a98586a <=( (not A267)  and  (not A266) );
 a98589a <=( A269  and  (not A268) );
 a98590a <=( a98589a  and  a98586a );
 a98593a <=( A299  and  (not A298) );
 a98596a <=( A301  and  A300 );
 a98597a <=( a98596a  and  a98593a );
 a98598a <=( a98597a  and  a98590a );
 a98601a <=( (not A168)  and  A169 );
 a98604a <=( (not A200)  and  A199 );
 a98605a <=( a98604a  and  a98601a );
 a98608a <=( (not A202)  and  (not A201) );
 a98611a <=( A265  and  A203 );
 a98612a <=( a98611a  and  a98608a );
 a98613a <=( a98612a  and  a98605a );
 a98616a <=( (not A267)  and  (not A266) );
 a98619a <=( A269  and  (not A268) );
 a98620a <=( a98619a  and  a98616a );
 a98623a <=( A299  and  (not A298) );
 a98626a <=( (not A302)  and  A300 );
 a98627a <=( a98626a  and  a98623a );
 a98628a <=( a98627a  and  a98620a );
 a98631a <=( (not A169)  and  (not A170) );
 a98634a <=( (not A199)  and  A168 );
 a98635a <=( a98634a  and  a98631a );
 a98638a <=( A201  and  A200 );
 a98641a <=( (not A265)  and  A202 );
 a98642a <=( a98641a  and  a98638a );
 a98643a <=( a98642a  and  a98635a );
 a98646a <=( A267  and  A266 );
 a98649a <=( A298  and  A268 );
 a98650a <=( a98649a  and  a98646a );
 a98653a <=( (not A300)  and  (not A299) );
 a98656a <=( A302  and  (not A301) );
 a98657a <=( a98656a  and  a98653a );
 a98658a <=( a98657a  and  a98650a );
 a98661a <=( (not A169)  and  (not A170) );
 a98664a <=( (not A199)  and  A168 );
 a98665a <=( a98664a  and  a98661a );
 a98668a <=( A201  and  A200 );
 a98671a <=( (not A265)  and  A202 );
 a98672a <=( a98671a  and  a98668a );
 a98673a <=( a98672a  and  a98665a );
 a98676a <=( A267  and  A266 );
 a98679a <=( (not A298)  and  A268 );
 a98680a <=( a98679a  and  a98676a );
 a98683a <=( (not A300)  and  A299 );
 a98686a <=( A302  and  (not A301) );
 a98687a <=( a98686a  and  a98683a );
 a98688a <=( a98687a  and  a98680a );
 a98691a <=( (not A169)  and  (not A170) );
 a98694a <=( (not A199)  and  A168 );
 a98695a <=( a98694a  and  a98691a );
 a98698a <=( A201  and  A200 );
 a98701a <=( (not A265)  and  A202 );
 a98702a <=( a98701a  and  a98698a );
 a98703a <=( a98702a  and  a98695a );
 a98706a <=( A267  and  A266 );
 a98709a <=( A298  and  (not A269) );
 a98710a <=( a98709a  and  a98706a );
 a98713a <=( (not A300)  and  (not A299) );
 a98716a <=( A302  and  (not A301) );
 a98717a <=( a98716a  and  a98713a );
 a98718a <=( a98717a  and  a98710a );
 a98721a <=( (not A169)  and  (not A170) );
 a98724a <=( (not A199)  and  A168 );
 a98725a <=( a98724a  and  a98721a );
 a98728a <=( A201  and  A200 );
 a98731a <=( (not A265)  and  A202 );
 a98732a <=( a98731a  and  a98728a );
 a98733a <=( a98732a  and  a98725a );
 a98736a <=( A267  and  A266 );
 a98739a <=( (not A298)  and  (not A269) );
 a98740a <=( a98739a  and  a98736a );
 a98743a <=( (not A300)  and  A299 );
 a98746a <=( A302  and  (not A301) );
 a98747a <=( a98746a  and  a98743a );
 a98748a <=( a98747a  and  a98740a );
 a98751a <=( (not A169)  and  (not A170) );
 a98754a <=( (not A199)  and  A168 );
 a98755a <=( a98754a  and  a98751a );
 a98758a <=( A201  and  A200 );
 a98761a <=( (not A265)  and  A202 );
 a98762a <=( a98761a  and  a98758a );
 a98763a <=( a98762a  and  a98755a );
 a98766a <=( (not A267)  and  A266 );
 a98769a <=( A269  and  (not A268) );
 a98770a <=( a98769a  and  a98766a );
 a98773a <=( (not A299)  and  A298 );
 a98776a <=( A301  and  A300 );
 a98777a <=( a98776a  and  a98773a );
 a98778a <=( a98777a  and  a98770a );
 a98781a <=( (not A169)  and  (not A170) );
 a98784a <=( (not A199)  and  A168 );
 a98785a <=( a98784a  and  a98781a );
 a98788a <=( A201  and  A200 );
 a98791a <=( (not A265)  and  A202 );
 a98792a <=( a98791a  and  a98788a );
 a98793a <=( a98792a  and  a98785a );
 a98796a <=( (not A267)  and  A266 );
 a98799a <=( A269  and  (not A268) );
 a98800a <=( a98799a  and  a98796a );
 a98803a <=( (not A299)  and  A298 );
 a98806a <=( (not A302)  and  A300 );
 a98807a <=( a98806a  and  a98803a );
 a98808a <=( a98807a  and  a98800a );
 a98811a <=( (not A169)  and  (not A170) );
 a98814a <=( (not A199)  and  A168 );
 a98815a <=( a98814a  and  a98811a );
 a98818a <=( A201  and  A200 );
 a98821a <=( (not A265)  and  A202 );
 a98822a <=( a98821a  and  a98818a );
 a98823a <=( a98822a  and  a98815a );
 a98826a <=( (not A267)  and  A266 );
 a98829a <=( A269  and  (not A268) );
 a98830a <=( a98829a  and  a98826a );
 a98833a <=( A299  and  (not A298) );
 a98836a <=( A301  and  A300 );
 a98837a <=( a98836a  and  a98833a );
 a98838a <=( a98837a  and  a98830a );
 a98841a <=( (not A169)  and  (not A170) );
 a98844a <=( (not A199)  and  A168 );
 a98845a <=( a98844a  and  a98841a );
 a98848a <=( A201  and  A200 );
 a98851a <=( (not A265)  and  A202 );
 a98852a <=( a98851a  and  a98848a );
 a98853a <=( a98852a  and  a98845a );
 a98856a <=( (not A267)  and  A266 );
 a98859a <=( A269  and  (not A268) );
 a98860a <=( a98859a  and  a98856a );
 a98863a <=( A299  and  (not A298) );
 a98866a <=( (not A302)  and  A300 );
 a98867a <=( a98866a  and  a98863a );
 a98868a <=( a98867a  and  a98860a );
 a98871a <=( (not A169)  and  (not A170) );
 a98874a <=( (not A199)  and  A168 );
 a98875a <=( a98874a  and  a98871a );
 a98878a <=( A201  and  A200 );
 a98881a <=( A265  and  A202 );
 a98882a <=( a98881a  and  a98878a );
 a98883a <=( a98882a  and  a98875a );
 a98886a <=( A267  and  (not A266) );
 a98889a <=( A298  and  A268 );
 a98890a <=( a98889a  and  a98886a );
 a98893a <=( (not A300)  and  (not A299) );
 a98896a <=( A302  and  (not A301) );
 a98897a <=( a98896a  and  a98893a );
 a98898a <=( a98897a  and  a98890a );
 a98901a <=( (not A169)  and  (not A170) );
 a98904a <=( (not A199)  and  A168 );
 a98905a <=( a98904a  and  a98901a );
 a98908a <=( A201  and  A200 );
 a98911a <=( A265  and  A202 );
 a98912a <=( a98911a  and  a98908a );
 a98913a <=( a98912a  and  a98905a );
 a98916a <=( A267  and  (not A266) );
 a98919a <=( (not A298)  and  A268 );
 a98920a <=( a98919a  and  a98916a );
 a98923a <=( (not A300)  and  A299 );
 a98926a <=( A302  and  (not A301) );
 a98927a <=( a98926a  and  a98923a );
 a98928a <=( a98927a  and  a98920a );
 a98931a <=( (not A169)  and  (not A170) );
 a98934a <=( (not A199)  and  A168 );
 a98935a <=( a98934a  and  a98931a );
 a98938a <=( A201  and  A200 );
 a98941a <=( A265  and  A202 );
 a98942a <=( a98941a  and  a98938a );
 a98943a <=( a98942a  and  a98935a );
 a98946a <=( A267  and  (not A266) );
 a98949a <=( A298  and  (not A269) );
 a98950a <=( a98949a  and  a98946a );
 a98953a <=( (not A300)  and  (not A299) );
 a98956a <=( A302  and  (not A301) );
 a98957a <=( a98956a  and  a98953a );
 a98958a <=( a98957a  and  a98950a );
 a98961a <=( (not A169)  and  (not A170) );
 a98964a <=( (not A199)  and  A168 );
 a98965a <=( a98964a  and  a98961a );
 a98968a <=( A201  and  A200 );
 a98971a <=( A265  and  A202 );
 a98972a <=( a98971a  and  a98968a );
 a98973a <=( a98972a  and  a98965a );
 a98976a <=( A267  and  (not A266) );
 a98979a <=( (not A298)  and  (not A269) );
 a98980a <=( a98979a  and  a98976a );
 a98983a <=( (not A300)  and  A299 );
 a98986a <=( A302  and  (not A301) );
 a98987a <=( a98986a  and  a98983a );
 a98988a <=( a98987a  and  a98980a );
 a98991a <=( (not A169)  and  (not A170) );
 a98994a <=( (not A199)  and  A168 );
 a98995a <=( a98994a  and  a98991a );
 a98998a <=( A201  and  A200 );
 a99001a <=( A265  and  A202 );
 a99002a <=( a99001a  and  a98998a );
 a99003a <=( a99002a  and  a98995a );
 a99006a <=( (not A267)  and  (not A266) );
 a99009a <=( A269  and  (not A268) );
 a99010a <=( a99009a  and  a99006a );
 a99013a <=( (not A299)  and  A298 );
 a99016a <=( A301  and  A300 );
 a99017a <=( a99016a  and  a99013a );
 a99018a <=( a99017a  and  a99010a );
 a99021a <=( (not A169)  and  (not A170) );
 a99024a <=( (not A199)  and  A168 );
 a99025a <=( a99024a  and  a99021a );
 a99028a <=( A201  and  A200 );
 a99031a <=( A265  and  A202 );
 a99032a <=( a99031a  and  a99028a );
 a99033a <=( a99032a  and  a99025a );
 a99036a <=( (not A267)  and  (not A266) );
 a99039a <=( A269  and  (not A268) );
 a99040a <=( a99039a  and  a99036a );
 a99043a <=( (not A299)  and  A298 );
 a99046a <=( (not A302)  and  A300 );
 a99047a <=( a99046a  and  a99043a );
 a99048a <=( a99047a  and  a99040a );
 a99051a <=( (not A169)  and  (not A170) );
 a99054a <=( (not A199)  and  A168 );
 a99055a <=( a99054a  and  a99051a );
 a99058a <=( A201  and  A200 );
 a99061a <=( A265  and  A202 );
 a99062a <=( a99061a  and  a99058a );
 a99063a <=( a99062a  and  a99055a );
 a99066a <=( (not A267)  and  (not A266) );
 a99069a <=( A269  and  (not A268) );
 a99070a <=( a99069a  and  a99066a );
 a99073a <=( A299  and  (not A298) );
 a99076a <=( A301  and  A300 );
 a99077a <=( a99076a  and  a99073a );
 a99078a <=( a99077a  and  a99070a );
 a99081a <=( (not A169)  and  (not A170) );
 a99084a <=( (not A199)  and  A168 );
 a99085a <=( a99084a  and  a99081a );
 a99088a <=( A201  and  A200 );
 a99091a <=( A265  and  A202 );
 a99092a <=( a99091a  and  a99088a );
 a99093a <=( a99092a  and  a99085a );
 a99096a <=( (not A267)  and  (not A266) );
 a99099a <=( A269  and  (not A268) );
 a99100a <=( a99099a  and  a99096a );
 a99103a <=( A299  and  (not A298) );
 a99106a <=( (not A302)  and  A300 );
 a99107a <=( a99106a  and  a99103a );
 a99108a <=( a99107a  and  a99100a );
 a99111a <=( (not A169)  and  (not A170) );
 a99114a <=( (not A199)  and  A168 );
 a99115a <=( a99114a  and  a99111a );
 a99118a <=( A201  and  A200 );
 a99121a <=( (not A265)  and  (not A203) );
 a99122a <=( a99121a  and  a99118a );
 a99123a <=( a99122a  and  a99115a );
 a99126a <=( A267  and  A266 );
 a99129a <=( A298  and  A268 );
 a99130a <=( a99129a  and  a99126a );
 a99133a <=( (not A300)  and  (not A299) );
 a99136a <=( A302  and  (not A301) );
 a99137a <=( a99136a  and  a99133a );
 a99138a <=( a99137a  and  a99130a );
 a99141a <=( (not A169)  and  (not A170) );
 a99144a <=( (not A199)  and  A168 );
 a99145a <=( a99144a  and  a99141a );
 a99148a <=( A201  and  A200 );
 a99151a <=( (not A265)  and  (not A203) );
 a99152a <=( a99151a  and  a99148a );
 a99153a <=( a99152a  and  a99145a );
 a99156a <=( A267  and  A266 );
 a99159a <=( (not A298)  and  A268 );
 a99160a <=( a99159a  and  a99156a );
 a99163a <=( (not A300)  and  A299 );
 a99166a <=( A302  and  (not A301) );
 a99167a <=( a99166a  and  a99163a );
 a99168a <=( a99167a  and  a99160a );
 a99171a <=( (not A169)  and  (not A170) );
 a99174a <=( (not A199)  and  A168 );
 a99175a <=( a99174a  and  a99171a );
 a99178a <=( A201  and  A200 );
 a99181a <=( (not A265)  and  (not A203) );
 a99182a <=( a99181a  and  a99178a );
 a99183a <=( a99182a  and  a99175a );
 a99186a <=( A267  and  A266 );
 a99189a <=( A298  and  (not A269) );
 a99190a <=( a99189a  and  a99186a );
 a99193a <=( (not A300)  and  (not A299) );
 a99196a <=( A302  and  (not A301) );
 a99197a <=( a99196a  and  a99193a );
 a99198a <=( a99197a  and  a99190a );
 a99201a <=( (not A169)  and  (not A170) );
 a99204a <=( (not A199)  and  A168 );
 a99205a <=( a99204a  and  a99201a );
 a99208a <=( A201  and  A200 );
 a99211a <=( (not A265)  and  (not A203) );
 a99212a <=( a99211a  and  a99208a );
 a99213a <=( a99212a  and  a99205a );
 a99216a <=( A267  and  A266 );
 a99219a <=( (not A298)  and  (not A269) );
 a99220a <=( a99219a  and  a99216a );
 a99223a <=( (not A300)  and  A299 );
 a99226a <=( A302  and  (not A301) );
 a99227a <=( a99226a  and  a99223a );
 a99228a <=( a99227a  and  a99220a );
 a99231a <=( (not A169)  and  (not A170) );
 a99234a <=( (not A199)  and  A168 );
 a99235a <=( a99234a  and  a99231a );
 a99238a <=( A201  and  A200 );
 a99241a <=( (not A265)  and  (not A203) );
 a99242a <=( a99241a  and  a99238a );
 a99243a <=( a99242a  and  a99235a );
 a99246a <=( (not A267)  and  A266 );
 a99249a <=( A269  and  (not A268) );
 a99250a <=( a99249a  and  a99246a );
 a99253a <=( (not A299)  and  A298 );
 a99256a <=( A301  and  A300 );
 a99257a <=( a99256a  and  a99253a );
 a99258a <=( a99257a  and  a99250a );
 a99261a <=( (not A169)  and  (not A170) );
 a99264a <=( (not A199)  and  A168 );
 a99265a <=( a99264a  and  a99261a );
 a99268a <=( A201  and  A200 );
 a99271a <=( (not A265)  and  (not A203) );
 a99272a <=( a99271a  and  a99268a );
 a99273a <=( a99272a  and  a99265a );
 a99276a <=( (not A267)  and  A266 );
 a99279a <=( A269  and  (not A268) );
 a99280a <=( a99279a  and  a99276a );
 a99283a <=( (not A299)  and  A298 );
 a99286a <=( (not A302)  and  A300 );
 a99287a <=( a99286a  and  a99283a );
 a99288a <=( a99287a  and  a99280a );
 a99291a <=( (not A169)  and  (not A170) );
 a99294a <=( (not A199)  and  A168 );
 a99295a <=( a99294a  and  a99291a );
 a99298a <=( A201  and  A200 );
 a99301a <=( (not A265)  and  (not A203) );
 a99302a <=( a99301a  and  a99298a );
 a99303a <=( a99302a  and  a99295a );
 a99306a <=( (not A267)  and  A266 );
 a99309a <=( A269  and  (not A268) );
 a99310a <=( a99309a  and  a99306a );
 a99313a <=( A299  and  (not A298) );
 a99316a <=( A301  and  A300 );
 a99317a <=( a99316a  and  a99313a );
 a99318a <=( a99317a  and  a99310a );
 a99321a <=( (not A169)  and  (not A170) );
 a99324a <=( (not A199)  and  A168 );
 a99325a <=( a99324a  and  a99321a );
 a99328a <=( A201  and  A200 );
 a99331a <=( (not A265)  and  (not A203) );
 a99332a <=( a99331a  and  a99328a );
 a99333a <=( a99332a  and  a99325a );
 a99336a <=( (not A267)  and  A266 );
 a99339a <=( A269  and  (not A268) );
 a99340a <=( a99339a  and  a99336a );
 a99343a <=( A299  and  (not A298) );
 a99346a <=( (not A302)  and  A300 );
 a99347a <=( a99346a  and  a99343a );
 a99348a <=( a99347a  and  a99340a );
 a99351a <=( (not A169)  and  (not A170) );
 a99354a <=( (not A199)  and  A168 );
 a99355a <=( a99354a  and  a99351a );
 a99358a <=( A201  and  A200 );
 a99361a <=( A265  and  (not A203) );
 a99362a <=( a99361a  and  a99358a );
 a99363a <=( a99362a  and  a99355a );
 a99366a <=( A267  and  (not A266) );
 a99369a <=( A298  and  A268 );
 a99370a <=( a99369a  and  a99366a );
 a99373a <=( (not A300)  and  (not A299) );
 a99376a <=( A302  and  (not A301) );
 a99377a <=( a99376a  and  a99373a );
 a99378a <=( a99377a  and  a99370a );
 a99381a <=( (not A169)  and  (not A170) );
 a99384a <=( (not A199)  and  A168 );
 a99385a <=( a99384a  and  a99381a );
 a99388a <=( A201  and  A200 );
 a99391a <=( A265  and  (not A203) );
 a99392a <=( a99391a  and  a99388a );
 a99393a <=( a99392a  and  a99385a );
 a99396a <=( A267  and  (not A266) );
 a99399a <=( (not A298)  and  A268 );
 a99400a <=( a99399a  and  a99396a );
 a99403a <=( (not A300)  and  A299 );
 a99406a <=( A302  and  (not A301) );
 a99407a <=( a99406a  and  a99403a );
 a99408a <=( a99407a  and  a99400a );
 a99411a <=( (not A169)  and  (not A170) );
 a99414a <=( (not A199)  and  A168 );
 a99415a <=( a99414a  and  a99411a );
 a99418a <=( A201  and  A200 );
 a99421a <=( A265  and  (not A203) );
 a99422a <=( a99421a  and  a99418a );
 a99423a <=( a99422a  and  a99415a );
 a99426a <=( A267  and  (not A266) );
 a99429a <=( A298  and  (not A269) );
 a99430a <=( a99429a  and  a99426a );
 a99433a <=( (not A300)  and  (not A299) );
 a99436a <=( A302  and  (not A301) );
 a99437a <=( a99436a  and  a99433a );
 a99438a <=( a99437a  and  a99430a );
 a99441a <=( (not A169)  and  (not A170) );
 a99444a <=( (not A199)  and  A168 );
 a99445a <=( a99444a  and  a99441a );
 a99448a <=( A201  and  A200 );
 a99451a <=( A265  and  (not A203) );
 a99452a <=( a99451a  and  a99448a );
 a99453a <=( a99452a  and  a99445a );
 a99456a <=( A267  and  (not A266) );
 a99459a <=( (not A298)  and  (not A269) );
 a99460a <=( a99459a  and  a99456a );
 a99463a <=( (not A300)  and  A299 );
 a99466a <=( A302  and  (not A301) );
 a99467a <=( a99466a  and  a99463a );
 a99468a <=( a99467a  and  a99460a );
 a99471a <=( (not A169)  and  (not A170) );
 a99474a <=( (not A199)  and  A168 );
 a99475a <=( a99474a  and  a99471a );
 a99478a <=( A201  and  A200 );
 a99481a <=( A265  and  (not A203) );
 a99482a <=( a99481a  and  a99478a );
 a99483a <=( a99482a  and  a99475a );
 a99486a <=( (not A267)  and  (not A266) );
 a99489a <=( A269  and  (not A268) );
 a99490a <=( a99489a  and  a99486a );
 a99493a <=( (not A299)  and  A298 );
 a99496a <=( A301  and  A300 );
 a99497a <=( a99496a  and  a99493a );
 a99498a <=( a99497a  and  a99490a );
 a99501a <=( (not A169)  and  (not A170) );
 a99504a <=( (not A199)  and  A168 );
 a99505a <=( a99504a  and  a99501a );
 a99508a <=( A201  and  A200 );
 a99511a <=( A265  and  (not A203) );
 a99512a <=( a99511a  and  a99508a );
 a99513a <=( a99512a  and  a99505a );
 a99516a <=( (not A267)  and  (not A266) );
 a99519a <=( A269  and  (not A268) );
 a99520a <=( a99519a  and  a99516a );
 a99523a <=( (not A299)  and  A298 );
 a99526a <=( (not A302)  and  A300 );
 a99527a <=( a99526a  and  a99523a );
 a99528a <=( a99527a  and  a99520a );
 a99531a <=( (not A169)  and  (not A170) );
 a99534a <=( (not A199)  and  A168 );
 a99535a <=( a99534a  and  a99531a );
 a99538a <=( A201  and  A200 );
 a99541a <=( A265  and  (not A203) );
 a99542a <=( a99541a  and  a99538a );
 a99543a <=( a99542a  and  a99535a );
 a99546a <=( (not A267)  and  (not A266) );
 a99549a <=( A269  and  (not A268) );
 a99550a <=( a99549a  and  a99546a );
 a99553a <=( A299  and  (not A298) );
 a99556a <=( A301  and  A300 );
 a99557a <=( a99556a  and  a99553a );
 a99558a <=( a99557a  and  a99550a );
 a99561a <=( (not A169)  and  (not A170) );
 a99564a <=( (not A199)  and  A168 );
 a99565a <=( a99564a  and  a99561a );
 a99568a <=( A201  and  A200 );
 a99571a <=( A265  and  (not A203) );
 a99572a <=( a99571a  and  a99568a );
 a99573a <=( a99572a  and  a99565a );
 a99576a <=( (not A267)  and  (not A266) );
 a99579a <=( A269  and  (not A268) );
 a99580a <=( a99579a  and  a99576a );
 a99583a <=( A299  and  (not A298) );
 a99586a <=( (not A302)  and  A300 );
 a99587a <=( a99586a  and  a99583a );
 a99588a <=( a99587a  and  a99580a );
 a99591a <=( (not A169)  and  (not A170) );
 a99594a <=( (not A199)  and  A168 );
 a99595a <=( a99594a  and  a99591a );
 a99598a <=( (not A201)  and  A200 );
 a99601a <=( A203  and  (not A202) );
 a99602a <=( a99601a  and  a99598a );
 a99603a <=( a99602a  and  a99595a );
 a99606a <=( A266  and  (not A265) );
 a99609a <=( A268  and  A267 );
 a99610a <=( a99609a  and  a99606a );
 a99613a <=( (not A299)  and  A298 );
 a99616a <=( A301  and  A300 );
 a99617a <=( a99616a  and  a99613a );
 a99618a <=( a99617a  and  a99610a );
 a99621a <=( (not A169)  and  (not A170) );
 a99624a <=( (not A199)  and  A168 );
 a99625a <=( a99624a  and  a99621a );
 a99628a <=( (not A201)  and  A200 );
 a99631a <=( A203  and  (not A202) );
 a99632a <=( a99631a  and  a99628a );
 a99633a <=( a99632a  and  a99625a );
 a99636a <=( A266  and  (not A265) );
 a99639a <=( A268  and  A267 );
 a99640a <=( a99639a  and  a99636a );
 a99643a <=( (not A299)  and  A298 );
 a99646a <=( (not A302)  and  A300 );
 a99647a <=( a99646a  and  a99643a );
 a99648a <=( a99647a  and  a99640a );
 a99651a <=( (not A169)  and  (not A170) );
 a99654a <=( (not A199)  and  A168 );
 a99655a <=( a99654a  and  a99651a );
 a99658a <=( (not A201)  and  A200 );
 a99661a <=( A203  and  (not A202) );
 a99662a <=( a99661a  and  a99658a );
 a99663a <=( a99662a  and  a99655a );
 a99666a <=( A266  and  (not A265) );
 a99669a <=( A268  and  A267 );
 a99670a <=( a99669a  and  a99666a );
 a99673a <=( A299  and  (not A298) );
 a99676a <=( A301  and  A300 );
 a99677a <=( a99676a  and  a99673a );
 a99678a <=( a99677a  and  a99670a );
 a99681a <=( (not A169)  and  (not A170) );
 a99684a <=( (not A199)  and  A168 );
 a99685a <=( a99684a  and  a99681a );
 a99688a <=( (not A201)  and  A200 );
 a99691a <=( A203  and  (not A202) );
 a99692a <=( a99691a  and  a99688a );
 a99693a <=( a99692a  and  a99685a );
 a99696a <=( A266  and  (not A265) );
 a99699a <=( A268  and  A267 );
 a99700a <=( a99699a  and  a99696a );
 a99703a <=( A299  and  (not A298) );
 a99706a <=( (not A302)  and  A300 );
 a99707a <=( a99706a  and  a99703a );
 a99708a <=( a99707a  and  a99700a );
 a99711a <=( (not A169)  and  (not A170) );
 a99714a <=( (not A199)  and  A168 );
 a99715a <=( a99714a  and  a99711a );
 a99718a <=( (not A201)  and  A200 );
 a99721a <=( A203  and  (not A202) );
 a99722a <=( a99721a  and  a99718a );
 a99723a <=( a99722a  and  a99715a );
 a99726a <=( A266  and  (not A265) );
 a99729a <=( (not A269)  and  A267 );
 a99730a <=( a99729a  and  a99726a );
 a99733a <=( (not A299)  and  A298 );
 a99736a <=( A301  and  A300 );
 a99737a <=( a99736a  and  a99733a );
 a99738a <=( a99737a  and  a99730a );
 a99741a <=( (not A169)  and  (not A170) );
 a99744a <=( (not A199)  and  A168 );
 a99745a <=( a99744a  and  a99741a );
 a99748a <=( (not A201)  and  A200 );
 a99751a <=( A203  and  (not A202) );
 a99752a <=( a99751a  and  a99748a );
 a99753a <=( a99752a  and  a99745a );
 a99756a <=( A266  and  (not A265) );
 a99759a <=( (not A269)  and  A267 );
 a99760a <=( a99759a  and  a99756a );
 a99763a <=( (not A299)  and  A298 );
 a99766a <=( (not A302)  and  A300 );
 a99767a <=( a99766a  and  a99763a );
 a99768a <=( a99767a  and  a99760a );
 a99771a <=( (not A169)  and  (not A170) );
 a99774a <=( (not A199)  and  A168 );
 a99775a <=( a99774a  and  a99771a );
 a99778a <=( (not A201)  and  A200 );
 a99781a <=( A203  and  (not A202) );
 a99782a <=( a99781a  and  a99778a );
 a99783a <=( a99782a  and  a99775a );
 a99786a <=( A266  and  (not A265) );
 a99789a <=( (not A269)  and  A267 );
 a99790a <=( a99789a  and  a99786a );
 a99793a <=( A299  and  (not A298) );
 a99796a <=( A301  and  A300 );
 a99797a <=( a99796a  and  a99793a );
 a99798a <=( a99797a  and  a99790a );
 a99801a <=( (not A169)  and  (not A170) );
 a99804a <=( (not A199)  and  A168 );
 a99805a <=( a99804a  and  a99801a );
 a99808a <=( (not A201)  and  A200 );
 a99811a <=( A203  and  (not A202) );
 a99812a <=( a99811a  and  a99808a );
 a99813a <=( a99812a  and  a99805a );
 a99816a <=( A266  and  (not A265) );
 a99819a <=( (not A269)  and  A267 );
 a99820a <=( a99819a  and  a99816a );
 a99823a <=( A299  and  (not A298) );
 a99826a <=( (not A302)  and  A300 );
 a99827a <=( a99826a  and  a99823a );
 a99828a <=( a99827a  and  a99820a );
 a99831a <=( (not A169)  and  (not A170) );
 a99834a <=( (not A199)  and  A168 );
 a99835a <=( a99834a  and  a99831a );
 a99838a <=( (not A201)  and  A200 );
 a99841a <=( A203  and  (not A202) );
 a99842a <=( a99841a  and  a99838a );
 a99843a <=( a99842a  and  a99835a );
 a99846a <=( (not A266)  and  A265 );
 a99849a <=( A268  and  A267 );
 a99850a <=( a99849a  and  a99846a );
 a99853a <=( (not A299)  and  A298 );
 a99856a <=( A301  and  A300 );
 a99857a <=( a99856a  and  a99853a );
 a99858a <=( a99857a  and  a99850a );
 a99861a <=( (not A169)  and  (not A170) );
 a99864a <=( (not A199)  and  A168 );
 a99865a <=( a99864a  and  a99861a );
 a99868a <=( (not A201)  and  A200 );
 a99871a <=( A203  and  (not A202) );
 a99872a <=( a99871a  and  a99868a );
 a99873a <=( a99872a  and  a99865a );
 a99876a <=( (not A266)  and  A265 );
 a99879a <=( A268  and  A267 );
 a99880a <=( a99879a  and  a99876a );
 a99883a <=( (not A299)  and  A298 );
 a99886a <=( (not A302)  and  A300 );
 a99887a <=( a99886a  and  a99883a );
 a99888a <=( a99887a  and  a99880a );
 a99891a <=( (not A169)  and  (not A170) );
 a99894a <=( (not A199)  and  A168 );
 a99895a <=( a99894a  and  a99891a );
 a99898a <=( (not A201)  and  A200 );
 a99901a <=( A203  and  (not A202) );
 a99902a <=( a99901a  and  a99898a );
 a99903a <=( a99902a  and  a99895a );
 a99906a <=( (not A266)  and  A265 );
 a99909a <=( A268  and  A267 );
 a99910a <=( a99909a  and  a99906a );
 a99913a <=( A299  and  (not A298) );
 a99916a <=( A301  and  A300 );
 a99917a <=( a99916a  and  a99913a );
 a99918a <=( a99917a  and  a99910a );
 a99921a <=( (not A169)  and  (not A170) );
 a99924a <=( (not A199)  and  A168 );
 a99925a <=( a99924a  and  a99921a );
 a99928a <=( (not A201)  and  A200 );
 a99931a <=( A203  and  (not A202) );
 a99932a <=( a99931a  and  a99928a );
 a99933a <=( a99932a  and  a99925a );
 a99936a <=( (not A266)  and  A265 );
 a99939a <=( A268  and  A267 );
 a99940a <=( a99939a  and  a99936a );
 a99943a <=( A299  and  (not A298) );
 a99946a <=( (not A302)  and  A300 );
 a99947a <=( a99946a  and  a99943a );
 a99948a <=( a99947a  and  a99940a );
 a99951a <=( (not A169)  and  (not A170) );
 a99954a <=( (not A199)  and  A168 );
 a99955a <=( a99954a  and  a99951a );
 a99958a <=( (not A201)  and  A200 );
 a99961a <=( A203  and  (not A202) );
 a99962a <=( a99961a  and  a99958a );
 a99963a <=( a99962a  and  a99955a );
 a99966a <=( (not A266)  and  A265 );
 a99969a <=( (not A269)  and  A267 );
 a99970a <=( a99969a  and  a99966a );
 a99973a <=( (not A299)  and  A298 );
 a99976a <=( A301  and  A300 );
 a99977a <=( a99976a  and  a99973a );
 a99978a <=( a99977a  and  a99970a );
 a99981a <=( (not A169)  and  (not A170) );
 a99984a <=( (not A199)  and  A168 );
 a99985a <=( a99984a  and  a99981a );
 a99988a <=( (not A201)  and  A200 );
 a99991a <=( A203  and  (not A202) );
 a99992a <=( a99991a  and  a99988a );
 a99993a <=( a99992a  and  a99985a );
 a99996a <=( (not A266)  and  A265 );
 a99999a <=( (not A269)  and  A267 );
 a100000a <=( a99999a  and  a99996a );
 a100003a <=( (not A299)  and  A298 );
 a100006a <=( (not A302)  and  A300 );
 a100007a <=( a100006a  and  a100003a );
 a100008a <=( a100007a  and  a100000a );
 a100011a <=( (not A169)  and  (not A170) );
 a100014a <=( (not A199)  and  A168 );
 a100015a <=( a100014a  and  a100011a );
 a100018a <=( (not A201)  and  A200 );
 a100021a <=( A203  and  (not A202) );
 a100022a <=( a100021a  and  a100018a );
 a100023a <=( a100022a  and  a100015a );
 a100026a <=( (not A266)  and  A265 );
 a100029a <=( (not A269)  and  A267 );
 a100030a <=( a100029a  and  a100026a );
 a100033a <=( A299  and  (not A298) );
 a100036a <=( A301  and  A300 );
 a100037a <=( a100036a  and  a100033a );
 a100038a <=( a100037a  and  a100030a );
 a100041a <=( (not A169)  and  (not A170) );
 a100044a <=( (not A199)  and  A168 );
 a100045a <=( a100044a  and  a100041a );
 a100048a <=( (not A201)  and  A200 );
 a100051a <=( A203  and  (not A202) );
 a100052a <=( a100051a  and  a100048a );
 a100053a <=( a100052a  and  a100045a );
 a100056a <=( (not A266)  and  A265 );
 a100059a <=( (not A269)  and  A267 );
 a100060a <=( a100059a  and  a100056a );
 a100063a <=( A299  and  (not A298) );
 a100066a <=( (not A302)  and  A300 );
 a100067a <=( a100066a  and  a100063a );
 a100068a <=( a100067a  and  a100060a );
 a100071a <=( (not A169)  and  (not A170) );
 a100074a <=( A199  and  A168 );
 a100075a <=( a100074a  and  a100071a );
 a100078a <=( A201  and  (not A200) );
 a100081a <=( (not A265)  and  A202 );
 a100082a <=( a100081a  and  a100078a );
 a100083a <=( a100082a  and  a100075a );
 a100086a <=( A267  and  A266 );
 a100089a <=( A298  and  A268 );
 a100090a <=( a100089a  and  a100086a );
 a100093a <=( (not A300)  and  (not A299) );
 a100096a <=( A302  and  (not A301) );
 a100097a <=( a100096a  and  a100093a );
 a100098a <=( a100097a  and  a100090a );
 a100101a <=( (not A169)  and  (not A170) );
 a100104a <=( A199  and  A168 );
 a100105a <=( a100104a  and  a100101a );
 a100108a <=( A201  and  (not A200) );
 a100111a <=( (not A265)  and  A202 );
 a100112a <=( a100111a  and  a100108a );
 a100113a <=( a100112a  and  a100105a );
 a100116a <=( A267  and  A266 );
 a100119a <=( (not A298)  and  A268 );
 a100120a <=( a100119a  and  a100116a );
 a100123a <=( (not A300)  and  A299 );
 a100126a <=( A302  and  (not A301) );
 a100127a <=( a100126a  and  a100123a );
 a100128a <=( a100127a  and  a100120a );
 a100131a <=( (not A169)  and  (not A170) );
 a100134a <=( A199  and  A168 );
 a100135a <=( a100134a  and  a100131a );
 a100138a <=( A201  and  (not A200) );
 a100141a <=( (not A265)  and  A202 );
 a100142a <=( a100141a  and  a100138a );
 a100143a <=( a100142a  and  a100135a );
 a100146a <=( A267  and  A266 );
 a100149a <=( A298  and  (not A269) );
 a100150a <=( a100149a  and  a100146a );
 a100153a <=( (not A300)  and  (not A299) );
 a100156a <=( A302  and  (not A301) );
 a100157a <=( a100156a  and  a100153a );
 a100158a <=( a100157a  and  a100150a );
 a100161a <=( (not A169)  and  (not A170) );
 a100164a <=( A199  and  A168 );
 a100165a <=( a100164a  and  a100161a );
 a100168a <=( A201  and  (not A200) );
 a100171a <=( (not A265)  and  A202 );
 a100172a <=( a100171a  and  a100168a );
 a100173a <=( a100172a  and  a100165a );
 a100176a <=( A267  and  A266 );
 a100179a <=( (not A298)  and  (not A269) );
 a100180a <=( a100179a  and  a100176a );
 a100183a <=( (not A300)  and  A299 );
 a100186a <=( A302  and  (not A301) );
 a100187a <=( a100186a  and  a100183a );
 a100188a <=( a100187a  and  a100180a );
 a100191a <=( (not A169)  and  (not A170) );
 a100194a <=( A199  and  A168 );
 a100195a <=( a100194a  and  a100191a );
 a100198a <=( A201  and  (not A200) );
 a100201a <=( (not A265)  and  A202 );
 a100202a <=( a100201a  and  a100198a );
 a100203a <=( a100202a  and  a100195a );
 a100206a <=( (not A267)  and  A266 );
 a100209a <=( A269  and  (not A268) );
 a100210a <=( a100209a  and  a100206a );
 a100213a <=( (not A299)  and  A298 );
 a100216a <=( A301  and  A300 );
 a100217a <=( a100216a  and  a100213a );
 a100218a <=( a100217a  and  a100210a );
 a100221a <=( (not A169)  and  (not A170) );
 a100224a <=( A199  and  A168 );
 a100225a <=( a100224a  and  a100221a );
 a100228a <=( A201  and  (not A200) );
 a100231a <=( (not A265)  and  A202 );
 a100232a <=( a100231a  and  a100228a );
 a100233a <=( a100232a  and  a100225a );
 a100236a <=( (not A267)  and  A266 );
 a100239a <=( A269  and  (not A268) );
 a100240a <=( a100239a  and  a100236a );
 a100243a <=( (not A299)  and  A298 );
 a100246a <=( (not A302)  and  A300 );
 a100247a <=( a100246a  and  a100243a );
 a100248a <=( a100247a  and  a100240a );
 a100251a <=( (not A169)  and  (not A170) );
 a100254a <=( A199  and  A168 );
 a100255a <=( a100254a  and  a100251a );
 a100258a <=( A201  and  (not A200) );
 a100261a <=( (not A265)  and  A202 );
 a100262a <=( a100261a  and  a100258a );
 a100263a <=( a100262a  and  a100255a );
 a100266a <=( (not A267)  and  A266 );
 a100269a <=( A269  and  (not A268) );
 a100270a <=( a100269a  and  a100266a );
 a100273a <=( A299  and  (not A298) );
 a100276a <=( A301  and  A300 );
 a100277a <=( a100276a  and  a100273a );
 a100278a <=( a100277a  and  a100270a );
 a100281a <=( (not A169)  and  (not A170) );
 a100284a <=( A199  and  A168 );
 a100285a <=( a100284a  and  a100281a );
 a100288a <=( A201  and  (not A200) );
 a100291a <=( (not A265)  and  A202 );
 a100292a <=( a100291a  and  a100288a );
 a100293a <=( a100292a  and  a100285a );
 a100296a <=( (not A267)  and  A266 );
 a100299a <=( A269  and  (not A268) );
 a100300a <=( a100299a  and  a100296a );
 a100303a <=( A299  and  (not A298) );
 a100306a <=( (not A302)  and  A300 );
 a100307a <=( a100306a  and  a100303a );
 a100308a <=( a100307a  and  a100300a );
 a100311a <=( (not A169)  and  (not A170) );
 a100314a <=( A199  and  A168 );
 a100315a <=( a100314a  and  a100311a );
 a100318a <=( A201  and  (not A200) );
 a100321a <=( A265  and  A202 );
 a100322a <=( a100321a  and  a100318a );
 a100323a <=( a100322a  and  a100315a );
 a100326a <=( A267  and  (not A266) );
 a100329a <=( A298  and  A268 );
 a100330a <=( a100329a  and  a100326a );
 a100333a <=( (not A300)  and  (not A299) );
 a100336a <=( A302  and  (not A301) );
 a100337a <=( a100336a  and  a100333a );
 a100338a <=( a100337a  and  a100330a );
 a100341a <=( (not A169)  and  (not A170) );
 a100344a <=( A199  and  A168 );
 a100345a <=( a100344a  and  a100341a );
 a100348a <=( A201  and  (not A200) );
 a100351a <=( A265  and  A202 );
 a100352a <=( a100351a  and  a100348a );
 a100353a <=( a100352a  and  a100345a );
 a100356a <=( A267  and  (not A266) );
 a100359a <=( (not A298)  and  A268 );
 a100360a <=( a100359a  and  a100356a );
 a100363a <=( (not A300)  and  A299 );
 a100366a <=( A302  and  (not A301) );
 a100367a <=( a100366a  and  a100363a );
 a100368a <=( a100367a  and  a100360a );
 a100371a <=( (not A169)  and  (not A170) );
 a100374a <=( A199  and  A168 );
 a100375a <=( a100374a  and  a100371a );
 a100378a <=( A201  and  (not A200) );
 a100381a <=( A265  and  A202 );
 a100382a <=( a100381a  and  a100378a );
 a100383a <=( a100382a  and  a100375a );
 a100386a <=( A267  and  (not A266) );
 a100389a <=( A298  and  (not A269) );
 a100390a <=( a100389a  and  a100386a );
 a100393a <=( (not A300)  and  (not A299) );
 a100396a <=( A302  and  (not A301) );
 a100397a <=( a100396a  and  a100393a );
 a100398a <=( a100397a  and  a100390a );
 a100401a <=( (not A169)  and  (not A170) );
 a100404a <=( A199  and  A168 );
 a100405a <=( a100404a  and  a100401a );
 a100408a <=( A201  and  (not A200) );
 a100411a <=( A265  and  A202 );
 a100412a <=( a100411a  and  a100408a );
 a100413a <=( a100412a  and  a100405a );
 a100416a <=( A267  and  (not A266) );
 a100419a <=( (not A298)  and  (not A269) );
 a100420a <=( a100419a  and  a100416a );
 a100423a <=( (not A300)  and  A299 );
 a100426a <=( A302  and  (not A301) );
 a100427a <=( a100426a  and  a100423a );
 a100428a <=( a100427a  and  a100420a );
 a100431a <=( (not A169)  and  (not A170) );
 a100434a <=( A199  and  A168 );
 a100435a <=( a100434a  and  a100431a );
 a100438a <=( A201  and  (not A200) );
 a100441a <=( A265  and  A202 );
 a100442a <=( a100441a  and  a100438a );
 a100443a <=( a100442a  and  a100435a );
 a100446a <=( (not A267)  and  (not A266) );
 a100449a <=( A269  and  (not A268) );
 a100450a <=( a100449a  and  a100446a );
 a100453a <=( (not A299)  and  A298 );
 a100456a <=( A301  and  A300 );
 a100457a <=( a100456a  and  a100453a );
 a100458a <=( a100457a  and  a100450a );
 a100461a <=( (not A169)  and  (not A170) );
 a100464a <=( A199  and  A168 );
 a100465a <=( a100464a  and  a100461a );
 a100468a <=( A201  and  (not A200) );
 a100471a <=( A265  and  A202 );
 a100472a <=( a100471a  and  a100468a );
 a100473a <=( a100472a  and  a100465a );
 a100476a <=( (not A267)  and  (not A266) );
 a100479a <=( A269  and  (not A268) );
 a100480a <=( a100479a  and  a100476a );
 a100483a <=( (not A299)  and  A298 );
 a100486a <=( (not A302)  and  A300 );
 a100487a <=( a100486a  and  a100483a );
 a100488a <=( a100487a  and  a100480a );
 a100491a <=( (not A169)  and  (not A170) );
 a100494a <=( A199  and  A168 );
 a100495a <=( a100494a  and  a100491a );
 a100498a <=( A201  and  (not A200) );
 a100501a <=( A265  and  A202 );
 a100502a <=( a100501a  and  a100498a );
 a100503a <=( a100502a  and  a100495a );
 a100506a <=( (not A267)  and  (not A266) );
 a100509a <=( A269  and  (not A268) );
 a100510a <=( a100509a  and  a100506a );
 a100513a <=( A299  and  (not A298) );
 a100516a <=( A301  and  A300 );
 a100517a <=( a100516a  and  a100513a );
 a100518a <=( a100517a  and  a100510a );
 a100521a <=( (not A169)  and  (not A170) );
 a100524a <=( A199  and  A168 );
 a100525a <=( a100524a  and  a100521a );
 a100528a <=( A201  and  (not A200) );
 a100531a <=( A265  and  A202 );
 a100532a <=( a100531a  and  a100528a );
 a100533a <=( a100532a  and  a100525a );
 a100536a <=( (not A267)  and  (not A266) );
 a100539a <=( A269  and  (not A268) );
 a100540a <=( a100539a  and  a100536a );
 a100543a <=( A299  and  (not A298) );
 a100546a <=( (not A302)  and  A300 );
 a100547a <=( a100546a  and  a100543a );
 a100548a <=( a100547a  and  a100540a );
 a100551a <=( (not A169)  and  (not A170) );
 a100554a <=( A199  and  A168 );
 a100555a <=( a100554a  and  a100551a );
 a100558a <=( A201  and  (not A200) );
 a100561a <=( (not A265)  and  (not A203) );
 a100562a <=( a100561a  and  a100558a );
 a100563a <=( a100562a  and  a100555a );
 a100566a <=( A267  and  A266 );
 a100569a <=( A298  and  A268 );
 a100570a <=( a100569a  and  a100566a );
 a100573a <=( (not A300)  and  (not A299) );
 a100576a <=( A302  and  (not A301) );
 a100577a <=( a100576a  and  a100573a );
 a100578a <=( a100577a  and  a100570a );
 a100581a <=( (not A169)  and  (not A170) );
 a100584a <=( A199  and  A168 );
 a100585a <=( a100584a  and  a100581a );
 a100588a <=( A201  and  (not A200) );
 a100591a <=( (not A265)  and  (not A203) );
 a100592a <=( a100591a  and  a100588a );
 a100593a <=( a100592a  and  a100585a );
 a100596a <=( A267  and  A266 );
 a100599a <=( (not A298)  and  A268 );
 a100600a <=( a100599a  and  a100596a );
 a100603a <=( (not A300)  and  A299 );
 a100606a <=( A302  and  (not A301) );
 a100607a <=( a100606a  and  a100603a );
 a100608a <=( a100607a  and  a100600a );
 a100611a <=( (not A169)  and  (not A170) );
 a100614a <=( A199  and  A168 );
 a100615a <=( a100614a  and  a100611a );
 a100618a <=( A201  and  (not A200) );
 a100621a <=( (not A265)  and  (not A203) );
 a100622a <=( a100621a  and  a100618a );
 a100623a <=( a100622a  and  a100615a );
 a100626a <=( A267  and  A266 );
 a100629a <=( A298  and  (not A269) );
 a100630a <=( a100629a  and  a100626a );
 a100633a <=( (not A300)  and  (not A299) );
 a100636a <=( A302  and  (not A301) );
 a100637a <=( a100636a  and  a100633a );
 a100638a <=( a100637a  and  a100630a );
 a100641a <=( (not A169)  and  (not A170) );
 a100644a <=( A199  and  A168 );
 a100645a <=( a100644a  and  a100641a );
 a100648a <=( A201  and  (not A200) );
 a100651a <=( (not A265)  and  (not A203) );
 a100652a <=( a100651a  and  a100648a );
 a100653a <=( a100652a  and  a100645a );
 a100656a <=( A267  and  A266 );
 a100659a <=( (not A298)  and  (not A269) );
 a100660a <=( a100659a  and  a100656a );
 a100663a <=( (not A300)  and  A299 );
 a100666a <=( A302  and  (not A301) );
 a100667a <=( a100666a  and  a100663a );
 a100668a <=( a100667a  and  a100660a );
 a100671a <=( (not A169)  and  (not A170) );
 a100674a <=( A199  and  A168 );
 a100675a <=( a100674a  and  a100671a );
 a100678a <=( A201  and  (not A200) );
 a100681a <=( (not A265)  and  (not A203) );
 a100682a <=( a100681a  and  a100678a );
 a100683a <=( a100682a  and  a100675a );
 a100686a <=( (not A267)  and  A266 );
 a100689a <=( A269  and  (not A268) );
 a100690a <=( a100689a  and  a100686a );
 a100693a <=( (not A299)  and  A298 );
 a100696a <=( A301  and  A300 );
 a100697a <=( a100696a  and  a100693a );
 a100698a <=( a100697a  and  a100690a );
 a100701a <=( (not A169)  and  (not A170) );
 a100704a <=( A199  and  A168 );
 a100705a <=( a100704a  and  a100701a );
 a100708a <=( A201  and  (not A200) );
 a100711a <=( (not A265)  and  (not A203) );
 a100712a <=( a100711a  and  a100708a );
 a100713a <=( a100712a  and  a100705a );
 a100716a <=( (not A267)  and  A266 );
 a100719a <=( A269  and  (not A268) );
 a100720a <=( a100719a  and  a100716a );
 a100723a <=( (not A299)  and  A298 );
 a100726a <=( (not A302)  and  A300 );
 a100727a <=( a100726a  and  a100723a );
 a100728a <=( a100727a  and  a100720a );
 a100731a <=( (not A169)  and  (not A170) );
 a100734a <=( A199  and  A168 );
 a100735a <=( a100734a  and  a100731a );
 a100738a <=( A201  and  (not A200) );
 a100741a <=( (not A265)  and  (not A203) );
 a100742a <=( a100741a  and  a100738a );
 a100743a <=( a100742a  and  a100735a );
 a100746a <=( (not A267)  and  A266 );
 a100749a <=( A269  and  (not A268) );
 a100750a <=( a100749a  and  a100746a );
 a100753a <=( A299  and  (not A298) );
 a100756a <=( A301  and  A300 );
 a100757a <=( a100756a  and  a100753a );
 a100758a <=( a100757a  and  a100750a );
 a100761a <=( (not A169)  and  (not A170) );
 a100764a <=( A199  and  A168 );
 a100765a <=( a100764a  and  a100761a );
 a100768a <=( A201  and  (not A200) );
 a100771a <=( (not A265)  and  (not A203) );
 a100772a <=( a100771a  and  a100768a );
 a100773a <=( a100772a  and  a100765a );
 a100776a <=( (not A267)  and  A266 );
 a100779a <=( A269  and  (not A268) );
 a100780a <=( a100779a  and  a100776a );
 a100783a <=( A299  and  (not A298) );
 a100786a <=( (not A302)  and  A300 );
 a100787a <=( a100786a  and  a100783a );
 a100788a <=( a100787a  and  a100780a );
 a100791a <=( (not A169)  and  (not A170) );
 a100794a <=( A199  and  A168 );
 a100795a <=( a100794a  and  a100791a );
 a100798a <=( A201  and  (not A200) );
 a100801a <=( A265  and  (not A203) );
 a100802a <=( a100801a  and  a100798a );
 a100803a <=( a100802a  and  a100795a );
 a100806a <=( A267  and  (not A266) );
 a100809a <=( A298  and  A268 );
 a100810a <=( a100809a  and  a100806a );
 a100813a <=( (not A300)  and  (not A299) );
 a100816a <=( A302  and  (not A301) );
 a100817a <=( a100816a  and  a100813a );
 a100818a <=( a100817a  and  a100810a );
 a100821a <=( (not A169)  and  (not A170) );
 a100824a <=( A199  and  A168 );
 a100825a <=( a100824a  and  a100821a );
 a100828a <=( A201  and  (not A200) );
 a100831a <=( A265  and  (not A203) );
 a100832a <=( a100831a  and  a100828a );
 a100833a <=( a100832a  and  a100825a );
 a100836a <=( A267  and  (not A266) );
 a100839a <=( (not A298)  and  A268 );
 a100840a <=( a100839a  and  a100836a );
 a100843a <=( (not A300)  and  A299 );
 a100846a <=( A302  and  (not A301) );
 a100847a <=( a100846a  and  a100843a );
 a100848a <=( a100847a  and  a100840a );
 a100851a <=( (not A169)  and  (not A170) );
 a100854a <=( A199  and  A168 );
 a100855a <=( a100854a  and  a100851a );
 a100858a <=( A201  and  (not A200) );
 a100861a <=( A265  and  (not A203) );
 a100862a <=( a100861a  and  a100858a );
 a100863a <=( a100862a  and  a100855a );
 a100866a <=( A267  and  (not A266) );
 a100869a <=( A298  and  (not A269) );
 a100870a <=( a100869a  and  a100866a );
 a100873a <=( (not A300)  and  (not A299) );
 a100876a <=( A302  and  (not A301) );
 a100877a <=( a100876a  and  a100873a );
 a100878a <=( a100877a  and  a100870a );
 a100881a <=( (not A169)  and  (not A170) );
 a100884a <=( A199  and  A168 );
 a100885a <=( a100884a  and  a100881a );
 a100888a <=( A201  and  (not A200) );
 a100891a <=( A265  and  (not A203) );
 a100892a <=( a100891a  and  a100888a );
 a100893a <=( a100892a  and  a100885a );
 a100896a <=( A267  and  (not A266) );
 a100899a <=( (not A298)  and  (not A269) );
 a100900a <=( a100899a  and  a100896a );
 a100903a <=( (not A300)  and  A299 );
 a100906a <=( A302  and  (not A301) );
 a100907a <=( a100906a  and  a100903a );
 a100908a <=( a100907a  and  a100900a );
 a100911a <=( (not A169)  and  (not A170) );
 a100914a <=( A199  and  A168 );
 a100915a <=( a100914a  and  a100911a );
 a100918a <=( A201  and  (not A200) );
 a100921a <=( A265  and  (not A203) );
 a100922a <=( a100921a  and  a100918a );
 a100923a <=( a100922a  and  a100915a );
 a100926a <=( (not A267)  and  (not A266) );
 a100929a <=( A269  and  (not A268) );
 a100930a <=( a100929a  and  a100926a );
 a100933a <=( (not A299)  and  A298 );
 a100936a <=( A301  and  A300 );
 a100937a <=( a100936a  and  a100933a );
 a100938a <=( a100937a  and  a100930a );
 a100941a <=( (not A169)  and  (not A170) );
 a100944a <=( A199  and  A168 );
 a100945a <=( a100944a  and  a100941a );
 a100948a <=( A201  and  (not A200) );
 a100951a <=( A265  and  (not A203) );
 a100952a <=( a100951a  and  a100948a );
 a100953a <=( a100952a  and  a100945a );
 a100956a <=( (not A267)  and  (not A266) );
 a100959a <=( A269  and  (not A268) );
 a100960a <=( a100959a  and  a100956a );
 a100963a <=( (not A299)  and  A298 );
 a100966a <=( (not A302)  and  A300 );
 a100967a <=( a100966a  and  a100963a );
 a100968a <=( a100967a  and  a100960a );
 a100971a <=( (not A169)  and  (not A170) );
 a100974a <=( A199  and  A168 );
 a100975a <=( a100974a  and  a100971a );
 a100978a <=( A201  and  (not A200) );
 a100981a <=( A265  and  (not A203) );
 a100982a <=( a100981a  and  a100978a );
 a100983a <=( a100982a  and  a100975a );
 a100986a <=( (not A267)  and  (not A266) );
 a100989a <=( A269  and  (not A268) );
 a100990a <=( a100989a  and  a100986a );
 a100993a <=( A299  and  (not A298) );
 a100996a <=( A301  and  A300 );
 a100997a <=( a100996a  and  a100993a );
 a100998a <=( a100997a  and  a100990a );
 a101001a <=( (not A169)  and  (not A170) );
 a101004a <=( A199  and  A168 );
 a101005a <=( a101004a  and  a101001a );
 a101008a <=( A201  and  (not A200) );
 a101011a <=( A265  and  (not A203) );
 a101012a <=( a101011a  and  a101008a );
 a101013a <=( a101012a  and  a101005a );
 a101016a <=( (not A267)  and  (not A266) );
 a101019a <=( A269  and  (not A268) );
 a101020a <=( a101019a  and  a101016a );
 a101023a <=( A299  and  (not A298) );
 a101026a <=( (not A302)  and  A300 );
 a101027a <=( a101026a  and  a101023a );
 a101028a <=( a101027a  and  a101020a );
 a101031a <=( (not A169)  and  (not A170) );
 a101034a <=( A199  and  A168 );
 a101035a <=( a101034a  and  a101031a );
 a101038a <=( (not A201)  and  (not A200) );
 a101041a <=( A203  and  (not A202) );
 a101042a <=( a101041a  and  a101038a );
 a101043a <=( a101042a  and  a101035a );
 a101046a <=( A266  and  (not A265) );
 a101049a <=( A268  and  A267 );
 a101050a <=( a101049a  and  a101046a );
 a101053a <=( (not A299)  and  A298 );
 a101056a <=( A301  and  A300 );
 a101057a <=( a101056a  and  a101053a );
 a101058a <=( a101057a  and  a101050a );
 a101061a <=( (not A169)  and  (not A170) );
 a101064a <=( A199  and  A168 );
 a101065a <=( a101064a  and  a101061a );
 a101068a <=( (not A201)  and  (not A200) );
 a101071a <=( A203  and  (not A202) );
 a101072a <=( a101071a  and  a101068a );
 a101073a <=( a101072a  and  a101065a );
 a101076a <=( A266  and  (not A265) );
 a101079a <=( A268  and  A267 );
 a101080a <=( a101079a  and  a101076a );
 a101083a <=( (not A299)  and  A298 );
 a101086a <=( (not A302)  and  A300 );
 a101087a <=( a101086a  and  a101083a );
 a101088a <=( a101087a  and  a101080a );
 a101091a <=( (not A169)  and  (not A170) );
 a101094a <=( A199  and  A168 );
 a101095a <=( a101094a  and  a101091a );
 a101098a <=( (not A201)  and  (not A200) );
 a101101a <=( A203  and  (not A202) );
 a101102a <=( a101101a  and  a101098a );
 a101103a <=( a101102a  and  a101095a );
 a101106a <=( A266  and  (not A265) );
 a101109a <=( A268  and  A267 );
 a101110a <=( a101109a  and  a101106a );
 a101113a <=( A299  and  (not A298) );
 a101116a <=( A301  and  A300 );
 a101117a <=( a101116a  and  a101113a );
 a101118a <=( a101117a  and  a101110a );
 a101121a <=( (not A169)  and  (not A170) );
 a101124a <=( A199  and  A168 );
 a101125a <=( a101124a  and  a101121a );
 a101128a <=( (not A201)  and  (not A200) );
 a101131a <=( A203  and  (not A202) );
 a101132a <=( a101131a  and  a101128a );
 a101133a <=( a101132a  and  a101125a );
 a101136a <=( A266  and  (not A265) );
 a101139a <=( A268  and  A267 );
 a101140a <=( a101139a  and  a101136a );
 a101143a <=( A299  and  (not A298) );
 a101146a <=( (not A302)  and  A300 );
 a101147a <=( a101146a  and  a101143a );
 a101148a <=( a101147a  and  a101140a );
 a101151a <=( (not A169)  and  (not A170) );
 a101154a <=( A199  and  A168 );
 a101155a <=( a101154a  and  a101151a );
 a101158a <=( (not A201)  and  (not A200) );
 a101161a <=( A203  and  (not A202) );
 a101162a <=( a101161a  and  a101158a );
 a101163a <=( a101162a  and  a101155a );
 a101166a <=( A266  and  (not A265) );
 a101169a <=( (not A269)  and  A267 );
 a101170a <=( a101169a  and  a101166a );
 a101173a <=( (not A299)  and  A298 );
 a101176a <=( A301  and  A300 );
 a101177a <=( a101176a  and  a101173a );
 a101178a <=( a101177a  and  a101170a );
 a101181a <=( (not A169)  and  (not A170) );
 a101184a <=( A199  and  A168 );
 a101185a <=( a101184a  and  a101181a );
 a101188a <=( (not A201)  and  (not A200) );
 a101191a <=( A203  and  (not A202) );
 a101192a <=( a101191a  and  a101188a );
 a101193a <=( a101192a  and  a101185a );
 a101196a <=( A266  and  (not A265) );
 a101199a <=( (not A269)  and  A267 );
 a101200a <=( a101199a  and  a101196a );
 a101203a <=( (not A299)  and  A298 );
 a101206a <=( (not A302)  and  A300 );
 a101207a <=( a101206a  and  a101203a );
 a101208a <=( a101207a  and  a101200a );
 a101211a <=( (not A169)  and  (not A170) );
 a101214a <=( A199  and  A168 );
 a101215a <=( a101214a  and  a101211a );
 a101218a <=( (not A201)  and  (not A200) );
 a101221a <=( A203  and  (not A202) );
 a101222a <=( a101221a  and  a101218a );
 a101223a <=( a101222a  and  a101215a );
 a101226a <=( A266  and  (not A265) );
 a101229a <=( (not A269)  and  A267 );
 a101230a <=( a101229a  and  a101226a );
 a101233a <=( A299  and  (not A298) );
 a101236a <=( A301  and  A300 );
 a101237a <=( a101236a  and  a101233a );
 a101238a <=( a101237a  and  a101230a );
 a101241a <=( (not A169)  and  (not A170) );
 a101244a <=( A199  and  A168 );
 a101245a <=( a101244a  and  a101241a );
 a101248a <=( (not A201)  and  (not A200) );
 a101251a <=( A203  and  (not A202) );
 a101252a <=( a101251a  and  a101248a );
 a101253a <=( a101252a  and  a101245a );
 a101256a <=( A266  and  (not A265) );
 a101259a <=( (not A269)  and  A267 );
 a101260a <=( a101259a  and  a101256a );
 a101263a <=( A299  and  (not A298) );
 a101266a <=( (not A302)  and  A300 );
 a101267a <=( a101266a  and  a101263a );
 a101268a <=( a101267a  and  a101260a );
 a101271a <=( (not A169)  and  (not A170) );
 a101274a <=( A199  and  A168 );
 a101275a <=( a101274a  and  a101271a );
 a101278a <=( (not A201)  and  (not A200) );
 a101281a <=( A203  and  (not A202) );
 a101282a <=( a101281a  and  a101278a );
 a101283a <=( a101282a  and  a101275a );
 a101286a <=( (not A266)  and  A265 );
 a101289a <=( A268  and  A267 );
 a101290a <=( a101289a  and  a101286a );
 a101293a <=( (not A299)  and  A298 );
 a101296a <=( A301  and  A300 );
 a101297a <=( a101296a  and  a101293a );
 a101298a <=( a101297a  and  a101290a );
 a101301a <=( (not A169)  and  (not A170) );
 a101304a <=( A199  and  A168 );
 a101305a <=( a101304a  and  a101301a );
 a101308a <=( (not A201)  and  (not A200) );
 a101311a <=( A203  and  (not A202) );
 a101312a <=( a101311a  and  a101308a );
 a101313a <=( a101312a  and  a101305a );
 a101316a <=( (not A266)  and  A265 );
 a101319a <=( A268  and  A267 );
 a101320a <=( a101319a  and  a101316a );
 a101323a <=( (not A299)  and  A298 );
 a101326a <=( (not A302)  and  A300 );
 a101327a <=( a101326a  and  a101323a );
 a101328a <=( a101327a  and  a101320a );
 a101331a <=( (not A169)  and  (not A170) );
 a101334a <=( A199  and  A168 );
 a101335a <=( a101334a  and  a101331a );
 a101338a <=( (not A201)  and  (not A200) );
 a101341a <=( A203  and  (not A202) );
 a101342a <=( a101341a  and  a101338a );
 a101343a <=( a101342a  and  a101335a );
 a101346a <=( (not A266)  and  A265 );
 a101349a <=( A268  and  A267 );
 a101350a <=( a101349a  and  a101346a );
 a101353a <=( A299  and  (not A298) );
 a101356a <=( A301  and  A300 );
 a101357a <=( a101356a  and  a101353a );
 a101358a <=( a101357a  and  a101350a );
 a101361a <=( (not A169)  and  (not A170) );
 a101364a <=( A199  and  A168 );
 a101365a <=( a101364a  and  a101361a );
 a101368a <=( (not A201)  and  (not A200) );
 a101371a <=( A203  and  (not A202) );
 a101372a <=( a101371a  and  a101368a );
 a101373a <=( a101372a  and  a101365a );
 a101376a <=( (not A266)  and  A265 );
 a101379a <=( A268  and  A267 );
 a101380a <=( a101379a  and  a101376a );
 a101383a <=( A299  and  (not A298) );
 a101386a <=( (not A302)  and  A300 );
 a101387a <=( a101386a  and  a101383a );
 a101388a <=( a101387a  and  a101380a );
 a101391a <=( (not A169)  and  (not A170) );
 a101394a <=( A199  and  A168 );
 a101395a <=( a101394a  and  a101391a );
 a101398a <=( (not A201)  and  (not A200) );
 a101401a <=( A203  and  (not A202) );
 a101402a <=( a101401a  and  a101398a );
 a101403a <=( a101402a  and  a101395a );
 a101406a <=( (not A266)  and  A265 );
 a101409a <=( (not A269)  and  A267 );
 a101410a <=( a101409a  and  a101406a );
 a101413a <=( (not A299)  and  A298 );
 a101416a <=( A301  and  A300 );
 a101417a <=( a101416a  and  a101413a );
 a101418a <=( a101417a  and  a101410a );
 a101421a <=( (not A169)  and  (not A170) );
 a101424a <=( A199  and  A168 );
 a101425a <=( a101424a  and  a101421a );
 a101428a <=( (not A201)  and  (not A200) );
 a101431a <=( A203  and  (not A202) );
 a101432a <=( a101431a  and  a101428a );
 a101433a <=( a101432a  and  a101425a );
 a101436a <=( (not A266)  and  A265 );
 a101439a <=( (not A269)  and  A267 );
 a101440a <=( a101439a  and  a101436a );
 a101443a <=( (not A299)  and  A298 );
 a101446a <=( (not A302)  and  A300 );
 a101447a <=( a101446a  and  a101443a );
 a101448a <=( a101447a  and  a101440a );
 a101451a <=( (not A169)  and  (not A170) );
 a101454a <=( A199  and  A168 );
 a101455a <=( a101454a  and  a101451a );
 a101458a <=( (not A201)  and  (not A200) );
 a101461a <=( A203  and  (not A202) );
 a101462a <=( a101461a  and  a101458a );
 a101463a <=( a101462a  and  a101455a );
 a101466a <=( (not A266)  and  A265 );
 a101469a <=( (not A269)  and  A267 );
 a101470a <=( a101469a  and  a101466a );
 a101473a <=( A299  and  (not A298) );
 a101476a <=( A301  and  A300 );
 a101477a <=( a101476a  and  a101473a );
 a101478a <=( a101477a  and  a101470a );
 a101481a <=( (not A169)  and  (not A170) );
 a101484a <=( A199  and  A168 );
 a101485a <=( a101484a  and  a101481a );
 a101488a <=( (not A201)  and  (not A200) );
 a101491a <=( A203  and  (not A202) );
 a101492a <=( a101491a  and  a101488a );
 a101493a <=( a101492a  and  a101485a );
 a101496a <=( (not A266)  and  A265 );
 a101499a <=( (not A269)  and  A267 );
 a101500a <=( a101499a  and  a101496a );
 a101503a <=( A299  and  (not A298) );
 a101506a <=( (not A302)  and  A300 );
 a101507a <=( a101506a  and  a101503a );
 a101508a <=( a101507a  and  a101500a );
 a101511a <=( (not A169)  and  (not A170) );
 a101514a <=( A167  and  (not A168) );
 a101515a <=( a101514a  and  a101511a );
 a101518a <=( A201  and  (not A166) );
 a101521a <=( A203  and  (not A202) );
 a101522a <=( a101521a  and  a101518a );
 a101523a <=( a101522a  and  a101515a );
 a101526a <=( (not A268)  and  A267 );
 a101529a <=( A298  and  A269 );
 a101530a <=( a101529a  and  a101526a );
 a101533a <=( (not A300)  and  (not A299) );
 a101536a <=( A302  and  (not A301) );
 a101537a <=( a101536a  and  a101533a );
 a101538a <=( a101537a  and  a101530a );
 a101541a <=( (not A169)  and  (not A170) );
 a101544a <=( A167  and  (not A168) );
 a101545a <=( a101544a  and  a101541a );
 a101548a <=( A201  and  (not A166) );
 a101551a <=( A203  and  (not A202) );
 a101552a <=( a101551a  and  a101548a );
 a101553a <=( a101552a  and  a101545a );
 a101556a <=( (not A268)  and  A267 );
 a101559a <=( (not A298)  and  A269 );
 a101560a <=( a101559a  and  a101556a );
 a101563a <=( (not A300)  and  A299 );
 a101566a <=( A302  and  (not A301) );
 a101567a <=( a101566a  and  a101563a );
 a101568a <=( a101567a  and  a101560a );
 a101571a <=( (not A169)  and  (not A170) );
 a101574a <=( A167  and  (not A168) );
 a101575a <=( a101574a  and  a101571a );
 a101578a <=( A201  and  (not A166) );
 a101581a <=( A203  and  (not A202) );
 a101582a <=( a101581a  and  a101578a );
 a101583a <=( a101582a  and  a101575a );
 a101586a <=( A266  and  (not A265) );
 a101589a <=( (not A268)  and  (not A267) );
 a101590a <=( a101589a  and  a101586a );
 a101593a <=( A300  and  A269 );
 a101596a <=( A302  and  (not A301) );
 a101597a <=( a101596a  and  a101593a );
 a101598a <=( a101597a  and  a101590a );
 a101601a <=( (not A169)  and  (not A170) );
 a101604a <=( A167  and  (not A168) );
 a101605a <=( a101604a  and  a101601a );
 a101608a <=( A201  and  (not A166) );
 a101611a <=( A203  and  (not A202) );
 a101612a <=( a101611a  and  a101608a );
 a101613a <=( a101612a  and  a101605a );
 a101616a <=( (not A266)  and  A265 );
 a101619a <=( (not A268)  and  (not A267) );
 a101620a <=( a101619a  and  a101616a );
 a101623a <=( A300  and  A269 );
 a101626a <=( A302  and  (not A301) );
 a101627a <=( a101626a  and  a101623a );
 a101628a <=( a101627a  and  a101620a );
 a101631a <=( (not A169)  and  (not A170) );
 a101634a <=( (not A167)  and  (not A168) );
 a101635a <=( a101634a  and  a101631a );
 a101638a <=( A201  and  A166 );
 a101641a <=( A203  and  (not A202) );
 a101642a <=( a101641a  and  a101638a );
 a101643a <=( a101642a  and  a101635a );
 a101646a <=( (not A268)  and  A267 );
 a101649a <=( A298  and  A269 );
 a101650a <=( a101649a  and  a101646a );
 a101653a <=( (not A300)  and  (not A299) );
 a101656a <=( A302  and  (not A301) );
 a101657a <=( a101656a  and  a101653a );
 a101658a <=( a101657a  and  a101650a );
 a101661a <=( (not A169)  and  (not A170) );
 a101664a <=( (not A167)  and  (not A168) );
 a101665a <=( a101664a  and  a101661a );
 a101668a <=( A201  and  A166 );
 a101671a <=( A203  and  (not A202) );
 a101672a <=( a101671a  and  a101668a );
 a101673a <=( a101672a  and  a101665a );
 a101676a <=( (not A268)  and  A267 );
 a101679a <=( (not A298)  and  A269 );
 a101680a <=( a101679a  and  a101676a );
 a101683a <=( (not A300)  and  A299 );
 a101686a <=( A302  and  (not A301) );
 a101687a <=( a101686a  and  a101683a );
 a101688a <=( a101687a  and  a101680a );
 a101691a <=( (not A169)  and  (not A170) );
 a101694a <=( (not A167)  and  (not A168) );
 a101695a <=( a101694a  and  a101691a );
 a101698a <=( A201  and  A166 );
 a101701a <=( A203  and  (not A202) );
 a101702a <=( a101701a  and  a101698a );
 a101703a <=( a101702a  and  a101695a );
 a101706a <=( A266  and  (not A265) );
 a101709a <=( (not A268)  and  (not A267) );
 a101710a <=( a101709a  and  a101706a );
 a101713a <=( A300  and  A269 );
 a101716a <=( A302  and  (not A301) );
 a101717a <=( a101716a  and  a101713a );
 a101718a <=( a101717a  and  a101710a );
 a101721a <=( (not A169)  and  (not A170) );
 a101724a <=( (not A167)  and  (not A168) );
 a101725a <=( a101724a  and  a101721a );
 a101728a <=( A201  and  A166 );
 a101731a <=( A203  and  (not A202) );
 a101732a <=( a101731a  and  a101728a );
 a101733a <=( a101732a  and  a101725a );
 a101736a <=( (not A266)  and  A265 );
 a101739a <=( (not A268)  and  (not A267) );
 a101740a <=( a101739a  and  a101736a );
 a101743a <=( A300  and  A269 );
 a101746a <=( A302  and  (not A301) );
 a101747a <=( a101746a  and  a101743a );
 a101748a <=( a101747a  and  a101740a );
 a101751a <=( A166  and  A167 );
 a101754a <=( A200  and  (not A199) );
 a101755a <=( a101754a  and  a101751a );
 a101758a <=( (not A202)  and  (not A201) );
 a101761a <=( (not A265)  and  A203 );
 a101762a <=( a101761a  and  a101758a );
 a101763a <=( a101762a  and  a101755a );
 a101766a <=( (not A267)  and  A266 );
 a101769a <=( A269  and  (not A268) );
 a101770a <=( a101769a  and  a101766a );
 a101773a <=( (not A299)  and  A298 );
 a101777a <=( A302  and  (not A301) );
 a101778a <=( (not A300)  and  a101777a );
 a101779a <=( a101778a  and  a101773a );
 a101780a <=( a101779a  and  a101770a );
 a101783a <=( A166  and  A167 );
 a101786a <=( A200  and  (not A199) );
 a101787a <=( a101786a  and  a101783a );
 a101790a <=( (not A202)  and  (not A201) );
 a101793a <=( (not A265)  and  A203 );
 a101794a <=( a101793a  and  a101790a );
 a101795a <=( a101794a  and  a101787a );
 a101798a <=( (not A267)  and  A266 );
 a101801a <=( A269  and  (not A268) );
 a101802a <=( a101801a  and  a101798a );
 a101805a <=( A299  and  (not A298) );
 a101809a <=( A302  and  (not A301) );
 a101810a <=( (not A300)  and  a101809a );
 a101811a <=( a101810a  and  a101805a );
 a101812a <=( a101811a  and  a101802a );
 a101815a <=( A166  and  A167 );
 a101818a <=( A200  and  (not A199) );
 a101819a <=( a101818a  and  a101815a );
 a101822a <=( (not A202)  and  (not A201) );
 a101825a <=( A265  and  A203 );
 a101826a <=( a101825a  and  a101822a );
 a101827a <=( a101826a  and  a101819a );
 a101830a <=( (not A267)  and  (not A266) );
 a101833a <=( A269  and  (not A268) );
 a101834a <=( a101833a  and  a101830a );
 a101837a <=( (not A299)  and  A298 );
 a101841a <=( A302  and  (not A301) );
 a101842a <=( (not A300)  and  a101841a );
 a101843a <=( a101842a  and  a101837a );
 a101844a <=( a101843a  and  a101834a );
 a101847a <=( A166  and  A167 );
 a101850a <=( A200  and  (not A199) );
 a101851a <=( a101850a  and  a101847a );
 a101854a <=( (not A202)  and  (not A201) );
 a101857a <=( A265  and  A203 );
 a101858a <=( a101857a  and  a101854a );
 a101859a <=( a101858a  and  a101851a );
 a101862a <=( (not A267)  and  (not A266) );
 a101865a <=( A269  and  (not A268) );
 a101866a <=( a101865a  and  a101862a );
 a101869a <=( A299  and  (not A298) );
 a101873a <=( A302  and  (not A301) );
 a101874a <=( (not A300)  and  a101873a );
 a101875a <=( a101874a  and  a101869a );
 a101876a <=( a101875a  and  a101866a );
 a101879a <=( A166  and  A167 );
 a101882a <=( (not A200)  and  A199 );
 a101883a <=( a101882a  and  a101879a );
 a101886a <=( (not A202)  and  (not A201) );
 a101889a <=( (not A265)  and  A203 );
 a101890a <=( a101889a  and  a101886a );
 a101891a <=( a101890a  and  a101883a );
 a101894a <=( (not A267)  and  A266 );
 a101897a <=( A269  and  (not A268) );
 a101898a <=( a101897a  and  a101894a );
 a101901a <=( (not A299)  and  A298 );
 a101905a <=( A302  and  (not A301) );
 a101906a <=( (not A300)  and  a101905a );
 a101907a <=( a101906a  and  a101901a );
 a101908a <=( a101907a  and  a101898a );
 a101911a <=( A166  and  A167 );
 a101914a <=( (not A200)  and  A199 );
 a101915a <=( a101914a  and  a101911a );
 a101918a <=( (not A202)  and  (not A201) );
 a101921a <=( (not A265)  and  A203 );
 a101922a <=( a101921a  and  a101918a );
 a101923a <=( a101922a  and  a101915a );
 a101926a <=( (not A267)  and  A266 );
 a101929a <=( A269  and  (not A268) );
 a101930a <=( a101929a  and  a101926a );
 a101933a <=( A299  and  (not A298) );
 a101937a <=( A302  and  (not A301) );
 a101938a <=( (not A300)  and  a101937a );
 a101939a <=( a101938a  and  a101933a );
 a101940a <=( a101939a  and  a101930a );
 a101943a <=( A166  and  A167 );
 a101946a <=( (not A200)  and  A199 );
 a101947a <=( a101946a  and  a101943a );
 a101950a <=( (not A202)  and  (not A201) );
 a101953a <=( A265  and  A203 );
 a101954a <=( a101953a  and  a101950a );
 a101955a <=( a101954a  and  a101947a );
 a101958a <=( (not A267)  and  (not A266) );
 a101961a <=( A269  and  (not A268) );
 a101962a <=( a101961a  and  a101958a );
 a101965a <=( (not A299)  and  A298 );
 a101969a <=( A302  and  (not A301) );
 a101970a <=( (not A300)  and  a101969a );
 a101971a <=( a101970a  and  a101965a );
 a101972a <=( a101971a  and  a101962a );
 a101975a <=( A166  and  A167 );
 a101978a <=( (not A200)  and  A199 );
 a101979a <=( a101978a  and  a101975a );
 a101982a <=( (not A202)  and  (not A201) );
 a101985a <=( A265  and  A203 );
 a101986a <=( a101985a  and  a101982a );
 a101987a <=( a101986a  and  a101979a );
 a101990a <=( (not A267)  and  (not A266) );
 a101993a <=( A269  and  (not A268) );
 a101994a <=( a101993a  and  a101990a );
 a101997a <=( A299  and  (not A298) );
 a102001a <=( A302  and  (not A301) );
 a102002a <=( (not A300)  and  a102001a );
 a102003a <=( a102002a  and  a101997a );
 a102004a <=( a102003a  and  a101994a );
 a102007a <=( (not A166)  and  (not A167) );
 a102010a <=( A200  and  (not A199) );
 a102011a <=( a102010a  and  a102007a );
 a102014a <=( (not A202)  and  (not A201) );
 a102017a <=( (not A265)  and  A203 );
 a102018a <=( a102017a  and  a102014a );
 a102019a <=( a102018a  and  a102011a );
 a102022a <=( (not A267)  and  A266 );
 a102025a <=( A269  and  (not A268) );
 a102026a <=( a102025a  and  a102022a );
 a102029a <=( (not A299)  and  A298 );
 a102033a <=( A302  and  (not A301) );
 a102034a <=( (not A300)  and  a102033a );
 a102035a <=( a102034a  and  a102029a );
 a102036a <=( a102035a  and  a102026a );
 a102039a <=( (not A166)  and  (not A167) );
 a102042a <=( A200  and  (not A199) );
 a102043a <=( a102042a  and  a102039a );
 a102046a <=( (not A202)  and  (not A201) );
 a102049a <=( (not A265)  and  A203 );
 a102050a <=( a102049a  and  a102046a );
 a102051a <=( a102050a  and  a102043a );
 a102054a <=( (not A267)  and  A266 );
 a102057a <=( A269  and  (not A268) );
 a102058a <=( a102057a  and  a102054a );
 a102061a <=( A299  and  (not A298) );
 a102065a <=( A302  and  (not A301) );
 a102066a <=( (not A300)  and  a102065a );
 a102067a <=( a102066a  and  a102061a );
 a102068a <=( a102067a  and  a102058a );
 a102071a <=( (not A166)  and  (not A167) );
 a102074a <=( A200  and  (not A199) );
 a102075a <=( a102074a  and  a102071a );
 a102078a <=( (not A202)  and  (not A201) );
 a102081a <=( A265  and  A203 );
 a102082a <=( a102081a  and  a102078a );
 a102083a <=( a102082a  and  a102075a );
 a102086a <=( (not A267)  and  (not A266) );
 a102089a <=( A269  and  (not A268) );
 a102090a <=( a102089a  and  a102086a );
 a102093a <=( (not A299)  and  A298 );
 a102097a <=( A302  and  (not A301) );
 a102098a <=( (not A300)  and  a102097a );
 a102099a <=( a102098a  and  a102093a );
 a102100a <=( a102099a  and  a102090a );
 a102103a <=( (not A166)  and  (not A167) );
 a102106a <=( A200  and  (not A199) );
 a102107a <=( a102106a  and  a102103a );
 a102110a <=( (not A202)  and  (not A201) );
 a102113a <=( A265  and  A203 );
 a102114a <=( a102113a  and  a102110a );
 a102115a <=( a102114a  and  a102107a );
 a102118a <=( (not A267)  and  (not A266) );
 a102121a <=( A269  and  (not A268) );
 a102122a <=( a102121a  and  a102118a );
 a102125a <=( A299  and  (not A298) );
 a102129a <=( A302  and  (not A301) );
 a102130a <=( (not A300)  and  a102129a );
 a102131a <=( a102130a  and  a102125a );
 a102132a <=( a102131a  and  a102122a );
 a102135a <=( (not A166)  and  (not A167) );
 a102138a <=( (not A200)  and  A199 );
 a102139a <=( a102138a  and  a102135a );
 a102142a <=( (not A202)  and  (not A201) );
 a102145a <=( (not A265)  and  A203 );
 a102146a <=( a102145a  and  a102142a );
 a102147a <=( a102146a  and  a102139a );
 a102150a <=( (not A267)  and  A266 );
 a102153a <=( A269  and  (not A268) );
 a102154a <=( a102153a  and  a102150a );
 a102157a <=( (not A299)  and  A298 );
 a102161a <=( A302  and  (not A301) );
 a102162a <=( (not A300)  and  a102161a );
 a102163a <=( a102162a  and  a102157a );
 a102164a <=( a102163a  and  a102154a );
 a102167a <=( (not A166)  and  (not A167) );
 a102170a <=( (not A200)  and  A199 );
 a102171a <=( a102170a  and  a102167a );
 a102174a <=( (not A202)  and  (not A201) );
 a102177a <=( (not A265)  and  A203 );
 a102178a <=( a102177a  and  a102174a );
 a102179a <=( a102178a  and  a102171a );
 a102182a <=( (not A267)  and  A266 );
 a102185a <=( A269  and  (not A268) );
 a102186a <=( a102185a  and  a102182a );
 a102189a <=( A299  and  (not A298) );
 a102193a <=( A302  and  (not A301) );
 a102194a <=( (not A300)  and  a102193a );
 a102195a <=( a102194a  and  a102189a );
 a102196a <=( a102195a  and  a102186a );
 a102199a <=( (not A166)  and  (not A167) );
 a102202a <=( (not A200)  and  A199 );
 a102203a <=( a102202a  and  a102199a );
 a102206a <=( (not A202)  and  (not A201) );
 a102209a <=( A265  and  A203 );
 a102210a <=( a102209a  and  a102206a );
 a102211a <=( a102210a  and  a102203a );
 a102214a <=( (not A267)  and  (not A266) );
 a102217a <=( A269  and  (not A268) );
 a102218a <=( a102217a  and  a102214a );
 a102221a <=( (not A299)  and  A298 );
 a102225a <=( A302  and  (not A301) );
 a102226a <=( (not A300)  and  a102225a );
 a102227a <=( a102226a  and  a102221a );
 a102228a <=( a102227a  and  a102218a );
 a102231a <=( (not A166)  and  (not A167) );
 a102234a <=( (not A200)  and  A199 );
 a102235a <=( a102234a  and  a102231a );
 a102238a <=( (not A202)  and  (not A201) );
 a102241a <=( A265  and  A203 );
 a102242a <=( a102241a  and  a102238a );
 a102243a <=( a102242a  and  a102235a );
 a102246a <=( (not A267)  and  (not A266) );
 a102249a <=( A269  and  (not A268) );
 a102250a <=( a102249a  and  a102246a );
 a102253a <=( A299  and  (not A298) );
 a102257a <=( A302  and  (not A301) );
 a102258a <=( (not A300)  and  a102257a );
 a102259a <=( a102258a  and  a102253a );
 a102260a <=( a102259a  and  a102250a );
 a102263a <=( (not A168)  and  A170 );
 a102266a <=( A200  and  (not A199) );
 a102267a <=( a102266a  and  a102263a );
 a102270a <=( (not A202)  and  (not A201) );
 a102273a <=( (not A265)  and  A203 );
 a102274a <=( a102273a  and  a102270a );
 a102275a <=( a102274a  and  a102267a );
 a102278a <=( (not A267)  and  A266 );
 a102281a <=( A269  and  (not A268) );
 a102282a <=( a102281a  and  a102278a );
 a102285a <=( (not A299)  and  A298 );
 a102289a <=( A302  and  (not A301) );
 a102290a <=( (not A300)  and  a102289a );
 a102291a <=( a102290a  and  a102285a );
 a102292a <=( a102291a  and  a102282a );
 a102295a <=( (not A168)  and  A170 );
 a102298a <=( A200  and  (not A199) );
 a102299a <=( a102298a  and  a102295a );
 a102302a <=( (not A202)  and  (not A201) );
 a102305a <=( (not A265)  and  A203 );
 a102306a <=( a102305a  and  a102302a );
 a102307a <=( a102306a  and  a102299a );
 a102310a <=( (not A267)  and  A266 );
 a102313a <=( A269  and  (not A268) );
 a102314a <=( a102313a  and  a102310a );
 a102317a <=( A299  and  (not A298) );
 a102321a <=( A302  and  (not A301) );
 a102322a <=( (not A300)  and  a102321a );
 a102323a <=( a102322a  and  a102317a );
 a102324a <=( a102323a  and  a102314a );
 a102327a <=( (not A168)  and  A170 );
 a102330a <=( A200  and  (not A199) );
 a102331a <=( a102330a  and  a102327a );
 a102334a <=( (not A202)  and  (not A201) );
 a102337a <=( A265  and  A203 );
 a102338a <=( a102337a  and  a102334a );
 a102339a <=( a102338a  and  a102331a );
 a102342a <=( (not A267)  and  (not A266) );
 a102345a <=( A269  and  (not A268) );
 a102346a <=( a102345a  and  a102342a );
 a102349a <=( (not A299)  and  A298 );
 a102353a <=( A302  and  (not A301) );
 a102354a <=( (not A300)  and  a102353a );
 a102355a <=( a102354a  and  a102349a );
 a102356a <=( a102355a  and  a102346a );
 a102359a <=( (not A168)  and  A170 );
 a102362a <=( A200  and  (not A199) );
 a102363a <=( a102362a  and  a102359a );
 a102366a <=( (not A202)  and  (not A201) );
 a102369a <=( A265  and  A203 );
 a102370a <=( a102369a  and  a102366a );
 a102371a <=( a102370a  and  a102363a );
 a102374a <=( (not A267)  and  (not A266) );
 a102377a <=( A269  and  (not A268) );
 a102378a <=( a102377a  and  a102374a );
 a102381a <=( A299  and  (not A298) );
 a102385a <=( A302  and  (not A301) );
 a102386a <=( (not A300)  and  a102385a );
 a102387a <=( a102386a  and  a102381a );
 a102388a <=( a102387a  and  a102378a );
 a102391a <=( (not A168)  and  A170 );
 a102394a <=( (not A200)  and  A199 );
 a102395a <=( a102394a  and  a102391a );
 a102398a <=( (not A202)  and  (not A201) );
 a102401a <=( (not A265)  and  A203 );
 a102402a <=( a102401a  and  a102398a );
 a102403a <=( a102402a  and  a102395a );
 a102406a <=( (not A267)  and  A266 );
 a102409a <=( A269  and  (not A268) );
 a102410a <=( a102409a  and  a102406a );
 a102413a <=( (not A299)  and  A298 );
 a102417a <=( A302  and  (not A301) );
 a102418a <=( (not A300)  and  a102417a );
 a102419a <=( a102418a  and  a102413a );
 a102420a <=( a102419a  and  a102410a );
 a102423a <=( (not A168)  and  A170 );
 a102426a <=( (not A200)  and  A199 );
 a102427a <=( a102426a  and  a102423a );
 a102430a <=( (not A202)  and  (not A201) );
 a102433a <=( (not A265)  and  A203 );
 a102434a <=( a102433a  and  a102430a );
 a102435a <=( a102434a  and  a102427a );
 a102438a <=( (not A267)  and  A266 );
 a102441a <=( A269  and  (not A268) );
 a102442a <=( a102441a  and  a102438a );
 a102445a <=( A299  and  (not A298) );
 a102449a <=( A302  and  (not A301) );
 a102450a <=( (not A300)  and  a102449a );
 a102451a <=( a102450a  and  a102445a );
 a102452a <=( a102451a  and  a102442a );
 a102455a <=( (not A168)  and  A170 );
 a102458a <=( (not A200)  and  A199 );
 a102459a <=( a102458a  and  a102455a );
 a102462a <=( (not A202)  and  (not A201) );
 a102465a <=( A265  and  A203 );
 a102466a <=( a102465a  and  a102462a );
 a102467a <=( a102466a  and  a102459a );
 a102470a <=( (not A267)  and  (not A266) );
 a102473a <=( A269  and  (not A268) );
 a102474a <=( a102473a  and  a102470a );
 a102477a <=( (not A299)  and  A298 );
 a102481a <=( A302  and  (not A301) );
 a102482a <=( (not A300)  and  a102481a );
 a102483a <=( a102482a  and  a102477a );
 a102484a <=( a102483a  and  a102474a );
 a102487a <=( (not A168)  and  A170 );
 a102490a <=( (not A200)  and  A199 );
 a102491a <=( a102490a  and  a102487a );
 a102494a <=( (not A202)  and  (not A201) );
 a102497a <=( A265  and  A203 );
 a102498a <=( a102497a  and  a102494a );
 a102499a <=( a102498a  and  a102491a );
 a102502a <=( (not A267)  and  (not A266) );
 a102505a <=( A269  and  (not A268) );
 a102506a <=( a102505a  and  a102502a );
 a102509a <=( A299  and  (not A298) );
 a102513a <=( A302  and  (not A301) );
 a102514a <=( (not A300)  and  a102513a );
 a102515a <=( a102514a  and  a102509a );
 a102516a <=( a102515a  and  a102506a );
 a102519a <=( (not A168)  and  A169 );
 a102522a <=( A200  and  (not A199) );
 a102523a <=( a102522a  and  a102519a );
 a102526a <=( (not A202)  and  (not A201) );
 a102529a <=( (not A265)  and  A203 );
 a102530a <=( a102529a  and  a102526a );
 a102531a <=( a102530a  and  a102523a );
 a102534a <=( (not A267)  and  A266 );
 a102537a <=( A269  and  (not A268) );
 a102538a <=( a102537a  and  a102534a );
 a102541a <=( (not A299)  and  A298 );
 a102545a <=( A302  and  (not A301) );
 a102546a <=( (not A300)  and  a102545a );
 a102547a <=( a102546a  and  a102541a );
 a102548a <=( a102547a  and  a102538a );
 a102551a <=( (not A168)  and  A169 );
 a102554a <=( A200  and  (not A199) );
 a102555a <=( a102554a  and  a102551a );
 a102558a <=( (not A202)  and  (not A201) );
 a102561a <=( (not A265)  and  A203 );
 a102562a <=( a102561a  and  a102558a );
 a102563a <=( a102562a  and  a102555a );
 a102566a <=( (not A267)  and  A266 );
 a102569a <=( A269  and  (not A268) );
 a102570a <=( a102569a  and  a102566a );
 a102573a <=( A299  and  (not A298) );
 a102577a <=( A302  and  (not A301) );
 a102578a <=( (not A300)  and  a102577a );
 a102579a <=( a102578a  and  a102573a );
 a102580a <=( a102579a  and  a102570a );
 a102583a <=( (not A168)  and  A169 );
 a102586a <=( A200  and  (not A199) );
 a102587a <=( a102586a  and  a102583a );
 a102590a <=( (not A202)  and  (not A201) );
 a102593a <=( A265  and  A203 );
 a102594a <=( a102593a  and  a102590a );
 a102595a <=( a102594a  and  a102587a );
 a102598a <=( (not A267)  and  (not A266) );
 a102601a <=( A269  and  (not A268) );
 a102602a <=( a102601a  and  a102598a );
 a102605a <=( (not A299)  and  A298 );
 a102609a <=( A302  and  (not A301) );
 a102610a <=( (not A300)  and  a102609a );
 a102611a <=( a102610a  and  a102605a );
 a102612a <=( a102611a  and  a102602a );
 a102615a <=( (not A168)  and  A169 );
 a102618a <=( A200  and  (not A199) );
 a102619a <=( a102618a  and  a102615a );
 a102622a <=( (not A202)  and  (not A201) );
 a102625a <=( A265  and  A203 );
 a102626a <=( a102625a  and  a102622a );
 a102627a <=( a102626a  and  a102619a );
 a102630a <=( (not A267)  and  (not A266) );
 a102633a <=( A269  and  (not A268) );
 a102634a <=( a102633a  and  a102630a );
 a102637a <=( A299  and  (not A298) );
 a102641a <=( A302  and  (not A301) );
 a102642a <=( (not A300)  and  a102641a );
 a102643a <=( a102642a  and  a102637a );
 a102644a <=( a102643a  and  a102634a );
 a102647a <=( (not A168)  and  A169 );
 a102650a <=( (not A200)  and  A199 );
 a102651a <=( a102650a  and  a102647a );
 a102654a <=( (not A202)  and  (not A201) );
 a102657a <=( (not A265)  and  A203 );
 a102658a <=( a102657a  and  a102654a );
 a102659a <=( a102658a  and  a102651a );
 a102662a <=( (not A267)  and  A266 );
 a102665a <=( A269  and  (not A268) );
 a102666a <=( a102665a  and  a102662a );
 a102669a <=( (not A299)  and  A298 );
 a102673a <=( A302  and  (not A301) );
 a102674a <=( (not A300)  and  a102673a );
 a102675a <=( a102674a  and  a102669a );
 a102676a <=( a102675a  and  a102666a );
 a102679a <=( (not A168)  and  A169 );
 a102682a <=( (not A200)  and  A199 );
 a102683a <=( a102682a  and  a102679a );
 a102686a <=( (not A202)  and  (not A201) );
 a102689a <=( (not A265)  and  A203 );
 a102690a <=( a102689a  and  a102686a );
 a102691a <=( a102690a  and  a102683a );
 a102694a <=( (not A267)  and  A266 );
 a102697a <=( A269  and  (not A268) );
 a102698a <=( a102697a  and  a102694a );
 a102701a <=( A299  and  (not A298) );
 a102705a <=( A302  and  (not A301) );
 a102706a <=( (not A300)  and  a102705a );
 a102707a <=( a102706a  and  a102701a );
 a102708a <=( a102707a  and  a102698a );
 a102711a <=( (not A168)  and  A169 );
 a102714a <=( (not A200)  and  A199 );
 a102715a <=( a102714a  and  a102711a );
 a102718a <=( (not A202)  and  (not A201) );
 a102721a <=( A265  and  A203 );
 a102722a <=( a102721a  and  a102718a );
 a102723a <=( a102722a  and  a102715a );
 a102726a <=( (not A267)  and  (not A266) );
 a102729a <=( A269  and  (not A268) );
 a102730a <=( a102729a  and  a102726a );
 a102733a <=( (not A299)  and  A298 );
 a102737a <=( A302  and  (not A301) );
 a102738a <=( (not A300)  and  a102737a );
 a102739a <=( a102738a  and  a102733a );
 a102740a <=( a102739a  and  a102730a );
 a102743a <=( (not A168)  and  A169 );
 a102746a <=( (not A200)  and  A199 );
 a102747a <=( a102746a  and  a102743a );
 a102750a <=( (not A202)  and  (not A201) );
 a102753a <=( A265  and  A203 );
 a102754a <=( a102753a  and  a102750a );
 a102755a <=( a102754a  and  a102747a );
 a102758a <=( (not A267)  and  (not A266) );
 a102761a <=( A269  and  (not A268) );
 a102762a <=( a102761a  and  a102758a );
 a102765a <=( A299  and  (not A298) );
 a102769a <=( A302  and  (not A301) );
 a102770a <=( (not A300)  and  a102769a );
 a102771a <=( a102770a  and  a102765a );
 a102772a <=( a102771a  and  a102762a );
 a102775a <=( (not A169)  and  (not A170) );
 a102778a <=( (not A199)  and  A168 );
 a102779a <=( a102778a  and  a102775a );
 a102782a <=( A201  and  A200 );
 a102785a <=( (not A265)  and  A202 );
 a102786a <=( a102785a  and  a102782a );
 a102787a <=( a102786a  and  a102779a );
 a102790a <=( (not A267)  and  A266 );
 a102793a <=( A269  and  (not A268) );
 a102794a <=( a102793a  and  a102790a );
 a102797a <=( (not A299)  and  A298 );
 a102801a <=( A302  and  (not A301) );
 a102802a <=( (not A300)  and  a102801a );
 a102803a <=( a102802a  and  a102797a );
 a102804a <=( a102803a  and  a102794a );
 a102807a <=( (not A169)  and  (not A170) );
 a102810a <=( (not A199)  and  A168 );
 a102811a <=( a102810a  and  a102807a );
 a102814a <=( A201  and  A200 );
 a102817a <=( (not A265)  and  A202 );
 a102818a <=( a102817a  and  a102814a );
 a102819a <=( a102818a  and  a102811a );
 a102822a <=( (not A267)  and  A266 );
 a102825a <=( A269  and  (not A268) );
 a102826a <=( a102825a  and  a102822a );
 a102829a <=( A299  and  (not A298) );
 a102833a <=( A302  and  (not A301) );
 a102834a <=( (not A300)  and  a102833a );
 a102835a <=( a102834a  and  a102829a );
 a102836a <=( a102835a  and  a102826a );
 a102839a <=( (not A169)  and  (not A170) );
 a102842a <=( (not A199)  and  A168 );
 a102843a <=( a102842a  and  a102839a );
 a102846a <=( A201  and  A200 );
 a102849a <=( A265  and  A202 );
 a102850a <=( a102849a  and  a102846a );
 a102851a <=( a102850a  and  a102843a );
 a102854a <=( (not A267)  and  (not A266) );
 a102857a <=( A269  and  (not A268) );
 a102858a <=( a102857a  and  a102854a );
 a102861a <=( (not A299)  and  A298 );
 a102865a <=( A302  and  (not A301) );
 a102866a <=( (not A300)  and  a102865a );
 a102867a <=( a102866a  and  a102861a );
 a102868a <=( a102867a  and  a102858a );
 a102871a <=( (not A169)  and  (not A170) );
 a102874a <=( (not A199)  and  A168 );
 a102875a <=( a102874a  and  a102871a );
 a102878a <=( A201  and  A200 );
 a102881a <=( A265  and  A202 );
 a102882a <=( a102881a  and  a102878a );
 a102883a <=( a102882a  and  a102875a );
 a102886a <=( (not A267)  and  (not A266) );
 a102889a <=( A269  and  (not A268) );
 a102890a <=( a102889a  and  a102886a );
 a102893a <=( A299  and  (not A298) );
 a102897a <=( A302  and  (not A301) );
 a102898a <=( (not A300)  and  a102897a );
 a102899a <=( a102898a  and  a102893a );
 a102900a <=( a102899a  and  a102890a );
 a102903a <=( (not A169)  and  (not A170) );
 a102906a <=( (not A199)  and  A168 );
 a102907a <=( a102906a  and  a102903a );
 a102910a <=( A201  and  A200 );
 a102913a <=( (not A265)  and  (not A203) );
 a102914a <=( a102913a  and  a102910a );
 a102915a <=( a102914a  and  a102907a );
 a102918a <=( (not A267)  and  A266 );
 a102921a <=( A269  and  (not A268) );
 a102922a <=( a102921a  and  a102918a );
 a102925a <=( (not A299)  and  A298 );
 a102929a <=( A302  and  (not A301) );
 a102930a <=( (not A300)  and  a102929a );
 a102931a <=( a102930a  and  a102925a );
 a102932a <=( a102931a  and  a102922a );
 a102935a <=( (not A169)  and  (not A170) );
 a102938a <=( (not A199)  and  A168 );
 a102939a <=( a102938a  and  a102935a );
 a102942a <=( A201  and  A200 );
 a102945a <=( (not A265)  and  (not A203) );
 a102946a <=( a102945a  and  a102942a );
 a102947a <=( a102946a  and  a102939a );
 a102950a <=( (not A267)  and  A266 );
 a102953a <=( A269  and  (not A268) );
 a102954a <=( a102953a  and  a102950a );
 a102957a <=( A299  and  (not A298) );
 a102961a <=( A302  and  (not A301) );
 a102962a <=( (not A300)  and  a102961a );
 a102963a <=( a102962a  and  a102957a );
 a102964a <=( a102963a  and  a102954a );
 a102967a <=( (not A169)  and  (not A170) );
 a102970a <=( (not A199)  and  A168 );
 a102971a <=( a102970a  and  a102967a );
 a102974a <=( A201  and  A200 );
 a102977a <=( A265  and  (not A203) );
 a102978a <=( a102977a  and  a102974a );
 a102979a <=( a102978a  and  a102971a );
 a102982a <=( (not A267)  and  (not A266) );
 a102985a <=( A269  and  (not A268) );
 a102986a <=( a102985a  and  a102982a );
 a102989a <=( (not A299)  and  A298 );
 a102993a <=( A302  and  (not A301) );
 a102994a <=( (not A300)  and  a102993a );
 a102995a <=( a102994a  and  a102989a );
 a102996a <=( a102995a  and  a102986a );
 a102999a <=( (not A169)  and  (not A170) );
 a103002a <=( (not A199)  and  A168 );
 a103003a <=( a103002a  and  a102999a );
 a103006a <=( A201  and  A200 );
 a103009a <=( A265  and  (not A203) );
 a103010a <=( a103009a  and  a103006a );
 a103011a <=( a103010a  and  a103003a );
 a103014a <=( (not A267)  and  (not A266) );
 a103017a <=( A269  and  (not A268) );
 a103018a <=( a103017a  and  a103014a );
 a103021a <=( A299  and  (not A298) );
 a103025a <=( A302  and  (not A301) );
 a103026a <=( (not A300)  and  a103025a );
 a103027a <=( a103026a  and  a103021a );
 a103028a <=( a103027a  and  a103018a );
 a103031a <=( (not A169)  and  (not A170) );
 a103034a <=( (not A199)  and  A168 );
 a103035a <=( a103034a  and  a103031a );
 a103038a <=( (not A201)  and  A200 );
 a103041a <=( A203  and  (not A202) );
 a103042a <=( a103041a  and  a103038a );
 a103043a <=( a103042a  and  a103035a );
 a103046a <=( A266  and  (not A265) );
 a103049a <=( A268  and  A267 );
 a103050a <=( a103049a  and  a103046a );
 a103053a <=( (not A299)  and  A298 );
 a103057a <=( A302  and  (not A301) );
 a103058a <=( (not A300)  and  a103057a );
 a103059a <=( a103058a  and  a103053a );
 a103060a <=( a103059a  and  a103050a );
 a103063a <=( (not A169)  and  (not A170) );
 a103066a <=( (not A199)  and  A168 );
 a103067a <=( a103066a  and  a103063a );
 a103070a <=( (not A201)  and  A200 );
 a103073a <=( A203  and  (not A202) );
 a103074a <=( a103073a  and  a103070a );
 a103075a <=( a103074a  and  a103067a );
 a103078a <=( A266  and  (not A265) );
 a103081a <=( A268  and  A267 );
 a103082a <=( a103081a  and  a103078a );
 a103085a <=( A299  and  (not A298) );
 a103089a <=( A302  and  (not A301) );
 a103090a <=( (not A300)  and  a103089a );
 a103091a <=( a103090a  and  a103085a );
 a103092a <=( a103091a  and  a103082a );
 a103095a <=( (not A169)  and  (not A170) );
 a103098a <=( (not A199)  and  A168 );
 a103099a <=( a103098a  and  a103095a );
 a103102a <=( (not A201)  and  A200 );
 a103105a <=( A203  and  (not A202) );
 a103106a <=( a103105a  and  a103102a );
 a103107a <=( a103106a  and  a103099a );
 a103110a <=( A266  and  (not A265) );
 a103113a <=( (not A269)  and  A267 );
 a103114a <=( a103113a  and  a103110a );
 a103117a <=( (not A299)  and  A298 );
 a103121a <=( A302  and  (not A301) );
 a103122a <=( (not A300)  and  a103121a );
 a103123a <=( a103122a  and  a103117a );
 a103124a <=( a103123a  and  a103114a );
 a103127a <=( (not A169)  and  (not A170) );
 a103130a <=( (not A199)  and  A168 );
 a103131a <=( a103130a  and  a103127a );
 a103134a <=( (not A201)  and  A200 );
 a103137a <=( A203  and  (not A202) );
 a103138a <=( a103137a  and  a103134a );
 a103139a <=( a103138a  and  a103131a );
 a103142a <=( A266  and  (not A265) );
 a103145a <=( (not A269)  and  A267 );
 a103146a <=( a103145a  and  a103142a );
 a103149a <=( A299  and  (not A298) );
 a103153a <=( A302  and  (not A301) );
 a103154a <=( (not A300)  and  a103153a );
 a103155a <=( a103154a  and  a103149a );
 a103156a <=( a103155a  and  a103146a );
 a103159a <=( (not A169)  and  (not A170) );
 a103162a <=( (not A199)  and  A168 );
 a103163a <=( a103162a  and  a103159a );
 a103166a <=( (not A201)  and  A200 );
 a103169a <=( A203  and  (not A202) );
 a103170a <=( a103169a  and  a103166a );
 a103171a <=( a103170a  and  a103163a );
 a103174a <=( A266  and  (not A265) );
 a103177a <=( (not A268)  and  (not A267) );
 a103178a <=( a103177a  and  a103174a );
 a103181a <=( A298  and  A269 );
 a103185a <=( A301  and  A300 );
 a103186a <=( (not A299)  and  a103185a );
 a103187a <=( a103186a  and  a103181a );
 a103188a <=( a103187a  and  a103178a );
 a103191a <=( (not A169)  and  (not A170) );
 a103194a <=( (not A199)  and  A168 );
 a103195a <=( a103194a  and  a103191a );
 a103198a <=( (not A201)  and  A200 );
 a103201a <=( A203  and  (not A202) );
 a103202a <=( a103201a  and  a103198a );
 a103203a <=( a103202a  and  a103195a );
 a103206a <=( A266  and  (not A265) );
 a103209a <=( (not A268)  and  (not A267) );
 a103210a <=( a103209a  and  a103206a );
 a103213a <=( A298  and  A269 );
 a103217a <=( (not A302)  and  A300 );
 a103218a <=( (not A299)  and  a103217a );
 a103219a <=( a103218a  and  a103213a );
 a103220a <=( a103219a  and  a103210a );
 a103223a <=( (not A169)  and  (not A170) );
 a103226a <=( (not A199)  and  A168 );
 a103227a <=( a103226a  and  a103223a );
 a103230a <=( (not A201)  and  A200 );
 a103233a <=( A203  and  (not A202) );
 a103234a <=( a103233a  and  a103230a );
 a103235a <=( a103234a  and  a103227a );
 a103238a <=( A266  and  (not A265) );
 a103241a <=( (not A268)  and  (not A267) );
 a103242a <=( a103241a  and  a103238a );
 a103245a <=( (not A298)  and  A269 );
 a103249a <=( A301  and  A300 );
 a103250a <=( A299  and  a103249a );
 a103251a <=( a103250a  and  a103245a );
 a103252a <=( a103251a  and  a103242a );
 a103255a <=( (not A169)  and  (not A170) );
 a103258a <=( (not A199)  and  A168 );
 a103259a <=( a103258a  and  a103255a );
 a103262a <=( (not A201)  and  A200 );
 a103265a <=( A203  and  (not A202) );
 a103266a <=( a103265a  and  a103262a );
 a103267a <=( a103266a  and  a103259a );
 a103270a <=( A266  and  (not A265) );
 a103273a <=( (not A268)  and  (not A267) );
 a103274a <=( a103273a  and  a103270a );
 a103277a <=( (not A298)  and  A269 );
 a103281a <=( (not A302)  and  A300 );
 a103282a <=( A299  and  a103281a );
 a103283a <=( a103282a  and  a103277a );
 a103284a <=( a103283a  and  a103274a );
 a103287a <=( (not A169)  and  (not A170) );
 a103290a <=( (not A199)  and  A168 );
 a103291a <=( a103290a  and  a103287a );
 a103294a <=( (not A201)  and  A200 );
 a103297a <=( A203  and  (not A202) );
 a103298a <=( a103297a  and  a103294a );
 a103299a <=( a103298a  and  a103291a );
 a103302a <=( (not A266)  and  A265 );
 a103305a <=( A268  and  A267 );
 a103306a <=( a103305a  and  a103302a );
 a103309a <=( (not A299)  and  A298 );
 a103313a <=( A302  and  (not A301) );
 a103314a <=( (not A300)  and  a103313a );
 a103315a <=( a103314a  and  a103309a );
 a103316a <=( a103315a  and  a103306a );
 a103319a <=( (not A169)  and  (not A170) );
 a103322a <=( (not A199)  and  A168 );
 a103323a <=( a103322a  and  a103319a );
 a103326a <=( (not A201)  and  A200 );
 a103329a <=( A203  and  (not A202) );
 a103330a <=( a103329a  and  a103326a );
 a103331a <=( a103330a  and  a103323a );
 a103334a <=( (not A266)  and  A265 );
 a103337a <=( A268  and  A267 );
 a103338a <=( a103337a  and  a103334a );
 a103341a <=( A299  and  (not A298) );
 a103345a <=( A302  and  (not A301) );
 a103346a <=( (not A300)  and  a103345a );
 a103347a <=( a103346a  and  a103341a );
 a103348a <=( a103347a  and  a103338a );
 a103351a <=( (not A169)  and  (not A170) );
 a103354a <=( (not A199)  and  A168 );
 a103355a <=( a103354a  and  a103351a );
 a103358a <=( (not A201)  and  A200 );
 a103361a <=( A203  and  (not A202) );
 a103362a <=( a103361a  and  a103358a );
 a103363a <=( a103362a  and  a103355a );
 a103366a <=( (not A266)  and  A265 );
 a103369a <=( (not A269)  and  A267 );
 a103370a <=( a103369a  and  a103366a );
 a103373a <=( (not A299)  and  A298 );
 a103377a <=( A302  and  (not A301) );
 a103378a <=( (not A300)  and  a103377a );
 a103379a <=( a103378a  and  a103373a );
 a103380a <=( a103379a  and  a103370a );
 a103383a <=( (not A169)  and  (not A170) );
 a103386a <=( (not A199)  and  A168 );
 a103387a <=( a103386a  and  a103383a );
 a103390a <=( (not A201)  and  A200 );
 a103393a <=( A203  and  (not A202) );
 a103394a <=( a103393a  and  a103390a );
 a103395a <=( a103394a  and  a103387a );
 a103398a <=( (not A266)  and  A265 );
 a103401a <=( (not A269)  and  A267 );
 a103402a <=( a103401a  and  a103398a );
 a103405a <=( A299  and  (not A298) );
 a103409a <=( A302  and  (not A301) );
 a103410a <=( (not A300)  and  a103409a );
 a103411a <=( a103410a  and  a103405a );
 a103412a <=( a103411a  and  a103402a );
 a103415a <=( (not A169)  and  (not A170) );
 a103418a <=( (not A199)  and  A168 );
 a103419a <=( a103418a  and  a103415a );
 a103422a <=( (not A201)  and  A200 );
 a103425a <=( A203  and  (not A202) );
 a103426a <=( a103425a  and  a103422a );
 a103427a <=( a103426a  and  a103419a );
 a103430a <=( (not A266)  and  A265 );
 a103433a <=( (not A268)  and  (not A267) );
 a103434a <=( a103433a  and  a103430a );
 a103437a <=( A298  and  A269 );
 a103441a <=( A301  and  A300 );
 a103442a <=( (not A299)  and  a103441a );
 a103443a <=( a103442a  and  a103437a );
 a103444a <=( a103443a  and  a103434a );
 a103447a <=( (not A169)  and  (not A170) );
 a103450a <=( (not A199)  and  A168 );
 a103451a <=( a103450a  and  a103447a );
 a103454a <=( (not A201)  and  A200 );
 a103457a <=( A203  and  (not A202) );
 a103458a <=( a103457a  and  a103454a );
 a103459a <=( a103458a  and  a103451a );
 a103462a <=( (not A266)  and  A265 );
 a103465a <=( (not A268)  and  (not A267) );
 a103466a <=( a103465a  and  a103462a );
 a103469a <=( A298  and  A269 );
 a103473a <=( (not A302)  and  A300 );
 a103474a <=( (not A299)  and  a103473a );
 a103475a <=( a103474a  and  a103469a );
 a103476a <=( a103475a  and  a103466a );
 a103479a <=( (not A169)  and  (not A170) );
 a103482a <=( (not A199)  and  A168 );
 a103483a <=( a103482a  and  a103479a );
 a103486a <=( (not A201)  and  A200 );
 a103489a <=( A203  and  (not A202) );
 a103490a <=( a103489a  and  a103486a );
 a103491a <=( a103490a  and  a103483a );
 a103494a <=( (not A266)  and  A265 );
 a103497a <=( (not A268)  and  (not A267) );
 a103498a <=( a103497a  and  a103494a );
 a103501a <=( (not A298)  and  A269 );
 a103505a <=( A301  and  A300 );
 a103506a <=( A299  and  a103505a );
 a103507a <=( a103506a  and  a103501a );
 a103508a <=( a103507a  and  a103498a );
 a103511a <=( (not A169)  and  (not A170) );
 a103514a <=( (not A199)  and  A168 );
 a103515a <=( a103514a  and  a103511a );
 a103518a <=( (not A201)  and  A200 );
 a103521a <=( A203  and  (not A202) );
 a103522a <=( a103521a  and  a103518a );
 a103523a <=( a103522a  and  a103515a );
 a103526a <=( (not A266)  and  A265 );
 a103529a <=( (not A268)  and  (not A267) );
 a103530a <=( a103529a  and  a103526a );
 a103533a <=( (not A298)  and  A269 );
 a103537a <=( (not A302)  and  A300 );
 a103538a <=( A299  and  a103537a );
 a103539a <=( a103538a  and  a103533a );
 a103540a <=( a103539a  and  a103530a );
 a103543a <=( (not A169)  and  (not A170) );
 a103546a <=( A199  and  A168 );
 a103547a <=( a103546a  and  a103543a );
 a103550a <=( A201  and  (not A200) );
 a103553a <=( (not A265)  and  A202 );
 a103554a <=( a103553a  and  a103550a );
 a103555a <=( a103554a  and  a103547a );
 a103558a <=( (not A267)  and  A266 );
 a103561a <=( A269  and  (not A268) );
 a103562a <=( a103561a  and  a103558a );
 a103565a <=( (not A299)  and  A298 );
 a103569a <=( A302  and  (not A301) );
 a103570a <=( (not A300)  and  a103569a );
 a103571a <=( a103570a  and  a103565a );
 a103572a <=( a103571a  and  a103562a );
 a103575a <=( (not A169)  and  (not A170) );
 a103578a <=( A199  and  A168 );
 a103579a <=( a103578a  and  a103575a );
 a103582a <=( A201  and  (not A200) );
 a103585a <=( (not A265)  and  A202 );
 a103586a <=( a103585a  and  a103582a );
 a103587a <=( a103586a  and  a103579a );
 a103590a <=( (not A267)  and  A266 );
 a103593a <=( A269  and  (not A268) );
 a103594a <=( a103593a  and  a103590a );
 a103597a <=( A299  and  (not A298) );
 a103601a <=( A302  and  (not A301) );
 a103602a <=( (not A300)  and  a103601a );
 a103603a <=( a103602a  and  a103597a );
 a103604a <=( a103603a  and  a103594a );
 a103607a <=( (not A169)  and  (not A170) );
 a103610a <=( A199  and  A168 );
 a103611a <=( a103610a  and  a103607a );
 a103614a <=( A201  and  (not A200) );
 a103617a <=( A265  and  A202 );
 a103618a <=( a103617a  and  a103614a );
 a103619a <=( a103618a  and  a103611a );
 a103622a <=( (not A267)  and  (not A266) );
 a103625a <=( A269  and  (not A268) );
 a103626a <=( a103625a  and  a103622a );
 a103629a <=( (not A299)  and  A298 );
 a103633a <=( A302  and  (not A301) );
 a103634a <=( (not A300)  and  a103633a );
 a103635a <=( a103634a  and  a103629a );
 a103636a <=( a103635a  and  a103626a );
 a103639a <=( (not A169)  and  (not A170) );
 a103642a <=( A199  and  A168 );
 a103643a <=( a103642a  and  a103639a );
 a103646a <=( A201  and  (not A200) );
 a103649a <=( A265  and  A202 );
 a103650a <=( a103649a  and  a103646a );
 a103651a <=( a103650a  and  a103643a );
 a103654a <=( (not A267)  and  (not A266) );
 a103657a <=( A269  and  (not A268) );
 a103658a <=( a103657a  and  a103654a );
 a103661a <=( A299  and  (not A298) );
 a103665a <=( A302  and  (not A301) );
 a103666a <=( (not A300)  and  a103665a );
 a103667a <=( a103666a  and  a103661a );
 a103668a <=( a103667a  and  a103658a );
 a103671a <=( (not A169)  and  (not A170) );
 a103674a <=( A199  and  A168 );
 a103675a <=( a103674a  and  a103671a );
 a103678a <=( A201  and  (not A200) );
 a103681a <=( (not A265)  and  (not A203) );
 a103682a <=( a103681a  and  a103678a );
 a103683a <=( a103682a  and  a103675a );
 a103686a <=( (not A267)  and  A266 );
 a103689a <=( A269  and  (not A268) );
 a103690a <=( a103689a  and  a103686a );
 a103693a <=( (not A299)  and  A298 );
 a103697a <=( A302  and  (not A301) );
 a103698a <=( (not A300)  and  a103697a );
 a103699a <=( a103698a  and  a103693a );
 a103700a <=( a103699a  and  a103690a );
 a103703a <=( (not A169)  and  (not A170) );
 a103706a <=( A199  and  A168 );
 a103707a <=( a103706a  and  a103703a );
 a103710a <=( A201  and  (not A200) );
 a103713a <=( (not A265)  and  (not A203) );
 a103714a <=( a103713a  and  a103710a );
 a103715a <=( a103714a  and  a103707a );
 a103718a <=( (not A267)  and  A266 );
 a103721a <=( A269  and  (not A268) );
 a103722a <=( a103721a  and  a103718a );
 a103725a <=( A299  and  (not A298) );
 a103729a <=( A302  and  (not A301) );
 a103730a <=( (not A300)  and  a103729a );
 a103731a <=( a103730a  and  a103725a );
 a103732a <=( a103731a  and  a103722a );
 a103735a <=( (not A169)  and  (not A170) );
 a103738a <=( A199  and  A168 );
 a103739a <=( a103738a  and  a103735a );
 a103742a <=( A201  and  (not A200) );
 a103745a <=( A265  and  (not A203) );
 a103746a <=( a103745a  and  a103742a );
 a103747a <=( a103746a  and  a103739a );
 a103750a <=( (not A267)  and  (not A266) );
 a103753a <=( A269  and  (not A268) );
 a103754a <=( a103753a  and  a103750a );
 a103757a <=( (not A299)  and  A298 );
 a103761a <=( A302  and  (not A301) );
 a103762a <=( (not A300)  and  a103761a );
 a103763a <=( a103762a  and  a103757a );
 a103764a <=( a103763a  and  a103754a );
 a103767a <=( (not A169)  and  (not A170) );
 a103770a <=( A199  and  A168 );
 a103771a <=( a103770a  and  a103767a );
 a103774a <=( A201  and  (not A200) );
 a103777a <=( A265  and  (not A203) );
 a103778a <=( a103777a  and  a103774a );
 a103779a <=( a103778a  and  a103771a );
 a103782a <=( (not A267)  and  (not A266) );
 a103785a <=( A269  and  (not A268) );
 a103786a <=( a103785a  and  a103782a );
 a103789a <=( A299  and  (not A298) );
 a103793a <=( A302  and  (not A301) );
 a103794a <=( (not A300)  and  a103793a );
 a103795a <=( a103794a  and  a103789a );
 a103796a <=( a103795a  and  a103786a );
 a103799a <=( (not A169)  and  (not A170) );
 a103802a <=( A199  and  A168 );
 a103803a <=( a103802a  and  a103799a );
 a103806a <=( (not A201)  and  (not A200) );
 a103809a <=( A203  and  (not A202) );
 a103810a <=( a103809a  and  a103806a );
 a103811a <=( a103810a  and  a103803a );
 a103814a <=( A266  and  (not A265) );
 a103817a <=( A268  and  A267 );
 a103818a <=( a103817a  and  a103814a );
 a103821a <=( (not A299)  and  A298 );
 a103825a <=( A302  and  (not A301) );
 a103826a <=( (not A300)  and  a103825a );
 a103827a <=( a103826a  and  a103821a );
 a103828a <=( a103827a  and  a103818a );
 a103831a <=( (not A169)  and  (not A170) );
 a103834a <=( A199  and  A168 );
 a103835a <=( a103834a  and  a103831a );
 a103838a <=( (not A201)  and  (not A200) );
 a103841a <=( A203  and  (not A202) );
 a103842a <=( a103841a  and  a103838a );
 a103843a <=( a103842a  and  a103835a );
 a103846a <=( A266  and  (not A265) );
 a103849a <=( A268  and  A267 );
 a103850a <=( a103849a  and  a103846a );
 a103853a <=( A299  and  (not A298) );
 a103857a <=( A302  and  (not A301) );
 a103858a <=( (not A300)  and  a103857a );
 a103859a <=( a103858a  and  a103853a );
 a103860a <=( a103859a  and  a103850a );
 a103863a <=( (not A169)  and  (not A170) );
 a103866a <=( A199  and  A168 );
 a103867a <=( a103866a  and  a103863a );
 a103870a <=( (not A201)  and  (not A200) );
 a103873a <=( A203  and  (not A202) );
 a103874a <=( a103873a  and  a103870a );
 a103875a <=( a103874a  and  a103867a );
 a103878a <=( A266  and  (not A265) );
 a103881a <=( (not A269)  and  A267 );
 a103882a <=( a103881a  and  a103878a );
 a103885a <=( (not A299)  and  A298 );
 a103889a <=( A302  and  (not A301) );
 a103890a <=( (not A300)  and  a103889a );
 a103891a <=( a103890a  and  a103885a );
 a103892a <=( a103891a  and  a103882a );
 a103895a <=( (not A169)  and  (not A170) );
 a103898a <=( A199  and  A168 );
 a103899a <=( a103898a  and  a103895a );
 a103902a <=( (not A201)  and  (not A200) );
 a103905a <=( A203  and  (not A202) );
 a103906a <=( a103905a  and  a103902a );
 a103907a <=( a103906a  and  a103899a );
 a103910a <=( A266  and  (not A265) );
 a103913a <=( (not A269)  and  A267 );
 a103914a <=( a103913a  and  a103910a );
 a103917a <=( A299  and  (not A298) );
 a103921a <=( A302  and  (not A301) );
 a103922a <=( (not A300)  and  a103921a );
 a103923a <=( a103922a  and  a103917a );
 a103924a <=( a103923a  and  a103914a );
 a103927a <=( (not A169)  and  (not A170) );
 a103930a <=( A199  and  A168 );
 a103931a <=( a103930a  and  a103927a );
 a103934a <=( (not A201)  and  (not A200) );
 a103937a <=( A203  and  (not A202) );
 a103938a <=( a103937a  and  a103934a );
 a103939a <=( a103938a  and  a103931a );
 a103942a <=( A266  and  (not A265) );
 a103945a <=( (not A268)  and  (not A267) );
 a103946a <=( a103945a  and  a103942a );
 a103949a <=( A298  and  A269 );
 a103953a <=( A301  and  A300 );
 a103954a <=( (not A299)  and  a103953a );
 a103955a <=( a103954a  and  a103949a );
 a103956a <=( a103955a  and  a103946a );
 a103959a <=( (not A169)  and  (not A170) );
 a103962a <=( A199  and  A168 );
 a103963a <=( a103962a  and  a103959a );
 a103966a <=( (not A201)  and  (not A200) );
 a103969a <=( A203  and  (not A202) );
 a103970a <=( a103969a  and  a103966a );
 a103971a <=( a103970a  and  a103963a );
 a103974a <=( A266  and  (not A265) );
 a103977a <=( (not A268)  and  (not A267) );
 a103978a <=( a103977a  and  a103974a );
 a103981a <=( A298  and  A269 );
 a103985a <=( (not A302)  and  A300 );
 a103986a <=( (not A299)  and  a103985a );
 a103987a <=( a103986a  and  a103981a );
 a103988a <=( a103987a  and  a103978a );
 a103991a <=( (not A169)  and  (not A170) );
 a103994a <=( A199  and  A168 );
 a103995a <=( a103994a  and  a103991a );
 a103998a <=( (not A201)  and  (not A200) );
 a104001a <=( A203  and  (not A202) );
 a104002a <=( a104001a  and  a103998a );
 a104003a <=( a104002a  and  a103995a );
 a104006a <=( A266  and  (not A265) );
 a104009a <=( (not A268)  and  (not A267) );
 a104010a <=( a104009a  and  a104006a );
 a104013a <=( (not A298)  and  A269 );
 a104017a <=( A301  and  A300 );
 a104018a <=( A299  and  a104017a );
 a104019a <=( a104018a  and  a104013a );
 a104020a <=( a104019a  and  a104010a );
 a104023a <=( (not A169)  and  (not A170) );
 a104026a <=( A199  and  A168 );
 a104027a <=( a104026a  and  a104023a );
 a104030a <=( (not A201)  and  (not A200) );
 a104033a <=( A203  and  (not A202) );
 a104034a <=( a104033a  and  a104030a );
 a104035a <=( a104034a  and  a104027a );
 a104038a <=( A266  and  (not A265) );
 a104041a <=( (not A268)  and  (not A267) );
 a104042a <=( a104041a  and  a104038a );
 a104045a <=( (not A298)  and  A269 );
 a104049a <=( (not A302)  and  A300 );
 a104050a <=( A299  and  a104049a );
 a104051a <=( a104050a  and  a104045a );
 a104052a <=( a104051a  and  a104042a );
 a104055a <=( (not A169)  and  (not A170) );
 a104058a <=( A199  and  A168 );
 a104059a <=( a104058a  and  a104055a );
 a104062a <=( (not A201)  and  (not A200) );
 a104065a <=( A203  and  (not A202) );
 a104066a <=( a104065a  and  a104062a );
 a104067a <=( a104066a  and  a104059a );
 a104070a <=( (not A266)  and  A265 );
 a104073a <=( A268  and  A267 );
 a104074a <=( a104073a  and  a104070a );
 a104077a <=( (not A299)  and  A298 );
 a104081a <=( A302  and  (not A301) );
 a104082a <=( (not A300)  and  a104081a );
 a104083a <=( a104082a  and  a104077a );
 a104084a <=( a104083a  and  a104074a );
 a104087a <=( (not A169)  and  (not A170) );
 a104090a <=( A199  and  A168 );
 a104091a <=( a104090a  and  a104087a );
 a104094a <=( (not A201)  and  (not A200) );
 a104097a <=( A203  and  (not A202) );
 a104098a <=( a104097a  and  a104094a );
 a104099a <=( a104098a  and  a104091a );
 a104102a <=( (not A266)  and  A265 );
 a104105a <=( A268  and  A267 );
 a104106a <=( a104105a  and  a104102a );
 a104109a <=( A299  and  (not A298) );
 a104113a <=( A302  and  (not A301) );
 a104114a <=( (not A300)  and  a104113a );
 a104115a <=( a104114a  and  a104109a );
 a104116a <=( a104115a  and  a104106a );
 a104119a <=( (not A169)  and  (not A170) );
 a104122a <=( A199  and  A168 );
 a104123a <=( a104122a  and  a104119a );
 a104126a <=( (not A201)  and  (not A200) );
 a104129a <=( A203  and  (not A202) );
 a104130a <=( a104129a  and  a104126a );
 a104131a <=( a104130a  and  a104123a );
 a104134a <=( (not A266)  and  A265 );
 a104137a <=( (not A269)  and  A267 );
 a104138a <=( a104137a  and  a104134a );
 a104141a <=( (not A299)  and  A298 );
 a104145a <=( A302  and  (not A301) );
 a104146a <=( (not A300)  and  a104145a );
 a104147a <=( a104146a  and  a104141a );
 a104148a <=( a104147a  and  a104138a );
 a104151a <=( (not A169)  and  (not A170) );
 a104154a <=( A199  and  A168 );
 a104155a <=( a104154a  and  a104151a );
 a104158a <=( (not A201)  and  (not A200) );
 a104161a <=( A203  and  (not A202) );
 a104162a <=( a104161a  and  a104158a );
 a104163a <=( a104162a  and  a104155a );
 a104166a <=( (not A266)  and  A265 );
 a104169a <=( (not A269)  and  A267 );
 a104170a <=( a104169a  and  a104166a );
 a104173a <=( A299  and  (not A298) );
 a104177a <=( A302  and  (not A301) );
 a104178a <=( (not A300)  and  a104177a );
 a104179a <=( a104178a  and  a104173a );
 a104180a <=( a104179a  and  a104170a );
 a104183a <=( (not A169)  and  (not A170) );
 a104186a <=( A199  and  A168 );
 a104187a <=( a104186a  and  a104183a );
 a104190a <=( (not A201)  and  (not A200) );
 a104193a <=( A203  and  (not A202) );
 a104194a <=( a104193a  and  a104190a );
 a104195a <=( a104194a  and  a104187a );
 a104198a <=( (not A266)  and  A265 );
 a104201a <=( (not A268)  and  (not A267) );
 a104202a <=( a104201a  and  a104198a );
 a104205a <=( A298  and  A269 );
 a104209a <=( A301  and  A300 );
 a104210a <=( (not A299)  and  a104209a );
 a104211a <=( a104210a  and  a104205a );
 a104212a <=( a104211a  and  a104202a );
 a104215a <=( (not A169)  and  (not A170) );
 a104218a <=( A199  and  A168 );
 a104219a <=( a104218a  and  a104215a );
 a104222a <=( (not A201)  and  (not A200) );
 a104225a <=( A203  and  (not A202) );
 a104226a <=( a104225a  and  a104222a );
 a104227a <=( a104226a  and  a104219a );
 a104230a <=( (not A266)  and  A265 );
 a104233a <=( (not A268)  and  (not A267) );
 a104234a <=( a104233a  and  a104230a );
 a104237a <=( A298  and  A269 );
 a104241a <=( (not A302)  and  A300 );
 a104242a <=( (not A299)  and  a104241a );
 a104243a <=( a104242a  and  a104237a );
 a104244a <=( a104243a  and  a104234a );
 a104247a <=( (not A169)  and  (not A170) );
 a104250a <=( A199  and  A168 );
 a104251a <=( a104250a  and  a104247a );
 a104254a <=( (not A201)  and  (not A200) );
 a104257a <=( A203  and  (not A202) );
 a104258a <=( a104257a  and  a104254a );
 a104259a <=( a104258a  and  a104251a );
 a104262a <=( (not A266)  and  A265 );
 a104265a <=( (not A268)  and  (not A267) );
 a104266a <=( a104265a  and  a104262a );
 a104269a <=( (not A298)  and  A269 );
 a104273a <=( A301  and  A300 );
 a104274a <=( A299  and  a104273a );
 a104275a <=( a104274a  and  a104269a );
 a104276a <=( a104275a  and  a104266a );
 a104279a <=( (not A169)  and  (not A170) );
 a104282a <=( A199  and  A168 );
 a104283a <=( a104282a  and  a104279a );
 a104286a <=( (not A201)  and  (not A200) );
 a104289a <=( A203  and  (not A202) );
 a104290a <=( a104289a  and  a104286a );
 a104291a <=( a104290a  and  a104283a );
 a104294a <=( (not A266)  and  A265 );
 a104297a <=( (not A268)  and  (not A267) );
 a104298a <=( a104297a  and  a104294a );
 a104301a <=( (not A298)  and  A269 );
 a104305a <=( (not A302)  and  A300 );
 a104306a <=( A299  and  a104305a );
 a104307a <=( a104306a  and  a104301a );
 a104308a <=( a104307a  and  a104298a );
 a104311a <=( (not A169)  and  (not A170) );
 a104314a <=( (not A199)  and  A168 );
 a104315a <=( a104314a  and  a104311a );
 a104318a <=( (not A201)  and  A200 );
 a104322a <=( (not A265)  and  A203 );
 a104323a <=( (not A202)  and  a104322a );
 a104324a <=( a104323a  and  a104318a );
 a104325a <=( a104324a  and  a104315a );
 a104328a <=( (not A267)  and  A266 );
 a104331a <=( A269  and  (not A268) );
 a104332a <=( a104331a  and  a104328a );
 a104335a <=( (not A299)  and  A298 );
 a104339a <=( A302  and  (not A301) );
 a104340a <=( (not A300)  and  a104339a );
 a104341a <=( a104340a  and  a104335a );
 a104342a <=( a104341a  and  a104332a );
 a104345a <=( (not A169)  and  (not A170) );
 a104348a <=( (not A199)  and  A168 );
 a104349a <=( a104348a  and  a104345a );
 a104352a <=( (not A201)  and  A200 );
 a104356a <=( (not A265)  and  A203 );
 a104357a <=( (not A202)  and  a104356a );
 a104358a <=( a104357a  and  a104352a );
 a104359a <=( a104358a  and  a104349a );
 a104362a <=( (not A267)  and  A266 );
 a104365a <=( A269  and  (not A268) );
 a104366a <=( a104365a  and  a104362a );
 a104369a <=( A299  and  (not A298) );
 a104373a <=( A302  and  (not A301) );
 a104374a <=( (not A300)  and  a104373a );
 a104375a <=( a104374a  and  a104369a );
 a104376a <=( a104375a  and  a104366a );
 a104379a <=( (not A169)  and  (not A170) );
 a104382a <=( (not A199)  and  A168 );
 a104383a <=( a104382a  and  a104379a );
 a104386a <=( (not A201)  and  A200 );
 a104390a <=( A265  and  A203 );
 a104391a <=( (not A202)  and  a104390a );
 a104392a <=( a104391a  and  a104386a );
 a104393a <=( a104392a  and  a104383a );
 a104396a <=( (not A267)  and  (not A266) );
 a104399a <=( A269  and  (not A268) );
 a104400a <=( a104399a  and  a104396a );
 a104403a <=( (not A299)  and  A298 );
 a104407a <=( A302  and  (not A301) );
 a104408a <=( (not A300)  and  a104407a );
 a104409a <=( a104408a  and  a104403a );
 a104410a <=( a104409a  and  a104400a );
 a104413a <=( (not A169)  and  (not A170) );
 a104416a <=( (not A199)  and  A168 );
 a104417a <=( a104416a  and  a104413a );
 a104420a <=( (not A201)  and  A200 );
 a104424a <=( A265  and  A203 );
 a104425a <=( (not A202)  and  a104424a );
 a104426a <=( a104425a  and  a104420a );
 a104427a <=( a104426a  and  a104417a );
 a104430a <=( (not A267)  and  (not A266) );
 a104433a <=( A269  and  (not A268) );
 a104434a <=( a104433a  and  a104430a );
 a104437a <=( A299  and  (not A298) );
 a104441a <=( A302  and  (not A301) );
 a104442a <=( (not A300)  and  a104441a );
 a104443a <=( a104442a  and  a104437a );
 a104444a <=( a104443a  and  a104434a );
 a104447a <=( (not A169)  and  (not A170) );
 a104450a <=( A199  and  A168 );
 a104451a <=( a104450a  and  a104447a );
 a104454a <=( (not A201)  and  (not A200) );
 a104458a <=( (not A265)  and  A203 );
 a104459a <=( (not A202)  and  a104458a );
 a104460a <=( a104459a  and  a104454a );
 a104461a <=( a104460a  and  a104451a );
 a104464a <=( (not A267)  and  A266 );
 a104467a <=( A269  and  (not A268) );
 a104468a <=( a104467a  and  a104464a );
 a104471a <=( (not A299)  and  A298 );
 a104475a <=( A302  and  (not A301) );
 a104476a <=( (not A300)  and  a104475a );
 a104477a <=( a104476a  and  a104471a );
 a104478a <=( a104477a  and  a104468a );
 a104481a <=( (not A169)  and  (not A170) );
 a104484a <=( A199  and  A168 );
 a104485a <=( a104484a  and  a104481a );
 a104488a <=( (not A201)  and  (not A200) );
 a104492a <=( (not A265)  and  A203 );
 a104493a <=( (not A202)  and  a104492a );
 a104494a <=( a104493a  and  a104488a );
 a104495a <=( a104494a  and  a104485a );
 a104498a <=( (not A267)  and  A266 );
 a104501a <=( A269  and  (not A268) );
 a104502a <=( a104501a  and  a104498a );
 a104505a <=( A299  and  (not A298) );
 a104509a <=( A302  and  (not A301) );
 a104510a <=( (not A300)  and  a104509a );
 a104511a <=( a104510a  and  a104505a );
 a104512a <=( a104511a  and  a104502a );
 a104515a <=( (not A169)  and  (not A170) );
 a104518a <=( A199  and  A168 );
 a104519a <=( a104518a  and  a104515a );
 a104522a <=( (not A201)  and  (not A200) );
 a104526a <=( A265  and  A203 );
 a104527a <=( (not A202)  and  a104526a );
 a104528a <=( a104527a  and  a104522a );
 a104529a <=( a104528a  and  a104519a );
 a104532a <=( (not A267)  and  (not A266) );
 a104535a <=( A269  and  (not A268) );
 a104536a <=( a104535a  and  a104532a );
 a104539a <=( (not A299)  and  A298 );
 a104543a <=( A302  and  (not A301) );
 a104544a <=( (not A300)  and  a104543a );
 a104545a <=( a104544a  and  a104539a );
 a104546a <=( a104545a  and  a104536a );
 a104549a <=( (not A169)  and  (not A170) );
 a104552a <=( A199  and  A168 );
 a104553a <=( a104552a  and  a104549a );
 a104556a <=( (not A201)  and  (not A200) );
 a104560a <=( A265  and  A203 );
 a104561a <=( (not A202)  and  a104560a );
 a104562a <=( a104561a  and  a104556a );
 a104563a <=( a104562a  and  a104553a );
 a104566a <=( (not A267)  and  (not A266) );
 a104569a <=( A269  and  (not A268) );
 a104570a <=( a104569a  and  a104566a );
 a104573a <=( A299  and  (not A298) );
 a104577a <=( A302  and  (not A301) );
 a104578a <=( (not A300)  and  a104577a );
 a104579a <=( a104578a  and  a104573a );
 a104580a <=( a104579a  and  a104570a );


end x25_22x_behav;
