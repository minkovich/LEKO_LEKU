Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_9x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A106: buffer std_logic
);
end x25_9x;

architecture x25_9x_behav of x25_9x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1122a,a1125a,a1126a,a1129a,a1132a,a1133a,a1134a,a1137a,a1140a,a1141a,a1144a,a1148a,a1149a,a1150a,a1151a,a1152a,a1155a,a1158a,a1159a,a1162a,a1165a,a1166a,a1167a,a1170a,a1173a,a1174a,a1177a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1189a,a1192a,a1193a,a1196a,a1199a,a1200a,a1201a,a1204a,a1207a,a1208a,a1211a,a1215a,a1216a,a1217a,a1218a,a1219a,a1222a,a1225a,a1226a,a1229a,a1233a,a1234a,a1235a,a1236a,a1239a,a1242a,a1243a,a1246a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1259a,a1262a,a1263a,a1266a,a1269a,a1270a,a1271a,a1274a,a1277a,a1278a,a1281a,a1285a,a1286a,a1287a,a1288a,a1289a,a1292a,a1295a,a1296a,a1299a,a1303a,a1304a,a1305a,a1306a,a1309a,a1312a,a1313a,a1316a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1328a,a1331a,a1332a,a1335a,a1338a,a1339a,a1340a,a1343a,a1346a,a1347a,a1350a,a1354a,a1355a,a1356a,a1357a,a1358a,a1361a,a1364a,a1365a,a1368a,a1372a,a1373a,a1374a,a1375a,a1378a,a1381a,a1382a,a1385a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1399a,a1402a,a1403a,a1406a,a1409a,a1410a,a1411a,a1414a,a1417a,a1418a,a1421a,a1425a,a1426a,a1427a,a1428a,a1429a,a1432a,a1435a,a1436a,a1439a,a1443a,a1444a,a1445a,a1446a,a1449a,a1452a,a1453a,a1456a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1468a,a1471a,a1472a,a1475a,a1478a,a1479a,a1480a,a1483a,a1486a,a1487a,a1490a,a1494a,a1495a,a1496a,a1497a,a1498a,a1501a,a1504a,a1505a,a1508a,a1512a,a1513a,a1514a,a1515a,a1518a,a1521a,a1522a,a1525a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1538a,a1541a,a1542a,a1545a,a1548a,a1549a,a1550a,a1553a,a1556a,a1557a,a1560a,a1564a,a1565a,a1566a,a1567a,a1568a,a1571a,a1574a,a1575a,a1578a,a1582a,a1583a,a1584a,a1585a,a1588a,a1591a,a1592a,a1595a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1607a,a1610a,a1611a,a1614a,a1617a,a1618a,a1619a,a1622a,a1625a,a1626a,a1629a,a1633a,a1634a,a1635a,a1636a,a1637a,a1640a,a1643a,a1644a,a1647a,a1651a,a1652a,a1653a,a1654a,a1657a,a1660a,a1661a,a1664a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1679a,a1682a,a1683a,a1686a,a1689a,a1690a,a1691a,a1694a,a1697a,a1698a,a1701a,a1705a,a1706a,a1707a,a1708a,a1709a,a1712a,a1715a,a1716a,a1719a,a1723a,a1724a,a1725a,a1726a,a1729a,a1732a,a1733a,a1736a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1748a,a1751a,a1752a,a1755a,a1758a,a1759a,a1760a,a1763a,a1766a,a1767a,a1770a,a1774a,a1775a,a1776a,a1777a,a1778a,a1781a,a1784a,a1785a,a1788a,a1792a,a1793a,a1794a,a1795a,a1798a,a1801a,a1802a,a1805a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1818a,a1821a,a1822a,a1825a,a1828a,a1829a,a1830a,a1833a,a1836a,a1837a,a1840a,a1844a,a1845a,a1846a,a1847a,a1848a,a1851a,a1854a,a1855a,a1858a,a1862a,a1863a,a1864a,a1865a,a1868a,a1871a,a1872a,a1875a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1887a,a1890a,a1891a,a1894a,a1897a,a1898a,a1899a,a1902a,a1905a,a1906a,a1909a,a1913a,a1914a,a1915a,a1916a,a1917a,a1920a,a1923a,a1924a,a1927a,a1931a,a1932a,a1933a,a1934a,a1937a,a1940a,a1941a,a1944a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1958a,a1961a,a1962a,a1965a,a1968a,a1969a,a1970a,a1973a,a1976a,a1977a,a1980a,a1984a,a1985a,a1986a,a1987a,a1988a,a1991a,a1994a,a1995a,a1998a,a2002a,a2003a,a2004a,a2005a,a2008a,a2011a,a2012a,a2015a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2027a,a2030a,a2031a,a2034a,a2037a,a2038a,a2039a,a2042a,a2045a,a2046a,a2049a,a2053a,a2054a,a2055a,a2056a,a2057a,a2060a,a2063a,a2064a,a2067a,a2071a,a2072a,a2073a,a2074a,a2077a,a2080a,a2081a,a2084a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2097a,a2100a,a2101a,a2104a,a2107a,a2108a,a2109a,a2112a,a2115a,a2116a,a2119a,a2123a,a2124a,a2125a,a2126a,a2127a,a2130a,a2133a,a2134a,a2137a,a2141a,a2142a,a2143a,a2144a,a2147a,a2150a,a2151a,a2154a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2166a,a2169a,a2170a,a2173a,a2176a,a2177a,a2178a,a2181a,a2184a,a2185a,a2188a,a2192a,a2193a,a2194a,a2195a,a2196a,a2199a,a2202a,a2203a,a2206a,a2210a,a2211a,a2212a,a2213a,a2216a,a2219a,a2220a,a2223a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2239a,a2242a,a2243a,a2246a,a2249a,a2250a,a2251a,a2254a,a2257a,a2258a,a2261a,a2265a,a2266a,a2267a,a2268a,a2269a,a2272a,a2275a,a2276a,a2279a,a2283a,a2284a,a2285a,a2286a,a2289a,a2292a,a2293a,a2296a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2308a,a2311a,a2312a,a2315a,a2318a,a2319a,a2320a,a2323a,a2326a,a2327a,a2330a,a2334a,a2335a,a2336a,a2337a,a2338a,a2341a,a2344a,a2345a,a2348a,a2352a,a2353a,a2354a,a2355a,a2358a,a2361a,a2362a,a2365a,a2369a,a2370a,a2371a,a2372a,a2373a,a2374a,a2375a,a2378a,a2381a,a2382a,a2385a,a2388a,a2389a,a2390a,a2393a,a2396a,a2397a,a2400a,a2404a,a2405a,a2406a,a2407a,a2408a,a2411a,a2414a,a2415a,a2418a,a2422a,a2423a,a2424a,a2425a,a2428a,a2431a,a2432a,a2435a,a2439a,a2440a,a2441a,a2442a,a2443a,a2444a,a2447a,a2450a,a2451a,a2454a,a2457a,a2458a,a2459a,a2462a,a2465a,a2466a,a2469a,a2473a,a2474a,a2475a,a2476a,a2477a,a2480a,a2483a,a2484a,a2487a,a2491a,a2492a,a2493a,a2494a,a2497a,a2500a,a2501a,a2504a,a2508a,a2509a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2518a,a2521a,a2522a,a2525a,a2528a,a2529a,a2530a,a2533a,a2536a,a2537a,a2540a,a2544a,a2545a,a2546a,a2547a,a2548a,a2551a,a2554a,a2555a,a2558a,a2562a,a2563a,a2564a,a2565a,a2568a,a2571a,a2572a,a2575a,a2579a,a2580a,a2581a,a2582a,a2583a,a2584a,a2587a,a2590a,a2591a,a2594a,a2597a,a2598a,a2599a,a2602a,a2605a,a2606a,a2609a,a2613a,a2614a,a2615a,a2616a,a2617a,a2620a,a2623a,a2624a,a2627a,a2631a,a2632a,a2633a,a2634a,a2637a,a2640a,a2641a,a2644a,a2648a,a2649a,a2650a,a2651a,a2652a,a2653a,a2654a,a2657a,a2660a,a2661a,a2664a,a2667a,a2668a,a2669a,a2672a,a2675a,a2676a,a2679a,a2683a,a2684a,a2685a,a2686a,a2687a,a2690a,a2693a,a2694a,a2697a,a2701a,a2702a,a2703a,a2704a,a2707a,a2710a,a2711a,a2714a,a2718a,a2719a,a2720a,a2721a,a2722a,a2723a,a2726a,a2729a,a2730a,a2733a,a2736a,a2737a,a2738a,a2741a,a2744a,a2745a,a2748a,a2752a,a2753a,a2754a,a2755a,a2756a,a2759a,a2762a,a2763a,a2766a,a2770a,a2771a,a2772a,a2773a,a2776a,a2779a,a2780a,a2783a,a2787a,a2788a,a2789a,a2790a,a2791a,a2792a,a2793a,a2794a,a2795a,a2798a,a2801a,a2802a,a2805a,a2808a,a2809a,a2810a,a2813a,a2816a,a2817a,a2820a,a2824a,a2825a,a2826a,a2827a,a2828a,a2831a,a2834a,a2835a,a2838a,a2842a,a2843a,a2844a,a2845a,a2848a,a2851a,a2852a,a2855a,a2859a,a2860a,a2861a,a2862a,a2863a,a2864a,a2867a,a2870a,a2871a,a2874a,a2877a,a2878a,a2879a,a2882a,a2885a,a2886a,a2889a,a2893a,a2894a,a2895a,a2896a,a2897a,a2900a,a2903a,a2904a,a2907a,a2911a,a2912a,a2913a,a2914a,a2917a,a2920a,a2921a,a2924a,a2928a,a2929a,a2930a,a2931a,a2932a,a2933a,a2934a,a2937a,a2940a,a2941a,a2944a,a2947a,a2948a,a2949a,a2952a,a2955a,a2956a,a2959a,a2963a,a2964a,a2965a,a2966a,a2967a,a2970a,a2973a,a2974a,a2977a,a2981a,a2982a,a2983a,a2984a,a2987a,a2990a,a2991a,a2994a,a2998a,a2999a,a3000a,a3001a,a3002a,a3003a,a3006a,a3009a,a3010a,a3013a,a3016a,a3017a,a3018a,a3021a,a3024a,a3025a,a3028a,a3032a,a3033a,a3034a,a3035a,a3036a,a3039a,a3042a,a3043a,a3046a,a3050a,a3051a,a3052a,a3053a,a3056a,a3059a,a3060a,a3063a,a3067a,a3068a,a3069a,a3070a,a3071a,a3072a,a3073a,a3074a,a3077a,a3080a,a3081a,a3084a,a3087a,a3088a,a3089a,a3092a,a3095a,a3096a,a3099a,a3103a,a3104a,a3105a,a3106a,a3107a,a3110a,a3113a,a3114a,a3117a,a3121a,a3122a,a3123a,a3124a,a3127a,a3130a,a3131a,a3134a,a3138a,a3139a,a3140a,a3141a,a3142a,a3143a,a3146a,a3149a,a3150a,a3153a,a3156a,a3157a,a3158a,a3161a,a3164a,a3165a,a3168a,a3172a,a3173a,a3174a,a3175a,a3176a,a3179a,a3182a,a3183a,a3186a,a3190a,a3191a,a3192a,a3193a,a3196a,a3199a,a3200a,a3203a,a3207a,a3208a,a3209a,a3210a,a3211a,a3212a,a3213a,a3216a,a3219a,a3220a,a3223a,a3226a,a3227a,a3228a,a3231a,a3234a,a3235a,a3238a,a3242a,a3243a,a3244a,a3245a,a3246a,a3249a,a3252a,a3253a,a3256a,a3260a,a3261a,a3262a,a3263a,a3266a,a3269a,a3270a,a3273a,a3277a,a3278a,a3279a,a3280a,a3281a,a3282a,a3285a,a3288a,a3289a,a3292a,a3295a,a3296a,a3297a,a3300a,a3303a,a3304a,a3307a,a3311a,a3312a,a3313a,a3314a,a3315a,a3318a,a3321a,a3322a,a3325a,a3329a,a3330a,a3331a,a3332a,a3335a,a3338a,a3339a,a3342a,a3346a,a3347a,a3348a,a3349a,a3350a,a3351a,a3352a,a3353a,a3354a,a3355a,a3358a,a3361a,a3364a,a3367a,a3370a,a3373a,a3377a,a3378a,a3382a,a3383a,a3387a,a3388a,a3392a,a3393a,a3397a,a3398a,a3402a,a3403a,a3407a,a3408a,a3412a,a3413a,a3417a,a3418a,a3422a,a3423a,a3427a,a3428a,a3432a,a3433a,a3437a,a3438a,a3442a,a3443a,a3447a,a3448a,a3452a,a3453a,a3457a,a3458a,a3462a,a3463a,a3467a,a3468a,a3472a,a3473a,a3477a,a3478a,a3482a,a3483a,a3487a,a3488a,a3492a,a3493a,a3496a,a3499a,a3500a,a3503a,a3506a,a3507a,a3510a,a3513a,a3514a,a3517a,a3520a,a3521a,a3524a,a3527a,a3528a,a3531a,a3534a,a3535a,a3538a,a3541a,a3542a,a3545a,a3548a,a3549a,a3552a,a3555a,a3556a,a3559a,a3562a,a3563a,a3566a,a3569a,a3570a,a3573a,a3576a,a3577a,a3580a,a3583a,a3584a,a3587a,a3590a,a3591a,a3594a,a3597a,a3598a,a3601a,a3604a,a3605a,a3608a,a3611a,a3612a,a3615a,a3618a,a3619a,a3622a,a3625a,a3626a,a3629a,a3632a,a3633a,a3636a,a3639a,a3640a,a3643a,a3646a,a3647a,a3650a,a3653a,a3654a,a3657a,a3660a,a3661a,a3664a,a3667a,a3668a,a3671a,a3674a,a3675a,a3678a,a3681a,a3682a,a3685a,a3688a,a3689a,a3692a,a3695a,a3696a,a3699a,a3702a,a3703a,a3706a,a3709a,a3710a,a3713a,a3716a,a3717a,a3720a,a3723a,a3724a,a3727a,a3730a,a3731a,a3734a,a3737a,a3738a,a3741a,a3744a,a3745a,a3748a,a3751a,a3752a,a3755a,a3758a,a3759a,a3762a,a3765a,a3766a,a3769a,a3772a,a3773a,a3776a,a3779a,a3780a,a3783a,a3786a,a3787a,a3790a,a3793a,a3794a,a3797a,a3800a,a3801a,a3804a,a3807a,a3808a,a3811a,a3814a,a3815a,a3818a,a3821a,a3822a,a3825a,a3828a,a3829a,a3832a,a3835a,a3836a,a3839a,a3842a,a3843a,a3846a,a3849a,a3850a,a3853a,a3856a,a3857a,a3860a,a3863a,a3864a,a3867a,a3870a,a3871a,a3874a,a3877a,a3878a,a3881a,a3884a,a3885a,a3888a,a3891a,a3892a,a3895a,a3898a,a3899a,a3902a,a3905a,a3906a,a3909a,a3912a,a3913a,a3916a,a3919a,a3920a,a3923a,a3926a,a3927a,a3930a,a3933a,a3934a,a3937a,a3940a,a3941a,a3944a,a3947a,a3948a,a3951a,a3954a,a3955a,a3958a,a3961a,a3962a,a3965a,a3968a,a3969a,a3972a,a3975a,a3976a,a3979a,a3982a,a3983a,a3986a,a3989a,a3990a,a3993a,a3996a,a3997a,a4000a,a4003a,a4004a,a4007a,a4011a,a4012a,a4013a,a4016a,a4019a,a4020a,a4023a,a4027a,a4028a,a4029a,a4032a,a4035a,a4036a,a4039a,a4043a,a4044a,a4045a,a4048a,a4051a,a4052a,a4055a,a4059a,a4060a,a4061a,a4064a,a4067a,a4068a,a4071a,a4075a,a4076a,a4077a,a4080a,a4083a,a4084a,a4087a,a4091a,a4092a,a4093a,a4096a,a4099a,a4100a,a4103a,a4107a,a4108a,a4109a,a4112a,a4115a,a4116a,a4119a,a4123a,a4124a,a4125a,a4128a,a4131a,a4132a,a4135a,a4139a,a4140a,a4141a,a4144a,a4147a,a4148a,a4151a,a4155a,a4156a,a4157a,a4160a,a4163a,a4164a,a4167a,a4171a,a4172a,a4173a,a4176a,a4179a,a4180a,a4183a,a4187a,a4188a,a4189a,a4192a,a4195a,a4196a,a4199a,a4203a,a4204a,a4205a,a4208a,a4211a,a4212a,a4215a,a4219a,a4220a,a4221a,a4224a,a4227a,a4228a,a4231a,a4235a,a4236a,a4237a,a4240a,a4243a,a4244a,a4247a,a4251a,a4252a,a4253a,a4256a,a4259a,a4260a,a4263a,a4267a,a4268a,a4269a,a4272a,a4275a,a4276a,a4279a,a4283a,a4284a,a4285a,a4288a,a4291a,a4292a,a4295a,a4299a,a4300a,a4301a,a4304a,a4307a,a4308a,a4311a,a4315a,a4316a,a4317a,a4320a,a4323a,a4324a,a4327a,a4331a,a4332a,a4333a,a4336a,a4339a,a4340a,a4343a,a4347a,a4348a,a4349a,a4352a,a4355a,a4356a,a4359a,a4363a,a4364a,a4365a,a4368a,a4371a,a4372a,a4375a,a4379a,a4380a,a4381a,a4384a,a4387a,a4388a,a4391a,a4395a,a4396a,a4397a,a4400a,a4403a,a4404a,a4407a,a4411a,a4412a,a4413a,a4416a,a4419a,a4420a,a4423a,a4427a,a4428a,a4429a,a4432a,a4435a,a4436a,a4439a,a4443a,a4444a,a4445a,a4448a,a4451a,a4452a,a4455a,a4459a,a4460a,a4461a,a4464a,a4467a,a4468a,a4471a,a4475a,a4476a,a4477a,a4480a,a4483a,a4484a,a4487a,a4491a,a4492a,a4493a,a4496a,a4499a,a4500a,a4503a,a4507a,a4508a,a4509a,a4512a,a4515a,a4516a,a4519a,a4523a,a4524a,a4525a,a4528a,a4531a,a4532a,a4535a,a4539a,a4540a,a4541a,a4544a,a4547a,a4548a,a4551a,a4555a,a4556a,a4557a,a4560a,a4563a,a4564a,a4567a,a4571a,a4572a,a4573a,a4576a,a4579a,a4580a,a4583a,a4587a,a4588a,a4589a,a4592a,a4595a,a4596a,a4599a,a4603a,a4604a,a4605a,a4608a,a4611a,a4612a,a4615a,a4619a,a4620a,a4621a,a4624a,a4627a,a4628a,a4631a,a4635a,a4636a,a4637a,a4640a,a4643a,a4644a,a4647a,a4651a,a4652a,a4653a,a4656a,a4659a,a4660a,a4663a,a4667a,a4668a,a4669a,a4672a,a4675a,a4676a,a4679a,a4683a,a4684a,a4685a,a4688a,a4691a,a4692a,a4695a,a4699a,a4700a,a4701a,a4704a,a4707a,a4708a,a4711a,a4715a,a4716a,a4717a,a4720a,a4723a,a4724a,a4727a,a4731a,a4732a,a4733a,a4736a,a4739a,a4740a,a4743a,a4747a,a4748a,a4749a,a4752a,a4755a,a4756a,a4759a,a4763a,a4764a,a4765a,a4768a,a4771a,a4772a,a4775a,a4779a,a4780a,a4781a,a4784a,a4787a,a4788a,a4791a,a4795a,a4796a,a4797a,a4800a,a4803a,a4804a,a4807a,a4811a,a4812a,a4813a,a4816a,a4819a,a4820a,a4823a,a4827a,a4828a,a4829a,a4832a,a4835a,a4836a,a4839a,a4843a,a4844a,a4845a,a4848a,a4851a,a4852a,a4855a,a4859a,a4860a,a4861a,a4864a,a4867a,a4868a,a4871a,a4875a,a4876a,a4877a,a4880a,a4883a,a4884a,a4887a,a4891a,a4892a,a4893a,a4896a,a4899a,a4900a,a4903a,a4907a,a4908a,a4909a,a4912a,a4915a,a4916a,a4919a,a4923a,a4924a,a4925a,a4928a,a4931a,a4932a,a4935a,a4939a,a4940a,a4941a,a4944a,a4947a,a4948a,a4951a,a4955a,a4956a,a4957a,a4960a,a4963a,a4964a,a4967a,a4971a,a4972a,a4973a,a4976a,a4979a,a4980a,a4983a,a4987a,a4988a,a4989a,a4992a,a4996a,a4997a,a4998a,a5001a,a5005a,a5006a,a5007a,a5010a,a5014a,a5015a,a5016a,a5019a,a5023a,a5024a,a5025a,a5028a,a5032a,a5033a,a5034a,a5037a,a5041a,a5042a,a5043a,a5046a,a5050a,a5051a,a5052a,a5055a,a5059a,a5060a,a5061a,a5064a,a5068a,a5069a,a5070a,a5073a,a5077a,a5078a,a5079a,a5082a,a5086a,a5087a,a5088a,a5091a,a5095a,a5096a,a5097a,a5100a,a5104a,a5105a,a5106a,a5109a,a5113a,a5114a,a5115a,a5118a,a5122a,a5123a,a5124a,a5127a,a5131a,a5132a,a5133a,a5136a,a5140a,a5141a,a5142a,a5145a,a5149a,a5150a,a5151a,a5154a,a5158a,a5159a,a5160a,a5163a,a5167a,a5168a,a5169a,a5172a,a5176a,a5177a,a5178a,a5181a,a5185a,a5186a,a5187a,a5190a,a5194a,a5195a,a5196a,a5199a,a5203a,a5204a,a5205a,a5208a,a5212a,a5213a,a5214a,a5217a,a5221a,a5222a,a5223a,a5226a,a5230a,a5231a,a5232a,a5235a,a5239a,a5240a,a5241a,a5244a,a5248a,a5249a,a5250a,a5253a,a5257a,a5258a,a5259a,a5262a,a5266a,a5267a,a5268a,a5271a,a5275a,a5276a,a5277a,a5280a,a5284a,a5285a,a5286a,a5289a,a5293a,a5294a,a5295a,a5298a,a5302a,a5303a,a5304a,a5307a,a5311a,a5312a,a5313a,a5316a,a5320a,a5321a,a5322a,a5325a,a5329a,a5330a,a5331a,a5334a,a5338a,a5339a,a5340a,a5343a,a5347a,a5348a,a5349a,a5352a,a5356a,a5357a,a5358a,a5361a,a5365a,a5366a,a5367a,a5370a,a5374a,a5375a,a5376a,a5379a,a5383a,a5384a,a5385a,a5388a,a5392a,a5393a,a5394a,a5397a,a5401a,a5402a,a5403a,a5406a,a5410a,a5411a,a5412a,a5415a,a5419a,a5420a,a5421a,a5424a,a5428a,a5429a,a5430a,a5433a,a5437a,a5438a,a5439a,a5442a,a5446a,a5447a,a5448a,a5451a,a5455a,a5456a,a5457a,a5460a,a5464a,a5465a,a5466a,a5469a,a5473a,a5474a,a5475a,a5478a,a5482a,a5483a,a5484a,a5487a,a5491a,a5492a,a5493a,a5496a,a5500a,a5501a,a5502a,a5505a,a5509a,a5510a,a5511a,a5514a,a5518a,a5519a,a5520a,a5523a,a5527a,a5528a,a5529a,a5532a,a5536a,a5537a,a5538a,a5541a,a5545a,a5546a,a5547a,a5550a,a5554a,a5555a,a5556a,a5559a,a5563a,a5564a,a5565a,a5568a,a5572a,a5573a,a5574a,a5577a,a5581a,a5582a,a5583a,a5586a,a5590a,a5591a,a5592a,a5595a,a5599a,a5600a,a5601a,a5604a,a5608a,a5609a,a5610a,a5613a,a5617a,a5618a,a5619a,a5622a,a5626a,a5627a,a5628a,a5631a,a5635a,a5636a,a5637a,a5640a,a5644a,a5645a,a5646a,a5649a,a5653a,a5654a,a5655a,a5658a,a5662a,a5663a,a5664a,a5667a,a5671a,a5672a,a5673a,a5676a,a5680a,a5681a,a5682a,a5685a,a5689a,a5690a,a5691a,a5694a,a5698a,a5699a,a5700a,a5703a,a5707a,a5708a,a5709a,a5712a,a5716a,a5717a,a5718a,a5721a,a5725a,a5726a,a5727a,a5730a,a5734a,a5735a,a5736a,a5739a,a5743a,a5744a,a5745a,a5748a,a5752a,a5753a,a5754a,a5757a,a5761a,a5762a,a5763a,a5766a,a5770a,a5771a,a5772a,a5775a,a5779a,a5780a,a5781a,a5784a,a5788a,a5789a,a5790a,a5793a,a5797a,a5798a,a5799a,a5802a,a5806a,a5807a,a5808a,a5811a,a5815a,a5816a,a5817a,a5820a,a5824a,a5825a,a5826a,a5829a,a5833a,a5834a,a5835a,a5838a,a5842a,a5843a,a5844a,a5847a,a5851a,a5852a,a5853a,a5856a,a5860a,a5861a,a5862a,a5865a,a5869a,a5870a,a5871a,a5874a,a5878a,a5879a,a5880a,a5883a,a5887a,a5888a,a5889a,a5892a,a5896a,a5897a,a5898a,a5901a,a5905a,a5906a,a5907a,a5910a,a5914a,a5915a,a5916a,a5919a,a5923a,a5924a,a5925a,a5928a,a5932a,a5933a,a5934a,a5937a,a5941a,a5942a,a5943a,a5946a,a5950a,a5951a,a5952a,a5955a,a5959a,a5960a,a5961a,a5964a,a5968a,a5969a,a5970a,a5973a,a5977a,a5978a,a5979a,a5982a,a5986a,a5987a,a5988a,a5991a,a5995a,a5996a,a5997a,a6000a,a6004a,a6005a,a6006a,a6009a,a6013a,a6014a,a6015a,a6018a,a6022a,a6023a,a6024a,a6027a,a6031a,a6032a,a6033a,a6036a,a6040a,a6041a,a6042a,a6045a,a6049a,a6050a,a6051a,a6054a,a6058a,a6059a,a6060a,a6063a,a6067a,a6068a,a6069a,a6072a,a6076a,a6077a,a6078a,a6081a,a6085a,a6086a,a6087a,a6090a,a6094a,a6095a,a6096a,a6099a,a6103a,a6104a,a6105a,a6108a,a6112a,a6113a,a6114a,a6117a,a6121a,a6122a,a6123a,a6126a,a6130a,a6131a,a6132a,a6135a,a6139a,a6140a,a6141a,a6144a,a6148a,a6149a,a6150a,a6153a,a6157a,a6158a,a6159a,a6162a,a6166a,a6167a,a6168a,a6171a,a6175a,a6176a,a6177a,a6180a,a6184a,a6185a,a6186a,a6189a,a6193a,a6194a,a6195a,a6198a,a6202a,a6203a,a6204a,a6207a,a6211a,a6212a,a6213a,a6216a,a6220a,a6221a,a6222a,a6225a,a6229a,a6230a,a6231a,a6234a,a6238a,a6239a,a6240a,a6243a,a6247a,a6248a,a6249a,a6252a,a6256a,a6257a,a6258a,a6261a,a6265a,a6266a,a6267a,a6270a,a6274a,a6275a,a6276a,a6279a,a6283a,a6284a,a6285a,a6288a,a6292a,a6293a,a6294a,a6297a,a6301a,a6302a,a6303a,a6306a,a6310a,a6311a,a6312a,a6315a,a6319a,a6320a,a6321a,a6324a,a6328a,a6329a,a6330a,a6333a,a6337a,a6338a,a6339a,a6342a,a6346a,a6347a,a6348a,a6351a,a6355a,a6356a,a6357a,a6360a,a6364a,a6365a,a6366a,a6369a,a6373a,a6374a,a6375a,a6378a,a6382a,a6383a,a6384a,a6387a,a6391a,a6392a,a6393a,a6396a,a6400a,a6401a,a6402a,a6405a,a6409a,a6410a,a6411a,a6414a,a6418a,a6419a,a6420a,a6423a,a6427a,a6428a,a6429a,a6432a,a6436a,a6437a,a6438a,a6441a,a6445a,a6446a,a6447a,a6450a,a6454a,a6455a,a6456a,a6459a,a6463a,a6464a,a6465a,a6468a,a6472a,a6473a,a6474a,a6477a,a6481a,a6482a,a6483a,a6486a,a6490a,a6491a,a6492a,a6495a,a6499a,a6500a,a6501a,a6504a,a6508a,a6509a,a6510a,a6513a,a6517a,a6518a,a6519a,a6522a,a6526a,a6527a,a6528a,a6531a,a6535a,a6536a,a6537a,a6540a,a6544a,a6545a,a6546a,a6549a,a6553a,a6554a,a6555a,a6558a,a6562a,a6563a,a6564a,a6567a,a6571a,a6572a,a6573a,a6576a,a6580a,a6581a,a6582a,a6585a,a6589a,a6590a,a6591a,a6594a,a6598a,a6599a,a6600a,a6603a,a6607a,a6608a,a6609a,a6612a,a6616a,a6617a,a6618a,a6621a,a6625a,a6626a,a6627a,a6630a,a6634a,a6635a,a6636a,a6639a,a6643a,a6644a,a6645a,a6648a,a6652a,a6653a,a6654a,a6657a,a6661a,a6662a,a6663a,a6666a,a6670a,a6671a,a6672a,a6675a,a6679a,a6680a,a6681a,a6684a,a6688a,a6689a,a6690a,a6693a,a6697a,a6698a,a6699a,a6702a,a6706a,a6707a,a6708a,a6711a,a6715a,a6716a,a6717a,a6720a,a6724a,a6725a,a6726a,a6729a,a6733a,a6734a,a6735a,a6738a,a6742a,a6743a,a6744a,a6747a,a6751a,a6752a,a6753a,a6756a,a6760a,a6761a,a6762a,a6765a,a6769a,a6770a,a6771a,a6774a,a6778a,a6779a,a6780a,a6783a,a6787a,a6788a,a6789a,a6792a,a6796a,a6797a,a6798a,a6801a,a6805a,a6806a,a6807a,a6810a,a6814a,a6815a,a6816a,a6819a,a6823a,a6824a,a6825a,a6828a,a6832a,a6833a,a6834a,a6837a,a6841a,a6842a,a6843a,a6846a,a6850a,a6851a,a6852a,a6855a,a6859a,a6860a,a6861a,a6864a,a6868a,a6869a,a6870a,a6873a,a6877a,a6878a,a6879a,a6882a,a6886a,a6887a,a6888a,a6891a,a6895a,a6896a,a6897a,a6900a,a6904a,a6905a,a6906a,a6909a,a6913a,a6914a,a6915a,a6918a,a6922a,a6923a,a6924a,a6927a,a6931a,a6932a,a6933a,a6936a,a6940a,a6941a,a6942a,a6945a,a6949a,a6950a,a6951a,a6954a,a6958a,a6959a,a6960a,a6963a,a6967a,a6968a,a6969a,a6972a,a6976a,a6977a,a6978a,a6981a,a6985a,a6986a,a6987a,a6990a,a6994a,a6995a,a6996a,a6999a,a7003a,a7004a,a7005a,a7008a,a7012a,a7013a,a7014a,a7017a,a7021a,a7022a,a7023a,a7026a,a7030a,a7031a,a7032a,a7035a,a7039a,a7040a,a7041a,a7044a,a7048a,a7049a,a7050a,a7053a,a7057a,a7058a,a7059a,a7062a,a7066a,a7067a,a7068a,a7071a,a7075a,a7076a,a7077a,a7080a,a7084a,a7085a,a7086a,a7089a,a7093a,a7094a,a7095a,a7098a,a7102a,a7103a,a7104a,a7107a,a7111a,a7112a,a7113a,a7116a,a7120a,a7121a,a7122a,a7125a,a7129a,a7130a,a7131a,a7134a,a7138a,a7139a,a7140a,a7143a,a7147a,a7148a,a7149a,a7152a,a7156a,a7157a,a7158a,a7161a,a7165a,a7166a,a7167a,a7170a,a7174a,a7175a,a7176a,a7179a,a7183a,a7184a,a7185a,a7188a,a7192a,a7193a,a7194a,a7197a,a7201a,a7202a,a7203a,a7206a,a7210a,a7211a,a7212a,a7215a,a7219a,a7220a,a7221a,a7224a,a7228a,a7229a,a7230a,a7233a,a7237a,a7238a,a7239a,a7242a,a7246a,a7247a,a7248a,a7251a,a7255a,a7256a,a7257a,a7260a,a7264a,a7265a,a7266a,a7269a,a7273a,a7274a,a7275a,a7278a,a7282a,a7283a,a7284a,a7287a,a7291a,a7292a,a7293a,a7296a,a7300a,a7301a,a7302a,a7305a,a7309a,a7310a,a7311a,a7314a,a7318a,a7319a,a7320a,a7323a,a7327a,a7328a,a7329a,a7332a,a7336a,a7337a,a7338a,a7341a,a7345a,a7346a,a7347a,a7350a,a7354a,a7355a,a7356a,a7359a,a7363a,a7364a,a7365a,a7368a,a7372a,a7373a,a7374a,a7377a,a7381a,a7382a,a7383a,a7386a,a7390a,a7391a,a7392a,a7395a,a7399a,a7400a,a7401a,a7404a,a7408a,a7409a,a7410a,a7413a,a7417a,a7418a,a7419a,a7422a,a7426a,a7427a,a7428a,a7431a,a7435a,a7436a,a7437a,a7440a,a7444a,a7445a,a7446a,a7449a,a7453a,a7454a,a7455a,a7458a,a7462a,a7463a,a7464a,a7467a,a7471a,a7472a,a7473a,a7476a,a7480a,a7481a,a7482a,a7485a,a7489a,a7490a,a7491a,a7494a,a7498a,a7499a,a7500a,a7503a,a7507a,a7508a,a7509a,a7512a,a7516a,a7517a,a7518a,a7521a,a7525a,a7526a,a7527a,a7530a,a7534a,a7535a,a7536a,a7539a,a7543a,a7544a,a7545a,a7548a,a7552a,a7553a,a7554a,a7557a,a7561a,a7562a,a7563a,a7566a,a7570a,a7571a,a7572a,a7575a,a7579a,a7580a,a7581a,a7584a,a7588a,a7589a,a7590a,a7593a,a7597a,a7598a,a7599a,a7602a,a7606a,a7607a,a7608a,a7611a,a7615a,a7616a,a7617a,a7620a,a7624a,a7625a,a7626a,a7629a,a7633a,a7634a,a7635a,a7638a,a7642a,a7643a,a7644a,a7647a,a7651a,a7652a,a7653a,a7656a,a7660a,a7661a,a7662a,a7665a,a7669a,a7670a,a7671a,a7674a,a7678a,a7679a,a7680a,a7683a,a7687a,a7688a,a7689a,a7692a,a7696a,a7697a,a7698a,a7701a,a7705a,a7706a,a7707a,a7710a,a7714a,a7715a,a7716a,a7719a,a7723a,a7724a,a7725a,a7728a,a7732a,a7733a,a7734a,a7737a,a7741a,a7742a,a7743a,a7746a,a7750a,a7751a,a7752a,a7755a,a7759a,a7760a,a7761a,a7764a,a7768a,a7769a,a7770a,a7773a,a7777a,a7778a,a7779a,a7782a,a7786a,a7787a,a7788a,a7791a,a7795a,a7796a,a7797a,a7800a,a7804a,a7805a,a7806a,a7809a,a7813a,a7814a,a7815a,a7818a,a7822a,a7823a,a7824a,a7827a,a7831a,a7832a,a7833a,a7836a,a7840a,a7841a,a7842a,a7845a,a7849a,a7850a,a7851a,a7854a,a7858a,a7859a,a7860a,a7863a,a7867a,a7868a,a7869a,a7872a,a7876a,a7877a,a7878a,a7881a,a7885a,a7886a,a7887a,a7890a,a7894a,a7895a,a7896a,a7899a,a7903a,a7904a,a7905a,a7908a,a7912a,a7913a,a7914a,a7917a,a7921a,a7922a,a7923a,a7926a,a7930a,a7931a,a7932a,a7935a,a7939a,a7940a,a7941a,a7944a,a7948a,a7949a,a7950a,a7953a,a7957a,a7958a,a7959a,a7962a,a7966a,a7967a,a7968a,a7971a,a7975a,a7976a,a7977a,a7980a,a7984a,a7985a,a7986a,a7989a,a7993a,a7994a,a7995a,a7998a,a8002a,a8003a,a8004a,a8007a,a8011a,a8012a,a8013a,a8016a,a8020a,a8021a,a8022a,a8025a,a8029a,a8030a,a8031a,a8034a,a8038a,a8039a,a8040a,a8043a,a8047a,a8048a,a8049a,a8052a,a8056a,a8057a,a8058a,a8061a,a8065a,a8066a,a8067a,a8070a,a8074a,a8075a,a8076a,a8079a,a8083a,a8084a,a8085a,a8088a,a8092a,a8093a,a8094a,a8097a,a8101a,a8102a,a8103a,a8106a,a8110a,a8111a,a8112a,a8115a,a8119a,a8120a,a8121a,a8124a,a8128a,a8129a,a8130a,a8134a,a8135a,a8139a,a8140a,a8141a,a8144a,a8148a,a8149a,a8150a,a8154a,a8155a,a8159a,a8160a,a8161a,a8164a,a8168a,a8169a,a8170a,a8174a,a8175a,a8179a,a8180a,a8181a,a8184a,a8188a,a8189a,a8190a,a8194a,a8195a,a8199a,a8200a,a8201a,a8204a,a8208a,a8209a,a8210a,a8214a,a8215a,a8219a,a8220a,a8221a,a8224a,a8228a,a8229a,a8230a,a8234a,a8235a,a8239a,a8240a,a8241a,a8244a,a8248a,a8249a,a8250a,a8254a,a8255a,a8259a,a8260a,a8261a,a8264a,a8268a,a8269a,a8270a,a8274a,a8275a,a8279a,a8280a,a8281a,a8284a,a8288a,a8289a,a8290a,a8294a,a8295a,a8299a,a8300a,a8301a,a8304a,a8308a,a8309a,a8310a,a8314a,a8315a,a8319a,a8320a,a8321a,a8324a,a8328a,a8329a,a8330a,a8334a,a8335a,a8339a,a8340a,a8341a,a8344a,a8348a,a8349a,a8350a,a8354a,a8355a,a8359a,a8360a,a8361a,a8364a,a8368a,a8369a,a8370a,a8374a,a8375a,a8379a,a8380a,a8381a,a8384a,a8388a,a8389a,a8390a,a8394a,a8395a,a8399a,a8400a,a8401a,a8404a,a8408a,a8409a,a8410a,a8414a,a8415a,a8419a,a8420a,a8421a,a8424a,a8428a,a8429a,a8430a,a8434a,a8435a,a8439a,a8440a,a8441a,a8444a,a8448a,a8449a,a8450a,a8454a,a8455a,a8459a,a8460a,a8461a,a8464a,a8468a,a8469a,a8470a,a8474a,a8475a,a8479a,a8480a,a8481a,a8484a,a8488a,a8489a,a8490a,a8494a,a8495a,a8499a,a8500a,a8501a,a8504a,a8508a,a8509a,a8510a,a8514a,a8515a,a8519a,a8520a,a8521a,a8524a,a8528a,a8529a,a8530a,a8534a,a8535a,a8539a,a8540a,a8541a,a8544a,a8548a,a8549a,a8550a,a8554a,a8555a,a8559a,a8560a,a8561a,a8564a,a8568a,a8569a,a8570a,a8574a,a8575a,a8579a,a8580a,a8581a,a8584a,a8588a,a8589a,a8590a,a8594a,a8595a,a8599a,a8600a,a8601a,a8604a,a8608a,a8609a,a8610a,a8614a,a8615a,a8619a,a8620a,a8621a,a8624a,a8628a,a8629a,a8630a,a8634a,a8635a,a8639a,a8640a,a8641a,a8644a,a8648a,a8649a,a8650a,a8654a,a8655a,a8659a,a8660a,a8661a,a8664a,a8668a,a8669a,a8670a,a8674a,a8675a,a8679a,a8680a,a8681a,a8684a,a8688a,a8689a,a8690a,a8694a,a8695a,a8699a,a8700a,a8701a,a8704a,a8708a,a8709a,a8710a,a8714a,a8715a,a8719a,a8720a,a8721a,a8724a,a8728a,a8729a,a8730a,a8734a,a8735a,a8739a,a8740a,a8741a,a8744a,a8748a,a8749a,a8750a,a8754a,a8755a,a8759a,a8760a,a8761a,a8764a,a8768a,a8769a,a8770a,a8774a,a8775a,a8779a,a8780a,a8781a,a8784a,a8788a,a8789a,a8790a,a8794a,a8795a,a8799a,a8800a,a8801a,a8804a,a8808a,a8809a,a8810a,a8814a,a8815a,a8819a,a8820a,a8821a,a8824a,a8828a,a8829a,a8830a,a8834a,a8835a,a8839a,a8840a,a8841a,a8844a,a8848a,a8849a,a8850a,a8854a,a8855a,a8859a,a8860a,a8861a,a8864a,a8868a,a8869a,a8870a,a8874a,a8875a,a8879a,a8880a,a8881a,a8884a,a8888a,a8889a,a8890a,a8894a,a8895a,a8899a,a8900a,a8901a,a8904a,a8908a,a8909a,a8910a,a8914a,a8915a,a8919a,a8920a,a8921a,a8924a,a8928a,a8929a,a8930a,a8934a,a8935a,a8939a,a8940a,a8941a,a8944a,a8948a,a8949a,a8950a,a8954a,a8955a,a8959a,a8960a,a8961a,a8964a,a8968a,a8969a,a8970a,a8974a,a8975a,a8979a,a8980a,a8981a,a8984a,a8988a,a8989a,a8990a,a8994a,a8995a,a8999a,a9000a,a9001a,a9004a,a9008a,a9009a,a9010a,a9014a,a9015a,a9019a,a9020a,a9021a,a9024a,a9028a,a9029a,a9030a,a9034a,a9035a,a9039a,a9040a,a9041a,a9044a,a9048a,a9049a,a9050a,a9054a,a9055a,a9059a,a9060a,a9061a,a9064a,a9068a,a9069a,a9070a,a9074a,a9075a,a9079a,a9080a,a9081a,a9084a,a9088a,a9089a,a9090a,a9094a,a9095a,a9099a,a9100a,a9101a,a9104a,a9108a,a9109a,a9110a,a9114a,a9115a,a9119a,a9120a,a9121a,a9124a,a9128a,a9129a,a9130a,a9134a,a9135a,a9139a,a9140a,a9141a,a9144a,a9148a,a9149a,a9150a,a9154a,a9155a,a9159a,a9160a,a9161a,a9164a,a9168a,a9169a,a9170a,a9174a,a9175a,a9179a,a9180a,a9181a,a9184a,a9188a,a9189a,a9190a,a9194a,a9195a,a9199a,a9200a,a9201a,a9204a,a9208a,a9209a,a9210a,a9214a,a9215a,a9219a,a9220a,a9221a,a9224a,a9228a,a9229a,a9230a,a9234a,a9235a,a9239a,a9240a,a9241a,a9244a,a9248a,a9249a,a9250a,a9254a,a9255a,a9259a,a9260a,a9261a,a9264a,a9268a,a9269a,a9270a,a9274a,a9275a,a9279a,a9280a,a9281a,a9284a,a9288a,a9289a,a9290a,a9294a,a9295a,a9299a,a9300a,a9301a,a9304a,a9308a,a9309a,a9310a,a9314a,a9315a,a9319a,a9320a,a9321a,a9324a,a9328a,a9329a,a9330a,a9334a,a9335a,a9339a,a9340a,a9341a,a9344a,a9348a,a9349a,a9350a,a9354a,a9355a,a9359a,a9360a,a9361a,a9364a,a9368a,a9369a,a9370a,a9374a,a9375a,a9379a,a9380a,a9381a,a9384a,a9388a,a9389a,a9390a,a9394a,a9395a,a9399a,a9400a,a9401a,a9404a,a9408a,a9409a,a9410a,a9414a,a9415a,a9419a,a9420a,a9421a,a9424a,a9428a,a9429a,a9430a,a9434a,a9435a,a9439a,a9440a,a9441a,a9444a,a9448a,a9449a,a9450a,a9454a,a9455a,a9459a,a9460a,a9461a,a9464a,a9468a,a9469a,a9470a,a9474a,a9475a,a9479a,a9480a,a9481a,a9484a,a9488a,a9489a,a9490a,a9494a,a9495a,a9499a,a9500a,a9501a,a9504a,a9508a,a9509a,a9510a,a9514a,a9515a,a9519a,a9520a,a9521a,a9524a,a9528a,a9529a,a9530a,a9534a,a9535a,a9539a,a9540a,a9541a,a9544a,a9548a,a9549a,a9550a,a9554a,a9555a,a9559a,a9560a,a9561a,a9564a,a9568a,a9569a,a9570a,a9574a,a9575a,a9579a,a9580a,a9581a,a9584a,a9588a,a9589a,a9590a,a9594a,a9595a,a9599a,a9600a,a9601a,a9604a,a9608a,a9609a,a9610a,a9614a,a9615a,a9619a,a9620a,a9621a,a9624a,a9628a,a9629a,a9630a,a9634a,a9635a,a9639a,a9640a,a9641a,a9644a,a9648a,a9649a,a9650a,a9654a,a9655a,a9659a,a9660a,a9661a,a9664a,a9668a,a9669a,a9670a,a9674a,a9675a,a9679a,a9680a,a9681a,a9684a,a9688a,a9689a,a9690a,a9694a,a9695a,a9699a,a9700a,a9701a,a9704a,a9708a,a9709a,a9710a,a9714a,a9715a,a9719a,a9720a,a9721a,a9724a,a9728a,a9729a,a9730a,a9734a,a9735a,a9739a,a9740a,a9741a,a9744a,a9748a,a9749a,a9750a,a9754a,a9755a,a9759a,a9760a,a9761a,a9764a,a9768a,a9769a,a9770a,a9774a,a9775a,a9779a,a9780a,a9781a,a9784a,a9788a,a9789a,a9790a,a9794a,a9795a,a9799a,a9800a,a9801a,a9804a,a9808a,a9809a,a9810a,a9814a,a9815a,a9819a,a9820a,a9821a,a9824a,a9828a,a9829a,a9830a,a9834a,a9835a,a9839a,a9840a,a9841a,a9844a,a9848a,a9849a,a9850a,a9854a,a9855a,a9859a,a9860a,a9861a,a9864a,a9868a,a9869a,a9870a,a9874a,a9875a,a9879a,a9880a,a9881a,a9884a,a9888a,a9889a,a9890a,a9894a,a9895a,a9899a,a9900a,a9901a,a9904a,a9908a,a9909a,a9910a,a9914a,a9915a,a9919a,a9920a,a9921a,a9924a,a9928a,a9929a,a9930a,a9934a,a9935a,a9939a,a9940a,a9941a,a9944a,a9948a,a9949a,a9950a,a9954a,a9955a,a9959a,a9960a,a9961a,a9964a,a9968a,a9969a,a9970a,a9974a,a9975a,a9979a,a9980a,a9981a,a9984a,a9988a,a9989a,a9990a,a9994a,a9995a,a9999a,a10000a,a10001a,a10004a,a10008a,a10009a,a10010a,a10014a,a10015a,a10019a,a10020a,a10021a,a10024a,a10028a,a10029a,a10030a,a10034a,a10035a,a10039a,a10040a,a10041a,a10044a,a10048a,a10049a,a10050a,a10054a,a10055a,a10059a,a10060a,a10061a,a10064a,a10068a,a10069a,a10070a,a10074a,a10075a,a10079a,a10080a,a10081a,a10084a,a10088a,a10089a,a10090a,a10094a,a10095a,a10099a,a10100a,a10101a,a10104a,a10108a,a10109a,a10110a,a10114a,a10115a,a10119a,a10120a,a10121a,a10124a,a10128a,a10129a,a10130a,a10134a,a10135a,a10139a,a10140a,a10141a,a10144a,a10148a,a10149a,a10150a,a10154a,a10155a,a10159a,a10160a,a10161a,a10164a,a10168a,a10169a,a10170a,a10174a,a10175a,a10179a,a10180a,a10181a,a10184a,a10188a,a10189a,a10190a,a10194a,a10195a,a10199a,a10200a,a10201a,a10204a,a10208a,a10209a,a10210a,a10214a,a10215a,a10219a,a10220a,a10221a,a10224a,a10228a,a10229a,a10230a,a10234a,a10235a,a10239a,a10240a,a10241a,a10244a,a10248a,a10249a,a10250a,a10254a,a10255a,a10259a,a10260a,a10261a,a10264a,a10268a,a10269a,a10270a,a10274a,a10275a,a10279a,a10280a,a10281a,a10284a,a10288a,a10289a,a10290a,a10294a,a10295a,a10299a,a10300a,a10301a,a10304a,a10308a,a10309a,a10310a,a10314a,a10315a,a10319a,a10320a,a10321a,a10324a,a10328a,a10329a,a10330a,a10334a,a10335a,a10339a,a10340a,a10341a,a10344a,a10348a,a10349a,a10350a,a10354a,a10355a,a10359a,a10360a,a10361a,a10364a,a10368a,a10369a,a10370a,a10374a,a10375a,a10379a,a10380a,a10381a,a10384a,a10388a,a10389a,a10390a,a10394a,a10395a,a10399a,a10400a,a10401a,a10404a,a10408a,a10409a,a10410a,a10414a,a10415a,a10419a,a10420a,a10421a,a10424a,a10428a,a10429a,a10430a,a10434a,a10435a,a10439a,a10440a,a10441a,a10444a,a10448a,a10449a,a10450a,a10454a,a10455a,a10459a,a10460a,a10461a,a10464a,a10468a,a10469a,a10470a,a10474a,a10475a,a10479a,a10480a,a10481a,a10484a,a10488a,a10489a,a10490a,a10494a,a10495a,a10499a,a10500a,a10501a,a10504a,a10508a,a10509a,a10510a,a10514a,a10515a,a10519a,a10520a,a10521a,a10524a,a10528a,a10529a,a10530a,a10534a,a10535a,a10539a,a10540a,a10541a,a10544a,a10548a,a10549a,a10550a,a10554a,a10555a,a10559a,a10560a,a10561a,a10564a,a10568a,a10569a,a10570a,a10574a,a10575a,a10579a,a10580a,a10581a,a10584a,a10588a,a10589a,a10590a,a10594a,a10595a,a10599a,a10600a,a10601a,a10604a,a10608a,a10609a,a10610a,a10614a,a10615a,a10619a,a10620a,a10621a,a10624a,a10628a,a10629a,a10630a,a10634a,a10635a,a10639a,a10640a,a10641a,a10644a,a10648a,a10649a,a10650a,a10654a,a10655a,a10659a,a10660a,a10661a,a10664a,a10668a,a10669a,a10670a,a10674a,a10675a,a10679a,a10680a,a10681a,a10684a,a10688a,a10689a,a10690a,a10694a,a10695a,a10699a,a10700a,a10701a,a10704a,a10708a,a10709a,a10710a,a10714a,a10715a,a10719a,a10720a,a10721a,a10724a,a10728a,a10729a,a10730a,a10734a,a10735a,a10739a,a10740a,a10741a,a10744a,a10748a,a10749a,a10750a,a10754a,a10755a,a10759a,a10760a,a10761a,a10764a,a10768a,a10769a,a10770a,a10774a,a10775a,a10779a,a10780a,a10781a,a10784a,a10788a,a10789a,a10790a,a10794a,a10795a,a10799a,a10800a,a10801a,a10804a,a10808a,a10809a,a10810a,a10814a,a10815a,a10819a,a10820a,a10821a,a10824a,a10828a,a10829a,a10830a,a10834a,a10835a,a10839a,a10840a,a10841a,a10844a,a10848a,a10849a,a10850a,a10854a,a10855a,a10859a,a10860a,a10861a,a10864a,a10868a,a10869a,a10870a,a10874a,a10875a,a10879a,a10880a,a10881a,a10884a,a10888a,a10889a,a10890a,a10894a,a10895a,a10899a,a10900a,a10901a,a10904a,a10908a,a10909a,a10910a,a10914a,a10915a,a10919a,a10920a,a10921a,a10924a,a10928a,a10929a,a10930a,a10934a,a10935a,a10939a,a10940a,a10941a,a10944a,a10948a,a10949a,a10950a,a10954a,a10955a,a10959a,a10960a,a10961a,a10964a,a10968a,a10969a,a10970a,a10974a,a10975a,a10979a,a10980a,a10981a,a10984a,a10988a,a10989a,a10990a,a10994a,a10995a,a10999a,a11000a,a11001a,a11004a,a11008a,a11009a,a11010a,a11014a,a11015a,a11019a,a11020a,a11021a,a11024a,a11028a,a11029a,a11030a,a11034a,a11035a,a11039a,a11040a,a11041a,a11044a,a11048a,a11049a,a11050a,a11054a,a11055a,a11059a,a11060a,a11061a,a11064a,a11068a,a11069a,a11070a,a11074a,a11075a,a11079a,a11080a,a11081a,a11084a,a11088a,a11089a,a11090a,a11094a,a11095a,a11099a,a11100a,a11101a,a11104a,a11108a,a11109a,a11110a,a11114a,a11115a,a11119a,a11120a,a11121a,a11124a,a11128a,a11129a,a11130a,a11134a,a11135a,a11139a,a11140a,a11141a,a11144a,a11148a,a11149a,a11150a,a11154a,a11155a,a11159a,a11160a,a11161a,a11164a,a11168a,a11169a,a11170a,a11174a,a11175a,a11179a,a11180a,a11181a,a11184a,a11188a,a11189a,a11190a,a11194a,a11195a,a11199a,a11200a,a11201a,a11204a,a11208a,a11209a,a11210a,a11214a,a11215a,a11219a,a11220a,a11221a,a11224a,a11228a,a11229a,a11230a,a11234a,a11235a,a11239a,a11240a,a11241a,a11244a,a11248a,a11249a,a11250a,a11254a,a11255a,a11259a,a11260a,a11261a,a11264a,a11268a,a11269a,a11270a,a11274a,a11275a,a11279a,a11280a,a11281a,a11284a,a11288a,a11289a,a11290a,a11294a,a11295a,a11299a,a11300a,a11301a,a11304a,a11308a,a11309a,a11310a,a11314a,a11315a,a11319a,a11320a,a11321a,a11324a,a11328a,a11329a,a11330a,a11334a,a11335a,a11339a,a11340a,a11341a,a11344a,a11348a,a11349a,a11350a,a11354a,a11355a,a11359a,a11360a,a11361a,a11364a,a11368a,a11369a,a11370a,a11374a,a11375a,a11379a,a11380a,a11381a,a11384a,a11388a,a11389a,a11390a,a11394a,a11395a,a11399a,a11400a,a11401a,a11404a,a11408a,a11409a,a11410a,a11414a,a11415a,a11419a,a11420a,a11421a,a11424a,a11428a,a11429a,a11430a,a11434a,a11435a,a11439a,a11440a,a11441a,a11444a,a11448a,a11449a,a11450a,a11454a,a11455a,a11459a,a11460a,a11461a,a11464a,a11468a,a11469a,a11470a,a11474a,a11475a,a11479a,a11480a,a11481a,a11484a,a11488a,a11489a,a11490a,a11494a,a11495a,a11499a,a11500a,a11501a,a11504a,a11508a,a11509a,a11510a,a11514a,a11515a,a11519a,a11520a,a11521a,a11524a,a11528a,a11529a,a11530a,a11534a,a11535a,a11539a,a11540a,a11541a,a11544a,a11548a,a11549a,a11550a,a11554a,a11555a,a11559a,a11560a,a11561a,a11564a,a11568a,a11569a,a11570a,a11574a,a11575a,a11579a,a11580a,a11581a,a11584a,a11588a,a11589a,a11590a,a11594a,a11595a,a11599a,a11600a,a11601a,a11604a,a11608a,a11609a,a11610a,a11614a,a11615a,a11619a,a11620a,a11621a,a11624a,a11628a,a11629a,a11630a,a11634a,a11635a,a11639a,a11640a,a11641a,a11644a,a11648a,a11649a,a11650a,a11654a,a11655a,a11659a,a11660a,a11661a,a11664a,a11668a,a11669a,a11670a,a11674a,a11675a,a11679a,a11680a,a11681a,a11684a,a11688a,a11689a,a11690a,a11694a,a11695a,a11699a,a11700a,a11701a,a11704a,a11708a,a11709a,a11710a,a11714a,a11715a,a11719a,a11720a,a11721a,a11724a,a11728a,a11729a,a11730a,a11734a,a11735a,a11739a,a11740a,a11741a,a11744a,a11748a,a11749a,a11750a,a11754a,a11755a,a11759a,a11760a,a11761a,a11764a,a11768a,a11769a,a11770a,a11774a,a11775a,a11779a,a11780a,a11781a,a11784a,a11788a,a11789a,a11790a,a11794a,a11795a,a11799a,a11800a,a11801a,a11804a,a11808a,a11809a,a11810a,a11814a,a11815a,a11819a,a11820a,a11821a,a11824a,a11828a,a11829a,a11830a,a11834a,a11835a,a11839a,a11840a,a11841a,a11844a,a11848a,a11849a,a11850a,a11854a,a11855a,a11859a,a11860a,a11861a,a11864a,a11868a,a11869a,a11870a,a11874a,a11875a,a11879a,a11880a,a11881a,a11884a,a11888a,a11889a,a11890a,a11894a,a11895a,a11899a,a11900a,a11901a,a11904a,a11908a,a11909a,a11910a,a11914a,a11915a,a11919a,a11920a,a11921a,a11924a,a11928a,a11929a,a11930a,a11934a,a11935a,a11939a,a11940a,a11941a,a11944a,a11948a,a11949a,a11950a,a11954a,a11955a,a11959a,a11960a,a11961a,a11964a,a11968a,a11969a,a11970a,a11974a,a11975a,a11979a,a11980a,a11981a,a11984a,a11988a,a11989a,a11990a,a11994a,a11995a,a11999a,a12000a,a12001a,a12004a,a12008a,a12009a,a12010a,a12014a,a12015a,a12019a,a12020a,a12021a,a12024a,a12028a,a12029a,a12030a,a12034a,a12035a,a12039a,a12040a,a12041a,a12044a,a12048a,a12049a,a12050a,a12054a,a12055a,a12059a,a12060a,a12061a,a12064a,a12068a,a12069a,a12070a,a12074a,a12075a,a12079a,a12080a,a12081a,a12084a,a12088a,a12089a,a12090a,a12094a,a12095a,a12099a,a12100a,a12101a,a12104a,a12108a,a12109a,a12110a,a12114a,a12115a,a12119a,a12120a,a12121a,a12124a,a12128a,a12129a,a12130a,a12134a,a12135a,a12139a,a12140a,a12141a,a12144a,a12148a,a12149a,a12150a,a12154a,a12155a,a12159a,a12160a,a12161a,a12164a,a12168a,a12169a,a12170a,a12174a,a12175a,a12179a,a12180a,a12181a,a12184a,a12188a,a12189a,a12190a,a12194a,a12195a,a12199a,a12200a,a12201a,a12204a,a12208a,a12209a,a12210a,a12214a,a12215a,a12219a,a12220a,a12221a,a12225a,a12226a,a12230a,a12231a,a12232a,a12236a,a12237a,a12241a,a12242a,a12243a,a12247a,a12248a,a12252a,a12253a,a12254a,a12258a,a12259a,a12263a,a12264a,a12265a,a12269a,a12270a,a12274a,a12275a,a12276a,a12280a,a12281a,a12285a,a12286a,a12287a,a12291a,a12292a,a12296a,a12297a,a12298a,a12302a,a12303a,a12307a,a12308a,a12309a,a12313a,a12314a,a12318a,a12319a,a12320a,a12324a,a12325a,a12329a,a12330a,a12331a,a12335a,a12336a,a12340a,a12341a,a12342a,a12346a,a12347a,a12351a,a12352a,a12353a,a12357a,a12358a,a12362a,a12363a,a12364a,a12368a,a12369a,a12373a,a12374a,a12375a,a12379a,a12380a,a12384a,a12385a,a12386a,a12390a,a12391a,a12395a,a12396a,a12397a,a12401a,a12402a,a12406a,a12407a,a12408a,a12412a,a12413a,a12417a,a12418a,a12419a,a12423a,a12424a,a12428a,a12429a,a12430a,a12434a,a12435a,a12439a,a12440a,a12441a,a12445a,a12446a,a12450a,a12451a,a12452a,a12456a,a12457a,a12461a,a12462a,a12463a,a12467a,a12468a,a12472a,a12473a,a12474a,a12478a,a12479a,a12483a,a12484a,a12485a,a12489a,a12490a,a12494a,a12495a,a12496a,a12500a,a12501a,a12505a,a12506a,a12507a,a12511a,a12512a,a12516a,a12517a,a12518a,a12522a,a12523a,a12527a,a12528a,a12529a,a12533a,a12534a,a12538a,a12539a,a12540a,a12544a,a12545a,a12549a,a12550a,a12551a,a12555a,a12556a,a12560a,a12561a,a12562a,a12566a,a12567a,a12571a,a12572a,a12573a,a12577a,a12578a,a12582a,a12583a,a12584a,a12588a,a12589a,a12593a,a12594a,a12595a,a12599a,a12600a,a12604a,a12605a,a12606a,a12610a,a12611a,a12615a,a12616a,a12617a,a12621a,a12622a,a12626a,a12627a,a12628a,a12632a,a12633a,a12637a,a12638a,a12639a,a12643a,a12644a,a12648a,a12649a,a12650a,a12654a,a12655a,a12659a,a12660a,a12661a,a12665a,a12666a,a12670a,a12671a,a12672a,a12676a,a12677a,a12681a,a12682a,a12683a,a12687a,a12688a,a12692a,a12693a,a12694a,a12698a,a12699a,a12703a,a12704a,a12705a,a12709a,a12710a,a12714a,a12715a,a12716a,a12720a,a12721a,a12725a,a12726a,a12727a,a12731a,a12732a,a12736a,a12737a,a12738a,a12742a,a12743a,a12747a,a12748a,a12749a,a12753a,a12754a,a12758a,a12759a,a12760a,a12764a,a12765a,a12769a,a12770a,a12771a,a12775a,a12776a,a12780a,a12781a,a12782a,a12786a,a12787a,a12791a,a12792a,a12793a,a12797a,a12798a,a12802a,a12803a,a12804a,a12808a,a12809a,a12813a,a12814a,a12815a,a12819a,a12820a,a12824a,a12825a,a12826a,a12830a,a12831a,a12835a,a12836a,a12837a,a12841a,a12842a,a12846a,a12847a,a12848a,a12852a,a12853a,a12857a,a12858a,a12859a,a12863a,a12864a,a12868a,a12869a,a12870a,a12874a,a12875a,a12879a,a12880a,a12881a,a12885a,a12886a,a12890a,a12891a,a12892a,a12896a,a12897a,a12901a,a12902a,a12903a,a12907a,a12908a,a12912a,a12913a,a12914a,a12918a,a12919a,a12923a,a12924a,a12925a,a12929a,a12930a,a12934a,a12935a,a12936a,a12940a,a12941a,a12945a,a12946a,a12947a,a12951a,a12952a,a12956a,a12957a,a12958a,a12962a,a12963a,a12967a,a12968a,a12969a,a12973a,a12974a,a12978a,a12979a,a12980a,a12984a,a12985a,a12989a,a12990a,a12991a,a12995a,a12996a,a13000a,a13001a,a13002a,a13006a,a13007a,a13011a,a13012a,a13013a,a13017a,a13018a,a13022a,a13023a,a13024a,a13028a,a13029a,a13033a,a13034a,a13035a,a13039a,a13040a,a13044a,a13045a,a13046a,a13050a,a13051a,a13055a,a13056a,a13057a,a13061a,a13062a,a13066a,a13067a,a13068a,a13072a,a13073a,a13077a,a13078a,a13079a,a13083a,a13084a,a13088a,a13089a,a13090a,a13094a,a13095a,a13099a,a13100a,a13101a,a13105a,a13106a,a13110a,a13111a,a13112a,a13116a,a13117a,a13121a,a13122a,a13123a,a13127a,a13128a,a13132a,a13133a,a13134a,a13138a,a13139a,a13143a,a13144a,a13145a,a13149a,a13150a,a13154a,a13155a,a13156a,a13160a,a13161a,a13165a,a13166a,a13167a,a13171a,a13172a,a13176a,a13177a,a13178a,a13182a,a13183a,a13187a,a13188a,a13189a,a13193a,a13194a,a13198a,a13199a,a13200a,a13204a,a13205a,a13209a,a13210a,a13211a,a13215a,a13216a,a13220a,a13221a,a13222a,a13226a,a13227a,a13231a,a13232a,a13233a,a13237a,a13238a,a13242a,a13243a,a13244a,a13248a,a13249a,a13253a,a13254a,a13255a,a13259a,a13260a,a13264a,a13265a,a13266a,a13270a,a13271a,a13275a,a13276a,a13277a,a13281a,a13282a,a13286a,a13287a,a13288a,a13292a,a13293a,a13297a,a13298a,a13299a,a13303a,a13304a,a13308a,a13309a,a13310a,a13314a,a13315a,a13319a,a13320a,a13321a,a13325a,a13326a,a13330a,a13331a,a13332a,a13336a,a13337a,a13341a,a13342a,a13343a,a13347a,a13348a,a13352a,a13353a,a13354a,a13358a,a13359a,a13363a,a13364a,a13365a,a13369a,a13370a,a13374a,a13375a,a13376a,a13380a,a13381a,a13385a,a13386a,a13387a,a13391a,a13392a,a13396a,a13397a,a13398a,a13402a,a13403a,a13407a,a13408a,a13409a,a13413a,a13414a,a13418a,a13419a,a13420a,a13424a,a13425a,a13429a,a13430a,a13431a,a13435a,a13436a,a13440a,a13441a,a13442a,a13446a,a13447a,a13451a,a13452a,a13453a,a13457a,a13458a,a13462a,a13463a,a13464a,a13468a,a13469a,a13473a,a13474a,a13475a,a13479a,a13480a,a13484a,a13485a,a13486a,a13490a,a13491a,a13495a,a13496a,a13497a,a13501a,a13502a,a13506a,a13507a,a13508a,a13512a,a13513a,a13517a,a13518a,a13519a,a13523a,a13524a,a13528a,a13529a,a13530a,a13534a,a13535a,a13539a,a13540a,a13541a,a13545a,a13546a,a13550a,a13551a,a13552a,a13556a,a13557a,a13561a,a13562a,a13563a,a13567a,a13568a,a13572a,a13573a,a13574a,a13578a,a13579a,a13583a,a13584a,a13585a,a13589a,a13590a,a13594a,a13595a,a13596a,a13600a,a13601a,a13605a,a13606a,a13607a,a13611a,a13612a,a13616a,a13617a,a13618a,a13622a,a13623a,a13627a,a13628a,a13629a,a13633a,a13634a,a13638a,a13639a,a13640a,a13644a,a13645a,a13649a,a13650a,a13651a,a13655a,a13656a,a13660a,a13661a,a13662a,a13666a,a13667a,a13671a,a13672a,a13673a,a13677a,a13678a,a13682a,a13683a,a13684a,a13688a,a13689a,a13693a,a13694a,a13695a,a13699a,a13700a,a13704a,a13705a,a13706a,a13710a,a13711a,a13715a,a13716a,a13717a,a13721a,a13722a,a13726a,a13727a,a13728a,a13732a,a13733a,a13737a,a13738a,a13739a,a13743a,a13744a,a13748a,a13749a,a13750a,a13754a,a13755a,a13759a,a13760a,a13761a,a13765a,a13766a,a13770a,a13771a,a13772a,a13776a,a13777a,a13781a,a13782a,a13783a,a13787a,a13788a,a13792a,a13793a,a13794a,a13798a,a13799a,a13803a,a13804a,a13805a,a13809a,a13810a,a13814a,a13815a,a13816a,a13820a,a13821a,a13825a,a13826a,a13827a,a13831a,a13832a,a13836a,a13837a,a13838a,a13842a,a13843a,a13847a,a13848a,a13849a,a13853a,a13854a,a13858a,a13859a,a13860a,a13864a,a13865a,a13869a,a13870a,a13871a,a13875a,a13876a,a13880a,a13881a,a13882a,a13886a,a13887a,a13891a,a13892a,a13893a,a13897a,a13898a,a13902a,a13903a,a13904a,a13908a,a13909a,a13913a,a13914a,a13915a,a13919a,a13920a,a13924a,a13925a,a13926a,a13930a,a13931a,a13935a,a13936a,a13937a,a13941a,a13942a,a13946a,a13947a,a13948a,a13952a,a13953a,a13957a,a13958a,a13959a,a13963a,a13964a,a13968a,a13969a,a13970a,a13974a,a13975a,a13979a,a13980a,a13981a,a13985a,a13986a,a13990a,a13991a,a13992a,a13996a,a13997a,a14001a,a14002a,a14003a,a14007a,a14008a,a14012a,a14013a,a14014a,a14018a,a14019a,a14023a,a14024a,a14025a,a14029a,a14030a,a14034a,a14035a,a14036a,a14040a,a14041a,a14045a,a14046a,a14047a,a14051a,a14052a,a14056a,a14057a,a14058a,a14062a,a14063a,a14067a,a14068a,a14069a,a14073a,a14074a,a14078a,a14079a,a14080a,a14084a,a14085a,a14089a,a14090a,a14091a,a14095a,a14096a,a14100a,a14101a,a14102a,a14106a,a14107a,a14111a,a14112a,a14113a,a14117a,a14118a,a14122a,a14123a,a14124a,a14128a,a14129a,a14133a,a14134a,a14135a,a14139a,a14140a,a14144a,a14145a,a14146a,a14150a,a14151a,a14155a,a14156a,a14157a,a14161a,a14162a,a14166a,a14167a,a14168a,a14172a,a14173a,a14177a,a14178a,a14179a,a14183a,a14184a,a14188a,a14189a,a14190a,a14194a,a14195a,a14199a,a14200a,a14201a,a14205a,a14206a,a14210a,a14211a,a14212a,a14216a,a14217a,a14221a,a14222a,a14223a,a14227a,a14228a,a14232a,a14233a,a14234a,a14238a,a14239a,a14243a,a14244a,a14245a,a14249a,a14250a,a14254a,a14255a,a14256a,a14260a,a14261a,a14265a,a14266a,a14267a,a14271a,a14272a,a14276a,a14277a,a14278a,a14282a,a14283a,a14287a,a14288a,a14289a,a14293a,a14294a,a14298a,a14299a,a14300a,a14304a,a14305a,a14309a,a14310a,a14311a,a14315a,a14316a,a14320a,a14321a,a14322a,a14326a,a14327a,a14331a,a14332a,a14333a,a14337a,a14338a,a14342a,a14343a,a14344a,a14348a,a14349a,a14353a,a14354a,a14355a,a14359a,a14360a,a14364a,a14365a,a14366a,a14370a,a14371a,a14375a,a14376a,a14377a,a14381a,a14382a,a14386a,a14387a,a14388a,a14392a,a14393a,a14397a,a14398a,a14399a,a14403a,a14404a,a14408a,a14409a,a14410a,a14414a,a14415a,a14419a,a14420a,a14421a,a14425a,a14426a,a14430a,a14431a,a14432a,a14436a,a14437a,a14441a,a14442a,a14443a,a14447a,a14448a,a14452a,a14453a,a14454a,a14458a,a14459a,a14463a,a14464a,a14465a,a14469a,a14470a,a14474a,a14475a,a14476a,a14480a,a14481a,a14485a,a14486a,a14487a,a14491a,a14492a,a14496a,a14497a,a14498a,a14502a,a14503a,a14507a,a14508a,a14509a,a14513a,a14514a,a14518a,a14519a,a14520a,a14524a,a14525a,a14529a,a14530a,a14531a,a14535a,a14536a,a14540a,a14541a,a14542a,a14546a,a14547a,a14551a,a14552a,a14553a,a14557a,a14558a,a14562a,a14563a,a14564a,a14568a,a14569a,a14573a,a14574a,a14575a,a14579a,a14580a,a14584a,a14585a,a14586a,a14590a,a14591a,a14595a,a14596a,a14597a,a14601a,a14602a,a14606a,a14607a,a14608a,a14612a,a14613a,a14617a,a14618a,a14619a,a14623a,a14624a,a14628a,a14629a,a14630a,a14634a,a14635a,a14639a,a14640a,a14641a,a14645a,a14646a,a14650a,a14651a,a14652a,a14656a,a14657a,a14661a,a14662a,a14663a,a14667a,a14668a,a14672a,a14673a,a14674a,a14678a,a14679a,a14683a,a14684a,a14685a,a14689a,a14690a,a14694a,a14695a,a14696a,a14700a,a14701a,a14705a,a14706a,a14707a,a14711a,a14712a,a14716a,a14717a,a14718a,a14722a,a14723a,a14727a,a14728a,a14729a,a14733a,a14734a,a14738a,a14739a,a14740a,a14744a,a14745a,a14749a,a14750a,a14751a,a14755a,a14756a,a14760a,a14761a,a14762a,a14766a,a14767a,a14771a,a14772a,a14773a,a14777a,a14778a,a14782a,a14783a,a14784a,a14788a,a14789a,a14793a,a14794a,a14795a,a14799a,a14800a,a14804a,a14805a,a14806a,a14810a,a14811a,a14815a,a14816a,a14817a,a14821a,a14822a,a14826a,a14827a,a14828a,a14832a,a14833a,a14837a,a14838a,a14839a,a14843a,a14844a,a14848a,a14849a,a14850a,a14854a,a14855a,a14859a,a14860a,a14861a,a14865a,a14866a,a14870a,a14871a,a14872a,a14876a,a14877a,a14881a,a14882a,a14883a,a14887a,a14888a,a14892a,a14893a,a14894a,a14898a,a14899a,a14903a,a14904a,a14905a,a14909a,a14910a,a14914a,a14915a,a14916a,a14920a,a14921a,a14925a,a14926a,a14927a,a14931a,a14932a,a14936a,a14937a,a14938a,a14942a,a14943a,a14947a,a14948a,a14949a,a14953a,a14954a,a14958a,a14959a,a14960a,a14964a,a14965a,a14969a,a14970a,a14971a,a14975a,a14976a,a14980a,a14981a,a14982a,a14986a,a14987a,a14991a,a14992a,a14993a,a14997a,a14998a,a15002a,a15003a,a15004a,a15008a,a15009a,a15013a,a15014a,a15015a,a15019a,a15020a,a15024a,a15025a,a15026a,a15030a,a15031a,a15035a,a15036a,a15037a,a15041a,a15042a,a15046a,a15047a,a15048a,a15052a,a15053a,a15057a,a15058a,a15059a,a15063a,a15064a,a15068a,a15069a,a15070a,a15074a,a15075a,a15079a,a15080a,a15081a,a15085a,a15086a,a15090a,a15091a,a15092a,a15096a,a15097a,a15101a,a15102a,a15103a,a15107a,a15108a,a15112a,a15113a,a15114a,a15118a,a15119a,a15123a,a15124a,a15125a,a15129a,a15130a,a15134a,a15135a,a15136a,a15140a,a15141a,a15145a,a15146a,a15147a,a15151a,a15152a,a15156a,a15157a,a15158a,a15162a,a15163a,a15167a,a15168a,a15169a,a15173a,a15174a,a15178a,a15179a,a15180a,a15184a,a15185a,a15189a,a15190a,a15191a,a15195a,a15196a,a15200a,a15201a,a15202a,a15206a,a15207a,a15211a,a15212a,a15213a,a15217a,a15218a,a15222a,a15223a,a15224a,a15228a,a15229a,a15233a,a15234a,a15235a,a15239a,a15240a,a15244a,a15245a,a15246a,a15250a,a15251a,a15255a,a15256a,a15257a,a15261a,a15262a,a15266a,a15267a,a15268a,a15272a,a15273a,a15277a,a15278a,a15279a,a15283a,a15284a,a15288a,a15289a,a15290a,a15294a,a15295a,a15299a,a15300a,a15301a,a15305a,a15306a,a15310a,a15311a,a15312a,a15316a,a15317a,a15321a,a15322a,a15323a,a15327a,a15328a,a15332a,a15333a,a15334a,a15338a,a15339a,a15343a,a15344a,a15345a,a15349a,a15350a,a15354a,a15355a,a15356a,a15360a,a15361a,a15365a,a15366a,a15367a,a15371a,a15372a,a15376a,a15377a,a15378a,a15382a,a15383a,a15387a,a15388a,a15389a,a15393a,a15394a,a15398a,a15399a,a15400a,a15404a,a15405a,a15409a,a15410a,a15411a,a15415a,a15416a,a15420a,a15421a,a15422a,a15426a,a15427a,a15431a,a15432a,a15433a,a15437a,a15438a,a15442a,a15443a,a15444a,a15448a,a15449a,a15453a,a15454a,a15455a,a15459a,a15460a,a15464a,a15465a,a15466a,a15470a,a15471a,a15475a,a15476a,a15477a,a15481a,a15482a,a15486a,a15487a,a15488a,a15492a,a15493a,a15497a,a15498a,a15499a,a15503a,a15504a,a15508a,a15509a,a15510a,a15514a,a15515a,a15519a,a15520a,a15521a,a15525a,a15526a,a15530a,a15531a,a15532a,a15536a,a15537a,a15541a,a15542a,a15543a,a15547a,a15548a,a15552a,a15553a,a15554a,a15558a,a15559a,a15563a,a15564a,a15565a,a15569a,a15570a,a15574a,a15575a,a15576a,a15580a,a15581a,a15585a,a15586a,a15587a,a15591a,a15592a,a15596a,a15597a,a15598a,a15602a,a15603a,a15607a,a15608a,a15609a,a15613a,a15614a,a15618a,a15619a,a15620a,a15624a,a15625a,a15629a,a15630a,a15631a,a15635a,a15636a,a15640a,a15641a,a15642a,a15646a,a15647a,a15651a,a15652a,a15653a,a15657a,a15658a,a15662a,a15663a,a15664a,a15668a,a15669a,a15673a,a15674a,a15675a,a15679a,a15680a,a15684a,a15685a,a15686a,a15690a,a15691a,a15695a,a15696a,a15697a,a15701a,a15702a,a15706a,a15707a,a15708a,a15712a,a15713a,a15717a,a15718a,a15719a,a15723a,a15724a,a15728a,a15729a,a15730a,a15734a,a15735a,a15739a,a15740a,a15741a,a15745a,a15746a,a15750a,a15751a,a15752a,a15756a,a15757a,a15761a,a15762a,a15763a,a15767a,a15768a,a15772a,a15773a,a15774a,a15778a,a15779a,a15783a,a15784a,a15785a,a15789a,a15790a,a15794a,a15795a,a15796a,a15800a,a15801a,a15805a,a15806a,a15807a,a15811a,a15812a,a15816a,a15817a,a15818a,a15822a,a15823a,a15827a,a15828a,a15829a,a15833a,a15834a,a15838a,a15839a,a15840a,a15844a,a15845a,a15849a,a15850a,a15851a,a15855a,a15856a,a15860a,a15861a,a15862a,a15866a,a15867a,a15871a,a15872a,a15873a,a15877a,a15878a,a15882a,a15883a,a15884a,a15888a,a15889a,a15893a,a15894a,a15895a,a15899a,a15900a,a15904a,a15905a,a15906a,a15910a,a15911a,a15915a,a15916a,a15917a,a15921a,a15922a,a15926a,a15927a,a15928a,a15932a,a15933a,a15937a,a15938a,a15939a,a15943a,a15944a,a15948a,a15949a,a15950a,a15954a,a15955a,a15959a,a15960a,a15961a,a15965a,a15966a,a15970a,a15971a,a15972a,a15976a,a15977a,a15981a,a15982a,a15983a,a15987a,a15988a,a15992a,a15993a,a15994a,a15998a,a15999a,a16003a,a16004a,a16005a,a16009a,a16010a,a16014a,a16015a,a16016a,a16020a,a16021a,a16025a,a16026a,a16027a,a16031a,a16032a,a16036a,a16037a,a16038a,a16042a,a16043a,a16047a,a16048a,a16049a,a16053a,a16054a,a16058a,a16059a,a16060a,a16064a,a16065a,a16069a,a16070a,a16071a,a16075a,a16076a,a16080a,a16081a,a16082a,a16086a,a16087a,a16091a,a16092a,a16093a,a16097a,a16098a,a16102a,a16103a,a16104a,a16108a,a16109a,a16113a,a16114a,a16115a,a16119a,a16120a,a16124a,a16125a,a16126a,a16130a,a16131a,a16135a,a16136a,a16137a,a16141a,a16142a,a16146a,a16147a,a16148a,a16152a,a16153a,a16157a,a16158a,a16159a,a16163a,a16164a,a16168a,a16169a,a16170a,a16174a,a16175a,a16179a,a16180a,a16181a,a16185a,a16186a,a16190a,a16191a,a16192a,a16196a,a16197a,a16201a,a16202a,a16203a,a16207a,a16208a,a16212a,a16213a,a16214a,a16218a,a16219a,a16223a,a16224a,a16225a,a16229a,a16230a,a16234a,a16235a,a16236a,a16240a,a16241a,a16245a,a16246a,a16247a,a16251a,a16252a,a16256a,a16257a,a16258a,a16262a,a16263a,a16267a,a16268a,a16269a,a16273a,a16274a,a16278a,a16279a,a16280a,a16284a,a16285a,a16289a,a16290a,a16291a,a16295a,a16296a,a16300a,a16301a,a16302a,a16306a,a16307a,a16311a,a16312a,a16313a,a16317a,a16318a,a16322a,a16323a,a16324a,a16328a,a16329a,a16333a,a16334a,a16335a,a16339a,a16340a,a16344a,a16345a,a16346a,a16350a,a16351a,a16355a,a16356a,a16357a,a16361a,a16362a,a16366a,a16367a,a16368a,a16372a,a16373a,a16377a,a16378a,a16379a,a16383a,a16384a,a16388a,a16389a,a16390a,a16394a,a16395a,a16399a,a16400a,a16401a,a16405a,a16406a,a16410a,a16411a,a16412a,a16416a,a16417a,a16421a,a16422a,a16423a,a16427a,a16428a,a16432a,a16433a,a16434a,a16438a,a16439a,a16443a,a16444a,a16445a,a16449a,a16450a,a16454a,a16455a,a16456a,a16460a,a16461a,a16465a,a16466a,a16467a,a16471a,a16472a,a16476a,a16477a,a16478a,a16482a,a16483a,a16487a,a16488a,a16489a,a16493a,a16494a,a16498a,a16499a,a16500a,a16504a,a16505a,a16509a,a16510a,a16511a,a16515a,a16516a,a16520a,a16521a,a16522a,a16526a,a16527a,a16531a,a16532a,a16533a,a16537a,a16538a,a16542a,a16543a,a16544a,a16548a,a16549a,a16553a,a16554a,a16555a,a16559a,a16560a,a16564a,a16565a,a16566a,a16570a,a16571a,a16575a,a16576a,a16577a,a16581a,a16582a,a16586a,a16587a,a16588a,a16592a,a16593a,a16597a,a16598a,a16599a,a16603a,a16604a,a16608a,a16609a,a16610a,a16614a,a16615a,a16619a,a16620a,a16621a,a16625a,a16626a,a16630a,a16631a,a16632a,a16636a,a16637a,a16641a,a16642a,a16643a,a16647a,a16648a,a16652a,a16653a,a16654a,a16658a,a16659a,a16663a,a16664a,a16665a,a16669a,a16670a,a16674a,a16675a,a16676a,a16680a,a16681a,a16685a,a16686a,a16687a,a16691a,a16692a,a16696a,a16697a,a16698a,a16702a,a16703a,a16707a,a16708a,a16709a,a16713a,a16714a,a16718a,a16719a,a16720a,a16724a,a16725a,a16729a,a16730a,a16731a,a16735a,a16736a,a16740a,a16741a,a16742a,a16746a,a16747a,a16751a,a16752a,a16753a,a16757a,a16758a,a16762a,a16763a,a16764a,a16768a,a16769a,a16773a,a16774a,a16775a,a16779a,a16780a,a16784a,a16785a,a16786a,a16790a,a16791a,a16795a,a16796a,a16797a,a16801a,a16802a,a16806a,a16807a,a16808a,a16812a,a16813a,a16817a,a16818a,a16819a,a16823a,a16824a,a16828a,a16829a,a16830a,a16834a,a16835a,a16839a,a16840a,a16841a,a16845a,a16846a,a16850a,a16851a,a16852a,a16856a,a16857a,a16861a,a16862a,a16863a,a16867a,a16868a,a16872a,a16873a,a16874a,a16878a,a16879a,a16883a,a16884a,a16885a,a16889a,a16890a,a16894a,a16895a,a16896a,a16900a,a16901a,a16905a,a16906a,a16907a,a16911a,a16912a,a16916a,a16917a,a16918a,a16922a,a16923a,a16927a,a16928a,a16929a,a16933a,a16934a,a16938a,a16939a,a16940a,a16944a,a16945a,a16949a,a16950a,a16951a,a16955a,a16956a,a16960a,a16961a,a16962a,a16966a,a16967a,a16971a,a16972a,a16973a,a16977a,a16978a,a16982a,a16983a,a16984a,a16988a,a16989a,a16993a,a16994a,a16995a,a16999a,a17000a,a17004a,a17005a,a17006a,a17010a,a17011a,a17015a,a17016a,a17017a,a17021a,a17022a,a17026a,a17027a,a17028a,a17032a,a17033a,a17037a,a17038a,a17039a,a17043a,a17044a,a17048a,a17049a,a17050a,a17054a,a17055a,a17059a,a17060a,a17061a,a17065a,a17066a,a17070a,a17071a,a17072a,a17076a,a17077a,a17081a,a17082a,a17083a,a17087a,a17088a,a17092a,a17093a,a17094a,a17098a,a17099a,a17103a,a17104a,a17105a,a17109a,a17110a,a17114a,a17115a,a17116a,a17120a,a17121a,a17125a,a17126a,a17127a,a17131a,a17132a,a17136a,a17137a,a17138a,a17142a,a17143a,a17147a,a17148a,a17149a,a17153a,a17154a,a17158a,a17159a,a17160a,a17164a,a17165a,a17169a,a17170a,a17171a,a17175a,a17176a,a17180a,a17181a,a17182a,a17186a,a17187a,a17191a,a17192a,a17193a,a17197a,a17198a,a17202a,a17203a,a17204a,a17208a,a17209a,a17213a,a17214a,a17215a,a17219a,a17220a,a17224a,a17225a,a17226a,a17230a,a17231a,a17235a,a17236a,a17237a,a17241a,a17242a,a17246a,a17247a,a17248a,a17252a,a17253a,a17257a,a17258a,a17259a,a17263a,a17264a,a17268a,a17269a,a17270a,a17274a,a17275a,a17279a,a17280a,a17281a,a17285a,a17286a,a17290a,a17291a,a17292a,a17296a,a17297a,a17301a,a17302a,a17303a,a17307a,a17308a,a17312a,a17313a,a17314a,a17318a,a17319a,a17323a,a17324a,a17325a,a17329a,a17330a,a17334a,a17335a,a17336a,a17340a,a17341a,a17345a,a17346a,a17347a,a17351a,a17352a,a17356a,a17357a,a17358a,a17362a,a17363a,a17367a,a17368a,a17369a,a17373a,a17374a,a17378a,a17379a,a17380a,a17384a,a17385a,a17389a,a17390a,a17391a,a17395a,a17396a,a17400a,a17401a,a17402a,a17406a,a17407a,a17411a,a17412a,a17413a,a17417a,a17418a,a17422a,a17423a,a17424a,a17428a,a17429a,a17433a,a17434a,a17435a,a17439a,a17440a,a17444a,a17445a,a17446a,a17450a,a17451a,a17455a,a17456a,a17457a,a17461a,a17462a,a17466a,a17467a,a17468a,a17472a,a17473a,a17477a,a17478a,a17479a,a17483a,a17484a,a17488a,a17489a,a17490a,a17494a,a17495a,a17499a,a17500a,a17501a,a17505a,a17506a,a17510a,a17511a,a17512a,a17516a,a17517a,a17521a,a17522a,a17523a,a17527a,a17528a,a17532a,a17533a,a17534a,a17538a,a17539a,a17543a,a17544a,a17545a,a17549a,a17550a,a17554a,a17555a,a17556a,a17560a,a17561a,a17565a,a17566a,a17567a,a17571a,a17572a,a17576a,a17577a,a17578a,a17582a,a17583a,a17587a,a17588a,a17589a,a17593a,a17594a,a17598a,a17599a,a17600a,a17604a,a17605a,a17609a,a17610a,a17611a,a17615a,a17616a,a17620a,a17621a,a17622a,a17626a,a17627a,a17631a,a17632a,a17633a,a17637a,a17638a,a17642a,a17643a,a17644a,a17648a,a17649a,a17653a,a17654a,a17655a,a17659a,a17660a,a17664a,a17665a,a17666a,a17670a,a17671a,a17675a,a17676a,a17677a,a17681a,a17682a,a17686a,a17687a,a17688a,a17692a,a17693a,a17697a,a17698a,a17699a,a17703a,a17704a,a17708a,a17709a,a17710a,a17714a,a17715a,a17719a,a17720a,a17721a,a17725a,a17726a,a17730a,a17731a,a17732a,a17736a,a17737a,a17741a,a17742a,a17743a,a17747a,a17748a,a17752a,a17753a,a17754a,a17758a,a17759a,a17763a,a17764a,a17765a,a17769a,a17770a,a17774a,a17775a,a17776a,a17780a,a17781a,a17785a,a17786a,a17787a,a17791a,a17792a,a17796a,a17797a,a17798a,a17802a,a17803a,a17807a,a17808a,a17809a,a17813a,a17814a,a17818a,a17819a,a17820a,a17824a,a17825a,a17829a,a17830a,a17831a,a17835a,a17836a,a17840a,a17841a,a17842a,a17846a,a17847a,a17851a,a17852a,a17853a,a17857a,a17858a,a17862a,a17863a,a17864a,a17868a,a17869a,a17873a,a17874a,a17875a,a17879a,a17880a,a17884a,a17885a,a17886a,a17890a,a17891a,a17895a,a17896a,a17897a,a17901a,a17902a,a17906a,a17907a,a17908a,a17912a,a17913a,a17917a,a17918a,a17919a,a17923a,a17924a,a17928a,a17929a,a17930a,a17934a,a17935a,a17939a,a17940a,a17941a,a17945a,a17946a,a17950a,a17951a,a17952a,a17956a,a17957a,a17961a,a17962a,a17963a,a17967a,a17968a,a17972a,a17973a,a17974a,a17978a,a17979a,a17983a,a17984a,a17985a,a17989a,a17990a,a17994a,a17995a,a17996a,a18000a,a18001a,a18005a,a18006a,a18007a,a18011a,a18012a,a18016a,a18017a,a18018a,a18022a,a18023a,a18027a,a18028a,a18029a,a18033a,a18034a,a18038a,a18039a,a18040a,a18044a,a18045a,a18049a,a18050a,a18051a,a18055a,a18056a,a18060a,a18061a,a18062a,a18066a,a18067a,a18071a,a18072a,a18073a,a18077a,a18078a,a18082a,a18083a,a18084a,a18088a,a18089a,a18093a,a18094a,a18095a,a18099a,a18100a,a18104a,a18105a,a18106a,a18110a,a18111a,a18115a,a18116a,a18117a,a18121a,a18122a,a18126a,a18127a,a18128a,a18132a,a18133a,a18137a,a18138a,a18139a,a18143a,a18144a,a18148a,a18149a,a18150a,a18154a,a18155a,a18159a,a18160a,a18161a,a18165a,a18166a,a18170a,a18171a,a18172a,a18176a,a18177a,a18181a,a18182a,a18183a,a18187a,a18188a,a18192a,a18193a,a18194a,a18198a,a18199a,a18203a,a18204a,a18205a,a18209a,a18210a,a18214a,a18215a,a18216a,a18220a,a18221a,a18225a,a18226a,a18227a,a18231a,a18232a,a18236a,a18237a,a18238a,a18242a,a18243a,a18247a,a18248a,a18249a,a18253a,a18254a,a18258a,a18259a,a18260a,a18264a,a18265a,a18269a,a18270a,a18271a,a18275a,a18276a,a18280a,a18281a,a18282a,a18286a,a18287a,a18291a,a18292a,a18293a,a18297a,a18298a,a18302a,a18303a,a18304a,a18308a,a18309a,a18313a,a18314a,a18315a,a18319a,a18320a,a18324a,a18325a,a18326a,a18330a,a18331a,a18335a,a18336a,a18337a,a18341a,a18342a,a18346a,a18347a,a18348a,a18352a,a18353a,a18357a,a18358a,a18359a,a18363a,a18364a,a18368a,a18369a,a18370a,a18374a,a18375a,a18379a,a18380a,a18381a,a18385a,a18386a,a18390a,a18391a,a18392a,a18396a,a18397a,a18401a,a18402a,a18403a,a18407a,a18408a,a18412a,a18413a,a18414a,a18418a,a18419a,a18423a,a18424a,a18425a,a18429a,a18430a,a18434a,a18435a,a18436a,a18440a,a18441a,a18445a,a18446a,a18447a,a18451a,a18452a,a18456a,a18457a,a18458a,a18462a,a18463a,a18467a,a18468a,a18469a,a18473a,a18474a,a18478a,a18479a,a18480a,a18484a,a18485a,a18489a,a18490a,a18491a,a18495a,a18496a,a18500a,a18501a,a18502a,a18506a,a18507a,a18511a,a18512a,a18513a,a18517a,a18518a,a18522a,a18523a,a18524a,a18528a,a18529a,a18533a,a18534a,a18535a,a18539a,a18540a,a18544a,a18545a,a18546a,a18550a,a18551a,a18555a,a18556a,a18557a,a18561a,a18562a,a18566a,a18567a,a18568a,a18572a,a18573a,a18577a,a18578a,a18579a,a18583a,a18584a,a18588a,a18589a,a18590a,a18594a,a18595a,a18599a,a18600a,a18601a,a18605a,a18606a,a18610a,a18611a,a18612a,a18616a,a18617a,a18621a,a18622a,a18623a,a18627a,a18628a,a18632a,a18633a,a18634a,a18638a,a18639a,a18643a,a18644a,a18645a,a18649a,a18650a,a18654a,a18655a,a18656a,a18660a,a18661a,a18665a,a18666a,a18667a,a18671a,a18672a,a18676a,a18677a,a18678a,a18682a,a18683a,a18687a,a18688a,a18689a,a18693a,a18694a,a18698a,a18699a,a18700a,a18704a,a18705a,a18709a,a18710a,a18711a,a18715a,a18716a,a18720a,a18721a,a18722a,a18726a,a18727a,a18731a,a18732a,a18733a,a18737a,a18738a,a18742a,a18743a,a18744a,a18748a,a18749a,a18753a,a18754a,a18755a,a18759a,a18760a,a18764a,a18765a,a18766a,a18770a,a18771a,a18775a,a18776a,a18777a,a18781a,a18782a,a18786a,a18787a,a18788a,a18792a,a18793a,a18797a,a18798a,a18799a,a18803a,a18804a,a18808a,a18809a,a18810a,a18814a,a18815a,a18819a,a18820a,a18821a,a18825a,a18826a,a18830a,a18831a,a18832a,a18836a,a18837a,a18841a,a18842a,a18843a,a18847a,a18848a,a18852a,a18853a,a18854a,a18858a,a18859a,a18863a,a18864a,a18865a,a18869a,a18870a,a18874a,a18875a,a18876a,a18880a,a18881a,a18885a,a18886a,a18887a,a18891a,a18892a,a18896a,a18897a,a18898a,a18902a,a18903a,a18907a,a18908a,a18909a,a18913a,a18914a,a18918a,a18919a,a18920a,a18924a,a18925a,a18929a,a18930a,a18931a,a18935a,a18936a,a18940a,a18941a,a18942a,a18946a,a18947a,a18951a,a18952a,a18953a,a18957a,a18958a,a18962a,a18963a,a18964a,a18968a,a18969a,a18973a,a18974a,a18975a,a18979a,a18980a,a18984a,a18985a,a18986a,a18990a,a18991a,a18995a,a18996a,a18997a,a19001a,a19002a,a19006a,a19007a,a19008a,a19012a,a19013a,a19017a,a19018a,a19019a,a19023a,a19024a,a19028a,a19029a,a19030a,a19034a,a19035a,a19038a,a19041a,a19042a,a19043a,a19047a,a19048a,a19052a,a19053a,a19054a,a19058a,a19059a,a19062a,a19065a,a19066a,a19067a,a19071a,a19072a,a19076a,a19077a,a19078a,a19082a,a19083a,a19086a,a19089a,a19090a,a19091a,a19095a,a19096a,a19100a,a19101a,a19102a,a19106a,a19107a,a19110a,a19113a,a19114a,a19115a,a19119a,a19120a,a19124a,a19125a,a19126a,a19130a,a19131a,a19134a,a19137a,a19138a,a19139a,a19143a,a19144a,a19148a,a19149a,a19150a,a19154a,a19155a,a19158a,a19161a,a19162a,a19163a,a19167a,a19168a,a19172a,a19173a,a19174a,a19178a,a19179a,a19182a,a19185a,a19186a,a19187a,a19191a,a19192a,a19196a,a19197a,a19198a,a19202a,a19203a,a19206a,a19209a,a19210a,a19211a,a19215a,a19216a,a19220a,a19221a,a19222a,a19226a,a19227a,a19230a,a19233a,a19234a,a19235a,a19239a,a19240a,a19244a,a19245a,a19246a,a19250a,a19251a,a19254a,a19257a,a19258a,a19259a,a19263a,a19264a,a19268a,a19269a,a19270a,a19274a,a19275a,a19278a,a19281a,a19282a,a19283a,a19287a,a19288a,a19292a,a19293a,a19294a,a19298a,a19299a,a19302a,a19305a,a19306a,a19307a,a19311a,a19312a,a19316a,a19317a,a19318a,a19322a,a19323a,a19326a,a19329a,a19330a,a19331a,a19335a,a19336a,a19340a,a19341a,a19342a,a19346a,a19347a,a19350a,a19353a,a19354a,a19355a,a19359a,a19360a,a19364a,a19365a,a19366a,a19370a,a19371a,a19374a,a19377a,a19378a,a19379a,a19383a,a19384a,a19388a,a19389a,a19390a,a19394a,a19395a,a19398a,a19401a,a19402a,a19403a,a19407a,a19408a,a19412a,a19413a,a19414a,a19418a,a19419a,a19422a,a19425a,a19426a,a19427a,a19431a,a19432a,a19436a,a19437a,a19438a,a19442a,a19443a,a19446a,a19449a,a19450a,a19451a,a19455a,a19456a,a19460a,a19461a,a19462a,a19466a,a19467a,a19470a,a19473a,a19474a,a19475a,a19479a,a19480a,a19484a,a19485a,a19486a,a19490a,a19491a,a19494a,a19497a,a19498a,a19499a,a19503a,a19504a,a19508a,a19509a,a19510a,a19514a,a19515a,a19518a,a19521a,a19522a,a19523a,a19527a,a19528a,a19532a,a19533a,a19534a,a19538a,a19539a,a19542a,a19545a,a19546a,a19547a,a19551a,a19552a,a19556a,a19557a,a19558a,a19562a,a19563a,a19566a,a19569a,a19570a,a19571a,a19575a,a19576a,a19580a,a19581a,a19582a,a19586a,a19587a,a19590a,a19593a,a19594a,a19595a,a19599a,a19600a,a19604a,a19605a,a19606a,a19610a,a19611a,a19614a,a19617a,a19618a,a19619a,a19623a,a19624a,a19628a,a19629a,a19630a,a19634a,a19635a,a19638a,a19641a,a19642a,a19643a,a19647a,a19648a,a19652a,a19653a,a19654a,a19658a,a19659a,a19662a,a19665a,a19666a,a19667a,a19671a,a19672a,a19676a,a19677a,a19678a,a19682a,a19683a,a19686a,a19689a,a19690a,a19691a,a19695a,a19696a,a19700a,a19701a,a19702a,a19706a,a19707a,a19710a,a19713a,a19714a,a19715a,a19719a,a19720a,a19724a,a19725a,a19726a,a19730a,a19731a,a19734a,a19737a,a19738a,a19739a,a19743a,a19744a,a19748a,a19749a,a19750a,a19754a,a19755a,a19758a,a19761a,a19762a,a19763a,a19767a,a19768a,a19772a,a19773a,a19774a,a19778a,a19779a,a19782a,a19785a,a19786a,a19787a,a19791a,a19792a,a19796a,a19797a,a19798a,a19802a,a19803a,a19806a,a19809a,a19810a,a19811a,a19815a,a19816a,a19820a,a19821a,a19822a,a19826a,a19827a,a19830a,a19833a,a19834a,a19835a,a19839a,a19840a,a19844a,a19845a,a19846a,a19850a,a19851a,a19854a,a19857a,a19858a,a19859a,a19863a,a19864a,a19868a,a19869a,a19870a,a19874a,a19875a,a19878a,a19881a,a19882a,a19883a,a19887a,a19888a,a19892a,a19893a,a19894a,a19898a,a19899a,a19902a,a19905a,a19906a,a19907a,a19911a,a19912a,a19916a,a19917a,a19918a,a19922a,a19923a,a19926a,a19929a,a19930a,a19931a,a19935a,a19936a,a19940a,a19941a,a19942a,a19946a,a19947a,a19950a,a19953a,a19954a,a19955a,a19959a,a19960a,a19964a,a19965a,a19966a,a19970a,a19971a,a19974a,a19977a,a19978a,a19979a,a19983a,a19984a,a19988a,a19989a,a19990a,a19994a,a19995a,a19998a,a20001a,a20002a,a20003a,a20007a,a20008a,a20012a,a20013a,a20014a,a20018a,a20019a,a20022a,a20025a,a20026a,a20027a,a20031a,a20032a,a20036a,a20037a,a20038a,a20042a,a20043a,a20046a,a20049a,a20050a,a20051a,a20055a,a20056a,a20060a,a20061a,a20062a,a20066a,a20067a,a20070a,a20073a,a20074a,a20075a,a20079a,a20080a,a20084a,a20085a,a20086a,a20090a,a20091a,a20094a,a20097a,a20098a,a20099a,a20103a,a20104a,a20108a,a20109a,a20110a,a20114a,a20115a,a20118a,a20121a,a20122a,a20123a,a20127a,a20128a,a20132a,a20133a,a20134a,a20138a,a20139a,a20142a,a20145a,a20146a,a20147a,a20151a,a20152a,a20156a,a20157a,a20158a,a20162a,a20163a,a20166a,a20169a,a20170a,a20171a,a20175a,a20176a,a20180a,a20181a,a20182a,a20186a,a20187a,a20190a,a20193a,a20194a,a20195a,a20199a,a20200a,a20204a,a20205a,a20206a,a20210a,a20211a,a20214a,a20217a,a20218a,a20219a,a20223a,a20224a,a20228a,a20229a,a20230a,a20234a,a20235a,a20238a,a20241a,a20242a,a20243a,a20247a,a20248a,a20252a,a20253a,a20254a,a20258a,a20259a,a20262a,a20265a,a20266a,a20267a,a20271a,a20272a,a20276a,a20277a,a20278a,a20282a,a20283a,a20286a,a20289a,a20290a,a20291a,a20295a,a20296a,a20300a,a20301a,a20302a,a20306a,a20307a,a20310a,a20313a,a20314a,a20315a,a20319a,a20320a,a20324a,a20325a,a20326a,a20330a,a20331a,a20334a,a20337a,a20338a,a20339a,a20343a,a20344a,a20348a,a20349a,a20350a,a20354a,a20355a,a20358a,a20361a,a20362a,a20363a,a20367a,a20368a,a20372a,a20373a,a20374a,a20378a,a20379a,a20382a,a20385a,a20386a,a20387a,a20391a,a20392a,a20396a,a20397a,a20398a,a20402a,a20403a,a20406a,a20409a,a20410a,a20411a,a20415a,a20416a,a20420a,a20421a,a20422a,a20426a,a20427a,a20430a,a20433a,a20434a,a20435a,a20439a,a20440a,a20444a,a20445a,a20446a,a20450a,a20451a,a20454a,a20457a,a20458a,a20459a,a20463a,a20464a,a20468a,a20469a,a20470a,a20474a,a20475a,a20478a,a20481a,a20482a,a20483a,a20487a,a20488a,a20492a,a20493a,a20494a,a20498a,a20499a,a20502a,a20505a,a20506a,a20507a,a20511a,a20512a,a20516a,a20517a,a20518a,a20522a,a20523a,a20526a,a20529a,a20530a,a20531a,a20535a,a20536a,a20540a,a20541a,a20542a,a20546a,a20547a,a20550a,a20553a,a20554a,a20555a,a20559a,a20560a,a20564a,a20565a,a20566a,a20570a,a20571a,a20574a,a20577a,a20578a,a20579a,a20583a,a20584a,a20588a,a20589a,a20590a,a20594a,a20595a,a20598a,a20601a,a20602a,a20603a,a20607a,a20608a,a20612a,a20613a,a20614a,a20618a,a20619a,a20622a,a20625a,a20626a,a20627a,a20631a,a20632a,a20636a,a20637a,a20638a,a20642a,a20643a,a20646a,a20649a,a20650a,a20651a,a20655a,a20656a,a20660a,a20661a,a20662a,a20666a,a20667a,a20670a,a20673a,a20674a,a20675a,a20679a,a20680a,a20684a,a20685a,a20686a,a20690a,a20691a,a20694a,a20697a,a20698a,a20699a,a20703a,a20704a,a20708a,a20709a,a20710a,a20714a,a20715a,a20718a,a20721a,a20722a,a20723a,a20727a,a20728a,a20732a,a20733a,a20734a,a20738a,a20739a,a20742a,a20745a,a20746a,a20747a,a20751a,a20752a,a20756a,a20757a,a20758a,a20762a,a20763a,a20766a,a20769a,a20770a,a20771a,a20775a,a20776a,a20780a,a20781a,a20782a,a20786a,a20787a,a20790a,a20793a,a20794a,a20795a,a20799a,a20800a,a20804a,a20805a,a20806a,a20810a,a20811a,a20814a,a20817a,a20818a,a20819a,a20823a,a20824a,a20828a,a20829a,a20830a,a20834a,a20835a,a20838a,a20841a,a20842a,a20843a,a20847a,a20848a,a20852a,a20853a,a20854a,a20858a,a20859a,a20862a,a20865a,a20866a,a20867a,a20871a,a20872a,a20876a,a20877a,a20878a,a20882a,a20883a,a20886a,a20889a,a20890a,a20891a,a20895a,a20896a,a20900a,a20901a,a20902a,a20906a,a20907a,a20910a,a20913a,a20914a,a20915a,a20919a,a20920a,a20924a,a20925a,a20926a,a20930a,a20931a,a20934a,a20937a,a20938a,a20939a,a20943a,a20944a,a20948a,a20949a,a20950a,a20954a,a20955a,a20958a,a20961a,a20962a,a20963a,a20967a,a20968a,a20972a,a20973a,a20974a,a20978a,a20979a,a20982a,a20985a,a20986a,a20987a,a20991a,a20992a,a20996a,a20997a,a20998a,a21002a,a21003a,a21006a,a21009a,a21010a,a21011a,a21015a,a21016a,a21020a,a21021a,a21022a,a21026a,a21027a,a21030a,a21033a,a21034a,a21035a,a21039a,a21040a,a21044a,a21045a,a21046a,a21050a,a21051a,a21054a,a21057a,a21058a,a21059a,a21063a,a21064a,a21068a,a21069a,a21070a,a21074a,a21075a,a21078a,a21081a,a21082a,a21083a,a21087a,a21088a,a21092a,a21093a,a21094a,a21098a,a21099a,a21102a,a21105a,a21106a,a21107a,a21111a,a21112a,a21116a,a21117a,a21118a,a21122a,a21123a,a21126a,a21129a,a21130a,a21131a,a21135a,a21136a,a21140a,a21141a,a21142a,a21146a,a21147a,a21150a,a21153a,a21154a,a21155a,a21159a,a21160a,a21164a,a21165a,a21166a,a21170a,a21171a,a21174a,a21177a,a21178a,a21179a,a21183a,a21184a,a21188a,a21189a,a21190a,a21194a,a21195a,a21198a,a21201a,a21202a,a21203a,a21207a,a21208a,a21212a,a21213a,a21214a,a21218a,a21219a,a21222a,a21225a,a21226a,a21227a,a21231a,a21232a,a21236a,a21237a,a21238a,a21242a,a21243a,a21246a,a21249a,a21250a,a21251a,a21255a,a21256a,a21260a,a21261a,a21262a,a21266a,a21267a,a21270a,a21273a,a21274a,a21275a,a21279a,a21280a,a21284a,a21285a,a21286a,a21290a,a21291a,a21294a,a21297a,a21298a,a21299a,a21303a,a21304a,a21308a,a21309a,a21310a,a21314a,a21315a,a21318a,a21321a,a21322a,a21323a,a21327a,a21328a,a21332a,a21333a,a21334a,a21338a,a21339a,a21342a,a21345a,a21346a,a21347a,a21351a,a21352a,a21356a,a21357a,a21358a,a21362a,a21363a,a21366a,a21369a,a21370a,a21371a,a21375a,a21376a,a21380a,a21381a,a21382a,a21386a,a21387a,a21390a,a21393a,a21394a,a21395a,a21399a,a21400a,a21404a,a21405a,a21406a,a21410a,a21411a,a21414a,a21417a,a21418a,a21419a,a21423a,a21424a,a21428a,a21429a,a21430a,a21434a,a21435a,a21438a,a21441a,a21442a,a21443a,a21447a,a21448a,a21452a,a21453a,a21454a,a21458a,a21459a,a21462a,a21465a,a21466a,a21467a,a21471a,a21472a,a21476a,a21477a,a21478a,a21482a,a21483a,a21486a,a21489a,a21490a,a21491a,a21495a,a21496a,a21500a,a21501a,a21502a,a21506a,a21507a,a21510a,a21513a,a21514a,a21515a,a21519a,a21520a,a21524a,a21525a,a21526a,a21530a,a21531a,a21534a,a21537a,a21538a,a21539a,a21543a,a21544a,a21548a,a21549a,a21550a,a21554a,a21555a,a21558a,a21561a,a21562a,a21563a,a21567a,a21568a,a21572a,a21573a,a21574a,a21578a,a21579a,a21582a,a21585a,a21586a,a21587a,a21591a,a21592a,a21596a,a21597a,a21598a,a21602a,a21603a,a21606a,a21609a,a21610a,a21611a,a21615a,a21616a,a21620a,a21621a,a21622a,a21626a,a21627a,a21630a,a21633a,a21634a,a21635a,a21639a,a21640a,a21644a,a21645a,a21646a,a21650a,a21651a,a21654a,a21657a,a21658a,a21659a,a21663a,a21664a,a21668a,a21669a,a21670a,a21674a,a21675a,a21678a,a21681a,a21682a,a21683a,a21687a,a21688a,a21692a,a21693a,a21694a,a21698a,a21699a,a21702a,a21705a,a21706a,a21707a,a21711a,a21712a,a21716a,a21717a,a21718a,a21722a,a21723a,a21726a,a21729a,a21730a,a21731a,a21735a,a21736a,a21740a,a21741a,a21742a,a21746a,a21747a,a21750a,a21753a,a21754a,a21755a,a21759a,a21760a,a21764a,a21765a,a21766a,a21770a,a21771a,a21774a,a21777a,a21778a,a21779a,a21783a,a21784a,a21788a,a21789a,a21790a,a21794a,a21795a,a21798a,a21801a,a21802a,a21803a,a21807a,a21808a,a21812a,a21813a,a21814a,a21818a,a21819a,a21822a,a21825a,a21826a,a21827a,a21831a,a21832a,a21836a,a21837a,a21838a,a21842a,a21843a,a21846a,a21849a,a21850a,a21851a,a21855a,a21856a,a21860a,a21861a,a21862a,a21866a,a21867a,a21870a,a21873a,a21874a,a21875a,a21879a,a21880a,a21884a,a21885a,a21886a,a21890a,a21891a,a21894a,a21897a,a21898a,a21899a,a21903a,a21904a,a21908a,a21909a,a21910a,a21914a,a21915a,a21918a,a21921a,a21922a,a21923a,a21927a,a21928a,a21932a,a21933a,a21934a,a21938a,a21939a,a21942a,a21945a,a21946a,a21947a,a21951a,a21952a,a21956a,a21957a,a21958a,a21962a,a21963a,a21966a,a21969a,a21970a,a21971a,a21975a,a21976a,a21980a,a21981a,a21982a,a21986a,a21987a,a21990a,a21993a,a21994a,a21995a,a21999a,a22000a,a22004a,a22005a,a22006a,a22010a,a22011a,a22014a,a22017a,a22018a,a22019a,a22023a,a22024a,a22028a,a22029a,a22030a,a22034a,a22035a,a22038a,a22041a,a22042a,a22043a,a22047a,a22048a,a22052a,a22053a,a22054a,a22058a,a22059a,a22062a,a22065a,a22066a,a22067a,a22071a,a22072a,a22076a,a22077a,a22078a,a22082a,a22083a,a22086a,a22089a,a22090a,a22091a,a22095a,a22096a,a22100a,a22101a,a22102a,a22106a,a22107a,a22110a,a22113a,a22114a,a22115a,a22119a,a22120a,a22124a,a22125a,a22126a,a22130a,a22131a,a22134a,a22137a,a22138a,a22139a,a22143a,a22144a,a22148a,a22149a,a22150a,a22154a,a22155a,a22158a,a22161a,a22162a,a22163a,a22167a,a22168a,a22172a,a22173a,a22174a,a22178a,a22179a,a22182a,a22185a,a22186a,a22187a,a22191a,a22192a,a22196a,a22197a,a22198a,a22202a,a22203a,a22206a,a22209a,a22210a,a22211a,a22215a,a22216a,a22220a,a22221a,a22222a,a22226a,a22227a,a22230a,a22233a,a22234a,a22235a,a22239a,a22240a,a22244a,a22245a,a22246a,a22250a,a22251a,a22254a,a22257a,a22258a,a22259a,a22263a,a22264a,a22268a,a22269a,a22270a,a22274a,a22275a,a22278a,a22281a,a22282a,a22283a,a22287a,a22288a,a22292a,a22293a,a22294a,a22298a,a22299a,a22302a,a22305a,a22306a,a22307a,a22311a,a22312a,a22316a,a22317a,a22318a,a22322a,a22323a,a22326a,a22329a,a22330a,a22331a,a22335a,a22336a,a22340a,a22341a,a22342a,a22346a,a22347a,a22350a,a22353a,a22354a,a22355a,a22359a,a22360a,a22364a,a22365a,a22366a,a22370a,a22371a,a22374a,a22377a,a22378a,a22379a,a22383a,a22384a,a22388a,a22389a,a22390a,a22394a,a22395a,a22398a,a22401a,a22402a,a22403a,a22407a,a22408a,a22412a,a22413a,a22414a,a22418a,a22419a,a22422a,a22425a,a22426a,a22427a,a22431a,a22432a,a22436a,a22437a,a22438a,a22442a,a22443a,a22446a,a22449a,a22450a,a22451a,a22455a,a22456a,a22460a,a22461a,a22462a,a22466a,a22467a,a22470a,a22473a,a22474a,a22475a,a22479a,a22480a,a22484a,a22485a,a22486a,a22490a,a22491a,a22494a,a22497a,a22498a,a22499a,a22503a,a22504a,a22508a,a22509a,a22510a,a22514a,a22515a,a22518a,a22521a,a22522a,a22523a,a22527a,a22528a,a22532a,a22533a,a22534a,a22538a,a22539a,a22542a,a22545a,a22546a,a22547a,a22551a,a22552a,a22556a,a22557a,a22558a,a22562a,a22563a,a22566a,a22569a,a22570a,a22571a,a22575a,a22576a,a22580a,a22581a,a22582a,a22586a,a22587a,a22590a,a22593a,a22594a,a22595a,a22599a,a22600a,a22604a,a22605a,a22606a,a22610a,a22611a,a22614a,a22617a,a22618a,a22619a,a22623a,a22624a,a22628a,a22629a,a22630a,a22634a,a22635a,a22638a,a22641a,a22642a,a22643a,a22647a,a22648a,a22652a,a22653a,a22654a,a22658a,a22659a,a22662a,a22665a,a22666a,a22667a,a22671a,a22672a,a22676a,a22677a,a22678a,a22682a,a22683a,a22686a,a22689a,a22690a,a22691a,a22695a,a22696a,a22700a,a22701a,a22702a,a22706a,a22707a,a22710a,a22713a,a22714a,a22715a,a22719a,a22720a,a22724a,a22725a,a22726a,a22730a,a22731a,a22734a,a22737a,a22738a,a22739a,a22743a,a22744a,a22748a,a22749a,a22750a,a22754a,a22755a,a22758a,a22761a,a22762a,a22763a,a22767a,a22768a,a22772a,a22773a,a22774a,a22778a,a22779a,a22782a,a22785a,a22786a,a22787a,a22791a,a22792a,a22796a,a22797a,a22798a,a22802a,a22803a,a22806a,a22809a,a22810a,a22811a,a22815a,a22816a,a22820a,a22821a,a22822a,a22826a,a22827a,a22830a,a22833a,a22834a,a22835a,a22839a,a22840a,a22844a,a22845a,a22846a,a22850a,a22851a,a22854a,a22857a,a22858a,a22859a,a22863a,a22864a,a22868a,a22869a,a22870a,a22874a,a22875a,a22878a,a22881a,a22882a,a22883a,a22887a,a22888a,a22892a,a22893a,a22894a,a22898a,a22899a,a22902a,a22905a,a22906a,a22907a,a22911a,a22912a,a22916a,a22917a,a22918a,a22922a,a22923a,a22926a,a22929a,a22930a,a22931a,a22935a,a22936a,a22940a,a22941a,a22942a,a22946a,a22947a,a22950a,a22953a,a22954a,a22955a,a22959a,a22960a,a22964a,a22965a,a22966a,a22970a,a22971a,a22974a,a22977a,a22978a,a22979a,a22983a,a22984a,a22988a,a22989a,a22990a,a22994a,a22995a,a22998a,a23001a,a23002a,a23003a,a23007a,a23008a,a23012a,a23013a,a23014a,a23018a,a23019a,a23022a,a23025a,a23026a,a23027a,a23031a,a23032a,a23036a,a23037a,a23038a,a23042a,a23043a,a23046a,a23049a,a23050a,a23051a,a23055a,a23056a,a23060a,a23061a,a23062a,a23066a,a23067a,a23070a,a23073a,a23074a,a23075a,a23079a,a23080a,a23084a,a23085a,a23086a,a23090a,a23091a,a23094a,a23097a,a23098a,a23099a,a23103a,a23104a,a23108a,a23109a,a23110a,a23114a,a23115a,a23118a,a23121a,a23122a,a23123a,a23127a,a23128a,a23132a,a23133a,a23134a,a23138a,a23139a,a23142a,a23145a,a23146a,a23147a,a23151a,a23152a,a23156a,a23157a,a23158a,a23162a,a23163a,a23166a,a23169a,a23170a,a23171a,a23175a,a23176a,a23180a,a23181a,a23182a,a23186a,a23187a,a23190a,a23193a,a23194a,a23195a,a23199a,a23200a,a23204a,a23205a,a23206a,a23210a,a23211a,a23214a,a23217a,a23218a,a23219a,a23223a,a23224a,a23228a,a23229a,a23230a,a23234a,a23235a,a23238a,a23241a,a23242a,a23243a,a23247a,a23248a,a23251a,a23254a,a23255a,a23256a,a23260a,a23261a,a23264a,a23267a,a23268a,a23269a,a23273a,a23274a,a23277a,a23280a,a23281a,a23282a,a23286a,a23287a,a23290a,a23293a,a23294a,a23295a,a23299a,a23300a,a23303a,a23306a,a23307a,a23308a,a23312a,a23313a,a23316a,a23319a,a23320a,a23321a,a23325a,a23326a,a23329a,a23332a,a23333a,a23334a,a23338a,a23339a,a23342a,a23345a,a23346a,a23347a,a23351a,a23352a,a23355a,a23358a,a23359a,a23360a,a23364a,a23365a,a23368a,a23371a,a23372a,a23373a,a23377a,a23378a,a23381a,a23384a,a23385a,a23386a,a23390a,a23391a,a23394a,a23397a,a23398a,a23399a,a23403a,a23404a,a23407a,a23410a,a23411a,a23412a,a23416a,a23417a,a23420a,a23423a,a23424a,a23425a,a23429a,a23430a,a23433a,a23436a,a23437a,a23438a,a23442a,a23443a,a23446a,a23449a,a23450a,a23451a,a23455a,a23456a,a23459a,a23462a,a23463a,a23464a,a23468a,a23469a,a23472a,a23475a,a23476a,a23477a,a23481a,a23482a,a23485a,a23488a,a23489a,a23490a,a23494a,a23495a,a23498a,a23501a,a23502a,a23503a,a23507a,a23508a,a23511a,a23514a,a23515a,a23516a,a23520a,a23521a,a23524a,a23527a,a23528a,a23529a,a23533a,a23534a,a23537a,a23540a,a23541a,a23542a,a23546a,a23547a,a23550a,a23553a,a23554a,a23555a,a23559a,a23560a,a23563a,a23566a,a23567a,a23568a,a23572a,a23573a,a23576a,a23579a,a23580a,a23581a,a23585a,a23586a,a23589a,a23592a,a23593a,a23594a,a23598a,a23599a,a23602a,a23605a,a23606a,a23607a,a23611a,a23612a,a23615a,a23618a,a23619a,a23620a,a23624a,a23625a,a23628a,a23631a,a23632a,a23633a,a23637a,a23638a,a23641a,a23644a,a23645a,a23646a,a23650a,a23651a,a23654a,a23657a,a23658a,a23659a,a23663a,a23664a,a23667a,a23670a,a23671a,a23672a,a23676a,a23677a,a23680a,a23683a,a23684a,a23685a,a23689a,a23690a,a23693a,a23696a,a23697a,a23698a,a23702a,a23703a,a23706a,a23709a,a23710a,a23711a,a23715a,a23716a,a23719a,a23722a,a23723a,a23724a,a23728a,a23729a,a23732a,a23735a,a23736a,a23737a,a23741a,a23742a,a23745a,a23748a,a23749a,a23750a,a23754a,a23755a,a23758a,a23761a,a23762a,a23763a,a23767a,a23768a,a23771a,a23774a,a23775a,a23776a,a23780a,a23781a,a23784a,a23787a,a23788a,a23789a,a23793a,a23794a,a23797a,a23800a,a23801a,a23802a,a23806a,a23807a,a23810a,a23813a,a23814a,a23815a,a23819a,a23820a,a23823a,a23826a,a23827a,a23828a,a23832a,a23833a,a23836a,a23839a,a23840a,a23841a,a23845a,a23846a,a23849a,a23852a,a23853a,a23854a,a23858a,a23859a,a23862a,a23865a,a23866a,a23867a,a23871a,a23872a,a23875a,a23878a,a23879a,a23880a,a23884a,a23885a,a23888a,a23891a,a23892a,a23893a,a23897a,a23898a,a23901a,a23904a,a23905a,a23906a,a23910a,a23911a,a23914a,a23917a,a23918a,a23919a,a23923a,a23924a,a23927a,a23930a,a23931a,a23932a,a23936a,a23937a,a23940a,a23943a,a23944a,a23945a,a23949a,a23950a,a23953a,a23956a,a23957a,a23958a,a23962a,a23963a,a23966a,a23969a,a23970a,a23971a,a23975a,a23976a,a23979a,a23982a,a23983a,a23984a,a23988a,a23989a,a23992a,a23995a,a23996a,a23997a,a24001a,a24002a,a24005a,a24008a,a24009a,a24010a,a24014a,a24015a,a24018a,a24021a,a24022a,a24023a,a24027a,a24028a,a24031a,a24034a,a24035a,a24036a,a24040a,a24041a,a24044a,a24047a,a24048a,a24049a,a24053a,a24054a,a24057a,a24060a,a24061a,a24062a,a24066a,a24067a,a24070a,a24073a,a24074a,a24075a,a24079a,a24080a,a24083a,a24086a,a24087a,a24088a,a24092a,a24093a,a24096a,a24099a,a24100a,a24101a,a24105a,a24106a,a24109a,a24112a,a24113a,a24114a,a24118a,a24119a,a24122a,a24125a,a24126a,a24127a,a24131a,a24132a,a24135a,a24138a,a24139a,a24140a,a24144a,a24145a,a24148a,a24151a,a24152a,a24153a,a24157a,a24158a,a24161a,a24164a,a24165a,a24166a,a24170a,a24171a,a24174a,a24177a,a24178a,a24179a,a24183a,a24184a,a24187a,a24190a,a24191a,a24192a,a24196a,a24197a,a24200a,a24203a,a24204a,a24205a,a24209a,a24210a,a24213a,a24216a,a24217a,a24218a,a24222a,a24223a,a24226a,a24229a,a24230a,a24231a,a24235a,a24236a,a24239a,a24242a,a24243a,a24244a,a24248a,a24249a,a24252a,a24255a,a24256a,a24257a,a24261a,a24262a,a24265a,a24268a,a24269a,a24270a,a24274a,a24275a,a24278a,a24281a,a24282a,a24283a,a24287a,a24288a,a24291a,a24294a,a24295a,a24296a,a24300a,a24301a,a24304a,a24307a,a24308a,a24309a,a24313a,a24314a,a24317a,a24320a,a24321a,a24322a,a24326a,a24327a,a24330a,a24333a,a24334a,a24335a,a24339a,a24340a,a24343a,a24346a,a24347a,a24348a,a24352a,a24353a,a24356a,a24359a,a24360a,a24361a,a24365a,a24366a,a24369a,a24372a,a24373a,a24374a,a24378a,a24379a,a24382a,a24385a,a24386a,a24387a,a24391a,a24392a,a24395a,a24398a,a24399a,a24400a,a24404a,a24405a,a24408a,a24411a,a24412a,a24413a,a24417a,a24418a,a24421a,a24424a,a24425a,a24426a,a24430a,a24431a,a24434a,a24437a,a24438a,a24439a,a24443a,a24444a,a24447a,a24450a,a24451a,a24452a,a24456a,a24457a,a24460a,a24463a,a24464a,a24465a,a24469a,a24470a,a24473a,a24476a,a24477a,a24478a,a24482a,a24483a,a24486a,a24489a,a24490a,a24491a,a24495a,a24496a,a24499a,a24502a,a24503a,a24504a,a24508a,a24509a,a24512a,a24515a,a24516a,a24517a,a24521a,a24522a,a24525a,a24528a,a24529a,a24530a,a24534a,a24535a,a24538a,a24541a,a24542a,a24543a,a24547a,a24548a,a24551a,a24554a,a24555a,a24556a,a24560a,a24561a,a24564a,a24567a,a24568a,a24569a,a24573a,a24574a,a24577a,a24580a,a24581a,a24582a,a24586a,a24587a,a24590a,a24593a,a24594a,a24595a,a24599a,a24600a,a24603a,a24606a,a24607a,a24608a,a24612a,a24613a,a24616a,a24619a,a24620a,a24621a,a24625a,a24626a,a24629a,a24632a,a24633a,a24634a,a24638a,a24639a,a24642a,a24645a,a24646a,a24647a,a24651a,a24652a,a24655a,a24658a,a24659a,a24660a,a24664a,a24665a,a24668a,a24671a,a24672a,a24673a,a24677a,a24678a,a24681a,a24684a,a24685a,a24686a,a24690a,a24691a,a24694a,a24697a,a24698a,a24699a,a24703a,a24704a,a24707a,a24710a,a24711a,a24712a,a24716a,a24717a,a24720a,a24723a,a24724a,a24725a,a24729a,a24730a,a24733a,a24736a,a24737a,a24738a,a24742a,a24743a,a24746a,a24749a,a24750a,a24751a,a24755a,a24756a,a24759a,a24762a,a24763a,a24764a,a24768a,a24769a,a24772a,a24775a,a24776a,a24777a,a24781a,a24782a,a24785a,a24788a,a24789a,a24790a,a24794a,a24795a,a24798a,a24801a,a24802a,a24803a,a24807a,a24808a,a24811a,a24814a,a24815a,a24816a,a24820a,a24821a,a24824a,a24827a,a24828a,a24829a,a24833a,a24834a,a24837a,a24840a,a24841a,a24842a,a24846a,a24847a,a24850a,a24853a,a24854a,a24855a,a24859a,a24860a,a24863a,a24866a,a24867a,a24868a,a24872a,a24873a,a24876a,a24879a,a24880a,a24881a,a24885a,a24886a,a24889a,a24892a,a24893a,a24894a,a24898a,a24899a,a24902a,a24905a,a24906a,a24907a,a24911a,a24912a,a24915a,a24918a,a24919a,a24920a,a24924a,a24925a,a24928a,a24931a,a24932a,a24933a,a24937a,a24938a,a24941a,a24944a,a24945a,a24946a,a24950a,a24951a,a24954a,a24957a,a24958a,a24959a,a24963a,a24964a,a24967a,a24970a,a24971a,a24972a,a24976a,a24977a,a24980a,a24983a,a24984a,a24985a,a24989a,a24990a,a24993a,a24996a,a24997a,a24998a,a25002a,a25003a,a25006a,a25009a,a25010a,a25011a,a25015a,a25016a,a25019a,a25022a,a25023a,a25024a,a25028a,a25029a,a25032a,a25035a,a25036a,a25037a,a25041a,a25042a,a25045a,a25048a,a25049a,a25050a,a25054a,a25055a,a25058a,a25061a,a25062a,a25063a,a25067a,a25068a,a25071a,a25074a,a25075a,a25076a,a25080a,a25081a,a25084a,a25087a,a25088a,a25089a,a25093a,a25094a,a25097a,a25100a,a25101a,a25102a,a25106a,a25107a,a25110a,a25113a,a25114a,a25115a,a25119a,a25120a,a25123a,a25126a,a25127a,a25128a,a25132a,a25133a,a25136a,a25139a,a25140a,a25141a,a25145a,a25146a,a25149a,a25152a,a25153a,a25154a,a25158a,a25159a,a25162a,a25165a,a25166a,a25167a,a25171a,a25172a,a25175a,a25178a,a25179a,a25180a,a25184a,a25185a,a25188a,a25191a,a25192a,a25193a,a25197a,a25198a,a25201a,a25204a,a25205a,a25206a,a25210a,a25211a,a25214a,a25217a,a25218a,a25219a,a25223a,a25224a,a25227a,a25230a,a25231a,a25232a,a25236a,a25237a,a25240a,a25243a,a25244a,a25245a,a25249a,a25250a,a25253a,a25256a,a25257a,a25258a,a25262a,a25263a,a25266a,a25269a,a25270a,a25271a,a25275a,a25276a,a25279a,a25282a,a25283a,a25284a,a25288a,a25289a,a25292a,a25295a,a25296a,a25297a,a25301a,a25302a,a25305a,a25308a,a25309a,a25310a,a25314a,a25315a,a25318a,a25321a,a25322a,a25323a,a25327a,a25328a,a25331a,a25334a,a25335a,a25336a,a25340a,a25341a,a25344a,a25347a,a25348a,a25349a,a25353a,a25354a,a25357a,a25360a,a25361a,a25362a,a25366a,a25367a,a25370a,a25373a,a25374a,a25375a,a25379a,a25380a,a25383a,a25386a,a25387a,a25388a,a25392a,a25393a,a25396a,a25399a,a25400a,a25401a,a25405a,a25406a,a25409a,a25412a,a25413a,a25414a,a25418a,a25419a,a25422a,a25425a,a25426a,a25427a,a25431a,a25432a,a25435a,a25438a,a25439a,a25440a,a25444a,a25445a,a25448a,a25451a,a25452a,a25453a,a25457a,a25458a,a25461a,a25464a,a25465a,a25466a,a25470a,a25471a,a25474a,a25477a,a25478a,a25479a,a25483a,a25484a,a25487a,a25490a,a25491a,a25492a,a25496a,a25497a,a25500a,a25503a,a25504a,a25505a,a25509a,a25510a,a25513a,a25516a,a25517a,a25518a,a25522a,a25523a,a25526a,a25529a,a25530a,a25531a,a25535a,a25536a,a25539a,a25542a,a25543a,a25544a,a25548a,a25549a,a25552a,a25555a,a25556a,a25557a,a25561a,a25562a,a25565a,a25568a,a25569a,a25570a,a25574a,a25575a,a25578a,a25581a,a25582a,a25583a,a25587a,a25588a,a25591a,a25594a,a25595a,a25596a,a25600a,a25601a,a25604a,a25607a,a25608a,a25609a,a25613a,a25614a,a25617a,a25620a,a25621a,a25622a,a25626a,a25627a,a25630a,a25633a,a25634a,a25635a,a25639a,a25640a,a25643a,a25646a,a25647a,a25648a,a25652a,a25653a,a25656a,a25659a,a25660a,a25661a,a25665a,a25666a,a25669a,a25672a,a25673a,a25674a,a25678a,a25679a,a25682a,a25685a,a25686a,a25687a,a25691a,a25692a,a25695a,a25698a,a25699a,a25700a,a25704a,a25705a,a25708a,a25711a,a25712a,a25713a,a25717a,a25718a,a25721a,a25724a,a25725a,a25726a,a25730a,a25731a,a25734a,a25737a,a25738a,a25739a,a25743a,a25744a,a25747a,a25750a,a25751a,a25752a,a25756a,a25757a,a25760a,a25763a,a25764a,a25765a,a25769a,a25770a,a25773a,a25776a,a25777a,a25778a,a25782a,a25783a,a25786a,a25789a,a25790a,a25791a,a25795a,a25796a,a25799a,a25802a,a25803a,a25804a,a25808a,a25809a,a25812a,a25815a,a25816a,a25817a,a25821a,a25822a,a25825a,a25828a,a25829a,a25830a,a25834a,a25835a,a25838a,a25841a,a25842a,a25843a,a25847a,a25848a,a25851a,a25854a,a25855a,a25856a,a25860a,a25861a,a25864a,a25867a,a25868a,a25869a,a25873a,a25874a,a25877a,a25880a,a25881a,a25882a,a25886a,a25887a,a25890a,a25893a,a25894a,a25895a,a25899a,a25900a,a25903a,a25906a,a25907a,a25908a,a25912a,a25913a,a25916a,a25919a,a25920a,a25921a,a25925a,a25926a,a25929a,a25932a,a25933a,a25934a,a25938a,a25939a,a25942a,a25945a,a25946a,a25947a,a25951a,a25952a,a25955a,a25958a,a25959a,a25960a,a25964a,a25965a,a25968a,a25971a,a25972a,a25973a,a25977a,a25978a,a25981a,a25984a,a25985a,a25986a,a25990a,a25991a,a25994a,a25997a,a25998a,a25999a,a26003a,a26004a,a26007a,a26010a,a26011a,a26012a,a26016a,a26017a,a26020a,a26023a,a26024a,a26025a,a26029a,a26030a,a26033a,a26036a,a26037a,a26038a,a26042a,a26043a,a26046a,a26049a,a26050a,a26051a,a26055a,a26056a,a26059a,a26062a,a26063a,a26064a,a26068a,a26069a,a26072a,a26075a,a26076a,a26077a,a26081a,a26082a,a26085a,a26088a,a26089a,a26090a,a26094a,a26095a,a26098a,a26101a,a26102a,a26103a,a26107a,a26108a,a26111a,a26114a,a26115a,a26116a,a26120a,a26121a,a26124a,a26127a,a26128a,a26129a,a26133a,a26134a,a26137a,a26140a,a26141a,a26142a,a26146a,a26147a,a26150a,a26153a,a26154a,a26155a,a26159a,a26160a,a26163a,a26166a,a26167a,a26168a,a26172a,a26173a,a26176a,a26179a,a26180a,a26181a,a26185a,a26186a,a26189a,a26192a,a26193a,a26194a,a26198a,a26199a,a26202a,a26205a,a26206a,a26207a,a26211a,a26212a,a26215a,a26218a,a26219a,a26220a,a26223a,a26226a,a26227a,a26230a,a26233a,a26234a,a26235a,a26239a,a26240a,a26243a,a26246a,a26247a,a26248a,a26251a,a26254a,a26255a,a26258a,a26261a,a26262a,a26263a,a26267a,a26268a,a26271a,a26274a,a26275a,a26276a,a26279a,a26282a,a26283a,a26286a,a26289a,a26290a,a26291a,a26295a,a26296a,a26299a,a26302a,a26303a,a26304a,a26307a,a26310a,a26311a,a26314a,a26317a,a26318a,a26319a,a26323a,a26324a,a26327a,a26330a,a26331a,a26332a,a26335a,a26338a,a26339a,a26342a,a26345a,a26346a,a26347a,a26351a,a26352a,a26355a,a26358a,a26359a,a26360a,a26363a,a26366a,a26367a,a26370a,a26373a,a26374a,a26375a,a26379a,a26380a,a26383a,a26386a,a26387a,a26388a,a26391a,a26394a,a26395a,a26398a,a26401a,a26402a,a26403a,a26407a,a26408a,a26411a,a26414a,a26415a,a26416a,a26419a,a26422a,a26423a,a26426a,a26429a,a26430a,a26431a,a26435a,a26436a,a26439a,a26442a,a26443a,a26444a,a26447a,a26450a,a26451a,a26454a,a26457a,a26458a,a26459a,a26463a,a26464a,a26467a,a26470a,a26471a,a26472a,a26475a,a26478a,a26479a,a26482a,a26485a,a26486a,a26487a,a26491a,a26492a,a26495a,a26498a,a26499a,a26500a,a26503a,a26506a,a26507a,a26510a,a26513a,a26514a,a26515a,a26519a,a26520a,a26523a,a26526a,a26527a,a26528a,a26531a,a26534a,a26535a,a26538a,a26541a,a26542a,a26543a,a26547a,a26548a,a26551a,a26554a,a26555a,a26556a,a26559a,a26562a,a26563a,a26566a,a26569a,a26570a,a26571a,a26575a,a26576a,a26579a,a26582a,a26583a,a26584a,a26587a,a26590a,a26591a,a26594a,a26597a,a26598a,a26599a,a26603a,a26604a,a26607a,a26610a,a26611a,a26612a,a26615a,a26618a,a26619a,a26622a,a26625a,a26626a,a26627a,a26631a,a26632a,a26635a,a26638a,a26639a,a26640a,a26643a,a26646a,a26647a,a26650a,a26653a,a26654a,a26655a,a26659a,a26660a,a26663a,a26666a,a26667a,a26668a,a26671a,a26674a,a26675a,a26678a,a26681a,a26682a,a26683a,a26687a,a26688a,a26691a,a26694a,a26695a,a26696a,a26699a,a26702a,a26703a,a26706a,a26709a,a26710a,a26711a,a26715a,a26716a,a26719a,a26722a,a26723a,a26724a,a26727a,a26730a,a26731a,a26734a,a26737a,a26738a,a26739a,a26743a,a26744a,a26747a,a26750a,a26751a,a26752a,a26755a,a26758a,a26759a,a26762a,a26765a,a26766a,a26767a,a26771a,a26772a,a26775a,a26778a,a26779a,a26780a,a26783a,a26786a,a26787a,a26790a,a26793a,a26794a,a26795a,a26799a,a26800a,a26803a,a26806a,a26807a,a26808a,a26811a,a26814a,a26815a,a26818a,a26821a,a26822a,a26823a,a26827a,a26828a,a26831a,a26834a,a26835a,a26836a,a26839a,a26842a,a26843a,a26846a,a26849a,a26850a,a26851a,a26855a,a26856a,a26859a,a26862a,a26863a,a26864a,a26867a,a26870a,a26871a,a26874a,a26877a,a26878a,a26879a,a26883a,a26884a,a26887a,a26890a,a26891a,a26892a,a26895a,a26898a,a26899a,a26902a,a26905a,a26906a,a26907a,a26911a,a26912a,a26915a,a26918a,a26919a,a26920a,a26923a,a26926a,a26927a,a26930a,a26933a,a26934a,a26935a,a26939a,a26940a,a26943a,a26946a,a26947a,a26948a,a26951a,a26954a,a26955a,a26958a,a26961a,a26962a,a26963a,a26967a,a26968a,a26971a,a26974a,a26975a,a26976a,a26979a,a26982a,a26983a,a26986a,a26989a,a26990a,a26991a: std_logic;
begin

A106 <=( a3355a ) or ( a2236a );
 a1a <=( a26991a  and  a26976a );
 a2a <=( a26963a  and  a26948a );
 a3a <=( a26935a  and  a26920a );
 a4a <=( a26907a  and  a26892a );
 a5a <=( a26879a  and  a26864a );
 a6a <=( a26851a  and  a26836a );
 a7a <=( a26823a  and  a26808a );
 a8a <=( a26795a  and  a26780a );
 a9a <=( a26767a  and  a26752a );
 a10a <=( a26739a  and  a26724a );
 a11a <=( a26711a  and  a26696a );
 a12a <=( a26683a  and  a26668a );
 a13a <=( a26655a  and  a26640a );
 a14a <=( a26627a  and  a26612a );
 a15a <=( a26599a  and  a26584a );
 a16a <=( a26571a  and  a26556a );
 a17a <=( a26543a  and  a26528a );
 a18a <=( a26515a  and  a26500a );
 a19a <=( a26487a  and  a26472a );
 a20a <=( a26459a  and  a26444a );
 a21a <=( a26431a  and  a26416a );
 a22a <=( a26403a  and  a26388a );
 a23a <=( a26375a  and  a26360a );
 a24a <=( a26347a  and  a26332a );
 a25a <=( a26319a  and  a26304a );
 a26a <=( a26291a  and  a26276a );
 a27a <=( a26263a  and  a26248a );
 a28a <=( a26235a  and  a26220a );
 a29a <=( a26207a  and  a26194a );
 a30a <=( a26181a  and  a26168a );
 a31a <=( a26155a  and  a26142a );
 a32a <=( a26129a  and  a26116a );
 a33a <=( a26103a  and  a26090a );
 a34a <=( a26077a  and  a26064a );
 a35a <=( a26051a  and  a26038a );
 a36a <=( a26025a  and  a26012a );
 a37a <=( a25999a  and  a25986a );
 a38a <=( a25973a  and  a25960a );
 a39a <=( a25947a  and  a25934a );
 a40a <=( a25921a  and  a25908a );
 a41a <=( a25895a  and  a25882a );
 a42a <=( a25869a  and  a25856a );
 a43a <=( a25843a  and  a25830a );
 a44a <=( a25817a  and  a25804a );
 a45a <=( a25791a  and  a25778a );
 a46a <=( a25765a  and  a25752a );
 a47a <=( a25739a  and  a25726a );
 a48a <=( a25713a  and  a25700a );
 a49a <=( a25687a  and  a25674a );
 a50a <=( a25661a  and  a25648a );
 a51a <=( a25635a  and  a25622a );
 a52a <=( a25609a  and  a25596a );
 a53a <=( a25583a  and  a25570a );
 a54a <=( a25557a  and  a25544a );
 a55a <=( a25531a  and  a25518a );
 a56a <=( a25505a  and  a25492a );
 a57a <=( a25479a  and  a25466a );
 a58a <=( a25453a  and  a25440a );
 a59a <=( a25427a  and  a25414a );
 a60a <=( a25401a  and  a25388a );
 a61a <=( a25375a  and  a25362a );
 a62a <=( a25349a  and  a25336a );
 a63a <=( a25323a  and  a25310a );
 a64a <=( a25297a  and  a25284a );
 a65a <=( a25271a  and  a25258a );
 a66a <=( a25245a  and  a25232a );
 a67a <=( a25219a  and  a25206a );
 a68a <=( a25193a  and  a25180a );
 a69a <=( a25167a  and  a25154a );
 a70a <=( a25141a  and  a25128a );
 a71a <=( a25115a  and  a25102a );
 a72a <=( a25089a  and  a25076a );
 a73a <=( a25063a  and  a25050a );
 a74a <=( a25037a  and  a25024a );
 a75a <=( a25011a  and  a24998a );
 a76a <=( a24985a  and  a24972a );
 a77a <=( a24959a  and  a24946a );
 a78a <=( a24933a  and  a24920a );
 a79a <=( a24907a  and  a24894a );
 a80a <=( a24881a  and  a24868a );
 a81a <=( a24855a  and  a24842a );
 a82a <=( a24829a  and  a24816a );
 a83a <=( a24803a  and  a24790a );
 a84a <=( a24777a  and  a24764a );
 a85a <=( a24751a  and  a24738a );
 a86a <=( a24725a  and  a24712a );
 a87a <=( a24699a  and  a24686a );
 a88a <=( a24673a  and  a24660a );
 a89a <=( a24647a  and  a24634a );
 a90a <=( a24621a  and  a24608a );
 a91a <=( a24595a  and  a24582a );
 a92a <=( a24569a  and  a24556a );
 a93a <=( a24543a  and  a24530a );
 a94a <=( a24517a  and  a24504a );
 a95a <=( a24491a  and  a24478a );
 a96a <=( a24465a  and  a24452a );
 a97a <=( a24439a  and  a24426a );
 a98a <=( a24413a  and  a24400a );
 a99a <=( a24387a  and  a24374a );
 a100a <=( a24361a  and  a24348a );
 a101a <=( a24335a  and  a24322a );
 a102a <=( a24309a  and  a24296a );
 a103a <=( a24283a  and  a24270a );
 a104a <=( a24257a  and  a24244a );
 a105a <=( a24231a  and  a24218a );
 a106a <=( a24205a  and  a24192a );
 a107a <=( a24179a  and  a24166a );
 a108a <=( a24153a  and  a24140a );
 a109a <=( a24127a  and  a24114a );
 a110a <=( a24101a  and  a24088a );
 a111a <=( a24075a  and  a24062a );
 a112a <=( a24049a  and  a24036a );
 a113a <=( a24023a  and  a24010a );
 a114a <=( a23997a  and  a23984a );
 a115a <=( a23971a  and  a23958a );
 a116a <=( a23945a  and  a23932a );
 a117a <=( a23919a  and  a23906a );
 a118a <=( a23893a  and  a23880a );
 a119a <=( a23867a  and  a23854a );
 a120a <=( a23841a  and  a23828a );
 a121a <=( a23815a  and  a23802a );
 a122a <=( a23789a  and  a23776a );
 a123a <=( a23763a  and  a23750a );
 a124a <=( a23737a  and  a23724a );
 a125a <=( a23711a  and  a23698a );
 a126a <=( a23685a  and  a23672a );
 a127a <=( a23659a  and  a23646a );
 a128a <=( a23633a  and  a23620a );
 a129a <=( a23607a  and  a23594a );
 a130a <=( a23581a  and  a23568a );
 a131a <=( a23555a  and  a23542a );
 a132a <=( a23529a  and  a23516a );
 a133a <=( a23503a  and  a23490a );
 a134a <=( a23477a  and  a23464a );
 a135a <=( a23451a  and  a23438a );
 a136a <=( a23425a  and  a23412a );
 a137a <=( a23399a  and  a23386a );
 a138a <=( a23373a  and  a23360a );
 a139a <=( a23347a  and  a23334a );
 a140a <=( a23321a  and  a23308a );
 a141a <=( a23295a  and  a23282a );
 a142a <=( a23269a  and  a23256a );
 a143a <=( a23243a  and  a23230a );
 a144a <=( a23219a  and  a23206a );
 a145a <=( a23195a  and  a23182a );
 a146a <=( a23171a  and  a23158a );
 a147a <=( a23147a  and  a23134a );
 a148a <=( a23123a  and  a23110a );
 a149a <=( a23099a  and  a23086a );
 a150a <=( a23075a  and  a23062a );
 a151a <=( a23051a  and  a23038a );
 a152a <=( a23027a  and  a23014a );
 a153a <=( a23003a  and  a22990a );
 a154a <=( a22979a  and  a22966a );
 a155a <=( a22955a  and  a22942a );
 a156a <=( a22931a  and  a22918a );
 a157a <=( a22907a  and  a22894a );
 a158a <=( a22883a  and  a22870a );
 a159a <=( a22859a  and  a22846a );
 a160a <=( a22835a  and  a22822a );
 a161a <=( a22811a  and  a22798a );
 a162a <=( a22787a  and  a22774a );
 a163a <=( a22763a  and  a22750a );
 a164a <=( a22739a  and  a22726a );
 a165a <=( a22715a  and  a22702a );
 a166a <=( a22691a  and  a22678a );
 a167a <=( a22667a  and  a22654a );
 a168a <=( a22643a  and  a22630a );
 a169a <=( a22619a  and  a22606a );
 a170a <=( a22595a  and  a22582a );
 a171a <=( a22571a  and  a22558a );
 a172a <=( a22547a  and  a22534a );
 a173a <=( a22523a  and  a22510a );
 a174a <=( a22499a  and  a22486a );
 a175a <=( a22475a  and  a22462a );
 a176a <=( a22451a  and  a22438a );
 a177a <=( a22427a  and  a22414a );
 a178a <=( a22403a  and  a22390a );
 a179a <=( a22379a  and  a22366a );
 a180a <=( a22355a  and  a22342a );
 a181a <=( a22331a  and  a22318a );
 a182a <=( a22307a  and  a22294a );
 a183a <=( a22283a  and  a22270a );
 a184a <=( a22259a  and  a22246a );
 a185a <=( a22235a  and  a22222a );
 a186a <=( a22211a  and  a22198a );
 a187a <=( a22187a  and  a22174a );
 a188a <=( a22163a  and  a22150a );
 a189a <=( a22139a  and  a22126a );
 a190a <=( a22115a  and  a22102a );
 a191a <=( a22091a  and  a22078a );
 a192a <=( a22067a  and  a22054a );
 a193a <=( a22043a  and  a22030a );
 a194a <=( a22019a  and  a22006a );
 a195a <=( a21995a  and  a21982a );
 a196a <=( a21971a  and  a21958a );
 a197a <=( a21947a  and  a21934a );
 a198a <=( a21923a  and  a21910a );
 a199a <=( a21899a  and  a21886a );
 a200a <=( a21875a  and  a21862a );
 a201a <=( a21851a  and  a21838a );
 a202a <=( a21827a  and  a21814a );
 a203a <=( a21803a  and  a21790a );
 a204a <=( a21779a  and  a21766a );
 a205a <=( a21755a  and  a21742a );
 a206a <=( a21731a  and  a21718a );
 a207a <=( a21707a  and  a21694a );
 a208a <=( a21683a  and  a21670a );
 a209a <=( a21659a  and  a21646a );
 a210a <=( a21635a  and  a21622a );
 a211a <=( a21611a  and  a21598a );
 a212a <=( a21587a  and  a21574a );
 a213a <=( a21563a  and  a21550a );
 a214a <=( a21539a  and  a21526a );
 a215a <=( a21515a  and  a21502a );
 a216a <=( a21491a  and  a21478a );
 a217a <=( a21467a  and  a21454a );
 a218a <=( a21443a  and  a21430a );
 a219a <=( a21419a  and  a21406a );
 a220a <=( a21395a  and  a21382a );
 a221a <=( a21371a  and  a21358a );
 a222a <=( a21347a  and  a21334a );
 a223a <=( a21323a  and  a21310a );
 a224a <=( a21299a  and  a21286a );
 a225a <=( a21275a  and  a21262a );
 a226a <=( a21251a  and  a21238a );
 a227a <=( a21227a  and  a21214a );
 a228a <=( a21203a  and  a21190a );
 a229a <=( a21179a  and  a21166a );
 a230a <=( a21155a  and  a21142a );
 a231a <=( a21131a  and  a21118a );
 a232a <=( a21107a  and  a21094a );
 a233a <=( a21083a  and  a21070a );
 a234a <=( a21059a  and  a21046a );
 a235a <=( a21035a  and  a21022a );
 a236a <=( a21011a  and  a20998a );
 a237a <=( a20987a  and  a20974a );
 a238a <=( a20963a  and  a20950a );
 a239a <=( a20939a  and  a20926a );
 a240a <=( a20915a  and  a20902a );
 a241a <=( a20891a  and  a20878a );
 a242a <=( a20867a  and  a20854a );
 a243a <=( a20843a  and  a20830a );
 a244a <=( a20819a  and  a20806a );
 a245a <=( a20795a  and  a20782a );
 a246a <=( a20771a  and  a20758a );
 a247a <=( a20747a  and  a20734a );
 a248a <=( a20723a  and  a20710a );
 a249a <=( a20699a  and  a20686a );
 a250a <=( a20675a  and  a20662a );
 a251a <=( a20651a  and  a20638a );
 a252a <=( a20627a  and  a20614a );
 a253a <=( a20603a  and  a20590a );
 a254a <=( a20579a  and  a20566a );
 a255a <=( a20555a  and  a20542a );
 a256a <=( a20531a  and  a20518a );
 a257a <=( a20507a  and  a20494a );
 a258a <=( a20483a  and  a20470a );
 a259a <=( a20459a  and  a20446a );
 a260a <=( a20435a  and  a20422a );
 a261a <=( a20411a  and  a20398a );
 a262a <=( a20387a  and  a20374a );
 a263a <=( a20363a  and  a20350a );
 a264a <=( a20339a  and  a20326a );
 a265a <=( a20315a  and  a20302a );
 a266a <=( a20291a  and  a20278a );
 a267a <=( a20267a  and  a20254a );
 a268a <=( a20243a  and  a20230a );
 a269a <=( a20219a  and  a20206a );
 a270a <=( a20195a  and  a20182a );
 a271a <=( a20171a  and  a20158a );
 a272a <=( a20147a  and  a20134a );
 a273a <=( a20123a  and  a20110a );
 a274a <=( a20099a  and  a20086a );
 a275a <=( a20075a  and  a20062a );
 a276a <=( a20051a  and  a20038a );
 a277a <=( a20027a  and  a20014a );
 a278a <=( a20003a  and  a19990a );
 a279a <=( a19979a  and  a19966a );
 a280a <=( a19955a  and  a19942a );
 a281a <=( a19931a  and  a19918a );
 a282a <=( a19907a  and  a19894a );
 a283a <=( a19883a  and  a19870a );
 a284a <=( a19859a  and  a19846a );
 a285a <=( a19835a  and  a19822a );
 a286a <=( a19811a  and  a19798a );
 a287a <=( a19787a  and  a19774a );
 a288a <=( a19763a  and  a19750a );
 a289a <=( a19739a  and  a19726a );
 a290a <=( a19715a  and  a19702a );
 a291a <=( a19691a  and  a19678a );
 a292a <=( a19667a  and  a19654a );
 a293a <=( a19643a  and  a19630a );
 a294a <=( a19619a  and  a19606a );
 a295a <=( a19595a  and  a19582a );
 a296a <=( a19571a  and  a19558a );
 a297a <=( a19547a  and  a19534a );
 a298a <=( a19523a  and  a19510a );
 a299a <=( a19499a  and  a19486a );
 a300a <=( a19475a  and  a19462a );
 a301a <=( a19451a  and  a19438a );
 a302a <=( a19427a  and  a19414a );
 a303a <=( a19403a  and  a19390a );
 a304a <=( a19379a  and  a19366a );
 a305a <=( a19355a  and  a19342a );
 a306a <=( a19331a  and  a19318a );
 a307a <=( a19307a  and  a19294a );
 a308a <=( a19283a  and  a19270a );
 a309a <=( a19259a  and  a19246a );
 a310a <=( a19235a  and  a19222a );
 a311a <=( a19211a  and  a19198a );
 a312a <=( a19187a  and  a19174a );
 a313a <=( a19163a  and  a19150a );
 a314a <=( a19139a  and  a19126a );
 a315a <=( a19115a  and  a19102a );
 a316a <=( a19091a  and  a19078a );
 a317a <=( a19067a  and  a19054a );
 a318a <=( a19043a  and  a19030a );
 a319a <=( a19019a  and  a19008a );
 a320a <=( a18997a  and  a18986a );
 a321a <=( a18975a  and  a18964a );
 a322a <=( a18953a  and  a18942a );
 a323a <=( a18931a  and  a18920a );
 a324a <=( a18909a  and  a18898a );
 a325a <=( a18887a  and  a18876a );
 a326a <=( a18865a  and  a18854a );
 a327a <=( a18843a  and  a18832a );
 a328a <=( a18821a  and  a18810a );
 a329a <=( a18799a  and  a18788a );
 a330a <=( a18777a  and  a18766a );
 a331a <=( a18755a  and  a18744a );
 a332a <=( a18733a  and  a18722a );
 a333a <=( a18711a  and  a18700a );
 a334a <=( a18689a  and  a18678a );
 a335a <=( a18667a  and  a18656a );
 a336a <=( a18645a  and  a18634a );
 a337a <=( a18623a  and  a18612a );
 a338a <=( a18601a  and  a18590a );
 a339a <=( a18579a  and  a18568a );
 a340a <=( a18557a  and  a18546a );
 a341a <=( a18535a  and  a18524a );
 a342a <=( a18513a  and  a18502a );
 a343a <=( a18491a  and  a18480a );
 a344a <=( a18469a  and  a18458a );
 a345a <=( a18447a  and  a18436a );
 a346a <=( a18425a  and  a18414a );
 a347a <=( a18403a  and  a18392a );
 a348a <=( a18381a  and  a18370a );
 a349a <=( a18359a  and  a18348a );
 a350a <=( a18337a  and  a18326a );
 a351a <=( a18315a  and  a18304a );
 a352a <=( a18293a  and  a18282a );
 a353a <=( a18271a  and  a18260a );
 a354a <=( a18249a  and  a18238a );
 a355a <=( a18227a  and  a18216a );
 a356a <=( a18205a  and  a18194a );
 a357a <=( a18183a  and  a18172a );
 a358a <=( a18161a  and  a18150a );
 a359a <=( a18139a  and  a18128a );
 a360a <=( a18117a  and  a18106a );
 a361a <=( a18095a  and  a18084a );
 a362a <=( a18073a  and  a18062a );
 a363a <=( a18051a  and  a18040a );
 a364a <=( a18029a  and  a18018a );
 a365a <=( a18007a  and  a17996a );
 a366a <=( a17985a  and  a17974a );
 a367a <=( a17963a  and  a17952a );
 a368a <=( a17941a  and  a17930a );
 a369a <=( a17919a  and  a17908a );
 a370a <=( a17897a  and  a17886a );
 a371a <=( a17875a  and  a17864a );
 a372a <=( a17853a  and  a17842a );
 a373a <=( a17831a  and  a17820a );
 a374a <=( a17809a  and  a17798a );
 a375a <=( a17787a  and  a17776a );
 a376a <=( a17765a  and  a17754a );
 a377a <=( a17743a  and  a17732a );
 a378a <=( a17721a  and  a17710a );
 a379a <=( a17699a  and  a17688a );
 a380a <=( a17677a  and  a17666a );
 a381a <=( a17655a  and  a17644a );
 a382a <=( a17633a  and  a17622a );
 a383a <=( a17611a  and  a17600a );
 a384a <=( a17589a  and  a17578a );
 a385a <=( a17567a  and  a17556a );
 a386a <=( a17545a  and  a17534a );
 a387a <=( a17523a  and  a17512a );
 a388a <=( a17501a  and  a17490a );
 a389a <=( a17479a  and  a17468a );
 a390a <=( a17457a  and  a17446a );
 a391a <=( a17435a  and  a17424a );
 a392a <=( a17413a  and  a17402a );
 a393a <=( a17391a  and  a17380a );
 a394a <=( a17369a  and  a17358a );
 a395a <=( a17347a  and  a17336a );
 a396a <=( a17325a  and  a17314a );
 a397a <=( a17303a  and  a17292a );
 a398a <=( a17281a  and  a17270a );
 a399a <=( a17259a  and  a17248a );
 a400a <=( a17237a  and  a17226a );
 a401a <=( a17215a  and  a17204a );
 a402a <=( a17193a  and  a17182a );
 a403a <=( a17171a  and  a17160a );
 a404a <=( a17149a  and  a17138a );
 a405a <=( a17127a  and  a17116a );
 a406a <=( a17105a  and  a17094a );
 a407a <=( a17083a  and  a17072a );
 a408a <=( a17061a  and  a17050a );
 a409a <=( a17039a  and  a17028a );
 a410a <=( a17017a  and  a17006a );
 a411a <=( a16995a  and  a16984a );
 a412a <=( a16973a  and  a16962a );
 a413a <=( a16951a  and  a16940a );
 a414a <=( a16929a  and  a16918a );
 a415a <=( a16907a  and  a16896a );
 a416a <=( a16885a  and  a16874a );
 a417a <=( a16863a  and  a16852a );
 a418a <=( a16841a  and  a16830a );
 a419a <=( a16819a  and  a16808a );
 a420a <=( a16797a  and  a16786a );
 a421a <=( a16775a  and  a16764a );
 a422a <=( a16753a  and  a16742a );
 a423a <=( a16731a  and  a16720a );
 a424a <=( a16709a  and  a16698a );
 a425a <=( a16687a  and  a16676a );
 a426a <=( a16665a  and  a16654a );
 a427a <=( a16643a  and  a16632a );
 a428a <=( a16621a  and  a16610a );
 a429a <=( a16599a  and  a16588a );
 a430a <=( a16577a  and  a16566a );
 a431a <=( a16555a  and  a16544a );
 a432a <=( a16533a  and  a16522a );
 a433a <=( a16511a  and  a16500a );
 a434a <=( a16489a  and  a16478a );
 a435a <=( a16467a  and  a16456a );
 a436a <=( a16445a  and  a16434a );
 a437a <=( a16423a  and  a16412a );
 a438a <=( a16401a  and  a16390a );
 a439a <=( a16379a  and  a16368a );
 a440a <=( a16357a  and  a16346a );
 a441a <=( a16335a  and  a16324a );
 a442a <=( a16313a  and  a16302a );
 a443a <=( a16291a  and  a16280a );
 a444a <=( a16269a  and  a16258a );
 a445a <=( a16247a  and  a16236a );
 a446a <=( a16225a  and  a16214a );
 a447a <=( a16203a  and  a16192a );
 a448a <=( a16181a  and  a16170a );
 a449a <=( a16159a  and  a16148a );
 a450a <=( a16137a  and  a16126a );
 a451a <=( a16115a  and  a16104a );
 a452a <=( a16093a  and  a16082a );
 a453a <=( a16071a  and  a16060a );
 a454a <=( a16049a  and  a16038a );
 a455a <=( a16027a  and  a16016a );
 a456a <=( a16005a  and  a15994a );
 a457a <=( a15983a  and  a15972a );
 a458a <=( a15961a  and  a15950a );
 a459a <=( a15939a  and  a15928a );
 a460a <=( a15917a  and  a15906a );
 a461a <=( a15895a  and  a15884a );
 a462a <=( a15873a  and  a15862a );
 a463a <=( a15851a  and  a15840a );
 a464a <=( a15829a  and  a15818a );
 a465a <=( a15807a  and  a15796a );
 a466a <=( a15785a  and  a15774a );
 a467a <=( a15763a  and  a15752a );
 a468a <=( a15741a  and  a15730a );
 a469a <=( a15719a  and  a15708a );
 a470a <=( a15697a  and  a15686a );
 a471a <=( a15675a  and  a15664a );
 a472a <=( a15653a  and  a15642a );
 a473a <=( a15631a  and  a15620a );
 a474a <=( a15609a  and  a15598a );
 a475a <=( a15587a  and  a15576a );
 a476a <=( a15565a  and  a15554a );
 a477a <=( a15543a  and  a15532a );
 a478a <=( a15521a  and  a15510a );
 a479a <=( a15499a  and  a15488a );
 a480a <=( a15477a  and  a15466a );
 a481a <=( a15455a  and  a15444a );
 a482a <=( a15433a  and  a15422a );
 a483a <=( a15411a  and  a15400a );
 a484a <=( a15389a  and  a15378a );
 a485a <=( a15367a  and  a15356a );
 a486a <=( a15345a  and  a15334a );
 a487a <=( a15323a  and  a15312a );
 a488a <=( a15301a  and  a15290a );
 a489a <=( a15279a  and  a15268a );
 a490a <=( a15257a  and  a15246a );
 a491a <=( a15235a  and  a15224a );
 a492a <=( a15213a  and  a15202a );
 a493a <=( a15191a  and  a15180a );
 a494a <=( a15169a  and  a15158a );
 a495a <=( a15147a  and  a15136a );
 a496a <=( a15125a  and  a15114a );
 a497a <=( a15103a  and  a15092a );
 a498a <=( a15081a  and  a15070a );
 a499a <=( a15059a  and  a15048a );
 a500a <=( a15037a  and  a15026a );
 a501a <=( a15015a  and  a15004a );
 a502a <=( a14993a  and  a14982a );
 a503a <=( a14971a  and  a14960a );
 a504a <=( a14949a  and  a14938a );
 a505a <=( a14927a  and  a14916a );
 a506a <=( a14905a  and  a14894a );
 a507a <=( a14883a  and  a14872a );
 a508a <=( a14861a  and  a14850a );
 a509a <=( a14839a  and  a14828a );
 a510a <=( a14817a  and  a14806a );
 a511a <=( a14795a  and  a14784a );
 a512a <=( a14773a  and  a14762a );
 a513a <=( a14751a  and  a14740a );
 a514a <=( a14729a  and  a14718a );
 a515a <=( a14707a  and  a14696a );
 a516a <=( a14685a  and  a14674a );
 a517a <=( a14663a  and  a14652a );
 a518a <=( a14641a  and  a14630a );
 a519a <=( a14619a  and  a14608a );
 a520a <=( a14597a  and  a14586a );
 a521a <=( a14575a  and  a14564a );
 a522a <=( a14553a  and  a14542a );
 a523a <=( a14531a  and  a14520a );
 a524a <=( a14509a  and  a14498a );
 a525a <=( a14487a  and  a14476a );
 a526a <=( a14465a  and  a14454a );
 a527a <=( a14443a  and  a14432a );
 a528a <=( a14421a  and  a14410a );
 a529a <=( a14399a  and  a14388a );
 a530a <=( a14377a  and  a14366a );
 a531a <=( a14355a  and  a14344a );
 a532a <=( a14333a  and  a14322a );
 a533a <=( a14311a  and  a14300a );
 a534a <=( a14289a  and  a14278a );
 a535a <=( a14267a  and  a14256a );
 a536a <=( a14245a  and  a14234a );
 a537a <=( a14223a  and  a14212a );
 a538a <=( a14201a  and  a14190a );
 a539a <=( a14179a  and  a14168a );
 a540a <=( a14157a  and  a14146a );
 a541a <=( a14135a  and  a14124a );
 a542a <=( a14113a  and  a14102a );
 a543a <=( a14091a  and  a14080a );
 a544a <=( a14069a  and  a14058a );
 a545a <=( a14047a  and  a14036a );
 a546a <=( a14025a  and  a14014a );
 a547a <=( a14003a  and  a13992a );
 a548a <=( a13981a  and  a13970a );
 a549a <=( a13959a  and  a13948a );
 a550a <=( a13937a  and  a13926a );
 a551a <=( a13915a  and  a13904a );
 a552a <=( a13893a  and  a13882a );
 a553a <=( a13871a  and  a13860a );
 a554a <=( a13849a  and  a13838a );
 a555a <=( a13827a  and  a13816a );
 a556a <=( a13805a  and  a13794a );
 a557a <=( a13783a  and  a13772a );
 a558a <=( a13761a  and  a13750a );
 a559a <=( a13739a  and  a13728a );
 a560a <=( a13717a  and  a13706a );
 a561a <=( a13695a  and  a13684a );
 a562a <=( a13673a  and  a13662a );
 a563a <=( a13651a  and  a13640a );
 a564a <=( a13629a  and  a13618a );
 a565a <=( a13607a  and  a13596a );
 a566a <=( a13585a  and  a13574a );
 a567a <=( a13563a  and  a13552a );
 a568a <=( a13541a  and  a13530a );
 a569a <=( a13519a  and  a13508a );
 a570a <=( a13497a  and  a13486a );
 a571a <=( a13475a  and  a13464a );
 a572a <=( a13453a  and  a13442a );
 a573a <=( a13431a  and  a13420a );
 a574a <=( a13409a  and  a13398a );
 a575a <=( a13387a  and  a13376a );
 a576a <=( a13365a  and  a13354a );
 a577a <=( a13343a  and  a13332a );
 a578a <=( a13321a  and  a13310a );
 a579a <=( a13299a  and  a13288a );
 a580a <=( a13277a  and  a13266a );
 a581a <=( a13255a  and  a13244a );
 a582a <=( a13233a  and  a13222a );
 a583a <=( a13211a  and  a13200a );
 a584a <=( a13189a  and  a13178a );
 a585a <=( a13167a  and  a13156a );
 a586a <=( a13145a  and  a13134a );
 a587a <=( a13123a  and  a13112a );
 a588a <=( a13101a  and  a13090a );
 a589a <=( a13079a  and  a13068a );
 a590a <=( a13057a  and  a13046a );
 a591a <=( a13035a  and  a13024a );
 a592a <=( a13013a  and  a13002a );
 a593a <=( a12991a  and  a12980a );
 a594a <=( a12969a  and  a12958a );
 a595a <=( a12947a  and  a12936a );
 a596a <=( a12925a  and  a12914a );
 a597a <=( a12903a  and  a12892a );
 a598a <=( a12881a  and  a12870a );
 a599a <=( a12859a  and  a12848a );
 a600a <=( a12837a  and  a12826a );
 a601a <=( a12815a  and  a12804a );
 a602a <=( a12793a  and  a12782a );
 a603a <=( a12771a  and  a12760a );
 a604a <=( a12749a  and  a12738a );
 a605a <=( a12727a  and  a12716a );
 a606a <=( a12705a  and  a12694a );
 a607a <=( a12683a  and  a12672a );
 a608a <=( a12661a  and  a12650a );
 a609a <=( a12639a  and  a12628a );
 a610a <=( a12617a  and  a12606a );
 a611a <=( a12595a  and  a12584a );
 a612a <=( a12573a  and  a12562a );
 a613a <=( a12551a  and  a12540a );
 a614a <=( a12529a  and  a12518a );
 a615a <=( a12507a  and  a12496a );
 a616a <=( a12485a  and  a12474a );
 a617a <=( a12463a  and  a12452a );
 a618a <=( a12441a  and  a12430a );
 a619a <=( a12419a  and  a12408a );
 a620a <=( a12397a  and  a12386a );
 a621a <=( a12375a  and  a12364a );
 a622a <=( a12353a  and  a12342a );
 a623a <=( a12331a  and  a12320a );
 a624a <=( a12309a  and  a12298a );
 a625a <=( a12287a  and  a12276a );
 a626a <=( a12265a  and  a12254a );
 a627a <=( a12243a  and  a12232a );
 a628a <=( a12221a  and  a12210a );
 a629a <=( a12201a  and  a12190a );
 a630a <=( a12181a  and  a12170a );
 a631a <=( a12161a  and  a12150a );
 a632a <=( a12141a  and  a12130a );
 a633a <=( a12121a  and  a12110a );
 a634a <=( a12101a  and  a12090a );
 a635a <=( a12081a  and  a12070a );
 a636a <=( a12061a  and  a12050a );
 a637a <=( a12041a  and  a12030a );
 a638a <=( a12021a  and  a12010a );
 a639a <=( a12001a  and  a11990a );
 a640a <=( a11981a  and  a11970a );
 a641a <=( a11961a  and  a11950a );
 a642a <=( a11941a  and  a11930a );
 a643a <=( a11921a  and  a11910a );
 a644a <=( a11901a  and  a11890a );
 a645a <=( a11881a  and  a11870a );
 a646a <=( a11861a  and  a11850a );
 a647a <=( a11841a  and  a11830a );
 a648a <=( a11821a  and  a11810a );
 a649a <=( a11801a  and  a11790a );
 a650a <=( a11781a  and  a11770a );
 a651a <=( a11761a  and  a11750a );
 a652a <=( a11741a  and  a11730a );
 a653a <=( a11721a  and  a11710a );
 a654a <=( a11701a  and  a11690a );
 a655a <=( a11681a  and  a11670a );
 a656a <=( a11661a  and  a11650a );
 a657a <=( a11641a  and  a11630a );
 a658a <=( a11621a  and  a11610a );
 a659a <=( a11601a  and  a11590a );
 a660a <=( a11581a  and  a11570a );
 a661a <=( a11561a  and  a11550a );
 a662a <=( a11541a  and  a11530a );
 a663a <=( a11521a  and  a11510a );
 a664a <=( a11501a  and  a11490a );
 a665a <=( a11481a  and  a11470a );
 a666a <=( a11461a  and  a11450a );
 a667a <=( a11441a  and  a11430a );
 a668a <=( a11421a  and  a11410a );
 a669a <=( a11401a  and  a11390a );
 a670a <=( a11381a  and  a11370a );
 a671a <=( a11361a  and  a11350a );
 a672a <=( a11341a  and  a11330a );
 a673a <=( a11321a  and  a11310a );
 a674a <=( a11301a  and  a11290a );
 a675a <=( a11281a  and  a11270a );
 a676a <=( a11261a  and  a11250a );
 a677a <=( a11241a  and  a11230a );
 a678a <=( a11221a  and  a11210a );
 a679a <=( a11201a  and  a11190a );
 a680a <=( a11181a  and  a11170a );
 a681a <=( a11161a  and  a11150a );
 a682a <=( a11141a  and  a11130a );
 a683a <=( a11121a  and  a11110a );
 a684a <=( a11101a  and  a11090a );
 a685a <=( a11081a  and  a11070a );
 a686a <=( a11061a  and  a11050a );
 a687a <=( a11041a  and  a11030a );
 a688a <=( a11021a  and  a11010a );
 a689a <=( a11001a  and  a10990a );
 a690a <=( a10981a  and  a10970a );
 a691a <=( a10961a  and  a10950a );
 a692a <=( a10941a  and  a10930a );
 a693a <=( a10921a  and  a10910a );
 a694a <=( a10901a  and  a10890a );
 a695a <=( a10881a  and  a10870a );
 a696a <=( a10861a  and  a10850a );
 a697a <=( a10841a  and  a10830a );
 a698a <=( a10821a  and  a10810a );
 a699a <=( a10801a  and  a10790a );
 a700a <=( a10781a  and  a10770a );
 a701a <=( a10761a  and  a10750a );
 a702a <=( a10741a  and  a10730a );
 a703a <=( a10721a  and  a10710a );
 a704a <=( a10701a  and  a10690a );
 a705a <=( a10681a  and  a10670a );
 a706a <=( a10661a  and  a10650a );
 a707a <=( a10641a  and  a10630a );
 a708a <=( a10621a  and  a10610a );
 a709a <=( a10601a  and  a10590a );
 a710a <=( a10581a  and  a10570a );
 a711a <=( a10561a  and  a10550a );
 a712a <=( a10541a  and  a10530a );
 a713a <=( a10521a  and  a10510a );
 a714a <=( a10501a  and  a10490a );
 a715a <=( a10481a  and  a10470a );
 a716a <=( a10461a  and  a10450a );
 a717a <=( a10441a  and  a10430a );
 a718a <=( a10421a  and  a10410a );
 a719a <=( a10401a  and  a10390a );
 a720a <=( a10381a  and  a10370a );
 a721a <=( a10361a  and  a10350a );
 a722a <=( a10341a  and  a10330a );
 a723a <=( a10321a  and  a10310a );
 a724a <=( a10301a  and  a10290a );
 a725a <=( a10281a  and  a10270a );
 a726a <=( a10261a  and  a10250a );
 a727a <=( a10241a  and  a10230a );
 a728a <=( a10221a  and  a10210a );
 a729a <=( a10201a  and  a10190a );
 a730a <=( a10181a  and  a10170a );
 a731a <=( a10161a  and  a10150a );
 a732a <=( a10141a  and  a10130a );
 a733a <=( a10121a  and  a10110a );
 a734a <=( a10101a  and  a10090a );
 a735a <=( a10081a  and  a10070a );
 a736a <=( a10061a  and  a10050a );
 a737a <=( a10041a  and  a10030a );
 a738a <=( a10021a  and  a10010a );
 a739a <=( a10001a  and  a9990a );
 a740a <=( a9981a  and  a9970a );
 a741a <=( a9961a  and  a9950a );
 a742a <=( a9941a  and  a9930a );
 a743a <=( a9921a  and  a9910a );
 a744a <=( a9901a  and  a9890a );
 a745a <=( a9881a  and  a9870a );
 a746a <=( a9861a  and  a9850a );
 a747a <=( a9841a  and  a9830a );
 a748a <=( a9821a  and  a9810a );
 a749a <=( a9801a  and  a9790a );
 a750a <=( a9781a  and  a9770a );
 a751a <=( a9761a  and  a9750a );
 a752a <=( a9741a  and  a9730a );
 a753a <=( a9721a  and  a9710a );
 a754a <=( a9701a  and  a9690a );
 a755a <=( a9681a  and  a9670a );
 a756a <=( a9661a  and  a9650a );
 a757a <=( a9641a  and  a9630a );
 a758a <=( a9621a  and  a9610a );
 a759a <=( a9601a  and  a9590a );
 a760a <=( a9581a  and  a9570a );
 a761a <=( a9561a  and  a9550a );
 a762a <=( a9541a  and  a9530a );
 a763a <=( a9521a  and  a9510a );
 a764a <=( a9501a  and  a9490a );
 a765a <=( a9481a  and  a9470a );
 a766a <=( a9461a  and  a9450a );
 a767a <=( a9441a  and  a9430a );
 a768a <=( a9421a  and  a9410a );
 a769a <=( a9401a  and  a9390a );
 a770a <=( a9381a  and  a9370a );
 a771a <=( a9361a  and  a9350a );
 a772a <=( a9341a  and  a9330a );
 a773a <=( a9321a  and  a9310a );
 a774a <=( a9301a  and  a9290a );
 a775a <=( a9281a  and  a9270a );
 a776a <=( a9261a  and  a9250a );
 a777a <=( a9241a  and  a9230a );
 a778a <=( a9221a  and  a9210a );
 a779a <=( a9201a  and  a9190a );
 a780a <=( a9181a  and  a9170a );
 a781a <=( a9161a  and  a9150a );
 a782a <=( a9141a  and  a9130a );
 a783a <=( a9121a  and  a9110a );
 a784a <=( a9101a  and  a9090a );
 a785a <=( a9081a  and  a9070a );
 a786a <=( a9061a  and  a9050a );
 a787a <=( a9041a  and  a9030a );
 a788a <=( a9021a  and  a9010a );
 a789a <=( a9001a  and  a8990a );
 a790a <=( a8981a  and  a8970a );
 a791a <=( a8961a  and  a8950a );
 a792a <=( a8941a  and  a8930a );
 a793a <=( a8921a  and  a8910a );
 a794a <=( a8901a  and  a8890a );
 a795a <=( a8881a  and  a8870a );
 a796a <=( a8861a  and  a8850a );
 a797a <=( a8841a  and  a8830a );
 a798a <=( a8821a  and  a8810a );
 a799a <=( a8801a  and  a8790a );
 a800a <=( a8781a  and  a8770a );
 a801a <=( a8761a  and  a8750a );
 a802a <=( a8741a  and  a8730a );
 a803a <=( a8721a  and  a8710a );
 a804a <=( a8701a  and  a8690a );
 a805a <=( a8681a  and  a8670a );
 a806a <=( a8661a  and  a8650a );
 a807a <=( a8641a  and  a8630a );
 a808a <=( a8621a  and  a8610a );
 a809a <=( a8601a  and  a8590a );
 a810a <=( a8581a  and  a8570a );
 a811a <=( a8561a  and  a8550a );
 a812a <=( a8541a  and  a8530a );
 a813a <=( a8521a  and  a8510a );
 a814a <=( a8501a  and  a8490a );
 a815a <=( a8481a  and  a8470a );
 a816a <=( a8461a  and  a8450a );
 a817a <=( a8441a  and  a8430a );
 a818a <=( a8421a  and  a8410a );
 a819a <=( a8401a  and  a8390a );
 a820a <=( a8381a  and  a8370a );
 a821a <=( a8361a  and  a8350a );
 a822a <=( a8341a  and  a8330a );
 a823a <=( a8321a  and  a8310a );
 a824a <=( a8301a  and  a8290a );
 a825a <=( a8281a  and  a8270a );
 a826a <=( a8261a  and  a8250a );
 a827a <=( a8241a  and  a8230a );
 a828a <=( a8221a  and  a8210a );
 a829a <=( a8201a  and  a8190a );
 a830a <=( a8181a  and  a8170a );
 a831a <=( a8161a  and  a8150a );
 a832a <=( a8141a  and  a8130a );
 a833a <=( a8121a  and  a8112a );
 a834a <=( a8103a  and  a8094a );
 a835a <=( a8085a  and  a8076a );
 a836a <=( a8067a  and  a8058a );
 a837a <=( a8049a  and  a8040a );
 a838a <=( a8031a  and  a8022a );
 a839a <=( a8013a  and  a8004a );
 a840a <=( a7995a  and  a7986a );
 a841a <=( a7977a  and  a7968a );
 a842a <=( a7959a  and  a7950a );
 a843a <=( a7941a  and  a7932a );
 a844a <=( a7923a  and  a7914a );
 a845a <=( a7905a  and  a7896a );
 a846a <=( a7887a  and  a7878a );
 a847a <=( a7869a  and  a7860a );
 a848a <=( a7851a  and  a7842a );
 a849a <=( a7833a  and  a7824a );
 a850a <=( a7815a  and  a7806a );
 a851a <=( a7797a  and  a7788a );
 a852a <=( a7779a  and  a7770a );
 a853a <=( a7761a  and  a7752a );
 a854a <=( a7743a  and  a7734a );
 a855a <=( a7725a  and  a7716a );
 a856a <=( a7707a  and  a7698a );
 a857a <=( a7689a  and  a7680a );
 a858a <=( a7671a  and  a7662a );
 a859a <=( a7653a  and  a7644a );
 a860a <=( a7635a  and  a7626a );
 a861a <=( a7617a  and  a7608a );
 a862a <=( a7599a  and  a7590a );
 a863a <=( a7581a  and  a7572a );
 a864a <=( a7563a  and  a7554a );
 a865a <=( a7545a  and  a7536a );
 a866a <=( a7527a  and  a7518a );
 a867a <=( a7509a  and  a7500a );
 a868a <=( a7491a  and  a7482a );
 a869a <=( a7473a  and  a7464a );
 a870a <=( a7455a  and  a7446a );
 a871a <=( a7437a  and  a7428a );
 a872a <=( a7419a  and  a7410a );
 a873a <=( a7401a  and  a7392a );
 a874a <=( a7383a  and  a7374a );
 a875a <=( a7365a  and  a7356a );
 a876a <=( a7347a  and  a7338a );
 a877a <=( a7329a  and  a7320a );
 a878a <=( a7311a  and  a7302a );
 a879a <=( a7293a  and  a7284a );
 a880a <=( a7275a  and  a7266a );
 a881a <=( a7257a  and  a7248a );
 a882a <=( a7239a  and  a7230a );
 a883a <=( a7221a  and  a7212a );
 a884a <=( a7203a  and  a7194a );
 a885a <=( a7185a  and  a7176a );
 a886a <=( a7167a  and  a7158a );
 a887a <=( a7149a  and  a7140a );
 a888a <=( a7131a  and  a7122a );
 a889a <=( a7113a  and  a7104a );
 a890a <=( a7095a  and  a7086a );
 a891a <=( a7077a  and  a7068a );
 a892a <=( a7059a  and  a7050a );
 a893a <=( a7041a  and  a7032a );
 a894a <=( a7023a  and  a7014a );
 a895a <=( a7005a  and  a6996a );
 a896a <=( a6987a  and  a6978a );
 a897a <=( a6969a  and  a6960a );
 a898a <=( a6951a  and  a6942a );
 a899a <=( a6933a  and  a6924a );
 a900a <=( a6915a  and  a6906a );
 a901a <=( a6897a  and  a6888a );
 a902a <=( a6879a  and  a6870a );
 a903a <=( a6861a  and  a6852a );
 a904a <=( a6843a  and  a6834a );
 a905a <=( a6825a  and  a6816a );
 a906a <=( a6807a  and  a6798a );
 a907a <=( a6789a  and  a6780a );
 a908a <=( a6771a  and  a6762a );
 a909a <=( a6753a  and  a6744a );
 a910a <=( a6735a  and  a6726a );
 a911a <=( a6717a  and  a6708a );
 a912a <=( a6699a  and  a6690a );
 a913a <=( a6681a  and  a6672a );
 a914a <=( a6663a  and  a6654a );
 a915a <=( a6645a  and  a6636a );
 a916a <=( a6627a  and  a6618a );
 a917a <=( a6609a  and  a6600a );
 a918a <=( a6591a  and  a6582a );
 a919a <=( a6573a  and  a6564a );
 a920a <=( a6555a  and  a6546a );
 a921a <=( a6537a  and  a6528a );
 a922a <=( a6519a  and  a6510a );
 a923a <=( a6501a  and  a6492a );
 a924a <=( a6483a  and  a6474a );
 a925a <=( a6465a  and  a6456a );
 a926a <=( a6447a  and  a6438a );
 a927a <=( a6429a  and  a6420a );
 a928a <=( a6411a  and  a6402a );
 a929a <=( a6393a  and  a6384a );
 a930a <=( a6375a  and  a6366a );
 a931a <=( a6357a  and  a6348a );
 a932a <=( a6339a  and  a6330a );
 a933a <=( a6321a  and  a6312a );
 a934a <=( a6303a  and  a6294a );
 a935a <=( a6285a  and  a6276a );
 a936a <=( a6267a  and  a6258a );
 a937a <=( a6249a  and  a6240a );
 a938a <=( a6231a  and  a6222a );
 a939a <=( a6213a  and  a6204a );
 a940a <=( a6195a  and  a6186a );
 a941a <=( a6177a  and  a6168a );
 a942a <=( a6159a  and  a6150a );
 a943a <=( a6141a  and  a6132a );
 a944a <=( a6123a  and  a6114a );
 a945a <=( a6105a  and  a6096a );
 a946a <=( a6087a  and  a6078a );
 a947a <=( a6069a  and  a6060a );
 a948a <=( a6051a  and  a6042a );
 a949a <=( a6033a  and  a6024a );
 a950a <=( a6015a  and  a6006a );
 a951a <=( a5997a  and  a5988a );
 a952a <=( a5979a  and  a5970a );
 a953a <=( a5961a  and  a5952a );
 a954a <=( a5943a  and  a5934a );
 a955a <=( a5925a  and  a5916a );
 a956a <=( a5907a  and  a5898a );
 a957a <=( a5889a  and  a5880a );
 a958a <=( a5871a  and  a5862a );
 a959a <=( a5853a  and  a5844a );
 a960a <=( a5835a  and  a5826a );
 a961a <=( a5817a  and  a5808a );
 a962a <=( a5799a  and  a5790a );
 a963a <=( a5781a  and  a5772a );
 a964a <=( a5763a  and  a5754a );
 a965a <=( a5745a  and  a5736a );
 a966a <=( a5727a  and  a5718a );
 a967a <=( a5709a  and  a5700a );
 a968a <=( a5691a  and  a5682a );
 a969a <=( a5673a  and  a5664a );
 a970a <=( a5655a  and  a5646a );
 a971a <=( a5637a  and  a5628a );
 a972a <=( a5619a  and  a5610a );
 a973a <=( a5601a  and  a5592a );
 a974a <=( a5583a  and  a5574a );
 a975a <=( a5565a  and  a5556a );
 a976a <=( a5547a  and  a5538a );
 a977a <=( a5529a  and  a5520a );
 a978a <=( a5511a  and  a5502a );
 a979a <=( a5493a  and  a5484a );
 a980a <=( a5475a  and  a5466a );
 a981a <=( a5457a  and  a5448a );
 a982a <=( a5439a  and  a5430a );
 a983a <=( a5421a  and  a5412a );
 a984a <=( a5403a  and  a5394a );
 a985a <=( a5385a  and  a5376a );
 a986a <=( a5367a  and  a5358a );
 a987a <=( a5349a  and  a5340a );
 a988a <=( a5331a  and  a5322a );
 a989a <=( a5313a  and  a5304a );
 a990a <=( a5295a  and  a5286a );
 a991a <=( a5277a  and  a5268a );
 a992a <=( a5259a  and  a5250a );
 a993a <=( a5241a  and  a5232a );
 a994a <=( a5223a  and  a5214a );
 a995a <=( a5205a  and  a5196a );
 a996a <=( a5187a  and  a5178a );
 a997a <=( a5169a  and  a5160a );
 a998a <=( a5151a  and  a5142a );
 a999a <=( a5133a  and  a5124a );
 a1000a <=( a5115a  and  a5106a );
 a1001a <=( a5097a  and  a5088a );
 a1002a <=( a5079a  and  a5070a );
 a1003a <=( a5061a  and  a5052a );
 a1004a <=( a5043a  and  a5034a );
 a1005a <=( a5025a  and  a5016a );
 a1006a <=( a5007a  and  a4998a );
 a1007a <=( a4989a  and  a4980a );
 a1008a <=( a4973a  and  a4964a );
 a1009a <=( a4957a  and  a4948a );
 a1010a <=( a4941a  and  a4932a );
 a1011a <=( a4925a  and  a4916a );
 a1012a <=( a4909a  and  a4900a );
 a1013a <=( a4893a  and  a4884a );
 a1014a <=( a4877a  and  a4868a );
 a1015a <=( a4861a  and  a4852a );
 a1016a <=( a4845a  and  a4836a );
 a1017a <=( a4829a  and  a4820a );
 a1018a <=( a4813a  and  a4804a );
 a1019a <=( a4797a  and  a4788a );
 a1020a <=( a4781a  and  a4772a );
 a1021a <=( a4765a  and  a4756a );
 a1022a <=( a4749a  and  a4740a );
 a1023a <=( a4733a  and  a4724a );
 a1024a <=( a4717a  and  a4708a );
 a1025a <=( a4701a  and  a4692a );
 a1026a <=( a4685a  and  a4676a );
 a1027a <=( a4669a  and  a4660a );
 a1028a <=( a4653a  and  a4644a );
 a1029a <=( a4637a  and  a4628a );
 a1030a <=( a4621a  and  a4612a );
 a1031a <=( a4605a  and  a4596a );
 a1032a <=( a4589a  and  a4580a );
 a1033a <=( a4573a  and  a4564a );
 a1034a <=( a4557a  and  a4548a );
 a1035a <=( a4541a  and  a4532a );
 a1036a <=( a4525a  and  a4516a );
 a1037a <=( a4509a  and  a4500a );
 a1038a <=( a4493a  and  a4484a );
 a1039a <=( a4477a  and  a4468a );
 a1040a <=( a4461a  and  a4452a );
 a1041a <=( a4445a  and  a4436a );
 a1042a <=( a4429a  and  a4420a );
 a1043a <=( a4413a  and  a4404a );
 a1044a <=( a4397a  and  a4388a );
 a1045a <=( a4381a  and  a4372a );
 a1046a <=( a4365a  and  a4356a );
 a1047a <=( a4349a  and  a4340a );
 a1048a <=( a4333a  and  a4324a );
 a1049a <=( a4317a  and  a4308a );
 a1050a <=( a4301a  and  a4292a );
 a1051a <=( a4285a  and  a4276a );
 a1052a <=( a4269a  and  a4260a );
 a1053a <=( a4253a  and  a4244a );
 a1054a <=( a4237a  and  a4228a );
 a1055a <=( a4221a  and  a4212a );
 a1056a <=( a4205a  and  a4196a );
 a1057a <=( a4189a  and  a4180a );
 a1058a <=( a4173a  and  a4164a );
 a1059a <=( a4157a  and  a4148a );
 a1060a <=( a4141a  and  a4132a );
 a1061a <=( a4125a  and  a4116a );
 a1062a <=( a4109a  and  a4100a );
 a1063a <=( a4093a  and  a4084a );
 a1064a <=( a4077a  and  a4068a );
 a1065a <=( a4061a  and  a4052a );
 a1066a <=( a4045a  and  a4036a );
 a1067a <=( a4029a  and  a4020a );
 a1068a <=( a4013a  and  a4004a );
 a1069a <=( a3997a  and  a3990a );
 a1070a <=( a3983a  and  a3976a );
 a1071a <=( a3969a  and  a3962a );
 a1072a <=( a3955a  and  a3948a );
 a1073a <=( a3941a  and  a3934a );
 a1074a <=( a3927a  and  a3920a );
 a1075a <=( a3913a  and  a3906a );
 a1076a <=( a3899a  and  a3892a );
 a1077a <=( a3885a  and  a3878a );
 a1078a <=( a3871a  and  a3864a );
 a1079a <=( a3857a  and  a3850a );
 a1080a <=( a3843a  and  a3836a );
 a1081a <=( a3829a  and  a3822a );
 a1082a <=( a3815a  and  a3808a );
 a1083a <=( a3801a  and  a3794a );
 a1084a <=( a3787a  and  a3780a );
 a1085a <=( a3773a  and  a3766a );
 a1086a <=( a3759a  and  a3752a );
 a1087a <=( a3745a  and  a3738a );
 a1088a <=( a3731a  and  a3724a );
 a1089a <=( a3717a  and  a3710a );
 a1090a <=( a3703a  and  a3696a );
 a1091a <=( a3689a  and  a3682a );
 a1092a <=( a3675a  and  a3668a );
 a1093a <=( a3661a  and  a3654a );
 a1094a <=( a3647a  and  a3640a );
 a1095a <=( a3633a  and  a3626a );
 a1096a <=( a3619a  and  a3612a );
 a1097a <=( a3605a  and  a3598a );
 a1098a <=( a3591a  and  a3584a );
 a1099a <=( a3577a  and  a3570a );
 a1100a <=( a3563a  and  a3556a );
 a1101a <=( a3549a  and  a3542a );
 a1102a <=( a3535a  and  a3528a );
 a1103a <=( a3521a  and  a3514a );
 a1104a <=( a3507a  and  a3500a );
 a1105a <=( a3493a  and  a3488a );
 a1106a <=( a3483a  and  a3478a );
 a1107a <=( a3473a  and  a3468a );
 a1108a <=( a3463a  and  a3458a );
 a1109a <=( a3453a  and  a3448a );
 a1110a <=( a3443a  and  a3438a );
 a1111a <=( a3433a  and  a3428a );
 a1112a <=( a3423a  and  a3418a );
 a1113a <=( a3413a  and  a3408a );
 a1114a <=( a3403a  and  a3398a );
 a1115a <=( a3393a  and  a3388a );
 a1116a <=( a3383a  and  a3378a );
 a1117a <=( a3373a  and  a3370a );
 a1118a <=( a3367a  and  a3364a );
 a1119a <=( a3361a  and  a3358a );
 a1122a <=( a1118a ) or ( a1119a );
 a1125a <=( a1116a ) or ( a1117a );
 a1126a <=( a1125a ) or ( a1122a );
 a1129a <=( a1114a ) or ( a1115a );
 a1132a <=( a1112a ) or ( a1113a );
 a1133a <=( a1132a ) or ( a1129a );
 a1134a <=( a1133a ) or ( a1126a );
 a1137a <=( a1110a ) or ( a1111a );
 a1140a <=( a1108a ) or ( a1109a );
 a1141a <=( a1140a ) or ( a1137a );
 a1144a <=( a1106a ) or ( a1107a );
 a1148a <=( a1103a ) or ( a1104a );
 a1149a <=( a1105a ) or ( a1148a );
 a1150a <=( a1149a ) or ( a1144a );
 a1151a <=( a1150a ) or ( a1141a );
 a1152a <=( a1151a ) or ( a1134a );
 a1155a <=( a1101a ) or ( a1102a );
 a1158a <=( a1099a ) or ( a1100a );
 a1159a <=( a1158a ) or ( a1155a );
 a1162a <=( a1097a ) or ( a1098a );
 a1165a <=( a1095a ) or ( a1096a );
 a1166a <=( a1165a ) or ( a1162a );
 a1167a <=( a1166a ) or ( a1159a );
 a1170a <=( a1093a ) or ( a1094a );
 a1173a <=( a1091a ) or ( a1092a );
 a1174a <=( a1173a ) or ( a1170a );
 a1177a <=( a1089a ) or ( a1090a );
 a1181a <=( a1086a ) or ( a1087a );
 a1182a <=( a1088a ) or ( a1181a );
 a1183a <=( a1182a ) or ( a1177a );
 a1184a <=( a1183a ) or ( a1174a );
 a1185a <=( a1184a ) or ( a1167a );
 a1186a <=( a1185a ) or ( a1152a );
 a1189a <=( a1084a ) or ( a1085a );
 a1192a <=( a1082a ) or ( a1083a );
 a1193a <=( a1192a ) or ( a1189a );
 a1196a <=( a1080a ) or ( a1081a );
 a1199a <=( a1078a ) or ( a1079a );
 a1200a <=( a1199a ) or ( a1196a );
 a1201a <=( a1200a ) or ( a1193a );
 a1204a <=( a1076a ) or ( a1077a );
 a1207a <=( a1074a ) or ( a1075a );
 a1208a <=( a1207a ) or ( a1204a );
 a1211a <=( a1072a ) or ( a1073a );
 a1215a <=( a1069a ) or ( a1070a );
 a1216a <=( a1071a ) or ( a1215a );
 a1217a <=( a1216a ) or ( a1211a );
 a1218a <=( a1217a ) or ( a1208a );
 a1219a <=( a1218a ) or ( a1201a );
 a1222a <=( a1067a ) or ( a1068a );
 a1225a <=( a1065a ) or ( a1066a );
 a1226a <=( a1225a ) or ( a1222a );
 a1229a <=( a1063a ) or ( a1064a );
 a1233a <=( a1060a ) or ( a1061a );
 a1234a <=( a1062a ) or ( a1233a );
 a1235a <=( a1234a ) or ( a1229a );
 a1236a <=( a1235a ) or ( a1226a );
 a1239a <=( a1058a ) or ( a1059a );
 a1242a <=( a1056a ) or ( a1057a );
 a1243a <=( a1242a ) or ( a1239a );
 a1246a <=( a1054a ) or ( a1055a );
 a1250a <=( a1051a ) or ( a1052a );
 a1251a <=( a1053a ) or ( a1250a );
 a1252a <=( a1251a ) or ( a1246a );
 a1253a <=( a1252a ) or ( a1243a );
 a1254a <=( a1253a ) or ( a1236a );
 a1255a <=( a1254a ) or ( a1219a );
 a1256a <=( a1255a ) or ( a1186a );
 a1259a <=( a1049a ) or ( a1050a );
 a1262a <=( a1047a ) or ( a1048a );
 a1263a <=( a1262a ) or ( a1259a );
 a1266a <=( a1045a ) or ( a1046a );
 a1269a <=( a1043a ) or ( a1044a );
 a1270a <=( a1269a ) or ( a1266a );
 a1271a <=( a1270a ) or ( a1263a );
 a1274a <=( a1041a ) or ( a1042a );
 a1277a <=( a1039a ) or ( a1040a );
 a1278a <=( a1277a ) or ( a1274a );
 a1281a <=( a1037a ) or ( a1038a );
 a1285a <=( a1034a ) or ( a1035a );
 a1286a <=( a1036a ) or ( a1285a );
 a1287a <=( a1286a ) or ( a1281a );
 a1288a <=( a1287a ) or ( a1278a );
 a1289a <=( a1288a ) or ( a1271a );
 a1292a <=( a1032a ) or ( a1033a );
 a1295a <=( a1030a ) or ( a1031a );
 a1296a <=( a1295a ) or ( a1292a );
 a1299a <=( a1028a ) or ( a1029a );
 a1303a <=( a1025a ) or ( a1026a );
 a1304a <=( a1027a ) or ( a1303a );
 a1305a <=( a1304a ) or ( a1299a );
 a1306a <=( a1305a ) or ( a1296a );
 a1309a <=( a1023a ) or ( a1024a );
 a1312a <=( a1021a ) or ( a1022a );
 a1313a <=( a1312a ) or ( a1309a );
 a1316a <=( a1019a ) or ( a1020a );
 a1320a <=( a1016a ) or ( a1017a );
 a1321a <=( a1018a ) or ( a1320a );
 a1322a <=( a1321a ) or ( a1316a );
 a1323a <=( a1322a ) or ( a1313a );
 a1324a <=( a1323a ) or ( a1306a );
 a1325a <=( a1324a ) or ( a1289a );
 a1328a <=( a1014a ) or ( a1015a );
 a1331a <=( a1012a ) or ( a1013a );
 a1332a <=( a1331a ) or ( a1328a );
 a1335a <=( a1010a ) or ( a1011a );
 a1338a <=( a1008a ) or ( a1009a );
 a1339a <=( a1338a ) or ( a1335a );
 a1340a <=( a1339a ) or ( a1332a );
 a1343a <=( a1006a ) or ( a1007a );
 a1346a <=( a1004a ) or ( a1005a );
 a1347a <=( a1346a ) or ( a1343a );
 a1350a <=( a1002a ) or ( a1003a );
 a1354a <=( a999a ) or ( a1000a );
 a1355a <=( a1001a ) or ( a1354a );
 a1356a <=( a1355a ) or ( a1350a );
 a1357a <=( a1356a ) or ( a1347a );
 a1358a <=( a1357a ) or ( a1340a );
 a1361a <=( a997a ) or ( a998a );
 a1364a <=( a995a ) or ( a996a );
 a1365a <=( a1364a ) or ( a1361a );
 a1368a <=( a993a ) or ( a994a );
 a1372a <=( a990a ) or ( a991a );
 a1373a <=( a992a ) or ( a1372a );
 a1374a <=( a1373a ) or ( a1368a );
 a1375a <=( a1374a ) or ( a1365a );
 a1378a <=( a988a ) or ( a989a );
 a1381a <=( a986a ) or ( a987a );
 a1382a <=( a1381a ) or ( a1378a );
 a1385a <=( a984a ) or ( a985a );
 a1389a <=( a981a ) or ( a982a );
 a1390a <=( a983a ) or ( a1389a );
 a1391a <=( a1390a ) or ( a1385a );
 a1392a <=( a1391a ) or ( a1382a );
 a1393a <=( a1392a ) or ( a1375a );
 a1394a <=( a1393a ) or ( a1358a );
 a1395a <=( a1394a ) or ( a1325a );
 a1396a <=( a1395a ) or ( a1256a );
 a1399a <=( a979a ) or ( a980a );
 a1402a <=( a977a ) or ( a978a );
 a1403a <=( a1402a ) or ( a1399a );
 a1406a <=( a975a ) or ( a976a );
 a1409a <=( a973a ) or ( a974a );
 a1410a <=( a1409a ) or ( a1406a );
 a1411a <=( a1410a ) or ( a1403a );
 a1414a <=( a971a ) or ( a972a );
 a1417a <=( a969a ) or ( a970a );
 a1418a <=( a1417a ) or ( a1414a );
 a1421a <=( a967a ) or ( a968a );
 a1425a <=( a964a ) or ( a965a );
 a1426a <=( a966a ) or ( a1425a );
 a1427a <=( a1426a ) or ( a1421a );
 a1428a <=( a1427a ) or ( a1418a );
 a1429a <=( a1428a ) or ( a1411a );
 a1432a <=( a962a ) or ( a963a );
 a1435a <=( a960a ) or ( a961a );
 a1436a <=( a1435a ) or ( a1432a );
 a1439a <=( a958a ) or ( a959a );
 a1443a <=( a955a ) or ( a956a );
 a1444a <=( a957a ) or ( a1443a );
 a1445a <=( a1444a ) or ( a1439a );
 a1446a <=( a1445a ) or ( a1436a );
 a1449a <=( a953a ) or ( a954a );
 a1452a <=( a951a ) or ( a952a );
 a1453a <=( a1452a ) or ( a1449a );
 a1456a <=( a949a ) or ( a950a );
 a1460a <=( a946a ) or ( a947a );
 a1461a <=( a948a ) or ( a1460a );
 a1462a <=( a1461a ) or ( a1456a );
 a1463a <=( a1462a ) or ( a1453a );
 a1464a <=( a1463a ) or ( a1446a );
 a1465a <=( a1464a ) or ( a1429a );
 a1468a <=( a944a ) or ( a945a );
 a1471a <=( a942a ) or ( a943a );
 a1472a <=( a1471a ) or ( a1468a );
 a1475a <=( a940a ) or ( a941a );
 a1478a <=( a938a ) or ( a939a );
 a1479a <=( a1478a ) or ( a1475a );
 a1480a <=( a1479a ) or ( a1472a );
 a1483a <=( a936a ) or ( a937a );
 a1486a <=( a934a ) or ( a935a );
 a1487a <=( a1486a ) or ( a1483a );
 a1490a <=( a932a ) or ( a933a );
 a1494a <=( a929a ) or ( a930a );
 a1495a <=( a931a ) or ( a1494a );
 a1496a <=( a1495a ) or ( a1490a );
 a1497a <=( a1496a ) or ( a1487a );
 a1498a <=( a1497a ) or ( a1480a );
 a1501a <=( a927a ) or ( a928a );
 a1504a <=( a925a ) or ( a926a );
 a1505a <=( a1504a ) or ( a1501a );
 a1508a <=( a923a ) or ( a924a );
 a1512a <=( a920a ) or ( a921a );
 a1513a <=( a922a ) or ( a1512a );
 a1514a <=( a1513a ) or ( a1508a );
 a1515a <=( a1514a ) or ( a1505a );
 a1518a <=( a918a ) or ( a919a );
 a1521a <=( a916a ) or ( a917a );
 a1522a <=( a1521a ) or ( a1518a );
 a1525a <=( a914a ) or ( a915a );
 a1529a <=( a911a ) or ( a912a );
 a1530a <=( a913a ) or ( a1529a );
 a1531a <=( a1530a ) or ( a1525a );
 a1532a <=( a1531a ) or ( a1522a );
 a1533a <=( a1532a ) or ( a1515a );
 a1534a <=( a1533a ) or ( a1498a );
 a1535a <=( a1534a ) or ( a1465a );
 a1538a <=( a909a ) or ( a910a );
 a1541a <=( a907a ) or ( a908a );
 a1542a <=( a1541a ) or ( a1538a );
 a1545a <=( a905a ) or ( a906a );
 a1548a <=( a903a ) or ( a904a );
 a1549a <=( a1548a ) or ( a1545a );
 a1550a <=( a1549a ) or ( a1542a );
 a1553a <=( a901a ) or ( a902a );
 a1556a <=( a899a ) or ( a900a );
 a1557a <=( a1556a ) or ( a1553a );
 a1560a <=( a897a ) or ( a898a );
 a1564a <=( a894a ) or ( a895a );
 a1565a <=( a896a ) or ( a1564a );
 a1566a <=( a1565a ) or ( a1560a );
 a1567a <=( a1566a ) or ( a1557a );
 a1568a <=( a1567a ) or ( a1550a );
 a1571a <=( a892a ) or ( a893a );
 a1574a <=( a890a ) or ( a891a );
 a1575a <=( a1574a ) or ( a1571a );
 a1578a <=( a888a ) or ( a889a );
 a1582a <=( a885a ) or ( a886a );
 a1583a <=( a887a ) or ( a1582a );
 a1584a <=( a1583a ) or ( a1578a );
 a1585a <=( a1584a ) or ( a1575a );
 a1588a <=( a883a ) or ( a884a );
 a1591a <=( a881a ) or ( a882a );
 a1592a <=( a1591a ) or ( a1588a );
 a1595a <=( a879a ) or ( a880a );
 a1599a <=( a876a ) or ( a877a );
 a1600a <=( a878a ) or ( a1599a );
 a1601a <=( a1600a ) or ( a1595a );
 a1602a <=( a1601a ) or ( a1592a );
 a1603a <=( a1602a ) or ( a1585a );
 a1604a <=( a1603a ) or ( a1568a );
 a1607a <=( a874a ) or ( a875a );
 a1610a <=( a872a ) or ( a873a );
 a1611a <=( a1610a ) or ( a1607a );
 a1614a <=( a870a ) or ( a871a );
 a1617a <=( a868a ) or ( a869a );
 a1618a <=( a1617a ) or ( a1614a );
 a1619a <=( a1618a ) or ( a1611a );
 a1622a <=( a866a ) or ( a867a );
 a1625a <=( a864a ) or ( a865a );
 a1626a <=( a1625a ) or ( a1622a );
 a1629a <=( a862a ) or ( a863a );
 a1633a <=( a859a ) or ( a860a );
 a1634a <=( a861a ) or ( a1633a );
 a1635a <=( a1634a ) or ( a1629a );
 a1636a <=( a1635a ) or ( a1626a );
 a1637a <=( a1636a ) or ( a1619a );
 a1640a <=( a857a ) or ( a858a );
 a1643a <=( a855a ) or ( a856a );
 a1644a <=( a1643a ) or ( a1640a );
 a1647a <=( a853a ) or ( a854a );
 a1651a <=( a850a ) or ( a851a );
 a1652a <=( a852a ) or ( a1651a );
 a1653a <=( a1652a ) or ( a1647a );
 a1654a <=( a1653a ) or ( a1644a );
 a1657a <=( a848a ) or ( a849a );
 a1660a <=( a846a ) or ( a847a );
 a1661a <=( a1660a ) or ( a1657a );
 a1664a <=( a844a ) or ( a845a );
 a1668a <=( a841a ) or ( a842a );
 a1669a <=( a843a ) or ( a1668a );
 a1670a <=( a1669a ) or ( a1664a );
 a1671a <=( a1670a ) or ( a1661a );
 a1672a <=( a1671a ) or ( a1654a );
 a1673a <=( a1672a ) or ( a1637a );
 a1674a <=( a1673a ) or ( a1604a );
 a1675a <=( a1674a ) or ( a1535a );
 a1676a <=( a1675a ) or ( a1396a );
 a1679a <=( a839a ) or ( a840a );
 a1682a <=( a837a ) or ( a838a );
 a1683a <=( a1682a ) or ( a1679a );
 a1686a <=( a835a ) or ( a836a );
 a1689a <=( a833a ) or ( a834a );
 a1690a <=( a1689a ) or ( a1686a );
 a1691a <=( a1690a ) or ( a1683a );
 a1694a <=( a831a ) or ( a832a );
 a1697a <=( a829a ) or ( a830a );
 a1698a <=( a1697a ) or ( a1694a );
 a1701a <=( a827a ) or ( a828a );
 a1705a <=( a824a ) or ( a825a );
 a1706a <=( a826a ) or ( a1705a );
 a1707a <=( a1706a ) or ( a1701a );
 a1708a <=( a1707a ) or ( a1698a );
 a1709a <=( a1708a ) or ( a1691a );
 a1712a <=( a822a ) or ( a823a );
 a1715a <=( a820a ) or ( a821a );
 a1716a <=( a1715a ) or ( a1712a );
 a1719a <=( a818a ) or ( a819a );
 a1723a <=( a815a ) or ( a816a );
 a1724a <=( a817a ) or ( a1723a );
 a1725a <=( a1724a ) or ( a1719a );
 a1726a <=( a1725a ) or ( a1716a );
 a1729a <=( a813a ) or ( a814a );
 a1732a <=( a811a ) or ( a812a );
 a1733a <=( a1732a ) or ( a1729a );
 a1736a <=( a809a ) or ( a810a );
 a1740a <=( a806a ) or ( a807a );
 a1741a <=( a808a ) or ( a1740a );
 a1742a <=( a1741a ) or ( a1736a );
 a1743a <=( a1742a ) or ( a1733a );
 a1744a <=( a1743a ) or ( a1726a );
 a1745a <=( a1744a ) or ( a1709a );
 a1748a <=( a804a ) or ( a805a );
 a1751a <=( a802a ) or ( a803a );
 a1752a <=( a1751a ) or ( a1748a );
 a1755a <=( a800a ) or ( a801a );
 a1758a <=( a798a ) or ( a799a );
 a1759a <=( a1758a ) or ( a1755a );
 a1760a <=( a1759a ) or ( a1752a );
 a1763a <=( a796a ) or ( a797a );
 a1766a <=( a794a ) or ( a795a );
 a1767a <=( a1766a ) or ( a1763a );
 a1770a <=( a792a ) or ( a793a );
 a1774a <=( a789a ) or ( a790a );
 a1775a <=( a791a ) or ( a1774a );
 a1776a <=( a1775a ) or ( a1770a );
 a1777a <=( a1776a ) or ( a1767a );
 a1778a <=( a1777a ) or ( a1760a );
 a1781a <=( a787a ) or ( a788a );
 a1784a <=( a785a ) or ( a786a );
 a1785a <=( a1784a ) or ( a1781a );
 a1788a <=( a783a ) or ( a784a );
 a1792a <=( a780a ) or ( a781a );
 a1793a <=( a782a ) or ( a1792a );
 a1794a <=( a1793a ) or ( a1788a );
 a1795a <=( a1794a ) or ( a1785a );
 a1798a <=( a778a ) or ( a779a );
 a1801a <=( a776a ) or ( a777a );
 a1802a <=( a1801a ) or ( a1798a );
 a1805a <=( a774a ) or ( a775a );
 a1809a <=( a771a ) or ( a772a );
 a1810a <=( a773a ) or ( a1809a );
 a1811a <=( a1810a ) or ( a1805a );
 a1812a <=( a1811a ) or ( a1802a );
 a1813a <=( a1812a ) or ( a1795a );
 a1814a <=( a1813a ) or ( a1778a );
 a1815a <=( a1814a ) or ( a1745a );
 a1818a <=( a769a ) or ( a770a );
 a1821a <=( a767a ) or ( a768a );
 a1822a <=( a1821a ) or ( a1818a );
 a1825a <=( a765a ) or ( a766a );
 a1828a <=( a763a ) or ( a764a );
 a1829a <=( a1828a ) or ( a1825a );
 a1830a <=( a1829a ) or ( a1822a );
 a1833a <=( a761a ) or ( a762a );
 a1836a <=( a759a ) or ( a760a );
 a1837a <=( a1836a ) or ( a1833a );
 a1840a <=( a757a ) or ( a758a );
 a1844a <=( a754a ) or ( a755a );
 a1845a <=( a756a ) or ( a1844a );
 a1846a <=( a1845a ) or ( a1840a );
 a1847a <=( a1846a ) or ( a1837a );
 a1848a <=( a1847a ) or ( a1830a );
 a1851a <=( a752a ) or ( a753a );
 a1854a <=( a750a ) or ( a751a );
 a1855a <=( a1854a ) or ( a1851a );
 a1858a <=( a748a ) or ( a749a );
 a1862a <=( a745a ) or ( a746a );
 a1863a <=( a747a ) or ( a1862a );
 a1864a <=( a1863a ) or ( a1858a );
 a1865a <=( a1864a ) or ( a1855a );
 a1868a <=( a743a ) or ( a744a );
 a1871a <=( a741a ) or ( a742a );
 a1872a <=( a1871a ) or ( a1868a );
 a1875a <=( a739a ) or ( a740a );
 a1879a <=( a736a ) or ( a737a );
 a1880a <=( a738a ) or ( a1879a );
 a1881a <=( a1880a ) or ( a1875a );
 a1882a <=( a1881a ) or ( a1872a );
 a1883a <=( a1882a ) or ( a1865a );
 a1884a <=( a1883a ) or ( a1848a );
 a1887a <=( a734a ) or ( a735a );
 a1890a <=( a732a ) or ( a733a );
 a1891a <=( a1890a ) or ( a1887a );
 a1894a <=( a730a ) or ( a731a );
 a1897a <=( a728a ) or ( a729a );
 a1898a <=( a1897a ) or ( a1894a );
 a1899a <=( a1898a ) or ( a1891a );
 a1902a <=( a726a ) or ( a727a );
 a1905a <=( a724a ) or ( a725a );
 a1906a <=( a1905a ) or ( a1902a );
 a1909a <=( a722a ) or ( a723a );
 a1913a <=( a719a ) or ( a720a );
 a1914a <=( a721a ) or ( a1913a );
 a1915a <=( a1914a ) or ( a1909a );
 a1916a <=( a1915a ) or ( a1906a );
 a1917a <=( a1916a ) or ( a1899a );
 a1920a <=( a717a ) or ( a718a );
 a1923a <=( a715a ) or ( a716a );
 a1924a <=( a1923a ) or ( a1920a );
 a1927a <=( a713a ) or ( a714a );
 a1931a <=( a710a ) or ( a711a );
 a1932a <=( a712a ) or ( a1931a );
 a1933a <=( a1932a ) or ( a1927a );
 a1934a <=( a1933a ) or ( a1924a );
 a1937a <=( a708a ) or ( a709a );
 a1940a <=( a706a ) or ( a707a );
 a1941a <=( a1940a ) or ( a1937a );
 a1944a <=( a704a ) or ( a705a );
 a1948a <=( a701a ) or ( a702a );
 a1949a <=( a703a ) or ( a1948a );
 a1950a <=( a1949a ) or ( a1944a );
 a1951a <=( a1950a ) or ( a1941a );
 a1952a <=( a1951a ) or ( a1934a );
 a1953a <=( a1952a ) or ( a1917a );
 a1954a <=( a1953a ) or ( a1884a );
 a1955a <=( a1954a ) or ( a1815a );
 a1958a <=( a699a ) or ( a700a );
 a1961a <=( a697a ) or ( a698a );
 a1962a <=( a1961a ) or ( a1958a );
 a1965a <=( a695a ) or ( a696a );
 a1968a <=( a693a ) or ( a694a );
 a1969a <=( a1968a ) or ( a1965a );
 a1970a <=( a1969a ) or ( a1962a );
 a1973a <=( a691a ) or ( a692a );
 a1976a <=( a689a ) or ( a690a );
 a1977a <=( a1976a ) or ( a1973a );
 a1980a <=( a687a ) or ( a688a );
 a1984a <=( a684a ) or ( a685a );
 a1985a <=( a686a ) or ( a1984a );
 a1986a <=( a1985a ) or ( a1980a );
 a1987a <=( a1986a ) or ( a1977a );
 a1988a <=( a1987a ) or ( a1970a );
 a1991a <=( a682a ) or ( a683a );
 a1994a <=( a680a ) or ( a681a );
 a1995a <=( a1994a ) or ( a1991a );
 a1998a <=( a678a ) or ( a679a );
 a2002a <=( a675a ) or ( a676a );
 a2003a <=( a677a ) or ( a2002a );
 a2004a <=( a2003a ) or ( a1998a );
 a2005a <=( a2004a ) or ( a1995a );
 a2008a <=( a673a ) or ( a674a );
 a2011a <=( a671a ) or ( a672a );
 a2012a <=( a2011a ) or ( a2008a );
 a2015a <=( a669a ) or ( a670a );
 a2019a <=( a666a ) or ( a667a );
 a2020a <=( a668a ) or ( a2019a );
 a2021a <=( a2020a ) or ( a2015a );
 a2022a <=( a2021a ) or ( a2012a );
 a2023a <=( a2022a ) or ( a2005a );
 a2024a <=( a2023a ) or ( a1988a );
 a2027a <=( a664a ) or ( a665a );
 a2030a <=( a662a ) or ( a663a );
 a2031a <=( a2030a ) or ( a2027a );
 a2034a <=( a660a ) or ( a661a );
 a2037a <=( a658a ) or ( a659a );
 a2038a <=( a2037a ) or ( a2034a );
 a2039a <=( a2038a ) or ( a2031a );
 a2042a <=( a656a ) or ( a657a );
 a2045a <=( a654a ) or ( a655a );
 a2046a <=( a2045a ) or ( a2042a );
 a2049a <=( a652a ) or ( a653a );
 a2053a <=( a649a ) or ( a650a );
 a2054a <=( a651a ) or ( a2053a );
 a2055a <=( a2054a ) or ( a2049a );
 a2056a <=( a2055a ) or ( a2046a );
 a2057a <=( a2056a ) or ( a2039a );
 a2060a <=( a647a ) or ( a648a );
 a2063a <=( a645a ) or ( a646a );
 a2064a <=( a2063a ) or ( a2060a );
 a2067a <=( a643a ) or ( a644a );
 a2071a <=( a640a ) or ( a641a );
 a2072a <=( a642a ) or ( a2071a );
 a2073a <=( a2072a ) or ( a2067a );
 a2074a <=( a2073a ) or ( a2064a );
 a2077a <=( a638a ) or ( a639a );
 a2080a <=( a636a ) or ( a637a );
 a2081a <=( a2080a ) or ( a2077a );
 a2084a <=( a634a ) or ( a635a );
 a2088a <=( a631a ) or ( a632a );
 a2089a <=( a633a ) or ( a2088a );
 a2090a <=( a2089a ) or ( a2084a );
 a2091a <=( a2090a ) or ( a2081a );
 a2092a <=( a2091a ) or ( a2074a );
 a2093a <=( a2092a ) or ( a2057a );
 a2094a <=( a2093a ) or ( a2024a );
 a2097a <=( a629a ) or ( a630a );
 a2100a <=( a627a ) or ( a628a );
 a2101a <=( a2100a ) or ( a2097a );
 a2104a <=( a625a ) or ( a626a );
 a2107a <=( a623a ) or ( a624a );
 a2108a <=( a2107a ) or ( a2104a );
 a2109a <=( a2108a ) or ( a2101a );
 a2112a <=( a621a ) or ( a622a );
 a2115a <=( a619a ) or ( a620a );
 a2116a <=( a2115a ) or ( a2112a );
 a2119a <=( a617a ) or ( a618a );
 a2123a <=( a614a ) or ( a615a );
 a2124a <=( a616a ) or ( a2123a );
 a2125a <=( a2124a ) or ( a2119a );
 a2126a <=( a2125a ) or ( a2116a );
 a2127a <=( a2126a ) or ( a2109a );
 a2130a <=( a612a ) or ( a613a );
 a2133a <=( a610a ) or ( a611a );
 a2134a <=( a2133a ) or ( a2130a );
 a2137a <=( a608a ) or ( a609a );
 a2141a <=( a605a ) or ( a606a );
 a2142a <=( a607a ) or ( a2141a );
 a2143a <=( a2142a ) or ( a2137a );
 a2144a <=( a2143a ) or ( a2134a );
 a2147a <=( a603a ) or ( a604a );
 a2150a <=( a601a ) or ( a602a );
 a2151a <=( a2150a ) or ( a2147a );
 a2154a <=( a599a ) or ( a600a );
 a2158a <=( a596a ) or ( a597a );
 a2159a <=( a598a ) or ( a2158a );
 a2160a <=( a2159a ) or ( a2154a );
 a2161a <=( a2160a ) or ( a2151a );
 a2162a <=( a2161a ) or ( a2144a );
 a2163a <=( a2162a ) or ( a2127a );
 a2166a <=( a594a ) or ( a595a );
 a2169a <=( a592a ) or ( a593a );
 a2170a <=( a2169a ) or ( a2166a );
 a2173a <=( a590a ) or ( a591a );
 a2176a <=( a588a ) or ( a589a );
 a2177a <=( a2176a ) or ( a2173a );
 a2178a <=( a2177a ) or ( a2170a );
 a2181a <=( a586a ) or ( a587a );
 a2184a <=( a584a ) or ( a585a );
 a2185a <=( a2184a ) or ( a2181a );
 a2188a <=( a582a ) or ( a583a );
 a2192a <=( a579a ) or ( a580a );
 a2193a <=( a581a ) or ( a2192a );
 a2194a <=( a2193a ) or ( a2188a );
 a2195a <=( a2194a ) or ( a2185a );
 a2196a <=( a2195a ) or ( a2178a );
 a2199a <=( a577a ) or ( a578a );
 a2202a <=( a575a ) or ( a576a );
 a2203a <=( a2202a ) or ( a2199a );
 a2206a <=( a573a ) or ( a574a );
 a2210a <=( a570a ) or ( a571a );
 a2211a <=( a572a ) or ( a2210a );
 a2212a <=( a2211a ) or ( a2206a );
 a2213a <=( a2212a ) or ( a2203a );
 a2216a <=( a568a ) or ( a569a );
 a2219a <=( a566a ) or ( a567a );
 a2220a <=( a2219a ) or ( a2216a );
 a2223a <=( a564a ) or ( a565a );
 a2227a <=( a561a ) or ( a562a );
 a2228a <=( a563a ) or ( a2227a );
 a2229a <=( a2228a ) or ( a2223a );
 a2230a <=( a2229a ) or ( a2220a );
 a2231a <=( a2230a ) or ( a2213a );
 a2232a <=( a2231a ) or ( a2196a );
 a2233a <=( a2232a ) or ( a2163a );
 a2234a <=( a2233a ) or ( a2094a );
 a2235a <=( a2234a ) or ( a1955a );
 a2236a <=( a2235a ) or ( a1676a );
 a2239a <=( a559a ) or ( a560a );
 a2242a <=( a557a ) or ( a558a );
 a2243a <=( a2242a ) or ( a2239a );
 a2246a <=( a555a ) or ( a556a );
 a2249a <=( a553a ) or ( a554a );
 a2250a <=( a2249a ) or ( a2246a );
 a2251a <=( a2250a ) or ( a2243a );
 a2254a <=( a551a ) or ( a552a );
 a2257a <=( a549a ) or ( a550a );
 a2258a <=( a2257a ) or ( a2254a );
 a2261a <=( a547a ) or ( a548a );
 a2265a <=( a544a ) or ( a545a );
 a2266a <=( a546a ) or ( a2265a );
 a2267a <=( a2266a ) or ( a2261a );
 a2268a <=( a2267a ) or ( a2258a );
 a2269a <=( a2268a ) or ( a2251a );
 a2272a <=( a542a ) or ( a543a );
 a2275a <=( a540a ) or ( a541a );
 a2276a <=( a2275a ) or ( a2272a );
 a2279a <=( a538a ) or ( a539a );
 a2283a <=( a535a ) or ( a536a );
 a2284a <=( a537a ) or ( a2283a );
 a2285a <=( a2284a ) or ( a2279a );
 a2286a <=( a2285a ) or ( a2276a );
 a2289a <=( a533a ) or ( a534a );
 a2292a <=( a531a ) or ( a532a );
 a2293a <=( a2292a ) or ( a2289a );
 a2296a <=( a529a ) or ( a530a );
 a2300a <=( a526a ) or ( a527a );
 a2301a <=( a528a ) or ( a2300a );
 a2302a <=( a2301a ) or ( a2296a );
 a2303a <=( a2302a ) or ( a2293a );
 a2304a <=( a2303a ) or ( a2286a );
 a2305a <=( a2304a ) or ( a2269a );
 a2308a <=( a524a ) or ( a525a );
 a2311a <=( a522a ) or ( a523a );
 a2312a <=( a2311a ) or ( a2308a );
 a2315a <=( a520a ) or ( a521a );
 a2318a <=( a518a ) or ( a519a );
 a2319a <=( a2318a ) or ( a2315a );
 a2320a <=( a2319a ) or ( a2312a );
 a2323a <=( a516a ) or ( a517a );
 a2326a <=( a514a ) or ( a515a );
 a2327a <=( a2326a ) or ( a2323a );
 a2330a <=( a512a ) or ( a513a );
 a2334a <=( a509a ) or ( a510a );
 a2335a <=( a511a ) or ( a2334a );
 a2336a <=( a2335a ) or ( a2330a );
 a2337a <=( a2336a ) or ( a2327a );
 a2338a <=( a2337a ) or ( a2320a );
 a2341a <=( a507a ) or ( a508a );
 a2344a <=( a505a ) or ( a506a );
 a2345a <=( a2344a ) or ( a2341a );
 a2348a <=( a503a ) or ( a504a );
 a2352a <=( a500a ) or ( a501a );
 a2353a <=( a502a ) or ( a2352a );
 a2354a <=( a2353a ) or ( a2348a );
 a2355a <=( a2354a ) or ( a2345a );
 a2358a <=( a498a ) or ( a499a );
 a2361a <=( a496a ) or ( a497a );
 a2362a <=( a2361a ) or ( a2358a );
 a2365a <=( a494a ) or ( a495a );
 a2369a <=( a491a ) or ( a492a );
 a2370a <=( a493a ) or ( a2369a );
 a2371a <=( a2370a ) or ( a2365a );
 a2372a <=( a2371a ) or ( a2362a );
 a2373a <=( a2372a ) or ( a2355a );
 a2374a <=( a2373a ) or ( a2338a );
 a2375a <=( a2374a ) or ( a2305a );
 a2378a <=( a489a ) or ( a490a );
 a2381a <=( a487a ) or ( a488a );
 a2382a <=( a2381a ) or ( a2378a );
 a2385a <=( a485a ) or ( a486a );
 a2388a <=( a483a ) or ( a484a );
 a2389a <=( a2388a ) or ( a2385a );
 a2390a <=( a2389a ) or ( a2382a );
 a2393a <=( a481a ) or ( a482a );
 a2396a <=( a479a ) or ( a480a );
 a2397a <=( a2396a ) or ( a2393a );
 a2400a <=( a477a ) or ( a478a );
 a2404a <=( a474a ) or ( a475a );
 a2405a <=( a476a ) or ( a2404a );
 a2406a <=( a2405a ) or ( a2400a );
 a2407a <=( a2406a ) or ( a2397a );
 a2408a <=( a2407a ) or ( a2390a );
 a2411a <=( a472a ) or ( a473a );
 a2414a <=( a470a ) or ( a471a );
 a2415a <=( a2414a ) or ( a2411a );
 a2418a <=( a468a ) or ( a469a );
 a2422a <=( a465a ) or ( a466a );
 a2423a <=( a467a ) or ( a2422a );
 a2424a <=( a2423a ) or ( a2418a );
 a2425a <=( a2424a ) or ( a2415a );
 a2428a <=( a463a ) or ( a464a );
 a2431a <=( a461a ) or ( a462a );
 a2432a <=( a2431a ) or ( a2428a );
 a2435a <=( a459a ) or ( a460a );
 a2439a <=( a456a ) or ( a457a );
 a2440a <=( a458a ) or ( a2439a );
 a2441a <=( a2440a ) or ( a2435a );
 a2442a <=( a2441a ) or ( a2432a );
 a2443a <=( a2442a ) or ( a2425a );
 a2444a <=( a2443a ) or ( a2408a );
 a2447a <=( a454a ) or ( a455a );
 a2450a <=( a452a ) or ( a453a );
 a2451a <=( a2450a ) or ( a2447a );
 a2454a <=( a450a ) or ( a451a );
 a2457a <=( a448a ) or ( a449a );
 a2458a <=( a2457a ) or ( a2454a );
 a2459a <=( a2458a ) or ( a2451a );
 a2462a <=( a446a ) or ( a447a );
 a2465a <=( a444a ) or ( a445a );
 a2466a <=( a2465a ) or ( a2462a );
 a2469a <=( a442a ) or ( a443a );
 a2473a <=( a439a ) or ( a440a );
 a2474a <=( a441a ) or ( a2473a );
 a2475a <=( a2474a ) or ( a2469a );
 a2476a <=( a2475a ) or ( a2466a );
 a2477a <=( a2476a ) or ( a2459a );
 a2480a <=( a437a ) or ( a438a );
 a2483a <=( a435a ) or ( a436a );
 a2484a <=( a2483a ) or ( a2480a );
 a2487a <=( a433a ) or ( a434a );
 a2491a <=( a430a ) or ( a431a );
 a2492a <=( a432a ) or ( a2491a );
 a2493a <=( a2492a ) or ( a2487a );
 a2494a <=( a2493a ) or ( a2484a );
 a2497a <=( a428a ) or ( a429a );
 a2500a <=( a426a ) or ( a427a );
 a2501a <=( a2500a ) or ( a2497a );
 a2504a <=( a424a ) or ( a425a );
 a2508a <=( a421a ) or ( a422a );
 a2509a <=( a423a ) or ( a2508a );
 a2510a <=( a2509a ) or ( a2504a );
 a2511a <=( a2510a ) or ( a2501a );
 a2512a <=( a2511a ) or ( a2494a );
 a2513a <=( a2512a ) or ( a2477a );
 a2514a <=( a2513a ) or ( a2444a );
 a2515a <=( a2514a ) or ( a2375a );
 a2518a <=( a419a ) or ( a420a );
 a2521a <=( a417a ) or ( a418a );
 a2522a <=( a2521a ) or ( a2518a );
 a2525a <=( a415a ) or ( a416a );
 a2528a <=( a413a ) or ( a414a );
 a2529a <=( a2528a ) or ( a2525a );
 a2530a <=( a2529a ) or ( a2522a );
 a2533a <=( a411a ) or ( a412a );
 a2536a <=( a409a ) or ( a410a );
 a2537a <=( a2536a ) or ( a2533a );
 a2540a <=( a407a ) or ( a408a );
 a2544a <=( a404a ) or ( a405a );
 a2545a <=( a406a ) or ( a2544a );
 a2546a <=( a2545a ) or ( a2540a );
 a2547a <=( a2546a ) or ( a2537a );
 a2548a <=( a2547a ) or ( a2530a );
 a2551a <=( a402a ) or ( a403a );
 a2554a <=( a400a ) or ( a401a );
 a2555a <=( a2554a ) or ( a2551a );
 a2558a <=( a398a ) or ( a399a );
 a2562a <=( a395a ) or ( a396a );
 a2563a <=( a397a ) or ( a2562a );
 a2564a <=( a2563a ) or ( a2558a );
 a2565a <=( a2564a ) or ( a2555a );
 a2568a <=( a393a ) or ( a394a );
 a2571a <=( a391a ) or ( a392a );
 a2572a <=( a2571a ) or ( a2568a );
 a2575a <=( a389a ) or ( a390a );
 a2579a <=( a386a ) or ( a387a );
 a2580a <=( a388a ) or ( a2579a );
 a2581a <=( a2580a ) or ( a2575a );
 a2582a <=( a2581a ) or ( a2572a );
 a2583a <=( a2582a ) or ( a2565a );
 a2584a <=( a2583a ) or ( a2548a );
 a2587a <=( a384a ) or ( a385a );
 a2590a <=( a382a ) or ( a383a );
 a2591a <=( a2590a ) or ( a2587a );
 a2594a <=( a380a ) or ( a381a );
 a2597a <=( a378a ) or ( a379a );
 a2598a <=( a2597a ) or ( a2594a );
 a2599a <=( a2598a ) or ( a2591a );
 a2602a <=( a376a ) or ( a377a );
 a2605a <=( a374a ) or ( a375a );
 a2606a <=( a2605a ) or ( a2602a );
 a2609a <=( a372a ) or ( a373a );
 a2613a <=( a369a ) or ( a370a );
 a2614a <=( a371a ) or ( a2613a );
 a2615a <=( a2614a ) or ( a2609a );
 a2616a <=( a2615a ) or ( a2606a );
 a2617a <=( a2616a ) or ( a2599a );
 a2620a <=( a367a ) or ( a368a );
 a2623a <=( a365a ) or ( a366a );
 a2624a <=( a2623a ) or ( a2620a );
 a2627a <=( a363a ) or ( a364a );
 a2631a <=( a360a ) or ( a361a );
 a2632a <=( a362a ) or ( a2631a );
 a2633a <=( a2632a ) or ( a2627a );
 a2634a <=( a2633a ) or ( a2624a );
 a2637a <=( a358a ) or ( a359a );
 a2640a <=( a356a ) or ( a357a );
 a2641a <=( a2640a ) or ( a2637a );
 a2644a <=( a354a ) or ( a355a );
 a2648a <=( a351a ) or ( a352a );
 a2649a <=( a353a ) or ( a2648a );
 a2650a <=( a2649a ) or ( a2644a );
 a2651a <=( a2650a ) or ( a2641a );
 a2652a <=( a2651a ) or ( a2634a );
 a2653a <=( a2652a ) or ( a2617a );
 a2654a <=( a2653a ) or ( a2584a );
 a2657a <=( a349a ) or ( a350a );
 a2660a <=( a347a ) or ( a348a );
 a2661a <=( a2660a ) or ( a2657a );
 a2664a <=( a345a ) or ( a346a );
 a2667a <=( a343a ) or ( a344a );
 a2668a <=( a2667a ) or ( a2664a );
 a2669a <=( a2668a ) or ( a2661a );
 a2672a <=( a341a ) or ( a342a );
 a2675a <=( a339a ) or ( a340a );
 a2676a <=( a2675a ) or ( a2672a );
 a2679a <=( a337a ) or ( a338a );
 a2683a <=( a334a ) or ( a335a );
 a2684a <=( a336a ) or ( a2683a );
 a2685a <=( a2684a ) or ( a2679a );
 a2686a <=( a2685a ) or ( a2676a );
 a2687a <=( a2686a ) or ( a2669a );
 a2690a <=( a332a ) or ( a333a );
 a2693a <=( a330a ) or ( a331a );
 a2694a <=( a2693a ) or ( a2690a );
 a2697a <=( a328a ) or ( a329a );
 a2701a <=( a325a ) or ( a326a );
 a2702a <=( a327a ) or ( a2701a );
 a2703a <=( a2702a ) or ( a2697a );
 a2704a <=( a2703a ) or ( a2694a );
 a2707a <=( a323a ) or ( a324a );
 a2710a <=( a321a ) or ( a322a );
 a2711a <=( a2710a ) or ( a2707a );
 a2714a <=( a319a ) or ( a320a );
 a2718a <=( a316a ) or ( a317a );
 a2719a <=( a318a ) or ( a2718a );
 a2720a <=( a2719a ) or ( a2714a );
 a2721a <=( a2720a ) or ( a2711a );
 a2722a <=( a2721a ) or ( a2704a );
 a2723a <=( a2722a ) or ( a2687a );
 a2726a <=( a314a ) or ( a315a );
 a2729a <=( a312a ) or ( a313a );
 a2730a <=( a2729a ) or ( a2726a );
 a2733a <=( a310a ) or ( a311a );
 a2736a <=( a308a ) or ( a309a );
 a2737a <=( a2736a ) or ( a2733a );
 a2738a <=( a2737a ) or ( a2730a );
 a2741a <=( a306a ) or ( a307a );
 a2744a <=( a304a ) or ( a305a );
 a2745a <=( a2744a ) or ( a2741a );
 a2748a <=( a302a ) or ( a303a );
 a2752a <=( a299a ) or ( a300a );
 a2753a <=( a301a ) or ( a2752a );
 a2754a <=( a2753a ) or ( a2748a );
 a2755a <=( a2754a ) or ( a2745a );
 a2756a <=( a2755a ) or ( a2738a );
 a2759a <=( a297a ) or ( a298a );
 a2762a <=( a295a ) or ( a296a );
 a2763a <=( a2762a ) or ( a2759a );
 a2766a <=( a293a ) or ( a294a );
 a2770a <=( a290a ) or ( a291a );
 a2771a <=( a292a ) or ( a2770a );
 a2772a <=( a2771a ) or ( a2766a );
 a2773a <=( a2772a ) or ( a2763a );
 a2776a <=( a288a ) or ( a289a );
 a2779a <=( a286a ) or ( a287a );
 a2780a <=( a2779a ) or ( a2776a );
 a2783a <=( a284a ) or ( a285a );
 a2787a <=( a281a ) or ( a282a );
 a2788a <=( a283a ) or ( a2787a );
 a2789a <=( a2788a ) or ( a2783a );
 a2790a <=( a2789a ) or ( a2780a );
 a2791a <=( a2790a ) or ( a2773a );
 a2792a <=( a2791a ) or ( a2756a );
 a2793a <=( a2792a ) or ( a2723a );
 a2794a <=( a2793a ) or ( a2654a );
 a2795a <=( a2794a ) or ( a2515a );
 a2798a <=( a279a ) or ( a280a );
 a2801a <=( a277a ) or ( a278a );
 a2802a <=( a2801a ) or ( a2798a );
 a2805a <=( a275a ) or ( a276a );
 a2808a <=( a273a ) or ( a274a );
 a2809a <=( a2808a ) or ( a2805a );
 a2810a <=( a2809a ) or ( a2802a );
 a2813a <=( a271a ) or ( a272a );
 a2816a <=( a269a ) or ( a270a );
 a2817a <=( a2816a ) or ( a2813a );
 a2820a <=( a267a ) or ( a268a );
 a2824a <=( a264a ) or ( a265a );
 a2825a <=( a266a ) or ( a2824a );
 a2826a <=( a2825a ) or ( a2820a );
 a2827a <=( a2826a ) or ( a2817a );
 a2828a <=( a2827a ) or ( a2810a );
 a2831a <=( a262a ) or ( a263a );
 a2834a <=( a260a ) or ( a261a );
 a2835a <=( a2834a ) or ( a2831a );
 a2838a <=( a258a ) or ( a259a );
 a2842a <=( a255a ) or ( a256a );
 a2843a <=( a257a ) or ( a2842a );
 a2844a <=( a2843a ) or ( a2838a );
 a2845a <=( a2844a ) or ( a2835a );
 a2848a <=( a253a ) or ( a254a );
 a2851a <=( a251a ) or ( a252a );
 a2852a <=( a2851a ) or ( a2848a );
 a2855a <=( a249a ) or ( a250a );
 a2859a <=( a246a ) or ( a247a );
 a2860a <=( a248a ) or ( a2859a );
 a2861a <=( a2860a ) or ( a2855a );
 a2862a <=( a2861a ) or ( a2852a );
 a2863a <=( a2862a ) or ( a2845a );
 a2864a <=( a2863a ) or ( a2828a );
 a2867a <=( a244a ) or ( a245a );
 a2870a <=( a242a ) or ( a243a );
 a2871a <=( a2870a ) or ( a2867a );
 a2874a <=( a240a ) or ( a241a );
 a2877a <=( a238a ) or ( a239a );
 a2878a <=( a2877a ) or ( a2874a );
 a2879a <=( a2878a ) or ( a2871a );
 a2882a <=( a236a ) or ( a237a );
 a2885a <=( a234a ) or ( a235a );
 a2886a <=( a2885a ) or ( a2882a );
 a2889a <=( a232a ) or ( a233a );
 a2893a <=( a229a ) or ( a230a );
 a2894a <=( a231a ) or ( a2893a );
 a2895a <=( a2894a ) or ( a2889a );
 a2896a <=( a2895a ) or ( a2886a );
 a2897a <=( a2896a ) or ( a2879a );
 a2900a <=( a227a ) or ( a228a );
 a2903a <=( a225a ) or ( a226a );
 a2904a <=( a2903a ) or ( a2900a );
 a2907a <=( a223a ) or ( a224a );
 a2911a <=( a220a ) or ( a221a );
 a2912a <=( a222a ) or ( a2911a );
 a2913a <=( a2912a ) or ( a2907a );
 a2914a <=( a2913a ) or ( a2904a );
 a2917a <=( a218a ) or ( a219a );
 a2920a <=( a216a ) or ( a217a );
 a2921a <=( a2920a ) or ( a2917a );
 a2924a <=( a214a ) or ( a215a );
 a2928a <=( a211a ) or ( a212a );
 a2929a <=( a213a ) or ( a2928a );
 a2930a <=( a2929a ) or ( a2924a );
 a2931a <=( a2930a ) or ( a2921a );
 a2932a <=( a2931a ) or ( a2914a );
 a2933a <=( a2932a ) or ( a2897a );
 a2934a <=( a2933a ) or ( a2864a );
 a2937a <=( a209a ) or ( a210a );
 a2940a <=( a207a ) or ( a208a );
 a2941a <=( a2940a ) or ( a2937a );
 a2944a <=( a205a ) or ( a206a );
 a2947a <=( a203a ) or ( a204a );
 a2948a <=( a2947a ) or ( a2944a );
 a2949a <=( a2948a ) or ( a2941a );
 a2952a <=( a201a ) or ( a202a );
 a2955a <=( a199a ) or ( a200a );
 a2956a <=( a2955a ) or ( a2952a );
 a2959a <=( a197a ) or ( a198a );
 a2963a <=( a194a ) or ( a195a );
 a2964a <=( a196a ) or ( a2963a );
 a2965a <=( a2964a ) or ( a2959a );
 a2966a <=( a2965a ) or ( a2956a );
 a2967a <=( a2966a ) or ( a2949a );
 a2970a <=( a192a ) or ( a193a );
 a2973a <=( a190a ) or ( a191a );
 a2974a <=( a2973a ) or ( a2970a );
 a2977a <=( a188a ) or ( a189a );
 a2981a <=( a185a ) or ( a186a );
 a2982a <=( a187a ) or ( a2981a );
 a2983a <=( a2982a ) or ( a2977a );
 a2984a <=( a2983a ) or ( a2974a );
 a2987a <=( a183a ) or ( a184a );
 a2990a <=( a181a ) or ( a182a );
 a2991a <=( a2990a ) or ( a2987a );
 a2994a <=( a179a ) or ( a180a );
 a2998a <=( a176a ) or ( a177a );
 a2999a <=( a178a ) or ( a2998a );
 a3000a <=( a2999a ) or ( a2994a );
 a3001a <=( a3000a ) or ( a2991a );
 a3002a <=( a3001a ) or ( a2984a );
 a3003a <=( a3002a ) or ( a2967a );
 a3006a <=( a174a ) or ( a175a );
 a3009a <=( a172a ) or ( a173a );
 a3010a <=( a3009a ) or ( a3006a );
 a3013a <=( a170a ) or ( a171a );
 a3016a <=( a168a ) or ( a169a );
 a3017a <=( a3016a ) or ( a3013a );
 a3018a <=( a3017a ) or ( a3010a );
 a3021a <=( a166a ) or ( a167a );
 a3024a <=( a164a ) or ( a165a );
 a3025a <=( a3024a ) or ( a3021a );
 a3028a <=( a162a ) or ( a163a );
 a3032a <=( a159a ) or ( a160a );
 a3033a <=( a161a ) or ( a3032a );
 a3034a <=( a3033a ) or ( a3028a );
 a3035a <=( a3034a ) or ( a3025a );
 a3036a <=( a3035a ) or ( a3018a );
 a3039a <=( a157a ) or ( a158a );
 a3042a <=( a155a ) or ( a156a );
 a3043a <=( a3042a ) or ( a3039a );
 a3046a <=( a153a ) or ( a154a );
 a3050a <=( a150a ) or ( a151a );
 a3051a <=( a152a ) or ( a3050a );
 a3052a <=( a3051a ) or ( a3046a );
 a3053a <=( a3052a ) or ( a3043a );
 a3056a <=( a148a ) or ( a149a );
 a3059a <=( a146a ) or ( a147a );
 a3060a <=( a3059a ) or ( a3056a );
 a3063a <=( a144a ) or ( a145a );
 a3067a <=( a141a ) or ( a142a );
 a3068a <=( a143a ) or ( a3067a );
 a3069a <=( a3068a ) or ( a3063a );
 a3070a <=( a3069a ) or ( a3060a );
 a3071a <=( a3070a ) or ( a3053a );
 a3072a <=( a3071a ) or ( a3036a );
 a3073a <=( a3072a ) or ( a3003a );
 a3074a <=( a3073a ) or ( a2934a );
 a3077a <=( a139a ) or ( a140a );
 a3080a <=( a137a ) or ( a138a );
 a3081a <=( a3080a ) or ( a3077a );
 a3084a <=( a135a ) or ( a136a );
 a3087a <=( a133a ) or ( a134a );
 a3088a <=( a3087a ) or ( a3084a );
 a3089a <=( a3088a ) or ( a3081a );
 a3092a <=( a131a ) or ( a132a );
 a3095a <=( a129a ) or ( a130a );
 a3096a <=( a3095a ) or ( a3092a );
 a3099a <=( a127a ) or ( a128a );
 a3103a <=( a124a ) or ( a125a );
 a3104a <=( a126a ) or ( a3103a );
 a3105a <=( a3104a ) or ( a3099a );
 a3106a <=( a3105a ) or ( a3096a );
 a3107a <=( a3106a ) or ( a3089a );
 a3110a <=( a122a ) or ( a123a );
 a3113a <=( a120a ) or ( a121a );
 a3114a <=( a3113a ) or ( a3110a );
 a3117a <=( a118a ) or ( a119a );
 a3121a <=( a115a ) or ( a116a );
 a3122a <=( a117a ) or ( a3121a );
 a3123a <=( a3122a ) or ( a3117a );
 a3124a <=( a3123a ) or ( a3114a );
 a3127a <=( a113a ) or ( a114a );
 a3130a <=( a111a ) or ( a112a );
 a3131a <=( a3130a ) or ( a3127a );
 a3134a <=( a109a ) or ( a110a );
 a3138a <=( a106a ) or ( a107a );
 a3139a <=( a108a ) or ( a3138a );
 a3140a <=( a3139a ) or ( a3134a );
 a3141a <=( a3140a ) or ( a3131a );
 a3142a <=( a3141a ) or ( a3124a );
 a3143a <=( a3142a ) or ( a3107a );
 a3146a <=( a104a ) or ( a105a );
 a3149a <=( a102a ) or ( a103a );
 a3150a <=( a3149a ) or ( a3146a );
 a3153a <=( a100a ) or ( a101a );
 a3156a <=( a98a ) or ( a99a );
 a3157a <=( a3156a ) or ( a3153a );
 a3158a <=( a3157a ) or ( a3150a );
 a3161a <=( a96a ) or ( a97a );
 a3164a <=( a94a ) or ( a95a );
 a3165a <=( a3164a ) or ( a3161a );
 a3168a <=( a92a ) or ( a93a );
 a3172a <=( a89a ) or ( a90a );
 a3173a <=( a91a ) or ( a3172a );
 a3174a <=( a3173a ) or ( a3168a );
 a3175a <=( a3174a ) or ( a3165a );
 a3176a <=( a3175a ) or ( a3158a );
 a3179a <=( a87a ) or ( a88a );
 a3182a <=( a85a ) or ( a86a );
 a3183a <=( a3182a ) or ( a3179a );
 a3186a <=( a83a ) or ( a84a );
 a3190a <=( a80a ) or ( a81a );
 a3191a <=( a82a ) or ( a3190a );
 a3192a <=( a3191a ) or ( a3186a );
 a3193a <=( a3192a ) or ( a3183a );
 a3196a <=( a78a ) or ( a79a );
 a3199a <=( a76a ) or ( a77a );
 a3200a <=( a3199a ) or ( a3196a );
 a3203a <=( a74a ) or ( a75a );
 a3207a <=( a71a ) or ( a72a );
 a3208a <=( a73a ) or ( a3207a );
 a3209a <=( a3208a ) or ( a3203a );
 a3210a <=( a3209a ) or ( a3200a );
 a3211a <=( a3210a ) or ( a3193a );
 a3212a <=( a3211a ) or ( a3176a );
 a3213a <=( a3212a ) or ( a3143a );
 a3216a <=( a69a ) or ( a70a );
 a3219a <=( a67a ) or ( a68a );
 a3220a <=( a3219a ) or ( a3216a );
 a3223a <=( a65a ) or ( a66a );
 a3226a <=( a63a ) or ( a64a );
 a3227a <=( a3226a ) or ( a3223a );
 a3228a <=( a3227a ) or ( a3220a );
 a3231a <=( a61a ) or ( a62a );
 a3234a <=( a59a ) or ( a60a );
 a3235a <=( a3234a ) or ( a3231a );
 a3238a <=( a57a ) or ( a58a );
 a3242a <=( a54a ) or ( a55a );
 a3243a <=( a56a ) or ( a3242a );
 a3244a <=( a3243a ) or ( a3238a );
 a3245a <=( a3244a ) or ( a3235a );
 a3246a <=( a3245a ) or ( a3228a );
 a3249a <=( a52a ) or ( a53a );
 a3252a <=( a50a ) or ( a51a );
 a3253a <=( a3252a ) or ( a3249a );
 a3256a <=( a48a ) or ( a49a );
 a3260a <=( a45a ) or ( a46a );
 a3261a <=( a47a ) or ( a3260a );
 a3262a <=( a3261a ) or ( a3256a );
 a3263a <=( a3262a ) or ( a3253a );
 a3266a <=( a43a ) or ( a44a );
 a3269a <=( a41a ) or ( a42a );
 a3270a <=( a3269a ) or ( a3266a );
 a3273a <=( a39a ) or ( a40a );
 a3277a <=( a36a ) or ( a37a );
 a3278a <=( a38a ) or ( a3277a );
 a3279a <=( a3278a ) or ( a3273a );
 a3280a <=( a3279a ) or ( a3270a );
 a3281a <=( a3280a ) or ( a3263a );
 a3282a <=( a3281a ) or ( a3246a );
 a3285a <=( a34a ) or ( a35a );
 a3288a <=( a32a ) or ( a33a );
 a3289a <=( a3288a ) or ( a3285a );
 a3292a <=( a30a ) or ( a31a );
 a3295a <=( a28a ) or ( a29a );
 a3296a <=( a3295a ) or ( a3292a );
 a3297a <=( a3296a ) or ( a3289a );
 a3300a <=( a26a ) or ( a27a );
 a3303a <=( a24a ) or ( a25a );
 a3304a <=( a3303a ) or ( a3300a );
 a3307a <=( a22a ) or ( a23a );
 a3311a <=( a19a ) or ( a20a );
 a3312a <=( a21a ) or ( a3311a );
 a3313a <=( a3312a ) or ( a3307a );
 a3314a <=( a3313a ) or ( a3304a );
 a3315a <=( a3314a ) or ( a3297a );
 a3318a <=( a17a ) or ( a18a );
 a3321a <=( a15a ) or ( a16a );
 a3322a <=( a3321a ) or ( a3318a );
 a3325a <=( a13a ) or ( a14a );
 a3329a <=( a10a ) or ( a11a );
 a3330a <=( a12a ) or ( a3329a );
 a3331a <=( a3330a ) or ( a3325a );
 a3332a <=( a3331a ) or ( a3322a );
 a3335a <=( a8a ) or ( a9a );
 a3338a <=( a6a ) or ( a7a );
 a3339a <=( a3338a ) or ( a3335a );
 a3342a <=( a4a ) or ( a5a );
 a3346a <=( a1a ) or ( a2a );
 a3347a <=( a3a ) or ( a3346a );
 a3348a <=( a3347a ) or ( a3342a );
 a3349a <=( a3348a ) or ( a3339a );
 a3350a <=( a3349a ) or ( a3332a );
 a3351a <=( a3350a ) or ( a3315a );
 a3352a <=( a3351a ) or ( a3282a );
 a3353a <=( a3352a ) or ( a3213a );
 a3354a <=( a3353a ) or ( a3074a );
 a3355a <=( a3354a ) or ( a2795a );
 a3358a <=( A200  and  (not A199) );
 a3361a <=( A233  and  (not A232) );
 a3364a <=( A166  and  A168 );
 a3367a <=( A233  and  (not A232) );
 a3370a <=( A167  and  A168 );
 a3373a <=( A233  and  (not A232) );
 a3377a <=( A232  and  A200 );
 a3378a <=( (not A199)  and  a3377a );
 a3382a <=( A235  and  A234 );
 a3383a <=( (not A233)  and  a3382a );
 a3387a <=( A232  and  A200 );
 a3388a <=( (not A199)  and  a3387a );
 a3392a <=( A236  and  A234 );
 a3393a <=( (not A233)  and  a3392a );
 a3397a <=( A201  and  (not A200) );
 a3398a <=( A199  and  a3397a );
 a3402a <=( A233  and  (not A232) );
 a3403a <=( A202  and  a3402a );
 a3407a <=( A201  and  (not A200) );
 a3408a <=( A199  and  a3407a );
 a3412a <=( A233  and  (not A232) );
 a3413a <=( A203  and  a3412a );
 a3417a <=( A232  and  A166 );
 a3418a <=( A168  and  a3417a );
 a3422a <=( A235  and  A234 );
 a3423a <=( (not A233)  and  a3422a );
 a3427a <=( A232  and  A166 );
 a3428a <=( A168  and  a3427a );
 a3432a <=( A236  and  A234 );
 a3433a <=( (not A233)  and  a3432a );
 a3437a <=( A232  and  A167 );
 a3438a <=( A168  and  a3437a );
 a3442a <=( A235  and  A234 );
 a3443a <=( (not A233)  and  a3442a );
 a3447a <=( A232  and  A167 );
 a3448a <=( A168  and  a3447a );
 a3452a <=( A236  and  A234 );
 a3453a <=( (not A233)  and  a3452a );
 a3457a <=( A167  and  A169 );
 a3458a <=( (not A170)  and  a3457a );
 a3462a <=( A233  and  (not A232) );
 a3463a <=( A166  and  a3462a );
 a3467a <=( (not A167)  and  A169 );
 a3468a <=( (not A170)  and  a3467a );
 a3472a <=( A233  and  (not A232) );
 a3473a <=( (not A166)  and  a3472a );
 a3477a <=( A167  and  (not A169) );
 a3478a <=( A170  and  a3477a );
 a3482a <=( A233  and  (not A232) );
 a3483a <=( (not A166)  and  a3482a );
 a3487a <=( (not A167)  and  (not A169) );
 a3488a <=( A170  and  a3487a );
 a3492a <=( A233  and  (not A232) );
 a3493a <=( A166  and  a3492a );
 a3496a <=( (not A200)  and  A199 );
 a3499a <=( A202  and  A201 );
 a3500a <=( a3499a  and  a3496a );
 a3503a <=( (not A233)  and  A232 );
 a3506a <=( A235  and  A234 );
 a3507a <=( a3506a  and  a3503a );
 a3510a <=( (not A200)  and  A199 );
 a3513a <=( A202  and  A201 );
 a3514a <=( a3513a  and  a3510a );
 a3517a <=( (not A233)  and  A232 );
 a3520a <=( A236  and  A234 );
 a3521a <=( a3520a  and  a3517a );
 a3524a <=( (not A200)  and  A199 );
 a3527a <=( A203  and  A201 );
 a3528a <=( a3527a  and  a3524a );
 a3531a <=( (not A233)  and  A232 );
 a3534a <=( A235  and  A234 );
 a3535a <=( a3534a  and  a3531a );
 a3538a <=( (not A200)  and  A199 );
 a3541a <=( A203  and  A201 );
 a3542a <=( a3541a  and  a3538a );
 a3545a <=( (not A233)  and  A232 );
 a3548a <=( A236  and  A234 );
 a3549a <=( a3548a  and  a3545a );
 a3552a <=( A166  and  A168 );
 a3555a <=( A200  and  A199 );
 a3556a <=( a3555a  and  a3552a );
 a3559a <=( A266  and  A265 );
 a3562a <=( A299  and  (not A298) );
 a3563a <=( a3562a  and  a3559a );
 a3566a <=( A166  and  A168 );
 a3569a <=( A200  and  A199 );
 a3570a <=( a3569a  and  a3566a );
 a3573a <=( (not A267)  and  (not A266) );
 a3576a <=( A299  and  (not A298) );
 a3577a <=( a3576a  and  a3573a );
 a3580a <=( A166  and  A168 );
 a3583a <=( A200  and  A199 );
 a3584a <=( a3583a  and  a3580a );
 a3587a <=( (not A266)  and  (not A265) );
 a3590a <=( A299  and  (not A298) );
 a3591a <=( a3590a  and  a3587a );
 a3594a <=( A166  and  A168 );
 a3597a <=( A200  and  (not A199) );
 a3598a <=( a3597a  and  a3594a );
 a3601a <=( A266  and  (not A265) );
 a3604a <=( (not A300)  and  A298 );
 a3605a <=( a3604a  and  a3601a );
 a3608a <=( A166  and  A168 );
 a3611a <=( A200  and  (not A199) );
 a3612a <=( a3611a  and  a3608a );
 a3615a <=( A266  and  (not A265) );
 a3618a <=( A299  and  A298 );
 a3619a <=( a3618a  and  a3615a );
 a3622a <=( A166  and  A168 );
 a3625a <=( A200  and  (not A199) );
 a3626a <=( a3625a  and  a3622a );
 a3629a <=( A266  and  (not A265) );
 a3632a <=( (not A299)  and  (not A298) );
 a3633a <=( a3632a  and  a3629a );
 a3636a <=( A166  and  A168 );
 a3639a <=( (not A201)  and  (not A200) );
 a3640a <=( a3639a  and  a3636a );
 a3643a <=( A266  and  A265 );
 a3646a <=( A299  and  (not A298) );
 a3647a <=( a3646a  and  a3643a );
 a3650a <=( A166  and  A168 );
 a3653a <=( (not A201)  and  (not A200) );
 a3654a <=( a3653a  and  a3650a );
 a3657a <=( (not A267)  and  (not A266) );
 a3660a <=( A299  and  (not A298) );
 a3661a <=( a3660a  and  a3657a );
 a3664a <=( A166  and  A168 );
 a3667a <=( (not A201)  and  (not A200) );
 a3668a <=( a3667a  and  a3664a );
 a3671a <=( (not A266)  and  (not A265) );
 a3674a <=( A299  and  (not A298) );
 a3675a <=( a3674a  and  a3671a );
 a3678a <=( A166  and  A168 );
 a3681a <=( (not A200)  and  (not A199) );
 a3682a <=( a3681a  and  a3678a );
 a3685a <=( A266  and  A265 );
 a3688a <=( A299  and  (not A298) );
 a3689a <=( a3688a  and  a3685a );
 a3692a <=( A166  and  A168 );
 a3695a <=( (not A200)  and  (not A199) );
 a3696a <=( a3695a  and  a3692a );
 a3699a <=( (not A267)  and  (not A266) );
 a3702a <=( A299  and  (not A298) );
 a3703a <=( a3702a  and  a3699a );
 a3706a <=( A166  and  A168 );
 a3709a <=( (not A200)  and  (not A199) );
 a3710a <=( a3709a  and  a3706a );
 a3713a <=( (not A266)  and  (not A265) );
 a3716a <=( A299  and  (not A298) );
 a3717a <=( a3716a  and  a3713a );
 a3720a <=( A167  and  A168 );
 a3723a <=( A200  and  A199 );
 a3724a <=( a3723a  and  a3720a );
 a3727a <=( A266  and  A265 );
 a3730a <=( A299  and  (not A298) );
 a3731a <=( a3730a  and  a3727a );
 a3734a <=( A167  and  A168 );
 a3737a <=( A200  and  A199 );
 a3738a <=( a3737a  and  a3734a );
 a3741a <=( (not A267)  and  (not A266) );
 a3744a <=( A299  and  (not A298) );
 a3745a <=( a3744a  and  a3741a );
 a3748a <=( A167  and  A168 );
 a3751a <=( A200  and  A199 );
 a3752a <=( a3751a  and  a3748a );
 a3755a <=( (not A266)  and  (not A265) );
 a3758a <=( A299  and  (not A298) );
 a3759a <=( a3758a  and  a3755a );
 a3762a <=( A167  and  A168 );
 a3765a <=( A200  and  (not A199) );
 a3766a <=( a3765a  and  a3762a );
 a3769a <=( A266  and  (not A265) );
 a3772a <=( (not A300)  and  A298 );
 a3773a <=( a3772a  and  a3769a );
 a3776a <=( A167  and  A168 );
 a3779a <=( A200  and  (not A199) );
 a3780a <=( a3779a  and  a3776a );
 a3783a <=( A266  and  (not A265) );
 a3786a <=( A299  and  A298 );
 a3787a <=( a3786a  and  a3783a );
 a3790a <=( A167  and  A168 );
 a3793a <=( A200  and  (not A199) );
 a3794a <=( a3793a  and  a3790a );
 a3797a <=( A266  and  (not A265) );
 a3800a <=( (not A299)  and  (not A298) );
 a3801a <=( a3800a  and  a3797a );
 a3804a <=( A167  and  A168 );
 a3807a <=( (not A201)  and  (not A200) );
 a3808a <=( a3807a  and  a3804a );
 a3811a <=( A266  and  A265 );
 a3814a <=( A299  and  (not A298) );
 a3815a <=( a3814a  and  a3811a );
 a3818a <=( A167  and  A168 );
 a3821a <=( (not A201)  and  (not A200) );
 a3822a <=( a3821a  and  a3818a );
 a3825a <=( (not A267)  and  (not A266) );
 a3828a <=( A299  and  (not A298) );
 a3829a <=( a3828a  and  a3825a );
 a3832a <=( A167  and  A168 );
 a3835a <=( (not A201)  and  (not A200) );
 a3836a <=( a3835a  and  a3832a );
 a3839a <=( (not A266)  and  (not A265) );
 a3842a <=( A299  and  (not A298) );
 a3843a <=( a3842a  and  a3839a );
 a3846a <=( A167  and  A168 );
 a3849a <=( (not A200)  and  (not A199) );
 a3850a <=( a3849a  and  a3846a );
 a3853a <=( A266  and  A265 );
 a3856a <=( A299  and  (not A298) );
 a3857a <=( a3856a  and  a3853a );
 a3860a <=( A167  and  A168 );
 a3863a <=( (not A200)  and  (not A199) );
 a3864a <=( a3863a  and  a3860a );
 a3867a <=( (not A267)  and  (not A266) );
 a3870a <=( A299  and  (not A298) );
 a3871a <=( a3870a  and  a3867a );
 a3874a <=( A167  and  A168 );
 a3877a <=( (not A200)  and  (not A199) );
 a3878a <=( a3877a  and  a3874a );
 a3881a <=( (not A266)  and  (not A265) );
 a3884a <=( A299  and  (not A298) );
 a3885a <=( a3884a  and  a3881a );
 a3888a <=( A169  and  (not A170) );
 a3891a <=( A166  and  A167 );
 a3892a <=( a3891a  and  a3888a );
 a3895a <=( (not A233)  and  A232 );
 a3898a <=( A235  and  A234 );
 a3899a <=( a3898a  and  a3895a );
 a3902a <=( A169  and  (not A170) );
 a3905a <=( A166  and  A167 );
 a3906a <=( a3905a  and  a3902a );
 a3909a <=( (not A233)  and  A232 );
 a3912a <=( A236  and  A234 );
 a3913a <=( a3912a  and  a3909a );
 a3916a <=( A169  and  (not A170) );
 a3919a <=( (not A166)  and  (not A167) );
 a3920a <=( a3919a  and  a3916a );
 a3923a <=( (not A233)  and  A232 );
 a3926a <=( A235  and  A234 );
 a3927a <=( a3926a  and  a3923a );
 a3930a <=( A169  and  (not A170) );
 a3933a <=( (not A166)  and  (not A167) );
 a3934a <=( a3933a  and  a3930a );
 a3937a <=( (not A233)  and  A232 );
 a3940a <=( A236  and  A234 );
 a3941a <=( a3940a  and  a3937a );
 a3944a <=( (not A169)  and  A170 );
 a3947a <=( (not A166)  and  A167 );
 a3948a <=( a3947a  and  a3944a );
 a3951a <=( (not A233)  and  A232 );
 a3954a <=( A235  and  A234 );
 a3955a <=( a3954a  and  a3951a );
 a3958a <=( (not A169)  and  A170 );
 a3961a <=( (not A166)  and  A167 );
 a3962a <=( a3961a  and  a3958a );
 a3965a <=( (not A233)  and  A232 );
 a3968a <=( A236  and  A234 );
 a3969a <=( a3968a  and  a3965a );
 a3972a <=( (not A169)  and  A170 );
 a3975a <=( A166  and  (not A167) );
 a3976a <=( a3975a  and  a3972a );
 a3979a <=( (not A233)  and  A232 );
 a3982a <=( A235  and  A234 );
 a3983a <=( a3982a  and  a3979a );
 a3986a <=( (not A169)  and  A170 );
 a3989a <=( A166  and  (not A167) );
 a3990a <=( a3989a  and  a3986a );
 a3993a <=( (not A233)  and  A232 );
 a3996a <=( A236  and  A234 );
 a3997a <=( a3996a  and  a3993a );
 a4000a <=( A166  and  A168 );
 a4003a <=( A200  and  A199 );
 a4004a <=( a4003a  and  a4000a );
 a4007a <=( (not A268)  and  (not A266) );
 a4011a <=( A299  and  (not A298) );
 a4012a <=( (not A269)  and  a4011a );
 a4013a <=( a4012a  and  a4007a );
 a4016a <=( A166  and  A168 );
 a4019a <=( A200  and  (not A199) );
 a4020a <=( a4019a  and  a4016a );
 a4023a <=( A266  and  (not A265) );
 a4027a <=( (not A302)  and  (not A301) );
 a4028a <=( A298  and  a4027a );
 a4029a <=( a4028a  and  a4023a );
 a4032a <=( A166  and  A168 );
 a4035a <=( (not A202)  and  (not A200) );
 a4036a <=( a4035a  and  a4032a );
 a4039a <=( A265  and  (not A203) );
 a4043a <=( A299  and  (not A298) );
 a4044a <=( A266  and  a4043a );
 a4045a <=( a4044a  and  a4039a );
 a4048a <=( A166  and  A168 );
 a4051a <=( (not A202)  and  (not A200) );
 a4052a <=( a4051a  and  a4048a );
 a4055a <=( (not A266)  and  (not A203) );
 a4059a <=( A299  and  (not A298) );
 a4060a <=( (not A267)  and  a4059a );
 a4061a <=( a4060a  and  a4055a );
 a4064a <=( A166  and  A168 );
 a4067a <=( (not A202)  and  (not A200) );
 a4068a <=( a4067a  and  a4064a );
 a4071a <=( (not A265)  and  (not A203) );
 a4075a <=( A299  and  (not A298) );
 a4076a <=( (not A266)  and  a4075a );
 a4077a <=( a4076a  and  a4071a );
 a4080a <=( A166  and  A168 );
 a4083a <=( (not A201)  and  (not A200) );
 a4084a <=( a4083a  and  a4080a );
 a4087a <=( (not A268)  and  (not A266) );
 a4091a <=( A299  and  (not A298) );
 a4092a <=( (not A269)  and  a4091a );
 a4093a <=( a4092a  and  a4087a );
 a4096a <=( A166  and  A168 );
 a4099a <=( (not A200)  and  (not A199) );
 a4100a <=( a4099a  and  a4096a );
 a4103a <=( (not A268)  and  (not A266) );
 a4107a <=( A299  and  (not A298) );
 a4108a <=( (not A269)  and  a4107a );
 a4109a <=( a4108a  and  a4103a );
 a4112a <=( A167  and  A168 );
 a4115a <=( A200  and  A199 );
 a4116a <=( a4115a  and  a4112a );
 a4119a <=( (not A268)  and  (not A266) );
 a4123a <=( A299  and  (not A298) );
 a4124a <=( (not A269)  and  a4123a );
 a4125a <=( a4124a  and  a4119a );
 a4128a <=( A167  and  A168 );
 a4131a <=( A200  and  (not A199) );
 a4132a <=( a4131a  and  a4128a );
 a4135a <=( A266  and  (not A265) );
 a4139a <=( (not A302)  and  (not A301) );
 a4140a <=( A298  and  a4139a );
 a4141a <=( a4140a  and  a4135a );
 a4144a <=( A167  and  A168 );
 a4147a <=( (not A202)  and  (not A200) );
 a4148a <=( a4147a  and  a4144a );
 a4151a <=( A265  and  (not A203) );
 a4155a <=( A299  and  (not A298) );
 a4156a <=( A266  and  a4155a );
 a4157a <=( a4156a  and  a4151a );
 a4160a <=( A167  and  A168 );
 a4163a <=( (not A202)  and  (not A200) );
 a4164a <=( a4163a  and  a4160a );
 a4167a <=( (not A266)  and  (not A203) );
 a4171a <=( A299  and  (not A298) );
 a4172a <=( (not A267)  and  a4171a );
 a4173a <=( a4172a  and  a4167a );
 a4176a <=( A167  and  A168 );
 a4179a <=( (not A202)  and  (not A200) );
 a4180a <=( a4179a  and  a4176a );
 a4183a <=( (not A265)  and  (not A203) );
 a4187a <=( A299  and  (not A298) );
 a4188a <=( (not A266)  and  a4187a );
 a4189a <=( a4188a  and  a4183a );
 a4192a <=( A167  and  A168 );
 a4195a <=( (not A201)  and  (not A200) );
 a4196a <=( a4195a  and  a4192a );
 a4199a <=( (not A268)  and  (not A266) );
 a4203a <=( A299  and  (not A298) );
 a4204a <=( (not A269)  and  a4203a );
 a4205a <=( a4204a  and  a4199a );
 a4208a <=( A167  and  A168 );
 a4211a <=( (not A200)  and  (not A199) );
 a4212a <=( a4211a  and  a4208a );
 a4215a <=( (not A268)  and  (not A266) );
 a4219a <=( A299  and  (not A298) );
 a4220a <=( (not A269)  and  a4219a );
 a4221a <=( a4220a  and  a4215a );
 a4224a <=( (not A167)  and  A170 );
 a4227a <=( A199  and  (not A166) );
 a4228a <=( a4227a  and  a4224a );
 a4231a <=( (not A265)  and  A200 );
 a4235a <=( (not A300)  and  A298 );
 a4236a <=( A266  and  a4235a );
 a4237a <=( a4236a  and  a4231a );
 a4240a <=( (not A167)  and  A170 );
 a4243a <=( A199  and  (not A166) );
 a4244a <=( a4243a  and  a4240a );
 a4247a <=( (not A265)  and  A200 );
 a4251a <=( A299  and  A298 );
 a4252a <=( A266  and  a4251a );
 a4253a <=( a4252a  and  a4247a );
 a4256a <=( (not A167)  and  A170 );
 a4259a <=( A199  and  (not A166) );
 a4260a <=( a4259a  and  a4256a );
 a4263a <=( (not A265)  and  A200 );
 a4267a <=( (not A299)  and  (not A298) );
 a4268a <=( A266  and  a4267a );
 a4269a <=( a4268a  and  a4263a );
 a4272a <=( (not A167)  and  A170 );
 a4275a <=( (not A199)  and  (not A166) );
 a4276a <=( a4275a  and  a4272a );
 a4279a <=( A265  and  A200 );
 a4283a <=( A299  and  (not A298) );
 a4284a <=( A266  and  a4283a );
 a4285a <=( a4284a  and  a4279a );
 a4288a <=( (not A167)  and  A170 );
 a4291a <=( (not A199)  and  (not A166) );
 a4292a <=( a4291a  and  a4288a );
 a4295a <=( (not A266)  and  A200 );
 a4299a <=( A299  and  (not A298) );
 a4300a <=( (not A267)  and  a4299a );
 a4301a <=( a4300a  and  a4295a );
 a4304a <=( (not A167)  and  A170 );
 a4307a <=( (not A199)  and  (not A166) );
 a4308a <=( a4307a  and  a4304a );
 a4311a <=( (not A265)  and  A200 );
 a4315a <=( A299  and  (not A298) );
 a4316a <=( (not A266)  and  a4315a );
 a4317a <=( a4316a  and  a4311a );
 a4320a <=( (not A167)  and  A170 );
 a4323a <=( (not A200)  and  (not A166) );
 a4324a <=( a4323a  and  a4320a );
 a4327a <=( (not A265)  and  (not A201) );
 a4331a <=( (not A300)  and  A298 );
 a4332a <=( A266  and  a4331a );
 a4333a <=( a4332a  and  a4327a );
 a4336a <=( (not A167)  and  A170 );
 a4339a <=( (not A200)  and  (not A166) );
 a4340a <=( a4339a  and  a4336a );
 a4343a <=( (not A265)  and  (not A201) );
 a4347a <=( A299  and  A298 );
 a4348a <=( A266  and  a4347a );
 a4349a <=( a4348a  and  a4343a );
 a4352a <=( (not A167)  and  A170 );
 a4355a <=( (not A200)  and  (not A166) );
 a4356a <=( a4355a  and  a4352a );
 a4359a <=( (not A265)  and  (not A201) );
 a4363a <=( (not A299)  and  (not A298) );
 a4364a <=( A266  and  a4363a );
 a4365a <=( a4364a  and  a4359a );
 a4368a <=( (not A167)  and  A170 );
 a4371a <=( (not A199)  and  (not A166) );
 a4372a <=( a4371a  and  a4368a );
 a4375a <=( (not A265)  and  (not A200) );
 a4379a <=( (not A300)  and  A298 );
 a4380a <=( A266  and  a4379a );
 a4381a <=( a4380a  and  a4375a );
 a4384a <=( (not A167)  and  A170 );
 a4387a <=( (not A199)  and  (not A166) );
 a4388a <=( a4387a  and  a4384a );
 a4391a <=( (not A265)  and  (not A200) );
 a4395a <=( A299  and  A298 );
 a4396a <=( A266  and  a4395a );
 a4397a <=( a4396a  and  a4391a );
 a4400a <=( (not A167)  and  A170 );
 a4403a <=( (not A199)  and  (not A166) );
 a4404a <=( a4403a  and  a4400a );
 a4407a <=( (not A265)  and  (not A200) );
 a4411a <=( (not A299)  and  (not A298) );
 a4412a <=( A266  and  a4411a );
 a4413a <=( a4412a  and  a4407a );
 a4416a <=( A169  and  A170 );
 a4419a <=( A199  and  (not A168) );
 a4420a <=( a4419a  and  a4416a );
 a4423a <=( (not A265)  and  A200 );
 a4427a <=( (not A300)  and  A298 );
 a4428a <=( A266  and  a4427a );
 a4429a <=( a4428a  and  a4423a );
 a4432a <=( A169  and  A170 );
 a4435a <=( A199  and  (not A168) );
 a4436a <=( a4435a  and  a4432a );
 a4439a <=( (not A265)  and  A200 );
 a4443a <=( A299  and  A298 );
 a4444a <=( A266  and  a4443a );
 a4445a <=( a4444a  and  a4439a );
 a4448a <=( A169  and  A170 );
 a4451a <=( A199  and  (not A168) );
 a4452a <=( a4451a  and  a4448a );
 a4455a <=( (not A265)  and  A200 );
 a4459a <=( (not A299)  and  (not A298) );
 a4460a <=( A266  and  a4459a );
 a4461a <=( a4460a  and  a4455a );
 a4464a <=( A169  and  A170 );
 a4467a <=( (not A199)  and  (not A168) );
 a4468a <=( a4467a  and  a4464a );
 a4471a <=( A265  and  A200 );
 a4475a <=( A299  and  (not A298) );
 a4476a <=( A266  and  a4475a );
 a4477a <=( a4476a  and  a4471a );
 a4480a <=( A169  and  A170 );
 a4483a <=( (not A199)  and  (not A168) );
 a4484a <=( a4483a  and  a4480a );
 a4487a <=( (not A266)  and  A200 );
 a4491a <=( A299  and  (not A298) );
 a4492a <=( (not A267)  and  a4491a );
 a4493a <=( a4492a  and  a4487a );
 a4496a <=( A169  and  A170 );
 a4499a <=( (not A199)  and  (not A168) );
 a4500a <=( a4499a  and  a4496a );
 a4503a <=( (not A265)  and  A200 );
 a4507a <=( A299  and  (not A298) );
 a4508a <=( (not A266)  and  a4507a );
 a4509a <=( a4508a  and  a4503a );
 a4512a <=( A169  and  A170 );
 a4515a <=( (not A200)  and  (not A168) );
 a4516a <=( a4515a  and  a4512a );
 a4519a <=( (not A265)  and  (not A201) );
 a4523a <=( (not A300)  and  A298 );
 a4524a <=( A266  and  a4523a );
 a4525a <=( a4524a  and  a4519a );
 a4528a <=( A169  and  A170 );
 a4531a <=( (not A200)  and  (not A168) );
 a4532a <=( a4531a  and  a4528a );
 a4535a <=( (not A265)  and  (not A201) );
 a4539a <=( A299  and  A298 );
 a4540a <=( A266  and  a4539a );
 a4541a <=( a4540a  and  a4535a );
 a4544a <=( A169  and  A170 );
 a4547a <=( (not A200)  and  (not A168) );
 a4548a <=( a4547a  and  a4544a );
 a4551a <=( (not A265)  and  (not A201) );
 a4555a <=( (not A299)  and  (not A298) );
 a4556a <=( A266  and  a4555a );
 a4557a <=( a4556a  and  a4551a );
 a4560a <=( A169  and  A170 );
 a4563a <=( (not A199)  and  (not A168) );
 a4564a <=( a4563a  and  a4560a );
 a4567a <=( (not A265)  and  (not A200) );
 a4571a <=( (not A300)  and  A298 );
 a4572a <=( A266  and  a4571a );
 a4573a <=( a4572a  and  a4567a );
 a4576a <=( A169  and  A170 );
 a4579a <=( (not A199)  and  (not A168) );
 a4580a <=( a4579a  and  a4576a );
 a4583a <=( (not A265)  and  (not A200) );
 a4587a <=( A299  and  A298 );
 a4588a <=( A266  and  a4587a );
 a4589a <=( a4588a  and  a4583a );
 a4592a <=( A169  and  A170 );
 a4595a <=( (not A199)  and  (not A168) );
 a4596a <=( a4595a  and  a4592a );
 a4599a <=( (not A265)  and  (not A200) );
 a4603a <=( (not A299)  and  (not A298) );
 a4604a <=( A266  and  a4603a );
 a4605a <=( a4604a  and  a4599a );
 a4608a <=( (not A167)  and  (not A169) );
 a4611a <=( A199  and  (not A166) );
 a4612a <=( a4611a  and  a4608a );
 a4615a <=( (not A265)  and  A200 );
 a4619a <=( (not A300)  and  A298 );
 a4620a <=( A266  and  a4619a );
 a4621a <=( a4620a  and  a4615a );
 a4624a <=( (not A167)  and  (not A169) );
 a4627a <=( A199  and  (not A166) );
 a4628a <=( a4627a  and  a4624a );
 a4631a <=( (not A265)  and  A200 );
 a4635a <=( A299  and  A298 );
 a4636a <=( A266  and  a4635a );
 a4637a <=( a4636a  and  a4631a );
 a4640a <=( (not A167)  and  (not A169) );
 a4643a <=( A199  and  (not A166) );
 a4644a <=( a4643a  and  a4640a );
 a4647a <=( (not A265)  and  A200 );
 a4651a <=( (not A299)  and  (not A298) );
 a4652a <=( A266  and  a4651a );
 a4653a <=( a4652a  and  a4647a );
 a4656a <=( (not A167)  and  (not A169) );
 a4659a <=( (not A199)  and  (not A166) );
 a4660a <=( a4659a  and  a4656a );
 a4663a <=( A265  and  A200 );
 a4667a <=( A299  and  (not A298) );
 a4668a <=( A266  and  a4667a );
 a4669a <=( a4668a  and  a4663a );
 a4672a <=( (not A167)  and  (not A169) );
 a4675a <=( (not A199)  and  (not A166) );
 a4676a <=( a4675a  and  a4672a );
 a4679a <=( (not A266)  and  A200 );
 a4683a <=( A299  and  (not A298) );
 a4684a <=( (not A267)  and  a4683a );
 a4685a <=( a4684a  and  a4679a );
 a4688a <=( (not A167)  and  (not A169) );
 a4691a <=( (not A199)  and  (not A166) );
 a4692a <=( a4691a  and  a4688a );
 a4695a <=( (not A265)  and  A200 );
 a4699a <=( A299  and  (not A298) );
 a4700a <=( (not A266)  and  a4699a );
 a4701a <=( a4700a  and  a4695a );
 a4704a <=( (not A167)  and  (not A169) );
 a4707a <=( (not A200)  and  (not A166) );
 a4708a <=( a4707a  and  a4704a );
 a4711a <=( (not A265)  and  (not A201) );
 a4715a <=( (not A300)  and  A298 );
 a4716a <=( A266  and  a4715a );
 a4717a <=( a4716a  and  a4711a );
 a4720a <=( (not A167)  and  (not A169) );
 a4723a <=( (not A200)  and  (not A166) );
 a4724a <=( a4723a  and  a4720a );
 a4727a <=( (not A265)  and  (not A201) );
 a4731a <=( A299  and  A298 );
 a4732a <=( A266  and  a4731a );
 a4733a <=( a4732a  and  a4727a );
 a4736a <=( (not A167)  and  (not A169) );
 a4739a <=( (not A200)  and  (not A166) );
 a4740a <=( a4739a  and  a4736a );
 a4743a <=( (not A265)  and  (not A201) );
 a4747a <=( (not A299)  and  (not A298) );
 a4748a <=( A266  and  a4747a );
 a4749a <=( a4748a  and  a4743a );
 a4752a <=( (not A167)  and  (not A169) );
 a4755a <=( (not A199)  and  (not A166) );
 a4756a <=( a4755a  and  a4752a );
 a4759a <=( (not A265)  and  (not A200) );
 a4763a <=( (not A300)  and  A298 );
 a4764a <=( A266  and  a4763a );
 a4765a <=( a4764a  and  a4759a );
 a4768a <=( (not A167)  and  (not A169) );
 a4771a <=( (not A199)  and  (not A166) );
 a4772a <=( a4771a  and  a4768a );
 a4775a <=( (not A265)  and  (not A200) );
 a4779a <=( A299  and  A298 );
 a4780a <=( A266  and  a4779a );
 a4781a <=( a4780a  and  a4775a );
 a4784a <=( (not A167)  and  (not A169) );
 a4787a <=( (not A199)  and  (not A166) );
 a4788a <=( a4787a  and  a4784a );
 a4791a <=( (not A265)  and  (not A200) );
 a4795a <=( (not A299)  and  (not A298) );
 a4796a <=( A266  and  a4795a );
 a4797a <=( a4796a  and  a4791a );
 a4800a <=( (not A169)  and  (not A170) );
 a4803a <=( A199  and  (not A168) );
 a4804a <=( a4803a  and  a4800a );
 a4807a <=( (not A265)  and  A200 );
 a4811a <=( (not A300)  and  A298 );
 a4812a <=( A266  and  a4811a );
 a4813a <=( a4812a  and  a4807a );
 a4816a <=( (not A169)  and  (not A170) );
 a4819a <=( A199  and  (not A168) );
 a4820a <=( a4819a  and  a4816a );
 a4823a <=( (not A265)  and  A200 );
 a4827a <=( A299  and  A298 );
 a4828a <=( A266  and  a4827a );
 a4829a <=( a4828a  and  a4823a );
 a4832a <=( (not A169)  and  (not A170) );
 a4835a <=( A199  and  (not A168) );
 a4836a <=( a4835a  and  a4832a );
 a4839a <=( (not A265)  and  A200 );
 a4843a <=( (not A299)  and  (not A298) );
 a4844a <=( A266  and  a4843a );
 a4845a <=( a4844a  and  a4839a );
 a4848a <=( (not A169)  and  (not A170) );
 a4851a <=( (not A199)  and  (not A168) );
 a4852a <=( a4851a  and  a4848a );
 a4855a <=( A265  and  A200 );
 a4859a <=( A299  and  (not A298) );
 a4860a <=( A266  and  a4859a );
 a4861a <=( a4860a  and  a4855a );
 a4864a <=( (not A169)  and  (not A170) );
 a4867a <=( (not A199)  and  (not A168) );
 a4868a <=( a4867a  and  a4864a );
 a4871a <=( (not A266)  and  A200 );
 a4875a <=( A299  and  (not A298) );
 a4876a <=( (not A267)  and  a4875a );
 a4877a <=( a4876a  and  a4871a );
 a4880a <=( (not A169)  and  (not A170) );
 a4883a <=( (not A199)  and  (not A168) );
 a4884a <=( a4883a  and  a4880a );
 a4887a <=( (not A265)  and  A200 );
 a4891a <=( A299  and  (not A298) );
 a4892a <=( (not A266)  and  a4891a );
 a4893a <=( a4892a  and  a4887a );
 a4896a <=( (not A169)  and  (not A170) );
 a4899a <=( (not A200)  and  (not A168) );
 a4900a <=( a4899a  and  a4896a );
 a4903a <=( (not A265)  and  (not A201) );
 a4907a <=( (not A300)  and  A298 );
 a4908a <=( A266  and  a4907a );
 a4909a <=( a4908a  and  a4903a );
 a4912a <=( (not A169)  and  (not A170) );
 a4915a <=( (not A200)  and  (not A168) );
 a4916a <=( a4915a  and  a4912a );
 a4919a <=( (not A265)  and  (not A201) );
 a4923a <=( A299  and  A298 );
 a4924a <=( A266  and  a4923a );
 a4925a <=( a4924a  and  a4919a );
 a4928a <=( (not A169)  and  (not A170) );
 a4931a <=( (not A200)  and  (not A168) );
 a4932a <=( a4931a  and  a4928a );
 a4935a <=( (not A265)  and  (not A201) );
 a4939a <=( (not A299)  and  (not A298) );
 a4940a <=( A266  and  a4939a );
 a4941a <=( a4940a  and  a4935a );
 a4944a <=( (not A169)  and  (not A170) );
 a4947a <=( (not A199)  and  (not A168) );
 a4948a <=( a4947a  and  a4944a );
 a4951a <=( (not A265)  and  (not A200) );
 a4955a <=( (not A300)  and  A298 );
 a4956a <=( A266  and  a4955a );
 a4957a <=( a4956a  and  a4951a );
 a4960a <=( (not A169)  and  (not A170) );
 a4963a <=( (not A199)  and  (not A168) );
 a4964a <=( a4963a  and  a4960a );
 a4967a <=( (not A265)  and  (not A200) );
 a4971a <=( A299  and  A298 );
 a4972a <=( A266  and  a4971a );
 a4973a <=( a4972a  and  a4967a );
 a4976a <=( (not A169)  and  (not A170) );
 a4979a <=( (not A199)  and  (not A168) );
 a4980a <=( a4979a  and  a4976a );
 a4983a <=( (not A265)  and  (not A200) );
 a4987a <=( (not A299)  and  (not A298) );
 a4988a <=( A266  and  a4987a );
 a4989a <=( a4988a  and  a4983a );
 a4992a <=( A166  and  A168 );
 a4996a <=( A265  and  A200 );
 a4997a <=( A199  and  a4996a );
 a4998a <=( a4997a  and  a4992a );
 a5001a <=( A298  and  A266 );
 a5005a <=( A301  and  A300 );
 a5006a <=( (not A299)  and  a5005a );
 a5007a <=( a5006a  and  a5001a );
 a5010a <=( A166  and  A168 );
 a5014a <=( A265  and  A200 );
 a5015a <=( A199  and  a5014a );
 a5016a <=( a5015a  and  a5010a );
 a5019a <=( A298  and  A266 );
 a5023a <=( A302  and  A300 );
 a5024a <=( (not A299)  and  a5023a );
 a5025a <=( a5024a  and  a5019a );
 a5028a <=( A166  and  A168 );
 a5032a <=( (not A266)  and  A200 );
 a5033a <=( A199  and  a5032a );
 a5034a <=( a5033a  and  a5028a );
 a5037a <=( A298  and  (not A267) );
 a5041a <=( A301  and  A300 );
 a5042a <=( (not A299)  and  a5041a );
 a5043a <=( a5042a  and  a5037a );
 a5046a <=( A166  and  A168 );
 a5050a <=( (not A266)  and  A200 );
 a5051a <=( A199  and  a5050a );
 a5052a <=( a5051a  and  a5046a );
 a5055a <=( A298  and  (not A267) );
 a5059a <=( A302  and  A300 );
 a5060a <=( (not A299)  and  a5059a );
 a5061a <=( a5060a  and  a5055a );
 a5064a <=( A166  and  A168 );
 a5068a <=( (not A265)  and  A200 );
 a5069a <=( A199  and  a5068a );
 a5070a <=( a5069a  and  a5064a );
 a5073a <=( A298  and  (not A266) );
 a5077a <=( A301  and  A300 );
 a5078a <=( (not A299)  and  a5077a );
 a5079a <=( a5078a  and  a5073a );
 a5082a <=( A166  and  A168 );
 a5086a <=( (not A265)  and  A200 );
 a5087a <=( A199  and  a5086a );
 a5088a <=( a5087a  and  a5082a );
 a5091a <=( A298  and  (not A266) );
 a5095a <=( A302  and  A300 );
 a5096a <=( (not A299)  and  a5095a );
 a5097a <=( a5096a  and  a5091a );
 a5100a <=( A166  and  A168 );
 a5104a <=( A265  and  A200 );
 a5105a <=( (not A199)  and  a5104a );
 a5106a <=( a5105a  and  a5100a );
 a5109a <=( A267  and  (not A266) );
 a5113a <=( (not A300)  and  A298 );
 a5114a <=( A268  and  a5113a );
 a5115a <=( a5114a  and  a5109a );
 a5118a <=( A166  and  A168 );
 a5122a <=( A265  and  A200 );
 a5123a <=( (not A199)  and  a5122a );
 a5124a <=( a5123a  and  a5118a );
 a5127a <=( A267  and  (not A266) );
 a5131a <=( A299  and  A298 );
 a5132a <=( A268  and  a5131a );
 a5133a <=( a5132a  and  a5127a );
 a5136a <=( A166  and  A168 );
 a5140a <=( A265  and  A200 );
 a5141a <=( (not A199)  and  a5140a );
 a5142a <=( a5141a  and  a5136a );
 a5145a <=( A267  and  (not A266) );
 a5149a <=( (not A299)  and  (not A298) );
 a5150a <=( A268  and  a5149a );
 a5151a <=( a5150a  and  a5145a );
 a5154a <=( A166  and  A168 );
 a5158a <=( A265  and  A200 );
 a5159a <=( (not A199)  and  a5158a );
 a5160a <=( a5159a  and  a5154a );
 a5163a <=( A267  and  (not A266) );
 a5167a <=( (not A300)  and  A298 );
 a5168a <=( A269  and  a5167a );
 a5169a <=( a5168a  and  a5163a );
 a5172a <=( A166  and  A168 );
 a5176a <=( A265  and  A200 );
 a5177a <=( (not A199)  and  a5176a );
 a5178a <=( a5177a  and  a5172a );
 a5181a <=( A267  and  (not A266) );
 a5185a <=( A299  and  A298 );
 a5186a <=( A269  and  a5185a );
 a5187a <=( a5186a  and  a5181a );
 a5190a <=( A166  and  A168 );
 a5194a <=( A265  and  A200 );
 a5195a <=( (not A199)  and  a5194a );
 a5196a <=( a5195a  and  a5190a );
 a5199a <=( A267  and  (not A266) );
 a5203a <=( (not A299)  and  (not A298) );
 a5204a <=( A269  and  a5203a );
 a5205a <=( a5204a  and  a5199a );
 a5208a <=( A166  and  A168 );
 a5212a <=( (not A203)  and  (not A202) );
 a5213a <=( (not A200)  and  a5212a );
 a5214a <=( a5213a  and  a5208a );
 a5217a <=( (not A268)  and  (not A266) );
 a5221a <=( A299  and  (not A298) );
 a5222a <=( (not A269)  and  a5221a );
 a5223a <=( a5222a  and  a5217a );
 a5226a <=( A166  and  A168 );
 a5230a <=( A265  and  (not A201) );
 a5231a <=( (not A200)  and  a5230a );
 a5232a <=( a5231a  and  a5226a );
 a5235a <=( A298  and  A266 );
 a5239a <=( A301  and  A300 );
 a5240a <=( (not A299)  and  a5239a );
 a5241a <=( a5240a  and  a5235a );
 a5244a <=( A166  and  A168 );
 a5248a <=( A265  and  (not A201) );
 a5249a <=( (not A200)  and  a5248a );
 a5250a <=( a5249a  and  a5244a );
 a5253a <=( A298  and  A266 );
 a5257a <=( A302  and  A300 );
 a5258a <=( (not A299)  and  a5257a );
 a5259a <=( a5258a  and  a5253a );
 a5262a <=( A166  and  A168 );
 a5266a <=( (not A266)  and  (not A201) );
 a5267a <=( (not A200)  and  a5266a );
 a5268a <=( a5267a  and  a5262a );
 a5271a <=( A298  and  (not A267) );
 a5275a <=( A301  and  A300 );
 a5276a <=( (not A299)  and  a5275a );
 a5277a <=( a5276a  and  a5271a );
 a5280a <=( A166  and  A168 );
 a5284a <=( (not A266)  and  (not A201) );
 a5285a <=( (not A200)  and  a5284a );
 a5286a <=( a5285a  and  a5280a );
 a5289a <=( A298  and  (not A267) );
 a5293a <=( A302  and  A300 );
 a5294a <=( (not A299)  and  a5293a );
 a5295a <=( a5294a  and  a5289a );
 a5298a <=( A166  and  A168 );
 a5302a <=( (not A265)  and  (not A201) );
 a5303a <=( (not A200)  and  a5302a );
 a5304a <=( a5303a  and  a5298a );
 a5307a <=( A298  and  (not A266) );
 a5311a <=( A301  and  A300 );
 a5312a <=( (not A299)  and  a5311a );
 a5313a <=( a5312a  and  a5307a );
 a5316a <=( A166  and  A168 );
 a5320a <=( (not A265)  and  (not A201) );
 a5321a <=( (not A200)  and  a5320a );
 a5322a <=( a5321a  and  a5316a );
 a5325a <=( A298  and  (not A266) );
 a5329a <=( A302  and  A300 );
 a5330a <=( (not A299)  and  a5329a );
 a5331a <=( a5330a  and  a5325a );
 a5334a <=( A166  and  A168 );
 a5338a <=( A201  and  (not A200) );
 a5339a <=( A199  and  a5338a );
 a5340a <=( a5339a  and  a5334a );
 a5343a <=( (not A265)  and  A202 );
 a5347a <=( (not A300)  and  A298 );
 a5348a <=( A266  and  a5347a );
 a5349a <=( a5348a  and  a5343a );
 a5352a <=( A166  and  A168 );
 a5356a <=( A201  and  (not A200) );
 a5357a <=( A199  and  a5356a );
 a5358a <=( a5357a  and  a5352a );
 a5361a <=( (not A265)  and  A202 );
 a5365a <=( A299  and  A298 );
 a5366a <=( A266  and  a5365a );
 a5367a <=( a5366a  and  a5361a );
 a5370a <=( A166  and  A168 );
 a5374a <=( A201  and  (not A200) );
 a5375a <=( A199  and  a5374a );
 a5376a <=( a5375a  and  a5370a );
 a5379a <=( (not A265)  and  A202 );
 a5383a <=( (not A299)  and  (not A298) );
 a5384a <=( A266  and  a5383a );
 a5385a <=( a5384a  and  a5379a );
 a5388a <=( A166  and  A168 );
 a5392a <=( A201  and  (not A200) );
 a5393a <=( A199  and  a5392a );
 a5394a <=( a5393a  and  a5388a );
 a5397a <=( (not A265)  and  A203 );
 a5401a <=( (not A300)  and  A298 );
 a5402a <=( A266  and  a5401a );
 a5403a <=( a5402a  and  a5397a );
 a5406a <=( A166  and  A168 );
 a5410a <=( A201  and  (not A200) );
 a5411a <=( A199  and  a5410a );
 a5412a <=( a5411a  and  a5406a );
 a5415a <=( (not A265)  and  A203 );
 a5419a <=( A299  and  A298 );
 a5420a <=( A266  and  a5419a );
 a5421a <=( a5420a  and  a5415a );
 a5424a <=( A166  and  A168 );
 a5428a <=( A201  and  (not A200) );
 a5429a <=( A199  and  a5428a );
 a5430a <=( a5429a  and  a5424a );
 a5433a <=( (not A265)  and  A203 );
 a5437a <=( (not A299)  and  (not A298) );
 a5438a <=( A266  and  a5437a );
 a5439a <=( a5438a  and  a5433a );
 a5442a <=( A166  and  A168 );
 a5446a <=( A265  and  (not A200) );
 a5447a <=( (not A199)  and  a5446a );
 a5448a <=( a5447a  and  a5442a );
 a5451a <=( A298  and  A266 );
 a5455a <=( A301  and  A300 );
 a5456a <=( (not A299)  and  a5455a );
 a5457a <=( a5456a  and  a5451a );
 a5460a <=( A166  and  A168 );
 a5464a <=( A265  and  (not A200) );
 a5465a <=( (not A199)  and  a5464a );
 a5466a <=( a5465a  and  a5460a );
 a5469a <=( A298  and  A266 );
 a5473a <=( A302  and  A300 );
 a5474a <=( (not A299)  and  a5473a );
 a5475a <=( a5474a  and  a5469a );
 a5478a <=( A166  and  A168 );
 a5482a <=( (not A266)  and  (not A200) );
 a5483a <=( (not A199)  and  a5482a );
 a5484a <=( a5483a  and  a5478a );
 a5487a <=( A298  and  (not A267) );
 a5491a <=( A301  and  A300 );
 a5492a <=( (not A299)  and  a5491a );
 a5493a <=( a5492a  and  a5487a );
 a5496a <=( A166  and  A168 );
 a5500a <=( (not A266)  and  (not A200) );
 a5501a <=( (not A199)  and  a5500a );
 a5502a <=( a5501a  and  a5496a );
 a5505a <=( A298  and  (not A267) );
 a5509a <=( A302  and  A300 );
 a5510a <=( (not A299)  and  a5509a );
 a5511a <=( a5510a  and  a5505a );
 a5514a <=( A166  and  A168 );
 a5518a <=( (not A265)  and  (not A200) );
 a5519a <=( (not A199)  and  a5518a );
 a5520a <=( a5519a  and  a5514a );
 a5523a <=( A298  and  (not A266) );
 a5527a <=( A301  and  A300 );
 a5528a <=( (not A299)  and  a5527a );
 a5529a <=( a5528a  and  a5523a );
 a5532a <=( A166  and  A168 );
 a5536a <=( (not A265)  and  (not A200) );
 a5537a <=( (not A199)  and  a5536a );
 a5538a <=( a5537a  and  a5532a );
 a5541a <=( A298  and  (not A266) );
 a5545a <=( A302  and  A300 );
 a5546a <=( (not A299)  and  a5545a );
 a5547a <=( a5546a  and  a5541a );
 a5550a <=( A167  and  A168 );
 a5554a <=( A265  and  A200 );
 a5555a <=( A199  and  a5554a );
 a5556a <=( a5555a  and  a5550a );
 a5559a <=( A298  and  A266 );
 a5563a <=( A301  and  A300 );
 a5564a <=( (not A299)  and  a5563a );
 a5565a <=( a5564a  and  a5559a );
 a5568a <=( A167  and  A168 );
 a5572a <=( A265  and  A200 );
 a5573a <=( A199  and  a5572a );
 a5574a <=( a5573a  and  a5568a );
 a5577a <=( A298  and  A266 );
 a5581a <=( A302  and  A300 );
 a5582a <=( (not A299)  and  a5581a );
 a5583a <=( a5582a  and  a5577a );
 a5586a <=( A167  and  A168 );
 a5590a <=( (not A266)  and  A200 );
 a5591a <=( A199  and  a5590a );
 a5592a <=( a5591a  and  a5586a );
 a5595a <=( A298  and  (not A267) );
 a5599a <=( A301  and  A300 );
 a5600a <=( (not A299)  and  a5599a );
 a5601a <=( a5600a  and  a5595a );
 a5604a <=( A167  and  A168 );
 a5608a <=( (not A266)  and  A200 );
 a5609a <=( A199  and  a5608a );
 a5610a <=( a5609a  and  a5604a );
 a5613a <=( A298  and  (not A267) );
 a5617a <=( A302  and  A300 );
 a5618a <=( (not A299)  and  a5617a );
 a5619a <=( a5618a  and  a5613a );
 a5622a <=( A167  and  A168 );
 a5626a <=( (not A265)  and  A200 );
 a5627a <=( A199  and  a5626a );
 a5628a <=( a5627a  and  a5622a );
 a5631a <=( A298  and  (not A266) );
 a5635a <=( A301  and  A300 );
 a5636a <=( (not A299)  and  a5635a );
 a5637a <=( a5636a  and  a5631a );
 a5640a <=( A167  and  A168 );
 a5644a <=( (not A265)  and  A200 );
 a5645a <=( A199  and  a5644a );
 a5646a <=( a5645a  and  a5640a );
 a5649a <=( A298  and  (not A266) );
 a5653a <=( A302  and  A300 );
 a5654a <=( (not A299)  and  a5653a );
 a5655a <=( a5654a  and  a5649a );
 a5658a <=( A167  and  A168 );
 a5662a <=( A265  and  A200 );
 a5663a <=( (not A199)  and  a5662a );
 a5664a <=( a5663a  and  a5658a );
 a5667a <=( A267  and  (not A266) );
 a5671a <=( (not A300)  and  A298 );
 a5672a <=( A268  and  a5671a );
 a5673a <=( a5672a  and  a5667a );
 a5676a <=( A167  and  A168 );
 a5680a <=( A265  and  A200 );
 a5681a <=( (not A199)  and  a5680a );
 a5682a <=( a5681a  and  a5676a );
 a5685a <=( A267  and  (not A266) );
 a5689a <=( A299  and  A298 );
 a5690a <=( A268  and  a5689a );
 a5691a <=( a5690a  and  a5685a );
 a5694a <=( A167  and  A168 );
 a5698a <=( A265  and  A200 );
 a5699a <=( (not A199)  and  a5698a );
 a5700a <=( a5699a  and  a5694a );
 a5703a <=( A267  and  (not A266) );
 a5707a <=( (not A299)  and  (not A298) );
 a5708a <=( A268  and  a5707a );
 a5709a <=( a5708a  and  a5703a );
 a5712a <=( A167  and  A168 );
 a5716a <=( A265  and  A200 );
 a5717a <=( (not A199)  and  a5716a );
 a5718a <=( a5717a  and  a5712a );
 a5721a <=( A267  and  (not A266) );
 a5725a <=( (not A300)  and  A298 );
 a5726a <=( A269  and  a5725a );
 a5727a <=( a5726a  and  a5721a );
 a5730a <=( A167  and  A168 );
 a5734a <=( A265  and  A200 );
 a5735a <=( (not A199)  and  a5734a );
 a5736a <=( a5735a  and  a5730a );
 a5739a <=( A267  and  (not A266) );
 a5743a <=( A299  and  A298 );
 a5744a <=( A269  and  a5743a );
 a5745a <=( a5744a  and  a5739a );
 a5748a <=( A167  and  A168 );
 a5752a <=( A265  and  A200 );
 a5753a <=( (not A199)  and  a5752a );
 a5754a <=( a5753a  and  a5748a );
 a5757a <=( A267  and  (not A266) );
 a5761a <=( (not A299)  and  (not A298) );
 a5762a <=( A269  and  a5761a );
 a5763a <=( a5762a  and  a5757a );
 a5766a <=( A167  and  A168 );
 a5770a <=( (not A203)  and  (not A202) );
 a5771a <=( (not A200)  and  a5770a );
 a5772a <=( a5771a  and  a5766a );
 a5775a <=( (not A268)  and  (not A266) );
 a5779a <=( A299  and  (not A298) );
 a5780a <=( (not A269)  and  a5779a );
 a5781a <=( a5780a  and  a5775a );
 a5784a <=( A167  and  A168 );
 a5788a <=( A265  and  (not A201) );
 a5789a <=( (not A200)  and  a5788a );
 a5790a <=( a5789a  and  a5784a );
 a5793a <=( A298  and  A266 );
 a5797a <=( A301  and  A300 );
 a5798a <=( (not A299)  and  a5797a );
 a5799a <=( a5798a  and  a5793a );
 a5802a <=( A167  and  A168 );
 a5806a <=( A265  and  (not A201) );
 a5807a <=( (not A200)  and  a5806a );
 a5808a <=( a5807a  and  a5802a );
 a5811a <=( A298  and  A266 );
 a5815a <=( A302  and  A300 );
 a5816a <=( (not A299)  and  a5815a );
 a5817a <=( a5816a  and  a5811a );
 a5820a <=( A167  and  A168 );
 a5824a <=( (not A266)  and  (not A201) );
 a5825a <=( (not A200)  and  a5824a );
 a5826a <=( a5825a  and  a5820a );
 a5829a <=( A298  and  (not A267) );
 a5833a <=( A301  and  A300 );
 a5834a <=( (not A299)  and  a5833a );
 a5835a <=( a5834a  and  a5829a );
 a5838a <=( A167  and  A168 );
 a5842a <=( (not A266)  and  (not A201) );
 a5843a <=( (not A200)  and  a5842a );
 a5844a <=( a5843a  and  a5838a );
 a5847a <=( A298  and  (not A267) );
 a5851a <=( A302  and  A300 );
 a5852a <=( (not A299)  and  a5851a );
 a5853a <=( a5852a  and  a5847a );
 a5856a <=( A167  and  A168 );
 a5860a <=( (not A265)  and  (not A201) );
 a5861a <=( (not A200)  and  a5860a );
 a5862a <=( a5861a  and  a5856a );
 a5865a <=( A298  and  (not A266) );
 a5869a <=( A301  and  A300 );
 a5870a <=( (not A299)  and  a5869a );
 a5871a <=( a5870a  and  a5865a );
 a5874a <=( A167  and  A168 );
 a5878a <=( (not A265)  and  (not A201) );
 a5879a <=( (not A200)  and  a5878a );
 a5880a <=( a5879a  and  a5874a );
 a5883a <=( A298  and  (not A266) );
 a5887a <=( A302  and  A300 );
 a5888a <=( (not A299)  and  a5887a );
 a5889a <=( a5888a  and  a5883a );
 a5892a <=( A167  and  A168 );
 a5896a <=( A201  and  (not A200) );
 a5897a <=( A199  and  a5896a );
 a5898a <=( a5897a  and  a5892a );
 a5901a <=( (not A265)  and  A202 );
 a5905a <=( (not A300)  and  A298 );
 a5906a <=( A266  and  a5905a );
 a5907a <=( a5906a  and  a5901a );
 a5910a <=( A167  and  A168 );
 a5914a <=( A201  and  (not A200) );
 a5915a <=( A199  and  a5914a );
 a5916a <=( a5915a  and  a5910a );
 a5919a <=( (not A265)  and  A202 );
 a5923a <=( A299  and  A298 );
 a5924a <=( A266  and  a5923a );
 a5925a <=( a5924a  and  a5919a );
 a5928a <=( A167  and  A168 );
 a5932a <=( A201  and  (not A200) );
 a5933a <=( A199  and  a5932a );
 a5934a <=( a5933a  and  a5928a );
 a5937a <=( (not A265)  and  A202 );
 a5941a <=( (not A299)  and  (not A298) );
 a5942a <=( A266  and  a5941a );
 a5943a <=( a5942a  and  a5937a );
 a5946a <=( A167  and  A168 );
 a5950a <=( A201  and  (not A200) );
 a5951a <=( A199  and  a5950a );
 a5952a <=( a5951a  and  a5946a );
 a5955a <=( (not A265)  and  A203 );
 a5959a <=( (not A300)  and  A298 );
 a5960a <=( A266  and  a5959a );
 a5961a <=( a5960a  and  a5955a );
 a5964a <=( A167  and  A168 );
 a5968a <=( A201  and  (not A200) );
 a5969a <=( A199  and  a5968a );
 a5970a <=( a5969a  and  a5964a );
 a5973a <=( (not A265)  and  A203 );
 a5977a <=( A299  and  A298 );
 a5978a <=( A266  and  a5977a );
 a5979a <=( a5978a  and  a5973a );
 a5982a <=( A167  and  A168 );
 a5986a <=( A201  and  (not A200) );
 a5987a <=( A199  and  a5986a );
 a5988a <=( a5987a  and  a5982a );
 a5991a <=( (not A265)  and  A203 );
 a5995a <=( (not A299)  and  (not A298) );
 a5996a <=( A266  and  a5995a );
 a5997a <=( a5996a  and  a5991a );
 a6000a <=( A167  and  A168 );
 a6004a <=( A265  and  (not A200) );
 a6005a <=( (not A199)  and  a6004a );
 a6006a <=( a6005a  and  a6000a );
 a6009a <=( A298  and  A266 );
 a6013a <=( A301  and  A300 );
 a6014a <=( (not A299)  and  a6013a );
 a6015a <=( a6014a  and  a6009a );
 a6018a <=( A167  and  A168 );
 a6022a <=( A265  and  (not A200) );
 a6023a <=( (not A199)  and  a6022a );
 a6024a <=( a6023a  and  a6018a );
 a6027a <=( A298  and  A266 );
 a6031a <=( A302  and  A300 );
 a6032a <=( (not A299)  and  a6031a );
 a6033a <=( a6032a  and  a6027a );
 a6036a <=( A167  and  A168 );
 a6040a <=( (not A266)  and  (not A200) );
 a6041a <=( (not A199)  and  a6040a );
 a6042a <=( a6041a  and  a6036a );
 a6045a <=( A298  and  (not A267) );
 a6049a <=( A301  and  A300 );
 a6050a <=( (not A299)  and  a6049a );
 a6051a <=( a6050a  and  a6045a );
 a6054a <=( A167  and  A168 );
 a6058a <=( (not A266)  and  (not A200) );
 a6059a <=( (not A199)  and  a6058a );
 a6060a <=( a6059a  and  a6054a );
 a6063a <=( A298  and  (not A267) );
 a6067a <=( A302  and  A300 );
 a6068a <=( (not A299)  and  a6067a );
 a6069a <=( a6068a  and  a6063a );
 a6072a <=( A167  and  A168 );
 a6076a <=( (not A265)  and  (not A200) );
 a6077a <=( (not A199)  and  a6076a );
 a6078a <=( a6077a  and  a6072a );
 a6081a <=( A298  and  (not A266) );
 a6085a <=( A301  and  A300 );
 a6086a <=( (not A299)  and  a6085a );
 a6087a <=( a6086a  and  a6081a );
 a6090a <=( A167  and  A168 );
 a6094a <=( (not A265)  and  (not A200) );
 a6095a <=( (not A199)  and  a6094a );
 a6096a <=( a6095a  and  a6090a );
 a6099a <=( A298  and  (not A266) );
 a6103a <=( A302  and  A300 );
 a6104a <=( (not A299)  and  a6103a );
 a6105a <=( a6104a  and  a6099a );
 a6108a <=( (not A167)  and  A170 );
 a6112a <=( A200  and  A199 );
 a6113a <=( (not A166)  and  a6112a );
 a6114a <=( a6113a  and  a6108a );
 a6117a <=( A266  and  (not A265) );
 a6121a <=( (not A302)  and  (not A301) );
 a6122a <=( A298  and  a6121a );
 a6123a <=( a6122a  and  a6117a );
 a6126a <=( (not A167)  and  A170 );
 a6130a <=( A200  and  (not A199) );
 a6131a <=( (not A166)  and  a6130a );
 a6132a <=( a6131a  and  a6126a );
 a6135a <=( (not A268)  and  (not A266) );
 a6139a <=( A299  and  (not A298) );
 a6140a <=( (not A269)  and  a6139a );
 a6141a <=( a6140a  and  a6135a );
 a6144a <=( (not A167)  and  A170 );
 a6148a <=( (not A202)  and  (not A200) );
 a6149a <=( (not A166)  and  a6148a );
 a6150a <=( a6149a  and  a6144a );
 a6153a <=( (not A265)  and  (not A203) );
 a6157a <=( (not A300)  and  A298 );
 a6158a <=( A266  and  a6157a );
 a6159a <=( a6158a  and  a6153a );
 a6162a <=( (not A167)  and  A170 );
 a6166a <=( (not A202)  and  (not A200) );
 a6167a <=( (not A166)  and  a6166a );
 a6168a <=( a6167a  and  a6162a );
 a6171a <=( (not A265)  and  (not A203) );
 a6175a <=( A299  and  A298 );
 a6176a <=( A266  and  a6175a );
 a6177a <=( a6176a  and  a6171a );
 a6180a <=( (not A167)  and  A170 );
 a6184a <=( (not A202)  and  (not A200) );
 a6185a <=( (not A166)  and  a6184a );
 a6186a <=( a6185a  and  a6180a );
 a6189a <=( (not A265)  and  (not A203) );
 a6193a <=( (not A299)  and  (not A298) );
 a6194a <=( A266  and  a6193a );
 a6195a <=( a6194a  and  a6189a );
 a6198a <=( (not A167)  and  A170 );
 a6202a <=( (not A201)  and  (not A200) );
 a6203a <=( (not A166)  and  a6202a );
 a6204a <=( a6203a  and  a6198a );
 a6207a <=( A266  and  (not A265) );
 a6211a <=( (not A302)  and  (not A301) );
 a6212a <=( A298  and  a6211a );
 a6213a <=( a6212a  and  a6207a );
 a6216a <=( (not A167)  and  A170 );
 a6220a <=( (not A200)  and  (not A199) );
 a6221a <=( (not A166)  and  a6220a );
 a6222a <=( a6221a  and  a6216a );
 a6225a <=( A266  and  (not A265) );
 a6229a <=( (not A302)  and  (not A301) );
 a6230a <=( A298  and  a6229a );
 a6231a <=( a6230a  and  a6225a );
 a6234a <=( (not A168)  and  A169 );
 a6238a <=( A199  and  (not A166) );
 a6239a <=( A167  and  a6238a );
 a6240a <=( a6239a  and  a6234a );
 a6243a <=( (not A265)  and  A200 );
 a6247a <=( (not A300)  and  A298 );
 a6248a <=( A266  and  a6247a );
 a6249a <=( a6248a  and  a6243a );
 a6252a <=( (not A168)  and  A169 );
 a6256a <=( A199  and  (not A166) );
 a6257a <=( A167  and  a6256a );
 a6258a <=( a6257a  and  a6252a );
 a6261a <=( (not A265)  and  A200 );
 a6265a <=( A299  and  A298 );
 a6266a <=( A266  and  a6265a );
 a6267a <=( a6266a  and  a6261a );
 a6270a <=( (not A168)  and  A169 );
 a6274a <=( A199  and  (not A166) );
 a6275a <=( A167  and  a6274a );
 a6276a <=( a6275a  and  a6270a );
 a6279a <=( (not A265)  and  A200 );
 a6283a <=( (not A299)  and  (not A298) );
 a6284a <=( A266  and  a6283a );
 a6285a <=( a6284a  and  a6279a );
 a6288a <=( (not A168)  and  A169 );
 a6292a <=( (not A199)  and  (not A166) );
 a6293a <=( A167  and  a6292a );
 a6294a <=( a6293a  and  a6288a );
 a6297a <=( A265  and  A200 );
 a6301a <=( A299  and  (not A298) );
 a6302a <=( A266  and  a6301a );
 a6303a <=( a6302a  and  a6297a );
 a6306a <=( (not A168)  and  A169 );
 a6310a <=( (not A199)  and  (not A166) );
 a6311a <=( A167  and  a6310a );
 a6312a <=( a6311a  and  a6306a );
 a6315a <=( (not A266)  and  A200 );
 a6319a <=( A299  and  (not A298) );
 a6320a <=( (not A267)  and  a6319a );
 a6321a <=( a6320a  and  a6315a );
 a6324a <=( (not A168)  and  A169 );
 a6328a <=( (not A199)  and  (not A166) );
 a6329a <=( A167  and  a6328a );
 a6330a <=( a6329a  and  a6324a );
 a6333a <=( (not A265)  and  A200 );
 a6337a <=( A299  and  (not A298) );
 a6338a <=( (not A266)  and  a6337a );
 a6339a <=( a6338a  and  a6333a );
 a6342a <=( (not A168)  and  A169 );
 a6346a <=( (not A200)  and  (not A166) );
 a6347a <=( A167  and  a6346a );
 a6348a <=( a6347a  and  a6342a );
 a6351a <=( (not A265)  and  (not A201) );
 a6355a <=( (not A300)  and  A298 );
 a6356a <=( A266  and  a6355a );
 a6357a <=( a6356a  and  a6351a );
 a6360a <=( (not A168)  and  A169 );
 a6364a <=( (not A200)  and  (not A166) );
 a6365a <=( A167  and  a6364a );
 a6366a <=( a6365a  and  a6360a );
 a6369a <=( (not A265)  and  (not A201) );
 a6373a <=( A299  and  A298 );
 a6374a <=( A266  and  a6373a );
 a6375a <=( a6374a  and  a6369a );
 a6378a <=( (not A168)  and  A169 );
 a6382a <=( (not A200)  and  (not A166) );
 a6383a <=( A167  and  a6382a );
 a6384a <=( a6383a  and  a6378a );
 a6387a <=( (not A265)  and  (not A201) );
 a6391a <=( (not A299)  and  (not A298) );
 a6392a <=( A266  and  a6391a );
 a6393a <=( a6392a  and  a6387a );
 a6396a <=( (not A168)  and  A169 );
 a6400a <=( (not A199)  and  (not A166) );
 a6401a <=( A167  and  a6400a );
 a6402a <=( a6401a  and  a6396a );
 a6405a <=( (not A265)  and  (not A200) );
 a6409a <=( (not A300)  and  A298 );
 a6410a <=( A266  and  a6409a );
 a6411a <=( a6410a  and  a6405a );
 a6414a <=( (not A168)  and  A169 );
 a6418a <=( (not A199)  and  (not A166) );
 a6419a <=( A167  and  a6418a );
 a6420a <=( a6419a  and  a6414a );
 a6423a <=( (not A265)  and  (not A200) );
 a6427a <=( A299  and  A298 );
 a6428a <=( A266  and  a6427a );
 a6429a <=( a6428a  and  a6423a );
 a6432a <=( (not A168)  and  A169 );
 a6436a <=( (not A199)  and  (not A166) );
 a6437a <=( A167  and  a6436a );
 a6438a <=( a6437a  and  a6432a );
 a6441a <=( (not A265)  and  (not A200) );
 a6445a <=( (not A299)  and  (not A298) );
 a6446a <=( A266  and  a6445a );
 a6447a <=( a6446a  and  a6441a );
 a6450a <=( (not A168)  and  A169 );
 a6454a <=( A199  and  A166 );
 a6455a <=( (not A167)  and  a6454a );
 a6456a <=( a6455a  and  a6450a );
 a6459a <=( (not A265)  and  A200 );
 a6463a <=( (not A300)  and  A298 );
 a6464a <=( A266  and  a6463a );
 a6465a <=( a6464a  and  a6459a );
 a6468a <=( (not A168)  and  A169 );
 a6472a <=( A199  and  A166 );
 a6473a <=( (not A167)  and  a6472a );
 a6474a <=( a6473a  and  a6468a );
 a6477a <=( (not A265)  and  A200 );
 a6481a <=( A299  and  A298 );
 a6482a <=( A266  and  a6481a );
 a6483a <=( a6482a  and  a6477a );
 a6486a <=( (not A168)  and  A169 );
 a6490a <=( A199  and  A166 );
 a6491a <=( (not A167)  and  a6490a );
 a6492a <=( a6491a  and  a6486a );
 a6495a <=( (not A265)  and  A200 );
 a6499a <=( (not A299)  and  (not A298) );
 a6500a <=( A266  and  a6499a );
 a6501a <=( a6500a  and  a6495a );
 a6504a <=( (not A168)  and  A169 );
 a6508a <=( (not A199)  and  A166 );
 a6509a <=( (not A167)  and  a6508a );
 a6510a <=( a6509a  and  a6504a );
 a6513a <=( A265  and  A200 );
 a6517a <=( A299  and  (not A298) );
 a6518a <=( A266  and  a6517a );
 a6519a <=( a6518a  and  a6513a );
 a6522a <=( (not A168)  and  A169 );
 a6526a <=( (not A199)  and  A166 );
 a6527a <=( (not A167)  and  a6526a );
 a6528a <=( a6527a  and  a6522a );
 a6531a <=( (not A266)  and  A200 );
 a6535a <=( A299  and  (not A298) );
 a6536a <=( (not A267)  and  a6535a );
 a6537a <=( a6536a  and  a6531a );
 a6540a <=( (not A168)  and  A169 );
 a6544a <=( (not A199)  and  A166 );
 a6545a <=( (not A167)  and  a6544a );
 a6546a <=( a6545a  and  a6540a );
 a6549a <=( (not A265)  and  A200 );
 a6553a <=( A299  and  (not A298) );
 a6554a <=( (not A266)  and  a6553a );
 a6555a <=( a6554a  and  a6549a );
 a6558a <=( (not A168)  and  A169 );
 a6562a <=( (not A200)  and  A166 );
 a6563a <=( (not A167)  and  a6562a );
 a6564a <=( a6563a  and  a6558a );
 a6567a <=( (not A265)  and  (not A201) );
 a6571a <=( (not A300)  and  A298 );
 a6572a <=( A266  and  a6571a );
 a6573a <=( a6572a  and  a6567a );
 a6576a <=( (not A168)  and  A169 );
 a6580a <=( (not A200)  and  A166 );
 a6581a <=( (not A167)  and  a6580a );
 a6582a <=( a6581a  and  a6576a );
 a6585a <=( (not A265)  and  (not A201) );
 a6589a <=( A299  and  A298 );
 a6590a <=( A266  and  a6589a );
 a6591a <=( a6590a  and  a6585a );
 a6594a <=( (not A168)  and  A169 );
 a6598a <=( (not A200)  and  A166 );
 a6599a <=( (not A167)  and  a6598a );
 a6600a <=( a6599a  and  a6594a );
 a6603a <=( (not A265)  and  (not A201) );
 a6607a <=( (not A299)  and  (not A298) );
 a6608a <=( A266  and  a6607a );
 a6609a <=( a6608a  and  a6603a );
 a6612a <=( (not A168)  and  A169 );
 a6616a <=( (not A199)  and  A166 );
 a6617a <=( (not A167)  and  a6616a );
 a6618a <=( a6617a  and  a6612a );
 a6621a <=( (not A265)  and  (not A200) );
 a6625a <=( (not A300)  and  A298 );
 a6626a <=( A266  and  a6625a );
 a6627a <=( a6626a  and  a6621a );
 a6630a <=( (not A168)  and  A169 );
 a6634a <=( (not A199)  and  A166 );
 a6635a <=( (not A167)  and  a6634a );
 a6636a <=( a6635a  and  a6630a );
 a6639a <=( (not A265)  and  (not A200) );
 a6643a <=( A299  and  A298 );
 a6644a <=( A266  and  a6643a );
 a6645a <=( a6644a  and  a6639a );
 a6648a <=( (not A168)  and  A169 );
 a6652a <=( (not A199)  and  A166 );
 a6653a <=( (not A167)  and  a6652a );
 a6654a <=( a6653a  and  a6648a );
 a6657a <=( (not A265)  and  (not A200) );
 a6661a <=( (not A299)  and  (not A298) );
 a6662a <=( A266  and  a6661a );
 a6663a <=( a6662a  and  a6657a );
 a6666a <=( A169  and  A170 );
 a6670a <=( A200  and  A199 );
 a6671a <=( (not A168)  and  a6670a );
 a6672a <=( a6671a  and  a6666a );
 a6675a <=( A266  and  (not A265) );
 a6679a <=( (not A302)  and  (not A301) );
 a6680a <=( A298  and  a6679a );
 a6681a <=( a6680a  and  a6675a );
 a6684a <=( A169  and  A170 );
 a6688a <=( A200  and  (not A199) );
 a6689a <=( (not A168)  and  a6688a );
 a6690a <=( a6689a  and  a6684a );
 a6693a <=( (not A268)  and  (not A266) );
 a6697a <=( A299  and  (not A298) );
 a6698a <=( (not A269)  and  a6697a );
 a6699a <=( a6698a  and  a6693a );
 a6702a <=( A169  and  A170 );
 a6706a <=( (not A202)  and  (not A200) );
 a6707a <=( (not A168)  and  a6706a );
 a6708a <=( a6707a  and  a6702a );
 a6711a <=( (not A265)  and  (not A203) );
 a6715a <=( (not A300)  and  A298 );
 a6716a <=( A266  and  a6715a );
 a6717a <=( a6716a  and  a6711a );
 a6720a <=( A169  and  A170 );
 a6724a <=( (not A202)  and  (not A200) );
 a6725a <=( (not A168)  and  a6724a );
 a6726a <=( a6725a  and  a6720a );
 a6729a <=( (not A265)  and  (not A203) );
 a6733a <=( A299  and  A298 );
 a6734a <=( A266  and  a6733a );
 a6735a <=( a6734a  and  a6729a );
 a6738a <=( A169  and  A170 );
 a6742a <=( (not A202)  and  (not A200) );
 a6743a <=( (not A168)  and  a6742a );
 a6744a <=( a6743a  and  a6738a );
 a6747a <=( (not A265)  and  (not A203) );
 a6751a <=( (not A299)  and  (not A298) );
 a6752a <=( A266  and  a6751a );
 a6753a <=( a6752a  and  a6747a );
 a6756a <=( A169  and  A170 );
 a6760a <=( (not A201)  and  (not A200) );
 a6761a <=( (not A168)  and  a6760a );
 a6762a <=( a6761a  and  a6756a );
 a6765a <=( A266  and  (not A265) );
 a6769a <=( (not A302)  and  (not A301) );
 a6770a <=( A298  and  a6769a );
 a6771a <=( a6770a  and  a6765a );
 a6774a <=( A169  and  A170 );
 a6778a <=( (not A200)  and  (not A199) );
 a6779a <=( (not A168)  and  a6778a );
 a6780a <=( a6779a  and  a6774a );
 a6783a <=( A266  and  (not A265) );
 a6787a <=( (not A302)  and  (not A301) );
 a6788a <=( A298  and  a6787a );
 a6789a <=( a6788a  and  a6783a );
 a6792a <=( A169  and  (not A170) );
 a6796a <=( A199  and  A166 );
 a6797a <=( A167  and  a6796a );
 a6798a <=( a6797a  and  a6792a );
 a6801a <=( A265  and  A200 );
 a6805a <=( A299  and  (not A298) );
 a6806a <=( A266  and  a6805a );
 a6807a <=( a6806a  and  a6801a );
 a6810a <=( A169  and  (not A170) );
 a6814a <=( A199  and  A166 );
 a6815a <=( A167  and  a6814a );
 a6816a <=( a6815a  and  a6810a );
 a6819a <=( (not A266)  and  A200 );
 a6823a <=( A299  and  (not A298) );
 a6824a <=( (not A267)  and  a6823a );
 a6825a <=( a6824a  and  a6819a );
 a6828a <=( A169  and  (not A170) );
 a6832a <=( A199  and  A166 );
 a6833a <=( A167  and  a6832a );
 a6834a <=( a6833a  and  a6828a );
 a6837a <=( (not A265)  and  A200 );
 a6841a <=( A299  and  (not A298) );
 a6842a <=( (not A266)  and  a6841a );
 a6843a <=( a6842a  and  a6837a );
 a6846a <=( A169  and  (not A170) );
 a6850a <=( (not A199)  and  A166 );
 a6851a <=( A167  and  a6850a );
 a6852a <=( a6851a  and  a6846a );
 a6855a <=( (not A265)  and  A200 );
 a6859a <=( (not A300)  and  A298 );
 a6860a <=( A266  and  a6859a );
 a6861a <=( a6860a  and  a6855a );
 a6864a <=( A169  and  (not A170) );
 a6868a <=( (not A199)  and  A166 );
 a6869a <=( A167  and  a6868a );
 a6870a <=( a6869a  and  a6864a );
 a6873a <=( (not A265)  and  A200 );
 a6877a <=( A299  and  A298 );
 a6878a <=( A266  and  a6877a );
 a6879a <=( a6878a  and  a6873a );
 a6882a <=( A169  and  (not A170) );
 a6886a <=( (not A199)  and  A166 );
 a6887a <=( A167  and  a6886a );
 a6888a <=( a6887a  and  a6882a );
 a6891a <=( (not A265)  and  A200 );
 a6895a <=( (not A299)  and  (not A298) );
 a6896a <=( A266  and  a6895a );
 a6897a <=( a6896a  and  a6891a );
 a6900a <=( A169  and  (not A170) );
 a6904a <=( (not A200)  and  A166 );
 a6905a <=( A167  and  a6904a );
 a6906a <=( a6905a  and  a6900a );
 a6909a <=( A265  and  (not A201) );
 a6913a <=( A299  and  (not A298) );
 a6914a <=( A266  and  a6913a );
 a6915a <=( a6914a  and  a6909a );
 a6918a <=( A169  and  (not A170) );
 a6922a <=( (not A200)  and  A166 );
 a6923a <=( A167  and  a6922a );
 a6924a <=( a6923a  and  a6918a );
 a6927a <=( (not A266)  and  (not A201) );
 a6931a <=( A299  and  (not A298) );
 a6932a <=( (not A267)  and  a6931a );
 a6933a <=( a6932a  and  a6927a );
 a6936a <=( A169  and  (not A170) );
 a6940a <=( (not A200)  and  A166 );
 a6941a <=( A167  and  a6940a );
 a6942a <=( a6941a  and  a6936a );
 a6945a <=( (not A265)  and  (not A201) );
 a6949a <=( A299  and  (not A298) );
 a6950a <=( (not A266)  and  a6949a );
 a6951a <=( a6950a  and  a6945a );
 a6954a <=( A169  and  (not A170) );
 a6958a <=( (not A199)  and  A166 );
 a6959a <=( A167  and  a6958a );
 a6960a <=( a6959a  and  a6954a );
 a6963a <=( A265  and  (not A200) );
 a6967a <=( A299  and  (not A298) );
 a6968a <=( A266  and  a6967a );
 a6969a <=( a6968a  and  a6963a );
 a6972a <=( A169  and  (not A170) );
 a6976a <=( (not A199)  and  A166 );
 a6977a <=( A167  and  a6976a );
 a6978a <=( a6977a  and  a6972a );
 a6981a <=( (not A266)  and  (not A200) );
 a6985a <=( A299  and  (not A298) );
 a6986a <=( (not A267)  and  a6985a );
 a6987a <=( a6986a  and  a6981a );
 a6990a <=( A169  and  (not A170) );
 a6994a <=( (not A199)  and  A166 );
 a6995a <=( A167  and  a6994a );
 a6996a <=( a6995a  and  a6990a );
 a6999a <=( (not A265)  and  (not A200) );
 a7003a <=( A299  and  (not A298) );
 a7004a <=( (not A266)  and  a7003a );
 a7005a <=( a7004a  and  a6999a );
 a7008a <=( A169  and  (not A170) );
 a7012a <=( A199  and  (not A166) );
 a7013a <=( (not A167)  and  a7012a );
 a7014a <=( a7013a  and  a7008a );
 a7017a <=( A265  and  A200 );
 a7021a <=( A299  and  (not A298) );
 a7022a <=( A266  and  a7021a );
 a7023a <=( a7022a  and  a7017a );
 a7026a <=( A169  and  (not A170) );
 a7030a <=( A199  and  (not A166) );
 a7031a <=( (not A167)  and  a7030a );
 a7032a <=( a7031a  and  a7026a );
 a7035a <=( (not A266)  and  A200 );
 a7039a <=( A299  and  (not A298) );
 a7040a <=( (not A267)  and  a7039a );
 a7041a <=( a7040a  and  a7035a );
 a7044a <=( A169  and  (not A170) );
 a7048a <=( A199  and  (not A166) );
 a7049a <=( (not A167)  and  a7048a );
 a7050a <=( a7049a  and  a7044a );
 a7053a <=( (not A265)  and  A200 );
 a7057a <=( A299  and  (not A298) );
 a7058a <=( (not A266)  and  a7057a );
 a7059a <=( a7058a  and  a7053a );
 a7062a <=( A169  and  (not A170) );
 a7066a <=( (not A199)  and  (not A166) );
 a7067a <=( (not A167)  and  a7066a );
 a7068a <=( a7067a  and  a7062a );
 a7071a <=( (not A265)  and  A200 );
 a7075a <=( (not A300)  and  A298 );
 a7076a <=( A266  and  a7075a );
 a7077a <=( a7076a  and  a7071a );
 a7080a <=( A169  and  (not A170) );
 a7084a <=( (not A199)  and  (not A166) );
 a7085a <=( (not A167)  and  a7084a );
 a7086a <=( a7085a  and  a7080a );
 a7089a <=( (not A265)  and  A200 );
 a7093a <=( A299  and  A298 );
 a7094a <=( A266  and  a7093a );
 a7095a <=( a7094a  and  a7089a );
 a7098a <=( A169  and  (not A170) );
 a7102a <=( (not A199)  and  (not A166) );
 a7103a <=( (not A167)  and  a7102a );
 a7104a <=( a7103a  and  a7098a );
 a7107a <=( (not A265)  and  A200 );
 a7111a <=( (not A299)  and  (not A298) );
 a7112a <=( A266  and  a7111a );
 a7113a <=( a7112a  and  a7107a );
 a7116a <=( A169  and  (not A170) );
 a7120a <=( (not A200)  and  (not A166) );
 a7121a <=( (not A167)  and  a7120a );
 a7122a <=( a7121a  and  a7116a );
 a7125a <=( A265  and  (not A201) );
 a7129a <=( A299  and  (not A298) );
 a7130a <=( A266  and  a7129a );
 a7131a <=( a7130a  and  a7125a );
 a7134a <=( A169  and  (not A170) );
 a7138a <=( (not A200)  and  (not A166) );
 a7139a <=( (not A167)  and  a7138a );
 a7140a <=( a7139a  and  a7134a );
 a7143a <=( (not A266)  and  (not A201) );
 a7147a <=( A299  and  (not A298) );
 a7148a <=( (not A267)  and  a7147a );
 a7149a <=( a7148a  and  a7143a );
 a7152a <=( A169  and  (not A170) );
 a7156a <=( (not A200)  and  (not A166) );
 a7157a <=( (not A167)  and  a7156a );
 a7158a <=( a7157a  and  a7152a );
 a7161a <=( (not A265)  and  (not A201) );
 a7165a <=( A299  and  (not A298) );
 a7166a <=( (not A266)  and  a7165a );
 a7167a <=( a7166a  and  a7161a );
 a7170a <=( A169  and  (not A170) );
 a7174a <=( (not A199)  and  (not A166) );
 a7175a <=( (not A167)  and  a7174a );
 a7176a <=( a7175a  and  a7170a );
 a7179a <=( A265  and  (not A200) );
 a7183a <=( A299  and  (not A298) );
 a7184a <=( A266  and  a7183a );
 a7185a <=( a7184a  and  a7179a );
 a7188a <=( A169  and  (not A170) );
 a7192a <=( (not A199)  and  (not A166) );
 a7193a <=( (not A167)  and  a7192a );
 a7194a <=( a7193a  and  a7188a );
 a7197a <=( (not A266)  and  (not A200) );
 a7201a <=( A299  and  (not A298) );
 a7202a <=( (not A267)  and  a7201a );
 a7203a <=( a7202a  and  a7197a );
 a7206a <=( A169  and  (not A170) );
 a7210a <=( (not A199)  and  (not A166) );
 a7211a <=( (not A167)  and  a7210a );
 a7212a <=( a7211a  and  a7206a );
 a7215a <=( (not A265)  and  (not A200) );
 a7219a <=( A299  and  (not A298) );
 a7220a <=( (not A266)  and  a7219a );
 a7221a <=( a7220a  and  a7215a );
 a7224a <=( (not A167)  and  (not A169) );
 a7228a <=( A200  and  A199 );
 a7229a <=( (not A166)  and  a7228a );
 a7230a <=( a7229a  and  a7224a );
 a7233a <=( A266  and  (not A265) );
 a7237a <=( (not A302)  and  (not A301) );
 a7238a <=( A298  and  a7237a );
 a7239a <=( a7238a  and  a7233a );
 a7242a <=( (not A167)  and  (not A169) );
 a7246a <=( A200  and  (not A199) );
 a7247a <=( (not A166)  and  a7246a );
 a7248a <=( a7247a  and  a7242a );
 a7251a <=( (not A268)  and  (not A266) );
 a7255a <=( A299  and  (not A298) );
 a7256a <=( (not A269)  and  a7255a );
 a7257a <=( a7256a  and  a7251a );
 a7260a <=( (not A167)  and  (not A169) );
 a7264a <=( (not A202)  and  (not A200) );
 a7265a <=( (not A166)  and  a7264a );
 a7266a <=( a7265a  and  a7260a );
 a7269a <=( (not A265)  and  (not A203) );
 a7273a <=( (not A300)  and  A298 );
 a7274a <=( A266  and  a7273a );
 a7275a <=( a7274a  and  a7269a );
 a7278a <=( (not A167)  and  (not A169) );
 a7282a <=( (not A202)  and  (not A200) );
 a7283a <=( (not A166)  and  a7282a );
 a7284a <=( a7283a  and  a7278a );
 a7287a <=( (not A265)  and  (not A203) );
 a7291a <=( A299  and  A298 );
 a7292a <=( A266  and  a7291a );
 a7293a <=( a7292a  and  a7287a );
 a7296a <=( (not A167)  and  (not A169) );
 a7300a <=( (not A202)  and  (not A200) );
 a7301a <=( (not A166)  and  a7300a );
 a7302a <=( a7301a  and  a7296a );
 a7305a <=( (not A265)  and  (not A203) );
 a7309a <=( (not A299)  and  (not A298) );
 a7310a <=( A266  and  a7309a );
 a7311a <=( a7310a  and  a7305a );
 a7314a <=( (not A167)  and  (not A169) );
 a7318a <=( (not A201)  and  (not A200) );
 a7319a <=( (not A166)  and  a7318a );
 a7320a <=( a7319a  and  a7314a );
 a7323a <=( A266  and  (not A265) );
 a7327a <=( (not A302)  and  (not A301) );
 a7328a <=( A298  and  a7327a );
 a7329a <=( a7328a  and  a7323a );
 a7332a <=( (not A167)  and  (not A169) );
 a7336a <=( (not A200)  and  (not A199) );
 a7337a <=( (not A166)  and  a7336a );
 a7338a <=( a7337a  and  a7332a );
 a7341a <=( A266  and  (not A265) );
 a7345a <=( (not A302)  and  (not A301) );
 a7346a <=( A298  and  a7345a );
 a7347a <=( a7346a  and  a7341a );
 a7350a <=( (not A168)  and  (not A169) );
 a7354a <=( A199  and  A166 );
 a7355a <=( A167  and  a7354a );
 a7356a <=( a7355a  and  a7350a );
 a7359a <=( (not A265)  and  A200 );
 a7363a <=( (not A300)  and  A298 );
 a7364a <=( A266  and  a7363a );
 a7365a <=( a7364a  and  a7359a );
 a7368a <=( (not A168)  and  (not A169) );
 a7372a <=( A199  and  A166 );
 a7373a <=( A167  and  a7372a );
 a7374a <=( a7373a  and  a7368a );
 a7377a <=( (not A265)  and  A200 );
 a7381a <=( A299  and  A298 );
 a7382a <=( A266  and  a7381a );
 a7383a <=( a7382a  and  a7377a );
 a7386a <=( (not A168)  and  (not A169) );
 a7390a <=( A199  and  A166 );
 a7391a <=( A167  and  a7390a );
 a7392a <=( a7391a  and  a7386a );
 a7395a <=( (not A265)  and  A200 );
 a7399a <=( (not A299)  and  (not A298) );
 a7400a <=( A266  and  a7399a );
 a7401a <=( a7400a  and  a7395a );
 a7404a <=( (not A168)  and  (not A169) );
 a7408a <=( (not A199)  and  A166 );
 a7409a <=( A167  and  a7408a );
 a7410a <=( a7409a  and  a7404a );
 a7413a <=( A265  and  A200 );
 a7417a <=( A299  and  (not A298) );
 a7418a <=( A266  and  a7417a );
 a7419a <=( a7418a  and  a7413a );
 a7422a <=( (not A168)  and  (not A169) );
 a7426a <=( (not A199)  and  A166 );
 a7427a <=( A167  and  a7426a );
 a7428a <=( a7427a  and  a7422a );
 a7431a <=( (not A266)  and  A200 );
 a7435a <=( A299  and  (not A298) );
 a7436a <=( (not A267)  and  a7435a );
 a7437a <=( a7436a  and  a7431a );
 a7440a <=( (not A168)  and  (not A169) );
 a7444a <=( (not A199)  and  A166 );
 a7445a <=( A167  and  a7444a );
 a7446a <=( a7445a  and  a7440a );
 a7449a <=( (not A265)  and  A200 );
 a7453a <=( A299  and  (not A298) );
 a7454a <=( (not A266)  and  a7453a );
 a7455a <=( a7454a  and  a7449a );
 a7458a <=( (not A168)  and  (not A169) );
 a7462a <=( (not A200)  and  A166 );
 a7463a <=( A167  and  a7462a );
 a7464a <=( a7463a  and  a7458a );
 a7467a <=( (not A265)  and  (not A201) );
 a7471a <=( (not A300)  and  A298 );
 a7472a <=( A266  and  a7471a );
 a7473a <=( a7472a  and  a7467a );
 a7476a <=( (not A168)  and  (not A169) );
 a7480a <=( (not A200)  and  A166 );
 a7481a <=( A167  and  a7480a );
 a7482a <=( a7481a  and  a7476a );
 a7485a <=( (not A265)  and  (not A201) );
 a7489a <=( A299  and  A298 );
 a7490a <=( A266  and  a7489a );
 a7491a <=( a7490a  and  a7485a );
 a7494a <=( (not A168)  and  (not A169) );
 a7498a <=( (not A200)  and  A166 );
 a7499a <=( A167  and  a7498a );
 a7500a <=( a7499a  and  a7494a );
 a7503a <=( (not A265)  and  (not A201) );
 a7507a <=( (not A299)  and  (not A298) );
 a7508a <=( A266  and  a7507a );
 a7509a <=( a7508a  and  a7503a );
 a7512a <=( (not A168)  and  (not A169) );
 a7516a <=( (not A199)  and  A166 );
 a7517a <=( A167  and  a7516a );
 a7518a <=( a7517a  and  a7512a );
 a7521a <=( (not A265)  and  (not A200) );
 a7525a <=( (not A300)  and  A298 );
 a7526a <=( A266  and  a7525a );
 a7527a <=( a7526a  and  a7521a );
 a7530a <=( (not A168)  and  (not A169) );
 a7534a <=( (not A199)  and  A166 );
 a7535a <=( A167  and  a7534a );
 a7536a <=( a7535a  and  a7530a );
 a7539a <=( (not A265)  and  (not A200) );
 a7543a <=( A299  and  A298 );
 a7544a <=( A266  and  a7543a );
 a7545a <=( a7544a  and  a7539a );
 a7548a <=( (not A168)  and  (not A169) );
 a7552a <=( (not A199)  and  A166 );
 a7553a <=( A167  and  a7552a );
 a7554a <=( a7553a  and  a7548a );
 a7557a <=( (not A265)  and  (not A200) );
 a7561a <=( (not A299)  and  (not A298) );
 a7562a <=( A266  and  a7561a );
 a7563a <=( a7562a  and  a7557a );
 a7566a <=( (not A169)  and  A170 );
 a7570a <=( A199  and  (not A166) );
 a7571a <=( A167  and  a7570a );
 a7572a <=( a7571a  and  a7566a );
 a7575a <=( A265  and  A200 );
 a7579a <=( A299  and  (not A298) );
 a7580a <=( A266  and  a7579a );
 a7581a <=( a7580a  and  a7575a );
 a7584a <=( (not A169)  and  A170 );
 a7588a <=( A199  and  (not A166) );
 a7589a <=( A167  and  a7588a );
 a7590a <=( a7589a  and  a7584a );
 a7593a <=( (not A266)  and  A200 );
 a7597a <=( A299  and  (not A298) );
 a7598a <=( (not A267)  and  a7597a );
 a7599a <=( a7598a  and  a7593a );
 a7602a <=( (not A169)  and  A170 );
 a7606a <=( A199  and  (not A166) );
 a7607a <=( A167  and  a7606a );
 a7608a <=( a7607a  and  a7602a );
 a7611a <=( (not A265)  and  A200 );
 a7615a <=( A299  and  (not A298) );
 a7616a <=( (not A266)  and  a7615a );
 a7617a <=( a7616a  and  a7611a );
 a7620a <=( (not A169)  and  A170 );
 a7624a <=( (not A199)  and  (not A166) );
 a7625a <=( A167  and  a7624a );
 a7626a <=( a7625a  and  a7620a );
 a7629a <=( (not A265)  and  A200 );
 a7633a <=( (not A300)  and  A298 );
 a7634a <=( A266  and  a7633a );
 a7635a <=( a7634a  and  a7629a );
 a7638a <=( (not A169)  and  A170 );
 a7642a <=( (not A199)  and  (not A166) );
 a7643a <=( A167  and  a7642a );
 a7644a <=( a7643a  and  a7638a );
 a7647a <=( (not A265)  and  A200 );
 a7651a <=( A299  and  A298 );
 a7652a <=( A266  and  a7651a );
 a7653a <=( a7652a  and  a7647a );
 a7656a <=( (not A169)  and  A170 );
 a7660a <=( (not A199)  and  (not A166) );
 a7661a <=( A167  and  a7660a );
 a7662a <=( a7661a  and  a7656a );
 a7665a <=( (not A265)  and  A200 );
 a7669a <=( (not A299)  and  (not A298) );
 a7670a <=( A266  and  a7669a );
 a7671a <=( a7670a  and  a7665a );
 a7674a <=( (not A169)  and  A170 );
 a7678a <=( (not A200)  and  (not A166) );
 a7679a <=( A167  and  a7678a );
 a7680a <=( a7679a  and  a7674a );
 a7683a <=( A265  and  (not A201) );
 a7687a <=( A299  and  (not A298) );
 a7688a <=( A266  and  a7687a );
 a7689a <=( a7688a  and  a7683a );
 a7692a <=( (not A169)  and  A170 );
 a7696a <=( (not A200)  and  (not A166) );
 a7697a <=( A167  and  a7696a );
 a7698a <=( a7697a  and  a7692a );
 a7701a <=( (not A266)  and  (not A201) );
 a7705a <=( A299  and  (not A298) );
 a7706a <=( (not A267)  and  a7705a );
 a7707a <=( a7706a  and  a7701a );
 a7710a <=( (not A169)  and  A170 );
 a7714a <=( (not A200)  and  (not A166) );
 a7715a <=( A167  and  a7714a );
 a7716a <=( a7715a  and  a7710a );
 a7719a <=( (not A265)  and  (not A201) );
 a7723a <=( A299  and  (not A298) );
 a7724a <=( (not A266)  and  a7723a );
 a7725a <=( a7724a  and  a7719a );
 a7728a <=( (not A169)  and  A170 );
 a7732a <=( (not A199)  and  (not A166) );
 a7733a <=( A167  and  a7732a );
 a7734a <=( a7733a  and  a7728a );
 a7737a <=( A265  and  (not A200) );
 a7741a <=( A299  and  (not A298) );
 a7742a <=( A266  and  a7741a );
 a7743a <=( a7742a  and  a7737a );
 a7746a <=( (not A169)  and  A170 );
 a7750a <=( (not A199)  and  (not A166) );
 a7751a <=( A167  and  a7750a );
 a7752a <=( a7751a  and  a7746a );
 a7755a <=( (not A266)  and  (not A200) );
 a7759a <=( A299  and  (not A298) );
 a7760a <=( (not A267)  and  a7759a );
 a7761a <=( a7760a  and  a7755a );
 a7764a <=( (not A169)  and  A170 );
 a7768a <=( (not A199)  and  (not A166) );
 a7769a <=( A167  and  a7768a );
 a7770a <=( a7769a  and  a7764a );
 a7773a <=( (not A265)  and  (not A200) );
 a7777a <=( A299  and  (not A298) );
 a7778a <=( (not A266)  and  a7777a );
 a7779a <=( a7778a  and  a7773a );
 a7782a <=( (not A169)  and  A170 );
 a7786a <=( A199  and  A166 );
 a7787a <=( (not A167)  and  a7786a );
 a7788a <=( a7787a  and  a7782a );
 a7791a <=( A265  and  A200 );
 a7795a <=( A299  and  (not A298) );
 a7796a <=( A266  and  a7795a );
 a7797a <=( a7796a  and  a7791a );
 a7800a <=( (not A169)  and  A170 );
 a7804a <=( A199  and  A166 );
 a7805a <=( (not A167)  and  a7804a );
 a7806a <=( a7805a  and  a7800a );
 a7809a <=( (not A266)  and  A200 );
 a7813a <=( A299  and  (not A298) );
 a7814a <=( (not A267)  and  a7813a );
 a7815a <=( a7814a  and  a7809a );
 a7818a <=( (not A169)  and  A170 );
 a7822a <=( A199  and  A166 );
 a7823a <=( (not A167)  and  a7822a );
 a7824a <=( a7823a  and  a7818a );
 a7827a <=( (not A265)  and  A200 );
 a7831a <=( A299  and  (not A298) );
 a7832a <=( (not A266)  and  a7831a );
 a7833a <=( a7832a  and  a7827a );
 a7836a <=( (not A169)  and  A170 );
 a7840a <=( (not A199)  and  A166 );
 a7841a <=( (not A167)  and  a7840a );
 a7842a <=( a7841a  and  a7836a );
 a7845a <=( (not A265)  and  A200 );
 a7849a <=( (not A300)  and  A298 );
 a7850a <=( A266  and  a7849a );
 a7851a <=( a7850a  and  a7845a );
 a7854a <=( (not A169)  and  A170 );
 a7858a <=( (not A199)  and  A166 );
 a7859a <=( (not A167)  and  a7858a );
 a7860a <=( a7859a  and  a7854a );
 a7863a <=( (not A265)  and  A200 );
 a7867a <=( A299  and  A298 );
 a7868a <=( A266  and  a7867a );
 a7869a <=( a7868a  and  a7863a );
 a7872a <=( (not A169)  and  A170 );
 a7876a <=( (not A199)  and  A166 );
 a7877a <=( (not A167)  and  a7876a );
 a7878a <=( a7877a  and  a7872a );
 a7881a <=( (not A265)  and  A200 );
 a7885a <=( (not A299)  and  (not A298) );
 a7886a <=( A266  and  a7885a );
 a7887a <=( a7886a  and  a7881a );
 a7890a <=( (not A169)  and  A170 );
 a7894a <=( (not A200)  and  A166 );
 a7895a <=( (not A167)  and  a7894a );
 a7896a <=( a7895a  and  a7890a );
 a7899a <=( A265  and  (not A201) );
 a7903a <=( A299  and  (not A298) );
 a7904a <=( A266  and  a7903a );
 a7905a <=( a7904a  and  a7899a );
 a7908a <=( (not A169)  and  A170 );
 a7912a <=( (not A200)  and  A166 );
 a7913a <=( (not A167)  and  a7912a );
 a7914a <=( a7913a  and  a7908a );
 a7917a <=( (not A266)  and  (not A201) );
 a7921a <=( A299  and  (not A298) );
 a7922a <=( (not A267)  and  a7921a );
 a7923a <=( a7922a  and  a7917a );
 a7926a <=( (not A169)  and  A170 );
 a7930a <=( (not A200)  and  A166 );
 a7931a <=( (not A167)  and  a7930a );
 a7932a <=( a7931a  and  a7926a );
 a7935a <=( (not A265)  and  (not A201) );
 a7939a <=( A299  and  (not A298) );
 a7940a <=( (not A266)  and  a7939a );
 a7941a <=( a7940a  and  a7935a );
 a7944a <=( (not A169)  and  A170 );
 a7948a <=( (not A199)  and  A166 );
 a7949a <=( (not A167)  and  a7948a );
 a7950a <=( a7949a  and  a7944a );
 a7953a <=( A265  and  (not A200) );
 a7957a <=( A299  and  (not A298) );
 a7958a <=( A266  and  a7957a );
 a7959a <=( a7958a  and  a7953a );
 a7962a <=( (not A169)  and  A170 );
 a7966a <=( (not A199)  and  A166 );
 a7967a <=( (not A167)  and  a7966a );
 a7968a <=( a7967a  and  a7962a );
 a7971a <=( (not A266)  and  (not A200) );
 a7975a <=( A299  and  (not A298) );
 a7976a <=( (not A267)  and  a7975a );
 a7977a <=( a7976a  and  a7971a );
 a7980a <=( (not A169)  and  A170 );
 a7984a <=( (not A199)  and  A166 );
 a7985a <=( (not A167)  and  a7984a );
 a7986a <=( a7985a  and  a7980a );
 a7989a <=( (not A265)  and  (not A200) );
 a7993a <=( A299  and  (not A298) );
 a7994a <=( (not A266)  and  a7993a );
 a7995a <=( a7994a  and  a7989a );
 a7998a <=( (not A169)  and  (not A170) );
 a8002a <=( A200  and  A199 );
 a8003a <=( (not A168)  and  a8002a );
 a8004a <=( a8003a  and  a7998a );
 a8007a <=( A266  and  (not A265) );
 a8011a <=( (not A302)  and  (not A301) );
 a8012a <=( A298  and  a8011a );
 a8013a <=( a8012a  and  a8007a );
 a8016a <=( (not A169)  and  (not A170) );
 a8020a <=( A200  and  (not A199) );
 a8021a <=( (not A168)  and  a8020a );
 a8022a <=( a8021a  and  a8016a );
 a8025a <=( (not A268)  and  (not A266) );
 a8029a <=( A299  and  (not A298) );
 a8030a <=( (not A269)  and  a8029a );
 a8031a <=( a8030a  and  a8025a );
 a8034a <=( (not A169)  and  (not A170) );
 a8038a <=( (not A202)  and  (not A200) );
 a8039a <=( (not A168)  and  a8038a );
 a8040a <=( a8039a  and  a8034a );
 a8043a <=( (not A265)  and  (not A203) );
 a8047a <=( (not A300)  and  A298 );
 a8048a <=( A266  and  a8047a );
 a8049a <=( a8048a  and  a8043a );
 a8052a <=( (not A169)  and  (not A170) );
 a8056a <=( (not A202)  and  (not A200) );
 a8057a <=( (not A168)  and  a8056a );
 a8058a <=( a8057a  and  a8052a );
 a8061a <=( (not A265)  and  (not A203) );
 a8065a <=( A299  and  A298 );
 a8066a <=( A266  and  a8065a );
 a8067a <=( a8066a  and  a8061a );
 a8070a <=( (not A169)  and  (not A170) );
 a8074a <=( (not A202)  and  (not A200) );
 a8075a <=( (not A168)  and  a8074a );
 a8076a <=( a8075a  and  a8070a );
 a8079a <=( (not A265)  and  (not A203) );
 a8083a <=( (not A299)  and  (not A298) );
 a8084a <=( A266  and  a8083a );
 a8085a <=( a8084a  and  a8079a );
 a8088a <=( (not A169)  and  (not A170) );
 a8092a <=( (not A201)  and  (not A200) );
 a8093a <=( (not A168)  and  a8092a );
 a8094a <=( a8093a  and  a8088a );
 a8097a <=( A266  and  (not A265) );
 a8101a <=( (not A302)  and  (not A301) );
 a8102a <=( A298  and  a8101a );
 a8103a <=( a8102a  and  a8097a );
 a8106a <=( (not A169)  and  (not A170) );
 a8110a <=( (not A200)  and  (not A199) );
 a8111a <=( (not A168)  and  a8110a );
 a8112a <=( a8111a  and  a8106a );
 a8115a <=( A266  and  (not A265) );
 a8119a <=( (not A302)  and  (not A301) );
 a8120a <=( A298  and  a8119a );
 a8121a <=( a8120a  and  a8115a );
 a8124a <=( A166  and  A168 );
 a8128a <=( (not A266)  and  A200 );
 a8129a <=( A199  and  a8128a );
 a8130a <=( a8129a  and  a8124a );
 a8134a <=( A298  and  (not A269) );
 a8135a <=( (not A268)  and  a8134a );
 a8139a <=( A301  and  A300 );
 a8140a <=( (not A299)  and  a8139a );
 a8141a <=( a8140a  and  a8135a );
 a8144a <=( A166  and  A168 );
 a8148a <=( (not A266)  and  A200 );
 a8149a <=( A199  and  a8148a );
 a8150a <=( a8149a  and  a8144a );
 a8154a <=( A298  and  (not A269) );
 a8155a <=( (not A268)  and  a8154a );
 a8159a <=( A302  and  A300 );
 a8160a <=( (not A299)  and  a8159a );
 a8161a <=( a8160a  and  a8155a );
 a8164a <=( A166  and  A168 );
 a8168a <=( A265  and  A200 );
 a8169a <=( (not A199)  and  a8168a );
 a8170a <=( a8169a  and  a8164a );
 a8174a <=( A268  and  A267 );
 a8175a <=( (not A266)  and  a8174a );
 a8179a <=( (not A302)  and  (not A301) );
 a8180a <=( A298  and  a8179a );
 a8181a <=( a8180a  and  a8175a );
 a8184a <=( A166  and  A168 );
 a8188a <=( A265  and  A200 );
 a8189a <=( (not A199)  and  a8188a );
 a8190a <=( a8189a  and  a8184a );
 a8194a <=( A269  and  A267 );
 a8195a <=( (not A266)  and  a8194a );
 a8199a <=( (not A302)  and  (not A301) );
 a8200a <=( A298  and  a8199a );
 a8201a <=( a8200a  and  a8195a );
 a8204a <=( A166  and  A168 );
 a8208a <=( (not A203)  and  (not A202) );
 a8209a <=( (not A200)  and  a8208a );
 a8210a <=( a8209a  and  a8204a );
 a8214a <=( A298  and  A266 );
 a8215a <=( A265  and  a8214a );
 a8219a <=( A301  and  A300 );
 a8220a <=( (not A299)  and  a8219a );
 a8221a <=( a8220a  and  a8215a );
 a8224a <=( A166  and  A168 );
 a8228a <=( (not A203)  and  (not A202) );
 a8229a <=( (not A200)  and  a8228a );
 a8230a <=( a8229a  and  a8224a );
 a8234a <=( A298  and  A266 );
 a8235a <=( A265  and  a8234a );
 a8239a <=( A302  and  A300 );
 a8240a <=( (not A299)  and  a8239a );
 a8241a <=( a8240a  and  a8235a );
 a8244a <=( A166  and  A168 );
 a8248a <=( (not A203)  and  (not A202) );
 a8249a <=( (not A200)  and  a8248a );
 a8250a <=( a8249a  and  a8244a );
 a8254a <=( A298  and  (not A267) );
 a8255a <=( (not A266)  and  a8254a );
 a8259a <=( A301  and  A300 );
 a8260a <=( (not A299)  and  a8259a );
 a8261a <=( a8260a  and  a8255a );
 a8264a <=( A166  and  A168 );
 a8268a <=( (not A203)  and  (not A202) );
 a8269a <=( (not A200)  and  a8268a );
 a8270a <=( a8269a  and  a8264a );
 a8274a <=( A298  and  (not A267) );
 a8275a <=( (not A266)  and  a8274a );
 a8279a <=( A302  and  A300 );
 a8280a <=( (not A299)  and  a8279a );
 a8281a <=( a8280a  and  a8275a );
 a8284a <=( A166  and  A168 );
 a8288a <=( (not A203)  and  (not A202) );
 a8289a <=( (not A200)  and  a8288a );
 a8290a <=( a8289a  and  a8284a );
 a8294a <=( A298  and  (not A266) );
 a8295a <=( (not A265)  and  a8294a );
 a8299a <=( A301  and  A300 );
 a8300a <=( (not A299)  and  a8299a );
 a8301a <=( a8300a  and  a8295a );
 a8304a <=( A166  and  A168 );
 a8308a <=( (not A203)  and  (not A202) );
 a8309a <=( (not A200)  and  a8308a );
 a8310a <=( a8309a  and  a8304a );
 a8314a <=( A298  and  (not A266) );
 a8315a <=( (not A265)  and  a8314a );
 a8319a <=( A302  and  A300 );
 a8320a <=( (not A299)  and  a8319a );
 a8321a <=( a8320a  and  a8315a );
 a8324a <=( A166  and  A168 );
 a8328a <=( (not A266)  and  (not A201) );
 a8329a <=( (not A200)  and  a8328a );
 a8330a <=( a8329a  and  a8324a );
 a8334a <=( A298  and  (not A269) );
 a8335a <=( (not A268)  and  a8334a );
 a8339a <=( A301  and  A300 );
 a8340a <=( (not A299)  and  a8339a );
 a8341a <=( a8340a  and  a8335a );
 a8344a <=( A166  and  A168 );
 a8348a <=( (not A266)  and  (not A201) );
 a8349a <=( (not A200)  and  a8348a );
 a8350a <=( a8349a  and  a8344a );
 a8354a <=( A298  and  (not A269) );
 a8355a <=( (not A268)  and  a8354a );
 a8359a <=( A302  and  A300 );
 a8360a <=( (not A299)  and  a8359a );
 a8361a <=( a8360a  and  a8355a );
 a8364a <=( A166  and  A168 );
 a8368a <=( A201  and  (not A200) );
 a8369a <=( A199  and  a8368a );
 a8370a <=( a8369a  and  a8364a );
 a8374a <=( A266  and  (not A265) );
 a8375a <=( A202  and  a8374a );
 a8379a <=( (not A302)  and  (not A301) );
 a8380a <=( A298  and  a8379a );
 a8381a <=( a8380a  and  a8375a );
 a8384a <=( A166  and  A168 );
 a8388a <=( A201  and  (not A200) );
 a8389a <=( A199  and  a8388a );
 a8390a <=( a8389a  and  a8384a );
 a8394a <=( A266  and  (not A265) );
 a8395a <=( A203  and  a8394a );
 a8399a <=( (not A302)  and  (not A301) );
 a8400a <=( A298  and  a8399a );
 a8401a <=( a8400a  and  a8395a );
 a8404a <=( A166  and  A168 );
 a8408a <=( (not A266)  and  (not A200) );
 a8409a <=( (not A199)  and  a8408a );
 a8410a <=( a8409a  and  a8404a );
 a8414a <=( A298  and  (not A269) );
 a8415a <=( (not A268)  and  a8414a );
 a8419a <=( A301  and  A300 );
 a8420a <=( (not A299)  and  a8419a );
 a8421a <=( a8420a  and  a8415a );
 a8424a <=( A166  and  A168 );
 a8428a <=( (not A266)  and  (not A200) );
 a8429a <=( (not A199)  and  a8428a );
 a8430a <=( a8429a  and  a8424a );
 a8434a <=( A298  and  (not A269) );
 a8435a <=( (not A268)  and  a8434a );
 a8439a <=( A302  and  A300 );
 a8440a <=( (not A299)  and  a8439a );
 a8441a <=( a8440a  and  a8435a );
 a8444a <=( A167  and  A168 );
 a8448a <=( (not A266)  and  A200 );
 a8449a <=( A199  and  a8448a );
 a8450a <=( a8449a  and  a8444a );
 a8454a <=( A298  and  (not A269) );
 a8455a <=( (not A268)  and  a8454a );
 a8459a <=( A301  and  A300 );
 a8460a <=( (not A299)  and  a8459a );
 a8461a <=( a8460a  and  a8455a );
 a8464a <=( A167  and  A168 );
 a8468a <=( (not A266)  and  A200 );
 a8469a <=( A199  and  a8468a );
 a8470a <=( a8469a  and  a8464a );
 a8474a <=( A298  and  (not A269) );
 a8475a <=( (not A268)  and  a8474a );
 a8479a <=( A302  and  A300 );
 a8480a <=( (not A299)  and  a8479a );
 a8481a <=( a8480a  and  a8475a );
 a8484a <=( A167  and  A168 );
 a8488a <=( A265  and  A200 );
 a8489a <=( (not A199)  and  a8488a );
 a8490a <=( a8489a  and  a8484a );
 a8494a <=( A268  and  A267 );
 a8495a <=( (not A266)  and  a8494a );
 a8499a <=( (not A302)  and  (not A301) );
 a8500a <=( A298  and  a8499a );
 a8501a <=( a8500a  and  a8495a );
 a8504a <=( A167  and  A168 );
 a8508a <=( A265  and  A200 );
 a8509a <=( (not A199)  and  a8508a );
 a8510a <=( a8509a  and  a8504a );
 a8514a <=( A269  and  A267 );
 a8515a <=( (not A266)  and  a8514a );
 a8519a <=( (not A302)  and  (not A301) );
 a8520a <=( A298  and  a8519a );
 a8521a <=( a8520a  and  a8515a );
 a8524a <=( A167  and  A168 );
 a8528a <=( (not A203)  and  (not A202) );
 a8529a <=( (not A200)  and  a8528a );
 a8530a <=( a8529a  and  a8524a );
 a8534a <=( A298  and  A266 );
 a8535a <=( A265  and  a8534a );
 a8539a <=( A301  and  A300 );
 a8540a <=( (not A299)  and  a8539a );
 a8541a <=( a8540a  and  a8535a );
 a8544a <=( A167  and  A168 );
 a8548a <=( (not A203)  and  (not A202) );
 a8549a <=( (not A200)  and  a8548a );
 a8550a <=( a8549a  and  a8544a );
 a8554a <=( A298  and  A266 );
 a8555a <=( A265  and  a8554a );
 a8559a <=( A302  and  A300 );
 a8560a <=( (not A299)  and  a8559a );
 a8561a <=( a8560a  and  a8555a );
 a8564a <=( A167  and  A168 );
 a8568a <=( (not A203)  and  (not A202) );
 a8569a <=( (not A200)  and  a8568a );
 a8570a <=( a8569a  and  a8564a );
 a8574a <=( A298  and  (not A267) );
 a8575a <=( (not A266)  and  a8574a );
 a8579a <=( A301  and  A300 );
 a8580a <=( (not A299)  and  a8579a );
 a8581a <=( a8580a  and  a8575a );
 a8584a <=( A167  and  A168 );
 a8588a <=( (not A203)  and  (not A202) );
 a8589a <=( (not A200)  and  a8588a );
 a8590a <=( a8589a  and  a8584a );
 a8594a <=( A298  and  (not A267) );
 a8595a <=( (not A266)  and  a8594a );
 a8599a <=( A302  and  A300 );
 a8600a <=( (not A299)  and  a8599a );
 a8601a <=( a8600a  and  a8595a );
 a8604a <=( A167  and  A168 );
 a8608a <=( (not A203)  and  (not A202) );
 a8609a <=( (not A200)  and  a8608a );
 a8610a <=( a8609a  and  a8604a );
 a8614a <=( A298  and  (not A266) );
 a8615a <=( (not A265)  and  a8614a );
 a8619a <=( A301  and  A300 );
 a8620a <=( (not A299)  and  a8619a );
 a8621a <=( a8620a  and  a8615a );
 a8624a <=( A167  and  A168 );
 a8628a <=( (not A203)  and  (not A202) );
 a8629a <=( (not A200)  and  a8628a );
 a8630a <=( a8629a  and  a8624a );
 a8634a <=( A298  and  (not A266) );
 a8635a <=( (not A265)  and  a8634a );
 a8639a <=( A302  and  A300 );
 a8640a <=( (not A299)  and  a8639a );
 a8641a <=( a8640a  and  a8635a );
 a8644a <=( A167  and  A168 );
 a8648a <=( (not A266)  and  (not A201) );
 a8649a <=( (not A200)  and  a8648a );
 a8650a <=( a8649a  and  a8644a );
 a8654a <=( A298  and  (not A269) );
 a8655a <=( (not A268)  and  a8654a );
 a8659a <=( A301  and  A300 );
 a8660a <=( (not A299)  and  a8659a );
 a8661a <=( a8660a  and  a8655a );
 a8664a <=( A167  and  A168 );
 a8668a <=( (not A266)  and  (not A201) );
 a8669a <=( (not A200)  and  a8668a );
 a8670a <=( a8669a  and  a8664a );
 a8674a <=( A298  and  (not A269) );
 a8675a <=( (not A268)  and  a8674a );
 a8679a <=( A302  and  A300 );
 a8680a <=( (not A299)  and  a8679a );
 a8681a <=( a8680a  and  a8675a );
 a8684a <=( A167  and  A168 );
 a8688a <=( A201  and  (not A200) );
 a8689a <=( A199  and  a8688a );
 a8690a <=( a8689a  and  a8684a );
 a8694a <=( A266  and  (not A265) );
 a8695a <=( A202  and  a8694a );
 a8699a <=( (not A302)  and  (not A301) );
 a8700a <=( A298  and  a8699a );
 a8701a <=( a8700a  and  a8695a );
 a8704a <=( A167  and  A168 );
 a8708a <=( A201  and  (not A200) );
 a8709a <=( A199  and  a8708a );
 a8710a <=( a8709a  and  a8704a );
 a8714a <=( A266  and  (not A265) );
 a8715a <=( A203  and  a8714a );
 a8719a <=( (not A302)  and  (not A301) );
 a8720a <=( A298  and  a8719a );
 a8721a <=( a8720a  and  a8715a );
 a8724a <=( A167  and  A168 );
 a8728a <=( (not A266)  and  (not A200) );
 a8729a <=( (not A199)  and  a8728a );
 a8730a <=( a8729a  and  a8724a );
 a8734a <=( A298  and  (not A269) );
 a8735a <=( (not A268)  and  a8734a );
 a8739a <=( A301  and  A300 );
 a8740a <=( (not A299)  and  a8739a );
 a8741a <=( a8740a  and  a8735a );
 a8744a <=( A167  and  A168 );
 a8748a <=( (not A266)  and  (not A200) );
 a8749a <=( (not A199)  and  a8748a );
 a8750a <=( a8749a  and  a8744a );
 a8754a <=( A298  and  (not A269) );
 a8755a <=( (not A268)  and  a8754a );
 a8759a <=( A302  and  A300 );
 a8760a <=( (not A299)  and  a8759a );
 a8761a <=( a8760a  and  a8755a );
 a8764a <=( (not A167)  and  A170 );
 a8768a <=( A200  and  A199 );
 a8769a <=( (not A166)  and  a8768a );
 a8770a <=( a8769a  and  a8764a );
 a8774a <=( A267  and  (not A266) );
 a8775a <=( A265  and  a8774a );
 a8779a <=( (not A300)  and  A298 );
 a8780a <=( A268  and  a8779a );
 a8781a <=( a8780a  and  a8775a );
 a8784a <=( (not A167)  and  A170 );
 a8788a <=( A200  and  A199 );
 a8789a <=( (not A166)  and  a8788a );
 a8790a <=( a8789a  and  a8784a );
 a8794a <=( A267  and  (not A266) );
 a8795a <=( A265  and  a8794a );
 a8799a <=( A299  and  A298 );
 a8800a <=( A268  and  a8799a );
 a8801a <=( a8800a  and  a8795a );
 a8804a <=( (not A167)  and  A170 );
 a8808a <=( A200  and  A199 );
 a8809a <=( (not A166)  and  a8808a );
 a8810a <=( a8809a  and  a8804a );
 a8814a <=( A267  and  (not A266) );
 a8815a <=( A265  and  a8814a );
 a8819a <=( (not A299)  and  (not A298) );
 a8820a <=( A268  and  a8819a );
 a8821a <=( a8820a  and  a8815a );
 a8824a <=( (not A167)  and  A170 );
 a8828a <=( A200  and  A199 );
 a8829a <=( (not A166)  and  a8828a );
 a8830a <=( a8829a  and  a8824a );
 a8834a <=( A267  and  (not A266) );
 a8835a <=( A265  and  a8834a );
 a8839a <=( (not A300)  and  A298 );
 a8840a <=( A269  and  a8839a );
 a8841a <=( a8840a  and  a8835a );
 a8844a <=( (not A167)  and  A170 );
 a8848a <=( A200  and  A199 );
 a8849a <=( (not A166)  and  a8848a );
 a8850a <=( a8849a  and  a8844a );
 a8854a <=( A267  and  (not A266) );
 a8855a <=( A265  and  a8854a );
 a8859a <=( A299  and  A298 );
 a8860a <=( A269  and  a8859a );
 a8861a <=( a8860a  and  a8855a );
 a8864a <=( (not A167)  and  A170 );
 a8868a <=( A200  and  A199 );
 a8869a <=( (not A166)  and  a8868a );
 a8870a <=( a8869a  and  a8864a );
 a8874a <=( A267  and  (not A266) );
 a8875a <=( A265  and  a8874a );
 a8879a <=( (not A299)  and  (not A298) );
 a8880a <=( A269  and  a8879a );
 a8881a <=( a8880a  and  a8875a );
 a8884a <=( (not A167)  and  A170 );
 a8888a <=( A200  and  (not A199) );
 a8889a <=( (not A166)  and  a8888a );
 a8890a <=( a8889a  and  a8884a );
 a8894a <=( A298  and  A266 );
 a8895a <=( A265  and  a8894a );
 a8899a <=( A301  and  A300 );
 a8900a <=( (not A299)  and  a8899a );
 a8901a <=( a8900a  and  a8895a );
 a8904a <=( (not A167)  and  A170 );
 a8908a <=( A200  and  (not A199) );
 a8909a <=( (not A166)  and  a8908a );
 a8910a <=( a8909a  and  a8904a );
 a8914a <=( A298  and  A266 );
 a8915a <=( A265  and  a8914a );
 a8919a <=( A302  and  A300 );
 a8920a <=( (not A299)  and  a8919a );
 a8921a <=( a8920a  and  a8915a );
 a8924a <=( (not A167)  and  A170 );
 a8928a <=( A200  and  (not A199) );
 a8929a <=( (not A166)  and  a8928a );
 a8930a <=( a8929a  and  a8924a );
 a8934a <=( A298  and  (not A267) );
 a8935a <=( (not A266)  and  a8934a );
 a8939a <=( A301  and  A300 );
 a8940a <=( (not A299)  and  a8939a );
 a8941a <=( a8940a  and  a8935a );
 a8944a <=( (not A167)  and  A170 );
 a8948a <=( A200  and  (not A199) );
 a8949a <=( (not A166)  and  a8948a );
 a8950a <=( a8949a  and  a8944a );
 a8954a <=( A298  and  (not A267) );
 a8955a <=( (not A266)  and  a8954a );
 a8959a <=( A302  and  A300 );
 a8960a <=( (not A299)  and  a8959a );
 a8961a <=( a8960a  and  a8955a );
 a8964a <=( (not A167)  and  A170 );
 a8968a <=( A200  and  (not A199) );
 a8969a <=( (not A166)  and  a8968a );
 a8970a <=( a8969a  and  a8964a );
 a8974a <=( A298  and  (not A266) );
 a8975a <=( (not A265)  and  a8974a );
 a8979a <=( A301  and  A300 );
 a8980a <=( (not A299)  and  a8979a );
 a8981a <=( a8980a  and  a8975a );
 a8984a <=( (not A167)  and  A170 );
 a8988a <=( A200  and  (not A199) );
 a8989a <=( (not A166)  and  a8988a );
 a8990a <=( a8989a  and  a8984a );
 a8994a <=( A298  and  (not A266) );
 a8995a <=( (not A265)  and  a8994a );
 a8999a <=( A302  and  A300 );
 a9000a <=( (not A299)  and  a8999a );
 a9001a <=( a9000a  and  a8995a );
 a9004a <=( (not A167)  and  A170 );
 a9008a <=( (not A202)  and  (not A200) );
 a9009a <=( (not A166)  and  a9008a );
 a9010a <=( a9009a  and  a9004a );
 a9014a <=( A266  and  (not A265) );
 a9015a <=( (not A203)  and  a9014a );
 a9019a <=( (not A302)  and  (not A301) );
 a9020a <=( A298  and  a9019a );
 a9021a <=( a9020a  and  a9015a );
 a9024a <=( (not A167)  and  A170 );
 a9028a <=( (not A201)  and  (not A200) );
 a9029a <=( (not A166)  and  a9028a );
 a9030a <=( a9029a  and  a9024a );
 a9034a <=( A267  and  (not A266) );
 a9035a <=( A265  and  a9034a );
 a9039a <=( (not A300)  and  A298 );
 a9040a <=( A268  and  a9039a );
 a9041a <=( a9040a  and  a9035a );
 a9044a <=( (not A167)  and  A170 );
 a9048a <=( (not A201)  and  (not A200) );
 a9049a <=( (not A166)  and  a9048a );
 a9050a <=( a9049a  and  a9044a );
 a9054a <=( A267  and  (not A266) );
 a9055a <=( A265  and  a9054a );
 a9059a <=( A299  and  A298 );
 a9060a <=( A268  and  a9059a );
 a9061a <=( a9060a  and  a9055a );
 a9064a <=( (not A167)  and  A170 );
 a9068a <=( (not A201)  and  (not A200) );
 a9069a <=( (not A166)  and  a9068a );
 a9070a <=( a9069a  and  a9064a );
 a9074a <=( A267  and  (not A266) );
 a9075a <=( A265  and  a9074a );
 a9079a <=( (not A299)  and  (not A298) );
 a9080a <=( A268  and  a9079a );
 a9081a <=( a9080a  and  a9075a );
 a9084a <=( (not A167)  and  A170 );
 a9088a <=( (not A201)  and  (not A200) );
 a9089a <=( (not A166)  and  a9088a );
 a9090a <=( a9089a  and  a9084a );
 a9094a <=( A267  and  (not A266) );
 a9095a <=( A265  and  a9094a );
 a9099a <=( (not A300)  and  A298 );
 a9100a <=( A269  and  a9099a );
 a9101a <=( a9100a  and  a9095a );
 a9104a <=( (not A167)  and  A170 );
 a9108a <=( (not A201)  and  (not A200) );
 a9109a <=( (not A166)  and  a9108a );
 a9110a <=( a9109a  and  a9104a );
 a9114a <=( A267  and  (not A266) );
 a9115a <=( A265  and  a9114a );
 a9119a <=( A299  and  A298 );
 a9120a <=( A269  and  a9119a );
 a9121a <=( a9120a  and  a9115a );
 a9124a <=( (not A167)  and  A170 );
 a9128a <=( (not A201)  and  (not A200) );
 a9129a <=( (not A166)  and  a9128a );
 a9130a <=( a9129a  and  a9124a );
 a9134a <=( A267  and  (not A266) );
 a9135a <=( A265  and  a9134a );
 a9139a <=( (not A299)  and  (not A298) );
 a9140a <=( A269  and  a9139a );
 a9141a <=( a9140a  and  a9135a );
 a9144a <=( (not A167)  and  A170 );
 a9148a <=( (not A200)  and  A199 );
 a9149a <=( (not A166)  and  a9148a );
 a9150a <=( a9149a  and  a9144a );
 a9154a <=( A265  and  A202 );
 a9155a <=( A201  and  a9154a );
 a9159a <=( A299  and  (not A298) );
 a9160a <=( A266  and  a9159a );
 a9161a <=( a9160a  and  a9155a );
 a9164a <=( (not A167)  and  A170 );
 a9168a <=( (not A200)  and  A199 );
 a9169a <=( (not A166)  and  a9168a );
 a9170a <=( a9169a  and  a9164a );
 a9174a <=( (not A266)  and  A202 );
 a9175a <=( A201  and  a9174a );
 a9179a <=( A299  and  (not A298) );
 a9180a <=( (not A267)  and  a9179a );
 a9181a <=( a9180a  and  a9175a );
 a9184a <=( (not A167)  and  A170 );
 a9188a <=( (not A200)  and  A199 );
 a9189a <=( (not A166)  and  a9188a );
 a9190a <=( a9189a  and  a9184a );
 a9194a <=( (not A265)  and  A202 );
 a9195a <=( A201  and  a9194a );
 a9199a <=( A299  and  (not A298) );
 a9200a <=( (not A266)  and  a9199a );
 a9201a <=( a9200a  and  a9195a );
 a9204a <=( (not A167)  and  A170 );
 a9208a <=( (not A200)  and  A199 );
 a9209a <=( (not A166)  and  a9208a );
 a9210a <=( a9209a  and  a9204a );
 a9214a <=( A265  and  A203 );
 a9215a <=( A201  and  a9214a );
 a9219a <=( A299  and  (not A298) );
 a9220a <=( A266  and  a9219a );
 a9221a <=( a9220a  and  a9215a );
 a9224a <=( (not A167)  and  A170 );
 a9228a <=( (not A200)  and  A199 );
 a9229a <=( (not A166)  and  a9228a );
 a9230a <=( a9229a  and  a9224a );
 a9234a <=( (not A266)  and  A203 );
 a9235a <=( A201  and  a9234a );
 a9239a <=( A299  and  (not A298) );
 a9240a <=( (not A267)  and  a9239a );
 a9241a <=( a9240a  and  a9235a );
 a9244a <=( (not A167)  and  A170 );
 a9248a <=( (not A200)  and  A199 );
 a9249a <=( (not A166)  and  a9248a );
 a9250a <=( a9249a  and  a9244a );
 a9254a <=( (not A265)  and  A203 );
 a9255a <=( A201  and  a9254a );
 a9259a <=( A299  and  (not A298) );
 a9260a <=( (not A266)  and  a9259a );
 a9261a <=( a9260a  and  a9255a );
 a9264a <=( (not A167)  and  A170 );
 a9268a <=( (not A200)  and  (not A199) );
 a9269a <=( (not A166)  and  a9268a );
 a9270a <=( a9269a  and  a9264a );
 a9274a <=( A267  and  (not A266) );
 a9275a <=( A265  and  a9274a );
 a9279a <=( (not A300)  and  A298 );
 a9280a <=( A268  and  a9279a );
 a9281a <=( a9280a  and  a9275a );
 a9284a <=( (not A167)  and  A170 );
 a9288a <=( (not A200)  and  (not A199) );
 a9289a <=( (not A166)  and  a9288a );
 a9290a <=( a9289a  and  a9284a );
 a9294a <=( A267  and  (not A266) );
 a9295a <=( A265  and  a9294a );
 a9299a <=( A299  and  A298 );
 a9300a <=( A268  and  a9299a );
 a9301a <=( a9300a  and  a9295a );
 a9304a <=( (not A167)  and  A170 );
 a9308a <=( (not A200)  and  (not A199) );
 a9309a <=( (not A166)  and  a9308a );
 a9310a <=( a9309a  and  a9304a );
 a9314a <=( A267  and  (not A266) );
 a9315a <=( A265  and  a9314a );
 a9319a <=( (not A299)  and  (not A298) );
 a9320a <=( A268  and  a9319a );
 a9321a <=( a9320a  and  a9315a );
 a9324a <=( (not A167)  and  A170 );
 a9328a <=( (not A200)  and  (not A199) );
 a9329a <=( (not A166)  and  a9328a );
 a9330a <=( a9329a  and  a9324a );
 a9334a <=( A267  and  (not A266) );
 a9335a <=( A265  and  a9334a );
 a9339a <=( (not A300)  and  A298 );
 a9340a <=( A269  and  a9339a );
 a9341a <=( a9340a  and  a9335a );
 a9344a <=( (not A167)  and  A170 );
 a9348a <=( (not A200)  and  (not A199) );
 a9349a <=( (not A166)  and  a9348a );
 a9350a <=( a9349a  and  a9344a );
 a9354a <=( A267  and  (not A266) );
 a9355a <=( A265  and  a9354a );
 a9359a <=( A299  and  A298 );
 a9360a <=( A269  and  a9359a );
 a9361a <=( a9360a  and  a9355a );
 a9364a <=( (not A167)  and  A170 );
 a9368a <=( (not A200)  and  (not A199) );
 a9369a <=( (not A166)  and  a9368a );
 a9370a <=( a9369a  and  a9364a );
 a9374a <=( A267  and  (not A266) );
 a9375a <=( A265  and  a9374a );
 a9379a <=( (not A299)  and  (not A298) );
 a9380a <=( A269  and  a9379a );
 a9381a <=( a9380a  and  a9375a );
 a9384a <=( (not A168)  and  A169 );
 a9388a <=( A199  and  (not A166) );
 a9389a <=( A167  and  a9388a );
 a9390a <=( a9389a  and  a9384a );
 a9394a <=( A266  and  (not A265) );
 a9395a <=( A200  and  a9394a );
 a9399a <=( (not A302)  and  (not A301) );
 a9400a <=( A298  and  a9399a );
 a9401a <=( a9400a  and  a9395a );
 a9404a <=( (not A168)  and  A169 );
 a9408a <=( (not A199)  and  (not A166) );
 a9409a <=( A167  and  a9408a );
 a9410a <=( a9409a  and  a9404a );
 a9414a <=( (not A268)  and  (not A266) );
 a9415a <=( A200  and  a9414a );
 a9419a <=( A299  and  (not A298) );
 a9420a <=( (not A269)  and  a9419a );
 a9421a <=( a9420a  and  a9415a );
 a9424a <=( (not A168)  and  A169 );
 a9428a <=( (not A200)  and  (not A166) );
 a9429a <=( A167  and  a9428a );
 a9430a <=( a9429a  and  a9424a );
 a9434a <=( (not A265)  and  (not A203) );
 a9435a <=( (not A202)  and  a9434a );
 a9439a <=( (not A300)  and  A298 );
 a9440a <=( A266  and  a9439a );
 a9441a <=( a9440a  and  a9435a );
 a9444a <=( (not A168)  and  A169 );
 a9448a <=( (not A200)  and  (not A166) );
 a9449a <=( A167  and  a9448a );
 a9450a <=( a9449a  and  a9444a );
 a9454a <=( (not A265)  and  (not A203) );
 a9455a <=( (not A202)  and  a9454a );
 a9459a <=( A299  and  A298 );
 a9460a <=( A266  and  a9459a );
 a9461a <=( a9460a  and  a9455a );
 a9464a <=( (not A168)  and  A169 );
 a9468a <=( (not A200)  and  (not A166) );
 a9469a <=( A167  and  a9468a );
 a9470a <=( a9469a  and  a9464a );
 a9474a <=( (not A265)  and  (not A203) );
 a9475a <=( (not A202)  and  a9474a );
 a9479a <=( (not A299)  and  (not A298) );
 a9480a <=( A266  and  a9479a );
 a9481a <=( a9480a  and  a9475a );
 a9484a <=( (not A168)  and  A169 );
 a9488a <=( (not A200)  and  (not A166) );
 a9489a <=( A167  and  a9488a );
 a9490a <=( a9489a  and  a9484a );
 a9494a <=( A266  and  (not A265) );
 a9495a <=( (not A201)  and  a9494a );
 a9499a <=( (not A302)  and  (not A301) );
 a9500a <=( A298  and  a9499a );
 a9501a <=( a9500a  and  a9495a );
 a9504a <=( (not A168)  and  A169 );
 a9508a <=( (not A199)  and  (not A166) );
 a9509a <=( A167  and  a9508a );
 a9510a <=( a9509a  and  a9504a );
 a9514a <=( A266  and  (not A265) );
 a9515a <=( (not A200)  and  a9514a );
 a9519a <=( (not A302)  and  (not A301) );
 a9520a <=( A298  and  a9519a );
 a9521a <=( a9520a  and  a9515a );
 a9524a <=( (not A168)  and  A169 );
 a9528a <=( A199  and  A166 );
 a9529a <=( (not A167)  and  a9528a );
 a9530a <=( a9529a  and  a9524a );
 a9534a <=( A266  and  (not A265) );
 a9535a <=( A200  and  a9534a );
 a9539a <=( (not A302)  and  (not A301) );
 a9540a <=( A298  and  a9539a );
 a9541a <=( a9540a  and  a9535a );
 a9544a <=( (not A168)  and  A169 );
 a9548a <=( (not A199)  and  A166 );
 a9549a <=( (not A167)  and  a9548a );
 a9550a <=( a9549a  and  a9544a );
 a9554a <=( (not A268)  and  (not A266) );
 a9555a <=( A200  and  a9554a );
 a9559a <=( A299  and  (not A298) );
 a9560a <=( (not A269)  and  a9559a );
 a9561a <=( a9560a  and  a9555a );
 a9564a <=( (not A168)  and  A169 );
 a9568a <=( (not A200)  and  A166 );
 a9569a <=( (not A167)  and  a9568a );
 a9570a <=( a9569a  and  a9564a );
 a9574a <=( (not A265)  and  (not A203) );
 a9575a <=( (not A202)  and  a9574a );
 a9579a <=( (not A300)  and  A298 );
 a9580a <=( A266  and  a9579a );
 a9581a <=( a9580a  and  a9575a );
 a9584a <=( (not A168)  and  A169 );
 a9588a <=( (not A200)  and  A166 );
 a9589a <=( (not A167)  and  a9588a );
 a9590a <=( a9589a  and  a9584a );
 a9594a <=( (not A265)  and  (not A203) );
 a9595a <=( (not A202)  and  a9594a );
 a9599a <=( A299  and  A298 );
 a9600a <=( A266  and  a9599a );
 a9601a <=( a9600a  and  a9595a );
 a9604a <=( (not A168)  and  A169 );
 a9608a <=( (not A200)  and  A166 );
 a9609a <=( (not A167)  and  a9608a );
 a9610a <=( a9609a  and  a9604a );
 a9614a <=( (not A265)  and  (not A203) );
 a9615a <=( (not A202)  and  a9614a );
 a9619a <=( (not A299)  and  (not A298) );
 a9620a <=( A266  and  a9619a );
 a9621a <=( a9620a  and  a9615a );
 a9624a <=( (not A168)  and  A169 );
 a9628a <=( (not A200)  and  A166 );
 a9629a <=( (not A167)  and  a9628a );
 a9630a <=( a9629a  and  a9624a );
 a9634a <=( A266  and  (not A265) );
 a9635a <=( (not A201)  and  a9634a );
 a9639a <=( (not A302)  and  (not A301) );
 a9640a <=( A298  and  a9639a );
 a9641a <=( a9640a  and  a9635a );
 a9644a <=( (not A168)  and  A169 );
 a9648a <=( (not A199)  and  A166 );
 a9649a <=( (not A167)  and  a9648a );
 a9650a <=( a9649a  and  a9644a );
 a9654a <=( A266  and  (not A265) );
 a9655a <=( (not A200)  and  a9654a );
 a9659a <=( (not A302)  and  (not A301) );
 a9660a <=( A298  and  a9659a );
 a9661a <=( a9660a  and  a9655a );
 a9664a <=( A169  and  A170 );
 a9668a <=( A200  and  A199 );
 a9669a <=( (not A168)  and  a9668a );
 a9670a <=( a9669a  and  a9664a );
 a9674a <=( A267  and  (not A266) );
 a9675a <=( A265  and  a9674a );
 a9679a <=( (not A300)  and  A298 );
 a9680a <=( A268  and  a9679a );
 a9681a <=( a9680a  and  a9675a );
 a9684a <=( A169  and  A170 );
 a9688a <=( A200  and  A199 );
 a9689a <=( (not A168)  and  a9688a );
 a9690a <=( a9689a  and  a9684a );
 a9694a <=( A267  and  (not A266) );
 a9695a <=( A265  and  a9694a );
 a9699a <=( A299  and  A298 );
 a9700a <=( A268  and  a9699a );
 a9701a <=( a9700a  and  a9695a );
 a9704a <=( A169  and  A170 );
 a9708a <=( A200  and  A199 );
 a9709a <=( (not A168)  and  a9708a );
 a9710a <=( a9709a  and  a9704a );
 a9714a <=( A267  and  (not A266) );
 a9715a <=( A265  and  a9714a );
 a9719a <=( (not A299)  and  (not A298) );
 a9720a <=( A268  and  a9719a );
 a9721a <=( a9720a  and  a9715a );
 a9724a <=( A169  and  A170 );
 a9728a <=( A200  and  A199 );
 a9729a <=( (not A168)  and  a9728a );
 a9730a <=( a9729a  and  a9724a );
 a9734a <=( A267  and  (not A266) );
 a9735a <=( A265  and  a9734a );
 a9739a <=( (not A300)  and  A298 );
 a9740a <=( A269  and  a9739a );
 a9741a <=( a9740a  and  a9735a );
 a9744a <=( A169  and  A170 );
 a9748a <=( A200  and  A199 );
 a9749a <=( (not A168)  and  a9748a );
 a9750a <=( a9749a  and  a9744a );
 a9754a <=( A267  and  (not A266) );
 a9755a <=( A265  and  a9754a );
 a9759a <=( A299  and  A298 );
 a9760a <=( A269  and  a9759a );
 a9761a <=( a9760a  and  a9755a );
 a9764a <=( A169  and  A170 );
 a9768a <=( A200  and  A199 );
 a9769a <=( (not A168)  and  a9768a );
 a9770a <=( a9769a  and  a9764a );
 a9774a <=( A267  and  (not A266) );
 a9775a <=( A265  and  a9774a );
 a9779a <=( (not A299)  and  (not A298) );
 a9780a <=( A269  and  a9779a );
 a9781a <=( a9780a  and  a9775a );
 a9784a <=( A169  and  A170 );
 a9788a <=( A200  and  (not A199) );
 a9789a <=( (not A168)  and  a9788a );
 a9790a <=( a9789a  and  a9784a );
 a9794a <=( A298  and  A266 );
 a9795a <=( A265  and  a9794a );
 a9799a <=( A301  and  A300 );
 a9800a <=( (not A299)  and  a9799a );
 a9801a <=( a9800a  and  a9795a );
 a9804a <=( A169  and  A170 );
 a9808a <=( A200  and  (not A199) );
 a9809a <=( (not A168)  and  a9808a );
 a9810a <=( a9809a  and  a9804a );
 a9814a <=( A298  and  A266 );
 a9815a <=( A265  and  a9814a );
 a9819a <=( A302  and  A300 );
 a9820a <=( (not A299)  and  a9819a );
 a9821a <=( a9820a  and  a9815a );
 a9824a <=( A169  and  A170 );
 a9828a <=( A200  and  (not A199) );
 a9829a <=( (not A168)  and  a9828a );
 a9830a <=( a9829a  and  a9824a );
 a9834a <=( A298  and  (not A267) );
 a9835a <=( (not A266)  and  a9834a );
 a9839a <=( A301  and  A300 );
 a9840a <=( (not A299)  and  a9839a );
 a9841a <=( a9840a  and  a9835a );
 a9844a <=( A169  and  A170 );
 a9848a <=( A200  and  (not A199) );
 a9849a <=( (not A168)  and  a9848a );
 a9850a <=( a9849a  and  a9844a );
 a9854a <=( A298  and  (not A267) );
 a9855a <=( (not A266)  and  a9854a );
 a9859a <=( A302  and  A300 );
 a9860a <=( (not A299)  and  a9859a );
 a9861a <=( a9860a  and  a9855a );
 a9864a <=( A169  and  A170 );
 a9868a <=( A200  and  (not A199) );
 a9869a <=( (not A168)  and  a9868a );
 a9870a <=( a9869a  and  a9864a );
 a9874a <=( A298  and  (not A266) );
 a9875a <=( (not A265)  and  a9874a );
 a9879a <=( A301  and  A300 );
 a9880a <=( (not A299)  and  a9879a );
 a9881a <=( a9880a  and  a9875a );
 a9884a <=( A169  and  A170 );
 a9888a <=( A200  and  (not A199) );
 a9889a <=( (not A168)  and  a9888a );
 a9890a <=( a9889a  and  a9884a );
 a9894a <=( A298  and  (not A266) );
 a9895a <=( (not A265)  and  a9894a );
 a9899a <=( A302  and  A300 );
 a9900a <=( (not A299)  and  a9899a );
 a9901a <=( a9900a  and  a9895a );
 a9904a <=( A169  and  A170 );
 a9908a <=( (not A202)  and  (not A200) );
 a9909a <=( (not A168)  and  a9908a );
 a9910a <=( a9909a  and  a9904a );
 a9914a <=( A266  and  (not A265) );
 a9915a <=( (not A203)  and  a9914a );
 a9919a <=( (not A302)  and  (not A301) );
 a9920a <=( A298  and  a9919a );
 a9921a <=( a9920a  and  a9915a );
 a9924a <=( A169  and  A170 );
 a9928a <=( (not A201)  and  (not A200) );
 a9929a <=( (not A168)  and  a9928a );
 a9930a <=( a9929a  and  a9924a );
 a9934a <=( A267  and  (not A266) );
 a9935a <=( A265  and  a9934a );
 a9939a <=( (not A300)  and  A298 );
 a9940a <=( A268  and  a9939a );
 a9941a <=( a9940a  and  a9935a );
 a9944a <=( A169  and  A170 );
 a9948a <=( (not A201)  and  (not A200) );
 a9949a <=( (not A168)  and  a9948a );
 a9950a <=( a9949a  and  a9944a );
 a9954a <=( A267  and  (not A266) );
 a9955a <=( A265  and  a9954a );
 a9959a <=( A299  and  A298 );
 a9960a <=( A268  and  a9959a );
 a9961a <=( a9960a  and  a9955a );
 a9964a <=( A169  and  A170 );
 a9968a <=( (not A201)  and  (not A200) );
 a9969a <=( (not A168)  and  a9968a );
 a9970a <=( a9969a  and  a9964a );
 a9974a <=( A267  and  (not A266) );
 a9975a <=( A265  and  a9974a );
 a9979a <=( (not A299)  and  (not A298) );
 a9980a <=( A268  and  a9979a );
 a9981a <=( a9980a  and  a9975a );
 a9984a <=( A169  and  A170 );
 a9988a <=( (not A201)  and  (not A200) );
 a9989a <=( (not A168)  and  a9988a );
 a9990a <=( a9989a  and  a9984a );
 a9994a <=( A267  and  (not A266) );
 a9995a <=( A265  and  a9994a );
 a9999a <=( (not A300)  and  A298 );
 a10000a <=( A269  and  a9999a );
 a10001a <=( a10000a  and  a9995a );
 a10004a <=( A169  and  A170 );
 a10008a <=( (not A201)  and  (not A200) );
 a10009a <=( (not A168)  and  a10008a );
 a10010a <=( a10009a  and  a10004a );
 a10014a <=( A267  and  (not A266) );
 a10015a <=( A265  and  a10014a );
 a10019a <=( A299  and  A298 );
 a10020a <=( A269  and  a10019a );
 a10021a <=( a10020a  and  a10015a );
 a10024a <=( A169  and  A170 );
 a10028a <=( (not A201)  and  (not A200) );
 a10029a <=( (not A168)  and  a10028a );
 a10030a <=( a10029a  and  a10024a );
 a10034a <=( A267  and  (not A266) );
 a10035a <=( A265  and  a10034a );
 a10039a <=( (not A299)  and  (not A298) );
 a10040a <=( A269  and  a10039a );
 a10041a <=( a10040a  and  a10035a );
 a10044a <=( A169  and  A170 );
 a10048a <=( (not A200)  and  A199 );
 a10049a <=( (not A168)  and  a10048a );
 a10050a <=( a10049a  and  a10044a );
 a10054a <=( A265  and  A202 );
 a10055a <=( A201  and  a10054a );
 a10059a <=( A299  and  (not A298) );
 a10060a <=( A266  and  a10059a );
 a10061a <=( a10060a  and  a10055a );
 a10064a <=( A169  and  A170 );
 a10068a <=( (not A200)  and  A199 );
 a10069a <=( (not A168)  and  a10068a );
 a10070a <=( a10069a  and  a10064a );
 a10074a <=( (not A266)  and  A202 );
 a10075a <=( A201  and  a10074a );
 a10079a <=( A299  and  (not A298) );
 a10080a <=( (not A267)  and  a10079a );
 a10081a <=( a10080a  and  a10075a );
 a10084a <=( A169  and  A170 );
 a10088a <=( (not A200)  and  A199 );
 a10089a <=( (not A168)  and  a10088a );
 a10090a <=( a10089a  and  a10084a );
 a10094a <=( (not A265)  and  A202 );
 a10095a <=( A201  and  a10094a );
 a10099a <=( A299  and  (not A298) );
 a10100a <=( (not A266)  and  a10099a );
 a10101a <=( a10100a  and  a10095a );
 a10104a <=( A169  and  A170 );
 a10108a <=( (not A200)  and  A199 );
 a10109a <=( (not A168)  and  a10108a );
 a10110a <=( a10109a  and  a10104a );
 a10114a <=( A265  and  A203 );
 a10115a <=( A201  and  a10114a );
 a10119a <=( A299  and  (not A298) );
 a10120a <=( A266  and  a10119a );
 a10121a <=( a10120a  and  a10115a );
 a10124a <=( A169  and  A170 );
 a10128a <=( (not A200)  and  A199 );
 a10129a <=( (not A168)  and  a10128a );
 a10130a <=( a10129a  and  a10124a );
 a10134a <=( (not A266)  and  A203 );
 a10135a <=( A201  and  a10134a );
 a10139a <=( A299  and  (not A298) );
 a10140a <=( (not A267)  and  a10139a );
 a10141a <=( a10140a  and  a10135a );
 a10144a <=( A169  and  A170 );
 a10148a <=( (not A200)  and  A199 );
 a10149a <=( (not A168)  and  a10148a );
 a10150a <=( a10149a  and  a10144a );
 a10154a <=( (not A265)  and  A203 );
 a10155a <=( A201  and  a10154a );
 a10159a <=( A299  and  (not A298) );
 a10160a <=( (not A266)  and  a10159a );
 a10161a <=( a10160a  and  a10155a );
 a10164a <=( A169  and  A170 );
 a10168a <=( (not A200)  and  (not A199) );
 a10169a <=( (not A168)  and  a10168a );
 a10170a <=( a10169a  and  a10164a );
 a10174a <=( A267  and  (not A266) );
 a10175a <=( A265  and  a10174a );
 a10179a <=( (not A300)  and  A298 );
 a10180a <=( A268  and  a10179a );
 a10181a <=( a10180a  and  a10175a );
 a10184a <=( A169  and  A170 );
 a10188a <=( (not A200)  and  (not A199) );
 a10189a <=( (not A168)  and  a10188a );
 a10190a <=( a10189a  and  a10184a );
 a10194a <=( A267  and  (not A266) );
 a10195a <=( A265  and  a10194a );
 a10199a <=( A299  and  A298 );
 a10200a <=( A268  and  a10199a );
 a10201a <=( a10200a  and  a10195a );
 a10204a <=( A169  and  A170 );
 a10208a <=( (not A200)  and  (not A199) );
 a10209a <=( (not A168)  and  a10208a );
 a10210a <=( a10209a  and  a10204a );
 a10214a <=( A267  and  (not A266) );
 a10215a <=( A265  and  a10214a );
 a10219a <=( (not A299)  and  (not A298) );
 a10220a <=( A268  and  a10219a );
 a10221a <=( a10220a  and  a10215a );
 a10224a <=( A169  and  A170 );
 a10228a <=( (not A200)  and  (not A199) );
 a10229a <=( (not A168)  and  a10228a );
 a10230a <=( a10229a  and  a10224a );
 a10234a <=( A267  and  (not A266) );
 a10235a <=( A265  and  a10234a );
 a10239a <=( (not A300)  and  A298 );
 a10240a <=( A269  and  a10239a );
 a10241a <=( a10240a  and  a10235a );
 a10244a <=( A169  and  A170 );
 a10248a <=( (not A200)  and  (not A199) );
 a10249a <=( (not A168)  and  a10248a );
 a10250a <=( a10249a  and  a10244a );
 a10254a <=( A267  and  (not A266) );
 a10255a <=( A265  and  a10254a );
 a10259a <=( A299  and  A298 );
 a10260a <=( A269  and  a10259a );
 a10261a <=( a10260a  and  a10255a );
 a10264a <=( A169  and  A170 );
 a10268a <=( (not A200)  and  (not A199) );
 a10269a <=( (not A168)  and  a10268a );
 a10270a <=( a10269a  and  a10264a );
 a10274a <=( A267  and  (not A266) );
 a10275a <=( A265  and  a10274a );
 a10279a <=( (not A299)  and  (not A298) );
 a10280a <=( A269  and  a10279a );
 a10281a <=( a10280a  and  a10275a );
 a10284a <=( A169  and  (not A170) );
 a10288a <=( A199  and  A166 );
 a10289a <=( A167  and  a10288a );
 a10290a <=( a10289a  and  a10284a );
 a10294a <=( (not A268)  and  (not A266) );
 a10295a <=( A200  and  a10294a );
 a10299a <=( A299  and  (not A298) );
 a10300a <=( (not A269)  and  a10299a );
 a10301a <=( a10300a  and  a10295a );
 a10304a <=( A169  and  (not A170) );
 a10308a <=( (not A199)  and  A166 );
 a10309a <=( A167  and  a10308a );
 a10310a <=( a10309a  and  a10304a );
 a10314a <=( A266  and  (not A265) );
 a10315a <=( A200  and  a10314a );
 a10319a <=( (not A302)  and  (not A301) );
 a10320a <=( A298  and  a10319a );
 a10321a <=( a10320a  and  a10315a );
 a10324a <=( A169  and  (not A170) );
 a10328a <=( (not A200)  and  A166 );
 a10329a <=( A167  and  a10328a );
 a10330a <=( a10329a  and  a10324a );
 a10334a <=( A265  and  (not A203) );
 a10335a <=( (not A202)  and  a10334a );
 a10339a <=( A299  and  (not A298) );
 a10340a <=( A266  and  a10339a );
 a10341a <=( a10340a  and  a10335a );
 a10344a <=( A169  and  (not A170) );
 a10348a <=( (not A200)  and  A166 );
 a10349a <=( A167  and  a10348a );
 a10350a <=( a10349a  and  a10344a );
 a10354a <=( (not A266)  and  (not A203) );
 a10355a <=( (not A202)  and  a10354a );
 a10359a <=( A299  and  (not A298) );
 a10360a <=( (not A267)  and  a10359a );
 a10361a <=( a10360a  and  a10355a );
 a10364a <=( A169  and  (not A170) );
 a10368a <=( (not A200)  and  A166 );
 a10369a <=( A167  and  a10368a );
 a10370a <=( a10369a  and  a10364a );
 a10374a <=( (not A265)  and  (not A203) );
 a10375a <=( (not A202)  and  a10374a );
 a10379a <=( A299  and  (not A298) );
 a10380a <=( (not A266)  and  a10379a );
 a10381a <=( a10380a  and  a10375a );
 a10384a <=( A169  and  (not A170) );
 a10388a <=( (not A200)  and  A166 );
 a10389a <=( A167  and  a10388a );
 a10390a <=( a10389a  and  a10384a );
 a10394a <=( (not A268)  and  (not A266) );
 a10395a <=( (not A201)  and  a10394a );
 a10399a <=( A299  and  (not A298) );
 a10400a <=( (not A269)  and  a10399a );
 a10401a <=( a10400a  and  a10395a );
 a10404a <=( A169  and  (not A170) );
 a10408a <=( (not A199)  and  A166 );
 a10409a <=( A167  and  a10408a );
 a10410a <=( a10409a  and  a10404a );
 a10414a <=( (not A268)  and  (not A266) );
 a10415a <=( (not A200)  and  a10414a );
 a10419a <=( A299  and  (not A298) );
 a10420a <=( (not A269)  and  a10419a );
 a10421a <=( a10420a  and  a10415a );
 a10424a <=( A169  and  (not A170) );
 a10428a <=( A199  and  (not A166) );
 a10429a <=( (not A167)  and  a10428a );
 a10430a <=( a10429a  and  a10424a );
 a10434a <=( (not A268)  and  (not A266) );
 a10435a <=( A200  and  a10434a );
 a10439a <=( A299  and  (not A298) );
 a10440a <=( (not A269)  and  a10439a );
 a10441a <=( a10440a  and  a10435a );
 a10444a <=( A169  and  (not A170) );
 a10448a <=( (not A199)  and  (not A166) );
 a10449a <=( (not A167)  and  a10448a );
 a10450a <=( a10449a  and  a10444a );
 a10454a <=( A266  and  (not A265) );
 a10455a <=( A200  and  a10454a );
 a10459a <=( (not A302)  and  (not A301) );
 a10460a <=( A298  and  a10459a );
 a10461a <=( a10460a  and  a10455a );
 a10464a <=( A169  and  (not A170) );
 a10468a <=( (not A200)  and  (not A166) );
 a10469a <=( (not A167)  and  a10468a );
 a10470a <=( a10469a  and  a10464a );
 a10474a <=( A265  and  (not A203) );
 a10475a <=( (not A202)  and  a10474a );
 a10479a <=( A299  and  (not A298) );
 a10480a <=( A266  and  a10479a );
 a10481a <=( a10480a  and  a10475a );
 a10484a <=( A169  and  (not A170) );
 a10488a <=( (not A200)  and  (not A166) );
 a10489a <=( (not A167)  and  a10488a );
 a10490a <=( a10489a  and  a10484a );
 a10494a <=( (not A266)  and  (not A203) );
 a10495a <=( (not A202)  and  a10494a );
 a10499a <=( A299  and  (not A298) );
 a10500a <=( (not A267)  and  a10499a );
 a10501a <=( a10500a  and  a10495a );
 a10504a <=( A169  and  (not A170) );
 a10508a <=( (not A200)  and  (not A166) );
 a10509a <=( (not A167)  and  a10508a );
 a10510a <=( a10509a  and  a10504a );
 a10514a <=( (not A265)  and  (not A203) );
 a10515a <=( (not A202)  and  a10514a );
 a10519a <=( A299  and  (not A298) );
 a10520a <=( (not A266)  and  a10519a );
 a10521a <=( a10520a  and  a10515a );
 a10524a <=( A169  and  (not A170) );
 a10528a <=( (not A200)  and  (not A166) );
 a10529a <=( (not A167)  and  a10528a );
 a10530a <=( a10529a  and  a10524a );
 a10534a <=( (not A268)  and  (not A266) );
 a10535a <=( (not A201)  and  a10534a );
 a10539a <=( A299  and  (not A298) );
 a10540a <=( (not A269)  and  a10539a );
 a10541a <=( a10540a  and  a10535a );
 a10544a <=( A169  and  (not A170) );
 a10548a <=( (not A199)  and  (not A166) );
 a10549a <=( (not A167)  and  a10548a );
 a10550a <=( a10549a  and  a10544a );
 a10554a <=( (not A268)  and  (not A266) );
 a10555a <=( (not A200)  and  a10554a );
 a10559a <=( A299  and  (not A298) );
 a10560a <=( (not A269)  and  a10559a );
 a10561a <=( a10560a  and  a10555a );
 a10564a <=( (not A167)  and  (not A169) );
 a10568a <=( A200  and  A199 );
 a10569a <=( (not A166)  and  a10568a );
 a10570a <=( a10569a  and  a10564a );
 a10574a <=( A267  and  (not A266) );
 a10575a <=( A265  and  a10574a );
 a10579a <=( (not A300)  and  A298 );
 a10580a <=( A268  and  a10579a );
 a10581a <=( a10580a  and  a10575a );
 a10584a <=( (not A167)  and  (not A169) );
 a10588a <=( A200  and  A199 );
 a10589a <=( (not A166)  and  a10588a );
 a10590a <=( a10589a  and  a10584a );
 a10594a <=( A267  and  (not A266) );
 a10595a <=( A265  and  a10594a );
 a10599a <=( A299  and  A298 );
 a10600a <=( A268  and  a10599a );
 a10601a <=( a10600a  and  a10595a );
 a10604a <=( (not A167)  and  (not A169) );
 a10608a <=( A200  and  A199 );
 a10609a <=( (not A166)  and  a10608a );
 a10610a <=( a10609a  and  a10604a );
 a10614a <=( A267  and  (not A266) );
 a10615a <=( A265  and  a10614a );
 a10619a <=( (not A299)  and  (not A298) );
 a10620a <=( A268  and  a10619a );
 a10621a <=( a10620a  and  a10615a );
 a10624a <=( (not A167)  and  (not A169) );
 a10628a <=( A200  and  A199 );
 a10629a <=( (not A166)  and  a10628a );
 a10630a <=( a10629a  and  a10624a );
 a10634a <=( A267  and  (not A266) );
 a10635a <=( A265  and  a10634a );
 a10639a <=( (not A300)  and  A298 );
 a10640a <=( A269  and  a10639a );
 a10641a <=( a10640a  and  a10635a );
 a10644a <=( (not A167)  and  (not A169) );
 a10648a <=( A200  and  A199 );
 a10649a <=( (not A166)  and  a10648a );
 a10650a <=( a10649a  and  a10644a );
 a10654a <=( A267  and  (not A266) );
 a10655a <=( A265  and  a10654a );
 a10659a <=( A299  and  A298 );
 a10660a <=( A269  and  a10659a );
 a10661a <=( a10660a  and  a10655a );
 a10664a <=( (not A167)  and  (not A169) );
 a10668a <=( A200  and  A199 );
 a10669a <=( (not A166)  and  a10668a );
 a10670a <=( a10669a  and  a10664a );
 a10674a <=( A267  and  (not A266) );
 a10675a <=( A265  and  a10674a );
 a10679a <=( (not A299)  and  (not A298) );
 a10680a <=( A269  and  a10679a );
 a10681a <=( a10680a  and  a10675a );
 a10684a <=( (not A167)  and  (not A169) );
 a10688a <=( A200  and  (not A199) );
 a10689a <=( (not A166)  and  a10688a );
 a10690a <=( a10689a  and  a10684a );
 a10694a <=( A298  and  A266 );
 a10695a <=( A265  and  a10694a );
 a10699a <=( A301  and  A300 );
 a10700a <=( (not A299)  and  a10699a );
 a10701a <=( a10700a  and  a10695a );
 a10704a <=( (not A167)  and  (not A169) );
 a10708a <=( A200  and  (not A199) );
 a10709a <=( (not A166)  and  a10708a );
 a10710a <=( a10709a  and  a10704a );
 a10714a <=( A298  and  A266 );
 a10715a <=( A265  and  a10714a );
 a10719a <=( A302  and  A300 );
 a10720a <=( (not A299)  and  a10719a );
 a10721a <=( a10720a  and  a10715a );
 a10724a <=( (not A167)  and  (not A169) );
 a10728a <=( A200  and  (not A199) );
 a10729a <=( (not A166)  and  a10728a );
 a10730a <=( a10729a  and  a10724a );
 a10734a <=( A298  and  (not A267) );
 a10735a <=( (not A266)  and  a10734a );
 a10739a <=( A301  and  A300 );
 a10740a <=( (not A299)  and  a10739a );
 a10741a <=( a10740a  and  a10735a );
 a10744a <=( (not A167)  and  (not A169) );
 a10748a <=( A200  and  (not A199) );
 a10749a <=( (not A166)  and  a10748a );
 a10750a <=( a10749a  and  a10744a );
 a10754a <=( A298  and  (not A267) );
 a10755a <=( (not A266)  and  a10754a );
 a10759a <=( A302  and  A300 );
 a10760a <=( (not A299)  and  a10759a );
 a10761a <=( a10760a  and  a10755a );
 a10764a <=( (not A167)  and  (not A169) );
 a10768a <=( A200  and  (not A199) );
 a10769a <=( (not A166)  and  a10768a );
 a10770a <=( a10769a  and  a10764a );
 a10774a <=( A298  and  (not A266) );
 a10775a <=( (not A265)  and  a10774a );
 a10779a <=( A301  and  A300 );
 a10780a <=( (not A299)  and  a10779a );
 a10781a <=( a10780a  and  a10775a );
 a10784a <=( (not A167)  and  (not A169) );
 a10788a <=( A200  and  (not A199) );
 a10789a <=( (not A166)  and  a10788a );
 a10790a <=( a10789a  and  a10784a );
 a10794a <=( A298  and  (not A266) );
 a10795a <=( (not A265)  and  a10794a );
 a10799a <=( A302  and  A300 );
 a10800a <=( (not A299)  and  a10799a );
 a10801a <=( a10800a  and  a10795a );
 a10804a <=( (not A167)  and  (not A169) );
 a10808a <=( (not A202)  and  (not A200) );
 a10809a <=( (not A166)  and  a10808a );
 a10810a <=( a10809a  and  a10804a );
 a10814a <=( A266  and  (not A265) );
 a10815a <=( (not A203)  and  a10814a );
 a10819a <=( (not A302)  and  (not A301) );
 a10820a <=( A298  and  a10819a );
 a10821a <=( a10820a  and  a10815a );
 a10824a <=( (not A167)  and  (not A169) );
 a10828a <=( (not A201)  and  (not A200) );
 a10829a <=( (not A166)  and  a10828a );
 a10830a <=( a10829a  and  a10824a );
 a10834a <=( A267  and  (not A266) );
 a10835a <=( A265  and  a10834a );
 a10839a <=( (not A300)  and  A298 );
 a10840a <=( A268  and  a10839a );
 a10841a <=( a10840a  and  a10835a );
 a10844a <=( (not A167)  and  (not A169) );
 a10848a <=( (not A201)  and  (not A200) );
 a10849a <=( (not A166)  and  a10848a );
 a10850a <=( a10849a  and  a10844a );
 a10854a <=( A267  and  (not A266) );
 a10855a <=( A265  and  a10854a );
 a10859a <=( A299  and  A298 );
 a10860a <=( A268  and  a10859a );
 a10861a <=( a10860a  and  a10855a );
 a10864a <=( (not A167)  and  (not A169) );
 a10868a <=( (not A201)  and  (not A200) );
 a10869a <=( (not A166)  and  a10868a );
 a10870a <=( a10869a  and  a10864a );
 a10874a <=( A267  and  (not A266) );
 a10875a <=( A265  and  a10874a );
 a10879a <=( (not A299)  and  (not A298) );
 a10880a <=( A268  and  a10879a );
 a10881a <=( a10880a  and  a10875a );
 a10884a <=( (not A167)  and  (not A169) );
 a10888a <=( (not A201)  and  (not A200) );
 a10889a <=( (not A166)  and  a10888a );
 a10890a <=( a10889a  and  a10884a );
 a10894a <=( A267  and  (not A266) );
 a10895a <=( A265  and  a10894a );
 a10899a <=( (not A300)  and  A298 );
 a10900a <=( A269  and  a10899a );
 a10901a <=( a10900a  and  a10895a );
 a10904a <=( (not A167)  and  (not A169) );
 a10908a <=( (not A201)  and  (not A200) );
 a10909a <=( (not A166)  and  a10908a );
 a10910a <=( a10909a  and  a10904a );
 a10914a <=( A267  and  (not A266) );
 a10915a <=( A265  and  a10914a );
 a10919a <=( A299  and  A298 );
 a10920a <=( A269  and  a10919a );
 a10921a <=( a10920a  and  a10915a );
 a10924a <=( (not A167)  and  (not A169) );
 a10928a <=( (not A201)  and  (not A200) );
 a10929a <=( (not A166)  and  a10928a );
 a10930a <=( a10929a  and  a10924a );
 a10934a <=( A267  and  (not A266) );
 a10935a <=( A265  and  a10934a );
 a10939a <=( (not A299)  and  (not A298) );
 a10940a <=( A269  and  a10939a );
 a10941a <=( a10940a  and  a10935a );
 a10944a <=( (not A167)  and  (not A169) );
 a10948a <=( (not A200)  and  A199 );
 a10949a <=( (not A166)  and  a10948a );
 a10950a <=( a10949a  and  a10944a );
 a10954a <=( A265  and  A202 );
 a10955a <=( A201  and  a10954a );
 a10959a <=( A299  and  (not A298) );
 a10960a <=( A266  and  a10959a );
 a10961a <=( a10960a  and  a10955a );
 a10964a <=( (not A167)  and  (not A169) );
 a10968a <=( (not A200)  and  A199 );
 a10969a <=( (not A166)  and  a10968a );
 a10970a <=( a10969a  and  a10964a );
 a10974a <=( (not A266)  and  A202 );
 a10975a <=( A201  and  a10974a );
 a10979a <=( A299  and  (not A298) );
 a10980a <=( (not A267)  and  a10979a );
 a10981a <=( a10980a  and  a10975a );
 a10984a <=( (not A167)  and  (not A169) );
 a10988a <=( (not A200)  and  A199 );
 a10989a <=( (not A166)  and  a10988a );
 a10990a <=( a10989a  and  a10984a );
 a10994a <=( (not A265)  and  A202 );
 a10995a <=( A201  and  a10994a );
 a10999a <=( A299  and  (not A298) );
 a11000a <=( (not A266)  and  a10999a );
 a11001a <=( a11000a  and  a10995a );
 a11004a <=( (not A167)  and  (not A169) );
 a11008a <=( (not A200)  and  A199 );
 a11009a <=( (not A166)  and  a11008a );
 a11010a <=( a11009a  and  a11004a );
 a11014a <=( A265  and  A203 );
 a11015a <=( A201  and  a11014a );
 a11019a <=( A299  and  (not A298) );
 a11020a <=( A266  and  a11019a );
 a11021a <=( a11020a  and  a11015a );
 a11024a <=( (not A167)  and  (not A169) );
 a11028a <=( (not A200)  and  A199 );
 a11029a <=( (not A166)  and  a11028a );
 a11030a <=( a11029a  and  a11024a );
 a11034a <=( (not A266)  and  A203 );
 a11035a <=( A201  and  a11034a );
 a11039a <=( A299  and  (not A298) );
 a11040a <=( (not A267)  and  a11039a );
 a11041a <=( a11040a  and  a11035a );
 a11044a <=( (not A167)  and  (not A169) );
 a11048a <=( (not A200)  and  A199 );
 a11049a <=( (not A166)  and  a11048a );
 a11050a <=( a11049a  and  a11044a );
 a11054a <=( (not A265)  and  A203 );
 a11055a <=( A201  and  a11054a );
 a11059a <=( A299  and  (not A298) );
 a11060a <=( (not A266)  and  a11059a );
 a11061a <=( a11060a  and  a11055a );
 a11064a <=( (not A167)  and  (not A169) );
 a11068a <=( (not A200)  and  (not A199) );
 a11069a <=( (not A166)  and  a11068a );
 a11070a <=( a11069a  and  a11064a );
 a11074a <=( A267  and  (not A266) );
 a11075a <=( A265  and  a11074a );
 a11079a <=( (not A300)  and  A298 );
 a11080a <=( A268  and  a11079a );
 a11081a <=( a11080a  and  a11075a );
 a11084a <=( (not A167)  and  (not A169) );
 a11088a <=( (not A200)  and  (not A199) );
 a11089a <=( (not A166)  and  a11088a );
 a11090a <=( a11089a  and  a11084a );
 a11094a <=( A267  and  (not A266) );
 a11095a <=( A265  and  a11094a );
 a11099a <=( A299  and  A298 );
 a11100a <=( A268  and  a11099a );
 a11101a <=( a11100a  and  a11095a );
 a11104a <=( (not A167)  and  (not A169) );
 a11108a <=( (not A200)  and  (not A199) );
 a11109a <=( (not A166)  and  a11108a );
 a11110a <=( a11109a  and  a11104a );
 a11114a <=( A267  and  (not A266) );
 a11115a <=( A265  and  a11114a );
 a11119a <=( (not A299)  and  (not A298) );
 a11120a <=( A268  and  a11119a );
 a11121a <=( a11120a  and  a11115a );
 a11124a <=( (not A167)  and  (not A169) );
 a11128a <=( (not A200)  and  (not A199) );
 a11129a <=( (not A166)  and  a11128a );
 a11130a <=( a11129a  and  a11124a );
 a11134a <=( A267  and  (not A266) );
 a11135a <=( A265  and  a11134a );
 a11139a <=( (not A300)  and  A298 );
 a11140a <=( A269  and  a11139a );
 a11141a <=( a11140a  and  a11135a );
 a11144a <=( (not A167)  and  (not A169) );
 a11148a <=( (not A200)  and  (not A199) );
 a11149a <=( (not A166)  and  a11148a );
 a11150a <=( a11149a  and  a11144a );
 a11154a <=( A267  and  (not A266) );
 a11155a <=( A265  and  a11154a );
 a11159a <=( A299  and  A298 );
 a11160a <=( A269  and  a11159a );
 a11161a <=( a11160a  and  a11155a );
 a11164a <=( (not A167)  and  (not A169) );
 a11168a <=( (not A200)  and  (not A199) );
 a11169a <=( (not A166)  and  a11168a );
 a11170a <=( a11169a  and  a11164a );
 a11174a <=( A267  and  (not A266) );
 a11175a <=( A265  and  a11174a );
 a11179a <=( (not A299)  and  (not A298) );
 a11180a <=( A269  and  a11179a );
 a11181a <=( a11180a  and  a11175a );
 a11184a <=( (not A168)  and  (not A169) );
 a11188a <=( A199  and  A166 );
 a11189a <=( A167  and  a11188a );
 a11190a <=( a11189a  and  a11184a );
 a11194a <=( A266  and  (not A265) );
 a11195a <=( A200  and  a11194a );
 a11199a <=( (not A302)  and  (not A301) );
 a11200a <=( A298  and  a11199a );
 a11201a <=( a11200a  and  a11195a );
 a11204a <=( (not A168)  and  (not A169) );
 a11208a <=( (not A199)  and  A166 );
 a11209a <=( A167  and  a11208a );
 a11210a <=( a11209a  and  a11204a );
 a11214a <=( (not A268)  and  (not A266) );
 a11215a <=( A200  and  a11214a );
 a11219a <=( A299  and  (not A298) );
 a11220a <=( (not A269)  and  a11219a );
 a11221a <=( a11220a  and  a11215a );
 a11224a <=( (not A168)  and  (not A169) );
 a11228a <=( (not A200)  and  A166 );
 a11229a <=( A167  and  a11228a );
 a11230a <=( a11229a  and  a11224a );
 a11234a <=( (not A265)  and  (not A203) );
 a11235a <=( (not A202)  and  a11234a );
 a11239a <=( (not A300)  and  A298 );
 a11240a <=( A266  and  a11239a );
 a11241a <=( a11240a  and  a11235a );
 a11244a <=( (not A168)  and  (not A169) );
 a11248a <=( (not A200)  and  A166 );
 a11249a <=( A167  and  a11248a );
 a11250a <=( a11249a  and  a11244a );
 a11254a <=( (not A265)  and  (not A203) );
 a11255a <=( (not A202)  and  a11254a );
 a11259a <=( A299  and  A298 );
 a11260a <=( A266  and  a11259a );
 a11261a <=( a11260a  and  a11255a );
 a11264a <=( (not A168)  and  (not A169) );
 a11268a <=( (not A200)  and  A166 );
 a11269a <=( A167  and  a11268a );
 a11270a <=( a11269a  and  a11264a );
 a11274a <=( (not A265)  and  (not A203) );
 a11275a <=( (not A202)  and  a11274a );
 a11279a <=( (not A299)  and  (not A298) );
 a11280a <=( A266  and  a11279a );
 a11281a <=( a11280a  and  a11275a );
 a11284a <=( (not A168)  and  (not A169) );
 a11288a <=( (not A200)  and  A166 );
 a11289a <=( A167  and  a11288a );
 a11290a <=( a11289a  and  a11284a );
 a11294a <=( A266  and  (not A265) );
 a11295a <=( (not A201)  and  a11294a );
 a11299a <=( (not A302)  and  (not A301) );
 a11300a <=( A298  and  a11299a );
 a11301a <=( a11300a  and  a11295a );
 a11304a <=( (not A168)  and  (not A169) );
 a11308a <=( (not A199)  and  A166 );
 a11309a <=( A167  and  a11308a );
 a11310a <=( a11309a  and  a11304a );
 a11314a <=( A266  and  (not A265) );
 a11315a <=( (not A200)  and  a11314a );
 a11319a <=( (not A302)  and  (not A301) );
 a11320a <=( A298  and  a11319a );
 a11321a <=( a11320a  and  a11315a );
 a11324a <=( (not A169)  and  A170 );
 a11328a <=( A199  and  (not A166) );
 a11329a <=( A167  and  a11328a );
 a11330a <=( a11329a  and  a11324a );
 a11334a <=( (not A268)  and  (not A266) );
 a11335a <=( A200  and  a11334a );
 a11339a <=( A299  and  (not A298) );
 a11340a <=( (not A269)  and  a11339a );
 a11341a <=( a11340a  and  a11335a );
 a11344a <=( (not A169)  and  A170 );
 a11348a <=( (not A199)  and  (not A166) );
 a11349a <=( A167  and  a11348a );
 a11350a <=( a11349a  and  a11344a );
 a11354a <=( A266  and  (not A265) );
 a11355a <=( A200  and  a11354a );
 a11359a <=( (not A302)  and  (not A301) );
 a11360a <=( A298  and  a11359a );
 a11361a <=( a11360a  and  a11355a );
 a11364a <=( (not A169)  and  A170 );
 a11368a <=( (not A200)  and  (not A166) );
 a11369a <=( A167  and  a11368a );
 a11370a <=( a11369a  and  a11364a );
 a11374a <=( A265  and  (not A203) );
 a11375a <=( (not A202)  and  a11374a );
 a11379a <=( A299  and  (not A298) );
 a11380a <=( A266  and  a11379a );
 a11381a <=( a11380a  and  a11375a );
 a11384a <=( (not A169)  and  A170 );
 a11388a <=( (not A200)  and  (not A166) );
 a11389a <=( A167  and  a11388a );
 a11390a <=( a11389a  and  a11384a );
 a11394a <=( (not A266)  and  (not A203) );
 a11395a <=( (not A202)  and  a11394a );
 a11399a <=( A299  and  (not A298) );
 a11400a <=( (not A267)  and  a11399a );
 a11401a <=( a11400a  and  a11395a );
 a11404a <=( (not A169)  and  A170 );
 a11408a <=( (not A200)  and  (not A166) );
 a11409a <=( A167  and  a11408a );
 a11410a <=( a11409a  and  a11404a );
 a11414a <=( (not A265)  and  (not A203) );
 a11415a <=( (not A202)  and  a11414a );
 a11419a <=( A299  and  (not A298) );
 a11420a <=( (not A266)  and  a11419a );
 a11421a <=( a11420a  and  a11415a );
 a11424a <=( (not A169)  and  A170 );
 a11428a <=( (not A200)  and  (not A166) );
 a11429a <=( A167  and  a11428a );
 a11430a <=( a11429a  and  a11424a );
 a11434a <=( (not A268)  and  (not A266) );
 a11435a <=( (not A201)  and  a11434a );
 a11439a <=( A299  and  (not A298) );
 a11440a <=( (not A269)  and  a11439a );
 a11441a <=( a11440a  and  a11435a );
 a11444a <=( (not A169)  and  A170 );
 a11448a <=( (not A199)  and  (not A166) );
 a11449a <=( A167  and  a11448a );
 a11450a <=( a11449a  and  a11444a );
 a11454a <=( (not A268)  and  (not A266) );
 a11455a <=( (not A200)  and  a11454a );
 a11459a <=( A299  and  (not A298) );
 a11460a <=( (not A269)  and  a11459a );
 a11461a <=( a11460a  and  a11455a );
 a11464a <=( (not A169)  and  A170 );
 a11468a <=( A199  and  A166 );
 a11469a <=( (not A167)  and  a11468a );
 a11470a <=( a11469a  and  a11464a );
 a11474a <=( (not A268)  and  (not A266) );
 a11475a <=( A200  and  a11474a );
 a11479a <=( A299  and  (not A298) );
 a11480a <=( (not A269)  and  a11479a );
 a11481a <=( a11480a  and  a11475a );
 a11484a <=( (not A169)  and  A170 );
 a11488a <=( (not A199)  and  A166 );
 a11489a <=( (not A167)  and  a11488a );
 a11490a <=( a11489a  and  a11484a );
 a11494a <=( A266  and  (not A265) );
 a11495a <=( A200  and  a11494a );
 a11499a <=( (not A302)  and  (not A301) );
 a11500a <=( A298  and  a11499a );
 a11501a <=( a11500a  and  a11495a );
 a11504a <=( (not A169)  and  A170 );
 a11508a <=( (not A200)  and  A166 );
 a11509a <=( (not A167)  and  a11508a );
 a11510a <=( a11509a  and  a11504a );
 a11514a <=( A265  and  (not A203) );
 a11515a <=( (not A202)  and  a11514a );
 a11519a <=( A299  and  (not A298) );
 a11520a <=( A266  and  a11519a );
 a11521a <=( a11520a  and  a11515a );
 a11524a <=( (not A169)  and  A170 );
 a11528a <=( (not A200)  and  A166 );
 a11529a <=( (not A167)  and  a11528a );
 a11530a <=( a11529a  and  a11524a );
 a11534a <=( (not A266)  and  (not A203) );
 a11535a <=( (not A202)  and  a11534a );
 a11539a <=( A299  and  (not A298) );
 a11540a <=( (not A267)  and  a11539a );
 a11541a <=( a11540a  and  a11535a );
 a11544a <=( (not A169)  and  A170 );
 a11548a <=( (not A200)  and  A166 );
 a11549a <=( (not A167)  and  a11548a );
 a11550a <=( a11549a  and  a11544a );
 a11554a <=( (not A265)  and  (not A203) );
 a11555a <=( (not A202)  and  a11554a );
 a11559a <=( A299  and  (not A298) );
 a11560a <=( (not A266)  and  a11559a );
 a11561a <=( a11560a  and  a11555a );
 a11564a <=( (not A169)  and  A170 );
 a11568a <=( (not A200)  and  A166 );
 a11569a <=( (not A167)  and  a11568a );
 a11570a <=( a11569a  and  a11564a );
 a11574a <=( (not A268)  and  (not A266) );
 a11575a <=( (not A201)  and  a11574a );
 a11579a <=( A299  and  (not A298) );
 a11580a <=( (not A269)  and  a11579a );
 a11581a <=( a11580a  and  a11575a );
 a11584a <=( (not A169)  and  A170 );
 a11588a <=( (not A199)  and  A166 );
 a11589a <=( (not A167)  and  a11588a );
 a11590a <=( a11589a  and  a11584a );
 a11594a <=( (not A268)  and  (not A266) );
 a11595a <=( (not A200)  and  a11594a );
 a11599a <=( A299  and  (not A298) );
 a11600a <=( (not A269)  and  a11599a );
 a11601a <=( a11600a  and  a11595a );
 a11604a <=( (not A169)  and  (not A170) );
 a11608a <=( A200  and  A199 );
 a11609a <=( (not A168)  and  a11608a );
 a11610a <=( a11609a  and  a11604a );
 a11614a <=( A267  and  (not A266) );
 a11615a <=( A265  and  a11614a );
 a11619a <=( (not A300)  and  A298 );
 a11620a <=( A268  and  a11619a );
 a11621a <=( a11620a  and  a11615a );
 a11624a <=( (not A169)  and  (not A170) );
 a11628a <=( A200  and  A199 );
 a11629a <=( (not A168)  and  a11628a );
 a11630a <=( a11629a  and  a11624a );
 a11634a <=( A267  and  (not A266) );
 a11635a <=( A265  and  a11634a );
 a11639a <=( A299  and  A298 );
 a11640a <=( A268  and  a11639a );
 a11641a <=( a11640a  and  a11635a );
 a11644a <=( (not A169)  and  (not A170) );
 a11648a <=( A200  and  A199 );
 a11649a <=( (not A168)  and  a11648a );
 a11650a <=( a11649a  and  a11644a );
 a11654a <=( A267  and  (not A266) );
 a11655a <=( A265  and  a11654a );
 a11659a <=( (not A299)  and  (not A298) );
 a11660a <=( A268  and  a11659a );
 a11661a <=( a11660a  and  a11655a );
 a11664a <=( (not A169)  and  (not A170) );
 a11668a <=( A200  and  A199 );
 a11669a <=( (not A168)  and  a11668a );
 a11670a <=( a11669a  and  a11664a );
 a11674a <=( A267  and  (not A266) );
 a11675a <=( A265  and  a11674a );
 a11679a <=( (not A300)  and  A298 );
 a11680a <=( A269  and  a11679a );
 a11681a <=( a11680a  and  a11675a );
 a11684a <=( (not A169)  and  (not A170) );
 a11688a <=( A200  and  A199 );
 a11689a <=( (not A168)  and  a11688a );
 a11690a <=( a11689a  and  a11684a );
 a11694a <=( A267  and  (not A266) );
 a11695a <=( A265  and  a11694a );
 a11699a <=( A299  and  A298 );
 a11700a <=( A269  and  a11699a );
 a11701a <=( a11700a  and  a11695a );
 a11704a <=( (not A169)  and  (not A170) );
 a11708a <=( A200  and  A199 );
 a11709a <=( (not A168)  and  a11708a );
 a11710a <=( a11709a  and  a11704a );
 a11714a <=( A267  and  (not A266) );
 a11715a <=( A265  and  a11714a );
 a11719a <=( (not A299)  and  (not A298) );
 a11720a <=( A269  and  a11719a );
 a11721a <=( a11720a  and  a11715a );
 a11724a <=( (not A169)  and  (not A170) );
 a11728a <=( A200  and  (not A199) );
 a11729a <=( (not A168)  and  a11728a );
 a11730a <=( a11729a  and  a11724a );
 a11734a <=( A298  and  A266 );
 a11735a <=( A265  and  a11734a );
 a11739a <=( A301  and  A300 );
 a11740a <=( (not A299)  and  a11739a );
 a11741a <=( a11740a  and  a11735a );
 a11744a <=( (not A169)  and  (not A170) );
 a11748a <=( A200  and  (not A199) );
 a11749a <=( (not A168)  and  a11748a );
 a11750a <=( a11749a  and  a11744a );
 a11754a <=( A298  and  A266 );
 a11755a <=( A265  and  a11754a );
 a11759a <=( A302  and  A300 );
 a11760a <=( (not A299)  and  a11759a );
 a11761a <=( a11760a  and  a11755a );
 a11764a <=( (not A169)  and  (not A170) );
 a11768a <=( A200  and  (not A199) );
 a11769a <=( (not A168)  and  a11768a );
 a11770a <=( a11769a  and  a11764a );
 a11774a <=( A298  and  (not A267) );
 a11775a <=( (not A266)  and  a11774a );
 a11779a <=( A301  and  A300 );
 a11780a <=( (not A299)  and  a11779a );
 a11781a <=( a11780a  and  a11775a );
 a11784a <=( (not A169)  and  (not A170) );
 a11788a <=( A200  and  (not A199) );
 a11789a <=( (not A168)  and  a11788a );
 a11790a <=( a11789a  and  a11784a );
 a11794a <=( A298  and  (not A267) );
 a11795a <=( (not A266)  and  a11794a );
 a11799a <=( A302  and  A300 );
 a11800a <=( (not A299)  and  a11799a );
 a11801a <=( a11800a  and  a11795a );
 a11804a <=( (not A169)  and  (not A170) );
 a11808a <=( A200  and  (not A199) );
 a11809a <=( (not A168)  and  a11808a );
 a11810a <=( a11809a  and  a11804a );
 a11814a <=( A298  and  (not A266) );
 a11815a <=( (not A265)  and  a11814a );
 a11819a <=( A301  and  A300 );
 a11820a <=( (not A299)  and  a11819a );
 a11821a <=( a11820a  and  a11815a );
 a11824a <=( (not A169)  and  (not A170) );
 a11828a <=( A200  and  (not A199) );
 a11829a <=( (not A168)  and  a11828a );
 a11830a <=( a11829a  and  a11824a );
 a11834a <=( A298  and  (not A266) );
 a11835a <=( (not A265)  and  a11834a );
 a11839a <=( A302  and  A300 );
 a11840a <=( (not A299)  and  a11839a );
 a11841a <=( a11840a  and  a11835a );
 a11844a <=( (not A169)  and  (not A170) );
 a11848a <=( (not A202)  and  (not A200) );
 a11849a <=( (not A168)  and  a11848a );
 a11850a <=( a11849a  and  a11844a );
 a11854a <=( A266  and  (not A265) );
 a11855a <=( (not A203)  and  a11854a );
 a11859a <=( (not A302)  and  (not A301) );
 a11860a <=( A298  and  a11859a );
 a11861a <=( a11860a  and  a11855a );
 a11864a <=( (not A169)  and  (not A170) );
 a11868a <=( (not A201)  and  (not A200) );
 a11869a <=( (not A168)  and  a11868a );
 a11870a <=( a11869a  and  a11864a );
 a11874a <=( A267  and  (not A266) );
 a11875a <=( A265  and  a11874a );
 a11879a <=( (not A300)  and  A298 );
 a11880a <=( A268  and  a11879a );
 a11881a <=( a11880a  and  a11875a );
 a11884a <=( (not A169)  and  (not A170) );
 a11888a <=( (not A201)  and  (not A200) );
 a11889a <=( (not A168)  and  a11888a );
 a11890a <=( a11889a  and  a11884a );
 a11894a <=( A267  and  (not A266) );
 a11895a <=( A265  and  a11894a );
 a11899a <=( A299  and  A298 );
 a11900a <=( A268  and  a11899a );
 a11901a <=( a11900a  and  a11895a );
 a11904a <=( (not A169)  and  (not A170) );
 a11908a <=( (not A201)  and  (not A200) );
 a11909a <=( (not A168)  and  a11908a );
 a11910a <=( a11909a  and  a11904a );
 a11914a <=( A267  and  (not A266) );
 a11915a <=( A265  and  a11914a );
 a11919a <=( (not A299)  and  (not A298) );
 a11920a <=( A268  and  a11919a );
 a11921a <=( a11920a  and  a11915a );
 a11924a <=( (not A169)  and  (not A170) );
 a11928a <=( (not A201)  and  (not A200) );
 a11929a <=( (not A168)  and  a11928a );
 a11930a <=( a11929a  and  a11924a );
 a11934a <=( A267  and  (not A266) );
 a11935a <=( A265  and  a11934a );
 a11939a <=( (not A300)  and  A298 );
 a11940a <=( A269  and  a11939a );
 a11941a <=( a11940a  and  a11935a );
 a11944a <=( (not A169)  and  (not A170) );
 a11948a <=( (not A201)  and  (not A200) );
 a11949a <=( (not A168)  and  a11948a );
 a11950a <=( a11949a  and  a11944a );
 a11954a <=( A267  and  (not A266) );
 a11955a <=( A265  and  a11954a );
 a11959a <=( A299  and  A298 );
 a11960a <=( A269  and  a11959a );
 a11961a <=( a11960a  and  a11955a );
 a11964a <=( (not A169)  and  (not A170) );
 a11968a <=( (not A201)  and  (not A200) );
 a11969a <=( (not A168)  and  a11968a );
 a11970a <=( a11969a  and  a11964a );
 a11974a <=( A267  and  (not A266) );
 a11975a <=( A265  and  a11974a );
 a11979a <=( (not A299)  and  (not A298) );
 a11980a <=( A269  and  a11979a );
 a11981a <=( a11980a  and  a11975a );
 a11984a <=( (not A169)  and  (not A170) );
 a11988a <=( (not A200)  and  A199 );
 a11989a <=( (not A168)  and  a11988a );
 a11990a <=( a11989a  and  a11984a );
 a11994a <=( A265  and  A202 );
 a11995a <=( A201  and  a11994a );
 a11999a <=( A299  and  (not A298) );
 a12000a <=( A266  and  a11999a );
 a12001a <=( a12000a  and  a11995a );
 a12004a <=( (not A169)  and  (not A170) );
 a12008a <=( (not A200)  and  A199 );
 a12009a <=( (not A168)  and  a12008a );
 a12010a <=( a12009a  and  a12004a );
 a12014a <=( (not A266)  and  A202 );
 a12015a <=( A201  and  a12014a );
 a12019a <=( A299  and  (not A298) );
 a12020a <=( (not A267)  and  a12019a );
 a12021a <=( a12020a  and  a12015a );
 a12024a <=( (not A169)  and  (not A170) );
 a12028a <=( (not A200)  and  A199 );
 a12029a <=( (not A168)  and  a12028a );
 a12030a <=( a12029a  and  a12024a );
 a12034a <=( (not A265)  and  A202 );
 a12035a <=( A201  and  a12034a );
 a12039a <=( A299  and  (not A298) );
 a12040a <=( (not A266)  and  a12039a );
 a12041a <=( a12040a  and  a12035a );
 a12044a <=( (not A169)  and  (not A170) );
 a12048a <=( (not A200)  and  A199 );
 a12049a <=( (not A168)  and  a12048a );
 a12050a <=( a12049a  and  a12044a );
 a12054a <=( A265  and  A203 );
 a12055a <=( A201  and  a12054a );
 a12059a <=( A299  and  (not A298) );
 a12060a <=( A266  and  a12059a );
 a12061a <=( a12060a  and  a12055a );
 a12064a <=( (not A169)  and  (not A170) );
 a12068a <=( (not A200)  and  A199 );
 a12069a <=( (not A168)  and  a12068a );
 a12070a <=( a12069a  and  a12064a );
 a12074a <=( (not A266)  and  A203 );
 a12075a <=( A201  and  a12074a );
 a12079a <=( A299  and  (not A298) );
 a12080a <=( (not A267)  and  a12079a );
 a12081a <=( a12080a  and  a12075a );
 a12084a <=( (not A169)  and  (not A170) );
 a12088a <=( (not A200)  and  A199 );
 a12089a <=( (not A168)  and  a12088a );
 a12090a <=( a12089a  and  a12084a );
 a12094a <=( (not A265)  and  A203 );
 a12095a <=( A201  and  a12094a );
 a12099a <=( A299  and  (not A298) );
 a12100a <=( (not A266)  and  a12099a );
 a12101a <=( a12100a  and  a12095a );
 a12104a <=( (not A169)  and  (not A170) );
 a12108a <=( (not A200)  and  (not A199) );
 a12109a <=( (not A168)  and  a12108a );
 a12110a <=( a12109a  and  a12104a );
 a12114a <=( A267  and  (not A266) );
 a12115a <=( A265  and  a12114a );
 a12119a <=( (not A300)  and  A298 );
 a12120a <=( A268  and  a12119a );
 a12121a <=( a12120a  and  a12115a );
 a12124a <=( (not A169)  and  (not A170) );
 a12128a <=( (not A200)  and  (not A199) );
 a12129a <=( (not A168)  and  a12128a );
 a12130a <=( a12129a  and  a12124a );
 a12134a <=( A267  and  (not A266) );
 a12135a <=( A265  and  a12134a );
 a12139a <=( A299  and  A298 );
 a12140a <=( A268  and  a12139a );
 a12141a <=( a12140a  and  a12135a );
 a12144a <=( (not A169)  and  (not A170) );
 a12148a <=( (not A200)  and  (not A199) );
 a12149a <=( (not A168)  and  a12148a );
 a12150a <=( a12149a  and  a12144a );
 a12154a <=( A267  and  (not A266) );
 a12155a <=( A265  and  a12154a );
 a12159a <=( (not A299)  and  (not A298) );
 a12160a <=( A268  and  a12159a );
 a12161a <=( a12160a  and  a12155a );
 a12164a <=( (not A169)  and  (not A170) );
 a12168a <=( (not A200)  and  (not A199) );
 a12169a <=( (not A168)  and  a12168a );
 a12170a <=( a12169a  and  a12164a );
 a12174a <=( A267  and  (not A266) );
 a12175a <=( A265  and  a12174a );
 a12179a <=( (not A300)  and  A298 );
 a12180a <=( A269  and  a12179a );
 a12181a <=( a12180a  and  a12175a );
 a12184a <=( (not A169)  and  (not A170) );
 a12188a <=( (not A200)  and  (not A199) );
 a12189a <=( (not A168)  and  a12188a );
 a12190a <=( a12189a  and  a12184a );
 a12194a <=( A267  and  (not A266) );
 a12195a <=( A265  and  a12194a );
 a12199a <=( A299  and  A298 );
 a12200a <=( A269  and  a12199a );
 a12201a <=( a12200a  and  a12195a );
 a12204a <=( (not A169)  and  (not A170) );
 a12208a <=( (not A200)  and  (not A199) );
 a12209a <=( (not A168)  and  a12208a );
 a12210a <=( a12209a  and  a12204a );
 a12214a <=( A267  and  (not A266) );
 a12215a <=( A265  and  a12214a );
 a12219a <=( (not A299)  and  (not A298) );
 a12220a <=( A269  and  a12219a );
 a12221a <=( a12220a  and  a12215a );
 a12225a <=( (not A200)  and  A166 );
 a12226a <=( A168  and  a12225a );
 a12230a <=( (not A266)  and  (not A203) );
 a12231a <=( (not A202)  and  a12230a );
 a12232a <=( a12231a  and  a12226a );
 a12236a <=( A298  and  (not A269) );
 a12237a <=( (not A268)  and  a12236a );
 a12241a <=( A301  and  A300 );
 a12242a <=( (not A299)  and  a12241a );
 a12243a <=( a12242a  and  a12237a );
 a12247a <=( (not A200)  and  A166 );
 a12248a <=( A168  and  a12247a );
 a12252a <=( (not A266)  and  (not A203) );
 a12253a <=( (not A202)  and  a12252a );
 a12254a <=( a12253a  and  a12248a );
 a12258a <=( A298  and  (not A269) );
 a12259a <=( (not A268)  and  a12258a );
 a12263a <=( A302  and  A300 );
 a12264a <=( (not A299)  and  a12263a );
 a12265a <=( a12264a  and  a12259a );
 a12269a <=( A199  and  A166 );
 a12270a <=( A168  and  a12269a );
 a12274a <=( A202  and  A201 );
 a12275a <=( (not A200)  and  a12274a );
 a12276a <=( a12275a  and  a12270a );
 a12280a <=( A267  and  (not A266) );
 a12281a <=( A265  and  a12280a );
 a12285a <=( (not A300)  and  A298 );
 a12286a <=( A268  and  a12285a );
 a12287a <=( a12286a  and  a12281a );
 a12291a <=( A199  and  A166 );
 a12292a <=( A168  and  a12291a );
 a12296a <=( A202  and  A201 );
 a12297a <=( (not A200)  and  a12296a );
 a12298a <=( a12297a  and  a12292a );
 a12302a <=( A267  and  (not A266) );
 a12303a <=( A265  and  a12302a );
 a12307a <=( A299  and  A298 );
 a12308a <=( A268  and  a12307a );
 a12309a <=( a12308a  and  a12303a );
 a12313a <=( A199  and  A166 );
 a12314a <=( A168  and  a12313a );
 a12318a <=( A202  and  A201 );
 a12319a <=( (not A200)  and  a12318a );
 a12320a <=( a12319a  and  a12314a );
 a12324a <=( A267  and  (not A266) );
 a12325a <=( A265  and  a12324a );
 a12329a <=( (not A299)  and  (not A298) );
 a12330a <=( A268  and  a12329a );
 a12331a <=( a12330a  and  a12325a );
 a12335a <=( A199  and  A166 );
 a12336a <=( A168  and  a12335a );
 a12340a <=( A202  and  A201 );
 a12341a <=( (not A200)  and  a12340a );
 a12342a <=( a12341a  and  a12336a );
 a12346a <=( A267  and  (not A266) );
 a12347a <=( A265  and  a12346a );
 a12351a <=( (not A300)  and  A298 );
 a12352a <=( A269  and  a12351a );
 a12353a <=( a12352a  and  a12347a );
 a12357a <=( A199  and  A166 );
 a12358a <=( A168  and  a12357a );
 a12362a <=( A202  and  A201 );
 a12363a <=( (not A200)  and  a12362a );
 a12364a <=( a12363a  and  a12358a );
 a12368a <=( A267  and  (not A266) );
 a12369a <=( A265  and  a12368a );
 a12373a <=( A299  and  A298 );
 a12374a <=( A269  and  a12373a );
 a12375a <=( a12374a  and  a12369a );
 a12379a <=( A199  and  A166 );
 a12380a <=( A168  and  a12379a );
 a12384a <=( A202  and  A201 );
 a12385a <=( (not A200)  and  a12384a );
 a12386a <=( a12385a  and  a12380a );
 a12390a <=( A267  and  (not A266) );
 a12391a <=( A265  and  a12390a );
 a12395a <=( (not A299)  and  (not A298) );
 a12396a <=( A269  and  a12395a );
 a12397a <=( a12396a  and  a12391a );
 a12401a <=( A199  and  A166 );
 a12402a <=( A168  and  a12401a );
 a12406a <=( A203  and  A201 );
 a12407a <=( (not A200)  and  a12406a );
 a12408a <=( a12407a  and  a12402a );
 a12412a <=( A267  and  (not A266) );
 a12413a <=( A265  and  a12412a );
 a12417a <=( (not A300)  and  A298 );
 a12418a <=( A268  and  a12417a );
 a12419a <=( a12418a  and  a12413a );
 a12423a <=( A199  and  A166 );
 a12424a <=( A168  and  a12423a );
 a12428a <=( A203  and  A201 );
 a12429a <=( (not A200)  and  a12428a );
 a12430a <=( a12429a  and  a12424a );
 a12434a <=( A267  and  (not A266) );
 a12435a <=( A265  and  a12434a );
 a12439a <=( A299  and  A298 );
 a12440a <=( A268  and  a12439a );
 a12441a <=( a12440a  and  a12435a );
 a12445a <=( A199  and  A166 );
 a12446a <=( A168  and  a12445a );
 a12450a <=( A203  and  A201 );
 a12451a <=( (not A200)  and  a12450a );
 a12452a <=( a12451a  and  a12446a );
 a12456a <=( A267  and  (not A266) );
 a12457a <=( A265  and  a12456a );
 a12461a <=( (not A299)  and  (not A298) );
 a12462a <=( A268  and  a12461a );
 a12463a <=( a12462a  and  a12457a );
 a12467a <=( A199  and  A166 );
 a12468a <=( A168  and  a12467a );
 a12472a <=( A203  and  A201 );
 a12473a <=( (not A200)  and  a12472a );
 a12474a <=( a12473a  and  a12468a );
 a12478a <=( A267  and  (not A266) );
 a12479a <=( A265  and  a12478a );
 a12483a <=( (not A300)  and  A298 );
 a12484a <=( A269  and  a12483a );
 a12485a <=( a12484a  and  a12479a );
 a12489a <=( A199  and  A166 );
 a12490a <=( A168  and  a12489a );
 a12494a <=( A203  and  A201 );
 a12495a <=( (not A200)  and  a12494a );
 a12496a <=( a12495a  and  a12490a );
 a12500a <=( A267  and  (not A266) );
 a12501a <=( A265  and  a12500a );
 a12505a <=( A299  and  A298 );
 a12506a <=( A269  and  a12505a );
 a12507a <=( a12506a  and  a12501a );
 a12511a <=( A199  and  A166 );
 a12512a <=( A168  and  a12511a );
 a12516a <=( A203  and  A201 );
 a12517a <=( (not A200)  and  a12516a );
 a12518a <=( a12517a  and  a12512a );
 a12522a <=( A267  and  (not A266) );
 a12523a <=( A265  and  a12522a );
 a12527a <=( (not A299)  and  (not A298) );
 a12528a <=( A269  and  a12527a );
 a12529a <=( a12528a  and  a12523a );
 a12533a <=( (not A200)  and  A167 );
 a12534a <=( A168  and  a12533a );
 a12538a <=( (not A266)  and  (not A203) );
 a12539a <=( (not A202)  and  a12538a );
 a12540a <=( a12539a  and  a12534a );
 a12544a <=( A298  and  (not A269) );
 a12545a <=( (not A268)  and  a12544a );
 a12549a <=( A301  and  A300 );
 a12550a <=( (not A299)  and  a12549a );
 a12551a <=( a12550a  and  a12545a );
 a12555a <=( (not A200)  and  A167 );
 a12556a <=( A168  and  a12555a );
 a12560a <=( (not A266)  and  (not A203) );
 a12561a <=( (not A202)  and  a12560a );
 a12562a <=( a12561a  and  a12556a );
 a12566a <=( A298  and  (not A269) );
 a12567a <=( (not A268)  and  a12566a );
 a12571a <=( A302  and  A300 );
 a12572a <=( (not A299)  and  a12571a );
 a12573a <=( a12572a  and  a12567a );
 a12577a <=( A199  and  A167 );
 a12578a <=( A168  and  a12577a );
 a12582a <=( A202  and  A201 );
 a12583a <=( (not A200)  and  a12582a );
 a12584a <=( a12583a  and  a12578a );
 a12588a <=( A267  and  (not A266) );
 a12589a <=( A265  and  a12588a );
 a12593a <=( (not A300)  and  A298 );
 a12594a <=( A268  and  a12593a );
 a12595a <=( a12594a  and  a12589a );
 a12599a <=( A199  and  A167 );
 a12600a <=( A168  and  a12599a );
 a12604a <=( A202  and  A201 );
 a12605a <=( (not A200)  and  a12604a );
 a12606a <=( a12605a  and  a12600a );
 a12610a <=( A267  and  (not A266) );
 a12611a <=( A265  and  a12610a );
 a12615a <=( A299  and  A298 );
 a12616a <=( A268  and  a12615a );
 a12617a <=( a12616a  and  a12611a );
 a12621a <=( A199  and  A167 );
 a12622a <=( A168  and  a12621a );
 a12626a <=( A202  and  A201 );
 a12627a <=( (not A200)  and  a12626a );
 a12628a <=( a12627a  and  a12622a );
 a12632a <=( A267  and  (not A266) );
 a12633a <=( A265  and  a12632a );
 a12637a <=( (not A299)  and  (not A298) );
 a12638a <=( A268  and  a12637a );
 a12639a <=( a12638a  and  a12633a );
 a12643a <=( A199  and  A167 );
 a12644a <=( A168  and  a12643a );
 a12648a <=( A202  and  A201 );
 a12649a <=( (not A200)  and  a12648a );
 a12650a <=( a12649a  and  a12644a );
 a12654a <=( A267  and  (not A266) );
 a12655a <=( A265  and  a12654a );
 a12659a <=( (not A300)  and  A298 );
 a12660a <=( A269  and  a12659a );
 a12661a <=( a12660a  and  a12655a );
 a12665a <=( A199  and  A167 );
 a12666a <=( A168  and  a12665a );
 a12670a <=( A202  and  A201 );
 a12671a <=( (not A200)  and  a12670a );
 a12672a <=( a12671a  and  a12666a );
 a12676a <=( A267  and  (not A266) );
 a12677a <=( A265  and  a12676a );
 a12681a <=( A299  and  A298 );
 a12682a <=( A269  and  a12681a );
 a12683a <=( a12682a  and  a12677a );
 a12687a <=( A199  and  A167 );
 a12688a <=( A168  and  a12687a );
 a12692a <=( A202  and  A201 );
 a12693a <=( (not A200)  and  a12692a );
 a12694a <=( a12693a  and  a12688a );
 a12698a <=( A267  and  (not A266) );
 a12699a <=( A265  and  a12698a );
 a12703a <=( (not A299)  and  (not A298) );
 a12704a <=( A269  and  a12703a );
 a12705a <=( a12704a  and  a12699a );
 a12709a <=( A199  and  A167 );
 a12710a <=( A168  and  a12709a );
 a12714a <=( A203  and  A201 );
 a12715a <=( (not A200)  and  a12714a );
 a12716a <=( a12715a  and  a12710a );
 a12720a <=( A267  and  (not A266) );
 a12721a <=( A265  and  a12720a );
 a12725a <=( (not A300)  and  A298 );
 a12726a <=( A268  and  a12725a );
 a12727a <=( a12726a  and  a12721a );
 a12731a <=( A199  and  A167 );
 a12732a <=( A168  and  a12731a );
 a12736a <=( A203  and  A201 );
 a12737a <=( (not A200)  and  a12736a );
 a12738a <=( a12737a  and  a12732a );
 a12742a <=( A267  and  (not A266) );
 a12743a <=( A265  and  a12742a );
 a12747a <=( A299  and  A298 );
 a12748a <=( A268  and  a12747a );
 a12749a <=( a12748a  and  a12743a );
 a12753a <=( A199  and  A167 );
 a12754a <=( A168  and  a12753a );
 a12758a <=( A203  and  A201 );
 a12759a <=( (not A200)  and  a12758a );
 a12760a <=( a12759a  and  a12754a );
 a12764a <=( A267  and  (not A266) );
 a12765a <=( A265  and  a12764a );
 a12769a <=( (not A299)  and  (not A298) );
 a12770a <=( A268  and  a12769a );
 a12771a <=( a12770a  and  a12765a );
 a12775a <=( A199  and  A167 );
 a12776a <=( A168  and  a12775a );
 a12780a <=( A203  and  A201 );
 a12781a <=( (not A200)  and  a12780a );
 a12782a <=( a12781a  and  a12776a );
 a12786a <=( A267  and  (not A266) );
 a12787a <=( A265  and  a12786a );
 a12791a <=( (not A300)  and  A298 );
 a12792a <=( A269  and  a12791a );
 a12793a <=( a12792a  and  a12787a );
 a12797a <=( A199  and  A167 );
 a12798a <=( A168  and  a12797a );
 a12802a <=( A203  and  A201 );
 a12803a <=( (not A200)  and  a12802a );
 a12804a <=( a12803a  and  a12798a );
 a12808a <=( A267  and  (not A266) );
 a12809a <=( A265  and  a12808a );
 a12813a <=( A299  and  A298 );
 a12814a <=( A269  and  a12813a );
 a12815a <=( a12814a  and  a12809a );
 a12819a <=( A199  and  A167 );
 a12820a <=( A168  and  a12819a );
 a12824a <=( A203  and  A201 );
 a12825a <=( (not A200)  and  a12824a );
 a12826a <=( a12825a  and  a12820a );
 a12830a <=( A267  and  (not A266) );
 a12831a <=( A265  and  a12830a );
 a12835a <=( (not A299)  and  (not A298) );
 a12836a <=( A269  and  a12835a );
 a12837a <=( a12836a  and  a12831a );
 a12841a <=( (not A166)  and  (not A167) );
 a12842a <=( A170  and  a12841a );
 a12846a <=( A265  and  A200 );
 a12847a <=( A199  and  a12846a );
 a12848a <=( a12847a  and  a12842a );
 a12852a <=( A268  and  A267 );
 a12853a <=( (not A266)  and  a12852a );
 a12857a <=( (not A302)  and  (not A301) );
 a12858a <=( A298  and  a12857a );
 a12859a <=( a12858a  and  a12853a );
 a12863a <=( (not A166)  and  (not A167) );
 a12864a <=( A170  and  a12863a );
 a12868a <=( A265  and  A200 );
 a12869a <=( A199  and  a12868a );
 a12870a <=( a12869a  and  a12864a );
 a12874a <=( A269  and  A267 );
 a12875a <=( (not A266)  and  a12874a );
 a12879a <=( (not A302)  and  (not A301) );
 a12880a <=( A298  and  a12879a );
 a12881a <=( a12880a  and  a12875a );
 a12885a <=( (not A166)  and  (not A167) );
 a12886a <=( A170  and  a12885a );
 a12890a <=( (not A266)  and  A200 );
 a12891a <=( (not A199)  and  a12890a );
 a12892a <=( a12891a  and  a12886a );
 a12896a <=( A298  and  (not A269) );
 a12897a <=( (not A268)  and  a12896a );
 a12901a <=( A301  and  A300 );
 a12902a <=( (not A299)  and  a12901a );
 a12903a <=( a12902a  and  a12897a );
 a12907a <=( (not A166)  and  (not A167) );
 a12908a <=( A170  and  a12907a );
 a12912a <=( (not A266)  and  A200 );
 a12913a <=( (not A199)  and  a12912a );
 a12914a <=( a12913a  and  a12908a );
 a12918a <=( A298  and  (not A269) );
 a12919a <=( (not A268)  and  a12918a );
 a12923a <=( A302  and  A300 );
 a12924a <=( (not A299)  and  a12923a );
 a12925a <=( a12924a  and  a12919a );
 a12929a <=( (not A166)  and  (not A167) );
 a12930a <=( A170  and  a12929a );
 a12934a <=( (not A203)  and  (not A202) );
 a12935a <=( (not A200)  and  a12934a );
 a12936a <=( a12935a  and  a12930a );
 a12940a <=( A267  and  (not A266) );
 a12941a <=( A265  and  a12940a );
 a12945a <=( (not A300)  and  A298 );
 a12946a <=( A268  and  a12945a );
 a12947a <=( a12946a  and  a12941a );
 a12951a <=( (not A166)  and  (not A167) );
 a12952a <=( A170  and  a12951a );
 a12956a <=( (not A203)  and  (not A202) );
 a12957a <=( (not A200)  and  a12956a );
 a12958a <=( a12957a  and  a12952a );
 a12962a <=( A267  and  (not A266) );
 a12963a <=( A265  and  a12962a );
 a12967a <=( A299  and  A298 );
 a12968a <=( A268  and  a12967a );
 a12969a <=( a12968a  and  a12963a );
 a12973a <=( (not A166)  and  (not A167) );
 a12974a <=( A170  and  a12973a );
 a12978a <=( (not A203)  and  (not A202) );
 a12979a <=( (not A200)  and  a12978a );
 a12980a <=( a12979a  and  a12974a );
 a12984a <=( A267  and  (not A266) );
 a12985a <=( A265  and  a12984a );
 a12989a <=( (not A299)  and  (not A298) );
 a12990a <=( A268  and  a12989a );
 a12991a <=( a12990a  and  a12985a );
 a12995a <=( (not A166)  and  (not A167) );
 a12996a <=( A170  and  a12995a );
 a13000a <=( (not A203)  and  (not A202) );
 a13001a <=( (not A200)  and  a13000a );
 a13002a <=( a13001a  and  a12996a );
 a13006a <=( A267  and  (not A266) );
 a13007a <=( A265  and  a13006a );
 a13011a <=( (not A300)  and  A298 );
 a13012a <=( A269  and  a13011a );
 a13013a <=( a13012a  and  a13007a );
 a13017a <=( (not A166)  and  (not A167) );
 a13018a <=( A170  and  a13017a );
 a13022a <=( (not A203)  and  (not A202) );
 a13023a <=( (not A200)  and  a13022a );
 a13024a <=( a13023a  and  a13018a );
 a13028a <=( A267  and  (not A266) );
 a13029a <=( A265  and  a13028a );
 a13033a <=( A299  and  A298 );
 a13034a <=( A269  and  a13033a );
 a13035a <=( a13034a  and  a13029a );
 a13039a <=( (not A166)  and  (not A167) );
 a13040a <=( A170  and  a13039a );
 a13044a <=( (not A203)  and  (not A202) );
 a13045a <=( (not A200)  and  a13044a );
 a13046a <=( a13045a  and  a13040a );
 a13050a <=( A267  and  (not A266) );
 a13051a <=( A265  and  a13050a );
 a13055a <=( (not A299)  and  (not A298) );
 a13056a <=( A269  and  a13055a );
 a13057a <=( a13056a  and  a13051a );
 a13061a <=( (not A166)  and  (not A167) );
 a13062a <=( A170  and  a13061a );
 a13066a <=( A265  and  (not A201) );
 a13067a <=( (not A200)  and  a13066a );
 a13068a <=( a13067a  and  a13062a );
 a13072a <=( A268  and  A267 );
 a13073a <=( (not A266)  and  a13072a );
 a13077a <=( (not A302)  and  (not A301) );
 a13078a <=( A298  and  a13077a );
 a13079a <=( a13078a  and  a13073a );
 a13083a <=( (not A166)  and  (not A167) );
 a13084a <=( A170  and  a13083a );
 a13088a <=( A265  and  (not A201) );
 a13089a <=( (not A200)  and  a13088a );
 a13090a <=( a13089a  and  a13084a );
 a13094a <=( A269  and  A267 );
 a13095a <=( (not A266)  and  a13094a );
 a13099a <=( (not A302)  and  (not A301) );
 a13100a <=( A298  and  a13099a );
 a13101a <=( a13100a  and  a13095a );
 a13105a <=( (not A166)  and  (not A167) );
 a13106a <=( A170  and  a13105a );
 a13110a <=( A201  and  (not A200) );
 a13111a <=( A199  and  a13110a );
 a13112a <=( a13111a  and  a13106a );
 a13116a <=( (not A268)  and  (not A266) );
 a13117a <=( A202  and  a13116a );
 a13121a <=( A299  and  (not A298) );
 a13122a <=( (not A269)  and  a13121a );
 a13123a <=( a13122a  and  a13117a );
 a13127a <=( (not A166)  and  (not A167) );
 a13128a <=( A170  and  a13127a );
 a13132a <=( A201  and  (not A200) );
 a13133a <=( A199  and  a13132a );
 a13134a <=( a13133a  and  a13128a );
 a13138a <=( (not A268)  and  (not A266) );
 a13139a <=( A203  and  a13138a );
 a13143a <=( A299  and  (not A298) );
 a13144a <=( (not A269)  and  a13143a );
 a13145a <=( a13144a  and  a13139a );
 a13149a <=( (not A166)  and  (not A167) );
 a13150a <=( A170  and  a13149a );
 a13154a <=( A265  and  (not A200) );
 a13155a <=( (not A199)  and  a13154a );
 a13156a <=( a13155a  and  a13150a );
 a13160a <=( A268  and  A267 );
 a13161a <=( (not A266)  and  a13160a );
 a13165a <=( (not A302)  and  (not A301) );
 a13166a <=( A298  and  a13165a );
 a13167a <=( a13166a  and  a13161a );
 a13171a <=( (not A166)  and  (not A167) );
 a13172a <=( A170  and  a13171a );
 a13176a <=( A265  and  (not A200) );
 a13177a <=( (not A199)  and  a13176a );
 a13178a <=( a13177a  and  a13172a );
 a13182a <=( A269  and  A267 );
 a13183a <=( (not A266)  and  a13182a );
 a13187a <=( (not A302)  and  (not A301) );
 a13188a <=( A298  and  a13187a );
 a13189a <=( a13188a  and  a13183a );
 a13193a <=( A167  and  (not A168) );
 a13194a <=( A169  and  a13193a );
 a13198a <=( A200  and  A199 );
 a13199a <=( (not A166)  and  a13198a );
 a13200a <=( a13199a  and  a13194a );
 a13204a <=( A267  and  (not A266) );
 a13205a <=( A265  and  a13204a );
 a13209a <=( (not A300)  and  A298 );
 a13210a <=( A268  and  a13209a );
 a13211a <=( a13210a  and  a13205a );
 a13215a <=( A167  and  (not A168) );
 a13216a <=( A169  and  a13215a );
 a13220a <=( A200  and  A199 );
 a13221a <=( (not A166)  and  a13220a );
 a13222a <=( a13221a  and  a13216a );
 a13226a <=( A267  and  (not A266) );
 a13227a <=( A265  and  a13226a );
 a13231a <=( A299  and  A298 );
 a13232a <=( A268  and  a13231a );
 a13233a <=( a13232a  and  a13227a );
 a13237a <=( A167  and  (not A168) );
 a13238a <=( A169  and  a13237a );
 a13242a <=( A200  and  A199 );
 a13243a <=( (not A166)  and  a13242a );
 a13244a <=( a13243a  and  a13238a );
 a13248a <=( A267  and  (not A266) );
 a13249a <=( A265  and  a13248a );
 a13253a <=( (not A299)  and  (not A298) );
 a13254a <=( A268  and  a13253a );
 a13255a <=( a13254a  and  a13249a );
 a13259a <=( A167  and  (not A168) );
 a13260a <=( A169  and  a13259a );
 a13264a <=( A200  and  A199 );
 a13265a <=( (not A166)  and  a13264a );
 a13266a <=( a13265a  and  a13260a );
 a13270a <=( A267  and  (not A266) );
 a13271a <=( A265  and  a13270a );
 a13275a <=( (not A300)  and  A298 );
 a13276a <=( A269  and  a13275a );
 a13277a <=( a13276a  and  a13271a );
 a13281a <=( A167  and  (not A168) );
 a13282a <=( A169  and  a13281a );
 a13286a <=( A200  and  A199 );
 a13287a <=( (not A166)  and  a13286a );
 a13288a <=( a13287a  and  a13282a );
 a13292a <=( A267  and  (not A266) );
 a13293a <=( A265  and  a13292a );
 a13297a <=( A299  and  A298 );
 a13298a <=( A269  and  a13297a );
 a13299a <=( a13298a  and  a13293a );
 a13303a <=( A167  and  (not A168) );
 a13304a <=( A169  and  a13303a );
 a13308a <=( A200  and  A199 );
 a13309a <=( (not A166)  and  a13308a );
 a13310a <=( a13309a  and  a13304a );
 a13314a <=( A267  and  (not A266) );
 a13315a <=( A265  and  a13314a );
 a13319a <=( (not A299)  and  (not A298) );
 a13320a <=( A269  and  a13319a );
 a13321a <=( a13320a  and  a13315a );
 a13325a <=( A167  and  (not A168) );
 a13326a <=( A169  and  a13325a );
 a13330a <=( A200  and  (not A199) );
 a13331a <=( (not A166)  and  a13330a );
 a13332a <=( a13331a  and  a13326a );
 a13336a <=( A298  and  A266 );
 a13337a <=( A265  and  a13336a );
 a13341a <=( A301  and  A300 );
 a13342a <=( (not A299)  and  a13341a );
 a13343a <=( a13342a  and  a13337a );
 a13347a <=( A167  and  (not A168) );
 a13348a <=( A169  and  a13347a );
 a13352a <=( A200  and  (not A199) );
 a13353a <=( (not A166)  and  a13352a );
 a13354a <=( a13353a  and  a13348a );
 a13358a <=( A298  and  A266 );
 a13359a <=( A265  and  a13358a );
 a13363a <=( A302  and  A300 );
 a13364a <=( (not A299)  and  a13363a );
 a13365a <=( a13364a  and  a13359a );
 a13369a <=( A167  and  (not A168) );
 a13370a <=( A169  and  a13369a );
 a13374a <=( A200  and  (not A199) );
 a13375a <=( (not A166)  and  a13374a );
 a13376a <=( a13375a  and  a13370a );
 a13380a <=( A298  and  (not A267) );
 a13381a <=( (not A266)  and  a13380a );
 a13385a <=( A301  and  A300 );
 a13386a <=( (not A299)  and  a13385a );
 a13387a <=( a13386a  and  a13381a );
 a13391a <=( A167  and  (not A168) );
 a13392a <=( A169  and  a13391a );
 a13396a <=( A200  and  (not A199) );
 a13397a <=( (not A166)  and  a13396a );
 a13398a <=( a13397a  and  a13392a );
 a13402a <=( A298  and  (not A267) );
 a13403a <=( (not A266)  and  a13402a );
 a13407a <=( A302  and  A300 );
 a13408a <=( (not A299)  and  a13407a );
 a13409a <=( a13408a  and  a13403a );
 a13413a <=( A167  and  (not A168) );
 a13414a <=( A169  and  a13413a );
 a13418a <=( A200  and  (not A199) );
 a13419a <=( (not A166)  and  a13418a );
 a13420a <=( a13419a  and  a13414a );
 a13424a <=( A298  and  (not A266) );
 a13425a <=( (not A265)  and  a13424a );
 a13429a <=( A301  and  A300 );
 a13430a <=( (not A299)  and  a13429a );
 a13431a <=( a13430a  and  a13425a );
 a13435a <=( A167  and  (not A168) );
 a13436a <=( A169  and  a13435a );
 a13440a <=( A200  and  (not A199) );
 a13441a <=( (not A166)  and  a13440a );
 a13442a <=( a13441a  and  a13436a );
 a13446a <=( A298  and  (not A266) );
 a13447a <=( (not A265)  and  a13446a );
 a13451a <=( A302  and  A300 );
 a13452a <=( (not A299)  and  a13451a );
 a13453a <=( a13452a  and  a13447a );
 a13457a <=( A167  and  (not A168) );
 a13458a <=( A169  and  a13457a );
 a13462a <=( (not A202)  and  (not A200) );
 a13463a <=( (not A166)  and  a13462a );
 a13464a <=( a13463a  and  a13458a );
 a13468a <=( A266  and  (not A265) );
 a13469a <=( (not A203)  and  a13468a );
 a13473a <=( (not A302)  and  (not A301) );
 a13474a <=( A298  and  a13473a );
 a13475a <=( a13474a  and  a13469a );
 a13479a <=( A167  and  (not A168) );
 a13480a <=( A169  and  a13479a );
 a13484a <=( (not A201)  and  (not A200) );
 a13485a <=( (not A166)  and  a13484a );
 a13486a <=( a13485a  and  a13480a );
 a13490a <=( A267  and  (not A266) );
 a13491a <=( A265  and  a13490a );
 a13495a <=( (not A300)  and  A298 );
 a13496a <=( A268  and  a13495a );
 a13497a <=( a13496a  and  a13491a );
 a13501a <=( A167  and  (not A168) );
 a13502a <=( A169  and  a13501a );
 a13506a <=( (not A201)  and  (not A200) );
 a13507a <=( (not A166)  and  a13506a );
 a13508a <=( a13507a  and  a13502a );
 a13512a <=( A267  and  (not A266) );
 a13513a <=( A265  and  a13512a );
 a13517a <=( A299  and  A298 );
 a13518a <=( A268  and  a13517a );
 a13519a <=( a13518a  and  a13513a );
 a13523a <=( A167  and  (not A168) );
 a13524a <=( A169  and  a13523a );
 a13528a <=( (not A201)  and  (not A200) );
 a13529a <=( (not A166)  and  a13528a );
 a13530a <=( a13529a  and  a13524a );
 a13534a <=( A267  and  (not A266) );
 a13535a <=( A265  and  a13534a );
 a13539a <=( (not A299)  and  (not A298) );
 a13540a <=( A268  and  a13539a );
 a13541a <=( a13540a  and  a13535a );
 a13545a <=( A167  and  (not A168) );
 a13546a <=( A169  and  a13545a );
 a13550a <=( (not A201)  and  (not A200) );
 a13551a <=( (not A166)  and  a13550a );
 a13552a <=( a13551a  and  a13546a );
 a13556a <=( A267  and  (not A266) );
 a13557a <=( A265  and  a13556a );
 a13561a <=( (not A300)  and  A298 );
 a13562a <=( A269  and  a13561a );
 a13563a <=( a13562a  and  a13557a );
 a13567a <=( A167  and  (not A168) );
 a13568a <=( A169  and  a13567a );
 a13572a <=( (not A201)  and  (not A200) );
 a13573a <=( (not A166)  and  a13572a );
 a13574a <=( a13573a  and  a13568a );
 a13578a <=( A267  and  (not A266) );
 a13579a <=( A265  and  a13578a );
 a13583a <=( A299  and  A298 );
 a13584a <=( A269  and  a13583a );
 a13585a <=( a13584a  and  a13579a );
 a13589a <=( A167  and  (not A168) );
 a13590a <=( A169  and  a13589a );
 a13594a <=( (not A201)  and  (not A200) );
 a13595a <=( (not A166)  and  a13594a );
 a13596a <=( a13595a  and  a13590a );
 a13600a <=( A267  and  (not A266) );
 a13601a <=( A265  and  a13600a );
 a13605a <=( (not A299)  and  (not A298) );
 a13606a <=( A269  and  a13605a );
 a13607a <=( a13606a  and  a13601a );
 a13611a <=( A167  and  (not A168) );
 a13612a <=( A169  and  a13611a );
 a13616a <=( (not A200)  and  A199 );
 a13617a <=( (not A166)  and  a13616a );
 a13618a <=( a13617a  and  a13612a );
 a13622a <=( A265  and  A202 );
 a13623a <=( A201  and  a13622a );
 a13627a <=( A299  and  (not A298) );
 a13628a <=( A266  and  a13627a );
 a13629a <=( a13628a  and  a13623a );
 a13633a <=( A167  and  (not A168) );
 a13634a <=( A169  and  a13633a );
 a13638a <=( (not A200)  and  A199 );
 a13639a <=( (not A166)  and  a13638a );
 a13640a <=( a13639a  and  a13634a );
 a13644a <=( (not A266)  and  A202 );
 a13645a <=( A201  and  a13644a );
 a13649a <=( A299  and  (not A298) );
 a13650a <=( (not A267)  and  a13649a );
 a13651a <=( a13650a  and  a13645a );
 a13655a <=( A167  and  (not A168) );
 a13656a <=( A169  and  a13655a );
 a13660a <=( (not A200)  and  A199 );
 a13661a <=( (not A166)  and  a13660a );
 a13662a <=( a13661a  and  a13656a );
 a13666a <=( (not A265)  and  A202 );
 a13667a <=( A201  and  a13666a );
 a13671a <=( A299  and  (not A298) );
 a13672a <=( (not A266)  and  a13671a );
 a13673a <=( a13672a  and  a13667a );
 a13677a <=( A167  and  (not A168) );
 a13678a <=( A169  and  a13677a );
 a13682a <=( (not A200)  and  A199 );
 a13683a <=( (not A166)  and  a13682a );
 a13684a <=( a13683a  and  a13678a );
 a13688a <=( A265  and  A203 );
 a13689a <=( A201  and  a13688a );
 a13693a <=( A299  and  (not A298) );
 a13694a <=( A266  and  a13693a );
 a13695a <=( a13694a  and  a13689a );
 a13699a <=( A167  and  (not A168) );
 a13700a <=( A169  and  a13699a );
 a13704a <=( (not A200)  and  A199 );
 a13705a <=( (not A166)  and  a13704a );
 a13706a <=( a13705a  and  a13700a );
 a13710a <=( (not A266)  and  A203 );
 a13711a <=( A201  and  a13710a );
 a13715a <=( A299  and  (not A298) );
 a13716a <=( (not A267)  and  a13715a );
 a13717a <=( a13716a  and  a13711a );
 a13721a <=( A167  and  (not A168) );
 a13722a <=( A169  and  a13721a );
 a13726a <=( (not A200)  and  A199 );
 a13727a <=( (not A166)  and  a13726a );
 a13728a <=( a13727a  and  a13722a );
 a13732a <=( (not A265)  and  A203 );
 a13733a <=( A201  and  a13732a );
 a13737a <=( A299  and  (not A298) );
 a13738a <=( (not A266)  and  a13737a );
 a13739a <=( a13738a  and  a13733a );
 a13743a <=( A167  and  (not A168) );
 a13744a <=( A169  and  a13743a );
 a13748a <=( (not A200)  and  (not A199) );
 a13749a <=( (not A166)  and  a13748a );
 a13750a <=( a13749a  and  a13744a );
 a13754a <=( A267  and  (not A266) );
 a13755a <=( A265  and  a13754a );
 a13759a <=( (not A300)  and  A298 );
 a13760a <=( A268  and  a13759a );
 a13761a <=( a13760a  and  a13755a );
 a13765a <=( A167  and  (not A168) );
 a13766a <=( A169  and  a13765a );
 a13770a <=( (not A200)  and  (not A199) );
 a13771a <=( (not A166)  and  a13770a );
 a13772a <=( a13771a  and  a13766a );
 a13776a <=( A267  and  (not A266) );
 a13777a <=( A265  and  a13776a );
 a13781a <=( A299  and  A298 );
 a13782a <=( A268  and  a13781a );
 a13783a <=( a13782a  and  a13777a );
 a13787a <=( A167  and  (not A168) );
 a13788a <=( A169  and  a13787a );
 a13792a <=( (not A200)  and  (not A199) );
 a13793a <=( (not A166)  and  a13792a );
 a13794a <=( a13793a  and  a13788a );
 a13798a <=( A267  and  (not A266) );
 a13799a <=( A265  and  a13798a );
 a13803a <=( (not A299)  and  (not A298) );
 a13804a <=( A268  and  a13803a );
 a13805a <=( a13804a  and  a13799a );
 a13809a <=( A167  and  (not A168) );
 a13810a <=( A169  and  a13809a );
 a13814a <=( (not A200)  and  (not A199) );
 a13815a <=( (not A166)  and  a13814a );
 a13816a <=( a13815a  and  a13810a );
 a13820a <=( A267  and  (not A266) );
 a13821a <=( A265  and  a13820a );
 a13825a <=( (not A300)  and  A298 );
 a13826a <=( A269  and  a13825a );
 a13827a <=( a13826a  and  a13821a );
 a13831a <=( A167  and  (not A168) );
 a13832a <=( A169  and  a13831a );
 a13836a <=( (not A200)  and  (not A199) );
 a13837a <=( (not A166)  and  a13836a );
 a13838a <=( a13837a  and  a13832a );
 a13842a <=( A267  and  (not A266) );
 a13843a <=( A265  and  a13842a );
 a13847a <=( A299  and  A298 );
 a13848a <=( A269  and  a13847a );
 a13849a <=( a13848a  and  a13843a );
 a13853a <=( A167  and  (not A168) );
 a13854a <=( A169  and  a13853a );
 a13858a <=( (not A200)  and  (not A199) );
 a13859a <=( (not A166)  and  a13858a );
 a13860a <=( a13859a  and  a13854a );
 a13864a <=( A267  and  (not A266) );
 a13865a <=( A265  and  a13864a );
 a13869a <=( (not A299)  and  (not A298) );
 a13870a <=( A269  and  a13869a );
 a13871a <=( a13870a  and  a13865a );
 a13875a <=( (not A167)  and  (not A168) );
 a13876a <=( A169  and  a13875a );
 a13880a <=( A200  and  A199 );
 a13881a <=( A166  and  a13880a );
 a13882a <=( a13881a  and  a13876a );
 a13886a <=( A267  and  (not A266) );
 a13887a <=( A265  and  a13886a );
 a13891a <=( (not A300)  and  A298 );
 a13892a <=( A268  and  a13891a );
 a13893a <=( a13892a  and  a13887a );
 a13897a <=( (not A167)  and  (not A168) );
 a13898a <=( A169  and  a13897a );
 a13902a <=( A200  and  A199 );
 a13903a <=( A166  and  a13902a );
 a13904a <=( a13903a  and  a13898a );
 a13908a <=( A267  and  (not A266) );
 a13909a <=( A265  and  a13908a );
 a13913a <=( A299  and  A298 );
 a13914a <=( A268  and  a13913a );
 a13915a <=( a13914a  and  a13909a );
 a13919a <=( (not A167)  and  (not A168) );
 a13920a <=( A169  and  a13919a );
 a13924a <=( A200  and  A199 );
 a13925a <=( A166  and  a13924a );
 a13926a <=( a13925a  and  a13920a );
 a13930a <=( A267  and  (not A266) );
 a13931a <=( A265  and  a13930a );
 a13935a <=( (not A299)  and  (not A298) );
 a13936a <=( A268  and  a13935a );
 a13937a <=( a13936a  and  a13931a );
 a13941a <=( (not A167)  and  (not A168) );
 a13942a <=( A169  and  a13941a );
 a13946a <=( A200  and  A199 );
 a13947a <=( A166  and  a13946a );
 a13948a <=( a13947a  and  a13942a );
 a13952a <=( A267  and  (not A266) );
 a13953a <=( A265  and  a13952a );
 a13957a <=( (not A300)  and  A298 );
 a13958a <=( A269  and  a13957a );
 a13959a <=( a13958a  and  a13953a );
 a13963a <=( (not A167)  and  (not A168) );
 a13964a <=( A169  and  a13963a );
 a13968a <=( A200  and  A199 );
 a13969a <=( A166  and  a13968a );
 a13970a <=( a13969a  and  a13964a );
 a13974a <=( A267  and  (not A266) );
 a13975a <=( A265  and  a13974a );
 a13979a <=( A299  and  A298 );
 a13980a <=( A269  and  a13979a );
 a13981a <=( a13980a  and  a13975a );
 a13985a <=( (not A167)  and  (not A168) );
 a13986a <=( A169  and  a13985a );
 a13990a <=( A200  and  A199 );
 a13991a <=( A166  and  a13990a );
 a13992a <=( a13991a  and  a13986a );
 a13996a <=( A267  and  (not A266) );
 a13997a <=( A265  and  a13996a );
 a14001a <=( (not A299)  and  (not A298) );
 a14002a <=( A269  and  a14001a );
 a14003a <=( a14002a  and  a13997a );
 a14007a <=( (not A167)  and  (not A168) );
 a14008a <=( A169  and  a14007a );
 a14012a <=( A200  and  (not A199) );
 a14013a <=( A166  and  a14012a );
 a14014a <=( a14013a  and  a14008a );
 a14018a <=( A298  and  A266 );
 a14019a <=( A265  and  a14018a );
 a14023a <=( A301  and  A300 );
 a14024a <=( (not A299)  and  a14023a );
 a14025a <=( a14024a  and  a14019a );
 a14029a <=( (not A167)  and  (not A168) );
 a14030a <=( A169  and  a14029a );
 a14034a <=( A200  and  (not A199) );
 a14035a <=( A166  and  a14034a );
 a14036a <=( a14035a  and  a14030a );
 a14040a <=( A298  and  A266 );
 a14041a <=( A265  and  a14040a );
 a14045a <=( A302  and  A300 );
 a14046a <=( (not A299)  and  a14045a );
 a14047a <=( a14046a  and  a14041a );
 a14051a <=( (not A167)  and  (not A168) );
 a14052a <=( A169  and  a14051a );
 a14056a <=( A200  and  (not A199) );
 a14057a <=( A166  and  a14056a );
 a14058a <=( a14057a  and  a14052a );
 a14062a <=( A298  and  (not A267) );
 a14063a <=( (not A266)  and  a14062a );
 a14067a <=( A301  and  A300 );
 a14068a <=( (not A299)  and  a14067a );
 a14069a <=( a14068a  and  a14063a );
 a14073a <=( (not A167)  and  (not A168) );
 a14074a <=( A169  and  a14073a );
 a14078a <=( A200  and  (not A199) );
 a14079a <=( A166  and  a14078a );
 a14080a <=( a14079a  and  a14074a );
 a14084a <=( A298  and  (not A267) );
 a14085a <=( (not A266)  and  a14084a );
 a14089a <=( A302  and  A300 );
 a14090a <=( (not A299)  and  a14089a );
 a14091a <=( a14090a  and  a14085a );
 a14095a <=( (not A167)  and  (not A168) );
 a14096a <=( A169  and  a14095a );
 a14100a <=( A200  and  (not A199) );
 a14101a <=( A166  and  a14100a );
 a14102a <=( a14101a  and  a14096a );
 a14106a <=( A298  and  (not A266) );
 a14107a <=( (not A265)  and  a14106a );
 a14111a <=( A301  and  A300 );
 a14112a <=( (not A299)  and  a14111a );
 a14113a <=( a14112a  and  a14107a );
 a14117a <=( (not A167)  and  (not A168) );
 a14118a <=( A169  and  a14117a );
 a14122a <=( A200  and  (not A199) );
 a14123a <=( A166  and  a14122a );
 a14124a <=( a14123a  and  a14118a );
 a14128a <=( A298  and  (not A266) );
 a14129a <=( (not A265)  and  a14128a );
 a14133a <=( A302  and  A300 );
 a14134a <=( (not A299)  and  a14133a );
 a14135a <=( a14134a  and  a14129a );
 a14139a <=( (not A167)  and  (not A168) );
 a14140a <=( A169  and  a14139a );
 a14144a <=( (not A202)  and  (not A200) );
 a14145a <=( A166  and  a14144a );
 a14146a <=( a14145a  and  a14140a );
 a14150a <=( A266  and  (not A265) );
 a14151a <=( (not A203)  and  a14150a );
 a14155a <=( (not A302)  and  (not A301) );
 a14156a <=( A298  and  a14155a );
 a14157a <=( a14156a  and  a14151a );
 a14161a <=( (not A167)  and  (not A168) );
 a14162a <=( A169  and  a14161a );
 a14166a <=( (not A201)  and  (not A200) );
 a14167a <=( A166  and  a14166a );
 a14168a <=( a14167a  and  a14162a );
 a14172a <=( A267  and  (not A266) );
 a14173a <=( A265  and  a14172a );
 a14177a <=( (not A300)  and  A298 );
 a14178a <=( A268  and  a14177a );
 a14179a <=( a14178a  and  a14173a );
 a14183a <=( (not A167)  and  (not A168) );
 a14184a <=( A169  and  a14183a );
 a14188a <=( (not A201)  and  (not A200) );
 a14189a <=( A166  and  a14188a );
 a14190a <=( a14189a  and  a14184a );
 a14194a <=( A267  and  (not A266) );
 a14195a <=( A265  and  a14194a );
 a14199a <=( A299  and  A298 );
 a14200a <=( A268  and  a14199a );
 a14201a <=( a14200a  and  a14195a );
 a14205a <=( (not A167)  and  (not A168) );
 a14206a <=( A169  and  a14205a );
 a14210a <=( (not A201)  and  (not A200) );
 a14211a <=( A166  and  a14210a );
 a14212a <=( a14211a  and  a14206a );
 a14216a <=( A267  and  (not A266) );
 a14217a <=( A265  and  a14216a );
 a14221a <=( (not A299)  and  (not A298) );
 a14222a <=( A268  and  a14221a );
 a14223a <=( a14222a  and  a14217a );
 a14227a <=( (not A167)  and  (not A168) );
 a14228a <=( A169  and  a14227a );
 a14232a <=( (not A201)  and  (not A200) );
 a14233a <=( A166  and  a14232a );
 a14234a <=( a14233a  and  a14228a );
 a14238a <=( A267  and  (not A266) );
 a14239a <=( A265  and  a14238a );
 a14243a <=( (not A300)  and  A298 );
 a14244a <=( A269  and  a14243a );
 a14245a <=( a14244a  and  a14239a );
 a14249a <=( (not A167)  and  (not A168) );
 a14250a <=( A169  and  a14249a );
 a14254a <=( (not A201)  and  (not A200) );
 a14255a <=( A166  and  a14254a );
 a14256a <=( a14255a  and  a14250a );
 a14260a <=( A267  and  (not A266) );
 a14261a <=( A265  and  a14260a );
 a14265a <=( A299  and  A298 );
 a14266a <=( A269  and  a14265a );
 a14267a <=( a14266a  and  a14261a );
 a14271a <=( (not A167)  and  (not A168) );
 a14272a <=( A169  and  a14271a );
 a14276a <=( (not A201)  and  (not A200) );
 a14277a <=( A166  and  a14276a );
 a14278a <=( a14277a  and  a14272a );
 a14282a <=( A267  and  (not A266) );
 a14283a <=( A265  and  a14282a );
 a14287a <=( (not A299)  and  (not A298) );
 a14288a <=( A269  and  a14287a );
 a14289a <=( a14288a  and  a14283a );
 a14293a <=( (not A167)  and  (not A168) );
 a14294a <=( A169  and  a14293a );
 a14298a <=( (not A200)  and  A199 );
 a14299a <=( A166  and  a14298a );
 a14300a <=( a14299a  and  a14294a );
 a14304a <=( A265  and  A202 );
 a14305a <=( A201  and  a14304a );
 a14309a <=( A299  and  (not A298) );
 a14310a <=( A266  and  a14309a );
 a14311a <=( a14310a  and  a14305a );
 a14315a <=( (not A167)  and  (not A168) );
 a14316a <=( A169  and  a14315a );
 a14320a <=( (not A200)  and  A199 );
 a14321a <=( A166  and  a14320a );
 a14322a <=( a14321a  and  a14316a );
 a14326a <=( (not A266)  and  A202 );
 a14327a <=( A201  and  a14326a );
 a14331a <=( A299  and  (not A298) );
 a14332a <=( (not A267)  and  a14331a );
 a14333a <=( a14332a  and  a14327a );
 a14337a <=( (not A167)  and  (not A168) );
 a14338a <=( A169  and  a14337a );
 a14342a <=( (not A200)  and  A199 );
 a14343a <=( A166  and  a14342a );
 a14344a <=( a14343a  and  a14338a );
 a14348a <=( (not A265)  and  A202 );
 a14349a <=( A201  and  a14348a );
 a14353a <=( A299  and  (not A298) );
 a14354a <=( (not A266)  and  a14353a );
 a14355a <=( a14354a  and  a14349a );
 a14359a <=( (not A167)  and  (not A168) );
 a14360a <=( A169  and  a14359a );
 a14364a <=( (not A200)  and  A199 );
 a14365a <=( A166  and  a14364a );
 a14366a <=( a14365a  and  a14360a );
 a14370a <=( A265  and  A203 );
 a14371a <=( A201  and  a14370a );
 a14375a <=( A299  and  (not A298) );
 a14376a <=( A266  and  a14375a );
 a14377a <=( a14376a  and  a14371a );
 a14381a <=( (not A167)  and  (not A168) );
 a14382a <=( A169  and  a14381a );
 a14386a <=( (not A200)  and  A199 );
 a14387a <=( A166  and  a14386a );
 a14388a <=( a14387a  and  a14382a );
 a14392a <=( (not A266)  and  A203 );
 a14393a <=( A201  and  a14392a );
 a14397a <=( A299  and  (not A298) );
 a14398a <=( (not A267)  and  a14397a );
 a14399a <=( a14398a  and  a14393a );
 a14403a <=( (not A167)  and  (not A168) );
 a14404a <=( A169  and  a14403a );
 a14408a <=( (not A200)  and  A199 );
 a14409a <=( A166  and  a14408a );
 a14410a <=( a14409a  and  a14404a );
 a14414a <=( (not A265)  and  A203 );
 a14415a <=( A201  and  a14414a );
 a14419a <=( A299  and  (not A298) );
 a14420a <=( (not A266)  and  a14419a );
 a14421a <=( a14420a  and  a14415a );
 a14425a <=( (not A167)  and  (not A168) );
 a14426a <=( A169  and  a14425a );
 a14430a <=( (not A200)  and  (not A199) );
 a14431a <=( A166  and  a14430a );
 a14432a <=( a14431a  and  a14426a );
 a14436a <=( A267  and  (not A266) );
 a14437a <=( A265  and  a14436a );
 a14441a <=( (not A300)  and  A298 );
 a14442a <=( A268  and  a14441a );
 a14443a <=( a14442a  and  a14437a );
 a14447a <=( (not A167)  and  (not A168) );
 a14448a <=( A169  and  a14447a );
 a14452a <=( (not A200)  and  (not A199) );
 a14453a <=( A166  and  a14452a );
 a14454a <=( a14453a  and  a14448a );
 a14458a <=( A267  and  (not A266) );
 a14459a <=( A265  and  a14458a );
 a14463a <=( A299  and  A298 );
 a14464a <=( A268  and  a14463a );
 a14465a <=( a14464a  and  a14459a );
 a14469a <=( (not A167)  and  (not A168) );
 a14470a <=( A169  and  a14469a );
 a14474a <=( (not A200)  and  (not A199) );
 a14475a <=( A166  and  a14474a );
 a14476a <=( a14475a  and  a14470a );
 a14480a <=( A267  and  (not A266) );
 a14481a <=( A265  and  a14480a );
 a14485a <=( (not A299)  and  (not A298) );
 a14486a <=( A268  and  a14485a );
 a14487a <=( a14486a  and  a14481a );
 a14491a <=( (not A167)  and  (not A168) );
 a14492a <=( A169  and  a14491a );
 a14496a <=( (not A200)  and  (not A199) );
 a14497a <=( A166  and  a14496a );
 a14498a <=( a14497a  and  a14492a );
 a14502a <=( A267  and  (not A266) );
 a14503a <=( A265  and  a14502a );
 a14507a <=( (not A300)  and  A298 );
 a14508a <=( A269  and  a14507a );
 a14509a <=( a14508a  and  a14503a );
 a14513a <=( (not A167)  and  (not A168) );
 a14514a <=( A169  and  a14513a );
 a14518a <=( (not A200)  and  (not A199) );
 a14519a <=( A166  and  a14518a );
 a14520a <=( a14519a  and  a14514a );
 a14524a <=( A267  and  (not A266) );
 a14525a <=( A265  and  a14524a );
 a14529a <=( A299  and  A298 );
 a14530a <=( A269  and  a14529a );
 a14531a <=( a14530a  and  a14525a );
 a14535a <=( (not A167)  and  (not A168) );
 a14536a <=( A169  and  a14535a );
 a14540a <=( (not A200)  and  (not A199) );
 a14541a <=( A166  and  a14540a );
 a14542a <=( a14541a  and  a14536a );
 a14546a <=( A267  and  (not A266) );
 a14547a <=( A265  and  a14546a );
 a14551a <=( (not A299)  and  (not A298) );
 a14552a <=( A269  and  a14551a );
 a14553a <=( a14552a  and  a14547a );
 a14557a <=( (not A168)  and  A169 );
 a14558a <=( A170  and  a14557a );
 a14562a <=( A265  and  A200 );
 a14563a <=( A199  and  a14562a );
 a14564a <=( a14563a  and  a14558a );
 a14568a <=( A268  and  A267 );
 a14569a <=( (not A266)  and  a14568a );
 a14573a <=( (not A302)  and  (not A301) );
 a14574a <=( A298  and  a14573a );
 a14575a <=( a14574a  and  a14569a );
 a14579a <=( (not A168)  and  A169 );
 a14580a <=( A170  and  a14579a );
 a14584a <=( A265  and  A200 );
 a14585a <=( A199  and  a14584a );
 a14586a <=( a14585a  and  a14580a );
 a14590a <=( A269  and  A267 );
 a14591a <=( (not A266)  and  a14590a );
 a14595a <=( (not A302)  and  (not A301) );
 a14596a <=( A298  and  a14595a );
 a14597a <=( a14596a  and  a14591a );
 a14601a <=( (not A168)  and  A169 );
 a14602a <=( A170  and  a14601a );
 a14606a <=( (not A266)  and  A200 );
 a14607a <=( (not A199)  and  a14606a );
 a14608a <=( a14607a  and  a14602a );
 a14612a <=( A298  and  (not A269) );
 a14613a <=( (not A268)  and  a14612a );
 a14617a <=( A301  and  A300 );
 a14618a <=( (not A299)  and  a14617a );
 a14619a <=( a14618a  and  a14613a );
 a14623a <=( (not A168)  and  A169 );
 a14624a <=( A170  and  a14623a );
 a14628a <=( (not A266)  and  A200 );
 a14629a <=( (not A199)  and  a14628a );
 a14630a <=( a14629a  and  a14624a );
 a14634a <=( A298  and  (not A269) );
 a14635a <=( (not A268)  and  a14634a );
 a14639a <=( A302  and  A300 );
 a14640a <=( (not A299)  and  a14639a );
 a14641a <=( a14640a  and  a14635a );
 a14645a <=( (not A168)  and  A169 );
 a14646a <=( A170  and  a14645a );
 a14650a <=( (not A203)  and  (not A202) );
 a14651a <=( (not A200)  and  a14650a );
 a14652a <=( a14651a  and  a14646a );
 a14656a <=( A267  and  (not A266) );
 a14657a <=( A265  and  a14656a );
 a14661a <=( (not A300)  and  A298 );
 a14662a <=( A268  and  a14661a );
 a14663a <=( a14662a  and  a14657a );
 a14667a <=( (not A168)  and  A169 );
 a14668a <=( A170  and  a14667a );
 a14672a <=( (not A203)  and  (not A202) );
 a14673a <=( (not A200)  and  a14672a );
 a14674a <=( a14673a  and  a14668a );
 a14678a <=( A267  and  (not A266) );
 a14679a <=( A265  and  a14678a );
 a14683a <=( A299  and  A298 );
 a14684a <=( A268  and  a14683a );
 a14685a <=( a14684a  and  a14679a );
 a14689a <=( (not A168)  and  A169 );
 a14690a <=( A170  and  a14689a );
 a14694a <=( (not A203)  and  (not A202) );
 a14695a <=( (not A200)  and  a14694a );
 a14696a <=( a14695a  and  a14690a );
 a14700a <=( A267  and  (not A266) );
 a14701a <=( A265  and  a14700a );
 a14705a <=( (not A299)  and  (not A298) );
 a14706a <=( A268  and  a14705a );
 a14707a <=( a14706a  and  a14701a );
 a14711a <=( (not A168)  and  A169 );
 a14712a <=( A170  and  a14711a );
 a14716a <=( (not A203)  and  (not A202) );
 a14717a <=( (not A200)  and  a14716a );
 a14718a <=( a14717a  and  a14712a );
 a14722a <=( A267  and  (not A266) );
 a14723a <=( A265  and  a14722a );
 a14727a <=( (not A300)  and  A298 );
 a14728a <=( A269  and  a14727a );
 a14729a <=( a14728a  and  a14723a );
 a14733a <=( (not A168)  and  A169 );
 a14734a <=( A170  and  a14733a );
 a14738a <=( (not A203)  and  (not A202) );
 a14739a <=( (not A200)  and  a14738a );
 a14740a <=( a14739a  and  a14734a );
 a14744a <=( A267  and  (not A266) );
 a14745a <=( A265  and  a14744a );
 a14749a <=( A299  and  A298 );
 a14750a <=( A269  and  a14749a );
 a14751a <=( a14750a  and  a14745a );
 a14755a <=( (not A168)  and  A169 );
 a14756a <=( A170  and  a14755a );
 a14760a <=( (not A203)  and  (not A202) );
 a14761a <=( (not A200)  and  a14760a );
 a14762a <=( a14761a  and  a14756a );
 a14766a <=( A267  and  (not A266) );
 a14767a <=( A265  and  a14766a );
 a14771a <=( (not A299)  and  (not A298) );
 a14772a <=( A269  and  a14771a );
 a14773a <=( a14772a  and  a14767a );
 a14777a <=( (not A168)  and  A169 );
 a14778a <=( A170  and  a14777a );
 a14782a <=( A265  and  (not A201) );
 a14783a <=( (not A200)  and  a14782a );
 a14784a <=( a14783a  and  a14778a );
 a14788a <=( A268  and  A267 );
 a14789a <=( (not A266)  and  a14788a );
 a14793a <=( (not A302)  and  (not A301) );
 a14794a <=( A298  and  a14793a );
 a14795a <=( a14794a  and  a14789a );
 a14799a <=( (not A168)  and  A169 );
 a14800a <=( A170  and  a14799a );
 a14804a <=( A265  and  (not A201) );
 a14805a <=( (not A200)  and  a14804a );
 a14806a <=( a14805a  and  a14800a );
 a14810a <=( A269  and  A267 );
 a14811a <=( (not A266)  and  a14810a );
 a14815a <=( (not A302)  and  (not A301) );
 a14816a <=( A298  and  a14815a );
 a14817a <=( a14816a  and  a14811a );
 a14821a <=( (not A168)  and  A169 );
 a14822a <=( A170  and  a14821a );
 a14826a <=( A201  and  (not A200) );
 a14827a <=( A199  and  a14826a );
 a14828a <=( a14827a  and  a14822a );
 a14832a <=( (not A268)  and  (not A266) );
 a14833a <=( A202  and  a14832a );
 a14837a <=( A299  and  (not A298) );
 a14838a <=( (not A269)  and  a14837a );
 a14839a <=( a14838a  and  a14833a );
 a14843a <=( (not A168)  and  A169 );
 a14844a <=( A170  and  a14843a );
 a14848a <=( A201  and  (not A200) );
 a14849a <=( A199  and  a14848a );
 a14850a <=( a14849a  and  a14844a );
 a14854a <=( (not A268)  and  (not A266) );
 a14855a <=( A203  and  a14854a );
 a14859a <=( A299  and  (not A298) );
 a14860a <=( (not A269)  and  a14859a );
 a14861a <=( a14860a  and  a14855a );
 a14865a <=( (not A168)  and  A169 );
 a14866a <=( A170  and  a14865a );
 a14870a <=( A265  and  (not A200) );
 a14871a <=( (not A199)  and  a14870a );
 a14872a <=( a14871a  and  a14866a );
 a14876a <=( A268  and  A267 );
 a14877a <=( (not A266)  and  a14876a );
 a14881a <=( (not A302)  and  (not A301) );
 a14882a <=( A298  and  a14881a );
 a14883a <=( a14882a  and  a14877a );
 a14887a <=( (not A168)  and  A169 );
 a14888a <=( A170  and  a14887a );
 a14892a <=( A265  and  (not A200) );
 a14893a <=( (not A199)  and  a14892a );
 a14894a <=( a14893a  and  a14888a );
 a14898a <=( A269  and  A267 );
 a14899a <=( (not A266)  and  a14898a );
 a14903a <=( (not A302)  and  (not A301) );
 a14904a <=( A298  and  a14903a );
 a14905a <=( a14904a  and  a14899a );
 a14909a <=( A167  and  A169 );
 a14910a <=( (not A170)  and  a14909a );
 a14914a <=( A200  and  A199 );
 a14915a <=( A166  and  a14914a );
 a14916a <=( a14915a  and  a14910a );
 a14920a <=( A298  and  A266 );
 a14921a <=( A265  and  a14920a );
 a14925a <=( A301  and  A300 );
 a14926a <=( (not A299)  and  a14925a );
 a14927a <=( a14926a  and  a14921a );
 a14931a <=( A167  and  A169 );
 a14932a <=( (not A170)  and  a14931a );
 a14936a <=( A200  and  A199 );
 a14937a <=( A166  and  a14936a );
 a14938a <=( a14937a  and  a14932a );
 a14942a <=( A298  and  A266 );
 a14943a <=( A265  and  a14942a );
 a14947a <=( A302  and  A300 );
 a14948a <=( (not A299)  and  a14947a );
 a14949a <=( a14948a  and  a14943a );
 a14953a <=( A167  and  A169 );
 a14954a <=( (not A170)  and  a14953a );
 a14958a <=( A200  and  A199 );
 a14959a <=( A166  and  a14958a );
 a14960a <=( a14959a  and  a14954a );
 a14964a <=( A298  and  (not A267) );
 a14965a <=( (not A266)  and  a14964a );
 a14969a <=( A301  and  A300 );
 a14970a <=( (not A299)  and  a14969a );
 a14971a <=( a14970a  and  a14965a );
 a14975a <=( A167  and  A169 );
 a14976a <=( (not A170)  and  a14975a );
 a14980a <=( A200  and  A199 );
 a14981a <=( A166  and  a14980a );
 a14982a <=( a14981a  and  a14976a );
 a14986a <=( A298  and  (not A267) );
 a14987a <=( (not A266)  and  a14986a );
 a14991a <=( A302  and  A300 );
 a14992a <=( (not A299)  and  a14991a );
 a14993a <=( a14992a  and  a14987a );
 a14997a <=( A167  and  A169 );
 a14998a <=( (not A170)  and  a14997a );
 a15002a <=( A200  and  A199 );
 a15003a <=( A166  and  a15002a );
 a15004a <=( a15003a  and  a14998a );
 a15008a <=( A298  and  (not A266) );
 a15009a <=( (not A265)  and  a15008a );
 a15013a <=( A301  and  A300 );
 a15014a <=( (not A299)  and  a15013a );
 a15015a <=( a15014a  and  a15009a );
 a15019a <=( A167  and  A169 );
 a15020a <=( (not A170)  and  a15019a );
 a15024a <=( A200  and  A199 );
 a15025a <=( A166  and  a15024a );
 a15026a <=( a15025a  and  a15020a );
 a15030a <=( A298  and  (not A266) );
 a15031a <=( (not A265)  and  a15030a );
 a15035a <=( A302  and  A300 );
 a15036a <=( (not A299)  and  a15035a );
 a15037a <=( a15036a  and  a15031a );
 a15041a <=( A167  and  A169 );
 a15042a <=( (not A170)  and  a15041a );
 a15046a <=( A200  and  (not A199) );
 a15047a <=( A166  and  a15046a );
 a15048a <=( a15047a  and  a15042a );
 a15052a <=( A267  and  (not A266) );
 a15053a <=( A265  and  a15052a );
 a15057a <=( (not A300)  and  A298 );
 a15058a <=( A268  and  a15057a );
 a15059a <=( a15058a  and  a15053a );
 a15063a <=( A167  and  A169 );
 a15064a <=( (not A170)  and  a15063a );
 a15068a <=( A200  and  (not A199) );
 a15069a <=( A166  and  a15068a );
 a15070a <=( a15069a  and  a15064a );
 a15074a <=( A267  and  (not A266) );
 a15075a <=( A265  and  a15074a );
 a15079a <=( A299  and  A298 );
 a15080a <=( A268  and  a15079a );
 a15081a <=( a15080a  and  a15075a );
 a15085a <=( A167  and  A169 );
 a15086a <=( (not A170)  and  a15085a );
 a15090a <=( A200  and  (not A199) );
 a15091a <=( A166  and  a15090a );
 a15092a <=( a15091a  and  a15086a );
 a15096a <=( A267  and  (not A266) );
 a15097a <=( A265  and  a15096a );
 a15101a <=( (not A299)  and  (not A298) );
 a15102a <=( A268  and  a15101a );
 a15103a <=( a15102a  and  a15097a );
 a15107a <=( A167  and  A169 );
 a15108a <=( (not A170)  and  a15107a );
 a15112a <=( A200  and  (not A199) );
 a15113a <=( A166  and  a15112a );
 a15114a <=( a15113a  and  a15108a );
 a15118a <=( A267  and  (not A266) );
 a15119a <=( A265  and  a15118a );
 a15123a <=( (not A300)  and  A298 );
 a15124a <=( A269  and  a15123a );
 a15125a <=( a15124a  and  a15119a );
 a15129a <=( A167  and  A169 );
 a15130a <=( (not A170)  and  a15129a );
 a15134a <=( A200  and  (not A199) );
 a15135a <=( A166  and  a15134a );
 a15136a <=( a15135a  and  a15130a );
 a15140a <=( A267  and  (not A266) );
 a15141a <=( A265  and  a15140a );
 a15145a <=( A299  and  A298 );
 a15146a <=( A269  and  a15145a );
 a15147a <=( a15146a  and  a15141a );
 a15151a <=( A167  and  A169 );
 a15152a <=( (not A170)  and  a15151a );
 a15156a <=( A200  and  (not A199) );
 a15157a <=( A166  and  a15156a );
 a15158a <=( a15157a  and  a15152a );
 a15162a <=( A267  and  (not A266) );
 a15163a <=( A265  and  a15162a );
 a15167a <=( (not A299)  and  (not A298) );
 a15168a <=( A269  and  a15167a );
 a15169a <=( a15168a  and  a15163a );
 a15173a <=( A167  and  A169 );
 a15174a <=( (not A170)  and  a15173a );
 a15178a <=( (not A202)  and  (not A200) );
 a15179a <=( A166  and  a15178a );
 a15180a <=( a15179a  and  a15174a );
 a15184a <=( (not A268)  and  (not A266) );
 a15185a <=( (not A203)  and  a15184a );
 a15189a <=( A299  and  (not A298) );
 a15190a <=( (not A269)  and  a15189a );
 a15191a <=( a15190a  and  a15185a );
 a15195a <=( A167  and  A169 );
 a15196a <=( (not A170)  and  a15195a );
 a15200a <=( (not A201)  and  (not A200) );
 a15201a <=( A166  and  a15200a );
 a15202a <=( a15201a  and  a15196a );
 a15206a <=( A298  and  A266 );
 a15207a <=( A265  and  a15206a );
 a15211a <=( A301  and  A300 );
 a15212a <=( (not A299)  and  a15211a );
 a15213a <=( a15212a  and  a15207a );
 a15217a <=( A167  and  A169 );
 a15218a <=( (not A170)  and  a15217a );
 a15222a <=( (not A201)  and  (not A200) );
 a15223a <=( A166  and  a15222a );
 a15224a <=( a15223a  and  a15218a );
 a15228a <=( A298  and  A266 );
 a15229a <=( A265  and  a15228a );
 a15233a <=( A302  and  A300 );
 a15234a <=( (not A299)  and  a15233a );
 a15235a <=( a15234a  and  a15229a );
 a15239a <=( A167  and  A169 );
 a15240a <=( (not A170)  and  a15239a );
 a15244a <=( (not A201)  and  (not A200) );
 a15245a <=( A166  and  a15244a );
 a15246a <=( a15245a  and  a15240a );
 a15250a <=( A298  and  (not A267) );
 a15251a <=( (not A266)  and  a15250a );
 a15255a <=( A301  and  A300 );
 a15256a <=( (not A299)  and  a15255a );
 a15257a <=( a15256a  and  a15251a );
 a15261a <=( A167  and  A169 );
 a15262a <=( (not A170)  and  a15261a );
 a15266a <=( (not A201)  and  (not A200) );
 a15267a <=( A166  and  a15266a );
 a15268a <=( a15267a  and  a15262a );
 a15272a <=( A298  and  (not A267) );
 a15273a <=( (not A266)  and  a15272a );
 a15277a <=( A302  and  A300 );
 a15278a <=( (not A299)  and  a15277a );
 a15279a <=( a15278a  and  a15273a );
 a15283a <=( A167  and  A169 );
 a15284a <=( (not A170)  and  a15283a );
 a15288a <=( (not A201)  and  (not A200) );
 a15289a <=( A166  and  a15288a );
 a15290a <=( a15289a  and  a15284a );
 a15294a <=( A298  and  (not A266) );
 a15295a <=( (not A265)  and  a15294a );
 a15299a <=( A301  and  A300 );
 a15300a <=( (not A299)  and  a15299a );
 a15301a <=( a15300a  and  a15295a );
 a15305a <=( A167  and  A169 );
 a15306a <=( (not A170)  and  a15305a );
 a15310a <=( (not A201)  and  (not A200) );
 a15311a <=( A166  and  a15310a );
 a15312a <=( a15311a  and  a15306a );
 a15316a <=( A298  and  (not A266) );
 a15317a <=( (not A265)  and  a15316a );
 a15321a <=( A302  and  A300 );
 a15322a <=( (not A299)  and  a15321a );
 a15323a <=( a15322a  and  a15317a );
 a15327a <=( A167  and  A169 );
 a15328a <=( (not A170)  and  a15327a );
 a15332a <=( (not A200)  and  A199 );
 a15333a <=( A166  and  a15332a );
 a15334a <=( a15333a  and  a15328a );
 a15338a <=( (not A265)  and  A202 );
 a15339a <=( A201  and  a15338a );
 a15343a <=( (not A300)  and  A298 );
 a15344a <=( A266  and  a15343a );
 a15345a <=( a15344a  and  a15339a );
 a15349a <=( A167  and  A169 );
 a15350a <=( (not A170)  and  a15349a );
 a15354a <=( (not A200)  and  A199 );
 a15355a <=( A166  and  a15354a );
 a15356a <=( a15355a  and  a15350a );
 a15360a <=( (not A265)  and  A202 );
 a15361a <=( A201  and  a15360a );
 a15365a <=( A299  and  A298 );
 a15366a <=( A266  and  a15365a );
 a15367a <=( a15366a  and  a15361a );
 a15371a <=( A167  and  A169 );
 a15372a <=( (not A170)  and  a15371a );
 a15376a <=( (not A200)  and  A199 );
 a15377a <=( A166  and  a15376a );
 a15378a <=( a15377a  and  a15372a );
 a15382a <=( (not A265)  and  A202 );
 a15383a <=( A201  and  a15382a );
 a15387a <=( (not A299)  and  (not A298) );
 a15388a <=( A266  and  a15387a );
 a15389a <=( a15388a  and  a15383a );
 a15393a <=( A167  and  A169 );
 a15394a <=( (not A170)  and  a15393a );
 a15398a <=( (not A200)  and  A199 );
 a15399a <=( A166  and  a15398a );
 a15400a <=( a15399a  and  a15394a );
 a15404a <=( (not A265)  and  A203 );
 a15405a <=( A201  and  a15404a );
 a15409a <=( (not A300)  and  A298 );
 a15410a <=( A266  and  a15409a );
 a15411a <=( a15410a  and  a15405a );
 a15415a <=( A167  and  A169 );
 a15416a <=( (not A170)  and  a15415a );
 a15420a <=( (not A200)  and  A199 );
 a15421a <=( A166  and  a15420a );
 a15422a <=( a15421a  and  a15416a );
 a15426a <=( (not A265)  and  A203 );
 a15427a <=( A201  and  a15426a );
 a15431a <=( A299  and  A298 );
 a15432a <=( A266  and  a15431a );
 a15433a <=( a15432a  and  a15427a );
 a15437a <=( A167  and  A169 );
 a15438a <=( (not A170)  and  a15437a );
 a15442a <=( (not A200)  and  A199 );
 a15443a <=( A166  and  a15442a );
 a15444a <=( a15443a  and  a15438a );
 a15448a <=( (not A265)  and  A203 );
 a15449a <=( A201  and  a15448a );
 a15453a <=( (not A299)  and  (not A298) );
 a15454a <=( A266  and  a15453a );
 a15455a <=( a15454a  and  a15449a );
 a15459a <=( A167  and  A169 );
 a15460a <=( (not A170)  and  a15459a );
 a15464a <=( (not A200)  and  (not A199) );
 a15465a <=( A166  and  a15464a );
 a15466a <=( a15465a  and  a15460a );
 a15470a <=( A298  and  A266 );
 a15471a <=( A265  and  a15470a );
 a15475a <=( A301  and  A300 );
 a15476a <=( (not A299)  and  a15475a );
 a15477a <=( a15476a  and  a15471a );
 a15481a <=( A167  and  A169 );
 a15482a <=( (not A170)  and  a15481a );
 a15486a <=( (not A200)  and  (not A199) );
 a15487a <=( A166  and  a15486a );
 a15488a <=( a15487a  and  a15482a );
 a15492a <=( A298  and  A266 );
 a15493a <=( A265  and  a15492a );
 a15497a <=( A302  and  A300 );
 a15498a <=( (not A299)  and  a15497a );
 a15499a <=( a15498a  and  a15493a );
 a15503a <=( A167  and  A169 );
 a15504a <=( (not A170)  and  a15503a );
 a15508a <=( (not A200)  and  (not A199) );
 a15509a <=( A166  and  a15508a );
 a15510a <=( a15509a  and  a15504a );
 a15514a <=( A298  and  (not A267) );
 a15515a <=( (not A266)  and  a15514a );
 a15519a <=( A301  and  A300 );
 a15520a <=( (not A299)  and  a15519a );
 a15521a <=( a15520a  and  a15515a );
 a15525a <=( A167  and  A169 );
 a15526a <=( (not A170)  and  a15525a );
 a15530a <=( (not A200)  and  (not A199) );
 a15531a <=( A166  and  a15530a );
 a15532a <=( a15531a  and  a15526a );
 a15536a <=( A298  and  (not A267) );
 a15537a <=( (not A266)  and  a15536a );
 a15541a <=( A302  and  A300 );
 a15542a <=( (not A299)  and  a15541a );
 a15543a <=( a15542a  and  a15537a );
 a15547a <=( A167  and  A169 );
 a15548a <=( (not A170)  and  a15547a );
 a15552a <=( (not A200)  and  (not A199) );
 a15553a <=( A166  and  a15552a );
 a15554a <=( a15553a  and  a15548a );
 a15558a <=( A298  and  (not A266) );
 a15559a <=( (not A265)  and  a15558a );
 a15563a <=( A301  and  A300 );
 a15564a <=( (not A299)  and  a15563a );
 a15565a <=( a15564a  and  a15559a );
 a15569a <=( A167  and  A169 );
 a15570a <=( (not A170)  and  a15569a );
 a15574a <=( (not A200)  and  (not A199) );
 a15575a <=( A166  and  a15574a );
 a15576a <=( a15575a  and  a15570a );
 a15580a <=( A298  and  (not A266) );
 a15581a <=( (not A265)  and  a15580a );
 a15585a <=( A302  and  A300 );
 a15586a <=( (not A299)  and  a15585a );
 a15587a <=( a15586a  and  a15581a );
 a15591a <=( (not A167)  and  A169 );
 a15592a <=( (not A170)  and  a15591a );
 a15596a <=( A200  and  A199 );
 a15597a <=( (not A166)  and  a15596a );
 a15598a <=( a15597a  and  a15592a );
 a15602a <=( A298  and  A266 );
 a15603a <=( A265  and  a15602a );
 a15607a <=( A301  and  A300 );
 a15608a <=( (not A299)  and  a15607a );
 a15609a <=( a15608a  and  a15603a );
 a15613a <=( (not A167)  and  A169 );
 a15614a <=( (not A170)  and  a15613a );
 a15618a <=( A200  and  A199 );
 a15619a <=( (not A166)  and  a15618a );
 a15620a <=( a15619a  and  a15614a );
 a15624a <=( A298  and  A266 );
 a15625a <=( A265  and  a15624a );
 a15629a <=( A302  and  A300 );
 a15630a <=( (not A299)  and  a15629a );
 a15631a <=( a15630a  and  a15625a );
 a15635a <=( (not A167)  and  A169 );
 a15636a <=( (not A170)  and  a15635a );
 a15640a <=( A200  and  A199 );
 a15641a <=( (not A166)  and  a15640a );
 a15642a <=( a15641a  and  a15636a );
 a15646a <=( A298  and  (not A267) );
 a15647a <=( (not A266)  and  a15646a );
 a15651a <=( A301  and  A300 );
 a15652a <=( (not A299)  and  a15651a );
 a15653a <=( a15652a  and  a15647a );
 a15657a <=( (not A167)  and  A169 );
 a15658a <=( (not A170)  and  a15657a );
 a15662a <=( A200  and  A199 );
 a15663a <=( (not A166)  and  a15662a );
 a15664a <=( a15663a  and  a15658a );
 a15668a <=( A298  and  (not A267) );
 a15669a <=( (not A266)  and  a15668a );
 a15673a <=( A302  and  A300 );
 a15674a <=( (not A299)  and  a15673a );
 a15675a <=( a15674a  and  a15669a );
 a15679a <=( (not A167)  and  A169 );
 a15680a <=( (not A170)  and  a15679a );
 a15684a <=( A200  and  A199 );
 a15685a <=( (not A166)  and  a15684a );
 a15686a <=( a15685a  and  a15680a );
 a15690a <=( A298  and  (not A266) );
 a15691a <=( (not A265)  and  a15690a );
 a15695a <=( A301  and  A300 );
 a15696a <=( (not A299)  and  a15695a );
 a15697a <=( a15696a  and  a15691a );
 a15701a <=( (not A167)  and  A169 );
 a15702a <=( (not A170)  and  a15701a );
 a15706a <=( A200  and  A199 );
 a15707a <=( (not A166)  and  a15706a );
 a15708a <=( a15707a  and  a15702a );
 a15712a <=( A298  and  (not A266) );
 a15713a <=( (not A265)  and  a15712a );
 a15717a <=( A302  and  A300 );
 a15718a <=( (not A299)  and  a15717a );
 a15719a <=( a15718a  and  a15713a );
 a15723a <=( (not A167)  and  A169 );
 a15724a <=( (not A170)  and  a15723a );
 a15728a <=( A200  and  (not A199) );
 a15729a <=( (not A166)  and  a15728a );
 a15730a <=( a15729a  and  a15724a );
 a15734a <=( A267  and  (not A266) );
 a15735a <=( A265  and  a15734a );
 a15739a <=( (not A300)  and  A298 );
 a15740a <=( A268  and  a15739a );
 a15741a <=( a15740a  and  a15735a );
 a15745a <=( (not A167)  and  A169 );
 a15746a <=( (not A170)  and  a15745a );
 a15750a <=( A200  and  (not A199) );
 a15751a <=( (not A166)  and  a15750a );
 a15752a <=( a15751a  and  a15746a );
 a15756a <=( A267  and  (not A266) );
 a15757a <=( A265  and  a15756a );
 a15761a <=( A299  and  A298 );
 a15762a <=( A268  and  a15761a );
 a15763a <=( a15762a  and  a15757a );
 a15767a <=( (not A167)  and  A169 );
 a15768a <=( (not A170)  and  a15767a );
 a15772a <=( A200  and  (not A199) );
 a15773a <=( (not A166)  and  a15772a );
 a15774a <=( a15773a  and  a15768a );
 a15778a <=( A267  and  (not A266) );
 a15779a <=( A265  and  a15778a );
 a15783a <=( (not A299)  and  (not A298) );
 a15784a <=( A268  and  a15783a );
 a15785a <=( a15784a  and  a15779a );
 a15789a <=( (not A167)  and  A169 );
 a15790a <=( (not A170)  and  a15789a );
 a15794a <=( A200  and  (not A199) );
 a15795a <=( (not A166)  and  a15794a );
 a15796a <=( a15795a  and  a15790a );
 a15800a <=( A267  and  (not A266) );
 a15801a <=( A265  and  a15800a );
 a15805a <=( (not A300)  and  A298 );
 a15806a <=( A269  and  a15805a );
 a15807a <=( a15806a  and  a15801a );
 a15811a <=( (not A167)  and  A169 );
 a15812a <=( (not A170)  and  a15811a );
 a15816a <=( A200  and  (not A199) );
 a15817a <=( (not A166)  and  a15816a );
 a15818a <=( a15817a  and  a15812a );
 a15822a <=( A267  and  (not A266) );
 a15823a <=( A265  and  a15822a );
 a15827a <=( A299  and  A298 );
 a15828a <=( A269  and  a15827a );
 a15829a <=( a15828a  and  a15823a );
 a15833a <=( (not A167)  and  A169 );
 a15834a <=( (not A170)  and  a15833a );
 a15838a <=( A200  and  (not A199) );
 a15839a <=( (not A166)  and  a15838a );
 a15840a <=( a15839a  and  a15834a );
 a15844a <=( A267  and  (not A266) );
 a15845a <=( A265  and  a15844a );
 a15849a <=( (not A299)  and  (not A298) );
 a15850a <=( A269  and  a15849a );
 a15851a <=( a15850a  and  a15845a );
 a15855a <=( (not A167)  and  A169 );
 a15856a <=( (not A170)  and  a15855a );
 a15860a <=( (not A202)  and  (not A200) );
 a15861a <=( (not A166)  and  a15860a );
 a15862a <=( a15861a  and  a15856a );
 a15866a <=( (not A268)  and  (not A266) );
 a15867a <=( (not A203)  and  a15866a );
 a15871a <=( A299  and  (not A298) );
 a15872a <=( (not A269)  and  a15871a );
 a15873a <=( a15872a  and  a15867a );
 a15877a <=( (not A167)  and  A169 );
 a15878a <=( (not A170)  and  a15877a );
 a15882a <=( (not A201)  and  (not A200) );
 a15883a <=( (not A166)  and  a15882a );
 a15884a <=( a15883a  and  a15878a );
 a15888a <=( A298  and  A266 );
 a15889a <=( A265  and  a15888a );
 a15893a <=( A301  and  A300 );
 a15894a <=( (not A299)  and  a15893a );
 a15895a <=( a15894a  and  a15889a );
 a15899a <=( (not A167)  and  A169 );
 a15900a <=( (not A170)  and  a15899a );
 a15904a <=( (not A201)  and  (not A200) );
 a15905a <=( (not A166)  and  a15904a );
 a15906a <=( a15905a  and  a15900a );
 a15910a <=( A298  and  A266 );
 a15911a <=( A265  and  a15910a );
 a15915a <=( A302  and  A300 );
 a15916a <=( (not A299)  and  a15915a );
 a15917a <=( a15916a  and  a15911a );
 a15921a <=( (not A167)  and  A169 );
 a15922a <=( (not A170)  and  a15921a );
 a15926a <=( (not A201)  and  (not A200) );
 a15927a <=( (not A166)  and  a15926a );
 a15928a <=( a15927a  and  a15922a );
 a15932a <=( A298  and  (not A267) );
 a15933a <=( (not A266)  and  a15932a );
 a15937a <=( A301  and  A300 );
 a15938a <=( (not A299)  and  a15937a );
 a15939a <=( a15938a  and  a15933a );
 a15943a <=( (not A167)  and  A169 );
 a15944a <=( (not A170)  and  a15943a );
 a15948a <=( (not A201)  and  (not A200) );
 a15949a <=( (not A166)  and  a15948a );
 a15950a <=( a15949a  and  a15944a );
 a15954a <=( A298  and  (not A267) );
 a15955a <=( (not A266)  and  a15954a );
 a15959a <=( A302  and  A300 );
 a15960a <=( (not A299)  and  a15959a );
 a15961a <=( a15960a  and  a15955a );
 a15965a <=( (not A167)  and  A169 );
 a15966a <=( (not A170)  and  a15965a );
 a15970a <=( (not A201)  and  (not A200) );
 a15971a <=( (not A166)  and  a15970a );
 a15972a <=( a15971a  and  a15966a );
 a15976a <=( A298  and  (not A266) );
 a15977a <=( (not A265)  and  a15976a );
 a15981a <=( A301  and  A300 );
 a15982a <=( (not A299)  and  a15981a );
 a15983a <=( a15982a  and  a15977a );
 a15987a <=( (not A167)  and  A169 );
 a15988a <=( (not A170)  and  a15987a );
 a15992a <=( (not A201)  and  (not A200) );
 a15993a <=( (not A166)  and  a15992a );
 a15994a <=( a15993a  and  a15988a );
 a15998a <=( A298  and  (not A266) );
 a15999a <=( (not A265)  and  a15998a );
 a16003a <=( A302  and  A300 );
 a16004a <=( (not A299)  and  a16003a );
 a16005a <=( a16004a  and  a15999a );
 a16009a <=( (not A167)  and  A169 );
 a16010a <=( (not A170)  and  a16009a );
 a16014a <=( (not A200)  and  A199 );
 a16015a <=( (not A166)  and  a16014a );
 a16016a <=( a16015a  and  a16010a );
 a16020a <=( (not A265)  and  A202 );
 a16021a <=( A201  and  a16020a );
 a16025a <=( (not A300)  and  A298 );
 a16026a <=( A266  and  a16025a );
 a16027a <=( a16026a  and  a16021a );
 a16031a <=( (not A167)  and  A169 );
 a16032a <=( (not A170)  and  a16031a );
 a16036a <=( (not A200)  and  A199 );
 a16037a <=( (not A166)  and  a16036a );
 a16038a <=( a16037a  and  a16032a );
 a16042a <=( (not A265)  and  A202 );
 a16043a <=( A201  and  a16042a );
 a16047a <=( A299  and  A298 );
 a16048a <=( A266  and  a16047a );
 a16049a <=( a16048a  and  a16043a );
 a16053a <=( (not A167)  and  A169 );
 a16054a <=( (not A170)  and  a16053a );
 a16058a <=( (not A200)  and  A199 );
 a16059a <=( (not A166)  and  a16058a );
 a16060a <=( a16059a  and  a16054a );
 a16064a <=( (not A265)  and  A202 );
 a16065a <=( A201  and  a16064a );
 a16069a <=( (not A299)  and  (not A298) );
 a16070a <=( A266  and  a16069a );
 a16071a <=( a16070a  and  a16065a );
 a16075a <=( (not A167)  and  A169 );
 a16076a <=( (not A170)  and  a16075a );
 a16080a <=( (not A200)  and  A199 );
 a16081a <=( (not A166)  and  a16080a );
 a16082a <=( a16081a  and  a16076a );
 a16086a <=( (not A265)  and  A203 );
 a16087a <=( A201  and  a16086a );
 a16091a <=( (not A300)  and  A298 );
 a16092a <=( A266  and  a16091a );
 a16093a <=( a16092a  and  a16087a );
 a16097a <=( (not A167)  and  A169 );
 a16098a <=( (not A170)  and  a16097a );
 a16102a <=( (not A200)  and  A199 );
 a16103a <=( (not A166)  and  a16102a );
 a16104a <=( a16103a  and  a16098a );
 a16108a <=( (not A265)  and  A203 );
 a16109a <=( A201  and  a16108a );
 a16113a <=( A299  and  A298 );
 a16114a <=( A266  and  a16113a );
 a16115a <=( a16114a  and  a16109a );
 a16119a <=( (not A167)  and  A169 );
 a16120a <=( (not A170)  and  a16119a );
 a16124a <=( (not A200)  and  A199 );
 a16125a <=( (not A166)  and  a16124a );
 a16126a <=( a16125a  and  a16120a );
 a16130a <=( (not A265)  and  A203 );
 a16131a <=( A201  and  a16130a );
 a16135a <=( (not A299)  and  (not A298) );
 a16136a <=( A266  and  a16135a );
 a16137a <=( a16136a  and  a16131a );
 a16141a <=( (not A167)  and  A169 );
 a16142a <=( (not A170)  and  a16141a );
 a16146a <=( (not A200)  and  (not A199) );
 a16147a <=( (not A166)  and  a16146a );
 a16148a <=( a16147a  and  a16142a );
 a16152a <=( A298  and  A266 );
 a16153a <=( A265  and  a16152a );
 a16157a <=( A301  and  A300 );
 a16158a <=( (not A299)  and  a16157a );
 a16159a <=( a16158a  and  a16153a );
 a16163a <=( (not A167)  and  A169 );
 a16164a <=( (not A170)  and  a16163a );
 a16168a <=( (not A200)  and  (not A199) );
 a16169a <=( (not A166)  and  a16168a );
 a16170a <=( a16169a  and  a16164a );
 a16174a <=( A298  and  A266 );
 a16175a <=( A265  and  a16174a );
 a16179a <=( A302  and  A300 );
 a16180a <=( (not A299)  and  a16179a );
 a16181a <=( a16180a  and  a16175a );
 a16185a <=( (not A167)  and  A169 );
 a16186a <=( (not A170)  and  a16185a );
 a16190a <=( (not A200)  and  (not A199) );
 a16191a <=( (not A166)  and  a16190a );
 a16192a <=( a16191a  and  a16186a );
 a16196a <=( A298  and  (not A267) );
 a16197a <=( (not A266)  and  a16196a );
 a16201a <=( A301  and  A300 );
 a16202a <=( (not A299)  and  a16201a );
 a16203a <=( a16202a  and  a16197a );
 a16207a <=( (not A167)  and  A169 );
 a16208a <=( (not A170)  and  a16207a );
 a16212a <=( (not A200)  and  (not A199) );
 a16213a <=( (not A166)  and  a16212a );
 a16214a <=( a16213a  and  a16208a );
 a16218a <=( A298  and  (not A267) );
 a16219a <=( (not A266)  and  a16218a );
 a16223a <=( A302  and  A300 );
 a16224a <=( (not A299)  and  a16223a );
 a16225a <=( a16224a  and  a16219a );
 a16229a <=( (not A167)  and  A169 );
 a16230a <=( (not A170)  and  a16229a );
 a16234a <=( (not A200)  and  (not A199) );
 a16235a <=( (not A166)  and  a16234a );
 a16236a <=( a16235a  and  a16230a );
 a16240a <=( A298  and  (not A266) );
 a16241a <=( (not A265)  and  a16240a );
 a16245a <=( A301  and  A300 );
 a16246a <=( (not A299)  and  a16245a );
 a16247a <=( a16246a  and  a16241a );
 a16251a <=( (not A167)  and  A169 );
 a16252a <=( (not A170)  and  a16251a );
 a16256a <=( (not A200)  and  (not A199) );
 a16257a <=( (not A166)  and  a16256a );
 a16258a <=( a16257a  and  a16252a );
 a16262a <=( A298  and  (not A266) );
 a16263a <=( (not A265)  and  a16262a );
 a16267a <=( A302  and  A300 );
 a16268a <=( (not A299)  and  a16267a );
 a16269a <=( a16268a  and  a16263a );
 a16273a <=( (not A166)  and  (not A167) );
 a16274a <=( (not A169)  and  a16273a );
 a16278a <=( A265  and  A200 );
 a16279a <=( A199  and  a16278a );
 a16280a <=( a16279a  and  a16274a );
 a16284a <=( A268  and  A267 );
 a16285a <=( (not A266)  and  a16284a );
 a16289a <=( (not A302)  and  (not A301) );
 a16290a <=( A298  and  a16289a );
 a16291a <=( a16290a  and  a16285a );
 a16295a <=( (not A166)  and  (not A167) );
 a16296a <=( (not A169)  and  a16295a );
 a16300a <=( A265  and  A200 );
 a16301a <=( A199  and  a16300a );
 a16302a <=( a16301a  and  a16296a );
 a16306a <=( A269  and  A267 );
 a16307a <=( (not A266)  and  a16306a );
 a16311a <=( (not A302)  and  (not A301) );
 a16312a <=( A298  and  a16311a );
 a16313a <=( a16312a  and  a16307a );
 a16317a <=( (not A166)  and  (not A167) );
 a16318a <=( (not A169)  and  a16317a );
 a16322a <=( (not A266)  and  A200 );
 a16323a <=( (not A199)  and  a16322a );
 a16324a <=( a16323a  and  a16318a );
 a16328a <=( A298  and  (not A269) );
 a16329a <=( (not A268)  and  a16328a );
 a16333a <=( A301  and  A300 );
 a16334a <=( (not A299)  and  a16333a );
 a16335a <=( a16334a  and  a16329a );
 a16339a <=( (not A166)  and  (not A167) );
 a16340a <=( (not A169)  and  a16339a );
 a16344a <=( (not A266)  and  A200 );
 a16345a <=( (not A199)  and  a16344a );
 a16346a <=( a16345a  and  a16340a );
 a16350a <=( A298  and  (not A269) );
 a16351a <=( (not A268)  and  a16350a );
 a16355a <=( A302  and  A300 );
 a16356a <=( (not A299)  and  a16355a );
 a16357a <=( a16356a  and  a16351a );
 a16361a <=( (not A166)  and  (not A167) );
 a16362a <=( (not A169)  and  a16361a );
 a16366a <=( (not A203)  and  (not A202) );
 a16367a <=( (not A200)  and  a16366a );
 a16368a <=( a16367a  and  a16362a );
 a16372a <=( A267  and  (not A266) );
 a16373a <=( A265  and  a16372a );
 a16377a <=( (not A300)  and  A298 );
 a16378a <=( A268  and  a16377a );
 a16379a <=( a16378a  and  a16373a );
 a16383a <=( (not A166)  and  (not A167) );
 a16384a <=( (not A169)  and  a16383a );
 a16388a <=( (not A203)  and  (not A202) );
 a16389a <=( (not A200)  and  a16388a );
 a16390a <=( a16389a  and  a16384a );
 a16394a <=( A267  and  (not A266) );
 a16395a <=( A265  and  a16394a );
 a16399a <=( A299  and  A298 );
 a16400a <=( A268  and  a16399a );
 a16401a <=( a16400a  and  a16395a );
 a16405a <=( (not A166)  and  (not A167) );
 a16406a <=( (not A169)  and  a16405a );
 a16410a <=( (not A203)  and  (not A202) );
 a16411a <=( (not A200)  and  a16410a );
 a16412a <=( a16411a  and  a16406a );
 a16416a <=( A267  and  (not A266) );
 a16417a <=( A265  and  a16416a );
 a16421a <=( (not A299)  and  (not A298) );
 a16422a <=( A268  and  a16421a );
 a16423a <=( a16422a  and  a16417a );
 a16427a <=( (not A166)  and  (not A167) );
 a16428a <=( (not A169)  and  a16427a );
 a16432a <=( (not A203)  and  (not A202) );
 a16433a <=( (not A200)  and  a16432a );
 a16434a <=( a16433a  and  a16428a );
 a16438a <=( A267  and  (not A266) );
 a16439a <=( A265  and  a16438a );
 a16443a <=( (not A300)  and  A298 );
 a16444a <=( A269  and  a16443a );
 a16445a <=( a16444a  and  a16439a );
 a16449a <=( (not A166)  and  (not A167) );
 a16450a <=( (not A169)  and  a16449a );
 a16454a <=( (not A203)  and  (not A202) );
 a16455a <=( (not A200)  and  a16454a );
 a16456a <=( a16455a  and  a16450a );
 a16460a <=( A267  and  (not A266) );
 a16461a <=( A265  and  a16460a );
 a16465a <=( A299  and  A298 );
 a16466a <=( A269  and  a16465a );
 a16467a <=( a16466a  and  a16461a );
 a16471a <=( (not A166)  and  (not A167) );
 a16472a <=( (not A169)  and  a16471a );
 a16476a <=( (not A203)  and  (not A202) );
 a16477a <=( (not A200)  and  a16476a );
 a16478a <=( a16477a  and  a16472a );
 a16482a <=( A267  and  (not A266) );
 a16483a <=( A265  and  a16482a );
 a16487a <=( (not A299)  and  (not A298) );
 a16488a <=( A269  and  a16487a );
 a16489a <=( a16488a  and  a16483a );
 a16493a <=( (not A166)  and  (not A167) );
 a16494a <=( (not A169)  and  a16493a );
 a16498a <=( A265  and  (not A201) );
 a16499a <=( (not A200)  and  a16498a );
 a16500a <=( a16499a  and  a16494a );
 a16504a <=( A268  and  A267 );
 a16505a <=( (not A266)  and  a16504a );
 a16509a <=( (not A302)  and  (not A301) );
 a16510a <=( A298  and  a16509a );
 a16511a <=( a16510a  and  a16505a );
 a16515a <=( (not A166)  and  (not A167) );
 a16516a <=( (not A169)  and  a16515a );
 a16520a <=( A265  and  (not A201) );
 a16521a <=( (not A200)  and  a16520a );
 a16522a <=( a16521a  and  a16516a );
 a16526a <=( A269  and  A267 );
 a16527a <=( (not A266)  and  a16526a );
 a16531a <=( (not A302)  and  (not A301) );
 a16532a <=( A298  and  a16531a );
 a16533a <=( a16532a  and  a16527a );
 a16537a <=( (not A166)  and  (not A167) );
 a16538a <=( (not A169)  and  a16537a );
 a16542a <=( A201  and  (not A200) );
 a16543a <=( A199  and  a16542a );
 a16544a <=( a16543a  and  a16538a );
 a16548a <=( (not A268)  and  (not A266) );
 a16549a <=( A202  and  a16548a );
 a16553a <=( A299  and  (not A298) );
 a16554a <=( (not A269)  and  a16553a );
 a16555a <=( a16554a  and  a16549a );
 a16559a <=( (not A166)  and  (not A167) );
 a16560a <=( (not A169)  and  a16559a );
 a16564a <=( A201  and  (not A200) );
 a16565a <=( A199  and  a16564a );
 a16566a <=( a16565a  and  a16560a );
 a16570a <=( (not A268)  and  (not A266) );
 a16571a <=( A203  and  a16570a );
 a16575a <=( A299  and  (not A298) );
 a16576a <=( (not A269)  and  a16575a );
 a16577a <=( a16576a  and  a16571a );
 a16581a <=( (not A166)  and  (not A167) );
 a16582a <=( (not A169)  and  a16581a );
 a16586a <=( A265  and  (not A200) );
 a16587a <=( (not A199)  and  a16586a );
 a16588a <=( a16587a  and  a16582a );
 a16592a <=( A268  and  A267 );
 a16593a <=( (not A266)  and  a16592a );
 a16597a <=( (not A302)  and  (not A301) );
 a16598a <=( A298  and  a16597a );
 a16599a <=( a16598a  and  a16593a );
 a16603a <=( (not A166)  and  (not A167) );
 a16604a <=( (not A169)  and  a16603a );
 a16608a <=( A265  and  (not A200) );
 a16609a <=( (not A199)  and  a16608a );
 a16610a <=( a16609a  and  a16604a );
 a16614a <=( A269  and  A267 );
 a16615a <=( (not A266)  and  a16614a );
 a16619a <=( (not A302)  and  (not A301) );
 a16620a <=( A298  and  a16619a );
 a16621a <=( a16620a  and  a16615a );
 a16625a <=( A167  and  (not A168) );
 a16626a <=( (not A169)  and  a16625a );
 a16630a <=( A200  and  A199 );
 a16631a <=( A166  and  a16630a );
 a16632a <=( a16631a  and  a16626a );
 a16636a <=( A267  and  (not A266) );
 a16637a <=( A265  and  a16636a );
 a16641a <=( (not A300)  and  A298 );
 a16642a <=( A268  and  a16641a );
 a16643a <=( a16642a  and  a16637a );
 a16647a <=( A167  and  (not A168) );
 a16648a <=( (not A169)  and  a16647a );
 a16652a <=( A200  and  A199 );
 a16653a <=( A166  and  a16652a );
 a16654a <=( a16653a  and  a16648a );
 a16658a <=( A267  and  (not A266) );
 a16659a <=( A265  and  a16658a );
 a16663a <=( A299  and  A298 );
 a16664a <=( A268  and  a16663a );
 a16665a <=( a16664a  and  a16659a );
 a16669a <=( A167  and  (not A168) );
 a16670a <=( (not A169)  and  a16669a );
 a16674a <=( A200  and  A199 );
 a16675a <=( A166  and  a16674a );
 a16676a <=( a16675a  and  a16670a );
 a16680a <=( A267  and  (not A266) );
 a16681a <=( A265  and  a16680a );
 a16685a <=( (not A299)  and  (not A298) );
 a16686a <=( A268  and  a16685a );
 a16687a <=( a16686a  and  a16681a );
 a16691a <=( A167  and  (not A168) );
 a16692a <=( (not A169)  and  a16691a );
 a16696a <=( A200  and  A199 );
 a16697a <=( A166  and  a16696a );
 a16698a <=( a16697a  and  a16692a );
 a16702a <=( A267  and  (not A266) );
 a16703a <=( A265  and  a16702a );
 a16707a <=( (not A300)  and  A298 );
 a16708a <=( A269  and  a16707a );
 a16709a <=( a16708a  and  a16703a );
 a16713a <=( A167  and  (not A168) );
 a16714a <=( (not A169)  and  a16713a );
 a16718a <=( A200  and  A199 );
 a16719a <=( A166  and  a16718a );
 a16720a <=( a16719a  and  a16714a );
 a16724a <=( A267  and  (not A266) );
 a16725a <=( A265  and  a16724a );
 a16729a <=( A299  and  A298 );
 a16730a <=( A269  and  a16729a );
 a16731a <=( a16730a  and  a16725a );
 a16735a <=( A167  and  (not A168) );
 a16736a <=( (not A169)  and  a16735a );
 a16740a <=( A200  and  A199 );
 a16741a <=( A166  and  a16740a );
 a16742a <=( a16741a  and  a16736a );
 a16746a <=( A267  and  (not A266) );
 a16747a <=( A265  and  a16746a );
 a16751a <=( (not A299)  and  (not A298) );
 a16752a <=( A269  and  a16751a );
 a16753a <=( a16752a  and  a16747a );
 a16757a <=( A167  and  (not A168) );
 a16758a <=( (not A169)  and  a16757a );
 a16762a <=( A200  and  (not A199) );
 a16763a <=( A166  and  a16762a );
 a16764a <=( a16763a  and  a16758a );
 a16768a <=( A298  and  A266 );
 a16769a <=( A265  and  a16768a );
 a16773a <=( A301  and  A300 );
 a16774a <=( (not A299)  and  a16773a );
 a16775a <=( a16774a  and  a16769a );
 a16779a <=( A167  and  (not A168) );
 a16780a <=( (not A169)  and  a16779a );
 a16784a <=( A200  and  (not A199) );
 a16785a <=( A166  and  a16784a );
 a16786a <=( a16785a  and  a16780a );
 a16790a <=( A298  and  A266 );
 a16791a <=( A265  and  a16790a );
 a16795a <=( A302  and  A300 );
 a16796a <=( (not A299)  and  a16795a );
 a16797a <=( a16796a  and  a16791a );
 a16801a <=( A167  and  (not A168) );
 a16802a <=( (not A169)  and  a16801a );
 a16806a <=( A200  and  (not A199) );
 a16807a <=( A166  and  a16806a );
 a16808a <=( a16807a  and  a16802a );
 a16812a <=( A298  and  (not A267) );
 a16813a <=( (not A266)  and  a16812a );
 a16817a <=( A301  and  A300 );
 a16818a <=( (not A299)  and  a16817a );
 a16819a <=( a16818a  and  a16813a );
 a16823a <=( A167  and  (not A168) );
 a16824a <=( (not A169)  and  a16823a );
 a16828a <=( A200  and  (not A199) );
 a16829a <=( A166  and  a16828a );
 a16830a <=( a16829a  and  a16824a );
 a16834a <=( A298  and  (not A267) );
 a16835a <=( (not A266)  and  a16834a );
 a16839a <=( A302  and  A300 );
 a16840a <=( (not A299)  and  a16839a );
 a16841a <=( a16840a  and  a16835a );
 a16845a <=( A167  and  (not A168) );
 a16846a <=( (not A169)  and  a16845a );
 a16850a <=( A200  and  (not A199) );
 a16851a <=( A166  and  a16850a );
 a16852a <=( a16851a  and  a16846a );
 a16856a <=( A298  and  (not A266) );
 a16857a <=( (not A265)  and  a16856a );
 a16861a <=( A301  and  A300 );
 a16862a <=( (not A299)  and  a16861a );
 a16863a <=( a16862a  and  a16857a );
 a16867a <=( A167  and  (not A168) );
 a16868a <=( (not A169)  and  a16867a );
 a16872a <=( A200  and  (not A199) );
 a16873a <=( A166  and  a16872a );
 a16874a <=( a16873a  and  a16868a );
 a16878a <=( A298  and  (not A266) );
 a16879a <=( (not A265)  and  a16878a );
 a16883a <=( A302  and  A300 );
 a16884a <=( (not A299)  and  a16883a );
 a16885a <=( a16884a  and  a16879a );
 a16889a <=( A167  and  (not A168) );
 a16890a <=( (not A169)  and  a16889a );
 a16894a <=( (not A202)  and  (not A200) );
 a16895a <=( A166  and  a16894a );
 a16896a <=( a16895a  and  a16890a );
 a16900a <=( A266  and  (not A265) );
 a16901a <=( (not A203)  and  a16900a );
 a16905a <=( (not A302)  and  (not A301) );
 a16906a <=( A298  and  a16905a );
 a16907a <=( a16906a  and  a16901a );
 a16911a <=( A167  and  (not A168) );
 a16912a <=( (not A169)  and  a16911a );
 a16916a <=( (not A201)  and  (not A200) );
 a16917a <=( A166  and  a16916a );
 a16918a <=( a16917a  and  a16912a );
 a16922a <=( A267  and  (not A266) );
 a16923a <=( A265  and  a16922a );
 a16927a <=( (not A300)  and  A298 );
 a16928a <=( A268  and  a16927a );
 a16929a <=( a16928a  and  a16923a );
 a16933a <=( A167  and  (not A168) );
 a16934a <=( (not A169)  and  a16933a );
 a16938a <=( (not A201)  and  (not A200) );
 a16939a <=( A166  and  a16938a );
 a16940a <=( a16939a  and  a16934a );
 a16944a <=( A267  and  (not A266) );
 a16945a <=( A265  and  a16944a );
 a16949a <=( A299  and  A298 );
 a16950a <=( A268  and  a16949a );
 a16951a <=( a16950a  and  a16945a );
 a16955a <=( A167  and  (not A168) );
 a16956a <=( (not A169)  and  a16955a );
 a16960a <=( (not A201)  and  (not A200) );
 a16961a <=( A166  and  a16960a );
 a16962a <=( a16961a  and  a16956a );
 a16966a <=( A267  and  (not A266) );
 a16967a <=( A265  and  a16966a );
 a16971a <=( (not A299)  and  (not A298) );
 a16972a <=( A268  and  a16971a );
 a16973a <=( a16972a  and  a16967a );
 a16977a <=( A167  and  (not A168) );
 a16978a <=( (not A169)  and  a16977a );
 a16982a <=( (not A201)  and  (not A200) );
 a16983a <=( A166  and  a16982a );
 a16984a <=( a16983a  and  a16978a );
 a16988a <=( A267  and  (not A266) );
 a16989a <=( A265  and  a16988a );
 a16993a <=( (not A300)  and  A298 );
 a16994a <=( A269  and  a16993a );
 a16995a <=( a16994a  and  a16989a );
 a16999a <=( A167  and  (not A168) );
 a17000a <=( (not A169)  and  a16999a );
 a17004a <=( (not A201)  and  (not A200) );
 a17005a <=( A166  and  a17004a );
 a17006a <=( a17005a  and  a17000a );
 a17010a <=( A267  and  (not A266) );
 a17011a <=( A265  and  a17010a );
 a17015a <=( A299  and  A298 );
 a17016a <=( A269  and  a17015a );
 a17017a <=( a17016a  and  a17011a );
 a17021a <=( A167  and  (not A168) );
 a17022a <=( (not A169)  and  a17021a );
 a17026a <=( (not A201)  and  (not A200) );
 a17027a <=( A166  and  a17026a );
 a17028a <=( a17027a  and  a17022a );
 a17032a <=( A267  and  (not A266) );
 a17033a <=( A265  and  a17032a );
 a17037a <=( (not A299)  and  (not A298) );
 a17038a <=( A269  and  a17037a );
 a17039a <=( a17038a  and  a17033a );
 a17043a <=( A167  and  (not A168) );
 a17044a <=( (not A169)  and  a17043a );
 a17048a <=( (not A200)  and  A199 );
 a17049a <=( A166  and  a17048a );
 a17050a <=( a17049a  and  a17044a );
 a17054a <=( A265  and  A202 );
 a17055a <=( A201  and  a17054a );
 a17059a <=( A299  and  (not A298) );
 a17060a <=( A266  and  a17059a );
 a17061a <=( a17060a  and  a17055a );
 a17065a <=( A167  and  (not A168) );
 a17066a <=( (not A169)  and  a17065a );
 a17070a <=( (not A200)  and  A199 );
 a17071a <=( A166  and  a17070a );
 a17072a <=( a17071a  and  a17066a );
 a17076a <=( (not A266)  and  A202 );
 a17077a <=( A201  and  a17076a );
 a17081a <=( A299  and  (not A298) );
 a17082a <=( (not A267)  and  a17081a );
 a17083a <=( a17082a  and  a17077a );
 a17087a <=( A167  and  (not A168) );
 a17088a <=( (not A169)  and  a17087a );
 a17092a <=( (not A200)  and  A199 );
 a17093a <=( A166  and  a17092a );
 a17094a <=( a17093a  and  a17088a );
 a17098a <=( (not A265)  and  A202 );
 a17099a <=( A201  and  a17098a );
 a17103a <=( A299  and  (not A298) );
 a17104a <=( (not A266)  and  a17103a );
 a17105a <=( a17104a  and  a17099a );
 a17109a <=( A167  and  (not A168) );
 a17110a <=( (not A169)  and  a17109a );
 a17114a <=( (not A200)  and  A199 );
 a17115a <=( A166  and  a17114a );
 a17116a <=( a17115a  and  a17110a );
 a17120a <=( A265  and  A203 );
 a17121a <=( A201  and  a17120a );
 a17125a <=( A299  and  (not A298) );
 a17126a <=( A266  and  a17125a );
 a17127a <=( a17126a  and  a17121a );
 a17131a <=( A167  and  (not A168) );
 a17132a <=( (not A169)  and  a17131a );
 a17136a <=( (not A200)  and  A199 );
 a17137a <=( A166  and  a17136a );
 a17138a <=( a17137a  and  a17132a );
 a17142a <=( (not A266)  and  A203 );
 a17143a <=( A201  and  a17142a );
 a17147a <=( A299  and  (not A298) );
 a17148a <=( (not A267)  and  a17147a );
 a17149a <=( a17148a  and  a17143a );
 a17153a <=( A167  and  (not A168) );
 a17154a <=( (not A169)  and  a17153a );
 a17158a <=( (not A200)  and  A199 );
 a17159a <=( A166  and  a17158a );
 a17160a <=( a17159a  and  a17154a );
 a17164a <=( (not A265)  and  A203 );
 a17165a <=( A201  and  a17164a );
 a17169a <=( A299  and  (not A298) );
 a17170a <=( (not A266)  and  a17169a );
 a17171a <=( a17170a  and  a17165a );
 a17175a <=( A167  and  (not A168) );
 a17176a <=( (not A169)  and  a17175a );
 a17180a <=( (not A200)  and  (not A199) );
 a17181a <=( A166  and  a17180a );
 a17182a <=( a17181a  and  a17176a );
 a17186a <=( A267  and  (not A266) );
 a17187a <=( A265  and  a17186a );
 a17191a <=( (not A300)  and  A298 );
 a17192a <=( A268  and  a17191a );
 a17193a <=( a17192a  and  a17187a );
 a17197a <=( A167  and  (not A168) );
 a17198a <=( (not A169)  and  a17197a );
 a17202a <=( (not A200)  and  (not A199) );
 a17203a <=( A166  and  a17202a );
 a17204a <=( a17203a  and  a17198a );
 a17208a <=( A267  and  (not A266) );
 a17209a <=( A265  and  a17208a );
 a17213a <=( A299  and  A298 );
 a17214a <=( A268  and  a17213a );
 a17215a <=( a17214a  and  a17209a );
 a17219a <=( A167  and  (not A168) );
 a17220a <=( (not A169)  and  a17219a );
 a17224a <=( (not A200)  and  (not A199) );
 a17225a <=( A166  and  a17224a );
 a17226a <=( a17225a  and  a17220a );
 a17230a <=( A267  and  (not A266) );
 a17231a <=( A265  and  a17230a );
 a17235a <=( (not A299)  and  (not A298) );
 a17236a <=( A268  and  a17235a );
 a17237a <=( a17236a  and  a17231a );
 a17241a <=( A167  and  (not A168) );
 a17242a <=( (not A169)  and  a17241a );
 a17246a <=( (not A200)  and  (not A199) );
 a17247a <=( A166  and  a17246a );
 a17248a <=( a17247a  and  a17242a );
 a17252a <=( A267  and  (not A266) );
 a17253a <=( A265  and  a17252a );
 a17257a <=( (not A300)  and  A298 );
 a17258a <=( A269  and  a17257a );
 a17259a <=( a17258a  and  a17253a );
 a17263a <=( A167  and  (not A168) );
 a17264a <=( (not A169)  and  a17263a );
 a17268a <=( (not A200)  and  (not A199) );
 a17269a <=( A166  and  a17268a );
 a17270a <=( a17269a  and  a17264a );
 a17274a <=( A267  and  (not A266) );
 a17275a <=( A265  and  a17274a );
 a17279a <=( A299  and  A298 );
 a17280a <=( A269  and  a17279a );
 a17281a <=( a17280a  and  a17275a );
 a17285a <=( A167  and  (not A168) );
 a17286a <=( (not A169)  and  a17285a );
 a17290a <=( (not A200)  and  (not A199) );
 a17291a <=( A166  and  a17290a );
 a17292a <=( a17291a  and  a17286a );
 a17296a <=( A267  and  (not A266) );
 a17297a <=( A265  and  a17296a );
 a17301a <=( (not A299)  and  (not A298) );
 a17302a <=( A269  and  a17301a );
 a17303a <=( a17302a  and  a17297a );
 a17307a <=( A167  and  (not A169) );
 a17308a <=( A170  and  a17307a );
 a17312a <=( A200  and  A199 );
 a17313a <=( (not A166)  and  a17312a );
 a17314a <=( a17313a  and  a17308a );
 a17318a <=( A298  and  A266 );
 a17319a <=( A265  and  a17318a );
 a17323a <=( A301  and  A300 );
 a17324a <=( (not A299)  and  a17323a );
 a17325a <=( a17324a  and  a17319a );
 a17329a <=( A167  and  (not A169) );
 a17330a <=( A170  and  a17329a );
 a17334a <=( A200  and  A199 );
 a17335a <=( (not A166)  and  a17334a );
 a17336a <=( a17335a  and  a17330a );
 a17340a <=( A298  and  A266 );
 a17341a <=( A265  and  a17340a );
 a17345a <=( A302  and  A300 );
 a17346a <=( (not A299)  and  a17345a );
 a17347a <=( a17346a  and  a17341a );
 a17351a <=( A167  and  (not A169) );
 a17352a <=( A170  and  a17351a );
 a17356a <=( A200  and  A199 );
 a17357a <=( (not A166)  and  a17356a );
 a17358a <=( a17357a  and  a17352a );
 a17362a <=( A298  and  (not A267) );
 a17363a <=( (not A266)  and  a17362a );
 a17367a <=( A301  and  A300 );
 a17368a <=( (not A299)  and  a17367a );
 a17369a <=( a17368a  and  a17363a );
 a17373a <=( A167  and  (not A169) );
 a17374a <=( A170  and  a17373a );
 a17378a <=( A200  and  A199 );
 a17379a <=( (not A166)  and  a17378a );
 a17380a <=( a17379a  and  a17374a );
 a17384a <=( A298  and  (not A267) );
 a17385a <=( (not A266)  and  a17384a );
 a17389a <=( A302  and  A300 );
 a17390a <=( (not A299)  and  a17389a );
 a17391a <=( a17390a  and  a17385a );
 a17395a <=( A167  and  (not A169) );
 a17396a <=( A170  and  a17395a );
 a17400a <=( A200  and  A199 );
 a17401a <=( (not A166)  and  a17400a );
 a17402a <=( a17401a  and  a17396a );
 a17406a <=( A298  and  (not A266) );
 a17407a <=( (not A265)  and  a17406a );
 a17411a <=( A301  and  A300 );
 a17412a <=( (not A299)  and  a17411a );
 a17413a <=( a17412a  and  a17407a );
 a17417a <=( A167  and  (not A169) );
 a17418a <=( A170  and  a17417a );
 a17422a <=( A200  and  A199 );
 a17423a <=( (not A166)  and  a17422a );
 a17424a <=( a17423a  and  a17418a );
 a17428a <=( A298  and  (not A266) );
 a17429a <=( (not A265)  and  a17428a );
 a17433a <=( A302  and  A300 );
 a17434a <=( (not A299)  and  a17433a );
 a17435a <=( a17434a  and  a17429a );
 a17439a <=( A167  and  (not A169) );
 a17440a <=( A170  and  a17439a );
 a17444a <=( A200  and  (not A199) );
 a17445a <=( (not A166)  and  a17444a );
 a17446a <=( a17445a  and  a17440a );
 a17450a <=( A267  and  (not A266) );
 a17451a <=( A265  and  a17450a );
 a17455a <=( (not A300)  and  A298 );
 a17456a <=( A268  and  a17455a );
 a17457a <=( a17456a  and  a17451a );
 a17461a <=( A167  and  (not A169) );
 a17462a <=( A170  and  a17461a );
 a17466a <=( A200  and  (not A199) );
 a17467a <=( (not A166)  and  a17466a );
 a17468a <=( a17467a  and  a17462a );
 a17472a <=( A267  and  (not A266) );
 a17473a <=( A265  and  a17472a );
 a17477a <=( A299  and  A298 );
 a17478a <=( A268  and  a17477a );
 a17479a <=( a17478a  and  a17473a );
 a17483a <=( A167  and  (not A169) );
 a17484a <=( A170  and  a17483a );
 a17488a <=( A200  and  (not A199) );
 a17489a <=( (not A166)  and  a17488a );
 a17490a <=( a17489a  and  a17484a );
 a17494a <=( A267  and  (not A266) );
 a17495a <=( A265  and  a17494a );
 a17499a <=( (not A299)  and  (not A298) );
 a17500a <=( A268  and  a17499a );
 a17501a <=( a17500a  and  a17495a );
 a17505a <=( A167  and  (not A169) );
 a17506a <=( A170  and  a17505a );
 a17510a <=( A200  and  (not A199) );
 a17511a <=( (not A166)  and  a17510a );
 a17512a <=( a17511a  and  a17506a );
 a17516a <=( A267  and  (not A266) );
 a17517a <=( A265  and  a17516a );
 a17521a <=( (not A300)  and  A298 );
 a17522a <=( A269  and  a17521a );
 a17523a <=( a17522a  and  a17517a );
 a17527a <=( A167  and  (not A169) );
 a17528a <=( A170  and  a17527a );
 a17532a <=( A200  and  (not A199) );
 a17533a <=( (not A166)  and  a17532a );
 a17534a <=( a17533a  and  a17528a );
 a17538a <=( A267  and  (not A266) );
 a17539a <=( A265  and  a17538a );
 a17543a <=( A299  and  A298 );
 a17544a <=( A269  and  a17543a );
 a17545a <=( a17544a  and  a17539a );
 a17549a <=( A167  and  (not A169) );
 a17550a <=( A170  and  a17549a );
 a17554a <=( A200  and  (not A199) );
 a17555a <=( (not A166)  and  a17554a );
 a17556a <=( a17555a  and  a17550a );
 a17560a <=( A267  and  (not A266) );
 a17561a <=( A265  and  a17560a );
 a17565a <=( (not A299)  and  (not A298) );
 a17566a <=( A269  and  a17565a );
 a17567a <=( a17566a  and  a17561a );
 a17571a <=( A167  and  (not A169) );
 a17572a <=( A170  and  a17571a );
 a17576a <=( (not A202)  and  (not A200) );
 a17577a <=( (not A166)  and  a17576a );
 a17578a <=( a17577a  and  a17572a );
 a17582a <=( (not A268)  and  (not A266) );
 a17583a <=( (not A203)  and  a17582a );
 a17587a <=( A299  and  (not A298) );
 a17588a <=( (not A269)  and  a17587a );
 a17589a <=( a17588a  and  a17583a );
 a17593a <=( A167  and  (not A169) );
 a17594a <=( A170  and  a17593a );
 a17598a <=( (not A201)  and  (not A200) );
 a17599a <=( (not A166)  and  a17598a );
 a17600a <=( a17599a  and  a17594a );
 a17604a <=( A298  and  A266 );
 a17605a <=( A265  and  a17604a );
 a17609a <=( A301  and  A300 );
 a17610a <=( (not A299)  and  a17609a );
 a17611a <=( a17610a  and  a17605a );
 a17615a <=( A167  and  (not A169) );
 a17616a <=( A170  and  a17615a );
 a17620a <=( (not A201)  and  (not A200) );
 a17621a <=( (not A166)  and  a17620a );
 a17622a <=( a17621a  and  a17616a );
 a17626a <=( A298  and  A266 );
 a17627a <=( A265  and  a17626a );
 a17631a <=( A302  and  A300 );
 a17632a <=( (not A299)  and  a17631a );
 a17633a <=( a17632a  and  a17627a );
 a17637a <=( A167  and  (not A169) );
 a17638a <=( A170  and  a17637a );
 a17642a <=( (not A201)  and  (not A200) );
 a17643a <=( (not A166)  and  a17642a );
 a17644a <=( a17643a  and  a17638a );
 a17648a <=( A298  and  (not A267) );
 a17649a <=( (not A266)  and  a17648a );
 a17653a <=( A301  and  A300 );
 a17654a <=( (not A299)  and  a17653a );
 a17655a <=( a17654a  and  a17649a );
 a17659a <=( A167  and  (not A169) );
 a17660a <=( A170  and  a17659a );
 a17664a <=( (not A201)  and  (not A200) );
 a17665a <=( (not A166)  and  a17664a );
 a17666a <=( a17665a  and  a17660a );
 a17670a <=( A298  and  (not A267) );
 a17671a <=( (not A266)  and  a17670a );
 a17675a <=( A302  and  A300 );
 a17676a <=( (not A299)  and  a17675a );
 a17677a <=( a17676a  and  a17671a );
 a17681a <=( A167  and  (not A169) );
 a17682a <=( A170  and  a17681a );
 a17686a <=( (not A201)  and  (not A200) );
 a17687a <=( (not A166)  and  a17686a );
 a17688a <=( a17687a  and  a17682a );
 a17692a <=( A298  and  (not A266) );
 a17693a <=( (not A265)  and  a17692a );
 a17697a <=( A301  and  A300 );
 a17698a <=( (not A299)  and  a17697a );
 a17699a <=( a17698a  and  a17693a );
 a17703a <=( A167  and  (not A169) );
 a17704a <=( A170  and  a17703a );
 a17708a <=( (not A201)  and  (not A200) );
 a17709a <=( (not A166)  and  a17708a );
 a17710a <=( a17709a  and  a17704a );
 a17714a <=( A298  and  (not A266) );
 a17715a <=( (not A265)  and  a17714a );
 a17719a <=( A302  and  A300 );
 a17720a <=( (not A299)  and  a17719a );
 a17721a <=( a17720a  and  a17715a );
 a17725a <=( A167  and  (not A169) );
 a17726a <=( A170  and  a17725a );
 a17730a <=( (not A200)  and  A199 );
 a17731a <=( (not A166)  and  a17730a );
 a17732a <=( a17731a  and  a17726a );
 a17736a <=( (not A265)  and  A202 );
 a17737a <=( A201  and  a17736a );
 a17741a <=( (not A300)  and  A298 );
 a17742a <=( A266  and  a17741a );
 a17743a <=( a17742a  and  a17737a );
 a17747a <=( A167  and  (not A169) );
 a17748a <=( A170  and  a17747a );
 a17752a <=( (not A200)  and  A199 );
 a17753a <=( (not A166)  and  a17752a );
 a17754a <=( a17753a  and  a17748a );
 a17758a <=( (not A265)  and  A202 );
 a17759a <=( A201  and  a17758a );
 a17763a <=( A299  and  A298 );
 a17764a <=( A266  and  a17763a );
 a17765a <=( a17764a  and  a17759a );
 a17769a <=( A167  and  (not A169) );
 a17770a <=( A170  and  a17769a );
 a17774a <=( (not A200)  and  A199 );
 a17775a <=( (not A166)  and  a17774a );
 a17776a <=( a17775a  and  a17770a );
 a17780a <=( (not A265)  and  A202 );
 a17781a <=( A201  and  a17780a );
 a17785a <=( (not A299)  and  (not A298) );
 a17786a <=( A266  and  a17785a );
 a17787a <=( a17786a  and  a17781a );
 a17791a <=( A167  and  (not A169) );
 a17792a <=( A170  and  a17791a );
 a17796a <=( (not A200)  and  A199 );
 a17797a <=( (not A166)  and  a17796a );
 a17798a <=( a17797a  and  a17792a );
 a17802a <=( (not A265)  and  A203 );
 a17803a <=( A201  and  a17802a );
 a17807a <=( (not A300)  and  A298 );
 a17808a <=( A266  and  a17807a );
 a17809a <=( a17808a  and  a17803a );
 a17813a <=( A167  and  (not A169) );
 a17814a <=( A170  and  a17813a );
 a17818a <=( (not A200)  and  A199 );
 a17819a <=( (not A166)  and  a17818a );
 a17820a <=( a17819a  and  a17814a );
 a17824a <=( (not A265)  and  A203 );
 a17825a <=( A201  and  a17824a );
 a17829a <=( A299  and  A298 );
 a17830a <=( A266  and  a17829a );
 a17831a <=( a17830a  and  a17825a );
 a17835a <=( A167  and  (not A169) );
 a17836a <=( A170  and  a17835a );
 a17840a <=( (not A200)  and  A199 );
 a17841a <=( (not A166)  and  a17840a );
 a17842a <=( a17841a  and  a17836a );
 a17846a <=( (not A265)  and  A203 );
 a17847a <=( A201  and  a17846a );
 a17851a <=( (not A299)  and  (not A298) );
 a17852a <=( A266  and  a17851a );
 a17853a <=( a17852a  and  a17847a );
 a17857a <=( A167  and  (not A169) );
 a17858a <=( A170  and  a17857a );
 a17862a <=( (not A200)  and  (not A199) );
 a17863a <=( (not A166)  and  a17862a );
 a17864a <=( a17863a  and  a17858a );
 a17868a <=( A298  and  A266 );
 a17869a <=( A265  and  a17868a );
 a17873a <=( A301  and  A300 );
 a17874a <=( (not A299)  and  a17873a );
 a17875a <=( a17874a  and  a17869a );
 a17879a <=( A167  and  (not A169) );
 a17880a <=( A170  and  a17879a );
 a17884a <=( (not A200)  and  (not A199) );
 a17885a <=( (not A166)  and  a17884a );
 a17886a <=( a17885a  and  a17880a );
 a17890a <=( A298  and  A266 );
 a17891a <=( A265  and  a17890a );
 a17895a <=( A302  and  A300 );
 a17896a <=( (not A299)  and  a17895a );
 a17897a <=( a17896a  and  a17891a );
 a17901a <=( A167  and  (not A169) );
 a17902a <=( A170  and  a17901a );
 a17906a <=( (not A200)  and  (not A199) );
 a17907a <=( (not A166)  and  a17906a );
 a17908a <=( a17907a  and  a17902a );
 a17912a <=( A298  and  (not A267) );
 a17913a <=( (not A266)  and  a17912a );
 a17917a <=( A301  and  A300 );
 a17918a <=( (not A299)  and  a17917a );
 a17919a <=( a17918a  and  a17913a );
 a17923a <=( A167  and  (not A169) );
 a17924a <=( A170  and  a17923a );
 a17928a <=( (not A200)  and  (not A199) );
 a17929a <=( (not A166)  and  a17928a );
 a17930a <=( a17929a  and  a17924a );
 a17934a <=( A298  and  (not A267) );
 a17935a <=( (not A266)  and  a17934a );
 a17939a <=( A302  and  A300 );
 a17940a <=( (not A299)  and  a17939a );
 a17941a <=( a17940a  and  a17935a );
 a17945a <=( A167  and  (not A169) );
 a17946a <=( A170  and  a17945a );
 a17950a <=( (not A200)  and  (not A199) );
 a17951a <=( (not A166)  and  a17950a );
 a17952a <=( a17951a  and  a17946a );
 a17956a <=( A298  and  (not A266) );
 a17957a <=( (not A265)  and  a17956a );
 a17961a <=( A301  and  A300 );
 a17962a <=( (not A299)  and  a17961a );
 a17963a <=( a17962a  and  a17957a );
 a17967a <=( A167  and  (not A169) );
 a17968a <=( A170  and  a17967a );
 a17972a <=( (not A200)  and  (not A199) );
 a17973a <=( (not A166)  and  a17972a );
 a17974a <=( a17973a  and  a17968a );
 a17978a <=( A298  and  (not A266) );
 a17979a <=( (not A265)  and  a17978a );
 a17983a <=( A302  and  A300 );
 a17984a <=( (not A299)  and  a17983a );
 a17985a <=( a17984a  and  a17979a );
 a17989a <=( (not A167)  and  (not A169) );
 a17990a <=( A170  and  a17989a );
 a17994a <=( A200  and  A199 );
 a17995a <=( A166  and  a17994a );
 a17996a <=( a17995a  and  a17990a );
 a18000a <=( A298  and  A266 );
 a18001a <=( A265  and  a18000a );
 a18005a <=( A301  and  A300 );
 a18006a <=( (not A299)  and  a18005a );
 a18007a <=( a18006a  and  a18001a );
 a18011a <=( (not A167)  and  (not A169) );
 a18012a <=( A170  and  a18011a );
 a18016a <=( A200  and  A199 );
 a18017a <=( A166  and  a18016a );
 a18018a <=( a18017a  and  a18012a );
 a18022a <=( A298  and  A266 );
 a18023a <=( A265  and  a18022a );
 a18027a <=( A302  and  A300 );
 a18028a <=( (not A299)  and  a18027a );
 a18029a <=( a18028a  and  a18023a );
 a18033a <=( (not A167)  and  (not A169) );
 a18034a <=( A170  and  a18033a );
 a18038a <=( A200  and  A199 );
 a18039a <=( A166  and  a18038a );
 a18040a <=( a18039a  and  a18034a );
 a18044a <=( A298  and  (not A267) );
 a18045a <=( (not A266)  and  a18044a );
 a18049a <=( A301  and  A300 );
 a18050a <=( (not A299)  and  a18049a );
 a18051a <=( a18050a  and  a18045a );
 a18055a <=( (not A167)  and  (not A169) );
 a18056a <=( A170  and  a18055a );
 a18060a <=( A200  and  A199 );
 a18061a <=( A166  and  a18060a );
 a18062a <=( a18061a  and  a18056a );
 a18066a <=( A298  and  (not A267) );
 a18067a <=( (not A266)  and  a18066a );
 a18071a <=( A302  and  A300 );
 a18072a <=( (not A299)  and  a18071a );
 a18073a <=( a18072a  and  a18067a );
 a18077a <=( (not A167)  and  (not A169) );
 a18078a <=( A170  and  a18077a );
 a18082a <=( A200  and  A199 );
 a18083a <=( A166  and  a18082a );
 a18084a <=( a18083a  and  a18078a );
 a18088a <=( A298  and  (not A266) );
 a18089a <=( (not A265)  and  a18088a );
 a18093a <=( A301  and  A300 );
 a18094a <=( (not A299)  and  a18093a );
 a18095a <=( a18094a  and  a18089a );
 a18099a <=( (not A167)  and  (not A169) );
 a18100a <=( A170  and  a18099a );
 a18104a <=( A200  and  A199 );
 a18105a <=( A166  and  a18104a );
 a18106a <=( a18105a  and  a18100a );
 a18110a <=( A298  and  (not A266) );
 a18111a <=( (not A265)  and  a18110a );
 a18115a <=( A302  and  A300 );
 a18116a <=( (not A299)  and  a18115a );
 a18117a <=( a18116a  and  a18111a );
 a18121a <=( (not A167)  and  (not A169) );
 a18122a <=( A170  and  a18121a );
 a18126a <=( A200  and  (not A199) );
 a18127a <=( A166  and  a18126a );
 a18128a <=( a18127a  and  a18122a );
 a18132a <=( A267  and  (not A266) );
 a18133a <=( A265  and  a18132a );
 a18137a <=( (not A300)  and  A298 );
 a18138a <=( A268  and  a18137a );
 a18139a <=( a18138a  and  a18133a );
 a18143a <=( (not A167)  and  (not A169) );
 a18144a <=( A170  and  a18143a );
 a18148a <=( A200  and  (not A199) );
 a18149a <=( A166  and  a18148a );
 a18150a <=( a18149a  and  a18144a );
 a18154a <=( A267  and  (not A266) );
 a18155a <=( A265  and  a18154a );
 a18159a <=( A299  and  A298 );
 a18160a <=( A268  and  a18159a );
 a18161a <=( a18160a  and  a18155a );
 a18165a <=( (not A167)  and  (not A169) );
 a18166a <=( A170  and  a18165a );
 a18170a <=( A200  and  (not A199) );
 a18171a <=( A166  and  a18170a );
 a18172a <=( a18171a  and  a18166a );
 a18176a <=( A267  and  (not A266) );
 a18177a <=( A265  and  a18176a );
 a18181a <=( (not A299)  and  (not A298) );
 a18182a <=( A268  and  a18181a );
 a18183a <=( a18182a  and  a18177a );
 a18187a <=( (not A167)  and  (not A169) );
 a18188a <=( A170  and  a18187a );
 a18192a <=( A200  and  (not A199) );
 a18193a <=( A166  and  a18192a );
 a18194a <=( a18193a  and  a18188a );
 a18198a <=( A267  and  (not A266) );
 a18199a <=( A265  and  a18198a );
 a18203a <=( (not A300)  and  A298 );
 a18204a <=( A269  and  a18203a );
 a18205a <=( a18204a  and  a18199a );
 a18209a <=( (not A167)  and  (not A169) );
 a18210a <=( A170  and  a18209a );
 a18214a <=( A200  and  (not A199) );
 a18215a <=( A166  and  a18214a );
 a18216a <=( a18215a  and  a18210a );
 a18220a <=( A267  and  (not A266) );
 a18221a <=( A265  and  a18220a );
 a18225a <=( A299  and  A298 );
 a18226a <=( A269  and  a18225a );
 a18227a <=( a18226a  and  a18221a );
 a18231a <=( (not A167)  and  (not A169) );
 a18232a <=( A170  and  a18231a );
 a18236a <=( A200  and  (not A199) );
 a18237a <=( A166  and  a18236a );
 a18238a <=( a18237a  and  a18232a );
 a18242a <=( A267  and  (not A266) );
 a18243a <=( A265  and  a18242a );
 a18247a <=( (not A299)  and  (not A298) );
 a18248a <=( A269  and  a18247a );
 a18249a <=( a18248a  and  a18243a );
 a18253a <=( (not A167)  and  (not A169) );
 a18254a <=( A170  and  a18253a );
 a18258a <=( (not A202)  and  (not A200) );
 a18259a <=( A166  and  a18258a );
 a18260a <=( a18259a  and  a18254a );
 a18264a <=( (not A268)  and  (not A266) );
 a18265a <=( (not A203)  and  a18264a );
 a18269a <=( A299  and  (not A298) );
 a18270a <=( (not A269)  and  a18269a );
 a18271a <=( a18270a  and  a18265a );
 a18275a <=( (not A167)  and  (not A169) );
 a18276a <=( A170  and  a18275a );
 a18280a <=( (not A201)  and  (not A200) );
 a18281a <=( A166  and  a18280a );
 a18282a <=( a18281a  and  a18276a );
 a18286a <=( A298  and  A266 );
 a18287a <=( A265  and  a18286a );
 a18291a <=( A301  and  A300 );
 a18292a <=( (not A299)  and  a18291a );
 a18293a <=( a18292a  and  a18287a );
 a18297a <=( (not A167)  and  (not A169) );
 a18298a <=( A170  and  a18297a );
 a18302a <=( (not A201)  and  (not A200) );
 a18303a <=( A166  and  a18302a );
 a18304a <=( a18303a  and  a18298a );
 a18308a <=( A298  and  A266 );
 a18309a <=( A265  and  a18308a );
 a18313a <=( A302  and  A300 );
 a18314a <=( (not A299)  and  a18313a );
 a18315a <=( a18314a  and  a18309a );
 a18319a <=( (not A167)  and  (not A169) );
 a18320a <=( A170  and  a18319a );
 a18324a <=( (not A201)  and  (not A200) );
 a18325a <=( A166  and  a18324a );
 a18326a <=( a18325a  and  a18320a );
 a18330a <=( A298  and  (not A267) );
 a18331a <=( (not A266)  and  a18330a );
 a18335a <=( A301  and  A300 );
 a18336a <=( (not A299)  and  a18335a );
 a18337a <=( a18336a  and  a18331a );
 a18341a <=( (not A167)  and  (not A169) );
 a18342a <=( A170  and  a18341a );
 a18346a <=( (not A201)  and  (not A200) );
 a18347a <=( A166  and  a18346a );
 a18348a <=( a18347a  and  a18342a );
 a18352a <=( A298  and  (not A267) );
 a18353a <=( (not A266)  and  a18352a );
 a18357a <=( A302  and  A300 );
 a18358a <=( (not A299)  and  a18357a );
 a18359a <=( a18358a  and  a18353a );
 a18363a <=( (not A167)  and  (not A169) );
 a18364a <=( A170  and  a18363a );
 a18368a <=( (not A201)  and  (not A200) );
 a18369a <=( A166  and  a18368a );
 a18370a <=( a18369a  and  a18364a );
 a18374a <=( A298  and  (not A266) );
 a18375a <=( (not A265)  and  a18374a );
 a18379a <=( A301  and  A300 );
 a18380a <=( (not A299)  and  a18379a );
 a18381a <=( a18380a  and  a18375a );
 a18385a <=( (not A167)  and  (not A169) );
 a18386a <=( A170  and  a18385a );
 a18390a <=( (not A201)  and  (not A200) );
 a18391a <=( A166  and  a18390a );
 a18392a <=( a18391a  and  a18386a );
 a18396a <=( A298  and  (not A266) );
 a18397a <=( (not A265)  and  a18396a );
 a18401a <=( A302  and  A300 );
 a18402a <=( (not A299)  and  a18401a );
 a18403a <=( a18402a  and  a18397a );
 a18407a <=( (not A167)  and  (not A169) );
 a18408a <=( A170  and  a18407a );
 a18412a <=( (not A200)  and  A199 );
 a18413a <=( A166  and  a18412a );
 a18414a <=( a18413a  and  a18408a );
 a18418a <=( (not A265)  and  A202 );
 a18419a <=( A201  and  a18418a );
 a18423a <=( (not A300)  and  A298 );
 a18424a <=( A266  and  a18423a );
 a18425a <=( a18424a  and  a18419a );
 a18429a <=( (not A167)  and  (not A169) );
 a18430a <=( A170  and  a18429a );
 a18434a <=( (not A200)  and  A199 );
 a18435a <=( A166  and  a18434a );
 a18436a <=( a18435a  and  a18430a );
 a18440a <=( (not A265)  and  A202 );
 a18441a <=( A201  and  a18440a );
 a18445a <=( A299  and  A298 );
 a18446a <=( A266  and  a18445a );
 a18447a <=( a18446a  and  a18441a );
 a18451a <=( (not A167)  and  (not A169) );
 a18452a <=( A170  and  a18451a );
 a18456a <=( (not A200)  and  A199 );
 a18457a <=( A166  and  a18456a );
 a18458a <=( a18457a  and  a18452a );
 a18462a <=( (not A265)  and  A202 );
 a18463a <=( A201  and  a18462a );
 a18467a <=( (not A299)  and  (not A298) );
 a18468a <=( A266  and  a18467a );
 a18469a <=( a18468a  and  a18463a );
 a18473a <=( (not A167)  and  (not A169) );
 a18474a <=( A170  and  a18473a );
 a18478a <=( (not A200)  and  A199 );
 a18479a <=( A166  and  a18478a );
 a18480a <=( a18479a  and  a18474a );
 a18484a <=( (not A265)  and  A203 );
 a18485a <=( A201  and  a18484a );
 a18489a <=( (not A300)  and  A298 );
 a18490a <=( A266  and  a18489a );
 a18491a <=( a18490a  and  a18485a );
 a18495a <=( (not A167)  and  (not A169) );
 a18496a <=( A170  and  a18495a );
 a18500a <=( (not A200)  and  A199 );
 a18501a <=( A166  and  a18500a );
 a18502a <=( a18501a  and  a18496a );
 a18506a <=( (not A265)  and  A203 );
 a18507a <=( A201  and  a18506a );
 a18511a <=( A299  and  A298 );
 a18512a <=( A266  and  a18511a );
 a18513a <=( a18512a  and  a18507a );
 a18517a <=( (not A167)  and  (not A169) );
 a18518a <=( A170  and  a18517a );
 a18522a <=( (not A200)  and  A199 );
 a18523a <=( A166  and  a18522a );
 a18524a <=( a18523a  and  a18518a );
 a18528a <=( (not A265)  and  A203 );
 a18529a <=( A201  and  a18528a );
 a18533a <=( (not A299)  and  (not A298) );
 a18534a <=( A266  and  a18533a );
 a18535a <=( a18534a  and  a18529a );
 a18539a <=( (not A167)  and  (not A169) );
 a18540a <=( A170  and  a18539a );
 a18544a <=( (not A200)  and  (not A199) );
 a18545a <=( A166  and  a18544a );
 a18546a <=( a18545a  and  a18540a );
 a18550a <=( A298  and  A266 );
 a18551a <=( A265  and  a18550a );
 a18555a <=( A301  and  A300 );
 a18556a <=( (not A299)  and  a18555a );
 a18557a <=( a18556a  and  a18551a );
 a18561a <=( (not A167)  and  (not A169) );
 a18562a <=( A170  and  a18561a );
 a18566a <=( (not A200)  and  (not A199) );
 a18567a <=( A166  and  a18566a );
 a18568a <=( a18567a  and  a18562a );
 a18572a <=( A298  and  A266 );
 a18573a <=( A265  and  a18572a );
 a18577a <=( A302  and  A300 );
 a18578a <=( (not A299)  and  a18577a );
 a18579a <=( a18578a  and  a18573a );
 a18583a <=( (not A167)  and  (not A169) );
 a18584a <=( A170  and  a18583a );
 a18588a <=( (not A200)  and  (not A199) );
 a18589a <=( A166  and  a18588a );
 a18590a <=( a18589a  and  a18584a );
 a18594a <=( A298  and  (not A267) );
 a18595a <=( (not A266)  and  a18594a );
 a18599a <=( A301  and  A300 );
 a18600a <=( (not A299)  and  a18599a );
 a18601a <=( a18600a  and  a18595a );
 a18605a <=( (not A167)  and  (not A169) );
 a18606a <=( A170  and  a18605a );
 a18610a <=( (not A200)  and  (not A199) );
 a18611a <=( A166  and  a18610a );
 a18612a <=( a18611a  and  a18606a );
 a18616a <=( A298  and  (not A267) );
 a18617a <=( (not A266)  and  a18616a );
 a18621a <=( A302  and  A300 );
 a18622a <=( (not A299)  and  a18621a );
 a18623a <=( a18622a  and  a18617a );
 a18627a <=( (not A167)  and  (not A169) );
 a18628a <=( A170  and  a18627a );
 a18632a <=( (not A200)  and  (not A199) );
 a18633a <=( A166  and  a18632a );
 a18634a <=( a18633a  and  a18628a );
 a18638a <=( A298  and  (not A266) );
 a18639a <=( (not A265)  and  a18638a );
 a18643a <=( A301  and  A300 );
 a18644a <=( (not A299)  and  a18643a );
 a18645a <=( a18644a  and  a18639a );
 a18649a <=( (not A167)  and  (not A169) );
 a18650a <=( A170  and  a18649a );
 a18654a <=( (not A200)  and  (not A199) );
 a18655a <=( A166  and  a18654a );
 a18656a <=( a18655a  and  a18650a );
 a18660a <=( A298  and  (not A266) );
 a18661a <=( (not A265)  and  a18660a );
 a18665a <=( A302  and  A300 );
 a18666a <=( (not A299)  and  a18665a );
 a18667a <=( a18666a  and  a18661a );
 a18671a <=( (not A168)  and  (not A169) );
 a18672a <=( (not A170)  and  a18671a );
 a18676a <=( A265  and  A200 );
 a18677a <=( A199  and  a18676a );
 a18678a <=( a18677a  and  a18672a );
 a18682a <=( A268  and  A267 );
 a18683a <=( (not A266)  and  a18682a );
 a18687a <=( (not A302)  and  (not A301) );
 a18688a <=( A298  and  a18687a );
 a18689a <=( a18688a  and  a18683a );
 a18693a <=( (not A168)  and  (not A169) );
 a18694a <=( (not A170)  and  a18693a );
 a18698a <=( A265  and  A200 );
 a18699a <=( A199  and  a18698a );
 a18700a <=( a18699a  and  a18694a );
 a18704a <=( A269  and  A267 );
 a18705a <=( (not A266)  and  a18704a );
 a18709a <=( (not A302)  and  (not A301) );
 a18710a <=( A298  and  a18709a );
 a18711a <=( a18710a  and  a18705a );
 a18715a <=( (not A168)  and  (not A169) );
 a18716a <=( (not A170)  and  a18715a );
 a18720a <=( (not A266)  and  A200 );
 a18721a <=( (not A199)  and  a18720a );
 a18722a <=( a18721a  and  a18716a );
 a18726a <=( A298  and  (not A269) );
 a18727a <=( (not A268)  and  a18726a );
 a18731a <=( A301  and  A300 );
 a18732a <=( (not A299)  and  a18731a );
 a18733a <=( a18732a  and  a18727a );
 a18737a <=( (not A168)  and  (not A169) );
 a18738a <=( (not A170)  and  a18737a );
 a18742a <=( (not A266)  and  A200 );
 a18743a <=( (not A199)  and  a18742a );
 a18744a <=( a18743a  and  a18738a );
 a18748a <=( A298  and  (not A269) );
 a18749a <=( (not A268)  and  a18748a );
 a18753a <=( A302  and  A300 );
 a18754a <=( (not A299)  and  a18753a );
 a18755a <=( a18754a  and  a18749a );
 a18759a <=( (not A168)  and  (not A169) );
 a18760a <=( (not A170)  and  a18759a );
 a18764a <=( (not A203)  and  (not A202) );
 a18765a <=( (not A200)  and  a18764a );
 a18766a <=( a18765a  and  a18760a );
 a18770a <=( A267  and  (not A266) );
 a18771a <=( A265  and  a18770a );
 a18775a <=( (not A300)  and  A298 );
 a18776a <=( A268  and  a18775a );
 a18777a <=( a18776a  and  a18771a );
 a18781a <=( (not A168)  and  (not A169) );
 a18782a <=( (not A170)  and  a18781a );
 a18786a <=( (not A203)  and  (not A202) );
 a18787a <=( (not A200)  and  a18786a );
 a18788a <=( a18787a  and  a18782a );
 a18792a <=( A267  and  (not A266) );
 a18793a <=( A265  and  a18792a );
 a18797a <=( A299  and  A298 );
 a18798a <=( A268  and  a18797a );
 a18799a <=( a18798a  and  a18793a );
 a18803a <=( (not A168)  and  (not A169) );
 a18804a <=( (not A170)  and  a18803a );
 a18808a <=( (not A203)  and  (not A202) );
 a18809a <=( (not A200)  and  a18808a );
 a18810a <=( a18809a  and  a18804a );
 a18814a <=( A267  and  (not A266) );
 a18815a <=( A265  and  a18814a );
 a18819a <=( (not A299)  and  (not A298) );
 a18820a <=( A268  and  a18819a );
 a18821a <=( a18820a  and  a18815a );
 a18825a <=( (not A168)  and  (not A169) );
 a18826a <=( (not A170)  and  a18825a );
 a18830a <=( (not A203)  and  (not A202) );
 a18831a <=( (not A200)  and  a18830a );
 a18832a <=( a18831a  and  a18826a );
 a18836a <=( A267  and  (not A266) );
 a18837a <=( A265  and  a18836a );
 a18841a <=( (not A300)  and  A298 );
 a18842a <=( A269  and  a18841a );
 a18843a <=( a18842a  and  a18837a );
 a18847a <=( (not A168)  and  (not A169) );
 a18848a <=( (not A170)  and  a18847a );
 a18852a <=( (not A203)  and  (not A202) );
 a18853a <=( (not A200)  and  a18852a );
 a18854a <=( a18853a  and  a18848a );
 a18858a <=( A267  and  (not A266) );
 a18859a <=( A265  and  a18858a );
 a18863a <=( A299  and  A298 );
 a18864a <=( A269  and  a18863a );
 a18865a <=( a18864a  and  a18859a );
 a18869a <=( (not A168)  and  (not A169) );
 a18870a <=( (not A170)  and  a18869a );
 a18874a <=( (not A203)  and  (not A202) );
 a18875a <=( (not A200)  and  a18874a );
 a18876a <=( a18875a  and  a18870a );
 a18880a <=( A267  and  (not A266) );
 a18881a <=( A265  and  a18880a );
 a18885a <=( (not A299)  and  (not A298) );
 a18886a <=( A269  and  a18885a );
 a18887a <=( a18886a  and  a18881a );
 a18891a <=( (not A168)  and  (not A169) );
 a18892a <=( (not A170)  and  a18891a );
 a18896a <=( A265  and  (not A201) );
 a18897a <=( (not A200)  and  a18896a );
 a18898a <=( a18897a  and  a18892a );
 a18902a <=( A268  and  A267 );
 a18903a <=( (not A266)  and  a18902a );
 a18907a <=( (not A302)  and  (not A301) );
 a18908a <=( A298  and  a18907a );
 a18909a <=( a18908a  and  a18903a );
 a18913a <=( (not A168)  and  (not A169) );
 a18914a <=( (not A170)  and  a18913a );
 a18918a <=( A265  and  (not A201) );
 a18919a <=( (not A200)  and  a18918a );
 a18920a <=( a18919a  and  a18914a );
 a18924a <=( A269  and  A267 );
 a18925a <=( (not A266)  and  a18924a );
 a18929a <=( (not A302)  and  (not A301) );
 a18930a <=( A298  and  a18929a );
 a18931a <=( a18930a  and  a18925a );
 a18935a <=( (not A168)  and  (not A169) );
 a18936a <=( (not A170)  and  a18935a );
 a18940a <=( A201  and  (not A200) );
 a18941a <=( A199  and  a18940a );
 a18942a <=( a18941a  and  a18936a );
 a18946a <=( (not A268)  and  (not A266) );
 a18947a <=( A202  and  a18946a );
 a18951a <=( A299  and  (not A298) );
 a18952a <=( (not A269)  and  a18951a );
 a18953a <=( a18952a  and  a18947a );
 a18957a <=( (not A168)  and  (not A169) );
 a18958a <=( (not A170)  and  a18957a );
 a18962a <=( A201  and  (not A200) );
 a18963a <=( A199  and  a18962a );
 a18964a <=( a18963a  and  a18958a );
 a18968a <=( (not A268)  and  (not A266) );
 a18969a <=( A203  and  a18968a );
 a18973a <=( A299  and  (not A298) );
 a18974a <=( (not A269)  and  a18973a );
 a18975a <=( a18974a  and  a18969a );
 a18979a <=( (not A168)  and  (not A169) );
 a18980a <=( (not A170)  and  a18979a );
 a18984a <=( A265  and  (not A200) );
 a18985a <=( (not A199)  and  a18984a );
 a18986a <=( a18985a  and  a18980a );
 a18990a <=( A268  and  A267 );
 a18991a <=( (not A266)  and  a18990a );
 a18995a <=( (not A302)  and  (not A301) );
 a18996a <=( A298  and  a18995a );
 a18997a <=( a18996a  and  a18991a );
 a19001a <=( (not A168)  and  (not A169) );
 a19002a <=( (not A170)  and  a19001a );
 a19006a <=( A265  and  (not A200) );
 a19007a <=( (not A199)  and  a19006a );
 a19008a <=( a19007a  and  a19002a );
 a19012a <=( A269  and  A267 );
 a19013a <=( (not A266)  and  a19012a );
 a19017a <=( (not A302)  and  (not A301) );
 a19018a <=( A298  and  a19017a );
 a19019a <=( a19018a  and  a19013a );
 a19023a <=( A199  and  A166 );
 a19024a <=( A168  and  a19023a );
 a19028a <=( A202  and  A201 );
 a19029a <=( (not A200)  and  a19028a );
 a19030a <=( a19029a  and  a19024a );
 a19034a <=( A267  and  (not A266) );
 a19035a <=( A265  and  a19034a );
 a19038a <=( A298  and  A268 );
 a19041a <=( (not A302)  and  (not A301) );
 a19042a <=( a19041a  and  a19038a );
 a19043a <=( a19042a  and  a19035a );
 a19047a <=( A199  and  A166 );
 a19048a <=( A168  and  a19047a );
 a19052a <=( A202  and  A201 );
 a19053a <=( (not A200)  and  a19052a );
 a19054a <=( a19053a  and  a19048a );
 a19058a <=( A267  and  (not A266) );
 a19059a <=( A265  and  a19058a );
 a19062a <=( A298  and  A269 );
 a19065a <=( (not A302)  and  (not A301) );
 a19066a <=( a19065a  and  a19062a );
 a19067a <=( a19066a  and  a19059a );
 a19071a <=( A199  and  A166 );
 a19072a <=( A168  and  a19071a );
 a19076a <=( A203  and  A201 );
 a19077a <=( (not A200)  and  a19076a );
 a19078a <=( a19077a  and  a19072a );
 a19082a <=( A267  and  (not A266) );
 a19083a <=( A265  and  a19082a );
 a19086a <=( A298  and  A268 );
 a19089a <=( (not A302)  and  (not A301) );
 a19090a <=( a19089a  and  a19086a );
 a19091a <=( a19090a  and  a19083a );
 a19095a <=( A199  and  A166 );
 a19096a <=( A168  and  a19095a );
 a19100a <=( A203  and  A201 );
 a19101a <=( (not A200)  and  a19100a );
 a19102a <=( a19101a  and  a19096a );
 a19106a <=( A267  and  (not A266) );
 a19107a <=( A265  and  a19106a );
 a19110a <=( A298  and  A269 );
 a19113a <=( (not A302)  and  (not A301) );
 a19114a <=( a19113a  and  a19110a );
 a19115a <=( a19114a  and  a19107a );
 a19119a <=( A199  and  A167 );
 a19120a <=( A168  and  a19119a );
 a19124a <=( A202  and  A201 );
 a19125a <=( (not A200)  and  a19124a );
 a19126a <=( a19125a  and  a19120a );
 a19130a <=( A267  and  (not A266) );
 a19131a <=( A265  and  a19130a );
 a19134a <=( A298  and  A268 );
 a19137a <=( (not A302)  and  (not A301) );
 a19138a <=( a19137a  and  a19134a );
 a19139a <=( a19138a  and  a19131a );
 a19143a <=( A199  and  A167 );
 a19144a <=( A168  and  a19143a );
 a19148a <=( A202  and  A201 );
 a19149a <=( (not A200)  and  a19148a );
 a19150a <=( a19149a  and  a19144a );
 a19154a <=( A267  and  (not A266) );
 a19155a <=( A265  and  a19154a );
 a19158a <=( A298  and  A269 );
 a19161a <=( (not A302)  and  (not A301) );
 a19162a <=( a19161a  and  a19158a );
 a19163a <=( a19162a  and  a19155a );
 a19167a <=( A199  and  A167 );
 a19168a <=( A168  and  a19167a );
 a19172a <=( A203  and  A201 );
 a19173a <=( (not A200)  and  a19172a );
 a19174a <=( a19173a  and  a19168a );
 a19178a <=( A267  and  (not A266) );
 a19179a <=( A265  and  a19178a );
 a19182a <=( A298  and  A268 );
 a19185a <=( (not A302)  and  (not A301) );
 a19186a <=( a19185a  and  a19182a );
 a19187a <=( a19186a  and  a19179a );
 a19191a <=( A199  and  A167 );
 a19192a <=( A168  and  a19191a );
 a19196a <=( A203  and  A201 );
 a19197a <=( (not A200)  and  a19196a );
 a19198a <=( a19197a  and  a19192a );
 a19202a <=( A267  and  (not A266) );
 a19203a <=( A265  and  a19202a );
 a19206a <=( A298  and  A269 );
 a19209a <=( (not A302)  and  (not A301) );
 a19210a <=( a19209a  and  a19206a );
 a19211a <=( a19210a  and  a19203a );
 a19215a <=( (not A166)  and  (not A167) );
 a19216a <=( A170  and  a19215a );
 a19220a <=( (not A203)  and  (not A202) );
 a19221a <=( (not A200)  and  a19220a );
 a19222a <=( a19221a  and  a19216a );
 a19226a <=( A267  and  (not A266) );
 a19227a <=( A265  and  a19226a );
 a19230a <=( A298  and  A268 );
 a19233a <=( (not A302)  and  (not A301) );
 a19234a <=( a19233a  and  a19230a );
 a19235a <=( a19234a  and  a19227a );
 a19239a <=( (not A166)  and  (not A167) );
 a19240a <=( A170  and  a19239a );
 a19244a <=( (not A203)  and  (not A202) );
 a19245a <=( (not A200)  and  a19244a );
 a19246a <=( a19245a  and  a19240a );
 a19250a <=( A267  and  (not A266) );
 a19251a <=( A265  and  a19250a );
 a19254a <=( A298  and  A269 );
 a19257a <=( (not A302)  and  (not A301) );
 a19258a <=( a19257a  and  a19254a );
 a19259a <=( a19258a  and  a19251a );
 a19263a <=( (not A166)  and  (not A167) );
 a19264a <=( A170  and  a19263a );
 a19268a <=( A201  and  (not A200) );
 a19269a <=( A199  and  a19268a );
 a19270a <=( a19269a  and  a19264a );
 a19274a <=( A266  and  A265 );
 a19275a <=( A202  and  a19274a );
 a19278a <=( (not A299)  and  A298 );
 a19281a <=( A301  and  A300 );
 a19282a <=( a19281a  and  a19278a );
 a19283a <=( a19282a  and  a19275a );
 a19287a <=( (not A166)  and  (not A167) );
 a19288a <=( A170  and  a19287a );
 a19292a <=( A201  and  (not A200) );
 a19293a <=( A199  and  a19292a );
 a19294a <=( a19293a  and  a19288a );
 a19298a <=( A266  and  A265 );
 a19299a <=( A202  and  a19298a );
 a19302a <=( (not A299)  and  A298 );
 a19305a <=( A302  and  A300 );
 a19306a <=( a19305a  and  a19302a );
 a19307a <=( a19306a  and  a19299a );
 a19311a <=( (not A166)  and  (not A167) );
 a19312a <=( A170  and  a19311a );
 a19316a <=( A201  and  (not A200) );
 a19317a <=( A199  and  a19316a );
 a19318a <=( a19317a  and  a19312a );
 a19322a <=( (not A267)  and  (not A266) );
 a19323a <=( A202  and  a19322a );
 a19326a <=( (not A299)  and  A298 );
 a19329a <=( A301  and  A300 );
 a19330a <=( a19329a  and  a19326a );
 a19331a <=( a19330a  and  a19323a );
 a19335a <=( (not A166)  and  (not A167) );
 a19336a <=( A170  and  a19335a );
 a19340a <=( A201  and  (not A200) );
 a19341a <=( A199  and  a19340a );
 a19342a <=( a19341a  and  a19336a );
 a19346a <=( (not A267)  and  (not A266) );
 a19347a <=( A202  and  a19346a );
 a19350a <=( (not A299)  and  A298 );
 a19353a <=( A302  and  A300 );
 a19354a <=( a19353a  and  a19350a );
 a19355a <=( a19354a  and  a19347a );
 a19359a <=( (not A166)  and  (not A167) );
 a19360a <=( A170  and  a19359a );
 a19364a <=( A201  and  (not A200) );
 a19365a <=( A199  and  a19364a );
 a19366a <=( a19365a  and  a19360a );
 a19370a <=( (not A266)  and  (not A265) );
 a19371a <=( A202  and  a19370a );
 a19374a <=( (not A299)  and  A298 );
 a19377a <=( A301  and  A300 );
 a19378a <=( a19377a  and  a19374a );
 a19379a <=( a19378a  and  a19371a );
 a19383a <=( (not A166)  and  (not A167) );
 a19384a <=( A170  and  a19383a );
 a19388a <=( A201  and  (not A200) );
 a19389a <=( A199  and  a19388a );
 a19390a <=( a19389a  and  a19384a );
 a19394a <=( (not A266)  and  (not A265) );
 a19395a <=( A202  and  a19394a );
 a19398a <=( (not A299)  and  A298 );
 a19401a <=( A302  and  A300 );
 a19402a <=( a19401a  and  a19398a );
 a19403a <=( a19402a  and  a19395a );
 a19407a <=( (not A166)  and  (not A167) );
 a19408a <=( A170  and  a19407a );
 a19412a <=( A201  and  (not A200) );
 a19413a <=( A199  and  a19412a );
 a19414a <=( a19413a  and  a19408a );
 a19418a <=( A266  and  A265 );
 a19419a <=( A203  and  a19418a );
 a19422a <=( (not A299)  and  A298 );
 a19425a <=( A301  and  A300 );
 a19426a <=( a19425a  and  a19422a );
 a19427a <=( a19426a  and  a19419a );
 a19431a <=( (not A166)  and  (not A167) );
 a19432a <=( A170  and  a19431a );
 a19436a <=( A201  and  (not A200) );
 a19437a <=( A199  and  a19436a );
 a19438a <=( a19437a  and  a19432a );
 a19442a <=( A266  and  A265 );
 a19443a <=( A203  and  a19442a );
 a19446a <=( (not A299)  and  A298 );
 a19449a <=( A302  and  A300 );
 a19450a <=( a19449a  and  a19446a );
 a19451a <=( a19450a  and  a19443a );
 a19455a <=( (not A166)  and  (not A167) );
 a19456a <=( A170  and  a19455a );
 a19460a <=( A201  and  (not A200) );
 a19461a <=( A199  and  a19460a );
 a19462a <=( a19461a  and  a19456a );
 a19466a <=( (not A267)  and  (not A266) );
 a19467a <=( A203  and  a19466a );
 a19470a <=( (not A299)  and  A298 );
 a19473a <=( A301  and  A300 );
 a19474a <=( a19473a  and  a19470a );
 a19475a <=( a19474a  and  a19467a );
 a19479a <=( (not A166)  and  (not A167) );
 a19480a <=( A170  and  a19479a );
 a19484a <=( A201  and  (not A200) );
 a19485a <=( A199  and  a19484a );
 a19486a <=( a19485a  and  a19480a );
 a19490a <=( (not A267)  and  (not A266) );
 a19491a <=( A203  and  a19490a );
 a19494a <=( (not A299)  and  A298 );
 a19497a <=( A302  and  A300 );
 a19498a <=( a19497a  and  a19494a );
 a19499a <=( a19498a  and  a19491a );
 a19503a <=( (not A166)  and  (not A167) );
 a19504a <=( A170  and  a19503a );
 a19508a <=( A201  and  (not A200) );
 a19509a <=( A199  and  a19508a );
 a19510a <=( a19509a  and  a19504a );
 a19514a <=( (not A266)  and  (not A265) );
 a19515a <=( A203  and  a19514a );
 a19518a <=( (not A299)  and  A298 );
 a19521a <=( A301  and  A300 );
 a19522a <=( a19521a  and  a19518a );
 a19523a <=( a19522a  and  a19515a );
 a19527a <=( (not A166)  and  (not A167) );
 a19528a <=( A170  and  a19527a );
 a19532a <=( A201  and  (not A200) );
 a19533a <=( A199  and  a19532a );
 a19534a <=( a19533a  and  a19528a );
 a19538a <=( (not A266)  and  (not A265) );
 a19539a <=( A203  and  a19538a );
 a19542a <=( (not A299)  and  A298 );
 a19545a <=( A302  and  A300 );
 a19546a <=( a19545a  and  a19542a );
 a19547a <=( a19546a  and  a19539a );
 a19551a <=( A167  and  (not A168) );
 a19552a <=( A169  and  a19551a );
 a19556a <=( A200  and  A199 );
 a19557a <=( (not A166)  and  a19556a );
 a19558a <=( a19557a  and  a19552a );
 a19562a <=( A267  and  (not A266) );
 a19563a <=( A265  and  a19562a );
 a19566a <=( A298  and  A268 );
 a19569a <=( (not A302)  and  (not A301) );
 a19570a <=( a19569a  and  a19566a );
 a19571a <=( a19570a  and  a19563a );
 a19575a <=( A167  and  (not A168) );
 a19576a <=( A169  and  a19575a );
 a19580a <=( A200  and  A199 );
 a19581a <=( (not A166)  and  a19580a );
 a19582a <=( a19581a  and  a19576a );
 a19586a <=( A267  and  (not A266) );
 a19587a <=( A265  and  a19586a );
 a19590a <=( A298  and  A269 );
 a19593a <=( (not A302)  and  (not A301) );
 a19594a <=( a19593a  and  a19590a );
 a19595a <=( a19594a  and  a19587a );
 a19599a <=( A167  and  (not A168) );
 a19600a <=( A169  and  a19599a );
 a19604a <=( A200  and  (not A199) );
 a19605a <=( (not A166)  and  a19604a );
 a19606a <=( a19605a  and  a19600a );
 a19610a <=( (not A269)  and  (not A268) );
 a19611a <=( (not A266)  and  a19610a );
 a19614a <=( (not A299)  and  A298 );
 a19617a <=( A301  and  A300 );
 a19618a <=( a19617a  and  a19614a );
 a19619a <=( a19618a  and  a19611a );
 a19623a <=( A167  and  (not A168) );
 a19624a <=( A169  and  a19623a );
 a19628a <=( A200  and  (not A199) );
 a19629a <=( (not A166)  and  a19628a );
 a19630a <=( a19629a  and  a19624a );
 a19634a <=( (not A269)  and  (not A268) );
 a19635a <=( (not A266)  and  a19634a );
 a19638a <=( (not A299)  and  A298 );
 a19641a <=( A302  and  A300 );
 a19642a <=( a19641a  and  a19638a );
 a19643a <=( a19642a  and  a19635a );
 a19647a <=( A167  and  (not A168) );
 a19648a <=( A169  and  a19647a );
 a19652a <=( (not A202)  and  (not A200) );
 a19653a <=( (not A166)  and  a19652a );
 a19654a <=( a19653a  and  a19648a );
 a19658a <=( (not A266)  and  A265 );
 a19659a <=( (not A203)  and  a19658a );
 a19662a <=( A268  and  A267 );
 a19665a <=( (not A300)  and  A298 );
 a19666a <=( a19665a  and  a19662a );
 a19667a <=( a19666a  and  a19659a );
 a19671a <=( A167  and  (not A168) );
 a19672a <=( A169  and  a19671a );
 a19676a <=( (not A202)  and  (not A200) );
 a19677a <=( (not A166)  and  a19676a );
 a19678a <=( a19677a  and  a19672a );
 a19682a <=( (not A266)  and  A265 );
 a19683a <=( (not A203)  and  a19682a );
 a19686a <=( A268  and  A267 );
 a19689a <=( A299  and  A298 );
 a19690a <=( a19689a  and  a19686a );
 a19691a <=( a19690a  and  a19683a );
 a19695a <=( A167  and  (not A168) );
 a19696a <=( A169  and  a19695a );
 a19700a <=( (not A202)  and  (not A200) );
 a19701a <=( (not A166)  and  a19700a );
 a19702a <=( a19701a  and  a19696a );
 a19706a <=( (not A266)  and  A265 );
 a19707a <=( (not A203)  and  a19706a );
 a19710a <=( A268  and  A267 );
 a19713a <=( (not A299)  and  (not A298) );
 a19714a <=( a19713a  and  a19710a );
 a19715a <=( a19714a  and  a19707a );
 a19719a <=( A167  and  (not A168) );
 a19720a <=( A169  and  a19719a );
 a19724a <=( (not A202)  and  (not A200) );
 a19725a <=( (not A166)  and  a19724a );
 a19726a <=( a19725a  and  a19720a );
 a19730a <=( (not A266)  and  A265 );
 a19731a <=( (not A203)  and  a19730a );
 a19734a <=( A269  and  A267 );
 a19737a <=( (not A300)  and  A298 );
 a19738a <=( a19737a  and  a19734a );
 a19739a <=( a19738a  and  a19731a );
 a19743a <=( A167  and  (not A168) );
 a19744a <=( A169  and  a19743a );
 a19748a <=( (not A202)  and  (not A200) );
 a19749a <=( (not A166)  and  a19748a );
 a19750a <=( a19749a  and  a19744a );
 a19754a <=( (not A266)  and  A265 );
 a19755a <=( (not A203)  and  a19754a );
 a19758a <=( A269  and  A267 );
 a19761a <=( A299  and  A298 );
 a19762a <=( a19761a  and  a19758a );
 a19763a <=( a19762a  and  a19755a );
 a19767a <=( A167  and  (not A168) );
 a19768a <=( A169  and  a19767a );
 a19772a <=( (not A202)  and  (not A200) );
 a19773a <=( (not A166)  and  a19772a );
 a19774a <=( a19773a  and  a19768a );
 a19778a <=( (not A266)  and  A265 );
 a19779a <=( (not A203)  and  a19778a );
 a19782a <=( A269  and  A267 );
 a19785a <=( (not A299)  and  (not A298) );
 a19786a <=( a19785a  and  a19782a );
 a19787a <=( a19786a  and  a19779a );
 a19791a <=( A167  and  (not A168) );
 a19792a <=( A169  and  a19791a );
 a19796a <=( (not A201)  and  (not A200) );
 a19797a <=( (not A166)  and  a19796a );
 a19798a <=( a19797a  and  a19792a );
 a19802a <=( A267  and  (not A266) );
 a19803a <=( A265  and  a19802a );
 a19806a <=( A298  and  A268 );
 a19809a <=( (not A302)  and  (not A301) );
 a19810a <=( a19809a  and  a19806a );
 a19811a <=( a19810a  and  a19803a );
 a19815a <=( A167  and  (not A168) );
 a19816a <=( A169  and  a19815a );
 a19820a <=( (not A201)  and  (not A200) );
 a19821a <=( (not A166)  and  a19820a );
 a19822a <=( a19821a  and  a19816a );
 a19826a <=( A267  and  (not A266) );
 a19827a <=( A265  and  a19826a );
 a19830a <=( A298  and  A269 );
 a19833a <=( (not A302)  and  (not A301) );
 a19834a <=( a19833a  and  a19830a );
 a19835a <=( a19834a  and  a19827a );
 a19839a <=( A167  and  (not A168) );
 a19840a <=( A169  and  a19839a );
 a19844a <=( (not A200)  and  A199 );
 a19845a <=( (not A166)  and  a19844a );
 a19846a <=( a19845a  and  a19840a );
 a19850a <=( (not A266)  and  A202 );
 a19851a <=( A201  and  a19850a );
 a19854a <=( (not A269)  and  (not A268) );
 a19857a <=( A299  and  (not A298) );
 a19858a <=( a19857a  and  a19854a );
 a19859a <=( a19858a  and  a19851a );
 a19863a <=( A167  and  (not A168) );
 a19864a <=( A169  and  a19863a );
 a19868a <=( (not A200)  and  A199 );
 a19869a <=( (not A166)  and  a19868a );
 a19870a <=( a19869a  and  a19864a );
 a19874a <=( (not A266)  and  A203 );
 a19875a <=( A201  and  a19874a );
 a19878a <=( (not A269)  and  (not A268) );
 a19881a <=( A299  and  (not A298) );
 a19882a <=( a19881a  and  a19878a );
 a19883a <=( a19882a  and  a19875a );
 a19887a <=( A167  and  (not A168) );
 a19888a <=( A169  and  a19887a );
 a19892a <=( (not A200)  and  (not A199) );
 a19893a <=( (not A166)  and  a19892a );
 a19894a <=( a19893a  and  a19888a );
 a19898a <=( A267  and  (not A266) );
 a19899a <=( A265  and  a19898a );
 a19902a <=( A298  and  A268 );
 a19905a <=( (not A302)  and  (not A301) );
 a19906a <=( a19905a  and  a19902a );
 a19907a <=( a19906a  and  a19899a );
 a19911a <=( A167  and  (not A168) );
 a19912a <=( A169  and  a19911a );
 a19916a <=( (not A200)  and  (not A199) );
 a19917a <=( (not A166)  and  a19916a );
 a19918a <=( a19917a  and  a19912a );
 a19922a <=( A267  and  (not A266) );
 a19923a <=( A265  and  a19922a );
 a19926a <=( A298  and  A269 );
 a19929a <=( (not A302)  and  (not A301) );
 a19930a <=( a19929a  and  a19926a );
 a19931a <=( a19930a  and  a19923a );
 a19935a <=( (not A167)  and  (not A168) );
 a19936a <=( A169  and  a19935a );
 a19940a <=( A200  and  A199 );
 a19941a <=( A166  and  a19940a );
 a19942a <=( a19941a  and  a19936a );
 a19946a <=( A267  and  (not A266) );
 a19947a <=( A265  and  a19946a );
 a19950a <=( A298  and  A268 );
 a19953a <=( (not A302)  and  (not A301) );
 a19954a <=( a19953a  and  a19950a );
 a19955a <=( a19954a  and  a19947a );
 a19959a <=( (not A167)  and  (not A168) );
 a19960a <=( A169  and  a19959a );
 a19964a <=( A200  and  A199 );
 a19965a <=( A166  and  a19964a );
 a19966a <=( a19965a  and  a19960a );
 a19970a <=( A267  and  (not A266) );
 a19971a <=( A265  and  a19970a );
 a19974a <=( A298  and  A269 );
 a19977a <=( (not A302)  and  (not A301) );
 a19978a <=( a19977a  and  a19974a );
 a19979a <=( a19978a  and  a19971a );
 a19983a <=( (not A167)  and  (not A168) );
 a19984a <=( A169  and  a19983a );
 a19988a <=( A200  and  (not A199) );
 a19989a <=( A166  and  a19988a );
 a19990a <=( a19989a  and  a19984a );
 a19994a <=( (not A269)  and  (not A268) );
 a19995a <=( (not A266)  and  a19994a );
 a19998a <=( (not A299)  and  A298 );
 a20001a <=( A301  and  A300 );
 a20002a <=( a20001a  and  a19998a );
 a20003a <=( a20002a  and  a19995a );
 a20007a <=( (not A167)  and  (not A168) );
 a20008a <=( A169  and  a20007a );
 a20012a <=( A200  and  (not A199) );
 a20013a <=( A166  and  a20012a );
 a20014a <=( a20013a  and  a20008a );
 a20018a <=( (not A269)  and  (not A268) );
 a20019a <=( (not A266)  and  a20018a );
 a20022a <=( (not A299)  and  A298 );
 a20025a <=( A302  and  A300 );
 a20026a <=( a20025a  and  a20022a );
 a20027a <=( a20026a  and  a20019a );
 a20031a <=( (not A167)  and  (not A168) );
 a20032a <=( A169  and  a20031a );
 a20036a <=( (not A202)  and  (not A200) );
 a20037a <=( A166  and  a20036a );
 a20038a <=( a20037a  and  a20032a );
 a20042a <=( (not A266)  and  A265 );
 a20043a <=( (not A203)  and  a20042a );
 a20046a <=( A268  and  A267 );
 a20049a <=( (not A300)  and  A298 );
 a20050a <=( a20049a  and  a20046a );
 a20051a <=( a20050a  and  a20043a );
 a20055a <=( (not A167)  and  (not A168) );
 a20056a <=( A169  and  a20055a );
 a20060a <=( (not A202)  and  (not A200) );
 a20061a <=( A166  and  a20060a );
 a20062a <=( a20061a  and  a20056a );
 a20066a <=( (not A266)  and  A265 );
 a20067a <=( (not A203)  and  a20066a );
 a20070a <=( A268  and  A267 );
 a20073a <=( A299  and  A298 );
 a20074a <=( a20073a  and  a20070a );
 a20075a <=( a20074a  and  a20067a );
 a20079a <=( (not A167)  and  (not A168) );
 a20080a <=( A169  and  a20079a );
 a20084a <=( (not A202)  and  (not A200) );
 a20085a <=( A166  and  a20084a );
 a20086a <=( a20085a  and  a20080a );
 a20090a <=( (not A266)  and  A265 );
 a20091a <=( (not A203)  and  a20090a );
 a20094a <=( A268  and  A267 );
 a20097a <=( (not A299)  and  (not A298) );
 a20098a <=( a20097a  and  a20094a );
 a20099a <=( a20098a  and  a20091a );
 a20103a <=( (not A167)  and  (not A168) );
 a20104a <=( A169  and  a20103a );
 a20108a <=( (not A202)  and  (not A200) );
 a20109a <=( A166  and  a20108a );
 a20110a <=( a20109a  and  a20104a );
 a20114a <=( (not A266)  and  A265 );
 a20115a <=( (not A203)  and  a20114a );
 a20118a <=( A269  and  A267 );
 a20121a <=( (not A300)  and  A298 );
 a20122a <=( a20121a  and  a20118a );
 a20123a <=( a20122a  and  a20115a );
 a20127a <=( (not A167)  and  (not A168) );
 a20128a <=( A169  and  a20127a );
 a20132a <=( (not A202)  and  (not A200) );
 a20133a <=( A166  and  a20132a );
 a20134a <=( a20133a  and  a20128a );
 a20138a <=( (not A266)  and  A265 );
 a20139a <=( (not A203)  and  a20138a );
 a20142a <=( A269  and  A267 );
 a20145a <=( A299  and  A298 );
 a20146a <=( a20145a  and  a20142a );
 a20147a <=( a20146a  and  a20139a );
 a20151a <=( (not A167)  and  (not A168) );
 a20152a <=( A169  and  a20151a );
 a20156a <=( (not A202)  and  (not A200) );
 a20157a <=( A166  and  a20156a );
 a20158a <=( a20157a  and  a20152a );
 a20162a <=( (not A266)  and  A265 );
 a20163a <=( (not A203)  and  a20162a );
 a20166a <=( A269  and  A267 );
 a20169a <=( (not A299)  and  (not A298) );
 a20170a <=( a20169a  and  a20166a );
 a20171a <=( a20170a  and  a20163a );
 a20175a <=( (not A167)  and  (not A168) );
 a20176a <=( A169  and  a20175a );
 a20180a <=( (not A201)  and  (not A200) );
 a20181a <=( A166  and  a20180a );
 a20182a <=( a20181a  and  a20176a );
 a20186a <=( A267  and  (not A266) );
 a20187a <=( A265  and  a20186a );
 a20190a <=( A298  and  A268 );
 a20193a <=( (not A302)  and  (not A301) );
 a20194a <=( a20193a  and  a20190a );
 a20195a <=( a20194a  and  a20187a );
 a20199a <=( (not A167)  and  (not A168) );
 a20200a <=( A169  and  a20199a );
 a20204a <=( (not A201)  and  (not A200) );
 a20205a <=( A166  and  a20204a );
 a20206a <=( a20205a  and  a20200a );
 a20210a <=( A267  and  (not A266) );
 a20211a <=( A265  and  a20210a );
 a20214a <=( A298  and  A269 );
 a20217a <=( (not A302)  and  (not A301) );
 a20218a <=( a20217a  and  a20214a );
 a20219a <=( a20218a  and  a20211a );
 a20223a <=( (not A167)  and  (not A168) );
 a20224a <=( A169  and  a20223a );
 a20228a <=( (not A200)  and  A199 );
 a20229a <=( A166  and  a20228a );
 a20230a <=( a20229a  and  a20224a );
 a20234a <=( (not A266)  and  A202 );
 a20235a <=( A201  and  a20234a );
 a20238a <=( (not A269)  and  (not A268) );
 a20241a <=( A299  and  (not A298) );
 a20242a <=( a20241a  and  a20238a );
 a20243a <=( a20242a  and  a20235a );
 a20247a <=( (not A167)  and  (not A168) );
 a20248a <=( A169  and  a20247a );
 a20252a <=( (not A200)  and  A199 );
 a20253a <=( A166  and  a20252a );
 a20254a <=( a20253a  and  a20248a );
 a20258a <=( (not A266)  and  A203 );
 a20259a <=( A201  and  a20258a );
 a20262a <=( (not A269)  and  (not A268) );
 a20265a <=( A299  and  (not A298) );
 a20266a <=( a20265a  and  a20262a );
 a20267a <=( a20266a  and  a20259a );
 a20271a <=( (not A167)  and  (not A168) );
 a20272a <=( A169  and  a20271a );
 a20276a <=( (not A200)  and  (not A199) );
 a20277a <=( A166  and  a20276a );
 a20278a <=( a20277a  and  a20272a );
 a20282a <=( A267  and  (not A266) );
 a20283a <=( A265  and  a20282a );
 a20286a <=( A298  and  A268 );
 a20289a <=( (not A302)  and  (not A301) );
 a20290a <=( a20289a  and  a20286a );
 a20291a <=( a20290a  and  a20283a );
 a20295a <=( (not A167)  and  (not A168) );
 a20296a <=( A169  and  a20295a );
 a20300a <=( (not A200)  and  (not A199) );
 a20301a <=( A166  and  a20300a );
 a20302a <=( a20301a  and  a20296a );
 a20306a <=( A267  and  (not A266) );
 a20307a <=( A265  and  a20306a );
 a20310a <=( A298  and  A269 );
 a20313a <=( (not A302)  and  (not A301) );
 a20314a <=( a20313a  and  a20310a );
 a20315a <=( a20314a  and  a20307a );
 a20319a <=( (not A168)  and  A169 );
 a20320a <=( A170  and  a20319a );
 a20324a <=( (not A203)  and  (not A202) );
 a20325a <=( (not A200)  and  a20324a );
 a20326a <=( a20325a  and  a20320a );
 a20330a <=( A267  and  (not A266) );
 a20331a <=( A265  and  a20330a );
 a20334a <=( A298  and  A268 );
 a20337a <=( (not A302)  and  (not A301) );
 a20338a <=( a20337a  and  a20334a );
 a20339a <=( a20338a  and  a20331a );
 a20343a <=( (not A168)  and  A169 );
 a20344a <=( A170  and  a20343a );
 a20348a <=( (not A203)  and  (not A202) );
 a20349a <=( (not A200)  and  a20348a );
 a20350a <=( a20349a  and  a20344a );
 a20354a <=( A267  and  (not A266) );
 a20355a <=( A265  and  a20354a );
 a20358a <=( A298  and  A269 );
 a20361a <=( (not A302)  and  (not A301) );
 a20362a <=( a20361a  and  a20358a );
 a20363a <=( a20362a  and  a20355a );
 a20367a <=( (not A168)  and  A169 );
 a20368a <=( A170  and  a20367a );
 a20372a <=( A201  and  (not A200) );
 a20373a <=( A199  and  a20372a );
 a20374a <=( a20373a  and  a20368a );
 a20378a <=( A266  and  A265 );
 a20379a <=( A202  and  a20378a );
 a20382a <=( (not A299)  and  A298 );
 a20385a <=( A301  and  A300 );
 a20386a <=( a20385a  and  a20382a );
 a20387a <=( a20386a  and  a20379a );
 a20391a <=( (not A168)  and  A169 );
 a20392a <=( A170  and  a20391a );
 a20396a <=( A201  and  (not A200) );
 a20397a <=( A199  and  a20396a );
 a20398a <=( a20397a  and  a20392a );
 a20402a <=( A266  and  A265 );
 a20403a <=( A202  and  a20402a );
 a20406a <=( (not A299)  and  A298 );
 a20409a <=( A302  and  A300 );
 a20410a <=( a20409a  and  a20406a );
 a20411a <=( a20410a  and  a20403a );
 a20415a <=( (not A168)  and  A169 );
 a20416a <=( A170  and  a20415a );
 a20420a <=( A201  and  (not A200) );
 a20421a <=( A199  and  a20420a );
 a20422a <=( a20421a  and  a20416a );
 a20426a <=( (not A267)  and  (not A266) );
 a20427a <=( A202  and  a20426a );
 a20430a <=( (not A299)  and  A298 );
 a20433a <=( A301  and  A300 );
 a20434a <=( a20433a  and  a20430a );
 a20435a <=( a20434a  and  a20427a );
 a20439a <=( (not A168)  and  A169 );
 a20440a <=( A170  and  a20439a );
 a20444a <=( A201  and  (not A200) );
 a20445a <=( A199  and  a20444a );
 a20446a <=( a20445a  and  a20440a );
 a20450a <=( (not A267)  and  (not A266) );
 a20451a <=( A202  and  a20450a );
 a20454a <=( (not A299)  and  A298 );
 a20457a <=( A302  and  A300 );
 a20458a <=( a20457a  and  a20454a );
 a20459a <=( a20458a  and  a20451a );
 a20463a <=( (not A168)  and  A169 );
 a20464a <=( A170  and  a20463a );
 a20468a <=( A201  and  (not A200) );
 a20469a <=( A199  and  a20468a );
 a20470a <=( a20469a  and  a20464a );
 a20474a <=( (not A266)  and  (not A265) );
 a20475a <=( A202  and  a20474a );
 a20478a <=( (not A299)  and  A298 );
 a20481a <=( A301  and  A300 );
 a20482a <=( a20481a  and  a20478a );
 a20483a <=( a20482a  and  a20475a );
 a20487a <=( (not A168)  and  A169 );
 a20488a <=( A170  and  a20487a );
 a20492a <=( A201  and  (not A200) );
 a20493a <=( A199  and  a20492a );
 a20494a <=( a20493a  and  a20488a );
 a20498a <=( (not A266)  and  (not A265) );
 a20499a <=( A202  and  a20498a );
 a20502a <=( (not A299)  and  A298 );
 a20505a <=( A302  and  A300 );
 a20506a <=( a20505a  and  a20502a );
 a20507a <=( a20506a  and  a20499a );
 a20511a <=( (not A168)  and  A169 );
 a20512a <=( A170  and  a20511a );
 a20516a <=( A201  and  (not A200) );
 a20517a <=( A199  and  a20516a );
 a20518a <=( a20517a  and  a20512a );
 a20522a <=( A266  and  A265 );
 a20523a <=( A203  and  a20522a );
 a20526a <=( (not A299)  and  A298 );
 a20529a <=( A301  and  A300 );
 a20530a <=( a20529a  and  a20526a );
 a20531a <=( a20530a  and  a20523a );
 a20535a <=( (not A168)  and  A169 );
 a20536a <=( A170  and  a20535a );
 a20540a <=( A201  and  (not A200) );
 a20541a <=( A199  and  a20540a );
 a20542a <=( a20541a  and  a20536a );
 a20546a <=( A266  and  A265 );
 a20547a <=( A203  and  a20546a );
 a20550a <=( (not A299)  and  A298 );
 a20553a <=( A302  and  A300 );
 a20554a <=( a20553a  and  a20550a );
 a20555a <=( a20554a  and  a20547a );
 a20559a <=( (not A168)  and  A169 );
 a20560a <=( A170  and  a20559a );
 a20564a <=( A201  and  (not A200) );
 a20565a <=( A199  and  a20564a );
 a20566a <=( a20565a  and  a20560a );
 a20570a <=( (not A267)  and  (not A266) );
 a20571a <=( A203  and  a20570a );
 a20574a <=( (not A299)  and  A298 );
 a20577a <=( A301  and  A300 );
 a20578a <=( a20577a  and  a20574a );
 a20579a <=( a20578a  and  a20571a );
 a20583a <=( (not A168)  and  A169 );
 a20584a <=( A170  and  a20583a );
 a20588a <=( A201  and  (not A200) );
 a20589a <=( A199  and  a20588a );
 a20590a <=( a20589a  and  a20584a );
 a20594a <=( (not A267)  and  (not A266) );
 a20595a <=( A203  and  a20594a );
 a20598a <=( (not A299)  and  A298 );
 a20601a <=( A302  and  A300 );
 a20602a <=( a20601a  and  a20598a );
 a20603a <=( a20602a  and  a20595a );
 a20607a <=( (not A168)  and  A169 );
 a20608a <=( A170  and  a20607a );
 a20612a <=( A201  and  (not A200) );
 a20613a <=( A199  and  a20612a );
 a20614a <=( a20613a  and  a20608a );
 a20618a <=( (not A266)  and  (not A265) );
 a20619a <=( A203  and  a20618a );
 a20622a <=( (not A299)  and  A298 );
 a20625a <=( A301  and  A300 );
 a20626a <=( a20625a  and  a20622a );
 a20627a <=( a20626a  and  a20619a );
 a20631a <=( (not A168)  and  A169 );
 a20632a <=( A170  and  a20631a );
 a20636a <=( A201  and  (not A200) );
 a20637a <=( A199  and  a20636a );
 a20638a <=( a20637a  and  a20632a );
 a20642a <=( (not A266)  and  (not A265) );
 a20643a <=( A203  and  a20642a );
 a20646a <=( (not A299)  and  A298 );
 a20649a <=( A302  and  A300 );
 a20650a <=( a20649a  and  a20646a );
 a20651a <=( a20650a  and  a20643a );
 a20655a <=( A167  and  A169 );
 a20656a <=( (not A170)  and  a20655a );
 a20660a <=( A200  and  A199 );
 a20661a <=( A166  and  a20660a );
 a20662a <=( a20661a  and  a20656a );
 a20666a <=( (not A269)  and  (not A268) );
 a20667a <=( (not A266)  and  a20666a );
 a20670a <=( (not A299)  and  A298 );
 a20673a <=( A301  and  A300 );
 a20674a <=( a20673a  and  a20670a );
 a20675a <=( a20674a  and  a20667a );
 a20679a <=( A167  and  A169 );
 a20680a <=( (not A170)  and  a20679a );
 a20684a <=( A200  and  A199 );
 a20685a <=( A166  and  a20684a );
 a20686a <=( a20685a  and  a20680a );
 a20690a <=( (not A269)  and  (not A268) );
 a20691a <=( (not A266)  and  a20690a );
 a20694a <=( (not A299)  and  A298 );
 a20697a <=( A302  and  A300 );
 a20698a <=( a20697a  and  a20694a );
 a20699a <=( a20698a  and  a20691a );
 a20703a <=( A167  and  A169 );
 a20704a <=( (not A170)  and  a20703a );
 a20708a <=( A200  and  (not A199) );
 a20709a <=( A166  and  a20708a );
 a20710a <=( a20709a  and  a20704a );
 a20714a <=( A267  and  (not A266) );
 a20715a <=( A265  and  a20714a );
 a20718a <=( A298  and  A268 );
 a20721a <=( (not A302)  and  (not A301) );
 a20722a <=( a20721a  and  a20718a );
 a20723a <=( a20722a  and  a20715a );
 a20727a <=( A167  and  A169 );
 a20728a <=( (not A170)  and  a20727a );
 a20732a <=( A200  and  (not A199) );
 a20733a <=( A166  and  a20732a );
 a20734a <=( a20733a  and  a20728a );
 a20738a <=( A267  and  (not A266) );
 a20739a <=( A265  and  a20738a );
 a20742a <=( A298  and  A269 );
 a20745a <=( (not A302)  and  (not A301) );
 a20746a <=( a20745a  and  a20742a );
 a20747a <=( a20746a  and  a20739a );
 a20751a <=( A167  and  A169 );
 a20752a <=( (not A170)  and  a20751a );
 a20756a <=( (not A202)  and  (not A200) );
 a20757a <=( A166  and  a20756a );
 a20758a <=( a20757a  and  a20752a );
 a20762a <=( A266  and  A265 );
 a20763a <=( (not A203)  and  a20762a );
 a20766a <=( (not A299)  and  A298 );
 a20769a <=( A301  and  A300 );
 a20770a <=( a20769a  and  a20766a );
 a20771a <=( a20770a  and  a20763a );
 a20775a <=( A167  and  A169 );
 a20776a <=( (not A170)  and  a20775a );
 a20780a <=( (not A202)  and  (not A200) );
 a20781a <=( A166  and  a20780a );
 a20782a <=( a20781a  and  a20776a );
 a20786a <=( A266  and  A265 );
 a20787a <=( (not A203)  and  a20786a );
 a20790a <=( (not A299)  and  A298 );
 a20793a <=( A302  and  A300 );
 a20794a <=( a20793a  and  a20790a );
 a20795a <=( a20794a  and  a20787a );
 a20799a <=( A167  and  A169 );
 a20800a <=( (not A170)  and  a20799a );
 a20804a <=( (not A202)  and  (not A200) );
 a20805a <=( A166  and  a20804a );
 a20806a <=( a20805a  and  a20800a );
 a20810a <=( (not A267)  and  (not A266) );
 a20811a <=( (not A203)  and  a20810a );
 a20814a <=( (not A299)  and  A298 );
 a20817a <=( A301  and  A300 );
 a20818a <=( a20817a  and  a20814a );
 a20819a <=( a20818a  and  a20811a );
 a20823a <=( A167  and  A169 );
 a20824a <=( (not A170)  and  a20823a );
 a20828a <=( (not A202)  and  (not A200) );
 a20829a <=( A166  and  a20828a );
 a20830a <=( a20829a  and  a20824a );
 a20834a <=( (not A267)  and  (not A266) );
 a20835a <=( (not A203)  and  a20834a );
 a20838a <=( (not A299)  and  A298 );
 a20841a <=( A302  and  A300 );
 a20842a <=( a20841a  and  a20838a );
 a20843a <=( a20842a  and  a20835a );
 a20847a <=( A167  and  A169 );
 a20848a <=( (not A170)  and  a20847a );
 a20852a <=( (not A202)  and  (not A200) );
 a20853a <=( A166  and  a20852a );
 a20854a <=( a20853a  and  a20848a );
 a20858a <=( (not A266)  and  (not A265) );
 a20859a <=( (not A203)  and  a20858a );
 a20862a <=( (not A299)  and  A298 );
 a20865a <=( A301  and  A300 );
 a20866a <=( a20865a  and  a20862a );
 a20867a <=( a20866a  and  a20859a );
 a20871a <=( A167  and  A169 );
 a20872a <=( (not A170)  and  a20871a );
 a20876a <=( (not A202)  and  (not A200) );
 a20877a <=( A166  and  a20876a );
 a20878a <=( a20877a  and  a20872a );
 a20882a <=( (not A266)  and  (not A265) );
 a20883a <=( (not A203)  and  a20882a );
 a20886a <=( (not A299)  and  A298 );
 a20889a <=( A302  and  A300 );
 a20890a <=( a20889a  and  a20886a );
 a20891a <=( a20890a  and  a20883a );
 a20895a <=( A167  and  A169 );
 a20896a <=( (not A170)  and  a20895a );
 a20900a <=( (not A201)  and  (not A200) );
 a20901a <=( A166  and  a20900a );
 a20902a <=( a20901a  and  a20896a );
 a20906a <=( (not A269)  and  (not A268) );
 a20907a <=( (not A266)  and  a20906a );
 a20910a <=( (not A299)  and  A298 );
 a20913a <=( A301  and  A300 );
 a20914a <=( a20913a  and  a20910a );
 a20915a <=( a20914a  and  a20907a );
 a20919a <=( A167  and  A169 );
 a20920a <=( (not A170)  and  a20919a );
 a20924a <=( (not A201)  and  (not A200) );
 a20925a <=( A166  and  a20924a );
 a20926a <=( a20925a  and  a20920a );
 a20930a <=( (not A269)  and  (not A268) );
 a20931a <=( (not A266)  and  a20930a );
 a20934a <=( (not A299)  and  A298 );
 a20937a <=( A302  and  A300 );
 a20938a <=( a20937a  and  a20934a );
 a20939a <=( a20938a  and  a20931a );
 a20943a <=( A167  and  A169 );
 a20944a <=( (not A170)  and  a20943a );
 a20948a <=( (not A200)  and  A199 );
 a20949a <=( A166  and  a20948a );
 a20950a <=( a20949a  and  a20944a );
 a20954a <=( (not A265)  and  A202 );
 a20955a <=( A201  and  a20954a );
 a20958a <=( A298  and  A266 );
 a20961a <=( (not A302)  and  (not A301) );
 a20962a <=( a20961a  and  a20958a );
 a20963a <=( a20962a  and  a20955a );
 a20967a <=( A167  and  A169 );
 a20968a <=( (not A170)  and  a20967a );
 a20972a <=( (not A200)  and  A199 );
 a20973a <=( A166  and  a20972a );
 a20974a <=( a20973a  and  a20968a );
 a20978a <=( (not A265)  and  A203 );
 a20979a <=( A201  and  a20978a );
 a20982a <=( A298  and  A266 );
 a20985a <=( (not A302)  and  (not A301) );
 a20986a <=( a20985a  and  a20982a );
 a20987a <=( a20986a  and  a20979a );
 a20991a <=( A167  and  A169 );
 a20992a <=( (not A170)  and  a20991a );
 a20996a <=( (not A200)  and  (not A199) );
 a20997a <=( A166  and  a20996a );
 a20998a <=( a20997a  and  a20992a );
 a21002a <=( (not A269)  and  (not A268) );
 a21003a <=( (not A266)  and  a21002a );
 a21006a <=( (not A299)  and  A298 );
 a21009a <=( A301  and  A300 );
 a21010a <=( a21009a  and  a21006a );
 a21011a <=( a21010a  and  a21003a );
 a21015a <=( A167  and  A169 );
 a21016a <=( (not A170)  and  a21015a );
 a21020a <=( (not A200)  and  (not A199) );
 a21021a <=( A166  and  a21020a );
 a21022a <=( a21021a  and  a21016a );
 a21026a <=( (not A269)  and  (not A268) );
 a21027a <=( (not A266)  and  a21026a );
 a21030a <=( (not A299)  and  A298 );
 a21033a <=( A302  and  A300 );
 a21034a <=( a21033a  and  a21030a );
 a21035a <=( a21034a  and  a21027a );
 a21039a <=( (not A167)  and  A169 );
 a21040a <=( (not A170)  and  a21039a );
 a21044a <=( A200  and  A199 );
 a21045a <=( (not A166)  and  a21044a );
 a21046a <=( a21045a  and  a21040a );
 a21050a <=( (not A269)  and  (not A268) );
 a21051a <=( (not A266)  and  a21050a );
 a21054a <=( (not A299)  and  A298 );
 a21057a <=( A301  and  A300 );
 a21058a <=( a21057a  and  a21054a );
 a21059a <=( a21058a  and  a21051a );
 a21063a <=( (not A167)  and  A169 );
 a21064a <=( (not A170)  and  a21063a );
 a21068a <=( A200  and  A199 );
 a21069a <=( (not A166)  and  a21068a );
 a21070a <=( a21069a  and  a21064a );
 a21074a <=( (not A269)  and  (not A268) );
 a21075a <=( (not A266)  and  a21074a );
 a21078a <=( (not A299)  and  A298 );
 a21081a <=( A302  and  A300 );
 a21082a <=( a21081a  and  a21078a );
 a21083a <=( a21082a  and  a21075a );
 a21087a <=( (not A167)  and  A169 );
 a21088a <=( (not A170)  and  a21087a );
 a21092a <=( A200  and  (not A199) );
 a21093a <=( (not A166)  and  a21092a );
 a21094a <=( a21093a  and  a21088a );
 a21098a <=( A267  and  (not A266) );
 a21099a <=( A265  and  a21098a );
 a21102a <=( A298  and  A268 );
 a21105a <=( (not A302)  and  (not A301) );
 a21106a <=( a21105a  and  a21102a );
 a21107a <=( a21106a  and  a21099a );
 a21111a <=( (not A167)  and  A169 );
 a21112a <=( (not A170)  and  a21111a );
 a21116a <=( A200  and  (not A199) );
 a21117a <=( (not A166)  and  a21116a );
 a21118a <=( a21117a  and  a21112a );
 a21122a <=( A267  and  (not A266) );
 a21123a <=( A265  and  a21122a );
 a21126a <=( A298  and  A269 );
 a21129a <=( (not A302)  and  (not A301) );
 a21130a <=( a21129a  and  a21126a );
 a21131a <=( a21130a  and  a21123a );
 a21135a <=( (not A167)  and  A169 );
 a21136a <=( (not A170)  and  a21135a );
 a21140a <=( (not A202)  and  (not A200) );
 a21141a <=( (not A166)  and  a21140a );
 a21142a <=( a21141a  and  a21136a );
 a21146a <=( A266  and  A265 );
 a21147a <=( (not A203)  and  a21146a );
 a21150a <=( (not A299)  and  A298 );
 a21153a <=( A301  and  A300 );
 a21154a <=( a21153a  and  a21150a );
 a21155a <=( a21154a  and  a21147a );
 a21159a <=( (not A167)  and  A169 );
 a21160a <=( (not A170)  and  a21159a );
 a21164a <=( (not A202)  and  (not A200) );
 a21165a <=( (not A166)  and  a21164a );
 a21166a <=( a21165a  and  a21160a );
 a21170a <=( A266  and  A265 );
 a21171a <=( (not A203)  and  a21170a );
 a21174a <=( (not A299)  and  A298 );
 a21177a <=( A302  and  A300 );
 a21178a <=( a21177a  and  a21174a );
 a21179a <=( a21178a  and  a21171a );
 a21183a <=( (not A167)  and  A169 );
 a21184a <=( (not A170)  and  a21183a );
 a21188a <=( (not A202)  and  (not A200) );
 a21189a <=( (not A166)  and  a21188a );
 a21190a <=( a21189a  and  a21184a );
 a21194a <=( (not A267)  and  (not A266) );
 a21195a <=( (not A203)  and  a21194a );
 a21198a <=( (not A299)  and  A298 );
 a21201a <=( A301  and  A300 );
 a21202a <=( a21201a  and  a21198a );
 a21203a <=( a21202a  and  a21195a );
 a21207a <=( (not A167)  and  A169 );
 a21208a <=( (not A170)  and  a21207a );
 a21212a <=( (not A202)  and  (not A200) );
 a21213a <=( (not A166)  and  a21212a );
 a21214a <=( a21213a  and  a21208a );
 a21218a <=( (not A267)  and  (not A266) );
 a21219a <=( (not A203)  and  a21218a );
 a21222a <=( (not A299)  and  A298 );
 a21225a <=( A302  and  A300 );
 a21226a <=( a21225a  and  a21222a );
 a21227a <=( a21226a  and  a21219a );
 a21231a <=( (not A167)  and  A169 );
 a21232a <=( (not A170)  and  a21231a );
 a21236a <=( (not A202)  and  (not A200) );
 a21237a <=( (not A166)  and  a21236a );
 a21238a <=( a21237a  and  a21232a );
 a21242a <=( (not A266)  and  (not A265) );
 a21243a <=( (not A203)  and  a21242a );
 a21246a <=( (not A299)  and  A298 );
 a21249a <=( A301  and  A300 );
 a21250a <=( a21249a  and  a21246a );
 a21251a <=( a21250a  and  a21243a );
 a21255a <=( (not A167)  and  A169 );
 a21256a <=( (not A170)  and  a21255a );
 a21260a <=( (not A202)  and  (not A200) );
 a21261a <=( (not A166)  and  a21260a );
 a21262a <=( a21261a  and  a21256a );
 a21266a <=( (not A266)  and  (not A265) );
 a21267a <=( (not A203)  and  a21266a );
 a21270a <=( (not A299)  and  A298 );
 a21273a <=( A302  and  A300 );
 a21274a <=( a21273a  and  a21270a );
 a21275a <=( a21274a  and  a21267a );
 a21279a <=( (not A167)  and  A169 );
 a21280a <=( (not A170)  and  a21279a );
 a21284a <=( (not A201)  and  (not A200) );
 a21285a <=( (not A166)  and  a21284a );
 a21286a <=( a21285a  and  a21280a );
 a21290a <=( (not A269)  and  (not A268) );
 a21291a <=( (not A266)  and  a21290a );
 a21294a <=( (not A299)  and  A298 );
 a21297a <=( A301  and  A300 );
 a21298a <=( a21297a  and  a21294a );
 a21299a <=( a21298a  and  a21291a );
 a21303a <=( (not A167)  and  A169 );
 a21304a <=( (not A170)  and  a21303a );
 a21308a <=( (not A201)  and  (not A200) );
 a21309a <=( (not A166)  and  a21308a );
 a21310a <=( a21309a  and  a21304a );
 a21314a <=( (not A269)  and  (not A268) );
 a21315a <=( (not A266)  and  a21314a );
 a21318a <=( (not A299)  and  A298 );
 a21321a <=( A302  and  A300 );
 a21322a <=( a21321a  and  a21318a );
 a21323a <=( a21322a  and  a21315a );
 a21327a <=( (not A167)  and  A169 );
 a21328a <=( (not A170)  and  a21327a );
 a21332a <=( (not A200)  and  A199 );
 a21333a <=( (not A166)  and  a21332a );
 a21334a <=( a21333a  and  a21328a );
 a21338a <=( (not A265)  and  A202 );
 a21339a <=( A201  and  a21338a );
 a21342a <=( A298  and  A266 );
 a21345a <=( (not A302)  and  (not A301) );
 a21346a <=( a21345a  and  a21342a );
 a21347a <=( a21346a  and  a21339a );
 a21351a <=( (not A167)  and  A169 );
 a21352a <=( (not A170)  and  a21351a );
 a21356a <=( (not A200)  and  A199 );
 a21357a <=( (not A166)  and  a21356a );
 a21358a <=( a21357a  and  a21352a );
 a21362a <=( (not A265)  and  A203 );
 a21363a <=( A201  and  a21362a );
 a21366a <=( A298  and  A266 );
 a21369a <=( (not A302)  and  (not A301) );
 a21370a <=( a21369a  and  a21366a );
 a21371a <=( a21370a  and  a21363a );
 a21375a <=( (not A167)  and  A169 );
 a21376a <=( (not A170)  and  a21375a );
 a21380a <=( (not A200)  and  (not A199) );
 a21381a <=( (not A166)  and  a21380a );
 a21382a <=( a21381a  and  a21376a );
 a21386a <=( (not A269)  and  (not A268) );
 a21387a <=( (not A266)  and  a21386a );
 a21390a <=( (not A299)  and  A298 );
 a21393a <=( A301  and  A300 );
 a21394a <=( a21393a  and  a21390a );
 a21395a <=( a21394a  and  a21387a );
 a21399a <=( (not A167)  and  A169 );
 a21400a <=( (not A170)  and  a21399a );
 a21404a <=( (not A200)  and  (not A199) );
 a21405a <=( (not A166)  and  a21404a );
 a21406a <=( a21405a  and  a21400a );
 a21410a <=( (not A269)  and  (not A268) );
 a21411a <=( (not A266)  and  a21410a );
 a21414a <=( (not A299)  and  A298 );
 a21417a <=( A302  and  A300 );
 a21418a <=( a21417a  and  a21414a );
 a21419a <=( a21418a  and  a21411a );
 a21423a <=( (not A166)  and  (not A167) );
 a21424a <=( (not A169)  and  a21423a );
 a21428a <=( (not A203)  and  (not A202) );
 a21429a <=( (not A200)  and  a21428a );
 a21430a <=( a21429a  and  a21424a );
 a21434a <=( A267  and  (not A266) );
 a21435a <=( A265  and  a21434a );
 a21438a <=( A298  and  A268 );
 a21441a <=( (not A302)  and  (not A301) );
 a21442a <=( a21441a  and  a21438a );
 a21443a <=( a21442a  and  a21435a );
 a21447a <=( (not A166)  and  (not A167) );
 a21448a <=( (not A169)  and  a21447a );
 a21452a <=( (not A203)  and  (not A202) );
 a21453a <=( (not A200)  and  a21452a );
 a21454a <=( a21453a  and  a21448a );
 a21458a <=( A267  and  (not A266) );
 a21459a <=( A265  and  a21458a );
 a21462a <=( A298  and  A269 );
 a21465a <=( (not A302)  and  (not A301) );
 a21466a <=( a21465a  and  a21462a );
 a21467a <=( a21466a  and  a21459a );
 a21471a <=( (not A166)  and  (not A167) );
 a21472a <=( (not A169)  and  a21471a );
 a21476a <=( A201  and  (not A200) );
 a21477a <=( A199  and  a21476a );
 a21478a <=( a21477a  and  a21472a );
 a21482a <=( A266  and  A265 );
 a21483a <=( A202  and  a21482a );
 a21486a <=( (not A299)  and  A298 );
 a21489a <=( A301  and  A300 );
 a21490a <=( a21489a  and  a21486a );
 a21491a <=( a21490a  and  a21483a );
 a21495a <=( (not A166)  and  (not A167) );
 a21496a <=( (not A169)  and  a21495a );
 a21500a <=( A201  and  (not A200) );
 a21501a <=( A199  and  a21500a );
 a21502a <=( a21501a  and  a21496a );
 a21506a <=( A266  and  A265 );
 a21507a <=( A202  and  a21506a );
 a21510a <=( (not A299)  and  A298 );
 a21513a <=( A302  and  A300 );
 a21514a <=( a21513a  and  a21510a );
 a21515a <=( a21514a  and  a21507a );
 a21519a <=( (not A166)  and  (not A167) );
 a21520a <=( (not A169)  and  a21519a );
 a21524a <=( A201  and  (not A200) );
 a21525a <=( A199  and  a21524a );
 a21526a <=( a21525a  and  a21520a );
 a21530a <=( (not A267)  and  (not A266) );
 a21531a <=( A202  and  a21530a );
 a21534a <=( (not A299)  and  A298 );
 a21537a <=( A301  and  A300 );
 a21538a <=( a21537a  and  a21534a );
 a21539a <=( a21538a  and  a21531a );
 a21543a <=( (not A166)  and  (not A167) );
 a21544a <=( (not A169)  and  a21543a );
 a21548a <=( A201  and  (not A200) );
 a21549a <=( A199  and  a21548a );
 a21550a <=( a21549a  and  a21544a );
 a21554a <=( (not A267)  and  (not A266) );
 a21555a <=( A202  and  a21554a );
 a21558a <=( (not A299)  and  A298 );
 a21561a <=( A302  and  A300 );
 a21562a <=( a21561a  and  a21558a );
 a21563a <=( a21562a  and  a21555a );
 a21567a <=( (not A166)  and  (not A167) );
 a21568a <=( (not A169)  and  a21567a );
 a21572a <=( A201  and  (not A200) );
 a21573a <=( A199  and  a21572a );
 a21574a <=( a21573a  and  a21568a );
 a21578a <=( (not A266)  and  (not A265) );
 a21579a <=( A202  and  a21578a );
 a21582a <=( (not A299)  and  A298 );
 a21585a <=( A301  and  A300 );
 a21586a <=( a21585a  and  a21582a );
 a21587a <=( a21586a  and  a21579a );
 a21591a <=( (not A166)  and  (not A167) );
 a21592a <=( (not A169)  and  a21591a );
 a21596a <=( A201  and  (not A200) );
 a21597a <=( A199  and  a21596a );
 a21598a <=( a21597a  and  a21592a );
 a21602a <=( (not A266)  and  (not A265) );
 a21603a <=( A202  and  a21602a );
 a21606a <=( (not A299)  and  A298 );
 a21609a <=( A302  and  A300 );
 a21610a <=( a21609a  and  a21606a );
 a21611a <=( a21610a  and  a21603a );
 a21615a <=( (not A166)  and  (not A167) );
 a21616a <=( (not A169)  and  a21615a );
 a21620a <=( A201  and  (not A200) );
 a21621a <=( A199  and  a21620a );
 a21622a <=( a21621a  and  a21616a );
 a21626a <=( A266  and  A265 );
 a21627a <=( A203  and  a21626a );
 a21630a <=( (not A299)  and  A298 );
 a21633a <=( A301  and  A300 );
 a21634a <=( a21633a  and  a21630a );
 a21635a <=( a21634a  and  a21627a );
 a21639a <=( (not A166)  and  (not A167) );
 a21640a <=( (not A169)  and  a21639a );
 a21644a <=( A201  and  (not A200) );
 a21645a <=( A199  and  a21644a );
 a21646a <=( a21645a  and  a21640a );
 a21650a <=( A266  and  A265 );
 a21651a <=( A203  and  a21650a );
 a21654a <=( (not A299)  and  A298 );
 a21657a <=( A302  and  A300 );
 a21658a <=( a21657a  and  a21654a );
 a21659a <=( a21658a  and  a21651a );
 a21663a <=( (not A166)  and  (not A167) );
 a21664a <=( (not A169)  and  a21663a );
 a21668a <=( A201  and  (not A200) );
 a21669a <=( A199  and  a21668a );
 a21670a <=( a21669a  and  a21664a );
 a21674a <=( (not A267)  and  (not A266) );
 a21675a <=( A203  and  a21674a );
 a21678a <=( (not A299)  and  A298 );
 a21681a <=( A301  and  A300 );
 a21682a <=( a21681a  and  a21678a );
 a21683a <=( a21682a  and  a21675a );
 a21687a <=( (not A166)  and  (not A167) );
 a21688a <=( (not A169)  and  a21687a );
 a21692a <=( A201  and  (not A200) );
 a21693a <=( A199  and  a21692a );
 a21694a <=( a21693a  and  a21688a );
 a21698a <=( (not A267)  and  (not A266) );
 a21699a <=( A203  and  a21698a );
 a21702a <=( (not A299)  and  A298 );
 a21705a <=( A302  and  A300 );
 a21706a <=( a21705a  and  a21702a );
 a21707a <=( a21706a  and  a21699a );
 a21711a <=( (not A166)  and  (not A167) );
 a21712a <=( (not A169)  and  a21711a );
 a21716a <=( A201  and  (not A200) );
 a21717a <=( A199  and  a21716a );
 a21718a <=( a21717a  and  a21712a );
 a21722a <=( (not A266)  and  (not A265) );
 a21723a <=( A203  and  a21722a );
 a21726a <=( (not A299)  and  A298 );
 a21729a <=( A301  and  A300 );
 a21730a <=( a21729a  and  a21726a );
 a21731a <=( a21730a  and  a21723a );
 a21735a <=( (not A166)  and  (not A167) );
 a21736a <=( (not A169)  and  a21735a );
 a21740a <=( A201  and  (not A200) );
 a21741a <=( A199  and  a21740a );
 a21742a <=( a21741a  and  a21736a );
 a21746a <=( (not A266)  and  (not A265) );
 a21747a <=( A203  and  a21746a );
 a21750a <=( (not A299)  and  A298 );
 a21753a <=( A302  and  A300 );
 a21754a <=( a21753a  and  a21750a );
 a21755a <=( a21754a  and  a21747a );
 a21759a <=( A167  and  (not A168) );
 a21760a <=( (not A169)  and  a21759a );
 a21764a <=( A200  and  A199 );
 a21765a <=( A166  and  a21764a );
 a21766a <=( a21765a  and  a21760a );
 a21770a <=( A267  and  (not A266) );
 a21771a <=( A265  and  a21770a );
 a21774a <=( A298  and  A268 );
 a21777a <=( (not A302)  and  (not A301) );
 a21778a <=( a21777a  and  a21774a );
 a21779a <=( a21778a  and  a21771a );
 a21783a <=( A167  and  (not A168) );
 a21784a <=( (not A169)  and  a21783a );
 a21788a <=( A200  and  A199 );
 a21789a <=( A166  and  a21788a );
 a21790a <=( a21789a  and  a21784a );
 a21794a <=( A267  and  (not A266) );
 a21795a <=( A265  and  a21794a );
 a21798a <=( A298  and  A269 );
 a21801a <=( (not A302)  and  (not A301) );
 a21802a <=( a21801a  and  a21798a );
 a21803a <=( a21802a  and  a21795a );
 a21807a <=( A167  and  (not A168) );
 a21808a <=( (not A169)  and  a21807a );
 a21812a <=( A200  and  (not A199) );
 a21813a <=( A166  and  a21812a );
 a21814a <=( a21813a  and  a21808a );
 a21818a <=( (not A269)  and  (not A268) );
 a21819a <=( (not A266)  and  a21818a );
 a21822a <=( (not A299)  and  A298 );
 a21825a <=( A301  and  A300 );
 a21826a <=( a21825a  and  a21822a );
 a21827a <=( a21826a  and  a21819a );
 a21831a <=( A167  and  (not A168) );
 a21832a <=( (not A169)  and  a21831a );
 a21836a <=( A200  and  (not A199) );
 a21837a <=( A166  and  a21836a );
 a21838a <=( a21837a  and  a21832a );
 a21842a <=( (not A269)  and  (not A268) );
 a21843a <=( (not A266)  and  a21842a );
 a21846a <=( (not A299)  and  A298 );
 a21849a <=( A302  and  A300 );
 a21850a <=( a21849a  and  a21846a );
 a21851a <=( a21850a  and  a21843a );
 a21855a <=( A167  and  (not A168) );
 a21856a <=( (not A169)  and  a21855a );
 a21860a <=( (not A202)  and  (not A200) );
 a21861a <=( A166  and  a21860a );
 a21862a <=( a21861a  and  a21856a );
 a21866a <=( (not A266)  and  A265 );
 a21867a <=( (not A203)  and  a21866a );
 a21870a <=( A268  and  A267 );
 a21873a <=( (not A300)  and  A298 );
 a21874a <=( a21873a  and  a21870a );
 a21875a <=( a21874a  and  a21867a );
 a21879a <=( A167  and  (not A168) );
 a21880a <=( (not A169)  and  a21879a );
 a21884a <=( (not A202)  and  (not A200) );
 a21885a <=( A166  and  a21884a );
 a21886a <=( a21885a  and  a21880a );
 a21890a <=( (not A266)  and  A265 );
 a21891a <=( (not A203)  and  a21890a );
 a21894a <=( A268  and  A267 );
 a21897a <=( A299  and  A298 );
 a21898a <=( a21897a  and  a21894a );
 a21899a <=( a21898a  and  a21891a );
 a21903a <=( A167  and  (not A168) );
 a21904a <=( (not A169)  and  a21903a );
 a21908a <=( (not A202)  and  (not A200) );
 a21909a <=( A166  and  a21908a );
 a21910a <=( a21909a  and  a21904a );
 a21914a <=( (not A266)  and  A265 );
 a21915a <=( (not A203)  and  a21914a );
 a21918a <=( A268  and  A267 );
 a21921a <=( (not A299)  and  (not A298) );
 a21922a <=( a21921a  and  a21918a );
 a21923a <=( a21922a  and  a21915a );
 a21927a <=( A167  and  (not A168) );
 a21928a <=( (not A169)  and  a21927a );
 a21932a <=( (not A202)  and  (not A200) );
 a21933a <=( A166  and  a21932a );
 a21934a <=( a21933a  and  a21928a );
 a21938a <=( (not A266)  and  A265 );
 a21939a <=( (not A203)  and  a21938a );
 a21942a <=( A269  and  A267 );
 a21945a <=( (not A300)  and  A298 );
 a21946a <=( a21945a  and  a21942a );
 a21947a <=( a21946a  and  a21939a );
 a21951a <=( A167  and  (not A168) );
 a21952a <=( (not A169)  and  a21951a );
 a21956a <=( (not A202)  and  (not A200) );
 a21957a <=( A166  and  a21956a );
 a21958a <=( a21957a  and  a21952a );
 a21962a <=( (not A266)  and  A265 );
 a21963a <=( (not A203)  and  a21962a );
 a21966a <=( A269  and  A267 );
 a21969a <=( A299  and  A298 );
 a21970a <=( a21969a  and  a21966a );
 a21971a <=( a21970a  and  a21963a );
 a21975a <=( A167  and  (not A168) );
 a21976a <=( (not A169)  and  a21975a );
 a21980a <=( (not A202)  and  (not A200) );
 a21981a <=( A166  and  a21980a );
 a21982a <=( a21981a  and  a21976a );
 a21986a <=( (not A266)  and  A265 );
 a21987a <=( (not A203)  and  a21986a );
 a21990a <=( A269  and  A267 );
 a21993a <=( (not A299)  and  (not A298) );
 a21994a <=( a21993a  and  a21990a );
 a21995a <=( a21994a  and  a21987a );
 a21999a <=( A167  and  (not A168) );
 a22000a <=( (not A169)  and  a21999a );
 a22004a <=( (not A201)  and  (not A200) );
 a22005a <=( A166  and  a22004a );
 a22006a <=( a22005a  and  a22000a );
 a22010a <=( A267  and  (not A266) );
 a22011a <=( A265  and  a22010a );
 a22014a <=( A298  and  A268 );
 a22017a <=( (not A302)  and  (not A301) );
 a22018a <=( a22017a  and  a22014a );
 a22019a <=( a22018a  and  a22011a );
 a22023a <=( A167  and  (not A168) );
 a22024a <=( (not A169)  and  a22023a );
 a22028a <=( (not A201)  and  (not A200) );
 a22029a <=( A166  and  a22028a );
 a22030a <=( a22029a  and  a22024a );
 a22034a <=( A267  and  (not A266) );
 a22035a <=( A265  and  a22034a );
 a22038a <=( A298  and  A269 );
 a22041a <=( (not A302)  and  (not A301) );
 a22042a <=( a22041a  and  a22038a );
 a22043a <=( a22042a  and  a22035a );
 a22047a <=( A167  and  (not A168) );
 a22048a <=( (not A169)  and  a22047a );
 a22052a <=( (not A200)  and  A199 );
 a22053a <=( A166  and  a22052a );
 a22054a <=( a22053a  and  a22048a );
 a22058a <=( (not A266)  and  A202 );
 a22059a <=( A201  and  a22058a );
 a22062a <=( (not A269)  and  (not A268) );
 a22065a <=( A299  and  (not A298) );
 a22066a <=( a22065a  and  a22062a );
 a22067a <=( a22066a  and  a22059a );
 a22071a <=( A167  and  (not A168) );
 a22072a <=( (not A169)  and  a22071a );
 a22076a <=( (not A200)  and  A199 );
 a22077a <=( A166  and  a22076a );
 a22078a <=( a22077a  and  a22072a );
 a22082a <=( (not A266)  and  A203 );
 a22083a <=( A201  and  a22082a );
 a22086a <=( (not A269)  and  (not A268) );
 a22089a <=( A299  and  (not A298) );
 a22090a <=( a22089a  and  a22086a );
 a22091a <=( a22090a  and  a22083a );
 a22095a <=( A167  and  (not A168) );
 a22096a <=( (not A169)  and  a22095a );
 a22100a <=( (not A200)  and  (not A199) );
 a22101a <=( A166  and  a22100a );
 a22102a <=( a22101a  and  a22096a );
 a22106a <=( A267  and  (not A266) );
 a22107a <=( A265  and  a22106a );
 a22110a <=( A298  and  A268 );
 a22113a <=( (not A302)  and  (not A301) );
 a22114a <=( a22113a  and  a22110a );
 a22115a <=( a22114a  and  a22107a );
 a22119a <=( A167  and  (not A168) );
 a22120a <=( (not A169)  and  a22119a );
 a22124a <=( (not A200)  and  (not A199) );
 a22125a <=( A166  and  a22124a );
 a22126a <=( a22125a  and  a22120a );
 a22130a <=( A267  and  (not A266) );
 a22131a <=( A265  and  a22130a );
 a22134a <=( A298  and  A269 );
 a22137a <=( (not A302)  and  (not A301) );
 a22138a <=( a22137a  and  a22134a );
 a22139a <=( a22138a  and  a22131a );
 a22143a <=( A167  and  (not A169) );
 a22144a <=( A170  and  a22143a );
 a22148a <=( A200  and  A199 );
 a22149a <=( (not A166)  and  a22148a );
 a22150a <=( a22149a  and  a22144a );
 a22154a <=( (not A269)  and  (not A268) );
 a22155a <=( (not A266)  and  a22154a );
 a22158a <=( (not A299)  and  A298 );
 a22161a <=( A301  and  A300 );
 a22162a <=( a22161a  and  a22158a );
 a22163a <=( a22162a  and  a22155a );
 a22167a <=( A167  and  (not A169) );
 a22168a <=( A170  and  a22167a );
 a22172a <=( A200  and  A199 );
 a22173a <=( (not A166)  and  a22172a );
 a22174a <=( a22173a  and  a22168a );
 a22178a <=( (not A269)  and  (not A268) );
 a22179a <=( (not A266)  and  a22178a );
 a22182a <=( (not A299)  and  A298 );
 a22185a <=( A302  and  A300 );
 a22186a <=( a22185a  and  a22182a );
 a22187a <=( a22186a  and  a22179a );
 a22191a <=( A167  and  (not A169) );
 a22192a <=( A170  and  a22191a );
 a22196a <=( A200  and  (not A199) );
 a22197a <=( (not A166)  and  a22196a );
 a22198a <=( a22197a  and  a22192a );
 a22202a <=( A267  and  (not A266) );
 a22203a <=( A265  and  a22202a );
 a22206a <=( A298  and  A268 );
 a22209a <=( (not A302)  and  (not A301) );
 a22210a <=( a22209a  and  a22206a );
 a22211a <=( a22210a  and  a22203a );
 a22215a <=( A167  and  (not A169) );
 a22216a <=( A170  and  a22215a );
 a22220a <=( A200  and  (not A199) );
 a22221a <=( (not A166)  and  a22220a );
 a22222a <=( a22221a  and  a22216a );
 a22226a <=( A267  and  (not A266) );
 a22227a <=( A265  and  a22226a );
 a22230a <=( A298  and  A269 );
 a22233a <=( (not A302)  and  (not A301) );
 a22234a <=( a22233a  and  a22230a );
 a22235a <=( a22234a  and  a22227a );
 a22239a <=( A167  and  (not A169) );
 a22240a <=( A170  and  a22239a );
 a22244a <=( (not A202)  and  (not A200) );
 a22245a <=( (not A166)  and  a22244a );
 a22246a <=( a22245a  and  a22240a );
 a22250a <=( A266  and  A265 );
 a22251a <=( (not A203)  and  a22250a );
 a22254a <=( (not A299)  and  A298 );
 a22257a <=( A301  and  A300 );
 a22258a <=( a22257a  and  a22254a );
 a22259a <=( a22258a  and  a22251a );
 a22263a <=( A167  and  (not A169) );
 a22264a <=( A170  and  a22263a );
 a22268a <=( (not A202)  and  (not A200) );
 a22269a <=( (not A166)  and  a22268a );
 a22270a <=( a22269a  and  a22264a );
 a22274a <=( A266  and  A265 );
 a22275a <=( (not A203)  and  a22274a );
 a22278a <=( (not A299)  and  A298 );
 a22281a <=( A302  and  A300 );
 a22282a <=( a22281a  and  a22278a );
 a22283a <=( a22282a  and  a22275a );
 a22287a <=( A167  and  (not A169) );
 a22288a <=( A170  and  a22287a );
 a22292a <=( (not A202)  and  (not A200) );
 a22293a <=( (not A166)  and  a22292a );
 a22294a <=( a22293a  and  a22288a );
 a22298a <=( (not A267)  and  (not A266) );
 a22299a <=( (not A203)  and  a22298a );
 a22302a <=( (not A299)  and  A298 );
 a22305a <=( A301  and  A300 );
 a22306a <=( a22305a  and  a22302a );
 a22307a <=( a22306a  and  a22299a );
 a22311a <=( A167  and  (not A169) );
 a22312a <=( A170  and  a22311a );
 a22316a <=( (not A202)  and  (not A200) );
 a22317a <=( (not A166)  and  a22316a );
 a22318a <=( a22317a  and  a22312a );
 a22322a <=( (not A267)  and  (not A266) );
 a22323a <=( (not A203)  and  a22322a );
 a22326a <=( (not A299)  and  A298 );
 a22329a <=( A302  and  A300 );
 a22330a <=( a22329a  and  a22326a );
 a22331a <=( a22330a  and  a22323a );
 a22335a <=( A167  and  (not A169) );
 a22336a <=( A170  and  a22335a );
 a22340a <=( (not A202)  and  (not A200) );
 a22341a <=( (not A166)  and  a22340a );
 a22342a <=( a22341a  and  a22336a );
 a22346a <=( (not A266)  and  (not A265) );
 a22347a <=( (not A203)  and  a22346a );
 a22350a <=( (not A299)  and  A298 );
 a22353a <=( A301  and  A300 );
 a22354a <=( a22353a  and  a22350a );
 a22355a <=( a22354a  and  a22347a );
 a22359a <=( A167  and  (not A169) );
 a22360a <=( A170  and  a22359a );
 a22364a <=( (not A202)  and  (not A200) );
 a22365a <=( (not A166)  and  a22364a );
 a22366a <=( a22365a  and  a22360a );
 a22370a <=( (not A266)  and  (not A265) );
 a22371a <=( (not A203)  and  a22370a );
 a22374a <=( (not A299)  and  A298 );
 a22377a <=( A302  and  A300 );
 a22378a <=( a22377a  and  a22374a );
 a22379a <=( a22378a  and  a22371a );
 a22383a <=( A167  and  (not A169) );
 a22384a <=( A170  and  a22383a );
 a22388a <=( (not A201)  and  (not A200) );
 a22389a <=( (not A166)  and  a22388a );
 a22390a <=( a22389a  and  a22384a );
 a22394a <=( (not A269)  and  (not A268) );
 a22395a <=( (not A266)  and  a22394a );
 a22398a <=( (not A299)  and  A298 );
 a22401a <=( A301  and  A300 );
 a22402a <=( a22401a  and  a22398a );
 a22403a <=( a22402a  and  a22395a );
 a22407a <=( A167  and  (not A169) );
 a22408a <=( A170  and  a22407a );
 a22412a <=( (not A201)  and  (not A200) );
 a22413a <=( (not A166)  and  a22412a );
 a22414a <=( a22413a  and  a22408a );
 a22418a <=( (not A269)  and  (not A268) );
 a22419a <=( (not A266)  and  a22418a );
 a22422a <=( (not A299)  and  A298 );
 a22425a <=( A302  and  A300 );
 a22426a <=( a22425a  and  a22422a );
 a22427a <=( a22426a  and  a22419a );
 a22431a <=( A167  and  (not A169) );
 a22432a <=( A170  and  a22431a );
 a22436a <=( (not A200)  and  A199 );
 a22437a <=( (not A166)  and  a22436a );
 a22438a <=( a22437a  and  a22432a );
 a22442a <=( (not A265)  and  A202 );
 a22443a <=( A201  and  a22442a );
 a22446a <=( A298  and  A266 );
 a22449a <=( (not A302)  and  (not A301) );
 a22450a <=( a22449a  and  a22446a );
 a22451a <=( a22450a  and  a22443a );
 a22455a <=( A167  and  (not A169) );
 a22456a <=( A170  and  a22455a );
 a22460a <=( (not A200)  and  A199 );
 a22461a <=( (not A166)  and  a22460a );
 a22462a <=( a22461a  and  a22456a );
 a22466a <=( (not A265)  and  A203 );
 a22467a <=( A201  and  a22466a );
 a22470a <=( A298  and  A266 );
 a22473a <=( (not A302)  and  (not A301) );
 a22474a <=( a22473a  and  a22470a );
 a22475a <=( a22474a  and  a22467a );
 a22479a <=( A167  and  (not A169) );
 a22480a <=( A170  and  a22479a );
 a22484a <=( (not A200)  and  (not A199) );
 a22485a <=( (not A166)  and  a22484a );
 a22486a <=( a22485a  and  a22480a );
 a22490a <=( (not A269)  and  (not A268) );
 a22491a <=( (not A266)  and  a22490a );
 a22494a <=( (not A299)  and  A298 );
 a22497a <=( A301  and  A300 );
 a22498a <=( a22497a  and  a22494a );
 a22499a <=( a22498a  and  a22491a );
 a22503a <=( A167  and  (not A169) );
 a22504a <=( A170  and  a22503a );
 a22508a <=( (not A200)  and  (not A199) );
 a22509a <=( (not A166)  and  a22508a );
 a22510a <=( a22509a  and  a22504a );
 a22514a <=( (not A269)  and  (not A268) );
 a22515a <=( (not A266)  and  a22514a );
 a22518a <=( (not A299)  and  A298 );
 a22521a <=( A302  and  A300 );
 a22522a <=( a22521a  and  a22518a );
 a22523a <=( a22522a  and  a22515a );
 a22527a <=( (not A167)  and  (not A169) );
 a22528a <=( A170  and  a22527a );
 a22532a <=( A200  and  A199 );
 a22533a <=( A166  and  a22532a );
 a22534a <=( a22533a  and  a22528a );
 a22538a <=( (not A269)  and  (not A268) );
 a22539a <=( (not A266)  and  a22538a );
 a22542a <=( (not A299)  and  A298 );
 a22545a <=( A301  and  A300 );
 a22546a <=( a22545a  and  a22542a );
 a22547a <=( a22546a  and  a22539a );
 a22551a <=( (not A167)  and  (not A169) );
 a22552a <=( A170  and  a22551a );
 a22556a <=( A200  and  A199 );
 a22557a <=( A166  and  a22556a );
 a22558a <=( a22557a  and  a22552a );
 a22562a <=( (not A269)  and  (not A268) );
 a22563a <=( (not A266)  and  a22562a );
 a22566a <=( (not A299)  and  A298 );
 a22569a <=( A302  and  A300 );
 a22570a <=( a22569a  and  a22566a );
 a22571a <=( a22570a  and  a22563a );
 a22575a <=( (not A167)  and  (not A169) );
 a22576a <=( A170  and  a22575a );
 a22580a <=( A200  and  (not A199) );
 a22581a <=( A166  and  a22580a );
 a22582a <=( a22581a  and  a22576a );
 a22586a <=( A267  and  (not A266) );
 a22587a <=( A265  and  a22586a );
 a22590a <=( A298  and  A268 );
 a22593a <=( (not A302)  and  (not A301) );
 a22594a <=( a22593a  and  a22590a );
 a22595a <=( a22594a  and  a22587a );
 a22599a <=( (not A167)  and  (not A169) );
 a22600a <=( A170  and  a22599a );
 a22604a <=( A200  and  (not A199) );
 a22605a <=( A166  and  a22604a );
 a22606a <=( a22605a  and  a22600a );
 a22610a <=( A267  and  (not A266) );
 a22611a <=( A265  and  a22610a );
 a22614a <=( A298  and  A269 );
 a22617a <=( (not A302)  and  (not A301) );
 a22618a <=( a22617a  and  a22614a );
 a22619a <=( a22618a  and  a22611a );
 a22623a <=( (not A167)  and  (not A169) );
 a22624a <=( A170  and  a22623a );
 a22628a <=( (not A202)  and  (not A200) );
 a22629a <=( A166  and  a22628a );
 a22630a <=( a22629a  and  a22624a );
 a22634a <=( A266  and  A265 );
 a22635a <=( (not A203)  and  a22634a );
 a22638a <=( (not A299)  and  A298 );
 a22641a <=( A301  and  A300 );
 a22642a <=( a22641a  and  a22638a );
 a22643a <=( a22642a  and  a22635a );
 a22647a <=( (not A167)  and  (not A169) );
 a22648a <=( A170  and  a22647a );
 a22652a <=( (not A202)  and  (not A200) );
 a22653a <=( A166  and  a22652a );
 a22654a <=( a22653a  and  a22648a );
 a22658a <=( A266  and  A265 );
 a22659a <=( (not A203)  and  a22658a );
 a22662a <=( (not A299)  and  A298 );
 a22665a <=( A302  and  A300 );
 a22666a <=( a22665a  and  a22662a );
 a22667a <=( a22666a  and  a22659a );
 a22671a <=( (not A167)  and  (not A169) );
 a22672a <=( A170  and  a22671a );
 a22676a <=( (not A202)  and  (not A200) );
 a22677a <=( A166  and  a22676a );
 a22678a <=( a22677a  and  a22672a );
 a22682a <=( (not A267)  and  (not A266) );
 a22683a <=( (not A203)  and  a22682a );
 a22686a <=( (not A299)  and  A298 );
 a22689a <=( A301  and  A300 );
 a22690a <=( a22689a  and  a22686a );
 a22691a <=( a22690a  and  a22683a );
 a22695a <=( (not A167)  and  (not A169) );
 a22696a <=( A170  and  a22695a );
 a22700a <=( (not A202)  and  (not A200) );
 a22701a <=( A166  and  a22700a );
 a22702a <=( a22701a  and  a22696a );
 a22706a <=( (not A267)  and  (not A266) );
 a22707a <=( (not A203)  and  a22706a );
 a22710a <=( (not A299)  and  A298 );
 a22713a <=( A302  and  A300 );
 a22714a <=( a22713a  and  a22710a );
 a22715a <=( a22714a  and  a22707a );
 a22719a <=( (not A167)  and  (not A169) );
 a22720a <=( A170  and  a22719a );
 a22724a <=( (not A202)  and  (not A200) );
 a22725a <=( A166  and  a22724a );
 a22726a <=( a22725a  and  a22720a );
 a22730a <=( (not A266)  and  (not A265) );
 a22731a <=( (not A203)  and  a22730a );
 a22734a <=( (not A299)  and  A298 );
 a22737a <=( A301  and  A300 );
 a22738a <=( a22737a  and  a22734a );
 a22739a <=( a22738a  and  a22731a );
 a22743a <=( (not A167)  and  (not A169) );
 a22744a <=( A170  and  a22743a );
 a22748a <=( (not A202)  and  (not A200) );
 a22749a <=( A166  and  a22748a );
 a22750a <=( a22749a  and  a22744a );
 a22754a <=( (not A266)  and  (not A265) );
 a22755a <=( (not A203)  and  a22754a );
 a22758a <=( (not A299)  and  A298 );
 a22761a <=( A302  and  A300 );
 a22762a <=( a22761a  and  a22758a );
 a22763a <=( a22762a  and  a22755a );
 a22767a <=( (not A167)  and  (not A169) );
 a22768a <=( A170  and  a22767a );
 a22772a <=( (not A201)  and  (not A200) );
 a22773a <=( A166  and  a22772a );
 a22774a <=( a22773a  and  a22768a );
 a22778a <=( (not A269)  and  (not A268) );
 a22779a <=( (not A266)  and  a22778a );
 a22782a <=( (not A299)  and  A298 );
 a22785a <=( A301  and  A300 );
 a22786a <=( a22785a  and  a22782a );
 a22787a <=( a22786a  and  a22779a );
 a22791a <=( (not A167)  and  (not A169) );
 a22792a <=( A170  and  a22791a );
 a22796a <=( (not A201)  and  (not A200) );
 a22797a <=( A166  and  a22796a );
 a22798a <=( a22797a  and  a22792a );
 a22802a <=( (not A269)  and  (not A268) );
 a22803a <=( (not A266)  and  a22802a );
 a22806a <=( (not A299)  and  A298 );
 a22809a <=( A302  and  A300 );
 a22810a <=( a22809a  and  a22806a );
 a22811a <=( a22810a  and  a22803a );
 a22815a <=( (not A167)  and  (not A169) );
 a22816a <=( A170  and  a22815a );
 a22820a <=( (not A200)  and  A199 );
 a22821a <=( A166  and  a22820a );
 a22822a <=( a22821a  and  a22816a );
 a22826a <=( (not A265)  and  A202 );
 a22827a <=( A201  and  a22826a );
 a22830a <=( A298  and  A266 );
 a22833a <=( (not A302)  and  (not A301) );
 a22834a <=( a22833a  and  a22830a );
 a22835a <=( a22834a  and  a22827a );
 a22839a <=( (not A167)  and  (not A169) );
 a22840a <=( A170  and  a22839a );
 a22844a <=( (not A200)  and  A199 );
 a22845a <=( A166  and  a22844a );
 a22846a <=( a22845a  and  a22840a );
 a22850a <=( (not A265)  and  A203 );
 a22851a <=( A201  and  a22850a );
 a22854a <=( A298  and  A266 );
 a22857a <=( (not A302)  and  (not A301) );
 a22858a <=( a22857a  and  a22854a );
 a22859a <=( a22858a  and  a22851a );
 a22863a <=( (not A167)  and  (not A169) );
 a22864a <=( A170  and  a22863a );
 a22868a <=( (not A200)  and  (not A199) );
 a22869a <=( A166  and  a22868a );
 a22870a <=( a22869a  and  a22864a );
 a22874a <=( (not A269)  and  (not A268) );
 a22875a <=( (not A266)  and  a22874a );
 a22878a <=( (not A299)  and  A298 );
 a22881a <=( A301  and  A300 );
 a22882a <=( a22881a  and  a22878a );
 a22883a <=( a22882a  and  a22875a );
 a22887a <=( (not A167)  and  (not A169) );
 a22888a <=( A170  and  a22887a );
 a22892a <=( (not A200)  and  (not A199) );
 a22893a <=( A166  and  a22892a );
 a22894a <=( a22893a  and  a22888a );
 a22898a <=( (not A269)  and  (not A268) );
 a22899a <=( (not A266)  and  a22898a );
 a22902a <=( (not A299)  and  A298 );
 a22905a <=( A302  and  A300 );
 a22906a <=( a22905a  and  a22902a );
 a22907a <=( a22906a  and  a22899a );
 a22911a <=( (not A168)  and  (not A169) );
 a22912a <=( (not A170)  and  a22911a );
 a22916a <=( (not A203)  and  (not A202) );
 a22917a <=( (not A200)  and  a22916a );
 a22918a <=( a22917a  and  a22912a );
 a22922a <=( A267  and  (not A266) );
 a22923a <=( A265  and  a22922a );
 a22926a <=( A298  and  A268 );
 a22929a <=( (not A302)  and  (not A301) );
 a22930a <=( a22929a  and  a22926a );
 a22931a <=( a22930a  and  a22923a );
 a22935a <=( (not A168)  and  (not A169) );
 a22936a <=( (not A170)  and  a22935a );
 a22940a <=( (not A203)  and  (not A202) );
 a22941a <=( (not A200)  and  a22940a );
 a22942a <=( a22941a  and  a22936a );
 a22946a <=( A267  and  (not A266) );
 a22947a <=( A265  and  a22946a );
 a22950a <=( A298  and  A269 );
 a22953a <=( (not A302)  and  (not A301) );
 a22954a <=( a22953a  and  a22950a );
 a22955a <=( a22954a  and  a22947a );
 a22959a <=( (not A168)  and  (not A169) );
 a22960a <=( (not A170)  and  a22959a );
 a22964a <=( A201  and  (not A200) );
 a22965a <=( A199  and  a22964a );
 a22966a <=( a22965a  and  a22960a );
 a22970a <=( A266  and  A265 );
 a22971a <=( A202  and  a22970a );
 a22974a <=( (not A299)  and  A298 );
 a22977a <=( A301  and  A300 );
 a22978a <=( a22977a  and  a22974a );
 a22979a <=( a22978a  and  a22971a );
 a22983a <=( (not A168)  and  (not A169) );
 a22984a <=( (not A170)  and  a22983a );
 a22988a <=( A201  and  (not A200) );
 a22989a <=( A199  and  a22988a );
 a22990a <=( a22989a  and  a22984a );
 a22994a <=( A266  and  A265 );
 a22995a <=( A202  and  a22994a );
 a22998a <=( (not A299)  and  A298 );
 a23001a <=( A302  and  A300 );
 a23002a <=( a23001a  and  a22998a );
 a23003a <=( a23002a  and  a22995a );
 a23007a <=( (not A168)  and  (not A169) );
 a23008a <=( (not A170)  and  a23007a );
 a23012a <=( A201  and  (not A200) );
 a23013a <=( A199  and  a23012a );
 a23014a <=( a23013a  and  a23008a );
 a23018a <=( (not A267)  and  (not A266) );
 a23019a <=( A202  and  a23018a );
 a23022a <=( (not A299)  and  A298 );
 a23025a <=( A301  and  A300 );
 a23026a <=( a23025a  and  a23022a );
 a23027a <=( a23026a  and  a23019a );
 a23031a <=( (not A168)  and  (not A169) );
 a23032a <=( (not A170)  and  a23031a );
 a23036a <=( A201  and  (not A200) );
 a23037a <=( A199  and  a23036a );
 a23038a <=( a23037a  and  a23032a );
 a23042a <=( (not A267)  and  (not A266) );
 a23043a <=( A202  and  a23042a );
 a23046a <=( (not A299)  and  A298 );
 a23049a <=( A302  and  A300 );
 a23050a <=( a23049a  and  a23046a );
 a23051a <=( a23050a  and  a23043a );
 a23055a <=( (not A168)  and  (not A169) );
 a23056a <=( (not A170)  and  a23055a );
 a23060a <=( A201  and  (not A200) );
 a23061a <=( A199  and  a23060a );
 a23062a <=( a23061a  and  a23056a );
 a23066a <=( (not A266)  and  (not A265) );
 a23067a <=( A202  and  a23066a );
 a23070a <=( (not A299)  and  A298 );
 a23073a <=( A301  and  A300 );
 a23074a <=( a23073a  and  a23070a );
 a23075a <=( a23074a  and  a23067a );
 a23079a <=( (not A168)  and  (not A169) );
 a23080a <=( (not A170)  and  a23079a );
 a23084a <=( A201  and  (not A200) );
 a23085a <=( A199  and  a23084a );
 a23086a <=( a23085a  and  a23080a );
 a23090a <=( (not A266)  and  (not A265) );
 a23091a <=( A202  and  a23090a );
 a23094a <=( (not A299)  and  A298 );
 a23097a <=( A302  and  A300 );
 a23098a <=( a23097a  and  a23094a );
 a23099a <=( a23098a  and  a23091a );
 a23103a <=( (not A168)  and  (not A169) );
 a23104a <=( (not A170)  and  a23103a );
 a23108a <=( A201  and  (not A200) );
 a23109a <=( A199  and  a23108a );
 a23110a <=( a23109a  and  a23104a );
 a23114a <=( A266  and  A265 );
 a23115a <=( A203  and  a23114a );
 a23118a <=( (not A299)  and  A298 );
 a23121a <=( A301  and  A300 );
 a23122a <=( a23121a  and  a23118a );
 a23123a <=( a23122a  and  a23115a );
 a23127a <=( (not A168)  and  (not A169) );
 a23128a <=( (not A170)  and  a23127a );
 a23132a <=( A201  and  (not A200) );
 a23133a <=( A199  and  a23132a );
 a23134a <=( a23133a  and  a23128a );
 a23138a <=( A266  and  A265 );
 a23139a <=( A203  and  a23138a );
 a23142a <=( (not A299)  and  A298 );
 a23145a <=( A302  and  A300 );
 a23146a <=( a23145a  and  a23142a );
 a23147a <=( a23146a  and  a23139a );
 a23151a <=( (not A168)  and  (not A169) );
 a23152a <=( (not A170)  and  a23151a );
 a23156a <=( A201  and  (not A200) );
 a23157a <=( A199  and  a23156a );
 a23158a <=( a23157a  and  a23152a );
 a23162a <=( (not A267)  and  (not A266) );
 a23163a <=( A203  and  a23162a );
 a23166a <=( (not A299)  and  A298 );
 a23169a <=( A301  and  A300 );
 a23170a <=( a23169a  and  a23166a );
 a23171a <=( a23170a  and  a23163a );
 a23175a <=( (not A168)  and  (not A169) );
 a23176a <=( (not A170)  and  a23175a );
 a23180a <=( A201  and  (not A200) );
 a23181a <=( A199  and  a23180a );
 a23182a <=( a23181a  and  a23176a );
 a23186a <=( (not A267)  and  (not A266) );
 a23187a <=( A203  and  a23186a );
 a23190a <=( (not A299)  and  A298 );
 a23193a <=( A302  and  A300 );
 a23194a <=( a23193a  and  a23190a );
 a23195a <=( a23194a  and  a23187a );
 a23199a <=( (not A168)  and  (not A169) );
 a23200a <=( (not A170)  and  a23199a );
 a23204a <=( A201  and  (not A200) );
 a23205a <=( A199  and  a23204a );
 a23206a <=( a23205a  and  a23200a );
 a23210a <=( (not A266)  and  (not A265) );
 a23211a <=( A203  and  a23210a );
 a23214a <=( (not A299)  and  A298 );
 a23217a <=( A301  and  A300 );
 a23218a <=( a23217a  and  a23214a );
 a23219a <=( a23218a  and  a23211a );
 a23223a <=( (not A168)  and  (not A169) );
 a23224a <=( (not A170)  and  a23223a );
 a23228a <=( A201  and  (not A200) );
 a23229a <=( A199  and  a23228a );
 a23230a <=( a23229a  and  a23224a );
 a23234a <=( (not A266)  and  (not A265) );
 a23235a <=( A203  and  a23234a );
 a23238a <=( (not A299)  and  A298 );
 a23241a <=( A302  and  A300 );
 a23242a <=( a23241a  and  a23238a );
 a23243a <=( a23242a  and  a23235a );
 a23247a <=( (not A166)  and  (not A167) );
 a23248a <=( A170  and  a23247a );
 a23251a <=( (not A200)  and  A199 );
 a23254a <=( A202  and  A201 );
 a23255a <=( a23254a  and  a23251a );
 a23256a <=( a23255a  and  a23248a );
 a23260a <=( (not A269)  and  (not A268) );
 a23261a <=( (not A266)  and  a23260a );
 a23264a <=( (not A299)  and  A298 );
 a23267a <=( A301  and  A300 );
 a23268a <=( a23267a  and  a23264a );
 a23269a <=( a23268a  and  a23261a );
 a23273a <=( (not A166)  and  (not A167) );
 a23274a <=( A170  and  a23273a );
 a23277a <=( (not A200)  and  A199 );
 a23280a <=( A202  and  A201 );
 a23281a <=( a23280a  and  a23277a );
 a23282a <=( a23281a  and  a23274a );
 a23286a <=( (not A269)  and  (not A268) );
 a23287a <=( (not A266)  and  a23286a );
 a23290a <=( (not A299)  and  A298 );
 a23293a <=( A302  and  A300 );
 a23294a <=( a23293a  and  a23290a );
 a23295a <=( a23294a  and  a23287a );
 a23299a <=( (not A166)  and  (not A167) );
 a23300a <=( A170  and  a23299a );
 a23303a <=( (not A200)  and  A199 );
 a23306a <=( A203  and  A201 );
 a23307a <=( a23306a  and  a23303a );
 a23308a <=( a23307a  and  a23300a );
 a23312a <=( (not A269)  and  (not A268) );
 a23313a <=( (not A266)  and  a23312a );
 a23316a <=( (not A299)  and  A298 );
 a23319a <=( A301  and  A300 );
 a23320a <=( a23319a  and  a23316a );
 a23321a <=( a23320a  and  a23313a );
 a23325a <=( (not A166)  and  (not A167) );
 a23326a <=( A170  and  a23325a );
 a23329a <=( (not A200)  and  A199 );
 a23332a <=( A203  and  A201 );
 a23333a <=( a23332a  and  a23329a );
 a23334a <=( a23333a  and  a23326a );
 a23338a <=( (not A269)  and  (not A268) );
 a23339a <=( (not A266)  and  a23338a );
 a23342a <=( (not A299)  and  A298 );
 a23345a <=( A302  and  A300 );
 a23346a <=( a23345a  and  a23342a );
 a23347a <=( a23346a  and  a23339a );
 a23351a <=( A167  and  (not A168) );
 a23352a <=( A169  and  a23351a );
 a23355a <=( (not A200)  and  (not A166) );
 a23358a <=( (not A203)  and  (not A202) );
 a23359a <=( a23358a  and  a23355a );
 a23360a <=( a23359a  and  a23352a );
 a23364a <=( A267  and  (not A266) );
 a23365a <=( A265  and  a23364a );
 a23368a <=( A298  and  A268 );
 a23371a <=( (not A302)  and  (not A301) );
 a23372a <=( a23371a  and  a23368a );
 a23373a <=( a23372a  and  a23365a );
 a23377a <=( A167  and  (not A168) );
 a23378a <=( A169  and  a23377a );
 a23381a <=( (not A200)  and  (not A166) );
 a23384a <=( (not A203)  and  (not A202) );
 a23385a <=( a23384a  and  a23381a );
 a23386a <=( a23385a  and  a23378a );
 a23390a <=( A267  and  (not A266) );
 a23391a <=( A265  and  a23390a );
 a23394a <=( A298  and  A269 );
 a23397a <=( (not A302)  and  (not A301) );
 a23398a <=( a23397a  and  a23394a );
 a23399a <=( a23398a  and  a23391a );
 a23403a <=( A167  and  (not A168) );
 a23404a <=( A169  and  a23403a );
 a23407a <=( A199  and  (not A166) );
 a23410a <=( A201  and  (not A200) );
 a23411a <=( a23410a  and  a23407a );
 a23412a <=( a23411a  and  a23404a );
 a23416a <=( A266  and  A265 );
 a23417a <=( A202  and  a23416a );
 a23420a <=( (not A299)  and  A298 );
 a23423a <=( A301  and  A300 );
 a23424a <=( a23423a  and  a23420a );
 a23425a <=( a23424a  and  a23417a );
 a23429a <=( A167  and  (not A168) );
 a23430a <=( A169  and  a23429a );
 a23433a <=( A199  and  (not A166) );
 a23436a <=( A201  and  (not A200) );
 a23437a <=( a23436a  and  a23433a );
 a23438a <=( a23437a  and  a23430a );
 a23442a <=( A266  and  A265 );
 a23443a <=( A202  and  a23442a );
 a23446a <=( (not A299)  and  A298 );
 a23449a <=( A302  and  A300 );
 a23450a <=( a23449a  and  a23446a );
 a23451a <=( a23450a  and  a23443a );
 a23455a <=( A167  and  (not A168) );
 a23456a <=( A169  and  a23455a );
 a23459a <=( A199  and  (not A166) );
 a23462a <=( A201  and  (not A200) );
 a23463a <=( a23462a  and  a23459a );
 a23464a <=( a23463a  and  a23456a );
 a23468a <=( (not A267)  and  (not A266) );
 a23469a <=( A202  and  a23468a );
 a23472a <=( (not A299)  and  A298 );
 a23475a <=( A301  and  A300 );
 a23476a <=( a23475a  and  a23472a );
 a23477a <=( a23476a  and  a23469a );
 a23481a <=( A167  and  (not A168) );
 a23482a <=( A169  and  a23481a );
 a23485a <=( A199  and  (not A166) );
 a23488a <=( A201  and  (not A200) );
 a23489a <=( a23488a  and  a23485a );
 a23490a <=( a23489a  and  a23482a );
 a23494a <=( (not A267)  and  (not A266) );
 a23495a <=( A202  and  a23494a );
 a23498a <=( (not A299)  and  A298 );
 a23501a <=( A302  and  A300 );
 a23502a <=( a23501a  and  a23498a );
 a23503a <=( a23502a  and  a23495a );
 a23507a <=( A167  and  (not A168) );
 a23508a <=( A169  and  a23507a );
 a23511a <=( A199  and  (not A166) );
 a23514a <=( A201  and  (not A200) );
 a23515a <=( a23514a  and  a23511a );
 a23516a <=( a23515a  and  a23508a );
 a23520a <=( (not A266)  and  (not A265) );
 a23521a <=( A202  and  a23520a );
 a23524a <=( (not A299)  and  A298 );
 a23527a <=( A301  and  A300 );
 a23528a <=( a23527a  and  a23524a );
 a23529a <=( a23528a  and  a23521a );
 a23533a <=( A167  and  (not A168) );
 a23534a <=( A169  and  a23533a );
 a23537a <=( A199  and  (not A166) );
 a23540a <=( A201  and  (not A200) );
 a23541a <=( a23540a  and  a23537a );
 a23542a <=( a23541a  and  a23534a );
 a23546a <=( (not A266)  and  (not A265) );
 a23547a <=( A202  and  a23546a );
 a23550a <=( (not A299)  and  A298 );
 a23553a <=( A302  and  A300 );
 a23554a <=( a23553a  and  a23550a );
 a23555a <=( a23554a  and  a23547a );
 a23559a <=( A167  and  (not A168) );
 a23560a <=( A169  and  a23559a );
 a23563a <=( A199  and  (not A166) );
 a23566a <=( A201  and  (not A200) );
 a23567a <=( a23566a  and  a23563a );
 a23568a <=( a23567a  and  a23560a );
 a23572a <=( A266  and  A265 );
 a23573a <=( A203  and  a23572a );
 a23576a <=( (not A299)  and  A298 );
 a23579a <=( A301  and  A300 );
 a23580a <=( a23579a  and  a23576a );
 a23581a <=( a23580a  and  a23573a );
 a23585a <=( A167  and  (not A168) );
 a23586a <=( A169  and  a23585a );
 a23589a <=( A199  and  (not A166) );
 a23592a <=( A201  and  (not A200) );
 a23593a <=( a23592a  and  a23589a );
 a23594a <=( a23593a  and  a23586a );
 a23598a <=( A266  and  A265 );
 a23599a <=( A203  and  a23598a );
 a23602a <=( (not A299)  and  A298 );
 a23605a <=( A302  and  A300 );
 a23606a <=( a23605a  and  a23602a );
 a23607a <=( a23606a  and  a23599a );
 a23611a <=( A167  and  (not A168) );
 a23612a <=( A169  and  a23611a );
 a23615a <=( A199  and  (not A166) );
 a23618a <=( A201  and  (not A200) );
 a23619a <=( a23618a  and  a23615a );
 a23620a <=( a23619a  and  a23612a );
 a23624a <=( (not A267)  and  (not A266) );
 a23625a <=( A203  and  a23624a );
 a23628a <=( (not A299)  and  A298 );
 a23631a <=( A301  and  A300 );
 a23632a <=( a23631a  and  a23628a );
 a23633a <=( a23632a  and  a23625a );
 a23637a <=( A167  and  (not A168) );
 a23638a <=( A169  and  a23637a );
 a23641a <=( A199  and  (not A166) );
 a23644a <=( A201  and  (not A200) );
 a23645a <=( a23644a  and  a23641a );
 a23646a <=( a23645a  and  a23638a );
 a23650a <=( (not A267)  and  (not A266) );
 a23651a <=( A203  and  a23650a );
 a23654a <=( (not A299)  and  A298 );
 a23657a <=( A302  and  A300 );
 a23658a <=( a23657a  and  a23654a );
 a23659a <=( a23658a  and  a23651a );
 a23663a <=( A167  and  (not A168) );
 a23664a <=( A169  and  a23663a );
 a23667a <=( A199  and  (not A166) );
 a23670a <=( A201  and  (not A200) );
 a23671a <=( a23670a  and  a23667a );
 a23672a <=( a23671a  and  a23664a );
 a23676a <=( (not A266)  and  (not A265) );
 a23677a <=( A203  and  a23676a );
 a23680a <=( (not A299)  and  A298 );
 a23683a <=( A301  and  A300 );
 a23684a <=( a23683a  and  a23680a );
 a23685a <=( a23684a  and  a23677a );
 a23689a <=( A167  and  (not A168) );
 a23690a <=( A169  and  a23689a );
 a23693a <=( A199  and  (not A166) );
 a23696a <=( A201  and  (not A200) );
 a23697a <=( a23696a  and  a23693a );
 a23698a <=( a23697a  and  a23690a );
 a23702a <=( (not A266)  and  (not A265) );
 a23703a <=( A203  and  a23702a );
 a23706a <=( (not A299)  and  A298 );
 a23709a <=( A302  and  A300 );
 a23710a <=( a23709a  and  a23706a );
 a23711a <=( a23710a  and  a23703a );
 a23715a <=( (not A167)  and  (not A168) );
 a23716a <=( A169  and  a23715a );
 a23719a <=( (not A200)  and  A166 );
 a23722a <=( (not A203)  and  (not A202) );
 a23723a <=( a23722a  and  a23719a );
 a23724a <=( a23723a  and  a23716a );
 a23728a <=( A267  and  (not A266) );
 a23729a <=( A265  and  a23728a );
 a23732a <=( A298  and  A268 );
 a23735a <=( (not A302)  and  (not A301) );
 a23736a <=( a23735a  and  a23732a );
 a23737a <=( a23736a  and  a23729a );
 a23741a <=( (not A167)  and  (not A168) );
 a23742a <=( A169  and  a23741a );
 a23745a <=( (not A200)  and  A166 );
 a23748a <=( (not A203)  and  (not A202) );
 a23749a <=( a23748a  and  a23745a );
 a23750a <=( a23749a  and  a23742a );
 a23754a <=( A267  and  (not A266) );
 a23755a <=( A265  and  a23754a );
 a23758a <=( A298  and  A269 );
 a23761a <=( (not A302)  and  (not A301) );
 a23762a <=( a23761a  and  a23758a );
 a23763a <=( a23762a  and  a23755a );
 a23767a <=( (not A167)  and  (not A168) );
 a23768a <=( A169  and  a23767a );
 a23771a <=( A199  and  A166 );
 a23774a <=( A201  and  (not A200) );
 a23775a <=( a23774a  and  a23771a );
 a23776a <=( a23775a  and  a23768a );
 a23780a <=( A266  and  A265 );
 a23781a <=( A202  and  a23780a );
 a23784a <=( (not A299)  and  A298 );
 a23787a <=( A301  and  A300 );
 a23788a <=( a23787a  and  a23784a );
 a23789a <=( a23788a  and  a23781a );
 a23793a <=( (not A167)  and  (not A168) );
 a23794a <=( A169  and  a23793a );
 a23797a <=( A199  and  A166 );
 a23800a <=( A201  and  (not A200) );
 a23801a <=( a23800a  and  a23797a );
 a23802a <=( a23801a  and  a23794a );
 a23806a <=( A266  and  A265 );
 a23807a <=( A202  and  a23806a );
 a23810a <=( (not A299)  and  A298 );
 a23813a <=( A302  and  A300 );
 a23814a <=( a23813a  and  a23810a );
 a23815a <=( a23814a  and  a23807a );
 a23819a <=( (not A167)  and  (not A168) );
 a23820a <=( A169  and  a23819a );
 a23823a <=( A199  and  A166 );
 a23826a <=( A201  and  (not A200) );
 a23827a <=( a23826a  and  a23823a );
 a23828a <=( a23827a  and  a23820a );
 a23832a <=( (not A267)  and  (not A266) );
 a23833a <=( A202  and  a23832a );
 a23836a <=( (not A299)  and  A298 );
 a23839a <=( A301  and  A300 );
 a23840a <=( a23839a  and  a23836a );
 a23841a <=( a23840a  and  a23833a );
 a23845a <=( (not A167)  and  (not A168) );
 a23846a <=( A169  and  a23845a );
 a23849a <=( A199  and  A166 );
 a23852a <=( A201  and  (not A200) );
 a23853a <=( a23852a  and  a23849a );
 a23854a <=( a23853a  and  a23846a );
 a23858a <=( (not A267)  and  (not A266) );
 a23859a <=( A202  and  a23858a );
 a23862a <=( (not A299)  and  A298 );
 a23865a <=( A302  and  A300 );
 a23866a <=( a23865a  and  a23862a );
 a23867a <=( a23866a  and  a23859a );
 a23871a <=( (not A167)  and  (not A168) );
 a23872a <=( A169  and  a23871a );
 a23875a <=( A199  and  A166 );
 a23878a <=( A201  and  (not A200) );
 a23879a <=( a23878a  and  a23875a );
 a23880a <=( a23879a  and  a23872a );
 a23884a <=( (not A266)  and  (not A265) );
 a23885a <=( A202  and  a23884a );
 a23888a <=( (not A299)  and  A298 );
 a23891a <=( A301  and  A300 );
 a23892a <=( a23891a  and  a23888a );
 a23893a <=( a23892a  and  a23885a );
 a23897a <=( (not A167)  and  (not A168) );
 a23898a <=( A169  and  a23897a );
 a23901a <=( A199  and  A166 );
 a23904a <=( A201  and  (not A200) );
 a23905a <=( a23904a  and  a23901a );
 a23906a <=( a23905a  and  a23898a );
 a23910a <=( (not A266)  and  (not A265) );
 a23911a <=( A202  and  a23910a );
 a23914a <=( (not A299)  and  A298 );
 a23917a <=( A302  and  A300 );
 a23918a <=( a23917a  and  a23914a );
 a23919a <=( a23918a  and  a23911a );
 a23923a <=( (not A167)  and  (not A168) );
 a23924a <=( A169  and  a23923a );
 a23927a <=( A199  and  A166 );
 a23930a <=( A201  and  (not A200) );
 a23931a <=( a23930a  and  a23927a );
 a23932a <=( a23931a  and  a23924a );
 a23936a <=( A266  and  A265 );
 a23937a <=( A203  and  a23936a );
 a23940a <=( (not A299)  and  A298 );
 a23943a <=( A301  and  A300 );
 a23944a <=( a23943a  and  a23940a );
 a23945a <=( a23944a  and  a23937a );
 a23949a <=( (not A167)  and  (not A168) );
 a23950a <=( A169  and  a23949a );
 a23953a <=( A199  and  A166 );
 a23956a <=( A201  and  (not A200) );
 a23957a <=( a23956a  and  a23953a );
 a23958a <=( a23957a  and  a23950a );
 a23962a <=( A266  and  A265 );
 a23963a <=( A203  and  a23962a );
 a23966a <=( (not A299)  and  A298 );
 a23969a <=( A302  and  A300 );
 a23970a <=( a23969a  and  a23966a );
 a23971a <=( a23970a  and  a23963a );
 a23975a <=( (not A167)  and  (not A168) );
 a23976a <=( A169  and  a23975a );
 a23979a <=( A199  and  A166 );
 a23982a <=( A201  and  (not A200) );
 a23983a <=( a23982a  and  a23979a );
 a23984a <=( a23983a  and  a23976a );
 a23988a <=( (not A267)  and  (not A266) );
 a23989a <=( A203  and  a23988a );
 a23992a <=( (not A299)  and  A298 );
 a23995a <=( A301  and  A300 );
 a23996a <=( a23995a  and  a23992a );
 a23997a <=( a23996a  and  a23989a );
 a24001a <=( (not A167)  and  (not A168) );
 a24002a <=( A169  and  a24001a );
 a24005a <=( A199  and  A166 );
 a24008a <=( A201  and  (not A200) );
 a24009a <=( a24008a  and  a24005a );
 a24010a <=( a24009a  and  a24002a );
 a24014a <=( (not A267)  and  (not A266) );
 a24015a <=( A203  and  a24014a );
 a24018a <=( (not A299)  and  A298 );
 a24021a <=( A302  and  A300 );
 a24022a <=( a24021a  and  a24018a );
 a24023a <=( a24022a  and  a24015a );
 a24027a <=( (not A167)  and  (not A168) );
 a24028a <=( A169  and  a24027a );
 a24031a <=( A199  and  A166 );
 a24034a <=( A201  and  (not A200) );
 a24035a <=( a24034a  and  a24031a );
 a24036a <=( a24035a  and  a24028a );
 a24040a <=( (not A266)  and  (not A265) );
 a24041a <=( A203  and  a24040a );
 a24044a <=( (not A299)  and  A298 );
 a24047a <=( A301  and  A300 );
 a24048a <=( a24047a  and  a24044a );
 a24049a <=( a24048a  and  a24041a );
 a24053a <=( (not A167)  and  (not A168) );
 a24054a <=( A169  and  a24053a );
 a24057a <=( A199  and  A166 );
 a24060a <=( A201  and  (not A200) );
 a24061a <=( a24060a  and  a24057a );
 a24062a <=( a24061a  and  a24054a );
 a24066a <=( (not A266)  and  (not A265) );
 a24067a <=( A203  and  a24066a );
 a24070a <=( (not A299)  and  A298 );
 a24073a <=( A302  and  A300 );
 a24074a <=( a24073a  and  a24070a );
 a24075a <=( a24074a  and  a24067a );
 a24079a <=( (not A168)  and  A169 );
 a24080a <=( A170  and  a24079a );
 a24083a <=( (not A200)  and  A199 );
 a24086a <=( A202  and  A201 );
 a24087a <=( a24086a  and  a24083a );
 a24088a <=( a24087a  and  a24080a );
 a24092a <=( (not A269)  and  (not A268) );
 a24093a <=( (not A266)  and  a24092a );
 a24096a <=( (not A299)  and  A298 );
 a24099a <=( A301  and  A300 );
 a24100a <=( a24099a  and  a24096a );
 a24101a <=( a24100a  and  a24093a );
 a24105a <=( (not A168)  and  A169 );
 a24106a <=( A170  and  a24105a );
 a24109a <=( (not A200)  and  A199 );
 a24112a <=( A202  and  A201 );
 a24113a <=( a24112a  and  a24109a );
 a24114a <=( a24113a  and  a24106a );
 a24118a <=( (not A269)  and  (not A268) );
 a24119a <=( (not A266)  and  a24118a );
 a24122a <=( (not A299)  and  A298 );
 a24125a <=( A302  and  A300 );
 a24126a <=( a24125a  and  a24122a );
 a24127a <=( a24126a  and  a24119a );
 a24131a <=( (not A168)  and  A169 );
 a24132a <=( A170  and  a24131a );
 a24135a <=( (not A200)  and  A199 );
 a24138a <=( A203  and  A201 );
 a24139a <=( a24138a  and  a24135a );
 a24140a <=( a24139a  and  a24132a );
 a24144a <=( (not A269)  and  (not A268) );
 a24145a <=( (not A266)  and  a24144a );
 a24148a <=( (not A299)  and  A298 );
 a24151a <=( A301  and  A300 );
 a24152a <=( a24151a  and  a24148a );
 a24153a <=( a24152a  and  a24145a );
 a24157a <=( (not A168)  and  A169 );
 a24158a <=( A170  and  a24157a );
 a24161a <=( (not A200)  and  A199 );
 a24164a <=( A203  and  A201 );
 a24165a <=( a24164a  and  a24161a );
 a24166a <=( a24165a  and  a24158a );
 a24170a <=( (not A269)  and  (not A268) );
 a24171a <=( (not A266)  and  a24170a );
 a24174a <=( (not A299)  and  A298 );
 a24177a <=( A302  and  A300 );
 a24178a <=( a24177a  and  a24174a );
 a24179a <=( a24178a  and  a24171a );
 a24183a <=( A167  and  A169 );
 a24184a <=( (not A170)  and  a24183a );
 a24187a <=( (not A200)  and  A166 );
 a24190a <=( (not A203)  and  (not A202) );
 a24191a <=( a24190a  and  a24187a );
 a24192a <=( a24191a  and  a24184a );
 a24196a <=( (not A269)  and  (not A268) );
 a24197a <=( (not A266)  and  a24196a );
 a24200a <=( (not A299)  and  A298 );
 a24203a <=( A301  and  A300 );
 a24204a <=( a24203a  and  a24200a );
 a24205a <=( a24204a  and  a24197a );
 a24209a <=( A167  and  A169 );
 a24210a <=( (not A170)  and  a24209a );
 a24213a <=( (not A200)  and  A166 );
 a24216a <=( (not A203)  and  (not A202) );
 a24217a <=( a24216a  and  a24213a );
 a24218a <=( a24217a  and  a24210a );
 a24222a <=( (not A269)  and  (not A268) );
 a24223a <=( (not A266)  and  a24222a );
 a24226a <=( (not A299)  and  A298 );
 a24229a <=( A302  and  A300 );
 a24230a <=( a24229a  and  a24226a );
 a24231a <=( a24230a  and  a24223a );
 a24235a <=( A167  and  A169 );
 a24236a <=( (not A170)  and  a24235a );
 a24239a <=( A199  and  A166 );
 a24242a <=( A201  and  (not A200) );
 a24243a <=( a24242a  and  a24239a );
 a24244a <=( a24243a  and  a24236a );
 a24248a <=( (not A266)  and  A265 );
 a24249a <=( A202  and  a24248a );
 a24252a <=( A268  and  A267 );
 a24255a <=( (not A300)  and  A298 );
 a24256a <=( a24255a  and  a24252a );
 a24257a <=( a24256a  and  a24249a );
 a24261a <=( A167  and  A169 );
 a24262a <=( (not A170)  and  a24261a );
 a24265a <=( A199  and  A166 );
 a24268a <=( A201  and  (not A200) );
 a24269a <=( a24268a  and  a24265a );
 a24270a <=( a24269a  and  a24262a );
 a24274a <=( (not A266)  and  A265 );
 a24275a <=( A202  and  a24274a );
 a24278a <=( A268  and  A267 );
 a24281a <=( A299  and  A298 );
 a24282a <=( a24281a  and  a24278a );
 a24283a <=( a24282a  and  a24275a );
 a24287a <=( A167  and  A169 );
 a24288a <=( (not A170)  and  a24287a );
 a24291a <=( A199  and  A166 );
 a24294a <=( A201  and  (not A200) );
 a24295a <=( a24294a  and  a24291a );
 a24296a <=( a24295a  and  a24288a );
 a24300a <=( (not A266)  and  A265 );
 a24301a <=( A202  and  a24300a );
 a24304a <=( A268  and  A267 );
 a24307a <=( (not A299)  and  (not A298) );
 a24308a <=( a24307a  and  a24304a );
 a24309a <=( a24308a  and  a24301a );
 a24313a <=( A167  and  A169 );
 a24314a <=( (not A170)  and  a24313a );
 a24317a <=( A199  and  A166 );
 a24320a <=( A201  and  (not A200) );
 a24321a <=( a24320a  and  a24317a );
 a24322a <=( a24321a  and  a24314a );
 a24326a <=( (not A266)  and  A265 );
 a24327a <=( A202  and  a24326a );
 a24330a <=( A269  and  A267 );
 a24333a <=( (not A300)  and  A298 );
 a24334a <=( a24333a  and  a24330a );
 a24335a <=( a24334a  and  a24327a );
 a24339a <=( A167  and  A169 );
 a24340a <=( (not A170)  and  a24339a );
 a24343a <=( A199  and  A166 );
 a24346a <=( A201  and  (not A200) );
 a24347a <=( a24346a  and  a24343a );
 a24348a <=( a24347a  and  a24340a );
 a24352a <=( (not A266)  and  A265 );
 a24353a <=( A202  and  a24352a );
 a24356a <=( A269  and  A267 );
 a24359a <=( A299  and  A298 );
 a24360a <=( a24359a  and  a24356a );
 a24361a <=( a24360a  and  a24353a );
 a24365a <=( A167  and  A169 );
 a24366a <=( (not A170)  and  a24365a );
 a24369a <=( A199  and  A166 );
 a24372a <=( A201  and  (not A200) );
 a24373a <=( a24372a  and  a24369a );
 a24374a <=( a24373a  and  a24366a );
 a24378a <=( (not A266)  and  A265 );
 a24379a <=( A202  and  a24378a );
 a24382a <=( A269  and  A267 );
 a24385a <=( (not A299)  and  (not A298) );
 a24386a <=( a24385a  and  a24382a );
 a24387a <=( a24386a  and  a24379a );
 a24391a <=( A167  and  A169 );
 a24392a <=( (not A170)  and  a24391a );
 a24395a <=( A199  and  A166 );
 a24398a <=( A201  and  (not A200) );
 a24399a <=( a24398a  and  a24395a );
 a24400a <=( a24399a  and  a24392a );
 a24404a <=( (not A266)  and  A265 );
 a24405a <=( A203  and  a24404a );
 a24408a <=( A268  and  A267 );
 a24411a <=( (not A300)  and  A298 );
 a24412a <=( a24411a  and  a24408a );
 a24413a <=( a24412a  and  a24405a );
 a24417a <=( A167  and  A169 );
 a24418a <=( (not A170)  and  a24417a );
 a24421a <=( A199  and  A166 );
 a24424a <=( A201  and  (not A200) );
 a24425a <=( a24424a  and  a24421a );
 a24426a <=( a24425a  and  a24418a );
 a24430a <=( (not A266)  and  A265 );
 a24431a <=( A203  and  a24430a );
 a24434a <=( A268  and  A267 );
 a24437a <=( A299  and  A298 );
 a24438a <=( a24437a  and  a24434a );
 a24439a <=( a24438a  and  a24431a );
 a24443a <=( A167  and  A169 );
 a24444a <=( (not A170)  and  a24443a );
 a24447a <=( A199  and  A166 );
 a24450a <=( A201  and  (not A200) );
 a24451a <=( a24450a  and  a24447a );
 a24452a <=( a24451a  and  a24444a );
 a24456a <=( (not A266)  and  A265 );
 a24457a <=( A203  and  a24456a );
 a24460a <=( A268  and  A267 );
 a24463a <=( (not A299)  and  (not A298) );
 a24464a <=( a24463a  and  a24460a );
 a24465a <=( a24464a  and  a24457a );
 a24469a <=( A167  and  A169 );
 a24470a <=( (not A170)  and  a24469a );
 a24473a <=( A199  and  A166 );
 a24476a <=( A201  and  (not A200) );
 a24477a <=( a24476a  and  a24473a );
 a24478a <=( a24477a  and  a24470a );
 a24482a <=( (not A266)  and  A265 );
 a24483a <=( A203  and  a24482a );
 a24486a <=( A269  and  A267 );
 a24489a <=( (not A300)  and  A298 );
 a24490a <=( a24489a  and  a24486a );
 a24491a <=( a24490a  and  a24483a );
 a24495a <=( A167  and  A169 );
 a24496a <=( (not A170)  and  a24495a );
 a24499a <=( A199  and  A166 );
 a24502a <=( A201  and  (not A200) );
 a24503a <=( a24502a  and  a24499a );
 a24504a <=( a24503a  and  a24496a );
 a24508a <=( (not A266)  and  A265 );
 a24509a <=( A203  and  a24508a );
 a24512a <=( A269  and  A267 );
 a24515a <=( A299  and  A298 );
 a24516a <=( a24515a  and  a24512a );
 a24517a <=( a24516a  and  a24509a );
 a24521a <=( A167  and  A169 );
 a24522a <=( (not A170)  and  a24521a );
 a24525a <=( A199  and  A166 );
 a24528a <=( A201  and  (not A200) );
 a24529a <=( a24528a  and  a24525a );
 a24530a <=( a24529a  and  a24522a );
 a24534a <=( (not A266)  and  A265 );
 a24535a <=( A203  and  a24534a );
 a24538a <=( A269  and  A267 );
 a24541a <=( (not A299)  and  (not A298) );
 a24542a <=( a24541a  and  a24538a );
 a24543a <=( a24542a  and  a24535a );
 a24547a <=( (not A167)  and  A169 );
 a24548a <=( (not A170)  and  a24547a );
 a24551a <=( (not A200)  and  (not A166) );
 a24554a <=( (not A203)  and  (not A202) );
 a24555a <=( a24554a  and  a24551a );
 a24556a <=( a24555a  and  a24548a );
 a24560a <=( (not A269)  and  (not A268) );
 a24561a <=( (not A266)  and  a24560a );
 a24564a <=( (not A299)  and  A298 );
 a24567a <=( A301  and  A300 );
 a24568a <=( a24567a  and  a24564a );
 a24569a <=( a24568a  and  a24561a );
 a24573a <=( (not A167)  and  A169 );
 a24574a <=( (not A170)  and  a24573a );
 a24577a <=( (not A200)  and  (not A166) );
 a24580a <=( (not A203)  and  (not A202) );
 a24581a <=( a24580a  and  a24577a );
 a24582a <=( a24581a  and  a24574a );
 a24586a <=( (not A269)  and  (not A268) );
 a24587a <=( (not A266)  and  a24586a );
 a24590a <=( (not A299)  and  A298 );
 a24593a <=( A302  and  A300 );
 a24594a <=( a24593a  and  a24590a );
 a24595a <=( a24594a  and  a24587a );
 a24599a <=( (not A167)  and  A169 );
 a24600a <=( (not A170)  and  a24599a );
 a24603a <=( A199  and  (not A166) );
 a24606a <=( A201  and  (not A200) );
 a24607a <=( a24606a  and  a24603a );
 a24608a <=( a24607a  and  a24600a );
 a24612a <=( (not A266)  and  A265 );
 a24613a <=( A202  and  a24612a );
 a24616a <=( A268  and  A267 );
 a24619a <=( (not A300)  and  A298 );
 a24620a <=( a24619a  and  a24616a );
 a24621a <=( a24620a  and  a24613a );
 a24625a <=( (not A167)  and  A169 );
 a24626a <=( (not A170)  and  a24625a );
 a24629a <=( A199  and  (not A166) );
 a24632a <=( A201  and  (not A200) );
 a24633a <=( a24632a  and  a24629a );
 a24634a <=( a24633a  and  a24626a );
 a24638a <=( (not A266)  and  A265 );
 a24639a <=( A202  and  a24638a );
 a24642a <=( A268  and  A267 );
 a24645a <=( A299  and  A298 );
 a24646a <=( a24645a  and  a24642a );
 a24647a <=( a24646a  and  a24639a );
 a24651a <=( (not A167)  and  A169 );
 a24652a <=( (not A170)  and  a24651a );
 a24655a <=( A199  and  (not A166) );
 a24658a <=( A201  and  (not A200) );
 a24659a <=( a24658a  and  a24655a );
 a24660a <=( a24659a  and  a24652a );
 a24664a <=( (not A266)  and  A265 );
 a24665a <=( A202  and  a24664a );
 a24668a <=( A268  and  A267 );
 a24671a <=( (not A299)  and  (not A298) );
 a24672a <=( a24671a  and  a24668a );
 a24673a <=( a24672a  and  a24665a );
 a24677a <=( (not A167)  and  A169 );
 a24678a <=( (not A170)  and  a24677a );
 a24681a <=( A199  and  (not A166) );
 a24684a <=( A201  and  (not A200) );
 a24685a <=( a24684a  and  a24681a );
 a24686a <=( a24685a  and  a24678a );
 a24690a <=( (not A266)  and  A265 );
 a24691a <=( A202  and  a24690a );
 a24694a <=( A269  and  A267 );
 a24697a <=( (not A300)  and  A298 );
 a24698a <=( a24697a  and  a24694a );
 a24699a <=( a24698a  and  a24691a );
 a24703a <=( (not A167)  and  A169 );
 a24704a <=( (not A170)  and  a24703a );
 a24707a <=( A199  and  (not A166) );
 a24710a <=( A201  and  (not A200) );
 a24711a <=( a24710a  and  a24707a );
 a24712a <=( a24711a  and  a24704a );
 a24716a <=( (not A266)  and  A265 );
 a24717a <=( A202  and  a24716a );
 a24720a <=( A269  and  A267 );
 a24723a <=( A299  and  A298 );
 a24724a <=( a24723a  and  a24720a );
 a24725a <=( a24724a  and  a24717a );
 a24729a <=( (not A167)  and  A169 );
 a24730a <=( (not A170)  and  a24729a );
 a24733a <=( A199  and  (not A166) );
 a24736a <=( A201  and  (not A200) );
 a24737a <=( a24736a  and  a24733a );
 a24738a <=( a24737a  and  a24730a );
 a24742a <=( (not A266)  and  A265 );
 a24743a <=( A202  and  a24742a );
 a24746a <=( A269  and  A267 );
 a24749a <=( (not A299)  and  (not A298) );
 a24750a <=( a24749a  and  a24746a );
 a24751a <=( a24750a  and  a24743a );
 a24755a <=( (not A167)  and  A169 );
 a24756a <=( (not A170)  and  a24755a );
 a24759a <=( A199  and  (not A166) );
 a24762a <=( A201  and  (not A200) );
 a24763a <=( a24762a  and  a24759a );
 a24764a <=( a24763a  and  a24756a );
 a24768a <=( (not A266)  and  A265 );
 a24769a <=( A203  and  a24768a );
 a24772a <=( A268  and  A267 );
 a24775a <=( (not A300)  and  A298 );
 a24776a <=( a24775a  and  a24772a );
 a24777a <=( a24776a  and  a24769a );
 a24781a <=( (not A167)  and  A169 );
 a24782a <=( (not A170)  and  a24781a );
 a24785a <=( A199  and  (not A166) );
 a24788a <=( A201  and  (not A200) );
 a24789a <=( a24788a  and  a24785a );
 a24790a <=( a24789a  and  a24782a );
 a24794a <=( (not A266)  and  A265 );
 a24795a <=( A203  and  a24794a );
 a24798a <=( A268  and  A267 );
 a24801a <=( A299  and  A298 );
 a24802a <=( a24801a  and  a24798a );
 a24803a <=( a24802a  and  a24795a );
 a24807a <=( (not A167)  and  A169 );
 a24808a <=( (not A170)  and  a24807a );
 a24811a <=( A199  and  (not A166) );
 a24814a <=( A201  and  (not A200) );
 a24815a <=( a24814a  and  a24811a );
 a24816a <=( a24815a  and  a24808a );
 a24820a <=( (not A266)  and  A265 );
 a24821a <=( A203  and  a24820a );
 a24824a <=( A268  and  A267 );
 a24827a <=( (not A299)  and  (not A298) );
 a24828a <=( a24827a  and  a24824a );
 a24829a <=( a24828a  and  a24821a );
 a24833a <=( (not A167)  and  A169 );
 a24834a <=( (not A170)  and  a24833a );
 a24837a <=( A199  and  (not A166) );
 a24840a <=( A201  and  (not A200) );
 a24841a <=( a24840a  and  a24837a );
 a24842a <=( a24841a  and  a24834a );
 a24846a <=( (not A266)  and  A265 );
 a24847a <=( A203  and  a24846a );
 a24850a <=( A269  and  A267 );
 a24853a <=( (not A300)  and  A298 );
 a24854a <=( a24853a  and  a24850a );
 a24855a <=( a24854a  and  a24847a );
 a24859a <=( (not A167)  and  A169 );
 a24860a <=( (not A170)  and  a24859a );
 a24863a <=( A199  and  (not A166) );
 a24866a <=( A201  and  (not A200) );
 a24867a <=( a24866a  and  a24863a );
 a24868a <=( a24867a  and  a24860a );
 a24872a <=( (not A266)  and  A265 );
 a24873a <=( A203  and  a24872a );
 a24876a <=( A269  and  A267 );
 a24879a <=( A299  and  A298 );
 a24880a <=( a24879a  and  a24876a );
 a24881a <=( a24880a  and  a24873a );
 a24885a <=( (not A167)  and  A169 );
 a24886a <=( (not A170)  and  a24885a );
 a24889a <=( A199  and  (not A166) );
 a24892a <=( A201  and  (not A200) );
 a24893a <=( a24892a  and  a24889a );
 a24894a <=( a24893a  and  a24886a );
 a24898a <=( (not A266)  and  A265 );
 a24899a <=( A203  and  a24898a );
 a24902a <=( A269  and  A267 );
 a24905a <=( (not A299)  and  (not A298) );
 a24906a <=( a24905a  and  a24902a );
 a24907a <=( a24906a  and  a24899a );
 a24911a <=( (not A166)  and  (not A167) );
 a24912a <=( (not A169)  and  a24911a );
 a24915a <=( (not A200)  and  A199 );
 a24918a <=( A202  and  A201 );
 a24919a <=( a24918a  and  a24915a );
 a24920a <=( a24919a  and  a24912a );
 a24924a <=( (not A269)  and  (not A268) );
 a24925a <=( (not A266)  and  a24924a );
 a24928a <=( (not A299)  and  A298 );
 a24931a <=( A301  and  A300 );
 a24932a <=( a24931a  and  a24928a );
 a24933a <=( a24932a  and  a24925a );
 a24937a <=( (not A166)  and  (not A167) );
 a24938a <=( (not A169)  and  a24937a );
 a24941a <=( (not A200)  and  A199 );
 a24944a <=( A202  and  A201 );
 a24945a <=( a24944a  and  a24941a );
 a24946a <=( a24945a  and  a24938a );
 a24950a <=( (not A269)  and  (not A268) );
 a24951a <=( (not A266)  and  a24950a );
 a24954a <=( (not A299)  and  A298 );
 a24957a <=( A302  and  A300 );
 a24958a <=( a24957a  and  a24954a );
 a24959a <=( a24958a  and  a24951a );
 a24963a <=( (not A166)  and  (not A167) );
 a24964a <=( (not A169)  and  a24963a );
 a24967a <=( (not A200)  and  A199 );
 a24970a <=( A203  and  A201 );
 a24971a <=( a24970a  and  a24967a );
 a24972a <=( a24971a  and  a24964a );
 a24976a <=( (not A269)  and  (not A268) );
 a24977a <=( (not A266)  and  a24976a );
 a24980a <=( (not A299)  and  A298 );
 a24983a <=( A301  and  A300 );
 a24984a <=( a24983a  and  a24980a );
 a24985a <=( a24984a  and  a24977a );
 a24989a <=( (not A166)  and  (not A167) );
 a24990a <=( (not A169)  and  a24989a );
 a24993a <=( (not A200)  and  A199 );
 a24996a <=( A203  and  A201 );
 a24997a <=( a24996a  and  a24993a );
 a24998a <=( a24997a  and  a24990a );
 a25002a <=( (not A269)  and  (not A268) );
 a25003a <=( (not A266)  and  a25002a );
 a25006a <=( (not A299)  and  A298 );
 a25009a <=( A302  and  A300 );
 a25010a <=( a25009a  and  a25006a );
 a25011a <=( a25010a  and  a25003a );
 a25015a <=( A167  and  (not A168) );
 a25016a <=( (not A169)  and  a25015a );
 a25019a <=( (not A200)  and  A166 );
 a25022a <=( (not A203)  and  (not A202) );
 a25023a <=( a25022a  and  a25019a );
 a25024a <=( a25023a  and  a25016a );
 a25028a <=( A267  and  (not A266) );
 a25029a <=( A265  and  a25028a );
 a25032a <=( A298  and  A268 );
 a25035a <=( (not A302)  and  (not A301) );
 a25036a <=( a25035a  and  a25032a );
 a25037a <=( a25036a  and  a25029a );
 a25041a <=( A167  and  (not A168) );
 a25042a <=( (not A169)  and  a25041a );
 a25045a <=( (not A200)  and  A166 );
 a25048a <=( (not A203)  and  (not A202) );
 a25049a <=( a25048a  and  a25045a );
 a25050a <=( a25049a  and  a25042a );
 a25054a <=( A267  and  (not A266) );
 a25055a <=( A265  and  a25054a );
 a25058a <=( A298  and  A269 );
 a25061a <=( (not A302)  and  (not A301) );
 a25062a <=( a25061a  and  a25058a );
 a25063a <=( a25062a  and  a25055a );
 a25067a <=( A167  and  (not A168) );
 a25068a <=( (not A169)  and  a25067a );
 a25071a <=( A199  and  A166 );
 a25074a <=( A201  and  (not A200) );
 a25075a <=( a25074a  and  a25071a );
 a25076a <=( a25075a  and  a25068a );
 a25080a <=( A266  and  A265 );
 a25081a <=( A202  and  a25080a );
 a25084a <=( (not A299)  and  A298 );
 a25087a <=( A301  and  A300 );
 a25088a <=( a25087a  and  a25084a );
 a25089a <=( a25088a  and  a25081a );
 a25093a <=( A167  and  (not A168) );
 a25094a <=( (not A169)  and  a25093a );
 a25097a <=( A199  and  A166 );
 a25100a <=( A201  and  (not A200) );
 a25101a <=( a25100a  and  a25097a );
 a25102a <=( a25101a  and  a25094a );
 a25106a <=( A266  and  A265 );
 a25107a <=( A202  and  a25106a );
 a25110a <=( (not A299)  and  A298 );
 a25113a <=( A302  and  A300 );
 a25114a <=( a25113a  and  a25110a );
 a25115a <=( a25114a  and  a25107a );
 a25119a <=( A167  and  (not A168) );
 a25120a <=( (not A169)  and  a25119a );
 a25123a <=( A199  and  A166 );
 a25126a <=( A201  and  (not A200) );
 a25127a <=( a25126a  and  a25123a );
 a25128a <=( a25127a  and  a25120a );
 a25132a <=( (not A267)  and  (not A266) );
 a25133a <=( A202  and  a25132a );
 a25136a <=( (not A299)  and  A298 );
 a25139a <=( A301  and  A300 );
 a25140a <=( a25139a  and  a25136a );
 a25141a <=( a25140a  and  a25133a );
 a25145a <=( A167  and  (not A168) );
 a25146a <=( (not A169)  and  a25145a );
 a25149a <=( A199  and  A166 );
 a25152a <=( A201  and  (not A200) );
 a25153a <=( a25152a  and  a25149a );
 a25154a <=( a25153a  and  a25146a );
 a25158a <=( (not A267)  and  (not A266) );
 a25159a <=( A202  and  a25158a );
 a25162a <=( (not A299)  and  A298 );
 a25165a <=( A302  and  A300 );
 a25166a <=( a25165a  and  a25162a );
 a25167a <=( a25166a  and  a25159a );
 a25171a <=( A167  and  (not A168) );
 a25172a <=( (not A169)  and  a25171a );
 a25175a <=( A199  and  A166 );
 a25178a <=( A201  and  (not A200) );
 a25179a <=( a25178a  and  a25175a );
 a25180a <=( a25179a  and  a25172a );
 a25184a <=( (not A266)  and  (not A265) );
 a25185a <=( A202  and  a25184a );
 a25188a <=( (not A299)  and  A298 );
 a25191a <=( A301  and  A300 );
 a25192a <=( a25191a  and  a25188a );
 a25193a <=( a25192a  and  a25185a );
 a25197a <=( A167  and  (not A168) );
 a25198a <=( (not A169)  and  a25197a );
 a25201a <=( A199  and  A166 );
 a25204a <=( A201  and  (not A200) );
 a25205a <=( a25204a  and  a25201a );
 a25206a <=( a25205a  and  a25198a );
 a25210a <=( (not A266)  and  (not A265) );
 a25211a <=( A202  and  a25210a );
 a25214a <=( (not A299)  and  A298 );
 a25217a <=( A302  and  A300 );
 a25218a <=( a25217a  and  a25214a );
 a25219a <=( a25218a  and  a25211a );
 a25223a <=( A167  and  (not A168) );
 a25224a <=( (not A169)  and  a25223a );
 a25227a <=( A199  and  A166 );
 a25230a <=( A201  and  (not A200) );
 a25231a <=( a25230a  and  a25227a );
 a25232a <=( a25231a  and  a25224a );
 a25236a <=( A266  and  A265 );
 a25237a <=( A203  and  a25236a );
 a25240a <=( (not A299)  and  A298 );
 a25243a <=( A301  and  A300 );
 a25244a <=( a25243a  and  a25240a );
 a25245a <=( a25244a  and  a25237a );
 a25249a <=( A167  and  (not A168) );
 a25250a <=( (not A169)  and  a25249a );
 a25253a <=( A199  and  A166 );
 a25256a <=( A201  and  (not A200) );
 a25257a <=( a25256a  and  a25253a );
 a25258a <=( a25257a  and  a25250a );
 a25262a <=( A266  and  A265 );
 a25263a <=( A203  and  a25262a );
 a25266a <=( (not A299)  and  A298 );
 a25269a <=( A302  and  A300 );
 a25270a <=( a25269a  and  a25266a );
 a25271a <=( a25270a  and  a25263a );
 a25275a <=( A167  and  (not A168) );
 a25276a <=( (not A169)  and  a25275a );
 a25279a <=( A199  and  A166 );
 a25282a <=( A201  and  (not A200) );
 a25283a <=( a25282a  and  a25279a );
 a25284a <=( a25283a  and  a25276a );
 a25288a <=( (not A267)  and  (not A266) );
 a25289a <=( A203  and  a25288a );
 a25292a <=( (not A299)  and  A298 );
 a25295a <=( A301  and  A300 );
 a25296a <=( a25295a  and  a25292a );
 a25297a <=( a25296a  and  a25289a );
 a25301a <=( A167  and  (not A168) );
 a25302a <=( (not A169)  and  a25301a );
 a25305a <=( A199  and  A166 );
 a25308a <=( A201  and  (not A200) );
 a25309a <=( a25308a  and  a25305a );
 a25310a <=( a25309a  and  a25302a );
 a25314a <=( (not A267)  and  (not A266) );
 a25315a <=( A203  and  a25314a );
 a25318a <=( (not A299)  and  A298 );
 a25321a <=( A302  and  A300 );
 a25322a <=( a25321a  and  a25318a );
 a25323a <=( a25322a  and  a25315a );
 a25327a <=( A167  and  (not A168) );
 a25328a <=( (not A169)  and  a25327a );
 a25331a <=( A199  and  A166 );
 a25334a <=( A201  and  (not A200) );
 a25335a <=( a25334a  and  a25331a );
 a25336a <=( a25335a  and  a25328a );
 a25340a <=( (not A266)  and  (not A265) );
 a25341a <=( A203  and  a25340a );
 a25344a <=( (not A299)  and  A298 );
 a25347a <=( A301  and  A300 );
 a25348a <=( a25347a  and  a25344a );
 a25349a <=( a25348a  and  a25341a );
 a25353a <=( A167  and  (not A168) );
 a25354a <=( (not A169)  and  a25353a );
 a25357a <=( A199  and  A166 );
 a25360a <=( A201  and  (not A200) );
 a25361a <=( a25360a  and  a25357a );
 a25362a <=( a25361a  and  a25354a );
 a25366a <=( (not A266)  and  (not A265) );
 a25367a <=( A203  and  a25366a );
 a25370a <=( (not A299)  and  A298 );
 a25373a <=( A302  and  A300 );
 a25374a <=( a25373a  and  a25370a );
 a25375a <=( a25374a  and  a25367a );
 a25379a <=( A167  and  (not A169) );
 a25380a <=( A170  and  a25379a );
 a25383a <=( (not A200)  and  (not A166) );
 a25386a <=( (not A203)  and  (not A202) );
 a25387a <=( a25386a  and  a25383a );
 a25388a <=( a25387a  and  a25380a );
 a25392a <=( (not A269)  and  (not A268) );
 a25393a <=( (not A266)  and  a25392a );
 a25396a <=( (not A299)  and  A298 );
 a25399a <=( A301  and  A300 );
 a25400a <=( a25399a  and  a25396a );
 a25401a <=( a25400a  and  a25393a );
 a25405a <=( A167  and  (not A169) );
 a25406a <=( A170  and  a25405a );
 a25409a <=( (not A200)  and  (not A166) );
 a25412a <=( (not A203)  and  (not A202) );
 a25413a <=( a25412a  and  a25409a );
 a25414a <=( a25413a  and  a25406a );
 a25418a <=( (not A269)  and  (not A268) );
 a25419a <=( (not A266)  and  a25418a );
 a25422a <=( (not A299)  and  A298 );
 a25425a <=( A302  and  A300 );
 a25426a <=( a25425a  and  a25422a );
 a25427a <=( a25426a  and  a25419a );
 a25431a <=( A167  and  (not A169) );
 a25432a <=( A170  and  a25431a );
 a25435a <=( A199  and  (not A166) );
 a25438a <=( A201  and  (not A200) );
 a25439a <=( a25438a  and  a25435a );
 a25440a <=( a25439a  and  a25432a );
 a25444a <=( (not A266)  and  A265 );
 a25445a <=( A202  and  a25444a );
 a25448a <=( A268  and  A267 );
 a25451a <=( (not A300)  and  A298 );
 a25452a <=( a25451a  and  a25448a );
 a25453a <=( a25452a  and  a25445a );
 a25457a <=( A167  and  (not A169) );
 a25458a <=( A170  and  a25457a );
 a25461a <=( A199  and  (not A166) );
 a25464a <=( A201  and  (not A200) );
 a25465a <=( a25464a  and  a25461a );
 a25466a <=( a25465a  and  a25458a );
 a25470a <=( (not A266)  and  A265 );
 a25471a <=( A202  and  a25470a );
 a25474a <=( A268  and  A267 );
 a25477a <=( A299  and  A298 );
 a25478a <=( a25477a  and  a25474a );
 a25479a <=( a25478a  and  a25471a );
 a25483a <=( A167  and  (not A169) );
 a25484a <=( A170  and  a25483a );
 a25487a <=( A199  and  (not A166) );
 a25490a <=( A201  and  (not A200) );
 a25491a <=( a25490a  and  a25487a );
 a25492a <=( a25491a  and  a25484a );
 a25496a <=( (not A266)  and  A265 );
 a25497a <=( A202  and  a25496a );
 a25500a <=( A268  and  A267 );
 a25503a <=( (not A299)  and  (not A298) );
 a25504a <=( a25503a  and  a25500a );
 a25505a <=( a25504a  and  a25497a );
 a25509a <=( A167  and  (not A169) );
 a25510a <=( A170  and  a25509a );
 a25513a <=( A199  and  (not A166) );
 a25516a <=( A201  and  (not A200) );
 a25517a <=( a25516a  and  a25513a );
 a25518a <=( a25517a  and  a25510a );
 a25522a <=( (not A266)  and  A265 );
 a25523a <=( A202  and  a25522a );
 a25526a <=( A269  and  A267 );
 a25529a <=( (not A300)  and  A298 );
 a25530a <=( a25529a  and  a25526a );
 a25531a <=( a25530a  and  a25523a );
 a25535a <=( A167  and  (not A169) );
 a25536a <=( A170  and  a25535a );
 a25539a <=( A199  and  (not A166) );
 a25542a <=( A201  and  (not A200) );
 a25543a <=( a25542a  and  a25539a );
 a25544a <=( a25543a  and  a25536a );
 a25548a <=( (not A266)  and  A265 );
 a25549a <=( A202  and  a25548a );
 a25552a <=( A269  and  A267 );
 a25555a <=( A299  and  A298 );
 a25556a <=( a25555a  and  a25552a );
 a25557a <=( a25556a  and  a25549a );
 a25561a <=( A167  and  (not A169) );
 a25562a <=( A170  and  a25561a );
 a25565a <=( A199  and  (not A166) );
 a25568a <=( A201  and  (not A200) );
 a25569a <=( a25568a  and  a25565a );
 a25570a <=( a25569a  and  a25562a );
 a25574a <=( (not A266)  and  A265 );
 a25575a <=( A202  and  a25574a );
 a25578a <=( A269  and  A267 );
 a25581a <=( (not A299)  and  (not A298) );
 a25582a <=( a25581a  and  a25578a );
 a25583a <=( a25582a  and  a25575a );
 a25587a <=( A167  and  (not A169) );
 a25588a <=( A170  and  a25587a );
 a25591a <=( A199  and  (not A166) );
 a25594a <=( A201  and  (not A200) );
 a25595a <=( a25594a  and  a25591a );
 a25596a <=( a25595a  and  a25588a );
 a25600a <=( (not A266)  and  A265 );
 a25601a <=( A203  and  a25600a );
 a25604a <=( A268  and  A267 );
 a25607a <=( (not A300)  and  A298 );
 a25608a <=( a25607a  and  a25604a );
 a25609a <=( a25608a  and  a25601a );
 a25613a <=( A167  and  (not A169) );
 a25614a <=( A170  and  a25613a );
 a25617a <=( A199  and  (not A166) );
 a25620a <=( A201  and  (not A200) );
 a25621a <=( a25620a  and  a25617a );
 a25622a <=( a25621a  and  a25614a );
 a25626a <=( (not A266)  and  A265 );
 a25627a <=( A203  and  a25626a );
 a25630a <=( A268  and  A267 );
 a25633a <=( A299  and  A298 );
 a25634a <=( a25633a  and  a25630a );
 a25635a <=( a25634a  and  a25627a );
 a25639a <=( A167  and  (not A169) );
 a25640a <=( A170  and  a25639a );
 a25643a <=( A199  and  (not A166) );
 a25646a <=( A201  and  (not A200) );
 a25647a <=( a25646a  and  a25643a );
 a25648a <=( a25647a  and  a25640a );
 a25652a <=( (not A266)  and  A265 );
 a25653a <=( A203  and  a25652a );
 a25656a <=( A268  and  A267 );
 a25659a <=( (not A299)  and  (not A298) );
 a25660a <=( a25659a  and  a25656a );
 a25661a <=( a25660a  and  a25653a );
 a25665a <=( A167  and  (not A169) );
 a25666a <=( A170  and  a25665a );
 a25669a <=( A199  and  (not A166) );
 a25672a <=( A201  and  (not A200) );
 a25673a <=( a25672a  and  a25669a );
 a25674a <=( a25673a  and  a25666a );
 a25678a <=( (not A266)  and  A265 );
 a25679a <=( A203  and  a25678a );
 a25682a <=( A269  and  A267 );
 a25685a <=( (not A300)  and  A298 );
 a25686a <=( a25685a  and  a25682a );
 a25687a <=( a25686a  and  a25679a );
 a25691a <=( A167  and  (not A169) );
 a25692a <=( A170  and  a25691a );
 a25695a <=( A199  and  (not A166) );
 a25698a <=( A201  and  (not A200) );
 a25699a <=( a25698a  and  a25695a );
 a25700a <=( a25699a  and  a25692a );
 a25704a <=( (not A266)  and  A265 );
 a25705a <=( A203  and  a25704a );
 a25708a <=( A269  and  A267 );
 a25711a <=( A299  and  A298 );
 a25712a <=( a25711a  and  a25708a );
 a25713a <=( a25712a  and  a25705a );
 a25717a <=( A167  and  (not A169) );
 a25718a <=( A170  and  a25717a );
 a25721a <=( A199  and  (not A166) );
 a25724a <=( A201  and  (not A200) );
 a25725a <=( a25724a  and  a25721a );
 a25726a <=( a25725a  and  a25718a );
 a25730a <=( (not A266)  and  A265 );
 a25731a <=( A203  and  a25730a );
 a25734a <=( A269  and  A267 );
 a25737a <=( (not A299)  and  (not A298) );
 a25738a <=( a25737a  and  a25734a );
 a25739a <=( a25738a  and  a25731a );
 a25743a <=( (not A167)  and  (not A169) );
 a25744a <=( A170  and  a25743a );
 a25747a <=( (not A200)  and  A166 );
 a25750a <=( (not A203)  and  (not A202) );
 a25751a <=( a25750a  and  a25747a );
 a25752a <=( a25751a  and  a25744a );
 a25756a <=( (not A269)  and  (not A268) );
 a25757a <=( (not A266)  and  a25756a );
 a25760a <=( (not A299)  and  A298 );
 a25763a <=( A301  and  A300 );
 a25764a <=( a25763a  and  a25760a );
 a25765a <=( a25764a  and  a25757a );
 a25769a <=( (not A167)  and  (not A169) );
 a25770a <=( A170  and  a25769a );
 a25773a <=( (not A200)  and  A166 );
 a25776a <=( (not A203)  and  (not A202) );
 a25777a <=( a25776a  and  a25773a );
 a25778a <=( a25777a  and  a25770a );
 a25782a <=( (not A269)  and  (not A268) );
 a25783a <=( (not A266)  and  a25782a );
 a25786a <=( (not A299)  and  A298 );
 a25789a <=( A302  and  A300 );
 a25790a <=( a25789a  and  a25786a );
 a25791a <=( a25790a  and  a25783a );
 a25795a <=( (not A167)  and  (not A169) );
 a25796a <=( A170  and  a25795a );
 a25799a <=( A199  and  A166 );
 a25802a <=( A201  and  (not A200) );
 a25803a <=( a25802a  and  a25799a );
 a25804a <=( a25803a  and  a25796a );
 a25808a <=( (not A266)  and  A265 );
 a25809a <=( A202  and  a25808a );
 a25812a <=( A268  and  A267 );
 a25815a <=( (not A300)  and  A298 );
 a25816a <=( a25815a  and  a25812a );
 a25817a <=( a25816a  and  a25809a );
 a25821a <=( (not A167)  and  (not A169) );
 a25822a <=( A170  and  a25821a );
 a25825a <=( A199  and  A166 );
 a25828a <=( A201  and  (not A200) );
 a25829a <=( a25828a  and  a25825a );
 a25830a <=( a25829a  and  a25822a );
 a25834a <=( (not A266)  and  A265 );
 a25835a <=( A202  and  a25834a );
 a25838a <=( A268  and  A267 );
 a25841a <=( A299  and  A298 );
 a25842a <=( a25841a  and  a25838a );
 a25843a <=( a25842a  and  a25835a );
 a25847a <=( (not A167)  and  (not A169) );
 a25848a <=( A170  and  a25847a );
 a25851a <=( A199  and  A166 );
 a25854a <=( A201  and  (not A200) );
 a25855a <=( a25854a  and  a25851a );
 a25856a <=( a25855a  and  a25848a );
 a25860a <=( (not A266)  and  A265 );
 a25861a <=( A202  and  a25860a );
 a25864a <=( A268  and  A267 );
 a25867a <=( (not A299)  and  (not A298) );
 a25868a <=( a25867a  and  a25864a );
 a25869a <=( a25868a  and  a25861a );
 a25873a <=( (not A167)  and  (not A169) );
 a25874a <=( A170  and  a25873a );
 a25877a <=( A199  and  A166 );
 a25880a <=( A201  and  (not A200) );
 a25881a <=( a25880a  and  a25877a );
 a25882a <=( a25881a  and  a25874a );
 a25886a <=( (not A266)  and  A265 );
 a25887a <=( A202  and  a25886a );
 a25890a <=( A269  and  A267 );
 a25893a <=( (not A300)  and  A298 );
 a25894a <=( a25893a  and  a25890a );
 a25895a <=( a25894a  and  a25887a );
 a25899a <=( (not A167)  and  (not A169) );
 a25900a <=( A170  and  a25899a );
 a25903a <=( A199  and  A166 );
 a25906a <=( A201  and  (not A200) );
 a25907a <=( a25906a  and  a25903a );
 a25908a <=( a25907a  and  a25900a );
 a25912a <=( (not A266)  and  A265 );
 a25913a <=( A202  and  a25912a );
 a25916a <=( A269  and  A267 );
 a25919a <=( A299  and  A298 );
 a25920a <=( a25919a  and  a25916a );
 a25921a <=( a25920a  and  a25913a );
 a25925a <=( (not A167)  and  (not A169) );
 a25926a <=( A170  and  a25925a );
 a25929a <=( A199  and  A166 );
 a25932a <=( A201  and  (not A200) );
 a25933a <=( a25932a  and  a25929a );
 a25934a <=( a25933a  and  a25926a );
 a25938a <=( (not A266)  and  A265 );
 a25939a <=( A202  and  a25938a );
 a25942a <=( A269  and  A267 );
 a25945a <=( (not A299)  and  (not A298) );
 a25946a <=( a25945a  and  a25942a );
 a25947a <=( a25946a  and  a25939a );
 a25951a <=( (not A167)  and  (not A169) );
 a25952a <=( A170  and  a25951a );
 a25955a <=( A199  and  A166 );
 a25958a <=( A201  and  (not A200) );
 a25959a <=( a25958a  and  a25955a );
 a25960a <=( a25959a  and  a25952a );
 a25964a <=( (not A266)  and  A265 );
 a25965a <=( A203  and  a25964a );
 a25968a <=( A268  and  A267 );
 a25971a <=( (not A300)  and  A298 );
 a25972a <=( a25971a  and  a25968a );
 a25973a <=( a25972a  and  a25965a );
 a25977a <=( (not A167)  and  (not A169) );
 a25978a <=( A170  and  a25977a );
 a25981a <=( A199  and  A166 );
 a25984a <=( A201  and  (not A200) );
 a25985a <=( a25984a  and  a25981a );
 a25986a <=( a25985a  and  a25978a );
 a25990a <=( (not A266)  and  A265 );
 a25991a <=( A203  and  a25990a );
 a25994a <=( A268  and  A267 );
 a25997a <=( A299  and  A298 );
 a25998a <=( a25997a  and  a25994a );
 a25999a <=( a25998a  and  a25991a );
 a26003a <=( (not A167)  and  (not A169) );
 a26004a <=( A170  and  a26003a );
 a26007a <=( A199  and  A166 );
 a26010a <=( A201  and  (not A200) );
 a26011a <=( a26010a  and  a26007a );
 a26012a <=( a26011a  and  a26004a );
 a26016a <=( (not A266)  and  A265 );
 a26017a <=( A203  and  a26016a );
 a26020a <=( A268  and  A267 );
 a26023a <=( (not A299)  and  (not A298) );
 a26024a <=( a26023a  and  a26020a );
 a26025a <=( a26024a  and  a26017a );
 a26029a <=( (not A167)  and  (not A169) );
 a26030a <=( A170  and  a26029a );
 a26033a <=( A199  and  A166 );
 a26036a <=( A201  and  (not A200) );
 a26037a <=( a26036a  and  a26033a );
 a26038a <=( a26037a  and  a26030a );
 a26042a <=( (not A266)  and  A265 );
 a26043a <=( A203  and  a26042a );
 a26046a <=( A269  and  A267 );
 a26049a <=( (not A300)  and  A298 );
 a26050a <=( a26049a  and  a26046a );
 a26051a <=( a26050a  and  a26043a );
 a26055a <=( (not A167)  and  (not A169) );
 a26056a <=( A170  and  a26055a );
 a26059a <=( A199  and  A166 );
 a26062a <=( A201  and  (not A200) );
 a26063a <=( a26062a  and  a26059a );
 a26064a <=( a26063a  and  a26056a );
 a26068a <=( (not A266)  and  A265 );
 a26069a <=( A203  and  a26068a );
 a26072a <=( A269  and  A267 );
 a26075a <=( A299  and  A298 );
 a26076a <=( a26075a  and  a26072a );
 a26077a <=( a26076a  and  a26069a );
 a26081a <=( (not A167)  and  (not A169) );
 a26082a <=( A170  and  a26081a );
 a26085a <=( A199  and  A166 );
 a26088a <=( A201  and  (not A200) );
 a26089a <=( a26088a  and  a26085a );
 a26090a <=( a26089a  and  a26082a );
 a26094a <=( (not A266)  and  A265 );
 a26095a <=( A203  and  a26094a );
 a26098a <=( A269  and  A267 );
 a26101a <=( (not A299)  and  (not A298) );
 a26102a <=( a26101a  and  a26098a );
 a26103a <=( a26102a  and  a26095a );
 a26107a <=( (not A168)  and  (not A169) );
 a26108a <=( (not A170)  and  a26107a );
 a26111a <=( (not A200)  and  A199 );
 a26114a <=( A202  and  A201 );
 a26115a <=( a26114a  and  a26111a );
 a26116a <=( a26115a  and  a26108a );
 a26120a <=( (not A269)  and  (not A268) );
 a26121a <=( (not A266)  and  a26120a );
 a26124a <=( (not A299)  and  A298 );
 a26127a <=( A301  and  A300 );
 a26128a <=( a26127a  and  a26124a );
 a26129a <=( a26128a  and  a26121a );
 a26133a <=( (not A168)  and  (not A169) );
 a26134a <=( (not A170)  and  a26133a );
 a26137a <=( (not A200)  and  A199 );
 a26140a <=( A202  and  A201 );
 a26141a <=( a26140a  and  a26137a );
 a26142a <=( a26141a  and  a26134a );
 a26146a <=( (not A269)  and  (not A268) );
 a26147a <=( (not A266)  and  a26146a );
 a26150a <=( (not A299)  and  A298 );
 a26153a <=( A302  and  A300 );
 a26154a <=( a26153a  and  a26150a );
 a26155a <=( a26154a  and  a26147a );
 a26159a <=( (not A168)  and  (not A169) );
 a26160a <=( (not A170)  and  a26159a );
 a26163a <=( (not A200)  and  A199 );
 a26166a <=( A203  and  A201 );
 a26167a <=( a26166a  and  a26163a );
 a26168a <=( a26167a  and  a26160a );
 a26172a <=( (not A269)  and  (not A268) );
 a26173a <=( (not A266)  and  a26172a );
 a26176a <=( (not A299)  and  A298 );
 a26179a <=( A301  and  A300 );
 a26180a <=( a26179a  and  a26176a );
 a26181a <=( a26180a  and  a26173a );
 a26185a <=( (not A168)  and  (not A169) );
 a26186a <=( (not A170)  and  a26185a );
 a26189a <=( (not A200)  and  A199 );
 a26192a <=( A203  and  A201 );
 a26193a <=( a26192a  and  a26189a );
 a26194a <=( a26193a  and  a26186a );
 a26198a <=( (not A269)  and  (not A268) );
 a26199a <=( (not A266)  and  a26198a );
 a26202a <=( (not A299)  and  A298 );
 a26205a <=( A302  and  A300 );
 a26206a <=( a26205a  and  a26202a );
 a26207a <=( a26206a  and  a26199a );
 a26211a <=( A167  and  (not A168) );
 a26212a <=( A169  and  a26211a );
 a26215a <=( A199  and  (not A166) );
 a26218a <=( A201  and  (not A200) );
 a26219a <=( a26218a  and  a26215a );
 a26220a <=( a26219a  and  a26212a );
 a26223a <=( (not A266)  and  A202 );
 a26226a <=( (not A269)  and  (not A268) );
 a26227a <=( a26226a  and  a26223a );
 a26230a <=( (not A299)  and  A298 );
 a26233a <=( A301  and  A300 );
 a26234a <=( a26233a  and  a26230a );
 a26235a <=( a26234a  and  a26227a );
 a26239a <=( A167  and  (not A168) );
 a26240a <=( A169  and  a26239a );
 a26243a <=( A199  and  (not A166) );
 a26246a <=( A201  and  (not A200) );
 a26247a <=( a26246a  and  a26243a );
 a26248a <=( a26247a  and  a26240a );
 a26251a <=( (not A266)  and  A202 );
 a26254a <=( (not A269)  and  (not A268) );
 a26255a <=( a26254a  and  a26251a );
 a26258a <=( (not A299)  and  A298 );
 a26261a <=( A302  and  A300 );
 a26262a <=( a26261a  and  a26258a );
 a26263a <=( a26262a  and  a26255a );
 a26267a <=( A167  and  (not A168) );
 a26268a <=( A169  and  a26267a );
 a26271a <=( A199  and  (not A166) );
 a26274a <=( A201  and  (not A200) );
 a26275a <=( a26274a  and  a26271a );
 a26276a <=( a26275a  and  a26268a );
 a26279a <=( (not A266)  and  A203 );
 a26282a <=( (not A269)  and  (not A268) );
 a26283a <=( a26282a  and  a26279a );
 a26286a <=( (not A299)  and  A298 );
 a26289a <=( A301  and  A300 );
 a26290a <=( a26289a  and  a26286a );
 a26291a <=( a26290a  and  a26283a );
 a26295a <=( A167  and  (not A168) );
 a26296a <=( A169  and  a26295a );
 a26299a <=( A199  and  (not A166) );
 a26302a <=( A201  and  (not A200) );
 a26303a <=( a26302a  and  a26299a );
 a26304a <=( a26303a  and  a26296a );
 a26307a <=( (not A266)  and  A203 );
 a26310a <=( (not A269)  and  (not A268) );
 a26311a <=( a26310a  and  a26307a );
 a26314a <=( (not A299)  and  A298 );
 a26317a <=( A302  and  A300 );
 a26318a <=( a26317a  and  a26314a );
 a26319a <=( a26318a  and  a26311a );
 a26323a <=( (not A167)  and  (not A168) );
 a26324a <=( A169  and  a26323a );
 a26327a <=( A199  and  A166 );
 a26330a <=( A201  and  (not A200) );
 a26331a <=( a26330a  and  a26327a );
 a26332a <=( a26331a  and  a26324a );
 a26335a <=( (not A266)  and  A202 );
 a26338a <=( (not A269)  and  (not A268) );
 a26339a <=( a26338a  and  a26335a );
 a26342a <=( (not A299)  and  A298 );
 a26345a <=( A301  and  A300 );
 a26346a <=( a26345a  and  a26342a );
 a26347a <=( a26346a  and  a26339a );
 a26351a <=( (not A167)  and  (not A168) );
 a26352a <=( A169  and  a26351a );
 a26355a <=( A199  and  A166 );
 a26358a <=( A201  and  (not A200) );
 a26359a <=( a26358a  and  a26355a );
 a26360a <=( a26359a  and  a26352a );
 a26363a <=( (not A266)  and  A202 );
 a26366a <=( (not A269)  and  (not A268) );
 a26367a <=( a26366a  and  a26363a );
 a26370a <=( (not A299)  and  A298 );
 a26373a <=( A302  and  A300 );
 a26374a <=( a26373a  and  a26370a );
 a26375a <=( a26374a  and  a26367a );
 a26379a <=( (not A167)  and  (not A168) );
 a26380a <=( A169  and  a26379a );
 a26383a <=( A199  and  A166 );
 a26386a <=( A201  and  (not A200) );
 a26387a <=( a26386a  and  a26383a );
 a26388a <=( a26387a  and  a26380a );
 a26391a <=( (not A266)  and  A203 );
 a26394a <=( (not A269)  and  (not A268) );
 a26395a <=( a26394a  and  a26391a );
 a26398a <=( (not A299)  and  A298 );
 a26401a <=( A301  and  A300 );
 a26402a <=( a26401a  and  a26398a );
 a26403a <=( a26402a  and  a26395a );
 a26407a <=( (not A167)  and  (not A168) );
 a26408a <=( A169  and  a26407a );
 a26411a <=( A199  and  A166 );
 a26414a <=( A201  and  (not A200) );
 a26415a <=( a26414a  and  a26411a );
 a26416a <=( a26415a  and  a26408a );
 a26419a <=( (not A266)  and  A203 );
 a26422a <=( (not A269)  and  (not A268) );
 a26423a <=( a26422a  and  a26419a );
 a26426a <=( (not A299)  and  A298 );
 a26429a <=( A302  and  A300 );
 a26430a <=( a26429a  and  a26426a );
 a26431a <=( a26430a  and  a26423a );
 a26435a <=( A167  and  A169 );
 a26436a <=( (not A170)  and  a26435a );
 a26439a <=( A199  and  A166 );
 a26442a <=( A201  and  (not A200) );
 a26443a <=( a26442a  and  a26439a );
 a26444a <=( a26443a  and  a26436a );
 a26447a <=( A265  and  A202 );
 a26450a <=( A267  and  (not A266) );
 a26451a <=( a26450a  and  a26447a );
 a26454a <=( A298  and  A268 );
 a26457a <=( (not A302)  and  (not A301) );
 a26458a <=( a26457a  and  a26454a );
 a26459a <=( a26458a  and  a26451a );
 a26463a <=( A167  and  A169 );
 a26464a <=( (not A170)  and  a26463a );
 a26467a <=( A199  and  A166 );
 a26470a <=( A201  and  (not A200) );
 a26471a <=( a26470a  and  a26467a );
 a26472a <=( a26471a  and  a26464a );
 a26475a <=( A265  and  A202 );
 a26478a <=( A267  and  (not A266) );
 a26479a <=( a26478a  and  a26475a );
 a26482a <=( A298  and  A269 );
 a26485a <=( (not A302)  and  (not A301) );
 a26486a <=( a26485a  and  a26482a );
 a26487a <=( a26486a  and  a26479a );
 a26491a <=( A167  and  A169 );
 a26492a <=( (not A170)  and  a26491a );
 a26495a <=( A199  and  A166 );
 a26498a <=( A201  and  (not A200) );
 a26499a <=( a26498a  and  a26495a );
 a26500a <=( a26499a  and  a26492a );
 a26503a <=( A265  and  A203 );
 a26506a <=( A267  and  (not A266) );
 a26507a <=( a26506a  and  a26503a );
 a26510a <=( A298  and  A268 );
 a26513a <=( (not A302)  and  (not A301) );
 a26514a <=( a26513a  and  a26510a );
 a26515a <=( a26514a  and  a26507a );
 a26519a <=( A167  and  A169 );
 a26520a <=( (not A170)  and  a26519a );
 a26523a <=( A199  and  A166 );
 a26526a <=( A201  and  (not A200) );
 a26527a <=( a26526a  and  a26523a );
 a26528a <=( a26527a  and  a26520a );
 a26531a <=( A265  and  A203 );
 a26534a <=( A267  and  (not A266) );
 a26535a <=( a26534a  and  a26531a );
 a26538a <=( A298  and  A269 );
 a26541a <=( (not A302)  and  (not A301) );
 a26542a <=( a26541a  and  a26538a );
 a26543a <=( a26542a  and  a26535a );
 a26547a <=( (not A167)  and  A169 );
 a26548a <=( (not A170)  and  a26547a );
 a26551a <=( A199  and  (not A166) );
 a26554a <=( A201  and  (not A200) );
 a26555a <=( a26554a  and  a26551a );
 a26556a <=( a26555a  and  a26548a );
 a26559a <=( A265  and  A202 );
 a26562a <=( A267  and  (not A266) );
 a26563a <=( a26562a  and  a26559a );
 a26566a <=( A298  and  A268 );
 a26569a <=( (not A302)  and  (not A301) );
 a26570a <=( a26569a  and  a26566a );
 a26571a <=( a26570a  and  a26563a );
 a26575a <=( (not A167)  and  A169 );
 a26576a <=( (not A170)  and  a26575a );
 a26579a <=( A199  and  (not A166) );
 a26582a <=( A201  and  (not A200) );
 a26583a <=( a26582a  and  a26579a );
 a26584a <=( a26583a  and  a26576a );
 a26587a <=( A265  and  A202 );
 a26590a <=( A267  and  (not A266) );
 a26591a <=( a26590a  and  a26587a );
 a26594a <=( A298  and  A269 );
 a26597a <=( (not A302)  and  (not A301) );
 a26598a <=( a26597a  and  a26594a );
 a26599a <=( a26598a  and  a26591a );
 a26603a <=( (not A167)  and  A169 );
 a26604a <=( (not A170)  and  a26603a );
 a26607a <=( A199  and  (not A166) );
 a26610a <=( A201  and  (not A200) );
 a26611a <=( a26610a  and  a26607a );
 a26612a <=( a26611a  and  a26604a );
 a26615a <=( A265  and  A203 );
 a26618a <=( A267  and  (not A266) );
 a26619a <=( a26618a  and  a26615a );
 a26622a <=( A298  and  A268 );
 a26625a <=( (not A302)  and  (not A301) );
 a26626a <=( a26625a  and  a26622a );
 a26627a <=( a26626a  and  a26619a );
 a26631a <=( (not A167)  and  A169 );
 a26632a <=( (not A170)  and  a26631a );
 a26635a <=( A199  and  (not A166) );
 a26638a <=( A201  and  (not A200) );
 a26639a <=( a26638a  and  a26635a );
 a26640a <=( a26639a  and  a26632a );
 a26643a <=( A265  and  A203 );
 a26646a <=( A267  and  (not A266) );
 a26647a <=( a26646a  and  a26643a );
 a26650a <=( A298  and  A269 );
 a26653a <=( (not A302)  and  (not A301) );
 a26654a <=( a26653a  and  a26650a );
 a26655a <=( a26654a  and  a26647a );
 a26659a <=( A167  and  (not A168) );
 a26660a <=( (not A169)  and  a26659a );
 a26663a <=( A199  and  A166 );
 a26666a <=( A201  and  (not A200) );
 a26667a <=( a26666a  and  a26663a );
 a26668a <=( a26667a  and  a26660a );
 a26671a <=( (not A266)  and  A202 );
 a26674a <=( (not A269)  and  (not A268) );
 a26675a <=( a26674a  and  a26671a );
 a26678a <=( (not A299)  and  A298 );
 a26681a <=( A301  and  A300 );
 a26682a <=( a26681a  and  a26678a );
 a26683a <=( a26682a  and  a26675a );
 a26687a <=( A167  and  (not A168) );
 a26688a <=( (not A169)  and  a26687a );
 a26691a <=( A199  and  A166 );
 a26694a <=( A201  and  (not A200) );
 a26695a <=( a26694a  and  a26691a );
 a26696a <=( a26695a  and  a26688a );
 a26699a <=( (not A266)  and  A202 );
 a26702a <=( (not A269)  and  (not A268) );
 a26703a <=( a26702a  and  a26699a );
 a26706a <=( (not A299)  and  A298 );
 a26709a <=( A302  and  A300 );
 a26710a <=( a26709a  and  a26706a );
 a26711a <=( a26710a  and  a26703a );
 a26715a <=( A167  and  (not A168) );
 a26716a <=( (not A169)  and  a26715a );
 a26719a <=( A199  and  A166 );
 a26722a <=( A201  and  (not A200) );
 a26723a <=( a26722a  and  a26719a );
 a26724a <=( a26723a  and  a26716a );
 a26727a <=( (not A266)  and  A203 );
 a26730a <=( (not A269)  and  (not A268) );
 a26731a <=( a26730a  and  a26727a );
 a26734a <=( (not A299)  and  A298 );
 a26737a <=( A301  and  A300 );
 a26738a <=( a26737a  and  a26734a );
 a26739a <=( a26738a  and  a26731a );
 a26743a <=( A167  and  (not A168) );
 a26744a <=( (not A169)  and  a26743a );
 a26747a <=( A199  and  A166 );
 a26750a <=( A201  and  (not A200) );
 a26751a <=( a26750a  and  a26747a );
 a26752a <=( a26751a  and  a26744a );
 a26755a <=( (not A266)  and  A203 );
 a26758a <=( (not A269)  and  (not A268) );
 a26759a <=( a26758a  and  a26755a );
 a26762a <=( (not A299)  and  A298 );
 a26765a <=( A302  and  A300 );
 a26766a <=( a26765a  and  a26762a );
 a26767a <=( a26766a  and  a26759a );
 a26771a <=( A167  and  (not A169) );
 a26772a <=( A170  and  a26771a );
 a26775a <=( A199  and  (not A166) );
 a26778a <=( A201  and  (not A200) );
 a26779a <=( a26778a  and  a26775a );
 a26780a <=( a26779a  and  a26772a );
 a26783a <=( A265  and  A202 );
 a26786a <=( A267  and  (not A266) );
 a26787a <=( a26786a  and  a26783a );
 a26790a <=( A298  and  A268 );
 a26793a <=( (not A302)  and  (not A301) );
 a26794a <=( a26793a  and  a26790a );
 a26795a <=( a26794a  and  a26787a );
 a26799a <=( A167  and  (not A169) );
 a26800a <=( A170  and  a26799a );
 a26803a <=( A199  and  (not A166) );
 a26806a <=( A201  and  (not A200) );
 a26807a <=( a26806a  and  a26803a );
 a26808a <=( a26807a  and  a26800a );
 a26811a <=( A265  and  A202 );
 a26814a <=( A267  and  (not A266) );
 a26815a <=( a26814a  and  a26811a );
 a26818a <=( A298  and  A269 );
 a26821a <=( (not A302)  and  (not A301) );
 a26822a <=( a26821a  and  a26818a );
 a26823a <=( a26822a  and  a26815a );
 a26827a <=( A167  and  (not A169) );
 a26828a <=( A170  and  a26827a );
 a26831a <=( A199  and  (not A166) );
 a26834a <=( A201  and  (not A200) );
 a26835a <=( a26834a  and  a26831a );
 a26836a <=( a26835a  and  a26828a );
 a26839a <=( A265  and  A203 );
 a26842a <=( A267  and  (not A266) );
 a26843a <=( a26842a  and  a26839a );
 a26846a <=( A298  and  A268 );
 a26849a <=( (not A302)  and  (not A301) );
 a26850a <=( a26849a  and  a26846a );
 a26851a <=( a26850a  and  a26843a );
 a26855a <=( A167  and  (not A169) );
 a26856a <=( A170  and  a26855a );
 a26859a <=( A199  and  (not A166) );
 a26862a <=( A201  and  (not A200) );
 a26863a <=( a26862a  and  a26859a );
 a26864a <=( a26863a  and  a26856a );
 a26867a <=( A265  and  A203 );
 a26870a <=( A267  and  (not A266) );
 a26871a <=( a26870a  and  a26867a );
 a26874a <=( A298  and  A269 );
 a26877a <=( (not A302)  and  (not A301) );
 a26878a <=( a26877a  and  a26874a );
 a26879a <=( a26878a  and  a26871a );
 a26883a <=( (not A167)  and  (not A169) );
 a26884a <=( A170  and  a26883a );
 a26887a <=( A199  and  A166 );
 a26890a <=( A201  and  (not A200) );
 a26891a <=( a26890a  and  a26887a );
 a26892a <=( a26891a  and  a26884a );
 a26895a <=( A265  and  A202 );
 a26898a <=( A267  and  (not A266) );
 a26899a <=( a26898a  and  a26895a );
 a26902a <=( A298  and  A268 );
 a26905a <=( (not A302)  and  (not A301) );
 a26906a <=( a26905a  and  a26902a );
 a26907a <=( a26906a  and  a26899a );
 a26911a <=( (not A167)  and  (not A169) );
 a26912a <=( A170  and  a26911a );
 a26915a <=( A199  and  A166 );
 a26918a <=( A201  and  (not A200) );
 a26919a <=( a26918a  and  a26915a );
 a26920a <=( a26919a  and  a26912a );
 a26923a <=( A265  and  A202 );
 a26926a <=( A267  and  (not A266) );
 a26927a <=( a26926a  and  a26923a );
 a26930a <=( A298  and  A269 );
 a26933a <=( (not A302)  and  (not A301) );
 a26934a <=( a26933a  and  a26930a );
 a26935a <=( a26934a  and  a26927a );
 a26939a <=( (not A167)  and  (not A169) );
 a26940a <=( A170  and  a26939a );
 a26943a <=( A199  and  A166 );
 a26946a <=( A201  and  (not A200) );
 a26947a <=( a26946a  and  a26943a );
 a26948a <=( a26947a  and  a26940a );
 a26951a <=( A265  and  A203 );
 a26954a <=( A267  and  (not A266) );
 a26955a <=( a26954a  and  a26951a );
 a26958a <=( A298  and  A268 );
 a26961a <=( (not A302)  and  (not A301) );
 a26962a <=( a26961a  and  a26958a );
 a26963a <=( a26962a  and  a26955a );
 a26967a <=( (not A167)  and  (not A169) );
 a26968a <=( A170  and  a26967a );
 a26971a <=( A199  and  A166 );
 a26974a <=( A201  and  (not A200) );
 a26975a <=( a26974a  and  a26971a );
 a26976a <=( a26975a  and  a26968a );
 a26979a <=( A265  and  A203 );
 a26982a <=( A267  and  (not A266) );
 a26983a <=( a26982a  and  a26979a );
 a26986a <=( A298  and  A269 );
 a26989a <=( (not A302)  and  (not A301) );
 a26990a <=( a26989a  and  a26986a );
 a26991a <=( a26990a  and  a26983a );


end x25_9x_behav;
