Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_16x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A39: buffer std_logic
);
end x25_16x;

architecture x25_16x_behav of x25_16x is
signal n_32,n_33,n_37,n_38,n_39,n_40,n_46,n_47,n_48,n_49,n_55,n_56,n_57,n_58,n_59,n_60,n_66,n_67,n_68,n_69,n_72,n_73,n_74,n_81,n_82,n_83,n_84,n_87,n_88,n_91,n_94,n_97,n_98,n_99,n_104,n_105,n_106,n_107,n_108,n_109,n_114,n_120,n_121,n_122,n_123,n_126,n_127,n_128,n_129,n_130,n_135,n_136,n_140,n_141,n_142,n_143,n_149,n_150,n_151,n_152,n_158,n_159,n_160,n_161,n_165,n_168,n_171,n_172,n_173,n_178,n_179,n_180,n_181,n_182,n_187,n_188,n_189,n_190,n_191,n_192,n_193,n_197,n_200,n_203,n_204,n_205,n_210,n_211,n_212,n_213,n_214,n_219,n_220,n_221,n_222,n_223,n_228,n_229,n_233,n_234,n_235,n_236,n_242,n_243,n_244,n_245,n_251,n_252,n_253,n_254,n_255,n_256,n_262,n_263,n_267,n_268,n_269,n_270,n_276,n_277,n_278,n_279,n_285,n_286,n_287,n_288,n_289,n_290,n_293,n_296,n_299,n_300,n_301,n_306,n_307,n_308,n_309,n_310,n_311,n_316,n_321,n_322,n_326,n_327,n_328,n_329,n_335,n_336,n_337,n_338,n_344,n_345,n_346,n_347,n_348,n_349,n_350,n_351,n_352,n_353,n_354,n_355,n_356,n_357,n_358: std_logic;
begin

A39 <=( (not n_358) );
 n_32 <=( (not A202)  and  A203 );
 n_33 <=( A200  and  n_32 );
 n_37 <=( A202  and  (not A203) );
 n_38 <=( (not A200)  and  n_37 );
 n_39 <=( n_38 ) or ( n_33 );
 n_40 <=( (not A199)  and  n_39 );
 n_46 <=( A202  and  (not A203) );
 n_47 <=( A199  and  n_46 );
 n_48 <=( n_47 ) or ( A201 );
 n_49 <=( A200  and  n_48 );
 n_55 <=( (not A202)  and  A203 );
 n_56 <=( (not A200)  and  n_55 );
 n_57 <=( n_56 ) or ( A201 );
 n_58 <=( A199  and  n_57 );
 n_59 <=( n_58 ) or ( n_49 );
 n_60 <=( n_59 ) or ( n_40 );
 n_66 <=( A170 ) or ( A169 );
 n_67 <=( A168  and  n_66 );
 n_68 <=( (not A167)  and  n_67 );
 n_69 <=( A166  and  n_68 );
 n_72 <=( (not A166)  and  A167 );
 n_73 <=( n_72 ) or ( n_69 );
 n_74 <=( n_60  and  n_73 );
 n_81 <=( (not A169)  and  (not A170) );
 n_82 <=( n_81 ) or ( (not A168) );
 n_83 <=( n_82 ) or ( (not A166) );
 n_84 <=( (not A167)  and  n_83 );
 n_87 <=( A166  and  A167 );
 n_88 <=( n_87 ) or ( n_84 );
 n_91 <=( (not A203) ) or ( A202 );
 n_94 <=( (not A199)  and  A200 );
 n_97 <=( A199  and  (not A200) );
 n_98 <=( n_97 ) or ( n_94 );
 n_99 <=( n_91  and  n_98 );
 n_104 <=( A203 ) or ( (not A202) );
 n_105 <=( A200  and  n_104 );
 n_106 <=( A199  and  n_105 );
 n_107 <=( n_106 ) or ( n_99 );
 n_108 <=( n_88  and  n_107 );
 n_109 <=( (not A201)  and  n_108 );
 n_114 <=( A203 ) or ( (not A202) );
 n_120 <=( (not A169)  and  (not A170) );
 n_121 <=( n_120 ) or ( (not A168) );
 n_122 <=( n_121 ) or ( (not A166) );
 n_123 <=( (not A167)  and  n_122 );
 n_126 <=( A166  and  A167 );
 n_127 <=( n_126 ) or ( n_123 );
 n_128 <=( n_114  and  n_127 );
 n_129 <=( (not A200)  and  n_128 );
 n_130 <=( (not A199)  and  n_129 );
 n_135 <=( (not A268)  and  A269 );
 n_136 <=( A266  and  n_135 );
 n_140 <=( A268  and  (not A269) );
 n_141 <=( (not A266)  and  n_140 );
 n_142 <=( n_141 ) or ( n_136 );
 n_143 <=( (not A265)  and  n_142 );
 n_149 <=( A268  and  (not A269) );
 n_150 <=( A265  and  n_149 );
 n_151 <=( n_150 ) or ( A267 );
 n_152 <=( A266  and  n_151 );
 n_158 <=( (not A268)  and  A269 );
 n_159 <=( (not A266)  and  n_158 );
 n_160 <=( n_159 ) or ( A267 );
 n_161 <=( A265  and  n_160 );
 n_165 <=( (not A302) ) or ( A301 );
 n_168 <=( (not A298)  and  A299 );
 n_171 <=( A298  and  (not A299) );
 n_172 <=( n_171 ) or ( n_168 );
 n_173 <=( n_165  and  n_172 );
 n_178 <=( A302 ) or ( (not A301) );
 n_179 <=( A299  and  n_178 );
 n_180 <=( A298  and  n_179 );
 n_181 <=( n_180 ) or ( n_173 );
 n_182 <=( (not A300)  and  n_181 );
 n_187 <=( A302 ) or ( (not A301) );
 n_188 <=( (not A299)  and  n_187 );
 n_189 <=( (not A298)  and  n_188 );
 n_190 <=( n_189 ) or ( n_182 );
 n_191 <=( n_190 ) or ( n_161 );
 n_192 <=( n_191 ) or ( n_152 );
 n_193 <=( n_192 ) or ( n_143 );
 n_197 <=( (not A236) ) or ( A235 );
 n_200 <=( (not A232)  and  A233 );
 n_203 <=( A232  and  (not A233) );
 n_204 <=( n_203 ) or ( n_200 );
 n_205 <=( n_197  and  n_204 );
 n_210 <=( A236 ) or ( (not A235) );
 n_211 <=( A233  and  n_210 );
 n_212 <=( A232  and  n_211 );
 n_213 <=( n_212 ) or ( n_205 );
 n_214 <=( (not A234)  and  n_213 );
 n_219 <=( A236 ) or ( (not A235) );
 n_220 <=( (not A233)  and  n_219 );
 n_221 <=( (not A232)  and  n_220 );
 n_222 <=( n_221 ) or ( n_214 );
 n_223 <=( n_193  and  n_222 );
 n_228 <=( (not A301)  and  A302 );
 n_229 <=( A299  and  n_228 );
 n_233 <=( A301  and  (not A302) );
 n_234 <=( (not A299)  and  n_233 );
 n_235 <=( n_234 ) or ( n_229 );
 n_236 <=( (not A298)  and  n_235 );
 n_242 <=( A301  and  (not A302) );
 n_243 <=( A298  and  n_242 );
 n_244 <=( n_243 ) or ( A300 );
 n_245 <=( A299  and  n_244 );
 n_251 <=( (not A301)  and  A302 );
 n_252 <=( (not A299)  and  n_251 );
 n_253 <=( n_252 ) or ( A300 );
 n_254 <=( A298  and  n_253 );
 n_255 <=( n_254 ) or ( n_245 );
 n_256 <=( n_255 ) or ( n_236 );
 n_262 <=( (not A235)  and  A236 );
 n_263 <=( A233  and  n_262 );
 n_267 <=( A235  and  (not A236) );
 n_268 <=( (not A233)  and  n_267 );
 n_269 <=( n_268 ) or ( n_263 );
 n_270 <=( (not A232)  and  n_269 );
 n_276 <=( A235  and  (not A236) );
 n_277 <=( A232  and  n_276 );
 n_278 <=( n_277 ) or ( A234 );
 n_279 <=( A233  and  n_278 );
 n_285 <=( (not A235)  and  A236 );
 n_286 <=( (not A233)  and  n_285 );
 n_287 <=( n_286 ) or ( A234 );
 n_288 <=( A232  and  n_287 );
 n_289 <=( n_288 ) or ( n_279 );
 n_290 <=( n_289 ) or ( n_270 );
 n_293 <=( (not A269) ) or ( A268 );
 n_296 <=( (not A265)  and  A266 );
 n_299 <=( A265  and  (not A266) );
 n_300 <=( n_299 ) or ( n_296 );
 n_301 <=( n_293  and  n_300 );
 n_306 <=( A269 ) or ( (not A268) );
 n_307 <=( A266  and  n_306 );
 n_308 <=( A265  and  n_307 );
 n_309 <=( n_308 ) or ( n_301 );
 n_310 <=( n_290  and  n_309 );
 n_311 <=( (not A267)  and  n_310 );
 n_316 <=( A269 ) or ( (not A268) );
 n_321 <=( (not A235)  and  A236 );
 n_322 <=( A233  and  n_321 );
 n_326 <=( A235  and  (not A236) );
 n_327 <=( (not A233)  and  n_326 );
 n_328 <=( n_327 ) or ( n_322 );
 n_329 <=( (not A232)  and  n_328 );
 n_335 <=( A235  and  (not A236) );
 n_336 <=( A232  and  n_335 );
 n_337 <=( n_336 ) or ( A234 );
 n_338 <=( A233  and  n_337 );
 n_344 <=( (not A235)  and  A236 );
 n_345 <=( (not A233)  and  n_344 );
 n_346 <=( n_345 ) or ( A234 );
 n_347 <=( A232  and  n_346 );
 n_348 <=( n_347 ) or ( n_338 );
 n_349 <=( n_348 ) or ( n_329 );
 n_350 <=( n_316  and  n_349 );
 n_351 <=( (not A266)  and  n_350 );
 n_352 <=( (not A265)  and  n_351 );
 n_353 <=( n_352 ) or ( n_311 );
 n_354 <=( n_256  and  n_353 );
 n_355 <=( n_354 ) or ( n_223 );
 n_356 <=( n_355 ) or ( n_130 );
 n_357 <=( n_356 ) or ( n_109 );
 n_358 <=( n_357 ) or ( n_74 );


end x25_16x_behav;
