Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_4x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A139: buffer std_logic
);
end x25_4x;

architecture x25_4x_behav of x25_4x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2196a,a2197a,a2198a,a2199a,a2200a,a2201a,a2202a,a2203a,a2204a,a2205a,a2206a,a2207a,a2208a,a2209a,a2210a,a2211a,a2212a,a2213a,a2214a,a2215a,a2216a,a2217a,a2218a,a2219a,a2220a,a2221a,a2222a,a2223a,a2224a,a2225a,a2226a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2237a,a2238a,a2239a,a2240a,a2241a,a2242a,a2243a,a2244a,a2245a,a2246a,a2247a,a2248a,a2249a,a2250a,a2251a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2258a,a2259a,a2260a,a2261a,a2262a,a2263a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2271a,a2272a,a2273a,a2274a,a2275a,a2276a,a2277a,a2278a,a2279a,a2280a,a2281a,a2282a,a2283a,a2284a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2297a,a2298a,a2299a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2306a,a2307a,a2308a,a2309a,a2310a,a2311a,a2312a,a2313a,a2314a,a2315a,a2316a,a2317a,a2318a,a2319a,a2320a,a2321a,a2322a,a2323a,a2324a,a2325a,a2326a,a2327a,a2328a,a2329a,a2330a,a2331a,a2332a,a2333a,a2334a,a2335a,a2336a,a2337a,a2338a,a2339a,a2340a,a2341a,a2342a,a2343a,a2344a,a2345a,a2346a,a2347a,a2348a,a2349a,a2350a,a2351a,a2352a,a2353a,a2354a,a2355a,a2356a,a2357a,a2358a,a2359a,a2360a,a2361a,a2362a,a2363a,a2364a,a2365a,a2366a,a2367a,a2368a,a2369a,a2370a,a2371a,a2372a,a2373a,a2374a,a2375a,a2376a,a2377a,a2378a,a2379a,a2380a,a2381a,a2382a,a2383a,a2384a,a2385a,a2386a,a2387a,a2388a,a2389a,a2390a,a2391a,a2392a,a2393a,a2394a,a2395a,a2396a,a2397a,a2398a,a2399a,a2400a,a2401a,a2402a,a2403a,a2404a,a2405a,a2406a,a2407a,a2408a,a2409a,a2410a,a2411a,a2412a,a2413a,a2414a,a2415a,a2416a,a2417a,a2418a,a2419a,a2420a,a2421a,a2422a,a2423a,a2424a,a2425a,a2426a,a2427a,a2428a,a2429a,a2430a,a2431a,a2432a,a2433a,a2434a,a2435a,a2436a,a2437a,a2438a,a2439a,a2440a,a2441a,a2442a,a2443a,a2444a,a2445a,a2446a,a2447a,a2448a,a2449a,a2450a,a2451a,a2452a,a2453a,a2454a,a2455a,a2456a,a2457a,a2458a,a2459a,a2460a,a2461a,a2462a,a2463a,a2464a,a2465a,a2466a,a2467a,a2468a,a2469a,a2470a,a2471a,a2472a,a2473a,a2474a,a2475a,a2476a,a2477a,a2478a,a2479a,a2480a,a2481a,a2482a,a2483a,a2484a,a2485a,a2486a,a2487a,a2488a,a2489a,a2490a,a2491a,a2492a,a2493a,a2494a,a2495a,a2496a,a2497a,a2498a,a2499a,a2500a,a2501a,a2502a,a2503a,a2504a,a2505a,a2506a,a2507a,a2508a,a2509a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2516a,a2517a,a2518a,a2519a,a2520a,a2521a,a2522a,a2523a,a2524a,a2525a,a2526a,a2527a,a2528a,a2529a,a2530a,a2531a,a2532a,a2533a,a2534a,a2535a,a2536a,a2537a,a2538a,a2539a,a2540a,a2541a,a2542a,a2543a,a2544a,a2545a,a2546a,a2547a,a2548a,a2549a,a2550a,a2551a,a2552a,a2553a,a2554a,a2555a,a2556a,a2557a,a2558a,a2559a,a2560a,a2561a,a2562a,a2563a,a2564a,a2565a,a2566a,a2567a,a2568a,a2569a,a2570a,a2571a,a2572a,a2573a,a2574a,a2575a,a2576a,a2577a,a2578a,a2579a,a2580a,a2581a,a2582a,a2583a,a2584a,a2585a,a2586a,a2587a,a2588a,a2589a,a2590a,a2591a,a2592a,a2593a,a2594a,a2595a,a2596a,a2597a,a2598a,a2599a,a2600a,a2601a,a2602a,a2603a,a2604a,a2605a,a2606a,a2607a,a2608a,a2609a,a2610a,a2611a,a2612a,a2613a,a2614a,a2615a,a2616a,a2617a,a2618a,a2619a,a2620a,a2621a,a2622a,a2623a,a2624a,a2625a,a2626a,a2627a,a2628a,a2629a,a2630a,a2631a,a2632a,a2633a,a2634a,a2635a,a2636a,a2637a,a2638a,a2639a,a2640a,a2641a,a2642a,a2643a,a2644a,a2645a,a2646a,a2647a,a2648a,a2649a,a2650a,a2651a,a2652a,a2653a,a2654a,a2655a,a2656a,a2657a,a2658a,a2659a,a2660a,a2661a,a2662a,a2663a,a2664a,a2665a,a2666a,a2667a,a2668a,a2669a,a2670a,a2671a,a2672a,a2673a,a2674a,a2675a,a2676a,a2677a,a2678a,a2679a,a2680a,a2681a,a2682a,a2683a,a2684a,a2685a,a2686a,a2687a,a2688a,a2689a,a2690a,a2691a,a2692a,a2693a,a2694a,a2695a,a2696a,a2697a,a2698a,a2699a,a2700a,a2701a,a2702a,a2703a,a2704a,a2705a,a2706a,a2707a,a2708a,a2709a,a2710a,a2711a,a2712a,a2713a,a2714a,a2715a,a2716a,a2717a,a2718a,a2719a,a2720a,a2721a,a2722a,a2723a,a2724a,a2725a,a2726a,a2727a,a2728a,a2729a,a2730a,a2731a,a2732a,a2733a,a2734a,a2735a,a2736a,a2737a,a2738a,a2739a,a2740a,a2741a,a2742a,a2743a,a2744a,a2745a,a2746a,a2747a,a2748a,a2749a,a2750a,a2751a,a2752a,a2753a,a2754a,a2755a,a2756a,a2757a,a2758a,a2759a,a2760a,a2761a,a2762a,a2763a,a2764a,a2765a,a2766a,a2767a,a2768a,a2769a,a2770a,a2771a,a2772a,a2773a,a2774a,a2775a,a2776a,a2777a,a2778a,a2779a,a2780a,a2781a,a2782a,a2783a,a2784a,a2785a,a2786a,a2787a,a2788a,a2789a,a2790a,a2791a,a2792a,a2793a,a2794a,a2795a,a2796a,a2797a,a2798a,a2799a,a2800a,a2801a,a2802a,a2803a,a2804a,a2805a,a2806a,a2807a,a2808a,a2809a,a2810a,a2811a,a2812a,a2813a,a2814a,a2815a,a2816a,a2817a,a2818a,a2819a,a2820a,a2821a,a2822a,a2823a,a2824a,a2825a,a2826a,a2827a,a2828a,a2829a,a2830a,a2831a,a2832a,a2833a,a2834a,a2835a,a2836a,a2837a,a2838a,a2839a,a2840a,a2841a,a2842a,a2843a,a2844a,a2845a,a2846a,a2847a,a2848a,a2849a,a2850a,a2851a,a2852a,a2853a,a2854a,a2855a,a2856a,a2857a,a2858a,a2859a,a2860a,a2861a,a2862a,a2863a,a2864a,a2865a,a2866a,a2867a,a2868a,a2869a,a2870a,a2871a,a2872a,a2873a,a2874a,a2875a,a2876a,a2877a,a2878a,a2879a,a2880a,a2881a,a2882a,a2883a,a2884a,a2885a,a2886a,a2887a,a2888a,a2889a,a2890a,a2891a,a2892a,a2893a,a2894a,a2895a,a2896a,a2897a,a2898a,a2899a,a2900a,a2901a,a2902a,a2903a,a2904a,a2905a,a2906a,a2907a,a2908a,a2909a,a2910a,a2911a,a2912a,a2913a,a2914a,a2915a,a2916a,a2917a,a2918a,a2919a,a2920a,a2921a,a2922a,a2923a,a2924a,a2925a,a2926a,a2927a,a2928a,a2929a,a2930a,a2931a,a2932a,a2933a,a2934a,a2935a,a2936a,a2937a,a2938a,a2939a,a2940a,a2941a,a2942a,a2943a,a2944a,a2945a,a2946a,a2947a,a2948a,a2949a,a2950a,a2951a,a2952a,a2953a,a2954a,a2955a,a2956a,a2957a,a2958a,a2959a,a2960a,a2961a,a2962a,a2963a,a2964a,a2965a,a2966a,a2967a,a2968a,a2969a,a2970a,a2971a,a2972a,a2973a,a2974a,a2975a,a2976a,a2977a,a2978a,a2979a,a2980a,a2981a,a2982a,a2983a,a2984a,a2985a,a2986a,a2987a,a2988a,a2989a,a2990a,a2991a,a2992a,a2993a,a2994a,a2995a,a2996a,a2997a,a2998a,a2999a,a3000a,a3001a,a3002a,a3003a,a3004a,a3005a,a3006a,a3007a,a3008a,a3009a,a3010a,a3011a,a3012a,a3013a,a3014a,a3015a,a3016a,a3017a,a3018a,a3019a,a3020a,a3021a,a3022a,a3023a,a3024a,a3025a,a3026a,a3027a,a3028a,a3029a,a3030a,a3031a,a3032a,a3033a,a3034a,a3035a,a3036a,a3037a,a3038a,a3039a,a3040a,a3041a,a3042a,a3043a,a3044a,a3045a,a3046a,a3047a,a3048a,a3049a,a3050a,a3051a,a3052a,a3053a,a3054a,a3055a,a3056a,a3057a,a3058a,a3059a,a3060a,a3061a,a3062a,a3063a,a3064a,a3065a,a3066a,a3067a,a3068a,a3069a,a3070a,a3071a,a3072a,a3073a,a3074a,a3075a,a3076a,a3077a,a3078a,a3079a,a3080a,a3081a,a3082a,a3083a,a3084a,a3085a,a3086a,a3087a,a3088a,a3089a,a3090a,a3091a,a3092a,a3093a,a3094a,a3095a,a3096a,a3097a,a3098a,a3099a,a3100a,a3101a,a3102a,a3103a,a3104a,a3105a,a3106a,a3107a,a3108a,a3109a,a3110a,a3111a,a3112a,a3113a,a3114a,a3115a,a3116a,a3117a,a3118a,a3119a,a3120a,a3121a,a3122a,a3123a,a3124a,a3125a,a3126a,a3127a,a3128a,a3129a,a3130a,a3131a,a3132a,a3133a,a3134a,a3135a,a3136a,a3137a,a3138a,a3139a,a3140a,a3141a,a3142a,a3143a,a3144a,a3145a,a3146a,a3147a,a3148a,a3149a,a3150a,a3151a,a3152a,a3153a,a3154a,a3155a,a3156a,a3157a,a3158a,a3159a,a3160a,a3161a,a3162a,a3163a,a3164a,a3165a,a3166a,a3167a,a3168a,a3169a,a3170a,a3171a,a3172a,a3173a,a3174a,a3175a,a3176a,a3177a,a3178a,a3179a,a3180a,a3181a,a3182a,a3183a,a3184a,a3185a,a3186a,a3187a,a3188a,a3189a,a3190a,a3191a,a3192a,a3193a,a3194a,a3195a,a3196a,a3197a,a3198a,a3199a,a3200a,a3201a,a3202a,a3203a,a3204a,a3205a,a3206a,a3207a,a3208a,a3209a,a3210a,a3211a,a3212a,a3213a,a3214a,a3215a,a3216a,a3217a,a3218a,a3219a,a3220a,a3221a,a3222a,a3223a,a3224a,a3225a,a3226a,a3227a,a3228a,a3229a,a3230a,a3231a,a3232a,a3233a,a3234a,a3235a,a3236a,a3237a,a3238a,a3239a,a3240a,a3241a,a3242a,a3243a,a3244a,a3245a,a3246a,a3247a,a3248a,a3249a,a3250a,a3251a,a3252a,a3253a,a3254a,a3255a,a3256a,a3257a,a3258a,a3259a,a3260a,a3261a,a3262a,a3263a,a3264a,a3265a,a3266a,a3267a,a3268a,a3269a,a3270a,a3271a,a3272a,a3273a,a3274a,a3275a,a3276a,a3277a,a3278a,a3279a,a3280a,a3281a,a3282a,a3283a,a3284a,a3285a,a3286a,a3287a,a3288a,a3289a,a3290a,a3291a,a3292a,a3293a,a3294a,a3295a,a3296a,a3297a,a3298a,a3299a,a3300a,a3301a,a3302a,a3303a,a3304a,a3305a,a3306a,a3307a,a3308a,a3309a,a3310a,a3311a,a3312a,a3313a,a3314a,a3315a,a3316a,a3317a,a3318a,a3319a,a3320a,a3321a,a3322a,a3323a,a3324a,a3325a,a3326a,a3327a,a3328a,a3329a,a3330a,a3331a,a3332a,a3333a,a3334a,a3335a,a3336a,a3337a,a3338a,a3339a,a3340a,a3341a,a3342a,a3343a,a3344a,a3345a,a3346a,a3347a,a3348a,a3349a,a3350a,a3351a,a3352a,a3353a,a3354a,a3355a,a3356a,a3357a,a3358a,a3359a,a3360a,a3361a,a3362a,a3363a,a3364a,a3365a,a3366a,a3367a,a3368a,a3369a,a3370a,a3371a,a3372a,a3373a,a3374a,a3375a,a3376a,a3377a,a3378a,a3379a,a3380a,a3381a,a3382a,a3383a,a3384a,a3385a,a3386a,a3387a,a3388a,a3389a,a3390a,a3391a,a3392a,a3393a,a3394a,a3395a,a3396a,a3397a,a3398a,a3399a,a3400a,a3401a,a3402a,a3403a,a3404a,a3405a,a3406a,a3407a,a3408a,a3409a,a3410a,a3411a,a3412a,a3413a,a3414a,a3415a,a3416a,a3417a,a3418a,a3419a,a3420a,a3421a,a3422a,a3423a,a3424a,a3425a,a3426a,a3427a,a3428a,a3429a,a3430a,a3431a,a3432a,a3433a,a3434a,a3435a,a3436a,a3437a,a3438a,a3439a,a3440a,a3441a,a3442a,a3443a,a3444a,a3445a,a3446a,a3447a,a3448a,a3449a,a3450a,a3451a,a3452a,a3453a,a3454a,a3455a,a3456a,a3457a,a3458a,a3459a,a3460a,a3461a,a3462a,a3463a,a3464a,a3465a,a3466a,a3467a,a3468a,a3469a,a3470a,a3471a,a3472a,a3473a,a3474a,a3475a,a3476a,a3477a,a3478a,a3479a,a3480a,a3481a,a3482a,a3483a,a3484a,a3485a,a3486a,a3487a,a3488a,a3489a,a3490a,a3491a,a3492a,a3493a,a3494a,a3495a,a3496a,a3497a,a3498a,a3499a,a3500a,a3501a,a3502a,a3503a,a3504a,a3505a,a3506a,a3507a,a3508a,a3509a,a3510a,a3511a,a3512a,a3513a,a3514a,a3515a,a3516a,a3517a,a3518a,a3519a,a3520a,a3521a,a3522a,a3523a,a3524a,a3525a,a3526a,a3527a,a3528a,a3529a,a3530a,a3531a,a3532a,a3533a,a3534a,a3535a,a3536a,a3537a,a3538a,a3539a,a3540a,a3541a,a3542a,a3543a,a3544a,a3545a,a3546a,a3547a,a3548a,a3549a,a3550a,a3551a,a3552a,a3553a,a3554a,a3555a,a3556a,a3557a,a3558a,a3559a,a3560a,a3561a,a3562a,a3563a,a3564a,a3565a,a3566a,a3567a,a3568a,a3569a,a3570a,a3571a,a3572a,a3573a,a3574a,a3575a,a3576a,a3577a,a3578a,a3579a,a3580a,a3581a,a3582a,a3583a,a3584a,a3585a,a3586a,a3587a,a3588a,a3589a,a3590a,a3591a,a3592a,a3593a,a3594a,a3595a,a3596a,a3597a,a3598a,a3599a,a3600a,a3601a,a3602a,a3603a,a3604a,a3605a,a3606a,a3607a,a3608a,a3609a,a3610a,a3611a,a3612a,a3613a,a3614a,a3615a,a3616a,a3617a,a3618a,a3619a,a3620a,a3621a,a3622a,a3623a,a3624a,a3625a,a3626a,a3627a,a3628a,a3629a,a3630a,a3631a,a3632a,a3633a,a3634a,a3635a,a3636a,a3637a,a3638a,a3639a,a3640a,a3641a,a3642a,a3643a,a3644a,a3645a,a3646a,a3647a,a3648a,a3649a,a3650a,a3651a,a3652a,a3653a,a3654a,a3655a,a3656a,a3657a,a3658a,a3659a,a3660a,a3661a,a3662a,a3663a,a3664a,a3665a,a3666a,a3667a,a3668a,a3669a,a3670a,a3671a,a3672a,a3673a,a3674a,a3675a,a3676a,a3677a,a3678a,a3679a,a3680a,a3681a,a3682a,a3683a,a3684a,a3685a,a3686a,a3687a,a3688a,a3689a,a3690a,a3691a,a3692a,a3693a,a3694a,a3695a,a3696a,a3697a,a3698a,a3699a,a3700a,a3701a,a3702a,a3706a,a3707a,a3710a,a3713a,a3714a,a3715a,a3719a,a3720a,a3723a,a3726a,a3727a,a3728a,a3729a,a3733a,a3734a,a3737a,a3740a,a3741a,a3742a,a3746a,a3747a,a3750a,a3753a,a3754a,a3755a,a3756a,a3757a,a3761a,a3762a,a3765a,a3768a,a3769a,a3770a,a3774a,a3775a,a3778a,a3781a,a3782a,a3783a,a3784a,a3788a,a3789a,a3792a,a3795a,a3796a,a3797a,a3800a,a3803a,a3804a,a3807a,a3810a,a3811a,a3812a,a3813a,a3814a,a3815a,a3819a,a3820a,a3823a,a3826a,a3827a,a3828a,a3832a,a3833a,a3836a,a3839a,a3840a,a3841a,a3842a,a3846a,a3847a,a3850a,a3853a,a3854a,a3855a,a3858a,a3861a,a3862a,a3865a,a3868a,a3869a,a3870a,a3871a,a3872a,a3876a,a3877a,a3880a,a3883a,a3884a,a3885a,a3889a,a3890a,a3893a,a3896a,a3897a,a3898a,a3899a,a3903a,a3904a,a3907a,a3910a,a3911a,a3912a,a3915a,a3918a,a3919a,a3922a,a3925a,a3926a,a3927a,a3928a,a3929a,a3930a,a3931a,a3935a,a3936a,a3939a,a3942a,a3943a,a3944a,a3948a,a3949a,a3952a,a3955a,a3956a,a3957a,a3958a,a3962a,a3963a,a3966a,a3969a,a3970a,a3971a,a3974a,a3977a,a3978a,a3981a,a3984a,a3985a,a3986a,a3987a,a3988a,a3992a,a3993a,a3996a,a3999a,a4000a,a4001a,a4005a,a4006a,a4009a,a4012a,a4013a,a4014a,a4015a,a4019a,a4020a,a4023a,a4026a,a4027a,a4028a,a4031a,a4034a,a4035a,a4038a,a4041a,a4042a,a4043a,a4044a,a4045a,a4046a,a4050a,a4051a,a4054a,a4057a,a4058a,a4059a,a4063a,a4064a,a4067a,a4070a,a4071a,a4072a,a4073a,a4077a,a4078a,a4081a,a4084a,a4085a,a4086a,a4089a,a4092a,a4093a,a4096a,a4099a,a4100a,a4101a,a4102a,a4103a,a4107a,a4108a,a4111a,a4114a,a4115a,a4116a,a4120a,a4121a,a4124a,a4127a,a4128a,a4129a,a4130a,a4134a,a4135a,a4138a,a4141a,a4142a,a4143a,a4146a,a4149a,a4150a,a4153a,a4156a,a4157a,a4158a,a4159a,a4160a,a4161a,a4162a,a4163a,a4167a,a4168a,a4171a,a4174a,a4175a,a4176a,a4180a,a4181a,a4184a,a4187a,a4188a,a4189a,a4190a,a4194a,a4195a,a4198a,a4201a,a4202a,a4203a,a4207a,a4208a,a4211a,a4214a,a4215a,a4216a,a4217a,a4218a,a4222a,a4223a,a4226a,a4229a,a4230a,a4231a,a4235a,a4236a,a4239a,a4242a,a4243a,a4244a,a4245a,a4249a,a4250a,a4253a,a4256a,a4257a,a4258a,a4261a,a4264a,a4265a,a4268a,a4271a,a4272a,a4273a,a4274a,a4275a,a4276a,a4280a,a4281a,a4284a,a4287a,a4288a,a4289a,a4293a,a4294a,a4297a,a4300a,a4301a,a4302a,a4303a,a4307a,a4308a,a4311a,a4314a,a4315a,a4316a,a4319a,a4322a,a4323a,a4326a,a4329a,a4330a,a4331a,a4332a,a4333a,a4337a,a4338a,a4341a,a4344a,a4345a,a4346a,a4350a,a4351a,a4354a,a4357a,a4358a,a4359a,a4360a,a4364a,a4365a,a4368a,a4371a,a4372a,a4373a,a4376a,a4379a,a4380a,a4383a,a4386a,a4387a,a4388a,a4389a,a4390a,a4391a,a4392a,a4396a,a4397a,a4400a,a4403a,a4404a,a4405a,a4409a,a4410a,a4413a,a4416a,a4417a,a4418a,a4419a,a4423a,a4424a,a4427a,a4430a,a4431a,a4432a,a4435a,a4438a,a4439a,a4442a,a4445a,a4446a,a4447a,a4448a,a4449a,a4453a,a4454a,a4457a,a4460a,a4461a,a4462a,a4466a,a4467a,a4470a,a4473a,a4474a,a4475a,a4476a,a4480a,a4481a,a4484a,a4487a,a4488a,a4489a,a4492a,a4495a,a4496a,a4499a,a4502a,a4503a,a4504a,a4505a,a4506a,a4507a,a4511a,a4512a,a4515a,a4518a,a4519a,a4520a,a4524a,a4525a,a4528a,a4531a,a4532a,a4533a,a4534a,a4538a,a4539a,a4542a,a4545a,a4546a,a4547a,a4550a,a4553a,a4554a,a4557a,a4560a,a4561a,a4562a,a4563a,a4564a,a4568a,a4569a,a4572a,a4575a,a4576a,a4577a,a4581a,a4582a,a4585a,a4588a,a4589a,a4590a,a4591a,a4595a,a4596a,a4599a,a4602a,a4603a,a4604a,a4607a,a4610a,a4611a,a4614a,a4617a,a4618a,a4619a,a4620a,a4621a,a4622a,a4623a,a4624a,a4625a,a4629a,a4630a,a4633a,a4636a,a4637a,a4638a,a4642a,a4643a,a4646a,a4649a,a4650a,a4651a,a4652a,a4656a,a4657a,a4660a,a4663a,a4664a,a4665a,a4669a,a4670a,a4673a,a4676a,a4677a,a4678a,a4679a,a4680a,a4684a,a4685a,a4688a,a4691a,a4692a,a4693a,a4697a,a4698a,a4701a,a4704a,a4705a,a4706a,a4707a,a4711a,a4712a,a4715a,a4718a,a4719a,a4720a,a4723a,a4726a,a4727a,a4730a,a4733a,a4734a,a4735a,a4736a,a4737a,a4738a,a4742a,a4743a,a4746a,a4749a,a4750a,a4751a,a4755a,a4756a,a4759a,a4762a,a4763a,a4764a,a4765a,a4769a,a4770a,a4773a,a4776a,a4777a,a4778a,a4781a,a4784a,a4785a,a4788a,a4791a,a4792a,a4793a,a4794a,a4795a,a4799a,a4800a,a4803a,a4806a,a4807a,a4808a,a4812a,a4813a,a4816a,a4819a,a4820a,a4821a,a4822a,a4826a,a4827a,a4830a,a4833a,a4834a,a4835a,a4838a,a4841a,a4842a,a4845a,a4848a,a4849a,a4850a,a4851a,a4852a,a4853a,a4854a,a4858a,a4859a,a4862a,a4865a,a4866a,a4867a,a4871a,a4872a,a4875a,a4878a,a4879a,a4880a,a4881a,a4885a,a4886a,a4889a,a4892a,a4893a,a4894a,a4897a,a4900a,a4901a,a4904a,a4907a,a4908a,a4909a,a4910a,a4911a,a4915a,a4916a,a4919a,a4922a,a4923a,a4924a,a4928a,a4929a,a4932a,a4935a,a4936a,a4937a,a4938a,a4942a,a4943a,a4946a,a4949a,a4950a,a4951a,a4954a,a4957a,a4958a,a4961a,a4964a,a4965a,a4966a,a4967a,a4968a,a4969a,a4973a,a4974a,a4977a,a4980a,a4981a,a4982a,a4986a,a4987a,a4990a,a4993a,a4994a,a4995a,a4996a,a5000a,a5001a,a5004a,a5007a,a5008a,a5009a,a5012a,a5015a,a5016a,a5019a,a5022a,a5023a,a5024a,a5025a,a5026a,a5030a,a5031a,a5034a,a5037a,a5038a,a5039a,a5043a,a5044a,a5047a,a5050a,a5051a,a5052a,a5053a,a5057a,a5058a,a5061a,a5064a,a5065a,a5066a,a5069a,a5072a,a5073a,a5076a,a5079a,a5080a,a5081a,a5082a,a5083a,a5084a,a5085a,a5086a,a5090a,a5091a,a5094a,a5097a,a5098a,a5099a,a5103a,a5104a,a5107a,a5110a,a5111a,a5112a,a5113a,a5117a,a5118a,a5121a,a5124a,a5125a,a5126a,a5129a,a5132a,a5133a,a5136a,a5139a,a5140a,a5141a,a5142a,a5143a,a5147a,a5148a,a5151a,a5154a,a5155a,a5156a,a5160a,a5161a,a5164a,a5167a,a5168a,a5169a,a5170a,a5174a,a5175a,a5178a,a5181a,a5182a,a5183a,a5186a,a5189a,a5190a,a5193a,a5196a,a5197a,a5198a,a5199a,a5200a,a5201a,a5205a,a5206a,a5209a,a5212a,a5213a,a5214a,a5218a,a5219a,a5222a,a5225a,a5226a,a5227a,a5228a,a5232a,a5233a,a5236a,a5239a,a5240a,a5241a,a5244a,a5247a,a5248a,a5251a,a5254a,a5255a,a5256a,a5257a,a5258a,a5262a,a5263a,a5266a,a5269a,a5270a,a5271a,a5275a,a5276a,a5279a,a5282a,a5283a,a5284a,a5285a,a5289a,a5290a,a5293a,a5296a,a5297a,a5298a,a5301a,a5304a,a5305a,a5308a,a5311a,a5312a,a5313a,a5314a,a5315a,a5316a,a5317a,a5321a,a5322a,a5325a,a5328a,a5329a,a5330a,a5334a,a5335a,a5338a,a5341a,a5342a,a5343a,a5344a,a5348a,a5349a,a5352a,a5355a,a5356a,a5357a,a5360a,a5363a,a5364a,a5367a,a5370a,a5371a,a5372a,a5373a,a5374a,a5378a,a5379a,a5382a,a5385a,a5386a,a5387a,a5391a,a5392a,a5395a,a5398a,a5399a,a5400a,a5401a,a5405a,a5406a,a5409a,a5412a,a5413a,a5414a,a5417a,a5420a,a5421a,a5424a,a5427a,a5428a,a5429a,a5430a,a5431a,a5432a,a5436a,a5437a,a5440a,a5443a,a5444a,a5445a,a5449a,a5450a,a5453a,a5456a,a5457a,a5458a,a5459a,a5463a,a5464a,a5467a,a5470a,a5471a,a5472a,a5475a,a5478a,a5479a,a5482a,a5485a,a5486a,a5487a,a5488a,a5489a,a5493a,a5494a,a5497a,a5500a,a5501a,a5502a,a5506a,a5507a,a5510a,a5513a,a5514a,a5515a,a5516a,a5520a,a5521a,a5524a,a5527a,a5528a,a5529a,a5532a,a5535a,a5536a,a5539a,a5542a,a5543a,a5544a,a5545a,a5546a,a5547a,a5548a,a5549a,a5550a,a5551a,a5555a,a5556a,a5559a,a5562a,a5563a,a5564a,a5568a,a5569a,a5572a,a5575a,a5576a,a5577a,a5578a,a5582a,a5583a,a5586a,a5589a,a5590a,a5591a,a5595a,a5596a,a5599a,a5602a,a5603a,a5604a,a5605a,a5606a,a5610a,a5611a,a5614a,a5617a,a5618a,a5619a,a5623a,a5624a,a5627a,a5630a,a5631a,a5632a,a5633a,a5637a,a5638a,a5641a,a5644a,a5645a,a5646a,a5649a,a5652a,a5653a,a5656a,a5659a,a5660a,a5661a,a5662a,a5663a,a5664a,a5668a,a5669a,a5672a,a5675a,a5676a,a5677a,a5681a,a5682a,a5685a,a5688a,a5689a,a5690a,a5691a,a5695a,a5696a,a5699a,a5702a,a5703a,a5704a,a5707a,a5710a,a5711a,a5714a,a5717a,a5718a,a5719a,a5720a,a5721a,a5725a,a5726a,a5729a,a5732a,a5733a,a5734a,a5738a,a5739a,a5742a,a5745a,a5746a,a5747a,a5748a,a5752a,a5753a,a5756a,a5759a,a5760a,a5761a,a5764a,a5767a,a5768a,a5771a,a5774a,a5775a,a5776a,a5777a,a5778a,a5779a,a5780a,a5784a,a5785a,a5788a,a5791a,a5792a,a5793a,a5797a,a5798a,a5801a,a5804a,a5805a,a5806a,a5807a,a5811a,a5812a,a5815a,a5818a,a5819a,a5820a,a5823a,a5826a,a5827a,a5830a,a5833a,a5834a,a5835a,a5836a,a5837a,a5841a,a5842a,a5845a,a5848a,a5849a,a5850a,a5854a,a5855a,a5858a,a5861a,a5862a,a5863a,a5864a,a5868a,a5869a,a5872a,a5875a,a5876a,a5877a,a5880a,a5883a,a5884a,a5887a,a5890a,a5891a,a5892a,a5893a,a5894a,a5895a,a5899a,a5900a,a5903a,a5906a,a5907a,a5908a,a5912a,a5913a,a5916a,a5919a,a5920a,a5921a,a5922a,a5926a,a5927a,a5930a,a5933a,a5934a,a5935a,a5938a,a5941a,a5942a,a5945a,a5948a,a5949a,a5950a,a5951a,a5952a,a5956a,a5957a,a5960a,a5963a,a5964a,a5965a,a5969a,a5970a,a5973a,a5976a,a5977a,a5978a,a5979a,a5983a,a5984a,a5987a,a5990a,a5991a,a5992a,a5995a,a5998a,a5999a,a6002a,a6005a,a6006a,a6007a,a6008a,a6009a,a6010a,a6011a,a6012a,a6016a,a6017a,a6020a,a6023a,a6024a,a6025a,a6029a,a6030a,a6033a,a6036a,a6037a,a6038a,a6039a,a6043a,a6044a,a6047a,a6050a,a6051a,a6052a,a6055a,a6058a,a6059a,a6062a,a6065a,a6066a,a6067a,a6068a,a6069a,a6073a,a6074a,a6077a,a6080a,a6081a,a6082a,a6086a,a6087a,a6090a,a6093a,a6094a,a6095a,a6096a,a6100a,a6101a,a6104a,a6107a,a6108a,a6109a,a6112a,a6115a,a6116a,a6119a,a6122a,a6123a,a6124a,a6125a,a6126a,a6127a,a6131a,a6132a,a6135a,a6138a,a6139a,a6140a,a6144a,a6145a,a6148a,a6151a,a6152a,a6153a,a6154a,a6158a,a6159a,a6162a,a6165a,a6166a,a6167a,a6170a,a6173a,a6174a,a6177a,a6180a,a6181a,a6182a,a6183a,a6184a,a6188a,a6189a,a6192a,a6195a,a6196a,a6197a,a6201a,a6202a,a6205a,a6208a,a6209a,a6210a,a6211a,a6215a,a6216a,a6219a,a6222a,a6223a,a6224a,a6227a,a6230a,a6231a,a6234a,a6237a,a6238a,a6239a,a6240a,a6241a,a6242a,a6243a,a6247a,a6248a,a6251a,a6254a,a6255a,a6256a,a6260a,a6261a,a6264a,a6267a,a6268a,a6269a,a6270a,a6274a,a6275a,a6278a,a6281a,a6282a,a6283a,a6286a,a6289a,a6290a,a6293a,a6296a,a6297a,a6298a,a6299a,a6300a,a6304a,a6305a,a6308a,a6311a,a6312a,a6313a,a6317a,a6318a,a6321a,a6324a,a6325a,a6326a,a6327a,a6331a,a6332a,a6335a,a6338a,a6339a,a6340a,a6343a,a6346a,a6347a,a6350a,a6353a,a6354a,a6355a,a6356a,a6357a,a6358a,a6362a,a6363a,a6366a,a6369a,a6370a,a6371a,a6375a,a6376a,a6379a,a6382a,a6383a,a6384a,a6385a,a6389a,a6390a,a6393a,a6396a,a6397a,a6398a,a6401a,a6404a,a6405a,a6408a,a6411a,a6412a,a6413a,a6414a,a6415a,a6419a,a6420a,a6423a,a6426a,a6427a,a6428a,a6432a,a6433a,a6436a,a6439a,a6440a,a6441a,a6442a,a6446a,a6447a,a6450a,a6453a,a6454a,a6455a,a6458a,a6461a,a6462a,a6465a,a6468a,a6469a,a6470a,a6471a,a6472a,a6473a,a6474a,a6475a,a6476a,a6480a,a6481a,a6484a,a6487a,a6488a,a6489a,a6493a,a6494a,a6497a,a6500a,a6501a,a6502a,a6503a,a6507a,a6508a,a6511a,a6514a,a6515a,a6516a,a6520a,a6521a,a6524a,a6527a,a6528a,a6529a,a6530a,a6531a,a6535a,a6536a,a6539a,a6542a,a6543a,a6544a,a6548a,a6549a,a6552a,a6555a,a6556a,a6557a,a6558a,a6562a,a6563a,a6566a,a6569a,a6570a,a6571a,a6574a,a6577a,a6578a,a6581a,a6584a,a6585a,a6586a,a6587a,a6588a,a6589a,a6593a,a6594a,a6597a,a6600a,a6601a,a6602a,a6606a,a6607a,a6610a,a6613a,a6614a,a6615a,a6616a,a6620a,a6621a,a6624a,a6627a,a6628a,a6629a,a6632a,a6635a,a6636a,a6639a,a6642a,a6643a,a6644a,a6645a,a6646a,a6650a,a6651a,a6654a,a6657a,a6658a,a6659a,a6663a,a6664a,a6667a,a6670a,a6671a,a6672a,a6673a,a6677a,a6678a,a6681a,a6684a,a6685a,a6686a,a6689a,a6692a,a6693a,a6696a,a6699a,a6700a,a6701a,a6702a,a6703a,a6704a,a6705a,a6709a,a6710a,a6713a,a6716a,a6717a,a6718a,a6722a,a6723a,a6726a,a6729a,a6730a,a6731a,a6732a,a6736a,a6737a,a6740a,a6743a,a6744a,a6745a,a6748a,a6751a,a6752a,a6755a,a6758a,a6759a,a6760a,a6761a,a6762a,a6766a,a6767a,a6770a,a6773a,a6774a,a6775a,a6779a,a6780a,a6783a,a6786a,a6787a,a6788a,a6789a,a6793a,a6794a,a6797a,a6800a,a6801a,a6802a,a6805a,a6808a,a6809a,a6812a,a6815a,a6816a,a6817a,a6818a,a6819a,a6820a,a6824a,a6825a,a6828a,a6831a,a6832a,a6833a,a6837a,a6838a,a6841a,a6844a,a6845a,a6846a,a6847a,a6851a,a6852a,a6855a,a6858a,a6859a,a6860a,a6863a,a6866a,a6867a,a6870a,a6873a,a6874a,a6875a,a6876a,a6877a,a6881a,a6882a,a6885a,a6888a,a6889a,a6890a,a6894a,a6895a,a6898a,a6901a,a6902a,a6903a,a6904a,a6908a,a6909a,a6912a,a6915a,a6916a,a6917a,a6920a,a6923a,a6924a,a6927a,a6930a,a6931a,a6932a,a6933a,a6934a,a6935a,a6936a,a6937a,a6941a,a6942a,a6945a,a6948a,a6949a,a6950a,a6954a,a6955a,a6958a,a6961a,a6962a,a6963a,a6964a,a6968a,a6969a,a6972a,a6975a,a6976a,a6977a,a6980a,a6983a,a6984a,a6987a,a6990a,a6991a,a6992a,a6993a,a6994a,a6998a,a6999a,a7002a,a7005a,a7006a,a7007a,a7011a,a7012a,a7015a,a7018a,a7019a,a7020a,a7021a,a7025a,a7026a,a7029a,a7032a,a7033a,a7034a,a7037a,a7040a,a7041a,a7044a,a7047a,a7048a,a7049a,a7050a,a7051a,a7052a,a7056a,a7057a,a7060a,a7063a,a7064a,a7065a,a7069a,a7070a,a7073a,a7076a,a7077a,a7078a,a7079a,a7083a,a7084a,a7087a,a7090a,a7091a,a7092a,a7095a,a7098a,a7099a,a7102a,a7105a,a7106a,a7107a,a7108a,a7109a,a7113a,a7114a,a7117a,a7120a,a7121a,a7122a,a7126a,a7127a,a7130a,a7133a,a7134a,a7135a,a7136a,a7140a,a7141a,a7144a,a7147a,a7148a,a7149a,a7152a,a7155a,a7156a,a7159a,a7162a,a7163a,a7164a,a7165a,a7166a,a7167a,a7168a,a7172a,a7173a,a7176a,a7179a,a7180a,a7181a,a7185a,a7186a,a7189a,a7192a,a7193a,a7194a,a7195a,a7199a,a7200a,a7203a,a7206a,a7207a,a7208a,a7211a,a7214a,a7215a,a7218a,a7221a,a7222a,a7223a,a7224a,a7225a,a7229a,a7230a,a7233a,a7236a,a7237a,a7238a,a7242a,a7243a,a7246a,a7249a,a7250a,a7251a,a7252a,a7256a,a7257a,a7260a,a7263a,a7264a,a7265a,a7268a,a7271a,a7272a,a7275a,a7278a,a7279a,a7280a,a7281a,a7282a,a7283a,a7287a,a7288a,a7291a,a7294a,a7295a,a7296a,a7300a,a7301a,a7304a,a7307a,a7308a,a7309a,a7310a,a7314a,a7315a,a7318a,a7321a,a7322a,a7323a,a7326a,a7329a,a7330a,a7333a,a7336a,a7337a,a7338a,a7339a,a7340a,a7344a,a7345a,a7348a,a7351a,a7352a,a7353a,a7357a,a7358a,a7361a,a7364a,a7365a,a7366a,a7367a,a7371a,a7372a,a7375a,a7378a,a7379a,a7380a,a7383a,a7386a,a7387a,a7390a,a7393a,a7394a,a7395a,a7396a,a7397a,a7398a,a7399a,a7400a,a7401a,a7402a,a7403a,a7407a,a7408a,a7411a,a7414a,a7415a,a7416a,a7420a,a7421a,a7424a,a7427a,a7428a,a7429a,a7430a,a7434a,a7435a,a7438a,a7441a,a7442a,a7443a,a7447a,a7448a,a7451a,a7454a,a7455a,a7456a,a7457a,a7458a,a7462a,a7463a,a7466a,a7469a,a7470a,a7471a,a7475a,a7476a,a7479a,a7482a,a7483a,a7484a,a7485a,a7489a,a7490a,a7493a,a7496a,a7497a,a7498a,a7501a,a7504a,a7505a,a7508a,a7511a,a7512a,a7513a,a7514a,a7515a,a7516a,a7520a,a7521a,a7524a,a7527a,a7528a,a7529a,a7533a,a7534a,a7537a,a7540a,a7541a,a7542a,a7543a,a7547a,a7548a,a7551a,a7554a,a7555a,a7556a,a7559a,a7562a,a7563a,a7566a,a7569a,a7570a,a7571a,a7572a,a7573a,a7577a,a7578a,a7581a,a7584a,a7585a,a7586a,a7590a,a7591a,a7594a,a7597a,a7598a,a7599a,a7600a,a7604a,a7605a,a7608a,a7611a,a7612a,a7613a,a7616a,a7619a,a7620a,a7623a,a7626a,a7627a,a7628a,a7629a,a7630a,a7631a,a7632a,a7636a,a7637a,a7640a,a7643a,a7644a,a7645a,a7649a,a7650a,a7653a,a7656a,a7657a,a7658a,a7659a,a7663a,a7664a,a7667a,a7670a,a7671a,a7672a,a7675a,a7678a,a7679a,a7682a,a7685a,a7686a,a7687a,a7688a,a7689a,a7693a,a7694a,a7697a,a7700a,a7701a,a7702a,a7706a,a7707a,a7710a,a7713a,a7714a,a7715a,a7716a,a7720a,a7721a,a7724a,a7727a,a7728a,a7729a,a7732a,a7735a,a7736a,a7739a,a7742a,a7743a,a7744a,a7745a,a7746a,a7747a,a7751a,a7752a,a7755a,a7758a,a7759a,a7760a,a7764a,a7765a,a7768a,a7771a,a7772a,a7773a,a7774a,a7778a,a7779a,a7782a,a7785a,a7786a,a7787a,a7790a,a7793a,a7794a,a7797a,a7800a,a7801a,a7802a,a7803a,a7804a,a7808a,a7809a,a7812a,a7815a,a7816a,a7817a,a7821a,a7822a,a7825a,a7828a,a7829a,a7830a,a7831a,a7835a,a7836a,a7839a,a7842a,a7843a,a7844a,a7847a,a7850a,a7851a,a7854a,a7857a,a7858a,a7859a,a7860a,a7861a,a7862a,a7863a,a7864a,a7868a,a7869a,a7872a,a7875a,a7876a,a7877a,a7881a,a7882a,a7885a,a7888a,a7889a,a7890a,a7891a,a7895a,a7896a,a7899a,a7902a,a7903a,a7904a,a7908a,a7909a,a7912a,a7915a,a7916a,a7917a,a7918a,a7919a,a7923a,a7924a,a7927a,a7930a,a7931a,a7932a,a7936a,a7937a,a7940a,a7943a,a7944a,a7945a,a7946a,a7950a,a7951a,a7954a,a7957a,a7958a,a7959a,a7962a,a7965a,a7966a,a7969a,a7972a,a7973a,a7974a,a7975a,a7976a,a7977a,a7981a,a7982a,a7985a,a7988a,a7989a,a7990a,a7994a,a7995a,a7998a,a8001a,a8002a,a8003a,a8004a,a8008a,a8009a,a8012a,a8015a,a8016a,a8017a,a8020a,a8023a,a8024a,a8027a,a8030a,a8031a,a8032a,a8033a,a8034a,a8038a,a8039a,a8042a,a8045a,a8046a,a8047a,a8051a,a8052a,a8055a,a8058a,a8059a,a8060a,a8061a,a8065a,a8066a,a8069a,a8072a,a8073a,a8074a,a8077a,a8080a,a8081a,a8084a,a8087a,a8088a,a8089a,a8090a,a8091a,a8092a,a8093a,a8097a,a8098a,a8101a,a8104a,a8105a,a8106a,a8110a,a8111a,a8114a,a8117a,a8118a,a8119a,a8120a,a8124a,a8125a,a8128a,a8131a,a8132a,a8133a,a8136a,a8139a,a8140a,a8143a,a8146a,a8147a,a8148a,a8149a,a8150a,a8154a,a8155a,a8158a,a8161a,a8162a,a8163a,a8167a,a8168a,a8171a,a8174a,a8175a,a8176a,a8177a,a8181a,a8182a,a8185a,a8188a,a8189a,a8190a,a8193a,a8196a,a8197a,a8200a,a8203a,a8204a,a8205a,a8206a,a8207a,a8208a,a8212a,a8213a,a8216a,a8219a,a8220a,a8221a,a8225a,a8226a,a8229a,a8232a,a8233a,a8234a,a8235a,a8239a,a8240a,a8243a,a8246a,a8247a,a8248a,a8251a,a8254a,a8255a,a8258a,a8261a,a8262a,a8263a,a8264a,a8265a,a8269a,a8270a,a8273a,a8276a,a8277a,a8278a,a8282a,a8283a,a8286a,a8289a,a8290a,a8291a,a8292a,a8296a,a8297a,a8300a,a8303a,a8304a,a8305a,a8308a,a8311a,a8312a,a8315a,a8318a,a8319a,a8320a,a8321a,a8322a,a8323a,a8324a,a8325a,a8326a,a8330a,a8331a,a8334a,a8337a,a8338a,a8339a,a8343a,a8344a,a8347a,a8350a,a8351a,a8352a,a8353a,a8357a,a8358a,a8361a,a8364a,a8365a,a8366a,a8370a,a8371a,a8374a,a8377a,a8378a,a8379a,a8380a,a8381a,a8385a,a8386a,a8389a,a8392a,a8393a,a8394a,a8398a,a8399a,a8402a,a8405a,a8406a,a8407a,a8408a,a8412a,a8413a,a8416a,a8419a,a8420a,a8421a,a8424a,a8427a,a8428a,a8431a,a8434a,a8435a,a8436a,a8437a,a8438a,a8439a,a8443a,a8444a,a8447a,a8450a,a8451a,a8452a,a8456a,a8457a,a8460a,a8463a,a8464a,a8465a,a8466a,a8470a,a8471a,a8474a,a8477a,a8478a,a8479a,a8482a,a8485a,a8486a,a8489a,a8492a,a8493a,a8494a,a8495a,a8496a,a8500a,a8501a,a8504a,a8507a,a8508a,a8509a,a8513a,a8514a,a8517a,a8520a,a8521a,a8522a,a8523a,a8527a,a8528a,a8531a,a8534a,a8535a,a8536a,a8539a,a8542a,a8543a,a8546a,a8549a,a8550a,a8551a,a8552a,a8553a,a8554a,a8555a,a8559a,a8560a,a8563a,a8566a,a8567a,a8568a,a8572a,a8573a,a8576a,a8579a,a8580a,a8581a,a8582a,a8586a,a8587a,a8590a,a8593a,a8594a,a8595a,a8598a,a8601a,a8602a,a8605a,a8608a,a8609a,a8610a,a8611a,a8612a,a8616a,a8617a,a8620a,a8623a,a8624a,a8625a,a8629a,a8630a,a8633a,a8636a,a8637a,a8638a,a8639a,a8643a,a8644a,a8647a,a8650a,a8651a,a8652a,a8655a,a8658a,a8659a,a8662a,a8665a,a8666a,a8667a,a8668a,a8669a,a8670a,a8674a,a8675a,a8678a,a8681a,a8682a,a8683a,a8687a,a8688a,a8691a,a8694a,a8695a,a8696a,a8697a,a8701a,a8702a,a8705a,a8708a,a8709a,a8710a,a8713a,a8716a,a8717a,a8720a,a8723a,a8724a,a8725a,a8726a,a8727a,a8731a,a8732a,a8735a,a8738a,a8739a,a8740a,a8744a,a8745a,a8748a,a8751a,a8752a,a8753a,a8754a,a8758a,a8759a,a8762a,a8765a,a8766a,a8767a,a8770a,a8773a,a8774a,a8777a,a8780a,a8781a,a8782a,a8783a,a8784a,a8785a,a8786a,a8787a,a8791a,a8792a,a8795a,a8798a,a8799a,a8800a,a8804a,a8805a,a8808a,a8811a,a8812a,a8813a,a8814a,a8818a,a8819a,a8822a,a8825a,a8826a,a8827a,a8830a,a8833a,a8834a,a8837a,a8840a,a8841a,a8842a,a8843a,a8844a,a8848a,a8849a,a8852a,a8855a,a8856a,a8857a,a8861a,a8862a,a8865a,a8868a,a8869a,a8870a,a8871a,a8875a,a8876a,a8879a,a8882a,a8883a,a8884a,a8887a,a8890a,a8891a,a8894a,a8897a,a8898a,a8899a,a8900a,a8901a,a8902a,a8906a,a8907a,a8910a,a8913a,a8914a,a8915a,a8919a,a8920a,a8923a,a8926a,a8927a,a8928a,a8929a,a8933a,a8934a,a8937a,a8940a,a8941a,a8942a,a8945a,a8948a,a8949a,a8952a,a8955a,a8956a,a8957a,a8958a,a8959a,a8963a,a8964a,a8967a,a8970a,a8971a,a8972a,a8976a,a8977a,a8980a,a8983a,a8984a,a8985a,a8986a,a8990a,a8991a,a8994a,a8997a,a8998a,a8999a,a9002a,a9005a,a9006a,a9009a,a9012a,a9013a,a9014a,a9015a,a9016a,a9017a,a9018a,a9022a,a9023a,a9026a,a9029a,a9030a,a9031a,a9035a,a9036a,a9039a,a9042a,a9043a,a9044a,a9045a,a9049a,a9050a,a9053a,a9056a,a9057a,a9058a,a9061a,a9064a,a9065a,a9068a,a9071a,a9072a,a9073a,a9074a,a9075a,a9079a,a9080a,a9083a,a9086a,a9087a,a9088a,a9092a,a9093a,a9096a,a9099a,a9100a,a9101a,a9102a,a9106a,a9107a,a9110a,a9113a,a9114a,a9115a,a9118a,a9121a,a9122a,a9125a,a9128a,a9129a,a9130a,a9131a,a9132a,a9133a,a9137a,a9138a,a9141a,a9144a,a9145a,a9146a,a9150a,a9151a,a9154a,a9157a,a9158a,a9159a,a9160a,a9164a,a9165a,a9168a,a9171a,a9172a,a9173a,a9176a,a9179a,a9180a,a9183a,a9186a,a9187a,a9188a,a9189a,a9190a,a9194a,a9195a,a9198a,a9201a,a9202a,a9203a,a9207a,a9208a,a9211a,a9214a,a9215a,a9216a,a9217a,a9221a,a9222a,a9225a,a9228a,a9229a,a9230a,a9233a,a9236a,a9237a,a9240a,a9243a,a9244a,a9245a,a9246a,a9247a,a9248a,a9249a,a9250a,a9251a,a9252a,a9256a,a9257a,a9260a,a9263a,a9264a,a9265a,a9269a,a9270a,a9273a,a9276a,a9277a,a9278a,a9279a,a9283a,a9284a,a9287a,a9290a,a9291a,a9292a,a9296a,a9297a,a9300a,a9303a,a9304a,a9305a,a9306a,a9307a,a9311a,a9312a,a9315a,a9318a,a9319a,a9320a,a9324a,a9325a,a9328a,a9331a,a9332a,a9333a,a9334a,a9338a,a9339a,a9342a,a9345a,a9346a,a9347a,a9350a,a9353a,a9354a,a9357a,a9360a,a9361a,a9362a,a9363a,a9364a,a9365a,a9369a,a9370a,a9373a,a9376a,a9377a,a9378a,a9382a,a9383a,a9386a,a9389a,a9390a,a9391a,a9392a,a9396a,a9397a,a9400a,a9403a,a9404a,a9405a,a9408a,a9411a,a9412a,a9415a,a9418a,a9419a,a9420a,a9421a,a9422a,a9426a,a9427a,a9430a,a9433a,a9434a,a9435a,a9439a,a9440a,a9443a,a9446a,a9447a,a9448a,a9449a,a9453a,a9454a,a9457a,a9460a,a9461a,a9462a,a9465a,a9468a,a9469a,a9472a,a9475a,a9476a,a9477a,a9478a,a9479a,a9480a,a9481a,a9485a,a9486a,a9489a,a9492a,a9493a,a9494a,a9498a,a9499a,a9502a,a9505a,a9506a,a9507a,a9508a,a9512a,a9513a,a9516a,a9519a,a9520a,a9521a,a9524a,a9527a,a9528a,a9531a,a9534a,a9535a,a9536a,a9537a,a9538a,a9542a,a9543a,a9546a,a9549a,a9550a,a9551a,a9555a,a9556a,a9559a,a9562a,a9563a,a9564a,a9565a,a9569a,a9570a,a9573a,a9576a,a9577a,a9578a,a9581a,a9584a,a9585a,a9588a,a9591a,a9592a,a9593a,a9594a,a9595a,a9596a,a9600a,a9601a,a9604a,a9607a,a9608a,a9609a,a9613a,a9614a,a9617a,a9620a,a9621a,a9622a,a9623a,a9627a,a9628a,a9631a,a9634a,a9635a,a9636a,a9639a,a9642a,a9643a,a9646a,a9649a,a9650a,a9651a,a9652a,a9653a,a9657a,a9658a,a9661a,a9664a,a9665a,a9666a,a9670a,a9671a,a9674a,a9677a,a9678a,a9679a,a9680a,a9684a,a9685a,a9688a,a9691a,a9692a,a9693a,a9696a,a9699a,a9700a,a9703a,a9706a,a9707a,a9708a,a9709a,a9710a,a9711a,a9712a,a9713a,a9717a,a9718a,a9721a,a9724a,a9725a,a9726a,a9730a,a9731a,a9734a,a9737a,a9738a,a9739a,a9740a,a9744a,a9745a,a9748a,a9751a,a9752a,a9753a,a9756a,a9759a,a9760a,a9763a,a9766a,a9767a,a9768a,a9769a,a9770a,a9774a,a9775a,a9778a,a9781a,a9782a,a9783a,a9787a,a9788a,a9791a,a9794a,a9795a,a9796a,a9797a,a9801a,a9802a,a9805a,a9808a,a9809a,a9810a,a9813a,a9816a,a9817a,a9820a,a9823a,a9824a,a9825a,a9826a,a9827a,a9828a,a9832a,a9833a,a9836a,a9839a,a9840a,a9841a,a9845a,a9846a,a9849a,a9852a,a9853a,a9854a,a9855a,a9859a,a9860a,a9863a,a9866a,a9867a,a9868a,a9871a,a9874a,a9875a,a9878a,a9881a,a9882a,a9883a,a9884a,a9885a,a9889a,a9890a,a9893a,a9896a,a9897a,a9898a,a9902a,a9903a,a9906a,a9909a,a9910a,a9911a,a9912a,a9916a,a9917a,a9920a,a9923a,a9924a,a9925a,a9928a,a9931a,a9932a,a9935a,a9938a,a9939a,a9940a,a9941a,a9942a,a9943a,a9944a,a9948a,a9949a,a9952a,a9955a,a9956a,a9957a,a9961a,a9962a,a9965a,a9968a,a9969a,a9970a,a9971a,a9975a,a9976a,a9979a,a9982a,a9983a,a9984a,a9987a,a9990a,a9991a,a9994a,a9997a,a9998a,a9999a,a10000a,a10001a,a10005a,a10006a,a10009a,a10012a,a10013a,a10014a,a10018a,a10019a,a10022a,a10025a,a10026a,a10027a,a10028a,a10032a,a10033a,a10036a,a10039a,a10040a,a10041a,a10044a,a10047a,a10048a,a10051a,a10054a,a10055a,a10056a,a10057a,a10058a,a10059a,a10063a,a10064a,a10067a,a10070a,a10071a,a10072a,a10076a,a10077a,a10080a,a10083a,a10084a,a10085a,a10086a,a10090a,a10091a,a10094a,a10097a,a10098a,a10099a,a10102a,a10105a,a10106a,a10109a,a10112a,a10113a,a10114a,a10115a,a10116a,a10120a,a10121a,a10124a,a10127a,a10128a,a10129a,a10133a,a10134a,a10137a,a10140a,a10141a,a10142a,a10143a,a10147a,a10148a,a10151a,a10154a,a10155a,a10156a,a10159a,a10162a,a10163a,a10166a,a10169a,a10170a,a10171a,a10172a,a10173a,a10174a,a10175a,a10176a,a10177a,a10181a,a10182a,a10185a,a10188a,a10189a,a10190a,a10194a,a10195a,a10198a,a10201a,a10202a,a10203a,a10204a,a10208a,a10209a,a10212a,a10215a,a10216a,a10217a,a10221a,a10222a,a10225a,a10228a,a10229a,a10230a,a10231a,a10232a,a10236a,a10237a,a10240a,a10243a,a10244a,a10245a,a10249a,a10250a,a10253a,a10256a,a10257a,a10258a,a10259a,a10263a,a10264a,a10267a,a10270a,a10271a,a10272a,a10275a,a10278a,a10279a,a10282a,a10285a,a10286a,a10287a,a10288a,a10289a,a10290a,a10294a,a10295a,a10298a,a10301a,a10302a,a10303a,a10307a,a10308a,a10311a,a10314a,a10315a,a10316a,a10317a,a10321a,a10322a,a10325a,a10328a,a10329a,a10330a,a10333a,a10336a,a10337a,a10340a,a10343a,a10344a,a10345a,a10346a,a10347a,a10351a,a10352a,a10355a,a10358a,a10359a,a10360a,a10364a,a10365a,a10368a,a10371a,a10372a,a10373a,a10374a,a10378a,a10379a,a10382a,a10385a,a10386a,a10387a,a10390a,a10393a,a10394a,a10397a,a10400a,a10401a,a10402a,a10403a,a10404a,a10405a,a10406a,a10410a,a10411a,a10414a,a10417a,a10418a,a10419a,a10423a,a10424a,a10427a,a10430a,a10431a,a10432a,a10433a,a10437a,a10438a,a10441a,a10444a,a10445a,a10446a,a10449a,a10452a,a10453a,a10456a,a10459a,a10460a,a10461a,a10462a,a10463a,a10467a,a10468a,a10471a,a10474a,a10475a,a10476a,a10480a,a10481a,a10484a,a10487a,a10488a,a10489a,a10490a,a10494a,a10495a,a10498a,a10501a,a10502a,a10503a,a10506a,a10509a,a10510a,a10513a,a10516a,a10517a,a10518a,a10519a,a10520a,a10521a,a10525a,a10526a,a10529a,a10532a,a10533a,a10534a,a10538a,a10539a,a10542a,a10545a,a10546a,a10547a,a10548a,a10552a,a10553a,a10556a,a10559a,a10560a,a10561a,a10564a,a10567a,a10568a,a10571a,a10574a,a10575a,a10576a,a10577a,a10578a,a10582a,a10583a,a10586a,a10589a,a10590a,a10591a,a10595a,a10596a,a10599a,a10602a,a10603a,a10604a,a10605a,a10609a,a10610a,a10613a,a10616a,a10617a,a10618a,a10621a,a10624a,a10625a,a10628a,a10631a,a10632a,a10633a,a10634a,a10635a,a10636a,a10637a,a10638a,a10642a,a10643a,a10646a,a10649a,a10650a,a10651a,a10655a,a10656a,a10659a,a10662a,a10663a,a10664a,a10665a,a10669a,a10670a,a10673a,a10676a,a10677a,a10678a,a10681a,a10684a,a10685a,a10688a,a10691a,a10692a,a10693a,a10694a,a10695a,a10699a,a10700a,a10703a,a10706a,a10707a,a10708a,a10712a,a10713a,a10716a,a10719a,a10720a,a10721a,a10722a,a10726a,a10727a,a10730a,a10733a,a10734a,a10735a,a10738a,a10741a,a10742a,a10745a,a10748a,a10749a,a10750a,a10751a,a10752a,a10753a,a10757a,a10758a,a10761a,a10764a,a10765a,a10766a,a10770a,a10771a,a10774a,a10777a,a10778a,a10779a,a10780a,a10784a,a10785a,a10788a,a10791a,a10792a,a10793a,a10796a,a10799a,a10800a,a10803a,a10806a,a10807a,a10808a,a10809a,a10810a,a10814a,a10815a,a10818a,a10821a,a10822a,a10823a,a10827a,a10828a,a10831a,a10834a,a10835a,a10836a,a10837a,a10841a,a10842a,a10845a,a10848a,a10849a,a10850a,a10853a,a10856a,a10857a,a10860a,a10863a,a10864a,a10865a,a10866a,a10867a,a10868a,a10869a,a10873a,a10874a,a10877a,a10880a,a10881a,a10882a,a10886a,a10887a,a10890a,a10893a,a10894a,a10895a,a10896a,a10900a,a10901a,a10904a,a10907a,a10908a,a10909a,a10912a,a10915a,a10916a,a10919a,a10922a,a10923a,a10924a,a10925a,a10926a,a10930a,a10931a,a10934a,a10937a,a10938a,a10939a,a10943a,a10944a,a10947a,a10950a,a10951a,a10952a,a10953a,a10957a,a10958a,a10961a,a10964a,a10965a,a10966a,a10969a,a10972a,a10973a,a10976a,a10979a,a10980a,a10981a,a10982a,a10983a,a10984a,a10988a,a10989a,a10992a,a10995a,a10996a,a10997a,a11001a,a11002a,a11005a,a11008a,a11009a,a11010a,a11011a,a11015a,a11016a,a11019a,a11022a,a11023a,a11024a,a11027a,a11030a,a11031a,a11034a,a11037a,a11038a,a11039a,a11040a,a11041a,a11045a,a11046a,a11049a,a11052a,a11053a,a11054a,a11058a,a11059a,a11062a,a11065a,a11066a,a11067a,a11068a,a11072a,a11073a,a11076a,a11079a,a11080a,a11081a,a11084a,a11087a,a11088a,a11091a,a11094a,a11095a,a11096a,a11097a,a11098a,a11099a,a11100a,a11101a,a11102a,a11103a,a11104a,a11107a,a11110a,a11111a,a11114a,a11117a,a11118a,a11121a,a11124a,a11125a,a11128a,a11131a,a11132a,a11135a,a11138a,a11139a,a11142a,a11145a,a11146a,a11149a,a11152a,a11153a,a11156a,a11159a,a11160a,a11163a,a11166a,a11167a,a11170a,a11173a,a11174a,a11177a,a11180a,a11181a,a11184a,a11187a,a11188a,a11191a,a11194a,a11195a,a11198a,a11201a,a11202a,a11205a,a11208a,a11209a,a11212a,a11215a,a11216a,a11219a,a11222a,a11223a,a11226a,a11229a,a11230a,a11233a,a11236a,a11237a,a11240a,a11243a,a11244a,a11247a,a11250a,a11251a,a11254a,a11257a,a11258a,a11261a,a11264a,a11265a,a11268a,a11271a,a11272a,a11275a,a11278a,a11279a,a11282a,a11285a,a11286a,a11289a,a11292a,a11293a,a11296a,a11299a,a11300a,a11303a,a11306a,a11307a,a11310a,a11313a,a11314a,a11317a,a11320a,a11321a,a11324a,a11327a,a11328a,a11331a,a11334a,a11335a,a11338a,a11341a,a11342a,a11345a,a11348a,a11349a,a11352a,a11355a,a11356a,a11359a,a11362a,a11363a,a11366a,a11369a,a11370a,a11373a,a11376a,a11377a,a11380a,a11383a,a11384a,a11387a,a11390a,a11391a,a11394a,a11397a,a11398a,a11401a,a11404a,a11405a,a11408a,a11411a,a11412a,a11415a,a11418a,a11419a,a11422a,a11425a,a11426a,a11429a,a11432a,a11433a,a11436a,a11439a,a11440a,a11443a,a11446a,a11447a,a11450a,a11453a,a11454a,a11457a,a11460a,a11461a,a11464a,a11467a,a11468a,a11471a,a11474a,a11475a,a11478a,a11481a,a11482a,a11485a,a11488a,a11489a,a11492a,a11495a,a11496a,a11499a,a11502a,a11503a,a11506a,a11509a,a11510a,a11513a,a11516a,a11517a,a11520a,a11523a,a11524a,a11527a,a11530a,a11531a,a11534a,a11537a,a11538a,a11541a,a11544a,a11545a,a11548a,a11551a,a11552a,a11555a,a11558a,a11559a,a11562a,a11566a,a11567a,a11568a,a11571a,a11574a,a11575a,a11578a,a11582a,a11583a,a11584a,a11587a,a11590a,a11591a,a11594a,a11598a,a11599a,a11600a,a11603a,a11606a,a11607a,a11610a,a11614a,a11615a,a11616a,a11619a,a11622a,a11623a,a11626a,a11630a,a11631a,a11632a,a11635a,a11638a,a11639a,a11642a,a11646a,a11647a,a11648a,a11651a,a11654a,a11655a,a11658a,a11662a,a11663a,a11664a,a11667a,a11670a,a11671a,a11674a,a11678a,a11679a,a11680a,a11683a,a11686a,a11687a,a11690a,a11694a,a11695a,a11696a,a11699a,a11702a,a11703a,a11706a,a11710a,a11711a,a11712a,a11715a,a11718a,a11719a,a11722a,a11726a,a11727a,a11728a,a11731a,a11734a,a11735a,a11738a,a11742a,a11743a,a11744a,a11747a,a11750a,a11751a,a11754a,a11758a,a11759a,a11760a,a11763a,a11766a,a11767a,a11770a,a11774a,a11775a,a11776a,a11779a,a11782a,a11783a,a11786a,a11790a,a11791a,a11792a,a11795a,a11798a,a11799a,a11802a,a11806a,a11807a,a11808a,a11811a,a11814a,a11815a,a11818a,a11822a,a11823a,a11824a,a11827a,a11830a,a11831a,a11834a,a11838a,a11839a,a11840a,a11843a,a11846a,a11847a,a11850a,a11854a,a11855a,a11856a,a11859a,a11862a,a11863a,a11866a,a11870a,a11871a,a11872a,a11875a,a11878a,a11879a,a11882a,a11886a,a11887a,a11888a,a11891a,a11894a,a11895a,a11898a,a11902a,a11903a,a11904a,a11907a,a11910a,a11911a,a11914a,a11918a,a11919a,a11920a,a11923a,a11926a,a11927a,a11930a,a11934a,a11935a,a11936a,a11939a,a11942a,a11943a,a11946a,a11950a,a11951a,a11952a,a11955a,a11958a,a11959a,a11962a,a11966a,a11967a,a11968a,a11971a,a11974a,a11975a,a11978a,a11982a,a11983a,a11984a,a11987a,a11990a,a11991a,a11994a,a11998a,a11999a,a12000a,a12003a,a12006a,a12007a,a12010a,a12014a,a12015a,a12016a,a12019a,a12022a,a12023a,a12026a,a12030a,a12031a,a12032a,a12035a,a12038a,a12039a,a12042a,a12046a,a12047a,a12048a,a12051a,a12054a,a12055a,a12058a,a12062a,a12063a,a12064a,a12067a,a12071a,a12072a,a12073a,a12076a,a12080a,a12081a,a12082a,a12085a,a12089a,a12090a,a12091a,a12094a,a12098a,a12099a,a12100a,a12103a,a12107a,a12108a,a12109a,a12112a,a12116a,a12117a,a12118a,a12121a,a12125a,a12126a,a12127a,a12130a,a12134a,a12135a,a12136a,a12139a,a12143a,a12144a,a12145a,a12148a,a12152a,a12153a,a12154a,a12157a,a12161a,a12162a,a12163a,a12166a,a12170a,a12171a,a12172a,a12175a,a12179a,a12180a,a12181a,a12184a,a12188a,a12189a,a12190a,a12193a,a12197a,a12198a,a12199a,a12202a,a12206a,a12207a,a12208a,a12211a,a12215a,a12216a,a12217a,a12220a,a12224a,a12225a,a12226a,a12229a,a12233a,a12234a,a12235a,a12238a,a12242a,a12243a,a12244a,a12247a,a12251a,a12252a,a12253a,a12256a,a12260a,a12261a,a12262a,a12265a,a12269a,a12270a,a12271a,a12274a,a12278a,a12279a,a12280a,a12283a,a12287a,a12288a,a12289a,a12292a,a12296a,a12297a,a12298a,a12301a,a12305a,a12306a,a12307a,a12310a,a12314a,a12315a,a12316a,a12319a,a12323a,a12324a,a12325a,a12328a,a12332a,a12333a,a12334a,a12337a,a12341a,a12342a,a12343a,a12346a,a12350a,a12351a,a12352a,a12355a,a12359a,a12360a,a12361a,a12364a,a12368a,a12369a,a12370a,a12373a,a12377a,a12378a,a12379a,a12382a,a12386a,a12387a,a12388a,a12391a,a12395a,a12396a,a12397a,a12400a,a12404a,a12405a,a12406a,a12409a,a12413a,a12414a,a12415a,a12418a,a12422a,a12423a,a12424a,a12427a,a12431a,a12432a,a12433a,a12436a,a12440a,a12441a,a12442a,a12445a,a12449a,a12450a,a12451a,a12454a,a12458a,a12459a,a12460a,a12463a,a12467a,a12468a,a12469a,a12472a,a12476a,a12477a,a12478a,a12481a,a12485a,a12486a,a12487a,a12490a,a12494a,a12495a,a12496a,a12499a,a12503a,a12504a,a12505a,a12508a,a12512a,a12513a,a12514a,a12517a,a12521a,a12522a,a12523a,a12526a,a12530a,a12531a,a12532a,a12535a,a12539a,a12540a,a12541a,a12544a,a12548a,a12549a,a12550a,a12553a,a12557a,a12558a,a12559a,a12562a,a12566a,a12567a,a12568a,a12571a,a12575a,a12576a,a12577a,a12580a,a12584a,a12585a,a12586a,a12589a,a12593a,a12594a,a12595a,a12598a,a12602a,a12603a,a12604a,a12607a,a12611a,a12612a,a12613a,a12616a,a12620a,a12621a,a12622a,a12625a,a12629a,a12630a,a12631a,a12634a,a12638a,a12639a,a12640a,a12643a,a12647a,a12648a,a12649a,a12652a,a12656a,a12657a,a12658a,a12661a,a12665a,a12666a,a12667a,a12670a,a12674a,a12675a,a12676a,a12679a,a12683a,a12684a,a12685a,a12688a,a12692a,a12693a,a12694a,a12697a,a12701a,a12702a,a12703a,a12706a,a12710a,a12711a,a12712a,a12715a,a12719a,a12720a,a12721a,a12724a,a12728a,a12729a,a12730a,a12733a,a12737a,a12738a,a12739a,a12742a,a12746a,a12747a,a12748a,a12751a,a12755a,a12756a,a12757a,a12760a,a12764a,a12765a,a12766a,a12769a,a12773a,a12774a,a12775a,a12778a,a12782a,a12783a,a12784a,a12787a,a12791a,a12792a,a12793a,a12796a,a12800a,a12801a,a12802a,a12805a,a12809a,a12810a,a12811a,a12814a,a12818a,a12819a,a12820a,a12823a,a12827a,a12828a,a12829a,a12832a,a12836a,a12837a,a12838a,a12841a,a12845a,a12846a,a12847a,a12850a,a12854a,a12855a,a12856a,a12859a,a12863a,a12864a,a12865a,a12868a,a12872a,a12873a,a12874a,a12877a,a12881a,a12882a,a12883a,a12886a,a12890a,a12891a,a12892a,a12895a,a12899a,a12900a,a12901a,a12904a,a12908a,a12909a,a12910a,a12913a,a12917a,a12918a,a12919a,a12922a,a12926a,a12927a,a12928a,a12931a,a12935a,a12936a,a12937a,a12940a,a12944a,a12945a,a12946a,a12949a,a12953a,a12954a,a12955a,a12958a,a12962a,a12963a,a12964a,a12967a,a12971a,a12972a,a12973a,a12976a,a12980a,a12981a,a12982a,a12985a,a12989a,a12990a,a12991a,a12994a,a12998a,a12999a,a13000a,a13003a,a13007a,a13008a,a13009a,a13012a,a13016a,a13017a,a13018a,a13021a,a13025a,a13026a,a13027a,a13030a,a13034a,a13035a,a13036a,a13039a,a13043a,a13044a,a13045a,a13048a,a13052a,a13053a,a13054a,a13057a,a13061a,a13062a,a13063a,a13066a,a13070a,a13071a,a13072a,a13075a,a13079a,a13080a,a13081a,a13084a,a13088a,a13089a,a13090a,a13093a,a13097a,a13098a,a13099a,a13102a,a13106a,a13107a,a13108a,a13111a,a13115a,a13116a,a13117a,a13120a,a13124a,a13125a,a13126a,a13129a,a13133a,a13134a,a13135a,a13138a,a13142a,a13143a,a13144a,a13147a,a13151a,a13152a,a13153a,a13156a,a13160a,a13161a,a13162a,a13165a,a13169a,a13170a,a13171a,a13174a,a13178a,a13179a,a13180a,a13183a,a13187a,a13188a,a13189a,a13192a,a13196a,a13197a,a13198a,a13201a,a13205a,a13206a,a13207a,a13210a,a13214a,a13215a,a13216a,a13219a,a13223a,a13224a,a13225a,a13228a,a13232a,a13233a,a13234a,a13237a,a13241a,a13242a,a13243a,a13246a,a13250a,a13251a,a13252a,a13255a,a13259a,a13260a,a13261a,a13264a,a13268a,a13269a,a13270a,a13273a,a13277a,a13278a,a13279a,a13282a,a13286a,a13287a,a13288a,a13291a,a13295a,a13296a,a13297a,a13300a,a13304a,a13305a,a13306a,a13309a,a13313a,a13314a,a13315a,a13318a,a13322a,a13323a,a13324a,a13327a,a13331a,a13332a,a13333a,a13336a,a13340a,a13341a,a13342a,a13345a,a13349a,a13350a,a13351a,a13354a,a13358a,a13359a,a13360a,a13363a,a13367a,a13368a,a13369a,a13372a,a13376a,a13377a,a13378a,a13381a,a13385a,a13386a,a13387a,a13390a,a13394a,a13395a,a13396a,a13399a,a13403a,a13404a,a13405a,a13408a,a13412a,a13413a,a13414a,a13417a,a13421a,a13422a,a13423a,a13426a,a13430a,a13431a,a13432a,a13435a,a13439a,a13440a,a13441a,a13444a,a13448a,a13449a,a13450a,a13453a,a13457a,a13458a,a13459a,a13462a,a13466a,a13467a,a13468a,a13471a,a13475a,a13476a,a13477a,a13480a,a13484a,a13485a,a13486a,a13489a,a13493a,a13494a,a13495a,a13498a,a13502a,a13503a,a13504a,a13507a,a13511a,a13512a,a13513a,a13516a,a13520a,a13521a,a13522a,a13525a,a13529a,a13530a,a13531a,a13534a,a13538a,a13539a,a13540a,a13543a,a13547a,a13548a,a13549a,a13552a,a13556a,a13557a,a13558a,a13561a,a13565a,a13566a,a13567a,a13570a,a13574a,a13575a,a13576a,a13579a,a13583a,a13584a,a13585a,a13588a,a13592a,a13593a,a13594a,a13597a,a13601a,a13602a,a13603a,a13606a,a13610a,a13611a,a13612a,a13615a,a13619a,a13620a,a13621a,a13624a,a13628a,a13629a,a13630a,a13633a,a13637a,a13638a,a13639a,a13642a,a13646a,a13647a,a13648a,a13651a,a13655a,a13656a,a13657a,a13660a,a13664a,a13665a,a13666a,a13669a,a13673a,a13674a,a13675a,a13678a,a13682a,a13683a,a13684a,a13687a,a13691a,a13692a,a13693a,a13696a,a13700a,a13701a,a13702a,a13705a,a13709a,a13710a,a13711a,a13714a,a13718a,a13719a,a13720a,a13723a,a13727a,a13728a,a13729a,a13732a,a13736a,a13737a,a13738a,a13741a,a13745a,a13746a,a13747a,a13750a,a13754a,a13755a,a13756a,a13759a,a13763a,a13764a,a13765a,a13768a,a13772a,a13773a,a13774a,a13777a,a13781a,a13782a,a13783a,a13786a,a13790a,a13791a,a13792a,a13795a,a13799a,a13800a,a13801a,a13804a,a13808a,a13809a,a13810a,a13813a,a13817a,a13818a,a13819a,a13822a,a13826a,a13827a,a13828a,a13831a,a13835a,a13836a,a13837a,a13840a,a13844a,a13845a,a13846a,a13849a,a13853a,a13854a,a13855a,a13858a,a13862a,a13863a,a13864a,a13867a,a13871a,a13872a,a13873a,a13876a,a13880a,a13881a,a13882a,a13885a,a13889a,a13890a,a13891a,a13894a,a13898a,a13899a,a13900a,a13903a,a13907a,a13908a,a13909a,a13912a,a13916a,a13917a,a13918a,a13921a,a13925a,a13926a,a13927a,a13930a,a13934a,a13935a,a13936a,a13939a,a13943a,a13944a,a13945a,a13948a,a13952a,a13953a,a13954a,a13957a,a13961a,a13962a,a13963a,a13966a,a13970a,a13971a,a13972a,a13975a,a13979a,a13980a,a13981a,a13984a,a13988a,a13989a,a13990a,a13993a,a13997a,a13998a,a13999a,a14002a,a14006a,a14007a,a14008a,a14011a,a14015a,a14016a,a14017a,a14020a,a14024a,a14025a,a14026a,a14029a,a14033a,a14034a,a14035a,a14038a,a14042a,a14043a,a14044a,a14047a,a14051a,a14052a,a14053a,a14056a,a14060a,a14061a,a14062a,a14065a,a14069a,a14070a,a14071a,a14074a,a14078a,a14079a,a14080a,a14083a,a14087a,a14088a,a14089a,a14092a,a14096a,a14097a,a14098a,a14101a,a14105a,a14106a,a14107a,a14110a,a14114a,a14115a,a14116a,a14119a,a14123a,a14124a,a14125a,a14128a,a14132a,a14133a,a14134a,a14137a,a14141a,a14142a,a14143a,a14146a,a14150a,a14151a,a14152a,a14155a,a14159a,a14160a,a14161a,a14164a,a14168a,a14169a,a14170a,a14173a,a14177a,a14178a,a14179a,a14182a,a14186a,a14187a,a14188a,a14191a,a14195a,a14196a,a14197a,a14200a,a14204a,a14205a,a14206a,a14209a,a14213a,a14214a,a14215a,a14218a,a14222a,a14223a,a14224a,a14227a,a14231a,a14232a,a14233a,a14236a,a14240a,a14241a,a14242a,a14245a,a14249a,a14250a,a14251a,a14254a,a14258a,a14259a,a14260a,a14263a,a14267a,a14268a,a14269a,a14272a,a14276a,a14277a,a14278a,a14281a,a14285a,a14286a,a14287a,a14290a,a14294a,a14295a,a14296a,a14299a,a14303a,a14304a,a14305a,a14308a,a14312a,a14313a,a14314a,a14317a,a14321a,a14322a,a14323a,a14326a,a14330a,a14331a,a14332a,a14335a,a14339a,a14340a,a14341a,a14344a,a14348a,a14349a,a14350a,a14353a,a14357a,a14358a,a14359a,a14362a,a14366a,a14367a,a14368a,a14371a,a14375a,a14376a,a14377a,a14380a,a14384a,a14385a,a14386a,a14389a,a14393a,a14394a,a14395a,a14398a,a14402a,a14403a,a14404a,a14407a,a14411a,a14412a,a14413a,a14416a,a14420a,a14421a,a14422a,a14425a,a14429a,a14430a,a14431a,a14434a,a14438a,a14439a,a14440a,a14443a,a14447a,a14448a,a14449a,a14452a,a14456a,a14457a,a14458a,a14461a,a14465a,a14466a,a14467a,a14470a,a14474a,a14475a,a14476a,a14479a,a14483a,a14484a,a14485a,a14488a,a14492a,a14493a,a14494a,a14497a,a14501a,a14502a,a14503a,a14506a,a14510a,a14511a,a14512a,a14515a,a14519a,a14520a,a14521a,a14524a,a14528a,a14529a,a14530a,a14533a,a14537a,a14538a,a14539a,a14542a,a14546a,a14547a,a14548a,a14551a,a14555a,a14556a,a14557a,a14560a,a14564a,a14565a,a14566a,a14569a,a14573a,a14574a,a14575a,a14578a,a14582a,a14583a,a14584a,a14587a,a14591a,a14592a,a14593a,a14596a,a14600a,a14601a,a14602a,a14605a,a14609a,a14610a,a14611a,a14614a,a14618a,a14619a,a14620a,a14623a,a14627a,a14628a,a14629a,a14632a,a14636a,a14637a,a14638a,a14641a,a14645a,a14646a,a14647a,a14650a,a14654a,a14655a,a14656a,a14659a,a14663a,a14664a,a14665a,a14668a,a14672a,a14673a,a14674a,a14677a,a14681a,a14682a,a14683a,a14686a,a14690a,a14691a,a14692a,a14695a,a14699a,a14700a,a14701a,a14704a,a14708a,a14709a,a14710a,a14713a,a14717a,a14718a,a14719a,a14722a,a14726a,a14727a,a14728a,a14731a,a14735a,a14736a,a14737a,a14740a,a14744a,a14745a,a14746a,a14749a,a14753a,a14754a,a14755a,a14758a,a14762a,a14763a,a14764a,a14767a,a14771a,a14772a,a14773a,a14776a,a14780a,a14781a,a14782a,a14785a,a14789a,a14790a,a14791a,a14794a,a14798a,a14799a,a14800a,a14803a,a14807a,a14808a,a14809a,a14812a,a14816a,a14817a,a14818a,a14821a,a14825a,a14826a,a14827a,a14830a,a14834a,a14835a,a14836a,a14839a,a14843a,a14844a,a14845a,a14848a,a14852a,a14853a,a14854a,a14857a,a14861a,a14862a,a14863a,a14866a,a14870a,a14871a,a14872a,a14875a,a14879a,a14880a,a14881a,a14884a,a14888a,a14889a,a14890a,a14893a,a14897a,a14898a,a14899a,a14902a,a14906a,a14907a,a14908a,a14911a,a14915a,a14916a,a14917a,a14920a,a14924a,a14925a,a14926a,a14929a,a14933a,a14934a,a14935a,a14938a,a14942a,a14943a,a14944a,a14947a,a14951a,a14952a,a14953a,a14956a,a14960a,a14961a,a14962a,a14965a,a14969a,a14970a,a14971a,a14974a,a14978a,a14979a,a14980a,a14983a,a14987a,a14988a,a14989a,a14992a,a14996a,a14997a,a14998a,a15001a,a15005a,a15006a,a15007a,a15010a,a15014a,a15015a,a15016a,a15019a,a15023a,a15024a,a15025a,a15028a,a15032a,a15033a,a15034a,a15037a,a15041a,a15042a,a15043a,a15046a,a15050a,a15051a,a15052a,a15055a,a15059a,a15060a,a15061a,a15064a,a15068a,a15069a,a15070a,a15073a,a15077a,a15078a,a15079a,a15082a,a15086a,a15087a,a15088a,a15091a,a15095a,a15096a,a15097a,a15100a,a15104a,a15105a,a15106a,a15109a,a15113a,a15114a,a15115a,a15118a,a15122a,a15123a,a15124a,a15127a,a15131a,a15132a,a15133a,a15136a,a15140a,a15141a,a15142a,a15145a,a15149a,a15150a,a15151a,a15154a,a15158a,a15159a,a15160a,a15163a,a15167a,a15168a,a15169a,a15172a,a15176a,a15177a,a15178a,a15181a,a15185a,a15186a,a15187a,a15190a,a15194a,a15195a,a15196a,a15199a,a15203a,a15204a,a15205a,a15208a,a15212a,a15213a,a15214a,a15217a,a15221a,a15222a,a15223a,a15226a,a15230a,a15231a,a15232a,a15235a,a15239a,a15240a,a15241a,a15244a,a15248a,a15249a,a15250a,a15253a,a15257a,a15258a,a15259a,a15262a,a15266a,a15267a,a15268a,a15271a,a15275a,a15276a,a15277a,a15280a,a15284a,a15285a,a15286a,a15289a,a15293a,a15294a,a15295a,a15298a,a15302a,a15303a,a15304a,a15307a,a15311a,a15312a,a15313a,a15316a,a15320a,a15321a,a15322a,a15325a,a15329a,a15330a,a15331a,a15334a,a15338a,a15339a,a15340a,a15343a,a15347a,a15348a,a15349a,a15352a,a15356a,a15357a,a15358a,a15361a,a15365a,a15366a,a15367a,a15370a,a15374a,a15375a,a15376a,a15379a,a15383a,a15384a,a15385a,a15388a,a15392a,a15393a,a15394a,a15397a,a15401a,a15402a,a15403a,a15406a,a15410a,a15411a,a15412a,a15415a,a15419a,a15420a,a15421a,a15424a,a15428a,a15429a,a15430a,a15433a,a15437a,a15438a,a15439a,a15442a,a15446a,a15447a,a15448a,a15451a,a15455a,a15456a,a15457a,a15460a,a15464a,a15465a,a15466a,a15469a,a15473a,a15474a,a15475a,a15478a,a15482a,a15483a,a15484a,a15487a,a15491a,a15492a,a15493a,a15496a,a15500a,a15501a,a15502a,a15505a,a15509a,a15510a,a15511a,a15514a,a15518a,a15519a,a15520a,a15523a,a15527a,a15528a,a15529a,a15532a,a15536a,a15537a,a15538a,a15541a,a15545a,a15546a,a15547a,a15550a,a15554a,a15555a,a15556a,a15559a,a15563a,a15564a,a15565a,a15568a,a15572a,a15573a,a15574a,a15577a,a15581a,a15582a,a15583a,a15586a,a15590a,a15591a,a15592a,a15595a,a15599a,a15600a,a15601a,a15604a,a15608a,a15609a,a15610a,a15613a,a15617a,a15618a,a15619a,a15622a,a15626a,a15627a,a15628a,a15631a,a15635a,a15636a,a15637a,a15640a,a15644a,a15645a,a15646a,a15649a,a15653a,a15654a,a15655a,a15658a,a15662a,a15663a,a15664a,a15667a,a15671a,a15672a,a15673a,a15676a,a15680a,a15681a,a15682a,a15685a,a15689a,a15690a,a15691a,a15694a,a15698a,a15699a,a15700a,a15703a,a15707a,a15708a,a15709a,a15712a,a15716a,a15717a,a15718a,a15721a,a15725a,a15726a,a15727a,a15730a,a15734a,a15735a,a15736a,a15739a,a15743a,a15744a,a15745a,a15748a,a15752a,a15753a,a15754a,a15757a,a15761a,a15762a,a15763a,a15766a,a15770a,a15771a,a15772a,a15775a,a15779a,a15780a,a15781a,a15784a,a15788a,a15789a,a15790a,a15793a,a15797a,a15798a,a15799a,a15802a,a15806a,a15807a,a15808a,a15811a,a15815a,a15816a,a15817a,a15820a,a15824a,a15825a,a15826a,a15829a,a15833a,a15834a,a15835a,a15838a,a15842a,a15843a,a15844a,a15847a,a15851a,a15852a,a15853a,a15856a,a15860a,a15861a,a15862a,a15865a,a15869a,a15870a,a15871a,a15874a,a15878a,a15879a,a15880a,a15883a,a15887a,a15888a,a15889a,a15892a,a15896a,a15897a,a15898a,a15901a,a15905a,a15906a,a15907a,a15910a,a15914a,a15915a,a15916a,a15919a,a15923a,a15924a,a15925a,a15928a,a15932a,a15933a,a15934a,a15937a,a15941a,a15942a,a15943a,a15946a,a15950a,a15951a,a15952a,a15955a,a15959a,a15960a,a15961a,a15964a,a15968a,a15969a,a15970a,a15973a,a15977a,a15978a,a15979a,a15982a,a15986a,a15987a,a15988a,a15991a,a15995a,a15996a,a15997a,a16000a,a16004a,a16005a,a16006a,a16009a,a16013a,a16014a,a16015a,a16018a,a16022a,a16023a,a16024a,a16027a,a16031a,a16032a,a16033a,a16036a,a16040a,a16041a,a16042a,a16045a,a16049a,a16050a,a16051a,a16054a,a16058a,a16059a,a16060a,a16063a,a16067a,a16068a,a16069a,a16072a,a16076a,a16077a,a16078a,a16081a,a16085a,a16086a,a16087a,a16090a,a16094a,a16095a,a16096a,a16099a,a16103a,a16104a,a16105a,a16108a,a16112a,a16113a,a16114a,a16117a,a16121a,a16122a,a16123a,a16126a,a16130a,a16131a,a16132a,a16135a,a16139a,a16140a,a16141a,a16144a,a16148a,a16149a,a16150a,a16153a,a16157a,a16158a,a16159a,a16162a,a16166a,a16167a,a16168a,a16171a,a16175a,a16176a,a16177a,a16180a,a16184a,a16185a,a16186a,a16189a,a16193a,a16194a,a16195a,a16198a,a16202a,a16203a,a16204a,a16207a,a16211a,a16212a,a16213a,a16216a,a16220a,a16221a,a16222a,a16225a,a16229a,a16230a,a16231a,a16234a,a16238a,a16239a,a16240a,a16243a,a16247a,a16248a,a16249a,a16252a,a16256a,a16257a,a16258a,a16261a,a16265a,a16266a,a16267a,a16270a,a16274a,a16275a,a16276a,a16279a,a16283a,a16284a,a16285a,a16288a,a16292a,a16293a,a16294a,a16297a,a16301a,a16302a,a16303a,a16306a,a16310a,a16311a,a16312a,a16315a,a16319a,a16320a,a16321a,a16324a,a16328a,a16329a,a16330a,a16333a,a16337a,a16338a,a16339a,a16342a,a16346a,a16347a,a16348a,a16351a,a16355a,a16356a,a16357a,a16360a,a16364a,a16365a,a16366a,a16369a,a16373a,a16374a,a16375a,a16378a,a16382a,a16383a,a16384a,a16387a,a16391a,a16392a,a16393a,a16396a,a16400a,a16401a,a16402a,a16405a,a16409a,a16410a,a16411a,a16414a,a16418a,a16419a,a16420a,a16423a,a16427a,a16428a,a16429a,a16432a,a16436a,a16437a,a16438a,a16441a,a16445a,a16446a,a16447a,a16450a,a16454a,a16455a,a16456a,a16459a,a16463a,a16464a,a16465a,a16468a,a16472a,a16473a,a16474a,a16477a,a16481a,a16482a,a16483a,a16486a,a16490a,a16491a,a16492a,a16495a,a16499a,a16500a,a16501a,a16504a,a16508a,a16509a,a16510a,a16513a,a16517a,a16518a,a16519a,a16522a,a16526a,a16527a,a16528a,a16531a,a16535a,a16536a,a16537a,a16540a,a16544a,a16545a,a16546a,a16549a,a16553a,a16554a,a16555a,a16558a,a16562a,a16563a,a16564a,a16567a,a16571a,a16572a,a16573a,a16576a,a16580a,a16581a,a16582a,a16585a,a16589a,a16590a,a16591a,a16594a,a16598a,a16599a,a16600a,a16603a,a16607a,a16608a,a16609a,a16612a,a16616a,a16617a,a16618a,a16621a,a16625a,a16626a,a16627a,a16630a,a16634a,a16635a,a16636a,a16639a,a16643a,a16644a,a16645a,a16648a,a16652a,a16653a,a16654a,a16657a,a16661a,a16662a,a16663a,a16666a,a16670a,a16671a,a16672a,a16675a,a16679a,a16680a,a16681a,a16684a,a16688a,a16689a,a16690a,a16693a,a16697a,a16698a,a16699a,a16702a,a16706a,a16707a,a16708a,a16711a,a16715a,a16716a,a16717a,a16720a,a16724a,a16725a,a16726a,a16729a,a16733a,a16734a,a16735a,a16738a,a16742a,a16743a,a16744a,a16747a,a16751a,a16752a,a16753a,a16756a,a16760a,a16761a,a16762a,a16765a,a16769a,a16770a,a16771a,a16774a,a16778a,a16779a,a16780a,a16783a,a16787a,a16788a,a16789a,a16792a,a16796a,a16797a,a16798a,a16801a,a16805a,a16806a,a16807a,a16810a,a16814a,a16815a,a16816a,a16819a,a16823a,a16824a,a16825a,a16829a,a16830a,a16834a,a16835a,a16836a,a16839a,a16843a,a16844a,a16845a,a16849a,a16850a,a16854a,a16855a,a16856a,a16859a,a16863a,a16864a,a16865a,a16869a,a16870a,a16874a,a16875a,a16876a,a16879a,a16883a,a16884a,a16885a,a16889a,a16890a,a16894a,a16895a,a16896a,a16899a,a16903a,a16904a,a16905a,a16909a,a16910a,a16914a,a16915a,a16916a,a16919a,a16923a,a16924a,a16925a,a16929a,a16930a,a16934a,a16935a,a16936a,a16939a,a16943a,a16944a,a16945a,a16949a,a16950a,a16954a,a16955a,a16956a,a16959a,a16963a,a16964a,a16965a,a16969a,a16970a,a16974a,a16975a,a16976a,a16979a,a16983a,a16984a,a16985a,a16989a,a16990a,a16994a,a16995a,a16996a,a16999a,a17003a,a17004a,a17005a,a17009a,a17010a,a17014a,a17015a,a17016a,a17019a,a17023a,a17024a,a17025a,a17029a,a17030a,a17034a,a17035a,a17036a,a17039a,a17043a,a17044a,a17045a,a17049a,a17050a,a17054a,a17055a,a17056a,a17059a,a17063a,a17064a,a17065a,a17069a,a17070a,a17074a,a17075a,a17076a,a17079a,a17083a,a17084a,a17085a,a17089a,a17090a,a17094a,a17095a,a17096a,a17099a,a17103a,a17104a,a17105a,a17109a,a17110a,a17114a,a17115a,a17116a,a17119a,a17123a,a17124a,a17125a,a17129a,a17130a,a17134a,a17135a,a17136a,a17139a,a17143a,a17144a,a17145a,a17149a,a17150a,a17154a,a17155a,a17156a,a17159a,a17163a,a17164a,a17165a,a17169a,a17170a,a17174a,a17175a,a17176a,a17179a,a17183a,a17184a,a17185a,a17189a,a17190a,a17194a,a17195a,a17196a,a17199a,a17203a,a17204a,a17205a,a17209a,a17210a,a17214a,a17215a,a17216a,a17219a,a17223a,a17224a,a17225a,a17229a,a17230a,a17234a,a17235a,a17236a,a17239a,a17243a,a17244a,a17245a,a17249a,a17250a,a17254a,a17255a,a17256a,a17259a,a17263a,a17264a,a17265a,a17269a,a17270a,a17274a,a17275a,a17276a,a17279a,a17283a,a17284a,a17285a,a17289a,a17290a,a17294a,a17295a,a17296a,a17299a,a17303a,a17304a,a17305a,a17309a,a17310a,a17314a,a17315a,a17316a,a17319a,a17323a,a17324a,a17325a,a17329a,a17330a,a17334a,a17335a,a17336a,a17339a,a17343a,a17344a,a17345a,a17349a,a17350a,a17354a,a17355a,a17356a,a17359a,a17363a,a17364a,a17365a,a17369a,a17370a,a17374a,a17375a,a17376a,a17379a,a17383a,a17384a,a17385a,a17389a,a17390a,a17394a,a17395a,a17396a,a17399a,a17403a,a17404a,a17405a,a17409a,a17410a,a17414a,a17415a,a17416a,a17419a,a17423a,a17424a,a17425a,a17429a,a17430a,a17434a,a17435a,a17436a,a17439a,a17443a,a17444a,a17445a,a17449a,a17450a,a17454a,a17455a,a17456a,a17459a,a17463a,a17464a,a17465a,a17469a,a17470a,a17474a,a17475a,a17476a,a17479a,a17483a,a17484a,a17485a,a17489a,a17490a,a17494a,a17495a,a17496a,a17499a,a17503a,a17504a,a17505a,a17509a,a17510a,a17514a,a17515a,a17516a,a17519a,a17523a,a17524a,a17525a,a17529a,a17530a,a17534a,a17535a,a17536a,a17539a,a17543a,a17544a,a17545a,a17549a,a17550a,a17554a,a17555a,a17556a,a17559a,a17563a,a17564a,a17565a,a17569a,a17570a,a17574a,a17575a,a17576a,a17579a,a17583a,a17584a,a17585a,a17589a,a17590a,a17594a,a17595a,a17596a,a17599a,a17603a,a17604a,a17605a,a17609a,a17610a,a17614a,a17615a,a17616a,a17619a,a17623a,a17624a,a17625a,a17629a,a17630a,a17634a,a17635a,a17636a,a17639a,a17643a,a17644a,a17645a,a17649a,a17650a,a17654a,a17655a,a17656a,a17659a,a17663a,a17664a,a17665a,a17669a,a17670a,a17674a,a17675a,a17676a,a17679a,a17683a,a17684a,a17685a,a17689a,a17690a,a17694a,a17695a,a17696a,a17699a,a17703a,a17704a,a17705a,a17709a,a17710a,a17714a,a17715a,a17716a,a17719a,a17723a,a17724a,a17725a,a17729a,a17730a,a17734a,a17735a,a17736a,a17739a,a17743a,a17744a,a17745a,a17749a,a17750a,a17754a,a17755a,a17756a,a17759a,a17763a,a17764a,a17765a,a17769a,a17770a,a17774a,a17775a,a17776a,a17779a,a17783a,a17784a,a17785a,a17789a,a17790a,a17794a,a17795a,a17796a,a17799a,a17803a,a17804a,a17805a,a17809a,a17810a,a17814a,a17815a,a17816a,a17819a,a17823a,a17824a,a17825a,a17829a,a17830a,a17834a,a17835a,a17836a,a17839a,a17843a,a17844a,a17845a,a17849a,a17850a,a17854a,a17855a,a17856a,a17859a,a17863a,a17864a,a17865a,a17869a,a17870a,a17874a,a17875a,a17876a,a17879a,a17883a,a17884a,a17885a,a17889a,a17890a,a17894a,a17895a,a17896a,a17899a,a17903a,a17904a,a17905a,a17909a,a17910a,a17914a,a17915a,a17916a,a17919a,a17923a,a17924a,a17925a,a17929a,a17930a,a17934a,a17935a,a17936a,a17939a,a17943a,a17944a,a17945a,a17949a,a17950a,a17954a,a17955a,a17956a,a17959a,a17963a,a17964a,a17965a,a17969a,a17970a,a17974a,a17975a,a17976a,a17979a,a17983a,a17984a,a17985a,a17989a,a17990a,a17994a,a17995a,a17996a,a17999a,a18003a,a18004a,a18005a,a18009a,a18010a,a18014a,a18015a,a18016a,a18019a,a18023a,a18024a,a18025a,a18029a,a18030a,a18034a,a18035a,a18036a,a18039a,a18043a,a18044a,a18045a,a18049a,a18050a,a18054a,a18055a,a18056a,a18059a,a18063a,a18064a,a18065a,a18069a,a18070a,a18074a,a18075a,a18076a,a18079a,a18083a,a18084a,a18085a,a18089a,a18090a,a18094a,a18095a,a18096a,a18099a,a18103a,a18104a,a18105a,a18109a,a18110a,a18114a,a18115a,a18116a,a18119a,a18123a,a18124a,a18125a,a18129a,a18130a,a18134a,a18135a,a18136a,a18139a,a18143a,a18144a,a18145a,a18149a,a18150a,a18154a,a18155a,a18156a,a18159a,a18163a,a18164a,a18165a,a18169a,a18170a,a18174a,a18175a,a18176a,a18179a,a18183a,a18184a,a18185a,a18189a,a18190a,a18194a,a18195a,a18196a,a18199a,a18203a,a18204a,a18205a,a18209a,a18210a,a18214a,a18215a,a18216a,a18219a,a18223a,a18224a,a18225a,a18229a,a18230a,a18234a,a18235a,a18236a,a18239a,a18243a,a18244a,a18245a,a18249a,a18250a,a18254a,a18255a,a18256a,a18259a,a18263a,a18264a,a18265a,a18269a,a18270a,a18274a,a18275a,a18276a,a18279a,a18283a,a18284a,a18285a,a18289a,a18290a,a18294a,a18295a,a18296a,a18299a,a18303a,a18304a,a18305a,a18309a,a18310a,a18314a,a18315a,a18316a,a18319a,a18323a,a18324a,a18325a,a18329a,a18330a,a18334a,a18335a,a18336a,a18339a,a18343a,a18344a,a18345a,a18349a,a18350a,a18354a,a18355a,a18356a,a18359a,a18363a,a18364a,a18365a,a18369a,a18370a,a18374a,a18375a,a18376a,a18379a,a18383a,a18384a,a18385a,a18389a,a18390a,a18394a,a18395a,a18396a,a18399a,a18403a,a18404a,a18405a,a18409a,a18410a,a18414a,a18415a,a18416a,a18419a,a18423a,a18424a,a18425a,a18429a,a18430a,a18434a,a18435a,a18436a,a18439a,a18443a,a18444a,a18445a,a18449a,a18450a,a18454a,a18455a,a18456a,a18459a,a18463a,a18464a,a18465a,a18469a,a18470a,a18474a,a18475a,a18476a,a18479a,a18483a,a18484a,a18485a,a18489a,a18490a,a18494a,a18495a,a18496a,a18499a,a18503a,a18504a,a18505a,a18509a,a18510a,a18514a,a18515a,a18516a,a18519a,a18523a,a18524a,a18525a,a18529a,a18530a,a18534a,a18535a,a18536a,a18539a,a18543a,a18544a,a18545a,a18549a,a18550a,a18554a,a18555a,a18556a,a18559a,a18563a,a18564a,a18565a,a18569a,a18570a,a18574a,a18575a,a18576a,a18579a,a18583a,a18584a,a18585a,a18589a,a18590a,a18594a,a18595a,a18596a,a18599a,a18603a,a18604a,a18605a,a18609a,a18610a,a18614a,a18615a,a18616a,a18619a,a18623a,a18624a,a18625a,a18629a,a18630a,a18634a,a18635a,a18636a,a18639a,a18643a,a18644a,a18645a,a18649a,a18650a,a18654a,a18655a,a18656a,a18659a,a18663a,a18664a,a18665a,a18669a,a18670a,a18674a,a18675a,a18676a,a18679a,a18683a,a18684a,a18685a,a18689a,a18690a,a18694a,a18695a,a18696a,a18699a,a18703a,a18704a,a18705a,a18709a,a18710a,a18714a,a18715a,a18716a,a18719a,a18723a,a18724a,a18725a,a18729a,a18730a,a18734a,a18735a,a18736a,a18739a,a18743a,a18744a,a18745a,a18749a,a18750a,a18754a,a18755a,a18756a,a18759a,a18763a,a18764a,a18765a,a18769a,a18770a,a18774a,a18775a,a18776a,a18779a,a18783a,a18784a,a18785a,a18789a,a18790a,a18794a,a18795a,a18796a,a18799a,a18803a,a18804a,a18805a,a18809a,a18810a,a18814a,a18815a,a18816a,a18819a,a18823a,a18824a,a18825a,a18829a,a18830a,a18834a,a18835a,a18836a,a18839a,a18843a,a18844a,a18845a,a18849a,a18850a,a18854a,a18855a,a18856a,a18859a,a18863a,a18864a,a18865a,a18869a,a18870a,a18874a,a18875a,a18876a,a18879a,a18883a,a18884a,a18885a,a18889a,a18890a,a18894a,a18895a,a18896a,a18899a,a18903a,a18904a,a18905a,a18909a,a18910a,a18914a,a18915a,a18916a,a18919a,a18923a,a18924a,a18925a,a18929a,a18930a,a18934a,a18935a,a18936a,a18939a,a18943a,a18944a,a18945a,a18949a,a18950a,a18954a,a18955a,a18956a,a18959a,a18963a,a18964a,a18965a,a18969a,a18970a,a18974a,a18975a,a18976a,a18979a,a18983a,a18984a,a18985a,a18989a,a18990a,a18994a,a18995a,a18996a,a18999a,a19003a,a19004a,a19005a,a19009a,a19010a,a19014a,a19015a,a19016a,a19019a,a19023a,a19024a,a19025a,a19029a,a19030a,a19034a,a19035a,a19036a,a19039a,a19043a,a19044a,a19045a,a19049a,a19050a,a19054a,a19055a,a19056a,a19059a,a19063a,a19064a,a19065a,a19069a,a19070a,a19074a,a19075a,a19076a,a19079a,a19083a,a19084a,a19085a,a19089a,a19090a,a19094a,a19095a,a19096a,a19099a,a19103a,a19104a,a19105a,a19109a,a19110a,a19114a,a19115a,a19116a,a19119a,a19123a,a19124a,a19125a,a19129a,a19130a,a19134a,a19135a,a19136a,a19139a,a19143a,a19144a,a19145a,a19149a,a19150a,a19154a,a19155a,a19156a,a19159a,a19163a,a19164a,a19165a,a19169a,a19170a,a19174a,a19175a,a19176a,a19179a,a19183a,a19184a,a19185a,a19189a,a19190a,a19194a,a19195a,a19196a,a19199a,a19203a,a19204a,a19205a,a19209a,a19210a,a19214a,a19215a,a19216a,a19219a,a19223a,a19224a,a19225a,a19229a,a19230a,a19234a,a19235a,a19236a,a19239a,a19243a,a19244a,a19245a,a19249a,a19250a,a19254a,a19255a,a19256a,a19259a,a19263a,a19264a,a19265a,a19269a,a19270a,a19274a,a19275a,a19276a,a19279a,a19283a,a19284a,a19285a,a19289a,a19290a,a19294a,a19295a,a19296a,a19299a,a19303a,a19304a,a19305a,a19309a,a19310a,a19314a,a19315a,a19316a,a19319a,a19323a,a19324a,a19325a,a19329a,a19330a,a19334a,a19335a,a19336a,a19339a,a19343a,a19344a,a19345a,a19349a,a19350a,a19354a,a19355a,a19356a,a19359a,a19363a,a19364a,a19365a,a19369a,a19370a,a19374a,a19375a,a19376a,a19379a,a19383a,a19384a,a19385a,a19389a,a19390a,a19394a,a19395a,a19396a,a19399a,a19403a,a19404a,a19405a,a19409a,a19410a,a19414a,a19415a,a19416a,a19419a,a19423a,a19424a,a19425a,a19429a,a19430a,a19434a,a19435a,a19436a,a19439a,a19443a,a19444a,a19445a,a19449a,a19450a,a19454a,a19455a,a19456a,a19459a,a19463a,a19464a,a19465a,a19469a,a19470a,a19474a,a19475a,a19476a,a19479a,a19483a,a19484a,a19485a,a19489a,a19490a,a19494a,a19495a,a19496a,a19499a,a19503a,a19504a,a19505a,a19509a,a19510a,a19514a,a19515a,a19516a,a19519a,a19523a,a19524a,a19525a,a19529a,a19530a,a19534a,a19535a,a19536a,a19539a,a19543a,a19544a,a19545a,a19549a,a19550a,a19554a,a19555a,a19556a,a19559a,a19563a,a19564a,a19565a,a19569a,a19570a,a19574a,a19575a,a19576a,a19579a,a19583a,a19584a,a19585a,a19589a,a19590a,a19594a,a19595a,a19596a,a19599a,a19603a,a19604a,a19605a,a19609a,a19610a,a19614a,a19615a,a19616a,a19619a,a19623a,a19624a,a19625a,a19629a,a19630a,a19634a,a19635a,a19636a,a19639a,a19643a,a19644a,a19645a,a19649a,a19650a,a19654a,a19655a,a19656a,a19659a,a19663a,a19664a,a19665a,a19669a,a19670a,a19674a,a19675a,a19676a,a19679a,a19683a,a19684a,a19685a,a19689a,a19690a,a19694a,a19695a,a19696a,a19699a,a19703a,a19704a,a19705a,a19709a,a19710a,a19714a,a19715a,a19716a,a19719a,a19723a,a19724a,a19725a,a19729a,a19730a,a19734a,a19735a,a19736a,a19739a,a19743a,a19744a,a19745a,a19749a,a19750a,a19754a,a19755a,a19756a,a19759a,a19763a,a19764a,a19765a,a19769a,a19770a,a19774a,a19775a,a19776a,a19779a,a19783a,a19784a,a19785a,a19789a,a19790a,a19794a,a19795a,a19796a,a19799a,a19803a,a19804a,a19805a,a19809a,a19810a,a19814a,a19815a,a19816a,a19819a,a19823a,a19824a,a19825a,a19829a,a19830a,a19834a,a19835a,a19836a,a19839a,a19843a,a19844a,a19845a,a19849a,a19850a,a19854a,a19855a,a19856a,a19859a,a19863a,a19864a,a19865a,a19869a,a19870a,a19874a,a19875a,a19876a,a19879a,a19883a,a19884a,a19885a,a19889a,a19890a,a19894a,a19895a,a19896a,a19899a,a19903a,a19904a,a19905a,a19909a,a19910a,a19914a,a19915a,a19916a,a19919a,a19923a,a19924a,a19925a,a19929a,a19930a,a19934a,a19935a,a19936a,a19939a,a19943a,a19944a,a19945a,a19949a,a19950a,a19954a,a19955a,a19956a,a19959a,a19963a,a19964a,a19965a,a19969a,a19970a,a19974a,a19975a,a19976a,a19979a,a19983a,a19984a,a19985a,a19989a,a19990a,a19994a,a19995a,a19996a,a19999a,a20003a,a20004a,a20005a,a20009a,a20010a,a20014a,a20015a,a20016a,a20019a,a20023a,a20024a,a20025a,a20029a,a20030a,a20034a,a20035a,a20036a,a20039a,a20043a,a20044a,a20045a,a20049a,a20050a,a20054a,a20055a,a20056a,a20059a,a20063a,a20064a,a20065a,a20069a,a20070a,a20074a,a20075a,a20076a,a20079a,a20083a,a20084a,a20085a,a20089a,a20090a,a20094a,a20095a,a20096a,a20099a,a20103a,a20104a,a20105a,a20109a,a20110a,a20114a,a20115a,a20116a,a20119a,a20123a,a20124a,a20125a,a20129a,a20130a,a20134a,a20135a,a20136a,a20139a,a20143a,a20144a,a20145a,a20149a,a20150a,a20154a,a20155a,a20156a,a20159a,a20163a,a20164a,a20165a,a20169a,a20170a,a20174a,a20175a,a20176a,a20179a,a20183a,a20184a,a20185a,a20189a,a20190a,a20194a,a20195a,a20196a,a20199a,a20203a,a20204a,a20205a,a20209a,a20210a,a20214a,a20215a,a20216a,a20219a,a20223a,a20224a,a20225a,a20229a,a20230a,a20234a,a20235a,a20236a,a20239a,a20243a,a20244a,a20245a,a20249a,a20250a,a20254a,a20255a,a20256a,a20259a,a20263a,a20264a,a20265a,a20269a,a20270a,a20274a,a20275a,a20276a,a20279a,a20283a,a20284a,a20285a,a20289a,a20290a,a20294a,a20295a,a20296a,a20299a,a20303a,a20304a,a20305a,a20309a,a20310a,a20314a,a20315a,a20316a,a20319a,a20323a,a20324a,a20325a,a20329a,a20330a,a20334a,a20335a,a20336a,a20339a,a20343a,a20344a,a20345a,a20349a,a20350a,a20354a,a20355a,a20356a,a20359a,a20363a,a20364a,a20365a,a20369a,a20370a,a20374a,a20375a,a20376a,a20379a,a20383a,a20384a,a20385a,a20389a,a20390a,a20394a,a20395a,a20396a,a20399a,a20403a,a20404a,a20405a,a20409a,a20410a,a20414a,a20415a,a20416a,a20419a,a20423a,a20424a,a20425a,a20429a,a20430a,a20434a,a20435a,a20436a,a20439a,a20443a,a20444a,a20445a,a20449a,a20450a,a20454a,a20455a,a20456a,a20459a,a20463a,a20464a,a20465a,a20469a,a20470a,a20474a,a20475a,a20476a,a20479a,a20483a,a20484a,a20485a,a20489a,a20490a,a20494a,a20495a,a20496a,a20499a,a20503a,a20504a,a20505a,a20509a,a20510a,a20514a,a20515a,a20516a,a20519a,a20523a,a20524a,a20525a,a20529a,a20530a,a20534a,a20535a,a20536a,a20539a,a20543a,a20544a,a20545a,a20549a,a20550a,a20554a,a20555a,a20556a,a20559a,a20563a,a20564a,a20565a,a20569a,a20570a,a20574a,a20575a,a20576a,a20579a,a20583a,a20584a,a20585a,a20589a,a20590a,a20594a,a20595a,a20596a,a20599a,a20603a,a20604a,a20605a,a20609a,a20610a,a20614a,a20615a,a20616a,a20619a,a20623a,a20624a,a20625a,a20629a,a20630a,a20634a,a20635a,a20636a,a20639a,a20643a,a20644a,a20645a,a20649a,a20650a,a20654a,a20655a,a20656a,a20659a,a20663a,a20664a,a20665a,a20669a,a20670a,a20674a,a20675a,a20676a,a20679a,a20683a,a20684a,a20685a,a20689a,a20690a,a20694a,a20695a,a20696a,a20699a,a20703a,a20704a,a20705a,a20709a,a20710a,a20714a,a20715a,a20716a,a20719a,a20723a,a20724a,a20725a,a20729a,a20730a,a20734a,a20735a,a20736a,a20739a,a20743a,a20744a,a20745a,a20749a,a20750a,a20754a,a20755a,a20756a,a20759a,a20763a,a20764a,a20765a,a20769a,a20770a,a20774a,a20775a,a20776a,a20779a,a20783a,a20784a,a20785a,a20789a,a20790a,a20794a,a20795a,a20796a,a20799a,a20803a,a20804a,a20805a,a20809a,a20810a,a20814a,a20815a,a20816a,a20819a,a20823a,a20824a,a20825a,a20829a,a20830a,a20834a,a20835a,a20836a,a20839a,a20843a,a20844a,a20845a,a20849a,a20850a,a20854a,a20855a,a20856a,a20859a,a20863a,a20864a,a20865a,a20869a,a20870a,a20874a,a20875a,a20876a,a20879a,a20883a,a20884a,a20885a,a20889a,a20890a,a20894a,a20895a,a20896a,a20899a,a20903a,a20904a,a20905a,a20909a,a20910a,a20914a,a20915a,a20916a,a20919a,a20923a,a20924a,a20925a,a20929a,a20930a,a20934a,a20935a,a20936a,a20939a,a20943a,a20944a,a20945a,a20949a,a20950a,a20954a,a20955a,a20956a,a20959a,a20963a,a20964a,a20965a,a20969a,a20970a,a20974a,a20975a,a20976a,a20979a,a20983a,a20984a,a20985a,a20989a,a20990a,a20994a,a20995a,a20996a,a20999a,a21003a,a21004a,a21005a,a21009a,a21010a,a21014a,a21015a,a21016a,a21019a,a21023a,a21024a,a21025a,a21029a,a21030a,a21034a,a21035a,a21036a,a21039a,a21043a,a21044a,a21045a,a21049a,a21050a,a21054a,a21055a,a21056a,a21059a,a21063a,a21064a,a21065a,a21069a,a21070a,a21074a,a21075a,a21076a,a21079a,a21083a,a21084a,a21085a,a21089a,a21090a,a21094a,a21095a,a21096a,a21099a,a21103a,a21104a,a21105a,a21109a,a21110a,a21114a,a21115a,a21116a,a21119a,a21123a,a21124a,a21125a,a21129a,a21130a,a21134a,a21135a,a21136a,a21139a,a21143a,a21144a,a21145a,a21149a,a21150a,a21154a,a21155a,a21156a,a21159a,a21163a,a21164a,a21165a,a21169a,a21170a,a21174a,a21175a,a21176a,a21179a,a21183a,a21184a,a21185a,a21189a,a21190a,a21194a,a21195a,a21196a,a21199a,a21203a,a21204a,a21205a,a21209a,a21210a,a21214a,a21215a,a21216a,a21219a,a21223a,a21224a,a21225a,a21229a,a21230a,a21234a,a21235a,a21236a,a21239a,a21243a,a21244a,a21245a,a21249a,a21250a,a21254a,a21255a,a21256a,a21259a,a21263a,a21264a,a21265a,a21269a,a21270a,a21274a,a21275a,a21276a,a21279a,a21283a,a21284a,a21285a,a21289a,a21290a,a21294a,a21295a,a21296a,a21299a,a21303a,a21304a,a21305a,a21309a,a21310a,a21314a,a21315a,a21316a,a21319a,a21323a,a21324a,a21325a,a21329a,a21330a,a21334a,a21335a,a21336a,a21339a,a21343a,a21344a,a21345a,a21349a,a21350a,a21354a,a21355a,a21356a,a21359a,a21363a,a21364a,a21365a,a21369a,a21370a,a21374a,a21375a,a21376a,a21379a,a21383a,a21384a,a21385a,a21389a,a21390a,a21394a,a21395a,a21396a,a21399a,a21403a,a21404a,a21405a,a21409a,a21410a,a21414a,a21415a,a21416a,a21419a,a21423a,a21424a,a21425a,a21429a,a21430a,a21434a,a21435a,a21436a,a21439a,a21443a,a21444a,a21445a,a21449a,a21450a,a21454a,a21455a,a21456a,a21459a,a21463a,a21464a,a21465a,a21469a,a21470a,a21474a,a21475a,a21476a,a21479a,a21483a,a21484a,a21485a,a21489a,a21490a,a21494a,a21495a,a21496a,a21499a,a21503a,a21504a,a21505a,a21509a,a21510a,a21514a,a21515a,a21516a,a21519a,a21523a,a21524a,a21525a,a21529a,a21530a,a21534a,a21535a,a21536a,a21539a,a21543a,a21544a,a21545a,a21549a,a21550a,a21554a,a21555a,a21556a,a21559a,a21563a,a21564a,a21565a,a21569a,a21570a,a21574a,a21575a,a21576a,a21579a,a21583a,a21584a,a21585a,a21589a,a21590a,a21594a,a21595a,a21596a,a21599a,a21603a,a21604a,a21605a,a21609a,a21610a,a21614a,a21615a,a21616a,a21619a,a21623a,a21624a,a21625a,a21629a,a21630a,a21634a,a21635a,a21636a,a21639a,a21643a,a21644a,a21645a,a21649a,a21650a,a21654a,a21655a,a21656a,a21659a,a21663a,a21664a,a21665a,a21669a,a21670a,a21674a,a21675a,a21676a,a21679a,a21683a,a21684a,a21685a,a21689a,a21690a,a21694a,a21695a,a21696a,a21699a,a21703a,a21704a,a21705a,a21709a,a21710a,a21714a,a21715a,a21716a,a21719a,a21723a,a21724a,a21725a,a21729a,a21730a,a21734a,a21735a,a21736a,a21739a,a21743a,a21744a,a21745a,a21749a,a21750a,a21754a,a21755a,a21756a,a21759a,a21763a,a21764a,a21765a,a21769a,a21770a,a21774a,a21775a,a21776a,a21779a,a21783a,a21784a,a21785a,a21789a,a21790a,a21794a,a21795a,a21796a,a21799a,a21803a,a21804a,a21805a,a21809a,a21810a,a21814a,a21815a,a21816a,a21819a,a21823a,a21824a,a21825a,a21829a,a21830a,a21834a,a21835a,a21836a,a21839a,a21843a,a21844a,a21845a,a21849a,a21850a,a21854a,a21855a,a21856a,a21859a,a21863a,a21864a,a21865a,a21869a,a21870a,a21874a,a21875a,a21876a,a21879a,a21883a,a21884a,a21885a,a21889a,a21890a,a21894a,a21895a,a21896a,a21899a,a21903a,a21904a,a21905a,a21909a,a21910a,a21914a,a21915a,a21916a,a21919a,a21923a,a21924a,a21925a,a21929a,a21930a,a21934a,a21935a,a21936a,a21939a,a21943a,a21944a,a21945a,a21949a,a21950a,a21954a,a21955a,a21956a,a21959a,a21963a,a21964a,a21965a,a21969a,a21970a,a21974a,a21975a,a21976a,a21979a,a21983a,a21984a,a21985a,a21989a,a21990a,a21994a,a21995a,a21996a,a21999a,a22003a,a22004a,a22005a,a22009a,a22010a,a22014a,a22015a,a22016a,a22019a,a22023a,a22024a,a22025a,a22029a,a22030a,a22034a,a22035a,a22036a,a22039a,a22043a,a22044a,a22045a,a22049a,a22050a,a22054a,a22055a,a22056a,a22059a,a22063a,a22064a,a22065a,a22069a,a22070a,a22074a,a22075a,a22076a,a22079a,a22083a,a22084a,a22085a,a22089a,a22090a,a22094a,a22095a,a22096a,a22099a,a22103a,a22104a,a22105a,a22109a,a22110a,a22114a,a22115a,a22116a,a22119a,a22123a,a22124a,a22125a,a22129a,a22130a,a22134a,a22135a,a22136a,a22139a,a22143a,a22144a,a22145a,a22149a,a22150a,a22154a,a22155a,a22156a,a22159a,a22163a,a22164a,a22165a,a22169a,a22170a,a22174a,a22175a,a22176a,a22179a,a22183a,a22184a,a22185a,a22189a,a22190a,a22194a,a22195a,a22196a,a22199a,a22203a,a22204a,a22205a,a22209a,a22210a,a22214a,a22215a,a22216a,a22219a,a22223a,a22224a,a22225a,a22229a,a22230a,a22234a,a22235a,a22236a,a22239a,a22243a,a22244a,a22245a,a22249a,a22250a,a22254a,a22255a,a22256a,a22259a,a22263a,a22264a,a22265a,a22269a,a22270a,a22274a,a22275a,a22276a,a22279a,a22283a,a22284a,a22285a,a22289a,a22290a,a22294a,a22295a,a22296a,a22299a,a22303a,a22304a,a22305a,a22309a,a22310a,a22314a,a22315a,a22316a,a22319a,a22323a,a22324a,a22325a,a22329a,a22330a,a22334a,a22335a,a22336a,a22339a,a22343a,a22344a,a22345a,a22349a,a22350a,a22354a,a22355a,a22356a,a22359a,a22363a,a22364a,a22365a,a22369a,a22370a,a22374a,a22375a,a22376a,a22379a,a22383a,a22384a,a22385a,a22389a,a22390a,a22394a,a22395a,a22396a,a22399a,a22403a,a22404a,a22405a,a22409a,a22410a,a22414a,a22415a,a22416a,a22419a,a22423a,a22424a,a22425a,a22429a,a22430a,a22434a,a22435a,a22436a,a22439a,a22443a,a22444a,a22445a,a22449a,a22450a,a22454a,a22455a,a22456a,a22459a,a22463a,a22464a,a22465a,a22469a,a22470a,a22474a,a22475a,a22476a,a22479a,a22483a,a22484a,a22485a,a22489a,a22490a,a22494a,a22495a,a22496a,a22499a,a22503a,a22504a,a22505a,a22509a,a22510a,a22514a,a22515a,a22516a,a22519a,a22523a,a22524a,a22525a,a22529a,a22530a,a22534a,a22535a,a22536a,a22539a,a22543a,a22544a,a22545a,a22549a,a22550a,a22554a,a22555a,a22556a,a22559a,a22563a,a22564a,a22565a,a22569a,a22570a,a22574a,a22575a,a22576a,a22579a,a22583a,a22584a,a22585a,a22589a,a22590a,a22594a,a22595a,a22596a,a22599a,a22603a,a22604a,a22605a,a22609a,a22610a,a22614a,a22615a,a22616a,a22619a,a22623a,a22624a,a22625a,a22629a,a22630a,a22634a,a22635a,a22636a,a22639a,a22643a,a22644a,a22645a,a22649a,a22650a,a22654a,a22655a,a22656a,a22659a,a22663a,a22664a,a22665a,a22669a,a22670a,a22674a,a22675a,a22676a,a22679a,a22683a,a22684a,a22685a,a22689a,a22690a,a22694a,a22695a,a22696a,a22699a,a22703a,a22704a,a22705a,a22709a,a22710a,a22714a,a22715a,a22716a,a22719a,a22723a,a22724a,a22725a,a22729a,a22730a,a22734a,a22735a,a22736a,a22739a,a22743a,a22744a,a22745a,a22749a,a22750a,a22754a,a22755a,a22756a,a22759a,a22763a,a22764a,a22765a,a22769a,a22770a,a22774a,a22775a,a22776a,a22779a,a22783a,a22784a,a22785a,a22789a,a22790a,a22794a,a22795a,a22796a,a22799a,a22803a,a22804a,a22805a,a22809a,a22810a,a22814a,a22815a,a22816a,a22819a,a22823a,a22824a,a22825a,a22829a,a22830a,a22834a,a22835a,a22836a,a22839a,a22843a,a22844a,a22845a,a22849a,a22850a,a22854a,a22855a,a22856a,a22859a,a22863a,a22864a,a22865a,a22869a,a22870a,a22874a,a22875a,a22876a,a22879a,a22883a,a22884a,a22885a,a22889a,a22890a,a22894a,a22895a,a22896a,a22899a,a22903a,a22904a,a22905a,a22909a,a22910a,a22914a,a22915a,a22916a,a22919a,a22923a,a22924a,a22925a,a22929a,a22930a,a22934a,a22935a,a22936a,a22939a,a22943a,a22944a,a22945a,a22949a,a22950a,a22954a,a22955a,a22956a,a22959a,a22963a,a22964a,a22965a,a22969a,a22970a,a22974a,a22975a,a22976a,a22979a,a22983a,a22984a,a22985a,a22989a,a22990a,a22994a,a22995a,a22996a,a22999a,a23003a,a23004a,a23005a,a23009a,a23010a,a23014a,a23015a,a23016a,a23019a,a23023a,a23024a,a23025a,a23029a,a23030a,a23034a,a23035a,a23036a,a23039a,a23043a,a23044a,a23045a,a23049a,a23050a,a23054a,a23055a,a23056a,a23059a,a23063a,a23064a,a23065a,a23069a,a23070a,a23074a,a23075a,a23076a,a23079a,a23083a,a23084a,a23085a,a23089a,a23090a,a23094a,a23095a,a23096a,a23099a,a23103a,a23104a,a23105a,a23109a,a23110a,a23114a,a23115a,a23116a,a23119a,a23123a,a23124a,a23125a,a23129a,a23130a,a23134a,a23135a,a23136a,a23139a,a23143a,a23144a,a23145a,a23149a,a23150a,a23154a,a23155a,a23156a,a23159a,a23163a,a23164a,a23165a,a23169a,a23170a,a23174a,a23175a,a23176a,a23179a,a23183a,a23184a,a23185a,a23189a,a23190a,a23194a,a23195a,a23196a,a23199a,a23203a,a23204a,a23205a,a23209a,a23210a,a23214a,a23215a,a23216a,a23220a,a23221a,a23225a,a23226a,a23227a,a23231a,a23232a,a23236a,a23237a,a23238a,a23242a,a23243a,a23247a,a23248a,a23249a,a23253a,a23254a,a23258a,a23259a,a23260a,a23264a,a23265a,a23269a,a23270a,a23271a,a23275a,a23276a,a23280a,a23281a,a23282a,a23286a,a23287a,a23291a,a23292a,a23293a,a23297a,a23298a,a23302a,a23303a,a23304a,a23308a,a23309a,a23313a,a23314a,a23315a,a23319a,a23320a,a23324a,a23325a,a23326a,a23330a,a23331a,a23335a,a23336a,a23337a,a23341a,a23342a,a23346a,a23347a,a23348a,a23352a,a23353a,a23357a,a23358a,a23359a,a23363a,a23364a,a23368a,a23369a,a23370a,a23374a,a23375a,a23379a,a23380a,a23381a,a23385a,a23386a,a23390a,a23391a,a23392a,a23396a,a23397a,a23401a,a23402a,a23403a,a23407a,a23408a,a23412a,a23413a,a23414a,a23418a,a23419a,a23423a,a23424a,a23425a,a23429a,a23430a,a23434a,a23435a,a23436a,a23440a,a23441a,a23445a,a23446a,a23447a,a23451a,a23452a,a23456a,a23457a,a23458a,a23462a,a23463a,a23467a,a23468a,a23469a,a23473a,a23474a,a23478a,a23479a,a23480a,a23484a,a23485a,a23489a,a23490a,a23491a,a23495a,a23496a,a23500a,a23501a,a23502a,a23506a,a23507a,a23511a,a23512a,a23513a,a23517a,a23518a,a23522a,a23523a,a23524a,a23528a,a23529a,a23533a,a23534a,a23535a,a23539a,a23540a,a23544a,a23545a,a23546a,a23550a,a23551a,a23555a,a23556a,a23557a,a23561a,a23562a,a23566a,a23567a,a23568a,a23572a,a23573a,a23577a,a23578a,a23579a,a23583a,a23584a,a23588a,a23589a,a23590a,a23594a,a23595a,a23599a,a23600a,a23601a,a23605a,a23606a,a23610a,a23611a,a23612a,a23616a,a23617a,a23621a,a23622a,a23623a,a23627a,a23628a,a23632a,a23633a,a23634a,a23638a,a23639a,a23643a,a23644a,a23645a,a23649a,a23650a,a23654a,a23655a,a23656a,a23660a,a23661a,a23665a,a23666a,a23667a,a23671a,a23672a,a23676a,a23677a,a23678a,a23682a,a23683a,a23687a,a23688a,a23689a,a23693a,a23694a,a23698a,a23699a,a23700a,a23704a,a23705a,a23709a,a23710a,a23711a,a23715a,a23716a,a23720a,a23721a,a23722a,a23726a,a23727a,a23731a,a23732a,a23733a,a23737a,a23738a,a23742a,a23743a,a23744a,a23748a,a23749a,a23753a,a23754a,a23755a,a23759a,a23760a,a23764a,a23765a,a23766a,a23770a,a23771a,a23775a,a23776a,a23777a,a23781a,a23782a,a23786a,a23787a,a23788a,a23792a,a23793a,a23797a,a23798a,a23799a,a23803a,a23804a,a23808a,a23809a,a23810a,a23814a,a23815a,a23819a,a23820a,a23821a,a23825a,a23826a,a23830a,a23831a,a23832a,a23836a,a23837a,a23841a,a23842a,a23843a,a23847a,a23848a,a23852a,a23853a,a23854a,a23858a,a23859a,a23863a,a23864a,a23865a,a23869a,a23870a,a23874a,a23875a,a23876a,a23880a,a23881a,a23885a,a23886a,a23887a,a23891a,a23892a,a23896a,a23897a,a23898a,a23902a,a23903a,a23907a,a23908a,a23909a,a23913a,a23914a,a23918a,a23919a,a23920a,a23924a,a23925a,a23929a,a23930a,a23931a,a23935a,a23936a,a23940a,a23941a,a23942a,a23946a,a23947a,a23951a,a23952a,a23953a,a23957a,a23958a,a23962a,a23963a,a23964a,a23968a,a23969a,a23973a,a23974a,a23975a,a23979a,a23980a,a23984a,a23985a,a23986a,a23990a,a23991a,a23995a,a23996a,a23997a,a24001a,a24002a,a24006a,a24007a,a24008a,a24012a,a24013a,a24017a,a24018a,a24019a,a24023a,a24024a,a24028a,a24029a,a24030a,a24034a,a24035a,a24039a,a24040a,a24041a,a24045a,a24046a,a24050a,a24051a,a24052a,a24056a,a24057a,a24061a,a24062a,a24063a,a24067a,a24068a,a24072a,a24073a,a24074a,a24078a,a24079a,a24083a,a24084a,a24085a,a24089a,a24090a,a24094a,a24095a,a24096a,a24100a,a24101a,a24105a,a24106a,a24107a,a24111a,a24112a,a24116a,a24117a,a24118a,a24122a,a24123a,a24127a,a24128a,a24129a,a24133a,a24134a,a24138a,a24139a,a24140a,a24144a,a24145a,a24149a,a24150a,a24151a,a24155a,a24156a,a24160a,a24161a,a24162a,a24166a,a24167a,a24171a,a24172a,a24173a,a24177a,a24178a,a24182a,a24183a,a24184a,a24188a,a24189a,a24193a,a24194a,a24195a,a24199a,a24200a,a24204a,a24205a,a24206a,a24210a,a24211a,a24215a,a24216a,a24217a,a24221a,a24222a,a24226a,a24227a,a24228a,a24232a,a24233a,a24237a,a24238a,a24239a,a24243a,a24244a,a24248a,a24249a,a24250a,a24254a,a24255a,a24259a,a24260a,a24261a,a24265a,a24266a,a24270a,a24271a,a24272a,a24276a,a24277a,a24281a,a24282a,a24283a,a24287a,a24288a,a24292a,a24293a,a24294a,a24298a,a24299a,a24303a,a24304a,a24305a,a24309a,a24310a,a24314a,a24315a,a24316a,a24320a,a24321a,a24325a,a24326a,a24327a,a24331a,a24332a,a24336a,a24337a,a24338a,a24342a,a24343a,a24347a,a24348a,a24349a,a24353a,a24354a,a24358a,a24359a,a24360a,a24364a,a24365a,a24369a,a24370a,a24371a,a24375a,a24376a,a24380a,a24381a,a24382a,a24386a,a24387a,a24391a,a24392a,a24393a,a24397a,a24398a,a24402a,a24403a,a24404a,a24408a,a24409a,a24413a,a24414a,a24415a,a24419a,a24420a,a24424a,a24425a,a24426a,a24430a,a24431a,a24435a,a24436a,a24437a,a24441a,a24442a,a24446a,a24447a,a24448a,a24452a,a24453a,a24457a,a24458a,a24459a,a24463a,a24464a,a24468a,a24469a,a24470a,a24474a,a24475a,a24479a,a24480a,a24481a,a24485a,a24486a,a24490a,a24491a,a24492a,a24496a,a24497a,a24501a,a24502a,a24503a,a24507a,a24508a,a24512a,a24513a,a24514a,a24518a,a24519a,a24523a,a24524a,a24525a,a24529a,a24530a,a24534a,a24535a,a24536a,a24540a,a24541a,a24545a,a24546a,a24547a,a24551a,a24552a,a24556a,a24557a,a24558a,a24562a,a24563a,a24567a,a24568a,a24569a,a24573a,a24574a,a24578a,a24579a,a24580a,a24584a,a24585a,a24589a,a24590a,a24591a,a24595a,a24596a,a24600a,a24601a,a24602a,a24606a,a24607a,a24611a,a24612a,a24613a,a24617a,a24618a,a24622a,a24623a,a24624a,a24628a,a24629a,a24633a,a24634a,a24635a,a24639a,a24640a,a24644a,a24645a,a24646a,a24650a,a24651a,a24655a,a24656a,a24657a,a24661a,a24662a,a24666a,a24667a,a24668a,a24672a,a24673a,a24677a,a24678a,a24679a,a24683a,a24684a,a24688a,a24689a,a24690a,a24694a,a24695a,a24699a,a24700a,a24701a,a24705a,a24706a,a24710a,a24711a,a24712a,a24716a,a24717a,a24721a,a24722a,a24723a,a24727a,a24728a,a24732a,a24733a,a24734a,a24738a,a24739a,a24743a,a24744a,a24745a,a24749a,a24750a,a24754a,a24755a,a24756a,a24760a,a24761a,a24765a,a24766a,a24767a,a24771a,a24772a,a24776a,a24777a,a24778a,a24782a,a24783a,a24787a,a24788a,a24789a,a24793a,a24794a,a24798a,a24799a,a24800a,a24804a,a24805a,a24809a,a24810a,a24811a,a24815a,a24816a,a24820a,a24821a,a24822a,a24826a,a24827a,a24831a,a24832a,a24833a,a24837a,a24838a,a24842a,a24843a,a24844a,a24848a,a24849a,a24853a,a24854a,a24855a,a24859a,a24860a,a24864a,a24865a,a24866a,a24870a,a24871a,a24875a,a24876a,a24877a,a24881a,a24882a,a24886a,a24887a,a24888a,a24892a,a24893a,a24897a,a24898a,a24899a,a24903a,a24904a,a24908a,a24909a,a24910a,a24914a,a24915a,a24919a,a24920a,a24921a,a24925a,a24926a,a24930a,a24931a,a24932a,a24936a,a24937a,a24941a,a24942a,a24943a,a24947a,a24948a,a24952a,a24953a,a24954a,a24958a,a24959a,a24963a,a24964a,a24965a,a24969a,a24970a,a24974a,a24975a,a24976a,a24980a,a24981a,a24985a,a24986a,a24987a,a24991a,a24992a,a24996a,a24997a,a24998a,a25002a,a25003a,a25007a,a25008a,a25009a,a25013a,a25014a,a25018a,a25019a,a25020a,a25024a,a25025a,a25029a,a25030a,a25031a,a25035a,a25036a,a25040a,a25041a,a25042a,a25046a,a25047a,a25051a,a25052a,a25053a,a25057a,a25058a,a25062a,a25063a,a25064a,a25068a,a25069a,a25073a,a25074a,a25075a,a25079a,a25080a,a25084a,a25085a,a25086a,a25090a,a25091a,a25095a,a25096a,a25097a,a25101a,a25102a,a25106a,a25107a,a25108a,a25112a,a25113a,a25117a,a25118a,a25119a,a25123a,a25124a,a25128a,a25129a,a25130a,a25134a,a25135a,a25139a,a25140a,a25141a,a25145a,a25146a,a25150a,a25151a,a25152a,a25156a,a25157a,a25161a,a25162a,a25163a,a25167a,a25168a,a25172a,a25173a,a25174a,a25178a,a25179a,a25183a,a25184a,a25185a,a25189a,a25190a,a25194a,a25195a,a25196a,a25200a,a25201a,a25205a,a25206a,a25207a,a25211a,a25212a,a25216a,a25217a,a25218a,a25222a,a25223a,a25227a,a25228a,a25229a,a25233a,a25234a,a25238a,a25239a,a25240a,a25244a,a25245a,a25249a,a25250a,a25251a,a25255a,a25256a,a25260a,a25261a,a25262a,a25266a,a25267a,a25271a,a25272a,a25273a,a25277a,a25278a,a25282a,a25283a,a25284a,a25288a,a25289a,a25293a,a25294a,a25295a,a25299a,a25300a,a25304a,a25305a,a25306a,a25310a,a25311a,a25315a,a25316a,a25317a,a25321a,a25322a,a25326a,a25327a,a25328a,a25332a,a25333a,a25337a,a25338a,a25339a,a25343a,a25344a,a25348a,a25349a,a25350a,a25354a,a25355a,a25359a,a25360a,a25361a,a25365a,a25366a,a25370a,a25371a,a25372a,a25376a,a25377a,a25381a,a25382a,a25383a,a25387a,a25388a,a25392a,a25393a,a25394a,a25398a,a25399a,a25403a,a25404a,a25405a,a25409a,a25410a,a25414a,a25415a,a25416a,a25420a,a25421a,a25425a,a25426a,a25427a,a25431a,a25432a,a25436a,a25437a,a25438a,a25442a,a25443a,a25447a,a25448a,a25449a,a25453a,a25454a,a25458a,a25459a,a25460a,a25464a,a25465a,a25469a,a25470a,a25471a,a25475a,a25476a,a25480a,a25481a,a25482a,a25486a,a25487a,a25491a,a25492a,a25493a,a25497a,a25498a,a25502a,a25503a,a25504a,a25508a,a25509a,a25513a,a25514a,a25515a,a25519a,a25520a,a25524a,a25525a,a25526a,a25530a,a25531a,a25535a,a25536a,a25537a,a25541a,a25542a,a25546a,a25547a,a25548a,a25552a,a25553a,a25557a,a25558a,a25559a,a25563a,a25564a,a25568a,a25569a,a25570a,a25574a,a25575a,a25579a,a25580a,a25581a,a25585a,a25586a,a25590a,a25591a,a25592a,a25596a,a25597a,a25601a,a25602a,a25603a,a25607a,a25608a,a25612a,a25613a,a25614a,a25618a,a25619a,a25623a,a25624a,a25625a,a25629a,a25630a,a25634a,a25635a,a25636a,a25640a,a25641a,a25645a,a25646a,a25647a,a25651a,a25652a,a25656a,a25657a,a25658a,a25662a,a25663a,a25667a,a25668a,a25669a,a25673a,a25674a,a25678a,a25679a,a25680a,a25684a,a25685a,a25689a,a25690a,a25691a,a25695a,a25696a,a25700a,a25701a,a25702a,a25706a,a25707a,a25711a,a25712a,a25713a,a25717a,a25718a,a25722a,a25723a,a25724a,a25728a,a25729a,a25733a,a25734a,a25735a,a25739a,a25740a,a25744a,a25745a,a25746a,a25750a,a25751a,a25755a,a25756a,a25757a,a25761a,a25762a,a25766a,a25767a,a25768a,a25772a,a25773a,a25777a,a25778a,a25779a,a25783a,a25784a,a25788a,a25789a,a25790a,a25794a,a25795a,a25799a,a25800a,a25801a,a25805a,a25806a,a25810a,a25811a,a25812a,a25816a,a25817a,a25821a,a25822a,a25823a,a25827a,a25828a,a25832a,a25833a,a25834a,a25838a,a25839a,a25843a,a25844a,a25845a,a25849a,a25850a,a25854a,a25855a,a25856a,a25860a,a25861a,a25865a,a25866a,a25867a,a25871a,a25872a,a25876a,a25877a,a25878a,a25882a,a25883a,a25887a,a25888a,a25889a,a25893a,a25894a,a25898a,a25899a,a25900a,a25904a,a25905a,a25909a,a25910a,a25911a,a25915a,a25916a,a25920a,a25921a,a25922a,a25926a,a25927a,a25931a,a25932a,a25933a,a25937a,a25938a,a25942a,a25943a,a25944a,a25948a,a25949a,a25953a,a25954a,a25955a,a25959a,a25960a,a25964a,a25965a,a25966a,a25970a,a25971a,a25975a,a25976a,a25977a,a25981a,a25982a,a25986a,a25987a,a25988a,a25992a,a25993a,a25997a,a25998a,a25999a,a26003a,a26004a,a26008a,a26009a,a26010a,a26014a,a26015a,a26019a,a26020a,a26021a,a26025a,a26026a,a26030a,a26031a,a26032a,a26036a,a26037a,a26041a,a26042a,a26043a,a26047a,a26048a,a26052a,a26053a,a26054a,a26058a,a26059a,a26063a,a26064a,a26065a,a26069a,a26070a,a26074a,a26075a,a26076a,a26080a,a26081a,a26085a,a26086a,a26087a,a26091a,a26092a,a26096a,a26097a,a26098a,a26102a,a26103a,a26107a,a26108a,a26109a,a26113a,a26114a,a26118a,a26119a,a26120a,a26124a,a26125a,a26129a,a26130a,a26131a,a26135a,a26136a,a26140a,a26141a,a26142a,a26146a,a26147a,a26151a,a26152a,a26153a,a26157a,a26158a,a26162a,a26163a,a26164a,a26168a,a26169a,a26173a,a26174a,a26175a,a26179a,a26180a,a26184a,a26185a,a26186a,a26190a,a26191a,a26195a,a26196a,a26197a,a26201a,a26202a,a26206a,a26207a,a26208a,a26212a,a26213a,a26217a,a26218a,a26219a,a26223a,a26224a,a26228a,a26229a,a26230a,a26234a,a26235a,a26239a,a26240a,a26241a,a26245a,a26246a,a26250a,a26251a,a26252a,a26256a,a26257a,a26261a,a26262a,a26263a,a26267a,a26268a,a26272a,a26273a,a26274a,a26278a,a26279a,a26283a,a26284a,a26285a,a26289a,a26290a,a26294a,a26295a,a26296a,a26300a,a26301a,a26305a,a26306a,a26307a,a26311a,a26312a,a26316a,a26317a,a26318a,a26322a,a26323a,a26327a,a26328a,a26329a,a26333a,a26334a,a26338a,a26339a,a26340a,a26344a,a26345a,a26349a,a26350a,a26351a,a26355a,a26356a,a26360a,a26361a,a26362a,a26366a,a26367a,a26371a,a26372a,a26373a,a26377a,a26378a,a26382a,a26383a,a26384a,a26388a,a26389a,a26393a,a26394a,a26395a,a26399a,a26400a,a26404a,a26405a,a26406a,a26410a,a26411a,a26415a,a26416a,a26417a,a26421a,a26422a,a26426a,a26427a,a26428a,a26432a,a26433a,a26437a,a26438a,a26439a,a26443a,a26444a,a26448a,a26449a,a26450a,a26454a,a26455a,a26459a,a26460a,a26461a,a26465a,a26466a,a26470a,a26471a,a26472a,a26476a,a26477a,a26481a,a26482a,a26483a,a26487a,a26488a,a26492a,a26493a,a26494a,a26498a,a26499a,a26503a,a26504a,a26505a,a26509a,a26510a,a26514a,a26515a,a26516a,a26520a,a26521a,a26525a,a26526a,a26527a,a26531a,a26532a,a26536a,a26537a,a26538a,a26542a,a26543a,a26547a,a26548a,a26549a,a26553a,a26554a,a26558a,a26559a,a26560a,a26564a,a26565a,a26569a,a26570a,a26571a,a26575a,a26576a,a26580a,a26581a,a26582a,a26586a,a26587a,a26591a,a26592a,a26593a,a26597a,a26598a,a26602a,a26603a,a26604a,a26608a,a26609a,a26613a,a26614a,a26615a,a26619a,a26620a,a26624a,a26625a,a26626a,a26630a,a26631a,a26635a,a26636a,a26637a,a26641a,a26642a,a26646a,a26647a,a26648a,a26652a,a26653a,a26657a,a26658a,a26659a,a26663a,a26664a,a26668a,a26669a,a26670a,a26674a,a26675a,a26679a,a26680a,a26681a,a26685a,a26686a,a26690a,a26691a,a26692a,a26696a,a26697a,a26701a,a26702a,a26703a,a26707a,a26708a,a26712a,a26713a,a26714a,a26718a,a26719a,a26723a,a26724a,a26725a,a26729a,a26730a,a26734a,a26735a,a26736a,a26740a,a26741a,a26745a,a26746a,a26747a,a26751a,a26752a,a26756a,a26757a,a26758a,a26762a,a26763a,a26767a,a26768a,a26769a,a26773a,a26774a,a26778a,a26779a,a26780a,a26784a,a26785a,a26789a,a26790a,a26791a,a26795a,a26796a,a26800a,a26801a,a26802a,a26806a,a26807a,a26811a,a26812a,a26813a,a26817a,a26818a,a26822a,a26823a,a26824a,a26828a,a26829a,a26833a,a26834a,a26835a,a26839a,a26840a,a26844a,a26845a,a26846a,a26850a,a26851a,a26855a,a26856a,a26857a,a26861a,a26862a,a26866a,a26867a,a26868a,a26872a,a26873a,a26877a,a26878a,a26879a,a26883a,a26884a,a26888a,a26889a,a26890a,a26894a,a26895a,a26899a,a26900a,a26901a,a26905a,a26906a,a26910a,a26911a,a26912a,a26916a,a26917a,a26921a,a26922a,a26923a,a26927a,a26928a,a26932a,a26933a,a26934a,a26938a,a26939a,a26943a,a26944a,a26945a,a26949a,a26950a,a26954a,a26955a,a26956a,a26960a,a26961a,a26965a,a26966a,a26967a,a26971a,a26972a,a26976a,a26977a,a26978a,a26982a,a26983a,a26987a,a26988a,a26989a,a26993a,a26994a,a26998a,a26999a,a27000a,a27004a,a27005a,a27009a,a27010a,a27011a,a27015a,a27016a,a27020a,a27021a,a27022a,a27026a,a27027a,a27031a,a27032a,a27033a,a27037a,a27038a,a27042a,a27043a,a27044a,a27048a,a27049a,a27053a,a27054a,a27055a,a27059a,a27060a,a27064a,a27065a,a27066a,a27070a,a27071a,a27075a,a27076a,a27077a,a27081a,a27082a,a27086a,a27087a,a27088a,a27092a,a27093a,a27097a,a27098a,a27099a,a27103a,a27104a,a27108a,a27109a,a27110a,a27114a,a27115a,a27119a,a27120a,a27121a,a27125a,a27126a,a27130a,a27131a,a27132a,a27136a,a27137a,a27141a,a27142a,a27143a,a27147a,a27148a,a27152a,a27153a,a27154a,a27158a,a27159a,a27163a,a27164a,a27165a,a27169a,a27170a,a27174a,a27175a,a27176a,a27180a,a27181a,a27185a,a27186a,a27187a,a27191a,a27192a,a27196a,a27197a,a27198a,a27202a,a27203a,a27207a,a27208a,a27209a,a27213a,a27214a,a27218a,a27219a,a27220a,a27224a,a27225a,a27229a,a27230a,a27231a,a27235a,a27236a,a27240a,a27241a,a27242a,a27246a,a27247a,a27251a,a27252a,a27253a,a27257a,a27258a,a27262a,a27263a,a27264a,a27268a,a27269a,a27273a,a27274a,a27275a,a27279a,a27280a,a27284a,a27285a,a27286a,a27290a,a27291a,a27295a,a27296a,a27297a,a27301a,a27302a,a27306a,a27307a,a27308a,a27312a,a27313a,a27317a,a27318a,a27319a,a27323a,a27324a,a27328a,a27329a,a27330a,a27334a,a27335a,a27339a,a27340a,a27341a,a27345a,a27346a,a27350a,a27351a,a27352a,a27356a,a27357a,a27361a,a27362a,a27363a,a27367a,a27368a,a27372a,a27373a,a27374a,a27378a,a27379a,a27383a,a27384a,a27385a,a27389a,a27390a,a27394a,a27395a,a27396a,a27400a,a27401a,a27405a,a27406a,a27407a,a27411a,a27412a,a27416a,a27417a,a27418a,a27422a,a27423a,a27427a,a27428a,a27429a,a27433a,a27434a,a27438a,a27439a,a27440a,a27444a,a27445a,a27449a,a27450a,a27451a,a27455a,a27456a,a27460a,a27461a,a27462a,a27466a,a27467a,a27471a,a27472a,a27473a,a27477a,a27478a,a27482a,a27483a,a27484a,a27488a,a27489a,a27493a,a27494a,a27495a,a27499a,a27500a,a27504a,a27505a,a27506a,a27510a,a27511a,a27515a,a27516a,a27517a,a27521a,a27522a,a27526a,a27527a,a27528a,a27532a,a27533a,a27537a,a27538a,a27539a,a27543a,a27544a,a27548a,a27549a,a27550a,a27554a,a27555a,a27559a,a27560a,a27561a,a27565a,a27566a,a27570a,a27571a,a27572a,a27576a,a27577a,a27581a,a27582a,a27583a,a27587a,a27588a,a27592a,a27593a,a27594a,a27598a,a27599a,a27603a,a27604a,a27605a,a27609a,a27610a,a27614a,a27615a,a27616a,a27620a,a27621a,a27625a,a27626a,a27627a,a27631a,a27632a,a27636a,a27637a,a27638a,a27642a,a27643a,a27647a,a27648a,a27649a,a27653a,a27654a,a27658a,a27659a,a27660a,a27664a,a27665a,a27669a,a27670a,a27671a,a27675a,a27676a,a27680a,a27681a,a27682a,a27686a,a27687a,a27691a,a27692a,a27693a,a27697a,a27698a,a27702a,a27703a,a27704a,a27708a,a27709a,a27713a,a27714a,a27715a,a27719a,a27720a,a27724a,a27725a,a27726a,a27730a,a27731a,a27735a,a27736a,a27737a,a27741a,a27742a,a27746a,a27747a,a27748a,a27752a,a27753a,a27757a,a27758a,a27759a,a27763a,a27764a,a27768a,a27769a,a27770a,a27774a,a27775a,a27779a,a27780a,a27781a,a27785a,a27786a,a27790a,a27791a,a27792a,a27796a,a27797a,a27801a,a27802a,a27803a,a27807a,a27808a,a27812a,a27813a,a27814a,a27818a,a27819a,a27823a,a27824a,a27825a,a27829a,a27830a,a27834a,a27835a,a27836a,a27840a,a27841a,a27845a,a27846a,a27847a,a27851a,a27852a,a27856a,a27857a,a27858a,a27862a,a27863a,a27867a,a27868a,a27869a,a27873a,a27874a,a27878a,a27879a,a27880a,a27884a,a27885a,a27889a,a27890a,a27891a,a27895a,a27896a,a27900a,a27901a,a27902a,a27906a,a27907a,a27911a,a27912a,a27913a,a27917a,a27918a,a27922a,a27923a,a27924a,a27928a,a27929a,a27933a,a27934a,a27935a,a27939a,a27940a,a27944a,a27945a,a27946a,a27950a,a27951a,a27955a,a27956a,a27957a,a27961a,a27962a,a27966a,a27967a,a27968a,a27972a,a27973a,a27977a,a27978a,a27979a,a27983a,a27984a,a27988a,a27989a,a27990a,a27994a,a27995a,a27999a,a28000a,a28001a,a28005a,a28006a,a28010a,a28011a,a28012a,a28016a,a28017a,a28021a,a28022a,a28023a,a28027a,a28028a,a28032a,a28033a,a28034a,a28038a,a28039a,a28043a,a28044a,a28045a,a28049a,a28050a,a28054a,a28055a,a28056a,a28060a,a28061a,a28065a,a28066a,a28067a,a28071a,a28072a,a28076a,a28077a,a28078a,a28082a,a28083a,a28087a,a28088a,a28089a,a28093a,a28094a,a28098a,a28099a,a28100a,a28104a,a28105a,a28109a,a28110a,a28111a,a28115a,a28116a,a28120a,a28121a,a28122a,a28126a,a28127a,a28131a,a28132a,a28133a,a28137a,a28138a,a28142a,a28143a,a28144a,a28148a,a28149a,a28153a,a28154a,a28155a,a28159a,a28160a,a28164a,a28165a,a28166a,a28170a,a28171a,a28175a,a28176a,a28177a,a28181a,a28182a,a28186a,a28187a,a28188a,a28192a,a28193a,a28197a,a28198a,a28199a,a28203a,a28204a,a28208a,a28209a,a28210a,a28214a,a28215a,a28219a,a28220a,a28221a,a28225a,a28226a,a28230a,a28231a,a28232a,a28236a,a28237a,a28241a,a28242a,a28243a,a28247a,a28248a,a28252a,a28253a,a28254a,a28258a,a28259a,a28263a,a28264a,a28265a,a28269a,a28270a,a28274a,a28275a,a28276a,a28280a,a28281a,a28285a,a28286a,a28287a,a28291a,a28292a,a28296a,a28297a,a28298a,a28302a,a28303a,a28307a,a28308a,a28309a,a28313a,a28314a,a28318a,a28319a,a28320a,a28324a,a28325a,a28329a,a28330a,a28331a,a28335a,a28336a,a28340a,a28341a,a28342a,a28346a,a28347a,a28351a,a28352a,a28353a,a28357a,a28358a,a28362a,a28363a,a28364a,a28368a,a28369a,a28373a,a28374a,a28375a,a28379a,a28380a,a28384a,a28385a,a28386a,a28390a,a28391a,a28395a,a28396a,a28397a,a28401a,a28402a,a28406a,a28407a,a28408a,a28412a,a28413a,a28417a,a28418a,a28419a,a28423a,a28424a,a28428a,a28429a,a28430a,a28434a,a28435a,a28439a,a28440a,a28441a,a28445a,a28446a,a28450a,a28451a,a28452a,a28456a,a28457a,a28461a,a28462a,a28463a,a28467a,a28468a,a28472a,a28473a,a28474a,a28478a,a28479a,a28483a,a28484a,a28485a,a28489a,a28490a,a28494a,a28495a,a28496a,a28500a,a28501a,a28505a,a28506a,a28507a,a28511a,a28512a,a28516a,a28517a,a28518a,a28522a,a28523a,a28527a,a28528a,a28529a,a28533a,a28534a,a28538a,a28539a,a28540a,a28544a,a28545a,a28549a,a28550a,a28551a,a28555a,a28556a,a28560a,a28561a,a28562a,a28566a,a28567a,a28571a,a28572a,a28573a,a28577a,a28578a,a28582a,a28583a,a28584a,a28588a,a28589a,a28593a,a28594a,a28595a,a28599a,a28600a,a28604a,a28605a,a28606a,a28610a,a28611a,a28615a,a28616a,a28617a,a28621a,a28622a,a28626a,a28627a,a28628a,a28632a,a28633a,a28637a,a28638a,a28639a,a28643a,a28644a,a28648a,a28649a,a28650a,a28654a,a28655a,a28659a,a28660a,a28661a,a28665a,a28666a,a28670a,a28671a,a28672a,a28676a,a28677a,a28681a,a28682a,a28683a,a28687a,a28688a,a28692a,a28693a,a28694a,a28698a,a28699a,a28703a,a28704a,a28705a,a28709a,a28710a,a28714a,a28715a,a28716a,a28720a,a28721a,a28725a,a28726a,a28727a,a28731a,a28732a,a28736a,a28737a,a28738a,a28742a,a28743a,a28747a,a28748a,a28749a,a28753a,a28754a,a28758a,a28759a,a28760a,a28764a,a28765a,a28769a,a28770a,a28771a,a28775a,a28776a,a28780a,a28781a,a28782a,a28786a,a28787a,a28791a,a28792a,a28793a,a28797a,a28798a,a28802a,a28803a,a28804a,a28808a,a28809a,a28813a,a28814a,a28815a,a28819a,a28820a,a28824a,a28825a,a28826a,a28830a,a28831a,a28835a,a28836a,a28837a,a28841a,a28842a,a28846a,a28847a,a28848a,a28852a,a28853a,a28857a,a28858a,a28859a,a28863a,a28864a,a28868a,a28869a,a28870a,a28874a,a28875a,a28879a,a28880a,a28881a,a28885a,a28886a,a28890a,a28891a,a28892a,a28896a,a28897a,a28901a,a28902a,a28903a,a28907a,a28908a,a28912a,a28913a,a28914a,a28918a,a28919a,a28923a,a28924a,a28925a,a28929a,a28930a,a28934a,a28935a,a28936a,a28940a,a28941a,a28945a,a28946a,a28947a,a28951a,a28952a,a28956a,a28957a,a28958a,a28962a,a28963a,a28967a,a28968a,a28969a,a28973a,a28974a,a28978a,a28979a,a28980a,a28984a,a28985a,a28989a,a28990a,a28991a,a28995a,a28996a,a29000a,a29001a,a29002a,a29006a,a29007a,a29011a,a29012a,a29013a,a29017a,a29018a,a29022a,a29023a,a29024a,a29028a,a29029a,a29033a,a29034a,a29035a,a29039a,a29040a,a29044a,a29045a,a29046a,a29050a,a29051a,a29055a,a29056a,a29057a,a29061a,a29062a,a29066a,a29067a,a29068a,a29072a,a29073a,a29077a,a29078a,a29079a,a29083a,a29084a,a29088a,a29089a,a29090a,a29094a,a29095a,a29099a,a29100a,a29101a,a29105a,a29106a,a29110a,a29111a,a29112a,a29116a,a29117a,a29121a,a29122a,a29123a,a29127a,a29128a,a29132a,a29133a,a29134a,a29138a,a29139a,a29143a,a29144a,a29145a,a29149a,a29150a,a29154a,a29155a,a29156a,a29160a,a29161a,a29165a,a29166a,a29167a,a29171a,a29172a,a29176a,a29177a,a29178a,a29182a,a29183a,a29187a,a29188a,a29189a,a29193a,a29194a,a29198a,a29199a,a29200a,a29204a,a29205a,a29209a,a29210a,a29211a,a29215a,a29216a,a29220a,a29221a,a29222a,a29226a,a29227a,a29231a,a29232a,a29233a,a29237a,a29238a,a29242a,a29243a,a29244a,a29248a,a29249a,a29253a,a29254a,a29255a,a29259a,a29260a,a29264a,a29265a,a29266a,a29270a,a29271a,a29275a,a29276a,a29277a,a29281a,a29282a,a29286a,a29287a,a29288a,a29292a,a29293a,a29297a,a29298a,a29299a,a29303a,a29304a,a29308a,a29309a,a29310a,a29314a,a29315a,a29319a,a29320a,a29321a,a29325a,a29326a,a29330a,a29331a,a29332a,a29336a,a29337a,a29341a,a29342a,a29343a,a29347a,a29348a,a29352a,a29353a,a29354a,a29358a,a29359a,a29363a,a29364a,a29365a,a29369a,a29370a,a29374a,a29375a,a29376a,a29380a,a29381a,a29385a,a29386a,a29387a,a29391a,a29392a,a29396a,a29397a,a29398a,a29402a,a29403a,a29407a,a29408a,a29409a,a29413a,a29414a,a29418a,a29419a,a29420a,a29424a,a29425a,a29429a,a29430a,a29431a,a29435a,a29436a,a29440a,a29441a,a29442a,a29446a,a29447a,a29451a,a29452a,a29453a,a29457a,a29458a,a29462a,a29463a,a29464a,a29468a,a29469a,a29473a,a29474a,a29475a,a29479a,a29480a,a29484a,a29485a,a29486a,a29490a,a29491a,a29495a,a29496a,a29497a,a29501a,a29502a,a29506a,a29507a,a29508a,a29512a,a29513a,a29517a,a29518a,a29519a,a29523a,a29524a,a29528a,a29529a,a29530a,a29534a,a29535a,a29539a,a29540a,a29541a,a29545a,a29546a,a29550a,a29551a,a29552a,a29556a,a29557a,a29561a,a29562a,a29563a,a29567a,a29568a,a29572a,a29573a,a29574a,a29578a,a29579a,a29583a,a29584a,a29585a,a29589a,a29590a,a29594a,a29595a,a29596a,a29600a,a29601a,a29605a,a29606a,a29607a,a29611a,a29612a,a29616a,a29617a,a29618a,a29622a,a29623a,a29627a,a29628a,a29629a,a29633a,a29634a,a29638a,a29639a,a29640a,a29644a,a29645a,a29649a,a29650a,a29651a,a29655a,a29656a,a29660a,a29661a,a29662a,a29666a,a29667a,a29671a,a29672a,a29673a,a29677a,a29678a,a29682a,a29683a,a29684a,a29688a,a29689a,a29693a,a29694a,a29695a,a29699a,a29700a,a29704a,a29705a,a29706a,a29710a,a29711a,a29715a,a29716a,a29717a,a29721a,a29722a,a29726a,a29727a,a29728a,a29732a,a29733a,a29737a,a29738a,a29739a,a29743a,a29744a,a29748a,a29749a,a29750a,a29754a,a29755a,a29759a,a29760a,a29761a,a29765a,a29766a,a29770a,a29771a,a29772a,a29776a,a29777a,a29781a,a29782a,a29783a,a29787a,a29788a,a29792a,a29793a,a29794a,a29798a,a29799a,a29803a,a29804a,a29805a,a29809a,a29810a,a29814a,a29815a,a29816a,a29820a,a29821a,a29825a,a29826a,a29827a,a29831a,a29832a,a29836a,a29837a,a29838a,a29842a,a29843a,a29847a,a29848a,a29849a,a29853a,a29854a,a29858a,a29859a,a29860a,a29864a,a29865a,a29869a,a29870a,a29871a,a29875a,a29876a,a29880a,a29881a,a29882a,a29886a,a29887a,a29891a,a29892a,a29893a,a29897a,a29898a,a29902a,a29903a,a29904a,a29908a,a29909a,a29913a,a29914a,a29915a,a29919a,a29920a,a29924a,a29925a,a29926a,a29930a,a29931a,a29935a,a29936a,a29937a,a29941a,a29942a,a29946a,a29947a,a29948a,a29952a,a29953a,a29957a,a29958a,a29959a,a29963a,a29964a,a29968a,a29969a,a29970a,a29974a,a29975a,a29979a,a29980a,a29981a,a29985a,a29986a,a29990a,a29991a,a29992a,a29996a,a29997a,a30001a,a30002a,a30003a,a30007a,a30008a,a30012a,a30013a,a30014a,a30018a,a30019a,a30023a,a30024a,a30025a,a30029a,a30030a,a30034a,a30035a,a30036a,a30040a,a30041a,a30045a,a30046a,a30047a,a30051a,a30052a,a30056a,a30057a,a30058a,a30062a,a30063a,a30067a,a30068a,a30069a,a30073a,a30074a,a30078a,a30079a,a30080a,a30084a,a30085a,a30089a,a30090a,a30091a,a30095a,a30096a,a30100a,a30101a,a30102a,a30106a,a30107a,a30111a,a30112a,a30113a,a30117a,a30118a,a30122a,a30123a,a30124a,a30128a,a30129a,a30133a,a30134a,a30135a,a30139a,a30140a,a30144a,a30145a,a30146a,a30150a,a30151a,a30155a,a30156a,a30157a,a30161a,a30162a,a30166a,a30167a,a30168a,a30172a,a30173a,a30177a,a30178a,a30179a,a30183a,a30184a,a30188a,a30189a,a30190a,a30194a,a30195a,a30199a,a30200a,a30201a,a30205a,a30206a,a30210a,a30211a,a30212a,a30216a,a30217a,a30221a,a30222a,a30223a,a30227a,a30228a,a30232a,a30233a,a30234a,a30238a,a30239a,a30243a,a30244a,a30245a,a30249a,a30250a,a30254a,a30255a,a30256a,a30260a,a30261a,a30265a,a30266a,a30267a,a30271a,a30272a,a30276a,a30277a,a30278a,a30282a,a30283a,a30287a,a30288a,a30289a,a30293a,a30294a,a30298a,a30299a,a30300a,a30304a,a30305a,a30309a,a30310a,a30311a,a30315a,a30316a,a30320a,a30321a,a30322a,a30326a,a30327a,a30331a,a30332a,a30333a,a30337a,a30338a,a30342a,a30343a,a30344a,a30348a,a30349a,a30353a,a30354a,a30355a,a30359a,a30360a,a30364a,a30365a,a30366a,a30370a,a30371a,a30375a,a30376a,a30377a,a30381a,a30382a,a30386a,a30387a,a30388a,a30392a,a30393a,a30397a,a30398a,a30399a,a30403a,a30404a,a30408a,a30409a,a30410a,a30414a,a30415a,a30419a,a30420a,a30421a,a30425a,a30426a,a30430a,a30431a,a30432a,a30436a,a30437a,a30441a,a30442a,a30443a,a30447a,a30448a,a30452a,a30453a,a30454a,a30458a,a30459a,a30463a,a30464a,a30465a,a30469a,a30470a,a30474a,a30475a,a30476a,a30480a,a30481a,a30485a,a30486a,a30487a,a30491a,a30492a,a30496a,a30497a,a30498a,a30502a,a30503a,a30507a,a30508a,a30509a,a30513a,a30514a,a30518a,a30519a,a30520a,a30524a,a30525a,a30529a,a30530a,a30531a,a30535a,a30536a,a30540a,a30541a,a30542a,a30546a,a30547a,a30551a,a30552a,a30553a,a30557a,a30558a,a30562a,a30563a,a30564a,a30568a,a30569a,a30573a,a30574a,a30575a,a30579a,a30580a,a30584a,a30585a,a30586a,a30590a,a30591a,a30595a,a30596a,a30597a,a30601a,a30602a,a30606a,a30607a,a30608a,a30612a,a30613a,a30617a,a30618a,a30619a,a30623a,a30624a,a30628a,a30629a,a30630a,a30634a,a30635a,a30639a,a30640a,a30641a,a30645a,a30646a,a30650a,a30651a,a30652a,a30656a,a30657a,a30661a,a30662a,a30663a,a30667a,a30668a,a30672a,a30673a,a30674a,a30678a,a30679a,a30683a,a30684a,a30685a,a30689a,a30690a,a30694a,a30695a,a30696a,a30700a,a30701a,a30705a,a30706a,a30707a,a30711a,a30712a,a30716a,a30717a,a30718a,a30722a,a30723a,a30727a,a30728a,a30729a,a30733a,a30734a,a30738a,a30739a,a30740a,a30744a,a30745a,a30749a,a30750a,a30751a,a30755a,a30756a,a30760a,a30761a,a30762a,a30766a,a30767a,a30771a,a30772a,a30773a,a30777a,a30778a,a30782a,a30783a,a30784a,a30788a,a30789a,a30793a,a30794a,a30795a,a30799a,a30800a,a30804a,a30805a,a30806a,a30810a,a30811a,a30815a,a30816a,a30817a,a30821a,a30822a,a30826a,a30827a,a30828a,a30832a,a30833a,a30837a,a30838a,a30839a,a30843a,a30844a,a30848a,a30849a,a30850a,a30854a,a30855a,a30859a,a30860a,a30861a,a30865a,a30866a,a30870a,a30871a,a30872a,a30876a,a30877a,a30881a,a30882a,a30883a,a30887a,a30888a,a30892a,a30893a,a30894a,a30898a,a30899a,a30903a,a30904a,a30905a,a30909a,a30910a,a30914a,a30915a,a30916a,a30920a,a30921a,a30925a,a30926a,a30927a,a30931a,a30932a,a30936a,a30937a,a30938a,a30942a,a30943a,a30947a,a30948a,a30949a,a30953a,a30954a,a30958a,a30959a,a30960a,a30964a,a30965a,a30969a,a30970a,a30971a,a30975a,a30976a,a30980a,a30981a,a30982a,a30986a,a30987a,a30991a,a30992a,a30993a,a30997a,a30998a,a31002a,a31003a,a31004a,a31008a,a31009a,a31013a,a31014a,a31015a,a31019a,a31020a,a31024a,a31025a,a31026a,a31030a,a31031a,a31035a,a31036a,a31037a,a31041a,a31042a,a31046a,a31047a,a31048a,a31052a,a31053a,a31057a,a31058a,a31059a,a31063a,a31064a,a31068a,a31069a,a31070a,a31074a,a31075a,a31079a,a31080a,a31081a,a31085a,a31086a,a31090a,a31091a,a31092a,a31096a,a31097a,a31101a,a31102a,a31103a,a31107a,a31108a,a31112a,a31113a,a31114a,a31118a,a31119a,a31123a,a31124a,a31125a,a31129a,a31130a,a31134a,a31135a,a31136a,a31140a,a31141a,a31145a,a31146a,a31147a,a31151a,a31152a,a31156a,a31157a,a31158a,a31162a,a31163a,a31167a,a31168a,a31169a,a31173a,a31174a,a31178a,a31179a,a31180a,a31184a,a31185a,a31189a,a31190a,a31191a,a31195a,a31196a,a31200a,a31201a,a31202a,a31206a,a31207a,a31211a,a31212a,a31213a,a31217a,a31218a,a31222a,a31223a,a31224a,a31228a,a31229a,a31233a,a31234a,a31235a,a31239a,a31240a,a31244a,a31245a,a31246a,a31250a,a31251a,a31255a,a31256a,a31257a,a31261a,a31262a,a31266a,a31267a,a31268a,a31272a,a31273a,a31277a,a31278a,a31279a,a31283a,a31284a,a31288a,a31289a,a31290a,a31294a,a31295a,a31299a,a31300a,a31301a,a31305a,a31306a,a31310a,a31311a,a31312a,a31316a,a31317a,a31321a,a31322a,a31323a,a31327a,a31328a,a31332a,a31333a,a31334a,a31338a,a31339a,a31343a,a31344a,a31345a,a31349a,a31350a,a31354a,a31355a,a31356a,a31360a,a31361a,a31365a,a31366a,a31367a,a31371a,a31372a,a31376a,a31377a,a31378a,a31382a,a31383a,a31387a,a31388a,a31389a,a31393a,a31394a,a31398a,a31399a,a31400a,a31404a,a31405a,a31409a,a31410a,a31411a,a31415a,a31416a,a31420a,a31421a,a31422a,a31426a,a31427a,a31431a,a31432a,a31433a,a31437a,a31438a,a31442a,a31443a,a31444a,a31448a,a31449a,a31453a,a31454a,a31455a,a31459a,a31460a,a31464a,a31465a,a31466a,a31470a,a31471a,a31475a,a31476a,a31477a,a31481a,a31482a,a31486a,a31487a,a31488a,a31492a,a31493a,a31497a,a31498a,a31499a,a31503a,a31504a,a31508a,a31509a,a31510a,a31514a,a31515a,a31519a,a31520a,a31521a,a31525a,a31526a,a31530a,a31531a,a31532a,a31536a,a31537a,a31541a,a31542a,a31543a,a31547a,a31548a,a31552a,a31553a,a31554a,a31558a,a31559a,a31563a,a31564a,a31565a,a31569a,a31570a,a31574a,a31575a,a31576a,a31580a,a31581a,a31585a,a31586a,a31587a,a31591a,a31592a,a31596a,a31597a,a31598a,a31602a,a31603a,a31607a,a31608a,a31609a,a31613a,a31614a,a31618a,a31619a,a31620a,a31624a,a31625a,a31629a,a31630a,a31631a,a31635a,a31636a,a31640a,a31641a,a31642a,a31646a,a31647a,a31651a,a31652a,a31653a,a31657a,a31658a,a31662a,a31663a,a31664a,a31668a,a31669a,a31673a,a31674a,a31675a,a31679a,a31680a,a31684a,a31685a,a31686a,a31690a,a31691a,a31695a,a31696a,a31697a,a31701a,a31702a,a31706a,a31707a,a31708a,a31712a,a31713a,a31717a,a31718a,a31719a,a31723a,a31724a,a31728a,a31729a,a31730a,a31734a,a31735a,a31739a,a31740a,a31741a,a31745a,a31746a,a31750a,a31751a,a31752a,a31756a,a31757a,a31761a,a31762a,a31763a,a31767a,a31768a,a31772a,a31773a,a31774a,a31778a,a31779a,a31783a,a31784a,a31785a,a31789a,a31790a,a31794a,a31795a,a31796a,a31800a,a31801a,a31805a,a31806a,a31807a,a31811a,a31812a,a31816a,a31817a,a31818a,a31822a,a31823a,a31827a,a31828a,a31829a,a31833a,a31834a,a31838a,a31839a,a31840a,a31844a,a31845a,a31849a,a31850a,a31851a,a31855a,a31856a,a31860a,a31861a,a31862a,a31866a,a31867a,a31871a,a31872a,a31873a,a31877a,a31878a,a31882a,a31883a,a31884a,a31888a,a31889a,a31893a,a31894a,a31895a,a31899a,a31900a,a31904a,a31905a,a31906a,a31910a,a31911a,a31915a,a31916a,a31917a,a31921a,a31922a,a31926a,a31927a,a31928a,a31932a,a31933a,a31937a,a31938a,a31939a,a31943a,a31944a,a31948a,a31949a,a31950a,a31954a,a31955a,a31959a,a31960a,a31961a,a31965a,a31966a,a31970a,a31971a,a31972a,a31976a,a31977a,a31981a,a31982a,a31983a,a31987a,a31988a,a31992a,a31993a,a31994a,a31998a,a31999a,a32003a,a32004a,a32005a,a32009a,a32010a,a32014a,a32015a,a32016a,a32020a,a32021a,a32025a,a32026a,a32027a,a32031a,a32032a,a32036a,a32037a,a32038a,a32042a,a32043a,a32047a,a32048a,a32049a,a32053a,a32054a,a32058a,a32059a,a32060a,a32064a,a32065a,a32069a,a32070a,a32071a,a32075a,a32076a,a32080a,a32081a,a32082a,a32086a,a32087a,a32091a,a32092a,a32093a,a32097a,a32098a,a32102a,a32103a,a32104a,a32108a,a32109a,a32113a,a32114a,a32115a,a32119a,a32120a,a32124a,a32125a,a32126a,a32130a,a32131a,a32135a,a32136a,a32137a,a32141a,a32142a,a32146a,a32147a,a32148a,a32152a,a32153a,a32157a,a32158a,a32159a,a32163a,a32164a,a32168a,a32169a,a32170a,a32174a,a32175a,a32179a,a32180a,a32181a,a32185a,a32186a,a32190a,a32191a,a32192a,a32196a,a32197a,a32201a,a32202a,a32203a,a32207a,a32208a,a32212a,a32213a,a32214a,a32218a,a32219a,a32223a,a32224a,a32225a,a32229a,a32230a,a32234a,a32235a,a32236a,a32240a,a32241a,a32245a,a32246a,a32247a,a32251a,a32252a,a32256a,a32257a,a32258a,a32262a,a32263a,a32267a,a32268a,a32269a,a32273a,a32274a,a32278a,a32279a,a32280a,a32284a,a32285a,a32289a,a32290a,a32291a,a32295a,a32296a,a32300a,a32301a,a32302a,a32306a,a32307a,a32311a,a32312a,a32313a,a32317a,a32318a,a32322a,a32323a,a32324a,a32328a,a32329a,a32333a,a32334a,a32335a,a32339a,a32340a,a32344a,a32345a,a32346a,a32350a,a32351a,a32355a,a32356a,a32357a,a32361a,a32362a,a32366a,a32367a,a32368a,a32372a,a32373a,a32377a,a32378a,a32379a,a32383a,a32384a,a32388a,a32389a,a32390a,a32394a,a32395a,a32399a,a32400a,a32401a,a32405a,a32406a,a32410a,a32411a,a32412a,a32416a,a32417a,a32421a,a32422a,a32423a,a32427a,a32428a,a32432a,a32433a,a32434a,a32438a,a32439a,a32443a,a32444a,a32445a,a32449a,a32450a,a32454a,a32455a,a32456a,a32460a,a32461a,a32465a,a32466a,a32467a,a32471a,a32472a,a32476a,a32477a,a32478a,a32482a,a32483a,a32487a,a32488a,a32489a,a32493a,a32494a,a32498a,a32499a,a32500a,a32504a,a32505a,a32509a,a32510a,a32511a,a32515a,a32516a,a32520a,a32521a,a32522a,a32526a,a32527a,a32531a,a32532a,a32533a,a32537a,a32538a,a32542a,a32543a,a32544a,a32548a,a32549a,a32553a,a32554a,a32555a,a32559a,a32560a,a32564a,a32565a,a32566a,a32570a,a32571a,a32575a,a32576a,a32577a,a32581a,a32582a,a32586a,a32587a,a32588a,a32592a,a32593a,a32597a,a32598a,a32599a,a32603a,a32604a,a32608a,a32609a,a32610a,a32614a,a32615a,a32619a,a32620a,a32621a,a32625a,a32626a,a32630a,a32631a,a32632a,a32636a,a32637a,a32641a,a32642a,a32643a,a32647a,a32648a,a32652a,a32653a,a32654a,a32658a,a32659a,a32663a,a32664a,a32665a,a32669a,a32670a,a32674a,a32675a,a32676a,a32680a,a32681a,a32685a,a32686a,a32687a,a32691a,a32692a,a32696a,a32697a,a32698a,a32702a,a32703a,a32707a,a32708a,a32709a,a32713a,a32714a,a32718a,a32719a,a32720a,a32724a,a32725a,a32729a,a32730a,a32731a,a32735a,a32736a,a32740a,a32741a,a32742a,a32746a,a32747a,a32751a,a32752a,a32753a,a32757a,a32758a,a32762a,a32763a,a32764a,a32768a,a32769a,a32773a,a32774a,a32775a,a32779a,a32780a,a32784a,a32785a,a32786a,a32790a,a32791a,a32795a,a32796a,a32797a,a32801a,a32802a,a32806a,a32807a,a32808a,a32812a,a32813a,a32817a,a32818a,a32819a,a32823a,a32824a,a32828a,a32829a,a32830a,a32834a,a32835a,a32839a,a32840a,a32841a,a32845a,a32846a,a32850a,a32851a,a32852a,a32856a,a32857a,a32861a,a32862a,a32863a,a32867a,a32868a,a32872a,a32873a,a32874a,a32878a,a32879a,a32883a,a32884a,a32885a,a32889a,a32890a,a32894a,a32895a,a32896a,a32900a,a32901a,a32905a,a32906a,a32907a,a32911a,a32912a,a32916a,a32917a,a32918a,a32922a,a32923a,a32927a,a32928a,a32929a,a32933a,a32934a,a32938a,a32939a,a32940a,a32944a,a32945a,a32949a,a32950a,a32951a,a32955a,a32956a,a32960a,a32961a,a32962a,a32966a,a32967a,a32971a,a32972a,a32973a,a32977a,a32978a,a32982a,a32983a,a32984a,a32988a,a32989a,a32993a,a32994a,a32995a,a32999a,a33000a,a33004a,a33005a,a33006a,a33010a,a33011a,a33015a,a33016a,a33017a,a33021a,a33022a,a33026a,a33027a,a33028a,a33032a,a33033a,a33037a,a33038a,a33039a,a33043a,a33044a,a33048a,a33049a,a33050a,a33054a,a33055a,a33059a,a33060a,a33061a,a33065a,a33066a,a33070a,a33071a,a33072a,a33076a,a33077a,a33081a,a33082a,a33083a,a33087a,a33088a,a33092a,a33093a,a33094a,a33098a,a33099a,a33103a,a33104a,a33105a,a33109a,a33110a,a33114a,a33115a,a33116a,a33120a,a33121a,a33125a,a33126a,a33127a,a33131a,a33132a,a33136a,a33137a,a33138a,a33142a,a33143a,a33147a,a33148a,a33149a,a33153a,a33154a,a33158a,a33159a,a33160a,a33164a,a33165a,a33169a,a33170a,a33171a,a33175a,a33176a,a33180a,a33181a,a33182a,a33186a,a33187a,a33191a,a33192a,a33193a,a33197a,a33198a,a33202a,a33203a,a33204a,a33208a,a33209a,a33213a,a33214a,a33215a,a33219a,a33220a,a33224a,a33225a,a33226a,a33230a,a33231a,a33235a,a33236a,a33237a,a33241a,a33242a,a33246a,a33247a,a33248a,a33252a,a33253a,a33257a,a33258a,a33259a,a33263a,a33264a,a33268a,a33269a,a33270a,a33274a,a33275a,a33279a,a33280a,a33281a,a33285a,a33286a,a33290a,a33291a,a33292a,a33296a,a33297a,a33301a,a33302a,a33303a,a33307a,a33308a,a33312a,a33313a,a33314a,a33318a,a33319a,a33323a,a33324a,a33325a,a33329a,a33330a,a33334a,a33335a,a33336a,a33340a,a33341a,a33345a,a33346a,a33347a,a33351a,a33352a,a33356a,a33357a,a33358a,a33362a,a33363a,a33367a,a33368a,a33369a,a33373a,a33374a,a33378a,a33379a,a33380a,a33384a,a33385a,a33389a,a33390a,a33391a,a33395a,a33396a,a33400a,a33401a,a33402a,a33406a,a33407a,a33411a,a33412a,a33413a,a33417a,a33418a,a33422a,a33423a,a33424a,a33428a,a33429a,a33433a,a33434a,a33435a,a33439a,a33440a,a33444a,a33445a,a33446a,a33450a,a33451a,a33455a,a33456a,a33457a,a33461a,a33462a,a33466a,a33467a,a33468a,a33472a,a33473a,a33477a,a33478a,a33479a,a33483a,a33484a,a33488a,a33489a,a33490a,a33494a,a33495a,a33499a,a33500a,a33501a,a33505a,a33506a,a33510a,a33511a,a33512a,a33516a,a33517a,a33521a,a33522a,a33523a,a33527a,a33528a,a33532a,a33533a,a33534a,a33538a,a33539a,a33543a,a33544a,a33545a,a33549a,a33550a,a33554a,a33555a,a33556a,a33560a,a33561a,a33565a,a33566a,a33567a,a33571a,a33572a,a33576a,a33577a,a33578a,a33582a,a33583a,a33587a,a33588a,a33589a,a33593a,a33594a,a33598a,a33599a,a33600a,a33604a,a33605a,a33609a,a33610a,a33611a,a33615a,a33616a,a33620a,a33621a,a33622a,a33626a,a33627a,a33631a,a33632a,a33633a,a33637a,a33638a,a33642a,a33643a,a33644a,a33648a,a33649a,a33653a,a33654a,a33655a,a33659a,a33660a,a33664a,a33665a,a33666a,a33670a,a33671a,a33675a,a33676a,a33677a,a33681a,a33682a,a33686a,a33687a,a33688a,a33692a,a33693a,a33697a,a33698a,a33699a,a33703a,a33704a,a33708a,a33709a,a33710a,a33714a,a33715a,a33719a,a33720a,a33721a,a33725a,a33726a,a33730a,a33731a,a33732a,a33736a,a33737a,a33741a,a33742a,a33743a,a33747a,a33748a,a33752a,a33753a,a33754a,a33758a,a33759a,a33763a,a33764a,a33765a,a33769a,a33770a,a33774a,a33775a,a33776a,a33780a,a33781a,a33785a,a33786a,a33787a,a33791a,a33792a,a33796a,a33797a,a33798a,a33802a,a33803a,a33807a,a33808a,a33809a,a33813a,a33814a,a33818a,a33819a,a33820a,a33824a,a33825a,a33829a,a33830a,a33831a,a33835a,a33836a,a33840a,a33841a,a33842a,a33846a,a33847a,a33851a,a33852a,a33853a,a33857a,a33858a,a33862a,a33863a,a33864a,a33868a,a33869a,a33873a,a33874a,a33875a,a33879a,a33880a,a33884a,a33885a,a33886a,a33890a,a33891a,a33895a,a33896a,a33897a,a33901a,a33902a,a33906a,a33907a,a33908a,a33912a,a33913a,a33917a,a33918a,a33919a,a33923a,a33924a,a33928a,a33929a,a33930a,a33934a,a33935a,a33939a,a33940a,a33941a,a33945a,a33946a,a33950a,a33951a,a33952a,a33956a,a33957a,a33961a,a33962a,a33963a,a33967a,a33968a,a33972a,a33973a,a33974a,a33978a,a33979a,a33983a,a33984a,a33985a,a33989a,a33990a,a33994a,a33995a,a33996a,a34000a,a34001a,a34005a,a34006a,a34007a,a34011a,a34012a,a34016a,a34017a,a34018a,a34022a,a34023a,a34027a,a34028a,a34029a,a34033a,a34034a,a34038a,a34039a,a34040a,a34044a,a34045a,a34049a,a34050a,a34051a,a34055a,a34056a,a34060a,a34061a,a34062a,a34066a,a34067a,a34071a,a34072a,a34073a,a34077a,a34078a,a34082a,a34083a,a34084a,a34088a,a34089a,a34093a,a34094a,a34095a,a34099a,a34100a,a34104a,a34105a,a34106a,a34110a,a34111a,a34115a,a34116a,a34117a,a34121a,a34122a,a34126a,a34127a,a34128a,a34132a,a34133a,a34137a,a34138a,a34139a,a34143a,a34144a,a34148a,a34149a,a34150a,a34154a,a34155a,a34159a,a34160a,a34161a,a34165a,a34166a,a34170a,a34171a,a34172a,a34176a,a34177a,a34181a,a34182a,a34183a,a34187a,a34188a,a34192a,a34193a,a34194a,a34198a,a34199a,a34203a,a34204a,a34205a,a34209a,a34210a,a34214a,a34215a,a34216a,a34220a,a34221a,a34225a,a34226a,a34227a,a34231a,a34232a,a34236a,a34237a,a34238a,a34242a,a34243a,a34247a,a34248a,a34249a,a34253a,a34254a,a34258a,a34259a,a34260a,a34264a,a34265a,a34269a,a34270a,a34271a,a34275a,a34276a,a34280a,a34281a,a34282a,a34286a,a34287a,a34291a,a34292a,a34293a,a34297a,a34298a,a34302a,a34303a,a34304a,a34308a,a34309a,a34313a,a34314a,a34315a,a34319a,a34320a,a34324a,a34325a,a34326a,a34330a,a34331a,a34335a,a34336a,a34337a,a34341a,a34342a,a34346a,a34347a,a34348a,a34352a,a34353a,a34357a,a34358a,a34359a,a34363a,a34364a,a34368a,a34369a,a34370a,a34374a,a34375a,a34379a,a34380a,a34381a,a34385a,a34386a,a34390a,a34391a,a34392a,a34396a,a34397a,a34401a,a34402a,a34403a,a34407a,a34408a,a34412a,a34413a,a34414a,a34418a,a34419a,a34423a,a34424a,a34425a,a34429a,a34430a,a34434a,a34435a,a34436a,a34440a,a34441a,a34445a,a34446a,a34447a,a34451a,a34452a,a34456a,a34457a,a34458a,a34462a,a34463a,a34467a,a34468a,a34469a,a34473a,a34474a,a34478a,a34479a,a34480a,a34484a,a34485a,a34489a,a34490a,a34491a,a34495a,a34496a,a34500a,a34501a,a34502a,a34506a,a34507a,a34511a,a34512a,a34513a,a34517a,a34518a,a34522a,a34523a,a34524a,a34528a,a34529a,a34533a,a34534a,a34535a,a34539a,a34540a,a34544a,a34545a,a34546a,a34550a,a34551a,a34555a,a34556a,a34557a,a34561a,a34562a,a34566a,a34567a,a34568a,a34572a,a34573a,a34577a,a34578a,a34579a,a34583a,a34584a,a34588a,a34589a,a34590a,a34594a,a34595a,a34599a,a34600a,a34601a,a34605a,a34606a,a34610a,a34611a,a34612a,a34616a,a34617a,a34621a,a34622a,a34623a,a34627a,a34628a,a34632a,a34633a,a34634a,a34638a,a34639a,a34643a,a34644a,a34645a,a34649a,a34650a,a34654a,a34655a,a34656a,a34660a,a34661a,a34665a,a34666a,a34667a,a34671a,a34672a,a34676a,a34677a,a34678a,a34682a,a34683a,a34687a,a34688a,a34689a,a34693a,a34694a,a34698a,a34699a,a34700a,a34704a,a34705a,a34709a,a34710a,a34711a,a34715a,a34716a,a34720a,a34721a,a34722a,a34726a,a34727a,a34731a,a34732a,a34733a,a34737a,a34738a,a34742a,a34743a,a34744a,a34748a,a34749a,a34753a,a34754a,a34755a,a34759a,a34760a,a34764a,a34765a,a34766a,a34770a,a34771a,a34775a,a34776a,a34777a,a34781a,a34782a,a34786a,a34787a,a34788a,a34792a,a34793a,a34797a,a34798a,a34799a,a34803a,a34804a,a34808a,a34809a,a34810a,a34814a,a34815a,a34819a,a34820a,a34821a,a34825a,a34826a,a34830a,a34831a,a34832a,a34836a,a34837a,a34841a,a34842a,a34843a,a34847a,a34848a,a34852a,a34853a,a34854a,a34858a,a34859a,a34863a,a34864a,a34865a,a34869a,a34870a,a34874a,a34875a,a34876a,a34880a,a34881a,a34885a,a34886a,a34887a,a34891a,a34892a,a34896a,a34897a,a34898a,a34902a,a34903a,a34907a,a34908a,a34909a,a34913a,a34914a,a34918a,a34919a,a34920a,a34924a,a34925a,a34929a,a34930a,a34931a,a34935a,a34936a,a34940a,a34941a,a34942a,a34946a,a34947a,a34951a,a34952a,a34953a,a34957a,a34958a,a34962a,a34963a,a34964a,a34968a,a34969a,a34973a,a34974a,a34975a,a34979a,a34980a,a34984a,a34985a,a34986a,a34990a,a34991a,a34995a,a34996a,a34997a,a35001a,a35002a,a35006a,a35007a,a35008a,a35012a,a35013a,a35017a,a35018a,a35019a,a35023a,a35024a,a35028a,a35029a,a35030a,a35034a,a35035a,a35039a,a35040a,a35041a,a35045a,a35046a,a35050a,a35051a,a35052a,a35056a,a35057a,a35061a,a35062a,a35063a,a35067a,a35068a,a35072a,a35073a,a35074a,a35078a,a35079a,a35083a,a35084a,a35085a,a35089a,a35090a,a35094a,a35095a,a35096a,a35100a,a35101a,a35105a,a35106a,a35107a,a35111a,a35112a,a35116a,a35117a,a35118a,a35122a,a35123a,a35127a,a35128a,a35129a,a35133a,a35134a,a35138a,a35139a,a35140a,a35144a,a35145a,a35149a,a35150a,a35151a,a35155a,a35156a,a35160a,a35161a,a35162a,a35166a,a35167a,a35171a,a35172a,a35173a,a35177a,a35178a,a35182a,a35183a,a35184a,a35188a,a35189a,a35193a,a35194a,a35195a,a35199a,a35200a,a35204a,a35205a,a35206a,a35210a,a35211a,a35215a,a35216a,a35217a,a35221a,a35222a,a35226a,a35227a,a35228a,a35232a,a35233a,a35237a,a35238a,a35239a,a35243a,a35244a,a35248a,a35249a,a35250a,a35254a,a35255a,a35259a,a35260a,a35261a,a35265a,a35266a,a35270a,a35271a,a35272a,a35276a,a35277a,a35281a,a35282a,a35283a,a35287a,a35288a,a35292a,a35293a,a35294a,a35298a,a35299a,a35303a,a35304a,a35305a,a35309a,a35310a,a35314a,a35315a,a35316a,a35320a,a35321a,a35325a,a35326a,a35327a,a35331a,a35332a,a35336a,a35337a,a35338a,a35342a,a35343a,a35347a,a35348a,a35349a,a35353a,a35354a,a35358a,a35359a,a35360a,a35364a,a35365a,a35369a,a35370a,a35371a,a35375a,a35376a,a35380a,a35381a,a35382a,a35386a,a35387a,a35391a,a35392a,a35393a,a35397a,a35398a,a35402a,a35403a,a35404a,a35408a,a35409a,a35413a,a35414a,a35415a,a35419a,a35420a,a35424a,a35425a,a35426a,a35430a,a35431a,a35435a,a35436a,a35437a,a35441a,a35442a,a35446a,a35447a,a35448a,a35452a,a35453a,a35457a,a35458a,a35459a,a35463a,a35464a,a35468a,a35469a,a35470a,a35474a,a35475a,a35479a,a35480a,a35481a,a35485a,a35486a,a35490a,a35491a,a35492a,a35496a,a35497a,a35501a,a35502a,a35503a,a35507a,a35508a,a35512a,a35513a,a35514a,a35518a,a35519a,a35523a,a35524a,a35525a,a35529a,a35530a,a35534a,a35535a,a35536a,a35540a,a35541a,a35545a,a35546a,a35547a,a35551a,a35552a,a35556a,a35557a,a35558a,a35562a,a35563a,a35567a,a35568a,a35569a,a35573a,a35574a,a35578a,a35579a,a35580a,a35584a,a35585a,a35589a,a35590a,a35591a,a35595a,a35596a,a35600a,a35601a,a35602a,a35606a,a35607a,a35611a,a35612a,a35613a,a35617a,a35618a,a35622a,a35623a,a35624a,a35628a,a35629a,a35633a,a35634a,a35635a,a35639a,a35640a,a35644a,a35645a,a35646a,a35650a,a35651a,a35655a,a35656a,a35657a,a35661a,a35662a,a35666a,a35667a,a35668a,a35672a,a35673a,a35677a,a35678a,a35679a,a35683a,a35684a,a35688a,a35689a,a35690a,a35694a,a35695a,a35699a,a35700a,a35701a,a35705a,a35706a,a35710a,a35711a,a35712a,a35716a,a35717a,a35721a,a35722a,a35723a,a35727a,a35728a,a35732a,a35733a,a35734a,a35738a,a35739a,a35743a,a35744a,a35745a,a35749a,a35750a,a35754a,a35755a,a35756a,a35760a,a35761a,a35765a,a35766a,a35767a,a35771a,a35772a,a35776a,a35777a,a35778a,a35782a,a35783a,a35787a,a35788a,a35789a,a35793a,a35794a,a35798a,a35799a,a35800a,a35804a,a35805a,a35809a,a35810a,a35811a,a35815a,a35816a,a35820a,a35821a,a35822a,a35826a,a35827a,a35831a,a35832a,a35833a,a35837a,a35838a,a35842a,a35843a,a35844a,a35848a,a35849a,a35853a,a35854a,a35855a,a35859a,a35860a,a35864a,a35865a,a35866a,a35870a,a35871a,a35875a,a35876a,a35877a,a35881a,a35882a,a35886a,a35887a,a35888a,a35892a,a35893a,a35897a,a35898a,a35899a,a35903a,a35904a,a35908a,a35909a,a35910a,a35914a,a35915a,a35919a,a35920a,a35921a,a35925a,a35926a,a35930a,a35931a,a35932a,a35936a,a35937a,a35941a,a35942a,a35943a,a35947a,a35948a,a35952a,a35953a,a35954a,a35958a,a35959a,a35963a,a35964a,a35965a,a35969a,a35970a,a35974a,a35975a,a35976a,a35980a,a35981a,a35985a,a35986a,a35987a,a35991a,a35992a,a35996a,a35997a,a35998a,a36002a,a36003a,a36007a,a36008a,a36009a,a36013a,a36014a,a36018a,a36019a,a36020a,a36024a,a36025a,a36029a,a36030a,a36031a,a36035a,a36036a,a36040a,a36041a,a36042a,a36046a,a36047a,a36051a,a36052a,a36053a,a36057a,a36058a,a36062a,a36063a,a36064a,a36068a,a36069a,a36073a,a36074a,a36075a,a36079a,a36080a,a36084a,a36085a,a36086a,a36090a,a36091a,a36095a,a36096a,a36097a,a36101a,a36102a,a36106a,a36107a,a36108a,a36112a,a36113a,a36117a,a36118a,a36119a,a36123a,a36124a,a36128a,a36129a,a36130a,a36134a,a36135a,a36139a,a36140a,a36141a,a36145a,a36146a,a36150a,a36151a,a36152a,a36156a,a36157a,a36161a,a36162a,a36163a,a36167a,a36168a,a36172a,a36173a,a36174a,a36178a,a36179a,a36183a,a36184a,a36185a,a36189a,a36190a,a36194a,a36195a,a36196a,a36200a,a36201a,a36205a,a36206a,a36207a,a36211a,a36212a,a36216a,a36217a,a36218a,a36222a,a36223a,a36227a,a36228a,a36229a,a36233a,a36234a,a36238a,a36239a,a36240a,a36244a,a36245a,a36249a,a36250a,a36251a,a36255a,a36256a,a36260a,a36261a,a36262a,a36266a,a36267a,a36271a,a36272a,a36273a,a36277a,a36278a,a36282a,a36283a,a36284a,a36288a,a36289a,a36293a,a36294a,a36295a,a36299a,a36300a,a36304a,a36305a,a36306a,a36310a,a36311a,a36315a,a36316a,a36317a,a36321a,a36322a,a36326a,a36327a,a36328a,a36332a,a36333a,a36337a,a36338a,a36339a,a36343a,a36344a,a36348a,a36349a,a36350a,a36354a,a36355a,a36359a,a36360a,a36361a,a36365a,a36366a,a36370a,a36371a,a36372a,a36376a,a36377a,a36381a,a36382a,a36383a,a36387a,a36388a,a36392a,a36393a,a36394a,a36398a,a36399a,a36403a,a36404a,a36405a,a36409a,a36410a,a36414a,a36415a,a36416a,a36420a,a36421a,a36425a,a36426a,a36427a,a36431a,a36432a,a36436a,a36437a,a36438a,a36442a,a36443a,a36447a,a36448a,a36449a,a36453a,a36454a,a36458a,a36459a,a36460a,a36464a,a36465a,a36469a,a36470a,a36471a,a36475a,a36476a,a36480a,a36481a,a36482a,a36486a,a36487a,a36491a,a36492a,a36493a,a36497a,a36498a,a36502a,a36503a,a36504a,a36508a,a36509a,a36513a,a36514a,a36515a,a36519a,a36520a,a36524a,a36525a,a36526a,a36530a,a36531a,a36535a,a36536a,a36537a,a36541a,a36542a,a36546a,a36547a,a36548a,a36552a,a36553a,a36557a,a36558a,a36559a,a36563a,a36564a,a36568a,a36569a,a36570a,a36574a,a36575a,a36579a,a36580a,a36581a,a36585a,a36586a,a36590a,a36591a,a36592a,a36596a,a36597a,a36601a,a36602a,a36603a,a36607a,a36608a,a36612a,a36613a,a36614a,a36618a,a36619a,a36623a,a36624a,a36625a,a36629a,a36630a,a36634a,a36635a,a36636a,a36640a,a36641a,a36645a,a36646a,a36647a,a36651a,a36652a,a36656a,a36657a,a36658a,a36662a,a36663a,a36667a,a36668a,a36669a,a36673a,a36674a,a36678a,a36679a,a36680a,a36684a,a36685a,a36689a,a36690a,a36691a,a36695a,a36696a,a36700a,a36701a,a36702a,a36706a,a36707a,a36711a,a36712a,a36713a,a36717a,a36718a,a36722a,a36723a,a36724a,a36728a,a36729a,a36733a,a36734a,a36735a,a36739a,a36740a,a36744a,a36745a,a36746a,a36750a,a36751a,a36755a,a36756a,a36757a,a36761a,a36762a,a36766a,a36767a,a36768a,a36772a,a36773a,a36777a,a36778a,a36779a,a36783a,a36784a,a36788a,a36789a,a36790a,a36794a,a36795a,a36799a,a36800a,a36801a,a36805a,a36806a,a36810a,a36811a,a36812a,a36816a,a36817a,a36821a,a36822a,a36823a,a36827a,a36828a,a36832a,a36833a,a36834a,a36838a,a36839a,a36843a,a36844a,a36845a,a36849a,a36850a,a36854a,a36855a,a36856a,a36860a,a36861a,a36865a,a36866a,a36867a,a36871a,a36872a,a36876a,a36877a,a36878a,a36882a,a36883a,a36887a,a36888a,a36889a,a36893a,a36894a,a36898a,a36899a,a36900a,a36904a,a36905a,a36909a,a36910a,a36911a,a36915a,a36916a,a36920a,a36921a,a36922a,a36926a,a36927a,a36931a,a36932a,a36933a,a36937a,a36938a,a36942a,a36943a,a36944a,a36948a,a36949a,a36953a,a36954a,a36955a,a36959a,a36960a,a36964a,a36965a,a36966a,a36970a,a36971a,a36975a,a36976a,a36977a,a36981a,a36982a,a36986a,a36987a,a36988a,a36992a,a36993a,a36997a,a36998a,a36999a,a37003a,a37004a,a37008a,a37009a,a37010a,a37014a,a37015a,a37019a,a37020a,a37021a,a37025a,a37026a,a37030a,a37031a,a37032a,a37036a,a37037a,a37041a,a37042a,a37043a,a37047a,a37048a,a37052a,a37053a,a37054a,a37058a,a37059a,a37063a,a37064a,a37065a,a37069a,a37070a,a37074a,a37075a,a37076a,a37080a,a37081a,a37085a,a37086a,a37087a,a37091a,a37092a,a37096a,a37097a,a37098a,a37102a,a37103a,a37107a,a37108a,a37109a,a37113a,a37114a,a37118a,a37119a,a37120a,a37124a,a37125a,a37129a,a37130a,a37131a,a37135a,a37136a,a37140a,a37141a,a37142a,a37146a,a37147a,a37151a,a37152a,a37153a,a37157a,a37158a,a37162a,a37163a,a37164a,a37168a,a37169a,a37173a,a37174a,a37175a,a37179a,a37180a,a37184a,a37185a,a37186a,a37190a,a37191a,a37195a,a37196a,a37197a,a37201a,a37202a,a37206a,a37207a,a37208a,a37212a,a37213a,a37217a,a37218a,a37219a,a37223a,a37224a,a37228a,a37229a,a37230a,a37234a,a37235a,a37239a,a37240a,a37241a,a37245a,a37246a,a37250a,a37251a,a37252a,a37256a,a37257a,a37261a,a37262a,a37263a,a37267a,a37268a,a37272a,a37273a,a37274a,a37278a,a37279a,a37283a,a37284a,a37285a,a37289a,a37290a,a37294a,a37295a,a37296a,a37300a,a37301a,a37305a,a37306a,a37307a,a37311a,a37312a,a37316a,a37317a,a37318a,a37322a,a37323a,a37327a,a37328a,a37329a,a37333a,a37334a,a37338a,a37339a,a37340a,a37344a,a37345a,a37349a,a37350a,a37351a,a37355a,a37356a,a37360a,a37361a,a37362a,a37366a,a37367a,a37371a,a37372a,a37373a,a37377a,a37378a,a37382a,a37383a,a37384a,a37388a,a37389a,a37393a,a37394a,a37395a,a37399a,a37400a,a37404a,a37405a,a37406a,a37410a,a37411a,a37415a,a37416a,a37417a,a37421a,a37422a,a37426a,a37427a,a37428a,a37432a,a37433a,a37437a,a37438a,a37439a,a37443a,a37444a,a37448a,a37449a,a37450a,a37454a,a37455a,a37459a,a37460a,a37461a,a37465a,a37466a,a37470a,a37471a,a37472a,a37476a,a37477a,a37481a,a37482a,a37483a,a37487a,a37488a,a37492a,a37493a,a37494a,a37498a,a37499a,a37503a,a37504a,a37505a,a37509a,a37510a,a37514a,a37515a,a37516a,a37520a,a37521a,a37525a,a37526a,a37527a,a37531a,a37532a,a37536a,a37537a,a37538a,a37542a,a37543a,a37547a,a37548a,a37549a,a37553a,a37554a,a37558a,a37559a,a37560a,a37564a,a37565a,a37569a,a37570a,a37571a,a37575a,a37576a,a37580a,a37581a,a37582a,a37586a,a37587a,a37591a,a37592a,a37593a,a37597a,a37598a,a37602a,a37603a,a37604a,a37608a,a37609a,a37613a,a37614a,a37615a,a37619a,a37620a,a37624a,a37625a,a37626a,a37630a,a37631a,a37635a,a37636a,a37637a,a37641a,a37642a,a37646a,a37647a,a37648a,a37652a,a37653a,a37657a,a37658a,a37659a,a37663a,a37664a,a37667a,a37670a,a37671a,a37672a,a37676a,a37677a,a37681a,a37682a,a37683a,a37687a,a37688a,a37691a,a37694a,a37695a,a37696a,a37700a,a37701a,a37705a,a37706a,a37707a,a37711a,a37712a,a37715a,a37718a,a37719a,a37720a,a37724a,a37725a,a37729a,a37730a,a37731a,a37735a,a37736a,a37739a,a37742a,a37743a,a37744a,a37748a,a37749a,a37753a,a37754a,a37755a,a37759a,a37760a,a37763a,a37766a,a37767a,a37768a,a37772a,a37773a,a37777a,a37778a,a37779a,a37783a,a37784a,a37787a,a37790a,a37791a,a37792a,a37796a,a37797a,a37801a,a37802a,a37803a,a37807a,a37808a,a37811a,a37814a,a37815a,a37816a,a37820a,a37821a,a37825a,a37826a,a37827a,a37831a,a37832a,a37835a,a37838a,a37839a,a37840a,a37844a,a37845a,a37849a,a37850a,a37851a,a37855a,a37856a,a37859a,a37862a,a37863a,a37864a,a37868a,a37869a,a37873a,a37874a,a37875a,a37879a,a37880a,a37883a,a37886a,a37887a,a37888a,a37892a,a37893a,a37897a,a37898a,a37899a,a37903a,a37904a,a37907a,a37910a,a37911a,a37912a,a37916a,a37917a,a37921a,a37922a,a37923a,a37927a,a37928a,a37931a,a37934a,a37935a,a37936a,a37940a,a37941a,a37945a,a37946a,a37947a,a37951a,a37952a,a37955a,a37958a,a37959a,a37960a,a37964a,a37965a,a37969a,a37970a,a37971a,a37975a,a37976a,a37979a,a37982a,a37983a,a37984a,a37988a,a37989a,a37993a,a37994a,a37995a,a37999a,a38000a,a38003a,a38006a,a38007a,a38008a,a38012a,a38013a,a38017a,a38018a,a38019a,a38023a,a38024a,a38027a,a38030a,a38031a,a38032a,a38036a,a38037a,a38041a,a38042a,a38043a,a38047a,a38048a,a38051a,a38054a,a38055a,a38056a,a38060a,a38061a,a38065a,a38066a,a38067a,a38071a,a38072a,a38075a,a38078a,a38079a,a38080a,a38084a,a38085a,a38089a,a38090a,a38091a,a38095a,a38096a,a38099a,a38102a,a38103a,a38104a,a38108a,a38109a,a38113a,a38114a,a38115a,a38119a,a38120a,a38123a,a38126a,a38127a,a38128a,a38132a,a38133a,a38137a,a38138a,a38139a,a38143a,a38144a,a38147a,a38150a,a38151a,a38152a,a38156a,a38157a,a38161a,a38162a,a38163a,a38167a,a38168a,a38171a,a38174a,a38175a,a38176a,a38180a,a38181a,a38185a,a38186a,a38187a,a38191a,a38192a,a38195a,a38198a,a38199a,a38200a,a38204a,a38205a,a38209a,a38210a,a38211a,a38215a,a38216a,a38219a,a38222a,a38223a,a38224a,a38228a,a38229a,a38233a,a38234a,a38235a,a38239a,a38240a,a38243a,a38246a,a38247a,a38248a,a38252a,a38253a,a38257a,a38258a,a38259a,a38263a,a38264a,a38267a,a38270a,a38271a,a38272a,a38276a,a38277a,a38281a,a38282a,a38283a,a38287a,a38288a,a38291a,a38294a,a38295a,a38296a,a38300a,a38301a,a38305a,a38306a,a38307a,a38311a,a38312a,a38315a,a38318a,a38319a,a38320a,a38324a,a38325a,a38329a,a38330a,a38331a,a38335a,a38336a,a38339a,a38342a,a38343a,a38344a,a38348a,a38349a,a38353a,a38354a,a38355a,a38359a,a38360a,a38363a,a38366a,a38367a,a38368a,a38372a,a38373a,a38377a,a38378a,a38379a,a38383a,a38384a,a38387a,a38390a,a38391a,a38392a,a38396a,a38397a,a38401a,a38402a,a38403a,a38407a,a38408a,a38411a,a38414a,a38415a,a38416a,a38420a,a38421a,a38425a,a38426a,a38427a,a38431a,a38432a,a38435a,a38438a,a38439a,a38440a,a38444a,a38445a,a38449a,a38450a,a38451a,a38455a,a38456a,a38459a,a38462a,a38463a,a38464a,a38468a,a38469a,a38473a,a38474a,a38475a,a38479a,a38480a,a38483a,a38486a,a38487a,a38488a,a38492a,a38493a,a38497a,a38498a,a38499a,a38503a,a38504a,a38507a,a38510a,a38511a,a38512a,a38516a,a38517a,a38521a,a38522a,a38523a,a38527a,a38528a,a38531a,a38534a,a38535a,a38536a,a38540a,a38541a,a38545a,a38546a,a38547a,a38551a,a38552a,a38555a,a38558a,a38559a,a38560a,a38564a,a38565a,a38569a,a38570a,a38571a,a38575a,a38576a,a38579a,a38582a,a38583a,a38584a,a38588a,a38589a,a38593a,a38594a,a38595a,a38599a,a38600a,a38603a,a38606a,a38607a,a38608a,a38612a,a38613a,a38617a,a38618a,a38619a,a38623a,a38624a,a38627a,a38630a,a38631a,a38632a,a38636a,a38637a,a38641a,a38642a,a38643a,a38647a,a38648a,a38651a,a38654a,a38655a,a38656a,a38660a,a38661a,a38665a,a38666a,a38667a,a38671a,a38672a,a38675a,a38678a,a38679a,a38680a,a38684a,a38685a,a38689a,a38690a,a38691a,a38695a,a38696a,a38699a,a38702a,a38703a,a38704a,a38708a,a38709a,a38713a,a38714a,a38715a,a38719a,a38720a,a38723a,a38726a,a38727a,a38728a,a38732a,a38733a,a38737a,a38738a,a38739a,a38743a,a38744a,a38747a,a38750a,a38751a,a38752a,a38756a,a38757a,a38761a,a38762a,a38763a,a38767a,a38768a,a38771a,a38774a,a38775a,a38776a,a38780a,a38781a,a38785a,a38786a,a38787a,a38791a,a38792a,a38795a,a38798a,a38799a,a38800a,a38804a,a38805a,a38809a,a38810a,a38811a,a38815a,a38816a,a38819a,a38822a,a38823a,a38824a,a38828a,a38829a,a38833a,a38834a,a38835a,a38839a,a38840a,a38843a,a38846a,a38847a,a38848a,a38852a,a38853a,a38857a,a38858a,a38859a,a38863a,a38864a,a38867a,a38870a,a38871a,a38872a,a38876a,a38877a,a38881a,a38882a,a38883a,a38887a,a38888a,a38891a,a38894a,a38895a,a38896a,a38900a,a38901a,a38905a,a38906a,a38907a,a38911a,a38912a,a38915a,a38918a,a38919a,a38920a,a38924a,a38925a,a38929a,a38930a,a38931a,a38935a,a38936a,a38939a,a38942a,a38943a,a38944a,a38948a,a38949a,a38953a,a38954a,a38955a,a38959a,a38960a,a38963a,a38966a,a38967a,a38968a,a38972a,a38973a,a38977a,a38978a,a38979a,a38983a,a38984a,a38987a,a38990a,a38991a,a38992a,a38996a,a38997a,a39001a,a39002a,a39003a,a39007a,a39008a,a39011a,a39014a,a39015a,a39016a,a39020a,a39021a,a39025a,a39026a,a39027a,a39031a,a39032a,a39035a,a39038a,a39039a,a39040a,a39044a,a39045a,a39049a,a39050a,a39051a,a39055a,a39056a,a39059a,a39062a,a39063a,a39064a,a39068a,a39069a,a39073a,a39074a,a39075a,a39079a,a39080a,a39083a,a39086a,a39087a,a39088a,a39092a,a39093a,a39097a,a39098a,a39099a,a39103a,a39104a,a39107a,a39110a,a39111a,a39112a,a39116a,a39117a,a39121a,a39122a,a39123a,a39127a,a39128a,a39131a,a39134a,a39135a,a39136a,a39140a,a39141a,a39145a,a39146a,a39147a,a39151a,a39152a,a39155a,a39158a,a39159a,a39160a,a39164a,a39165a,a39169a,a39170a,a39171a,a39175a,a39176a,a39179a,a39182a,a39183a,a39184a,a39188a,a39189a,a39193a,a39194a,a39195a,a39199a,a39200a,a39203a,a39206a,a39207a,a39208a,a39212a,a39213a,a39217a,a39218a,a39219a,a39223a,a39224a,a39227a,a39230a,a39231a,a39232a,a39236a,a39237a,a39241a,a39242a,a39243a,a39247a,a39248a,a39251a,a39254a,a39255a,a39256a,a39260a,a39261a,a39265a,a39266a,a39267a,a39271a,a39272a,a39275a,a39278a,a39279a,a39280a,a39284a,a39285a,a39289a,a39290a,a39291a,a39295a,a39296a,a39299a,a39302a,a39303a,a39304a,a39308a,a39309a,a39313a,a39314a,a39315a,a39319a,a39320a,a39323a,a39326a,a39327a,a39328a,a39332a,a39333a,a39337a,a39338a,a39339a,a39343a,a39344a,a39347a,a39350a,a39351a,a39352a,a39356a,a39357a,a39361a,a39362a,a39363a,a39367a,a39368a,a39371a,a39374a,a39375a,a39376a,a39380a,a39381a,a39385a,a39386a,a39387a,a39391a,a39392a,a39395a,a39398a,a39399a,a39400a,a39404a,a39405a,a39409a,a39410a,a39411a,a39415a,a39416a,a39419a,a39422a,a39423a,a39424a,a39428a,a39429a,a39433a,a39434a,a39435a,a39439a,a39440a,a39443a,a39446a,a39447a,a39448a,a39452a,a39453a,a39457a,a39458a,a39459a,a39463a,a39464a,a39467a,a39470a,a39471a,a39472a,a39476a,a39477a,a39481a,a39482a,a39483a,a39487a,a39488a,a39491a,a39494a,a39495a,a39496a,a39500a,a39501a,a39505a,a39506a,a39507a,a39511a,a39512a,a39515a,a39518a,a39519a,a39520a,a39524a,a39525a,a39529a,a39530a,a39531a,a39535a,a39536a,a39539a,a39542a,a39543a,a39544a,a39548a,a39549a,a39553a,a39554a,a39555a,a39559a,a39560a,a39563a,a39566a,a39567a,a39568a,a39572a,a39573a,a39577a,a39578a,a39579a,a39583a,a39584a,a39587a,a39590a,a39591a,a39592a,a39596a,a39597a,a39601a,a39602a,a39603a,a39607a,a39608a,a39611a,a39614a,a39615a,a39616a,a39620a,a39621a,a39625a,a39626a,a39627a,a39631a,a39632a,a39635a,a39638a,a39639a,a39640a,a39644a,a39645a,a39649a,a39650a,a39651a,a39655a,a39656a,a39659a,a39662a,a39663a,a39664a,a39668a,a39669a,a39673a,a39674a,a39675a,a39679a,a39680a,a39683a,a39686a,a39687a,a39688a,a39692a,a39693a,a39697a,a39698a,a39699a,a39703a,a39704a,a39707a,a39710a,a39711a,a39712a,a39716a,a39717a,a39721a,a39722a,a39723a,a39727a,a39728a,a39731a,a39734a,a39735a,a39736a,a39740a,a39741a,a39745a,a39746a,a39747a,a39751a,a39752a,a39755a,a39758a,a39759a,a39760a,a39764a,a39765a,a39769a,a39770a,a39771a,a39775a,a39776a,a39779a,a39782a,a39783a,a39784a,a39788a,a39789a,a39793a,a39794a,a39795a,a39799a,a39800a,a39803a,a39806a,a39807a,a39808a,a39812a,a39813a,a39817a,a39818a,a39819a,a39823a,a39824a,a39827a,a39830a,a39831a,a39832a,a39836a,a39837a,a39841a,a39842a,a39843a,a39847a,a39848a,a39851a,a39854a,a39855a,a39856a,a39860a,a39861a,a39865a,a39866a,a39867a,a39871a,a39872a,a39875a,a39878a,a39879a,a39880a,a39884a,a39885a,a39889a,a39890a,a39891a,a39895a,a39896a,a39899a,a39902a,a39903a,a39904a,a39908a,a39909a,a39913a,a39914a,a39915a,a39919a,a39920a,a39923a,a39926a,a39927a,a39928a,a39932a,a39933a,a39937a,a39938a,a39939a,a39943a,a39944a,a39947a,a39950a,a39951a,a39952a,a39956a,a39957a,a39961a,a39962a,a39963a,a39967a,a39968a,a39971a,a39974a,a39975a,a39976a,a39980a,a39981a,a39985a,a39986a,a39987a,a39991a,a39992a,a39995a,a39998a,a39999a,a40000a,a40004a,a40005a,a40009a,a40010a,a40011a,a40015a,a40016a,a40019a,a40022a,a40023a,a40024a,a40028a,a40029a,a40033a,a40034a,a40035a,a40039a,a40040a,a40043a,a40046a,a40047a,a40048a,a40052a,a40053a,a40057a,a40058a,a40059a,a40063a,a40064a,a40067a,a40070a,a40071a,a40072a,a40076a,a40077a,a40081a,a40082a,a40083a,a40087a,a40088a,a40091a,a40094a,a40095a,a40096a,a40100a,a40101a,a40105a,a40106a,a40107a,a40111a,a40112a,a40115a,a40118a,a40119a,a40120a,a40124a,a40125a,a40129a,a40130a,a40131a,a40135a,a40136a,a40139a,a40142a,a40143a,a40144a,a40148a,a40149a,a40153a,a40154a,a40155a,a40159a,a40160a,a40163a,a40166a,a40167a,a40168a,a40172a,a40173a,a40177a,a40178a,a40179a,a40183a,a40184a,a40187a,a40190a,a40191a,a40192a,a40196a,a40197a,a40201a,a40202a,a40203a,a40207a,a40208a,a40211a,a40214a,a40215a,a40216a,a40220a,a40221a,a40225a,a40226a,a40227a,a40231a,a40232a,a40235a,a40238a,a40239a,a40240a,a40244a,a40245a,a40249a,a40250a,a40251a,a40255a,a40256a,a40259a,a40262a,a40263a,a40264a,a40268a,a40269a,a40273a,a40274a,a40275a,a40279a,a40280a,a40283a,a40286a,a40287a,a40288a,a40292a,a40293a,a40297a,a40298a,a40299a,a40303a,a40304a,a40307a,a40310a,a40311a,a40312a,a40316a,a40317a,a40321a,a40322a,a40323a,a40327a,a40328a,a40331a,a40334a,a40335a,a40336a,a40340a,a40341a,a40345a,a40346a,a40347a,a40351a,a40352a,a40355a,a40358a,a40359a,a40360a,a40364a,a40365a,a40369a,a40370a,a40371a,a40375a,a40376a,a40379a,a40382a,a40383a,a40384a,a40388a,a40389a,a40393a,a40394a,a40395a,a40399a,a40400a,a40403a,a40406a,a40407a,a40408a,a40412a,a40413a,a40417a,a40418a,a40419a,a40423a,a40424a,a40427a,a40430a,a40431a,a40432a,a40436a,a40437a,a40441a,a40442a,a40443a,a40447a,a40448a,a40451a,a40454a,a40455a,a40456a,a40460a,a40461a,a40465a,a40466a,a40467a,a40471a,a40472a,a40475a,a40478a,a40479a,a40480a,a40484a,a40485a,a40489a,a40490a,a40491a,a40495a,a40496a,a40499a,a40502a,a40503a,a40504a,a40508a,a40509a,a40513a,a40514a,a40515a,a40519a,a40520a,a40523a,a40526a,a40527a,a40528a,a40532a,a40533a,a40537a,a40538a,a40539a,a40543a,a40544a,a40547a,a40550a,a40551a,a40552a,a40556a,a40557a,a40561a,a40562a,a40563a,a40567a,a40568a,a40571a,a40574a,a40575a,a40576a,a40580a,a40581a,a40585a,a40586a,a40587a,a40591a,a40592a,a40595a,a40598a,a40599a,a40600a,a40604a,a40605a,a40609a,a40610a,a40611a,a40615a,a40616a,a40619a,a40622a,a40623a,a40624a,a40628a,a40629a,a40633a,a40634a,a40635a,a40639a,a40640a,a40643a,a40646a,a40647a,a40648a,a40652a,a40653a,a40657a,a40658a,a40659a,a40663a,a40664a,a40667a,a40670a,a40671a,a40672a,a40676a,a40677a,a40681a,a40682a,a40683a,a40687a,a40688a,a40691a,a40694a,a40695a,a40696a,a40700a,a40701a,a40705a,a40706a,a40707a,a40711a,a40712a,a40715a,a40718a,a40719a,a40720a,a40724a,a40725a,a40729a,a40730a,a40731a,a40735a,a40736a,a40739a,a40742a,a40743a,a40744a,a40748a,a40749a,a40753a,a40754a,a40755a,a40759a,a40760a,a40763a,a40766a,a40767a,a40768a,a40772a,a40773a,a40777a,a40778a,a40779a,a40783a,a40784a,a40787a,a40790a,a40791a,a40792a,a40796a,a40797a,a40801a,a40802a,a40803a,a40807a,a40808a,a40811a,a40814a,a40815a,a40816a,a40820a,a40821a,a40825a,a40826a,a40827a,a40831a,a40832a,a40835a,a40838a,a40839a,a40840a,a40844a,a40845a,a40849a,a40850a,a40851a,a40855a,a40856a,a40859a,a40862a,a40863a,a40864a,a40868a,a40869a,a40873a,a40874a,a40875a,a40879a,a40880a,a40883a,a40886a,a40887a,a40888a,a40892a,a40893a,a40897a,a40898a,a40899a,a40903a,a40904a,a40907a,a40910a,a40911a,a40912a,a40916a,a40917a,a40921a,a40922a,a40923a,a40927a,a40928a,a40931a,a40934a,a40935a,a40936a,a40940a,a40941a,a40945a,a40946a,a40947a,a40951a,a40952a,a40955a,a40958a,a40959a,a40960a,a40964a,a40965a,a40969a,a40970a,a40971a,a40975a,a40976a,a40979a,a40982a,a40983a,a40984a,a40988a,a40989a,a40993a,a40994a,a40995a,a40999a,a41000a,a41003a,a41006a,a41007a,a41008a,a41012a,a41013a,a41017a,a41018a,a41019a,a41023a,a41024a,a41027a,a41030a,a41031a,a41032a,a41036a,a41037a,a41041a,a41042a,a41043a,a41047a,a41048a,a41051a,a41054a,a41055a,a41056a,a41060a,a41061a,a41065a,a41066a,a41067a,a41071a,a41072a,a41075a,a41078a,a41079a,a41080a,a41084a,a41085a,a41089a,a41090a,a41091a,a41095a,a41096a,a41099a,a41102a,a41103a,a41104a,a41108a,a41109a,a41113a,a41114a,a41115a,a41119a,a41120a,a41123a,a41126a,a41127a,a41128a,a41132a,a41133a,a41137a,a41138a,a41139a,a41143a,a41144a,a41147a,a41150a,a41151a,a41152a,a41156a,a41157a,a41161a,a41162a,a41163a,a41167a,a41168a,a41171a,a41174a,a41175a,a41176a,a41180a,a41181a,a41185a,a41186a,a41187a,a41191a,a41192a,a41195a,a41198a,a41199a,a41200a,a41204a,a41205a,a41209a,a41210a,a41211a,a41215a,a41216a,a41219a,a41222a,a41223a,a41224a,a41228a,a41229a,a41233a,a41234a,a41235a,a41239a,a41240a,a41243a,a41246a,a41247a,a41248a,a41252a,a41253a,a41257a,a41258a,a41259a,a41263a,a41264a,a41267a,a41270a,a41271a,a41272a,a41276a,a41277a,a41281a,a41282a,a41283a,a41287a,a41288a,a41291a,a41294a,a41295a,a41296a,a41300a,a41301a,a41305a,a41306a,a41307a,a41311a,a41312a,a41315a,a41318a,a41319a,a41320a,a41324a,a41325a,a41329a,a41330a,a41331a,a41335a,a41336a,a41339a,a41342a,a41343a,a41344a,a41348a,a41349a,a41353a,a41354a,a41355a,a41359a,a41360a,a41363a,a41366a,a41367a,a41368a,a41372a,a41373a,a41377a,a41378a,a41379a,a41383a,a41384a,a41387a,a41390a,a41391a,a41392a,a41396a,a41397a,a41401a,a41402a,a41403a,a41407a,a41408a,a41411a,a41414a,a41415a,a41416a,a41420a,a41421a,a41425a,a41426a,a41427a,a41431a,a41432a,a41435a,a41438a,a41439a,a41440a,a41444a,a41445a,a41449a,a41450a,a41451a,a41455a,a41456a,a41459a,a41462a,a41463a,a41464a,a41468a,a41469a,a41473a,a41474a,a41475a,a41479a,a41480a,a41483a,a41486a,a41487a,a41488a,a41492a,a41493a,a41497a,a41498a,a41499a,a41503a,a41504a,a41507a,a41510a,a41511a,a41512a,a41516a,a41517a,a41521a,a41522a,a41523a,a41527a,a41528a,a41531a,a41534a,a41535a,a41536a,a41540a,a41541a,a41545a,a41546a,a41547a,a41551a,a41552a,a41555a,a41558a,a41559a,a41560a,a41564a,a41565a,a41569a,a41570a,a41571a,a41575a,a41576a,a41579a,a41582a,a41583a,a41584a,a41588a,a41589a,a41593a,a41594a,a41595a,a41599a,a41600a,a41603a,a41606a,a41607a,a41608a,a41612a,a41613a,a41617a,a41618a,a41619a,a41623a,a41624a,a41627a,a41630a,a41631a,a41632a,a41636a,a41637a,a41641a,a41642a,a41643a,a41647a,a41648a,a41651a,a41654a,a41655a,a41656a,a41660a,a41661a,a41665a,a41666a,a41667a,a41671a,a41672a,a41675a,a41678a,a41679a,a41680a,a41684a,a41685a,a41689a,a41690a,a41691a,a41695a,a41696a,a41699a,a41702a,a41703a,a41704a,a41708a,a41709a,a41713a,a41714a,a41715a,a41719a,a41720a,a41723a,a41726a,a41727a,a41728a,a41732a,a41733a,a41737a,a41738a,a41739a,a41743a,a41744a,a41747a,a41750a,a41751a,a41752a,a41756a,a41757a,a41761a,a41762a,a41763a,a41767a,a41768a,a41771a,a41774a,a41775a,a41776a,a41780a,a41781a,a41785a,a41786a,a41787a,a41791a,a41792a,a41795a,a41798a,a41799a,a41800a,a41804a,a41805a,a41809a,a41810a,a41811a,a41815a,a41816a,a41819a,a41822a,a41823a,a41824a,a41828a,a41829a,a41833a,a41834a,a41835a,a41839a,a41840a,a41843a,a41846a,a41847a,a41848a,a41852a,a41853a,a41857a,a41858a,a41859a,a41863a,a41864a,a41867a,a41870a,a41871a,a41872a,a41876a,a41877a,a41881a,a41882a,a41883a,a41887a,a41888a,a41891a,a41894a,a41895a,a41896a,a41900a,a41901a,a41905a,a41906a,a41907a,a41911a,a41912a,a41915a,a41918a,a41919a,a41920a,a41924a,a41925a,a41929a,a41930a,a41931a,a41935a,a41936a,a41939a,a41942a,a41943a,a41944a,a41948a,a41949a,a41953a,a41954a,a41955a,a41959a,a41960a,a41963a,a41966a,a41967a,a41968a,a41972a,a41973a,a41977a,a41978a,a41979a,a41983a,a41984a,a41987a,a41990a,a41991a,a41992a,a41996a,a41997a,a42001a,a42002a,a42003a,a42007a,a42008a,a42011a,a42014a,a42015a,a42016a,a42020a,a42021a,a42025a,a42026a,a42027a,a42031a,a42032a,a42035a,a42038a,a42039a,a42040a,a42044a,a42045a,a42049a,a42050a,a42051a,a42055a,a42056a,a42059a,a42062a,a42063a,a42064a,a42068a,a42069a,a42073a,a42074a,a42075a,a42079a,a42080a,a42083a,a42086a,a42087a,a42088a,a42092a,a42093a,a42097a,a42098a,a42099a,a42103a,a42104a,a42107a,a42110a,a42111a,a42112a,a42116a,a42117a,a42121a,a42122a,a42123a,a42127a,a42128a,a42131a,a42134a,a42135a,a42136a,a42140a,a42141a,a42145a,a42146a,a42147a,a42151a,a42152a,a42155a,a42158a,a42159a,a42160a,a42164a,a42165a,a42169a,a42170a,a42171a,a42175a,a42176a,a42179a,a42182a,a42183a,a42184a,a42188a,a42189a,a42193a,a42194a,a42195a,a42199a,a42200a,a42203a,a42206a,a42207a,a42208a,a42212a,a42213a,a42217a,a42218a,a42219a,a42223a,a42224a,a42227a,a42230a,a42231a,a42232a,a42236a,a42237a,a42241a,a42242a,a42243a,a42247a,a42248a,a42251a,a42254a,a42255a,a42256a,a42260a,a42261a,a42265a,a42266a,a42267a,a42271a,a42272a,a42275a,a42278a,a42279a,a42280a,a42284a,a42285a,a42289a,a42290a,a42291a,a42295a,a42296a,a42299a,a42302a,a42303a,a42304a,a42308a,a42309a,a42313a,a42314a,a42315a,a42319a,a42320a,a42323a,a42326a,a42327a,a42328a,a42332a,a42333a,a42337a,a42338a,a42339a,a42343a,a42344a,a42347a,a42350a,a42351a,a42352a,a42356a,a42357a,a42361a,a42362a,a42363a,a42367a,a42368a,a42371a,a42374a,a42375a,a42376a,a42380a,a42381a,a42385a,a42386a,a42387a,a42391a,a42392a,a42395a,a42398a,a42399a,a42400a,a42404a,a42405a,a42409a,a42410a,a42411a,a42415a,a42416a,a42419a,a42422a,a42423a,a42424a,a42428a,a42429a,a42433a,a42434a,a42435a,a42439a,a42440a,a42443a,a42446a,a42447a,a42448a,a42452a,a42453a,a42457a,a42458a,a42459a,a42463a,a42464a,a42467a,a42470a,a42471a,a42472a,a42476a,a42477a,a42481a,a42482a,a42483a,a42487a,a42488a,a42491a,a42494a,a42495a,a42496a,a42500a,a42501a,a42505a,a42506a,a42507a,a42511a,a42512a,a42515a,a42518a,a42519a,a42520a,a42524a,a42525a,a42529a,a42530a,a42531a,a42535a,a42536a,a42539a,a42542a,a42543a,a42544a,a42548a,a42549a,a42553a,a42554a,a42555a,a42559a,a42560a,a42563a,a42566a,a42567a,a42568a,a42572a,a42573a,a42577a,a42578a,a42579a,a42583a,a42584a,a42587a,a42590a,a42591a,a42592a,a42596a,a42597a,a42601a,a42602a,a42603a,a42607a,a42608a,a42611a,a42614a,a42615a,a42616a,a42620a,a42621a,a42625a,a42626a,a42627a,a42631a,a42632a,a42635a,a42638a,a42639a,a42640a,a42644a,a42645a,a42649a,a42650a,a42651a,a42655a,a42656a,a42659a,a42662a,a42663a,a42664a,a42668a,a42669a,a42673a,a42674a,a42675a,a42679a,a42680a,a42683a,a42686a,a42687a,a42688a,a42692a,a42693a,a42697a,a42698a,a42699a,a42703a,a42704a,a42707a,a42710a,a42711a,a42712a,a42716a,a42717a,a42721a,a42722a,a42723a,a42727a,a42728a,a42731a,a42734a,a42735a,a42736a,a42740a,a42741a,a42745a,a42746a,a42747a,a42751a,a42752a,a42755a,a42758a,a42759a,a42760a,a42764a,a42765a,a42769a,a42770a,a42771a,a42775a,a42776a,a42779a,a42782a,a42783a,a42784a,a42788a,a42789a,a42793a,a42794a,a42795a,a42799a,a42800a,a42803a,a42806a,a42807a,a42808a,a42812a,a42813a,a42817a,a42818a,a42819a,a42823a,a42824a,a42827a,a42830a,a42831a,a42832a,a42836a,a42837a,a42841a,a42842a,a42843a,a42847a,a42848a,a42851a,a42854a,a42855a,a42856a,a42860a,a42861a,a42865a,a42866a,a42867a,a42871a,a42872a,a42875a,a42878a,a42879a,a42880a,a42884a,a42885a,a42889a,a42890a,a42891a,a42895a,a42896a,a42899a,a42902a,a42903a,a42904a,a42908a,a42909a,a42913a,a42914a,a42915a,a42919a,a42920a,a42923a,a42926a,a42927a,a42928a,a42932a,a42933a,a42937a,a42938a,a42939a,a42943a,a42944a,a42947a,a42950a,a42951a,a42952a,a42956a,a42957a,a42961a,a42962a,a42963a,a42967a,a42968a,a42971a,a42974a,a42975a,a42976a,a42980a,a42981a,a42985a,a42986a,a42987a,a42991a,a42992a,a42995a,a42998a,a42999a,a43000a,a43004a,a43005a,a43009a,a43010a,a43011a,a43015a,a43016a,a43019a,a43022a,a43023a,a43024a,a43028a,a43029a,a43033a,a43034a,a43035a,a43039a,a43040a,a43043a,a43046a,a43047a,a43048a,a43052a,a43053a,a43057a,a43058a,a43059a,a43063a,a43064a,a43067a,a43070a,a43071a,a43072a,a43076a,a43077a,a43081a,a43082a,a43083a,a43087a,a43088a,a43091a,a43094a,a43095a,a43096a,a43100a,a43101a,a43105a,a43106a,a43107a,a43111a,a43112a,a43115a,a43118a,a43119a,a43120a,a43124a,a43125a,a43129a,a43130a,a43131a,a43135a,a43136a,a43139a,a43142a,a43143a,a43144a,a43148a,a43149a,a43153a,a43154a,a43155a,a43159a,a43160a,a43163a,a43166a,a43167a,a43168a,a43172a,a43173a,a43177a,a43178a,a43179a,a43183a,a43184a,a43187a,a43190a,a43191a,a43192a,a43196a,a43197a,a43201a,a43202a,a43203a,a43207a,a43208a,a43211a,a43214a,a43215a,a43216a,a43220a,a43221a,a43225a,a43226a,a43227a,a43231a,a43232a,a43235a,a43238a,a43239a,a43240a,a43244a,a43245a,a43249a,a43250a,a43251a,a43255a,a43256a,a43259a,a43262a,a43263a,a43264a,a43268a,a43269a,a43273a,a43274a,a43275a,a43279a,a43280a,a43283a,a43286a,a43287a,a43288a,a43292a,a43293a,a43297a,a43298a,a43299a,a43303a,a43304a,a43307a,a43310a,a43311a,a43312a,a43316a,a43317a,a43321a,a43322a,a43323a,a43327a,a43328a,a43331a,a43334a,a43335a,a43336a,a43340a,a43341a,a43345a,a43346a,a43347a,a43351a,a43352a,a43355a,a43358a,a43359a,a43360a,a43364a,a43365a,a43369a,a43370a,a43371a,a43375a,a43376a,a43379a,a43382a,a43383a,a43384a,a43388a,a43389a,a43393a,a43394a,a43395a,a43399a,a43400a,a43403a,a43406a,a43407a,a43408a,a43412a,a43413a,a43417a,a43418a,a43419a,a43423a,a43424a,a43427a,a43430a,a43431a,a43432a,a43436a,a43437a,a43441a,a43442a,a43443a,a43447a,a43448a,a43451a,a43454a,a43455a,a43456a,a43460a,a43461a,a43465a,a43466a,a43467a,a43471a,a43472a,a43475a,a43478a,a43479a,a43480a,a43484a,a43485a,a43489a,a43490a,a43491a,a43495a,a43496a,a43499a,a43502a,a43503a,a43504a,a43508a,a43509a,a43513a,a43514a,a43515a,a43519a,a43520a,a43523a,a43526a,a43527a,a43528a,a43532a,a43533a,a43537a,a43538a,a43539a,a43543a,a43544a,a43547a,a43550a,a43551a,a43552a,a43556a,a43557a,a43561a,a43562a,a43563a,a43567a,a43568a,a43571a,a43574a,a43575a,a43576a,a43580a,a43581a,a43585a,a43586a,a43587a,a43591a,a43592a,a43595a,a43598a,a43599a,a43600a,a43604a,a43605a,a43609a,a43610a,a43611a,a43615a,a43616a,a43619a,a43622a,a43623a,a43624a,a43628a,a43629a,a43633a,a43634a,a43635a,a43639a,a43640a,a43643a,a43646a,a43647a,a43648a,a43652a,a43653a,a43657a,a43658a,a43659a,a43663a,a43664a,a43667a,a43670a,a43671a,a43672a,a43676a,a43677a,a43681a,a43682a,a43683a,a43687a,a43688a,a43691a,a43694a,a43695a,a43696a,a43700a,a43701a,a43705a,a43706a,a43707a,a43711a,a43712a,a43715a,a43718a,a43719a,a43720a,a43724a,a43725a,a43729a,a43730a,a43731a,a43735a,a43736a,a43739a,a43742a,a43743a,a43744a,a43748a,a43749a,a43753a,a43754a,a43755a,a43759a,a43760a,a43763a,a43766a,a43767a,a43768a,a43772a,a43773a,a43777a,a43778a,a43779a,a43783a,a43784a,a43787a,a43790a,a43791a,a43792a,a43796a,a43797a,a43801a,a43802a,a43803a,a43807a,a43808a,a43811a,a43814a,a43815a,a43816a,a43820a,a43821a,a43825a,a43826a,a43827a,a43831a,a43832a,a43835a,a43838a,a43839a,a43840a,a43844a,a43845a,a43849a,a43850a,a43851a,a43855a,a43856a,a43859a,a43862a,a43863a,a43864a,a43868a,a43869a,a43873a,a43874a,a43875a,a43879a,a43880a,a43883a,a43886a,a43887a,a43888a,a43892a,a43893a,a43897a,a43898a,a43899a,a43903a,a43904a,a43907a,a43910a,a43911a,a43912a,a43916a,a43917a,a43921a,a43922a,a43923a,a43927a,a43928a,a43931a,a43934a,a43935a,a43936a,a43940a,a43941a,a43945a,a43946a,a43947a,a43951a,a43952a,a43955a,a43958a,a43959a,a43960a,a43964a,a43965a,a43969a,a43970a,a43971a,a43975a,a43976a,a43979a,a43982a,a43983a,a43984a,a43988a,a43989a,a43993a,a43994a,a43995a,a43999a,a44000a,a44003a,a44006a,a44007a,a44008a,a44012a,a44013a,a44017a,a44018a,a44019a,a44023a,a44024a,a44027a,a44030a,a44031a,a44032a,a44036a,a44037a,a44041a,a44042a,a44043a,a44047a,a44048a,a44051a,a44054a,a44055a,a44056a,a44060a,a44061a,a44065a,a44066a,a44067a,a44071a,a44072a,a44075a,a44078a,a44079a,a44080a,a44084a,a44085a,a44089a,a44090a,a44091a,a44095a,a44096a,a44099a,a44102a,a44103a,a44104a,a44108a,a44109a,a44113a,a44114a,a44115a,a44119a,a44120a,a44123a,a44126a,a44127a,a44128a,a44132a,a44133a,a44137a,a44138a,a44139a,a44143a,a44144a,a44147a,a44150a,a44151a,a44152a,a44156a,a44157a,a44161a,a44162a,a44163a,a44167a,a44168a,a44171a,a44174a,a44175a,a44176a,a44180a,a44181a,a44185a,a44186a,a44187a,a44191a,a44192a,a44195a,a44198a,a44199a,a44200a,a44204a,a44205a,a44209a,a44210a,a44211a,a44215a,a44216a,a44219a,a44222a,a44223a,a44224a,a44228a,a44229a,a44233a,a44234a,a44235a,a44239a,a44240a,a44243a,a44246a,a44247a,a44248a,a44252a,a44253a,a44257a,a44258a,a44259a,a44263a,a44264a,a44267a,a44270a,a44271a,a44272a,a44276a,a44277a,a44281a,a44282a,a44283a,a44287a,a44288a,a44291a,a44294a,a44295a,a44296a,a44300a,a44301a,a44305a,a44306a,a44307a,a44311a,a44312a,a44315a,a44318a,a44319a,a44320a,a44324a,a44325a,a44329a,a44330a,a44331a,a44335a,a44336a,a44339a,a44342a,a44343a,a44344a,a44348a,a44349a,a44353a,a44354a,a44355a,a44359a,a44360a,a44363a,a44366a,a44367a,a44368a,a44372a,a44373a,a44377a,a44378a,a44379a,a44383a,a44384a,a44387a,a44390a,a44391a,a44392a,a44396a,a44397a,a44401a,a44402a,a44403a,a44407a,a44408a,a44411a,a44414a,a44415a,a44416a,a44420a,a44421a,a44425a,a44426a,a44427a,a44431a,a44432a,a44435a,a44438a,a44439a,a44440a,a44444a,a44445a,a44449a,a44450a,a44451a,a44455a,a44456a,a44459a,a44462a,a44463a,a44464a,a44468a,a44469a,a44473a,a44474a,a44475a,a44479a,a44480a,a44483a,a44486a,a44487a,a44488a,a44492a,a44493a,a44497a,a44498a,a44499a,a44503a,a44504a,a44507a,a44510a,a44511a,a44512a,a44516a,a44517a,a44521a,a44522a,a44523a,a44527a,a44528a,a44531a,a44534a,a44535a,a44536a,a44540a,a44541a,a44545a,a44546a,a44547a,a44551a,a44552a,a44555a,a44558a,a44559a,a44560a,a44564a,a44565a,a44569a,a44570a,a44571a,a44575a,a44576a,a44579a,a44582a,a44583a,a44584a,a44588a,a44589a,a44593a,a44594a,a44595a,a44599a,a44600a,a44603a,a44606a,a44607a,a44608a,a44612a,a44613a,a44617a,a44618a,a44619a,a44623a,a44624a,a44627a,a44630a,a44631a,a44632a,a44636a,a44637a,a44641a,a44642a,a44643a,a44647a,a44648a,a44651a,a44654a,a44655a,a44656a,a44660a,a44661a,a44665a,a44666a,a44667a,a44671a,a44672a,a44675a,a44678a,a44679a,a44680a,a44684a,a44685a,a44689a,a44690a,a44691a,a44695a,a44696a,a44699a,a44702a,a44703a,a44704a,a44708a,a44709a,a44713a,a44714a,a44715a,a44719a,a44720a,a44723a,a44726a,a44727a,a44728a,a44732a,a44733a,a44737a,a44738a,a44739a,a44743a,a44744a,a44747a,a44750a,a44751a,a44752a,a44756a,a44757a,a44761a,a44762a,a44763a,a44767a,a44768a,a44771a,a44774a,a44775a,a44776a,a44780a,a44781a,a44785a,a44786a,a44787a,a44791a,a44792a,a44795a,a44798a,a44799a,a44800a,a44804a,a44805a,a44809a,a44810a,a44811a,a44815a,a44816a,a44819a,a44822a,a44823a,a44824a,a44828a,a44829a,a44833a,a44834a,a44835a,a44839a,a44840a,a44843a,a44846a,a44847a,a44848a,a44852a,a44853a,a44857a,a44858a,a44859a,a44863a,a44864a,a44867a,a44870a,a44871a,a44872a,a44876a,a44877a,a44881a,a44882a,a44883a,a44887a,a44888a,a44891a,a44894a,a44895a,a44896a,a44900a,a44901a,a44905a,a44906a,a44907a,a44911a,a44912a,a44915a,a44918a,a44919a,a44920a,a44924a,a44925a,a44929a,a44930a,a44931a,a44935a,a44936a,a44939a,a44942a,a44943a,a44944a,a44948a,a44949a,a44953a,a44954a,a44955a,a44959a,a44960a,a44963a,a44966a,a44967a,a44968a,a44972a,a44973a,a44977a,a44978a,a44979a,a44983a,a44984a,a44987a,a44990a,a44991a,a44992a,a44996a,a44997a,a45001a,a45002a,a45003a,a45007a,a45008a,a45011a,a45014a,a45015a,a45016a,a45020a,a45021a,a45025a,a45026a,a45027a,a45031a,a45032a,a45035a,a45038a,a45039a,a45040a,a45044a,a45045a,a45049a,a45050a,a45051a,a45055a,a45056a,a45059a,a45062a,a45063a,a45064a,a45068a,a45069a,a45073a,a45074a,a45075a,a45079a,a45080a,a45083a,a45086a,a45087a,a45088a,a45092a,a45093a,a45097a,a45098a,a45099a,a45103a,a45104a,a45107a,a45110a,a45111a,a45112a,a45116a,a45117a,a45121a,a45122a,a45123a,a45127a,a45128a,a45131a,a45134a,a45135a,a45136a,a45140a,a45141a,a45145a,a45146a,a45147a,a45151a,a45152a,a45155a,a45158a,a45159a,a45160a,a45164a,a45165a,a45169a,a45170a,a45171a,a45175a,a45176a,a45179a,a45182a,a45183a,a45184a,a45188a,a45189a,a45193a,a45194a,a45195a,a45199a,a45200a,a45203a,a45206a,a45207a,a45208a,a45212a,a45213a,a45217a,a45218a,a45219a,a45223a,a45224a,a45227a,a45230a,a45231a,a45232a,a45236a,a45237a,a45241a,a45242a,a45243a,a45247a,a45248a,a45251a,a45254a,a45255a,a45256a,a45260a,a45261a,a45265a,a45266a,a45267a,a45271a,a45272a,a45275a,a45278a,a45279a,a45280a,a45284a,a45285a,a45289a,a45290a,a45291a,a45295a,a45296a,a45299a,a45302a,a45303a,a45304a,a45308a,a45309a,a45313a,a45314a,a45315a,a45319a,a45320a,a45323a,a45326a,a45327a,a45328a,a45332a,a45333a,a45337a,a45338a,a45339a,a45343a,a45344a,a45347a,a45350a,a45351a,a45352a,a45356a,a45357a,a45361a,a45362a,a45363a,a45367a,a45368a,a45371a,a45374a,a45375a,a45376a,a45380a,a45381a,a45385a,a45386a,a45387a,a45391a,a45392a,a45395a,a45398a,a45399a,a45400a,a45404a,a45405a,a45409a,a45410a,a45411a,a45415a,a45416a,a45419a,a45422a,a45423a,a45424a,a45428a,a45429a,a45433a,a45434a,a45435a,a45439a,a45440a,a45443a,a45446a,a45447a,a45448a,a45452a,a45453a,a45457a,a45458a,a45459a,a45463a,a45464a,a45467a,a45470a,a45471a,a45472a,a45476a,a45477a,a45481a,a45482a,a45483a,a45487a,a45488a,a45491a,a45494a,a45495a,a45496a,a45500a,a45501a,a45505a,a45506a,a45507a,a45511a,a45512a,a45515a,a45518a,a45519a,a45520a,a45524a,a45525a,a45529a,a45530a,a45531a,a45535a,a45536a,a45539a,a45542a,a45543a,a45544a,a45548a,a45549a,a45553a,a45554a,a45555a,a45559a,a45560a,a45563a,a45566a,a45567a,a45568a,a45572a,a45573a,a45577a,a45578a,a45579a,a45583a,a45584a,a45587a,a45590a,a45591a,a45592a,a45596a,a45597a,a45601a,a45602a,a45603a,a45607a,a45608a,a45611a,a45614a,a45615a,a45616a,a45620a,a45621a,a45625a,a45626a,a45627a,a45631a,a45632a,a45635a,a45638a,a45639a,a45640a,a45644a,a45645a,a45649a,a45650a,a45651a,a45655a,a45656a,a45659a,a45662a,a45663a,a45664a,a45668a,a45669a,a45673a,a45674a,a45675a,a45679a,a45680a,a45683a,a45686a,a45687a,a45688a,a45692a,a45693a,a45697a,a45698a,a45699a,a45703a,a45704a,a45707a,a45710a,a45711a,a45712a,a45716a,a45717a,a45721a,a45722a,a45723a,a45727a,a45728a,a45731a,a45734a,a45735a,a45736a,a45740a,a45741a,a45745a,a45746a,a45747a,a45751a,a45752a,a45755a,a45758a,a45759a,a45760a,a45764a,a45765a,a45769a,a45770a,a45771a,a45775a,a45776a,a45779a,a45782a,a45783a,a45784a,a45788a,a45789a,a45793a,a45794a,a45795a,a45799a,a45800a,a45803a,a45806a,a45807a,a45808a,a45812a,a45813a,a45817a,a45818a,a45819a,a45823a,a45824a,a45827a,a45830a,a45831a,a45832a,a45836a,a45837a,a45841a,a45842a,a45843a,a45847a,a45848a,a45851a,a45854a,a45855a,a45856a,a45860a,a45861a,a45865a,a45866a,a45867a,a45871a,a45872a,a45875a,a45878a,a45879a,a45880a,a45884a,a45885a,a45889a,a45890a,a45891a,a45895a,a45896a,a45899a,a45902a,a45903a,a45904a,a45908a,a45909a,a45913a,a45914a,a45915a,a45919a,a45920a,a45923a,a45926a,a45927a,a45928a,a45932a,a45933a,a45937a,a45938a,a45939a,a45943a,a45944a,a45947a,a45950a,a45951a,a45952a,a45956a,a45957a,a45961a,a45962a,a45963a,a45967a,a45968a,a45971a,a45974a,a45975a,a45976a,a45980a,a45981a,a45985a,a45986a,a45987a,a45991a,a45992a,a45995a,a45998a,a45999a,a46000a,a46004a,a46005a,a46009a,a46010a,a46011a,a46015a,a46016a,a46019a,a46022a,a46023a,a46024a,a46028a,a46029a,a46033a,a46034a,a46035a,a46039a,a46040a,a46043a,a46046a,a46047a,a46048a,a46052a,a46053a,a46057a,a46058a,a46059a,a46063a,a46064a,a46067a,a46070a,a46071a,a46072a,a46076a,a46077a,a46081a,a46082a,a46083a,a46087a,a46088a,a46091a,a46094a,a46095a,a46096a,a46100a,a46101a,a46105a,a46106a,a46107a,a46111a,a46112a,a46115a,a46118a,a46119a,a46120a,a46124a,a46125a,a46129a,a46130a,a46131a,a46135a,a46136a,a46139a,a46142a,a46143a,a46144a,a46148a,a46149a,a46153a,a46154a,a46155a,a46159a,a46160a,a46163a,a46166a,a46167a,a46168a,a46172a,a46173a,a46177a,a46178a,a46179a,a46183a,a46184a,a46187a,a46190a,a46191a,a46192a,a46196a,a46197a,a46201a,a46202a,a46203a,a46207a,a46208a,a46211a,a46214a,a46215a,a46216a,a46220a,a46221a,a46225a,a46226a,a46227a,a46231a,a46232a,a46235a,a46238a,a46239a,a46240a,a46244a,a46245a,a46249a,a46250a,a46251a,a46255a,a46256a,a46259a,a46262a,a46263a,a46264a,a46268a,a46269a,a46273a,a46274a,a46275a,a46279a,a46280a,a46283a,a46286a,a46287a,a46288a,a46292a,a46293a,a46297a,a46298a,a46299a,a46303a,a46304a,a46307a,a46310a,a46311a,a46312a,a46316a,a46317a,a46321a,a46322a,a46323a,a46327a,a46328a,a46331a,a46334a,a46335a,a46336a,a46340a,a46341a,a46345a,a46346a,a46347a,a46351a,a46352a,a46355a,a46358a,a46359a,a46360a,a46364a,a46365a,a46369a,a46370a,a46371a,a46375a,a46376a,a46379a,a46382a,a46383a,a46384a,a46388a,a46389a,a46393a,a46394a,a46395a,a46399a,a46400a,a46403a,a46406a,a46407a,a46408a,a46412a,a46413a,a46417a,a46418a,a46419a,a46423a,a46424a,a46427a,a46430a,a46431a,a46432a,a46436a,a46437a,a46441a,a46442a,a46443a,a46447a,a46448a,a46451a,a46454a,a46455a,a46456a,a46460a,a46461a,a46465a,a46466a,a46467a,a46471a,a46472a,a46475a,a46478a,a46479a,a46480a,a46484a,a46485a,a46489a,a46490a,a46491a,a46495a,a46496a,a46499a,a46502a,a46503a,a46504a,a46508a,a46509a,a46513a,a46514a,a46515a,a46519a,a46520a,a46523a,a46526a,a46527a,a46528a,a46532a,a46533a,a46537a,a46538a,a46539a,a46543a,a46544a,a46547a,a46550a,a46551a,a46552a,a46556a,a46557a,a46561a,a46562a,a46563a,a46567a,a46568a,a46571a,a46574a,a46575a,a46576a,a46580a,a46581a,a46585a,a46586a,a46587a,a46591a,a46592a,a46595a,a46598a,a46599a,a46600a,a46604a,a46605a,a46609a,a46610a,a46611a,a46615a,a46616a,a46619a,a46622a,a46623a,a46624a,a46628a,a46629a,a46633a,a46634a,a46635a,a46639a,a46640a,a46643a,a46646a,a46647a,a46648a,a46652a,a46653a,a46657a,a46658a,a46659a,a46663a,a46664a,a46667a,a46670a,a46671a,a46672a,a46676a,a46677a,a46681a,a46682a,a46683a,a46687a,a46688a,a46691a,a46694a,a46695a,a46696a,a46700a,a46701a,a46705a,a46706a,a46707a,a46711a,a46712a,a46715a,a46718a,a46719a,a46720a,a46724a,a46725a,a46729a,a46730a,a46731a,a46735a,a46736a,a46739a,a46742a,a46743a,a46744a,a46748a,a46749a,a46753a,a46754a,a46755a,a46759a,a46760a,a46763a,a46766a,a46767a,a46768a,a46772a,a46773a,a46777a,a46778a,a46779a,a46783a,a46784a,a46787a,a46790a,a46791a,a46792a,a46796a,a46797a,a46801a,a46802a,a46803a,a46807a,a46808a,a46811a,a46814a,a46815a,a46816a,a46820a,a46821a,a46825a,a46826a,a46827a,a46831a,a46832a,a46835a,a46838a,a46839a,a46840a,a46844a,a46845a,a46849a,a46850a,a46851a,a46855a,a46856a,a46859a,a46862a,a46863a,a46864a,a46868a,a46869a,a46873a,a46874a,a46875a,a46879a,a46880a,a46883a,a46886a,a46887a,a46888a,a46892a,a46893a,a46897a,a46898a,a46899a,a46903a,a46904a,a46907a,a46910a,a46911a,a46912a,a46916a,a46917a,a46921a,a46922a,a46923a,a46927a,a46928a,a46931a,a46934a,a46935a,a46936a,a46940a,a46941a,a46945a,a46946a,a46947a,a46951a,a46952a,a46955a,a46958a,a46959a,a46960a,a46964a,a46965a,a46969a,a46970a,a46971a,a46975a,a46976a,a46979a,a46982a,a46983a,a46984a,a46988a,a46989a,a46993a,a46994a,a46995a,a46999a,a47000a,a47003a,a47006a,a47007a,a47008a,a47012a,a47013a,a47017a,a47018a,a47019a,a47023a,a47024a,a47027a,a47030a,a47031a,a47032a,a47036a,a47037a,a47041a,a47042a,a47043a,a47047a,a47048a,a47051a,a47054a,a47055a,a47056a,a47060a,a47061a,a47065a,a47066a,a47067a,a47071a,a47072a,a47075a,a47078a,a47079a,a47080a,a47084a,a47085a,a47089a,a47090a,a47091a,a47095a,a47096a,a47099a,a47102a,a47103a,a47104a,a47108a,a47109a,a47113a,a47114a,a47115a,a47119a,a47120a,a47123a,a47126a,a47127a,a47128a,a47132a,a47133a,a47137a,a47138a,a47139a,a47143a,a47144a,a47147a,a47150a,a47151a,a47152a,a47156a,a47157a,a47161a,a47162a,a47163a,a47167a,a47168a,a47171a,a47174a,a47175a,a47176a,a47180a,a47181a,a47185a,a47186a,a47187a,a47191a,a47192a,a47195a,a47198a,a47199a,a47200a,a47204a,a47205a,a47209a,a47210a,a47211a,a47215a,a47216a,a47219a,a47222a,a47223a,a47224a,a47228a,a47229a,a47233a,a47234a,a47235a,a47239a,a47240a,a47243a,a47246a,a47247a,a47248a,a47252a,a47253a,a47257a,a47258a,a47259a,a47263a,a47264a,a47267a,a47270a,a47271a,a47272a,a47276a,a47277a,a47281a,a47282a,a47283a,a47287a,a47288a,a47291a,a47294a,a47295a,a47296a,a47300a,a47301a,a47305a,a47306a,a47307a,a47311a,a47312a,a47315a,a47318a,a47319a,a47320a,a47324a,a47325a,a47329a,a47330a,a47331a,a47335a,a47336a,a47339a,a47342a,a47343a,a47344a,a47348a,a47349a,a47353a,a47354a,a47355a,a47359a,a47360a,a47363a,a47366a,a47367a,a47368a,a47372a,a47373a,a47377a,a47378a,a47379a,a47383a,a47384a,a47387a,a47390a,a47391a,a47392a,a47396a,a47397a,a47401a,a47402a,a47403a,a47407a,a47408a,a47411a,a47414a,a47415a,a47416a,a47420a,a47421a,a47425a,a47426a,a47427a,a47431a,a47432a,a47435a,a47438a,a47439a,a47440a,a47444a,a47445a,a47449a,a47450a,a47451a,a47455a,a47456a,a47459a,a47462a,a47463a,a47464a,a47468a,a47469a,a47473a,a47474a,a47475a,a47479a,a47480a,a47483a,a47486a,a47487a,a47488a,a47492a,a47493a,a47497a,a47498a,a47499a,a47503a,a47504a,a47507a,a47510a,a47511a,a47512a,a47516a,a47517a,a47521a,a47522a,a47523a,a47527a,a47528a,a47531a,a47534a,a47535a,a47536a,a47540a,a47541a,a47545a,a47546a,a47547a,a47551a,a47552a,a47555a,a47558a,a47559a,a47560a,a47564a,a47565a,a47569a,a47570a,a47571a,a47575a,a47576a,a47579a,a47582a,a47583a,a47584a,a47588a,a47589a,a47593a,a47594a,a47595a,a47599a,a47600a,a47603a,a47606a,a47607a,a47608a,a47612a,a47613a,a47617a,a47618a,a47619a,a47623a,a47624a,a47627a,a47630a,a47631a,a47632a,a47636a,a47637a,a47641a,a47642a,a47643a,a47647a,a47648a,a47651a,a47654a,a47655a,a47656a,a47660a,a47661a,a47665a,a47666a,a47667a,a47671a,a47672a,a47675a,a47678a,a47679a,a47680a,a47684a,a47685a,a47689a,a47690a,a47691a,a47695a,a47696a,a47699a,a47702a,a47703a,a47704a,a47708a,a47709a,a47713a,a47714a,a47715a,a47719a,a47720a,a47723a,a47726a,a47727a,a47728a,a47732a,a47733a,a47737a,a47738a,a47739a,a47743a,a47744a,a47747a,a47750a,a47751a,a47752a,a47756a,a47757a,a47761a,a47762a,a47763a,a47767a,a47768a,a47771a,a47774a,a47775a,a47776a,a47780a,a47781a,a47785a,a47786a,a47787a,a47791a,a47792a,a47795a,a47798a,a47799a,a47800a,a47804a,a47805a,a47809a,a47810a,a47811a,a47815a,a47816a,a47819a,a47822a,a47823a,a47824a,a47828a,a47829a,a47833a,a47834a,a47835a,a47839a,a47840a,a47843a,a47846a,a47847a,a47848a,a47852a,a47853a,a47857a,a47858a,a47859a,a47863a,a47864a,a47867a,a47870a,a47871a,a47872a,a47876a,a47877a,a47881a,a47882a,a47883a,a47887a,a47888a,a47891a,a47894a,a47895a,a47896a,a47900a,a47901a,a47905a,a47906a,a47907a,a47911a,a47912a,a47915a,a47918a,a47919a,a47920a,a47924a,a47925a,a47929a,a47930a,a47931a,a47935a,a47936a,a47939a,a47942a,a47943a,a47944a,a47948a,a47949a,a47953a,a47954a,a47955a,a47959a,a47960a,a47963a,a47966a,a47967a,a47968a,a47972a,a47973a,a47977a,a47978a,a47979a,a47983a,a47984a,a47987a,a47990a,a47991a,a47992a,a47996a,a47997a,a48001a,a48002a,a48003a,a48007a,a48008a,a48011a,a48014a,a48015a,a48016a,a48020a,a48021a,a48025a,a48026a,a48027a,a48031a,a48032a,a48035a,a48038a,a48039a,a48040a,a48044a,a48045a,a48049a,a48050a,a48051a,a48055a,a48056a,a48059a,a48062a,a48063a,a48064a,a48068a,a48069a,a48073a,a48074a,a48075a,a48079a,a48080a,a48083a,a48086a,a48087a,a48088a,a48092a,a48093a,a48097a,a48098a,a48099a,a48103a,a48104a,a48107a,a48110a,a48111a,a48112a,a48116a,a48117a,a48121a,a48122a,a48123a,a48127a,a48128a,a48131a,a48134a,a48135a,a48136a,a48140a,a48141a,a48145a,a48146a,a48147a,a48151a,a48152a,a48155a,a48158a,a48159a,a48160a,a48164a,a48165a,a48169a,a48170a,a48171a,a48175a,a48176a,a48179a,a48182a,a48183a,a48184a,a48188a,a48189a,a48193a,a48194a,a48195a,a48199a,a48200a,a48203a,a48206a,a48207a,a48208a,a48212a,a48213a,a48217a,a48218a,a48219a,a48223a,a48224a,a48227a,a48230a,a48231a,a48232a,a48236a,a48237a,a48241a,a48242a,a48243a,a48247a,a48248a,a48251a,a48254a,a48255a,a48256a,a48260a,a48261a,a48265a,a48266a,a48267a,a48271a,a48272a,a48275a,a48278a,a48279a,a48280a,a48284a,a48285a,a48289a,a48290a,a48291a,a48295a,a48296a,a48299a,a48302a,a48303a,a48304a,a48308a,a48309a,a48313a,a48314a,a48315a,a48319a,a48320a,a48323a,a48326a,a48327a,a48328a,a48332a,a48333a,a48337a,a48338a,a48339a,a48343a,a48344a,a48347a,a48350a,a48351a,a48352a,a48356a,a48357a,a48361a,a48362a,a48363a,a48367a,a48368a,a48371a,a48374a,a48375a,a48376a,a48380a,a48381a,a48385a,a48386a,a48387a,a48391a,a48392a,a48395a,a48398a,a48399a,a48400a,a48404a,a48405a,a48409a,a48410a,a48411a,a48415a,a48416a,a48419a,a48422a,a48423a,a48424a,a48428a,a48429a,a48433a,a48434a,a48435a,a48439a,a48440a,a48443a,a48446a,a48447a,a48448a,a48452a,a48453a,a48457a,a48458a,a48459a,a48463a,a48464a,a48467a,a48470a,a48471a,a48472a,a48476a,a48477a,a48481a,a48482a,a48483a,a48487a,a48488a,a48491a,a48494a,a48495a,a48496a,a48500a,a48501a,a48505a,a48506a,a48507a,a48511a,a48512a,a48515a,a48518a,a48519a,a48520a,a48524a,a48525a,a48529a,a48530a,a48531a,a48535a,a48536a,a48539a,a48542a,a48543a,a48544a,a48548a,a48549a,a48553a,a48554a,a48555a,a48559a,a48560a,a48563a,a48566a,a48567a,a48568a,a48572a,a48573a,a48577a,a48578a,a48579a,a48583a,a48584a,a48587a,a48590a,a48591a,a48592a,a48596a,a48597a,a48601a,a48602a,a48603a,a48607a,a48608a,a48611a,a48614a,a48615a,a48616a,a48620a,a48621a,a48625a,a48626a,a48627a,a48631a,a48632a,a48635a,a48638a,a48639a,a48640a,a48644a,a48645a,a48649a,a48650a,a48651a,a48655a,a48656a,a48659a,a48662a,a48663a,a48664a,a48668a,a48669a,a48673a,a48674a,a48675a,a48679a,a48680a,a48683a,a48686a,a48687a,a48688a,a48692a,a48693a,a48697a,a48698a,a48699a,a48703a,a48704a,a48707a,a48710a,a48711a,a48712a,a48716a,a48717a,a48721a,a48722a,a48723a,a48727a,a48728a,a48731a,a48734a,a48735a,a48736a,a48740a,a48741a,a48745a,a48746a,a48747a,a48751a,a48752a,a48755a,a48758a,a48759a,a48760a,a48764a,a48765a,a48769a,a48770a,a48771a,a48775a,a48776a,a48779a,a48782a,a48783a,a48784a,a48788a,a48789a,a48793a,a48794a,a48795a,a48799a,a48800a,a48803a,a48806a,a48807a,a48808a,a48812a,a48813a,a48817a,a48818a,a48819a,a48823a,a48824a,a48827a,a48830a,a48831a,a48832a,a48836a,a48837a,a48841a,a48842a,a48843a,a48847a,a48848a,a48851a,a48854a,a48855a,a48856a,a48860a,a48861a,a48865a,a48866a,a48867a,a48871a,a48872a,a48875a,a48878a,a48879a,a48880a,a48884a,a48885a,a48889a,a48890a,a48891a,a48895a,a48896a,a48899a,a48902a,a48903a,a48904a,a48908a,a48909a,a48913a,a48914a,a48915a,a48919a,a48920a,a48923a,a48926a,a48927a,a48928a,a48932a,a48933a,a48937a,a48938a,a48939a,a48943a,a48944a,a48947a,a48950a,a48951a,a48952a,a48956a,a48957a,a48961a,a48962a,a48963a,a48967a,a48968a,a48971a,a48974a,a48975a,a48976a,a48980a,a48981a,a48985a,a48986a,a48987a,a48991a,a48992a,a48995a,a48998a,a48999a,a49000a,a49004a,a49005a,a49009a,a49010a,a49011a,a49015a,a49016a,a49019a,a49022a,a49023a,a49024a,a49028a,a49029a,a49033a,a49034a,a49035a,a49039a,a49040a,a49043a,a49046a,a49047a,a49048a,a49052a,a49053a,a49057a,a49058a,a49059a,a49063a,a49064a,a49067a,a49070a,a49071a,a49072a,a49076a,a49077a,a49081a,a49082a,a49083a,a49087a,a49088a,a49091a,a49094a,a49095a,a49096a,a49100a,a49101a,a49105a,a49106a,a49107a,a49111a,a49112a,a49115a,a49118a,a49119a,a49120a,a49124a,a49125a,a49129a,a49130a,a49131a,a49135a,a49136a,a49139a,a49142a,a49143a,a49144a,a49148a,a49149a,a49153a,a49154a,a49155a,a49159a,a49160a,a49163a,a49166a,a49167a,a49168a,a49172a,a49173a,a49177a,a49178a,a49179a,a49183a,a49184a,a49187a,a49190a,a49191a,a49192a,a49196a,a49197a,a49201a,a49202a,a49203a,a49207a,a49208a,a49211a,a49214a,a49215a,a49216a,a49220a,a49221a,a49225a,a49226a,a49227a,a49231a,a49232a,a49235a,a49238a,a49239a,a49240a,a49244a,a49245a,a49249a,a49250a,a49251a,a49255a,a49256a,a49259a,a49262a,a49263a,a49264a,a49268a,a49269a,a49273a,a49274a,a49275a,a49279a,a49280a,a49283a,a49286a,a49287a,a49288a,a49292a,a49293a,a49297a,a49298a,a49299a,a49303a,a49304a,a49307a,a49310a,a49311a,a49312a,a49316a,a49317a,a49321a,a49322a,a49323a,a49327a,a49328a,a49331a,a49334a,a49335a,a49336a,a49340a,a49341a,a49345a,a49346a,a49347a,a49351a,a49352a,a49355a,a49358a,a49359a,a49360a,a49364a,a49365a,a49369a,a49370a,a49371a,a49375a,a49376a,a49379a,a49382a,a49383a,a49384a,a49388a,a49389a,a49393a,a49394a,a49395a,a49399a,a49400a,a49403a,a49406a,a49407a,a49408a,a49412a,a49413a,a49417a,a49418a,a49419a,a49423a,a49424a,a49427a,a49430a,a49431a,a49432a,a49436a,a49437a,a49441a,a49442a,a49443a,a49447a,a49448a,a49451a,a49454a,a49455a,a49456a,a49460a,a49461a,a49465a,a49466a,a49467a,a49471a,a49472a,a49475a,a49478a,a49479a,a49480a,a49484a,a49485a,a49489a,a49490a,a49491a,a49495a,a49496a,a49499a,a49502a,a49503a,a49504a,a49508a,a49509a,a49513a,a49514a,a49515a,a49519a,a49520a,a49523a,a49526a,a49527a,a49528a,a49532a,a49533a,a49537a,a49538a,a49539a,a49543a,a49544a,a49547a,a49550a,a49551a,a49552a,a49556a,a49557a,a49561a,a49562a,a49563a,a49567a,a49568a,a49571a,a49574a,a49575a,a49576a,a49580a,a49581a,a49585a,a49586a,a49587a,a49591a,a49592a,a49595a,a49598a,a49599a,a49600a,a49604a,a49605a,a49609a,a49610a,a49611a,a49615a,a49616a,a49619a,a49622a,a49623a,a49624a,a49628a,a49629a,a49633a,a49634a,a49635a,a49639a,a49640a,a49643a,a49646a,a49647a,a49648a,a49652a,a49653a,a49657a,a49658a,a49659a,a49663a,a49664a,a49667a,a49670a,a49671a,a49672a,a49676a,a49677a,a49681a,a49682a,a49683a,a49687a,a49688a,a49691a,a49694a,a49695a,a49696a,a49700a,a49701a,a49705a,a49706a,a49707a,a49711a,a49712a,a49715a,a49718a,a49719a,a49720a,a49724a,a49725a,a49729a,a49730a,a49731a,a49735a,a49736a,a49739a,a49742a,a49743a,a49744a,a49748a,a49749a,a49753a,a49754a,a49755a,a49759a,a49760a,a49763a,a49766a,a49767a,a49768a,a49772a,a49773a,a49777a,a49778a,a49779a,a49783a,a49784a,a49787a,a49790a,a49791a,a49792a,a49796a,a49797a,a49801a,a49802a,a49803a,a49807a,a49808a,a49811a,a49814a,a49815a,a49816a,a49820a,a49821a,a49825a,a49826a,a49827a,a49831a,a49832a,a49835a,a49838a,a49839a,a49840a,a49844a,a49845a,a49849a,a49850a,a49851a,a49855a,a49856a,a49859a,a49862a,a49863a,a49864a,a49868a,a49869a,a49873a,a49874a,a49875a,a49879a,a49880a,a49883a,a49886a,a49887a,a49888a,a49892a,a49893a,a49897a,a49898a,a49899a,a49903a,a49904a,a49907a,a49910a,a49911a,a49912a,a49916a,a49917a,a49921a,a49922a,a49923a,a49927a,a49928a,a49931a,a49934a,a49935a,a49936a,a49940a,a49941a,a49945a,a49946a,a49947a,a49951a,a49952a,a49955a,a49958a,a49959a,a49960a,a49964a,a49965a,a49969a,a49970a,a49971a,a49975a,a49976a,a49979a,a49982a,a49983a,a49984a,a49988a,a49989a,a49993a,a49994a,a49995a,a49999a,a50000a,a50003a,a50006a,a50007a,a50008a,a50012a,a50013a,a50017a,a50018a,a50019a,a50023a,a50024a,a50027a,a50030a,a50031a,a50032a,a50036a,a50037a,a50041a,a50042a,a50043a,a50047a,a50048a,a50051a,a50054a,a50055a,a50056a,a50060a,a50061a,a50065a,a50066a,a50067a,a50071a,a50072a,a50075a,a50078a,a50079a,a50080a,a50084a,a50085a,a50089a,a50090a,a50091a,a50095a,a50096a,a50099a,a50102a,a50103a,a50104a,a50108a,a50109a,a50113a,a50114a,a50115a,a50119a,a50120a,a50123a,a50126a,a50127a,a50128a,a50132a,a50133a,a50137a,a50138a,a50139a,a50143a,a50144a,a50147a,a50150a,a50151a,a50152a,a50156a,a50157a,a50161a,a50162a,a50163a,a50167a,a50168a,a50171a,a50174a,a50175a,a50176a,a50180a,a50181a,a50185a,a50186a,a50187a,a50191a,a50192a,a50195a,a50198a,a50199a,a50200a,a50204a,a50205a,a50209a,a50210a,a50211a,a50215a,a50216a,a50219a,a50222a,a50223a,a50224a,a50228a,a50229a,a50233a,a50234a,a50235a,a50239a,a50240a,a50243a,a50246a,a50247a,a50248a,a50252a,a50253a,a50257a,a50258a,a50259a,a50263a,a50264a,a50267a,a50270a,a50271a,a50272a,a50276a,a50277a,a50281a,a50282a,a50283a,a50287a,a50288a,a50291a,a50294a,a50295a,a50296a,a50300a,a50301a,a50305a,a50306a,a50307a,a50311a,a50312a,a50315a,a50318a,a50319a,a50320a,a50324a,a50325a,a50329a,a50330a,a50331a,a50335a,a50336a,a50339a,a50342a,a50343a,a50344a,a50348a,a50349a,a50353a,a50354a,a50355a,a50359a,a50360a,a50363a,a50366a,a50367a,a50368a,a50372a,a50373a,a50377a,a50378a,a50379a,a50383a,a50384a,a50387a,a50390a,a50391a,a50392a,a50396a,a50397a,a50401a,a50402a,a50403a,a50407a,a50408a,a50411a,a50414a,a50415a,a50416a,a50420a,a50421a,a50425a,a50426a,a50427a,a50431a,a50432a,a50435a,a50438a,a50439a,a50440a,a50444a,a50445a,a50449a,a50450a,a50451a,a50455a,a50456a,a50459a,a50462a,a50463a,a50464a,a50468a,a50469a,a50473a,a50474a,a50475a,a50479a,a50480a,a50483a,a50486a,a50487a,a50488a,a50492a,a50493a,a50497a,a50498a,a50499a,a50503a,a50504a,a50507a,a50510a,a50511a,a50512a,a50516a,a50517a,a50521a,a50522a,a50523a,a50527a,a50528a,a50531a,a50534a,a50535a,a50536a,a50540a,a50541a,a50545a,a50546a,a50547a,a50551a,a50552a,a50555a,a50558a,a50559a,a50560a,a50564a,a50565a,a50569a,a50570a,a50571a,a50575a,a50576a,a50579a,a50582a,a50583a,a50584a,a50588a,a50589a,a50593a,a50594a,a50595a,a50599a,a50600a,a50603a,a50606a,a50607a,a50608a,a50612a,a50613a,a50617a,a50618a,a50619a,a50623a,a50624a,a50627a,a50630a,a50631a,a50632a,a50636a,a50637a,a50641a,a50642a,a50643a,a50647a,a50648a,a50651a,a50654a,a50655a,a50656a,a50660a,a50661a,a50665a,a50666a,a50667a,a50671a,a50672a,a50675a,a50678a,a50679a,a50680a,a50684a,a50685a,a50689a,a50690a,a50691a,a50695a,a50696a,a50699a,a50702a,a50703a,a50704a,a50708a,a50709a,a50713a,a50714a,a50715a,a50719a,a50720a,a50723a,a50726a,a50727a,a50728a,a50732a,a50733a,a50737a,a50738a,a50739a,a50743a,a50744a,a50747a,a50750a,a50751a,a50752a,a50756a,a50757a,a50761a,a50762a,a50763a,a50767a,a50768a,a50771a,a50774a,a50775a,a50776a,a50780a,a50781a,a50785a,a50786a,a50787a,a50791a,a50792a,a50795a,a50798a,a50799a,a50800a,a50804a,a50805a,a50809a,a50810a,a50811a,a50815a,a50816a,a50819a,a50822a,a50823a,a50824a,a50828a,a50829a,a50833a,a50834a,a50835a,a50839a,a50840a,a50843a,a50846a,a50847a,a50848a,a50852a,a50853a,a50857a,a50858a,a50859a,a50863a,a50864a,a50867a,a50870a,a50871a,a50872a,a50876a,a50877a,a50881a,a50882a,a50883a,a50887a,a50888a,a50891a,a50894a,a50895a,a50896a,a50900a,a50901a,a50905a,a50906a,a50907a,a50911a,a50912a,a50915a,a50918a,a50919a,a50920a,a50924a,a50925a,a50929a,a50930a,a50931a,a50935a,a50936a,a50939a,a50942a,a50943a,a50944a,a50948a,a50949a,a50953a,a50954a,a50955a,a50959a,a50960a,a50963a,a50966a,a50967a,a50968a,a50972a,a50973a,a50977a,a50978a,a50979a,a50983a,a50984a,a50987a,a50990a,a50991a,a50992a,a50996a,a50997a,a51001a,a51002a,a51003a,a51007a,a51008a,a51011a,a51014a,a51015a,a51016a,a51020a,a51021a,a51025a,a51026a,a51027a,a51031a,a51032a,a51035a,a51038a,a51039a,a51040a,a51044a,a51045a,a51049a,a51050a,a51051a,a51055a,a51056a,a51059a,a51062a,a51063a,a51064a,a51068a,a51069a,a51073a,a51074a,a51075a,a51079a,a51080a,a51083a,a51086a,a51087a,a51088a,a51092a,a51093a,a51097a,a51098a,a51099a,a51103a,a51104a,a51107a,a51110a,a51111a,a51112a,a51116a,a51117a,a51121a,a51122a,a51123a,a51127a,a51128a,a51131a,a51134a,a51135a,a51136a,a51140a,a51141a,a51145a,a51146a,a51147a,a51151a,a51152a,a51155a,a51158a,a51159a,a51160a,a51164a,a51165a,a51169a,a51170a,a51171a,a51175a,a51176a,a51179a,a51182a,a51183a,a51184a,a51188a,a51189a,a51193a,a51194a,a51195a,a51199a,a51200a,a51203a,a51206a,a51207a,a51208a,a51212a,a51213a,a51217a,a51218a,a51219a,a51223a,a51224a,a51227a,a51230a,a51231a,a51232a,a51236a,a51237a,a51241a,a51242a,a51243a,a51247a,a51248a,a51251a,a51254a,a51255a,a51256a,a51260a,a51261a,a51265a,a51266a,a51267a,a51271a,a51272a,a51275a,a51278a,a51279a,a51280a,a51284a,a51285a,a51289a,a51290a,a51291a,a51295a,a51296a,a51299a,a51302a,a51303a,a51304a,a51308a,a51309a,a51313a,a51314a,a51315a,a51319a,a51320a,a51323a,a51326a,a51327a,a51328a,a51332a,a51333a,a51337a,a51338a,a51339a,a51343a,a51344a,a51347a,a51350a,a51351a,a51352a,a51356a,a51357a,a51361a,a51362a,a51363a,a51367a,a51368a,a51371a,a51374a,a51375a,a51376a,a51380a,a51381a,a51385a,a51386a,a51387a,a51391a,a51392a,a51395a,a51398a,a51399a,a51400a,a51404a,a51405a,a51409a,a51410a,a51411a,a51415a,a51416a,a51419a,a51422a,a51423a,a51424a,a51428a,a51429a,a51433a,a51434a,a51435a,a51439a,a51440a,a51443a,a51446a,a51447a,a51448a,a51452a,a51453a,a51457a,a51458a,a51459a,a51463a,a51464a,a51467a,a51470a,a51471a,a51472a,a51476a,a51477a,a51481a,a51482a,a51483a,a51487a,a51488a,a51491a,a51494a,a51495a,a51496a,a51500a,a51501a,a51505a,a51506a,a51507a,a51511a,a51512a,a51515a,a51518a,a51519a,a51520a,a51524a,a51525a,a51529a,a51530a,a51531a,a51535a,a51536a,a51539a,a51542a,a51543a,a51544a,a51548a,a51549a,a51553a,a51554a,a51555a,a51559a,a51560a,a51563a,a51566a,a51567a,a51568a,a51572a,a51573a,a51577a,a51578a,a51579a,a51583a,a51584a,a51587a,a51590a,a51591a,a51592a,a51596a,a51597a,a51601a,a51602a,a51603a,a51607a,a51608a,a51611a,a51614a,a51615a,a51616a,a51620a,a51621a,a51625a,a51626a,a51627a,a51631a,a51632a,a51635a,a51638a,a51639a,a51640a,a51644a,a51645a,a51649a,a51650a,a51651a,a51655a,a51656a,a51659a,a51662a,a51663a,a51664a,a51668a,a51669a,a51673a,a51674a,a51675a,a51679a,a51680a,a51683a,a51686a,a51687a,a51688a,a51692a,a51693a,a51697a,a51698a,a51699a,a51703a,a51704a,a51707a,a51710a,a51711a,a51712a,a51716a,a51717a,a51721a,a51722a,a51723a,a51727a,a51728a,a51731a,a51734a,a51735a,a51736a,a51740a,a51741a,a51745a,a51746a,a51747a,a51751a,a51752a,a51755a,a51758a,a51759a,a51760a,a51764a,a51765a,a51769a,a51770a,a51771a,a51775a,a51776a,a51779a,a51782a,a51783a,a51784a,a51788a,a51789a,a51793a,a51794a,a51795a,a51799a,a51800a,a51803a,a51806a,a51807a,a51808a,a51812a,a51813a,a51817a,a51818a,a51819a,a51823a,a51824a,a51827a,a51830a,a51831a,a51832a,a51836a,a51837a,a51841a,a51842a,a51843a,a51847a,a51848a,a51851a,a51854a,a51855a,a51856a,a51860a,a51861a,a51865a,a51866a,a51867a,a51871a,a51872a,a51875a,a51878a,a51879a,a51880a,a51884a,a51885a,a51889a,a51890a,a51891a,a51895a,a51896a,a51899a,a51902a,a51903a,a51904a,a51908a,a51909a,a51913a,a51914a,a51915a,a51919a,a51920a,a51923a,a51926a,a51927a,a51928a,a51932a,a51933a,a51937a,a51938a,a51939a,a51943a,a51944a,a51947a,a51950a,a51951a,a51952a,a51956a,a51957a,a51961a,a51962a,a51963a,a51967a,a51968a,a51971a,a51974a,a51975a,a51976a,a51980a,a51981a,a51985a,a51986a,a51987a,a51991a,a51992a,a51995a,a51998a,a51999a,a52000a,a52004a,a52005a,a52009a,a52010a,a52011a,a52015a,a52016a,a52019a,a52022a,a52023a,a52024a,a52028a,a52029a,a52033a,a52034a,a52035a,a52039a,a52040a,a52043a,a52046a,a52047a,a52048a,a52052a,a52053a,a52057a,a52058a,a52059a,a52063a,a52064a,a52067a,a52070a,a52071a,a52072a,a52076a,a52077a,a52081a,a52082a,a52083a,a52087a,a52088a,a52091a,a52094a,a52095a,a52096a,a52100a,a52101a,a52105a,a52106a,a52107a,a52111a,a52112a,a52115a,a52118a,a52119a,a52120a,a52124a,a52125a,a52129a,a52130a,a52131a,a52135a,a52136a,a52139a,a52142a,a52143a,a52144a,a52148a,a52149a,a52153a,a52154a,a52155a,a52159a,a52160a,a52163a,a52166a,a52167a,a52168a,a52172a,a52173a,a52177a,a52178a,a52179a,a52183a,a52184a,a52187a,a52190a,a52191a,a52192a,a52196a,a52197a,a52201a,a52202a,a52203a,a52207a,a52208a,a52211a,a52214a,a52215a,a52216a,a52220a,a52221a,a52225a,a52226a,a52227a,a52231a,a52232a,a52235a,a52238a,a52239a,a52240a,a52244a,a52245a,a52249a,a52250a,a52251a,a52255a,a52256a,a52259a,a52262a,a52263a,a52264a,a52268a,a52269a,a52273a,a52274a,a52275a,a52279a,a52280a,a52283a,a52286a,a52287a,a52288a,a52292a,a52293a,a52297a,a52298a,a52299a,a52303a,a52304a,a52307a,a52310a,a52311a,a52312a,a52316a,a52317a,a52321a,a52322a,a52323a,a52327a,a52328a,a52331a,a52334a,a52335a,a52336a,a52340a,a52341a,a52345a,a52346a,a52347a,a52351a,a52352a,a52355a,a52358a,a52359a,a52360a,a52364a,a52365a,a52369a,a52370a,a52371a,a52375a,a52376a,a52379a,a52382a,a52383a,a52384a,a52388a,a52389a,a52393a,a52394a,a52395a,a52399a,a52400a,a52403a,a52406a,a52407a,a52408a,a52412a,a52413a,a52417a,a52418a,a52419a,a52423a,a52424a,a52427a,a52430a,a52431a,a52432a,a52436a,a52437a,a52441a,a52442a,a52443a,a52447a,a52448a,a52451a,a52454a,a52455a,a52456a,a52460a,a52461a,a52465a,a52466a,a52467a,a52471a,a52472a,a52475a,a52478a,a52479a,a52480a,a52484a,a52485a,a52489a,a52490a,a52491a,a52495a,a52496a,a52499a,a52502a,a52503a,a52504a,a52508a,a52509a,a52513a,a52514a,a52515a,a52519a,a52520a,a52523a,a52526a,a52527a,a52528a,a52532a,a52533a,a52537a,a52538a,a52539a,a52543a,a52544a,a52547a,a52550a,a52551a,a52552a,a52556a,a52557a,a52561a,a52562a,a52563a,a52567a,a52568a,a52571a,a52574a,a52575a,a52576a,a52580a,a52581a,a52585a,a52586a,a52587a,a52591a,a52592a,a52595a,a52598a,a52599a,a52600a,a52604a,a52605a,a52609a,a52610a,a52611a,a52615a,a52616a,a52619a,a52622a,a52623a,a52624a,a52628a,a52629a,a52633a,a52634a,a52635a,a52639a,a52640a,a52643a,a52646a,a52647a,a52648a,a52652a,a52653a,a52657a,a52658a,a52659a,a52663a,a52664a,a52667a,a52670a,a52671a,a52672a,a52676a,a52677a,a52681a,a52682a,a52683a,a52687a,a52688a,a52691a,a52694a,a52695a,a52696a,a52700a,a52701a,a52705a,a52706a,a52707a,a52711a,a52712a,a52715a,a52718a,a52719a,a52720a,a52724a,a52725a,a52729a,a52730a,a52731a,a52735a,a52736a,a52739a,a52742a,a52743a,a52744a,a52748a,a52749a,a52753a,a52754a,a52755a,a52759a,a52760a,a52763a,a52766a,a52767a,a52768a,a52772a,a52773a,a52777a,a52778a,a52779a,a52783a,a52784a,a52787a,a52790a,a52791a,a52792a,a52796a,a52797a,a52801a,a52802a,a52803a,a52807a,a52808a,a52811a,a52814a,a52815a,a52816a,a52820a,a52821a,a52825a,a52826a,a52827a,a52831a,a52832a,a52835a,a52838a,a52839a,a52840a,a52844a,a52845a,a52849a,a52850a,a52851a,a52855a,a52856a,a52859a,a52862a,a52863a,a52864a,a52868a,a52869a,a52873a,a52874a,a52875a,a52879a,a52880a,a52883a,a52886a,a52887a,a52888a,a52892a,a52893a,a52897a,a52898a,a52899a,a52903a,a52904a,a52907a,a52910a,a52911a,a52912a,a52916a,a52917a,a52921a,a52922a,a52923a,a52927a,a52928a,a52931a,a52934a,a52935a,a52936a,a52940a,a52941a,a52945a,a52946a,a52947a,a52951a,a52952a,a52955a,a52958a,a52959a,a52960a,a52964a,a52965a,a52969a,a52970a,a52971a,a52975a,a52976a,a52979a,a52982a,a52983a,a52984a,a52988a,a52989a,a52993a,a52994a,a52995a,a52999a,a53000a,a53003a,a53006a,a53007a,a53008a,a53012a,a53013a,a53017a,a53018a,a53019a,a53023a,a53024a,a53027a,a53030a,a53031a,a53032a,a53036a,a53037a,a53041a,a53042a,a53043a,a53047a,a53048a,a53051a,a53054a,a53055a,a53056a,a53060a,a53061a,a53065a,a53066a,a53067a,a53071a,a53072a,a53075a,a53078a,a53079a,a53080a,a53084a,a53085a,a53089a,a53090a,a53091a,a53095a,a53096a,a53099a,a53102a,a53103a,a53104a,a53108a,a53109a,a53113a,a53114a,a53115a,a53119a,a53120a,a53123a,a53126a,a53127a,a53128a,a53132a,a53133a,a53137a,a53138a,a53139a,a53143a,a53144a,a53147a,a53150a,a53151a,a53152a,a53156a,a53157a,a53161a,a53162a,a53163a,a53167a,a53168a,a53171a,a53174a,a53175a,a53176a,a53180a,a53181a,a53185a,a53186a,a53187a,a53191a,a53192a,a53195a,a53198a,a53199a,a53200a,a53204a,a53205a,a53209a,a53210a,a53211a,a53215a,a53216a,a53219a,a53222a,a53223a,a53224a,a53228a,a53229a,a53233a,a53234a,a53235a,a53239a,a53240a,a53243a,a53246a,a53247a,a53248a,a53252a,a53253a,a53257a,a53258a,a53259a,a53263a,a53264a,a53267a,a53270a,a53271a,a53272a,a53276a,a53277a,a53281a,a53282a,a53283a,a53287a,a53288a,a53291a,a53294a,a53295a,a53296a,a53300a,a53301a,a53305a,a53306a,a53307a,a53311a,a53312a,a53315a,a53318a,a53319a,a53320a,a53324a,a53325a,a53329a,a53330a,a53331a,a53335a,a53336a,a53339a,a53342a,a53343a,a53344a,a53348a,a53349a,a53353a,a53354a,a53355a,a53359a,a53360a,a53363a,a53366a,a53367a,a53368a,a53372a,a53373a,a53377a,a53378a,a53379a,a53383a,a53384a,a53387a,a53390a,a53391a,a53392a,a53396a,a53397a,a53401a,a53402a,a53403a,a53407a,a53408a,a53411a,a53414a,a53415a,a53416a,a53420a,a53421a,a53425a,a53426a,a53427a,a53431a,a53432a,a53435a,a53438a,a53439a,a53440a,a53444a,a53445a,a53449a,a53450a,a53451a,a53455a,a53456a,a53459a,a53462a,a53463a,a53464a,a53468a,a53469a,a53473a,a53474a,a53475a,a53479a,a53480a,a53483a,a53486a,a53487a,a53488a,a53492a,a53493a,a53497a,a53498a,a53499a,a53503a,a53504a,a53507a,a53510a,a53511a,a53512a,a53516a,a53517a,a53521a,a53522a,a53523a,a53527a,a53528a,a53531a,a53534a,a53535a,a53536a,a53540a,a53541a,a53545a,a53546a,a53547a,a53551a,a53552a,a53555a,a53558a,a53559a,a53560a,a53564a,a53565a,a53569a,a53570a,a53571a,a53575a,a53576a,a53579a,a53582a,a53583a,a53584a,a53588a,a53589a,a53593a,a53594a,a53595a,a53599a,a53600a,a53603a,a53606a,a53607a,a53608a,a53612a,a53613a,a53617a,a53618a,a53619a,a53623a,a53624a,a53627a,a53630a,a53631a,a53632a,a53636a,a53637a,a53641a,a53642a,a53643a,a53647a,a53648a,a53651a,a53654a,a53655a,a53656a,a53660a,a53661a,a53665a,a53666a,a53667a,a53671a,a53672a,a53675a,a53678a,a53679a,a53680a,a53684a,a53685a,a53689a,a53690a,a53691a,a53695a,a53696a,a53699a,a53702a,a53703a,a53704a,a53708a,a53709a,a53713a,a53714a,a53715a,a53719a,a53720a,a53723a,a53726a,a53727a,a53728a,a53732a,a53733a,a53737a,a53738a,a53739a,a53743a,a53744a,a53747a,a53750a,a53751a,a53752a,a53756a,a53757a,a53761a,a53762a,a53763a,a53767a,a53768a,a53771a,a53774a,a53775a,a53776a,a53780a,a53781a,a53785a,a53786a,a53787a,a53791a,a53792a,a53795a,a53798a,a53799a,a53800a,a53804a,a53805a,a53809a,a53810a,a53811a,a53815a,a53816a,a53819a,a53822a,a53823a,a53824a,a53828a,a53829a,a53833a,a53834a,a53835a,a53839a,a53840a,a53843a,a53846a,a53847a,a53848a,a53852a,a53853a,a53857a,a53858a,a53859a,a53863a,a53864a,a53867a,a53870a,a53871a,a53872a,a53876a,a53877a,a53881a,a53882a,a53883a,a53887a,a53888a,a53891a,a53894a,a53895a,a53896a,a53900a,a53901a,a53905a,a53906a,a53907a,a53911a,a53912a,a53915a,a53918a,a53919a,a53920a,a53924a,a53925a,a53929a,a53930a,a53931a,a53935a,a53936a,a53939a,a53942a,a53943a,a53944a,a53948a,a53949a,a53953a,a53954a,a53955a,a53959a,a53960a,a53963a,a53966a,a53967a,a53968a,a53972a,a53973a,a53977a,a53978a,a53979a,a53983a,a53984a,a53987a,a53990a,a53991a,a53992a,a53996a,a53997a,a54001a,a54002a,a54003a,a54007a,a54008a,a54011a,a54014a,a54015a,a54016a,a54020a,a54021a,a54025a,a54026a,a54027a,a54031a,a54032a,a54035a,a54038a,a54039a,a54040a,a54044a,a54045a,a54049a,a54050a,a54051a,a54055a,a54056a,a54059a,a54062a,a54063a,a54064a,a54068a,a54069a,a54073a,a54074a,a54075a,a54079a,a54080a,a54083a,a54086a,a54087a,a54088a,a54092a,a54093a,a54097a,a54098a,a54099a,a54103a,a54104a,a54107a,a54110a,a54111a,a54112a,a54116a,a54117a,a54121a,a54122a,a54123a,a54127a,a54128a,a54131a,a54134a,a54135a,a54136a,a54140a,a54141a,a54145a,a54146a,a54147a,a54151a,a54152a,a54155a,a54158a,a54159a,a54160a,a54164a,a54165a,a54169a,a54170a,a54171a,a54175a,a54176a,a54179a,a54182a,a54183a,a54184a,a54188a,a54189a,a54193a,a54194a,a54195a,a54199a,a54200a,a54203a,a54206a,a54207a,a54208a,a54212a,a54213a,a54217a,a54218a,a54219a,a54223a,a54224a,a54227a,a54230a,a54231a,a54232a,a54236a,a54237a,a54241a,a54242a,a54243a,a54247a,a54248a,a54251a,a54254a,a54255a,a54256a,a54260a,a54261a,a54265a,a54266a,a54267a,a54271a,a54272a,a54275a,a54278a,a54279a,a54280a,a54284a,a54285a,a54289a,a54290a,a54291a,a54295a,a54296a,a54299a,a54302a,a54303a,a54304a,a54308a,a54309a,a54313a,a54314a,a54315a,a54319a,a54320a,a54323a,a54326a,a54327a,a54328a,a54332a,a54333a,a54337a,a54338a,a54339a,a54343a,a54344a,a54347a,a54350a,a54351a,a54352a,a54356a,a54357a,a54361a,a54362a,a54363a,a54367a,a54368a,a54371a,a54374a,a54375a,a54376a,a54380a,a54381a,a54385a,a54386a,a54387a,a54391a,a54392a,a54395a,a54398a,a54399a,a54400a,a54404a,a54405a,a54409a,a54410a,a54411a,a54415a,a54416a,a54419a,a54422a,a54423a,a54424a,a54428a,a54429a,a54433a,a54434a,a54435a,a54439a,a54440a,a54443a,a54446a,a54447a,a54448a,a54452a,a54453a,a54457a,a54458a,a54459a,a54463a,a54464a,a54467a,a54470a,a54471a,a54472a,a54476a,a54477a,a54481a,a54482a,a54483a,a54487a,a54488a,a54491a,a54494a,a54495a,a54496a,a54500a,a54501a,a54505a,a54506a,a54507a,a54511a,a54512a,a54515a,a54518a,a54519a,a54520a,a54524a,a54525a,a54529a,a54530a,a54531a,a54535a,a54536a,a54539a,a54542a,a54543a,a54544a,a54548a,a54549a,a54553a,a54554a,a54555a,a54559a,a54560a,a54563a,a54566a,a54567a,a54568a,a54572a,a54573a,a54577a,a54578a,a54579a,a54583a,a54584a,a54587a,a54590a,a54591a,a54592a,a54596a,a54597a,a54601a,a54602a,a54603a,a54607a,a54608a,a54611a,a54614a,a54615a,a54616a,a54620a,a54621a,a54625a,a54626a,a54627a,a54631a,a54632a,a54635a,a54638a,a54639a,a54640a,a54644a,a54645a,a54649a,a54650a,a54651a,a54655a,a54656a,a54659a,a54662a,a54663a,a54664a,a54668a,a54669a,a54673a,a54674a,a54675a,a54679a,a54680a,a54683a,a54686a,a54687a,a54688a,a54692a,a54693a,a54697a,a54698a,a54699a,a54703a,a54704a,a54707a,a54710a,a54711a,a54712a,a54716a,a54717a,a54721a,a54722a,a54723a,a54727a,a54728a,a54731a,a54734a,a54735a,a54736a,a54740a,a54741a,a54745a,a54746a,a54747a,a54751a,a54752a,a54755a,a54758a,a54759a,a54760a,a54764a,a54765a,a54769a,a54770a,a54771a,a54775a,a54776a,a54779a,a54782a,a54783a,a54784a,a54788a,a54789a,a54793a,a54794a,a54795a,a54799a,a54800a,a54803a,a54806a,a54807a,a54808a,a54812a,a54813a,a54817a,a54818a,a54819a,a54823a,a54824a,a54827a,a54830a,a54831a,a54832a,a54836a,a54837a,a54841a,a54842a,a54843a,a54847a,a54848a,a54851a,a54854a,a54855a,a54856a,a54860a,a54861a,a54865a,a54866a,a54867a,a54871a,a54872a,a54875a,a54878a,a54879a,a54880a,a54884a,a54885a,a54889a,a54890a,a54891a,a54895a,a54896a,a54899a,a54902a,a54903a,a54904a,a54908a,a54909a,a54913a,a54914a,a54915a,a54919a,a54920a,a54923a,a54926a,a54927a,a54928a,a54932a,a54933a,a54937a,a54938a,a54939a,a54943a,a54944a,a54947a,a54950a,a54951a,a54952a,a54956a,a54957a,a54961a,a54962a,a54963a,a54967a,a54968a,a54971a,a54974a,a54975a,a54976a,a54980a,a54981a,a54985a,a54986a,a54987a,a54991a,a54992a,a54995a,a54998a,a54999a,a55000a,a55004a,a55005a,a55009a,a55010a,a55011a,a55015a,a55016a,a55019a,a55022a,a55023a,a55024a,a55028a,a55029a,a55033a,a55034a,a55035a,a55039a,a55040a,a55043a,a55046a,a55047a,a55048a,a55052a,a55053a,a55057a,a55058a,a55059a,a55063a,a55064a,a55067a,a55070a,a55071a,a55072a,a55076a,a55077a,a55081a,a55082a,a55083a,a55087a,a55088a,a55091a,a55094a,a55095a,a55096a,a55100a,a55101a,a55105a,a55106a,a55107a,a55111a,a55112a,a55115a,a55118a,a55119a,a55120a,a55124a,a55125a,a55129a,a55130a,a55131a,a55135a,a55136a,a55139a,a55142a,a55143a,a55144a,a55148a,a55149a,a55153a,a55154a,a55155a,a55159a,a55160a,a55163a,a55166a,a55167a,a55168a,a55172a,a55173a,a55177a,a55178a,a55179a,a55183a,a55184a,a55187a,a55190a,a55191a,a55192a,a55196a,a55197a,a55201a,a55202a,a55203a,a55207a,a55208a,a55211a,a55214a,a55215a,a55216a,a55220a,a55221a,a55225a,a55226a,a55227a,a55231a,a55232a,a55235a,a55238a,a55239a,a55240a,a55244a,a55245a,a55249a,a55250a,a55251a,a55255a,a55256a,a55259a,a55262a,a55263a,a55264a,a55268a,a55269a,a55273a,a55274a,a55275a,a55279a,a55280a,a55283a,a55286a,a55287a,a55288a,a55292a,a55293a,a55297a,a55298a,a55299a,a55303a,a55304a,a55307a,a55310a,a55311a,a55312a,a55316a,a55317a,a55321a,a55322a,a55323a,a55327a,a55328a,a55331a,a55334a,a55335a,a55336a,a55340a,a55341a,a55345a,a55346a,a55347a,a55351a,a55352a,a55355a,a55358a,a55359a,a55360a,a55364a,a55365a,a55369a,a55370a,a55371a,a55375a,a55376a,a55379a,a55382a,a55383a,a55384a,a55388a,a55389a,a55393a,a55394a,a55395a,a55399a,a55400a,a55403a,a55406a,a55407a,a55408a,a55412a,a55413a,a55417a,a55418a,a55419a,a55423a,a55424a,a55427a,a55430a,a55431a,a55432a,a55436a,a55437a,a55441a,a55442a,a55443a,a55447a,a55448a,a55451a,a55454a,a55455a,a55456a,a55460a,a55461a,a55465a,a55466a,a55467a,a55471a,a55472a,a55475a,a55478a,a55479a,a55480a,a55484a,a55485a,a55489a,a55490a,a55491a,a55495a,a55496a,a55499a,a55502a,a55503a,a55504a,a55508a,a55509a,a55513a,a55514a,a55515a,a55519a,a55520a,a55523a,a55526a,a55527a,a55528a,a55532a,a55533a,a55537a,a55538a,a55539a,a55543a,a55544a,a55547a,a55550a,a55551a,a55552a,a55556a,a55557a,a55561a,a55562a,a55563a,a55567a,a55568a,a55571a,a55574a,a55575a,a55576a,a55580a,a55581a,a55585a,a55586a,a55587a,a55591a,a55592a,a55595a,a55598a,a55599a,a55600a,a55604a,a55605a,a55609a,a55610a,a55611a,a55615a,a55616a,a55619a,a55622a,a55623a,a55624a,a55628a,a55629a,a55633a,a55634a,a55635a,a55639a,a55640a,a55643a,a55646a,a55647a,a55648a,a55652a,a55653a,a55657a,a55658a,a55659a,a55663a,a55664a,a55667a,a55670a,a55671a,a55672a,a55676a,a55677a,a55681a,a55682a,a55683a,a55687a,a55688a,a55691a,a55694a,a55695a,a55696a,a55700a,a55701a,a55705a,a55706a,a55707a,a55711a,a55712a,a55715a,a55718a,a55719a,a55720a,a55724a,a55725a,a55729a,a55730a,a55731a,a55735a,a55736a,a55739a,a55742a,a55743a,a55744a,a55748a,a55749a,a55753a,a55754a,a55755a,a55759a,a55760a,a55763a,a55766a,a55767a,a55768a,a55772a,a55773a,a55777a,a55778a,a55779a,a55783a,a55784a,a55787a,a55790a,a55791a,a55792a,a55796a,a55797a,a55801a,a55802a,a55803a,a55807a,a55808a,a55811a,a55814a,a55815a,a55816a,a55820a,a55821a,a55825a,a55826a,a55827a,a55831a,a55832a,a55835a,a55838a,a55839a,a55840a,a55844a,a55845a,a55849a,a55850a,a55851a,a55855a,a55856a,a55859a,a55862a,a55863a,a55864a,a55868a,a55869a,a55873a,a55874a,a55875a,a55879a,a55880a,a55883a,a55886a,a55887a,a55888a,a55892a,a55893a,a55897a,a55898a,a55899a,a55903a,a55904a,a55907a,a55910a,a55911a,a55912a,a55916a,a55917a,a55921a,a55922a,a55923a,a55927a,a55928a,a55931a,a55934a,a55935a,a55936a,a55940a,a55941a,a55945a,a55946a,a55947a,a55951a,a55952a,a55955a,a55958a,a55959a,a55960a,a55964a,a55965a,a55969a,a55970a,a55971a,a55975a,a55976a,a55979a,a55982a,a55983a,a55984a,a55988a,a55989a,a55993a,a55994a,a55995a,a55999a,a56000a,a56003a,a56006a,a56007a,a56008a,a56012a,a56013a,a56017a,a56018a,a56019a,a56023a,a56024a,a56027a,a56030a,a56031a,a56032a,a56036a,a56037a,a56041a,a56042a,a56043a,a56047a,a56048a,a56051a,a56054a,a56055a,a56056a,a56060a,a56061a,a56065a,a56066a,a56067a,a56071a,a56072a,a56075a,a56078a,a56079a,a56080a,a56084a,a56085a,a56089a,a56090a,a56091a,a56095a,a56096a,a56099a,a56102a,a56103a,a56104a,a56108a,a56109a,a56113a,a56114a,a56115a,a56119a,a56120a,a56123a,a56126a,a56127a,a56128a,a56132a,a56133a,a56137a,a56138a,a56139a,a56143a,a56144a,a56147a,a56150a,a56151a,a56152a,a56156a,a56157a,a56161a,a56162a,a56163a,a56167a,a56168a,a56171a,a56174a,a56175a,a56176a,a56180a,a56181a,a56185a,a56186a,a56187a,a56191a,a56192a,a56195a,a56198a,a56199a,a56200a,a56204a,a56205a,a56209a,a56210a,a56211a,a56215a,a56216a,a56219a,a56222a,a56223a,a56224a,a56228a,a56229a,a56233a,a56234a,a56235a,a56239a,a56240a,a56243a,a56246a,a56247a,a56248a,a56252a,a56253a,a56257a,a56258a,a56259a,a56263a,a56264a,a56267a,a56270a,a56271a,a56272a,a56276a,a56277a,a56281a,a56282a,a56283a,a56287a,a56288a,a56291a,a56294a,a56295a,a56296a,a56300a,a56301a,a56305a,a56306a,a56307a,a56311a,a56312a,a56315a,a56318a,a56319a,a56320a,a56324a,a56325a,a56329a,a56330a,a56331a,a56335a,a56336a,a56339a,a56342a,a56343a,a56344a,a56348a,a56349a,a56353a,a56354a,a56355a,a56359a,a56360a,a56363a,a56366a,a56367a,a56368a,a56372a,a56373a,a56377a,a56378a,a56379a,a56383a,a56384a,a56387a,a56390a,a56391a,a56392a,a56396a,a56397a,a56401a,a56402a,a56403a,a56407a,a56408a,a56411a,a56414a,a56415a,a56416a,a56420a,a56421a,a56425a,a56426a,a56427a,a56431a,a56432a,a56435a,a56438a,a56439a,a56440a,a56444a,a56445a,a56449a,a56450a,a56451a,a56455a,a56456a,a56459a,a56462a,a56463a,a56464a,a56468a,a56469a,a56473a,a56474a,a56475a,a56479a,a56480a,a56483a,a56486a,a56487a,a56488a,a56492a,a56493a,a56497a,a56498a,a56499a,a56503a,a56504a,a56507a,a56510a,a56511a,a56512a,a56516a,a56517a,a56521a,a56522a,a56523a,a56527a,a56528a,a56531a,a56534a,a56535a,a56536a,a56540a,a56541a,a56545a,a56546a,a56547a,a56551a,a56552a,a56555a,a56558a,a56559a,a56560a,a56564a,a56565a,a56569a,a56570a,a56571a,a56575a,a56576a,a56579a,a56582a,a56583a,a56584a,a56588a,a56589a,a56593a,a56594a,a56595a,a56599a,a56600a,a56603a,a56606a,a56607a,a56608a,a56612a,a56613a,a56617a,a56618a,a56619a,a56623a,a56624a,a56627a,a56630a,a56631a,a56632a,a56636a,a56637a,a56641a,a56642a,a56643a,a56647a,a56648a,a56651a,a56654a,a56655a,a56656a,a56660a,a56661a,a56665a,a56666a,a56667a,a56671a,a56672a,a56675a,a56678a,a56679a,a56680a,a56684a,a56685a,a56689a,a56690a,a56691a,a56695a,a56696a,a56699a,a56702a,a56703a,a56704a,a56708a,a56709a,a56713a,a56714a,a56715a,a56719a,a56720a,a56723a,a56726a,a56727a,a56728a,a56732a,a56733a,a56737a,a56738a,a56739a,a56743a,a56744a,a56747a,a56750a,a56751a,a56752a,a56756a,a56757a,a56760a,a56763a,a56764a,a56765a,a56769a,a56770a,a56773a,a56776a,a56777a,a56778a,a56782a,a56783a,a56786a,a56789a,a56790a,a56791a,a56795a,a56796a,a56799a,a56802a,a56803a,a56804a,a56808a,a56809a,a56812a,a56815a,a56816a,a56817a,a56821a,a56822a,a56825a,a56828a,a56829a,a56830a,a56834a,a56835a,a56838a,a56841a,a56842a,a56843a,a56847a,a56848a,a56851a,a56854a,a56855a,a56856a,a56860a,a56861a,a56864a,a56867a,a56868a,a56869a,a56873a,a56874a,a56877a,a56880a,a56881a,a56882a,a56886a,a56887a,a56890a,a56893a,a56894a,a56895a,a56899a,a56900a,a56903a,a56906a,a56907a,a56908a,a56912a,a56913a,a56916a,a56919a,a56920a,a56921a,a56925a,a56926a,a56929a,a56932a,a56933a,a56934a,a56938a,a56939a,a56942a,a56945a,a56946a,a56947a,a56951a,a56952a,a56955a,a56958a,a56959a,a56960a,a56964a,a56965a,a56968a,a56971a,a56972a,a56973a,a56977a,a56978a,a56981a,a56984a,a56985a,a56986a,a56990a,a56991a,a56994a,a56997a,a56998a,a56999a,a57003a,a57004a,a57007a,a57010a,a57011a,a57012a,a57016a,a57017a,a57020a,a57023a,a57024a,a57025a,a57029a,a57030a,a57033a,a57036a,a57037a,a57038a,a57042a,a57043a,a57046a,a57049a,a57050a,a57051a,a57055a,a57056a,a57059a,a57062a,a57063a,a57064a,a57068a,a57069a,a57072a,a57075a,a57076a,a57077a,a57081a,a57082a,a57085a,a57088a,a57089a,a57090a,a57094a,a57095a,a57098a,a57101a,a57102a,a57103a,a57107a,a57108a,a57111a,a57114a,a57115a,a57116a,a57120a,a57121a,a57124a,a57127a,a57128a,a57129a,a57133a,a57134a,a57137a,a57140a,a57141a,a57142a,a57146a,a57147a,a57150a,a57153a,a57154a,a57155a,a57159a,a57160a,a57163a,a57166a,a57167a,a57168a,a57172a,a57173a,a57176a,a57179a,a57180a,a57181a,a57185a,a57186a,a57189a,a57192a,a57193a,a57194a,a57198a,a57199a,a57202a,a57205a,a57206a,a57207a,a57211a,a57212a,a57215a,a57218a,a57219a,a57220a,a57224a,a57225a,a57228a,a57231a,a57232a,a57233a,a57237a,a57238a,a57241a,a57244a,a57245a,a57246a,a57250a,a57251a,a57254a,a57257a,a57258a,a57259a,a57263a,a57264a,a57267a,a57270a,a57271a,a57272a,a57276a,a57277a,a57280a,a57283a,a57284a,a57285a,a57289a,a57290a,a57293a,a57296a,a57297a,a57298a,a57302a,a57303a,a57306a,a57309a,a57310a,a57311a,a57315a,a57316a,a57319a,a57322a,a57323a,a57324a,a57328a,a57329a,a57332a,a57335a,a57336a,a57337a,a57341a,a57342a,a57345a,a57348a,a57349a,a57350a,a57354a,a57355a,a57358a,a57361a,a57362a,a57363a,a57367a,a57368a,a57371a,a57374a,a57375a,a57376a,a57380a,a57381a,a57384a,a57387a,a57388a,a57389a,a57393a,a57394a,a57397a,a57400a,a57401a,a57402a,a57406a,a57407a,a57410a,a57413a,a57414a,a57415a,a57419a,a57420a,a57423a,a57426a,a57427a,a57428a,a57432a,a57433a,a57436a,a57439a,a57440a,a57441a,a57445a,a57446a,a57449a,a57452a,a57453a,a57454a,a57458a,a57459a,a57462a,a57465a,a57466a,a57467a,a57471a,a57472a,a57475a,a57478a,a57479a,a57480a,a57484a,a57485a,a57488a,a57491a,a57492a,a57493a,a57497a,a57498a,a57501a,a57504a,a57505a,a57506a,a57510a,a57511a,a57514a,a57517a,a57518a,a57519a,a57523a,a57524a,a57527a,a57530a,a57531a,a57532a,a57536a,a57537a,a57540a,a57543a,a57544a,a57545a,a57549a,a57550a,a57553a,a57556a,a57557a,a57558a,a57562a,a57563a,a57566a,a57569a,a57570a,a57571a,a57575a,a57576a,a57579a,a57582a,a57583a,a57584a,a57588a,a57589a,a57592a,a57595a,a57596a,a57597a,a57601a,a57602a,a57605a,a57608a,a57609a,a57610a,a57614a,a57615a,a57618a,a57621a,a57622a,a57623a,a57627a,a57628a,a57631a,a57634a,a57635a,a57636a,a57640a,a57641a,a57644a,a57647a,a57648a,a57649a,a57653a,a57654a,a57657a,a57660a,a57661a,a57662a,a57666a,a57667a,a57670a,a57673a,a57674a,a57675a,a57679a,a57680a,a57683a,a57686a,a57687a,a57688a,a57692a,a57693a,a57696a,a57699a,a57700a,a57701a,a57705a,a57706a,a57709a,a57712a,a57713a,a57714a,a57718a,a57719a,a57722a,a57725a,a57726a,a57727a,a57731a,a57732a,a57735a,a57738a,a57739a,a57740a,a57744a,a57745a,a57748a,a57751a,a57752a,a57753a,a57757a,a57758a,a57761a,a57764a,a57765a,a57766a,a57770a,a57771a,a57774a,a57777a,a57778a,a57779a,a57783a,a57784a,a57787a,a57790a,a57791a,a57792a,a57796a,a57797a,a57800a,a57803a,a57804a,a57805a,a57809a,a57810a,a57813a,a57816a,a57817a,a57818a,a57822a,a57823a,a57826a,a57829a,a57830a,a57831a,a57835a,a57836a,a57839a,a57842a,a57843a,a57844a,a57848a,a57849a,a57852a,a57855a,a57856a,a57857a,a57861a,a57862a,a57865a,a57868a,a57869a,a57870a,a57874a,a57875a,a57878a,a57881a,a57882a,a57883a,a57887a,a57888a,a57891a,a57894a,a57895a,a57896a,a57900a,a57901a,a57904a,a57907a,a57908a,a57909a,a57913a,a57914a,a57917a,a57920a,a57921a,a57922a,a57926a,a57927a,a57930a,a57933a,a57934a,a57935a,a57939a,a57940a,a57943a,a57946a,a57947a,a57948a,a57952a,a57953a,a57956a,a57959a,a57960a,a57961a,a57965a,a57966a,a57969a,a57972a,a57973a,a57974a,a57978a,a57979a,a57982a,a57985a,a57986a,a57987a,a57991a,a57992a,a57995a,a57998a,a57999a,a58000a,a58004a,a58005a,a58008a,a58011a,a58012a,a58013a,a58017a,a58018a,a58021a,a58024a,a58025a,a58026a,a58030a,a58031a,a58034a,a58037a,a58038a,a58039a,a58043a,a58044a,a58047a,a58050a,a58051a,a58052a,a58056a,a58057a,a58060a,a58063a,a58064a,a58065a,a58069a,a58070a,a58073a,a58076a,a58077a,a58078a,a58082a,a58083a,a58086a,a58089a,a58090a,a58091a,a58095a,a58096a,a58099a,a58102a,a58103a,a58104a,a58108a,a58109a,a58112a,a58115a,a58116a,a58117a,a58121a,a58122a,a58125a,a58128a,a58129a,a58130a,a58134a,a58135a,a58138a,a58141a,a58142a,a58143a,a58147a,a58148a,a58151a,a58154a,a58155a,a58156a,a58160a,a58161a,a58164a,a58167a,a58168a,a58169a,a58173a,a58174a,a58177a,a58180a,a58181a,a58182a,a58186a,a58187a,a58190a,a58193a,a58194a,a58195a,a58199a,a58200a,a58203a,a58206a,a58207a,a58208a,a58212a,a58213a,a58216a,a58219a,a58220a,a58221a,a58225a,a58226a,a58229a,a58232a,a58233a,a58234a,a58238a,a58239a,a58242a,a58245a,a58246a,a58247a,a58251a,a58252a,a58255a,a58258a,a58259a,a58260a,a58264a,a58265a,a58268a,a58271a,a58272a,a58273a,a58277a,a58278a,a58281a,a58284a,a58285a,a58286a,a58290a,a58291a,a58294a,a58297a,a58298a,a58299a,a58303a,a58304a,a58307a,a58310a,a58311a,a58312a,a58316a,a58317a,a58320a,a58323a,a58324a,a58325a,a58329a,a58330a,a58333a,a58336a,a58337a,a58338a,a58342a,a58343a,a58346a,a58349a,a58350a,a58351a,a58355a,a58356a,a58359a,a58362a,a58363a,a58364a,a58368a,a58369a,a58372a,a58375a,a58376a,a58377a,a58381a,a58382a,a58385a,a58388a,a58389a,a58390a,a58394a,a58395a,a58398a,a58401a,a58402a,a58403a,a58407a,a58408a,a58411a,a58414a,a58415a,a58416a,a58420a,a58421a,a58424a,a58427a,a58428a,a58429a,a58433a,a58434a,a58437a,a58440a,a58441a,a58442a,a58446a,a58447a,a58450a,a58453a,a58454a,a58455a,a58459a,a58460a,a58463a,a58466a,a58467a,a58468a,a58472a,a58473a,a58476a,a58479a,a58480a,a58481a,a58485a,a58486a,a58489a,a58492a,a58493a,a58494a,a58498a,a58499a,a58502a,a58505a,a58506a,a58507a,a58511a,a58512a,a58515a,a58518a,a58519a,a58520a,a58524a,a58525a,a58528a,a58531a,a58532a,a58533a,a58537a,a58538a,a58541a,a58544a,a58545a,a58546a,a58550a,a58551a,a58554a,a58557a,a58558a,a58559a,a58563a,a58564a,a58567a,a58570a,a58571a,a58572a,a58576a,a58577a,a58580a,a58583a,a58584a,a58585a,a58589a,a58590a,a58593a,a58596a,a58597a,a58598a,a58602a,a58603a,a58606a,a58609a,a58610a,a58611a,a58615a,a58616a,a58619a,a58622a,a58623a,a58624a,a58628a,a58629a,a58632a,a58635a,a58636a,a58637a,a58641a,a58642a,a58645a,a58648a,a58649a,a58650a,a58654a,a58655a,a58658a,a58661a,a58662a,a58663a,a58667a,a58668a,a58671a,a58674a,a58675a,a58676a,a58680a,a58681a,a58684a,a58687a,a58688a,a58689a,a58693a,a58694a,a58697a,a58700a,a58701a,a58702a,a58706a,a58707a,a58710a,a58713a,a58714a,a58715a,a58719a,a58720a,a58723a,a58726a,a58727a,a58728a,a58732a,a58733a,a58736a,a58739a,a58740a,a58741a,a58745a,a58746a,a58749a,a58752a,a58753a,a58754a,a58758a,a58759a,a58762a,a58765a,a58766a,a58767a,a58771a,a58772a,a58775a,a58778a,a58779a,a58780a,a58784a,a58785a,a58788a,a58791a,a58792a,a58793a,a58797a,a58798a,a58801a,a58804a,a58805a,a58806a,a58810a,a58811a,a58814a,a58817a,a58818a,a58819a,a58823a,a58824a,a58827a,a58830a,a58831a,a58832a,a58836a,a58837a,a58840a,a58843a,a58844a,a58845a,a58849a,a58850a,a58853a,a58856a,a58857a,a58858a,a58862a,a58863a,a58866a,a58869a,a58870a,a58871a,a58875a,a58876a,a58879a,a58882a,a58883a,a58884a,a58888a,a58889a,a58892a,a58895a,a58896a,a58897a,a58901a,a58902a,a58905a,a58908a,a58909a,a58910a,a58914a,a58915a,a58918a,a58921a,a58922a,a58923a,a58927a,a58928a,a58931a,a58934a,a58935a,a58936a,a58940a,a58941a,a58944a,a58947a,a58948a,a58949a,a58953a,a58954a,a58957a,a58960a,a58961a,a58962a,a58966a,a58967a,a58970a,a58973a,a58974a,a58975a,a58979a,a58980a,a58983a,a58986a,a58987a,a58988a,a58992a,a58993a,a58996a,a58999a,a59000a,a59001a,a59005a,a59006a,a59009a,a59012a,a59013a,a59014a,a59018a,a59019a,a59022a,a59025a,a59026a,a59027a,a59031a,a59032a,a59035a,a59038a,a59039a,a59040a,a59044a,a59045a,a59048a,a59051a,a59052a,a59053a,a59057a,a59058a,a59061a,a59064a,a59065a,a59066a,a59070a,a59071a,a59074a,a59077a,a59078a,a59079a,a59083a,a59084a,a59087a,a59090a,a59091a,a59092a,a59096a,a59097a,a59100a,a59103a,a59104a,a59105a,a59109a,a59110a,a59113a,a59116a,a59117a,a59118a,a59122a,a59123a,a59126a,a59129a,a59130a,a59131a,a59135a,a59136a,a59139a,a59142a,a59143a,a59144a,a59148a,a59149a,a59152a,a59155a,a59156a,a59157a,a59161a,a59162a,a59165a,a59168a,a59169a,a59170a,a59174a,a59175a,a59178a,a59181a,a59182a,a59183a,a59187a,a59188a,a59191a,a59194a,a59195a,a59196a,a59200a,a59201a,a59204a,a59207a,a59208a,a59209a,a59213a,a59214a,a59217a,a59220a,a59221a,a59222a,a59226a,a59227a,a59230a,a59233a,a59234a,a59235a,a59239a,a59240a,a59243a,a59246a,a59247a,a59248a,a59252a,a59253a,a59256a,a59259a,a59260a,a59261a,a59265a,a59266a,a59269a,a59272a,a59273a,a59274a,a59278a,a59279a,a59282a,a59285a,a59286a,a59287a,a59291a,a59292a,a59295a,a59298a,a59299a,a59300a,a59304a,a59305a,a59308a,a59311a,a59312a,a59313a,a59317a,a59318a,a59321a,a59324a,a59325a,a59326a,a59330a,a59331a,a59334a,a59337a,a59338a,a59339a,a59343a,a59344a,a59347a,a59350a,a59351a,a59352a,a59356a,a59357a,a59360a,a59363a,a59364a,a59365a,a59369a,a59370a,a59373a,a59376a,a59377a,a59378a,a59382a,a59383a,a59386a,a59389a,a59390a,a59391a,a59395a,a59396a,a59399a,a59402a,a59403a,a59404a,a59408a,a59409a,a59412a,a59415a,a59416a,a59417a,a59421a,a59422a,a59425a,a59428a,a59429a,a59430a,a59434a,a59435a,a59438a,a59441a,a59442a,a59443a,a59447a,a59448a,a59451a,a59454a,a59455a,a59456a,a59460a,a59461a,a59464a,a59467a,a59468a,a59469a,a59473a,a59474a,a59477a,a59480a,a59481a,a59482a,a59486a,a59487a,a59490a,a59493a,a59494a,a59495a,a59499a,a59500a,a59503a,a59506a,a59507a,a59508a,a59512a,a59513a,a59516a,a59519a,a59520a,a59521a,a59525a,a59526a,a59529a,a59532a,a59533a,a59534a,a59538a,a59539a,a59542a,a59545a,a59546a,a59547a,a59551a,a59552a,a59555a,a59558a,a59559a,a59560a,a59564a,a59565a,a59568a,a59571a,a59572a,a59573a,a59577a,a59578a,a59581a,a59584a,a59585a,a59586a,a59590a,a59591a,a59594a,a59597a,a59598a,a59599a,a59603a,a59604a,a59607a,a59610a,a59611a,a59612a,a59616a,a59617a,a59620a,a59623a,a59624a,a59625a,a59629a,a59630a,a59633a,a59636a,a59637a,a59638a,a59642a,a59643a,a59646a,a59649a,a59650a,a59651a,a59655a,a59656a,a59659a,a59662a,a59663a,a59664a,a59668a,a59669a,a59672a,a59675a,a59676a,a59677a,a59681a,a59682a,a59685a,a59688a,a59689a,a59690a,a59694a,a59695a,a59698a,a59701a,a59702a,a59703a,a59707a,a59708a,a59711a,a59714a,a59715a,a59716a,a59720a,a59721a,a59724a,a59727a,a59728a,a59729a,a59733a,a59734a,a59737a,a59740a,a59741a,a59742a,a59746a,a59747a,a59750a,a59753a,a59754a,a59755a,a59759a,a59760a,a59763a,a59766a,a59767a,a59768a,a59772a,a59773a,a59776a,a59779a,a59780a,a59781a,a59785a,a59786a,a59789a,a59792a,a59793a,a59794a,a59798a,a59799a,a59802a,a59805a,a59806a,a59807a,a59811a,a59812a,a59815a,a59818a,a59819a,a59820a,a59824a,a59825a,a59828a,a59831a,a59832a,a59833a,a59837a,a59838a,a59841a,a59844a,a59845a,a59846a,a59850a,a59851a,a59854a,a59857a,a59858a,a59859a,a59863a,a59864a,a59867a,a59870a,a59871a,a59872a,a59876a,a59877a,a59880a,a59883a,a59884a,a59885a,a59889a,a59890a,a59893a,a59896a,a59897a,a59898a,a59902a,a59903a,a59906a,a59909a,a59910a,a59911a,a59915a,a59916a,a59919a,a59922a,a59923a,a59924a,a59928a,a59929a,a59932a,a59935a,a59936a,a59937a,a59941a,a59942a,a59945a,a59948a,a59949a,a59950a,a59954a,a59955a,a59958a,a59961a,a59962a,a59963a,a59967a,a59968a,a59971a,a59974a,a59975a,a59976a,a59980a,a59981a,a59984a,a59987a,a59988a,a59989a,a59993a,a59994a,a59997a,a60000a,a60001a,a60002a,a60006a,a60007a,a60010a,a60013a,a60014a,a60015a,a60019a,a60020a,a60023a,a60026a,a60027a,a60028a,a60032a,a60033a,a60036a,a60039a,a60040a,a60041a,a60045a,a60046a,a60049a,a60052a,a60053a,a60054a,a60058a,a60059a,a60062a,a60065a,a60066a,a60067a,a60071a,a60072a,a60075a,a60078a,a60079a,a60080a,a60084a,a60085a,a60088a,a60091a,a60092a,a60093a,a60097a,a60098a,a60101a,a60104a,a60105a,a60106a,a60110a,a60111a,a60114a,a60117a,a60118a,a60119a,a60123a,a60124a,a60127a,a60130a,a60131a,a60132a,a60136a,a60137a,a60140a,a60143a,a60144a,a60145a,a60149a,a60150a,a60153a,a60156a,a60157a,a60158a,a60162a,a60163a,a60166a,a60169a,a60170a,a60171a,a60175a,a60176a,a60179a,a60182a,a60183a,a60184a,a60188a,a60189a,a60192a,a60195a,a60196a,a60197a,a60201a,a60202a,a60205a,a60208a,a60209a,a60210a,a60214a,a60215a,a60218a,a60221a,a60222a,a60223a,a60227a,a60228a,a60231a,a60234a,a60235a,a60236a,a60240a,a60241a,a60244a,a60247a,a60248a,a60249a,a60253a,a60254a,a60257a,a60260a,a60261a,a60262a,a60266a,a60267a,a60270a,a60273a,a60274a,a60275a,a60279a,a60280a,a60283a,a60286a,a60287a,a60288a,a60292a,a60293a,a60296a,a60299a,a60300a,a60301a,a60305a,a60306a,a60309a,a60312a,a60313a,a60314a,a60318a,a60319a,a60322a,a60325a,a60326a,a60327a,a60331a,a60332a,a60335a,a60338a,a60339a,a60340a,a60344a,a60345a,a60348a,a60351a,a60352a,a60353a,a60357a,a60358a,a60361a,a60364a,a60365a,a60366a,a60370a,a60371a,a60374a,a60377a,a60378a,a60379a,a60383a,a60384a,a60387a,a60390a,a60391a,a60392a,a60396a,a60397a,a60400a,a60403a,a60404a,a60405a,a60409a,a60410a,a60413a,a60416a,a60417a,a60418a,a60422a,a60423a,a60426a,a60429a,a60430a,a60431a,a60435a,a60436a,a60439a,a60442a,a60443a,a60444a,a60448a,a60449a,a60452a,a60455a,a60456a,a60457a,a60461a,a60462a,a60465a,a60468a,a60469a,a60470a,a60474a,a60475a,a60478a,a60481a,a60482a,a60483a,a60487a,a60488a,a60491a,a60494a,a60495a,a60496a,a60500a,a60501a,a60504a,a60507a,a60508a,a60509a,a60513a,a60514a,a60517a,a60520a,a60521a,a60522a,a60526a,a60527a,a60530a,a60533a,a60534a,a60535a,a60539a,a60540a,a60543a,a60546a,a60547a,a60548a,a60552a,a60553a,a60556a,a60559a,a60560a,a60561a,a60565a,a60566a,a60569a,a60572a,a60573a,a60574a,a60578a,a60579a,a60582a,a60585a,a60586a,a60587a,a60591a,a60592a,a60595a,a60598a,a60599a,a60600a,a60604a,a60605a,a60608a,a60611a,a60612a,a60613a,a60617a,a60618a,a60621a,a60624a,a60625a,a60626a,a60630a,a60631a,a60634a,a60637a,a60638a,a60639a,a60643a,a60644a,a60647a,a60650a,a60651a,a60652a,a60656a,a60657a,a60660a,a60663a,a60664a,a60665a,a60669a,a60670a,a60673a,a60676a,a60677a,a60678a,a60682a,a60683a,a60686a,a60689a,a60690a,a60691a,a60695a,a60696a,a60699a,a60702a,a60703a,a60704a,a60708a,a60709a,a60712a,a60715a,a60716a,a60717a,a60721a,a60722a,a60725a,a60728a,a60729a,a60730a,a60734a,a60735a,a60738a,a60741a,a60742a,a60743a,a60747a,a60748a,a60751a,a60754a,a60755a,a60756a,a60760a,a60761a,a60764a,a60767a,a60768a,a60769a,a60773a,a60774a,a60777a,a60780a,a60781a,a60782a,a60786a,a60787a,a60790a,a60793a,a60794a,a60795a,a60799a,a60800a,a60803a,a60806a,a60807a,a60808a,a60812a,a60813a,a60816a,a60819a,a60820a,a60821a,a60825a,a60826a,a60829a,a60832a,a60833a,a60834a,a60838a,a60839a,a60842a,a60845a,a60846a,a60847a,a60851a,a60852a,a60855a,a60858a,a60859a,a60860a,a60864a,a60865a,a60868a,a60871a,a60872a,a60873a,a60877a,a60878a,a60881a,a60884a,a60885a,a60886a,a60890a,a60891a,a60894a,a60897a,a60898a,a60899a,a60903a,a60904a,a60907a,a60910a,a60911a,a60912a,a60916a,a60917a,a60920a,a60923a,a60924a,a60925a,a60929a,a60930a,a60933a,a60936a,a60937a,a60938a,a60942a,a60943a,a60946a,a60949a,a60950a,a60951a,a60955a,a60956a,a60959a,a60962a,a60963a,a60964a,a60968a,a60969a,a60972a,a60975a,a60976a,a60977a,a60981a,a60982a,a60985a,a60988a,a60989a,a60990a,a60994a,a60995a,a60998a,a61001a,a61002a,a61003a,a61007a,a61008a,a61011a,a61014a,a61015a,a61016a,a61020a,a61021a,a61024a,a61027a,a61028a,a61029a,a61033a,a61034a,a61037a,a61040a,a61041a,a61042a,a61046a,a61047a,a61050a,a61053a,a61054a,a61055a,a61059a,a61060a,a61063a,a61066a,a61067a,a61068a,a61072a,a61073a,a61076a,a61079a,a61080a,a61081a,a61085a,a61086a,a61089a,a61092a,a61093a,a61094a,a61098a,a61099a,a61102a,a61105a,a61106a,a61107a,a61111a,a61112a,a61115a,a61118a,a61119a,a61120a,a61124a,a61125a,a61128a,a61131a,a61132a,a61133a,a61137a,a61138a,a61141a,a61144a,a61145a,a61146a,a61150a,a61151a,a61154a,a61157a,a61158a,a61159a,a61163a,a61164a,a61167a,a61170a,a61171a,a61172a,a61176a,a61177a,a61180a,a61183a,a61184a,a61185a,a61189a,a61190a,a61193a,a61196a,a61197a,a61198a,a61202a,a61203a,a61206a,a61209a,a61210a,a61211a,a61215a,a61216a,a61219a,a61222a,a61223a,a61224a,a61228a,a61229a,a61232a,a61235a,a61236a,a61237a,a61241a,a61242a,a61245a,a61248a,a61249a,a61250a,a61254a,a61255a,a61258a,a61261a,a61262a,a61263a,a61267a,a61268a,a61271a,a61274a,a61275a,a61276a,a61280a,a61281a,a61284a,a61287a,a61288a,a61289a,a61293a,a61294a,a61297a,a61300a,a61301a,a61302a,a61306a,a61307a,a61310a,a61313a,a61314a,a61315a,a61319a,a61320a,a61323a,a61326a,a61327a,a61328a,a61332a,a61333a,a61336a,a61339a,a61340a,a61341a,a61345a,a61346a,a61349a,a61352a,a61353a,a61354a,a61358a,a61359a,a61362a,a61365a,a61366a,a61367a,a61371a,a61372a,a61375a,a61378a,a61379a,a61380a,a61384a,a61385a,a61388a,a61391a,a61392a,a61393a,a61397a,a61398a,a61401a,a61404a,a61405a,a61406a,a61410a,a61411a,a61414a,a61417a,a61418a,a61419a,a61423a,a61424a,a61427a,a61430a,a61431a,a61432a,a61436a,a61437a,a61440a,a61443a,a61444a,a61445a,a61449a,a61450a,a61453a,a61456a,a61457a,a61458a,a61462a,a61463a,a61466a,a61469a,a61470a,a61471a,a61475a,a61476a,a61479a,a61482a,a61483a,a61484a,a61488a,a61489a,a61492a,a61495a,a61496a,a61497a,a61501a,a61502a,a61505a,a61508a,a61509a,a61510a,a61514a,a61515a,a61518a,a61521a,a61522a,a61523a,a61527a,a61528a,a61531a,a61534a,a61535a,a61536a,a61540a,a61541a,a61544a,a61547a,a61548a,a61549a,a61553a,a61554a,a61557a,a61560a,a61561a,a61562a,a61566a,a61567a,a61570a,a61573a,a61574a,a61575a,a61579a,a61580a,a61583a,a61586a,a61587a,a61588a,a61592a,a61593a,a61596a,a61599a,a61600a,a61601a,a61605a,a61606a,a61609a,a61612a,a61613a,a61614a,a61618a,a61619a,a61622a,a61625a,a61626a,a61627a,a61631a,a61632a,a61635a,a61638a,a61639a,a61640a,a61644a,a61645a,a61648a,a61651a,a61652a,a61653a,a61657a,a61658a,a61661a,a61664a,a61665a,a61666a,a61670a,a61671a,a61674a,a61677a,a61678a,a61679a,a61683a,a61684a,a61687a,a61690a,a61691a,a61692a,a61696a,a61697a,a61700a,a61703a,a61704a,a61705a,a61709a,a61710a,a61713a,a61716a,a61717a,a61718a,a61722a,a61723a,a61726a,a61729a,a61730a,a61731a,a61735a,a61736a,a61739a,a61742a,a61743a,a61744a,a61748a,a61749a,a61752a,a61755a,a61756a,a61757a,a61761a,a61762a,a61765a,a61768a,a61769a,a61770a,a61774a,a61775a,a61778a,a61781a,a61782a,a61783a,a61787a,a61788a,a61791a,a61794a,a61795a,a61796a,a61800a,a61801a,a61804a,a61807a,a61808a,a61809a,a61813a,a61814a,a61817a,a61820a,a61821a,a61822a,a61826a,a61827a,a61830a,a61833a,a61834a,a61835a,a61839a,a61840a,a61843a,a61846a,a61847a,a61848a,a61852a,a61853a,a61856a,a61859a,a61860a,a61861a,a61865a,a61866a,a61869a,a61872a,a61873a,a61874a,a61878a,a61879a,a61882a,a61885a,a61886a,a61887a,a61891a,a61892a,a61895a,a61898a,a61899a,a61900a,a61904a,a61905a,a61908a,a61911a,a61912a,a61913a,a61917a,a61918a,a61921a,a61924a,a61925a,a61926a,a61930a,a61931a,a61934a,a61937a,a61938a,a61939a,a61943a,a61944a,a61947a,a61950a,a61951a,a61952a,a61956a,a61957a,a61960a,a61963a,a61964a,a61965a,a61969a,a61970a,a61973a,a61976a,a61977a,a61978a,a61982a,a61983a,a61986a,a61989a,a61990a,a61991a,a61995a,a61996a,a61999a,a62002a,a62003a,a62004a,a62008a,a62009a,a62012a,a62015a,a62016a,a62017a,a62021a,a62022a,a62025a,a62028a,a62029a,a62030a,a62034a,a62035a,a62038a,a62041a,a62042a,a62043a,a62047a,a62048a,a62051a,a62054a,a62055a,a62056a,a62060a,a62061a,a62064a,a62067a,a62068a,a62069a,a62073a,a62074a,a62077a,a62080a,a62081a,a62082a,a62086a,a62087a,a62090a,a62093a,a62094a,a62095a,a62099a,a62100a,a62103a,a62106a,a62107a,a62108a,a62112a,a62113a,a62116a,a62119a,a62120a,a62121a,a62125a,a62126a,a62129a,a62132a,a62133a,a62134a,a62138a,a62139a,a62142a,a62145a,a62146a,a62147a,a62151a,a62152a,a62155a,a62158a,a62159a,a62160a,a62164a,a62165a,a62168a,a62171a,a62172a,a62173a,a62177a,a62178a,a62181a,a62184a,a62185a,a62186a,a62190a,a62191a,a62194a,a62197a,a62198a,a62199a,a62203a,a62204a,a62207a,a62210a,a62211a,a62212a,a62216a,a62217a,a62220a,a62223a,a62224a,a62225a,a62229a,a62230a,a62233a,a62236a,a62237a,a62238a,a62242a,a62243a,a62246a,a62249a,a62250a,a62251a,a62255a,a62256a,a62259a,a62262a,a62263a,a62264a,a62268a,a62269a,a62272a,a62275a,a62276a,a62277a,a62281a,a62282a,a62285a,a62288a,a62289a,a62290a,a62294a,a62295a,a62298a,a62301a,a62302a,a62303a,a62307a,a62308a,a62311a,a62314a,a62315a,a62316a,a62320a,a62321a,a62324a,a62327a,a62328a,a62329a,a62333a,a62334a,a62337a,a62340a,a62341a,a62342a,a62346a,a62347a,a62350a,a62353a,a62354a,a62355a,a62359a,a62360a,a62363a,a62366a,a62367a,a62368a,a62372a,a62373a,a62376a,a62379a,a62380a,a62381a,a62385a,a62386a,a62389a,a62392a,a62393a,a62394a,a62398a,a62399a,a62402a,a62405a,a62406a,a62407a,a62411a,a62412a,a62415a,a62418a,a62419a,a62420a,a62424a,a62425a,a62428a,a62431a,a62432a,a62433a,a62437a,a62438a,a62441a,a62444a,a62445a,a62446a,a62450a,a62451a,a62454a,a62457a,a62458a,a62459a,a62463a,a62464a,a62467a,a62470a,a62471a,a62472a,a62476a,a62477a,a62480a,a62483a,a62484a,a62485a,a62489a,a62490a,a62493a,a62496a,a62497a,a62498a,a62502a,a62503a,a62506a,a62509a,a62510a,a62511a,a62515a,a62516a,a62519a,a62522a,a62523a,a62524a,a62528a,a62529a,a62532a,a62535a,a62536a,a62537a,a62541a,a62542a,a62545a,a62548a,a62549a,a62550a,a62554a,a62555a,a62558a,a62561a,a62562a,a62563a,a62567a,a62568a,a62571a,a62574a,a62575a,a62576a,a62580a,a62581a,a62584a,a62587a,a62588a,a62589a,a62593a,a62594a,a62597a,a62600a,a62601a,a62602a,a62606a,a62607a,a62610a,a62613a,a62614a,a62615a,a62619a,a62620a,a62623a,a62626a,a62627a,a62628a,a62632a,a62633a,a62636a,a62639a,a62640a,a62641a,a62645a,a62646a,a62649a,a62652a,a62653a,a62654a,a62658a,a62659a,a62662a,a62665a,a62666a,a62667a,a62671a,a62672a,a62675a,a62678a,a62679a,a62680a,a62684a,a62685a,a62688a,a62691a,a62692a,a62693a,a62697a,a62698a,a62701a,a62704a,a62705a,a62706a,a62710a,a62711a,a62714a,a62717a,a62718a,a62719a,a62723a,a62724a,a62727a,a62730a,a62731a,a62732a,a62736a,a62737a,a62740a,a62743a,a62744a,a62745a,a62749a,a62750a,a62753a,a62756a,a62757a,a62758a,a62762a,a62763a,a62766a,a62769a,a62770a,a62771a,a62775a,a62776a,a62779a,a62782a,a62783a,a62784a,a62788a,a62789a,a62792a,a62795a,a62796a,a62797a,a62801a,a62802a,a62805a,a62808a,a62809a,a62810a,a62814a,a62815a,a62818a,a62821a,a62822a,a62823a,a62827a,a62828a,a62831a,a62834a,a62835a,a62836a,a62840a,a62841a,a62844a,a62847a,a62848a,a62849a,a62853a,a62854a,a62857a,a62860a,a62861a,a62862a,a62866a,a62867a,a62870a,a62873a,a62874a,a62875a,a62879a,a62880a,a62883a,a62886a,a62887a,a62888a,a62892a,a62893a,a62896a,a62899a,a62900a,a62901a,a62905a,a62906a,a62909a,a62912a,a62913a,a62914a,a62918a,a62919a,a62922a,a62925a,a62926a,a62927a,a62931a,a62932a,a62935a,a62938a,a62939a,a62940a,a62944a,a62945a,a62948a,a62951a,a62952a,a62953a,a62957a,a62958a,a62961a,a62964a,a62965a,a62966a,a62970a,a62971a,a62974a,a62977a,a62978a,a62979a,a62983a,a62984a,a62987a,a62990a,a62991a,a62992a,a62996a,a62997a,a63000a,a63003a,a63004a,a63005a,a63009a,a63010a,a63013a,a63016a,a63017a,a63018a,a63022a,a63023a,a63026a,a63029a,a63030a,a63031a,a63035a,a63036a,a63039a,a63042a,a63043a,a63044a,a63048a,a63049a,a63052a,a63055a,a63056a,a63057a,a63061a,a63062a,a63065a,a63068a,a63069a,a63070a,a63074a,a63075a,a63078a,a63081a,a63082a,a63083a,a63087a,a63088a,a63091a,a63094a,a63095a,a63096a,a63100a,a63101a,a63104a,a63107a,a63108a,a63109a,a63113a,a63114a,a63117a,a63120a,a63121a,a63122a,a63126a,a63127a,a63130a,a63133a,a63134a,a63135a,a63139a,a63140a,a63143a,a63146a,a63147a,a63148a,a63152a,a63153a,a63156a,a63159a,a63160a,a63161a,a63165a,a63166a,a63169a,a63172a,a63173a,a63174a,a63178a,a63179a,a63182a,a63185a,a63186a,a63187a,a63191a,a63192a,a63195a,a63198a,a63199a,a63200a,a63204a,a63205a,a63208a,a63211a,a63212a,a63213a,a63217a,a63218a,a63221a,a63224a,a63225a,a63226a,a63230a,a63231a,a63234a,a63237a,a63238a,a63239a,a63243a,a63244a,a63247a,a63250a,a63251a,a63252a,a63256a,a63257a,a63260a,a63263a,a63264a,a63265a,a63269a,a63270a,a63273a,a63276a,a63277a,a63278a,a63282a,a63283a,a63286a,a63289a,a63290a,a63291a,a63295a,a63296a,a63299a,a63302a,a63303a,a63304a,a63308a,a63309a,a63312a,a63315a,a63316a,a63317a,a63321a,a63322a,a63325a,a63328a,a63329a,a63330a,a63334a,a63335a,a63338a,a63341a,a63342a,a63343a,a63347a,a63348a,a63351a,a63354a,a63355a,a63356a,a63360a,a63361a,a63364a,a63367a,a63368a,a63369a,a63373a,a63374a,a63377a,a63380a,a63381a,a63382a,a63386a,a63387a,a63390a,a63393a,a63394a,a63395a,a63399a,a63400a,a63403a,a63406a,a63407a,a63408a,a63412a,a63413a,a63416a,a63419a,a63420a,a63421a,a63425a,a63426a,a63429a,a63432a,a63433a,a63434a,a63438a,a63439a,a63442a,a63445a,a63446a,a63447a,a63451a,a63452a,a63455a,a63458a,a63459a,a63460a,a63464a,a63465a,a63468a,a63471a,a63472a,a63473a,a63477a,a63478a,a63481a,a63484a,a63485a,a63486a,a63490a,a63491a,a63494a,a63497a,a63498a,a63499a,a63503a,a63504a,a63507a,a63510a,a63511a,a63512a,a63516a,a63517a,a63520a,a63523a,a63524a,a63525a,a63529a,a63530a,a63533a,a63536a,a63537a,a63538a,a63542a,a63543a,a63546a,a63549a,a63550a,a63551a,a63555a,a63556a,a63559a,a63562a,a63563a,a63564a,a63568a,a63569a,a63572a,a63575a,a63576a,a63577a,a63581a,a63582a,a63585a,a63588a,a63589a,a63590a,a63594a,a63595a,a63598a,a63601a,a63602a,a63603a,a63607a,a63608a,a63611a,a63614a,a63615a,a63616a,a63620a,a63621a,a63624a,a63627a,a63628a,a63629a,a63633a,a63634a,a63637a,a63640a,a63641a,a63642a,a63646a,a63647a,a63650a,a63653a,a63654a,a63655a,a63659a,a63660a,a63663a,a63666a,a63667a,a63668a,a63672a,a63673a,a63676a,a63679a,a63680a,a63681a,a63685a,a63686a,a63689a,a63692a,a63693a,a63694a,a63698a,a63699a,a63702a,a63705a,a63706a,a63707a,a63711a,a63712a,a63715a,a63718a,a63719a,a63720a,a63724a,a63725a,a63728a,a63731a,a63732a,a63733a,a63737a,a63738a,a63741a,a63744a,a63745a,a63746a,a63750a,a63751a,a63754a,a63757a,a63758a,a63759a,a63763a,a63764a,a63767a,a63770a,a63771a,a63772a,a63776a,a63777a,a63780a,a63783a,a63784a,a63785a,a63789a,a63790a,a63793a,a63796a,a63797a,a63798a,a63802a,a63803a,a63806a,a63809a,a63810a,a63811a,a63815a,a63816a,a63819a,a63822a,a63823a,a63824a,a63828a,a63829a,a63832a,a63835a,a63836a,a63837a,a63841a,a63842a,a63845a,a63848a,a63849a,a63850a,a63854a,a63855a,a63858a,a63861a,a63862a,a63863a,a63867a,a63868a,a63871a,a63874a,a63875a,a63876a,a63880a,a63881a,a63884a,a63887a,a63888a,a63889a,a63893a,a63894a,a63897a,a63900a,a63901a,a63902a,a63906a,a63907a,a63910a,a63913a,a63914a,a63915a,a63919a,a63920a,a63923a,a63926a,a63927a,a63928a,a63932a,a63933a,a63936a,a63939a,a63940a,a63941a,a63945a,a63946a,a63949a,a63952a,a63953a,a63954a,a63958a,a63959a,a63962a,a63965a,a63966a,a63967a,a63971a,a63972a,a63975a,a63978a,a63979a,a63980a,a63984a,a63985a,a63988a,a63991a,a63992a,a63993a,a63997a,a63998a,a64001a,a64004a,a64005a,a64006a,a64010a,a64011a,a64014a,a64017a,a64018a,a64019a,a64023a,a64024a,a64027a,a64030a,a64031a,a64032a,a64036a,a64037a,a64040a,a64043a,a64044a,a64045a,a64049a,a64050a,a64053a,a64056a,a64057a,a64058a,a64062a,a64063a,a64066a,a64069a,a64070a,a64071a,a64075a,a64076a,a64079a,a64082a,a64083a,a64084a,a64088a,a64089a,a64092a,a64095a,a64096a,a64097a,a64101a,a64102a,a64105a,a64108a,a64109a,a64110a,a64114a,a64115a,a64118a,a64121a,a64122a,a64123a,a64127a,a64128a,a64131a,a64134a,a64135a,a64136a,a64140a,a64141a,a64144a,a64147a,a64148a,a64149a,a64153a,a64154a,a64157a,a64160a,a64161a,a64162a,a64166a,a64167a,a64170a,a64173a,a64174a,a64175a,a64179a,a64180a,a64183a,a64186a,a64187a,a64188a,a64192a,a64193a,a64196a,a64199a,a64200a,a64201a,a64205a,a64206a,a64209a,a64212a,a64213a,a64214a,a64218a,a64219a,a64222a,a64225a,a64226a,a64227a,a64231a,a64232a,a64235a,a64238a,a64239a,a64240a,a64244a,a64245a,a64248a,a64251a,a64252a,a64253a,a64257a,a64258a,a64261a,a64264a,a64265a,a64266a,a64270a,a64271a,a64274a,a64277a,a64278a,a64279a,a64283a,a64284a,a64287a,a64290a,a64291a,a64292a,a64296a,a64297a,a64300a,a64303a,a64304a,a64305a,a64309a,a64310a,a64313a,a64316a,a64317a,a64318a,a64322a,a64323a,a64326a,a64329a,a64330a,a64331a,a64335a,a64336a,a64339a,a64342a,a64343a,a64344a,a64348a,a64349a,a64352a,a64355a,a64356a,a64357a,a64361a,a64362a,a64365a,a64368a,a64369a,a64370a,a64374a,a64375a,a64378a,a64381a,a64382a,a64383a,a64387a,a64388a,a64391a,a64394a,a64395a,a64396a,a64400a,a64401a,a64404a,a64407a,a64408a,a64409a,a64413a,a64414a,a64417a,a64420a,a64421a,a64422a,a64426a,a64427a,a64430a,a64433a,a64434a,a64435a,a64439a,a64440a,a64443a,a64446a,a64447a,a64448a,a64452a,a64453a,a64456a,a64459a,a64460a,a64461a,a64465a,a64466a,a64469a,a64472a,a64473a,a64474a,a64478a,a64479a,a64482a,a64485a,a64486a,a64487a,a64491a,a64492a,a64495a,a64498a,a64499a,a64500a,a64504a,a64505a,a64508a,a64511a,a64512a,a64513a,a64517a,a64518a,a64521a,a64524a,a64525a,a64526a,a64530a,a64531a,a64534a,a64537a,a64538a,a64539a,a64543a,a64544a,a64547a,a64550a,a64551a,a64552a,a64556a,a64557a,a64560a,a64563a,a64564a,a64565a,a64569a,a64570a,a64573a,a64576a,a64577a,a64578a,a64582a,a64583a,a64586a,a64589a,a64590a,a64591a,a64595a,a64596a,a64599a,a64602a,a64603a,a64604a,a64608a,a64609a,a64612a,a64615a,a64616a,a64617a,a64621a,a64622a,a64625a,a64628a,a64629a,a64630a,a64634a,a64635a,a64638a,a64641a,a64642a,a64643a,a64647a,a64648a,a64651a,a64654a,a64655a,a64656a,a64660a,a64661a,a64664a,a64667a,a64668a,a64669a,a64673a,a64674a,a64677a,a64680a,a64681a,a64682a,a64686a,a64687a,a64690a,a64693a,a64694a,a64695a,a64699a,a64700a,a64703a,a64706a,a64707a,a64708a,a64712a,a64713a,a64716a,a64719a,a64720a,a64721a,a64725a,a64726a,a64729a,a64732a,a64733a,a64734a,a64738a,a64739a,a64742a,a64745a,a64746a,a64747a,a64751a,a64752a,a64755a,a64758a,a64759a,a64760a,a64764a,a64765a,a64768a,a64771a,a64772a,a64773a,a64777a,a64778a,a64781a,a64784a,a64785a,a64786a,a64790a,a64791a,a64794a,a64797a,a64798a,a64799a,a64803a,a64804a,a64807a,a64810a,a64811a,a64812a,a64816a,a64817a,a64820a,a64823a,a64824a,a64825a,a64829a,a64830a,a64833a,a64836a,a64837a,a64838a,a64842a,a64843a,a64846a,a64849a,a64850a,a64851a,a64855a,a64856a,a64859a,a64862a,a64863a,a64864a,a64868a,a64869a,a64872a,a64875a,a64876a,a64877a,a64881a,a64882a,a64885a,a64888a,a64889a,a64890a,a64894a,a64895a,a64898a,a64901a,a64902a,a64903a,a64907a,a64908a,a64911a,a64914a,a64915a,a64916a,a64920a,a64921a,a64924a,a64927a,a64928a,a64929a,a64933a,a64934a,a64937a,a64940a,a64941a,a64942a,a64946a,a64947a,a64950a,a64953a,a64954a,a64955a,a64959a,a64960a,a64963a,a64966a,a64967a,a64968a,a64972a,a64973a,a64976a,a64979a,a64980a,a64981a,a64985a,a64986a,a64989a,a64992a,a64993a,a64994a,a64998a,a64999a,a65002a,a65005a,a65006a,a65007a,a65011a,a65012a,a65015a,a65018a,a65019a,a65020a,a65024a,a65025a,a65028a,a65031a,a65032a,a65033a,a65037a,a65038a,a65041a,a65044a,a65045a,a65046a,a65050a,a65051a,a65054a,a65057a,a65058a,a65059a,a65063a,a65064a,a65067a,a65070a,a65071a,a65072a,a65076a,a65077a,a65080a,a65083a,a65084a,a65085a,a65089a,a65090a,a65093a,a65096a,a65097a,a65098a,a65102a,a65103a,a65106a,a65109a,a65110a,a65111a,a65115a,a65116a,a65119a,a65122a,a65123a,a65124a,a65128a,a65129a,a65132a,a65135a,a65136a,a65137a,a65141a,a65142a,a65145a,a65148a,a65149a,a65150a,a65154a,a65155a,a65158a,a65161a,a65162a,a65163a,a65167a,a65168a,a65171a,a65174a,a65175a,a65176a,a65180a,a65181a,a65184a,a65187a,a65188a,a65189a,a65193a,a65194a,a65197a,a65200a,a65201a,a65202a,a65206a,a65207a,a65210a,a65213a,a65214a,a65215a,a65219a,a65220a,a65223a,a65226a,a65227a,a65228a,a65232a,a65233a,a65236a,a65239a,a65240a,a65241a,a65245a,a65246a,a65249a,a65252a,a65253a,a65254a,a65258a,a65259a,a65262a,a65265a,a65266a,a65267a,a65271a,a65272a,a65275a,a65278a,a65279a,a65280a,a65284a,a65285a,a65288a,a65291a,a65292a,a65293a,a65297a,a65298a,a65301a,a65304a,a65305a,a65306a,a65310a,a65311a,a65314a,a65317a,a65318a,a65319a,a65323a,a65324a,a65327a,a65330a,a65331a,a65332a,a65336a,a65337a,a65340a,a65343a,a65344a,a65345a,a65349a,a65350a,a65353a,a65356a,a65357a,a65358a,a65362a,a65363a,a65366a,a65369a,a65370a,a65371a,a65375a,a65376a,a65379a,a65382a,a65383a,a65384a,a65388a,a65389a,a65392a,a65395a,a65396a,a65397a,a65401a,a65402a,a65405a,a65408a,a65409a,a65410a,a65414a,a65415a,a65418a,a65421a,a65422a,a65423a,a65427a,a65428a,a65431a,a65434a,a65435a,a65436a,a65440a,a65441a,a65444a,a65447a,a65448a,a65449a,a65453a,a65454a,a65457a,a65460a,a65461a,a65462a,a65466a,a65467a,a65470a,a65473a,a65474a,a65475a,a65479a,a65480a,a65483a,a65486a,a65487a,a65488a,a65492a,a65493a,a65496a,a65499a,a65500a,a65501a,a65505a,a65506a,a65509a,a65512a,a65513a,a65514a,a65518a,a65519a,a65522a,a65525a,a65526a,a65527a,a65531a,a65532a,a65535a,a65538a,a65539a,a65540a,a65544a,a65545a,a65548a,a65551a,a65552a,a65553a,a65557a,a65558a,a65561a,a65564a,a65565a,a65566a,a65570a,a65571a,a65574a,a65577a,a65578a,a65579a,a65583a,a65584a,a65587a,a65590a,a65591a,a65592a,a65596a,a65597a,a65600a,a65603a,a65604a,a65605a,a65609a,a65610a,a65613a,a65616a,a65617a,a65618a,a65622a,a65623a,a65626a,a65629a,a65630a,a65631a,a65635a,a65636a,a65639a,a65642a,a65643a,a65644a,a65648a,a65649a,a65652a,a65655a,a65656a,a65657a,a65661a,a65662a,a65665a,a65668a,a65669a,a65670a,a65674a,a65675a,a65678a,a65681a,a65682a,a65683a,a65687a,a65688a,a65691a,a65694a,a65695a,a65696a,a65700a,a65701a,a65704a,a65707a,a65708a,a65709a,a65713a,a65714a,a65717a,a65720a,a65721a,a65722a,a65726a,a65727a,a65730a,a65733a,a65734a,a65735a,a65739a,a65740a,a65743a,a65746a,a65747a,a65748a,a65752a,a65753a,a65756a,a65759a,a65760a,a65761a,a65765a,a65766a,a65769a,a65772a,a65773a,a65774a,a65778a,a65779a,a65782a,a65785a,a65786a,a65787a,a65791a,a65792a,a65795a,a65798a,a65799a,a65800a,a65804a,a65805a,a65808a,a65811a,a65812a,a65813a,a65817a,a65818a,a65821a,a65824a,a65825a,a65826a,a65830a,a65831a,a65834a,a65837a,a65838a,a65839a,a65843a,a65844a,a65847a,a65850a,a65851a,a65852a,a65856a,a65857a,a65860a,a65863a,a65864a,a65865a,a65869a,a65870a,a65873a,a65876a,a65877a,a65878a,a65882a,a65883a,a65886a,a65889a,a65890a,a65891a,a65895a,a65896a,a65899a,a65902a,a65903a,a65904a,a65908a,a65909a,a65912a,a65915a,a65916a,a65917a,a65921a,a65922a,a65925a,a65928a,a65929a,a65930a,a65934a,a65935a,a65938a,a65941a,a65942a,a65943a,a65947a,a65948a,a65951a,a65954a,a65955a,a65956a,a65960a,a65961a,a65964a,a65967a,a65968a,a65969a,a65973a,a65974a,a65977a,a65980a,a65981a,a65982a,a65986a,a65987a,a65990a,a65993a,a65994a,a65995a,a65999a,a66000a,a66003a,a66006a,a66007a,a66008a,a66012a,a66013a,a66016a,a66019a,a66020a,a66021a,a66025a,a66026a,a66029a,a66032a,a66033a,a66034a,a66038a,a66039a,a66042a,a66045a,a66046a,a66047a,a66051a,a66052a,a66055a,a66058a,a66059a,a66060a,a66064a,a66065a,a66068a,a66071a,a66072a,a66073a,a66077a,a66078a,a66081a,a66084a,a66085a,a66086a,a66090a,a66091a,a66094a,a66097a,a66098a,a66099a,a66103a,a66104a,a66107a,a66110a,a66111a,a66112a,a66116a,a66117a,a66120a,a66123a,a66124a,a66125a,a66129a,a66130a,a66133a,a66136a,a66137a,a66138a,a66142a,a66143a,a66146a,a66149a,a66150a,a66151a,a66155a,a66156a,a66159a,a66162a,a66163a,a66164a,a66168a,a66169a,a66172a,a66175a,a66176a,a66177a,a66181a,a66182a,a66185a,a66188a,a66189a,a66190a,a66194a,a66195a,a66198a,a66201a,a66202a,a66203a,a66207a,a66208a,a66211a,a66214a,a66215a,a66216a,a66220a,a66221a,a66224a,a66227a,a66228a,a66229a,a66233a,a66234a,a66237a,a66240a,a66241a,a66242a,a66246a,a66247a,a66250a,a66253a,a66254a,a66255a,a66259a,a66260a,a66263a,a66266a,a66267a,a66268a,a66272a,a66273a,a66276a,a66279a,a66280a,a66281a,a66285a,a66286a,a66289a,a66292a,a66293a,a66294a,a66298a,a66299a,a66302a,a66305a,a66306a,a66307a,a66311a,a66312a,a66315a,a66318a,a66319a,a66320a,a66324a,a66325a,a66328a,a66331a,a66332a,a66333a,a66337a,a66338a,a66341a,a66344a,a66345a,a66346a,a66350a,a66351a,a66354a,a66357a,a66358a,a66359a,a66363a,a66364a,a66367a,a66370a,a66371a,a66372a,a66376a,a66377a,a66380a,a66383a,a66384a,a66385a,a66389a,a66390a,a66393a,a66396a,a66397a,a66398a,a66402a,a66403a,a66406a,a66409a,a66410a,a66411a,a66415a,a66416a,a66419a,a66422a,a66423a,a66424a,a66428a,a66429a,a66432a,a66435a,a66436a,a66437a,a66441a,a66442a,a66445a,a66448a,a66449a,a66450a,a66454a,a66455a,a66458a,a66461a,a66462a,a66463a,a66467a,a66468a,a66471a,a66474a,a66475a,a66476a,a66480a,a66481a,a66484a,a66487a,a66488a,a66489a,a66493a,a66494a,a66497a,a66500a,a66501a,a66502a,a66506a,a66507a,a66510a,a66513a,a66514a,a66515a,a66519a,a66520a,a66523a,a66526a,a66527a,a66528a,a66532a,a66533a,a66536a,a66539a,a66540a,a66541a,a66545a,a66546a,a66549a,a66552a,a66553a,a66554a,a66558a,a66559a,a66562a,a66565a,a66566a,a66567a,a66571a,a66572a,a66575a,a66578a,a66579a,a66580a,a66584a,a66585a,a66588a,a66591a,a66592a,a66593a,a66597a,a66598a,a66601a,a66604a,a66605a,a66606a,a66610a,a66611a,a66614a,a66617a,a66618a,a66619a,a66623a,a66624a,a66627a,a66630a,a66631a,a66632a,a66636a,a66637a,a66640a,a66643a,a66644a,a66645a,a66649a,a66650a,a66653a,a66656a,a66657a,a66658a,a66662a,a66663a,a66666a,a66669a,a66670a,a66671a,a66675a,a66676a,a66679a,a66682a,a66683a,a66684a,a66688a,a66689a,a66692a,a66695a,a66696a,a66697a,a66701a,a66702a,a66705a,a66708a,a66709a,a66710a,a66714a,a66715a,a66718a,a66721a,a66722a,a66723a,a66727a,a66728a,a66731a,a66734a,a66735a,a66736a,a66740a,a66741a,a66744a,a66747a,a66748a,a66749a,a66753a,a66754a,a66757a,a66760a,a66761a,a66762a,a66766a,a66767a,a66770a,a66773a,a66774a,a66775a,a66779a,a66780a,a66783a,a66786a,a66787a,a66788a,a66792a,a66793a,a66796a,a66799a,a66800a,a66801a,a66805a,a66806a,a66809a,a66812a,a66813a,a66814a,a66818a,a66819a,a66822a,a66825a,a66826a,a66827a,a66831a,a66832a,a66835a,a66838a,a66839a,a66840a,a66844a,a66845a,a66848a,a66851a,a66852a,a66853a,a66857a,a66858a,a66861a,a66864a,a66865a,a66866a,a66870a,a66871a,a66874a,a66877a,a66878a,a66879a,a66883a,a66884a,a66887a,a66890a,a66891a,a66892a,a66896a,a66897a,a66900a,a66903a,a66904a,a66905a,a66909a,a66910a,a66913a,a66916a,a66917a,a66918a,a66922a,a66923a,a66926a,a66929a,a66930a,a66931a,a66935a,a66936a,a66939a,a66942a,a66943a,a66944a,a66948a,a66949a,a66952a,a66955a,a66956a,a66957a,a66961a,a66962a,a66965a,a66968a,a66969a,a66970a,a66974a,a66975a,a66978a,a66981a,a66982a,a66983a,a66987a,a66988a,a66991a,a66994a,a66995a,a66996a,a67000a,a67001a,a67004a,a67007a,a67008a,a67009a,a67013a,a67014a,a67017a,a67020a,a67021a,a67022a,a67026a,a67027a,a67030a,a67033a,a67034a,a67035a,a67039a,a67040a,a67043a,a67046a,a67047a,a67048a,a67052a,a67053a,a67056a,a67059a,a67060a,a67061a,a67065a,a67066a,a67069a,a67072a,a67073a,a67074a,a67078a,a67079a,a67082a,a67085a,a67086a,a67087a,a67091a,a67092a,a67095a,a67098a,a67099a,a67100a,a67104a,a67105a,a67108a,a67111a,a67112a,a67113a,a67117a,a67118a,a67121a,a67124a,a67125a,a67126a,a67130a,a67131a,a67134a,a67137a,a67138a,a67139a,a67143a,a67144a,a67147a,a67150a,a67151a,a67152a,a67156a,a67157a,a67160a,a67163a,a67164a,a67165a,a67169a,a67170a,a67173a,a67176a,a67177a,a67178a,a67182a,a67183a,a67186a,a67189a,a67190a,a67191a,a67195a,a67196a,a67199a,a67202a,a67203a,a67204a,a67208a,a67209a,a67212a,a67215a,a67216a,a67217a,a67221a,a67222a,a67225a,a67228a,a67229a,a67230a,a67234a,a67235a,a67238a,a67241a,a67242a,a67243a,a67247a,a67248a,a67251a,a67254a,a67255a,a67256a,a67260a,a67261a,a67264a,a67267a,a67268a,a67269a,a67273a,a67274a,a67277a,a67280a,a67281a,a67282a,a67286a,a67287a,a67290a,a67293a,a67294a,a67295a,a67299a,a67300a,a67303a,a67306a,a67307a,a67308a,a67312a,a67313a,a67316a,a67319a,a67320a,a67321a,a67325a,a67326a,a67329a,a67332a,a67333a,a67334a,a67338a,a67339a,a67342a,a67345a,a67346a,a67347a,a67351a,a67352a,a67355a,a67358a,a67359a,a67360a,a67364a,a67365a,a67368a,a67371a,a67372a,a67373a,a67377a,a67378a,a67381a,a67384a,a67385a,a67386a,a67390a,a67391a,a67394a,a67397a,a67398a,a67399a,a67403a,a67404a,a67407a,a67410a,a67411a,a67412a,a67416a,a67417a,a67420a,a67423a,a67424a,a67425a,a67429a,a67430a,a67433a,a67436a,a67437a,a67438a,a67442a,a67443a,a67446a,a67449a,a67450a,a67451a,a67455a,a67456a,a67459a,a67462a,a67463a,a67464a,a67468a,a67469a,a67472a,a67475a,a67476a,a67477a,a67481a,a67482a,a67485a,a67488a,a67489a,a67490a,a67494a,a67495a,a67498a,a67501a,a67502a,a67503a,a67507a,a67508a,a67511a,a67514a,a67515a,a67516a,a67520a,a67521a,a67524a,a67527a,a67528a,a67529a,a67533a,a67534a,a67537a,a67540a,a67541a,a67542a,a67546a,a67547a,a67550a,a67553a,a67554a,a67555a,a67559a,a67560a,a67563a,a67566a,a67567a,a67568a,a67572a,a67573a,a67576a,a67579a,a67580a,a67581a,a67585a,a67586a,a67589a,a67592a,a67593a,a67594a,a67598a,a67599a,a67602a,a67605a,a67606a,a67607a,a67611a,a67612a,a67615a,a67618a,a67619a,a67620a,a67624a,a67625a,a67628a,a67631a,a67632a,a67633a,a67637a,a67638a,a67641a,a67644a,a67645a,a67646a,a67650a,a67651a,a67654a,a67657a,a67658a,a67659a,a67663a,a67664a,a67667a,a67670a,a67671a,a67672a,a67676a,a67677a,a67680a,a67683a,a67684a,a67685a,a67689a,a67690a,a67693a,a67696a,a67697a,a67698a,a67702a,a67703a,a67706a,a67709a,a67710a,a67711a,a67715a,a67716a,a67719a,a67722a,a67723a,a67724a,a67728a,a67729a,a67732a,a67735a,a67736a,a67737a,a67741a,a67742a,a67745a,a67748a,a67749a,a67750a,a67754a,a67755a,a67758a,a67761a,a67762a,a67763a,a67767a,a67768a,a67771a,a67774a,a67775a,a67776a,a67780a,a67781a,a67784a,a67787a,a67788a,a67789a,a67793a,a67794a,a67797a,a67800a,a67801a,a67802a,a67806a,a67807a,a67810a,a67813a,a67814a,a67815a,a67819a,a67820a,a67823a,a67826a,a67827a,a67828a,a67832a,a67833a,a67836a,a67839a,a67840a,a67841a,a67845a,a67846a,a67849a,a67852a,a67853a,a67854a,a67858a,a67859a,a67862a,a67865a,a67866a,a67867a,a67871a,a67872a,a67875a,a67878a,a67879a,a67880a,a67884a,a67885a,a67888a,a67891a,a67892a,a67893a,a67897a,a67898a,a67901a,a67904a,a67905a,a67906a,a67910a,a67911a,a67914a,a67917a,a67918a,a67919a,a67923a,a67924a,a67927a,a67930a,a67931a,a67932a,a67936a,a67937a,a67940a,a67943a,a67944a,a67945a,a67949a,a67950a,a67953a,a67956a,a67957a,a67958a,a67962a,a67963a,a67966a,a67969a,a67970a,a67971a,a67975a,a67976a,a67979a,a67982a,a67983a,a67984a,a67988a,a67989a,a67992a,a67995a,a67996a,a67997a,a68001a,a68002a,a68005a,a68008a,a68009a,a68010a,a68014a,a68015a,a68018a,a68021a,a68022a,a68023a,a68027a,a68028a,a68031a,a68034a,a68035a,a68036a,a68040a,a68041a,a68044a,a68047a,a68048a,a68049a,a68053a,a68054a,a68057a,a68060a,a68061a,a68062a,a68066a,a68067a,a68070a,a68073a,a68074a,a68075a,a68079a,a68080a,a68083a,a68086a,a68087a,a68088a,a68092a,a68093a,a68096a,a68099a,a68100a,a68101a,a68105a,a68106a,a68109a,a68112a,a68113a,a68114a,a68118a,a68119a,a68122a,a68125a,a68126a,a68127a,a68131a,a68132a,a68135a,a68138a,a68139a,a68140a,a68144a,a68145a,a68148a,a68151a,a68152a,a68153a,a68157a,a68158a,a68161a,a68164a,a68165a,a68166a,a68170a,a68171a,a68174a,a68177a,a68178a,a68179a,a68183a,a68184a,a68187a,a68190a,a68191a,a68192a,a68196a,a68197a,a68200a,a68203a,a68204a,a68205a,a68209a,a68210a,a68213a,a68216a,a68217a,a68218a,a68222a,a68223a,a68226a,a68229a,a68230a,a68231a,a68235a,a68236a,a68239a,a68242a,a68243a,a68244a,a68248a,a68249a,a68252a,a68255a,a68256a,a68257a,a68261a,a68262a,a68265a,a68268a,a68269a,a68270a,a68274a,a68275a,a68278a,a68281a,a68282a,a68283a,a68287a,a68288a,a68291a,a68294a,a68295a,a68296a,a68300a,a68301a,a68304a,a68307a,a68308a,a68309a,a68313a,a68314a,a68317a,a68320a,a68321a,a68322a,a68326a,a68327a,a68330a,a68333a,a68334a,a68335a,a68339a,a68340a,a68343a,a68346a,a68347a,a68348a,a68352a,a68353a,a68356a,a68359a,a68360a,a68361a,a68365a,a68366a,a68369a,a68372a,a68373a,a68374a,a68378a,a68379a,a68382a,a68385a,a68386a,a68387a,a68391a,a68392a,a68395a,a68398a,a68399a,a68400a,a68404a,a68405a,a68408a,a68411a,a68412a,a68413a,a68417a,a68418a,a68421a,a68424a,a68425a,a68426a,a68430a,a68431a,a68434a,a68437a,a68438a,a68439a,a68443a,a68444a,a68447a,a68450a,a68451a,a68452a,a68456a,a68457a,a68460a,a68463a,a68464a,a68465a,a68469a,a68470a,a68473a,a68476a,a68477a,a68478a,a68482a,a68483a,a68486a,a68489a,a68490a,a68491a,a68495a,a68496a,a68499a,a68502a,a68503a,a68504a,a68508a,a68509a,a68512a,a68515a,a68516a,a68517a,a68521a,a68522a,a68525a,a68528a,a68529a,a68530a,a68534a,a68535a,a68538a,a68541a,a68542a,a68543a,a68547a,a68548a,a68551a,a68554a,a68555a,a68556a,a68560a,a68561a,a68564a,a68567a,a68568a,a68569a,a68573a,a68574a,a68577a,a68580a,a68581a,a68582a,a68586a,a68587a,a68590a,a68593a,a68594a,a68595a,a68599a,a68600a,a68603a,a68606a,a68607a,a68608a,a68612a,a68613a,a68616a,a68619a,a68620a,a68621a,a68625a,a68626a,a68629a,a68632a,a68633a,a68634a,a68638a,a68639a,a68642a,a68645a,a68646a,a68647a,a68651a,a68652a,a68655a,a68658a,a68659a,a68660a,a68664a,a68665a,a68668a,a68671a,a68672a,a68673a,a68677a,a68678a,a68681a,a68684a,a68685a,a68686a,a68690a,a68691a,a68694a,a68697a,a68698a,a68699a,a68703a,a68704a,a68707a,a68710a,a68711a,a68712a,a68716a,a68717a,a68720a,a68723a,a68724a,a68725a,a68729a,a68730a,a68733a,a68736a,a68737a,a68738a,a68742a,a68743a,a68746a,a68749a,a68750a,a68751a,a68755a,a68756a,a68759a,a68762a,a68763a,a68764a,a68768a,a68769a,a68772a,a68775a,a68776a,a68777a,a68781a,a68782a,a68785a,a68788a,a68789a,a68790a,a68794a,a68795a,a68798a,a68801a,a68802a,a68803a,a68807a,a68808a,a68811a,a68814a,a68815a,a68816a,a68820a,a68821a,a68824a,a68827a,a68828a,a68829a,a68833a,a68834a,a68837a,a68840a,a68841a,a68842a,a68846a,a68847a,a68850a,a68853a,a68854a,a68855a,a68859a,a68860a,a68863a,a68866a,a68867a,a68868a,a68872a,a68873a,a68876a,a68879a,a68880a,a68881a,a68885a,a68886a,a68889a,a68892a,a68893a,a68894a,a68898a,a68899a,a68902a,a68905a,a68906a,a68907a,a68911a,a68912a,a68915a,a68918a,a68919a,a68920a,a68924a,a68925a,a68928a,a68931a,a68932a,a68933a,a68937a,a68938a,a68941a,a68944a,a68945a,a68946a,a68950a,a68951a,a68954a,a68957a,a68958a,a68959a,a68963a,a68964a,a68967a,a68970a,a68971a,a68972a,a68976a,a68977a,a68980a,a68983a,a68984a,a68985a,a68989a,a68990a,a68993a,a68996a,a68997a,a68998a,a69002a,a69003a,a69006a,a69009a,a69010a,a69011a,a69015a,a69016a,a69019a,a69022a,a69023a,a69024a,a69028a,a69029a,a69032a,a69035a,a69036a,a69037a,a69041a,a69042a,a69045a,a69048a,a69049a,a69050a,a69054a,a69055a,a69058a,a69061a,a69062a,a69063a,a69067a,a69068a,a69071a,a69074a,a69075a,a69076a,a69080a,a69081a,a69084a,a69087a,a69088a,a69089a,a69093a,a69094a,a69097a,a69100a,a69101a,a69102a,a69106a,a69107a,a69110a,a69113a,a69114a,a69115a,a69119a,a69120a,a69123a,a69126a,a69127a,a69128a,a69132a,a69133a,a69136a,a69139a,a69140a,a69141a,a69145a,a69146a,a69149a,a69152a,a69153a,a69154a,a69158a,a69159a,a69162a,a69165a,a69166a,a69167a,a69171a,a69172a,a69175a,a69178a,a69179a,a69180a,a69184a,a69185a,a69188a,a69191a,a69192a,a69193a,a69197a,a69198a,a69201a,a69204a,a69205a,a69206a,a69210a,a69211a,a69214a,a69217a,a69218a,a69219a,a69223a,a69224a,a69227a,a69230a,a69231a,a69232a,a69236a,a69237a,a69240a,a69243a,a69244a,a69245a,a69249a,a69250a,a69253a,a69256a,a69257a,a69258a,a69262a,a69263a,a69266a,a69269a,a69270a,a69271a,a69275a,a69276a,a69279a,a69282a,a69283a,a69284a,a69288a,a69289a,a69292a,a69295a,a69296a,a69297a,a69301a,a69302a,a69305a,a69308a,a69309a,a69310a,a69314a,a69315a,a69318a,a69321a,a69322a,a69323a,a69327a,a69328a,a69331a,a69334a,a69335a,a69336a,a69340a,a69341a,a69344a,a69347a,a69348a,a69349a,a69353a,a69354a,a69357a,a69360a,a69361a,a69362a,a69366a,a69367a,a69370a,a69373a,a69374a,a69375a,a69379a,a69380a,a69383a,a69386a,a69387a,a69388a,a69392a,a69393a,a69396a,a69399a,a69400a,a69401a,a69405a,a69406a,a69409a,a69412a,a69413a,a69414a,a69418a,a69419a,a69422a,a69425a,a69426a,a69427a,a69431a,a69432a,a69435a,a69438a,a69439a,a69440a,a69444a,a69445a,a69448a,a69451a,a69452a,a69453a,a69457a,a69458a,a69461a,a69464a,a69465a,a69466a,a69470a,a69471a,a69474a,a69477a,a69478a,a69479a,a69483a,a69484a,a69487a,a69490a,a69491a,a69492a,a69496a,a69497a,a69500a,a69503a,a69504a,a69505a,a69509a,a69510a,a69513a,a69516a,a69517a,a69518a,a69522a,a69523a,a69526a,a69529a,a69530a,a69531a,a69535a,a69536a,a69539a,a69542a,a69543a,a69544a,a69548a,a69549a,a69552a,a69555a,a69556a,a69557a,a69561a,a69562a,a69565a,a69568a,a69569a,a69570a,a69574a,a69575a,a69578a,a69581a,a69582a,a69583a,a69587a,a69588a,a69591a,a69594a,a69595a,a69596a,a69600a,a69601a,a69604a,a69607a,a69608a,a69609a,a69613a,a69614a,a69617a,a69620a,a69621a,a69622a,a69626a,a69627a,a69630a,a69633a,a69634a,a69635a,a69639a,a69640a,a69643a,a69646a,a69647a,a69648a,a69652a,a69653a,a69656a,a69659a,a69660a,a69661a,a69665a,a69666a,a69669a,a69672a,a69673a,a69674a,a69678a,a69679a,a69682a,a69685a,a69686a,a69687a,a69691a,a69692a,a69695a,a69698a,a69699a,a69700a,a69704a,a69705a,a69708a,a69711a,a69712a,a69713a,a69717a,a69718a,a69721a,a69724a,a69725a,a69726a,a69730a,a69731a,a69734a,a69737a,a69738a,a69739a,a69743a,a69744a,a69747a,a69750a,a69751a,a69752a,a69756a,a69757a,a69760a,a69763a,a69764a,a69765a,a69769a,a69770a,a69773a,a69776a,a69777a,a69778a,a69782a,a69783a,a69786a,a69789a,a69790a,a69791a,a69795a,a69796a,a69799a,a69802a,a69803a,a69804a,a69808a,a69809a,a69812a,a69815a,a69816a,a69817a,a69821a,a69822a,a69825a,a69828a,a69829a,a69830a,a69834a,a69835a,a69838a,a69841a,a69842a,a69843a,a69847a,a69848a,a69851a,a69854a,a69855a,a69856a,a69860a,a69861a,a69864a,a69867a,a69868a,a69869a,a69873a,a69874a,a69877a,a69880a,a69881a,a69882a,a69886a,a69887a,a69890a,a69893a,a69894a,a69895a,a69899a,a69900a,a69903a,a69906a,a69907a,a69908a,a69912a,a69913a,a69916a,a69919a,a69920a,a69921a,a69925a,a69926a,a69929a,a69932a,a69933a,a69934a,a69938a,a69939a,a69942a,a69945a,a69946a,a69947a,a69951a,a69952a,a69955a,a69958a,a69959a,a69960a,a69964a,a69965a,a69968a,a69971a,a69972a,a69973a,a69977a,a69978a,a69981a,a69984a,a69985a,a69986a,a69990a,a69991a,a69994a,a69997a,a69998a,a69999a,a70003a,a70004a,a70007a,a70010a,a70011a,a70012a,a70016a,a70017a,a70020a,a70023a,a70024a,a70025a,a70029a,a70030a,a70033a,a70036a,a70037a,a70038a,a70042a,a70043a,a70046a,a70049a,a70050a,a70051a,a70055a,a70056a,a70059a,a70062a,a70063a,a70064a,a70068a,a70069a,a70072a,a70075a,a70076a,a70077a,a70081a,a70082a,a70085a,a70088a,a70089a,a70090a,a70094a,a70095a,a70098a,a70101a,a70102a,a70103a,a70107a,a70108a,a70111a,a70114a,a70115a,a70116a,a70120a,a70121a,a70124a,a70127a,a70128a,a70129a,a70133a,a70134a,a70137a,a70140a,a70141a,a70142a,a70146a,a70147a,a70150a,a70153a,a70154a,a70155a,a70159a,a70160a,a70163a,a70166a,a70167a,a70168a,a70172a,a70173a,a70176a,a70179a,a70180a,a70181a,a70185a,a70186a,a70189a,a70192a,a70193a,a70194a,a70198a,a70199a,a70202a,a70205a,a70206a,a70207a,a70211a,a70212a,a70215a,a70218a,a70219a,a70220a,a70224a,a70225a,a70228a,a70231a,a70232a,a70233a,a70237a,a70238a,a70241a,a70244a,a70245a,a70246a,a70250a,a70251a,a70254a,a70257a,a70258a,a70259a,a70263a,a70264a,a70267a,a70270a,a70271a,a70272a,a70276a,a70277a,a70280a,a70283a,a70284a,a70285a,a70289a,a70290a,a70293a,a70296a,a70297a,a70298a,a70302a,a70303a,a70306a,a70309a,a70310a,a70311a,a70315a,a70316a,a70319a,a70322a,a70323a,a70324a,a70328a,a70329a,a70332a,a70335a,a70336a,a70337a,a70341a,a70342a,a70345a,a70348a,a70349a,a70350a,a70354a,a70355a,a70358a,a70361a,a70362a,a70363a,a70367a,a70368a,a70371a,a70374a,a70375a,a70376a,a70380a,a70381a,a70384a,a70387a,a70388a,a70389a,a70393a,a70394a,a70397a,a70400a,a70401a,a70402a,a70406a,a70407a,a70410a,a70413a,a70414a,a70415a,a70419a,a70420a,a70423a,a70426a,a70427a,a70428a,a70432a,a70433a,a70436a,a70439a,a70440a,a70441a,a70445a,a70446a,a70449a,a70452a,a70453a,a70454a,a70458a,a70459a,a70462a,a70465a,a70466a,a70467a,a70471a,a70472a,a70475a,a70478a,a70479a,a70480a,a70484a,a70485a,a70488a,a70491a,a70492a,a70493a,a70497a,a70498a,a70501a,a70504a,a70505a,a70506a,a70510a,a70511a,a70514a,a70517a,a70518a,a70519a,a70523a,a70524a,a70527a,a70530a,a70531a,a70532a,a70536a,a70537a,a70540a,a70543a,a70544a,a70545a,a70549a,a70550a,a70553a,a70556a,a70557a,a70558a,a70562a,a70563a,a70566a,a70569a,a70570a,a70571a,a70575a,a70576a,a70579a,a70582a,a70583a,a70584a,a70588a,a70589a,a70592a,a70595a,a70596a,a70597a,a70601a,a70602a,a70605a,a70608a,a70609a,a70610a,a70614a,a70615a,a70618a,a70621a,a70622a,a70623a,a70627a,a70628a,a70631a,a70634a,a70635a,a70636a,a70640a,a70641a,a70644a,a70647a,a70648a,a70649a,a70653a,a70654a,a70657a,a70660a,a70661a,a70662a,a70666a,a70667a,a70670a,a70673a,a70674a,a70675a,a70679a,a70680a,a70683a,a70686a,a70687a,a70688a,a70692a,a70693a,a70696a,a70699a,a70700a,a70701a,a70705a,a70706a,a70709a,a70712a,a70713a,a70714a,a70718a,a70719a,a70722a,a70725a,a70726a,a70727a,a70731a,a70732a,a70735a,a70738a,a70739a,a70740a,a70744a,a70745a,a70748a,a70751a,a70752a,a70753a,a70757a,a70758a,a70761a,a70764a,a70765a,a70766a,a70770a,a70771a,a70774a,a70777a,a70778a,a70779a,a70783a,a70784a,a70787a,a70790a,a70791a,a70792a,a70796a,a70797a,a70800a,a70803a,a70804a,a70805a,a70809a,a70810a,a70813a,a70816a,a70817a,a70818a,a70822a,a70823a,a70826a,a70829a,a70830a,a70831a,a70835a,a70836a,a70839a,a70842a,a70843a,a70844a,a70848a,a70849a,a70852a,a70855a,a70856a,a70857a,a70861a,a70862a,a70865a,a70868a,a70869a,a70870a,a70874a,a70875a,a70878a,a70881a,a70882a,a70883a,a70887a,a70888a,a70891a,a70894a,a70895a,a70896a,a70900a,a70901a,a70904a,a70907a,a70908a,a70909a,a70913a,a70914a,a70917a,a70920a,a70921a,a70922a,a70926a,a70927a,a70930a,a70933a,a70934a,a70935a,a70939a,a70940a,a70943a,a70946a,a70947a,a70948a,a70952a,a70953a,a70956a,a70959a,a70960a,a70961a,a70965a,a70966a,a70969a,a70972a,a70973a,a70974a,a70978a,a70979a,a70982a,a70985a,a70986a,a70987a,a70991a,a70992a,a70995a,a70998a,a70999a,a71000a,a71004a,a71005a,a71008a,a71011a,a71012a,a71013a,a71017a,a71018a,a71021a,a71024a,a71025a,a71026a,a71030a,a71031a,a71034a,a71037a,a71038a,a71039a,a71043a,a71044a,a71047a,a71050a,a71051a,a71052a,a71056a,a71057a,a71060a,a71063a,a71064a,a71065a,a71069a,a71070a,a71073a,a71076a,a71077a,a71078a,a71082a,a71083a,a71086a,a71089a,a71090a,a71091a,a71095a,a71096a,a71099a,a71102a,a71103a,a71104a,a71108a,a71109a,a71112a,a71115a,a71116a,a71117a,a71121a,a71122a,a71125a,a71128a,a71129a,a71130a,a71134a,a71135a,a71138a,a71141a,a71142a,a71143a,a71147a,a71148a,a71151a,a71154a,a71155a,a71156a,a71160a,a71161a,a71164a,a71167a,a71168a,a71169a,a71173a,a71174a,a71177a,a71180a,a71181a,a71182a,a71186a,a71187a,a71190a,a71193a,a71194a,a71195a,a71199a,a71200a,a71203a,a71206a,a71207a,a71208a,a71212a,a71213a,a71216a,a71219a,a71220a,a71221a,a71225a,a71226a,a71229a,a71232a,a71233a,a71234a,a71238a,a71239a,a71242a,a71245a,a71246a,a71247a,a71251a,a71252a,a71255a,a71258a,a71259a,a71260a,a71264a,a71265a,a71268a,a71271a,a71272a,a71273a,a71277a,a71278a,a71281a,a71284a,a71285a,a71286a,a71290a,a71291a,a71294a,a71297a,a71298a,a71299a,a71303a,a71304a,a71307a,a71310a,a71311a,a71312a,a71316a,a71317a,a71320a,a71323a,a71324a,a71325a,a71329a,a71330a,a71333a,a71336a,a71337a,a71338a,a71342a,a71343a,a71346a,a71349a,a71350a,a71351a,a71355a,a71356a,a71359a,a71362a,a71363a,a71364a,a71368a,a71369a,a71372a,a71375a,a71376a,a71377a,a71381a,a71382a,a71385a,a71388a,a71389a,a71390a,a71394a,a71395a,a71398a,a71401a,a71402a,a71403a,a71407a,a71408a,a71411a,a71414a,a71415a,a71416a,a71420a,a71421a,a71424a,a71427a,a71428a,a71429a,a71433a,a71434a,a71437a,a71440a,a71441a,a71442a,a71446a,a71447a,a71450a,a71453a,a71454a,a71455a,a71459a,a71460a,a71463a,a71466a,a71467a,a71468a,a71472a,a71473a,a71476a,a71479a,a71480a,a71481a,a71485a,a71486a,a71489a,a71492a,a71493a,a71494a,a71498a,a71499a,a71502a,a71505a,a71506a,a71507a,a71511a,a71512a,a71515a,a71518a,a71519a,a71520a,a71524a,a71525a,a71528a,a71531a,a71532a,a71533a,a71537a,a71538a,a71541a,a71544a,a71545a,a71546a,a71550a,a71551a,a71554a,a71557a,a71558a,a71559a,a71563a,a71564a,a71567a,a71570a,a71571a,a71572a,a71576a,a71577a,a71580a,a71583a,a71584a,a71585a,a71589a,a71590a,a71593a,a71596a,a71597a,a71598a,a71602a,a71603a,a71606a,a71609a,a71610a,a71611a,a71615a,a71616a,a71619a,a71622a,a71623a,a71624a,a71628a,a71629a,a71632a,a71635a,a71636a,a71637a,a71641a,a71642a,a71645a,a71648a,a71649a,a71650a,a71654a,a71655a,a71658a,a71661a,a71662a,a71663a,a71667a,a71668a,a71671a,a71674a,a71675a,a71676a,a71680a,a71681a,a71684a,a71687a,a71688a,a71689a,a71693a,a71694a,a71697a,a71700a,a71701a,a71702a,a71706a,a71707a,a71710a,a71713a,a71714a,a71715a,a71719a,a71720a,a71723a,a71726a,a71727a,a71728a,a71732a,a71733a,a71736a,a71739a,a71740a,a71741a,a71745a,a71746a,a71749a,a71752a,a71753a,a71754a,a71758a,a71759a,a71762a,a71765a,a71766a,a71767a,a71771a,a71772a,a71775a,a71778a,a71779a,a71780a,a71784a,a71785a,a71788a,a71791a,a71792a,a71793a,a71797a,a71798a,a71801a,a71804a,a71805a,a71806a,a71810a,a71811a,a71814a,a71817a,a71818a,a71819a,a71823a,a71824a,a71827a,a71830a,a71831a,a71832a,a71836a,a71837a,a71840a,a71843a,a71844a,a71845a,a71849a,a71850a,a71853a,a71856a,a71857a,a71858a,a71862a,a71863a,a71866a,a71869a,a71870a,a71871a,a71875a,a71876a,a71879a,a71882a,a71883a,a71884a,a71888a,a71889a,a71892a,a71895a,a71896a,a71897a,a71901a,a71902a,a71905a,a71908a,a71909a,a71910a,a71914a,a71915a,a71918a,a71921a,a71922a,a71923a,a71927a,a71928a,a71931a,a71934a,a71935a,a71936a,a71940a,a71941a,a71944a,a71947a,a71948a,a71949a,a71953a,a71954a,a71957a,a71960a,a71961a,a71962a,a71966a,a71967a,a71970a,a71973a,a71974a,a71975a,a71979a,a71980a,a71983a,a71986a,a71987a,a71988a,a71992a,a71993a,a71996a,a71999a,a72000a,a72001a,a72005a,a72006a,a72009a,a72012a,a72013a,a72014a,a72018a,a72019a,a72022a,a72025a,a72026a,a72027a,a72031a,a72032a,a72035a,a72038a,a72039a,a72040a,a72044a,a72045a,a72048a,a72051a,a72052a,a72053a,a72057a,a72058a,a72061a,a72064a,a72065a,a72066a,a72070a,a72071a,a72074a,a72077a,a72078a,a72079a,a72083a,a72084a,a72087a,a72090a,a72091a,a72092a,a72096a,a72097a,a72100a,a72103a,a72104a,a72105a,a72109a,a72110a,a72113a,a72116a,a72117a,a72118a,a72122a,a72123a,a72126a,a72129a,a72130a,a72131a,a72135a,a72136a,a72139a,a72142a,a72143a,a72144a,a72148a,a72149a,a72152a,a72155a,a72156a,a72157a,a72161a,a72162a,a72165a,a72168a,a72169a,a72170a,a72174a,a72175a,a72178a,a72181a,a72182a,a72183a,a72187a,a72188a,a72191a,a72194a,a72195a,a72196a,a72200a,a72201a,a72204a,a72207a,a72208a,a72209a,a72213a,a72214a,a72217a,a72220a,a72221a,a72222a,a72226a,a72227a,a72230a,a72233a,a72234a,a72235a,a72239a,a72240a,a72243a,a72246a,a72247a,a72248a,a72252a,a72253a,a72256a,a72259a,a72260a,a72261a,a72265a,a72266a,a72269a,a72272a,a72273a,a72274a,a72278a,a72279a,a72282a,a72285a,a72286a,a72287a,a72291a,a72292a,a72295a,a72298a,a72299a,a72300a,a72304a,a72305a,a72308a,a72311a,a72312a,a72313a,a72317a,a72318a,a72321a,a72324a,a72325a,a72326a,a72330a,a72331a,a72334a,a72337a,a72338a,a72339a,a72343a,a72344a,a72347a,a72350a,a72351a,a72352a,a72356a,a72357a,a72360a,a72363a,a72364a,a72365a,a72369a,a72370a,a72373a,a72376a,a72377a,a72378a,a72382a,a72383a,a72386a,a72389a,a72390a,a72391a,a72395a,a72396a,a72399a,a72402a,a72403a,a72404a,a72408a,a72409a,a72412a,a72415a,a72416a,a72417a,a72421a,a72422a,a72425a,a72428a,a72429a,a72430a,a72434a,a72435a,a72438a,a72441a,a72442a,a72443a,a72447a,a72448a,a72451a,a72454a,a72455a,a72456a,a72460a,a72461a,a72464a,a72467a,a72468a,a72469a,a72473a,a72474a,a72477a,a72480a,a72481a,a72482a,a72486a,a72487a,a72490a,a72493a,a72494a,a72495a,a72499a,a72500a,a72503a,a72506a,a72507a,a72508a,a72512a,a72513a,a72516a,a72519a,a72520a,a72521a,a72525a,a72526a,a72529a,a72532a,a72533a,a72534a,a72538a,a72539a,a72542a,a72545a,a72546a,a72547a,a72551a,a72552a,a72555a,a72558a,a72559a,a72560a,a72564a,a72565a,a72568a,a72571a,a72572a,a72573a,a72577a,a72578a,a72581a,a72584a,a72585a,a72586a,a72590a,a72591a,a72594a,a72597a,a72598a,a72599a,a72603a,a72604a,a72607a,a72610a,a72611a,a72612a,a72616a,a72617a,a72620a,a72623a,a72624a,a72625a,a72629a,a72630a,a72633a,a72636a,a72637a,a72638a,a72642a,a72643a,a72646a,a72649a,a72650a,a72651a,a72655a,a72656a,a72659a,a72662a,a72663a,a72664a,a72668a,a72669a,a72672a,a72675a,a72676a,a72677a,a72681a,a72682a,a72685a,a72688a,a72689a,a72690a,a72694a,a72695a,a72698a,a72701a,a72702a,a72703a,a72707a,a72708a,a72711a,a72714a,a72715a,a72716a,a72720a,a72721a,a72724a,a72727a,a72728a,a72729a,a72733a,a72734a,a72737a,a72740a,a72741a,a72742a,a72746a,a72747a,a72750a,a72753a,a72754a,a72755a,a72759a,a72760a,a72763a,a72766a,a72767a,a72768a,a72772a,a72773a,a72776a,a72779a,a72780a,a72781a,a72785a,a72786a,a72789a,a72792a,a72793a,a72794a,a72798a,a72799a,a72802a,a72805a,a72806a,a72807a,a72811a,a72812a,a72815a,a72818a,a72819a,a72820a,a72824a,a72825a,a72828a,a72831a,a72832a,a72833a,a72837a,a72838a,a72841a,a72844a,a72845a,a72846a,a72850a,a72851a,a72854a,a72857a,a72858a,a72859a,a72863a,a72864a,a72867a,a72870a,a72871a,a72872a,a72876a,a72877a,a72880a,a72883a,a72884a,a72885a,a72889a,a72890a,a72893a,a72896a,a72897a,a72898a,a72902a,a72903a,a72906a,a72909a,a72910a,a72911a,a72915a,a72916a,a72919a,a72922a,a72923a,a72924a,a72928a,a72929a,a72932a,a72935a,a72936a,a72937a,a72941a,a72942a,a72945a,a72948a,a72949a,a72950a,a72954a,a72955a,a72958a,a72961a,a72962a,a72963a,a72967a,a72968a,a72971a,a72974a,a72975a,a72976a,a72980a,a72981a,a72984a,a72987a,a72988a,a72989a,a72993a,a72994a,a72997a,a73000a,a73001a,a73002a,a73006a,a73007a,a73010a,a73013a,a73014a,a73015a,a73019a,a73020a,a73023a,a73026a,a73027a,a73028a,a73032a,a73033a,a73036a,a73039a,a73040a,a73041a,a73045a,a73046a,a73049a,a73052a,a73053a,a73054a,a73058a,a73059a,a73062a,a73065a,a73066a,a73067a,a73071a,a73072a,a73075a,a73078a,a73079a,a73080a,a73084a,a73085a,a73088a,a73091a,a73092a,a73093a,a73097a,a73098a,a73101a,a73104a,a73105a,a73106a,a73110a,a73111a,a73114a,a73117a,a73118a,a73119a,a73123a,a73124a,a73127a,a73130a,a73131a,a73132a,a73136a,a73137a,a73140a,a73143a,a73144a,a73145a,a73149a,a73150a,a73153a,a73156a,a73157a,a73158a,a73162a,a73163a,a73166a,a73169a,a73170a,a73171a,a73175a,a73176a,a73179a,a73182a,a73183a,a73184a,a73188a,a73189a,a73192a,a73195a,a73196a,a73197a,a73201a,a73202a,a73205a,a73208a,a73209a,a73210a,a73214a,a73215a,a73218a,a73221a,a73222a,a73223a,a73227a,a73228a,a73231a,a73234a,a73235a,a73236a,a73240a,a73241a,a73244a,a73247a,a73248a,a73249a,a73253a,a73254a,a73257a,a73260a,a73261a,a73262a,a73266a,a73267a,a73270a,a73273a,a73274a,a73275a,a73279a,a73280a,a73283a,a73286a,a73287a,a73288a,a73292a,a73293a,a73296a,a73299a,a73300a,a73301a,a73305a,a73306a,a73309a,a73312a,a73313a,a73314a,a73318a,a73319a,a73322a,a73325a,a73326a,a73327a,a73331a,a73332a,a73335a,a73338a,a73339a,a73340a,a73344a,a73345a,a73348a,a73351a,a73352a,a73353a,a73357a,a73358a,a73361a,a73364a,a73365a,a73366a,a73370a,a73371a,a73374a,a73377a,a73378a,a73379a,a73383a,a73384a,a73387a,a73390a,a73391a,a73392a,a73396a,a73397a,a73400a,a73403a,a73404a,a73405a,a73409a,a73410a,a73413a,a73416a,a73417a,a73418a,a73422a,a73423a,a73426a,a73429a,a73430a,a73431a,a73435a,a73436a,a73439a,a73442a,a73443a,a73444a,a73448a,a73449a,a73452a,a73455a,a73456a,a73457a,a73461a,a73462a,a73465a,a73468a,a73469a,a73470a,a73474a,a73475a,a73478a,a73481a,a73482a,a73483a,a73487a,a73488a,a73491a,a73494a,a73495a,a73496a,a73500a,a73501a,a73504a,a73507a,a73508a,a73509a,a73513a,a73514a,a73517a,a73520a,a73521a,a73522a,a73526a,a73527a,a73530a,a73533a,a73534a,a73535a,a73539a,a73540a,a73543a,a73546a,a73547a,a73548a,a73552a,a73553a,a73556a,a73559a,a73560a,a73561a,a73565a,a73566a,a73569a,a73572a,a73573a,a73574a,a73578a,a73579a,a73582a,a73585a,a73586a,a73587a,a73591a,a73592a,a73595a,a73598a,a73599a,a73600a,a73604a,a73605a,a73608a,a73611a,a73612a,a73613a,a73617a,a73618a,a73621a,a73624a,a73625a,a73626a,a73630a,a73631a,a73634a,a73637a,a73638a,a73639a,a73643a,a73644a,a73647a,a73650a,a73651a,a73652a,a73656a,a73657a,a73660a,a73663a,a73664a,a73665a,a73669a,a73670a,a73673a,a73676a,a73677a,a73678a,a73682a,a73683a,a73686a,a73689a,a73690a,a73691a,a73695a,a73696a,a73699a,a73702a,a73703a,a73704a,a73708a,a73709a,a73712a,a73715a,a73716a,a73717a,a73721a,a73722a,a73725a,a73728a,a73729a,a73730a,a73734a,a73735a,a73738a,a73741a,a73742a,a73743a,a73747a,a73748a,a73751a,a73754a,a73755a,a73756a,a73760a,a73761a,a73764a,a73767a,a73768a,a73769a,a73773a,a73774a,a73777a,a73780a,a73781a,a73782a,a73786a,a73787a,a73790a,a73793a,a73794a,a73795a,a73799a,a73800a,a73803a,a73806a,a73807a,a73808a,a73812a,a73813a,a73816a,a73819a,a73820a,a73821a,a73825a,a73826a,a73829a,a73832a,a73833a,a73834a,a73838a,a73839a,a73842a,a73845a,a73846a,a73847a,a73851a,a73852a,a73855a,a73858a,a73859a,a73860a,a73864a,a73865a,a73868a,a73871a,a73872a,a73873a,a73877a,a73878a,a73881a,a73884a,a73885a,a73886a,a73890a,a73891a,a73894a,a73897a,a73898a,a73899a,a73903a,a73904a,a73907a,a73910a,a73911a,a73912a,a73916a,a73917a,a73920a,a73923a,a73924a,a73925a,a73929a,a73930a,a73933a,a73936a,a73937a,a73938a,a73942a,a73943a,a73946a,a73949a,a73950a,a73951a,a73955a,a73956a,a73959a,a73962a,a73963a,a73964a,a73968a,a73969a,a73972a,a73975a,a73976a,a73977a,a73981a,a73982a,a73985a,a73988a,a73989a,a73990a,a73994a,a73995a,a73998a,a74001a,a74002a,a74003a,a74007a,a74008a,a74011a,a74014a,a74015a,a74016a,a74020a,a74021a,a74024a,a74027a,a74028a,a74029a,a74033a,a74034a,a74037a,a74040a,a74041a,a74042a,a74046a,a74047a,a74050a,a74053a,a74054a,a74055a,a74059a,a74060a,a74063a,a74066a,a74067a,a74068a,a74072a,a74073a,a74076a,a74079a,a74080a,a74081a,a74085a,a74086a,a74089a,a74092a,a74093a,a74094a,a74098a,a74099a,a74102a,a74105a,a74106a,a74107a,a74111a,a74112a,a74115a,a74118a,a74119a,a74120a,a74124a,a74125a,a74128a,a74131a,a74132a,a74133a,a74137a,a74138a,a74141a,a74144a,a74145a,a74146a,a74150a,a74151a,a74154a,a74157a,a74158a,a74159a,a74163a,a74164a,a74167a,a74170a,a74171a,a74172a,a74176a,a74177a,a74180a,a74183a,a74184a,a74185a,a74189a,a74190a,a74193a,a74196a,a74197a,a74198a,a74202a,a74203a,a74206a,a74209a,a74210a,a74211a,a74215a,a74216a,a74219a,a74222a,a74223a,a74224a,a74228a,a74229a,a74232a,a74235a,a74236a,a74237a,a74241a,a74242a,a74245a,a74248a,a74249a,a74250a,a74254a,a74255a,a74258a,a74261a,a74262a,a74263a,a74267a,a74268a,a74271a,a74274a,a74275a,a74276a,a74280a,a74281a,a74284a,a74287a,a74288a,a74289a,a74292a,a74295a,a74296a,a74299a,a74302a,a74303a,a74304a,a74308a,a74309a,a74312a,a74315a,a74316a,a74317a,a74320a,a74323a,a74324a,a74327a,a74330a,a74331a,a74332a,a74336a,a74337a,a74340a,a74343a,a74344a,a74345a,a74348a,a74351a,a74352a,a74355a,a74358a,a74359a,a74360a,a74364a,a74365a,a74368a,a74371a,a74372a,a74373a,a74376a,a74379a,a74380a,a74383a,a74386a,a74387a,a74388a,a74392a,a74393a,a74396a,a74399a,a74400a,a74401a,a74404a,a74407a,a74408a,a74411a,a74414a,a74415a,a74416a,a74420a,a74421a,a74424a,a74427a,a74428a,a74429a,a74432a,a74435a,a74436a,a74439a,a74442a,a74443a,a74444a,a74448a,a74449a,a74452a,a74455a,a74456a,a74457a,a74460a,a74463a,a74464a,a74467a,a74470a,a74471a,a74472a,a74476a,a74477a,a74480a,a74483a,a74484a,a74485a,a74488a,a74491a,a74492a,a74495a,a74498a,a74499a,a74500a,a74504a,a74505a,a74508a,a74511a,a74512a,a74513a,a74516a,a74519a,a74520a,a74523a,a74526a,a74527a,a74528a,a74532a,a74533a,a74536a,a74539a,a74540a,a74541a,a74544a,a74547a,a74548a,a74551a,a74554a,a74555a,a74556a,a74560a,a74561a,a74564a,a74567a,a74568a,a74569a,a74572a,a74575a,a74576a,a74579a,a74582a,a74583a,a74584a,a74588a,a74589a,a74592a,a74595a,a74596a,a74597a,a74600a,a74603a,a74604a,a74607a,a74610a,a74611a,a74612a,a74616a,a74617a,a74620a,a74623a,a74624a,a74625a,a74628a,a74631a,a74632a,a74635a,a74638a,a74639a,a74640a,a74644a,a74645a,a74648a,a74651a,a74652a,a74653a,a74656a,a74659a,a74660a,a74663a,a74666a,a74667a,a74668a,a74672a,a74673a,a74676a,a74679a,a74680a,a74681a,a74684a,a74687a,a74688a,a74691a,a74694a,a74695a,a74696a,a74700a,a74701a,a74704a,a74707a,a74708a,a74709a,a74712a,a74715a,a74716a,a74719a,a74722a,a74723a,a74724a,a74728a,a74729a,a74732a,a74735a,a74736a,a74737a,a74740a,a74743a,a74744a,a74747a,a74750a,a74751a,a74752a,a74756a,a74757a,a74760a,a74763a,a74764a,a74765a,a74768a,a74771a,a74772a,a74775a,a74778a,a74779a,a74780a,a74784a,a74785a,a74788a,a74791a,a74792a,a74793a,a74796a,a74799a,a74800a,a74803a,a74806a,a74807a,a74808a,a74812a,a74813a,a74816a,a74819a,a74820a,a74821a,a74824a,a74827a,a74828a,a74831a,a74834a,a74835a,a74836a,a74840a,a74841a,a74844a,a74847a,a74848a,a74849a,a74852a,a74855a,a74856a,a74859a,a74862a,a74863a,a74864a,a74868a,a74869a,a74872a,a74875a,a74876a,a74877a,a74880a,a74883a,a74884a,a74887a,a74890a,a74891a,a74892a,a74896a,a74897a,a74900a,a74903a,a74904a,a74905a,a74908a,a74911a,a74912a,a74915a,a74918a,a74919a,a74920a,a74924a,a74925a,a74928a,a74931a,a74932a,a74933a,a74936a,a74939a,a74940a,a74943a,a74946a,a74947a,a74948a,a74952a,a74953a,a74956a,a74959a,a74960a,a74961a,a74964a,a74967a,a74968a,a74971a,a74974a,a74975a,a74976a,a74980a,a74981a,a74984a,a74987a,a74988a,a74989a,a74992a,a74995a,a74996a,a74999a,a75002a,a75003a,a75004a,a75008a,a75009a,a75012a,a75015a,a75016a,a75017a,a75020a,a75023a,a75024a,a75027a,a75030a,a75031a,a75032a,a75036a,a75037a,a75040a,a75043a,a75044a,a75045a,a75048a,a75051a,a75052a,a75055a,a75058a,a75059a,a75060a,a75064a,a75065a,a75068a,a75071a,a75072a,a75073a,a75076a,a75079a,a75080a,a75083a,a75086a,a75087a,a75088a,a75092a,a75093a,a75096a,a75099a,a75100a,a75101a,a75104a,a75107a,a75108a,a75111a,a75114a,a75115a,a75116a,a75120a,a75121a,a75124a,a75127a,a75128a,a75129a,a75132a,a75135a,a75136a,a75139a,a75142a,a75143a,a75144a,a75148a,a75149a,a75152a,a75155a,a75156a,a75157a,a75160a,a75163a,a75164a,a75167a,a75170a,a75171a,a75172a,a75176a,a75177a,a75180a,a75183a,a75184a,a75185a,a75188a,a75191a,a75192a,a75195a,a75198a,a75199a,a75200a,a75204a,a75205a,a75208a,a75211a,a75212a,a75213a,a75216a,a75219a,a75220a,a75223a,a75226a,a75227a,a75228a,a75232a,a75233a,a75236a,a75239a,a75240a,a75241a,a75244a,a75247a,a75248a,a75251a,a75254a,a75255a,a75256a,a75260a,a75261a,a75264a,a75267a,a75268a,a75269a,a75272a,a75275a,a75276a,a75279a,a75282a,a75283a,a75284a,a75288a,a75289a,a75292a,a75295a,a75296a,a75297a,a75300a,a75303a,a75304a,a75307a,a75310a,a75311a,a75312a,a75316a,a75317a,a75320a,a75323a,a75324a,a75325a,a75328a,a75331a,a75332a,a75335a,a75338a,a75339a,a75340a,a75344a,a75345a,a75348a,a75351a,a75352a,a75353a,a75356a,a75359a,a75360a,a75363a,a75366a,a75367a,a75368a,a75372a,a75373a,a75376a,a75379a,a75380a,a75381a,a75384a,a75387a,a75388a,a75391a,a75394a,a75395a,a75396a,a75400a,a75401a,a75404a,a75407a,a75408a,a75409a,a75412a,a75415a,a75416a,a75419a,a75422a,a75423a,a75424a,a75428a,a75429a,a75432a,a75435a,a75436a,a75437a,a75440a,a75443a,a75444a,a75447a,a75450a,a75451a,a75452a,a75456a,a75457a,a75460a,a75463a,a75464a,a75465a,a75468a,a75471a,a75472a,a75475a,a75478a,a75479a,a75480a,a75484a,a75485a,a75488a,a75491a,a75492a,a75493a,a75496a,a75499a,a75500a,a75503a,a75506a,a75507a,a75508a,a75512a,a75513a,a75516a,a75519a,a75520a,a75521a,a75524a,a75527a,a75528a,a75531a,a75534a,a75535a,a75536a,a75540a,a75541a,a75544a,a75547a,a75548a,a75549a,a75552a,a75555a,a75556a,a75559a,a75562a,a75563a,a75564a,a75568a,a75569a,a75572a,a75575a,a75576a,a75577a,a75580a,a75583a,a75584a,a75587a,a75590a,a75591a,a75592a,a75596a,a75597a,a75600a,a75603a,a75604a,a75605a,a75608a,a75611a,a75612a,a75615a,a75618a,a75619a,a75620a,a75624a,a75625a,a75628a,a75631a,a75632a,a75633a,a75636a,a75639a,a75640a,a75643a,a75646a,a75647a,a75648a,a75652a,a75653a,a75656a,a75659a,a75660a,a75661a,a75664a,a75667a,a75668a,a75671a,a75674a,a75675a,a75676a,a75680a,a75681a,a75684a,a75687a,a75688a,a75689a,a75692a,a75695a,a75696a,a75699a,a75702a,a75703a,a75704a,a75708a,a75709a,a75712a,a75715a,a75716a,a75717a,a75720a,a75723a,a75724a,a75727a,a75730a,a75731a,a75732a,a75736a,a75737a,a75740a,a75743a,a75744a,a75745a,a75748a,a75751a,a75752a,a75755a,a75758a,a75759a,a75760a,a75764a,a75765a,a75768a,a75771a,a75772a,a75773a,a75776a,a75779a,a75780a,a75783a,a75786a,a75787a,a75788a,a75792a,a75793a,a75796a,a75799a,a75800a,a75801a,a75804a,a75807a,a75808a,a75811a,a75814a,a75815a,a75816a,a75820a,a75821a,a75824a,a75827a,a75828a,a75829a,a75832a,a75835a,a75836a,a75839a,a75842a,a75843a,a75844a,a75848a,a75849a,a75852a,a75855a,a75856a,a75857a,a75860a,a75863a,a75864a,a75867a,a75870a,a75871a,a75872a,a75876a,a75877a,a75880a,a75883a,a75884a,a75885a,a75888a,a75891a,a75892a,a75895a,a75898a,a75899a,a75900a,a75904a,a75905a,a75908a,a75911a,a75912a,a75913a,a75916a,a75919a,a75920a,a75923a,a75926a,a75927a,a75928a,a75932a,a75933a,a75936a,a75939a,a75940a,a75941a,a75944a,a75947a,a75948a,a75951a,a75954a,a75955a,a75956a,a75960a,a75961a,a75964a,a75967a,a75968a,a75969a,a75972a,a75975a,a75976a,a75979a,a75982a,a75983a,a75984a,a75988a,a75989a,a75992a,a75995a,a75996a,a75997a,a76000a,a76003a,a76004a,a76007a,a76010a,a76011a,a76012a,a76016a,a76017a,a76020a,a76023a,a76024a,a76025a,a76028a,a76031a,a76032a,a76035a,a76038a,a76039a,a76040a,a76044a,a76045a,a76048a,a76051a,a76052a,a76053a,a76056a,a76059a,a76060a,a76063a,a76066a,a76067a,a76068a,a76072a,a76073a,a76076a,a76079a,a76080a,a76081a,a76084a,a76087a,a76088a,a76091a,a76094a,a76095a,a76096a,a76100a,a76101a,a76104a,a76107a,a76108a,a76109a,a76112a,a76115a,a76116a,a76119a,a76122a,a76123a,a76124a,a76128a,a76129a,a76132a,a76135a,a76136a,a76137a,a76140a,a76143a,a76144a,a76147a,a76150a,a76151a,a76152a,a76156a,a76157a,a76160a,a76163a,a76164a,a76165a,a76168a,a76171a,a76172a,a76175a,a76178a,a76179a,a76180a,a76184a,a76185a,a76188a,a76191a,a76192a,a76193a,a76196a,a76199a,a76200a,a76203a,a76206a,a76207a,a76208a,a76212a,a76213a,a76216a,a76219a,a76220a,a76221a,a76224a,a76227a,a76228a,a76231a,a76234a,a76235a,a76236a,a76240a,a76241a,a76244a,a76247a,a76248a,a76249a,a76252a,a76255a,a76256a,a76259a,a76262a,a76263a,a76264a,a76268a,a76269a,a76272a,a76275a,a76276a,a76277a,a76280a,a76283a,a76284a,a76287a,a76290a,a76291a,a76292a,a76296a,a76297a,a76300a,a76303a,a76304a,a76305a,a76308a,a76311a,a76312a,a76315a,a76318a,a76319a,a76320a,a76324a,a76325a,a76328a,a76331a,a76332a,a76333a,a76336a,a76339a,a76340a,a76343a,a76346a,a76347a,a76348a,a76352a,a76353a,a76356a,a76359a,a76360a,a76361a,a76364a,a76367a,a76368a,a76371a,a76374a,a76375a,a76376a,a76380a,a76381a,a76384a,a76387a,a76388a,a76389a,a76392a,a76395a,a76396a,a76399a,a76402a,a76403a,a76404a,a76408a,a76409a,a76412a,a76415a,a76416a,a76417a,a76420a,a76423a,a76424a,a76427a,a76430a,a76431a,a76432a,a76436a,a76437a,a76440a,a76443a,a76444a,a76445a,a76448a,a76451a,a76452a,a76455a,a76458a,a76459a,a76460a,a76464a,a76465a,a76468a,a76471a,a76472a,a76473a,a76476a,a76479a,a76480a,a76483a,a76486a,a76487a,a76488a,a76492a,a76493a,a76496a,a76499a,a76500a,a76501a,a76504a,a76507a,a76508a,a76511a,a76514a,a76515a,a76516a,a76520a,a76521a,a76524a,a76527a,a76528a,a76529a,a76532a,a76535a,a76536a,a76539a,a76542a,a76543a,a76544a,a76548a,a76549a,a76552a,a76555a,a76556a,a76557a,a76560a,a76563a,a76564a,a76567a,a76570a,a76571a,a76572a,a76576a,a76577a,a76580a,a76583a,a76584a,a76585a,a76588a,a76591a,a76592a,a76595a,a76598a,a76599a,a76600a,a76604a,a76605a,a76608a,a76611a,a76612a,a76613a,a76616a,a76619a,a76620a,a76623a,a76626a,a76627a,a76628a,a76632a,a76633a,a76636a,a76639a,a76640a,a76641a,a76644a,a76647a,a76648a,a76651a,a76654a,a76655a,a76656a,a76660a,a76661a,a76664a,a76667a,a76668a,a76669a,a76672a,a76675a,a76676a,a76679a,a76682a,a76683a,a76684a,a76688a,a76689a,a76692a,a76695a,a76696a,a76697a,a76700a,a76703a,a76704a,a76707a,a76710a,a76711a,a76712a,a76716a,a76717a,a76720a,a76723a,a76724a,a76725a,a76728a,a76731a,a76732a,a76735a,a76738a,a76739a,a76740a,a76744a,a76745a,a76748a,a76751a,a76752a,a76753a,a76756a,a76759a,a76760a,a76763a,a76766a,a76767a,a76768a,a76772a,a76773a,a76776a,a76779a,a76780a,a76781a,a76784a,a76787a,a76788a,a76791a,a76794a,a76795a,a76796a,a76800a,a76801a,a76804a,a76807a,a76808a,a76809a,a76812a,a76815a,a76816a,a76819a,a76822a,a76823a,a76824a,a76828a,a76829a,a76832a,a76835a,a76836a,a76837a,a76840a,a76843a,a76844a,a76847a,a76850a,a76851a,a76852a,a76856a,a76857a,a76860a,a76863a,a76864a,a76865a,a76868a,a76871a,a76872a,a76875a,a76878a,a76879a,a76880a,a76884a,a76885a,a76888a,a76891a,a76892a,a76893a,a76896a,a76899a,a76900a,a76903a,a76906a,a76907a,a76908a,a76912a,a76913a,a76916a,a76919a,a76920a,a76921a,a76924a,a76927a,a76928a,a76931a,a76934a,a76935a,a76936a,a76940a,a76941a,a76944a,a76947a,a76948a,a76949a,a76952a,a76955a,a76956a,a76959a,a76962a,a76963a,a76964a,a76968a,a76969a,a76972a,a76975a,a76976a,a76977a,a76980a,a76983a,a76984a,a76987a,a76990a,a76991a,a76992a,a76996a,a76997a,a77000a,a77003a,a77004a,a77005a,a77008a,a77011a,a77012a,a77015a,a77018a,a77019a,a77020a,a77024a,a77025a,a77028a,a77031a,a77032a,a77033a,a77036a,a77039a,a77040a,a77043a,a77046a,a77047a,a77048a,a77052a,a77053a,a77056a,a77059a,a77060a,a77061a,a77064a,a77067a,a77068a,a77071a,a77074a,a77075a,a77076a,a77080a,a77081a,a77084a,a77087a,a77088a,a77089a,a77092a,a77095a,a77096a,a77099a,a77102a,a77103a,a77104a,a77108a,a77109a,a77112a,a77115a,a77116a,a77117a,a77120a,a77123a,a77124a,a77127a,a77130a,a77131a,a77132a,a77136a,a77137a,a77140a,a77143a,a77144a,a77145a,a77148a,a77151a,a77152a,a77155a,a77158a,a77159a,a77160a,a77164a,a77165a,a77168a,a77171a,a77172a,a77173a,a77176a,a77179a,a77180a,a77183a,a77186a,a77187a,a77188a,a77192a,a77193a,a77196a,a77199a,a77200a,a77201a,a77204a,a77207a,a77208a,a77211a,a77214a,a77215a,a77216a,a77220a,a77221a,a77224a,a77227a,a77228a,a77229a,a77232a,a77235a,a77236a,a77239a,a77242a,a77243a,a77244a,a77248a,a77249a,a77252a,a77255a,a77256a,a77257a,a77260a,a77263a,a77264a,a77267a,a77270a,a77271a,a77272a,a77276a,a77277a,a77280a,a77283a,a77284a,a77285a,a77288a,a77291a,a77292a,a77295a,a77298a,a77299a,a77300a,a77304a,a77305a,a77308a,a77311a,a77312a,a77313a,a77316a,a77319a,a77320a,a77323a,a77326a,a77327a,a77328a,a77332a,a77333a,a77336a,a77339a,a77340a,a77341a,a77344a,a77347a,a77348a,a77351a,a77354a,a77355a,a77356a,a77360a,a77361a,a77364a,a77367a,a77368a,a77369a,a77372a,a77375a,a77376a,a77379a,a77382a,a77383a,a77384a,a77388a,a77389a,a77392a,a77395a,a77396a,a77397a,a77400a,a77403a,a77404a,a77407a,a77410a,a77411a,a77412a,a77416a,a77417a,a77420a,a77423a,a77424a,a77425a,a77428a,a77431a,a77432a,a77435a,a77438a,a77439a,a77440a,a77444a,a77445a,a77448a,a77451a,a77452a,a77453a,a77456a,a77459a,a77460a,a77463a,a77466a,a77467a,a77468a,a77472a,a77473a,a77476a,a77479a,a77480a,a77481a,a77484a,a77487a,a77488a,a77491a,a77494a,a77495a,a77496a,a77500a,a77501a,a77504a,a77507a,a77508a,a77509a,a77512a,a77515a,a77516a,a77519a,a77522a,a77523a,a77524a,a77528a,a77529a,a77532a,a77535a,a77536a,a77537a,a77540a,a77543a,a77544a,a77547a,a77550a,a77551a,a77552a,a77556a,a77557a,a77560a,a77563a,a77564a,a77565a,a77568a,a77571a,a77572a,a77575a,a77578a,a77579a,a77580a,a77584a,a77585a,a77588a,a77591a,a77592a,a77593a,a77596a,a77599a,a77600a,a77603a,a77606a,a77607a,a77608a,a77612a,a77613a,a77616a,a77619a,a77620a,a77621a,a77624a,a77627a,a77628a,a77631a,a77634a,a77635a,a77636a,a77640a,a77641a,a77644a,a77647a,a77648a,a77649a,a77652a,a77655a,a77656a,a77659a,a77662a,a77663a,a77664a,a77668a,a77669a,a77672a,a77675a,a77676a,a77677a,a77680a,a77683a,a77684a,a77687a,a77690a,a77691a,a77692a,a77696a,a77697a,a77700a,a77703a,a77704a,a77705a,a77708a,a77711a,a77712a,a77715a,a77718a,a77719a,a77720a,a77724a,a77725a,a77728a,a77731a,a77732a,a77733a,a77736a,a77739a,a77740a,a77743a,a77746a,a77747a,a77748a,a77752a,a77753a,a77756a,a77759a,a77760a,a77761a,a77764a,a77767a,a77768a,a77771a,a77774a,a77775a,a77776a,a77780a,a77781a,a77784a,a77787a,a77788a,a77789a,a77792a,a77795a,a77796a,a77799a,a77802a,a77803a,a77804a,a77808a,a77809a,a77812a,a77815a,a77816a,a77817a,a77820a,a77823a,a77824a,a77827a,a77830a,a77831a,a77832a,a77836a,a77837a,a77840a,a77843a,a77844a,a77845a,a77848a,a77851a,a77852a,a77855a,a77858a,a77859a,a77860a,a77864a,a77865a,a77868a,a77871a,a77872a,a77873a,a77876a,a77879a,a77880a,a77883a,a77886a,a77887a,a77888a,a77892a,a77893a,a77896a,a77899a,a77900a,a77901a,a77904a,a77907a,a77908a,a77911a,a77914a,a77915a,a77916a,a77920a,a77921a,a77924a,a77927a,a77928a,a77929a,a77932a,a77935a,a77936a,a77939a,a77942a,a77943a,a77944a,a77948a,a77949a,a77952a,a77955a,a77956a,a77957a,a77960a,a77963a,a77964a,a77967a,a77970a,a77971a,a77972a,a77976a,a77977a,a77980a,a77983a,a77984a,a77985a,a77988a,a77991a,a77992a,a77995a,a77998a,a77999a,a78000a,a78004a,a78005a,a78008a,a78011a,a78012a,a78013a,a78016a,a78019a,a78020a,a78023a,a78026a,a78027a,a78028a,a78032a,a78033a,a78036a,a78039a,a78040a,a78041a,a78044a,a78047a,a78048a,a78051a,a78054a,a78055a,a78056a,a78060a,a78061a,a78064a,a78067a,a78068a,a78069a,a78072a,a78075a,a78076a,a78079a,a78082a,a78083a,a78084a,a78088a,a78089a,a78092a,a78095a,a78096a,a78097a,a78100a,a78103a,a78104a,a78107a,a78110a,a78111a,a78112a,a78116a,a78117a,a78120a,a78123a,a78124a,a78125a,a78128a,a78131a,a78132a,a78135a,a78138a,a78139a,a78140a,a78144a,a78145a,a78148a,a78151a,a78152a,a78153a,a78156a,a78159a,a78160a,a78163a,a78166a,a78167a,a78168a,a78172a,a78173a,a78176a,a78179a,a78180a,a78181a,a78184a,a78187a,a78188a,a78191a,a78194a,a78195a,a78196a,a78200a,a78201a,a78204a,a78207a,a78208a,a78209a,a78212a,a78215a,a78216a,a78219a,a78222a,a78223a,a78224a,a78228a,a78229a,a78232a,a78235a,a78236a,a78237a,a78240a,a78243a,a78244a,a78247a,a78250a,a78251a,a78252a,a78256a,a78257a,a78260a,a78263a,a78264a,a78265a,a78268a,a78271a,a78272a,a78275a,a78278a,a78279a,a78280a,a78284a,a78285a,a78288a,a78291a,a78292a,a78293a,a78296a,a78299a,a78300a,a78303a,a78306a,a78307a,a78308a,a78312a,a78313a,a78316a,a78319a,a78320a,a78321a,a78324a,a78327a,a78328a,a78331a,a78334a,a78335a,a78336a,a78340a,a78341a,a78344a,a78347a,a78348a,a78349a,a78352a,a78355a,a78356a,a78359a,a78362a,a78363a,a78364a,a78368a,a78369a,a78372a,a78375a,a78376a,a78377a,a78380a,a78383a,a78384a,a78387a,a78390a,a78391a,a78392a,a78396a,a78397a,a78400a,a78403a,a78404a,a78405a,a78408a,a78411a,a78412a,a78415a,a78418a,a78419a,a78420a,a78424a,a78425a,a78428a,a78431a,a78432a,a78433a,a78436a,a78439a,a78440a,a78443a,a78446a,a78447a,a78448a,a78452a,a78453a,a78456a,a78459a,a78460a,a78461a,a78464a,a78467a,a78468a,a78471a,a78474a,a78475a,a78476a,a78480a,a78481a,a78484a,a78487a,a78488a,a78489a,a78492a,a78495a,a78496a,a78499a,a78502a,a78503a,a78504a,a78508a,a78509a,a78512a,a78515a,a78516a,a78517a,a78520a,a78523a,a78524a,a78527a,a78530a,a78531a,a78532a,a78536a,a78537a,a78540a,a78543a,a78544a,a78545a,a78548a,a78551a,a78552a,a78555a,a78558a,a78559a,a78560a,a78564a,a78565a,a78568a,a78571a,a78572a,a78573a,a78576a,a78579a,a78580a,a78583a,a78586a,a78587a,a78588a,a78592a,a78593a,a78596a,a78599a,a78600a,a78601a,a78604a,a78607a,a78608a,a78611a,a78614a,a78615a,a78616a,a78620a,a78621a,a78624a,a78627a,a78628a,a78629a,a78632a,a78635a,a78636a,a78639a,a78642a,a78643a,a78644a,a78648a,a78649a,a78652a,a78655a,a78656a,a78657a,a78660a,a78663a,a78664a,a78667a,a78670a,a78671a,a78672a,a78676a,a78677a,a78680a,a78683a,a78684a,a78685a,a78688a,a78691a,a78692a,a78695a,a78698a,a78699a,a78700a,a78704a,a78705a,a78708a,a78711a,a78712a,a78713a,a78716a,a78719a,a78720a,a78723a,a78726a,a78727a,a78728a,a78732a,a78733a,a78736a,a78739a,a78740a,a78741a,a78744a,a78747a,a78748a,a78751a,a78754a,a78755a,a78756a,a78760a,a78761a,a78764a,a78767a,a78768a,a78769a,a78772a,a78775a,a78776a,a78779a,a78782a,a78783a,a78784a,a78788a,a78789a,a78792a,a78795a,a78796a,a78797a,a78800a,a78803a,a78804a,a78807a,a78810a,a78811a,a78812a,a78816a,a78817a,a78820a,a78823a,a78824a,a78825a,a78828a,a78831a,a78832a,a78835a,a78838a,a78839a,a78840a,a78844a,a78845a,a78848a,a78851a,a78852a,a78853a,a78856a,a78859a,a78860a,a78863a,a78866a,a78867a,a78868a,a78872a,a78873a,a78876a,a78879a,a78880a,a78881a,a78884a,a78887a,a78888a,a78891a,a78894a,a78895a,a78896a,a78900a,a78901a,a78904a,a78907a,a78908a,a78909a,a78912a,a78915a,a78916a,a78919a,a78922a,a78923a,a78924a,a78928a,a78929a,a78932a,a78935a,a78936a,a78937a,a78940a,a78943a,a78944a,a78947a,a78950a,a78951a,a78952a,a78956a,a78957a,a78960a,a78963a,a78964a,a78965a,a78968a,a78971a,a78972a,a78975a,a78978a,a78979a,a78980a,a78984a,a78985a,a78988a,a78991a,a78992a,a78993a,a78996a,a78999a,a79000a,a79003a,a79006a,a79007a,a79008a,a79012a,a79013a,a79016a,a79019a,a79020a,a79021a,a79024a,a79027a,a79028a,a79031a,a79034a,a79035a,a79036a,a79040a,a79041a,a79044a,a79047a,a79048a,a79049a,a79052a,a79055a,a79056a,a79059a,a79062a,a79063a,a79064a,a79068a,a79069a,a79072a,a79075a,a79076a,a79077a,a79080a,a79083a,a79084a,a79087a,a79090a,a79091a,a79092a,a79096a,a79097a,a79100a,a79103a,a79104a,a79105a,a79108a,a79111a,a79112a,a79115a,a79118a,a79119a,a79120a,a79124a,a79125a,a79128a,a79131a,a79132a,a79133a,a79136a,a79139a,a79140a,a79143a,a79146a,a79147a,a79148a,a79152a,a79153a,a79156a,a79159a,a79160a,a79161a,a79164a,a79167a,a79168a,a79171a,a79174a,a79175a,a79176a,a79180a,a79181a,a79184a,a79187a,a79188a,a79189a,a79192a,a79195a,a79196a,a79199a,a79202a,a79203a,a79204a,a79208a,a79209a,a79212a,a79215a,a79216a,a79217a,a79220a,a79223a,a79224a,a79227a,a79230a,a79231a,a79232a,a79236a,a79237a,a79240a,a79243a,a79244a,a79245a,a79248a,a79251a,a79252a,a79255a,a79258a,a79259a,a79260a,a79264a,a79265a,a79268a,a79271a,a79272a,a79273a,a79276a,a79279a,a79280a,a79283a,a79286a,a79287a,a79288a,a79292a,a79293a,a79296a,a79299a,a79300a,a79301a,a79304a,a79307a,a79308a,a79311a,a79314a,a79315a,a79316a,a79320a,a79321a,a79324a,a79327a,a79328a,a79329a,a79332a,a79335a,a79336a,a79339a,a79342a,a79343a,a79344a,a79348a,a79349a,a79352a,a79355a,a79356a,a79357a,a79360a,a79363a,a79364a,a79367a,a79370a,a79371a,a79372a,a79376a,a79377a,a79380a,a79383a,a79384a,a79385a,a79388a,a79391a,a79392a,a79395a,a79398a,a79399a,a79400a,a79404a,a79405a,a79408a,a79411a,a79412a,a79413a,a79416a,a79419a,a79420a,a79423a,a79426a,a79427a,a79428a,a79432a,a79433a,a79436a,a79439a,a79440a,a79441a,a79444a,a79447a,a79448a,a79451a,a79454a,a79455a,a79456a,a79460a,a79461a,a79464a,a79467a,a79468a,a79469a,a79472a,a79475a,a79476a,a79479a,a79482a,a79483a,a79484a,a79488a,a79489a,a79492a,a79495a,a79496a,a79497a,a79500a,a79503a,a79504a,a79507a,a79510a,a79511a,a79512a,a79516a,a79517a,a79520a,a79523a,a79524a,a79525a,a79528a,a79531a,a79532a,a79535a,a79538a,a79539a,a79540a,a79544a,a79545a,a79548a,a79551a,a79552a,a79553a,a79556a,a79559a,a79560a,a79563a,a79566a,a79567a,a79568a,a79572a,a79573a,a79576a,a79579a,a79580a,a79581a,a79584a,a79587a,a79588a,a79591a,a79594a,a79595a,a79596a,a79600a,a79601a,a79604a,a79607a,a79608a,a79609a,a79612a,a79615a,a79616a,a79619a,a79622a,a79623a,a79624a,a79628a,a79629a,a79632a,a79635a,a79636a,a79637a,a79640a,a79643a,a79644a,a79647a,a79650a,a79651a,a79652a,a79656a,a79657a,a79660a,a79663a,a79664a,a79665a,a79668a,a79671a,a79672a,a79675a,a79678a,a79679a,a79680a,a79684a,a79685a,a79688a,a79691a,a79692a,a79693a,a79696a,a79699a,a79700a,a79703a,a79706a,a79707a,a79708a,a79712a,a79713a,a79716a,a79719a,a79720a,a79721a,a79724a,a79727a,a79728a,a79731a,a79734a,a79735a,a79736a,a79740a,a79741a,a79744a,a79747a,a79748a,a79749a,a79752a,a79755a,a79756a,a79759a,a79762a,a79763a,a79764a,a79768a,a79769a,a79772a,a79775a,a79776a,a79777a,a79780a,a79783a,a79784a,a79787a,a79790a,a79791a,a79792a,a79796a,a79797a,a79800a,a79803a,a79804a,a79805a,a79808a,a79811a,a79812a,a79815a,a79818a,a79819a,a79820a,a79824a,a79825a,a79828a,a79831a,a79832a,a79833a,a79836a,a79839a,a79840a,a79843a,a79846a,a79847a,a79848a,a79852a,a79853a,a79856a,a79859a,a79860a,a79861a,a79864a,a79867a,a79868a,a79871a,a79874a,a79875a,a79876a,a79880a,a79881a,a79884a,a79887a,a79888a,a79889a,a79892a,a79895a,a79896a,a79899a,a79902a,a79903a,a79904a,a79908a,a79909a,a79912a,a79915a,a79916a,a79917a,a79920a,a79923a,a79924a,a79927a,a79930a,a79931a,a79932a,a79936a,a79937a,a79940a,a79943a,a79944a,a79945a,a79948a,a79951a,a79952a,a79955a,a79958a,a79959a,a79960a,a79964a,a79965a,a79968a,a79971a,a79972a,a79973a,a79976a,a79979a,a79980a,a79983a,a79986a,a79987a,a79988a,a79992a,a79993a,a79996a,a79999a,a80000a,a80001a,a80004a,a80007a,a80008a,a80011a,a80014a,a80015a,a80016a,a80020a,a80021a,a80024a,a80027a,a80028a,a80029a,a80032a,a80035a,a80036a,a80039a,a80042a,a80043a,a80044a,a80048a,a80049a,a80052a,a80055a,a80056a,a80057a,a80060a,a80063a,a80064a,a80067a,a80070a,a80071a,a80072a,a80076a,a80077a,a80080a,a80083a,a80084a,a80085a,a80088a,a80091a,a80092a,a80095a,a80098a,a80099a,a80100a,a80104a,a80105a,a80108a,a80111a,a80112a,a80113a,a80116a,a80119a,a80120a,a80123a,a80126a,a80127a,a80128a,a80132a,a80133a,a80136a,a80139a,a80140a,a80141a,a80144a,a80147a,a80148a,a80151a,a80154a,a80155a,a80156a,a80160a,a80161a,a80164a,a80167a,a80168a,a80169a,a80172a,a80175a,a80176a,a80179a,a80182a,a80183a,a80184a,a80188a,a80189a,a80192a,a80195a,a80196a,a80197a,a80200a,a80203a,a80204a,a80207a,a80210a,a80211a,a80212a,a80216a,a80217a,a80220a,a80223a,a80224a,a80225a,a80228a,a80231a,a80232a,a80235a,a80238a,a80239a,a80240a,a80244a,a80245a,a80248a,a80251a,a80252a,a80253a,a80256a,a80259a,a80260a,a80263a,a80266a,a80267a,a80268a,a80272a,a80273a,a80276a,a80279a,a80280a,a80281a,a80284a,a80287a,a80288a,a80291a,a80294a,a80295a,a80296a,a80300a,a80301a,a80304a,a80307a,a80308a,a80309a,a80312a,a80315a,a80316a,a80319a,a80322a,a80323a,a80324a,a80328a,a80329a,a80332a,a80335a,a80336a,a80337a,a80340a,a80343a,a80344a,a80347a,a80350a,a80351a,a80352a,a80356a,a80357a,a80360a,a80363a,a80364a,a80365a,a80368a,a80371a,a80372a,a80375a,a80378a,a80379a,a80380a,a80384a,a80385a,a80388a,a80391a,a80392a,a80393a,a80396a,a80399a,a80400a,a80403a,a80406a,a80407a,a80408a,a80412a,a80413a,a80416a,a80419a,a80420a,a80421a,a80424a,a80427a,a80428a,a80431a,a80434a,a80435a,a80436a,a80440a,a80441a,a80444a,a80447a,a80448a,a80449a,a80452a,a80455a,a80456a,a80459a,a80462a,a80463a,a80464a,a80468a,a80469a,a80472a,a80475a,a80476a,a80477a,a80480a,a80483a,a80484a,a80487a,a80490a,a80491a,a80492a,a80496a,a80497a,a80500a,a80503a,a80504a,a80505a,a80508a,a80511a,a80512a,a80515a,a80518a,a80519a,a80520a,a80524a,a80525a,a80528a,a80531a,a80532a,a80533a,a80536a,a80539a,a80540a,a80543a,a80546a,a80547a,a80548a,a80552a,a80553a,a80556a,a80559a,a80560a,a80561a,a80564a,a80567a,a80568a,a80571a,a80574a,a80575a,a80576a,a80580a,a80581a,a80584a,a80587a,a80588a,a80589a,a80592a,a80595a,a80596a,a80599a,a80602a,a80603a,a80604a,a80608a,a80609a,a80612a,a80615a,a80616a,a80617a,a80620a,a80623a,a80624a,a80627a,a80630a,a80631a,a80632a,a80636a,a80637a,a80640a,a80643a,a80644a,a80645a,a80648a,a80651a,a80652a,a80655a,a80658a,a80659a,a80660a,a80664a,a80665a,a80668a,a80671a,a80672a,a80673a,a80676a,a80679a,a80680a,a80683a,a80686a,a80687a,a80688a,a80692a,a80693a,a80696a,a80699a,a80700a,a80701a,a80704a,a80707a,a80708a,a80711a,a80714a,a80715a,a80716a,a80720a,a80721a,a80724a,a80727a,a80728a,a80729a,a80732a,a80735a,a80736a,a80739a,a80742a,a80743a,a80744a,a80748a,a80749a,a80752a,a80755a,a80756a,a80757a,a80760a,a80763a,a80764a,a80767a,a80770a,a80771a,a80772a,a80776a,a80777a,a80780a,a80783a,a80784a,a80785a,a80788a,a80791a,a80792a,a80795a,a80798a,a80799a,a80800a,a80804a,a80805a,a80808a,a80811a,a80812a,a80813a,a80816a,a80819a,a80820a,a80823a,a80826a,a80827a,a80828a,a80832a,a80833a,a80836a,a80839a,a80840a,a80841a,a80844a,a80847a,a80848a,a80851a,a80854a,a80855a,a80856a,a80860a,a80861a,a80864a,a80867a,a80868a,a80869a,a80872a,a80875a,a80876a,a80879a,a80882a,a80883a,a80884a,a80888a,a80889a,a80892a,a80895a,a80896a,a80897a,a80900a,a80903a,a80904a,a80907a,a80910a,a80911a,a80912a,a80916a,a80917a,a80920a,a80923a,a80924a,a80925a,a80928a,a80931a,a80932a,a80935a,a80938a,a80939a,a80940a,a80944a,a80945a,a80948a,a80951a,a80952a,a80953a,a80956a,a80959a,a80960a,a80963a,a80966a,a80967a,a80968a,a80972a,a80973a,a80976a,a80979a,a80980a,a80981a,a80984a,a80987a,a80988a,a80991a,a80994a,a80995a,a80996a,a81000a,a81001a,a81004a,a81007a,a81008a,a81009a,a81012a,a81015a,a81016a,a81019a,a81022a,a81023a,a81024a,a81028a,a81029a,a81032a,a81035a,a81036a,a81037a,a81040a,a81043a,a81044a,a81047a,a81050a,a81051a,a81052a,a81056a,a81057a,a81060a,a81063a,a81064a,a81065a,a81068a,a81071a,a81072a,a81075a,a81078a,a81079a,a81080a,a81084a,a81085a,a81088a,a81091a,a81092a,a81093a,a81096a,a81099a,a81100a,a81103a,a81106a,a81107a,a81108a,a81112a,a81113a,a81116a,a81119a,a81120a,a81121a,a81124a,a81127a,a81128a,a81131a,a81134a,a81135a,a81136a,a81140a,a81141a,a81144a,a81147a,a81148a,a81149a,a81152a,a81155a,a81156a,a81159a,a81162a,a81163a,a81164a,a81168a,a81169a,a81172a,a81175a,a81176a,a81177a,a81180a,a81183a,a81184a,a81187a,a81190a,a81191a,a81192a,a81196a,a81197a,a81200a,a81203a,a81204a,a81205a,a81208a,a81211a,a81212a,a81215a,a81218a,a81219a,a81220a,a81224a,a81225a,a81228a,a81231a,a81232a,a81233a,a81236a,a81239a,a81240a,a81243a,a81246a,a81247a,a81248a,a81252a,a81253a,a81256a,a81259a,a81260a,a81261a,a81264a,a81267a,a81268a,a81271a,a81274a,a81275a,a81276a,a81280a,a81281a,a81284a,a81287a,a81288a,a81289a,a81292a,a81295a,a81296a,a81299a,a81302a,a81303a,a81304a,a81308a,a81309a,a81312a,a81315a,a81316a,a81317a,a81320a,a81323a,a81324a,a81327a,a81330a,a81331a,a81332a,a81336a,a81337a,a81340a,a81343a,a81344a,a81345a,a81348a,a81351a,a81352a,a81355a,a81358a,a81359a,a81360a,a81364a,a81365a,a81368a,a81371a,a81372a,a81373a,a81376a,a81379a,a81380a,a81383a,a81386a,a81387a,a81388a,a81392a,a81393a,a81396a,a81399a,a81400a,a81401a,a81404a,a81407a,a81408a,a81411a,a81414a,a81415a,a81416a,a81420a,a81421a,a81424a,a81427a,a81428a,a81429a,a81432a,a81435a,a81436a,a81439a,a81442a,a81443a,a81444a,a81448a,a81449a,a81452a,a81455a,a81456a,a81457a,a81460a,a81463a,a81464a,a81467a,a81470a,a81471a,a81472a,a81476a,a81477a,a81480a,a81483a,a81484a,a81485a,a81488a,a81491a,a81492a,a81495a,a81498a,a81499a,a81500a,a81504a,a81505a,a81508a,a81511a,a81512a,a81513a,a81516a,a81519a,a81520a,a81523a,a81526a,a81527a,a81528a,a81532a,a81533a,a81536a,a81539a,a81540a,a81541a,a81544a,a81547a,a81548a,a81551a,a81554a,a81555a,a81556a,a81560a,a81561a,a81564a,a81567a,a81568a,a81569a,a81572a,a81575a,a81576a,a81579a,a81582a,a81583a,a81584a,a81588a,a81589a,a81592a,a81595a,a81596a,a81597a,a81600a,a81603a,a81604a,a81607a,a81610a,a81611a,a81612a,a81616a,a81617a,a81620a,a81623a,a81624a,a81625a,a81628a,a81631a,a81632a,a81635a,a81638a,a81639a,a81640a,a81644a,a81645a,a81648a,a81651a,a81652a,a81653a,a81656a,a81659a,a81660a,a81663a,a81666a,a81667a,a81668a,a81672a,a81673a,a81676a,a81679a,a81680a,a81681a,a81684a,a81687a,a81688a,a81691a,a81694a,a81695a,a81696a,a81700a,a81701a,a81704a,a81707a,a81708a,a81709a,a81712a,a81715a,a81716a,a81719a,a81722a,a81723a,a81724a,a81728a,a81729a,a81732a,a81735a,a81736a,a81737a,a81740a,a81743a,a81744a,a81747a,a81750a,a81751a,a81752a,a81756a,a81757a,a81760a,a81763a,a81764a,a81765a,a81768a,a81771a,a81772a,a81775a,a81778a,a81779a,a81780a,a81784a,a81785a,a81788a,a81791a,a81792a,a81793a,a81796a,a81799a,a81800a,a81803a,a81806a,a81807a,a81808a,a81812a,a81813a,a81816a,a81819a,a81820a,a81821a,a81824a,a81827a,a81828a,a81831a,a81834a,a81835a,a81836a,a81840a,a81841a,a81844a,a81847a,a81848a,a81849a,a81852a,a81855a,a81856a,a81859a,a81862a,a81863a,a81864a,a81868a,a81869a,a81872a,a81875a,a81876a,a81877a,a81880a,a81883a,a81884a,a81887a,a81890a,a81891a,a81892a,a81896a,a81897a,a81900a,a81903a,a81904a,a81905a,a81908a,a81911a,a81912a,a81915a,a81918a,a81919a,a81920a,a81924a,a81925a,a81928a,a81931a,a81932a,a81933a,a81936a,a81939a,a81940a,a81943a,a81946a,a81947a,a81948a,a81952a,a81953a,a81956a,a81959a,a81960a,a81961a,a81964a,a81967a,a81968a,a81971a,a81974a,a81975a,a81976a,a81980a,a81981a,a81984a,a81987a,a81988a,a81989a,a81992a,a81995a,a81996a,a81999a,a82002a,a82003a,a82004a,a82008a,a82009a,a82012a,a82015a,a82016a,a82017a,a82020a,a82023a,a82024a,a82027a,a82030a,a82031a,a82032a,a82036a,a82037a,a82040a,a82043a,a82044a,a82045a,a82048a,a82051a,a82052a,a82055a,a82058a,a82059a,a82060a,a82064a,a82065a,a82068a,a82071a,a82072a,a82073a,a82076a,a82079a,a82080a,a82083a,a82086a,a82087a,a82088a,a82092a,a82093a,a82096a,a82099a,a82100a,a82101a,a82104a,a82107a,a82108a,a82111a,a82114a,a82115a,a82116a,a82120a,a82121a,a82124a,a82127a,a82128a,a82129a,a82132a,a82135a,a82136a,a82139a,a82142a,a82143a,a82144a,a82148a,a82149a,a82152a,a82155a,a82156a,a82157a,a82160a,a82163a,a82164a,a82167a,a82170a,a82171a,a82172a,a82176a,a82177a,a82180a,a82183a,a82184a,a82185a,a82188a,a82191a,a82192a,a82195a,a82198a,a82199a,a82200a,a82204a,a82205a,a82208a,a82211a,a82212a,a82213a,a82216a,a82219a,a82220a,a82223a,a82226a,a82227a,a82228a,a82232a,a82233a,a82236a,a82239a,a82240a,a82241a,a82244a,a82247a,a82248a,a82251a,a82254a,a82255a,a82256a,a82260a,a82261a,a82264a,a82267a,a82268a,a82269a,a82272a,a82275a,a82276a,a82279a,a82282a,a82283a,a82284a,a82288a,a82289a,a82292a,a82295a,a82296a,a82297a,a82300a,a82303a,a82304a,a82307a,a82310a,a82311a,a82312a,a82316a,a82317a,a82320a,a82323a,a82324a,a82325a,a82328a,a82331a,a82332a,a82335a,a82338a,a82339a,a82340a,a82344a,a82345a,a82348a,a82351a,a82352a,a82353a,a82356a,a82359a,a82360a,a82363a,a82366a,a82367a,a82368a,a82372a,a82373a,a82376a,a82379a,a82380a,a82381a,a82384a,a82387a,a82388a,a82391a,a82394a,a82395a,a82396a,a82400a,a82401a,a82404a,a82407a,a82408a,a82409a,a82412a,a82415a,a82416a,a82419a,a82422a,a82423a,a82424a,a82428a,a82429a,a82432a,a82435a,a82436a,a82437a,a82440a,a82443a,a82444a,a82447a,a82450a,a82451a,a82452a,a82456a,a82457a,a82460a,a82463a,a82464a,a82465a,a82468a,a82471a,a82472a,a82475a,a82478a,a82479a,a82480a,a82484a,a82485a,a82488a,a82491a,a82492a,a82493a,a82496a,a82499a,a82500a,a82503a,a82506a,a82507a,a82508a,a82512a,a82513a,a82516a,a82519a,a82520a,a82521a,a82524a,a82527a,a82528a,a82531a,a82534a,a82535a,a82536a,a82540a,a82541a,a82544a,a82547a,a82548a,a82549a,a82552a,a82555a,a82556a,a82559a,a82562a,a82563a,a82564a,a82568a,a82569a,a82572a,a82575a,a82576a,a82577a,a82580a,a82583a,a82584a,a82587a,a82590a,a82591a,a82592a,a82596a,a82597a,a82600a,a82603a,a82604a,a82605a,a82608a,a82611a,a82612a,a82615a,a82618a,a82619a,a82620a,a82624a,a82625a,a82628a,a82631a,a82632a,a82633a,a82636a,a82639a,a82640a,a82643a,a82646a,a82647a,a82648a,a82652a,a82653a,a82656a,a82659a,a82660a,a82661a,a82664a,a82667a,a82668a,a82671a,a82674a,a82675a,a82676a,a82680a,a82681a,a82684a,a82687a,a82688a,a82689a,a82692a,a82695a,a82696a,a82699a,a82702a,a82703a,a82704a,a82708a,a82709a,a82712a,a82715a,a82716a,a82717a,a82720a,a82723a,a82724a,a82727a,a82730a,a82731a,a82732a,a82736a,a82737a,a82740a,a82743a,a82744a,a82745a,a82748a,a82751a,a82752a,a82755a,a82758a,a82759a,a82760a,a82764a,a82765a,a82768a,a82771a,a82772a,a82773a,a82776a,a82779a,a82780a,a82783a,a82786a,a82787a,a82788a,a82792a,a82793a,a82796a,a82799a,a82800a,a82801a,a82804a,a82807a,a82808a,a82811a,a82814a,a82815a,a82816a,a82820a,a82821a,a82824a,a82827a,a82828a,a82829a,a82832a,a82835a,a82836a,a82839a,a82842a,a82843a,a82844a,a82848a,a82849a,a82852a,a82855a,a82856a,a82857a,a82860a,a82863a,a82864a,a82867a,a82870a,a82871a,a82872a,a82876a,a82877a,a82880a,a82883a,a82884a,a82885a,a82888a,a82891a,a82892a,a82895a,a82898a,a82899a,a82900a,a82904a,a82905a,a82908a,a82911a,a82912a,a82913a,a82916a,a82919a,a82920a,a82923a,a82926a,a82927a,a82928a,a82932a,a82933a,a82936a,a82939a,a82940a,a82941a,a82944a,a82947a,a82948a,a82951a,a82954a,a82955a,a82956a,a82960a,a82961a,a82964a,a82967a,a82968a,a82969a,a82972a,a82975a,a82976a,a82979a,a82982a,a82983a,a82984a,a82988a,a82989a,a82992a,a82995a,a82996a,a82997a,a83000a,a83003a,a83004a,a83007a,a83010a,a83011a,a83012a,a83016a,a83017a,a83020a,a83023a,a83024a,a83025a,a83028a,a83031a,a83032a,a83035a,a83038a,a83039a,a83040a,a83044a,a83045a,a83048a,a83051a,a83052a,a83053a,a83056a,a83059a,a83060a,a83063a,a83066a,a83067a,a83068a,a83072a,a83073a,a83076a,a83079a,a83080a,a83081a,a83084a,a83087a,a83088a,a83091a,a83094a,a83095a,a83096a,a83100a,a83101a,a83104a,a83107a,a83108a,a83109a,a83112a,a83115a,a83116a,a83119a,a83122a,a83123a,a83124a,a83128a,a83129a,a83132a,a83135a,a83136a,a83137a,a83140a,a83143a,a83144a,a83147a,a83150a,a83151a,a83152a,a83156a,a83157a,a83160a,a83163a,a83164a,a83165a,a83168a,a83171a,a83172a,a83175a,a83178a,a83179a,a83180a,a83184a,a83185a,a83188a,a83191a,a83192a,a83193a,a83196a,a83199a,a83200a,a83203a,a83206a,a83207a,a83208a,a83212a,a83213a,a83216a,a83219a,a83220a,a83221a,a83224a,a83227a,a83228a,a83231a,a83234a,a83235a,a83236a,a83240a,a83241a,a83244a,a83247a,a83248a,a83249a,a83252a,a83255a,a83256a,a83259a,a83262a,a83263a,a83264a,a83268a,a83269a,a83272a,a83275a,a83276a,a83277a,a83280a,a83283a,a83284a,a83287a,a83290a,a83291a,a83292a,a83296a,a83297a,a83300a,a83303a,a83304a,a83305a,a83308a,a83311a,a83312a,a83315a,a83318a,a83319a,a83320a,a83324a,a83325a,a83328a,a83331a,a83332a,a83333a,a83336a,a83339a,a83340a,a83343a,a83346a,a83347a,a83348a,a83352a,a83353a,a83356a,a83359a,a83360a,a83361a,a83364a,a83367a,a83368a,a83371a,a83374a,a83375a,a83376a,a83380a,a83381a,a83384a,a83387a,a83388a,a83389a,a83392a,a83395a,a83396a,a83399a,a83402a,a83403a,a83404a,a83408a,a83409a,a83412a,a83415a,a83416a,a83417a,a83420a,a83423a,a83424a,a83427a,a83430a,a83431a,a83432a,a83436a,a83437a,a83440a,a83443a,a83444a,a83445a,a83448a,a83451a,a83452a,a83455a,a83458a,a83459a,a83460a,a83464a,a83465a,a83468a,a83471a,a83472a,a83473a,a83476a,a83479a,a83480a,a83483a,a83486a,a83487a,a83488a,a83492a,a83493a,a83496a,a83499a,a83500a,a83501a,a83504a,a83507a,a83508a,a83511a,a83514a,a83515a,a83516a,a83520a,a83521a,a83524a,a83527a,a83528a,a83529a,a83532a,a83535a,a83536a,a83539a,a83542a,a83543a,a83544a,a83548a,a83549a,a83552a,a83555a,a83556a,a83557a,a83560a,a83563a,a83564a,a83567a,a83570a,a83571a,a83572a,a83576a,a83577a,a83580a,a83583a,a83584a,a83585a,a83588a,a83591a,a83592a,a83595a,a83598a,a83599a,a83600a,a83604a,a83605a,a83608a,a83611a,a83612a,a83613a,a83616a,a83619a,a83620a,a83623a,a83626a,a83627a,a83628a,a83632a,a83633a,a83636a,a83639a,a83640a,a83641a,a83644a,a83647a,a83648a,a83651a,a83654a,a83655a,a83656a,a83660a,a83661a,a83664a,a83667a,a83668a,a83669a,a83672a,a83675a,a83676a,a83679a,a83682a,a83683a,a83684a,a83688a,a83689a,a83692a,a83695a,a83696a,a83697a,a83700a,a83703a,a83704a,a83707a,a83710a,a83711a,a83712a,a83716a,a83717a,a83720a,a83723a,a83724a,a83725a,a83728a,a83731a,a83732a,a83735a,a83738a,a83739a,a83740a,a83744a,a83745a,a83748a,a83751a,a83752a,a83753a,a83756a,a83759a,a83760a,a83763a,a83766a,a83767a,a83768a,a83772a,a83773a,a83776a,a83779a,a83780a,a83781a,a83784a,a83787a,a83788a,a83791a,a83794a,a83795a,a83796a,a83800a,a83801a,a83804a,a83807a,a83808a,a83809a,a83812a,a83815a,a83816a,a83819a,a83822a,a83823a,a83824a,a83828a,a83829a,a83832a,a83835a,a83836a,a83837a,a83840a,a83843a,a83844a,a83847a,a83850a,a83851a,a83852a,a83856a,a83857a,a83860a,a83863a,a83864a,a83865a,a83868a,a83871a,a83872a,a83875a,a83878a,a83879a,a83880a,a83884a,a83885a,a83888a,a83891a,a83892a,a83893a,a83896a,a83899a,a83900a,a83903a,a83906a,a83907a,a83908a,a83912a,a83913a,a83916a,a83919a,a83920a,a83921a,a83924a,a83927a,a83928a,a83931a,a83934a,a83935a,a83936a,a83940a,a83941a,a83944a,a83947a,a83948a,a83949a,a83952a,a83955a,a83956a,a83959a,a83962a,a83963a,a83964a,a83968a,a83969a,a83972a,a83975a,a83976a,a83977a,a83980a,a83983a,a83984a,a83987a,a83990a,a83991a,a83992a,a83996a,a83997a,a84000a,a84003a,a84004a,a84005a,a84008a,a84011a,a84012a,a84015a,a84018a,a84019a,a84020a,a84024a,a84025a,a84028a,a84031a,a84032a,a84033a,a84036a,a84039a,a84040a,a84043a,a84046a,a84047a,a84048a,a84052a,a84053a,a84056a,a84059a,a84060a,a84061a,a84064a,a84067a,a84068a,a84071a,a84074a,a84075a,a84076a,a84080a,a84081a,a84084a,a84087a,a84088a,a84089a,a84092a,a84095a,a84096a,a84099a,a84102a,a84103a,a84104a,a84108a,a84109a,a84112a,a84115a,a84116a,a84117a,a84120a,a84123a,a84124a,a84127a,a84130a,a84131a,a84132a,a84136a,a84137a,a84140a,a84143a,a84144a,a84145a,a84148a,a84151a,a84152a,a84155a,a84158a,a84159a,a84160a,a84164a,a84165a,a84168a,a84171a,a84172a,a84173a,a84176a,a84179a,a84180a,a84183a,a84186a,a84187a,a84188a,a84192a,a84193a,a84196a,a84199a,a84200a,a84201a,a84204a,a84207a,a84208a,a84211a,a84214a,a84215a,a84216a,a84220a,a84221a,a84224a,a84227a,a84228a,a84229a,a84232a,a84235a,a84236a,a84239a,a84242a,a84243a,a84244a,a84248a,a84249a,a84252a,a84255a,a84256a,a84257a,a84260a,a84263a,a84264a,a84267a,a84270a,a84271a,a84272a,a84276a,a84277a,a84280a,a84283a,a84284a,a84285a,a84288a,a84291a,a84292a,a84295a,a84298a,a84299a,a84300a,a84304a,a84305a,a84308a,a84311a,a84312a,a84313a,a84316a,a84319a,a84320a,a84323a,a84326a,a84327a,a84328a,a84332a,a84333a,a84336a,a84339a,a84340a,a84341a,a84344a,a84347a,a84348a,a84351a,a84354a,a84355a,a84356a,a84360a,a84361a,a84364a,a84367a,a84368a,a84369a,a84372a,a84375a,a84376a,a84379a,a84382a,a84383a,a84384a,a84388a,a84389a,a84392a,a84395a,a84396a,a84397a,a84400a,a84403a,a84404a,a84407a,a84410a,a84411a,a84412a,a84416a,a84417a,a84420a,a84423a,a84424a,a84425a,a84428a,a84431a,a84432a,a84435a,a84438a,a84439a,a84440a,a84444a,a84445a,a84448a,a84451a,a84452a,a84453a,a84456a,a84459a,a84460a,a84463a,a84466a,a84467a,a84468a,a84472a,a84473a,a84476a,a84479a,a84480a,a84481a,a84484a,a84487a,a84488a,a84491a,a84494a,a84495a,a84496a,a84500a,a84501a,a84504a,a84507a,a84508a,a84509a,a84512a,a84515a,a84516a,a84519a,a84522a,a84523a,a84524a,a84528a,a84529a,a84532a,a84535a,a84536a,a84537a,a84540a,a84543a,a84544a,a84547a,a84550a,a84551a,a84552a,a84556a,a84557a,a84560a,a84563a,a84564a,a84565a,a84568a,a84571a,a84572a,a84575a,a84578a,a84579a,a84580a,a84584a,a84585a,a84588a,a84591a,a84592a,a84593a,a84596a,a84599a,a84600a,a84603a,a84606a,a84607a,a84608a,a84612a,a84613a,a84616a,a84619a,a84620a,a84621a,a84624a,a84627a,a84628a,a84631a,a84634a,a84635a,a84636a,a84640a,a84641a,a84644a,a84647a,a84648a,a84649a,a84652a,a84655a,a84656a,a84659a,a84662a,a84663a,a84664a,a84668a,a84669a,a84672a,a84675a,a84676a,a84677a,a84680a,a84683a,a84684a,a84687a,a84690a,a84691a,a84692a,a84696a,a84697a,a84700a,a84703a,a84704a,a84705a,a84708a,a84711a,a84712a,a84715a,a84718a,a84719a,a84720a,a84724a,a84725a,a84728a,a84731a,a84732a,a84733a,a84736a,a84739a,a84740a,a84743a,a84746a,a84747a,a84748a,a84752a,a84753a,a84756a,a84759a,a84760a,a84761a,a84764a,a84767a,a84768a,a84771a,a84774a,a84775a,a84776a,a84780a,a84781a,a84784a,a84787a,a84788a,a84789a,a84792a,a84795a,a84796a,a84799a,a84802a,a84803a,a84804a,a84808a,a84809a,a84812a,a84815a,a84816a,a84817a,a84820a,a84823a,a84824a,a84827a,a84830a,a84831a,a84832a,a84836a,a84837a,a84840a,a84843a,a84844a,a84845a,a84848a,a84851a,a84852a,a84855a,a84858a,a84859a,a84860a,a84864a,a84865a,a84868a,a84871a,a84872a,a84873a,a84876a,a84879a,a84880a,a84883a,a84886a,a84887a,a84888a,a84892a,a84893a,a84896a,a84899a,a84900a,a84901a,a84904a,a84907a,a84908a,a84911a,a84914a,a84915a,a84916a,a84920a,a84921a,a84924a,a84927a,a84928a,a84929a,a84932a,a84935a,a84936a,a84939a,a84942a,a84943a,a84944a,a84948a,a84949a,a84952a,a84955a,a84956a,a84957a,a84960a,a84963a,a84964a,a84967a,a84970a,a84971a,a84972a,a84976a,a84977a,a84980a,a84983a,a84984a,a84985a,a84988a,a84991a,a84992a,a84995a,a84998a,a84999a,a85000a,a85004a,a85005a,a85008a,a85011a,a85012a,a85013a,a85016a,a85019a,a85020a,a85023a,a85026a,a85027a,a85028a,a85032a,a85033a,a85036a,a85039a,a85040a,a85041a,a85044a,a85047a,a85048a,a85051a,a85054a,a85055a,a85056a,a85060a,a85061a,a85064a,a85067a,a85068a,a85069a,a85072a,a85075a,a85076a,a85079a,a85082a,a85083a,a85084a,a85088a,a85089a,a85092a,a85095a,a85096a,a85097a,a85100a,a85103a,a85104a,a85107a,a85110a,a85111a,a85112a,a85116a,a85117a,a85120a,a85123a,a85124a,a85125a,a85128a,a85131a,a85132a,a85135a,a85138a,a85139a,a85140a,a85144a,a85145a,a85148a,a85151a,a85152a,a85153a,a85156a,a85159a,a85160a,a85163a,a85166a,a85167a,a85168a,a85172a,a85173a,a85176a,a85179a,a85180a,a85181a,a85184a,a85187a,a85188a,a85191a,a85194a,a85195a,a85196a,a85200a,a85201a,a85204a,a85207a,a85208a,a85209a,a85212a,a85215a,a85216a,a85219a,a85222a,a85223a,a85224a,a85228a,a85229a,a85232a,a85235a,a85236a,a85237a,a85240a,a85243a,a85244a,a85247a,a85250a,a85251a,a85252a,a85256a,a85257a,a85260a,a85263a,a85264a,a85265a,a85268a,a85271a,a85272a,a85275a,a85278a,a85279a,a85280a,a85284a,a85285a,a85288a,a85291a,a85292a,a85293a,a85296a,a85299a,a85300a,a85303a,a85306a,a85307a,a85308a,a85312a,a85313a,a85316a,a85319a,a85320a,a85321a,a85324a,a85327a,a85328a,a85331a,a85334a,a85335a,a85336a,a85340a,a85341a,a85344a,a85347a,a85348a,a85349a,a85352a,a85355a,a85356a,a85359a,a85362a,a85363a,a85364a,a85368a,a85369a,a85372a,a85375a,a85376a,a85377a,a85380a,a85383a,a85384a,a85387a,a85390a,a85391a,a85392a,a85396a,a85397a,a85400a,a85403a,a85404a,a85405a,a85408a,a85411a,a85412a,a85415a,a85418a,a85419a,a85420a,a85424a,a85425a,a85428a,a85431a,a85432a,a85433a,a85436a,a85439a,a85440a,a85443a,a85446a,a85447a,a85448a,a85452a,a85453a,a85456a,a85459a,a85460a,a85461a,a85464a,a85467a,a85468a,a85471a,a85474a,a85475a,a85476a,a85480a,a85481a,a85484a,a85487a,a85488a,a85489a,a85492a,a85495a,a85496a,a85499a,a85502a,a85503a,a85504a,a85508a,a85509a,a85512a,a85515a,a85516a,a85517a,a85520a,a85523a,a85524a,a85527a,a85530a,a85531a,a85532a,a85536a,a85537a,a85540a,a85543a,a85544a,a85545a,a85548a,a85551a,a85552a,a85555a,a85558a,a85559a,a85560a,a85564a,a85565a,a85568a,a85571a,a85572a,a85573a,a85576a,a85579a,a85580a,a85583a,a85586a,a85587a,a85588a,a85592a,a85593a,a85596a,a85599a,a85600a,a85601a,a85604a,a85607a,a85608a,a85611a,a85614a,a85615a,a85616a,a85620a,a85621a,a85624a,a85627a,a85628a,a85629a,a85632a,a85635a,a85636a,a85639a,a85642a,a85643a,a85644a,a85648a,a85649a,a85652a,a85655a,a85656a,a85657a,a85660a,a85663a,a85664a,a85667a,a85670a,a85671a,a85672a,a85676a,a85677a,a85680a,a85683a,a85684a,a85685a,a85688a,a85691a,a85692a,a85695a,a85698a,a85699a,a85700a,a85704a,a85705a,a85708a,a85711a,a85712a,a85713a,a85716a,a85719a,a85720a,a85723a,a85726a,a85727a,a85728a,a85732a,a85733a,a85736a,a85739a,a85740a,a85741a,a85744a,a85747a,a85748a,a85751a,a85754a,a85755a,a85756a,a85760a,a85761a,a85764a,a85767a,a85768a,a85769a,a85772a,a85775a,a85776a,a85779a,a85782a,a85783a,a85784a,a85788a,a85789a,a85792a,a85795a,a85796a,a85797a,a85800a,a85803a,a85804a,a85807a,a85810a,a85811a,a85812a,a85816a,a85817a,a85820a,a85823a,a85824a,a85825a,a85828a,a85831a,a85832a,a85835a,a85838a,a85839a,a85840a,a85844a,a85845a,a85848a,a85851a,a85852a,a85853a,a85856a,a85859a,a85860a,a85863a,a85866a,a85867a,a85868a,a85872a,a85873a,a85876a,a85879a,a85880a,a85881a,a85884a,a85887a,a85888a,a85891a,a85894a,a85895a,a85896a,a85900a,a85901a,a85904a,a85907a,a85908a,a85909a,a85912a,a85915a,a85916a,a85919a,a85922a,a85923a,a85924a,a85928a,a85929a,a85932a,a85935a,a85936a,a85937a,a85940a,a85943a,a85944a,a85947a,a85950a,a85951a,a85952a,a85956a,a85957a,a85960a,a85963a,a85964a,a85965a,a85968a,a85971a,a85972a,a85975a,a85978a,a85979a,a85980a,a85984a,a85985a,a85988a,a85991a,a85992a,a85993a,a85996a,a85999a,a86000a,a86003a,a86006a,a86007a,a86008a,a86012a,a86013a,a86016a,a86019a,a86020a,a86021a,a86024a,a86027a,a86028a,a86031a,a86034a,a86035a,a86036a,a86040a,a86041a,a86044a,a86047a,a86048a,a86049a,a86052a,a86055a,a86056a,a86059a,a86062a,a86063a,a86064a,a86068a,a86069a,a86072a,a86075a,a86076a,a86077a,a86080a,a86083a,a86084a,a86087a,a86090a,a86091a,a86092a,a86096a,a86097a,a86100a,a86103a,a86104a,a86105a,a86108a,a86111a,a86112a,a86115a,a86118a,a86119a,a86120a,a86124a,a86125a,a86128a,a86131a,a86132a,a86133a,a86136a,a86139a,a86140a,a86143a,a86146a,a86147a,a86148a,a86152a,a86153a,a86156a,a86159a,a86160a,a86161a,a86164a,a86167a,a86168a,a86171a,a86174a,a86175a,a86176a,a86180a,a86181a,a86184a,a86187a,a86188a,a86189a,a86192a,a86195a,a86196a,a86199a,a86202a,a86203a,a86204a,a86208a,a86209a,a86212a,a86215a,a86216a,a86217a,a86220a,a86223a,a86224a,a86227a,a86230a,a86231a,a86232a,a86236a,a86237a,a86240a,a86243a,a86244a,a86245a,a86248a,a86251a,a86252a,a86255a,a86258a,a86259a,a86260a,a86264a,a86265a,a86268a,a86271a,a86272a,a86273a,a86276a,a86279a,a86280a,a86283a,a86286a,a86287a,a86288a,a86292a,a86293a,a86296a,a86299a,a86300a,a86301a,a86304a,a86307a,a86308a,a86311a,a86314a,a86315a,a86316a,a86320a,a86321a,a86324a,a86327a,a86328a,a86329a,a86332a,a86335a,a86336a,a86339a,a86342a,a86343a,a86344a,a86348a,a86349a,a86352a,a86355a,a86356a,a86357a,a86360a,a86363a,a86364a,a86367a,a86370a,a86371a,a86372a,a86376a,a86377a,a86380a,a86383a,a86384a,a86385a,a86388a,a86391a,a86392a,a86395a,a86398a,a86399a,a86400a,a86404a,a86405a,a86408a,a86411a,a86412a,a86413a,a86416a,a86419a,a86420a,a86423a,a86426a,a86427a,a86428a,a86432a,a86433a,a86436a,a86439a,a86440a,a86441a,a86444a,a86447a,a86448a,a86451a,a86454a,a86455a,a86456a,a86460a,a86461a,a86464a,a86467a,a86468a,a86469a,a86472a,a86475a,a86476a,a86479a,a86482a,a86483a,a86484a,a86488a,a86489a,a86492a,a86495a,a86496a,a86497a,a86500a,a86503a,a86504a,a86507a,a86510a,a86511a,a86512a,a86516a,a86517a,a86520a,a86523a,a86524a,a86525a,a86528a,a86531a,a86532a,a86535a,a86538a,a86539a,a86540a,a86544a,a86545a,a86548a,a86551a,a86552a,a86553a,a86556a,a86559a,a86560a,a86563a,a86566a,a86567a,a86568a,a86572a,a86573a,a86576a,a86579a,a86580a,a86581a,a86584a,a86587a,a86588a,a86591a,a86594a,a86595a,a86596a,a86600a,a86601a,a86604a,a86607a,a86608a,a86609a,a86612a,a86615a,a86616a,a86619a,a86622a,a86623a,a86624a,a86628a,a86629a,a86632a,a86635a,a86636a,a86637a,a86640a,a86643a,a86644a,a86647a,a86650a,a86651a,a86652a,a86656a,a86657a,a86660a,a86663a,a86664a,a86665a,a86668a,a86671a,a86672a,a86675a,a86678a,a86679a,a86680a,a86684a,a86685a,a86688a,a86691a,a86692a,a86693a,a86696a,a86699a,a86700a,a86703a,a86706a,a86707a,a86708a,a86712a,a86713a,a86716a,a86719a,a86720a,a86721a,a86724a,a86727a,a86728a,a86731a,a86734a,a86735a,a86736a,a86740a,a86741a,a86744a,a86747a,a86748a,a86749a,a86752a,a86755a,a86756a,a86759a,a86762a,a86763a,a86764a,a86768a,a86769a,a86772a,a86775a,a86776a,a86777a,a86780a,a86783a,a86784a,a86787a,a86790a,a86791a,a86792a,a86796a,a86797a,a86800a,a86803a,a86804a,a86805a,a86808a,a86811a,a86812a,a86815a,a86818a,a86819a,a86820a,a86824a,a86825a,a86828a,a86831a,a86832a,a86833a,a86836a,a86839a,a86840a,a86843a,a86846a,a86847a,a86848a,a86852a,a86853a,a86856a,a86859a,a86860a,a86861a,a86864a,a86867a,a86868a,a86871a,a86874a,a86875a,a86876a,a86880a,a86881a,a86884a,a86887a,a86888a,a86889a,a86892a,a86895a,a86896a,a86899a,a86902a,a86903a,a86904a,a86908a,a86909a,a86912a,a86915a,a86916a,a86917a,a86920a,a86923a,a86924a,a86927a,a86930a,a86931a,a86932a,a86936a,a86937a,a86940a,a86943a,a86944a,a86945a,a86948a,a86951a,a86952a,a86955a,a86958a,a86959a,a86960a,a86964a,a86965a,a86968a,a86971a,a86972a,a86973a,a86976a,a86979a,a86980a,a86983a,a86986a,a86987a,a86988a,a86992a,a86993a,a86996a,a86999a,a87000a,a87001a,a87004a,a87007a,a87008a,a87011a,a87014a,a87015a,a87016a,a87020a,a87021a,a87024a,a87027a,a87028a,a87029a,a87032a,a87035a,a87036a,a87039a,a87042a,a87043a,a87044a,a87048a,a87049a,a87052a,a87055a,a87056a,a87057a,a87060a,a87063a,a87064a,a87067a,a87070a,a87071a,a87072a,a87076a,a87077a,a87080a,a87083a,a87084a,a87085a,a87088a,a87091a,a87092a,a87095a,a87098a,a87099a,a87100a,a87104a,a87105a,a87108a,a87111a,a87112a,a87113a,a87116a,a87119a,a87120a,a87123a,a87126a,a87127a,a87128a,a87132a,a87133a,a87136a,a87139a,a87140a,a87141a,a87144a,a87147a,a87148a,a87151a,a87154a,a87155a,a87156a,a87160a,a87161a,a87164a,a87167a,a87168a,a87169a,a87172a,a87175a,a87176a,a87179a,a87182a,a87183a,a87184a,a87188a,a87189a,a87192a,a87195a,a87196a,a87197a,a87200a,a87203a,a87204a,a87207a,a87210a,a87211a,a87212a,a87216a,a87217a,a87220a,a87223a,a87224a,a87225a,a87228a,a87231a,a87232a,a87235a,a87238a,a87239a,a87240a,a87244a,a87245a,a87248a,a87251a,a87252a,a87253a,a87256a,a87259a,a87260a,a87263a,a87266a,a87267a,a87268a,a87272a,a87273a,a87276a,a87279a,a87280a,a87281a,a87284a,a87287a,a87288a,a87291a,a87294a,a87295a,a87296a,a87300a,a87301a,a87304a,a87307a,a87308a,a87309a,a87312a,a87315a,a87316a,a87319a,a87322a,a87323a,a87324a,a87328a,a87329a,a87332a,a87335a,a87336a,a87337a,a87340a,a87343a,a87344a,a87347a,a87350a,a87351a,a87352a,a87356a,a87357a,a87360a,a87363a,a87364a,a87365a,a87368a,a87371a,a87372a,a87375a,a87378a,a87379a,a87380a,a87384a,a87385a,a87388a,a87391a,a87392a,a87393a,a87396a,a87399a,a87400a,a87403a,a87406a,a87407a,a87408a,a87412a,a87413a,a87416a,a87419a,a87420a,a87421a,a87424a,a87427a,a87428a,a87431a,a87434a,a87435a,a87436a,a87440a,a87441a,a87444a,a87447a,a87448a,a87449a,a87452a,a87455a,a87456a,a87459a,a87462a,a87463a,a87464a,a87468a,a87469a,a87472a,a87475a,a87476a,a87477a,a87480a,a87483a,a87484a,a87487a,a87490a,a87491a,a87492a,a87496a,a87497a,a87500a,a87503a,a87504a,a87505a,a87508a,a87511a,a87512a,a87515a,a87518a,a87519a,a87520a,a87524a,a87525a,a87528a,a87531a,a87532a,a87533a,a87536a,a87539a,a87540a,a87543a,a87546a,a87547a,a87548a,a87552a,a87553a,a87556a,a87559a,a87560a,a87561a,a87564a,a87567a,a87568a,a87571a,a87574a,a87575a,a87576a,a87580a,a87581a,a87584a,a87587a,a87588a,a87589a,a87592a,a87595a,a87596a,a87599a,a87602a,a87603a,a87604a,a87608a,a87609a,a87612a,a87615a,a87616a,a87617a,a87620a,a87623a,a87624a,a87627a,a87630a,a87631a,a87632a,a87636a,a87637a,a87640a,a87643a,a87644a,a87645a,a87648a,a87651a,a87652a,a87655a,a87658a,a87659a,a87660a,a87664a,a87665a,a87668a,a87671a,a87672a,a87673a,a87676a,a87679a,a87680a,a87683a,a87686a,a87687a,a87688a,a87692a,a87693a,a87696a,a87699a,a87700a,a87701a,a87704a,a87707a,a87708a,a87711a,a87714a,a87715a,a87716a,a87720a,a87721a,a87724a,a87727a,a87728a,a87729a,a87732a,a87735a,a87736a,a87739a,a87742a,a87743a,a87744a,a87748a,a87749a,a87752a,a87755a,a87756a,a87757a,a87760a,a87763a,a87764a,a87767a,a87770a,a87771a,a87772a,a87776a,a87777a,a87780a,a87783a,a87784a,a87785a,a87788a,a87791a,a87792a,a87795a,a87798a,a87799a,a87800a,a87804a,a87805a,a87808a,a87811a,a87812a,a87813a,a87816a,a87819a,a87820a,a87823a,a87826a,a87827a,a87828a,a87832a,a87833a,a87836a,a87839a,a87840a,a87841a,a87844a,a87847a,a87848a,a87851a,a87854a,a87855a,a87856a,a87860a,a87861a,a87864a,a87867a,a87868a,a87869a,a87872a,a87875a,a87876a,a87879a,a87882a,a87883a,a87884a,a87888a,a87889a,a87892a,a87895a,a87896a,a87897a,a87900a,a87903a,a87904a,a87907a,a87910a,a87911a,a87912a,a87916a,a87917a,a87920a,a87923a,a87924a,a87925a,a87928a,a87931a,a87932a,a87935a,a87938a,a87939a,a87940a,a87944a,a87945a,a87948a,a87951a,a87952a,a87953a,a87956a,a87959a,a87960a,a87963a,a87966a,a87967a,a87968a,a87972a,a87973a,a87976a,a87979a,a87980a,a87981a,a87984a,a87987a,a87988a,a87991a,a87994a,a87995a,a87996a,a88000a,a88001a,a88004a,a88007a,a88008a,a88009a,a88012a,a88015a,a88016a,a88019a,a88022a,a88023a,a88024a,a88028a,a88029a,a88032a,a88035a,a88036a,a88037a,a88040a,a88043a,a88044a,a88047a,a88050a,a88051a,a88052a,a88056a,a88057a,a88060a,a88063a,a88064a,a88065a,a88068a,a88071a,a88072a,a88075a,a88078a,a88079a,a88080a,a88084a,a88085a,a88088a,a88091a,a88092a,a88093a,a88096a,a88099a,a88100a,a88103a,a88106a,a88107a,a88108a,a88112a,a88113a,a88116a,a88119a,a88120a,a88121a,a88124a,a88127a,a88128a,a88131a,a88134a,a88135a,a88136a,a88140a,a88141a,a88144a,a88147a,a88148a,a88149a,a88152a,a88155a,a88156a,a88159a,a88162a,a88163a,a88164a,a88168a,a88169a,a88172a,a88175a,a88176a,a88177a,a88180a,a88183a,a88184a,a88187a,a88190a,a88191a,a88192a,a88196a,a88197a,a88200a,a88203a,a88204a,a88205a,a88208a,a88211a,a88212a,a88215a,a88218a,a88219a,a88220a,a88224a,a88225a,a88228a,a88231a,a88232a,a88233a,a88236a,a88239a,a88240a,a88243a,a88246a,a88247a,a88248a,a88252a,a88253a,a88256a,a88259a,a88260a,a88261a,a88264a,a88267a,a88268a,a88271a,a88274a,a88275a,a88276a,a88280a,a88281a,a88284a,a88287a,a88288a,a88289a,a88292a,a88295a,a88296a,a88299a,a88302a,a88303a,a88304a,a88308a,a88309a,a88312a,a88315a,a88316a,a88317a,a88320a,a88323a,a88324a,a88327a,a88330a,a88331a,a88332a,a88336a,a88337a,a88340a,a88343a,a88344a,a88345a,a88348a,a88351a,a88352a,a88355a,a88358a,a88359a,a88360a,a88364a,a88365a,a88368a,a88371a,a88372a,a88373a,a88376a,a88379a,a88380a,a88383a,a88386a,a88387a,a88388a,a88392a,a88393a,a88396a,a88399a,a88400a,a88401a,a88404a,a88407a,a88408a,a88411a,a88414a,a88415a,a88416a,a88420a,a88421a,a88424a,a88427a,a88428a,a88429a,a88432a,a88435a,a88436a,a88439a,a88442a,a88443a,a88444a,a88448a,a88449a,a88452a,a88455a,a88456a,a88457a,a88460a,a88463a,a88464a,a88467a,a88470a,a88471a,a88472a,a88476a,a88477a,a88480a,a88483a,a88484a,a88485a,a88488a,a88491a,a88492a,a88495a,a88498a,a88499a,a88500a,a88504a,a88505a,a88508a,a88511a,a88512a,a88513a,a88516a,a88519a,a88520a,a88523a,a88526a,a88527a,a88528a,a88532a,a88533a,a88536a,a88539a,a88540a,a88541a,a88544a,a88547a,a88548a,a88551a,a88554a,a88555a,a88556a,a88560a,a88561a,a88564a,a88567a,a88568a,a88569a,a88572a,a88575a,a88576a,a88579a,a88582a,a88583a,a88584a,a88588a,a88589a,a88592a,a88595a,a88596a,a88597a,a88600a,a88603a,a88604a,a88607a,a88610a,a88611a,a88612a,a88616a,a88617a,a88620a,a88623a,a88624a,a88625a,a88628a,a88631a,a88632a,a88635a,a88638a,a88639a,a88640a,a88644a,a88645a,a88648a,a88651a,a88652a,a88653a,a88656a,a88659a,a88660a,a88663a,a88666a,a88667a,a88668a,a88672a,a88673a,a88676a,a88679a,a88680a,a88681a,a88684a,a88687a,a88688a,a88691a,a88694a,a88695a,a88696a,a88700a,a88701a,a88704a,a88707a,a88708a,a88709a,a88712a,a88715a,a88716a,a88719a,a88722a,a88723a,a88724a,a88728a,a88729a,a88732a,a88735a,a88736a,a88737a,a88740a,a88743a,a88744a,a88747a,a88750a,a88751a,a88752a,a88756a,a88757a,a88760a,a88763a,a88764a,a88765a,a88768a,a88771a,a88772a,a88775a,a88778a,a88779a,a88780a,a88784a,a88785a,a88788a,a88791a,a88792a,a88793a,a88796a,a88799a,a88800a,a88803a,a88806a,a88807a,a88808a,a88812a,a88813a,a88816a,a88819a,a88820a,a88821a,a88824a,a88827a,a88828a,a88831a,a88834a,a88835a,a88836a,a88840a,a88841a,a88844a,a88847a,a88848a,a88849a,a88852a,a88855a,a88856a,a88859a,a88862a,a88863a,a88864a,a88868a,a88869a,a88872a,a88875a,a88876a,a88877a,a88880a,a88883a,a88884a,a88887a,a88890a,a88891a,a88892a,a88896a,a88897a,a88900a,a88903a,a88904a,a88905a,a88908a,a88911a,a88912a,a88915a,a88918a,a88919a,a88920a,a88924a,a88925a,a88928a,a88931a,a88932a,a88933a,a88936a,a88939a,a88940a,a88943a,a88946a,a88947a,a88948a,a88952a,a88953a,a88956a,a88959a,a88960a,a88961a,a88964a,a88967a,a88968a,a88971a,a88974a,a88975a,a88976a,a88980a,a88981a,a88984a,a88987a,a88988a,a88989a,a88992a,a88995a,a88996a,a88999a,a89002a,a89003a,a89004a,a89008a,a89009a,a89012a,a89015a,a89016a,a89017a,a89020a,a89023a,a89024a,a89027a,a89030a,a89031a,a89032a,a89036a,a89037a,a89040a,a89043a,a89044a,a89045a,a89048a,a89051a,a89052a,a89055a,a89058a,a89059a,a89060a,a89064a,a89065a,a89068a,a89071a,a89072a,a89073a,a89076a,a89079a,a89080a,a89083a,a89086a,a89087a,a89088a,a89092a,a89093a,a89096a,a89099a,a89100a,a89101a,a89104a,a89107a,a89108a,a89111a,a89114a,a89115a,a89116a,a89120a,a89121a,a89124a,a89127a,a89128a,a89129a,a89132a,a89135a,a89136a,a89139a,a89142a,a89143a,a89144a,a89148a,a89149a,a89152a,a89155a,a89156a,a89157a,a89160a,a89163a,a89164a,a89167a,a89170a,a89171a,a89172a,a89176a,a89177a,a89180a,a89183a,a89184a,a89185a,a89188a,a89191a,a89192a,a89195a,a89198a,a89199a,a89200a,a89204a,a89205a,a89208a,a89211a,a89212a,a89213a,a89216a,a89219a,a89220a,a89223a,a89226a,a89227a,a89228a,a89232a,a89233a,a89236a,a89239a,a89240a,a89241a,a89244a,a89247a,a89248a,a89251a,a89254a,a89255a,a89256a,a89260a,a89261a,a89264a,a89267a,a89268a,a89269a,a89272a,a89275a,a89276a,a89279a,a89282a,a89283a,a89284a,a89288a,a89289a,a89292a,a89295a,a89296a,a89297a,a89300a,a89303a,a89304a,a89307a,a89310a,a89311a,a89312a,a89316a,a89317a,a89320a,a89323a,a89324a,a89325a,a89328a,a89331a,a89332a,a89335a,a89338a,a89339a,a89340a,a89344a,a89345a,a89348a,a89351a,a89352a,a89353a,a89356a,a89359a,a89360a,a89363a,a89366a,a89367a,a89368a,a89372a,a89373a,a89376a,a89379a,a89380a,a89381a,a89384a,a89387a,a89388a,a89391a,a89394a,a89395a,a89396a,a89400a,a89401a,a89404a,a89407a,a89408a,a89409a,a89412a,a89415a,a89416a,a89419a,a89422a,a89423a,a89424a,a89428a,a89429a,a89432a,a89435a,a89436a,a89437a,a89440a,a89443a,a89444a,a89447a,a89450a,a89451a,a89452a,a89456a,a89457a,a89460a,a89463a,a89464a,a89465a,a89468a,a89471a,a89472a,a89475a,a89478a,a89479a,a89480a,a89484a,a89485a,a89488a,a89491a,a89492a,a89493a,a89496a,a89499a,a89500a,a89503a,a89506a,a89507a,a89508a,a89511a,a89514a,a89515a,a89518a,a89521a,a89522a,a89523a,a89526a,a89529a,a89530a,a89533a,a89536a,a89537a,a89538a,a89541a,a89544a,a89545a,a89548a,a89551a,a89552a,a89553a,a89556a,a89559a,a89560a,a89563a,a89566a,a89567a,a89568a,a89571a,a89574a,a89575a,a89578a,a89581a,a89582a,a89583a,a89586a,a89589a,a89590a,a89593a,a89596a,a89597a,a89598a,a89601a,a89604a,a89605a,a89608a,a89611a,a89612a,a89613a,a89616a,a89619a,a89620a,a89623a,a89626a,a89627a,a89628a,a89631a,a89634a,a89635a,a89638a,a89641a,a89642a,a89643a,a89646a,a89649a,a89650a,a89653a,a89656a,a89657a,a89658a,a89661a,a89664a,a89665a,a89668a,a89671a,a89672a,a89673a,a89676a,a89679a,a89680a,a89683a,a89686a,a89687a,a89688a,a89691a,a89694a,a89695a,a89698a,a89701a,a89702a,a89703a,a89706a,a89709a,a89710a,a89713a,a89716a,a89717a,a89718a,a89721a,a89724a,a89725a,a89728a,a89731a,a89732a,a89733a,a89736a,a89739a,a89740a,a89743a,a89746a,a89747a,a89748a,a89751a,a89754a,a89755a,a89758a,a89761a,a89762a,a89763a,a89766a,a89769a,a89770a,a89773a,a89776a,a89777a,a89778a,a89781a,a89784a,a89785a,a89788a,a89791a,a89792a,a89793a,a89796a,a89799a,a89800a,a89803a,a89806a,a89807a,a89808a,a89811a,a89814a,a89815a,a89818a,a89821a,a89822a,a89823a,a89826a,a89829a,a89830a,a89833a,a89836a,a89837a,a89838a,a89841a,a89844a,a89845a,a89848a,a89851a,a89852a,a89853a,a89856a,a89859a,a89860a,a89863a,a89866a,a89867a,a89868a,a89871a,a89874a,a89875a,a89878a,a89881a,a89882a,a89883a,a89886a,a89889a,a89890a,a89893a,a89896a,a89897a,a89898a,a89901a,a89904a,a89905a,a89908a,a89911a,a89912a,a89913a,a89916a,a89919a,a89920a,a89923a,a89926a,a89927a,a89928a,a89931a,a89934a,a89935a,a89938a,a89941a,a89942a,a89943a,a89946a,a89949a,a89950a,a89953a,a89956a,a89957a,a89958a,a89961a,a89964a,a89965a,a89968a,a89971a,a89972a,a89973a,a89976a,a89979a,a89980a,a89983a,a89986a,a89987a,a89988a,a89991a,a89994a,a89995a,a89998a,a90001a,a90002a,a90003a,a90006a,a90009a,a90010a,a90013a,a90016a,a90017a,a90018a,a90021a,a90024a,a90025a,a90028a,a90031a,a90032a,a90033a,a90036a,a90039a,a90040a,a90043a,a90046a,a90047a,a90048a,a90051a,a90054a,a90055a,a90058a,a90061a,a90062a,a90063a,a90066a,a90069a,a90070a,a90073a,a90076a,a90077a,a90078a,a90081a,a90084a,a90085a,a90088a,a90091a,a90092a,a90093a,a90096a,a90099a,a90100a,a90103a,a90106a,a90107a,a90108a,a90111a,a90114a,a90115a,a90118a,a90121a,a90122a,a90123a,a90126a,a90129a,a90130a,a90133a,a90136a,a90137a,a90138a,a90141a,a90144a,a90145a,a90148a,a90151a,a90152a,a90153a,a90156a,a90159a,a90160a,a90163a,a90166a,a90167a,a90168a,a90171a,a90174a,a90175a,a90178a,a90181a,a90182a,a90183a,a90186a,a90189a,a90190a,a90193a,a90196a,a90197a,a90198a,a90201a,a90204a,a90205a,a90208a,a90211a,a90212a,a90213a,a90216a,a90219a,a90220a,a90223a,a90226a,a90227a,a90228a,a90231a,a90234a,a90235a,a90238a,a90241a,a90242a,a90243a,a90246a,a90249a,a90250a,a90253a,a90256a,a90257a,a90258a,a90261a,a90264a,a90265a,a90268a,a90271a,a90272a,a90273a,a90276a,a90279a,a90280a,a90283a,a90286a,a90287a,a90288a,a90291a,a90294a,a90295a,a90298a,a90301a,a90302a,a90303a,a90306a,a90309a,a90310a,a90313a,a90316a,a90317a,a90318a,a90321a,a90324a,a90325a,a90328a,a90331a,a90332a,a90333a,a90336a,a90339a,a90340a,a90343a,a90346a,a90347a,a90348a,a90351a,a90354a,a90355a,a90358a,a90361a,a90362a,a90363a,a90366a,a90369a,a90370a,a90373a,a90376a,a90377a,a90378a,a90381a,a90384a,a90385a,a90388a,a90391a,a90392a,a90393a,a90396a,a90399a,a90400a,a90403a,a90406a,a90407a,a90408a,a90411a,a90414a,a90415a,a90418a,a90421a,a90422a,a90423a,a90426a,a90429a,a90430a,a90433a,a90436a,a90437a,a90438a,a90441a,a90444a,a90445a,a90448a,a90451a,a90452a,a90453a,a90456a,a90459a,a90460a,a90463a,a90466a,a90467a,a90468a,a90471a,a90474a,a90475a,a90478a,a90481a,a90482a,a90483a,a90486a,a90489a,a90490a,a90493a,a90496a,a90497a,a90498a,a90501a,a90504a,a90505a,a90508a,a90511a,a90512a,a90513a,a90516a,a90519a,a90520a,a90523a,a90526a,a90527a,a90528a,a90531a,a90534a,a90535a,a90538a,a90541a,a90542a,a90543a,a90546a,a90549a,a90550a,a90553a,a90556a,a90557a,a90558a,a90561a,a90564a,a90565a,a90568a,a90571a,a90572a,a90573a,a90576a,a90579a,a90580a,a90583a,a90586a,a90587a,a90588a,a90591a,a90594a,a90595a,a90598a,a90601a,a90602a,a90603a,a90606a,a90609a,a90610a,a90613a,a90616a,a90617a,a90618a,a90621a,a90624a,a90625a,a90628a,a90631a,a90632a,a90633a,a90636a,a90639a,a90640a,a90643a,a90646a,a90647a,a90648a,a90651a,a90654a,a90655a,a90658a,a90661a,a90662a,a90663a,a90666a,a90669a,a90670a,a90673a,a90676a,a90677a,a90678a,a90681a,a90684a,a90685a,a90688a,a90691a,a90692a,a90693a,a90696a,a90699a,a90700a,a90703a,a90706a,a90707a,a90708a,a90711a,a90714a,a90715a,a90718a,a90721a,a90722a,a90723a,a90726a,a90729a,a90730a,a90733a,a90736a,a90737a,a90738a,a90741a,a90744a,a90745a,a90748a,a90751a,a90752a,a90753a,a90756a,a90759a,a90760a,a90763a,a90766a,a90767a,a90768a,a90771a,a90774a,a90775a,a90778a,a90781a,a90782a,a90783a,a90786a,a90789a,a90790a,a90793a,a90796a,a90797a,a90798a,a90801a,a90804a,a90805a,a90808a,a90811a,a90812a,a90813a,a90816a,a90819a,a90820a,a90823a,a90826a,a90827a,a90828a,a90831a,a90834a,a90835a,a90838a,a90841a,a90842a,a90843a,a90846a,a90849a,a90850a,a90853a,a90856a,a90857a,a90858a,a90861a,a90864a,a90865a,a90868a,a90871a,a90872a,a90873a,a90876a,a90879a,a90880a,a90883a,a90886a,a90887a,a90888a,a90891a,a90894a,a90895a,a90898a,a90901a,a90902a,a90903a,a90906a,a90909a,a90910a,a90913a,a90916a,a90917a,a90918a,a90921a,a90924a,a90925a,a90928a,a90931a,a90932a,a90933a,a90936a,a90939a,a90940a,a90943a,a90946a,a90947a,a90948a,a90951a,a90954a,a90955a,a90958a,a90961a,a90962a,a90963a,a90966a,a90969a,a90970a,a90973a,a90976a,a90977a,a90978a,a90981a,a90984a,a90985a,a90988a,a90991a,a90992a,a90993a,a90996a,a90999a,a91000a,a91003a,a91006a,a91007a,a91008a,a91011a,a91014a,a91015a,a91018a,a91021a,a91022a,a91023a,a91026a,a91029a,a91030a,a91033a,a91036a,a91037a,a91038a,a91041a,a91044a,a91045a,a91048a,a91051a,a91052a,a91053a,a91056a,a91059a,a91060a,a91063a,a91066a,a91067a,a91068a,a91071a,a91074a,a91075a,a91078a,a91081a,a91082a,a91083a,a91086a,a91089a,a91090a,a91093a,a91096a,a91097a,a91098a,a91101a,a91104a,a91105a,a91108a,a91111a,a91112a,a91113a,a91116a,a91119a,a91120a,a91123a,a91126a,a91127a,a91128a,a91131a,a91134a,a91135a,a91138a,a91141a,a91142a,a91143a,a91146a,a91149a,a91150a,a91153a,a91156a,a91157a,a91158a,a91161a,a91164a,a91165a,a91168a,a91171a,a91172a,a91173a,a91176a,a91179a,a91180a,a91183a,a91186a,a91187a,a91188a,a91191a,a91194a,a91195a,a91198a,a91201a,a91202a,a91203a,a91206a,a91209a,a91210a,a91213a,a91216a,a91217a,a91218a,a91221a,a91224a,a91225a,a91228a,a91231a,a91232a,a91233a,a91236a,a91239a,a91240a,a91243a,a91246a,a91247a,a91248a,a91251a,a91254a,a91255a,a91258a,a91261a,a91262a,a91263a,a91266a,a91269a,a91270a,a91273a,a91276a,a91277a,a91278a,a91281a,a91284a,a91285a,a91288a,a91291a,a91292a,a91293a,a91296a,a91299a,a91300a,a91303a,a91306a,a91307a,a91308a,a91311a,a91314a,a91315a,a91318a,a91321a,a91322a,a91323a,a91326a,a91329a,a91330a,a91333a,a91336a,a91337a,a91338a,a91341a,a91344a,a91345a,a91348a,a91351a,a91352a,a91353a,a91356a,a91359a,a91360a,a91363a,a91366a,a91367a,a91368a,a91371a,a91374a,a91375a,a91378a,a91381a,a91382a,a91383a,a91386a,a91389a,a91390a,a91393a,a91396a,a91397a,a91398a,a91401a,a91404a,a91405a,a91408a,a91411a,a91412a,a91413a,a91416a,a91419a,a91420a,a91423a,a91426a,a91427a,a91428a,a91431a,a91434a,a91435a,a91438a,a91441a,a91442a,a91443a,a91446a,a91449a,a91450a,a91453a,a91456a,a91457a,a91458a,a91461a,a91464a,a91465a,a91468a,a91471a,a91472a,a91473a,a91476a,a91479a,a91480a,a91483a,a91486a,a91487a,a91488a,a91491a,a91494a,a91495a,a91498a,a91501a,a91502a,a91503a,a91506a,a91509a,a91510a,a91513a,a91516a,a91517a,a91518a,a91521a,a91524a,a91525a,a91528a,a91531a,a91532a,a91533a,a91536a,a91539a,a91540a,a91543a,a91546a,a91547a,a91548a,a91551a,a91554a,a91555a,a91558a,a91561a,a91562a,a91563a,a91566a,a91569a,a91570a,a91573a,a91576a,a91577a,a91578a,a91581a,a91584a,a91585a,a91588a,a91591a,a91592a,a91593a,a91596a,a91599a,a91600a,a91603a,a91606a,a91607a,a91608a,a91611a,a91614a,a91615a,a91618a,a91621a,a91622a,a91623a,a91626a,a91629a,a91630a,a91633a,a91636a,a91637a,a91638a,a91641a,a91644a,a91645a,a91648a,a91651a,a91652a,a91653a,a91656a,a91659a,a91660a,a91663a,a91666a,a91667a,a91668a,a91671a,a91674a,a91675a,a91678a,a91681a,a91682a,a91683a,a91686a,a91689a,a91690a,a91693a,a91696a,a91697a,a91698a,a91701a,a91704a,a91705a,a91708a,a91711a,a91712a,a91713a,a91716a,a91719a,a91720a,a91723a,a91726a,a91727a,a91728a,a91731a,a91734a,a91735a,a91738a,a91741a,a91742a,a91743a,a91746a,a91749a,a91750a,a91753a,a91756a,a91757a,a91758a,a91761a,a91764a,a91765a,a91768a,a91771a,a91772a,a91773a,a91776a,a91779a,a91780a,a91783a,a91786a,a91787a,a91788a,a91791a,a91794a,a91795a,a91798a,a91801a,a91802a,a91803a,a91806a,a91809a,a91810a,a91813a,a91816a,a91817a,a91818a,a91821a,a91824a,a91825a,a91828a,a91831a,a91832a,a91833a,a91836a,a91839a,a91840a,a91843a,a91846a,a91847a,a91848a,a91851a,a91854a,a91855a,a91858a,a91861a,a91862a,a91863a,a91866a,a91869a,a91870a,a91873a,a91876a,a91877a,a91878a,a91881a,a91884a,a91885a,a91888a,a91891a,a91892a,a91893a,a91896a,a91899a,a91900a,a91903a,a91906a,a91907a,a91908a,a91911a,a91914a,a91915a,a91918a,a91921a,a91922a,a91923a,a91926a,a91929a,a91930a,a91933a,a91936a,a91937a,a91938a,a91941a,a91944a,a91945a,a91948a,a91951a,a91952a,a91953a,a91956a,a91959a,a91960a,a91963a,a91966a,a91967a,a91968a,a91971a,a91974a,a91975a,a91978a,a91981a,a91982a,a91983a,a91986a,a91989a,a91990a,a91993a,a91996a,a91997a,a91998a,a92001a,a92004a,a92005a,a92008a,a92011a,a92012a,a92013a,a92016a,a92019a,a92020a,a92023a,a92026a,a92027a,a92028a,a92031a,a92034a,a92035a,a92038a,a92041a,a92042a,a92043a,a92046a,a92049a,a92050a,a92053a,a92056a,a92057a,a92058a,a92061a,a92064a,a92065a,a92068a,a92071a,a92072a,a92073a,a92076a,a92079a,a92080a,a92083a,a92086a,a92087a,a92088a,a92091a,a92094a,a92095a,a92098a,a92101a,a92102a,a92103a,a92106a,a92109a,a92110a,a92113a,a92116a,a92117a,a92118a,a92121a,a92124a,a92125a,a92128a,a92131a,a92132a,a92133a,a92136a,a92139a,a92140a,a92143a,a92146a,a92147a,a92148a,a92151a,a92154a,a92155a,a92158a,a92161a,a92162a,a92163a,a92166a,a92169a,a92170a,a92173a,a92176a,a92177a,a92178a,a92181a,a92184a,a92185a,a92188a,a92191a,a92192a,a92193a,a92196a,a92199a,a92200a,a92203a,a92206a,a92207a,a92208a,a92211a,a92214a,a92215a,a92218a,a92221a,a92222a,a92223a,a92226a,a92229a,a92230a,a92233a,a92236a,a92237a,a92238a,a92241a,a92244a,a92245a,a92248a,a92251a,a92252a,a92253a,a92256a,a92259a,a92260a,a92263a,a92266a,a92267a,a92268a,a92271a,a92274a,a92275a,a92278a,a92281a,a92282a,a92283a,a92286a,a92289a,a92290a,a92293a,a92296a,a92297a,a92298a,a92301a,a92304a,a92305a,a92308a,a92311a,a92312a,a92313a,a92316a,a92319a,a92320a,a92323a,a92326a,a92327a,a92328a,a92331a,a92334a,a92335a,a92338a,a92341a,a92342a,a92343a,a92346a,a92349a,a92350a,a92353a,a92356a,a92357a,a92358a,a92361a,a92364a,a92365a,a92368a,a92371a,a92372a,a92373a,a92376a,a92379a,a92380a,a92383a,a92386a,a92387a,a92388a,a92391a,a92394a,a92395a,a92398a,a92401a,a92402a,a92403a,a92406a,a92409a,a92410a,a92413a,a92416a,a92417a,a92418a,a92421a,a92424a,a92425a,a92428a,a92431a,a92432a,a92433a,a92436a,a92439a,a92440a,a92443a,a92446a,a92447a,a92448a,a92451a,a92454a,a92455a,a92458a,a92461a,a92462a,a92463a,a92466a,a92469a,a92470a,a92473a,a92476a,a92477a,a92478a,a92481a,a92484a,a92485a,a92488a,a92491a,a92492a,a92493a,a92496a,a92499a,a92500a,a92503a,a92506a,a92507a,a92508a,a92511a,a92514a,a92515a,a92518a,a92521a,a92522a,a92523a,a92526a,a92529a,a92530a,a92533a,a92536a,a92537a,a92538a,a92541a,a92544a,a92545a,a92548a,a92551a,a92552a,a92553a,a92556a,a92559a,a92560a,a92563a,a92566a,a92567a,a92568a,a92571a,a92574a,a92575a,a92578a,a92581a,a92582a,a92583a,a92586a,a92589a,a92590a,a92593a,a92596a,a92597a,a92598a,a92601a,a92604a,a92605a,a92608a,a92611a,a92612a,a92613a,a92616a,a92619a,a92620a,a92623a,a92626a,a92627a,a92628a,a92631a,a92634a,a92635a,a92638a,a92641a,a92642a,a92643a,a92646a,a92649a,a92650a,a92653a,a92656a,a92657a,a92658a,a92661a,a92664a,a92665a,a92668a,a92671a,a92672a,a92673a,a92676a,a92679a,a92680a,a92683a,a92686a,a92687a,a92688a,a92691a,a92694a,a92695a,a92698a,a92701a,a92702a,a92703a,a92706a,a92709a,a92710a,a92713a,a92716a,a92717a,a92718a,a92721a,a92724a,a92725a,a92728a,a92731a,a92732a,a92733a,a92736a,a92739a,a92740a,a92743a,a92746a,a92747a,a92748a,a92751a,a92754a,a92755a,a92758a,a92761a,a92762a,a92763a,a92766a,a92769a,a92770a,a92773a,a92776a,a92777a,a92778a,a92781a,a92784a,a92785a,a92788a,a92791a,a92792a,a92793a,a92796a,a92799a,a92800a,a92803a,a92806a,a92807a,a92808a,a92811a,a92814a,a92815a,a92818a,a92821a,a92822a,a92823a,a92826a,a92829a,a92830a,a92833a,a92836a,a92837a,a92838a,a92841a,a92844a,a92845a,a92848a,a92851a,a92852a,a92853a,a92856a,a92859a,a92860a,a92863a,a92866a,a92867a,a92868a,a92871a,a92874a,a92875a,a92878a,a92881a,a92882a,a92883a,a92886a,a92889a,a92890a,a92893a,a92896a,a92897a,a92898a,a92901a,a92904a,a92905a,a92908a,a92911a,a92912a,a92913a,a92916a,a92919a,a92920a,a92923a,a92926a,a92927a,a92928a,a92931a,a92934a,a92935a,a92938a,a92941a,a92942a,a92943a,a92946a,a92949a,a92950a,a92953a,a92956a,a92957a,a92958a,a92961a,a92964a,a92965a,a92968a,a92971a,a92972a,a92973a,a92976a,a92979a,a92980a,a92983a,a92986a,a92987a,a92988a,a92991a,a92994a,a92995a,a92998a,a93001a,a93002a,a93003a,a93006a,a93009a,a93010a,a93013a,a93016a,a93017a,a93018a,a93021a,a93024a,a93025a,a93028a,a93031a,a93032a,a93033a,a93036a,a93039a,a93040a,a93043a,a93046a,a93047a,a93048a,a93051a,a93054a,a93055a,a93058a,a93061a,a93062a,a93063a,a93066a,a93069a,a93070a,a93073a,a93076a,a93077a,a93078a,a93081a,a93084a,a93085a,a93088a,a93091a,a93092a,a93093a,a93096a,a93099a,a93100a,a93103a,a93106a,a93107a,a93108a,a93111a,a93114a,a93115a,a93118a,a93121a,a93122a,a93123a,a93126a,a93129a,a93130a,a93133a,a93136a,a93137a,a93138a,a93141a,a93144a,a93145a,a93148a,a93151a,a93152a,a93153a,a93156a,a93159a,a93160a,a93163a,a93166a,a93167a,a93168a,a93171a,a93174a,a93175a,a93178a,a93181a,a93182a,a93183a,a93186a,a93189a,a93190a,a93193a,a93196a,a93197a,a93198a,a93201a,a93204a,a93205a,a93208a,a93211a,a93212a,a93213a,a93216a,a93219a,a93220a,a93223a,a93226a,a93227a,a93228a,a93231a,a93234a,a93235a,a93238a,a93241a,a93242a,a93243a,a93246a,a93249a,a93250a,a93253a,a93256a,a93257a,a93258a,a93261a,a93264a,a93265a,a93268a,a93271a,a93272a,a93273a,a93276a,a93279a,a93280a,a93283a,a93286a,a93287a,a93288a,a93291a,a93294a,a93295a,a93298a,a93301a,a93302a,a93303a,a93306a,a93309a,a93310a,a93313a,a93316a,a93317a,a93318a,a93321a,a93324a,a93325a,a93328a,a93331a,a93332a,a93333a,a93336a,a93339a,a93340a,a93343a,a93346a,a93347a,a93348a,a93351a,a93354a,a93355a,a93358a,a93361a,a93362a,a93363a,a93366a,a93369a,a93370a,a93373a,a93376a,a93377a,a93378a,a93381a,a93384a,a93385a,a93388a,a93391a,a93392a,a93393a,a93396a,a93399a,a93400a,a93403a,a93406a,a93407a,a93408a,a93411a,a93414a,a93415a,a93418a,a93421a,a93422a,a93423a,a93426a,a93429a,a93430a,a93433a,a93436a,a93437a,a93438a,a93441a,a93444a,a93445a,a93448a,a93451a,a93452a,a93453a,a93456a,a93459a,a93460a,a93463a,a93466a,a93467a,a93468a,a93471a,a93474a,a93475a,a93478a,a93481a,a93482a,a93483a,a93486a,a93489a,a93490a,a93493a,a93496a,a93497a,a93498a,a93501a,a93504a,a93505a,a93508a,a93511a,a93512a,a93513a,a93516a,a93519a,a93520a,a93523a,a93526a,a93527a,a93528a,a93531a,a93534a,a93535a,a93538a,a93541a,a93542a,a93543a,a93546a,a93549a,a93550a,a93553a,a93556a,a93557a,a93558a,a93561a,a93564a,a93565a,a93568a,a93571a,a93572a,a93573a,a93576a,a93579a,a93580a,a93583a,a93586a,a93587a,a93588a,a93591a,a93594a,a93595a,a93598a,a93601a,a93602a,a93603a,a93606a,a93609a,a93610a,a93613a,a93616a,a93617a,a93618a,a93621a,a93624a,a93625a,a93628a,a93631a,a93632a,a93633a,a93636a,a93639a,a93640a,a93643a,a93646a,a93647a,a93648a,a93651a,a93654a,a93655a,a93658a,a93661a,a93662a,a93663a,a93666a,a93669a,a93670a,a93673a,a93676a,a93677a,a93678a,a93681a,a93684a,a93685a,a93688a,a93691a,a93692a,a93693a,a93696a,a93699a,a93700a,a93703a,a93706a,a93707a,a93708a,a93711a,a93714a,a93715a,a93718a,a93721a,a93722a,a93723a,a93726a,a93729a,a93730a,a93733a,a93736a,a93737a,a93738a,a93741a,a93744a,a93745a,a93748a,a93751a,a93752a,a93753a,a93756a,a93759a,a93760a,a93763a,a93766a,a93767a,a93768a,a93771a,a93774a,a93775a,a93778a,a93781a,a93782a,a93783a,a93786a,a93789a,a93790a,a93793a,a93796a,a93797a,a93798a,a93801a,a93804a,a93805a,a93808a,a93811a,a93812a,a93813a,a93816a,a93819a,a93820a,a93823a,a93826a,a93827a,a93828a,a93831a,a93834a,a93835a,a93838a,a93841a,a93842a,a93843a,a93846a,a93849a,a93850a,a93853a,a93856a,a93857a,a93858a,a93861a,a93864a,a93865a,a93868a,a93871a,a93872a,a93873a,a93876a,a93879a,a93880a,a93883a,a93886a,a93887a,a93888a,a93891a,a93894a,a93895a,a93898a,a93901a,a93902a,a93903a,a93906a,a93909a,a93910a,a93913a,a93916a,a93917a,a93918a,a93921a,a93924a,a93925a,a93928a,a93931a,a93932a,a93933a,a93936a,a93939a,a93940a,a93943a,a93946a,a93947a,a93948a,a93951a,a93954a,a93955a,a93958a,a93961a,a93962a,a93963a,a93966a,a93969a,a93970a,a93973a,a93976a,a93977a,a93978a,a93981a,a93984a,a93985a,a93988a,a93991a,a93992a,a93993a,a93996a,a93999a,a94000a,a94003a,a94006a,a94007a,a94008a,a94011a,a94014a,a94015a,a94018a,a94021a,a94022a,a94023a,a94026a,a94029a,a94030a,a94033a,a94036a,a94037a,a94038a,a94041a,a94044a,a94045a,a94048a,a94051a,a94052a,a94053a,a94056a,a94059a,a94060a,a94063a,a94066a,a94067a,a94068a,a94071a,a94074a,a94075a,a94078a,a94081a,a94082a,a94083a,a94086a,a94089a,a94090a,a94093a,a94096a,a94097a,a94098a,a94101a,a94104a,a94105a,a94108a,a94111a,a94112a,a94113a,a94116a,a94119a,a94120a,a94123a,a94126a,a94127a,a94128a,a94131a,a94134a,a94135a,a94138a,a94141a,a94142a,a94143a,a94146a,a94149a,a94150a,a94153a,a94156a,a94157a,a94158a,a94161a,a94164a,a94165a,a94168a,a94171a,a94172a,a94173a,a94176a,a94179a,a94180a,a94183a,a94186a,a94187a,a94188a,a94191a,a94194a,a94195a,a94198a,a94201a,a94202a,a94203a,a94206a,a94209a,a94210a,a94213a,a94216a,a94217a,a94218a,a94221a,a94224a,a94225a,a94228a,a94231a,a94232a,a94233a,a94236a,a94239a,a94240a,a94243a,a94246a,a94247a,a94248a,a94251a,a94254a,a94255a,a94258a,a94261a,a94262a,a94263a,a94266a,a94269a,a94270a,a94273a,a94276a,a94277a,a94278a,a94281a,a94284a,a94285a,a94288a,a94291a,a94292a,a94293a,a94296a,a94299a,a94300a,a94303a,a94306a,a94307a,a94308a,a94311a,a94314a,a94315a,a94318a,a94321a,a94322a,a94323a,a94326a,a94329a,a94330a,a94333a,a94336a,a94337a,a94338a,a94341a,a94344a,a94345a,a94348a,a94351a,a94352a,a94353a,a94356a,a94359a,a94360a,a94363a,a94366a,a94367a,a94368a,a94371a,a94374a,a94375a,a94378a,a94381a,a94382a,a94383a,a94386a,a94389a,a94390a,a94393a,a94396a,a94397a,a94398a,a94401a,a94404a,a94405a,a94408a,a94411a,a94412a,a94413a,a94416a,a94419a,a94420a,a94423a,a94426a,a94427a,a94428a,a94431a,a94434a,a94435a,a94438a,a94441a,a94442a,a94443a,a94446a,a94449a,a94450a,a94453a,a94456a,a94457a,a94458a,a94461a,a94464a,a94465a,a94468a,a94471a,a94472a,a94473a,a94476a,a94479a,a94480a,a94483a,a94486a,a94487a,a94488a,a94491a,a94494a,a94495a,a94498a,a94501a,a94502a,a94503a,a94506a,a94509a,a94510a,a94513a,a94516a,a94517a,a94518a,a94521a,a94524a,a94525a,a94528a,a94531a,a94532a,a94533a,a94536a,a94539a,a94540a,a94543a,a94546a,a94547a,a94548a,a94551a,a94554a,a94555a,a94558a,a94561a,a94562a,a94563a,a94566a,a94569a,a94570a,a94573a,a94576a,a94577a,a94578a,a94581a,a94584a,a94585a,a94588a,a94591a,a94592a,a94593a,a94596a,a94599a,a94600a,a94603a,a94606a,a94607a,a94608a,a94611a,a94614a,a94615a,a94618a,a94621a,a94622a,a94623a,a94626a,a94629a,a94630a,a94633a,a94636a,a94637a,a94638a,a94641a,a94644a,a94645a,a94648a,a94651a,a94652a,a94653a,a94656a,a94659a,a94660a,a94663a,a94666a,a94667a,a94668a,a94671a,a94674a,a94675a,a94678a,a94681a,a94682a,a94683a,a94686a,a94689a,a94690a,a94693a,a94696a,a94697a,a94698a,a94701a,a94704a,a94705a,a94708a,a94711a,a94712a,a94713a,a94716a,a94719a,a94720a,a94723a,a94726a,a94727a,a94728a,a94731a,a94734a,a94735a,a94738a,a94741a,a94742a,a94743a,a94746a,a94749a,a94750a,a94753a,a94756a,a94757a,a94758a,a94761a,a94764a,a94765a,a94768a,a94771a,a94772a,a94773a,a94776a,a94779a,a94780a,a94783a,a94786a,a94787a,a94788a,a94791a,a94794a,a94795a,a94798a,a94801a,a94802a,a94803a,a94806a,a94809a,a94810a,a94813a,a94816a,a94817a,a94818a,a94821a,a94824a,a94825a,a94828a,a94831a,a94832a,a94833a,a94836a,a94839a,a94840a,a94843a,a94846a,a94847a,a94848a,a94851a,a94854a,a94855a,a94858a,a94861a,a94862a,a94863a,a94866a,a94869a,a94870a,a94873a,a94876a,a94877a,a94878a,a94881a,a94884a,a94885a,a94888a,a94891a,a94892a,a94893a,a94896a,a94899a,a94900a,a94903a,a94906a,a94907a,a94908a,a94911a,a94914a,a94915a,a94918a,a94921a,a94922a,a94923a,a94926a,a94929a,a94930a,a94933a,a94936a,a94937a,a94938a,a94941a,a94944a,a94945a,a94948a,a94951a,a94952a,a94953a,a94956a,a94959a,a94960a,a94963a,a94966a,a94967a,a94968a,a94971a,a94974a,a94975a,a94978a,a94981a,a94982a,a94983a,a94986a,a94989a,a94990a,a94993a,a94996a,a94997a,a94998a,a95001a,a95004a,a95005a,a95008a,a95011a,a95012a,a95013a,a95016a,a95019a,a95020a,a95023a,a95026a,a95027a,a95028a,a95031a,a95034a,a95035a,a95038a,a95041a,a95042a,a95043a,a95046a,a95049a,a95050a,a95053a,a95056a,a95057a,a95058a,a95061a,a95064a,a95065a,a95068a,a95071a,a95072a,a95073a,a95076a,a95079a,a95080a,a95083a,a95086a,a95087a,a95088a,a95091a,a95094a,a95095a,a95098a,a95101a,a95102a,a95103a,a95106a,a95109a,a95110a,a95113a,a95116a,a95117a,a95118a,a95121a,a95124a,a95125a,a95128a,a95131a,a95132a,a95133a,a95136a,a95139a,a95140a,a95143a,a95146a,a95147a,a95148a,a95151a,a95154a,a95155a,a95158a,a95161a,a95162a,a95163a,a95166a,a95169a,a95170a,a95173a,a95176a,a95177a,a95178a,a95181a,a95184a,a95185a,a95188a,a95191a,a95192a,a95193a,a95196a,a95199a,a95200a,a95203a,a95206a,a95207a,a95208a,a95211a,a95214a,a95215a,a95218a,a95221a,a95222a,a95223a,a95226a,a95229a,a95230a,a95233a,a95236a,a95237a,a95238a,a95241a,a95244a,a95245a,a95248a,a95251a,a95252a,a95253a,a95256a,a95259a,a95260a,a95263a,a95266a,a95267a,a95268a,a95271a,a95274a,a95275a,a95278a,a95281a,a95282a,a95283a,a95286a,a95289a,a95290a,a95293a,a95296a,a95297a,a95298a,a95301a,a95304a,a95305a,a95308a,a95311a,a95312a,a95313a,a95316a,a95319a,a95320a,a95323a,a95326a,a95327a,a95328a,a95331a,a95334a,a95335a,a95338a,a95341a,a95342a,a95343a,a95346a,a95349a,a95350a,a95353a,a95356a,a95357a,a95358a,a95361a,a95364a,a95365a,a95368a,a95371a,a95372a,a95373a,a95376a,a95379a,a95380a,a95383a,a95386a,a95387a,a95388a,a95391a,a95394a,a95395a,a95398a,a95401a,a95402a,a95403a,a95406a,a95409a,a95410a,a95413a,a95416a,a95417a,a95418a,a95421a,a95424a,a95425a,a95428a,a95431a,a95432a,a95433a,a95436a,a95439a,a95440a,a95443a,a95446a,a95447a,a95448a,a95451a,a95454a,a95455a,a95458a,a95461a,a95462a,a95463a,a95466a,a95469a,a95470a,a95473a,a95476a,a95477a,a95478a,a95481a,a95484a,a95485a,a95488a,a95491a,a95492a,a95493a,a95496a,a95499a,a95500a,a95503a,a95506a,a95507a,a95508a,a95511a,a95514a,a95515a,a95518a,a95521a,a95522a,a95523a,a95526a,a95529a,a95530a,a95533a,a95536a,a95537a,a95538a,a95541a,a95544a,a95545a,a95548a,a95551a,a95552a,a95553a,a95556a,a95559a,a95560a,a95563a,a95566a,a95567a,a95568a,a95571a,a95574a,a95575a,a95578a,a95581a,a95582a,a95583a,a95586a,a95589a,a95590a,a95593a,a95596a,a95597a,a95598a,a95601a,a95604a,a95605a,a95608a,a95611a,a95612a,a95613a,a95616a,a95619a,a95620a,a95623a,a95626a,a95627a,a95628a,a95631a,a95634a,a95635a,a95638a,a95641a,a95642a,a95643a,a95646a,a95649a,a95650a,a95653a,a95656a,a95657a,a95658a,a95661a,a95664a,a95665a,a95668a,a95671a,a95672a,a95673a,a95676a,a95679a,a95680a,a95683a,a95686a,a95687a,a95688a,a95691a,a95694a,a95695a,a95698a,a95701a,a95702a,a95703a,a95706a,a95709a,a95710a,a95713a,a95716a,a95717a,a95718a,a95721a,a95724a,a95725a,a95728a,a95731a,a95732a,a95733a,a95736a,a95739a,a95740a,a95743a,a95746a,a95747a,a95748a,a95751a,a95754a,a95755a,a95758a,a95761a,a95762a,a95763a,a95766a,a95769a,a95770a,a95773a,a95776a,a95777a,a95778a,a95781a,a95784a,a95785a,a95788a,a95791a,a95792a,a95793a,a95796a,a95799a,a95800a,a95803a,a95806a,a95807a,a95808a,a95811a,a95814a,a95815a,a95818a,a95821a,a95822a,a95823a,a95826a,a95829a,a95830a,a95833a,a95836a,a95837a,a95838a,a95841a,a95844a,a95845a,a95848a,a95851a,a95852a,a95853a,a95856a,a95859a,a95860a,a95863a,a95866a,a95867a,a95868a,a95871a,a95874a,a95875a,a95878a,a95881a,a95882a,a95883a,a95886a,a95889a,a95890a,a95893a,a95896a,a95897a,a95898a,a95901a,a95904a,a95905a,a95908a,a95911a,a95912a,a95913a,a95916a,a95919a,a95920a,a95923a,a95926a,a95927a,a95928a,a95931a,a95934a,a95935a,a95938a,a95941a,a95942a,a95943a,a95946a,a95949a,a95950a,a95953a,a95956a,a95957a,a95958a,a95961a,a95964a,a95965a,a95968a,a95971a,a95972a,a95973a,a95976a,a95979a,a95980a,a95983a,a95986a,a95987a,a95988a,a95991a,a95994a,a95995a,a95998a,a96001a,a96002a,a96003a,a96006a,a96009a,a96010a,a96013a,a96016a,a96017a,a96018a,a96021a,a96024a,a96025a,a96028a,a96031a,a96032a,a96033a,a96036a,a96039a,a96040a,a96043a,a96046a,a96047a,a96048a,a96051a,a96054a,a96055a,a96058a,a96061a,a96062a,a96063a,a96066a,a96069a,a96070a,a96073a,a96076a,a96077a,a96078a,a96081a,a96084a,a96085a,a96088a,a96091a,a96092a,a96093a,a96096a,a96099a,a96100a,a96103a,a96106a,a96107a,a96108a,a96111a,a96114a,a96115a,a96118a,a96121a,a96122a,a96123a,a96126a,a96129a,a96130a,a96133a,a96136a,a96137a,a96138a,a96141a,a96144a,a96145a,a96148a,a96151a,a96152a,a96153a,a96156a,a96159a,a96160a,a96163a,a96166a,a96167a,a96168a,a96171a,a96174a,a96175a,a96178a,a96181a,a96182a,a96183a,a96186a,a96189a,a96190a,a96193a,a96196a,a96197a,a96198a,a96201a,a96204a,a96205a,a96208a,a96211a,a96212a,a96213a,a96216a,a96219a,a96220a,a96223a,a96226a,a96227a,a96228a,a96231a,a96234a,a96235a,a96238a,a96241a,a96242a,a96243a,a96246a,a96249a,a96250a,a96253a,a96256a,a96257a,a96258a,a96261a,a96264a,a96265a,a96268a,a96271a,a96272a,a96273a,a96276a,a96279a,a96280a,a96283a,a96286a,a96287a,a96288a,a96291a,a96294a,a96295a,a96298a,a96301a,a96302a,a96303a,a96306a,a96309a,a96310a,a96313a,a96316a,a96317a,a96318a,a96321a,a96324a,a96325a,a96328a,a96331a,a96332a,a96333a,a96336a,a96339a,a96340a,a96343a,a96346a,a96347a,a96348a,a96351a,a96354a,a96355a,a96358a,a96361a,a96362a,a96363a,a96366a,a96369a,a96370a,a96373a,a96376a,a96377a,a96378a,a96381a,a96384a,a96385a,a96388a,a96391a,a96392a,a96393a,a96396a,a96399a,a96400a,a96403a,a96406a,a96407a,a96408a,a96411a,a96414a,a96415a,a96418a,a96421a,a96422a,a96423a,a96426a,a96429a,a96430a,a96433a,a96436a,a96437a,a96438a,a96441a,a96444a,a96445a,a96448a,a96451a,a96452a,a96453a,a96456a,a96459a,a96460a,a96463a,a96466a,a96467a,a96468a,a96471a,a96474a,a96475a,a96478a,a96481a,a96482a,a96483a,a96486a,a96489a,a96490a,a96493a,a96496a,a96497a,a96498a,a96501a,a96504a,a96505a,a96508a,a96511a,a96512a,a96513a,a96516a,a96519a,a96520a,a96523a,a96526a,a96527a,a96528a,a96531a,a96534a,a96535a,a96538a,a96541a,a96542a,a96543a,a96546a,a96549a,a96550a,a96553a,a96556a,a96557a,a96558a,a96561a,a96564a,a96565a,a96568a,a96571a,a96572a,a96573a,a96576a,a96579a,a96580a,a96583a,a96586a,a96587a,a96588a,a96591a,a96594a,a96595a,a96598a,a96601a,a96602a,a96603a,a96606a,a96609a,a96610a,a96613a,a96616a,a96617a,a96618a,a96621a,a96624a,a96625a,a96628a,a96631a,a96632a,a96633a,a96636a,a96639a,a96640a,a96643a,a96646a,a96647a,a96648a,a96651a,a96654a,a96655a,a96658a,a96661a,a96662a,a96663a,a96666a,a96669a,a96670a,a96673a,a96676a,a96677a,a96678a,a96681a,a96684a,a96685a,a96688a,a96691a,a96692a,a96693a,a96696a,a96699a,a96700a,a96703a,a96706a,a96707a,a96708a,a96711a,a96714a,a96715a,a96718a,a96721a,a96722a,a96723a,a96726a,a96729a,a96730a,a96733a,a96736a,a96737a,a96738a,a96741a,a96744a,a96745a,a96748a,a96751a,a96752a,a96753a,a96756a,a96759a,a96760a,a96763a,a96766a,a96767a,a96768a,a96771a,a96774a,a96775a,a96778a,a96781a,a96782a,a96783a,a96786a,a96789a,a96790a,a96793a,a96796a,a96797a,a96798a,a96801a,a96804a,a96805a,a96808a,a96811a,a96812a,a96813a,a96816a,a96819a,a96820a,a96823a,a96826a,a96827a,a96828a,a96831a,a96834a,a96835a,a96838a,a96841a,a96842a,a96843a,a96846a,a96849a,a96850a,a96853a,a96856a,a96857a,a96858a,a96861a,a96864a,a96865a,a96868a,a96871a,a96872a,a96873a,a96876a,a96879a,a96880a,a96883a,a96886a,a96887a,a96888a,a96891a,a96894a,a96895a,a96898a,a96901a,a96902a,a96903a,a96906a,a96909a,a96910a,a96913a,a96916a,a96917a,a96918a,a96921a,a96924a,a96925a,a96928a,a96931a,a96932a,a96933a,a96936a,a96939a,a96940a,a96943a,a96946a,a96947a,a96948a,a96951a,a96954a,a96955a,a96958a,a96961a,a96962a,a96963a,a96966a,a96969a,a96970a,a96973a,a96976a,a96977a,a96978a,a96981a,a96984a,a96985a,a96988a,a96991a,a96992a,a96993a,a96996a,a96999a,a97000a,a97003a,a97006a,a97007a,a97008a,a97011a,a97014a,a97015a,a97018a,a97021a,a97022a,a97023a,a97026a,a97029a,a97030a,a97033a,a97036a,a97037a,a97038a,a97041a,a97044a,a97045a,a97048a,a97051a,a97052a,a97053a,a97056a,a97059a,a97060a,a97063a,a97066a,a97067a,a97068a,a97071a,a97074a,a97075a,a97078a,a97081a,a97082a,a97083a,a97086a,a97089a,a97090a,a97093a,a97096a,a97097a,a97098a,a97101a,a97104a,a97105a,a97108a,a97111a,a97112a,a97113a,a97116a,a97119a,a97120a,a97123a,a97126a,a97127a,a97128a,a97131a,a97134a,a97135a,a97138a,a97141a,a97142a,a97143a,a97146a,a97149a,a97150a,a97153a,a97156a,a97157a,a97158a,a97161a,a97164a,a97165a,a97168a,a97171a,a97172a,a97173a,a97176a,a97179a,a97180a,a97183a,a97186a,a97187a,a97188a,a97191a,a97194a,a97195a,a97198a,a97201a,a97202a,a97203a,a97206a,a97209a,a97210a,a97213a,a97216a,a97217a,a97218a,a97221a,a97224a,a97225a,a97228a,a97231a,a97232a,a97233a,a97236a,a97239a,a97240a,a97243a,a97246a,a97247a,a97248a,a97251a,a97254a,a97255a,a97258a,a97261a,a97262a,a97263a,a97266a,a97269a,a97270a,a97273a,a97276a,a97277a,a97278a,a97281a,a97284a,a97285a,a97288a,a97291a,a97292a,a97293a,a97296a,a97299a,a97300a,a97303a,a97306a,a97307a,a97308a,a97311a,a97314a,a97315a,a97318a,a97321a,a97322a,a97323a,a97326a,a97329a,a97330a,a97333a,a97336a,a97337a,a97338a,a97341a,a97344a,a97345a,a97348a,a97351a,a97352a,a97353a,a97356a,a97359a,a97360a,a97363a,a97366a,a97367a,a97368a,a97371a,a97374a,a97375a,a97378a,a97381a,a97382a,a97383a,a97386a,a97389a,a97390a,a97393a,a97396a,a97397a,a97398a,a97401a,a97404a,a97405a,a97408a,a97411a,a97412a,a97413a,a97416a,a97419a,a97420a,a97423a,a97426a,a97427a,a97428a,a97431a,a97434a,a97435a,a97438a,a97441a,a97442a,a97443a,a97446a,a97449a,a97450a,a97453a,a97456a,a97457a,a97458a,a97461a,a97464a,a97465a,a97468a,a97471a,a97472a,a97473a,a97476a,a97479a,a97480a,a97483a,a97486a,a97487a,a97488a,a97491a,a97494a,a97495a,a97498a,a97501a,a97502a,a97503a,a97506a,a97509a,a97510a,a97513a,a97516a,a97517a,a97518a,a97521a,a97524a,a97525a,a97528a,a97531a,a97532a,a97533a,a97536a,a97539a,a97540a,a97543a,a97546a,a97547a,a97548a,a97551a,a97554a,a97555a,a97558a,a97561a,a97562a,a97563a,a97566a,a97569a,a97570a,a97573a,a97576a,a97577a,a97578a,a97581a,a97584a,a97585a,a97588a,a97591a,a97592a,a97593a,a97596a,a97599a,a97600a,a97603a,a97606a,a97607a,a97608a,a97611a,a97614a,a97615a,a97618a,a97621a,a97622a,a97623a,a97626a,a97629a,a97630a,a97633a,a97636a,a97637a,a97638a,a97641a,a97644a,a97645a,a97648a,a97651a,a97652a,a97653a,a97656a,a97659a,a97660a,a97663a,a97666a,a97667a,a97668a,a97671a,a97674a,a97675a,a97678a,a97681a,a97682a,a97683a,a97686a,a97689a,a97690a,a97693a,a97696a,a97697a,a97698a,a97701a,a97704a,a97705a,a97708a,a97711a,a97712a,a97713a,a97716a,a97719a,a97720a,a97723a,a97726a,a97727a,a97728a,a97731a,a97734a,a97735a,a97738a,a97741a,a97742a,a97743a,a97746a,a97749a,a97750a,a97753a,a97756a,a97757a,a97758a,a97761a,a97764a,a97765a,a97768a,a97771a,a97772a,a97773a,a97776a,a97779a,a97780a,a97783a,a97786a,a97787a,a97788a,a97791a,a97794a,a97795a,a97798a,a97801a,a97802a,a97803a,a97806a,a97809a,a97810a,a97813a,a97816a,a97817a,a97818a,a97821a,a97824a,a97825a,a97828a,a97831a,a97832a,a97833a,a97836a,a97839a,a97840a,a97843a,a97846a,a97847a,a97848a,a97851a,a97854a,a97855a,a97858a,a97861a,a97862a,a97863a,a97866a,a97869a,a97870a,a97873a,a97876a,a97877a,a97878a,a97881a,a97884a,a97885a,a97888a,a97891a,a97892a,a97893a,a97896a,a97899a,a97900a,a97903a,a97906a,a97907a,a97908a,a97911a,a97914a,a97915a,a97918a,a97921a,a97922a,a97923a,a97926a,a97929a,a97930a,a97933a,a97936a,a97937a,a97938a,a97941a,a97944a,a97945a,a97948a,a97951a,a97952a,a97953a,a97956a,a97959a,a97960a,a97963a,a97966a,a97967a,a97968a,a97971a,a97974a,a97975a,a97978a,a97981a,a97982a,a97983a,a97986a,a97989a,a97990a,a97993a,a97996a,a97997a,a97998a,a98001a,a98004a,a98005a,a98008a,a98011a,a98012a,a98013a,a98016a,a98019a,a98020a,a98023a,a98026a,a98027a,a98028a,a98031a,a98034a,a98035a,a98038a,a98041a,a98042a,a98043a,a98046a,a98049a,a98050a,a98053a,a98056a,a98057a,a98058a,a98061a,a98064a,a98065a,a98068a,a98071a,a98072a,a98073a,a98076a,a98079a,a98080a,a98083a,a98086a,a98087a,a98088a,a98091a,a98094a,a98095a,a98098a,a98101a,a98102a,a98103a,a98106a,a98109a,a98110a,a98113a,a98116a,a98117a,a98118a,a98121a,a98124a,a98125a,a98128a,a98131a,a98132a,a98133a,a98136a,a98139a,a98140a,a98143a,a98146a,a98147a,a98148a,a98151a,a98154a,a98155a,a98158a,a98161a,a98162a,a98163a,a98166a,a98169a,a98170a,a98173a,a98176a,a98177a,a98178a,a98181a,a98184a,a98185a,a98188a,a98191a,a98192a,a98193a,a98196a,a98199a,a98200a,a98203a,a98206a,a98207a,a98208a,a98211a,a98214a,a98215a,a98218a,a98221a,a98222a,a98223a,a98226a,a98229a,a98230a,a98233a,a98236a,a98237a,a98238a,a98241a,a98244a,a98245a,a98248a,a98251a,a98252a,a98253a,a98256a,a98259a,a98260a,a98263a,a98266a,a98267a,a98268a,a98271a,a98274a,a98275a,a98278a,a98281a,a98282a,a98283a,a98286a,a98289a,a98290a,a98293a,a98296a,a98297a,a98298a,a98301a,a98304a,a98305a,a98308a,a98311a,a98312a,a98313a,a98316a,a98319a,a98320a,a98323a,a98326a,a98327a,a98328a,a98331a,a98334a,a98335a,a98338a,a98341a,a98342a,a98343a,a98346a,a98349a,a98350a,a98353a,a98356a,a98357a,a98358a,a98361a,a98364a,a98365a,a98368a,a98371a,a98372a,a98373a,a98376a,a98379a,a98380a,a98383a,a98386a,a98387a,a98388a,a98391a,a98394a,a98395a,a98398a,a98401a,a98402a,a98403a,a98406a,a98409a,a98410a,a98413a,a98417a,a98418a,a98419a,a98420a,a98423a,a98426a,a98427a,a98430a,a98433a,a98434a,a98435a,a98438a,a98441a,a98442a,a98445a,a98449a,a98450a,a98451a,a98452a,a98455a,a98458a,a98459a,a98462a,a98465a,a98466a,a98467a,a98470a,a98473a,a98474a,a98477a,a98481a,a98482a,a98483a,a98484a,a98487a,a98490a,a98491a,a98494a,a98497a,a98498a,a98499a,a98502a,a98505a,a98506a,a98509a,a98513a,a98514a,a98515a,a98516a,a98519a,a98522a,a98523a,a98526a,a98529a,a98530a,a98531a,a98534a,a98537a,a98538a,a98541a,a98545a,a98546a,a98547a,a98548a,a98551a,a98554a,a98555a,a98558a,a98561a,a98562a,a98563a,a98566a,a98569a,a98570a,a98573a,a98577a,a98578a,a98579a,a98580a,a98583a,a98586a,a98587a,a98590a,a98593a,a98594a,a98595a,a98598a,a98601a,a98602a,a98605a,a98609a,a98610a,a98611a,a98612a,a98615a,a98618a,a98619a,a98622a,a98625a,a98626a,a98627a,a98630a,a98633a,a98634a,a98637a,a98641a,a98642a,a98643a,a98644a,a98647a,a98650a,a98651a,a98654a,a98657a,a98658a,a98659a,a98662a,a98665a,a98666a,a98669a,a98673a,a98674a,a98675a,a98676a,a98679a,a98682a,a98683a,a98686a,a98689a,a98690a,a98691a,a98694a,a98697a,a98698a,a98701a,a98705a,a98706a,a98707a,a98708a,a98711a,a98714a,a98715a,a98718a,a98721a,a98722a,a98723a,a98726a,a98729a,a98730a,a98733a,a98737a,a98738a,a98739a,a98740a,a98743a,a98746a,a98747a,a98750a,a98753a,a98754a,a98755a,a98758a,a98761a,a98762a,a98765a,a98769a,a98770a,a98771a,a98772a,a98775a,a98778a,a98779a,a98782a,a98785a,a98786a,a98787a,a98790a,a98793a,a98794a,a98797a,a98801a,a98802a,a98803a,a98804a,a98807a,a98810a,a98811a,a98814a,a98817a,a98818a,a98819a,a98822a,a98825a,a98826a,a98829a,a98833a,a98834a,a98835a,a98836a,a98839a,a98842a,a98843a,a98846a,a98849a,a98850a,a98851a,a98854a,a98857a,a98858a,a98861a,a98865a,a98866a,a98867a,a98868a,a98871a,a98874a,a98875a,a98878a,a98881a,a98882a,a98883a,a98886a,a98889a,a98890a,a98893a,a98897a,a98898a,a98899a,a98900a,a98903a,a98906a,a98907a,a98910a,a98913a,a98914a,a98915a,a98918a,a98921a,a98922a,a98925a,a98929a,a98930a,a98931a,a98932a,a98935a,a98938a,a98939a,a98942a,a98945a,a98946a,a98947a,a98950a,a98953a,a98954a,a98957a,a98961a,a98962a,a98963a,a98964a,a98967a,a98970a,a98971a,a98974a,a98977a,a98978a,a98979a,a98982a,a98985a,a98986a,a98989a,a98993a,a98994a,a98995a,a98996a,a98999a,a99002a,a99003a,a99006a,a99009a,a99010a,a99011a,a99014a,a99017a,a99018a,a99021a,a99025a,a99026a,a99027a,a99028a,a99031a,a99034a,a99035a,a99038a,a99041a,a99042a,a99043a,a99046a,a99049a,a99050a,a99053a,a99057a,a99058a,a99059a,a99060a,a99063a,a99066a,a99067a,a99070a,a99073a,a99074a,a99075a,a99078a,a99081a,a99082a,a99085a,a99089a,a99090a,a99091a,a99092a,a99095a,a99098a,a99099a,a99102a,a99105a,a99106a,a99107a,a99110a,a99113a,a99114a,a99117a,a99121a,a99122a,a99123a,a99124a,a99127a,a99130a,a99131a,a99134a,a99137a,a99138a,a99139a,a99142a,a99145a,a99146a,a99149a,a99153a,a99154a,a99155a,a99156a,a99159a,a99162a,a99163a,a99166a,a99169a,a99170a,a99171a,a99174a,a99177a,a99178a,a99181a,a99185a,a99186a,a99187a,a99188a,a99191a,a99194a,a99195a,a99198a,a99201a,a99202a,a99203a,a99206a,a99209a,a99210a,a99213a,a99217a,a99218a,a99219a,a99220a,a99223a,a99226a,a99227a,a99230a,a99233a,a99234a,a99235a,a99238a,a99241a,a99242a,a99245a,a99249a,a99250a,a99251a,a99252a,a99255a,a99258a,a99259a,a99262a,a99265a,a99266a,a99267a,a99270a,a99273a,a99274a,a99277a,a99281a,a99282a,a99283a,a99284a,a99287a,a99290a,a99291a,a99294a,a99297a,a99298a,a99299a,a99302a,a99305a,a99306a,a99309a,a99313a,a99314a,a99315a,a99316a,a99319a,a99322a,a99323a,a99326a,a99329a,a99330a,a99331a,a99334a,a99337a,a99338a,a99341a,a99345a,a99346a,a99347a,a99348a,a99351a,a99354a,a99355a,a99358a,a99361a,a99362a,a99363a,a99366a,a99369a,a99370a,a99373a,a99377a,a99378a,a99379a,a99380a,a99383a,a99386a,a99387a,a99390a,a99393a,a99394a,a99395a,a99398a,a99401a,a99402a,a99405a,a99409a,a99410a,a99411a,a99412a,a99415a,a99418a,a99419a,a99422a,a99425a,a99426a,a99427a,a99430a,a99433a,a99434a,a99437a,a99441a,a99442a,a99443a,a99444a,a99447a,a99450a,a99451a,a99454a,a99457a,a99458a,a99459a,a99462a,a99465a,a99466a,a99469a,a99473a,a99474a,a99475a,a99476a,a99479a,a99482a,a99483a,a99486a,a99489a,a99490a,a99491a,a99494a,a99497a,a99498a,a99501a,a99505a,a99506a,a99507a,a99508a,a99511a,a99514a,a99515a,a99518a,a99521a,a99522a,a99523a,a99526a,a99529a,a99530a,a99533a,a99537a,a99538a,a99539a,a99540a,a99543a,a99546a,a99547a,a99550a,a99553a,a99554a,a99555a,a99558a,a99561a,a99562a,a99565a,a99569a,a99570a,a99571a,a99572a,a99575a,a99578a,a99579a,a99582a,a99585a,a99586a,a99587a,a99590a,a99593a,a99594a,a99597a,a99601a,a99602a,a99603a,a99604a,a99607a,a99610a,a99611a,a99614a,a99617a,a99618a,a99619a,a99622a,a99625a,a99626a,a99629a,a99633a,a99634a,a99635a,a99636a,a99639a,a99642a,a99643a,a99646a,a99649a,a99650a,a99651a,a99654a,a99657a,a99658a,a99661a,a99665a,a99666a,a99667a,a99668a,a99671a,a99674a,a99675a,a99678a,a99681a,a99682a,a99683a,a99686a,a99689a,a99690a,a99693a,a99697a,a99698a,a99699a,a99700a,a99703a,a99706a,a99707a,a99710a,a99713a,a99714a,a99715a,a99718a,a99721a,a99722a,a99725a,a99729a,a99730a,a99731a,a99732a,a99735a,a99738a,a99739a,a99742a,a99745a,a99746a,a99747a,a99750a,a99753a,a99754a,a99757a,a99761a,a99762a,a99763a,a99764a,a99767a,a99770a,a99771a,a99774a,a99777a,a99778a,a99779a,a99782a,a99785a,a99786a,a99789a,a99793a,a99794a,a99795a,a99796a,a99799a,a99802a,a99803a,a99806a,a99809a,a99810a,a99811a,a99814a,a99817a,a99818a,a99821a,a99825a,a99826a,a99827a,a99828a,a99831a,a99834a,a99835a,a99838a,a99841a,a99842a,a99843a,a99846a,a99849a,a99850a,a99853a,a99857a,a99858a,a99859a,a99860a,a99863a,a99866a,a99867a,a99870a,a99873a,a99874a,a99875a,a99878a,a99881a,a99882a,a99885a,a99889a,a99890a,a99891a,a99892a,a99895a,a99898a,a99899a,a99902a,a99905a,a99906a,a99907a,a99910a,a99913a,a99914a,a99917a,a99921a,a99922a,a99923a,a99924a,a99927a,a99930a,a99931a,a99934a,a99937a,a99938a,a99939a,a99942a,a99945a,a99946a,a99949a,a99953a,a99954a,a99955a,a99956a,a99959a,a99962a,a99963a,a99966a,a99969a,a99970a,a99971a,a99974a,a99977a,a99978a,a99981a,a99985a,a99986a,a99987a,a99988a,a99991a,a99994a,a99995a,a99998a,a100001a,a100002a,a100003a,a100006a,a100009a,a100010a,a100013a,a100017a,a100018a,a100019a,a100020a,a100023a,a100026a,a100027a,a100030a,a100033a,a100034a,a100035a,a100038a,a100041a,a100042a,a100045a,a100049a,a100050a,a100051a,a100052a,a100055a,a100058a,a100059a,a100062a,a100065a,a100066a,a100067a,a100070a,a100073a,a100074a,a100077a,a100081a,a100082a,a100083a,a100084a,a100087a,a100090a,a100091a,a100094a,a100097a,a100098a,a100099a,a100102a,a100105a,a100106a,a100109a,a100113a,a100114a,a100115a,a100116a,a100119a,a100122a,a100123a,a100126a,a100129a,a100130a,a100131a,a100134a,a100137a,a100138a,a100141a,a100145a,a100146a,a100147a,a100148a,a100151a,a100154a,a100155a,a100158a,a100161a,a100162a,a100163a,a100166a,a100169a,a100170a,a100173a,a100177a,a100178a,a100179a,a100180a,a100183a,a100186a,a100187a,a100190a,a100193a,a100194a,a100195a,a100198a,a100201a,a100202a,a100205a,a100209a,a100210a,a100211a,a100212a,a100215a,a100218a,a100219a,a100222a,a100225a,a100226a,a100227a,a100230a,a100233a,a100234a,a100237a,a100241a,a100242a,a100243a,a100244a,a100247a,a100250a,a100251a,a100254a,a100257a,a100258a,a100259a,a100262a,a100265a,a100266a,a100269a,a100273a,a100274a,a100275a,a100276a,a100279a,a100282a,a100283a,a100286a,a100289a,a100290a,a100291a,a100294a,a100297a,a100298a,a100301a,a100305a,a100306a,a100307a,a100308a,a100311a,a100314a,a100315a,a100318a,a100321a,a100322a,a100323a,a100326a,a100329a,a100330a,a100333a,a100337a,a100338a,a100339a,a100340a,a100343a,a100346a,a100347a,a100350a,a100353a,a100354a,a100355a,a100358a,a100361a,a100362a,a100365a,a100369a,a100370a,a100371a,a100372a,a100375a,a100378a,a100379a,a100382a,a100385a,a100386a,a100387a,a100390a,a100393a,a100394a,a100397a,a100401a,a100402a,a100403a,a100404a,a100407a,a100410a,a100411a,a100414a,a100417a,a100418a,a100419a,a100422a,a100425a,a100426a,a100429a,a100433a,a100434a,a100435a,a100436a,a100439a,a100442a,a100443a,a100446a,a100449a,a100450a,a100451a,a100454a,a100457a,a100458a,a100461a,a100465a,a100466a,a100467a,a100468a,a100471a,a100474a,a100475a,a100478a,a100481a,a100482a,a100483a,a100486a,a100489a,a100490a,a100493a,a100497a,a100498a,a100499a,a100500a,a100503a,a100506a,a100507a,a100510a,a100513a,a100514a,a100515a,a100518a,a100521a,a100522a,a100525a,a100529a,a100530a,a100531a,a100532a,a100535a,a100538a,a100539a,a100542a,a100545a,a100546a,a100547a,a100550a,a100553a,a100554a,a100557a,a100561a,a100562a,a100563a,a100564a,a100567a,a100570a,a100571a,a100574a,a100577a,a100578a,a100579a,a100582a,a100585a,a100586a,a100589a,a100593a,a100594a,a100595a,a100596a,a100599a,a100602a,a100603a,a100606a,a100609a,a100610a,a100611a,a100614a,a100617a,a100618a,a100621a,a100625a,a100626a,a100627a,a100628a,a100631a,a100634a,a100635a,a100638a,a100641a,a100642a,a100643a,a100646a,a100649a,a100650a,a100653a,a100657a,a100658a,a100659a,a100660a,a100663a,a100666a,a100667a,a100670a,a100673a,a100674a,a100675a,a100678a,a100681a,a100682a,a100685a,a100689a,a100690a,a100691a,a100692a,a100695a,a100698a,a100699a,a100702a,a100705a,a100706a,a100707a,a100710a,a100713a,a100714a,a100717a,a100721a,a100722a,a100723a,a100724a,a100727a,a100730a,a100731a,a100734a,a100737a,a100738a,a100739a,a100742a,a100745a,a100746a,a100749a,a100753a,a100754a,a100755a,a100756a,a100759a,a100762a,a100763a,a100766a,a100769a,a100770a,a100771a,a100774a,a100777a,a100778a,a100781a,a100785a,a100786a,a100787a,a100788a,a100791a,a100794a,a100795a,a100798a,a100801a,a100802a,a100803a,a100806a,a100809a,a100810a,a100813a,a100817a,a100818a,a100819a,a100820a,a100823a,a100826a,a100827a,a100830a,a100833a,a100834a,a100835a,a100838a,a100841a,a100842a,a100845a,a100849a,a100850a,a100851a,a100852a,a100855a,a100858a,a100859a,a100862a,a100865a,a100866a,a100867a,a100870a,a100873a,a100874a,a100877a,a100881a,a100882a,a100883a,a100884a,a100887a,a100890a,a100891a,a100894a,a100897a,a100898a,a100899a,a100902a,a100905a,a100906a,a100909a,a100913a,a100914a,a100915a,a100916a,a100919a,a100922a,a100923a,a100926a,a100929a,a100930a,a100931a,a100934a,a100937a,a100938a,a100941a,a100945a,a100946a,a100947a,a100948a,a100951a,a100954a,a100955a,a100958a,a100962a,a100963a,a100964a,a100965a,a100968a,a100971a,a100972a,a100975a,a100979a,a100980a,a100981a,a100982a,a100985a,a100988a,a100989a,a100992a,a100996a,a100997a,a100998a,a100999a,a101002a,a101005a,a101006a,a101009a,a101013a,a101014a,a101015a,a101016a,a101019a,a101022a,a101023a,a101026a,a101030a,a101031a,a101032a,a101033a,a101036a,a101039a,a101040a,a101043a,a101047a,a101048a,a101049a,a101050a,a101053a,a101056a,a101057a,a101060a,a101064a,a101065a,a101066a,a101067a,a101070a,a101073a,a101074a,a101077a,a101081a,a101082a,a101083a,a101084a,a101087a,a101090a,a101091a,a101094a,a101098a,a101099a,a101100a,a101101a,a101104a,a101107a,a101108a,a101111a,a101115a,a101116a,a101117a,a101118a,a101121a,a101124a,a101125a,a101128a,a101132a,a101133a,a101134a,a101135a,a101138a,a101141a,a101142a,a101145a,a101149a,a101150a,a101151a,a101152a,a101155a,a101158a,a101159a,a101162a,a101166a,a101167a,a101168a,a101169a,a101172a,a101175a,a101176a,a101179a,a101183a,a101184a,a101185a,a101186a,a101189a,a101192a,a101193a,a101196a,a101200a,a101201a,a101202a,a101203a,a101206a,a101209a,a101210a,a101213a,a101217a,a101218a,a101219a,a101220a: std_logic;
begin

A139 <=( a11104a ) or ( a7403a );
 a1a <=( a101220a  and  a101203a );
 a2a <=( a101186a  and  a101169a );
 a3a <=( a101152a  and  a101135a );
 a4a <=( a101118a  and  a101101a );
 a5a <=( a101084a  and  a101067a );
 a6a <=( a101050a  and  a101033a );
 a7a <=( a101016a  and  a100999a );
 a8a <=( a100982a  and  a100965a );
 a9a <=( a100948a  and  a100931a );
 a10a <=( a100916a  and  a100899a );
 a11a <=( a100884a  and  a100867a );
 a12a <=( a100852a  and  a100835a );
 a13a <=( a100820a  and  a100803a );
 a14a <=( a100788a  and  a100771a );
 a15a <=( a100756a  and  a100739a );
 a16a <=( a100724a  and  a100707a );
 a17a <=( a100692a  and  a100675a );
 a18a <=( a100660a  and  a100643a );
 a19a <=( a100628a  and  a100611a );
 a20a <=( a100596a  and  a100579a );
 a21a <=( a100564a  and  a100547a );
 a22a <=( a100532a  and  a100515a );
 a23a <=( a100500a  and  a100483a );
 a24a <=( a100468a  and  a100451a );
 a25a <=( a100436a  and  a100419a );
 a26a <=( a100404a  and  a100387a );
 a27a <=( a100372a  and  a100355a );
 a28a <=( a100340a  and  a100323a );
 a29a <=( a100308a  and  a100291a );
 a30a <=( a100276a  and  a100259a );
 a31a <=( a100244a  and  a100227a );
 a32a <=( a100212a  and  a100195a );
 a33a <=( a100180a  and  a100163a );
 a34a <=( a100148a  and  a100131a );
 a35a <=( a100116a  and  a100099a );
 a36a <=( a100084a  and  a100067a );
 a37a <=( a100052a  and  a100035a );
 a38a <=( a100020a  and  a100003a );
 a39a <=( a99988a  and  a99971a );
 a40a <=( a99956a  and  a99939a );
 a41a <=( a99924a  and  a99907a );
 a42a <=( a99892a  and  a99875a );
 a43a <=( a99860a  and  a99843a );
 a44a <=( a99828a  and  a99811a );
 a45a <=( a99796a  and  a99779a );
 a46a <=( a99764a  and  a99747a );
 a47a <=( a99732a  and  a99715a );
 a48a <=( a99700a  and  a99683a );
 a49a <=( a99668a  and  a99651a );
 a50a <=( a99636a  and  a99619a );
 a51a <=( a99604a  and  a99587a );
 a52a <=( a99572a  and  a99555a );
 a53a <=( a99540a  and  a99523a );
 a54a <=( a99508a  and  a99491a );
 a55a <=( a99476a  and  a99459a );
 a56a <=( a99444a  and  a99427a );
 a57a <=( a99412a  and  a99395a );
 a58a <=( a99380a  and  a99363a );
 a59a <=( a99348a  and  a99331a );
 a60a <=( a99316a  and  a99299a );
 a61a <=( a99284a  and  a99267a );
 a62a <=( a99252a  and  a99235a );
 a63a <=( a99220a  and  a99203a );
 a64a <=( a99188a  and  a99171a );
 a65a <=( a99156a  and  a99139a );
 a66a <=( a99124a  and  a99107a );
 a67a <=( a99092a  and  a99075a );
 a68a <=( a99060a  and  a99043a );
 a69a <=( a99028a  and  a99011a );
 a70a <=( a98996a  and  a98979a );
 a71a <=( a98964a  and  a98947a );
 a72a <=( a98932a  and  a98915a );
 a73a <=( a98900a  and  a98883a );
 a74a <=( a98868a  and  a98851a );
 a75a <=( a98836a  and  a98819a );
 a76a <=( a98804a  and  a98787a );
 a77a <=( a98772a  and  a98755a );
 a78a <=( a98740a  and  a98723a );
 a79a <=( a98708a  and  a98691a );
 a80a <=( a98676a  and  a98659a );
 a81a <=( a98644a  and  a98627a );
 a82a <=( a98612a  and  a98595a );
 a83a <=( a98580a  and  a98563a );
 a84a <=( a98548a  and  a98531a );
 a85a <=( a98516a  and  a98499a );
 a86a <=( a98484a  and  a98467a );
 a87a <=( a98452a  and  a98435a );
 a88a <=( a98420a  and  a98403a );
 a89a <=( a98388a  and  a98373a );
 a90a <=( a98358a  and  a98343a );
 a91a <=( a98328a  and  a98313a );
 a92a <=( a98298a  and  a98283a );
 a93a <=( a98268a  and  a98253a );
 a94a <=( a98238a  and  a98223a );
 a95a <=( a98208a  and  a98193a );
 a96a <=( a98178a  and  a98163a );
 a97a <=( a98148a  and  a98133a );
 a98a <=( a98118a  and  a98103a );
 a99a <=( a98088a  and  a98073a );
 a100a <=( a98058a  and  a98043a );
 a101a <=( a98028a  and  a98013a );
 a102a <=( a97998a  and  a97983a );
 a103a <=( a97968a  and  a97953a );
 a104a <=( a97938a  and  a97923a );
 a105a <=( a97908a  and  a97893a );
 a106a <=( a97878a  and  a97863a );
 a107a <=( a97848a  and  a97833a );
 a108a <=( a97818a  and  a97803a );
 a109a <=( a97788a  and  a97773a );
 a110a <=( a97758a  and  a97743a );
 a111a <=( a97728a  and  a97713a );
 a112a <=( a97698a  and  a97683a );
 a113a <=( a97668a  and  a97653a );
 a114a <=( a97638a  and  a97623a );
 a115a <=( a97608a  and  a97593a );
 a116a <=( a97578a  and  a97563a );
 a117a <=( a97548a  and  a97533a );
 a118a <=( a97518a  and  a97503a );
 a119a <=( a97488a  and  a97473a );
 a120a <=( a97458a  and  a97443a );
 a121a <=( a97428a  and  a97413a );
 a122a <=( a97398a  and  a97383a );
 a123a <=( a97368a  and  a97353a );
 a124a <=( a97338a  and  a97323a );
 a125a <=( a97308a  and  a97293a );
 a126a <=( a97278a  and  a97263a );
 a127a <=( a97248a  and  a97233a );
 a128a <=( a97218a  and  a97203a );
 a129a <=( a97188a  and  a97173a );
 a130a <=( a97158a  and  a97143a );
 a131a <=( a97128a  and  a97113a );
 a132a <=( a97098a  and  a97083a );
 a133a <=( a97068a  and  a97053a );
 a134a <=( a97038a  and  a97023a );
 a135a <=( a97008a  and  a96993a );
 a136a <=( a96978a  and  a96963a );
 a137a <=( a96948a  and  a96933a );
 a138a <=( a96918a  and  a96903a );
 a139a <=( a96888a  and  a96873a );
 a140a <=( a96858a  and  a96843a );
 a141a <=( a96828a  and  a96813a );
 a142a <=( a96798a  and  a96783a );
 a143a <=( a96768a  and  a96753a );
 a144a <=( a96738a  and  a96723a );
 a145a <=( a96708a  and  a96693a );
 a146a <=( a96678a  and  a96663a );
 a147a <=( a96648a  and  a96633a );
 a148a <=( a96618a  and  a96603a );
 a149a <=( a96588a  and  a96573a );
 a150a <=( a96558a  and  a96543a );
 a151a <=( a96528a  and  a96513a );
 a152a <=( a96498a  and  a96483a );
 a153a <=( a96468a  and  a96453a );
 a154a <=( a96438a  and  a96423a );
 a155a <=( a96408a  and  a96393a );
 a156a <=( a96378a  and  a96363a );
 a157a <=( a96348a  and  a96333a );
 a158a <=( a96318a  and  a96303a );
 a159a <=( a96288a  and  a96273a );
 a160a <=( a96258a  and  a96243a );
 a161a <=( a96228a  and  a96213a );
 a162a <=( a96198a  and  a96183a );
 a163a <=( a96168a  and  a96153a );
 a164a <=( a96138a  and  a96123a );
 a165a <=( a96108a  and  a96093a );
 a166a <=( a96078a  and  a96063a );
 a167a <=( a96048a  and  a96033a );
 a168a <=( a96018a  and  a96003a );
 a169a <=( a95988a  and  a95973a );
 a170a <=( a95958a  and  a95943a );
 a171a <=( a95928a  and  a95913a );
 a172a <=( a95898a  and  a95883a );
 a173a <=( a95868a  and  a95853a );
 a174a <=( a95838a  and  a95823a );
 a175a <=( a95808a  and  a95793a );
 a176a <=( a95778a  and  a95763a );
 a177a <=( a95748a  and  a95733a );
 a178a <=( a95718a  and  a95703a );
 a179a <=( a95688a  and  a95673a );
 a180a <=( a95658a  and  a95643a );
 a181a <=( a95628a  and  a95613a );
 a182a <=( a95598a  and  a95583a );
 a183a <=( a95568a  and  a95553a );
 a184a <=( a95538a  and  a95523a );
 a185a <=( a95508a  and  a95493a );
 a186a <=( a95478a  and  a95463a );
 a187a <=( a95448a  and  a95433a );
 a188a <=( a95418a  and  a95403a );
 a189a <=( a95388a  and  a95373a );
 a190a <=( a95358a  and  a95343a );
 a191a <=( a95328a  and  a95313a );
 a192a <=( a95298a  and  a95283a );
 a193a <=( a95268a  and  a95253a );
 a194a <=( a95238a  and  a95223a );
 a195a <=( a95208a  and  a95193a );
 a196a <=( a95178a  and  a95163a );
 a197a <=( a95148a  and  a95133a );
 a198a <=( a95118a  and  a95103a );
 a199a <=( a95088a  and  a95073a );
 a200a <=( a95058a  and  a95043a );
 a201a <=( a95028a  and  a95013a );
 a202a <=( a94998a  and  a94983a );
 a203a <=( a94968a  and  a94953a );
 a204a <=( a94938a  and  a94923a );
 a205a <=( a94908a  and  a94893a );
 a206a <=( a94878a  and  a94863a );
 a207a <=( a94848a  and  a94833a );
 a208a <=( a94818a  and  a94803a );
 a209a <=( a94788a  and  a94773a );
 a210a <=( a94758a  and  a94743a );
 a211a <=( a94728a  and  a94713a );
 a212a <=( a94698a  and  a94683a );
 a213a <=( a94668a  and  a94653a );
 a214a <=( a94638a  and  a94623a );
 a215a <=( a94608a  and  a94593a );
 a216a <=( a94578a  and  a94563a );
 a217a <=( a94548a  and  a94533a );
 a218a <=( a94518a  and  a94503a );
 a219a <=( a94488a  and  a94473a );
 a220a <=( a94458a  and  a94443a );
 a221a <=( a94428a  and  a94413a );
 a222a <=( a94398a  and  a94383a );
 a223a <=( a94368a  and  a94353a );
 a224a <=( a94338a  and  a94323a );
 a225a <=( a94308a  and  a94293a );
 a226a <=( a94278a  and  a94263a );
 a227a <=( a94248a  and  a94233a );
 a228a <=( a94218a  and  a94203a );
 a229a <=( a94188a  and  a94173a );
 a230a <=( a94158a  and  a94143a );
 a231a <=( a94128a  and  a94113a );
 a232a <=( a94098a  and  a94083a );
 a233a <=( a94068a  and  a94053a );
 a234a <=( a94038a  and  a94023a );
 a235a <=( a94008a  and  a93993a );
 a236a <=( a93978a  and  a93963a );
 a237a <=( a93948a  and  a93933a );
 a238a <=( a93918a  and  a93903a );
 a239a <=( a93888a  and  a93873a );
 a240a <=( a93858a  and  a93843a );
 a241a <=( a93828a  and  a93813a );
 a242a <=( a93798a  and  a93783a );
 a243a <=( a93768a  and  a93753a );
 a244a <=( a93738a  and  a93723a );
 a245a <=( a93708a  and  a93693a );
 a246a <=( a93678a  and  a93663a );
 a247a <=( a93648a  and  a93633a );
 a248a <=( a93618a  and  a93603a );
 a249a <=( a93588a  and  a93573a );
 a250a <=( a93558a  and  a93543a );
 a251a <=( a93528a  and  a93513a );
 a252a <=( a93498a  and  a93483a );
 a253a <=( a93468a  and  a93453a );
 a254a <=( a93438a  and  a93423a );
 a255a <=( a93408a  and  a93393a );
 a256a <=( a93378a  and  a93363a );
 a257a <=( a93348a  and  a93333a );
 a258a <=( a93318a  and  a93303a );
 a259a <=( a93288a  and  a93273a );
 a260a <=( a93258a  and  a93243a );
 a261a <=( a93228a  and  a93213a );
 a262a <=( a93198a  and  a93183a );
 a263a <=( a93168a  and  a93153a );
 a264a <=( a93138a  and  a93123a );
 a265a <=( a93108a  and  a93093a );
 a266a <=( a93078a  and  a93063a );
 a267a <=( a93048a  and  a93033a );
 a268a <=( a93018a  and  a93003a );
 a269a <=( a92988a  and  a92973a );
 a270a <=( a92958a  and  a92943a );
 a271a <=( a92928a  and  a92913a );
 a272a <=( a92898a  and  a92883a );
 a273a <=( a92868a  and  a92853a );
 a274a <=( a92838a  and  a92823a );
 a275a <=( a92808a  and  a92793a );
 a276a <=( a92778a  and  a92763a );
 a277a <=( a92748a  and  a92733a );
 a278a <=( a92718a  and  a92703a );
 a279a <=( a92688a  and  a92673a );
 a280a <=( a92658a  and  a92643a );
 a281a <=( a92628a  and  a92613a );
 a282a <=( a92598a  and  a92583a );
 a283a <=( a92568a  and  a92553a );
 a284a <=( a92538a  and  a92523a );
 a285a <=( a92508a  and  a92493a );
 a286a <=( a92478a  and  a92463a );
 a287a <=( a92448a  and  a92433a );
 a288a <=( a92418a  and  a92403a );
 a289a <=( a92388a  and  a92373a );
 a290a <=( a92358a  and  a92343a );
 a291a <=( a92328a  and  a92313a );
 a292a <=( a92298a  and  a92283a );
 a293a <=( a92268a  and  a92253a );
 a294a <=( a92238a  and  a92223a );
 a295a <=( a92208a  and  a92193a );
 a296a <=( a92178a  and  a92163a );
 a297a <=( a92148a  and  a92133a );
 a298a <=( a92118a  and  a92103a );
 a299a <=( a92088a  and  a92073a );
 a300a <=( a92058a  and  a92043a );
 a301a <=( a92028a  and  a92013a );
 a302a <=( a91998a  and  a91983a );
 a303a <=( a91968a  and  a91953a );
 a304a <=( a91938a  and  a91923a );
 a305a <=( a91908a  and  a91893a );
 a306a <=( a91878a  and  a91863a );
 a307a <=( a91848a  and  a91833a );
 a308a <=( a91818a  and  a91803a );
 a309a <=( a91788a  and  a91773a );
 a310a <=( a91758a  and  a91743a );
 a311a <=( a91728a  and  a91713a );
 a312a <=( a91698a  and  a91683a );
 a313a <=( a91668a  and  a91653a );
 a314a <=( a91638a  and  a91623a );
 a315a <=( a91608a  and  a91593a );
 a316a <=( a91578a  and  a91563a );
 a317a <=( a91548a  and  a91533a );
 a318a <=( a91518a  and  a91503a );
 a319a <=( a91488a  and  a91473a );
 a320a <=( a91458a  and  a91443a );
 a321a <=( a91428a  and  a91413a );
 a322a <=( a91398a  and  a91383a );
 a323a <=( a91368a  and  a91353a );
 a324a <=( a91338a  and  a91323a );
 a325a <=( a91308a  and  a91293a );
 a326a <=( a91278a  and  a91263a );
 a327a <=( a91248a  and  a91233a );
 a328a <=( a91218a  and  a91203a );
 a329a <=( a91188a  and  a91173a );
 a330a <=( a91158a  and  a91143a );
 a331a <=( a91128a  and  a91113a );
 a332a <=( a91098a  and  a91083a );
 a333a <=( a91068a  and  a91053a );
 a334a <=( a91038a  and  a91023a );
 a335a <=( a91008a  and  a90993a );
 a336a <=( a90978a  and  a90963a );
 a337a <=( a90948a  and  a90933a );
 a338a <=( a90918a  and  a90903a );
 a339a <=( a90888a  and  a90873a );
 a340a <=( a90858a  and  a90843a );
 a341a <=( a90828a  and  a90813a );
 a342a <=( a90798a  and  a90783a );
 a343a <=( a90768a  and  a90753a );
 a344a <=( a90738a  and  a90723a );
 a345a <=( a90708a  and  a90693a );
 a346a <=( a90678a  and  a90663a );
 a347a <=( a90648a  and  a90633a );
 a348a <=( a90618a  and  a90603a );
 a349a <=( a90588a  and  a90573a );
 a350a <=( a90558a  and  a90543a );
 a351a <=( a90528a  and  a90513a );
 a352a <=( a90498a  and  a90483a );
 a353a <=( a90468a  and  a90453a );
 a354a <=( a90438a  and  a90423a );
 a355a <=( a90408a  and  a90393a );
 a356a <=( a90378a  and  a90363a );
 a357a <=( a90348a  and  a90333a );
 a358a <=( a90318a  and  a90303a );
 a359a <=( a90288a  and  a90273a );
 a360a <=( a90258a  and  a90243a );
 a361a <=( a90228a  and  a90213a );
 a362a <=( a90198a  and  a90183a );
 a363a <=( a90168a  and  a90153a );
 a364a <=( a90138a  and  a90123a );
 a365a <=( a90108a  and  a90093a );
 a366a <=( a90078a  and  a90063a );
 a367a <=( a90048a  and  a90033a );
 a368a <=( a90018a  and  a90003a );
 a369a <=( a89988a  and  a89973a );
 a370a <=( a89958a  and  a89943a );
 a371a <=( a89928a  and  a89913a );
 a372a <=( a89898a  and  a89883a );
 a373a <=( a89868a  and  a89853a );
 a374a <=( a89838a  and  a89823a );
 a375a <=( a89808a  and  a89793a );
 a376a <=( a89778a  and  a89763a );
 a377a <=( a89748a  and  a89733a );
 a378a <=( a89718a  and  a89703a );
 a379a <=( a89688a  and  a89673a );
 a380a <=( a89658a  and  a89643a );
 a381a <=( a89628a  and  a89613a );
 a382a <=( a89598a  and  a89583a );
 a383a <=( a89568a  and  a89553a );
 a384a <=( a89538a  and  a89523a );
 a385a <=( a89508a  and  a89493a );
 a386a <=( a89480a  and  a89465a );
 a387a <=( a89452a  and  a89437a );
 a388a <=( a89424a  and  a89409a );
 a389a <=( a89396a  and  a89381a );
 a390a <=( a89368a  and  a89353a );
 a391a <=( a89340a  and  a89325a );
 a392a <=( a89312a  and  a89297a );
 a393a <=( a89284a  and  a89269a );
 a394a <=( a89256a  and  a89241a );
 a395a <=( a89228a  and  a89213a );
 a396a <=( a89200a  and  a89185a );
 a397a <=( a89172a  and  a89157a );
 a398a <=( a89144a  and  a89129a );
 a399a <=( a89116a  and  a89101a );
 a400a <=( a89088a  and  a89073a );
 a401a <=( a89060a  and  a89045a );
 a402a <=( a89032a  and  a89017a );
 a403a <=( a89004a  and  a88989a );
 a404a <=( a88976a  and  a88961a );
 a405a <=( a88948a  and  a88933a );
 a406a <=( a88920a  and  a88905a );
 a407a <=( a88892a  and  a88877a );
 a408a <=( a88864a  and  a88849a );
 a409a <=( a88836a  and  a88821a );
 a410a <=( a88808a  and  a88793a );
 a411a <=( a88780a  and  a88765a );
 a412a <=( a88752a  and  a88737a );
 a413a <=( a88724a  and  a88709a );
 a414a <=( a88696a  and  a88681a );
 a415a <=( a88668a  and  a88653a );
 a416a <=( a88640a  and  a88625a );
 a417a <=( a88612a  and  a88597a );
 a418a <=( a88584a  and  a88569a );
 a419a <=( a88556a  and  a88541a );
 a420a <=( a88528a  and  a88513a );
 a421a <=( a88500a  and  a88485a );
 a422a <=( a88472a  and  a88457a );
 a423a <=( a88444a  and  a88429a );
 a424a <=( a88416a  and  a88401a );
 a425a <=( a88388a  and  a88373a );
 a426a <=( a88360a  and  a88345a );
 a427a <=( a88332a  and  a88317a );
 a428a <=( a88304a  and  a88289a );
 a429a <=( a88276a  and  a88261a );
 a430a <=( a88248a  and  a88233a );
 a431a <=( a88220a  and  a88205a );
 a432a <=( a88192a  and  a88177a );
 a433a <=( a88164a  and  a88149a );
 a434a <=( a88136a  and  a88121a );
 a435a <=( a88108a  and  a88093a );
 a436a <=( a88080a  and  a88065a );
 a437a <=( a88052a  and  a88037a );
 a438a <=( a88024a  and  a88009a );
 a439a <=( a87996a  and  a87981a );
 a440a <=( a87968a  and  a87953a );
 a441a <=( a87940a  and  a87925a );
 a442a <=( a87912a  and  a87897a );
 a443a <=( a87884a  and  a87869a );
 a444a <=( a87856a  and  a87841a );
 a445a <=( a87828a  and  a87813a );
 a446a <=( a87800a  and  a87785a );
 a447a <=( a87772a  and  a87757a );
 a448a <=( a87744a  and  a87729a );
 a449a <=( a87716a  and  a87701a );
 a450a <=( a87688a  and  a87673a );
 a451a <=( a87660a  and  a87645a );
 a452a <=( a87632a  and  a87617a );
 a453a <=( a87604a  and  a87589a );
 a454a <=( a87576a  and  a87561a );
 a455a <=( a87548a  and  a87533a );
 a456a <=( a87520a  and  a87505a );
 a457a <=( a87492a  and  a87477a );
 a458a <=( a87464a  and  a87449a );
 a459a <=( a87436a  and  a87421a );
 a460a <=( a87408a  and  a87393a );
 a461a <=( a87380a  and  a87365a );
 a462a <=( a87352a  and  a87337a );
 a463a <=( a87324a  and  a87309a );
 a464a <=( a87296a  and  a87281a );
 a465a <=( a87268a  and  a87253a );
 a466a <=( a87240a  and  a87225a );
 a467a <=( a87212a  and  a87197a );
 a468a <=( a87184a  and  a87169a );
 a469a <=( a87156a  and  a87141a );
 a470a <=( a87128a  and  a87113a );
 a471a <=( a87100a  and  a87085a );
 a472a <=( a87072a  and  a87057a );
 a473a <=( a87044a  and  a87029a );
 a474a <=( a87016a  and  a87001a );
 a475a <=( a86988a  and  a86973a );
 a476a <=( a86960a  and  a86945a );
 a477a <=( a86932a  and  a86917a );
 a478a <=( a86904a  and  a86889a );
 a479a <=( a86876a  and  a86861a );
 a480a <=( a86848a  and  a86833a );
 a481a <=( a86820a  and  a86805a );
 a482a <=( a86792a  and  a86777a );
 a483a <=( a86764a  and  a86749a );
 a484a <=( a86736a  and  a86721a );
 a485a <=( a86708a  and  a86693a );
 a486a <=( a86680a  and  a86665a );
 a487a <=( a86652a  and  a86637a );
 a488a <=( a86624a  and  a86609a );
 a489a <=( a86596a  and  a86581a );
 a490a <=( a86568a  and  a86553a );
 a491a <=( a86540a  and  a86525a );
 a492a <=( a86512a  and  a86497a );
 a493a <=( a86484a  and  a86469a );
 a494a <=( a86456a  and  a86441a );
 a495a <=( a86428a  and  a86413a );
 a496a <=( a86400a  and  a86385a );
 a497a <=( a86372a  and  a86357a );
 a498a <=( a86344a  and  a86329a );
 a499a <=( a86316a  and  a86301a );
 a500a <=( a86288a  and  a86273a );
 a501a <=( a86260a  and  a86245a );
 a502a <=( a86232a  and  a86217a );
 a503a <=( a86204a  and  a86189a );
 a504a <=( a86176a  and  a86161a );
 a505a <=( a86148a  and  a86133a );
 a506a <=( a86120a  and  a86105a );
 a507a <=( a86092a  and  a86077a );
 a508a <=( a86064a  and  a86049a );
 a509a <=( a86036a  and  a86021a );
 a510a <=( a86008a  and  a85993a );
 a511a <=( a85980a  and  a85965a );
 a512a <=( a85952a  and  a85937a );
 a513a <=( a85924a  and  a85909a );
 a514a <=( a85896a  and  a85881a );
 a515a <=( a85868a  and  a85853a );
 a516a <=( a85840a  and  a85825a );
 a517a <=( a85812a  and  a85797a );
 a518a <=( a85784a  and  a85769a );
 a519a <=( a85756a  and  a85741a );
 a520a <=( a85728a  and  a85713a );
 a521a <=( a85700a  and  a85685a );
 a522a <=( a85672a  and  a85657a );
 a523a <=( a85644a  and  a85629a );
 a524a <=( a85616a  and  a85601a );
 a525a <=( a85588a  and  a85573a );
 a526a <=( a85560a  and  a85545a );
 a527a <=( a85532a  and  a85517a );
 a528a <=( a85504a  and  a85489a );
 a529a <=( a85476a  and  a85461a );
 a530a <=( a85448a  and  a85433a );
 a531a <=( a85420a  and  a85405a );
 a532a <=( a85392a  and  a85377a );
 a533a <=( a85364a  and  a85349a );
 a534a <=( a85336a  and  a85321a );
 a535a <=( a85308a  and  a85293a );
 a536a <=( a85280a  and  a85265a );
 a537a <=( a85252a  and  a85237a );
 a538a <=( a85224a  and  a85209a );
 a539a <=( a85196a  and  a85181a );
 a540a <=( a85168a  and  a85153a );
 a541a <=( a85140a  and  a85125a );
 a542a <=( a85112a  and  a85097a );
 a543a <=( a85084a  and  a85069a );
 a544a <=( a85056a  and  a85041a );
 a545a <=( a85028a  and  a85013a );
 a546a <=( a85000a  and  a84985a );
 a547a <=( a84972a  and  a84957a );
 a548a <=( a84944a  and  a84929a );
 a549a <=( a84916a  and  a84901a );
 a550a <=( a84888a  and  a84873a );
 a551a <=( a84860a  and  a84845a );
 a552a <=( a84832a  and  a84817a );
 a553a <=( a84804a  and  a84789a );
 a554a <=( a84776a  and  a84761a );
 a555a <=( a84748a  and  a84733a );
 a556a <=( a84720a  and  a84705a );
 a557a <=( a84692a  and  a84677a );
 a558a <=( a84664a  and  a84649a );
 a559a <=( a84636a  and  a84621a );
 a560a <=( a84608a  and  a84593a );
 a561a <=( a84580a  and  a84565a );
 a562a <=( a84552a  and  a84537a );
 a563a <=( a84524a  and  a84509a );
 a564a <=( a84496a  and  a84481a );
 a565a <=( a84468a  and  a84453a );
 a566a <=( a84440a  and  a84425a );
 a567a <=( a84412a  and  a84397a );
 a568a <=( a84384a  and  a84369a );
 a569a <=( a84356a  and  a84341a );
 a570a <=( a84328a  and  a84313a );
 a571a <=( a84300a  and  a84285a );
 a572a <=( a84272a  and  a84257a );
 a573a <=( a84244a  and  a84229a );
 a574a <=( a84216a  and  a84201a );
 a575a <=( a84188a  and  a84173a );
 a576a <=( a84160a  and  a84145a );
 a577a <=( a84132a  and  a84117a );
 a578a <=( a84104a  and  a84089a );
 a579a <=( a84076a  and  a84061a );
 a580a <=( a84048a  and  a84033a );
 a581a <=( a84020a  and  a84005a );
 a582a <=( a83992a  and  a83977a );
 a583a <=( a83964a  and  a83949a );
 a584a <=( a83936a  and  a83921a );
 a585a <=( a83908a  and  a83893a );
 a586a <=( a83880a  and  a83865a );
 a587a <=( a83852a  and  a83837a );
 a588a <=( a83824a  and  a83809a );
 a589a <=( a83796a  and  a83781a );
 a590a <=( a83768a  and  a83753a );
 a591a <=( a83740a  and  a83725a );
 a592a <=( a83712a  and  a83697a );
 a593a <=( a83684a  and  a83669a );
 a594a <=( a83656a  and  a83641a );
 a595a <=( a83628a  and  a83613a );
 a596a <=( a83600a  and  a83585a );
 a597a <=( a83572a  and  a83557a );
 a598a <=( a83544a  and  a83529a );
 a599a <=( a83516a  and  a83501a );
 a600a <=( a83488a  and  a83473a );
 a601a <=( a83460a  and  a83445a );
 a602a <=( a83432a  and  a83417a );
 a603a <=( a83404a  and  a83389a );
 a604a <=( a83376a  and  a83361a );
 a605a <=( a83348a  and  a83333a );
 a606a <=( a83320a  and  a83305a );
 a607a <=( a83292a  and  a83277a );
 a608a <=( a83264a  and  a83249a );
 a609a <=( a83236a  and  a83221a );
 a610a <=( a83208a  and  a83193a );
 a611a <=( a83180a  and  a83165a );
 a612a <=( a83152a  and  a83137a );
 a613a <=( a83124a  and  a83109a );
 a614a <=( a83096a  and  a83081a );
 a615a <=( a83068a  and  a83053a );
 a616a <=( a83040a  and  a83025a );
 a617a <=( a83012a  and  a82997a );
 a618a <=( a82984a  and  a82969a );
 a619a <=( a82956a  and  a82941a );
 a620a <=( a82928a  and  a82913a );
 a621a <=( a82900a  and  a82885a );
 a622a <=( a82872a  and  a82857a );
 a623a <=( a82844a  and  a82829a );
 a624a <=( a82816a  and  a82801a );
 a625a <=( a82788a  and  a82773a );
 a626a <=( a82760a  and  a82745a );
 a627a <=( a82732a  and  a82717a );
 a628a <=( a82704a  and  a82689a );
 a629a <=( a82676a  and  a82661a );
 a630a <=( a82648a  and  a82633a );
 a631a <=( a82620a  and  a82605a );
 a632a <=( a82592a  and  a82577a );
 a633a <=( a82564a  and  a82549a );
 a634a <=( a82536a  and  a82521a );
 a635a <=( a82508a  and  a82493a );
 a636a <=( a82480a  and  a82465a );
 a637a <=( a82452a  and  a82437a );
 a638a <=( a82424a  and  a82409a );
 a639a <=( a82396a  and  a82381a );
 a640a <=( a82368a  and  a82353a );
 a641a <=( a82340a  and  a82325a );
 a642a <=( a82312a  and  a82297a );
 a643a <=( a82284a  and  a82269a );
 a644a <=( a82256a  and  a82241a );
 a645a <=( a82228a  and  a82213a );
 a646a <=( a82200a  and  a82185a );
 a647a <=( a82172a  and  a82157a );
 a648a <=( a82144a  and  a82129a );
 a649a <=( a82116a  and  a82101a );
 a650a <=( a82088a  and  a82073a );
 a651a <=( a82060a  and  a82045a );
 a652a <=( a82032a  and  a82017a );
 a653a <=( a82004a  and  a81989a );
 a654a <=( a81976a  and  a81961a );
 a655a <=( a81948a  and  a81933a );
 a656a <=( a81920a  and  a81905a );
 a657a <=( a81892a  and  a81877a );
 a658a <=( a81864a  and  a81849a );
 a659a <=( a81836a  and  a81821a );
 a660a <=( a81808a  and  a81793a );
 a661a <=( a81780a  and  a81765a );
 a662a <=( a81752a  and  a81737a );
 a663a <=( a81724a  and  a81709a );
 a664a <=( a81696a  and  a81681a );
 a665a <=( a81668a  and  a81653a );
 a666a <=( a81640a  and  a81625a );
 a667a <=( a81612a  and  a81597a );
 a668a <=( a81584a  and  a81569a );
 a669a <=( a81556a  and  a81541a );
 a670a <=( a81528a  and  a81513a );
 a671a <=( a81500a  and  a81485a );
 a672a <=( a81472a  and  a81457a );
 a673a <=( a81444a  and  a81429a );
 a674a <=( a81416a  and  a81401a );
 a675a <=( a81388a  and  a81373a );
 a676a <=( a81360a  and  a81345a );
 a677a <=( a81332a  and  a81317a );
 a678a <=( a81304a  and  a81289a );
 a679a <=( a81276a  and  a81261a );
 a680a <=( a81248a  and  a81233a );
 a681a <=( a81220a  and  a81205a );
 a682a <=( a81192a  and  a81177a );
 a683a <=( a81164a  and  a81149a );
 a684a <=( a81136a  and  a81121a );
 a685a <=( a81108a  and  a81093a );
 a686a <=( a81080a  and  a81065a );
 a687a <=( a81052a  and  a81037a );
 a688a <=( a81024a  and  a81009a );
 a689a <=( a80996a  and  a80981a );
 a690a <=( a80968a  and  a80953a );
 a691a <=( a80940a  and  a80925a );
 a692a <=( a80912a  and  a80897a );
 a693a <=( a80884a  and  a80869a );
 a694a <=( a80856a  and  a80841a );
 a695a <=( a80828a  and  a80813a );
 a696a <=( a80800a  and  a80785a );
 a697a <=( a80772a  and  a80757a );
 a698a <=( a80744a  and  a80729a );
 a699a <=( a80716a  and  a80701a );
 a700a <=( a80688a  and  a80673a );
 a701a <=( a80660a  and  a80645a );
 a702a <=( a80632a  and  a80617a );
 a703a <=( a80604a  and  a80589a );
 a704a <=( a80576a  and  a80561a );
 a705a <=( a80548a  and  a80533a );
 a706a <=( a80520a  and  a80505a );
 a707a <=( a80492a  and  a80477a );
 a708a <=( a80464a  and  a80449a );
 a709a <=( a80436a  and  a80421a );
 a710a <=( a80408a  and  a80393a );
 a711a <=( a80380a  and  a80365a );
 a712a <=( a80352a  and  a80337a );
 a713a <=( a80324a  and  a80309a );
 a714a <=( a80296a  and  a80281a );
 a715a <=( a80268a  and  a80253a );
 a716a <=( a80240a  and  a80225a );
 a717a <=( a80212a  and  a80197a );
 a718a <=( a80184a  and  a80169a );
 a719a <=( a80156a  and  a80141a );
 a720a <=( a80128a  and  a80113a );
 a721a <=( a80100a  and  a80085a );
 a722a <=( a80072a  and  a80057a );
 a723a <=( a80044a  and  a80029a );
 a724a <=( a80016a  and  a80001a );
 a725a <=( a79988a  and  a79973a );
 a726a <=( a79960a  and  a79945a );
 a727a <=( a79932a  and  a79917a );
 a728a <=( a79904a  and  a79889a );
 a729a <=( a79876a  and  a79861a );
 a730a <=( a79848a  and  a79833a );
 a731a <=( a79820a  and  a79805a );
 a732a <=( a79792a  and  a79777a );
 a733a <=( a79764a  and  a79749a );
 a734a <=( a79736a  and  a79721a );
 a735a <=( a79708a  and  a79693a );
 a736a <=( a79680a  and  a79665a );
 a737a <=( a79652a  and  a79637a );
 a738a <=( a79624a  and  a79609a );
 a739a <=( a79596a  and  a79581a );
 a740a <=( a79568a  and  a79553a );
 a741a <=( a79540a  and  a79525a );
 a742a <=( a79512a  and  a79497a );
 a743a <=( a79484a  and  a79469a );
 a744a <=( a79456a  and  a79441a );
 a745a <=( a79428a  and  a79413a );
 a746a <=( a79400a  and  a79385a );
 a747a <=( a79372a  and  a79357a );
 a748a <=( a79344a  and  a79329a );
 a749a <=( a79316a  and  a79301a );
 a750a <=( a79288a  and  a79273a );
 a751a <=( a79260a  and  a79245a );
 a752a <=( a79232a  and  a79217a );
 a753a <=( a79204a  and  a79189a );
 a754a <=( a79176a  and  a79161a );
 a755a <=( a79148a  and  a79133a );
 a756a <=( a79120a  and  a79105a );
 a757a <=( a79092a  and  a79077a );
 a758a <=( a79064a  and  a79049a );
 a759a <=( a79036a  and  a79021a );
 a760a <=( a79008a  and  a78993a );
 a761a <=( a78980a  and  a78965a );
 a762a <=( a78952a  and  a78937a );
 a763a <=( a78924a  and  a78909a );
 a764a <=( a78896a  and  a78881a );
 a765a <=( a78868a  and  a78853a );
 a766a <=( a78840a  and  a78825a );
 a767a <=( a78812a  and  a78797a );
 a768a <=( a78784a  and  a78769a );
 a769a <=( a78756a  and  a78741a );
 a770a <=( a78728a  and  a78713a );
 a771a <=( a78700a  and  a78685a );
 a772a <=( a78672a  and  a78657a );
 a773a <=( a78644a  and  a78629a );
 a774a <=( a78616a  and  a78601a );
 a775a <=( a78588a  and  a78573a );
 a776a <=( a78560a  and  a78545a );
 a777a <=( a78532a  and  a78517a );
 a778a <=( a78504a  and  a78489a );
 a779a <=( a78476a  and  a78461a );
 a780a <=( a78448a  and  a78433a );
 a781a <=( a78420a  and  a78405a );
 a782a <=( a78392a  and  a78377a );
 a783a <=( a78364a  and  a78349a );
 a784a <=( a78336a  and  a78321a );
 a785a <=( a78308a  and  a78293a );
 a786a <=( a78280a  and  a78265a );
 a787a <=( a78252a  and  a78237a );
 a788a <=( a78224a  and  a78209a );
 a789a <=( a78196a  and  a78181a );
 a790a <=( a78168a  and  a78153a );
 a791a <=( a78140a  and  a78125a );
 a792a <=( a78112a  and  a78097a );
 a793a <=( a78084a  and  a78069a );
 a794a <=( a78056a  and  a78041a );
 a795a <=( a78028a  and  a78013a );
 a796a <=( a78000a  and  a77985a );
 a797a <=( a77972a  and  a77957a );
 a798a <=( a77944a  and  a77929a );
 a799a <=( a77916a  and  a77901a );
 a800a <=( a77888a  and  a77873a );
 a801a <=( a77860a  and  a77845a );
 a802a <=( a77832a  and  a77817a );
 a803a <=( a77804a  and  a77789a );
 a804a <=( a77776a  and  a77761a );
 a805a <=( a77748a  and  a77733a );
 a806a <=( a77720a  and  a77705a );
 a807a <=( a77692a  and  a77677a );
 a808a <=( a77664a  and  a77649a );
 a809a <=( a77636a  and  a77621a );
 a810a <=( a77608a  and  a77593a );
 a811a <=( a77580a  and  a77565a );
 a812a <=( a77552a  and  a77537a );
 a813a <=( a77524a  and  a77509a );
 a814a <=( a77496a  and  a77481a );
 a815a <=( a77468a  and  a77453a );
 a816a <=( a77440a  and  a77425a );
 a817a <=( a77412a  and  a77397a );
 a818a <=( a77384a  and  a77369a );
 a819a <=( a77356a  and  a77341a );
 a820a <=( a77328a  and  a77313a );
 a821a <=( a77300a  and  a77285a );
 a822a <=( a77272a  and  a77257a );
 a823a <=( a77244a  and  a77229a );
 a824a <=( a77216a  and  a77201a );
 a825a <=( a77188a  and  a77173a );
 a826a <=( a77160a  and  a77145a );
 a827a <=( a77132a  and  a77117a );
 a828a <=( a77104a  and  a77089a );
 a829a <=( a77076a  and  a77061a );
 a830a <=( a77048a  and  a77033a );
 a831a <=( a77020a  and  a77005a );
 a832a <=( a76992a  and  a76977a );
 a833a <=( a76964a  and  a76949a );
 a834a <=( a76936a  and  a76921a );
 a835a <=( a76908a  and  a76893a );
 a836a <=( a76880a  and  a76865a );
 a837a <=( a76852a  and  a76837a );
 a838a <=( a76824a  and  a76809a );
 a839a <=( a76796a  and  a76781a );
 a840a <=( a76768a  and  a76753a );
 a841a <=( a76740a  and  a76725a );
 a842a <=( a76712a  and  a76697a );
 a843a <=( a76684a  and  a76669a );
 a844a <=( a76656a  and  a76641a );
 a845a <=( a76628a  and  a76613a );
 a846a <=( a76600a  and  a76585a );
 a847a <=( a76572a  and  a76557a );
 a848a <=( a76544a  and  a76529a );
 a849a <=( a76516a  and  a76501a );
 a850a <=( a76488a  and  a76473a );
 a851a <=( a76460a  and  a76445a );
 a852a <=( a76432a  and  a76417a );
 a853a <=( a76404a  and  a76389a );
 a854a <=( a76376a  and  a76361a );
 a855a <=( a76348a  and  a76333a );
 a856a <=( a76320a  and  a76305a );
 a857a <=( a76292a  and  a76277a );
 a858a <=( a76264a  and  a76249a );
 a859a <=( a76236a  and  a76221a );
 a860a <=( a76208a  and  a76193a );
 a861a <=( a76180a  and  a76165a );
 a862a <=( a76152a  and  a76137a );
 a863a <=( a76124a  and  a76109a );
 a864a <=( a76096a  and  a76081a );
 a865a <=( a76068a  and  a76053a );
 a866a <=( a76040a  and  a76025a );
 a867a <=( a76012a  and  a75997a );
 a868a <=( a75984a  and  a75969a );
 a869a <=( a75956a  and  a75941a );
 a870a <=( a75928a  and  a75913a );
 a871a <=( a75900a  and  a75885a );
 a872a <=( a75872a  and  a75857a );
 a873a <=( a75844a  and  a75829a );
 a874a <=( a75816a  and  a75801a );
 a875a <=( a75788a  and  a75773a );
 a876a <=( a75760a  and  a75745a );
 a877a <=( a75732a  and  a75717a );
 a878a <=( a75704a  and  a75689a );
 a879a <=( a75676a  and  a75661a );
 a880a <=( a75648a  and  a75633a );
 a881a <=( a75620a  and  a75605a );
 a882a <=( a75592a  and  a75577a );
 a883a <=( a75564a  and  a75549a );
 a884a <=( a75536a  and  a75521a );
 a885a <=( a75508a  and  a75493a );
 a886a <=( a75480a  and  a75465a );
 a887a <=( a75452a  and  a75437a );
 a888a <=( a75424a  and  a75409a );
 a889a <=( a75396a  and  a75381a );
 a890a <=( a75368a  and  a75353a );
 a891a <=( a75340a  and  a75325a );
 a892a <=( a75312a  and  a75297a );
 a893a <=( a75284a  and  a75269a );
 a894a <=( a75256a  and  a75241a );
 a895a <=( a75228a  and  a75213a );
 a896a <=( a75200a  and  a75185a );
 a897a <=( a75172a  and  a75157a );
 a898a <=( a75144a  and  a75129a );
 a899a <=( a75116a  and  a75101a );
 a900a <=( a75088a  and  a75073a );
 a901a <=( a75060a  and  a75045a );
 a902a <=( a75032a  and  a75017a );
 a903a <=( a75004a  and  a74989a );
 a904a <=( a74976a  and  a74961a );
 a905a <=( a74948a  and  a74933a );
 a906a <=( a74920a  and  a74905a );
 a907a <=( a74892a  and  a74877a );
 a908a <=( a74864a  and  a74849a );
 a909a <=( a74836a  and  a74821a );
 a910a <=( a74808a  and  a74793a );
 a911a <=( a74780a  and  a74765a );
 a912a <=( a74752a  and  a74737a );
 a913a <=( a74724a  and  a74709a );
 a914a <=( a74696a  and  a74681a );
 a915a <=( a74668a  and  a74653a );
 a916a <=( a74640a  and  a74625a );
 a917a <=( a74612a  and  a74597a );
 a918a <=( a74584a  and  a74569a );
 a919a <=( a74556a  and  a74541a );
 a920a <=( a74528a  and  a74513a );
 a921a <=( a74500a  and  a74485a );
 a922a <=( a74472a  and  a74457a );
 a923a <=( a74444a  and  a74429a );
 a924a <=( a74416a  and  a74401a );
 a925a <=( a74388a  and  a74373a );
 a926a <=( a74360a  and  a74345a );
 a927a <=( a74332a  and  a74317a );
 a928a <=( a74304a  and  a74289a );
 a929a <=( a74276a  and  a74263a );
 a930a <=( a74250a  and  a74237a );
 a931a <=( a74224a  and  a74211a );
 a932a <=( a74198a  and  a74185a );
 a933a <=( a74172a  and  a74159a );
 a934a <=( a74146a  and  a74133a );
 a935a <=( a74120a  and  a74107a );
 a936a <=( a74094a  and  a74081a );
 a937a <=( a74068a  and  a74055a );
 a938a <=( a74042a  and  a74029a );
 a939a <=( a74016a  and  a74003a );
 a940a <=( a73990a  and  a73977a );
 a941a <=( a73964a  and  a73951a );
 a942a <=( a73938a  and  a73925a );
 a943a <=( a73912a  and  a73899a );
 a944a <=( a73886a  and  a73873a );
 a945a <=( a73860a  and  a73847a );
 a946a <=( a73834a  and  a73821a );
 a947a <=( a73808a  and  a73795a );
 a948a <=( a73782a  and  a73769a );
 a949a <=( a73756a  and  a73743a );
 a950a <=( a73730a  and  a73717a );
 a951a <=( a73704a  and  a73691a );
 a952a <=( a73678a  and  a73665a );
 a953a <=( a73652a  and  a73639a );
 a954a <=( a73626a  and  a73613a );
 a955a <=( a73600a  and  a73587a );
 a956a <=( a73574a  and  a73561a );
 a957a <=( a73548a  and  a73535a );
 a958a <=( a73522a  and  a73509a );
 a959a <=( a73496a  and  a73483a );
 a960a <=( a73470a  and  a73457a );
 a961a <=( a73444a  and  a73431a );
 a962a <=( a73418a  and  a73405a );
 a963a <=( a73392a  and  a73379a );
 a964a <=( a73366a  and  a73353a );
 a965a <=( a73340a  and  a73327a );
 a966a <=( a73314a  and  a73301a );
 a967a <=( a73288a  and  a73275a );
 a968a <=( a73262a  and  a73249a );
 a969a <=( a73236a  and  a73223a );
 a970a <=( a73210a  and  a73197a );
 a971a <=( a73184a  and  a73171a );
 a972a <=( a73158a  and  a73145a );
 a973a <=( a73132a  and  a73119a );
 a974a <=( a73106a  and  a73093a );
 a975a <=( a73080a  and  a73067a );
 a976a <=( a73054a  and  a73041a );
 a977a <=( a73028a  and  a73015a );
 a978a <=( a73002a  and  a72989a );
 a979a <=( a72976a  and  a72963a );
 a980a <=( a72950a  and  a72937a );
 a981a <=( a72924a  and  a72911a );
 a982a <=( a72898a  and  a72885a );
 a983a <=( a72872a  and  a72859a );
 a984a <=( a72846a  and  a72833a );
 a985a <=( a72820a  and  a72807a );
 a986a <=( a72794a  and  a72781a );
 a987a <=( a72768a  and  a72755a );
 a988a <=( a72742a  and  a72729a );
 a989a <=( a72716a  and  a72703a );
 a990a <=( a72690a  and  a72677a );
 a991a <=( a72664a  and  a72651a );
 a992a <=( a72638a  and  a72625a );
 a993a <=( a72612a  and  a72599a );
 a994a <=( a72586a  and  a72573a );
 a995a <=( a72560a  and  a72547a );
 a996a <=( a72534a  and  a72521a );
 a997a <=( a72508a  and  a72495a );
 a998a <=( a72482a  and  a72469a );
 a999a <=( a72456a  and  a72443a );
 a1000a <=( a72430a  and  a72417a );
 a1001a <=( a72404a  and  a72391a );
 a1002a <=( a72378a  and  a72365a );
 a1003a <=( a72352a  and  a72339a );
 a1004a <=( a72326a  and  a72313a );
 a1005a <=( a72300a  and  a72287a );
 a1006a <=( a72274a  and  a72261a );
 a1007a <=( a72248a  and  a72235a );
 a1008a <=( a72222a  and  a72209a );
 a1009a <=( a72196a  and  a72183a );
 a1010a <=( a72170a  and  a72157a );
 a1011a <=( a72144a  and  a72131a );
 a1012a <=( a72118a  and  a72105a );
 a1013a <=( a72092a  and  a72079a );
 a1014a <=( a72066a  and  a72053a );
 a1015a <=( a72040a  and  a72027a );
 a1016a <=( a72014a  and  a72001a );
 a1017a <=( a71988a  and  a71975a );
 a1018a <=( a71962a  and  a71949a );
 a1019a <=( a71936a  and  a71923a );
 a1020a <=( a71910a  and  a71897a );
 a1021a <=( a71884a  and  a71871a );
 a1022a <=( a71858a  and  a71845a );
 a1023a <=( a71832a  and  a71819a );
 a1024a <=( a71806a  and  a71793a );
 a1025a <=( a71780a  and  a71767a );
 a1026a <=( a71754a  and  a71741a );
 a1027a <=( a71728a  and  a71715a );
 a1028a <=( a71702a  and  a71689a );
 a1029a <=( a71676a  and  a71663a );
 a1030a <=( a71650a  and  a71637a );
 a1031a <=( a71624a  and  a71611a );
 a1032a <=( a71598a  and  a71585a );
 a1033a <=( a71572a  and  a71559a );
 a1034a <=( a71546a  and  a71533a );
 a1035a <=( a71520a  and  a71507a );
 a1036a <=( a71494a  and  a71481a );
 a1037a <=( a71468a  and  a71455a );
 a1038a <=( a71442a  and  a71429a );
 a1039a <=( a71416a  and  a71403a );
 a1040a <=( a71390a  and  a71377a );
 a1041a <=( a71364a  and  a71351a );
 a1042a <=( a71338a  and  a71325a );
 a1043a <=( a71312a  and  a71299a );
 a1044a <=( a71286a  and  a71273a );
 a1045a <=( a71260a  and  a71247a );
 a1046a <=( a71234a  and  a71221a );
 a1047a <=( a71208a  and  a71195a );
 a1048a <=( a71182a  and  a71169a );
 a1049a <=( a71156a  and  a71143a );
 a1050a <=( a71130a  and  a71117a );
 a1051a <=( a71104a  and  a71091a );
 a1052a <=( a71078a  and  a71065a );
 a1053a <=( a71052a  and  a71039a );
 a1054a <=( a71026a  and  a71013a );
 a1055a <=( a71000a  and  a70987a );
 a1056a <=( a70974a  and  a70961a );
 a1057a <=( a70948a  and  a70935a );
 a1058a <=( a70922a  and  a70909a );
 a1059a <=( a70896a  and  a70883a );
 a1060a <=( a70870a  and  a70857a );
 a1061a <=( a70844a  and  a70831a );
 a1062a <=( a70818a  and  a70805a );
 a1063a <=( a70792a  and  a70779a );
 a1064a <=( a70766a  and  a70753a );
 a1065a <=( a70740a  and  a70727a );
 a1066a <=( a70714a  and  a70701a );
 a1067a <=( a70688a  and  a70675a );
 a1068a <=( a70662a  and  a70649a );
 a1069a <=( a70636a  and  a70623a );
 a1070a <=( a70610a  and  a70597a );
 a1071a <=( a70584a  and  a70571a );
 a1072a <=( a70558a  and  a70545a );
 a1073a <=( a70532a  and  a70519a );
 a1074a <=( a70506a  and  a70493a );
 a1075a <=( a70480a  and  a70467a );
 a1076a <=( a70454a  and  a70441a );
 a1077a <=( a70428a  and  a70415a );
 a1078a <=( a70402a  and  a70389a );
 a1079a <=( a70376a  and  a70363a );
 a1080a <=( a70350a  and  a70337a );
 a1081a <=( a70324a  and  a70311a );
 a1082a <=( a70298a  and  a70285a );
 a1083a <=( a70272a  and  a70259a );
 a1084a <=( a70246a  and  a70233a );
 a1085a <=( a70220a  and  a70207a );
 a1086a <=( a70194a  and  a70181a );
 a1087a <=( a70168a  and  a70155a );
 a1088a <=( a70142a  and  a70129a );
 a1089a <=( a70116a  and  a70103a );
 a1090a <=( a70090a  and  a70077a );
 a1091a <=( a70064a  and  a70051a );
 a1092a <=( a70038a  and  a70025a );
 a1093a <=( a70012a  and  a69999a );
 a1094a <=( a69986a  and  a69973a );
 a1095a <=( a69960a  and  a69947a );
 a1096a <=( a69934a  and  a69921a );
 a1097a <=( a69908a  and  a69895a );
 a1098a <=( a69882a  and  a69869a );
 a1099a <=( a69856a  and  a69843a );
 a1100a <=( a69830a  and  a69817a );
 a1101a <=( a69804a  and  a69791a );
 a1102a <=( a69778a  and  a69765a );
 a1103a <=( a69752a  and  a69739a );
 a1104a <=( a69726a  and  a69713a );
 a1105a <=( a69700a  and  a69687a );
 a1106a <=( a69674a  and  a69661a );
 a1107a <=( a69648a  and  a69635a );
 a1108a <=( a69622a  and  a69609a );
 a1109a <=( a69596a  and  a69583a );
 a1110a <=( a69570a  and  a69557a );
 a1111a <=( a69544a  and  a69531a );
 a1112a <=( a69518a  and  a69505a );
 a1113a <=( a69492a  and  a69479a );
 a1114a <=( a69466a  and  a69453a );
 a1115a <=( a69440a  and  a69427a );
 a1116a <=( a69414a  and  a69401a );
 a1117a <=( a69388a  and  a69375a );
 a1118a <=( a69362a  and  a69349a );
 a1119a <=( a69336a  and  a69323a );
 a1120a <=( a69310a  and  a69297a );
 a1121a <=( a69284a  and  a69271a );
 a1122a <=( a69258a  and  a69245a );
 a1123a <=( a69232a  and  a69219a );
 a1124a <=( a69206a  and  a69193a );
 a1125a <=( a69180a  and  a69167a );
 a1126a <=( a69154a  and  a69141a );
 a1127a <=( a69128a  and  a69115a );
 a1128a <=( a69102a  and  a69089a );
 a1129a <=( a69076a  and  a69063a );
 a1130a <=( a69050a  and  a69037a );
 a1131a <=( a69024a  and  a69011a );
 a1132a <=( a68998a  and  a68985a );
 a1133a <=( a68972a  and  a68959a );
 a1134a <=( a68946a  and  a68933a );
 a1135a <=( a68920a  and  a68907a );
 a1136a <=( a68894a  and  a68881a );
 a1137a <=( a68868a  and  a68855a );
 a1138a <=( a68842a  and  a68829a );
 a1139a <=( a68816a  and  a68803a );
 a1140a <=( a68790a  and  a68777a );
 a1141a <=( a68764a  and  a68751a );
 a1142a <=( a68738a  and  a68725a );
 a1143a <=( a68712a  and  a68699a );
 a1144a <=( a68686a  and  a68673a );
 a1145a <=( a68660a  and  a68647a );
 a1146a <=( a68634a  and  a68621a );
 a1147a <=( a68608a  and  a68595a );
 a1148a <=( a68582a  and  a68569a );
 a1149a <=( a68556a  and  a68543a );
 a1150a <=( a68530a  and  a68517a );
 a1151a <=( a68504a  and  a68491a );
 a1152a <=( a68478a  and  a68465a );
 a1153a <=( a68452a  and  a68439a );
 a1154a <=( a68426a  and  a68413a );
 a1155a <=( a68400a  and  a68387a );
 a1156a <=( a68374a  and  a68361a );
 a1157a <=( a68348a  and  a68335a );
 a1158a <=( a68322a  and  a68309a );
 a1159a <=( a68296a  and  a68283a );
 a1160a <=( a68270a  and  a68257a );
 a1161a <=( a68244a  and  a68231a );
 a1162a <=( a68218a  and  a68205a );
 a1163a <=( a68192a  and  a68179a );
 a1164a <=( a68166a  and  a68153a );
 a1165a <=( a68140a  and  a68127a );
 a1166a <=( a68114a  and  a68101a );
 a1167a <=( a68088a  and  a68075a );
 a1168a <=( a68062a  and  a68049a );
 a1169a <=( a68036a  and  a68023a );
 a1170a <=( a68010a  and  a67997a );
 a1171a <=( a67984a  and  a67971a );
 a1172a <=( a67958a  and  a67945a );
 a1173a <=( a67932a  and  a67919a );
 a1174a <=( a67906a  and  a67893a );
 a1175a <=( a67880a  and  a67867a );
 a1176a <=( a67854a  and  a67841a );
 a1177a <=( a67828a  and  a67815a );
 a1178a <=( a67802a  and  a67789a );
 a1179a <=( a67776a  and  a67763a );
 a1180a <=( a67750a  and  a67737a );
 a1181a <=( a67724a  and  a67711a );
 a1182a <=( a67698a  and  a67685a );
 a1183a <=( a67672a  and  a67659a );
 a1184a <=( a67646a  and  a67633a );
 a1185a <=( a67620a  and  a67607a );
 a1186a <=( a67594a  and  a67581a );
 a1187a <=( a67568a  and  a67555a );
 a1188a <=( a67542a  and  a67529a );
 a1189a <=( a67516a  and  a67503a );
 a1190a <=( a67490a  and  a67477a );
 a1191a <=( a67464a  and  a67451a );
 a1192a <=( a67438a  and  a67425a );
 a1193a <=( a67412a  and  a67399a );
 a1194a <=( a67386a  and  a67373a );
 a1195a <=( a67360a  and  a67347a );
 a1196a <=( a67334a  and  a67321a );
 a1197a <=( a67308a  and  a67295a );
 a1198a <=( a67282a  and  a67269a );
 a1199a <=( a67256a  and  a67243a );
 a1200a <=( a67230a  and  a67217a );
 a1201a <=( a67204a  and  a67191a );
 a1202a <=( a67178a  and  a67165a );
 a1203a <=( a67152a  and  a67139a );
 a1204a <=( a67126a  and  a67113a );
 a1205a <=( a67100a  and  a67087a );
 a1206a <=( a67074a  and  a67061a );
 a1207a <=( a67048a  and  a67035a );
 a1208a <=( a67022a  and  a67009a );
 a1209a <=( a66996a  and  a66983a );
 a1210a <=( a66970a  and  a66957a );
 a1211a <=( a66944a  and  a66931a );
 a1212a <=( a66918a  and  a66905a );
 a1213a <=( a66892a  and  a66879a );
 a1214a <=( a66866a  and  a66853a );
 a1215a <=( a66840a  and  a66827a );
 a1216a <=( a66814a  and  a66801a );
 a1217a <=( a66788a  and  a66775a );
 a1218a <=( a66762a  and  a66749a );
 a1219a <=( a66736a  and  a66723a );
 a1220a <=( a66710a  and  a66697a );
 a1221a <=( a66684a  and  a66671a );
 a1222a <=( a66658a  and  a66645a );
 a1223a <=( a66632a  and  a66619a );
 a1224a <=( a66606a  and  a66593a );
 a1225a <=( a66580a  and  a66567a );
 a1226a <=( a66554a  and  a66541a );
 a1227a <=( a66528a  and  a66515a );
 a1228a <=( a66502a  and  a66489a );
 a1229a <=( a66476a  and  a66463a );
 a1230a <=( a66450a  and  a66437a );
 a1231a <=( a66424a  and  a66411a );
 a1232a <=( a66398a  and  a66385a );
 a1233a <=( a66372a  and  a66359a );
 a1234a <=( a66346a  and  a66333a );
 a1235a <=( a66320a  and  a66307a );
 a1236a <=( a66294a  and  a66281a );
 a1237a <=( a66268a  and  a66255a );
 a1238a <=( a66242a  and  a66229a );
 a1239a <=( a66216a  and  a66203a );
 a1240a <=( a66190a  and  a66177a );
 a1241a <=( a66164a  and  a66151a );
 a1242a <=( a66138a  and  a66125a );
 a1243a <=( a66112a  and  a66099a );
 a1244a <=( a66086a  and  a66073a );
 a1245a <=( a66060a  and  a66047a );
 a1246a <=( a66034a  and  a66021a );
 a1247a <=( a66008a  and  a65995a );
 a1248a <=( a65982a  and  a65969a );
 a1249a <=( a65956a  and  a65943a );
 a1250a <=( a65930a  and  a65917a );
 a1251a <=( a65904a  and  a65891a );
 a1252a <=( a65878a  and  a65865a );
 a1253a <=( a65852a  and  a65839a );
 a1254a <=( a65826a  and  a65813a );
 a1255a <=( a65800a  and  a65787a );
 a1256a <=( a65774a  and  a65761a );
 a1257a <=( a65748a  and  a65735a );
 a1258a <=( a65722a  and  a65709a );
 a1259a <=( a65696a  and  a65683a );
 a1260a <=( a65670a  and  a65657a );
 a1261a <=( a65644a  and  a65631a );
 a1262a <=( a65618a  and  a65605a );
 a1263a <=( a65592a  and  a65579a );
 a1264a <=( a65566a  and  a65553a );
 a1265a <=( a65540a  and  a65527a );
 a1266a <=( a65514a  and  a65501a );
 a1267a <=( a65488a  and  a65475a );
 a1268a <=( a65462a  and  a65449a );
 a1269a <=( a65436a  and  a65423a );
 a1270a <=( a65410a  and  a65397a );
 a1271a <=( a65384a  and  a65371a );
 a1272a <=( a65358a  and  a65345a );
 a1273a <=( a65332a  and  a65319a );
 a1274a <=( a65306a  and  a65293a );
 a1275a <=( a65280a  and  a65267a );
 a1276a <=( a65254a  and  a65241a );
 a1277a <=( a65228a  and  a65215a );
 a1278a <=( a65202a  and  a65189a );
 a1279a <=( a65176a  and  a65163a );
 a1280a <=( a65150a  and  a65137a );
 a1281a <=( a65124a  and  a65111a );
 a1282a <=( a65098a  and  a65085a );
 a1283a <=( a65072a  and  a65059a );
 a1284a <=( a65046a  and  a65033a );
 a1285a <=( a65020a  and  a65007a );
 a1286a <=( a64994a  and  a64981a );
 a1287a <=( a64968a  and  a64955a );
 a1288a <=( a64942a  and  a64929a );
 a1289a <=( a64916a  and  a64903a );
 a1290a <=( a64890a  and  a64877a );
 a1291a <=( a64864a  and  a64851a );
 a1292a <=( a64838a  and  a64825a );
 a1293a <=( a64812a  and  a64799a );
 a1294a <=( a64786a  and  a64773a );
 a1295a <=( a64760a  and  a64747a );
 a1296a <=( a64734a  and  a64721a );
 a1297a <=( a64708a  and  a64695a );
 a1298a <=( a64682a  and  a64669a );
 a1299a <=( a64656a  and  a64643a );
 a1300a <=( a64630a  and  a64617a );
 a1301a <=( a64604a  and  a64591a );
 a1302a <=( a64578a  and  a64565a );
 a1303a <=( a64552a  and  a64539a );
 a1304a <=( a64526a  and  a64513a );
 a1305a <=( a64500a  and  a64487a );
 a1306a <=( a64474a  and  a64461a );
 a1307a <=( a64448a  and  a64435a );
 a1308a <=( a64422a  and  a64409a );
 a1309a <=( a64396a  and  a64383a );
 a1310a <=( a64370a  and  a64357a );
 a1311a <=( a64344a  and  a64331a );
 a1312a <=( a64318a  and  a64305a );
 a1313a <=( a64292a  and  a64279a );
 a1314a <=( a64266a  and  a64253a );
 a1315a <=( a64240a  and  a64227a );
 a1316a <=( a64214a  and  a64201a );
 a1317a <=( a64188a  and  a64175a );
 a1318a <=( a64162a  and  a64149a );
 a1319a <=( a64136a  and  a64123a );
 a1320a <=( a64110a  and  a64097a );
 a1321a <=( a64084a  and  a64071a );
 a1322a <=( a64058a  and  a64045a );
 a1323a <=( a64032a  and  a64019a );
 a1324a <=( a64006a  and  a63993a );
 a1325a <=( a63980a  and  a63967a );
 a1326a <=( a63954a  and  a63941a );
 a1327a <=( a63928a  and  a63915a );
 a1328a <=( a63902a  and  a63889a );
 a1329a <=( a63876a  and  a63863a );
 a1330a <=( a63850a  and  a63837a );
 a1331a <=( a63824a  and  a63811a );
 a1332a <=( a63798a  and  a63785a );
 a1333a <=( a63772a  and  a63759a );
 a1334a <=( a63746a  and  a63733a );
 a1335a <=( a63720a  and  a63707a );
 a1336a <=( a63694a  and  a63681a );
 a1337a <=( a63668a  and  a63655a );
 a1338a <=( a63642a  and  a63629a );
 a1339a <=( a63616a  and  a63603a );
 a1340a <=( a63590a  and  a63577a );
 a1341a <=( a63564a  and  a63551a );
 a1342a <=( a63538a  and  a63525a );
 a1343a <=( a63512a  and  a63499a );
 a1344a <=( a63486a  and  a63473a );
 a1345a <=( a63460a  and  a63447a );
 a1346a <=( a63434a  and  a63421a );
 a1347a <=( a63408a  and  a63395a );
 a1348a <=( a63382a  and  a63369a );
 a1349a <=( a63356a  and  a63343a );
 a1350a <=( a63330a  and  a63317a );
 a1351a <=( a63304a  and  a63291a );
 a1352a <=( a63278a  and  a63265a );
 a1353a <=( a63252a  and  a63239a );
 a1354a <=( a63226a  and  a63213a );
 a1355a <=( a63200a  and  a63187a );
 a1356a <=( a63174a  and  a63161a );
 a1357a <=( a63148a  and  a63135a );
 a1358a <=( a63122a  and  a63109a );
 a1359a <=( a63096a  and  a63083a );
 a1360a <=( a63070a  and  a63057a );
 a1361a <=( a63044a  and  a63031a );
 a1362a <=( a63018a  and  a63005a );
 a1363a <=( a62992a  and  a62979a );
 a1364a <=( a62966a  and  a62953a );
 a1365a <=( a62940a  and  a62927a );
 a1366a <=( a62914a  and  a62901a );
 a1367a <=( a62888a  and  a62875a );
 a1368a <=( a62862a  and  a62849a );
 a1369a <=( a62836a  and  a62823a );
 a1370a <=( a62810a  and  a62797a );
 a1371a <=( a62784a  and  a62771a );
 a1372a <=( a62758a  and  a62745a );
 a1373a <=( a62732a  and  a62719a );
 a1374a <=( a62706a  and  a62693a );
 a1375a <=( a62680a  and  a62667a );
 a1376a <=( a62654a  and  a62641a );
 a1377a <=( a62628a  and  a62615a );
 a1378a <=( a62602a  and  a62589a );
 a1379a <=( a62576a  and  a62563a );
 a1380a <=( a62550a  and  a62537a );
 a1381a <=( a62524a  and  a62511a );
 a1382a <=( a62498a  and  a62485a );
 a1383a <=( a62472a  and  a62459a );
 a1384a <=( a62446a  and  a62433a );
 a1385a <=( a62420a  and  a62407a );
 a1386a <=( a62394a  and  a62381a );
 a1387a <=( a62368a  and  a62355a );
 a1388a <=( a62342a  and  a62329a );
 a1389a <=( a62316a  and  a62303a );
 a1390a <=( a62290a  and  a62277a );
 a1391a <=( a62264a  and  a62251a );
 a1392a <=( a62238a  and  a62225a );
 a1393a <=( a62212a  and  a62199a );
 a1394a <=( a62186a  and  a62173a );
 a1395a <=( a62160a  and  a62147a );
 a1396a <=( a62134a  and  a62121a );
 a1397a <=( a62108a  and  a62095a );
 a1398a <=( a62082a  and  a62069a );
 a1399a <=( a62056a  and  a62043a );
 a1400a <=( a62030a  and  a62017a );
 a1401a <=( a62004a  and  a61991a );
 a1402a <=( a61978a  and  a61965a );
 a1403a <=( a61952a  and  a61939a );
 a1404a <=( a61926a  and  a61913a );
 a1405a <=( a61900a  and  a61887a );
 a1406a <=( a61874a  and  a61861a );
 a1407a <=( a61848a  and  a61835a );
 a1408a <=( a61822a  and  a61809a );
 a1409a <=( a61796a  and  a61783a );
 a1410a <=( a61770a  and  a61757a );
 a1411a <=( a61744a  and  a61731a );
 a1412a <=( a61718a  and  a61705a );
 a1413a <=( a61692a  and  a61679a );
 a1414a <=( a61666a  and  a61653a );
 a1415a <=( a61640a  and  a61627a );
 a1416a <=( a61614a  and  a61601a );
 a1417a <=( a61588a  and  a61575a );
 a1418a <=( a61562a  and  a61549a );
 a1419a <=( a61536a  and  a61523a );
 a1420a <=( a61510a  and  a61497a );
 a1421a <=( a61484a  and  a61471a );
 a1422a <=( a61458a  and  a61445a );
 a1423a <=( a61432a  and  a61419a );
 a1424a <=( a61406a  and  a61393a );
 a1425a <=( a61380a  and  a61367a );
 a1426a <=( a61354a  and  a61341a );
 a1427a <=( a61328a  and  a61315a );
 a1428a <=( a61302a  and  a61289a );
 a1429a <=( a61276a  and  a61263a );
 a1430a <=( a61250a  and  a61237a );
 a1431a <=( a61224a  and  a61211a );
 a1432a <=( a61198a  and  a61185a );
 a1433a <=( a61172a  and  a61159a );
 a1434a <=( a61146a  and  a61133a );
 a1435a <=( a61120a  and  a61107a );
 a1436a <=( a61094a  and  a61081a );
 a1437a <=( a61068a  and  a61055a );
 a1438a <=( a61042a  and  a61029a );
 a1439a <=( a61016a  and  a61003a );
 a1440a <=( a60990a  and  a60977a );
 a1441a <=( a60964a  and  a60951a );
 a1442a <=( a60938a  and  a60925a );
 a1443a <=( a60912a  and  a60899a );
 a1444a <=( a60886a  and  a60873a );
 a1445a <=( a60860a  and  a60847a );
 a1446a <=( a60834a  and  a60821a );
 a1447a <=( a60808a  and  a60795a );
 a1448a <=( a60782a  and  a60769a );
 a1449a <=( a60756a  and  a60743a );
 a1450a <=( a60730a  and  a60717a );
 a1451a <=( a60704a  and  a60691a );
 a1452a <=( a60678a  and  a60665a );
 a1453a <=( a60652a  and  a60639a );
 a1454a <=( a60626a  and  a60613a );
 a1455a <=( a60600a  and  a60587a );
 a1456a <=( a60574a  and  a60561a );
 a1457a <=( a60548a  and  a60535a );
 a1458a <=( a60522a  and  a60509a );
 a1459a <=( a60496a  and  a60483a );
 a1460a <=( a60470a  and  a60457a );
 a1461a <=( a60444a  and  a60431a );
 a1462a <=( a60418a  and  a60405a );
 a1463a <=( a60392a  and  a60379a );
 a1464a <=( a60366a  and  a60353a );
 a1465a <=( a60340a  and  a60327a );
 a1466a <=( a60314a  and  a60301a );
 a1467a <=( a60288a  and  a60275a );
 a1468a <=( a60262a  and  a60249a );
 a1469a <=( a60236a  and  a60223a );
 a1470a <=( a60210a  and  a60197a );
 a1471a <=( a60184a  and  a60171a );
 a1472a <=( a60158a  and  a60145a );
 a1473a <=( a60132a  and  a60119a );
 a1474a <=( a60106a  and  a60093a );
 a1475a <=( a60080a  and  a60067a );
 a1476a <=( a60054a  and  a60041a );
 a1477a <=( a60028a  and  a60015a );
 a1478a <=( a60002a  and  a59989a );
 a1479a <=( a59976a  and  a59963a );
 a1480a <=( a59950a  and  a59937a );
 a1481a <=( a59924a  and  a59911a );
 a1482a <=( a59898a  and  a59885a );
 a1483a <=( a59872a  and  a59859a );
 a1484a <=( a59846a  and  a59833a );
 a1485a <=( a59820a  and  a59807a );
 a1486a <=( a59794a  and  a59781a );
 a1487a <=( a59768a  and  a59755a );
 a1488a <=( a59742a  and  a59729a );
 a1489a <=( a59716a  and  a59703a );
 a1490a <=( a59690a  and  a59677a );
 a1491a <=( a59664a  and  a59651a );
 a1492a <=( a59638a  and  a59625a );
 a1493a <=( a59612a  and  a59599a );
 a1494a <=( a59586a  and  a59573a );
 a1495a <=( a59560a  and  a59547a );
 a1496a <=( a59534a  and  a59521a );
 a1497a <=( a59508a  and  a59495a );
 a1498a <=( a59482a  and  a59469a );
 a1499a <=( a59456a  and  a59443a );
 a1500a <=( a59430a  and  a59417a );
 a1501a <=( a59404a  and  a59391a );
 a1502a <=( a59378a  and  a59365a );
 a1503a <=( a59352a  and  a59339a );
 a1504a <=( a59326a  and  a59313a );
 a1505a <=( a59300a  and  a59287a );
 a1506a <=( a59274a  and  a59261a );
 a1507a <=( a59248a  and  a59235a );
 a1508a <=( a59222a  and  a59209a );
 a1509a <=( a59196a  and  a59183a );
 a1510a <=( a59170a  and  a59157a );
 a1511a <=( a59144a  and  a59131a );
 a1512a <=( a59118a  and  a59105a );
 a1513a <=( a59092a  and  a59079a );
 a1514a <=( a59066a  and  a59053a );
 a1515a <=( a59040a  and  a59027a );
 a1516a <=( a59014a  and  a59001a );
 a1517a <=( a58988a  and  a58975a );
 a1518a <=( a58962a  and  a58949a );
 a1519a <=( a58936a  and  a58923a );
 a1520a <=( a58910a  and  a58897a );
 a1521a <=( a58884a  and  a58871a );
 a1522a <=( a58858a  and  a58845a );
 a1523a <=( a58832a  and  a58819a );
 a1524a <=( a58806a  and  a58793a );
 a1525a <=( a58780a  and  a58767a );
 a1526a <=( a58754a  and  a58741a );
 a1527a <=( a58728a  and  a58715a );
 a1528a <=( a58702a  and  a58689a );
 a1529a <=( a58676a  and  a58663a );
 a1530a <=( a58650a  and  a58637a );
 a1531a <=( a58624a  and  a58611a );
 a1532a <=( a58598a  and  a58585a );
 a1533a <=( a58572a  and  a58559a );
 a1534a <=( a58546a  and  a58533a );
 a1535a <=( a58520a  and  a58507a );
 a1536a <=( a58494a  and  a58481a );
 a1537a <=( a58468a  and  a58455a );
 a1538a <=( a58442a  and  a58429a );
 a1539a <=( a58416a  and  a58403a );
 a1540a <=( a58390a  and  a58377a );
 a1541a <=( a58364a  and  a58351a );
 a1542a <=( a58338a  and  a58325a );
 a1543a <=( a58312a  and  a58299a );
 a1544a <=( a58286a  and  a58273a );
 a1545a <=( a58260a  and  a58247a );
 a1546a <=( a58234a  and  a58221a );
 a1547a <=( a58208a  and  a58195a );
 a1548a <=( a58182a  and  a58169a );
 a1549a <=( a58156a  and  a58143a );
 a1550a <=( a58130a  and  a58117a );
 a1551a <=( a58104a  and  a58091a );
 a1552a <=( a58078a  and  a58065a );
 a1553a <=( a58052a  and  a58039a );
 a1554a <=( a58026a  and  a58013a );
 a1555a <=( a58000a  and  a57987a );
 a1556a <=( a57974a  and  a57961a );
 a1557a <=( a57948a  and  a57935a );
 a1558a <=( a57922a  and  a57909a );
 a1559a <=( a57896a  and  a57883a );
 a1560a <=( a57870a  and  a57857a );
 a1561a <=( a57844a  and  a57831a );
 a1562a <=( a57818a  and  a57805a );
 a1563a <=( a57792a  and  a57779a );
 a1564a <=( a57766a  and  a57753a );
 a1565a <=( a57740a  and  a57727a );
 a1566a <=( a57714a  and  a57701a );
 a1567a <=( a57688a  and  a57675a );
 a1568a <=( a57662a  and  a57649a );
 a1569a <=( a57636a  and  a57623a );
 a1570a <=( a57610a  and  a57597a );
 a1571a <=( a57584a  and  a57571a );
 a1572a <=( a57558a  and  a57545a );
 a1573a <=( a57532a  and  a57519a );
 a1574a <=( a57506a  and  a57493a );
 a1575a <=( a57480a  and  a57467a );
 a1576a <=( a57454a  and  a57441a );
 a1577a <=( a57428a  and  a57415a );
 a1578a <=( a57402a  and  a57389a );
 a1579a <=( a57376a  and  a57363a );
 a1580a <=( a57350a  and  a57337a );
 a1581a <=( a57324a  and  a57311a );
 a1582a <=( a57298a  and  a57285a );
 a1583a <=( a57272a  and  a57259a );
 a1584a <=( a57246a  and  a57233a );
 a1585a <=( a57220a  and  a57207a );
 a1586a <=( a57194a  and  a57181a );
 a1587a <=( a57168a  and  a57155a );
 a1588a <=( a57142a  and  a57129a );
 a1589a <=( a57116a  and  a57103a );
 a1590a <=( a57090a  and  a57077a );
 a1591a <=( a57064a  and  a57051a );
 a1592a <=( a57038a  and  a57025a );
 a1593a <=( a57012a  and  a56999a );
 a1594a <=( a56986a  and  a56973a );
 a1595a <=( a56960a  and  a56947a );
 a1596a <=( a56934a  and  a56921a );
 a1597a <=( a56908a  and  a56895a );
 a1598a <=( a56882a  and  a56869a );
 a1599a <=( a56856a  and  a56843a );
 a1600a <=( a56830a  and  a56817a );
 a1601a <=( a56804a  and  a56791a );
 a1602a <=( a56778a  and  a56765a );
 a1603a <=( a56752a  and  a56739a );
 a1604a <=( a56728a  and  a56715a );
 a1605a <=( a56704a  and  a56691a );
 a1606a <=( a56680a  and  a56667a );
 a1607a <=( a56656a  and  a56643a );
 a1608a <=( a56632a  and  a56619a );
 a1609a <=( a56608a  and  a56595a );
 a1610a <=( a56584a  and  a56571a );
 a1611a <=( a56560a  and  a56547a );
 a1612a <=( a56536a  and  a56523a );
 a1613a <=( a56512a  and  a56499a );
 a1614a <=( a56488a  and  a56475a );
 a1615a <=( a56464a  and  a56451a );
 a1616a <=( a56440a  and  a56427a );
 a1617a <=( a56416a  and  a56403a );
 a1618a <=( a56392a  and  a56379a );
 a1619a <=( a56368a  and  a56355a );
 a1620a <=( a56344a  and  a56331a );
 a1621a <=( a56320a  and  a56307a );
 a1622a <=( a56296a  and  a56283a );
 a1623a <=( a56272a  and  a56259a );
 a1624a <=( a56248a  and  a56235a );
 a1625a <=( a56224a  and  a56211a );
 a1626a <=( a56200a  and  a56187a );
 a1627a <=( a56176a  and  a56163a );
 a1628a <=( a56152a  and  a56139a );
 a1629a <=( a56128a  and  a56115a );
 a1630a <=( a56104a  and  a56091a );
 a1631a <=( a56080a  and  a56067a );
 a1632a <=( a56056a  and  a56043a );
 a1633a <=( a56032a  and  a56019a );
 a1634a <=( a56008a  and  a55995a );
 a1635a <=( a55984a  and  a55971a );
 a1636a <=( a55960a  and  a55947a );
 a1637a <=( a55936a  and  a55923a );
 a1638a <=( a55912a  and  a55899a );
 a1639a <=( a55888a  and  a55875a );
 a1640a <=( a55864a  and  a55851a );
 a1641a <=( a55840a  and  a55827a );
 a1642a <=( a55816a  and  a55803a );
 a1643a <=( a55792a  and  a55779a );
 a1644a <=( a55768a  and  a55755a );
 a1645a <=( a55744a  and  a55731a );
 a1646a <=( a55720a  and  a55707a );
 a1647a <=( a55696a  and  a55683a );
 a1648a <=( a55672a  and  a55659a );
 a1649a <=( a55648a  and  a55635a );
 a1650a <=( a55624a  and  a55611a );
 a1651a <=( a55600a  and  a55587a );
 a1652a <=( a55576a  and  a55563a );
 a1653a <=( a55552a  and  a55539a );
 a1654a <=( a55528a  and  a55515a );
 a1655a <=( a55504a  and  a55491a );
 a1656a <=( a55480a  and  a55467a );
 a1657a <=( a55456a  and  a55443a );
 a1658a <=( a55432a  and  a55419a );
 a1659a <=( a55408a  and  a55395a );
 a1660a <=( a55384a  and  a55371a );
 a1661a <=( a55360a  and  a55347a );
 a1662a <=( a55336a  and  a55323a );
 a1663a <=( a55312a  and  a55299a );
 a1664a <=( a55288a  and  a55275a );
 a1665a <=( a55264a  and  a55251a );
 a1666a <=( a55240a  and  a55227a );
 a1667a <=( a55216a  and  a55203a );
 a1668a <=( a55192a  and  a55179a );
 a1669a <=( a55168a  and  a55155a );
 a1670a <=( a55144a  and  a55131a );
 a1671a <=( a55120a  and  a55107a );
 a1672a <=( a55096a  and  a55083a );
 a1673a <=( a55072a  and  a55059a );
 a1674a <=( a55048a  and  a55035a );
 a1675a <=( a55024a  and  a55011a );
 a1676a <=( a55000a  and  a54987a );
 a1677a <=( a54976a  and  a54963a );
 a1678a <=( a54952a  and  a54939a );
 a1679a <=( a54928a  and  a54915a );
 a1680a <=( a54904a  and  a54891a );
 a1681a <=( a54880a  and  a54867a );
 a1682a <=( a54856a  and  a54843a );
 a1683a <=( a54832a  and  a54819a );
 a1684a <=( a54808a  and  a54795a );
 a1685a <=( a54784a  and  a54771a );
 a1686a <=( a54760a  and  a54747a );
 a1687a <=( a54736a  and  a54723a );
 a1688a <=( a54712a  and  a54699a );
 a1689a <=( a54688a  and  a54675a );
 a1690a <=( a54664a  and  a54651a );
 a1691a <=( a54640a  and  a54627a );
 a1692a <=( a54616a  and  a54603a );
 a1693a <=( a54592a  and  a54579a );
 a1694a <=( a54568a  and  a54555a );
 a1695a <=( a54544a  and  a54531a );
 a1696a <=( a54520a  and  a54507a );
 a1697a <=( a54496a  and  a54483a );
 a1698a <=( a54472a  and  a54459a );
 a1699a <=( a54448a  and  a54435a );
 a1700a <=( a54424a  and  a54411a );
 a1701a <=( a54400a  and  a54387a );
 a1702a <=( a54376a  and  a54363a );
 a1703a <=( a54352a  and  a54339a );
 a1704a <=( a54328a  and  a54315a );
 a1705a <=( a54304a  and  a54291a );
 a1706a <=( a54280a  and  a54267a );
 a1707a <=( a54256a  and  a54243a );
 a1708a <=( a54232a  and  a54219a );
 a1709a <=( a54208a  and  a54195a );
 a1710a <=( a54184a  and  a54171a );
 a1711a <=( a54160a  and  a54147a );
 a1712a <=( a54136a  and  a54123a );
 a1713a <=( a54112a  and  a54099a );
 a1714a <=( a54088a  and  a54075a );
 a1715a <=( a54064a  and  a54051a );
 a1716a <=( a54040a  and  a54027a );
 a1717a <=( a54016a  and  a54003a );
 a1718a <=( a53992a  and  a53979a );
 a1719a <=( a53968a  and  a53955a );
 a1720a <=( a53944a  and  a53931a );
 a1721a <=( a53920a  and  a53907a );
 a1722a <=( a53896a  and  a53883a );
 a1723a <=( a53872a  and  a53859a );
 a1724a <=( a53848a  and  a53835a );
 a1725a <=( a53824a  and  a53811a );
 a1726a <=( a53800a  and  a53787a );
 a1727a <=( a53776a  and  a53763a );
 a1728a <=( a53752a  and  a53739a );
 a1729a <=( a53728a  and  a53715a );
 a1730a <=( a53704a  and  a53691a );
 a1731a <=( a53680a  and  a53667a );
 a1732a <=( a53656a  and  a53643a );
 a1733a <=( a53632a  and  a53619a );
 a1734a <=( a53608a  and  a53595a );
 a1735a <=( a53584a  and  a53571a );
 a1736a <=( a53560a  and  a53547a );
 a1737a <=( a53536a  and  a53523a );
 a1738a <=( a53512a  and  a53499a );
 a1739a <=( a53488a  and  a53475a );
 a1740a <=( a53464a  and  a53451a );
 a1741a <=( a53440a  and  a53427a );
 a1742a <=( a53416a  and  a53403a );
 a1743a <=( a53392a  and  a53379a );
 a1744a <=( a53368a  and  a53355a );
 a1745a <=( a53344a  and  a53331a );
 a1746a <=( a53320a  and  a53307a );
 a1747a <=( a53296a  and  a53283a );
 a1748a <=( a53272a  and  a53259a );
 a1749a <=( a53248a  and  a53235a );
 a1750a <=( a53224a  and  a53211a );
 a1751a <=( a53200a  and  a53187a );
 a1752a <=( a53176a  and  a53163a );
 a1753a <=( a53152a  and  a53139a );
 a1754a <=( a53128a  and  a53115a );
 a1755a <=( a53104a  and  a53091a );
 a1756a <=( a53080a  and  a53067a );
 a1757a <=( a53056a  and  a53043a );
 a1758a <=( a53032a  and  a53019a );
 a1759a <=( a53008a  and  a52995a );
 a1760a <=( a52984a  and  a52971a );
 a1761a <=( a52960a  and  a52947a );
 a1762a <=( a52936a  and  a52923a );
 a1763a <=( a52912a  and  a52899a );
 a1764a <=( a52888a  and  a52875a );
 a1765a <=( a52864a  and  a52851a );
 a1766a <=( a52840a  and  a52827a );
 a1767a <=( a52816a  and  a52803a );
 a1768a <=( a52792a  and  a52779a );
 a1769a <=( a52768a  and  a52755a );
 a1770a <=( a52744a  and  a52731a );
 a1771a <=( a52720a  and  a52707a );
 a1772a <=( a52696a  and  a52683a );
 a1773a <=( a52672a  and  a52659a );
 a1774a <=( a52648a  and  a52635a );
 a1775a <=( a52624a  and  a52611a );
 a1776a <=( a52600a  and  a52587a );
 a1777a <=( a52576a  and  a52563a );
 a1778a <=( a52552a  and  a52539a );
 a1779a <=( a52528a  and  a52515a );
 a1780a <=( a52504a  and  a52491a );
 a1781a <=( a52480a  and  a52467a );
 a1782a <=( a52456a  and  a52443a );
 a1783a <=( a52432a  and  a52419a );
 a1784a <=( a52408a  and  a52395a );
 a1785a <=( a52384a  and  a52371a );
 a1786a <=( a52360a  and  a52347a );
 a1787a <=( a52336a  and  a52323a );
 a1788a <=( a52312a  and  a52299a );
 a1789a <=( a52288a  and  a52275a );
 a1790a <=( a52264a  and  a52251a );
 a1791a <=( a52240a  and  a52227a );
 a1792a <=( a52216a  and  a52203a );
 a1793a <=( a52192a  and  a52179a );
 a1794a <=( a52168a  and  a52155a );
 a1795a <=( a52144a  and  a52131a );
 a1796a <=( a52120a  and  a52107a );
 a1797a <=( a52096a  and  a52083a );
 a1798a <=( a52072a  and  a52059a );
 a1799a <=( a52048a  and  a52035a );
 a1800a <=( a52024a  and  a52011a );
 a1801a <=( a52000a  and  a51987a );
 a1802a <=( a51976a  and  a51963a );
 a1803a <=( a51952a  and  a51939a );
 a1804a <=( a51928a  and  a51915a );
 a1805a <=( a51904a  and  a51891a );
 a1806a <=( a51880a  and  a51867a );
 a1807a <=( a51856a  and  a51843a );
 a1808a <=( a51832a  and  a51819a );
 a1809a <=( a51808a  and  a51795a );
 a1810a <=( a51784a  and  a51771a );
 a1811a <=( a51760a  and  a51747a );
 a1812a <=( a51736a  and  a51723a );
 a1813a <=( a51712a  and  a51699a );
 a1814a <=( a51688a  and  a51675a );
 a1815a <=( a51664a  and  a51651a );
 a1816a <=( a51640a  and  a51627a );
 a1817a <=( a51616a  and  a51603a );
 a1818a <=( a51592a  and  a51579a );
 a1819a <=( a51568a  and  a51555a );
 a1820a <=( a51544a  and  a51531a );
 a1821a <=( a51520a  and  a51507a );
 a1822a <=( a51496a  and  a51483a );
 a1823a <=( a51472a  and  a51459a );
 a1824a <=( a51448a  and  a51435a );
 a1825a <=( a51424a  and  a51411a );
 a1826a <=( a51400a  and  a51387a );
 a1827a <=( a51376a  and  a51363a );
 a1828a <=( a51352a  and  a51339a );
 a1829a <=( a51328a  and  a51315a );
 a1830a <=( a51304a  and  a51291a );
 a1831a <=( a51280a  and  a51267a );
 a1832a <=( a51256a  and  a51243a );
 a1833a <=( a51232a  and  a51219a );
 a1834a <=( a51208a  and  a51195a );
 a1835a <=( a51184a  and  a51171a );
 a1836a <=( a51160a  and  a51147a );
 a1837a <=( a51136a  and  a51123a );
 a1838a <=( a51112a  and  a51099a );
 a1839a <=( a51088a  and  a51075a );
 a1840a <=( a51064a  and  a51051a );
 a1841a <=( a51040a  and  a51027a );
 a1842a <=( a51016a  and  a51003a );
 a1843a <=( a50992a  and  a50979a );
 a1844a <=( a50968a  and  a50955a );
 a1845a <=( a50944a  and  a50931a );
 a1846a <=( a50920a  and  a50907a );
 a1847a <=( a50896a  and  a50883a );
 a1848a <=( a50872a  and  a50859a );
 a1849a <=( a50848a  and  a50835a );
 a1850a <=( a50824a  and  a50811a );
 a1851a <=( a50800a  and  a50787a );
 a1852a <=( a50776a  and  a50763a );
 a1853a <=( a50752a  and  a50739a );
 a1854a <=( a50728a  and  a50715a );
 a1855a <=( a50704a  and  a50691a );
 a1856a <=( a50680a  and  a50667a );
 a1857a <=( a50656a  and  a50643a );
 a1858a <=( a50632a  and  a50619a );
 a1859a <=( a50608a  and  a50595a );
 a1860a <=( a50584a  and  a50571a );
 a1861a <=( a50560a  and  a50547a );
 a1862a <=( a50536a  and  a50523a );
 a1863a <=( a50512a  and  a50499a );
 a1864a <=( a50488a  and  a50475a );
 a1865a <=( a50464a  and  a50451a );
 a1866a <=( a50440a  and  a50427a );
 a1867a <=( a50416a  and  a50403a );
 a1868a <=( a50392a  and  a50379a );
 a1869a <=( a50368a  and  a50355a );
 a1870a <=( a50344a  and  a50331a );
 a1871a <=( a50320a  and  a50307a );
 a1872a <=( a50296a  and  a50283a );
 a1873a <=( a50272a  and  a50259a );
 a1874a <=( a50248a  and  a50235a );
 a1875a <=( a50224a  and  a50211a );
 a1876a <=( a50200a  and  a50187a );
 a1877a <=( a50176a  and  a50163a );
 a1878a <=( a50152a  and  a50139a );
 a1879a <=( a50128a  and  a50115a );
 a1880a <=( a50104a  and  a50091a );
 a1881a <=( a50080a  and  a50067a );
 a1882a <=( a50056a  and  a50043a );
 a1883a <=( a50032a  and  a50019a );
 a1884a <=( a50008a  and  a49995a );
 a1885a <=( a49984a  and  a49971a );
 a1886a <=( a49960a  and  a49947a );
 a1887a <=( a49936a  and  a49923a );
 a1888a <=( a49912a  and  a49899a );
 a1889a <=( a49888a  and  a49875a );
 a1890a <=( a49864a  and  a49851a );
 a1891a <=( a49840a  and  a49827a );
 a1892a <=( a49816a  and  a49803a );
 a1893a <=( a49792a  and  a49779a );
 a1894a <=( a49768a  and  a49755a );
 a1895a <=( a49744a  and  a49731a );
 a1896a <=( a49720a  and  a49707a );
 a1897a <=( a49696a  and  a49683a );
 a1898a <=( a49672a  and  a49659a );
 a1899a <=( a49648a  and  a49635a );
 a1900a <=( a49624a  and  a49611a );
 a1901a <=( a49600a  and  a49587a );
 a1902a <=( a49576a  and  a49563a );
 a1903a <=( a49552a  and  a49539a );
 a1904a <=( a49528a  and  a49515a );
 a1905a <=( a49504a  and  a49491a );
 a1906a <=( a49480a  and  a49467a );
 a1907a <=( a49456a  and  a49443a );
 a1908a <=( a49432a  and  a49419a );
 a1909a <=( a49408a  and  a49395a );
 a1910a <=( a49384a  and  a49371a );
 a1911a <=( a49360a  and  a49347a );
 a1912a <=( a49336a  and  a49323a );
 a1913a <=( a49312a  and  a49299a );
 a1914a <=( a49288a  and  a49275a );
 a1915a <=( a49264a  and  a49251a );
 a1916a <=( a49240a  and  a49227a );
 a1917a <=( a49216a  and  a49203a );
 a1918a <=( a49192a  and  a49179a );
 a1919a <=( a49168a  and  a49155a );
 a1920a <=( a49144a  and  a49131a );
 a1921a <=( a49120a  and  a49107a );
 a1922a <=( a49096a  and  a49083a );
 a1923a <=( a49072a  and  a49059a );
 a1924a <=( a49048a  and  a49035a );
 a1925a <=( a49024a  and  a49011a );
 a1926a <=( a49000a  and  a48987a );
 a1927a <=( a48976a  and  a48963a );
 a1928a <=( a48952a  and  a48939a );
 a1929a <=( a48928a  and  a48915a );
 a1930a <=( a48904a  and  a48891a );
 a1931a <=( a48880a  and  a48867a );
 a1932a <=( a48856a  and  a48843a );
 a1933a <=( a48832a  and  a48819a );
 a1934a <=( a48808a  and  a48795a );
 a1935a <=( a48784a  and  a48771a );
 a1936a <=( a48760a  and  a48747a );
 a1937a <=( a48736a  and  a48723a );
 a1938a <=( a48712a  and  a48699a );
 a1939a <=( a48688a  and  a48675a );
 a1940a <=( a48664a  and  a48651a );
 a1941a <=( a48640a  and  a48627a );
 a1942a <=( a48616a  and  a48603a );
 a1943a <=( a48592a  and  a48579a );
 a1944a <=( a48568a  and  a48555a );
 a1945a <=( a48544a  and  a48531a );
 a1946a <=( a48520a  and  a48507a );
 a1947a <=( a48496a  and  a48483a );
 a1948a <=( a48472a  and  a48459a );
 a1949a <=( a48448a  and  a48435a );
 a1950a <=( a48424a  and  a48411a );
 a1951a <=( a48400a  and  a48387a );
 a1952a <=( a48376a  and  a48363a );
 a1953a <=( a48352a  and  a48339a );
 a1954a <=( a48328a  and  a48315a );
 a1955a <=( a48304a  and  a48291a );
 a1956a <=( a48280a  and  a48267a );
 a1957a <=( a48256a  and  a48243a );
 a1958a <=( a48232a  and  a48219a );
 a1959a <=( a48208a  and  a48195a );
 a1960a <=( a48184a  and  a48171a );
 a1961a <=( a48160a  and  a48147a );
 a1962a <=( a48136a  and  a48123a );
 a1963a <=( a48112a  and  a48099a );
 a1964a <=( a48088a  and  a48075a );
 a1965a <=( a48064a  and  a48051a );
 a1966a <=( a48040a  and  a48027a );
 a1967a <=( a48016a  and  a48003a );
 a1968a <=( a47992a  and  a47979a );
 a1969a <=( a47968a  and  a47955a );
 a1970a <=( a47944a  and  a47931a );
 a1971a <=( a47920a  and  a47907a );
 a1972a <=( a47896a  and  a47883a );
 a1973a <=( a47872a  and  a47859a );
 a1974a <=( a47848a  and  a47835a );
 a1975a <=( a47824a  and  a47811a );
 a1976a <=( a47800a  and  a47787a );
 a1977a <=( a47776a  and  a47763a );
 a1978a <=( a47752a  and  a47739a );
 a1979a <=( a47728a  and  a47715a );
 a1980a <=( a47704a  and  a47691a );
 a1981a <=( a47680a  and  a47667a );
 a1982a <=( a47656a  and  a47643a );
 a1983a <=( a47632a  and  a47619a );
 a1984a <=( a47608a  and  a47595a );
 a1985a <=( a47584a  and  a47571a );
 a1986a <=( a47560a  and  a47547a );
 a1987a <=( a47536a  and  a47523a );
 a1988a <=( a47512a  and  a47499a );
 a1989a <=( a47488a  and  a47475a );
 a1990a <=( a47464a  and  a47451a );
 a1991a <=( a47440a  and  a47427a );
 a1992a <=( a47416a  and  a47403a );
 a1993a <=( a47392a  and  a47379a );
 a1994a <=( a47368a  and  a47355a );
 a1995a <=( a47344a  and  a47331a );
 a1996a <=( a47320a  and  a47307a );
 a1997a <=( a47296a  and  a47283a );
 a1998a <=( a47272a  and  a47259a );
 a1999a <=( a47248a  and  a47235a );
 a2000a <=( a47224a  and  a47211a );
 a2001a <=( a47200a  and  a47187a );
 a2002a <=( a47176a  and  a47163a );
 a2003a <=( a47152a  and  a47139a );
 a2004a <=( a47128a  and  a47115a );
 a2005a <=( a47104a  and  a47091a );
 a2006a <=( a47080a  and  a47067a );
 a2007a <=( a47056a  and  a47043a );
 a2008a <=( a47032a  and  a47019a );
 a2009a <=( a47008a  and  a46995a );
 a2010a <=( a46984a  and  a46971a );
 a2011a <=( a46960a  and  a46947a );
 a2012a <=( a46936a  and  a46923a );
 a2013a <=( a46912a  and  a46899a );
 a2014a <=( a46888a  and  a46875a );
 a2015a <=( a46864a  and  a46851a );
 a2016a <=( a46840a  and  a46827a );
 a2017a <=( a46816a  and  a46803a );
 a2018a <=( a46792a  and  a46779a );
 a2019a <=( a46768a  and  a46755a );
 a2020a <=( a46744a  and  a46731a );
 a2021a <=( a46720a  and  a46707a );
 a2022a <=( a46696a  and  a46683a );
 a2023a <=( a46672a  and  a46659a );
 a2024a <=( a46648a  and  a46635a );
 a2025a <=( a46624a  and  a46611a );
 a2026a <=( a46600a  and  a46587a );
 a2027a <=( a46576a  and  a46563a );
 a2028a <=( a46552a  and  a46539a );
 a2029a <=( a46528a  and  a46515a );
 a2030a <=( a46504a  and  a46491a );
 a2031a <=( a46480a  and  a46467a );
 a2032a <=( a46456a  and  a46443a );
 a2033a <=( a46432a  and  a46419a );
 a2034a <=( a46408a  and  a46395a );
 a2035a <=( a46384a  and  a46371a );
 a2036a <=( a46360a  and  a46347a );
 a2037a <=( a46336a  and  a46323a );
 a2038a <=( a46312a  and  a46299a );
 a2039a <=( a46288a  and  a46275a );
 a2040a <=( a46264a  and  a46251a );
 a2041a <=( a46240a  and  a46227a );
 a2042a <=( a46216a  and  a46203a );
 a2043a <=( a46192a  and  a46179a );
 a2044a <=( a46168a  and  a46155a );
 a2045a <=( a46144a  and  a46131a );
 a2046a <=( a46120a  and  a46107a );
 a2047a <=( a46096a  and  a46083a );
 a2048a <=( a46072a  and  a46059a );
 a2049a <=( a46048a  and  a46035a );
 a2050a <=( a46024a  and  a46011a );
 a2051a <=( a46000a  and  a45987a );
 a2052a <=( a45976a  and  a45963a );
 a2053a <=( a45952a  and  a45939a );
 a2054a <=( a45928a  and  a45915a );
 a2055a <=( a45904a  and  a45891a );
 a2056a <=( a45880a  and  a45867a );
 a2057a <=( a45856a  and  a45843a );
 a2058a <=( a45832a  and  a45819a );
 a2059a <=( a45808a  and  a45795a );
 a2060a <=( a45784a  and  a45771a );
 a2061a <=( a45760a  and  a45747a );
 a2062a <=( a45736a  and  a45723a );
 a2063a <=( a45712a  and  a45699a );
 a2064a <=( a45688a  and  a45675a );
 a2065a <=( a45664a  and  a45651a );
 a2066a <=( a45640a  and  a45627a );
 a2067a <=( a45616a  and  a45603a );
 a2068a <=( a45592a  and  a45579a );
 a2069a <=( a45568a  and  a45555a );
 a2070a <=( a45544a  and  a45531a );
 a2071a <=( a45520a  and  a45507a );
 a2072a <=( a45496a  and  a45483a );
 a2073a <=( a45472a  and  a45459a );
 a2074a <=( a45448a  and  a45435a );
 a2075a <=( a45424a  and  a45411a );
 a2076a <=( a45400a  and  a45387a );
 a2077a <=( a45376a  and  a45363a );
 a2078a <=( a45352a  and  a45339a );
 a2079a <=( a45328a  and  a45315a );
 a2080a <=( a45304a  and  a45291a );
 a2081a <=( a45280a  and  a45267a );
 a2082a <=( a45256a  and  a45243a );
 a2083a <=( a45232a  and  a45219a );
 a2084a <=( a45208a  and  a45195a );
 a2085a <=( a45184a  and  a45171a );
 a2086a <=( a45160a  and  a45147a );
 a2087a <=( a45136a  and  a45123a );
 a2088a <=( a45112a  and  a45099a );
 a2089a <=( a45088a  and  a45075a );
 a2090a <=( a45064a  and  a45051a );
 a2091a <=( a45040a  and  a45027a );
 a2092a <=( a45016a  and  a45003a );
 a2093a <=( a44992a  and  a44979a );
 a2094a <=( a44968a  and  a44955a );
 a2095a <=( a44944a  and  a44931a );
 a2096a <=( a44920a  and  a44907a );
 a2097a <=( a44896a  and  a44883a );
 a2098a <=( a44872a  and  a44859a );
 a2099a <=( a44848a  and  a44835a );
 a2100a <=( a44824a  and  a44811a );
 a2101a <=( a44800a  and  a44787a );
 a2102a <=( a44776a  and  a44763a );
 a2103a <=( a44752a  and  a44739a );
 a2104a <=( a44728a  and  a44715a );
 a2105a <=( a44704a  and  a44691a );
 a2106a <=( a44680a  and  a44667a );
 a2107a <=( a44656a  and  a44643a );
 a2108a <=( a44632a  and  a44619a );
 a2109a <=( a44608a  and  a44595a );
 a2110a <=( a44584a  and  a44571a );
 a2111a <=( a44560a  and  a44547a );
 a2112a <=( a44536a  and  a44523a );
 a2113a <=( a44512a  and  a44499a );
 a2114a <=( a44488a  and  a44475a );
 a2115a <=( a44464a  and  a44451a );
 a2116a <=( a44440a  and  a44427a );
 a2117a <=( a44416a  and  a44403a );
 a2118a <=( a44392a  and  a44379a );
 a2119a <=( a44368a  and  a44355a );
 a2120a <=( a44344a  and  a44331a );
 a2121a <=( a44320a  and  a44307a );
 a2122a <=( a44296a  and  a44283a );
 a2123a <=( a44272a  and  a44259a );
 a2124a <=( a44248a  and  a44235a );
 a2125a <=( a44224a  and  a44211a );
 a2126a <=( a44200a  and  a44187a );
 a2127a <=( a44176a  and  a44163a );
 a2128a <=( a44152a  and  a44139a );
 a2129a <=( a44128a  and  a44115a );
 a2130a <=( a44104a  and  a44091a );
 a2131a <=( a44080a  and  a44067a );
 a2132a <=( a44056a  and  a44043a );
 a2133a <=( a44032a  and  a44019a );
 a2134a <=( a44008a  and  a43995a );
 a2135a <=( a43984a  and  a43971a );
 a2136a <=( a43960a  and  a43947a );
 a2137a <=( a43936a  and  a43923a );
 a2138a <=( a43912a  and  a43899a );
 a2139a <=( a43888a  and  a43875a );
 a2140a <=( a43864a  and  a43851a );
 a2141a <=( a43840a  and  a43827a );
 a2142a <=( a43816a  and  a43803a );
 a2143a <=( a43792a  and  a43779a );
 a2144a <=( a43768a  and  a43755a );
 a2145a <=( a43744a  and  a43731a );
 a2146a <=( a43720a  and  a43707a );
 a2147a <=( a43696a  and  a43683a );
 a2148a <=( a43672a  and  a43659a );
 a2149a <=( a43648a  and  a43635a );
 a2150a <=( a43624a  and  a43611a );
 a2151a <=( a43600a  and  a43587a );
 a2152a <=( a43576a  and  a43563a );
 a2153a <=( a43552a  and  a43539a );
 a2154a <=( a43528a  and  a43515a );
 a2155a <=( a43504a  and  a43491a );
 a2156a <=( a43480a  and  a43467a );
 a2157a <=( a43456a  and  a43443a );
 a2158a <=( a43432a  and  a43419a );
 a2159a <=( a43408a  and  a43395a );
 a2160a <=( a43384a  and  a43371a );
 a2161a <=( a43360a  and  a43347a );
 a2162a <=( a43336a  and  a43323a );
 a2163a <=( a43312a  and  a43299a );
 a2164a <=( a43288a  and  a43275a );
 a2165a <=( a43264a  and  a43251a );
 a2166a <=( a43240a  and  a43227a );
 a2167a <=( a43216a  and  a43203a );
 a2168a <=( a43192a  and  a43179a );
 a2169a <=( a43168a  and  a43155a );
 a2170a <=( a43144a  and  a43131a );
 a2171a <=( a43120a  and  a43107a );
 a2172a <=( a43096a  and  a43083a );
 a2173a <=( a43072a  and  a43059a );
 a2174a <=( a43048a  and  a43035a );
 a2175a <=( a43024a  and  a43011a );
 a2176a <=( a43000a  and  a42987a );
 a2177a <=( a42976a  and  a42963a );
 a2178a <=( a42952a  and  a42939a );
 a2179a <=( a42928a  and  a42915a );
 a2180a <=( a42904a  and  a42891a );
 a2181a <=( a42880a  and  a42867a );
 a2182a <=( a42856a  and  a42843a );
 a2183a <=( a42832a  and  a42819a );
 a2184a <=( a42808a  and  a42795a );
 a2185a <=( a42784a  and  a42771a );
 a2186a <=( a42760a  and  a42747a );
 a2187a <=( a42736a  and  a42723a );
 a2188a <=( a42712a  and  a42699a );
 a2189a <=( a42688a  and  a42675a );
 a2190a <=( a42664a  and  a42651a );
 a2191a <=( a42640a  and  a42627a );
 a2192a <=( a42616a  and  a42603a );
 a2193a <=( a42592a  and  a42579a );
 a2194a <=( a42568a  and  a42555a );
 a2195a <=( a42544a  and  a42531a );
 a2196a <=( a42520a  and  a42507a );
 a2197a <=( a42496a  and  a42483a );
 a2198a <=( a42472a  and  a42459a );
 a2199a <=( a42448a  and  a42435a );
 a2200a <=( a42424a  and  a42411a );
 a2201a <=( a42400a  and  a42387a );
 a2202a <=( a42376a  and  a42363a );
 a2203a <=( a42352a  and  a42339a );
 a2204a <=( a42328a  and  a42315a );
 a2205a <=( a42304a  and  a42291a );
 a2206a <=( a42280a  and  a42267a );
 a2207a <=( a42256a  and  a42243a );
 a2208a <=( a42232a  and  a42219a );
 a2209a <=( a42208a  and  a42195a );
 a2210a <=( a42184a  and  a42171a );
 a2211a <=( a42160a  and  a42147a );
 a2212a <=( a42136a  and  a42123a );
 a2213a <=( a42112a  and  a42099a );
 a2214a <=( a42088a  and  a42075a );
 a2215a <=( a42064a  and  a42051a );
 a2216a <=( a42040a  and  a42027a );
 a2217a <=( a42016a  and  a42003a );
 a2218a <=( a41992a  and  a41979a );
 a2219a <=( a41968a  and  a41955a );
 a2220a <=( a41944a  and  a41931a );
 a2221a <=( a41920a  and  a41907a );
 a2222a <=( a41896a  and  a41883a );
 a2223a <=( a41872a  and  a41859a );
 a2224a <=( a41848a  and  a41835a );
 a2225a <=( a41824a  and  a41811a );
 a2226a <=( a41800a  and  a41787a );
 a2227a <=( a41776a  and  a41763a );
 a2228a <=( a41752a  and  a41739a );
 a2229a <=( a41728a  and  a41715a );
 a2230a <=( a41704a  and  a41691a );
 a2231a <=( a41680a  and  a41667a );
 a2232a <=( a41656a  and  a41643a );
 a2233a <=( a41632a  and  a41619a );
 a2234a <=( a41608a  and  a41595a );
 a2235a <=( a41584a  and  a41571a );
 a2236a <=( a41560a  and  a41547a );
 a2237a <=( a41536a  and  a41523a );
 a2238a <=( a41512a  and  a41499a );
 a2239a <=( a41488a  and  a41475a );
 a2240a <=( a41464a  and  a41451a );
 a2241a <=( a41440a  and  a41427a );
 a2242a <=( a41416a  and  a41403a );
 a2243a <=( a41392a  and  a41379a );
 a2244a <=( a41368a  and  a41355a );
 a2245a <=( a41344a  and  a41331a );
 a2246a <=( a41320a  and  a41307a );
 a2247a <=( a41296a  and  a41283a );
 a2248a <=( a41272a  and  a41259a );
 a2249a <=( a41248a  and  a41235a );
 a2250a <=( a41224a  and  a41211a );
 a2251a <=( a41200a  and  a41187a );
 a2252a <=( a41176a  and  a41163a );
 a2253a <=( a41152a  and  a41139a );
 a2254a <=( a41128a  and  a41115a );
 a2255a <=( a41104a  and  a41091a );
 a2256a <=( a41080a  and  a41067a );
 a2257a <=( a41056a  and  a41043a );
 a2258a <=( a41032a  and  a41019a );
 a2259a <=( a41008a  and  a40995a );
 a2260a <=( a40984a  and  a40971a );
 a2261a <=( a40960a  and  a40947a );
 a2262a <=( a40936a  and  a40923a );
 a2263a <=( a40912a  and  a40899a );
 a2264a <=( a40888a  and  a40875a );
 a2265a <=( a40864a  and  a40851a );
 a2266a <=( a40840a  and  a40827a );
 a2267a <=( a40816a  and  a40803a );
 a2268a <=( a40792a  and  a40779a );
 a2269a <=( a40768a  and  a40755a );
 a2270a <=( a40744a  and  a40731a );
 a2271a <=( a40720a  and  a40707a );
 a2272a <=( a40696a  and  a40683a );
 a2273a <=( a40672a  and  a40659a );
 a2274a <=( a40648a  and  a40635a );
 a2275a <=( a40624a  and  a40611a );
 a2276a <=( a40600a  and  a40587a );
 a2277a <=( a40576a  and  a40563a );
 a2278a <=( a40552a  and  a40539a );
 a2279a <=( a40528a  and  a40515a );
 a2280a <=( a40504a  and  a40491a );
 a2281a <=( a40480a  and  a40467a );
 a2282a <=( a40456a  and  a40443a );
 a2283a <=( a40432a  and  a40419a );
 a2284a <=( a40408a  and  a40395a );
 a2285a <=( a40384a  and  a40371a );
 a2286a <=( a40360a  and  a40347a );
 a2287a <=( a40336a  and  a40323a );
 a2288a <=( a40312a  and  a40299a );
 a2289a <=( a40288a  and  a40275a );
 a2290a <=( a40264a  and  a40251a );
 a2291a <=( a40240a  and  a40227a );
 a2292a <=( a40216a  and  a40203a );
 a2293a <=( a40192a  and  a40179a );
 a2294a <=( a40168a  and  a40155a );
 a2295a <=( a40144a  and  a40131a );
 a2296a <=( a40120a  and  a40107a );
 a2297a <=( a40096a  and  a40083a );
 a2298a <=( a40072a  and  a40059a );
 a2299a <=( a40048a  and  a40035a );
 a2300a <=( a40024a  and  a40011a );
 a2301a <=( a40000a  and  a39987a );
 a2302a <=( a39976a  and  a39963a );
 a2303a <=( a39952a  and  a39939a );
 a2304a <=( a39928a  and  a39915a );
 a2305a <=( a39904a  and  a39891a );
 a2306a <=( a39880a  and  a39867a );
 a2307a <=( a39856a  and  a39843a );
 a2308a <=( a39832a  and  a39819a );
 a2309a <=( a39808a  and  a39795a );
 a2310a <=( a39784a  and  a39771a );
 a2311a <=( a39760a  and  a39747a );
 a2312a <=( a39736a  and  a39723a );
 a2313a <=( a39712a  and  a39699a );
 a2314a <=( a39688a  and  a39675a );
 a2315a <=( a39664a  and  a39651a );
 a2316a <=( a39640a  and  a39627a );
 a2317a <=( a39616a  and  a39603a );
 a2318a <=( a39592a  and  a39579a );
 a2319a <=( a39568a  and  a39555a );
 a2320a <=( a39544a  and  a39531a );
 a2321a <=( a39520a  and  a39507a );
 a2322a <=( a39496a  and  a39483a );
 a2323a <=( a39472a  and  a39459a );
 a2324a <=( a39448a  and  a39435a );
 a2325a <=( a39424a  and  a39411a );
 a2326a <=( a39400a  and  a39387a );
 a2327a <=( a39376a  and  a39363a );
 a2328a <=( a39352a  and  a39339a );
 a2329a <=( a39328a  and  a39315a );
 a2330a <=( a39304a  and  a39291a );
 a2331a <=( a39280a  and  a39267a );
 a2332a <=( a39256a  and  a39243a );
 a2333a <=( a39232a  and  a39219a );
 a2334a <=( a39208a  and  a39195a );
 a2335a <=( a39184a  and  a39171a );
 a2336a <=( a39160a  and  a39147a );
 a2337a <=( a39136a  and  a39123a );
 a2338a <=( a39112a  and  a39099a );
 a2339a <=( a39088a  and  a39075a );
 a2340a <=( a39064a  and  a39051a );
 a2341a <=( a39040a  and  a39027a );
 a2342a <=( a39016a  and  a39003a );
 a2343a <=( a38992a  and  a38979a );
 a2344a <=( a38968a  and  a38955a );
 a2345a <=( a38944a  and  a38931a );
 a2346a <=( a38920a  and  a38907a );
 a2347a <=( a38896a  and  a38883a );
 a2348a <=( a38872a  and  a38859a );
 a2349a <=( a38848a  and  a38835a );
 a2350a <=( a38824a  and  a38811a );
 a2351a <=( a38800a  and  a38787a );
 a2352a <=( a38776a  and  a38763a );
 a2353a <=( a38752a  and  a38739a );
 a2354a <=( a38728a  and  a38715a );
 a2355a <=( a38704a  and  a38691a );
 a2356a <=( a38680a  and  a38667a );
 a2357a <=( a38656a  and  a38643a );
 a2358a <=( a38632a  and  a38619a );
 a2359a <=( a38608a  and  a38595a );
 a2360a <=( a38584a  and  a38571a );
 a2361a <=( a38560a  and  a38547a );
 a2362a <=( a38536a  and  a38523a );
 a2363a <=( a38512a  and  a38499a );
 a2364a <=( a38488a  and  a38475a );
 a2365a <=( a38464a  and  a38451a );
 a2366a <=( a38440a  and  a38427a );
 a2367a <=( a38416a  and  a38403a );
 a2368a <=( a38392a  and  a38379a );
 a2369a <=( a38368a  and  a38355a );
 a2370a <=( a38344a  and  a38331a );
 a2371a <=( a38320a  and  a38307a );
 a2372a <=( a38296a  and  a38283a );
 a2373a <=( a38272a  and  a38259a );
 a2374a <=( a38248a  and  a38235a );
 a2375a <=( a38224a  and  a38211a );
 a2376a <=( a38200a  and  a38187a );
 a2377a <=( a38176a  and  a38163a );
 a2378a <=( a38152a  and  a38139a );
 a2379a <=( a38128a  and  a38115a );
 a2380a <=( a38104a  and  a38091a );
 a2381a <=( a38080a  and  a38067a );
 a2382a <=( a38056a  and  a38043a );
 a2383a <=( a38032a  and  a38019a );
 a2384a <=( a38008a  and  a37995a );
 a2385a <=( a37984a  and  a37971a );
 a2386a <=( a37960a  and  a37947a );
 a2387a <=( a37936a  and  a37923a );
 a2388a <=( a37912a  and  a37899a );
 a2389a <=( a37888a  and  a37875a );
 a2390a <=( a37864a  and  a37851a );
 a2391a <=( a37840a  and  a37827a );
 a2392a <=( a37816a  and  a37803a );
 a2393a <=( a37792a  and  a37779a );
 a2394a <=( a37768a  and  a37755a );
 a2395a <=( a37744a  and  a37731a );
 a2396a <=( a37720a  and  a37707a );
 a2397a <=( a37696a  and  a37683a );
 a2398a <=( a37672a  and  a37659a );
 a2399a <=( a37648a  and  a37637a );
 a2400a <=( a37626a  and  a37615a );
 a2401a <=( a37604a  and  a37593a );
 a2402a <=( a37582a  and  a37571a );
 a2403a <=( a37560a  and  a37549a );
 a2404a <=( a37538a  and  a37527a );
 a2405a <=( a37516a  and  a37505a );
 a2406a <=( a37494a  and  a37483a );
 a2407a <=( a37472a  and  a37461a );
 a2408a <=( a37450a  and  a37439a );
 a2409a <=( a37428a  and  a37417a );
 a2410a <=( a37406a  and  a37395a );
 a2411a <=( a37384a  and  a37373a );
 a2412a <=( a37362a  and  a37351a );
 a2413a <=( a37340a  and  a37329a );
 a2414a <=( a37318a  and  a37307a );
 a2415a <=( a37296a  and  a37285a );
 a2416a <=( a37274a  and  a37263a );
 a2417a <=( a37252a  and  a37241a );
 a2418a <=( a37230a  and  a37219a );
 a2419a <=( a37208a  and  a37197a );
 a2420a <=( a37186a  and  a37175a );
 a2421a <=( a37164a  and  a37153a );
 a2422a <=( a37142a  and  a37131a );
 a2423a <=( a37120a  and  a37109a );
 a2424a <=( a37098a  and  a37087a );
 a2425a <=( a37076a  and  a37065a );
 a2426a <=( a37054a  and  a37043a );
 a2427a <=( a37032a  and  a37021a );
 a2428a <=( a37010a  and  a36999a );
 a2429a <=( a36988a  and  a36977a );
 a2430a <=( a36966a  and  a36955a );
 a2431a <=( a36944a  and  a36933a );
 a2432a <=( a36922a  and  a36911a );
 a2433a <=( a36900a  and  a36889a );
 a2434a <=( a36878a  and  a36867a );
 a2435a <=( a36856a  and  a36845a );
 a2436a <=( a36834a  and  a36823a );
 a2437a <=( a36812a  and  a36801a );
 a2438a <=( a36790a  and  a36779a );
 a2439a <=( a36768a  and  a36757a );
 a2440a <=( a36746a  and  a36735a );
 a2441a <=( a36724a  and  a36713a );
 a2442a <=( a36702a  and  a36691a );
 a2443a <=( a36680a  and  a36669a );
 a2444a <=( a36658a  and  a36647a );
 a2445a <=( a36636a  and  a36625a );
 a2446a <=( a36614a  and  a36603a );
 a2447a <=( a36592a  and  a36581a );
 a2448a <=( a36570a  and  a36559a );
 a2449a <=( a36548a  and  a36537a );
 a2450a <=( a36526a  and  a36515a );
 a2451a <=( a36504a  and  a36493a );
 a2452a <=( a36482a  and  a36471a );
 a2453a <=( a36460a  and  a36449a );
 a2454a <=( a36438a  and  a36427a );
 a2455a <=( a36416a  and  a36405a );
 a2456a <=( a36394a  and  a36383a );
 a2457a <=( a36372a  and  a36361a );
 a2458a <=( a36350a  and  a36339a );
 a2459a <=( a36328a  and  a36317a );
 a2460a <=( a36306a  and  a36295a );
 a2461a <=( a36284a  and  a36273a );
 a2462a <=( a36262a  and  a36251a );
 a2463a <=( a36240a  and  a36229a );
 a2464a <=( a36218a  and  a36207a );
 a2465a <=( a36196a  and  a36185a );
 a2466a <=( a36174a  and  a36163a );
 a2467a <=( a36152a  and  a36141a );
 a2468a <=( a36130a  and  a36119a );
 a2469a <=( a36108a  and  a36097a );
 a2470a <=( a36086a  and  a36075a );
 a2471a <=( a36064a  and  a36053a );
 a2472a <=( a36042a  and  a36031a );
 a2473a <=( a36020a  and  a36009a );
 a2474a <=( a35998a  and  a35987a );
 a2475a <=( a35976a  and  a35965a );
 a2476a <=( a35954a  and  a35943a );
 a2477a <=( a35932a  and  a35921a );
 a2478a <=( a35910a  and  a35899a );
 a2479a <=( a35888a  and  a35877a );
 a2480a <=( a35866a  and  a35855a );
 a2481a <=( a35844a  and  a35833a );
 a2482a <=( a35822a  and  a35811a );
 a2483a <=( a35800a  and  a35789a );
 a2484a <=( a35778a  and  a35767a );
 a2485a <=( a35756a  and  a35745a );
 a2486a <=( a35734a  and  a35723a );
 a2487a <=( a35712a  and  a35701a );
 a2488a <=( a35690a  and  a35679a );
 a2489a <=( a35668a  and  a35657a );
 a2490a <=( a35646a  and  a35635a );
 a2491a <=( a35624a  and  a35613a );
 a2492a <=( a35602a  and  a35591a );
 a2493a <=( a35580a  and  a35569a );
 a2494a <=( a35558a  and  a35547a );
 a2495a <=( a35536a  and  a35525a );
 a2496a <=( a35514a  and  a35503a );
 a2497a <=( a35492a  and  a35481a );
 a2498a <=( a35470a  and  a35459a );
 a2499a <=( a35448a  and  a35437a );
 a2500a <=( a35426a  and  a35415a );
 a2501a <=( a35404a  and  a35393a );
 a2502a <=( a35382a  and  a35371a );
 a2503a <=( a35360a  and  a35349a );
 a2504a <=( a35338a  and  a35327a );
 a2505a <=( a35316a  and  a35305a );
 a2506a <=( a35294a  and  a35283a );
 a2507a <=( a35272a  and  a35261a );
 a2508a <=( a35250a  and  a35239a );
 a2509a <=( a35228a  and  a35217a );
 a2510a <=( a35206a  and  a35195a );
 a2511a <=( a35184a  and  a35173a );
 a2512a <=( a35162a  and  a35151a );
 a2513a <=( a35140a  and  a35129a );
 a2514a <=( a35118a  and  a35107a );
 a2515a <=( a35096a  and  a35085a );
 a2516a <=( a35074a  and  a35063a );
 a2517a <=( a35052a  and  a35041a );
 a2518a <=( a35030a  and  a35019a );
 a2519a <=( a35008a  and  a34997a );
 a2520a <=( a34986a  and  a34975a );
 a2521a <=( a34964a  and  a34953a );
 a2522a <=( a34942a  and  a34931a );
 a2523a <=( a34920a  and  a34909a );
 a2524a <=( a34898a  and  a34887a );
 a2525a <=( a34876a  and  a34865a );
 a2526a <=( a34854a  and  a34843a );
 a2527a <=( a34832a  and  a34821a );
 a2528a <=( a34810a  and  a34799a );
 a2529a <=( a34788a  and  a34777a );
 a2530a <=( a34766a  and  a34755a );
 a2531a <=( a34744a  and  a34733a );
 a2532a <=( a34722a  and  a34711a );
 a2533a <=( a34700a  and  a34689a );
 a2534a <=( a34678a  and  a34667a );
 a2535a <=( a34656a  and  a34645a );
 a2536a <=( a34634a  and  a34623a );
 a2537a <=( a34612a  and  a34601a );
 a2538a <=( a34590a  and  a34579a );
 a2539a <=( a34568a  and  a34557a );
 a2540a <=( a34546a  and  a34535a );
 a2541a <=( a34524a  and  a34513a );
 a2542a <=( a34502a  and  a34491a );
 a2543a <=( a34480a  and  a34469a );
 a2544a <=( a34458a  and  a34447a );
 a2545a <=( a34436a  and  a34425a );
 a2546a <=( a34414a  and  a34403a );
 a2547a <=( a34392a  and  a34381a );
 a2548a <=( a34370a  and  a34359a );
 a2549a <=( a34348a  and  a34337a );
 a2550a <=( a34326a  and  a34315a );
 a2551a <=( a34304a  and  a34293a );
 a2552a <=( a34282a  and  a34271a );
 a2553a <=( a34260a  and  a34249a );
 a2554a <=( a34238a  and  a34227a );
 a2555a <=( a34216a  and  a34205a );
 a2556a <=( a34194a  and  a34183a );
 a2557a <=( a34172a  and  a34161a );
 a2558a <=( a34150a  and  a34139a );
 a2559a <=( a34128a  and  a34117a );
 a2560a <=( a34106a  and  a34095a );
 a2561a <=( a34084a  and  a34073a );
 a2562a <=( a34062a  and  a34051a );
 a2563a <=( a34040a  and  a34029a );
 a2564a <=( a34018a  and  a34007a );
 a2565a <=( a33996a  and  a33985a );
 a2566a <=( a33974a  and  a33963a );
 a2567a <=( a33952a  and  a33941a );
 a2568a <=( a33930a  and  a33919a );
 a2569a <=( a33908a  and  a33897a );
 a2570a <=( a33886a  and  a33875a );
 a2571a <=( a33864a  and  a33853a );
 a2572a <=( a33842a  and  a33831a );
 a2573a <=( a33820a  and  a33809a );
 a2574a <=( a33798a  and  a33787a );
 a2575a <=( a33776a  and  a33765a );
 a2576a <=( a33754a  and  a33743a );
 a2577a <=( a33732a  and  a33721a );
 a2578a <=( a33710a  and  a33699a );
 a2579a <=( a33688a  and  a33677a );
 a2580a <=( a33666a  and  a33655a );
 a2581a <=( a33644a  and  a33633a );
 a2582a <=( a33622a  and  a33611a );
 a2583a <=( a33600a  and  a33589a );
 a2584a <=( a33578a  and  a33567a );
 a2585a <=( a33556a  and  a33545a );
 a2586a <=( a33534a  and  a33523a );
 a2587a <=( a33512a  and  a33501a );
 a2588a <=( a33490a  and  a33479a );
 a2589a <=( a33468a  and  a33457a );
 a2590a <=( a33446a  and  a33435a );
 a2591a <=( a33424a  and  a33413a );
 a2592a <=( a33402a  and  a33391a );
 a2593a <=( a33380a  and  a33369a );
 a2594a <=( a33358a  and  a33347a );
 a2595a <=( a33336a  and  a33325a );
 a2596a <=( a33314a  and  a33303a );
 a2597a <=( a33292a  and  a33281a );
 a2598a <=( a33270a  and  a33259a );
 a2599a <=( a33248a  and  a33237a );
 a2600a <=( a33226a  and  a33215a );
 a2601a <=( a33204a  and  a33193a );
 a2602a <=( a33182a  and  a33171a );
 a2603a <=( a33160a  and  a33149a );
 a2604a <=( a33138a  and  a33127a );
 a2605a <=( a33116a  and  a33105a );
 a2606a <=( a33094a  and  a33083a );
 a2607a <=( a33072a  and  a33061a );
 a2608a <=( a33050a  and  a33039a );
 a2609a <=( a33028a  and  a33017a );
 a2610a <=( a33006a  and  a32995a );
 a2611a <=( a32984a  and  a32973a );
 a2612a <=( a32962a  and  a32951a );
 a2613a <=( a32940a  and  a32929a );
 a2614a <=( a32918a  and  a32907a );
 a2615a <=( a32896a  and  a32885a );
 a2616a <=( a32874a  and  a32863a );
 a2617a <=( a32852a  and  a32841a );
 a2618a <=( a32830a  and  a32819a );
 a2619a <=( a32808a  and  a32797a );
 a2620a <=( a32786a  and  a32775a );
 a2621a <=( a32764a  and  a32753a );
 a2622a <=( a32742a  and  a32731a );
 a2623a <=( a32720a  and  a32709a );
 a2624a <=( a32698a  and  a32687a );
 a2625a <=( a32676a  and  a32665a );
 a2626a <=( a32654a  and  a32643a );
 a2627a <=( a32632a  and  a32621a );
 a2628a <=( a32610a  and  a32599a );
 a2629a <=( a32588a  and  a32577a );
 a2630a <=( a32566a  and  a32555a );
 a2631a <=( a32544a  and  a32533a );
 a2632a <=( a32522a  and  a32511a );
 a2633a <=( a32500a  and  a32489a );
 a2634a <=( a32478a  and  a32467a );
 a2635a <=( a32456a  and  a32445a );
 a2636a <=( a32434a  and  a32423a );
 a2637a <=( a32412a  and  a32401a );
 a2638a <=( a32390a  and  a32379a );
 a2639a <=( a32368a  and  a32357a );
 a2640a <=( a32346a  and  a32335a );
 a2641a <=( a32324a  and  a32313a );
 a2642a <=( a32302a  and  a32291a );
 a2643a <=( a32280a  and  a32269a );
 a2644a <=( a32258a  and  a32247a );
 a2645a <=( a32236a  and  a32225a );
 a2646a <=( a32214a  and  a32203a );
 a2647a <=( a32192a  and  a32181a );
 a2648a <=( a32170a  and  a32159a );
 a2649a <=( a32148a  and  a32137a );
 a2650a <=( a32126a  and  a32115a );
 a2651a <=( a32104a  and  a32093a );
 a2652a <=( a32082a  and  a32071a );
 a2653a <=( a32060a  and  a32049a );
 a2654a <=( a32038a  and  a32027a );
 a2655a <=( a32016a  and  a32005a );
 a2656a <=( a31994a  and  a31983a );
 a2657a <=( a31972a  and  a31961a );
 a2658a <=( a31950a  and  a31939a );
 a2659a <=( a31928a  and  a31917a );
 a2660a <=( a31906a  and  a31895a );
 a2661a <=( a31884a  and  a31873a );
 a2662a <=( a31862a  and  a31851a );
 a2663a <=( a31840a  and  a31829a );
 a2664a <=( a31818a  and  a31807a );
 a2665a <=( a31796a  and  a31785a );
 a2666a <=( a31774a  and  a31763a );
 a2667a <=( a31752a  and  a31741a );
 a2668a <=( a31730a  and  a31719a );
 a2669a <=( a31708a  and  a31697a );
 a2670a <=( a31686a  and  a31675a );
 a2671a <=( a31664a  and  a31653a );
 a2672a <=( a31642a  and  a31631a );
 a2673a <=( a31620a  and  a31609a );
 a2674a <=( a31598a  and  a31587a );
 a2675a <=( a31576a  and  a31565a );
 a2676a <=( a31554a  and  a31543a );
 a2677a <=( a31532a  and  a31521a );
 a2678a <=( a31510a  and  a31499a );
 a2679a <=( a31488a  and  a31477a );
 a2680a <=( a31466a  and  a31455a );
 a2681a <=( a31444a  and  a31433a );
 a2682a <=( a31422a  and  a31411a );
 a2683a <=( a31400a  and  a31389a );
 a2684a <=( a31378a  and  a31367a );
 a2685a <=( a31356a  and  a31345a );
 a2686a <=( a31334a  and  a31323a );
 a2687a <=( a31312a  and  a31301a );
 a2688a <=( a31290a  and  a31279a );
 a2689a <=( a31268a  and  a31257a );
 a2690a <=( a31246a  and  a31235a );
 a2691a <=( a31224a  and  a31213a );
 a2692a <=( a31202a  and  a31191a );
 a2693a <=( a31180a  and  a31169a );
 a2694a <=( a31158a  and  a31147a );
 a2695a <=( a31136a  and  a31125a );
 a2696a <=( a31114a  and  a31103a );
 a2697a <=( a31092a  and  a31081a );
 a2698a <=( a31070a  and  a31059a );
 a2699a <=( a31048a  and  a31037a );
 a2700a <=( a31026a  and  a31015a );
 a2701a <=( a31004a  and  a30993a );
 a2702a <=( a30982a  and  a30971a );
 a2703a <=( a30960a  and  a30949a );
 a2704a <=( a30938a  and  a30927a );
 a2705a <=( a30916a  and  a30905a );
 a2706a <=( a30894a  and  a30883a );
 a2707a <=( a30872a  and  a30861a );
 a2708a <=( a30850a  and  a30839a );
 a2709a <=( a30828a  and  a30817a );
 a2710a <=( a30806a  and  a30795a );
 a2711a <=( a30784a  and  a30773a );
 a2712a <=( a30762a  and  a30751a );
 a2713a <=( a30740a  and  a30729a );
 a2714a <=( a30718a  and  a30707a );
 a2715a <=( a30696a  and  a30685a );
 a2716a <=( a30674a  and  a30663a );
 a2717a <=( a30652a  and  a30641a );
 a2718a <=( a30630a  and  a30619a );
 a2719a <=( a30608a  and  a30597a );
 a2720a <=( a30586a  and  a30575a );
 a2721a <=( a30564a  and  a30553a );
 a2722a <=( a30542a  and  a30531a );
 a2723a <=( a30520a  and  a30509a );
 a2724a <=( a30498a  and  a30487a );
 a2725a <=( a30476a  and  a30465a );
 a2726a <=( a30454a  and  a30443a );
 a2727a <=( a30432a  and  a30421a );
 a2728a <=( a30410a  and  a30399a );
 a2729a <=( a30388a  and  a30377a );
 a2730a <=( a30366a  and  a30355a );
 a2731a <=( a30344a  and  a30333a );
 a2732a <=( a30322a  and  a30311a );
 a2733a <=( a30300a  and  a30289a );
 a2734a <=( a30278a  and  a30267a );
 a2735a <=( a30256a  and  a30245a );
 a2736a <=( a30234a  and  a30223a );
 a2737a <=( a30212a  and  a30201a );
 a2738a <=( a30190a  and  a30179a );
 a2739a <=( a30168a  and  a30157a );
 a2740a <=( a30146a  and  a30135a );
 a2741a <=( a30124a  and  a30113a );
 a2742a <=( a30102a  and  a30091a );
 a2743a <=( a30080a  and  a30069a );
 a2744a <=( a30058a  and  a30047a );
 a2745a <=( a30036a  and  a30025a );
 a2746a <=( a30014a  and  a30003a );
 a2747a <=( a29992a  and  a29981a );
 a2748a <=( a29970a  and  a29959a );
 a2749a <=( a29948a  and  a29937a );
 a2750a <=( a29926a  and  a29915a );
 a2751a <=( a29904a  and  a29893a );
 a2752a <=( a29882a  and  a29871a );
 a2753a <=( a29860a  and  a29849a );
 a2754a <=( a29838a  and  a29827a );
 a2755a <=( a29816a  and  a29805a );
 a2756a <=( a29794a  and  a29783a );
 a2757a <=( a29772a  and  a29761a );
 a2758a <=( a29750a  and  a29739a );
 a2759a <=( a29728a  and  a29717a );
 a2760a <=( a29706a  and  a29695a );
 a2761a <=( a29684a  and  a29673a );
 a2762a <=( a29662a  and  a29651a );
 a2763a <=( a29640a  and  a29629a );
 a2764a <=( a29618a  and  a29607a );
 a2765a <=( a29596a  and  a29585a );
 a2766a <=( a29574a  and  a29563a );
 a2767a <=( a29552a  and  a29541a );
 a2768a <=( a29530a  and  a29519a );
 a2769a <=( a29508a  and  a29497a );
 a2770a <=( a29486a  and  a29475a );
 a2771a <=( a29464a  and  a29453a );
 a2772a <=( a29442a  and  a29431a );
 a2773a <=( a29420a  and  a29409a );
 a2774a <=( a29398a  and  a29387a );
 a2775a <=( a29376a  and  a29365a );
 a2776a <=( a29354a  and  a29343a );
 a2777a <=( a29332a  and  a29321a );
 a2778a <=( a29310a  and  a29299a );
 a2779a <=( a29288a  and  a29277a );
 a2780a <=( a29266a  and  a29255a );
 a2781a <=( a29244a  and  a29233a );
 a2782a <=( a29222a  and  a29211a );
 a2783a <=( a29200a  and  a29189a );
 a2784a <=( a29178a  and  a29167a );
 a2785a <=( a29156a  and  a29145a );
 a2786a <=( a29134a  and  a29123a );
 a2787a <=( a29112a  and  a29101a );
 a2788a <=( a29090a  and  a29079a );
 a2789a <=( a29068a  and  a29057a );
 a2790a <=( a29046a  and  a29035a );
 a2791a <=( a29024a  and  a29013a );
 a2792a <=( a29002a  and  a28991a );
 a2793a <=( a28980a  and  a28969a );
 a2794a <=( a28958a  and  a28947a );
 a2795a <=( a28936a  and  a28925a );
 a2796a <=( a28914a  and  a28903a );
 a2797a <=( a28892a  and  a28881a );
 a2798a <=( a28870a  and  a28859a );
 a2799a <=( a28848a  and  a28837a );
 a2800a <=( a28826a  and  a28815a );
 a2801a <=( a28804a  and  a28793a );
 a2802a <=( a28782a  and  a28771a );
 a2803a <=( a28760a  and  a28749a );
 a2804a <=( a28738a  and  a28727a );
 a2805a <=( a28716a  and  a28705a );
 a2806a <=( a28694a  and  a28683a );
 a2807a <=( a28672a  and  a28661a );
 a2808a <=( a28650a  and  a28639a );
 a2809a <=( a28628a  and  a28617a );
 a2810a <=( a28606a  and  a28595a );
 a2811a <=( a28584a  and  a28573a );
 a2812a <=( a28562a  and  a28551a );
 a2813a <=( a28540a  and  a28529a );
 a2814a <=( a28518a  and  a28507a );
 a2815a <=( a28496a  and  a28485a );
 a2816a <=( a28474a  and  a28463a );
 a2817a <=( a28452a  and  a28441a );
 a2818a <=( a28430a  and  a28419a );
 a2819a <=( a28408a  and  a28397a );
 a2820a <=( a28386a  and  a28375a );
 a2821a <=( a28364a  and  a28353a );
 a2822a <=( a28342a  and  a28331a );
 a2823a <=( a28320a  and  a28309a );
 a2824a <=( a28298a  and  a28287a );
 a2825a <=( a28276a  and  a28265a );
 a2826a <=( a28254a  and  a28243a );
 a2827a <=( a28232a  and  a28221a );
 a2828a <=( a28210a  and  a28199a );
 a2829a <=( a28188a  and  a28177a );
 a2830a <=( a28166a  and  a28155a );
 a2831a <=( a28144a  and  a28133a );
 a2832a <=( a28122a  and  a28111a );
 a2833a <=( a28100a  and  a28089a );
 a2834a <=( a28078a  and  a28067a );
 a2835a <=( a28056a  and  a28045a );
 a2836a <=( a28034a  and  a28023a );
 a2837a <=( a28012a  and  a28001a );
 a2838a <=( a27990a  and  a27979a );
 a2839a <=( a27968a  and  a27957a );
 a2840a <=( a27946a  and  a27935a );
 a2841a <=( a27924a  and  a27913a );
 a2842a <=( a27902a  and  a27891a );
 a2843a <=( a27880a  and  a27869a );
 a2844a <=( a27858a  and  a27847a );
 a2845a <=( a27836a  and  a27825a );
 a2846a <=( a27814a  and  a27803a );
 a2847a <=( a27792a  and  a27781a );
 a2848a <=( a27770a  and  a27759a );
 a2849a <=( a27748a  and  a27737a );
 a2850a <=( a27726a  and  a27715a );
 a2851a <=( a27704a  and  a27693a );
 a2852a <=( a27682a  and  a27671a );
 a2853a <=( a27660a  and  a27649a );
 a2854a <=( a27638a  and  a27627a );
 a2855a <=( a27616a  and  a27605a );
 a2856a <=( a27594a  and  a27583a );
 a2857a <=( a27572a  and  a27561a );
 a2858a <=( a27550a  and  a27539a );
 a2859a <=( a27528a  and  a27517a );
 a2860a <=( a27506a  and  a27495a );
 a2861a <=( a27484a  and  a27473a );
 a2862a <=( a27462a  and  a27451a );
 a2863a <=( a27440a  and  a27429a );
 a2864a <=( a27418a  and  a27407a );
 a2865a <=( a27396a  and  a27385a );
 a2866a <=( a27374a  and  a27363a );
 a2867a <=( a27352a  and  a27341a );
 a2868a <=( a27330a  and  a27319a );
 a2869a <=( a27308a  and  a27297a );
 a2870a <=( a27286a  and  a27275a );
 a2871a <=( a27264a  and  a27253a );
 a2872a <=( a27242a  and  a27231a );
 a2873a <=( a27220a  and  a27209a );
 a2874a <=( a27198a  and  a27187a );
 a2875a <=( a27176a  and  a27165a );
 a2876a <=( a27154a  and  a27143a );
 a2877a <=( a27132a  and  a27121a );
 a2878a <=( a27110a  and  a27099a );
 a2879a <=( a27088a  and  a27077a );
 a2880a <=( a27066a  and  a27055a );
 a2881a <=( a27044a  and  a27033a );
 a2882a <=( a27022a  and  a27011a );
 a2883a <=( a27000a  and  a26989a );
 a2884a <=( a26978a  and  a26967a );
 a2885a <=( a26956a  and  a26945a );
 a2886a <=( a26934a  and  a26923a );
 a2887a <=( a26912a  and  a26901a );
 a2888a <=( a26890a  and  a26879a );
 a2889a <=( a26868a  and  a26857a );
 a2890a <=( a26846a  and  a26835a );
 a2891a <=( a26824a  and  a26813a );
 a2892a <=( a26802a  and  a26791a );
 a2893a <=( a26780a  and  a26769a );
 a2894a <=( a26758a  and  a26747a );
 a2895a <=( a26736a  and  a26725a );
 a2896a <=( a26714a  and  a26703a );
 a2897a <=( a26692a  and  a26681a );
 a2898a <=( a26670a  and  a26659a );
 a2899a <=( a26648a  and  a26637a );
 a2900a <=( a26626a  and  a26615a );
 a2901a <=( a26604a  and  a26593a );
 a2902a <=( a26582a  and  a26571a );
 a2903a <=( a26560a  and  a26549a );
 a2904a <=( a26538a  and  a26527a );
 a2905a <=( a26516a  and  a26505a );
 a2906a <=( a26494a  and  a26483a );
 a2907a <=( a26472a  and  a26461a );
 a2908a <=( a26450a  and  a26439a );
 a2909a <=( a26428a  and  a26417a );
 a2910a <=( a26406a  and  a26395a );
 a2911a <=( a26384a  and  a26373a );
 a2912a <=( a26362a  and  a26351a );
 a2913a <=( a26340a  and  a26329a );
 a2914a <=( a26318a  and  a26307a );
 a2915a <=( a26296a  and  a26285a );
 a2916a <=( a26274a  and  a26263a );
 a2917a <=( a26252a  and  a26241a );
 a2918a <=( a26230a  and  a26219a );
 a2919a <=( a26208a  and  a26197a );
 a2920a <=( a26186a  and  a26175a );
 a2921a <=( a26164a  and  a26153a );
 a2922a <=( a26142a  and  a26131a );
 a2923a <=( a26120a  and  a26109a );
 a2924a <=( a26098a  and  a26087a );
 a2925a <=( a26076a  and  a26065a );
 a2926a <=( a26054a  and  a26043a );
 a2927a <=( a26032a  and  a26021a );
 a2928a <=( a26010a  and  a25999a );
 a2929a <=( a25988a  and  a25977a );
 a2930a <=( a25966a  and  a25955a );
 a2931a <=( a25944a  and  a25933a );
 a2932a <=( a25922a  and  a25911a );
 a2933a <=( a25900a  and  a25889a );
 a2934a <=( a25878a  and  a25867a );
 a2935a <=( a25856a  and  a25845a );
 a2936a <=( a25834a  and  a25823a );
 a2937a <=( a25812a  and  a25801a );
 a2938a <=( a25790a  and  a25779a );
 a2939a <=( a25768a  and  a25757a );
 a2940a <=( a25746a  and  a25735a );
 a2941a <=( a25724a  and  a25713a );
 a2942a <=( a25702a  and  a25691a );
 a2943a <=( a25680a  and  a25669a );
 a2944a <=( a25658a  and  a25647a );
 a2945a <=( a25636a  and  a25625a );
 a2946a <=( a25614a  and  a25603a );
 a2947a <=( a25592a  and  a25581a );
 a2948a <=( a25570a  and  a25559a );
 a2949a <=( a25548a  and  a25537a );
 a2950a <=( a25526a  and  a25515a );
 a2951a <=( a25504a  and  a25493a );
 a2952a <=( a25482a  and  a25471a );
 a2953a <=( a25460a  and  a25449a );
 a2954a <=( a25438a  and  a25427a );
 a2955a <=( a25416a  and  a25405a );
 a2956a <=( a25394a  and  a25383a );
 a2957a <=( a25372a  and  a25361a );
 a2958a <=( a25350a  and  a25339a );
 a2959a <=( a25328a  and  a25317a );
 a2960a <=( a25306a  and  a25295a );
 a2961a <=( a25284a  and  a25273a );
 a2962a <=( a25262a  and  a25251a );
 a2963a <=( a25240a  and  a25229a );
 a2964a <=( a25218a  and  a25207a );
 a2965a <=( a25196a  and  a25185a );
 a2966a <=( a25174a  and  a25163a );
 a2967a <=( a25152a  and  a25141a );
 a2968a <=( a25130a  and  a25119a );
 a2969a <=( a25108a  and  a25097a );
 a2970a <=( a25086a  and  a25075a );
 a2971a <=( a25064a  and  a25053a );
 a2972a <=( a25042a  and  a25031a );
 a2973a <=( a25020a  and  a25009a );
 a2974a <=( a24998a  and  a24987a );
 a2975a <=( a24976a  and  a24965a );
 a2976a <=( a24954a  and  a24943a );
 a2977a <=( a24932a  and  a24921a );
 a2978a <=( a24910a  and  a24899a );
 a2979a <=( a24888a  and  a24877a );
 a2980a <=( a24866a  and  a24855a );
 a2981a <=( a24844a  and  a24833a );
 a2982a <=( a24822a  and  a24811a );
 a2983a <=( a24800a  and  a24789a );
 a2984a <=( a24778a  and  a24767a );
 a2985a <=( a24756a  and  a24745a );
 a2986a <=( a24734a  and  a24723a );
 a2987a <=( a24712a  and  a24701a );
 a2988a <=( a24690a  and  a24679a );
 a2989a <=( a24668a  and  a24657a );
 a2990a <=( a24646a  and  a24635a );
 a2991a <=( a24624a  and  a24613a );
 a2992a <=( a24602a  and  a24591a );
 a2993a <=( a24580a  and  a24569a );
 a2994a <=( a24558a  and  a24547a );
 a2995a <=( a24536a  and  a24525a );
 a2996a <=( a24514a  and  a24503a );
 a2997a <=( a24492a  and  a24481a );
 a2998a <=( a24470a  and  a24459a );
 a2999a <=( a24448a  and  a24437a );
 a3000a <=( a24426a  and  a24415a );
 a3001a <=( a24404a  and  a24393a );
 a3002a <=( a24382a  and  a24371a );
 a3003a <=( a24360a  and  a24349a );
 a3004a <=( a24338a  and  a24327a );
 a3005a <=( a24316a  and  a24305a );
 a3006a <=( a24294a  and  a24283a );
 a3007a <=( a24272a  and  a24261a );
 a3008a <=( a24250a  and  a24239a );
 a3009a <=( a24228a  and  a24217a );
 a3010a <=( a24206a  and  a24195a );
 a3011a <=( a24184a  and  a24173a );
 a3012a <=( a24162a  and  a24151a );
 a3013a <=( a24140a  and  a24129a );
 a3014a <=( a24118a  and  a24107a );
 a3015a <=( a24096a  and  a24085a );
 a3016a <=( a24074a  and  a24063a );
 a3017a <=( a24052a  and  a24041a );
 a3018a <=( a24030a  and  a24019a );
 a3019a <=( a24008a  and  a23997a );
 a3020a <=( a23986a  and  a23975a );
 a3021a <=( a23964a  and  a23953a );
 a3022a <=( a23942a  and  a23931a );
 a3023a <=( a23920a  and  a23909a );
 a3024a <=( a23898a  and  a23887a );
 a3025a <=( a23876a  and  a23865a );
 a3026a <=( a23854a  and  a23843a );
 a3027a <=( a23832a  and  a23821a );
 a3028a <=( a23810a  and  a23799a );
 a3029a <=( a23788a  and  a23777a );
 a3030a <=( a23766a  and  a23755a );
 a3031a <=( a23744a  and  a23733a );
 a3032a <=( a23722a  and  a23711a );
 a3033a <=( a23700a  and  a23689a );
 a3034a <=( a23678a  and  a23667a );
 a3035a <=( a23656a  and  a23645a );
 a3036a <=( a23634a  and  a23623a );
 a3037a <=( a23612a  and  a23601a );
 a3038a <=( a23590a  and  a23579a );
 a3039a <=( a23568a  and  a23557a );
 a3040a <=( a23546a  and  a23535a );
 a3041a <=( a23524a  and  a23513a );
 a3042a <=( a23502a  and  a23491a );
 a3043a <=( a23480a  and  a23469a );
 a3044a <=( a23458a  and  a23447a );
 a3045a <=( a23436a  and  a23425a );
 a3046a <=( a23414a  and  a23403a );
 a3047a <=( a23392a  and  a23381a );
 a3048a <=( a23370a  and  a23359a );
 a3049a <=( a23348a  and  a23337a );
 a3050a <=( a23326a  and  a23315a );
 a3051a <=( a23304a  and  a23293a );
 a3052a <=( a23282a  and  a23271a );
 a3053a <=( a23260a  and  a23249a );
 a3054a <=( a23238a  and  a23227a );
 a3055a <=( a23216a  and  a23205a );
 a3056a <=( a23196a  and  a23185a );
 a3057a <=( a23176a  and  a23165a );
 a3058a <=( a23156a  and  a23145a );
 a3059a <=( a23136a  and  a23125a );
 a3060a <=( a23116a  and  a23105a );
 a3061a <=( a23096a  and  a23085a );
 a3062a <=( a23076a  and  a23065a );
 a3063a <=( a23056a  and  a23045a );
 a3064a <=( a23036a  and  a23025a );
 a3065a <=( a23016a  and  a23005a );
 a3066a <=( a22996a  and  a22985a );
 a3067a <=( a22976a  and  a22965a );
 a3068a <=( a22956a  and  a22945a );
 a3069a <=( a22936a  and  a22925a );
 a3070a <=( a22916a  and  a22905a );
 a3071a <=( a22896a  and  a22885a );
 a3072a <=( a22876a  and  a22865a );
 a3073a <=( a22856a  and  a22845a );
 a3074a <=( a22836a  and  a22825a );
 a3075a <=( a22816a  and  a22805a );
 a3076a <=( a22796a  and  a22785a );
 a3077a <=( a22776a  and  a22765a );
 a3078a <=( a22756a  and  a22745a );
 a3079a <=( a22736a  and  a22725a );
 a3080a <=( a22716a  and  a22705a );
 a3081a <=( a22696a  and  a22685a );
 a3082a <=( a22676a  and  a22665a );
 a3083a <=( a22656a  and  a22645a );
 a3084a <=( a22636a  and  a22625a );
 a3085a <=( a22616a  and  a22605a );
 a3086a <=( a22596a  and  a22585a );
 a3087a <=( a22576a  and  a22565a );
 a3088a <=( a22556a  and  a22545a );
 a3089a <=( a22536a  and  a22525a );
 a3090a <=( a22516a  and  a22505a );
 a3091a <=( a22496a  and  a22485a );
 a3092a <=( a22476a  and  a22465a );
 a3093a <=( a22456a  and  a22445a );
 a3094a <=( a22436a  and  a22425a );
 a3095a <=( a22416a  and  a22405a );
 a3096a <=( a22396a  and  a22385a );
 a3097a <=( a22376a  and  a22365a );
 a3098a <=( a22356a  and  a22345a );
 a3099a <=( a22336a  and  a22325a );
 a3100a <=( a22316a  and  a22305a );
 a3101a <=( a22296a  and  a22285a );
 a3102a <=( a22276a  and  a22265a );
 a3103a <=( a22256a  and  a22245a );
 a3104a <=( a22236a  and  a22225a );
 a3105a <=( a22216a  and  a22205a );
 a3106a <=( a22196a  and  a22185a );
 a3107a <=( a22176a  and  a22165a );
 a3108a <=( a22156a  and  a22145a );
 a3109a <=( a22136a  and  a22125a );
 a3110a <=( a22116a  and  a22105a );
 a3111a <=( a22096a  and  a22085a );
 a3112a <=( a22076a  and  a22065a );
 a3113a <=( a22056a  and  a22045a );
 a3114a <=( a22036a  and  a22025a );
 a3115a <=( a22016a  and  a22005a );
 a3116a <=( a21996a  and  a21985a );
 a3117a <=( a21976a  and  a21965a );
 a3118a <=( a21956a  and  a21945a );
 a3119a <=( a21936a  and  a21925a );
 a3120a <=( a21916a  and  a21905a );
 a3121a <=( a21896a  and  a21885a );
 a3122a <=( a21876a  and  a21865a );
 a3123a <=( a21856a  and  a21845a );
 a3124a <=( a21836a  and  a21825a );
 a3125a <=( a21816a  and  a21805a );
 a3126a <=( a21796a  and  a21785a );
 a3127a <=( a21776a  and  a21765a );
 a3128a <=( a21756a  and  a21745a );
 a3129a <=( a21736a  and  a21725a );
 a3130a <=( a21716a  and  a21705a );
 a3131a <=( a21696a  and  a21685a );
 a3132a <=( a21676a  and  a21665a );
 a3133a <=( a21656a  and  a21645a );
 a3134a <=( a21636a  and  a21625a );
 a3135a <=( a21616a  and  a21605a );
 a3136a <=( a21596a  and  a21585a );
 a3137a <=( a21576a  and  a21565a );
 a3138a <=( a21556a  and  a21545a );
 a3139a <=( a21536a  and  a21525a );
 a3140a <=( a21516a  and  a21505a );
 a3141a <=( a21496a  and  a21485a );
 a3142a <=( a21476a  and  a21465a );
 a3143a <=( a21456a  and  a21445a );
 a3144a <=( a21436a  and  a21425a );
 a3145a <=( a21416a  and  a21405a );
 a3146a <=( a21396a  and  a21385a );
 a3147a <=( a21376a  and  a21365a );
 a3148a <=( a21356a  and  a21345a );
 a3149a <=( a21336a  and  a21325a );
 a3150a <=( a21316a  and  a21305a );
 a3151a <=( a21296a  and  a21285a );
 a3152a <=( a21276a  and  a21265a );
 a3153a <=( a21256a  and  a21245a );
 a3154a <=( a21236a  and  a21225a );
 a3155a <=( a21216a  and  a21205a );
 a3156a <=( a21196a  and  a21185a );
 a3157a <=( a21176a  and  a21165a );
 a3158a <=( a21156a  and  a21145a );
 a3159a <=( a21136a  and  a21125a );
 a3160a <=( a21116a  and  a21105a );
 a3161a <=( a21096a  and  a21085a );
 a3162a <=( a21076a  and  a21065a );
 a3163a <=( a21056a  and  a21045a );
 a3164a <=( a21036a  and  a21025a );
 a3165a <=( a21016a  and  a21005a );
 a3166a <=( a20996a  and  a20985a );
 a3167a <=( a20976a  and  a20965a );
 a3168a <=( a20956a  and  a20945a );
 a3169a <=( a20936a  and  a20925a );
 a3170a <=( a20916a  and  a20905a );
 a3171a <=( a20896a  and  a20885a );
 a3172a <=( a20876a  and  a20865a );
 a3173a <=( a20856a  and  a20845a );
 a3174a <=( a20836a  and  a20825a );
 a3175a <=( a20816a  and  a20805a );
 a3176a <=( a20796a  and  a20785a );
 a3177a <=( a20776a  and  a20765a );
 a3178a <=( a20756a  and  a20745a );
 a3179a <=( a20736a  and  a20725a );
 a3180a <=( a20716a  and  a20705a );
 a3181a <=( a20696a  and  a20685a );
 a3182a <=( a20676a  and  a20665a );
 a3183a <=( a20656a  and  a20645a );
 a3184a <=( a20636a  and  a20625a );
 a3185a <=( a20616a  and  a20605a );
 a3186a <=( a20596a  and  a20585a );
 a3187a <=( a20576a  and  a20565a );
 a3188a <=( a20556a  and  a20545a );
 a3189a <=( a20536a  and  a20525a );
 a3190a <=( a20516a  and  a20505a );
 a3191a <=( a20496a  and  a20485a );
 a3192a <=( a20476a  and  a20465a );
 a3193a <=( a20456a  and  a20445a );
 a3194a <=( a20436a  and  a20425a );
 a3195a <=( a20416a  and  a20405a );
 a3196a <=( a20396a  and  a20385a );
 a3197a <=( a20376a  and  a20365a );
 a3198a <=( a20356a  and  a20345a );
 a3199a <=( a20336a  and  a20325a );
 a3200a <=( a20316a  and  a20305a );
 a3201a <=( a20296a  and  a20285a );
 a3202a <=( a20276a  and  a20265a );
 a3203a <=( a20256a  and  a20245a );
 a3204a <=( a20236a  and  a20225a );
 a3205a <=( a20216a  and  a20205a );
 a3206a <=( a20196a  and  a20185a );
 a3207a <=( a20176a  and  a20165a );
 a3208a <=( a20156a  and  a20145a );
 a3209a <=( a20136a  and  a20125a );
 a3210a <=( a20116a  and  a20105a );
 a3211a <=( a20096a  and  a20085a );
 a3212a <=( a20076a  and  a20065a );
 a3213a <=( a20056a  and  a20045a );
 a3214a <=( a20036a  and  a20025a );
 a3215a <=( a20016a  and  a20005a );
 a3216a <=( a19996a  and  a19985a );
 a3217a <=( a19976a  and  a19965a );
 a3218a <=( a19956a  and  a19945a );
 a3219a <=( a19936a  and  a19925a );
 a3220a <=( a19916a  and  a19905a );
 a3221a <=( a19896a  and  a19885a );
 a3222a <=( a19876a  and  a19865a );
 a3223a <=( a19856a  and  a19845a );
 a3224a <=( a19836a  and  a19825a );
 a3225a <=( a19816a  and  a19805a );
 a3226a <=( a19796a  and  a19785a );
 a3227a <=( a19776a  and  a19765a );
 a3228a <=( a19756a  and  a19745a );
 a3229a <=( a19736a  and  a19725a );
 a3230a <=( a19716a  and  a19705a );
 a3231a <=( a19696a  and  a19685a );
 a3232a <=( a19676a  and  a19665a );
 a3233a <=( a19656a  and  a19645a );
 a3234a <=( a19636a  and  a19625a );
 a3235a <=( a19616a  and  a19605a );
 a3236a <=( a19596a  and  a19585a );
 a3237a <=( a19576a  and  a19565a );
 a3238a <=( a19556a  and  a19545a );
 a3239a <=( a19536a  and  a19525a );
 a3240a <=( a19516a  and  a19505a );
 a3241a <=( a19496a  and  a19485a );
 a3242a <=( a19476a  and  a19465a );
 a3243a <=( a19456a  and  a19445a );
 a3244a <=( a19436a  and  a19425a );
 a3245a <=( a19416a  and  a19405a );
 a3246a <=( a19396a  and  a19385a );
 a3247a <=( a19376a  and  a19365a );
 a3248a <=( a19356a  and  a19345a );
 a3249a <=( a19336a  and  a19325a );
 a3250a <=( a19316a  and  a19305a );
 a3251a <=( a19296a  and  a19285a );
 a3252a <=( a19276a  and  a19265a );
 a3253a <=( a19256a  and  a19245a );
 a3254a <=( a19236a  and  a19225a );
 a3255a <=( a19216a  and  a19205a );
 a3256a <=( a19196a  and  a19185a );
 a3257a <=( a19176a  and  a19165a );
 a3258a <=( a19156a  and  a19145a );
 a3259a <=( a19136a  and  a19125a );
 a3260a <=( a19116a  and  a19105a );
 a3261a <=( a19096a  and  a19085a );
 a3262a <=( a19076a  and  a19065a );
 a3263a <=( a19056a  and  a19045a );
 a3264a <=( a19036a  and  a19025a );
 a3265a <=( a19016a  and  a19005a );
 a3266a <=( a18996a  and  a18985a );
 a3267a <=( a18976a  and  a18965a );
 a3268a <=( a18956a  and  a18945a );
 a3269a <=( a18936a  and  a18925a );
 a3270a <=( a18916a  and  a18905a );
 a3271a <=( a18896a  and  a18885a );
 a3272a <=( a18876a  and  a18865a );
 a3273a <=( a18856a  and  a18845a );
 a3274a <=( a18836a  and  a18825a );
 a3275a <=( a18816a  and  a18805a );
 a3276a <=( a18796a  and  a18785a );
 a3277a <=( a18776a  and  a18765a );
 a3278a <=( a18756a  and  a18745a );
 a3279a <=( a18736a  and  a18725a );
 a3280a <=( a18716a  and  a18705a );
 a3281a <=( a18696a  and  a18685a );
 a3282a <=( a18676a  and  a18665a );
 a3283a <=( a18656a  and  a18645a );
 a3284a <=( a18636a  and  a18625a );
 a3285a <=( a18616a  and  a18605a );
 a3286a <=( a18596a  and  a18585a );
 a3287a <=( a18576a  and  a18565a );
 a3288a <=( a18556a  and  a18545a );
 a3289a <=( a18536a  and  a18525a );
 a3290a <=( a18516a  and  a18505a );
 a3291a <=( a18496a  and  a18485a );
 a3292a <=( a18476a  and  a18465a );
 a3293a <=( a18456a  and  a18445a );
 a3294a <=( a18436a  and  a18425a );
 a3295a <=( a18416a  and  a18405a );
 a3296a <=( a18396a  and  a18385a );
 a3297a <=( a18376a  and  a18365a );
 a3298a <=( a18356a  and  a18345a );
 a3299a <=( a18336a  and  a18325a );
 a3300a <=( a18316a  and  a18305a );
 a3301a <=( a18296a  and  a18285a );
 a3302a <=( a18276a  and  a18265a );
 a3303a <=( a18256a  and  a18245a );
 a3304a <=( a18236a  and  a18225a );
 a3305a <=( a18216a  and  a18205a );
 a3306a <=( a18196a  and  a18185a );
 a3307a <=( a18176a  and  a18165a );
 a3308a <=( a18156a  and  a18145a );
 a3309a <=( a18136a  and  a18125a );
 a3310a <=( a18116a  and  a18105a );
 a3311a <=( a18096a  and  a18085a );
 a3312a <=( a18076a  and  a18065a );
 a3313a <=( a18056a  and  a18045a );
 a3314a <=( a18036a  and  a18025a );
 a3315a <=( a18016a  and  a18005a );
 a3316a <=( a17996a  and  a17985a );
 a3317a <=( a17976a  and  a17965a );
 a3318a <=( a17956a  and  a17945a );
 a3319a <=( a17936a  and  a17925a );
 a3320a <=( a17916a  and  a17905a );
 a3321a <=( a17896a  and  a17885a );
 a3322a <=( a17876a  and  a17865a );
 a3323a <=( a17856a  and  a17845a );
 a3324a <=( a17836a  and  a17825a );
 a3325a <=( a17816a  and  a17805a );
 a3326a <=( a17796a  and  a17785a );
 a3327a <=( a17776a  and  a17765a );
 a3328a <=( a17756a  and  a17745a );
 a3329a <=( a17736a  and  a17725a );
 a3330a <=( a17716a  and  a17705a );
 a3331a <=( a17696a  and  a17685a );
 a3332a <=( a17676a  and  a17665a );
 a3333a <=( a17656a  and  a17645a );
 a3334a <=( a17636a  and  a17625a );
 a3335a <=( a17616a  and  a17605a );
 a3336a <=( a17596a  and  a17585a );
 a3337a <=( a17576a  and  a17565a );
 a3338a <=( a17556a  and  a17545a );
 a3339a <=( a17536a  and  a17525a );
 a3340a <=( a17516a  and  a17505a );
 a3341a <=( a17496a  and  a17485a );
 a3342a <=( a17476a  and  a17465a );
 a3343a <=( a17456a  and  a17445a );
 a3344a <=( a17436a  and  a17425a );
 a3345a <=( a17416a  and  a17405a );
 a3346a <=( a17396a  and  a17385a );
 a3347a <=( a17376a  and  a17365a );
 a3348a <=( a17356a  and  a17345a );
 a3349a <=( a17336a  and  a17325a );
 a3350a <=( a17316a  and  a17305a );
 a3351a <=( a17296a  and  a17285a );
 a3352a <=( a17276a  and  a17265a );
 a3353a <=( a17256a  and  a17245a );
 a3354a <=( a17236a  and  a17225a );
 a3355a <=( a17216a  and  a17205a );
 a3356a <=( a17196a  and  a17185a );
 a3357a <=( a17176a  and  a17165a );
 a3358a <=( a17156a  and  a17145a );
 a3359a <=( a17136a  and  a17125a );
 a3360a <=( a17116a  and  a17105a );
 a3361a <=( a17096a  and  a17085a );
 a3362a <=( a17076a  and  a17065a );
 a3363a <=( a17056a  and  a17045a );
 a3364a <=( a17036a  and  a17025a );
 a3365a <=( a17016a  and  a17005a );
 a3366a <=( a16996a  and  a16985a );
 a3367a <=( a16976a  and  a16965a );
 a3368a <=( a16956a  and  a16945a );
 a3369a <=( a16936a  and  a16925a );
 a3370a <=( a16916a  and  a16905a );
 a3371a <=( a16896a  and  a16885a );
 a3372a <=( a16876a  and  a16865a );
 a3373a <=( a16856a  and  a16845a );
 a3374a <=( a16836a  and  a16825a );
 a3375a <=( a16816a  and  a16807a );
 a3376a <=( a16798a  and  a16789a );
 a3377a <=( a16780a  and  a16771a );
 a3378a <=( a16762a  and  a16753a );
 a3379a <=( a16744a  and  a16735a );
 a3380a <=( a16726a  and  a16717a );
 a3381a <=( a16708a  and  a16699a );
 a3382a <=( a16690a  and  a16681a );
 a3383a <=( a16672a  and  a16663a );
 a3384a <=( a16654a  and  a16645a );
 a3385a <=( a16636a  and  a16627a );
 a3386a <=( a16618a  and  a16609a );
 a3387a <=( a16600a  and  a16591a );
 a3388a <=( a16582a  and  a16573a );
 a3389a <=( a16564a  and  a16555a );
 a3390a <=( a16546a  and  a16537a );
 a3391a <=( a16528a  and  a16519a );
 a3392a <=( a16510a  and  a16501a );
 a3393a <=( a16492a  and  a16483a );
 a3394a <=( a16474a  and  a16465a );
 a3395a <=( a16456a  and  a16447a );
 a3396a <=( a16438a  and  a16429a );
 a3397a <=( a16420a  and  a16411a );
 a3398a <=( a16402a  and  a16393a );
 a3399a <=( a16384a  and  a16375a );
 a3400a <=( a16366a  and  a16357a );
 a3401a <=( a16348a  and  a16339a );
 a3402a <=( a16330a  and  a16321a );
 a3403a <=( a16312a  and  a16303a );
 a3404a <=( a16294a  and  a16285a );
 a3405a <=( a16276a  and  a16267a );
 a3406a <=( a16258a  and  a16249a );
 a3407a <=( a16240a  and  a16231a );
 a3408a <=( a16222a  and  a16213a );
 a3409a <=( a16204a  and  a16195a );
 a3410a <=( a16186a  and  a16177a );
 a3411a <=( a16168a  and  a16159a );
 a3412a <=( a16150a  and  a16141a );
 a3413a <=( a16132a  and  a16123a );
 a3414a <=( a16114a  and  a16105a );
 a3415a <=( a16096a  and  a16087a );
 a3416a <=( a16078a  and  a16069a );
 a3417a <=( a16060a  and  a16051a );
 a3418a <=( a16042a  and  a16033a );
 a3419a <=( a16024a  and  a16015a );
 a3420a <=( a16006a  and  a15997a );
 a3421a <=( a15988a  and  a15979a );
 a3422a <=( a15970a  and  a15961a );
 a3423a <=( a15952a  and  a15943a );
 a3424a <=( a15934a  and  a15925a );
 a3425a <=( a15916a  and  a15907a );
 a3426a <=( a15898a  and  a15889a );
 a3427a <=( a15880a  and  a15871a );
 a3428a <=( a15862a  and  a15853a );
 a3429a <=( a15844a  and  a15835a );
 a3430a <=( a15826a  and  a15817a );
 a3431a <=( a15808a  and  a15799a );
 a3432a <=( a15790a  and  a15781a );
 a3433a <=( a15772a  and  a15763a );
 a3434a <=( a15754a  and  a15745a );
 a3435a <=( a15736a  and  a15727a );
 a3436a <=( a15718a  and  a15709a );
 a3437a <=( a15700a  and  a15691a );
 a3438a <=( a15682a  and  a15673a );
 a3439a <=( a15664a  and  a15655a );
 a3440a <=( a15646a  and  a15637a );
 a3441a <=( a15628a  and  a15619a );
 a3442a <=( a15610a  and  a15601a );
 a3443a <=( a15592a  and  a15583a );
 a3444a <=( a15574a  and  a15565a );
 a3445a <=( a15556a  and  a15547a );
 a3446a <=( a15538a  and  a15529a );
 a3447a <=( a15520a  and  a15511a );
 a3448a <=( a15502a  and  a15493a );
 a3449a <=( a15484a  and  a15475a );
 a3450a <=( a15466a  and  a15457a );
 a3451a <=( a15448a  and  a15439a );
 a3452a <=( a15430a  and  a15421a );
 a3453a <=( a15412a  and  a15403a );
 a3454a <=( a15394a  and  a15385a );
 a3455a <=( a15376a  and  a15367a );
 a3456a <=( a15358a  and  a15349a );
 a3457a <=( a15340a  and  a15331a );
 a3458a <=( a15322a  and  a15313a );
 a3459a <=( a15304a  and  a15295a );
 a3460a <=( a15286a  and  a15277a );
 a3461a <=( a15268a  and  a15259a );
 a3462a <=( a15250a  and  a15241a );
 a3463a <=( a15232a  and  a15223a );
 a3464a <=( a15214a  and  a15205a );
 a3465a <=( a15196a  and  a15187a );
 a3466a <=( a15178a  and  a15169a );
 a3467a <=( a15160a  and  a15151a );
 a3468a <=( a15142a  and  a15133a );
 a3469a <=( a15124a  and  a15115a );
 a3470a <=( a15106a  and  a15097a );
 a3471a <=( a15088a  and  a15079a );
 a3472a <=( a15070a  and  a15061a );
 a3473a <=( a15052a  and  a15043a );
 a3474a <=( a15034a  and  a15025a );
 a3475a <=( a15016a  and  a15007a );
 a3476a <=( a14998a  and  a14989a );
 a3477a <=( a14980a  and  a14971a );
 a3478a <=( a14962a  and  a14953a );
 a3479a <=( a14944a  and  a14935a );
 a3480a <=( a14926a  and  a14917a );
 a3481a <=( a14908a  and  a14899a );
 a3482a <=( a14890a  and  a14881a );
 a3483a <=( a14872a  and  a14863a );
 a3484a <=( a14854a  and  a14845a );
 a3485a <=( a14836a  and  a14827a );
 a3486a <=( a14818a  and  a14809a );
 a3487a <=( a14800a  and  a14791a );
 a3488a <=( a14782a  and  a14773a );
 a3489a <=( a14764a  and  a14755a );
 a3490a <=( a14746a  and  a14737a );
 a3491a <=( a14728a  and  a14719a );
 a3492a <=( a14710a  and  a14701a );
 a3493a <=( a14692a  and  a14683a );
 a3494a <=( a14674a  and  a14665a );
 a3495a <=( a14656a  and  a14647a );
 a3496a <=( a14638a  and  a14629a );
 a3497a <=( a14620a  and  a14611a );
 a3498a <=( a14602a  and  a14593a );
 a3499a <=( a14584a  and  a14575a );
 a3500a <=( a14566a  and  a14557a );
 a3501a <=( a14548a  and  a14539a );
 a3502a <=( a14530a  and  a14521a );
 a3503a <=( a14512a  and  a14503a );
 a3504a <=( a14494a  and  a14485a );
 a3505a <=( a14476a  and  a14467a );
 a3506a <=( a14458a  and  a14449a );
 a3507a <=( a14440a  and  a14431a );
 a3508a <=( a14422a  and  a14413a );
 a3509a <=( a14404a  and  a14395a );
 a3510a <=( a14386a  and  a14377a );
 a3511a <=( a14368a  and  a14359a );
 a3512a <=( a14350a  and  a14341a );
 a3513a <=( a14332a  and  a14323a );
 a3514a <=( a14314a  and  a14305a );
 a3515a <=( a14296a  and  a14287a );
 a3516a <=( a14278a  and  a14269a );
 a3517a <=( a14260a  and  a14251a );
 a3518a <=( a14242a  and  a14233a );
 a3519a <=( a14224a  and  a14215a );
 a3520a <=( a14206a  and  a14197a );
 a3521a <=( a14188a  and  a14179a );
 a3522a <=( a14170a  and  a14161a );
 a3523a <=( a14152a  and  a14143a );
 a3524a <=( a14134a  and  a14125a );
 a3525a <=( a14116a  and  a14107a );
 a3526a <=( a14098a  and  a14089a );
 a3527a <=( a14080a  and  a14071a );
 a3528a <=( a14062a  and  a14053a );
 a3529a <=( a14044a  and  a14035a );
 a3530a <=( a14026a  and  a14017a );
 a3531a <=( a14008a  and  a13999a );
 a3532a <=( a13990a  and  a13981a );
 a3533a <=( a13972a  and  a13963a );
 a3534a <=( a13954a  and  a13945a );
 a3535a <=( a13936a  and  a13927a );
 a3536a <=( a13918a  and  a13909a );
 a3537a <=( a13900a  and  a13891a );
 a3538a <=( a13882a  and  a13873a );
 a3539a <=( a13864a  and  a13855a );
 a3540a <=( a13846a  and  a13837a );
 a3541a <=( a13828a  and  a13819a );
 a3542a <=( a13810a  and  a13801a );
 a3543a <=( a13792a  and  a13783a );
 a3544a <=( a13774a  and  a13765a );
 a3545a <=( a13756a  and  a13747a );
 a3546a <=( a13738a  and  a13729a );
 a3547a <=( a13720a  and  a13711a );
 a3548a <=( a13702a  and  a13693a );
 a3549a <=( a13684a  and  a13675a );
 a3550a <=( a13666a  and  a13657a );
 a3551a <=( a13648a  and  a13639a );
 a3552a <=( a13630a  and  a13621a );
 a3553a <=( a13612a  and  a13603a );
 a3554a <=( a13594a  and  a13585a );
 a3555a <=( a13576a  and  a13567a );
 a3556a <=( a13558a  and  a13549a );
 a3557a <=( a13540a  and  a13531a );
 a3558a <=( a13522a  and  a13513a );
 a3559a <=( a13504a  and  a13495a );
 a3560a <=( a13486a  and  a13477a );
 a3561a <=( a13468a  and  a13459a );
 a3562a <=( a13450a  and  a13441a );
 a3563a <=( a13432a  and  a13423a );
 a3564a <=( a13414a  and  a13405a );
 a3565a <=( a13396a  and  a13387a );
 a3566a <=( a13378a  and  a13369a );
 a3567a <=( a13360a  and  a13351a );
 a3568a <=( a13342a  and  a13333a );
 a3569a <=( a13324a  and  a13315a );
 a3570a <=( a13306a  and  a13297a );
 a3571a <=( a13288a  and  a13279a );
 a3572a <=( a13270a  and  a13261a );
 a3573a <=( a13252a  and  a13243a );
 a3574a <=( a13234a  and  a13225a );
 a3575a <=( a13216a  and  a13207a );
 a3576a <=( a13198a  and  a13189a );
 a3577a <=( a13180a  and  a13171a );
 a3578a <=( a13162a  and  a13153a );
 a3579a <=( a13144a  and  a13135a );
 a3580a <=( a13126a  and  a13117a );
 a3581a <=( a13108a  and  a13099a );
 a3582a <=( a13090a  and  a13081a );
 a3583a <=( a13072a  and  a13063a );
 a3584a <=( a13054a  and  a13045a );
 a3585a <=( a13036a  and  a13027a );
 a3586a <=( a13018a  and  a13009a );
 a3587a <=( a13000a  and  a12991a );
 a3588a <=( a12982a  and  a12973a );
 a3589a <=( a12964a  and  a12955a );
 a3590a <=( a12946a  and  a12937a );
 a3591a <=( a12928a  and  a12919a );
 a3592a <=( a12910a  and  a12901a );
 a3593a <=( a12892a  and  a12883a );
 a3594a <=( a12874a  and  a12865a );
 a3595a <=( a12856a  and  a12847a );
 a3596a <=( a12838a  and  a12829a );
 a3597a <=( a12820a  and  a12811a );
 a3598a <=( a12802a  and  a12793a );
 a3599a <=( a12784a  and  a12775a );
 a3600a <=( a12766a  and  a12757a );
 a3601a <=( a12748a  and  a12739a );
 a3602a <=( a12730a  and  a12721a );
 a3603a <=( a12712a  and  a12703a );
 a3604a <=( a12694a  and  a12685a );
 a3605a <=( a12676a  and  a12667a );
 a3606a <=( a12658a  and  a12649a );
 a3607a <=( a12640a  and  a12631a );
 a3608a <=( a12622a  and  a12613a );
 a3609a <=( a12604a  and  a12595a );
 a3610a <=( a12586a  and  a12577a );
 a3611a <=( a12568a  and  a12559a );
 a3612a <=( a12550a  and  a12541a );
 a3613a <=( a12532a  and  a12523a );
 a3614a <=( a12514a  and  a12505a );
 a3615a <=( a12496a  and  a12487a );
 a3616a <=( a12478a  and  a12469a );
 a3617a <=( a12460a  and  a12451a );
 a3618a <=( a12442a  and  a12433a );
 a3619a <=( a12424a  and  a12415a );
 a3620a <=( a12406a  and  a12397a );
 a3621a <=( a12388a  and  a12379a );
 a3622a <=( a12370a  and  a12361a );
 a3623a <=( a12352a  and  a12343a );
 a3624a <=( a12334a  and  a12325a );
 a3625a <=( a12316a  and  a12307a );
 a3626a <=( a12298a  and  a12289a );
 a3627a <=( a12280a  and  a12271a );
 a3628a <=( a12262a  and  a12253a );
 a3629a <=( a12244a  and  a12235a );
 a3630a <=( a12226a  and  a12217a );
 a3631a <=( a12208a  and  a12199a );
 a3632a <=( a12190a  and  a12181a );
 a3633a <=( a12172a  and  a12163a );
 a3634a <=( a12154a  and  a12145a );
 a3635a <=( a12136a  and  a12127a );
 a3636a <=( a12118a  and  a12109a );
 a3637a <=( a12100a  and  a12091a );
 a3638a <=( a12082a  and  a12073a );
 a3639a <=( a12064a  and  a12055a );
 a3640a <=( a12048a  and  a12039a );
 a3641a <=( a12032a  and  a12023a );
 a3642a <=( a12016a  and  a12007a );
 a3643a <=( a12000a  and  a11991a );
 a3644a <=( a11984a  and  a11975a );
 a3645a <=( a11968a  and  a11959a );
 a3646a <=( a11952a  and  a11943a );
 a3647a <=( a11936a  and  a11927a );
 a3648a <=( a11920a  and  a11911a );
 a3649a <=( a11904a  and  a11895a );
 a3650a <=( a11888a  and  a11879a );
 a3651a <=( a11872a  and  a11863a );
 a3652a <=( a11856a  and  a11847a );
 a3653a <=( a11840a  and  a11831a );
 a3654a <=( a11824a  and  a11815a );
 a3655a <=( a11808a  and  a11799a );
 a3656a <=( a11792a  and  a11783a );
 a3657a <=( a11776a  and  a11767a );
 a3658a <=( a11760a  and  a11751a );
 a3659a <=( a11744a  and  a11735a );
 a3660a <=( a11728a  and  a11719a );
 a3661a <=( a11712a  and  a11703a );
 a3662a <=( a11696a  and  a11687a );
 a3663a <=( a11680a  and  a11671a );
 a3664a <=( a11664a  and  a11655a );
 a3665a <=( a11648a  and  a11639a );
 a3666a <=( a11632a  and  a11623a );
 a3667a <=( a11616a  and  a11607a );
 a3668a <=( a11600a  and  a11591a );
 a3669a <=( a11584a  and  a11575a );
 a3670a <=( a11568a  and  a11559a );
 a3671a <=( a11552a  and  a11545a );
 a3672a <=( a11538a  and  a11531a );
 a3673a <=( a11524a  and  a11517a );
 a3674a <=( a11510a  and  a11503a );
 a3675a <=( a11496a  and  a11489a );
 a3676a <=( a11482a  and  a11475a );
 a3677a <=( a11468a  and  a11461a );
 a3678a <=( a11454a  and  a11447a );
 a3679a <=( a11440a  and  a11433a );
 a3680a <=( a11426a  and  a11419a );
 a3681a <=( a11412a  and  a11405a );
 a3682a <=( a11398a  and  a11391a );
 a3683a <=( a11384a  and  a11377a );
 a3684a <=( a11370a  and  a11363a );
 a3685a <=( a11356a  and  a11349a );
 a3686a <=( a11342a  and  a11335a );
 a3687a <=( a11328a  and  a11321a );
 a3688a <=( a11314a  and  a11307a );
 a3689a <=( a11300a  and  a11293a );
 a3690a <=( a11286a  and  a11279a );
 a3691a <=( a11272a  and  a11265a );
 a3692a <=( a11258a  and  a11251a );
 a3693a <=( a11244a  and  a11237a );
 a3694a <=( a11230a  and  a11223a );
 a3695a <=( a11216a  and  a11209a );
 a3696a <=( a11202a  and  a11195a );
 a3697a <=( a11188a  and  a11181a );
 a3698a <=( a11174a  and  a11167a );
 a3699a <=( a11160a  and  a11153a );
 a3700a <=( a11146a  and  a11139a );
 a3701a <=( a11132a  and  a11125a );
 a3702a <=( a11118a  and  a11111a );
 a3706a <=( a3700a ) or ( a3701a );
 a3707a <=( a3702a ) or ( a3706a );
 a3710a <=( a3698a ) or ( a3699a );
 a3713a <=( a3696a ) or ( a3697a );
 a3714a <=( a3713a ) or ( a3710a );
 a3715a <=( a3714a ) or ( a3707a );
 a3719a <=( a3693a ) or ( a3694a );
 a3720a <=( a3695a ) or ( a3719a );
 a3723a <=( a3691a ) or ( a3692a );
 a3726a <=( a3689a ) or ( a3690a );
 a3727a <=( a3726a ) or ( a3723a );
 a3728a <=( a3727a ) or ( a3720a );
 a3729a <=( a3728a ) or ( a3715a );
 a3733a <=( a3686a ) or ( a3687a );
 a3734a <=( a3688a ) or ( a3733a );
 a3737a <=( a3684a ) or ( a3685a );
 a3740a <=( a3682a ) or ( a3683a );
 a3741a <=( a3740a ) or ( a3737a );
 a3742a <=( a3741a ) or ( a3734a );
 a3746a <=( a3679a ) or ( a3680a );
 a3747a <=( a3681a ) or ( a3746a );
 a3750a <=( a3677a ) or ( a3678a );
 a3753a <=( a3675a ) or ( a3676a );
 a3754a <=( a3753a ) or ( a3750a );
 a3755a <=( a3754a ) or ( a3747a );
 a3756a <=( a3755a ) or ( a3742a );
 a3757a <=( a3756a ) or ( a3729a );
 a3761a <=( a3672a ) or ( a3673a );
 a3762a <=( a3674a ) or ( a3761a );
 a3765a <=( a3670a ) or ( a3671a );
 a3768a <=( a3668a ) or ( a3669a );
 a3769a <=( a3768a ) or ( a3765a );
 a3770a <=( a3769a ) or ( a3762a );
 a3774a <=( a3665a ) or ( a3666a );
 a3775a <=( a3667a ) or ( a3774a );
 a3778a <=( a3663a ) or ( a3664a );
 a3781a <=( a3661a ) or ( a3662a );
 a3782a <=( a3781a ) or ( a3778a );
 a3783a <=( a3782a ) or ( a3775a );
 a3784a <=( a3783a ) or ( a3770a );
 a3788a <=( a3658a ) or ( a3659a );
 a3789a <=( a3660a ) or ( a3788a );
 a3792a <=( a3656a ) or ( a3657a );
 a3795a <=( a3654a ) or ( a3655a );
 a3796a <=( a3795a ) or ( a3792a );
 a3797a <=( a3796a ) or ( a3789a );
 a3800a <=( a3652a ) or ( a3653a );
 a3803a <=( a3650a ) or ( a3651a );
 a3804a <=( a3803a ) or ( a3800a );
 a3807a <=( a3648a ) or ( a3649a );
 a3810a <=( a3646a ) or ( a3647a );
 a3811a <=( a3810a ) or ( a3807a );
 a3812a <=( a3811a ) or ( a3804a );
 a3813a <=( a3812a ) or ( a3797a );
 a3814a <=( a3813a ) or ( a3784a );
 a3815a <=( a3814a ) or ( a3757a );
 a3819a <=( a3643a ) or ( a3644a );
 a3820a <=( a3645a ) or ( a3819a );
 a3823a <=( a3641a ) or ( a3642a );
 a3826a <=( a3639a ) or ( a3640a );
 a3827a <=( a3826a ) or ( a3823a );
 a3828a <=( a3827a ) or ( a3820a );
 a3832a <=( a3636a ) or ( a3637a );
 a3833a <=( a3638a ) or ( a3832a );
 a3836a <=( a3634a ) or ( a3635a );
 a3839a <=( a3632a ) or ( a3633a );
 a3840a <=( a3839a ) or ( a3836a );
 a3841a <=( a3840a ) or ( a3833a );
 a3842a <=( a3841a ) or ( a3828a );
 a3846a <=( a3629a ) or ( a3630a );
 a3847a <=( a3631a ) or ( a3846a );
 a3850a <=( a3627a ) or ( a3628a );
 a3853a <=( a3625a ) or ( a3626a );
 a3854a <=( a3853a ) or ( a3850a );
 a3855a <=( a3854a ) or ( a3847a );
 a3858a <=( a3623a ) or ( a3624a );
 a3861a <=( a3621a ) or ( a3622a );
 a3862a <=( a3861a ) or ( a3858a );
 a3865a <=( a3619a ) or ( a3620a );
 a3868a <=( a3617a ) or ( a3618a );
 a3869a <=( a3868a ) or ( a3865a );
 a3870a <=( a3869a ) or ( a3862a );
 a3871a <=( a3870a ) or ( a3855a );
 a3872a <=( a3871a ) or ( a3842a );
 a3876a <=( a3614a ) or ( a3615a );
 a3877a <=( a3616a ) or ( a3876a );
 a3880a <=( a3612a ) or ( a3613a );
 a3883a <=( a3610a ) or ( a3611a );
 a3884a <=( a3883a ) or ( a3880a );
 a3885a <=( a3884a ) or ( a3877a );
 a3889a <=( a3607a ) or ( a3608a );
 a3890a <=( a3609a ) or ( a3889a );
 a3893a <=( a3605a ) or ( a3606a );
 a3896a <=( a3603a ) or ( a3604a );
 a3897a <=( a3896a ) or ( a3893a );
 a3898a <=( a3897a ) or ( a3890a );
 a3899a <=( a3898a ) or ( a3885a );
 a3903a <=( a3600a ) or ( a3601a );
 a3904a <=( a3602a ) or ( a3903a );
 a3907a <=( a3598a ) or ( a3599a );
 a3910a <=( a3596a ) or ( a3597a );
 a3911a <=( a3910a ) or ( a3907a );
 a3912a <=( a3911a ) or ( a3904a );
 a3915a <=( a3594a ) or ( a3595a );
 a3918a <=( a3592a ) or ( a3593a );
 a3919a <=( a3918a ) or ( a3915a );
 a3922a <=( a3590a ) or ( a3591a );
 a3925a <=( a3588a ) or ( a3589a );
 a3926a <=( a3925a ) or ( a3922a );
 a3927a <=( a3926a ) or ( a3919a );
 a3928a <=( a3927a ) or ( a3912a );
 a3929a <=( a3928a ) or ( a3899a );
 a3930a <=( a3929a ) or ( a3872a );
 a3931a <=( a3930a ) or ( a3815a );
 a3935a <=( a3585a ) or ( a3586a );
 a3936a <=( a3587a ) or ( a3935a );
 a3939a <=( a3583a ) or ( a3584a );
 a3942a <=( a3581a ) or ( a3582a );
 a3943a <=( a3942a ) or ( a3939a );
 a3944a <=( a3943a ) or ( a3936a );
 a3948a <=( a3578a ) or ( a3579a );
 a3949a <=( a3580a ) or ( a3948a );
 a3952a <=( a3576a ) or ( a3577a );
 a3955a <=( a3574a ) or ( a3575a );
 a3956a <=( a3955a ) or ( a3952a );
 a3957a <=( a3956a ) or ( a3949a );
 a3958a <=( a3957a ) or ( a3944a );
 a3962a <=( a3571a ) or ( a3572a );
 a3963a <=( a3573a ) or ( a3962a );
 a3966a <=( a3569a ) or ( a3570a );
 a3969a <=( a3567a ) or ( a3568a );
 a3970a <=( a3969a ) or ( a3966a );
 a3971a <=( a3970a ) or ( a3963a );
 a3974a <=( a3565a ) or ( a3566a );
 a3977a <=( a3563a ) or ( a3564a );
 a3978a <=( a3977a ) or ( a3974a );
 a3981a <=( a3561a ) or ( a3562a );
 a3984a <=( a3559a ) or ( a3560a );
 a3985a <=( a3984a ) or ( a3981a );
 a3986a <=( a3985a ) or ( a3978a );
 a3987a <=( a3986a ) or ( a3971a );
 a3988a <=( a3987a ) or ( a3958a );
 a3992a <=( a3556a ) or ( a3557a );
 a3993a <=( a3558a ) or ( a3992a );
 a3996a <=( a3554a ) or ( a3555a );
 a3999a <=( a3552a ) or ( a3553a );
 a4000a <=( a3999a ) or ( a3996a );
 a4001a <=( a4000a ) or ( a3993a );
 a4005a <=( a3549a ) or ( a3550a );
 a4006a <=( a3551a ) or ( a4005a );
 a4009a <=( a3547a ) or ( a3548a );
 a4012a <=( a3545a ) or ( a3546a );
 a4013a <=( a4012a ) or ( a4009a );
 a4014a <=( a4013a ) or ( a4006a );
 a4015a <=( a4014a ) or ( a4001a );
 a4019a <=( a3542a ) or ( a3543a );
 a4020a <=( a3544a ) or ( a4019a );
 a4023a <=( a3540a ) or ( a3541a );
 a4026a <=( a3538a ) or ( a3539a );
 a4027a <=( a4026a ) or ( a4023a );
 a4028a <=( a4027a ) or ( a4020a );
 a4031a <=( a3536a ) or ( a3537a );
 a4034a <=( a3534a ) or ( a3535a );
 a4035a <=( a4034a ) or ( a4031a );
 a4038a <=( a3532a ) or ( a3533a );
 a4041a <=( a3530a ) or ( a3531a );
 a4042a <=( a4041a ) or ( a4038a );
 a4043a <=( a4042a ) or ( a4035a );
 a4044a <=( a4043a ) or ( a4028a );
 a4045a <=( a4044a ) or ( a4015a );
 a4046a <=( a4045a ) or ( a3988a );
 a4050a <=( a3527a ) or ( a3528a );
 a4051a <=( a3529a ) or ( a4050a );
 a4054a <=( a3525a ) or ( a3526a );
 a4057a <=( a3523a ) or ( a3524a );
 a4058a <=( a4057a ) or ( a4054a );
 a4059a <=( a4058a ) or ( a4051a );
 a4063a <=( a3520a ) or ( a3521a );
 a4064a <=( a3522a ) or ( a4063a );
 a4067a <=( a3518a ) or ( a3519a );
 a4070a <=( a3516a ) or ( a3517a );
 a4071a <=( a4070a ) or ( a4067a );
 a4072a <=( a4071a ) or ( a4064a );
 a4073a <=( a4072a ) or ( a4059a );
 a4077a <=( a3513a ) or ( a3514a );
 a4078a <=( a3515a ) or ( a4077a );
 a4081a <=( a3511a ) or ( a3512a );
 a4084a <=( a3509a ) or ( a3510a );
 a4085a <=( a4084a ) or ( a4081a );
 a4086a <=( a4085a ) or ( a4078a );
 a4089a <=( a3507a ) or ( a3508a );
 a4092a <=( a3505a ) or ( a3506a );
 a4093a <=( a4092a ) or ( a4089a );
 a4096a <=( a3503a ) or ( a3504a );
 a4099a <=( a3501a ) or ( a3502a );
 a4100a <=( a4099a ) or ( a4096a );
 a4101a <=( a4100a ) or ( a4093a );
 a4102a <=( a4101a ) or ( a4086a );
 a4103a <=( a4102a ) or ( a4073a );
 a4107a <=( a3498a ) or ( a3499a );
 a4108a <=( a3500a ) or ( a4107a );
 a4111a <=( a3496a ) or ( a3497a );
 a4114a <=( a3494a ) or ( a3495a );
 a4115a <=( a4114a ) or ( a4111a );
 a4116a <=( a4115a ) or ( a4108a );
 a4120a <=( a3491a ) or ( a3492a );
 a4121a <=( a3493a ) or ( a4120a );
 a4124a <=( a3489a ) or ( a3490a );
 a4127a <=( a3487a ) or ( a3488a );
 a4128a <=( a4127a ) or ( a4124a );
 a4129a <=( a4128a ) or ( a4121a );
 a4130a <=( a4129a ) or ( a4116a );
 a4134a <=( a3484a ) or ( a3485a );
 a4135a <=( a3486a ) or ( a4134a );
 a4138a <=( a3482a ) or ( a3483a );
 a4141a <=( a3480a ) or ( a3481a );
 a4142a <=( a4141a ) or ( a4138a );
 a4143a <=( a4142a ) or ( a4135a );
 a4146a <=( a3478a ) or ( a3479a );
 a4149a <=( a3476a ) or ( a3477a );
 a4150a <=( a4149a ) or ( a4146a );
 a4153a <=( a3474a ) or ( a3475a );
 a4156a <=( a3472a ) or ( a3473a );
 a4157a <=( a4156a ) or ( a4153a );
 a4158a <=( a4157a ) or ( a4150a );
 a4159a <=( a4158a ) or ( a4143a );
 a4160a <=( a4159a ) or ( a4130a );
 a4161a <=( a4160a ) or ( a4103a );
 a4162a <=( a4161a ) or ( a4046a );
 a4163a <=( a4162a ) or ( a3931a );
 a4167a <=( a3469a ) or ( a3470a );
 a4168a <=( a3471a ) or ( a4167a );
 a4171a <=( a3467a ) or ( a3468a );
 a4174a <=( a3465a ) or ( a3466a );
 a4175a <=( a4174a ) or ( a4171a );
 a4176a <=( a4175a ) or ( a4168a );
 a4180a <=( a3462a ) or ( a3463a );
 a4181a <=( a3464a ) or ( a4180a );
 a4184a <=( a3460a ) or ( a3461a );
 a4187a <=( a3458a ) or ( a3459a );
 a4188a <=( a4187a ) or ( a4184a );
 a4189a <=( a4188a ) or ( a4181a );
 a4190a <=( a4189a ) or ( a4176a );
 a4194a <=( a3455a ) or ( a3456a );
 a4195a <=( a3457a ) or ( a4194a );
 a4198a <=( a3453a ) or ( a3454a );
 a4201a <=( a3451a ) or ( a3452a );
 a4202a <=( a4201a ) or ( a4198a );
 a4203a <=( a4202a ) or ( a4195a );
 a4207a <=( a3448a ) or ( a3449a );
 a4208a <=( a3450a ) or ( a4207a );
 a4211a <=( a3446a ) or ( a3447a );
 a4214a <=( a3444a ) or ( a3445a );
 a4215a <=( a4214a ) or ( a4211a );
 a4216a <=( a4215a ) or ( a4208a );
 a4217a <=( a4216a ) or ( a4203a );
 a4218a <=( a4217a ) or ( a4190a );
 a4222a <=( a3441a ) or ( a3442a );
 a4223a <=( a3443a ) or ( a4222a );
 a4226a <=( a3439a ) or ( a3440a );
 a4229a <=( a3437a ) or ( a3438a );
 a4230a <=( a4229a ) or ( a4226a );
 a4231a <=( a4230a ) or ( a4223a );
 a4235a <=( a3434a ) or ( a3435a );
 a4236a <=( a3436a ) or ( a4235a );
 a4239a <=( a3432a ) or ( a3433a );
 a4242a <=( a3430a ) or ( a3431a );
 a4243a <=( a4242a ) or ( a4239a );
 a4244a <=( a4243a ) or ( a4236a );
 a4245a <=( a4244a ) or ( a4231a );
 a4249a <=( a3427a ) or ( a3428a );
 a4250a <=( a3429a ) or ( a4249a );
 a4253a <=( a3425a ) or ( a3426a );
 a4256a <=( a3423a ) or ( a3424a );
 a4257a <=( a4256a ) or ( a4253a );
 a4258a <=( a4257a ) or ( a4250a );
 a4261a <=( a3421a ) or ( a3422a );
 a4264a <=( a3419a ) or ( a3420a );
 a4265a <=( a4264a ) or ( a4261a );
 a4268a <=( a3417a ) or ( a3418a );
 a4271a <=( a3415a ) or ( a3416a );
 a4272a <=( a4271a ) or ( a4268a );
 a4273a <=( a4272a ) or ( a4265a );
 a4274a <=( a4273a ) or ( a4258a );
 a4275a <=( a4274a ) or ( a4245a );
 a4276a <=( a4275a ) or ( a4218a );
 a4280a <=( a3412a ) or ( a3413a );
 a4281a <=( a3414a ) or ( a4280a );
 a4284a <=( a3410a ) or ( a3411a );
 a4287a <=( a3408a ) or ( a3409a );
 a4288a <=( a4287a ) or ( a4284a );
 a4289a <=( a4288a ) or ( a4281a );
 a4293a <=( a3405a ) or ( a3406a );
 a4294a <=( a3407a ) or ( a4293a );
 a4297a <=( a3403a ) or ( a3404a );
 a4300a <=( a3401a ) or ( a3402a );
 a4301a <=( a4300a ) or ( a4297a );
 a4302a <=( a4301a ) or ( a4294a );
 a4303a <=( a4302a ) or ( a4289a );
 a4307a <=( a3398a ) or ( a3399a );
 a4308a <=( a3400a ) or ( a4307a );
 a4311a <=( a3396a ) or ( a3397a );
 a4314a <=( a3394a ) or ( a3395a );
 a4315a <=( a4314a ) or ( a4311a );
 a4316a <=( a4315a ) or ( a4308a );
 a4319a <=( a3392a ) or ( a3393a );
 a4322a <=( a3390a ) or ( a3391a );
 a4323a <=( a4322a ) or ( a4319a );
 a4326a <=( a3388a ) or ( a3389a );
 a4329a <=( a3386a ) or ( a3387a );
 a4330a <=( a4329a ) or ( a4326a );
 a4331a <=( a4330a ) or ( a4323a );
 a4332a <=( a4331a ) or ( a4316a );
 a4333a <=( a4332a ) or ( a4303a );
 a4337a <=( a3383a ) or ( a3384a );
 a4338a <=( a3385a ) or ( a4337a );
 a4341a <=( a3381a ) or ( a3382a );
 a4344a <=( a3379a ) or ( a3380a );
 a4345a <=( a4344a ) or ( a4341a );
 a4346a <=( a4345a ) or ( a4338a );
 a4350a <=( a3376a ) or ( a3377a );
 a4351a <=( a3378a ) or ( a4350a );
 a4354a <=( a3374a ) or ( a3375a );
 a4357a <=( a3372a ) or ( a3373a );
 a4358a <=( a4357a ) or ( a4354a );
 a4359a <=( a4358a ) or ( a4351a );
 a4360a <=( a4359a ) or ( a4346a );
 a4364a <=( a3369a ) or ( a3370a );
 a4365a <=( a3371a ) or ( a4364a );
 a4368a <=( a3367a ) or ( a3368a );
 a4371a <=( a3365a ) or ( a3366a );
 a4372a <=( a4371a ) or ( a4368a );
 a4373a <=( a4372a ) or ( a4365a );
 a4376a <=( a3363a ) or ( a3364a );
 a4379a <=( a3361a ) or ( a3362a );
 a4380a <=( a4379a ) or ( a4376a );
 a4383a <=( a3359a ) or ( a3360a );
 a4386a <=( a3357a ) or ( a3358a );
 a4387a <=( a4386a ) or ( a4383a );
 a4388a <=( a4387a ) or ( a4380a );
 a4389a <=( a4388a ) or ( a4373a );
 a4390a <=( a4389a ) or ( a4360a );
 a4391a <=( a4390a ) or ( a4333a );
 a4392a <=( a4391a ) or ( a4276a );
 a4396a <=( a3354a ) or ( a3355a );
 a4397a <=( a3356a ) or ( a4396a );
 a4400a <=( a3352a ) or ( a3353a );
 a4403a <=( a3350a ) or ( a3351a );
 a4404a <=( a4403a ) or ( a4400a );
 a4405a <=( a4404a ) or ( a4397a );
 a4409a <=( a3347a ) or ( a3348a );
 a4410a <=( a3349a ) or ( a4409a );
 a4413a <=( a3345a ) or ( a3346a );
 a4416a <=( a3343a ) or ( a3344a );
 a4417a <=( a4416a ) or ( a4413a );
 a4418a <=( a4417a ) or ( a4410a );
 a4419a <=( a4418a ) or ( a4405a );
 a4423a <=( a3340a ) or ( a3341a );
 a4424a <=( a3342a ) or ( a4423a );
 a4427a <=( a3338a ) or ( a3339a );
 a4430a <=( a3336a ) or ( a3337a );
 a4431a <=( a4430a ) or ( a4427a );
 a4432a <=( a4431a ) or ( a4424a );
 a4435a <=( a3334a ) or ( a3335a );
 a4438a <=( a3332a ) or ( a3333a );
 a4439a <=( a4438a ) or ( a4435a );
 a4442a <=( a3330a ) or ( a3331a );
 a4445a <=( a3328a ) or ( a3329a );
 a4446a <=( a4445a ) or ( a4442a );
 a4447a <=( a4446a ) or ( a4439a );
 a4448a <=( a4447a ) or ( a4432a );
 a4449a <=( a4448a ) or ( a4419a );
 a4453a <=( a3325a ) or ( a3326a );
 a4454a <=( a3327a ) or ( a4453a );
 a4457a <=( a3323a ) or ( a3324a );
 a4460a <=( a3321a ) or ( a3322a );
 a4461a <=( a4460a ) or ( a4457a );
 a4462a <=( a4461a ) or ( a4454a );
 a4466a <=( a3318a ) or ( a3319a );
 a4467a <=( a3320a ) or ( a4466a );
 a4470a <=( a3316a ) or ( a3317a );
 a4473a <=( a3314a ) or ( a3315a );
 a4474a <=( a4473a ) or ( a4470a );
 a4475a <=( a4474a ) or ( a4467a );
 a4476a <=( a4475a ) or ( a4462a );
 a4480a <=( a3311a ) or ( a3312a );
 a4481a <=( a3313a ) or ( a4480a );
 a4484a <=( a3309a ) or ( a3310a );
 a4487a <=( a3307a ) or ( a3308a );
 a4488a <=( a4487a ) or ( a4484a );
 a4489a <=( a4488a ) or ( a4481a );
 a4492a <=( a3305a ) or ( a3306a );
 a4495a <=( a3303a ) or ( a3304a );
 a4496a <=( a4495a ) or ( a4492a );
 a4499a <=( a3301a ) or ( a3302a );
 a4502a <=( a3299a ) or ( a3300a );
 a4503a <=( a4502a ) or ( a4499a );
 a4504a <=( a4503a ) or ( a4496a );
 a4505a <=( a4504a ) or ( a4489a );
 a4506a <=( a4505a ) or ( a4476a );
 a4507a <=( a4506a ) or ( a4449a );
 a4511a <=( a3296a ) or ( a3297a );
 a4512a <=( a3298a ) or ( a4511a );
 a4515a <=( a3294a ) or ( a3295a );
 a4518a <=( a3292a ) or ( a3293a );
 a4519a <=( a4518a ) or ( a4515a );
 a4520a <=( a4519a ) or ( a4512a );
 a4524a <=( a3289a ) or ( a3290a );
 a4525a <=( a3291a ) or ( a4524a );
 a4528a <=( a3287a ) or ( a3288a );
 a4531a <=( a3285a ) or ( a3286a );
 a4532a <=( a4531a ) or ( a4528a );
 a4533a <=( a4532a ) or ( a4525a );
 a4534a <=( a4533a ) or ( a4520a );
 a4538a <=( a3282a ) or ( a3283a );
 a4539a <=( a3284a ) or ( a4538a );
 a4542a <=( a3280a ) or ( a3281a );
 a4545a <=( a3278a ) or ( a3279a );
 a4546a <=( a4545a ) or ( a4542a );
 a4547a <=( a4546a ) or ( a4539a );
 a4550a <=( a3276a ) or ( a3277a );
 a4553a <=( a3274a ) or ( a3275a );
 a4554a <=( a4553a ) or ( a4550a );
 a4557a <=( a3272a ) or ( a3273a );
 a4560a <=( a3270a ) or ( a3271a );
 a4561a <=( a4560a ) or ( a4557a );
 a4562a <=( a4561a ) or ( a4554a );
 a4563a <=( a4562a ) or ( a4547a );
 a4564a <=( a4563a ) or ( a4534a );
 a4568a <=( a3267a ) or ( a3268a );
 a4569a <=( a3269a ) or ( a4568a );
 a4572a <=( a3265a ) or ( a3266a );
 a4575a <=( a3263a ) or ( a3264a );
 a4576a <=( a4575a ) or ( a4572a );
 a4577a <=( a4576a ) or ( a4569a );
 a4581a <=( a3260a ) or ( a3261a );
 a4582a <=( a3262a ) or ( a4581a );
 a4585a <=( a3258a ) or ( a3259a );
 a4588a <=( a3256a ) or ( a3257a );
 a4589a <=( a4588a ) or ( a4585a );
 a4590a <=( a4589a ) or ( a4582a );
 a4591a <=( a4590a ) or ( a4577a );
 a4595a <=( a3253a ) or ( a3254a );
 a4596a <=( a3255a ) or ( a4595a );
 a4599a <=( a3251a ) or ( a3252a );
 a4602a <=( a3249a ) or ( a3250a );
 a4603a <=( a4602a ) or ( a4599a );
 a4604a <=( a4603a ) or ( a4596a );
 a4607a <=( a3247a ) or ( a3248a );
 a4610a <=( a3245a ) or ( a3246a );
 a4611a <=( a4610a ) or ( a4607a );
 a4614a <=( a3243a ) or ( a3244a );
 a4617a <=( a3241a ) or ( a3242a );
 a4618a <=( a4617a ) or ( a4614a );
 a4619a <=( a4618a ) or ( a4611a );
 a4620a <=( a4619a ) or ( a4604a );
 a4621a <=( a4620a ) or ( a4591a );
 a4622a <=( a4621a ) or ( a4564a );
 a4623a <=( a4622a ) or ( a4507a );
 a4624a <=( a4623a ) or ( a4392a );
 a4625a <=( a4624a ) or ( a4163a );
 a4629a <=( a3238a ) or ( a3239a );
 a4630a <=( a3240a ) or ( a4629a );
 a4633a <=( a3236a ) or ( a3237a );
 a4636a <=( a3234a ) or ( a3235a );
 a4637a <=( a4636a ) or ( a4633a );
 a4638a <=( a4637a ) or ( a4630a );
 a4642a <=( a3231a ) or ( a3232a );
 a4643a <=( a3233a ) or ( a4642a );
 a4646a <=( a3229a ) or ( a3230a );
 a4649a <=( a3227a ) or ( a3228a );
 a4650a <=( a4649a ) or ( a4646a );
 a4651a <=( a4650a ) or ( a4643a );
 a4652a <=( a4651a ) or ( a4638a );
 a4656a <=( a3224a ) or ( a3225a );
 a4657a <=( a3226a ) or ( a4656a );
 a4660a <=( a3222a ) or ( a3223a );
 a4663a <=( a3220a ) or ( a3221a );
 a4664a <=( a4663a ) or ( a4660a );
 a4665a <=( a4664a ) or ( a4657a );
 a4669a <=( a3217a ) or ( a3218a );
 a4670a <=( a3219a ) or ( a4669a );
 a4673a <=( a3215a ) or ( a3216a );
 a4676a <=( a3213a ) or ( a3214a );
 a4677a <=( a4676a ) or ( a4673a );
 a4678a <=( a4677a ) or ( a4670a );
 a4679a <=( a4678a ) or ( a4665a );
 a4680a <=( a4679a ) or ( a4652a );
 a4684a <=( a3210a ) or ( a3211a );
 a4685a <=( a3212a ) or ( a4684a );
 a4688a <=( a3208a ) or ( a3209a );
 a4691a <=( a3206a ) or ( a3207a );
 a4692a <=( a4691a ) or ( a4688a );
 a4693a <=( a4692a ) or ( a4685a );
 a4697a <=( a3203a ) or ( a3204a );
 a4698a <=( a3205a ) or ( a4697a );
 a4701a <=( a3201a ) or ( a3202a );
 a4704a <=( a3199a ) or ( a3200a );
 a4705a <=( a4704a ) or ( a4701a );
 a4706a <=( a4705a ) or ( a4698a );
 a4707a <=( a4706a ) or ( a4693a );
 a4711a <=( a3196a ) or ( a3197a );
 a4712a <=( a3198a ) or ( a4711a );
 a4715a <=( a3194a ) or ( a3195a );
 a4718a <=( a3192a ) or ( a3193a );
 a4719a <=( a4718a ) or ( a4715a );
 a4720a <=( a4719a ) or ( a4712a );
 a4723a <=( a3190a ) or ( a3191a );
 a4726a <=( a3188a ) or ( a3189a );
 a4727a <=( a4726a ) or ( a4723a );
 a4730a <=( a3186a ) or ( a3187a );
 a4733a <=( a3184a ) or ( a3185a );
 a4734a <=( a4733a ) or ( a4730a );
 a4735a <=( a4734a ) or ( a4727a );
 a4736a <=( a4735a ) or ( a4720a );
 a4737a <=( a4736a ) or ( a4707a );
 a4738a <=( a4737a ) or ( a4680a );
 a4742a <=( a3181a ) or ( a3182a );
 a4743a <=( a3183a ) or ( a4742a );
 a4746a <=( a3179a ) or ( a3180a );
 a4749a <=( a3177a ) or ( a3178a );
 a4750a <=( a4749a ) or ( a4746a );
 a4751a <=( a4750a ) or ( a4743a );
 a4755a <=( a3174a ) or ( a3175a );
 a4756a <=( a3176a ) or ( a4755a );
 a4759a <=( a3172a ) or ( a3173a );
 a4762a <=( a3170a ) or ( a3171a );
 a4763a <=( a4762a ) or ( a4759a );
 a4764a <=( a4763a ) or ( a4756a );
 a4765a <=( a4764a ) or ( a4751a );
 a4769a <=( a3167a ) or ( a3168a );
 a4770a <=( a3169a ) or ( a4769a );
 a4773a <=( a3165a ) or ( a3166a );
 a4776a <=( a3163a ) or ( a3164a );
 a4777a <=( a4776a ) or ( a4773a );
 a4778a <=( a4777a ) or ( a4770a );
 a4781a <=( a3161a ) or ( a3162a );
 a4784a <=( a3159a ) or ( a3160a );
 a4785a <=( a4784a ) or ( a4781a );
 a4788a <=( a3157a ) or ( a3158a );
 a4791a <=( a3155a ) or ( a3156a );
 a4792a <=( a4791a ) or ( a4788a );
 a4793a <=( a4792a ) or ( a4785a );
 a4794a <=( a4793a ) or ( a4778a );
 a4795a <=( a4794a ) or ( a4765a );
 a4799a <=( a3152a ) or ( a3153a );
 a4800a <=( a3154a ) or ( a4799a );
 a4803a <=( a3150a ) or ( a3151a );
 a4806a <=( a3148a ) or ( a3149a );
 a4807a <=( a4806a ) or ( a4803a );
 a4808a <=( a4807a ) or ( a4800a );
 a4812a <=( a3145a ) or ( a3146a );
 a4813a <=( a3147a ) or ( a4812a );
 a4816a <=( a3143a ) or ( a3144a );
 a4819a <=( a3141a ) or ( a3142a );
 a4820a <=( a4819a ) or ( a4816a );
 a4821a <=( a4820a ) or ( a4813a );
 a4822a <=( a4821a ) or ( a4808a );
 a4826a <=( a3138a ) or ( a3139a );
 a4827a <=( a3140a ) or ( a4826a );
 a4830a <=( a3136a ) or ( a3137a );
 a4833a <=( a3134a ) or ( a3135a );
 a4834a <=( a4833a ) or ( a4830a );
 a4835a <=( a4834a ) or ( a4827a );
 a4838a <=( a3132a ) or ( a3133a );
 a4841a <=( a3130a ) or ( a3131a );
 a4842a <=( a4841a ) or ( a4838a );
 a4845a <=( a3128a ) or ( a3129a );
 a4848a <=( a3126a ) or ( a3127a );
 a4849a <=( a4848a ) or ( a4845a );
 a4850a <=( a4849a ) or ( a4842a );
 a4851a <=( a4850a ) or ( a4835a );
 a4852a <=( a4851a ) or ( a4822a );
 a4853a <=( a4852a ) or ( a4795a );
 a4854a <=( a4853a ) or ( a4738a );
 a4858a <=( a3123a ) or ( a3124a );
 a4859a <=( a3125a ) or ( a4858a );
 a4862a <=( a3121a ) or ( a3122a );
 a4865a <=( a3119a ) or ( a3120a );
 a4866a <=( a4865a ) or ( a4862a );
 a4867a <=( a4866a ) or ( a4859a );
 a4871a <=( a3116a ) or ( a3117a );
 a4872a <=( a3118a ) or ( a4871a );
 a4875a <=( a3114a ) or ( a3115a );
 a4878a <=( a3112a ) or ( a3113a );
 a4879a <=( a4878a ) or ( a4875a );
 a4880a <=( a4879a ) or ( a4872a );
 a4881a <=( a4880a ) or ( a4867a );
 a4885a <=( a3109a ) or ( a3110a );
 a4886a <=( a3111a ) or ( a4885a );
 a4889a <=( a3107a ) or ( a3108a );
 a4892a <=( a3105a ) or ( a3106a );
 a4893a <=( a4892a ) or ( a4889a );
 a4894a <=( a4893a ) or ( a4886a );
 a4897a <=( a3103a ) or ( a3104a );
 a4900a <=( a3101a ) or ( a3102a );
 a4901a <=( a4900a ) or ( a4897a );
 a4904a <=( a3099a ) or ( a3100a );
 a4907a <=( a3097a ) or ( a3098a );
 a4908a <=( a4907a ) or ( a4904a );
 a4909a <=( a4908a ) or ( a4901a );
 a4910a <=( a4909a ) or ( a4894a );
 a4911a <=( a4910a ) or ( a4881a );
 a4915a <=( a3094a ) or ( a3095a );
 a4916a <=( a3096a ) or ( a4915a );
 a4919a <=( a3092a ) or ( a3093a );
 a4922a <=( a3090a ) or ( a3091a );
 a4923a <=( a4922a ) or ( a4919a );
 a4924a <=( a4923a ) or ( a4916a );
 a4928a <=( a3087a ) or ( a3088a );
 a4929a <=( a3089a ) or ( a4928a );
 a4932a <=( a3085a ) or ( a3086a );
 a4935a <=( a3083a ) or ( a3084a );
 a4936a <=( a4935a ) or ( a4932a );
 a4937a <=( a4936a ) or ( a4929a );
 a4938a <=( a4937a ) or ( a4924a );
 a4942a <=( a3080a ) or ( a3081a );
 a4943a <=( a3082a ) or ( a4942a );
 a4946a <=( a3078a ) or ( a3079a );
 a4949a <=( a3076a ) or ( a3077a );
 a4950a <=( a4949a ) or ( a4946a );
 a4951a <=( a4950a ) or ( a4943a );
 a4954a <=( a3074a ) or ( a3075a );
 a4957a <=( a3072a ) or ( a3073a );
 a4958a <=( a4957a ) or ( a4954a );
 a4961a <=( a3070a ) or ( a3071a );
 a4964a <=( a3068a ) or ( a3069a );
 a4965a <=( a4964a ) or ( a4961a );
 a4966a <=( a4965a ) or ( a4958a );
 a4967a <=( a4966a ) or ( a4951a );
 a4968a <=( a4967a ) or ( a4938a );
 a4969a <=( a4968a ) or ( a4911a );
 a4973a <=( a3065a ) or ( a3066a );
 a4974a <=( a3067a ) or ( a4973a );
 a4977a <=( a3063a ) or ( a3064a );
 a4980a <=( a3061a ) or ( a3062a );
 a4981a <=( a4980a ) or ( a4977a );
 a4982a <=( a4981a ) or ( a4974a );
 a4986a <=( a3058a ) or ( a3059a );
 a4987a <=( a3060a ) or ( a4986a );
 a4990a <=( a3056a ) or ( a3057a );
 a4993a <=( a3054a ) or ( a3055a );
 a4994a <=( a4993a ) or ( a4990a );
 a4995a <=( a4994a ) or ( a4987a );
 a4996a <=( a4995a ) or ( a4982a );
 a5000a <=( a3051a ) or ( a3052a );
 a5001a <=( a3053a ) or ( a5000a );
 a5004a <=( a3049a ) or ( a3050a );
 a5007a <=( a3047a ) or ( a3048a );
 a5008a <=( a5007a ) or ( a5004a );
 a5009a <=( a5008a ) or ( a5001a );
 a5012a <=( a3045a ) or ( a3046a );
 a5015a <=( a3043a ) or ( a3044a );
 a5016a <=( a5015a ) or ( a5012a );
 a5019a <=( a3041a ) or ( a3042a );
 a5022a <=( a3039a ) or ( a3040a );
 a5023a <=( a5022a ) or ( a5019a );
 a5024a <=( a5023a ) or ( a5016a );
 a5025a <=( a5024a ) or ( a5009a );
 a5026a <=( a5025a ) or ( a4996a );
 a5030a <=( a3036a ) or ( a3037a );
 a5031a <=( a3038a ) or ( a5030a );
 a5034a <=( a3034a ) or ( a3035a );
 a5037a <=( a3032a ) or ( a3033a );
 a5038a <=( a5037a ) or ( a5034a );
 a5039a <=( a5038a ) or ( a5031a );
 a5043a <=( a3029a ) or ( a3030a );
 a5044a <=( a3031a ) or ( a5043a );
 a5047a <=( a3027a ) or ( a3028a );
 a5050a <=( a3025a ) or ( a3026a );
 a5051a <=( a5050a ) or ( a5047a );
 a5052a <=( a5051a ) or ( a5044a );
 a5053a <=( a5052a ) or ( a5039a );
 a5057a <=( a3022a ) or ( a3023a );
 a5058a <=( a3024a ) or ( a5057a );
 a5061a <=( a3020a ) or ( a3021a );
 a5064a <=( a3018a ) or ( a3019a );
 a5065a <=( a5064a ) or ( a5061a );
 a5066a <=( a5065a ) or ( a5058a );
 a5069a <=( a3016a ) or ( a3017a );
 a5072a <=( a3014a ) or ( a3015a );
 a5073a <=( a5072a ) or ( a5069a );
 a5076a <=( a3012a ) or ( a3013a );
 a5079a <=( a3010a ) or ( a3011a );
 a5080a <=( a5079a ) or ( a5076a );
 a5081a <=( a5080a ) or ( a5073a );
 a5082a <=( a5081a ) or ( a5066a );
 a5083a <=( a5082a ) or ( a5053a );
 a5084a <=( a5083a ) or ( a5026a );
 a5085a <=( a5084a ) or ( a4969a );
 a5086a <=( a5085a ) or ( a4854a );
 a5090a <=( a3007a ) or ( a3008a );
 a5091a <=( a3009a ) or ( a5090a );
 a5094a <=( a3005a ) or ( a3006a );
 a5097a <=( a3003a ) or ( a3004a );
 a5098a <=( a5097a ) or ( a5094a );
 a5099a <=( a5098a ) or ( a5091a );
 a5103a <=( a3000a ) or ( a3001a );
 a5104a <=( a3002a ) or ( a5103a );
 a5107a <=( a2998a ) or ( a2999a );
 a5110a <=( a2996a ) or ( a2997a );
 a5111a <=( a5110a ) or ( a5107a );
 a5112a <=( a5111a ) or ( a5104a );
 a5113a <=( a5112a ) or ( a5099a );
 a5117a <=( a2993a ) or ( a2994a );
 a5118a <=( a2995a ) or ( a5117a );
 a5121a <=( a2991a ) or ( a2992a );
 a5124a <=( a2989a ) or ( a2990a );
 a5125a <=( a5124a ) or ( a5121a );
 a5126a <=( a5125a ) or ( a5118a );
 a5129a <=( a2987a ) or ( a2988a );
 a5132a <=( a2985a ) or ( a2986a );
 a5133a <=( a5132a ) or ( a5129a );
 a5136a <=( a2983a ) or ( a2984a );
 a5139a <=( a2981a ) or ( a2982a );
 a5140a <=( a5139a ) or ( a5136a );
 a5141a <=( a5140a ) or ( a5133a );
 a5142a <=( a5141a ) or ( a5126a );
 a5143a <=( a5142a ) or ( a5113a );
 a5147a <=( a2978a ) or ( a2979a );
 a5148a <=( a2980a ) or ( a5147a );
 a5151a <=( a2976a ) or ( a2977a );
 a5154a <=( a2974a ) or ( a2975a );
 a5155a <=( a5154a ) or ( a5151a );
 a5156a <=( a5155a ) or ( a5148a );
 a5160a <=( a2971a ) or ( a2972a );
 a5161a <=( a2973a ) or ( a5160a );
 a5164a <=( a2969a ) or ( a2970a );
 a5167a <=( a2967a ) or ( a2968a );
 a5168a <=( a5167a ) or ( a5164a );
 a5169a <=( a5168a ) or ( a5161a );
 a5170a <=( a5169a ) or ( a5156a );
 a5174a <=( a2964a ) or ( a2965a );
 a5175a <=( a2966a ) or ( a5174a );
 a5178a <=( a2962a ) or ( a2963a );
 a5181a <=( a2960a ) or ( a2961a );
 a5182a <=( a5181a ) or ( a5178a );
 a5183a <=( a5182a ) or ( a5175a );
 a5186a <=( a2958a ) or ( a2959a );
 a5189a <=( a2956a ) or ( a2957a );
 a5190a <=( a5189a ) or ( a5186a );
 a5193a <=( a2954a ) or ( a2955a );
 a5196a <=( a2952a ) or ( a2953a );
 a5197a <=( a5196a ) or ( a5193a );
 a5198a <=( a5197a ) or ( a5190a );
 a5199a <=( a5198a ) or ( a5183a );
 a5200a <=( a5199a ) or ( a5170a );
 a5201a <=( a5200a ) or ( a5143a );
 a5205a <=( a2949a ) or ( a2950a );
 a5206a <=( a2951a ) or ( a5205a );
 a5209a <=( a2947a ) or ( a2948a );
 a5212a <=( a2945a ) or ( a2946a );
 a5213a <=( a5212a ) or ( a5209a );
 a5214a <=( a5213a ) or ( a5206a );
 a5218a <=( a2942a ) or ( a2943a );
 a5219a <=( a2944a ) or ( a5218a );
 a5222a <=( a2940a ) or ( a2941a );
 a5225a <=( a2938a ) or ( a2939a );
 a5226a <=( a5225a ) or ( a5222a );
 a5227a <=( a5226a ) or ( a5219a );
 a5228a <=( a5227a ) or ( a5214a );
 a5232a <=( a2935a ) or ( a2936a );
 a5233a <=( a2937a ) or ( a5232a );
 a5236a <=( a2933a ) or ( a2934a );
 a5239a <=( a2931a ) or ( a2932a );
 a5240a <=( a5239a ) or ( a5236a );
 a5241a <=( a5240a ) or ( a5233a );
 a5244a <=( a2929a ) or ( a2930a );
 a5247a <=( a2927a ) or ( a2928a );
 a5248a <=( a5247a ) or ( a5244a );
 a5251a <=( a2925a ) or ( a2926a );
 a5254a <=( a2923a ) or ( a2924a );
 a5255a <=( a5254a ) or ( a5251a );
 a5256a <=( a5255a ) or ( a5248a );
 a5257a <=( a5256a ) or ( a5241a );
 a5258a <=( a5257a ) or ( a5228a );
 a5262a <=( a2920a ) or ( a2921a );
 a5263a <=( a2922a ) or ( a5262a );
 a5266a <=( a2918a ) or ( a2919a );
 a5269a <=( a2916a ) or ( a2917a );
 a5270a <=( a5269a ) or ( a5266a );
 a5271a <=( a5270a ) or ( a5263a );
 a5275a <=( a2913a ) or ( a2914a );
 a5276a <=( a2915a ) or ( a5275a );
 a5279a <=( a2911a ) or ( a2912a );
 a5282a <=( a2909a ) or ( a2910a );
 a5283a <=( a5282a ) or ( a5279a );
 a5284a <=( a5283a ) or ( a5276a );
 a5285a <=( a5284a ) or ( a5271a );
 a5289a <=( a2906a ) or ( a2907a );
 a5290a <=( a2908a ) or ( a5289a );
 a5293a <=( a2904a ) or ( a2905a );
 a5296a <=( a2902a ) or ( a2903a );
 a5297a <=( a5296a ) or ( a5293a );
 a5298a <=( a5297a ) or ( a5290a );
 a5301a <=( a2900a ) or ( a2901a );
 a5304a <=( a2898a ) or ( a2899a );
 a5305a <=( a5304a ) or ( a5301a );
 a5308a <=( a2896a ) or ( a2897a );
 a5311a <=( a2894a ) or ( a2895a );
 a5312a <=( a5311a ) or ( a5308a );
 a5313a <=( a5312a ) or ( a5305a );
 a5314a <=( a5313a ) or ( a5298a );
 a5315a <=( a5314a ) or ( a5285a );
 a5316a <=( a5315a ) or ( a5258a );
 a5317a <=( a5316a ) or ( a5201a );
 a5321a <=( a2891a ) or ( a2892a );
 a5322a <=( a2893a ) or ( a5321a );
 a5325a <=( a2889a ) or ( a2890a );
 a5328a <=( a2887a ) or ( a2888a );
 a5329a <=( a5328a ) or ( a5325a );
 a5330a <=( a5329a ) or ( a5322a );
 a5334a <=( a2884a ) or ( a2885a );
 a5335a <=( a2886a ) or ( a5334a );
 a5338a <=( a2882a ) or ( a2883a );
 a5341a <=( a2880a ) or ( a2881a );
 a5342a <=( a5341a ) or ( a5338a );
 a5343a <=( a5342a ) or ( a5335a );
 a5344a <=( a5343a ) or ( a5330a );
 a5348a <=( a2877a ) or ( a2878a );
 a5349a <=( a2879a ) or ( a5348a );
 a5352a <=( a2875a ) or ( a2876a );
 a5355a <=( a2873a ) or ( a2874a );
 a5356a <=( a5355a ) or ( a5352a );
 a5357a <=( a5356a ) or ( a5349a );
 a5360a <=( a2871a ) or ( a2872a );
 a5363a <=( a2869a ) or ( a2870a );
 a5364a <=( a5363a ) or ( a5360a );
 a5367a <=( a2867a ) or ( a2868a );
 a5370a <=( a2865a ) or ( a2866a );
 a5371a <=( a5370a ) or ( a5367a );
 a5372a <=( a5371a ) or ( a5364a );
 a5373a <=( a5372a ) or ( a5357a );
 a5374a <=( a5373a ) or ( a5344a );
 a5378a <=( a2862a ) or ( a2863a );
 a5379a <=( a2864a ) or ( a5378a );
 a5382a <=( a2860a ) or ( a2861a );
 a5385a <=( a2858a ) or ( a2859a );
 a5386a <=( a5385a ) or ( a5382a );
 a5387a <=( a5386a ) or ( a5379a );
 a5391a <=( a2855a ) or ( a2856a );
 a5392a <=( a2857a ) or ( a5391a );
 a5395a <=( a2853a ) or ( a2854a );
 a5398a <=( a2851a ) or ( a2852a );
 a5399a <=( a5398a ) or ( a5395a );
 a5400a <=( a5399a ) or ( a5392a );
 a5401a <=( a5400a ) or ( a5387a );
 a5405a <=( a2848a ) or ( a2849a );
 a5406a <=( a2850a ) or ( a5405a );
 a5409a <=( a2846a ) or ( a2847a );
 a5412a <=( a2844a ) or ( a2845a );
 a5413a <=( a5412a ) or ( a5409a );
 a5414a <=( a5413a ) or ( a5406a );
 a5417a <=( a2842a ) or ( a2843a );
 a5420a <=( a2840a ) or ( a2841a );
 a5421a <=( a5420a ) or ( a5417a );
 a5424a <=( a2838a ) or ( a2839a );
 a5427a <=( a2836a ) or ( a2837a );
 a5428a <=( a5427a ) or ( a5424a );
 a5429a <=( a5428a ) or ( a5421a );
 a5430a <=( a5429a ) or ( a5414a );
 a5431a <=( a5430a ) or ( a5401a );
 a5432a <=( a5431a ) or ( a5374a );
 a5436a <=( a2833a ) or ( a2834a );
 a5437a <=( a2835a ) or ( a5436a );
 a5440a <=( a2831a ) or ( a2832a );
 a5443a <=( a2829a ) or ( a2830a );
 a5444a <=( a5443a ) or ( a5440a );
 a5445a <=( a5444a ) or ( a5437a );
 a5449a <=( a2826a ) or ( a2827a );
 a5450a <=( a2828a ) or ( a5449a );
 a5453a <=( a2824a ) or ( a2825a );
 a5456a <=( a2822a ) or ( a2823a );
 a5457a <=( a5456a ) or ( a5453a );
 a5458a <=( a5457a ) or ( a5450a );
 a5459a <=( a5458a ) or ( a5445a );
 a5463a <=( a2819a ) or ( a2820a );
 a5464a <=( a2821a ) or ( a5463a );
 a5467a <=( a2817a ) or ( a2818a );
 a5470a <=( a2815a ) or ( a2816a );
 a5471a <=( a5470a ) or ( a5467a );
 a5472a <=( a5471a ) or ( a5464a );
 a5475a <=( a2813a ) or ( a2814a );
 a5478a <=( a2811a ) or ( a2812a );
 a5479a <=( a5478a ) or ( a5475a );
 a5482a <=( a2809a ) or ( a2810a );
 a5485a <=( a2807a ) or ( a2808a );
 a5486a <=( a5485a ) or ( a5482a );
 a5487a <=( a5486a ) or ( a5479a );
 a5488a <=( a5487a ) or ( a5472a );
 a5489a <=( a5488a ) or ( a5459a );
 a5493a <=( a2804a ) or ( a2805a );
 a5494a <=( a2806a ) or ( a5493a );
 a5497a <=( a2802a ) or ( a2803a );
 a5500a <=( a2800a ) or ( a2801a );
 a5501a <=( a5500a ) or ( a5497a );
 a5502a <=( a5501a ) or ( a5494a );
 a5506a <=( a2797a ) or ( a2798a );
 a5507a <=( a2799a ) or ( a5506a );
 a5510a <=( a2795a ) or ( a2796a );
 a5513a <=( a2793a ) or ( a2794a );
 a5514a <=( a5513a ) or ( a5510a );
 a5515a <=( a5514a ) or ( a5507a );
 a5516a <=( a5515a ) or ( a5502a );
 a5520a <=( a2790a ) or ( a2791a );
 a5521a <=( a2792a ) or ( a5520a );
 a5524a <=( a2788a ) or ( a2789a );
 a5527a <=( a2786a ) or ( a2787a );
 a5528a <=( a5527a ) or ( a5524a );
 a5529a <=( a5528a ) or ( a5521a );
 a5532a <=( a2784a ) or ( a2785a );
 a5535a <=( a2782a ) or ( a2783a );
 a5536a <=( a5535a ) or ( a5532a );
 a5539a <=( a2780a ) or ( a2781a );
 a5542a <=( a2778a ) or ( a2779a );
 a5543a <=( a5542a ) or ( a5539a );
 a5544a <=( a5543a ) or ( a5536a );
 a5545a <=( a5544a ) or ( a5529a );
 a5546a <=( a5545a ) or ( a5516a );
 a5547a <=( a5546a ) or ( a5489a );
 a5548a <=( a5547a ) or ( a5432a );
 a5549a <=( a5548a ) or ( a5317a );
 a5550a <=( a5549a ) or ( a5086a );
 a5551a <=( a5550a ) or ( a4625a );
 a5555a <=( a2775a ) or ( a2776a );
 a5556a <=( a2777a ) or ( a5555a );
 a5559a <=( a2773a ) or ( a2774a );
 a5562a <=( a2771a ) or ( a2772a );
 a5563a <=( a5562a ) or ( a5559a );
 a5564a <=( a5563a ) or ( a5556a );
 a5568a <=( a2768a ) or ( a2769a );
 a5569a <=( a2770a ) or ( a5568a );
 a5572a <=( a2766a ) or ( a2767a );
 a5575a <=( a2764a ) or ( a2765a );
 a5576a <=( a5575a ) or ( a5572a );
 a5577a <=( a5576a ) or ( a5569a );
 a5578a <=( a5577a ) or ( a5564a );
 a5582a <=( a2761a ) or ( a2762a );
 a5583a <=( a2763a ) or ( a5582a );
 a5586a <=( a2759a ) or ( a2760a );
 a5589a <=( a2757a ) or ( a2758a );
 a5590a <=( a5589a ) or ( a5586a );
 a5591a <=( a5590a ) or ( a5583a );
 a5595a <=( a2754a ) or ( a2755a );
 a5596a <=( a2756a ) or ( a5595a );
 a5599a <=( a2752a ) or ( a2753a );
 a5602a <=( a2750a ) or ( a2751a );
 a5603a <=( a5602a ) or ( a5599a );
 a5604a <=( a5603a ) or ( a5596a );
 a5605a <=( a5604a ) or ( a5591a );
 a5606a <=( a5605a ) or ( a5578a );
 a5610a <=( a2747a ) or ( a2748a );
 a5611a <=( a2749a ) or ( a5610a );
 a5614a <=( a2745a ) or ( a2746a );
 a5617a <=( a2743a ) or ( a2744a );
 a5618a <=( a5617a ) or ( a5614a );
 a5619a <=( a5618a ) or ( a5611a );
 a5623a <=( a2740a ) or ( a2741a );
 a5624a <=( a2742a ) or ( a5623a );
 a5627a <=( a2738a ) or ( a2739a );
 a5630a <=( a2736a ) or ( a2737a );
 a5631a <=( a5630a ) or ( a5627a );
 a5632a <=( a5631a ) or ( a5624a );
 a5633a <=( a5632a ) or ( a5619a );
 a5637a <=( a2733a ) or ( a2734a );
 a5638a <=( a2735a ) or ( a5637a );
 a5641a <=( a2731a ) or ( a2732a );
 a5644a <=( a2729a ) or ( a2730a );
 a5645a <=( a5644a ) or ( a5641a );
 a5646a <=( a5645a ) or ( a5638a );
 a5649a <=( a2727a ) or ( a2728a );
 a5652a <=( a2725a ) or ( a2726a );
 a5653a <=( a5652a ) or ( a5649a );
 a5656a <=( a2723a ) or ( a2724a );
 a5659a <=( a2721a ) or ( a2722a );
 a5660a <=( a5659a ) or ( a5656a );
 a5661a <=( a5660a ) or ( a5653a );
 a5662a <=( a5661a ) or ( a5646a );
 a5663a <=( a5662a ) or ( a5633a );
 a5664a <=( a5663a ) or ( a5606a );
 a5668a <=( a2718a ) or ( a2719a );
 a5669a <=( a2720a ) or ( a5668a );
 a5672a <=( a2716a ) or ( a2717a );
 a5675a <=( a2714a ) or ( a2715a );
 a5676a <=( a5675a ) or ( a5672a );
 a5677a <=( a5676a ) or ( a5669a );
 a5681a <=( a2711a ) or ( a2712a );
 a5682a <=( a2713a ) or ( a5681a );
 a5685a <=( a2709a ) or ( a2710a );
 a5688a <=( a2707a ) or ( a2708a );
 a5689a <=( a5688a ) or ( a5685a );
 a5690a <=( a5689a ) or ( a5682a );
 a5691a <=( a5690a ) or ( a5677a );
 a5695a <=( a2704a ) or ( a2705a );
 a5696a <=( a2706a ) or ( a5695a );
 a5699a <=( a2702a ) or ( a2703a );
 a5702a <=( a2700a ) or ( a2701a );
 a5703a <=( a5702a ) or ( a5699a );
 a5704a <=( a5703a ) or ( a5696a );
 a5707a <=( a2698a ) or ( a2699a );
 a5710a <=( a2696a ) or ( a2697a );
 a5711a <=( a5710a ) or ( a5707a );
 a5714a <=( a2694a ) or ( a2695a );
 a5717a <=( a2692a ) or ( a2693a );
 a5718a <=( a5717a ) or ( a5714a );
 a5719a <=( a5718a ) or ( a5711a );
 a5720a <=( a5719a ) or ( a5704a );
 a5721a <=( a5720a ) or ( a5691a );
 a5725a <=( a2689a ) or ( a2690a );
 a5726a <=( a2691a ) or ( a5725a );
 a5729a <=( a2687a ) or ( a2688a );
 a5732a <=( a2685a ) or ( a2686a );
 a5733a <=( a5732a ) or ( a5729a );
 a5734a <=( a5733a ) or ( a5726a );
 a5738a <=( a2682a ) or ( a2683a );
 a5739a <=( a2684a ) or ( a5738a );
 a5742a <=( a2680a ) or ( a2681a );
 a5745a <=( a2678a ) or ( a2679a );
 a5746a <=( a5745a ) or ( a5742a );
 a5747a <=( a5746a ) or ( a5739a );
 a5748a <=( a5747a ) or ( a5734a );
 a5752a <=( a2675a ) or ( a2676a );
 a5753a <=( a2677a ) or ( a5752a );
 a5756a <=( a2673a ) or ( a2674a );
 a5759a <=( a2671a ) or ( a2672a );
 a5760a <=( a5759a ) or ( a5756a );
 a5761a <=( a5760a ) or ( a5753a );
 a5764a <=( a2669a ) or ( a2670a );
 a5767a <=( a2667a ) or ( a2668a );
 a5768a <=( a5767a ) or ( a5764a );
 a5771a <=( a2665a ) or ( a2666a );
 a5774a <=( a2663a ) or ( a2664a );
 a5775a <=( a5774a ) or ( a5771a );
 a5776a <=( a5775a ) or ( a5768a );
 a5777a <=( a5776a ) or ( a5761a );
 a5778a <=( a5777a ) or ( a5748a );
 a5779a <=( a5778a ) or ( a5721a );
 a5780a <=( a5779a ) or ( a5664a );
 a5784a <=( a2660a ) or ( a2661a );
 a5785a <=( a2662a ) or ( a5784a );
 a5788a <=( a2658a ) or ( a2659a );
 a5791a <=( a2656a ) or ( a2657a );
 a5792a <=( a5791a ) or ( a5788a );
 a5793a <=( a5792a ) or ( a5785a );
 a5797a <=( a2653a ) or ( a2654a );
 a5798a <=( a2655a ) or ( a5797a );
 a5801a <=( a2651a ) or ( a2652a );
 a5804a <=( a2649a ) or ( a2650a );
 a5805a <=( a5804a ) or ( a5801a );
 a5806a <=( a5805a ) or ( a5798a );
 a5807a <=( a5806a ) or ( a5793a );
 a5811a <=( a2646a ) or ( a2647a );
 a5812a <=( a2648a ) or ( a5811a );
 a5815a <=( a2644a ) or ( a2645a );
 a5818a <=( a2642a ) or ( a2643a );
 a5819a <=( a5818a ) or ( a5815a );
 a5820a <=( a5819a ) or ( a5812a );
 a5823a <=( a2640a ) or ( a2641a );
 a5826a <=( a2638a ) or ( a2639a );
 a5827a <=( a5826a ) or ( a5823a );
 a5830a <=( a2636a ) or ( a2637a );
 a5833a <=( a2634a ) or ( a2635a );
 a5834a <=( a5833a ) or ( a5830a );
 a5835a <=( a5834a ) or ( a5827a );
 a5836a <=( a5835a ) or ( a5820a );
 a5837a <=( a5836a ) or ( a5807a );
 a5841a <=( a2631a ) or ( a2632a );
 a5842a <=( a2633a ) or ( a5841a );
 a5845a <=( a2629a ) or ( a2630a );
 a5848a <=( a2627a ) or ( a2628a );
 a5849a <=( a5848a ) or ( a5845a );
 a5850a <=( a5849a ) or ( a5842a );
 a5854a <=( a2624a ) or ( a2625a );
 a5855a <=( a2626a ) or ( a5854a );
 a5858a <=( a2622a ) or ( a2623a );
 a5861a <=( a2620a ) or ( a2621a );
 a5862a <=( a5861a ) or ( a5858a );
 a5863a <=( a5862a ) or ( a5855a );
 a5864a <=( a5863a ) or ( a5850a );
 a5868a <=( a2617a ) or ( a2618a );
 a5869a <=( a2619a ) or ( a5868a );
 a5872a <=( a2615a ) or ( a2616a );
 a5875a <=( a2613a ) or ( a2614a );
 a5876a <=( a5875a ) or ( a5872a );
 a5877a <=( a5876a ) or ( a5869a );
 a5880a <=( a2611a ) or ( a2612a );
 a5883a <=( a2609a ) or ( a2610a );
 a5884a <=( a5883a ) or ( a5880a );
 a5887a <=( a2607a ) or ( a2608a );
 a5890a <=( a2605a ) or ( a2606a );
 a5891a <=( a5890a ) or ( a5887a );
 a5892a <=( a5891a ) or ( a5884a );
 a5893a <=( a5892a ) or ( a5877a );
 a5894a <=( a5893a ) or ( a5864a );
 a5895a <=( a5894a ) or ( a5837a );
 a5899a <=( a2602a ) or ( a2603a );
 a5900a <=( a2604a ) or ( a5899a );
 a5903a <=( a2600a ) or ( a2601a );
 a5906a <=( a2598a ) or ( a2599a );
 a5907a <=( a5906a ) or ( a5903a );
 a5908a <=( a5907a ) or ( a5900a );
 a5912a <=( a2595a ) or ( a2596a );
 a5913a <=( a2597a ) or ( a5912a );
 a5916a <=( a2593a ) or ( a2594a );
 a5919a <=( a2591a ) or ( a2592a );
 a5920a <=( a5919a ) or ( a5916a );
 a5921a <=( a5920a ) or ( a5913a );
 a5922a <=( a5921a ) or ( a5908a );
 a5926a <=( a2588a ) or ( a2589a );
 a5927a <=( a2590a ) or ( a5926a );
 a5930a <=( a2586a ) or ( a2587a );
 a5933a <=( a2584a ) or ( a2585a );
 a5934a <=( a5933a ) or ( a5930a );
 a5935a <=( a5934a ) or ( a5927a );
 a5938a <=( a2582a ) or ( a2583a );
 a5941a <=( a2580a ) or ( a2581a );
 a5942a <=( a5941a ) or ( a5938a );
 a5945a <=( a2578a ) or ( a2579a );
 a5948a <=( a2576a ) or ( a2577a );
 a5949a <=( a5948a ) or ( a5945a );
 a5950a <=( a5949a ) or ( a5942a );
 a5951a <=( a5950a ) or ( a5935a );
 a5952a <=( a5951a ) or ( a5922a );
 a5956a <=( a2573a ) or ( a2574a );
 a5957a <=( a2575a ) or ( a5956a );
 a5960a <=( a2571a ) or ( a2572a );
 a5963a <=( a2569a ) or ( a2570a );
 a5964a <=( a5963a ) or ( a5960a );
 a5965a <=( a5964a ) or ( a5957a );
 a5969a <=( a2566a ) or ( a2567a );
 a5970a <=( a2568a ) or ( a5969a );
 a5973a <=( a2564a ) or ( a2565a );
 a5976a <=( a2562a ) or ( a2563a );
 a5977a <=( a5976a ) or ( a5973a );
 a5978a <=( a5977a ) or ( a5970a );
 a5979a <=( a5978a ) or ( a5965a );
 a5983a <=( a2559a ) or ( a2560a );
 a5984a <=( a2561a ) or ( a5983a );
 a5987a <=( a2557a ) or ( a2558a );
 a5990a <=( a2555a ) or ( a2556a );
 a5991a <=( a5990a ) or ( a5987a );
 a5992a <=( a5991a ) or ( a5984a );
 a5995a <=( a2553a ) or ( a2554a );
 a5998a <=( a2551a ) or ( a2552a );
 a5999a <=( a5998a ) or ( a5995a );
 a6002a <=( a2549a ) or ( a2550a );
 a6005a <=( a2547a ) or ( a2548a );
 a6006a <=( a6005a ) or ( a6002a );
 a6007a <=( a6006a ) or ( a5999a );
 a6008a <=( a6007a ) or ( a5992a );
 a6009a <=( a6008a ) or ( a5979a );
 a6010a <=( a6009a ) or ( a5952a );
 a6011a <=( a6010a ) or ( a5895a );
 a6012a <=( a6011a ) or ( a5780a );
 a6016a <=( a2544a ) or ( a2545a );
 a6017a <=( a2546a ) or ( a6016a );
 a6020a <=( a2542a ) or ( a2543a );
 a6023a <=( a2540a ) or ( a2541a );
 a6024a <=( a6023a ) or ( a6020a );
 a6025a <=( a6024a ) or ( a6017a );
 a6029a <=( a2537a ) or ( a2538a );
 a6030a <=( a2539a ) or ( a6029a );
 a6033a <=( a2535a ) or ( a2536a );
 a6036a <=( a2533a ) or ( a2534a );
 a6037a <=( a6036a ) or ( a6033a );
 a6038a <=( a6037a ) or ( a6030a );
 a6039a <=( a6038a ) or ( a6025a );
 a6043a <=( a2530a ) or ( a2531a );
 a6044a <=( a2532a ) or ( a6043a );
 a6047a <=( a2528a ) or ( a2529a );
 a6050a <=( a2526a ) or ( a2527a );
 a6051a <=( a6050a ) or ( a6047a );
 a6052a <=( a6051a ) or ( a6044a );
 a6055a <=( a2524a ) or ( a2525a );
 a6058a <=( a2522a ) or ( a2523a );
 a6059a <=( a6058a ) or ( a6055a );
 a6062a <=( a2520a ) or ( a2521a );
 a6065a <=( a2518a ) or ( a2519a );
 a6066a <=( a6065a ) or ( a6062a );
 a6067a <=( a6066a ) or ( a6059a );
 a6068a <=( a6067a ) or ( a6052a );
 a6069a <=( a6068a ) or ( a6039a );
 a6073a <=( a2515a ) or ( a2516a );
 a6074a <=( a2517a ) or ( a6073a );
 a6077a <=( a2513a ) or ( a2514a );
 a6080a <=( a2511a ) or ( a2512a );
 a6081a <=( a6080a ) or ( a6077a );
 a6082a <=( a6081a ) or ( a6074a );
 a6086a <=( a2508a ) or ( a2509a );
 a6087a <=( a2510a ) or ( a6086a );
 a6090a <=( a2506a ) or ( a2507a );
 a6093a <=( a2504a ) or ( a2505a );
 a6094a <=( a6093a ) or ( a6090a );
 a6095a <=( a6094a ) or ( a6087a );
 a6096a <=( a6095a ) or ( a6082a );
 a6100a <=( a2501a ) or ( a2502a );
 a6101a <=( a2503a ) or ( a6100a );
 a6104a <=( a2499a ) or ( a2500a );
 a6107a <=( a2497a ) or ( a2498a );
 a6108a <=( a6107a ) or ( a6104a );
 a6109a <=( a6108a ) or ( a6101a );
 a6112a <=( a2495a ) or ( a2496a );
 a6115a <=( a2493a ) or ( a2494a );
 a6116a <=( a6115a ) or ( a6112a );
 a6119a <=( a2491a ) or ( a2492a );
 a6122a <=( a2489a ) or ( a2490a );
 a6123a <=( a6122a ) or ( a6119a );
 a6124a <=( a6123a ) or ( a6116a );
 a6125a <=( a6124a ) or ( a6109a );
 a6126a <=( a6125a ) or ( a6096a );
 a6127a <=( a6126a ) or ( a6069a );
 a6131a <=( a2486a ) or ( a2487a );
 a6132a <=( a2488a ) or ( a6131a );
 a6135a <=( a2484a ) or ( a2485a );
 a6138a <=( a2482a ) or ( a2483a );
 a6139a <=( a6138a ) or ( a6135a );
 a6140a <=( a6139a ) or ( a6132a );
 a6144a <=( a2479a ) or ( a2480a );
 a6145a <=( a2481a ) or ( a6144a );
 a6148a <=( a2477a ) or ( a2478a );
 a6151a <=( a2475a ) or ( a2476a );
 a6152a <=( a6151a ) or ( a6148a );
 a6153a <=( a6152a ) or ( a6145a );
 a6154a <=( a6153a ) or ( a6140a );
 a6158a <=( a2472a ) or ( a2473a );
 a6159a <=( a2474a ) or ( a6158a );
 a6162a <=( a2470a ) or ( a2471a );
 a6165a <=( a2468a ) or ( a2469a );
 a6166a <=( a6165a ) or ( a6162a );
 a6167a <=( a6166a ) or ( a6159a );
 a6170a <=( a2466a ) or ( a2467a );
 a6173a <=( a2464a ) or ( a2465a );
 a6174a <=( a6173a ) or ( a6170a );
 a6177a <=( a2462a ) or ( a2463a );
 a6180a <=( a2460a ) or ( a2461a );
 a6181a <=( a6180a ) or ( a6177a );
 a6182a <=( a6181a ) or ( a6174a );
 a6183a <=( a6182a ) or ( a6167a );
 a6184a <=( a6183a ) or ( a6154a );
 a6188a <=( a2457a ) or ( a2458a );
 a6189a <=( a2459a ) or ( a6188a );
 a6192a <=( a2455a ) or ( a2456a );
 a6195a <=( a2453a ) or ( a2454a );
 a6196a <=( a6195a ) or ( a6192a );
 a6197a <=( a6196a ) or ( a6189a );
 a6201a <=( a2450a ) or ( a2451a );
 a6202a <=( a2452a ) or ( a6201a );
 a6205a <=( a2448a ) or ( a2449a );
 a6208a <=( a2446a ) or ( a2447a );
 a6209a <=( a6208a ) or ( a6205a );
 a6210a <=( a6209a ) or ( a6202a );
 a6211a <=( a6210a ) or ( a6197a );
 a6215a <=( a2443a ) or ( a2444a );
 a6216a <=( a2445a ) or ( a6215a );
 a6219a <=( a2441a ) or ( a2442a );
 a6222a <=( a2439a ) or ( a2440a );
 a6223a <=( a6222a ) or ( a6219a );
 a6224a <=( a6223a ) or ( a6216a );
 a6227a <=( a2437a ) or ( a2438a );
 a6230a <=( a2435a ) or ( a2436a );
 a6231a <=( a6230a ) or ( a6227a );
 a6234a <=( a2433a ) or ( a2434a );
 a6237a <=( a2431a ) or ( a2432a );
 a6238a <=( a6237a ) or ( a6234a );
 a6239a <=( a6238a ) or ( a6231a );
 a6240a <=( a6239a ) or ( a6224a );
 a6241a <=( a6240a ) or ( a6211a );
 a6242a <=( a6241a ) or ( a6184a );
 a6243a <=( a6242a ) or ( a6127a );
 a6247a <=( a2428a ) or ( a2429a );
 a6248a <=( a2430a ) or ( a6247a );
 a6251a <=( a2426a ) or ( a2427a );
 a6254a <=( a2424a ) or ( a2425a );
 a6255a <=( a6254a ) or ( a6251a );
 a6256a <=( a6255a ) or ( a6248a );
 a6260a <=( a2421a ) or ( a2422a );
 a6261a <=( a2423a ) or ( a6260a );
 a6264a <=( a2419a ) or ( a2420a );
 a6267a <=( a2417a ) or ( a2418a );
 a6268a <=( a6267a ) or ( a6264a );
 a6269a <=( a6268a ) or ( a6261a );
 a6270a <=( a6269a ) or ( a6256a );
 a6274a <=( a2414a ) or ( a2415a );
 a6275a <=( a2416a ) or ( a6274a );
 a6278a <=( a2412a ) or ( a2413a );
 a6281a <=( a2410a ) or ( a2411a );
 a6282a <=( a6281a ) or ( a6278a );
 a6283a <=( a6282a ) or ( a6275a );
 a6286a <=( a2408a ) or ( a2409a );
 a6289a <=( a2406a ) or ( a2407a );
 a6290a <=( a6289a ) or ( a6286a );
 a6293a <=( a2404a ) or ( a2405a );
 a6296a <=( a2402a ) or ( a2403a );
 a6297a <=( a6296a ) or ( a6293a );
 a6298a <=( a6297a ) or ( a6290a );
 a6299a <=( a6298a ) or ( a6283a );
 a6300a <=( a6299a ) or ( a6270a );
 a6304a <=( a2399a ) or ( a2400a );
 a6305a <=( a2401a ) or ( a6304a );
 a6308a <=( a2397a ) or ( a2398a );
 a6311a <=( a2395a ) or ( a2396a );
 a6312a <=( a6311a ) or ( a6308a );
 a6313a <=( a6312a ) or ( a6305a );
 a6317a <=( a2392a ) or ( a2393a );
 a6318a <=( a2394a ) or ( a6317a );
 a6321a <=( a2390a ) or ( a2391a );
 a6324a <=( a2388a ) or ( a2389a );
 a6325a <=( a6324a ) or ( a6321a );
 a6326a <=( a6325a ) or ( a6318a );
 a6327a <=( a6326a ) or ( a6313a );
 a6331a <=( a2385a ) or ( a2386a );
 a6332a <=( a2387a ) or ( a6331a );
 a6335a <=( a2383a ) or ( a2384a );
 a6338a <=( a2381a ) or ( a2382a );
 a6339a <=( a6338a ) or ( a6335a );
 a6340a <=( a6339a ) or ( a6332a );
 a6343a <=( a2379a ) or ( a2380a );
 a6346a <=( a2377a ) or ( a2378a );
 a6347a <=( a6346a ) or ( a6343a );
 a6350a <=( a2375a ) or ( a2376a );
 a6353a <=( a2373a ) or ( a2374a );
 a6354a <=( a6353a ) or ( a6350a );
 a6355a <=( a6354a ) or ( a6347a );
 a6356a <=( a6355a ) or ( a6340a );
 a6357a <=( a6356a ) or ( a6327a );
 a6358a <=( a6357a ) or ( a6300a );
 a6362a <=( a2370a ) or ( a2371a );
 a6363a <=( a2372a ) or ( a6362a );
 a6366a <=( a2368a ) or ( a2369a );
 a6369a <=( a2366a ) or ( a2367a );
 a6370a <=( a6369a ) or ( a6366a );
 a6371a <=( a6370a ) or ( a6363a );
 a6375a <=( a2363a ) or ( a2364a );
 a6376a <=( a2365a ) or ( a6375a );
 a6379a <=( a2361a ) or ( a2362a );
 a6382a <=( a2359a ) or ( a2360a );
 a6383a <=( a6382a ) or ( a6379a );
 a6384a <=( a6383a ) or ( a6376a );
 a6385a <=( a6384a ) or ( a6371a );
 a6389a <=( a2356a ) or ( a2357a );
 a6390a <=( a2358a ) or ( a6389a );
 a6393a <=( a2354a ) or ( a2355a );
 a6396a <=( a2352a ) or ( a2353a );
 a6397a <=( a6396a ) or ( a6393a );
 a6398a <=( a6397a ) or ( a6390a );
 a6401a <=( a2350a ) or ( a2351a );
 a6404a <=( a2348a ) or ( a2349a );
 a6405a <=( a6404a ) or ( a6401a );
 a6408a <=( a2346a ) or ( a2347a );
 a6411a <=( a2344a ) or ( a2345a );
 a6412a <=( a6411a ) or ( a6408a );
 a6413a <=( a6412a ) or ( a6405a );
 a6414a <=( a6413a ) or ( a6398a );
 a6415a <=( a6414a ) or ( a6385a );
 a6419a <=( a2341a ) or ( a2342a );
 a6420a <=( a2343a ) or ( a6419a );
 a6423a <=( a2339a ) or ( a2340a );
 a6426a <=( a2337a ) or ( a2338a );
 a6427a <=( a6426a ) or ( a6423a );
 a6428a <=( a6427a ) or ( a6420a );
 a6432a <=( a2334a ) or ( a2335a );
 a6433a <=( a2336a ) or ( a6432a );
 a6436a <=( a2332a ) or ( a2333a );
 a6439a <=( a2330a ) or ( a2331a );
 a6440a <=( a6439a ) or ( a6436a );
 a6441a <=( a6440a ) or ( a6433a );
 a6442a <=( a6441a ) or ( a6428a );
 a6446a <=( a2327a ) or ( a2328a );
 a6447a <=( a2329a ) or ( a6446a );
 a6450a <=( a2325a ) or ( a2326a );
 a6453a <=( a2323a ) or ( a2324a );
 a6454a <=( a6453a ) or ( a6450a );
 a6455a <=( a6454a ) or ( a6447a );
 a6458a <=( a2321a ) or ( a2322a );
 a6461a <=( a2319a ) or ( a2320a );
 a6462a <=( a6461a ) or ( a6458a );
 a6465a <=( a2317a ) or ( a2318a );
 a6468a <=( a2315a ) or ( a2316a );
 a6469a <=( a6468a ) or ( a6465a );
 a6470a <=( a6469a ) or ( a6462a );
 a6471a <=( a6470a ) or ( a6455a );
 a6472a <=( a6471a ) or ( a6442a );
 a6473a <=( a6472a ) or ( a6415a );
 a6474a <=( a6473a ) or ( a6358a );
 a6475a <=( a6474a ) or ( a6243a );
 a6476a <=( a6475a ) or ( a6012a );
 a6480a <=( a2312a ) or ( a2313a );
 a6481a <=( a2314a ) or ( a6480a );
 a6484a <=( a2310a ) or ( a2311a );
 a6487a <=( a2308a ) or ( a2309a );
 a6488a <=( a6487a ) or ( a6484a );
 a6489a <=( a6488a ) or ( a6481a );
 a6493a <=( a2305a ) or ( a2306a );
 a6494a <=( a2307a ) or ( a6493a );
 a6497a <=( a2303a ) or ( a2304a );
 a6500a <=( a2301a ) or ( a2302a );
 a6501a <=( a6500a ) or ( a6497a );
 a6502a <=( a6501a ) or ( a6494a );
 a6503a <=( a6502a ) or ( a6489a );
 a6507a <=( a2298a ) or ( a2299a );
 a6508a <=( a2300a ) or ( a6507a );
 a6511a <=( a2296a ) or ( a2297a );
 a6514a <=( a2294a ) or ( a2295a );
 a6515a <=( a6514a ) or ( a6511a );
 a6516a <=( a6515a ) or ( a6508a );
 a6520a <=( a2291a ) or ( a2292a );
 a6521a <=( a2293a ) or ( a6520a );
 a6524a <=( a2289a ) or ( a2290a );
 a6527a <=( a2287a ) or ( a2288a );
 a6528a <=( a6527a ) or ( a6524a );
 a6529a <=( a6528a ) or ( a6521a );
 a6530a <=( a6529a ) or ( a6516a );
 a6531a <=( a6530a ) or ( a6503a );
 a6535a <=( a2284a ) or ( a2285a );
 a6536a <=( a2286a ) or ( a6535a );
 a6539a <=( a2282a ) or ( a2283a );
 a6542a <=( a2280a ) or ( a2281a );
 a6543a <=( a6542a ) or ( a6539a );
 a6544a <=( a6543a ) or ( a6536a );
 a6548a <=( a2277a ) or ( a2278a );
 a6549a <=( a2279a ) or ( a6548a );
 a6552a <=( a2275a ) or ( a2276a );
 a6555a <=( a2273a ) or ( a2274a );
 a6556a <=( a6555a ) or ( a6552a );
 a6557a <=( a6556a ) or ( a6549a );
 a6558a <=( a6557a ) or ( a6544a );
 a6562a <=( a2270a ) or ( a2271a );
 a6563a <=( a2272a ) or ( a6562a );
 a6566a <=( a2268a ) or ( a2269a );
 a6569a <=( a2266a ) or ( a2267a );
 a6570a <=( a6569a ) or ( a6566a );
 a6571a <=( a6570a ) or ( a6563a );
 a6574a <=( a2264a ) or ( a2265a );
 a6577a <=( a2262a ) or ( a2263a );
 a6578a <=( a6577a ) or ( a6574a );
 a6581a <=( a2260a ) or ( a2261a );
 a6584a <=( a2258a ) or ( a2259a );
 a6585a <=( a6584a ) or ( a6581a );
 a6586a <=( a6585a ) or ( a6578a );
 a6587a <=( a6586a ) or ( a6571a );
 a6588a <=( a6587a ) or ( a6558a );
 a6589a <=( a6588a ) or ( a6531a );
 a6593a <=( a2255a ) or ( a2256a );
 a6594a <=( a2257a ) or ( a6593a );
 a6597a <=( a2253a ) or ( a2254a );
 a6600a <=( a2251a ) or ( a2252a );
 a6601a <=( a6600a ) or ( a6597a );
 a6602a <=( a6601a ) or ( a6594a );
 a6606a <=( a2248a ) or ( a2249a );
 a6607a <=( a2250a ) or ( a6606a );
 a6610a <=( a2246a ) or ( a2247a );
 a6613a <=( a2244a ) or ( a2245a );
 a6614a <=( a6613a ) or ( a6610a );
 a6615a <=( a6614a ) or ( a6607a );
 a6616a <=( a6615a ) or ( a6602a );
 a6620a <=( a2241a ) or ( a2242a );
 a6621a <=( a2243a ) or ( a6620a );
 a6624a <=( a2239a ) or ( a2240a );
 a6627a <=( a2237a ) or ( a2238a );
 a6628a <=( a6627a ) or ( a6624a );
 a6629a <=( a6628a ) or ( a6621a );
 a6632a <=( a2235a ) or ( a2236a );
 a6635a <=( a2233a ) or ( a2234a );
 a6636a <=( a6635a ) or ( a6632a );
 a6639a <=( a2231a ) or ( a2232a );
 a6642a <=( a2229a ) or ( a2230a );
 a6643a <=( a6642a ) or ( a6639a );
 a6644a <=( a6643a ) or ( a6636a );
 a6645a <=( a6644a ) or ( a6629a );
 a6646a <=( a6645a ) or ( a6616a );
 a6650a <=( a2226a ) or ( a2227a );
 a6651a <=( a2228a ) or ( a6650a );
 a6654a <=( a2224a ) or ( a2225a );
 a6657a <=( a2222a ) or ( a2223a );
 a6658a <=( a6657a ) or ( a6654a );
 a6659a <=( a6658a ) or ( a6651a );
 a6663a <=( a2219a ) or ( a2220a );
 a6664a <=( a2221a ) or ( a6663a );
 a6667a <=( a2217a ) or ( a2218a );
 a6670a <=( a2215a ) or ( a2216a );
 a6671a <=( a6670a ) or ( a6667a );
 a6672a <=( a6671a ) or ( a6664a );
 a6673a <=( a6672a ) or ( a6659a );
 a6677a <=( a2212a ) or ( a2213a );
 a6678a <=( a2214a ) or ( a6677a );
 a6681a <=( a2210a ) or ( a2211a );
 a6684a <=( a2208a ) or ( a2209a );
 a6685a <=( a6684a ) or ( a6681a );
 a6686a <=( a6685a ) or ( a6678a );
 a6689a <=( a2206a ) or ( a2207a );
 a6692a <=( a2204a ) or ( a2205a );
 a6693a <=( a6692a ) or ( a6689a );
 a6696a <=( a2202a ) or ( a2203a );
 a6699a <=( a2200a ) or ( a2201a );
 a6700a <=( a6699a ) or ( a6696a );
 a6701a <=( a6700a ) or ( a6693a );
 a6702a <=( a6701a ) or ( a6686a );
 a6703a <=( a6702a ) or ( a6673a );
 a6704a <=( a6703a ) or ( a6646a );
 a6705a <=( a6704a ) or ( a6589a );
 a6709a <=( a2197a ) or ( a2198a );
 a6710a <=( a2199a ) or ( a6709a );
 a6713a <=( a2195a ) or ( a2196a );
 a6716a <=( a2193a ) or ( a2194a );
 a6717a <=( a6716a ) or ( a6713a );
 a6718a <=( a6717a ) or ( a6710a );
 a6722a <=( a2190a ) or ( a2191a );
 a6723a <=( a2192a ) or ( a6722a );
 a6726a <=( a2188a ) or ( a2189a );
 a6729a <=( a2186a ) or ( a2187a );
 a6730a <=( a6729a ) or ( a6726a );
 a6731a <=( a6730a ) or ( a6723a );
 a6732a <=( a6731a ) or ( a6718a );
 a6736a <=( a2183a ) or ( a2184a );
 a6737a <=( a2185a ) or ( a6736a );
 a6740a <=( a2181a ) or ( a2182a );
 a6743a <=( a2179a ) or ( a2180a );
 a6744a <=( a6743a ) or ( a6740a );
 a6745a <=( a6744a ) or ( a6737a );
 a6748a <=( a2177a ) or ( a2178a );
 a6751a <=( a2175a ) or ( a2176a );
 a6752a <=( a6751a ) or ( a6748a );
 a6755a <=( a2173a ) or ( a2174a );
 a6758a <=( a2171a ) or ( a2172a );
 a6759a <=( a6758a ) or ( a6755a );
 a6760a <=( a6759a ) or ( a6752a );
 a6761a <=( a6760a ) or ( a6745a );
 a6762a <=( a6761a ) or ( a6732a );
 a6766a <=( a2168a ) or ( a2169a );
 a6767a <=( a2170a ) or ( a6766a );
 a6770a <=( a2166a ) or ( a2167a );
 a6773a <=( a2164a ) or ( a2165a );
 a6774a <=( a6773a ) or ( a6770a );
 a6775a <=( a6774a ) or ( a6767a );
 a6779a <=( a2161a ) or ( a2162a );
 a6780a <=( a2163a ) or ( a6779a );
 a6783a <=( a2159a ) or ( a2160a );
 a6786a <=( a2157a ) or ( a2158a );
 a6787a <=( a6786a ) or ( a6783a );
 a6788a <=( a6787a ) or ( a6780a );
 a6789a <=( a6788a ) or ( a6775a );
 a6793a <=( a2154a ) or ( a2155a );
 a6794a <=( a2156a ) or ( a6793a );
 a6797a <=( a2152a ) or ( a2153a );
 a6800a <=( a2150a ) or ( a2151a );
 a6801a <=( a6800a ) or ( a6797a );
 a6802a <=( a6801a ) or ( a6794a );
 a6805a <=( a2148a ) or ( a2149a );
 a6808a <=( a2146a ) or ( a2147a );
 a6809a <=( a6808a ) or ( a6805a );
 a6812a <=( a2144a ) or ( a2145a );
 a6815a <=( a2142a ) or ( a2143a );
 a6816a <=( a6815a ) or ( a6812a );
 a6817a <=( a6816a ) or ( a6809a );
 a6818a <=( a6817a ) or ( a6802a );
 a6819a <=( a6818a ) or ( a6789a );
 a6820a <=( a6819a ) or ( a6762a );
 a6824a <=( a2139a ) or ( a2140a );
 a6825a <=( a2141a ) or ( a6824a );
 a6828a <=( a2137a ) or ( a2138a );
 a6831a <=( a2135a ) or ( a2136a );
 a6832a <=( a6831a ) or ( a6828a );
 a6833a <=( a6832a ) or ( a6825a );
 a6837a <=( a2132a ) or ( a2133a );
 a6838a <=( a2134a ) or ( a6837a );
 a6841a <=( a2130a ) or ( a2131a );
 a6844a <=( a2128a ) or ( a2129a );
 a6845a <=( a6844a ) or ( a6841a );
 a6846a <=( a6845a ) or ( a6838a );
 a6847a <=( a6846a ) or ( a6833a );
 a6851a <=( a2125a ) or ( a2126a );
 a6852a <=( a2127a ) or ( a6851a );
 a6855a <=( a2123a ) or ( a2124a );
 a6858a <=( a2121a ) or ( a2122a );
 a6859a <=( a6858a ) or ( a6855a );
 a6860a <=( a6859a ) or ( a6852a );
 a6863a <=( a2119a ) or ( a2120a );
 a6866a <=( a2117a ) or ( a2118a );
 a6867a <=( a6866a ) or ( a6863a );
 a6870a <=( a2115a ) or ( a2116a );
 a6873a <=( a2113a ) or ( a2114a );
 a6874a <=( a6873a ) or ( a6870a );
 a6875a <=( a6874a ) or ( a6867a );
 a6876a <=( a6875a ) or ( a6860a );
 a6877a <=( a6876a ) or ( a6847a );
 a6881a <=( a2110a ) or ( a2111a );
 a6882a <=( a2112a ) or ( a6881a );
 a6885a <=( a2108a ) or ( a2109a );
 a6888a <=( a2106a ) or ( a2107a );
 a6889a <=( a6888a ) or ( a6885a );
 a6890a <=( a6889a ) or ( a6882a );
 a6894a <=( a2103a ) or ( a2104a );
 a6895a <=( a2105a ) or ( a6894a );
 a6898a <=( a2101a ) or ( a2102a );
 a6901a <=( a2099a ) or ( a2100a );
 a6902a <=( a6901a ) or ( a6898a );
 a6903a <=( a6902a ) or ( a6895a );
 a6904a <=( a6903a ) or ( a6890a );
 a6908a <=( a2096a ) or ( a2097a );
 a6909a <=( a2098a ) or ( a6908a );
 a6912a <=( a2094a ) or ( a2095a );
 a6915a <=( a2092a ) or ( a2093a );
 a6916a <=( a6915a ) or ( a6912a );
 a6917a <=( a6916a ) or ( a6909a );
 a6920a <=( a2090a ) or ( a2091a );
 a6923a <=( a2088a ) or ( a2089a );
 a6924a <=( a6923a ) or ( a6920a );
 a6927a <=( a2086a ) or ( a2087a );
 a6930a <=( a2084a ) or ( a2085a );
 a6931a <=( a6930a ) or ( a6927a );
 a6932a <=( a6931a ) or ( a6924a );
 a6933a <=( a6932a ) or ( a6917a );
 a6934a <=( a6933a ) or ( a6904a );
 a6935a <=( a6934a ) or ( a6877a );
 a6936a <=( a6935a ) or ( a6820a );
 a6937a <=( a6936a ) or ( a6705a );
 a6941a <=( a2081a ) or ( a2082a );
 a6942a <=( a2083a ) or ( a6941a );
 a6945a <=( a2079a ) or ( a2080a );
 a6948a <=( a2077a ) or ( a2078a );
 a6949a <=( a6948a ) or ( a6945a );
 a6950a <=( a6949a ) or ( a6942a );
 a6954a <=( a2074a ) or ( a2075a );
 a6955a <=( a2076a ) or ( a6954a );
 a6958a <=( a2072a ) or ( a2073a );
 a6961a <=( a2070a ) or ( a2071a );
 a6962a <=( a6961a ) or ( a6958a );
 a6963a <=( a6962a ) or ( a6955a );
 a6964a <=( a6963a ) or ( a6950a );
 a6968a <=( a2067a ) or ( a2068a );
 a6969a <=( a2069a ) or ( a6968a );
 a6972a <=( a2065a ) or ( a2066a );
 a6975a <=( a2063a ) or ( a2064a );
 a6976a <=( a6975a ) or ( a6972a );
 a6977a <=( a6976a ) or ( a6969a );
 a6980a <=( a2061a ) or ( a2062a );
 a6983a <=( a2059a ) or ( a2060a );
 a6984a <=( a6983a ) or ( a6980a );
 a6987a <=( a2057a ) or ( a2058a );
 a6990a <=( a2055a ) or ( a2056a );
 a6991a <=( a6990a ) or ( a6987a );
 a6992a <=( a6991a ) or ( a6984a );
 a6993a <=( a6992a ) or ( a6977a );
 a6994a <=( a6993a ) or ( a6964a );
 a6998a <=( a2052a ) or ( a2053a );
 a6999a <=( a2054a ) or ( a6998a );
 a7002a <=( a2050a ) or ( a2051a );
 a7005a <=( a2048a ) or ( a2049a );
 a7006a <=( a7005a ) or ( a7002a );
 a7007a <=( a7006a ) or ( a6999a );
 a7011a <=( a2045a ) or ( a2046a );
 a7012a <=( a2047a ) or ( a7011a );
 a7015a <=( a2043a ) or ( a2044a );
 a7018a <=( a2041a ) or ( a2042a );
 a7019a <=( a7018a ) or ( a7015a );
 a7020a <=( a7019a ) or ( a7012a );
 a7021a <=( a7020a ) or ( a7007a );
 a7025a <=( a2038a ) or ( a2039a );
 a7026a <=( a2040a ) or ( a7025a );
 a7029a <=( a2036a ) or ( a2037a );
 a7032a <=( a2034a ) or ( a2035a );
 a7033a <=( a7032a ) or ( a7029a );
 a7034a <=( a7033a ) or ( a7026a );
 a7037a <=( a2032a ) or ( a2033a );
 a7040a <=( a2030a ) or ( a2031a );
 a7041a <=( a7040a ) or ( a7037a );
 a7044a <=( a2028a ) or ( a2029a );
 a7047a <=( a2026a ) or ( a2027a );
 a7048a <=( a7047a ) or ( a7044a );
 a7049a <=( a7048a ) or ( a7041a );
 a7050a <=( a7049a ) or ( a7034a );
 a7051a <=( a7050a ) or ( a7021a );
 a7052a <=( a7051a ) or ( a6994a );
 a7056a <=( a2023a ) or ( a2024a );
 a7057a <=( a2025a ) or ( a7056a );
 a7060a <=( a2021a ) or ( a2022a );
 a7063a <=( a2019a ) or ( a2020a );
 a7064a <=( a7063a ) or ( a7060a );
 a7065a <=( a7064a ) or ( a7057a );
 a7069a <=( a2016a ) or ( a2017a );
 a7070a <=( a2018a ) or ( a7069a );
 a7073a <=( a2014a ) or ( a2015a );
 a7076a <=( a2012a ) or ( a2013a );
 a7077a <=( a7076a ) or ( a7073a );
 a7078a <=( a7077a ) or ( a7070a );
 a7079a <=( a7078a ) or ( a7065a );
 a7083a <=( a2009a ) or ( a2010a );
 a7084a <=( a2011a ) or ( a7083a );
 a7087a <=( a2007a ) or ( a2008a );
 a7090a <=( a2005a ) or ( a2006a );
 a7091a <=( a7090a ) or ( a7087a );
 a7092a <=( a7091a ) or ( a7084a );
 a7095a <=( a2003a ) or ( a2004a );
 a7098a <=( a2001a ) or ( a2002a );
 a7099a <=( a7098a ) or ( a7095a );
 a7102a <=( a1999a ) or ( a2000a );
 a7105a <=( a1997a ) or ( a1998a );
 a7106a <=( a7105a ) or ( a7102a );
 a7107a <=( a7106a ) or ( a7099a );
 a7108a <=( a7107a ) or ( a7092a );
 a7109a <=( a7108a ) or ( a7079a );
 a7113a <=( a1994a ) or ( a1995a );
 a7114a <=( a1996a ) or ( a7113a );
 a7117a <=( a1992a ) or ( a1993a );
 a7120a <=( a1990a ) or ( a1991a );
 a7121a <=( a7120a ) or ( a7117a );
 a7122a <=( a7121a ) or ( a7114a );
 a7126a <=( a1987a ) or ( a1988a );
 a7127a <=( a1989a ) or ( a7126a );
 a7130a <=( a1985a ) or ( a1986a );
 a7133a <=( a1983a ) or ( a1984a );
 a7134a <=( a7133a ) or ( a7130a );
 a7135a <=( a7134a ) or ( a7127a );
 a7136a <=( a7135a ) or ( a7122a );
 a7140a <=( a1980a ) or ( a1981a );
 a7141a <=( a1982a ) or ( a7140a );
 a7144a <=( a1978a ) or ( a1979a );
 a7147a <=( a1976a ) or ( a1977a );
 a7148a <=( a7147a ) or ( a7144a );
 a7149a <=( a7148a ) or ( a7141a );
 a7152a <=( a1974a ) or ( a1975a );
 a7155a <=( a1972a ) or ( a1973a );
 a7156a <=( a7155a ) or ( a7152a );
 a7159a <=( a1970a ) or ( a1971a );
 a7162a <=( a1968a ) or ( a1969a );
 a7163a <=( a7162a ) or ( a7159a );
 a7164a <=( a7163a ) or ( a7156a );
 a7165a <=( a7164a ) or ( a7149a );
 a7166a <=( a7165a ) or ( a7136a );
 a7167a <=( a7166a ) or ( a7109a );
 a7168a <=( a7167a ) or ( a7052a );
 a7172a <=( a1965a ) or ( a1966a );
 a7173a <=( a1967a ) or ( a7172a );
 a7176a <=( a1963a ) or ( a1964a );
 a7179a <=( a1961a ) or ( a1962a );
 a7180a <=( a7179a ) or ( a7176a );
 a7181a <=( a7180a ) or ( a7173a );
 a7185a <=( a1958a ) or ( a1959a );
 a7186a <=( a1960a ) or ( a7185a );
 a7189a <=( a1956a ) or ( a1957a );
 a7192a <=( a1954a ) or ( a1955a );
 a7193a <=( a7192a ) or ( a7189a );
 a7194a <=( a7193a ) or ( a7186a );
 a7195a <=( a7194a ) or ( a7181a );
 a7199a <=( a1951a ) or ( a1952a );
 a7200a <=( a1953a ) or ( a7199a );
 a7203a <=( a1949a ) or ( a1950a );
 a7206a <=( a1947a ) or ( a1948a );
 a7207a <=( a7206a ) or ( a7203a );
 a7208a <=( a7207a ) or ( a7200a );
 a7211a <=( a1945a ) or ( a1946a );
 a7214a <=( a1943a ) or ( a1944a );
 a7215a <=( a7214a ) or ( a7211a );
 a7218a <=( a1941a ) or ( a1942a );
 a7221a <=( a1939a ) or ( a1940a );
 a7222a <=( a7221a ) or ( a7218a );
 a7223a <=( a7222a ) or ( a7215a );
 a7224a <=( a7223a ) or ( a7208a );
 a7225a <=( a7224a ) or ( a7195a );
 a7229a <=( a1936a ) or ( a1937a );
 a7230a <=( a1938a ) or ( a7229a );
 a7233a <=( a1934a ) or ( a1935a );
 a7236a <=( a1932a ) or ( a1933a );
 a7237a <=( a7236a ) or ( a7233a );
 a7238a <=( a7237a ) or ( a7230a );
 a7242a <=( a1929a ) or ( a1930a );
 a7243a <=( a1931a ) or ( a7242a );
 a7246a <=( a1927a ) or ( a1928a );
 a7249a <=( a1925a ) or ( a1926a );
 a7250a <=( a7249a ) or ( a7246a );
 a7251a <=( a7250a ) or ( a7243a );
 a7252a <=( a7251a ) or ( a7238a );
 a7256a <=( a1922a ) or ( a1923a );
 a7257a <=( a1924a ) or ( a7256a );
 a7260a <=( a1920a ) or ( a1921a );
 a7263a <=( a1918a ) or ( a1919a );
 a7264a <=( a7263a ) or ( a7260a );
 a7265a <=( a7264a ) or ( a7257a );
 a7268a <=( a1916a ) or ( a1917a );
 a7271a <=( a1914a ) or ( a1915a );
 a7272a <=( a7271a ) or ( a7268a );
 a7275a <=( a1912a ) or ( a1913a );
 a7278a <=( a1910a ) or ( a1911a );
 a7279a <=( a7278a ) or ( a7275a );
 a7280a <=( a7279a ) or ( a7272a );
 a7281a <=( a7280a ) or ( a7265a );
 a7282a <=( a7281a ) or ( a7252a );
 a7283a <=( a7282a ) or ( a7225a );
 a7287a <=( a1907a ) or ( a1908a );
 a7288a <=( a1909a ) or ( a7287a );
 a7291a <=( a1905a ) or ( a1906a );
 a7294a <=( a1903a ) or ( a1904a );
 a7295a <=( a7294a ) or ( a7291a );
 a7296a <=( a7295a ) or ( a7288a );
 a7300a <=( a1900a ) or ( a1901a );
 a7301a <=( a1902a ) or ( a7300a );
 a7304a <=( a1898a ) or ( a1899a );
 a7307a <=( a1896a ) or ( a1897a );
 a7308a <=( a7307a ) or ( a7304a );
 a7309a <=( a7308a ) or ( a7301a );
 a7310a <=( a7309a ) or ( a7296a );
 a7314a <=( a1893a ) or ( a1894a );
 a7315a <=( a1895a ) or ( a7314a );
 a7318a <=( a1891a ) or ( a1892a );
 a7321a <=( a1889a ) or ( a1890a );
 a7322a <=( a7321a ) or ( a7318a );
 a7323a <=( a7322a ) or ( a7315a );
 a7326a <=( a1887a ) or ( a1888a );
 a7329a <=( a1885a ) or ( a1886a );
 a7330a <=( a7329a ) or ( a7326a );
 a7333a <=( a1883a ) or ( a1884a );
 a7336a <=( a1881a ) or ( a1882a );
 a7337a <=( a7336a ) or ( a7333a );
 a7338a <=( a7337a ) or ( a7330a );
 a7339a <=( a7338a ) or ( a7323a );
 a7340a <=( a7339a ) or ( a7310a );
 a7344a <=( a1878a ) or ( a1879a );
 a7345a <=( a1880a ) or ( a7344a );
 a7348a <=( a1876a ) or ( a1877a );
 a7351a <=( a1874a ) or ( a1875a );
 a7352a <=( a7351a ) or ( a7348a );
 a7353a <=( a7352a ) or ( a7345a );
 a7357a <=( a1871a ) or ( a1872a );
 a7358a <=( a1873a ) or ( a7357a );
 a7361a <=( a1869a ) or ( a1870a );
 a7364a <=( a1867a ) or ( a1868a );
 a7365a <=( a7364a ) or ( a7361a );
 a7366a <=( a7365a ) or ( a7358a );
 a7367a <=( a7366a ) or ( a7353a );
 a7371a <=( a1864a ) or ( a1865a );
 a7372a <=( a1866a ) or ( a7371a );
 a7375a <=( a1862a ) or ( a1863a );
 a7378a <=( a1860a ) or ( a1861a );
 a7379a <=( a7378a ) or ( a7375a );
 a7380a <=( a7379a ) or ( a7372a );
 a7383a <=( a1858a ) or ( a1859a );
 a7386a <=( a1856a ) or ( a1857a );
 a7387a <=( a7386a ) or ( a7383a );
 a7390a <=( a1854a ) or ( a1855a );
 a7393a <=( a1852a ) or ( a1853a );
 a7394a <=( a7393a ) or ( a7390a );
 a7395a <=( a7394a ) or ( a7387a );
 a7396a <=( a7395a ) or ( a7380a );
 a7397a <=( a7396a ) or ( a7367a );
 a7398a <=( a7397a ) or ( a7340a );
 a7399a <=( a7398a ) or ( a7283a );
 a7400a <=( a7399a ) or ( a7168a );
 a7401a <=( a7400a ) or ( a6937a );
 a7402a <=( a7401a ) or ( a6476a );
 a7403a <=( a7402a ) or ( a5551a );
 a7407a <=( a1849a ) or ( a1850a );
 a7408a <=( a1851a ) or ( a7407a );
 a7411a <=( a1847a ) or ( a1848a );
 a7414a <=( a1845a ) or ( a1846a );
 a7415a <=( a7414a ) or ( a7411a );
 a7416a <=( a7415a ) or ( a7408a );
 a7420a <=( a1842a ) or ( a1843a );
 a7421a <=( a1844a ) or ( a7420a );
 a7424a <=( a1840a ) or ( a1841a );
 a7427a <=( a1838a ) or ( a1839a );
 a7428a <=( a7427a ) or ( a7424a );
 a7429a <=( a7428a ) or ( a7421a );
 a7430a <=( a7429a ) or ( a7416a );
 a7434a <=( a1835a ) or ( a1836a );
 a7435a <=( a1837a ) or ( a7434a );
 a7438a <=( a1833a ) or ( a1834a );
 a7441a <=( a1831a ) or ( a1832a );
 a7442a <=( a7441a ) or ( a7438a );
 a7443a <=( a7442a ) or ( a7435a );
 a7447a <=( a1828a ) or ( a1829a );
 a7448a <=( a1830a ) or ( a7447a );
 a7451a <=( a1826a ) or ( a1827a );
 a7454a <=( a1824a ) or ( a1825a );
 a7455a <=( a7454a ) or ( a7451a );
 a7456a <=( a7455a ) or ( a7448a );
 a7457a <=( a7456a ) or ( a7443a );
 a7458a <=( a7457a ) or ( a7430a );
 a7462a <=( a1821a ) or ( a1822a );
 a7463a <=( a1823a ) or ( a7462a );
 a7466a <=( a1819a ) or ( a1820a );
 a7469a <=( a1817a ) or ( a1818a );
 a7470a <=( a7469a ) or ( a7466a );
 a7471a <=( a7470a ) or ( a7463a );
 a7475a <=( a1814a ) or ( a1815a );
 a7476a <=( a1816a ) or ( a7475a );
 a7479a <=( a1812a ) or ( a1813a );
 a7482a <=( a1810a ) or ( a1811a );
 a7483a <=( a7482a ) or ( a7479a );
 a7484a <=( a7483a ) or ( a7476a );
 a7485a <=( a7484a ) or ( a7471a );
 a7489a <=( a1807a ) or ( a1808a );
 a7490a <=( a1809a ) or ( a7489a );
 a7493a <=( a1805a ) or ( a1806a );
 a7496a <=( a1803a ) or ( a1804a );
 a7497a <=( a7496a ) or ( a7493a );
 a7498a <=( a7497a ) or ( a7490a );
 a7501a <=( a1801a ) or ( a1802a );
 a7504a <=( a1799a ) or ( a1800a );
 a7505a <=( a7504a ) or ( a7501a );
 a7508a <=( a1797a ) or ( a1798a );
 a7511a <=( a1795a ) or ( a1796a );
 a7512a <=( a7511a ) or ( a7508a );
 a7513a <=( a7512a ) or ( a7505a );
 a7514a <=( a7513a ) or ( a7498a );
 a7515a <=( a7514a ) or ( a7485a );
 a7516a <=( a7515a ) or ( a7458a );
 a7520a <=( a1792a ) or ( a1793a );
 a7521a <=( a1794a ) or ( a7520a );
 a7524a <=( a1790a ) or ( a1791a );
 a7527a <=( a1788a ) or ( a1789a );
 a7528a <=( a7527a ) or ( a7524a );
 a7529a <=( a7528a ) or ( a7521a );
 a7533a <=( a1785a ) or ( a1786a );
 a7534a <=( a1787a ) or ( a7533a );
 a7537a <=( a1783a ) or ( a1784a );
 a7540a <=( a1781a ) or ( a1782a );
 a7541a <=( a7540a ) or ( a7537a );
 a7542a <=( a7541a ) or ( a7534a );
 a7543a <=( a7542a ) or ( a7529a );
 a7547a <=( a1778a ) or ( a1779a );
 a7548a <=( a1780a ) or ( a7547a );
 a7551a <=( a1776a ) or ( a1777a );
 a7554a <=( a1774a ) or ( a1775a );
 a7555a <=( a7554a ) or ( a7551a );
 a7556a <=( a7555a ) or ( a7548a );
 a7559a <=( a1772a ) or ( a1773a );
 a7562a <=( a1770a ) or ( a1771a );
 a7563a <=( a7562a ) or ( a7559a );
 a7566a <=( a1768a ) or ( a1769a );
 a7569a <=( a1766a ) or ( a1767a );
 a7570a <=( a7569a ) or ( a7566a );
 a7571a <=( a7570a ) or ( a7563a );
 a7572a <=( a7571a ) or ( a7556a );
 a7573a <=( a7572a ) or ( a7543a );
 a7577a <=( a1763a ) or ( a1764a );
 a7578a <=( a1765a ) or ( a7577a );
 a7581a <=( a1761a ) or ( a1762a );
 a7584a <=( a1759a ) or ( a1760a );
 a7585a <=( a7584a ) or ( a7581a );
 a7586a <=( a7585a ) or ( a7578a );
 a7590a <=( a1756a ) or ( a1757a );
 a7591a <=( a1758a ) or ( a7590a );
 a7594a <=( a1754a ) or ( a1755a );
 a7597a <=( a1752a ) or ( a1753a );
 a7598a <=( a7597a ) or ( a7594a );
 a7599a <=( a7598a ) or ( a7591a );
 a7600a <=( a7599a ) or ( a7586a );
 a7604a <=( a1749a ) or ( a1750a );
 a7605a <=( a1751a ) or ( a7604a );
 a7608a <=( a1747a ) or ( a1748a );
 a7611a <=( a1745a ) or ( a1746a );
 a7612a <=( a7611a ) or ( a7608a );
 a7613a <=( a7612a ) or ( a7605a );
 a7616a <=( a1743a ) or ( a1744a );
 a7619a <=( a1741a ) or ( a1742a );
 a7620a <=( a7619a ) or ( a7616a );
 a7623a <=( a1739a ) or ( a1740a );
 a7626a <=( a1737a ) or ( a1738a );
 a7627a <=( a7626a ) or ( a7623a );
 a7628a <=( a7627a ) or ( a7620a );
 a7629a <=( a7628a ) or ( a7613a );
 a7630a <=( a7629a ) or ( a7600a );
 a7631a <=( a7630a ) or ( a7573a );
 a7632a <=( a7631a ) or ( a7516a );
 a7636a <=( a1734a ) or ( a1735a );
 a7637a <=( a1736a ) or ( a7636a );
 a7640a <=( a1732a ) or ( a1733a );
 a7643a <=( a1730a ) or ( a1731a );
 a7644a <=( a7643a ) or ( a7640a );
 a7645a <=( a7644a ) or ( a7637a );
 a7649a <=( a1727a ) or ( a1728a );
 a7650a <=( a1729a ) or ( a7649a );
 a7653a <=( a1725a ) or ( a1726a );
 a7656a <=( a1723a ) or ( a1724a );
 a7657a <=( a7656a ) or ( a7653a );
 a7658a <=( a7657a ) or ( a7650a );
 a7659a <=( a7658a ) or ( a7645a );
 a7663a <=( a1720a ) or ( a1721a );
 a7664a <=( a1722a ) or ( a7663a );
 a7667a <=( a1718a ) or ( a1719a );
 a7670a <=( a1716a ) or ( a1717a );
 a7671a <=( a7670a ) or ( a7667a );
 a7672a <=( a7671a ) or ( a7664a );
 a7675a <=( a1714a ) or ( a1715a );
 a7678a <=( a1712a ) or ( a1713a );
 a7679a <=( a7678a ) or ( a7675a );
 a7682a <=( a1710a ) or ( a1711a );
 a7685a <=( a1708a ) or ( a1709a );
 a7686a <=( a7685a ) or ( a7682a );
 a7687a <=( a7686a ) or ( a7679a );
 a7688a <=( a7687a ) or ( a7672a );
 a7689a <=( a7688a ) or ( a7659a );
 a7693a <=( a1705a ) or ( a1706a );
 a7694a <=( a1707a ) or ( a7693a );
 a7697a <=( a1703a ) or ( a1704a );
 a7700a <=( a1701a ) or ( a1702a );
 a7701a <=( a7700a ) or ( a7697a );
 a7702a <=( a7701a ) or ( a7694a );
 a7706a <=( a1698a ) or ( a1699a );
 a7707a <=( a1700a ) or ( a7706a );
 a7710a <=( a1696a ) or ( a1697a );
 a7713a <=( a1694a ) or ( a1695a );
 a7714a <=( a7713a ) or ( a7710a );
 a7715a <=( a7714a ) or ( a7707a );
 a7716a <=( a7715a ) or ( a7702a );
 a7720a <=( a1691a ) or ( a1692a );
 a7721a <=( a1693a ) or ( a7720a );
 a7724a <=( a1689a ) or ( a1690a );
 a7727a <=( a1687a ) or ( a1688a );
 a7728a <=( a7727a ) or ( a7724a );
 a7729a <=( a7728a ) or ( a7721a );
 a7732a <=( a1685a ) or ( a1686a );
 a7735a <=( a1683a ) or ( a1684a );
 a7736a <=( a7735a ) or ( a7732a );
 a7739a <=( a1681a ) or ( a1682a );
 a7742a <=( a1679a ) or ( a1680a );
 a7743a <=( a7742a ) or ( a7739a );
 a7744a <=( a7743a ) or ( a7736a );
 a7745a <=( a7744a ) or ( a7729a );
 a7746a <=( a7745a ) or ( a7716a );
 a7747a <=( a7746a ) or ( a7689a );
 a7751a <=( a1676a ) or ( a1677a );
 a7752a <=( a1678a ) or ( a7751a );
 a7755a <=( a1674a ) or ( a1675a );
 a7758a <=( a1672a ) or ( a1673a );
 a7759a <=( a7758a ) or ( a7755a );
 a7760a <=( a7759a ) or ( a7752a );
 a7764a <=( a1669a ) or ( a1670a );
 a7765a <=( a1671a ) or ( a7764a );
 a7768a <=( a1667a ) or ( a1668a );
 a7771a <=( a1665a ) or ( a1666a );
 a7772a <=( a7771a ) or ( a7768a );
 a7773a <=( a7772a ) or ( a7765a );
 a7774a <=( a7773a ) or ( a7760a );
 a7778a <=( a1662a ) or ( a1663a );
 a7779a <=( a1664a ) or ( a7778a );
 a7782a <=( a1660a ) or ( a1661a );
 a7785a <=( a1658a ) or ( a1659a );
 a7786a <=( a7785a ) or ( a7782a );
 a7787a <=( a7786a ) or ( a7779a );
 a7790a <=( a1656a ) or ( a1657a );
 a7793a <=( a1654a ) or ( a1655a );
 a7794a <=( a7793a ) or ( a7790a );
 a7797a <=( a1652a ) or ( a1653a );
 a7800a <=( a1650a ) or ( a1651a );
 a7801a <=( a7800a ) or ( a7797a );
 a7802a <=( a7801a ) or ( a7794a );
 a7803a <=( a7802a ) or ( a7787a );
 a7804a <=( a7803a ) or ( a7774a );
 a7808a <=( a1647a ) or ( a1648a );
 a7809a <=( a1649a ) or ( a7808a );
 a7812a <=( a1645a ) or ( a1646a );
 a7815a <=( a1643a ) or ( a1644a );
 a7816a <=( a7815a ) or ( a7812a );
 a7817a <=( a7816a ) or ( a7809a );
 a7821a <=( a1640a ) or ( a1641a );
 a7822a <=( a1642a ) or ( a7821a );
 a7825a <=( a1638a ) or ( a1639a );
 a7828a <=( a1636a ) or ( a1637a );
 a7829a <=( a7828a ) or ( a7825a );
 a7830a <=( a7829a ) or ( a7822a );
 a7831a <=( a7830a ) or ( a7817a );
 a7835a <=( a1633a ) or ( a1634a );
 a7836a <=( a1635a ) or ( a7835a );
 a7839a <=( a1631a ) or ( a1632a );
 a7842a <=( a1629a ) or ( a1630a );
 a7843a <=( a7842a ) or ( a7839a );
 a7844a <=( a7843a ) or ( a7836a );
 a7847a <=( a1627a ) or ( a1628a );
 a7850a <=( a1625a ) or ( a1626a );
 a7851a <=( a7850a ) or ( a7847a );
 a7854a <=( a1623a ) or ( a1624a );
 a7857a <=( a1621a ) or ( a1622a );
 a7858a <=( a7857a ) or ( a7854a );
 a7859a <=( a7858a ) or ( a7851a );
 a7860a <=( a7859a ) or ( a7844a );
 a7861a <=( a7860a ) or ( a7831a );
 a7862a <=( a7861a ) or ( a7804a );
 a7863a <=( a7862a ) or ( a7747a );
 a7864a <=( a7863a ) or ( a7632a );
 a7868a <=( a1618a ) or ( a1619a );
 a7869a <=( a1620a ) or ( a7868a );
 a7872a <=( a1616a ) or ( a1617a );
 a7875a <=( a1614a ) or ( a1615a );
 a7876a <=( a7875a ) or ( a7872a );
 a7877a <=( a7876a ) or ( a7869a );
 a7881a <=( a1611a ) or ( a1612a );
 a7882a <=( a1613a ) or ( a7881a );
 a7885a <=( a1609a ) or ( a1610a );
 a7888a <=( a1607a ) or ( a1608a );
 a7889a <=( a7888a ) or ( a7885a );
 a7890a <=( a7889a ) or ( a7882a );
 a7891a <=( a7890a ) or ( a7877a );
 a7895a <=( a1604a ) or ( a1605a );
 a7896a <=( a1606a ) or ( a7895a );
 a7899a <=( a1602a ) or ( a1603a );
 a7902a <=( a1600a ) or ( a1601a );
 a7903a <=( a7902a ) or ( a7899a );
 a7904a <=( a7903a ) or ( a7896a );
 a7908a <=( a1597a ) or ( a1598a );
 a7909a <=( a1599a ) or ( a7908a );
 a7912a <=( a1595a ) or ( a1596a );
 a7915a <=( a1593a ) or ( a1594a );
 a7916a <=( a7915a ) or ( a7912a );
 a7917a <=( a7916a ) or ( a7909a );
 a7918a <=( a7917a ) or ( a7904a );
 a7919a <=( a7918a ) or ( a7891a );
 a7923a <=( a1590a ) or ( a1591a );
 a7924a <=( a1592a ) or ( a7923a );
 a7927a <=( a1588a ) or ( a1589a );
 a7930a <=( a1586a ) or ( a1587a );
 a7931a <=( a7930a ) or ( a7927a );
 a7932a <=( a7931a ) or ( a7924a );
 a7936a <=( a1583a ) or ( a1584a );
 a7937a <=( a1585a ) or ( a7936a );
 a7940a <=( a1581a ) or ( a1582a );
 a7943a <=( a1579a ) or ( a1580a );
 a7944a <=( a7943a ) or ( a7940a );
 a7945a <=( a7944a ) or ( a7937a );
 a7946a <=( a7945a ) or ( a7932a );
 a7950a <=( a1576a ) or ( a1577a );
 a7951a <=( a1578a ) or ( a7950a );
 a7954a <=( a1574a ) or ( a1575a );
 a7957a <=( a1572a ) or ( a1573a );
 a7958a <=( a7957a ) or ( a7954a );
 a7959a <=( a7958a ) or ( a7951a );
 a7962a <=( a1570a ) or ( a1571a );
 a7965a <=( a1568a ) or ( a1569a );
 a7966a <=( a7965a ) or ( a7962a );
 a7969a <=( a1566a ) or ( a1567a );
 a7972a <=( a1564a ) or ( a1565a );
 a7973a <=( a7972a ) or ( a7969a );
 a7974a <=( a7973a ) or ( a7966a );
 a7975a <=( a7974a ) or ( a7959a );
 a7976a <=( a7975a ) or ( a7946a );
 a7977a <=( a7976a ) or ( a7919a );
 a7981a <=( a1561a ) or ( a1562a );
 a7982a <=( a1563a ) or ( a7981a );
 a7985a <=( a1559a ) or ( a1560a );
 a7988a <=( a1557a ) or ( a1558a );
 a7989a <=( a7988a ) or ( a7985a );
 a7990a <=( a7989a ) or ( a7982a );
 a7994a <=( a1554a ) or ( a1555a );
 a7995a <=( a1556a ) or ( a7994a );
 a7998a <=( a1552a ) or ( a1553a );
 a8001a <=( a1550a ) or ( a1551a );
 a8002a <=( a8001a ) or ( a7998a );
 a8003a <=( a8002a ) or ( a7995a );
 a8004a <=( a8003a ) or ( a7990a );
 a8008a <=( a1547a ) or ( a1548a );
 a8009a <=( a1549a ) or ( a8008a );
 a8012a <=( a1545a ) or ( a1546a );
 a8015a <=( a1543a ) or ( a1544a );
 a8016a <=( a8015a ) or ( a8012a );
 a8017a <=( a8016a ) or ( a8009a );
 a8020a <=( a1541a ) or ( a1542a );
 a8023a <=( a1539a ) or ( a1540a );
 a8024a <=( a8023a ) or ( a8020a );
 a8027a <=( a1537a ) or ( a1538a );
 a8030a <=( a1535a ) or ( a1536a );
 a8031a <=( a8030a ) or ( a8027a );
 a8032a <=( a8031a ) or ( a8024a );
 a8033a <=( a8032a ) or ( a8017a );
 a8034a <=( a8033a ) or ( a8004a );
 a8038a <=( a1532a ) or ( a1533a );
 a8039a <=( a1534a ) or ( a8038a );
 a8042a <=( a1530a ) or ( a1531a );
 a8045a <=( a1528a ) or ( a1529a );
 a8046a <=( a8045a ) or ( a8042a );
 a8047a <=( a8046a ) or ( a8039a );
 a8051a <=( a1525a ) or ( a1526a );
 a8052a <=( a1527a ) or ( a8051a );
 a8055a <=( a1523a ) or ( a1524a );
 a8058a <=( a1521a ) or ( a1522a );
 a8059a <=( a8058a ) or ( a8055a );
 a8060a <=( a8059a ) or ( a8052a );
 a8061a <=( a8060a ) or ( a8047a );
 a8065a <=( a1518a ) or ( a1519a );
 a8066a <=( a1520a ) or ( a8065a );
 a8069a <=( a1516a ) or ( a1517a );
 a8072a <=( a1514a ) or ( a1515a );
 a8073a <=( a8072a ) or ( a8069a );
 a8074a <=( a8073a ) or ( a8066a );
 a8077a <=( a1512a ) or ( a1513a );
 a8080a <=( a1510a ) or ( a1511a );
 a8081a <=( a8080a ) or ( a8077a );
 a8084a <=( a1508a ) or ( a1509a );
 a8087a <=( a1506a ) or ( a1507a );
 a8088a <=( a8087a ) or ( a8084a );
 a8089a <=( a8088a ) or ( a8081a );
 a8090a <=( a8089a ) or ( a8074a );
 a8091a <=( a8090a ) or ( a8061a );
 a8092a <=( a8091a ) or ( a8034a );
 a8093a <=( a8092a ) or ( a7977a );
 a8097a <=( a1503a ) or ( a1504a );
 a8098a <=( a1505a ) or ( a8097a );
 a8101a <=( a1501a ) or ( a1502a );
 a8104a <=( a1499a ) or ( a1500a );
 a8105a <=( a8104a ) or ( a8101a );
 a8106a <=( a8105a ) or ( a8098a );
 a8110a <=( a1496a ) or ( a1497a );
 a8111a <=( a1498a ) or ( a8110a );
 a8114a <=( a1494a ) or ( a1495a );
 a8117a <=( a1492a ) or ( a1493a );
 a8118a <=( a8117a ) or ( a8114a );
 a8119a <=( a8118a ) or ( a8111a );
 a8120a <=( a8119a ) or ( a8106a );
 a8124a <=( a1489a ) or ( a1490a );
 a8125a <=( a1491a ) or ( a8124a );
 a8128a <=( a1487a ) or ( a1488a );
 a8131a <=( a1485a ) or ( a1486a );
 a8132a <=( a8131a ) or ( a8128a );
 a8133a <=( a8132a ) or ( a8125a );
 a8136a <=( a1483a ) or ( a1484a );
 a8139a <=( a1481a ) or ( a1482a );
 a8140a <=( a8139a ) or ( a8136a );
 a8143a <=( a1479a ) or ( a1480a );
 a8146a <=( a1477a ) or ( a1478a );
 a8147a <=( a8146a ) or ( a8143a );
 a8148a <=( a8147a ) or ( a8140a );
 a8149a <=( a8148a ) or ( a8133a );
 a8150a <=( a8149a ) or ( a8120a );
 a8154a <=( a1474a ) or ( a1475a );
 a8155a <=( a1476a ) or ( a8154a );
 a8158a <=( a1472a ) or ( a1473a );
 a8161a <=( a1470a ) or ( a1471a );
 a8162a <=( a8161a ) or ( a8158a );
 a8163a <=( a8162a ) or ( a8155a );
 a8167a <=( a1467a ) or ( a1468a );
 a8168a <=( a1469a ) or ( a8167a );
 a8171a <=( a1465a ) or ( a1466a );
 a8174a <=( a1463a ) or ( a1464a );
 a8175a <=( a8174a ) or ( a8171a );
 a8176a <=( a8175a ) or ( a8168a );
 a8177a <=( a8176a ) or ( a8163a );
 a8181a <=( a1460a ) or ( a1461a );
 a8182a <=( a1462a ) or ( a8181a );
 a8185a <=( a1458a ) or ( a1459a );
 a8188a <=( a1456a ) or ( a1457a );
 a8189a <=( a8188a ) or ( a8185a );
 a8190a <=( a8189a ) or ( a8182a );
 a8193a <=( a1454a ) or ( a1455a );
 a8196a <=( a1452a ) or ( a1453a );
 a8197a <=( a8196a ) or ( a8193a );
 a8200a <=( a1450a ) or ( a1451a );
 a8203a <=( a1448a ) or ( a1449a );
 a8204a <=( a8203a ) or ( a8200a );
 a8205a <=( a8204a ) or ( a8197a );
 a8206a <=( a8205a ) or ( a8190a );
 a8207a <=( a8206a ) or ( a8177a );
 a8208a <=( a8207a ) or ( a8150a );
 a8212a <=( a1445a ) or ( a1446a );
 a8213a <=( a1447a ) or ( a8212a );
 a8216a <=( a1443a ) or ( a1444a );
 a8219a <=( a1441a ) or ( a1442a );
 a8220a <=( a8219a ) or ( a8216a );
 a8221a <=( a8220a ) or ( a8213a );
 a8225a <=( a1438a ) or ( a1439a );
 a8226a <=( a1440a ) or ( a8225a );
 a8229a <=( a1436a ) or ( a1437a );
 a8232a <=( a1434a ) or ( a1435a );
 a8233a <=( a8232a ) or ( a8229a );
 a8234a <=( a8233a ) or ( a8226a );
 a8235a <=( a8234a ) or ( a8221a );
 a8239a <=( a1431a ) or ( a1432a );
 a8240a <=( a1433a ) or ( a8239a );
 a8243a <=( a1429a ) or ( a1430a );
 a8246a <=( a1427a ) or ( a1428a );
 a8247a <=( a8246a ) or ( a8243a );
 a8248a <=( a8247a ) or ( a8240a );
 a8251a <=( a1425a ) or ( a1426a );
 a8254a <=( a1423a ) or ( a1424a );
 a8255a <=( a8254a ) or ( a8251a );
 a8258a <=( a1421a ) or ( a1422a );
 a8261a <=( a1419a ) or ( a1420a );
 a8262a <=( a8261a ) or ( a8258a );
 a8263a <=( a8262a ) or ( a8255a );
 a8264a <=( a8263a ) or ( a8248a );
 a8265a <=( a8264a ) or ( a8235a );
 a8269a <=( a1416a ) or ( a1417a );
 a8270a <=( a1418a ) or ( a8269a );
 a8273a <=( a1414a ) or ( a1415a );
 a8276a <=( a1412a ) or ( a1413a );
 a8277a <=( a8276a ) or ( a8273a );
 a8278a <=( a8277a ) or ( a8270a );
 a8282a <=( a1409a ) or ( a1410a );
 a8283a <=( a1411a ) or ( a8282a );
 a8286a <=( a1407a ) or ( a1408a );
 a8289a <=( a1405a ) or ( a1406a );
 a8290a <=( a8289a ) or ( a8286a );
 a8291a <=( a8290a ) or ( a8283a );
 a8292a <=( a8291a ) or ( a8278a );
 a8296a <=( a1402a ) or ( a1403a );
 a8297a <=( a1404a ) or ( a8296a );
 a8300a <=( a1400a ) or ( a1401a );
 a8303a <=( a1398a ) or ( a1399a );
 a8304a <=( a8303a ) or ( a8300a );
 a8305a <=( a8304a ) or ( a8297a );
 a8308a <=( a1396a ) or ( a1397a );
 a8311a <=( a1394a ) or ( a1395a );
 a8312a <=( a8311a ) or ( a8308a );
 a8315a <=( a1392a ) or ( a1393a );
 a8318a <=( a1390a ) or ( a1391a );
 a8319a <=( a8318a ) or ( a8315a );
 a8320a <=( a8319a ) or ( a8312a );
 a8321a <=( a8320a ) or ( a8305a );
 a8322a <=( a8321a ) or ( a8292a );
 a8323a <=( a8322a ) or ( a8265a );
 a8324a <=( a8323a ) or ( a8208a );
 a8325a <=( a8324a ) or ( a8093a );
 a8326a <=( a8325a ) or ( a7864a );
 a8330a <=( a1387a ) or ( a1388a );
 a8331a <=( a1389a ) or ( a8330a );
 a8334a <=( a1385a ) or ( a1386a );
 a8337a <=( a1383a ) or ( a1384a );
 a8338a <=( a8337a ) or ( a8334a );
 a8339a <=( a8338a ) or ( a8331a );
 a8343a <=( a1380a ) or ( a1381a );
 a8344a <=( a1382a ) or ( a8343a );
 a8347a <=( a1378a ) or ( a1379a );
 a8350a <=( a1376a ) or ( a1377a );
 a8351a <=( a8350a ) or ( a8347a );
 a8352a <=( a8351a ) or ( a8344a );
 a8353a <=( a8352a ) or ( a8339a );
 a8357a <=( a1373a ) or ( a1374a );
 a8358a <=( a1375a ) or ( a8357a );
 a8361a <=( a1371a ) or ( a1372a );
 a8364a <=( a1369a ) or ( a1370a );
 a8365a <=( a8364a ) or ( a8361a );
 a8366a <=( a8365a ) or ( a8358a );
 a8370a <=( a1366a ) or ( a1367a );
 a8371a <=( a1368a ) or ( a8370a );
 a8374a <=( a1364a ) or ( a1365a );
 a8377a <=( a1362a ) or ( a1363a );
 a8378a <=( a8377a ) or ( a8374a );
 a8379a <=( a8378a ) or ( a8371a );
 a8380a <=( a8379a ) or ( a8366a );
 a8381a <=( a8380a ) or ( a8353a );
 a8385a <=( a1359a ) or ( a1360a );
 a8386a <=( a1361a ) or ( a8385a );
 a8389a <=( a1357a ) or ( a1358a );
 a8392a <=( a1355a ) or ( a1356a );
 a8393a <=( a8392a ) or ( a8389a );
 a8394a <=( a8393a ) or ( a8386a );
 a8398a <=( a1352a ) or ( a1353a );
 a8399a <=( a1354a ) or ( a8398a );
 a8402a <=( a1350a ) or ( a1351a );
 a8405a <=( a1348a ) or ( a1349a );
 a8406a <=( a8405a ) or ( a8402a );
 a8407a <=( a8406a ) or ( a8399a );
 a8408a <=( a8407a ) or ( a8394a );
 a8412a <=( a1345a ) or ( a1346a );
 a8413a <=( a1347a ) or ( a8412a );
 a8416a <=( a1343a ) or ( a1344a );
 a8419a <=( a1341a ) or ( a1342a );
 a8420a <=( a8419a ) or ( a8416a );
 a8421a <=( a8420a ) or ( a8413a );
 a8424a <=( a1339a ) or ( a1340a );
 a8427a <=( a1337a ) or ( a1338a );
 a8428a <=( a8427a ) or ( a8424a );
 a8431a <=( a1335a ) or ( a1336a );
 a8434a <=( a1333a ) or ( a1334a );
 a8435a <=( a8434a ) or ( a8431a );
 a8436a <=( a8435a ) or ( a8428a );
 a8437a <=( a8436a ) or ( a8421a );
 a8438a <=( a8437a ) or ( a8408a );
 a8439a <=( a8438a ) or ( a8381a );
 a8443a <=( a1330a ) or ( a1331a );
 a8444a <=( a1332a ) or ( a8443a );
 a8447a <=( a1328a ) or ( a1329a );
 a8450a <=( a1326a ) or ( a1327a );
 a8451a <=( a8450a ) or ( a8447a );
 a8452a <=( a8451a ) or ( a8444a );
 a8456a <=( a1323a ) or ( a1324a );
 a8457a <=( a1325a ) or ( a8456a );
 a8460a <=( a1321a ) or ( a1322a );
 a8463a <=( a1319a ) or ( a1320a );
 a8464a <=( a8463a ) or ( a8460a );
 a8465a <=( a8464a ) or ( a8457a );
 a8466a <=( a8465a ) or ( a8452a );
 a8470a <=( a1316a ) or ( a1317a );
 a8471a <=( a1318a ) or ( a8470a );
 a8474a <=( a1314a ) or ( a1315a );
 a8477a <=( a1312a ) or ( a1313a );
 a8478a <=( a8477a ) or ( a8474a );
 a8479a <=( a8478a ) or ( a8471a );
 a8482a <=( a1310a ) or ( a1311a );
 a8485a <=( a1308a ) or ( a1309a );
 a8486a <=( a8485a ) or ( a8482a );
 a8489a <=( a1306a ) or ( a1307a );
 a8492a <=( a1304a ) or ( a1305a );
 a8493a <=( a8492a ) or ( a8489a );
 a8494a <=( a8493a ) or ( a8486a );
 a8495a <=( a8494a ) or ( a8479a );
 a8496a <=( a8495a ) or ( a8466a );
 a8500a <=( a1301a ) or ( a1302a );
 a8501a <=( a1303a ) or ( a8500a );
 a8504a <=( a1299a ) or ( a1300a );
 a8507a <=( a1297a ) or ( a1298a );
 a8508a <=( a8507a ) or ( a8504a );
 a8509a <=( a8508a ) or ( a8501a );
 a8513a <=( a1294a ) or ( a1295a );
 a8514a <=( a1296a ) or ( a8513a );
 a8517a <=( a1292a ) or ( a1293a );
 a8520a <=( a1290a ) or ( a1291a );
 a8521a <=( a8520a ) or ( a8517a );
 a8522a <=( a8521a ) or ( a8514a );
 a8523a <=( a8522a ) or ( a8509a );
 a8527a <=( a1287a ) or ( a1288a );
 a8528a <=( a1289a ) or ( a8527a );
 a8531a <=( a1285a ) or ( a1286a );
 a8534a <=( a1283a ) or ( a1284a );
 a8535a <=( a8534a ) or ( a8531a );
 a8536a <=( a8535a ) or ( a8528a );
 a8539a <=( a1281a ) or ( a1282a );
 a8542a <=( a1279a ) or ( a1280a );
 a8543a <=( a8542a ) or ( a8539a );
 a8546a <=( a1277a ) or ( a1278a );
 a8549a <=( a1275a ) or ( a1276a );
 a8550a <=( a8549a ) or ( a8546a );
 a8551a <=( a8550a ) or ( a8543a );
 a8552a <=( a8551a ) or ( a8536a );
 a8553a <=( a8552a ) or ( a8523a );
 a8554a <=( a8553a ) or ( a8496a );
 a8555a <=( a8554a ) or ( a8439a );
 a8559a <=( a1272a ) or ( a1273a );
 a8560a <=( a1274a ) or ( a8559a );
 a8563a <=( a1270a ) or ( a1271a );
 a8566a <=( a1268a ) or ( a1269a );
 a8567a <=( a8566a ) or ( a8563a );
 a8568a <=( a8567a ) or ( a8560a );
 a8572a <=( a1265a ) or ( a1266a );
 a8573a <=( a1267a ) or ( a8572a );
 a8576a <=( a1263a ) or ( a1264a );
 a8579a <=( a1261a ) or ( a1262a );
 a8580a <=( a8579a ) or ( a8576a );
 a8581a <=( a8580a ) or ( a8573a );
 a8582a <=( a8581a ) or ( a8568a );
 a8586a <=( a1258a ) or ( a1259a );
 a8587a <=( a1260a ) or ( a8586a );
 a8590a <=( a1256a ) or ( a1257a );
 a8593a <=( a1254a ) or ( a1255a );
 a8594a <=( a8593a ) or ( a8590a );
 a8595a <=( a8594a ) or ( a8587a );
 a8598a <=( a1252a ) or ( a1253a );
 a8601a <=( a1250a ) or ( a1251a );
 a8602a <=( a8601a ) or ( a8598a );
 a8605a <=( a1248a ) or ( a1249a );
 a8608a <=( a1246a ) or ( a1247a );
 a8609a <=( a8608a ) or ( a8605a );
 a8610a <=( a8609a ) or ( a8602a );
 a8611a <=( a8610a ) or ( a8595a );
 a8612a <=( a8611a ) or ( a8582a );
 a8616a <=( a1243a ) or ( a1244a );
 a8617a <=( a1245a ) or ( a8616a );
 a8620a <=( a1241a ) or ( a1242a );
 a8623a <=( a1239a ) or ( a1240a );
 a8624a <=( a8623a ) or ( a8620a );
 a8625a <=( a8624a ) or ( a8617a );
 a8629a <=( a1236a ) or ( a1237a );
 a8630a <=( a1238a ) or ( a8629a );
 a8633a <=( a1234a ) or ( a1235a );
 a8636a <=( a1232a ) or ( a1233a );
 a8637a <=( a8636a ) or ( a8633a );
 a8638a <=( a8637a ) or ( a8630a );
 a8639a <=( a8638a ) or ( a8625a );
 a8643a <=( a1229a ) or ( a1230a );
 a8644a <=( a1231a ) or ( a8643a );
 a8647a <=( a1227a ) or ( a1228a );
 a8650a <=( a1225a ) or ( a1226a );
 a8651a <=( a8650a ) or ( a8647a );
 a8652a <=( a8651a ) or ( a8644a );
 a8655a <=( a1223a ) or ( a1224a );
 a8658a <=( a1221a ) or ( a1222a );
 a8659a <=( a8658a ) or ( a8655a );
 a8662a <=( a1219a ) or ( a1220a );
 a8665a <=( a1217a ) or ( a1218a );
 a8666a <=( a8665a ) or ( a8662a );
 a8667a <=( a8666a ) or ( a8659a );
 a8668a <=( a8667a ) or ( a8652a );
 a8669a <=( a8668a ) or ( a8639a );
 a8670a <=( a8669a ) or ( a8612a );
 a8674a <=( a1214a ) or ( a1215a );
 a8675a <=( a1216a ) or ( a8674a );
 a8678a <=( a1212a ) or ( a1213a );
 a8681a <=( a1210a ) or ( a1211a );
 a8682a <=( a8681a ) or ( a8678a );
 a8683a <=( a8682a ) or ( a8675a );
 a8687a <=( a1207a ) or ( a1208a );
 a8688a <=( a1209a ) or ( a8687a );
 a8691a <=( a1205a ) or ( a1206a );
 a8694a <=( a1203a ) or ( a1204a );
 a8695a <=( a8694a ) or ( a8691a );
 a8696a <=( a8695a ) or ( a8688a );
 a8697a <=( a8696a ) or ( a8683a );
 a8701a <=( a1200a ) or ( a1201a );
 a8702a <=( a1202a ) or ( a8701a );
 a8705a <=( a1198a ) or ( a1199a );
 a8708a <=( a1196a ) or ( a1197a );
 a8709a <=( a8708a ) or ( a8705a );
 a8710a <=( a8709a ) or ( a8702a );
 a8713a <=( a1194a ) or ( a1195a );
 a8716a <=( a1192a ) or ( a1193a );
 a8717a <=( a8716a ) or ( a8713a );
 a8720a <=( a1190a ) or ( a1191a );
 a8723a <=( a1188a ) or ( a1189a );
 a8724a <=( a8723a ) or ( a8720a );
 a8725a <=( a8724a ) or ( a8717a );
 a8726a <=( a8725a ) or ( a8710a );
 a8727a <=( a8726a ) or ( a8697a );
 a8731a <=( a1185a ) or ( a1186a );
 a8732a <=( a1187a ) or ( a8731a );
 a8735a <=( a1183a ) or ( a1184a );
 a8738a <=( a1181a ) or ( a1182a );
 a8739a <=( a8738a ) or ( a8735a );
 a8740a <=( a8739a ) or ( a8732a );
 a8744a <=( a1178a ) or ( a1179a );
 a8745a <=( a1180a ) or ( a8744a );
 a8748a <=( a1176a ) or ( a1177a );
 a8751a <=( a1174a ) or ( a1175a );
 a8752a <=( a8751a ) or ( a8748a );
 a8753a <=( a8752a ) or ( a8745a );
 a8754a <=( a8753a ) or ( a8740a );
 a8758a <=( a1171a ) or ( a1172a );
 a8759a <=( a1173a ) or ( a8758a );
 a8762a <=( a1169a ) or ( a1170a );
 a8765a <=( a1167a ) or ( a1168a );
 a8766a <=( a8765a ) or ( a8762a );
 a8767a <=( a8766a ) or ( a8759a );
 a8770a <=( a1165a ) or ( a1166a );
 a8773a <=( a1163a ) or ( a1164a );
 a8774a <=( a8773a ) or ( a8770a );
 a8777a <=( a1161a ) or ( a1162a );
 a8780a <=( a1159a ) or ( a1160a );
 a8781a <=( a8780a ) or ( a8777a );
 a8782a <=( a8781a ) or ( a8774a );
 a8783a <=( a8782a ) or ( a8767a );
 a8784a <=( a8783a ) or ( a8754a );
 a8785a <=( a8784a ) or ( a8727a );
 a8786a <=( a8785a ) or ( a8670a );
 a8787a <=( a8786a ) or ( a8555a );
 a8791a <=( a1156a ) or ( a1157a );
 a8792a <=( a1158a ) or ( a8791a );
 a8795a <=( a1154a ) or ( a1155a );
 a8798a <=( a1152a ) or ( a1153a );
 a8799a <=( a8798a ) or ( a8795a );
 a8800a <=( a8799a ) or ( a8792a );
 a8804a <=( a1149a ) or ( a1150a );
 a8805a <=( a1151a ) or ( a8804a );
 a8808a <=( a1147a ) or ( a1148a );
 a8811a <=( a1145a ) or ( a1146a );
 a8812a <=( a8811a ) or ( a8808a );
 a8813a <=( a8812a ) or ( a8805a );
 a8814a <=( a8813a ) or ( a8800a );
 a8818a <=( a1142a ) or ( a1143a );
 a8819a <=( a1144a ) or ( a8818a );
 a8822a <=( a1140a ) or ( a1141a );
 a8825a <=( a1138a ) or ( a1139a );
 a8826a <=( a8825a ) or ( a8822a );
 a8827a <=( a8826a ) or ( a8819a );
 a8830a <=( a1136a ) or ( a1137a );
 a8833a <=( a1134a ) or ( a1135a );
 a8834a <=( a8833a ) or ( a8830a );
 a8837a <=( a1132a ) or ( a1133a );
 a8840a <=( a1130a ) or ( a1131a );
 a8841a <=( a8840a ) or ( a8837a );
 a8842a <=( a8841a ) or ( a8834a );
 a8843a <=( a8842a ) or ( a8827a );
 a8844a <=( a8843a ) or ( a8814a );
 a8848a <=( a1127a ) or ( a1128a );
 a8849a <=( a1129a ) or ( a8848a );
 a8852a <=( a1125a ) or ( a1126a );
 a8855a <=( a1123a ) or ( a1124a );
 a8856a <=( a8855a ) or ( a8852a );
 a8857a <=( a8856a ) or ( a8849a );
 a8861a <=( a1120a ) or ( a1121a );
 a8862a <=( a1122a ) or ( a8861a );
 a8865a <=( a1118a ) or ( a1119a );
 a8868a <=( a1116a ) or ( a1117a );
 a8869a <=( a8868a ) or ( a8865a );
 a8870a <=( a8869a ) or ( a8862a );
 a8871a <=( a8870a ) or ( a8857a );
 a8875a <=( a1113a ) or ( a1114a );
 a8876a <=( a1115a ) or ( a8875a );
 a8879a <=( a1111a ) or ( a1112a );
 a8882a <=( a1109a ) or ( a1110a );
 a8883a <=( a8882a ) or ( a8879a );
 a8884a <=( a8883a ) or ( a8876a );
 a8887a <=( a1107a ) or ( a1108a );
 a8890a <=( a1105a ) or ( a1106a );
 a8891a <=( a8890a ) or ( a8887a );
 a8894a <=( a1103a ) or ( a1104a );
 a8897a <=( a1101a ) or ( a1102a );
 a8898a <=( a8897a ) or ( a8894a );
 a8899a <=( a8898a ) or ( a8891a );
 a8900a <=( a8899a ) or ( a8884a );
 a8901a <=( a8900a ) or ( a8871a );
 a8902a <=( a8901a ) or ( a8844a );
 a8906a <=( a1098a ) or ( a1099a );
 a8907a <=( a1100a ) or ( a8906a );
 a8910a <=( a1096a ) or ( a1097a );
 a8913a <=( a1094a ) or ( a1095a );
 a8914a <=( a8913a ) or ( a8910a );
 a8915a <=( a8914a ) or ( a8907a );
 a8919a <=( a1091a ) or ( a1092a );
 a8920a <=( a1093a ) or ( a8919a );
 a8923a <=( a1089a ) or ( a1090a );
 a8926a <=( a1087a ) or ( a1088a );
 a8927a <=( a8926a ) or ( a8923a );
 a8928a <=( a8927a ) or ( a8920a );
 a8929a <=( a8928a ) or ( a8915a );
 a8933a <=( a1084a ) or ( a1085a );
 a8934a <=( a1086a ) or ( a8933a );
 a8937a <=( a1082a ) or ( a1083a );
 a8940a <=( a1080a ) or ( a1081a );
 a8941a <=( a8940a ) or ( a8937a );
 a8942a <=( a8941a ) or ( a8934a );
 a8945a <=( a1078a ) or ( a1079a );
 a8948a <=( a1076a ) or ( a1077a );
 a8949a <=( a8948a ) or ( a8945a );
 a8952a <=( a1074a ) or ( a1075a );
 a8955a <=( a1072a ) or ( a1073a );
 a8956a <=( a8955a ) or ( a8952a );
 a8957a <=( a8956a ) or ( a8949a );
 a8958a <=( a8957a ) or ( a8942a );
 a8959a <=( a8958a ) or ( a8929a );
 a8963a <=( a1069a ) or ( a1070a );
 a8964a <=( a1071a ) or ( a8963a );
 a8967a <=( a1067a ) or ( a1068a );
 a8970a <=( a1065a ) or ( a1066a );
 a8971a <=( a8970a ) or ( a8967a );
 a8972a <=( a8971a ) or ( a8964a );
 a8976a <=( a1062a ) or ( a1063a );
 a8977a <=( a1064a ) or ( a8976a );
 a8980a <=( a1060a ) or ( a1061a );
 a8983a <=( a1058a ) or ( a1059a );
 a8984a <=( a8983a ) or ( a8980a );
 a8985a <=( a8984a ) or ( a8977a );
 a8986a <=( a8985a ) or ( a8972a );
 a8990a <=( a1055a ) or ( a1056a );
 a8991a <=( a1057a ) or ( a8990a );
 a8994a <=( a1053a ) or ( a1054a );
 a8997a <=( a1051a ) or ( a1052a );
 a8998a <=( a8997a ) or ( a8994a );
 a8999a <=( a8998a ) or ( a8991a );
 a9002a <=( a1049a ) or ( a1050a );
 a9005a <=( a1047a ) or ( a1048a );
 a9006a <=( a9005a ) or ( a9002a );
 a9009a <=( a1045a ) or ( a1046a );
 a9012a <=( a1043a ) or ( a1044a );
 a9013a <=( a9012a ) or ( a9009a );
 a9014a <=( a9013a ) or ( a9006a );
 a9015a <=( a9014a ) or ( a8999a );
 a9016a <=( a9015a ) or ( a8986a );
 a9017a <=( a9016a ) or ( a8959a );
 a9018a <=( a9017a ) or ( a8902a );
 a9022a <=( a1040a ) or ( a1041a );
 a9023a <=( a1042a ) or ( a9022a );
 a9026a <=( a1038a ) or ( a1039a );
 a9029a <=( a1036a ) or ( a1037a );
 a9030a <=( a9029a ) or ( a9026a );
 a9031a <=( a9030a ) or ( a9023a );
 a9035a <=( a1033a ) or ( a1034a );
 a9036a <=( a1035a ) or ( a9035a );
 a9039a <=( a1031a ) or ( a1032a );
 a9042a <=( a1029a ) or ( a1030a );
 a9043a <=( a9042a ) or ( a9039a );
 a9044a <=( a9043a ) or ( a9036a );
 a9045a <=( a9044a ) or ( a9031a );
 a9049a <=( a1026a ) or ( a1027a );
 a9050a <=( a1028a ) or ( a9049a );
 a9053a <=( a1024a ) or ( a1025a );
 a9056a <=( a1022a ) or ( a1023a );
 a9057a <=( a9056a ) or ( a9053a );
 a9058a <=( a9057a ) or ( a9050a );
 a9061a <=( a1020a ) or ( a1021a );
 a9064a <=( a1018a ) or ( a1019a );
 a9065a <=( a9064a ) or ( a9061a );
 a9068a <=( a1016a ) or ( a1017a );
 a9071a <=( a1014a ) or ( a1015a );
 a9072a <=( a9071a ) or ( a9068a );
 a9073a <=( a9072a ) or ( a9065a );
 a9074a <=( a9073a ) or ( a9058a );
 a9075a <=( a9074a ) or ( a9045a );
 a9079a <=( a1011a ) or ( a1012a );
 a9080a <=( a1013a ) or ( a9079a );
 a9083a <=( a1009a ) or ( a1010a );
 a9086a <=( a1007a ) or ( a1008a );
 a9087a <=( a9086a ) or ( a9083a );
 a9088a <=( a9087a ) or ( a9080a );
 a9092a <=( a1004a ) or ( a1005a );
 a9093a <=( a1006a ) or ( a9092a );
 a9096a <=( a1002a ) or ( a1003a );
 a9099a <=( a1000a ) or ( a1001a );
 a9100a <=( a9099a ) or ( a9096a );
 a9101a <=( a9100a ) or ( a9093a );
 a9102a <=( a9101a ) or ( a9088a );
 a9106a <=( a997a ) or ( a998a );
 a9107a <=( a999a ) or ( a9106a );
 a9110a <=( a995a ) or ( a996a );
 a9113a <=( a993a ) or ( a994a );
 a9114a <=( a9113a ) or ( a9110a );
 a9115a <=( a9114a ) or ( a9107a );
 a9118a <=( a991a ) or ( a992a );
 a9121a <=( a989a ) or ( a990a );
 a9122a <=( a9121a ) or ( a9118a );
 a9125a <=( a987a ) or ( a988a );
 a9128a <=( a985a ) or ( a986a );
 a9129a <=( a9128a ) or ( a9125a );
 a9130a <=( a9129a ) or ( a9122a );
 a9131a <=( a9130a ) or ( a9115a );
 a9132a <=( a9131a ) or ( a9102a );
 a9133a <=( a9132a ) or ( a9075a );
 a9137a <=( a982a ) or ( a983a );
 a9138a <=( a984a ) or ( a9137a );
 a9141a <=( a980a ) or ( a981a );
 a9144a <=( a978a ) or ( a979a );
 a9145a <=( a9144a ) or ( a9141a );
 a9146a <=( a9145a ) or ( a9138a );
 a9150a <=( a975a ) or ( a976a );
 a9151a <=( a977a ) or ( a9150a );
 a9154a <=( a973a ) or ( a974a );
 a9157a <=( a971a ) or ( a972a );
 a9158a <=( a9157a ) or ( a9154a );
 a9159a <=( a9158a ) or ( a9151a );
 a9160a <=( a9159a ) or ( a9146a );
 a9164a <=( a968a ) or ( a969a );
 a9165a <=( a970a ) or ( a9164a );
 a9168a <=( a966a ) or ( a967a );
 a9171a <=( a964a ) or ( a965a );
 a9172a <=( a9171a ) or ( a9168a );
 a9173a <=( a9172a ) or ( a9165a );
 a9176a <=( a962a ) or ( a963a );
 a9179a <=( a960a ) or ( a961a );
 a9180a <=( a9179a ) or ( a9176a );
 a9183a <=( a958a ) or ( a959a );
 a9186a <=( a956a ) or ( a957a );
 a9187a <=( a9186a ) or ( a9183a );
 a9188a <=( a9187a ) or ( a9180a );
 a9189a <=( a9188a ) or ( a9173a );
 a9190a <=( a9189a ) or ( a9160a );
 a9194a <=( a953a ) or ( a954a );
 a9195a <=( a955a ) or ( a9194a );
 a9198a <=( a951a ) or ( a952a );
 a9201a <=( a949a ) or ( a950a );
 a9202a <=( a9201a ) or ( a9198a );
 a9203a <=( a9202a ) or ( a9195a );
 a9207a <=( a946a ) or ( a947a );
 a9208a <=( a948a ) or ( a9207a );
 a9211a <=( a944a ) or ( a945a );
 a9214a <=( a942a ) or ( a943a );
 a9215a <=( a9214a ) or ( a9211a );
 a9216a <=( a9215a ) or ( a9208a );
 a9217a <=( a9216a ) or ( a9203a );
 a9221a <=( a939a ) or ( a940a );
 a9222a <=( a941a ) or ( a9221a );
 a9225a <=( a937a ) or ( a938a );
 a9228a <=( a935a ) or ( a936a );
 a9229a <=( a9228a ) or ( a9225a );
 a9230a <=( a9229a ) or ( a9222a );
 a9233a <=( a933a ) or ( a934a );
 a9236a <=( a931a ) or ( a932a );
 a9237a <=( a9236a ) or ( a9233a );
 a9240a <=( a929a ) or ( a930a );
 a9243a <=( a927a ) or ( a928a );
 a9244a <=( a9243a ) or ( a9240a );
 a9245a <=( a9244a ) or ( a9237a );
 a9246a <=( a9245a ) or ( a9230a );
 a9247a <=( a9246a ) or ( a9217a );
 a9248a <=( a9247a ) or ( a9190a );
 a9249a <=( a9248a ) or ( a9133a );
 a9250a <=( a9249a ) or ( a9018a );
 a9251a <=( a9250a ) or ( a8787a );
 a9252a <=( a9251a ) or ( a8326a );
 a9256a <=( a924a ) or ( a925a );
 a9257a <=( a926a ) or ( a9256a );
 a9260a <=( a922a ) or ( a923a );
 a9263a <=( a920a ) or ( a921a );
 a9264a <=( a9263a ) or ( a9260a );
 a9265a <=( a9264a ) or ( a9257a );
 a9269a <=( a917a ) or ( a918a );
 a9270a <=( a919a ) or ( a9269a );
 a9273a <=( a915a ) or ( a916a );
 a9276a <=( a913a ) or ( a914a );
 a9277a <=( a9276a ) or ( a9273a );
 a9278a <=( a9277a ) or ( a9270a );
 a9279a <=( a9278a ) or ( a9265a );
 a9283a <=( a910a ) or ( a911a );
 a9284a <=( a912a ) or ( a9283a );
 a9287a <=( a908a ) or ( a909a );
 a9290a <=( a906a ) or ( a907a );
 a9291a <=( a9290a ) or ( a9287a );
 a9292a <=( a9291a ) or ( a9284a );
 a9296a <=( a903a ) or ( a904a );
 a9297a <=( a905a ) or ( a9296a );
 a9300a <=( a901a ) or ( a902a );
 a9303a <=( a899a ) or ( a900a );
 a9304a <=( a9303a ) or ( a9300a );
 a9305a <=( a9304a ) or ( a9297a );
 a9306a <=( a9305a ) or ( a9292a );
 a9307a <=( a9306a ) or ( a9279a );
 a9311a <=( a896a ) or ( a897a );
 a9312a <=( a898a ) or ( a9311a );
 a9315a <=( a894a ) or ( a895a );
 a9318a <=( a892a ) or ( a893a );
 a9319a <=( a9318a ) or ( a9315a );
 a9320a <=( a9319a ) or ( a9312a );
 a9324a <=( a889a ) or ( a890a );
 a9325a <=( a891a ) or ( a9324a );
 a9328a <=( a887a ) or ( a888a );
 a9331a <=( a885a ) or ( a886a );
 a9332a <=( a9331a ) or ( a9328a );
 a9333a <=( a9332a ) or ( a9325a );
 a9334a <=( a9333a ) or ( a9320a );
 a9338a <=( a882a ) or ( a883a );
 a9339a <=( a884a ) or ( a9338a );
 a9342a <=( a880a ) or ( a881a );
 a9345a <=( a878a ) or ( a879a );
 a9346a <=( a9345a ) or ( a9342a );
 a9347a <=( a9346a ) or ( a9339a );
 a9350a <=( a876a ) or ( a877a );
 a9353a <=( a874a ) or ( a875a );
 a9354a <=( a9353a ) or ( a9350a );
 a9357a <=( a872a ) or ( a873a );
 a9360a <=( a870a ) or ( a871a );
 a9361a <=( a9360a ) or ( a9357a );
 a9362a <=( a9361a ) or ( a9354a );
 a9363a <=( a9362a ) or ( a9347a );
 a9364a <=( a9363a ) or ( a9334a );
 a9365a <=( a9364a ) or ( a9307a );
 a9369a <=( a867a ) or ( a868a );
 a9370a <=( a869a ) or ( a9369a );
 a9373a <=( a865a ) or ( a866a );
 a9376a <=( a863a ) or ( a864a );
 a9377a <=( a9376a ) or ( a9373a );
 a9378a <=( a9377a ) or ( a9370a );
 a9382a <=( a860a ) or ( a861a );
 a9383a <=( a862a ) or ( a9382a );
 a9386a <=( a858a ) or ( a859a );
 a9389a <=( a856a ) or ( a857a );
 a9390a <=( a9389a ) or ( a9386a );
 a9391a <=( a9390a ) or ( a9383a );
 a9392a <=( a9391a ) or ( a9378a );
 a9396a <=( a853a ) or ( a854a );
 a9397a <=( a855a ) or ( a9396a );
 a9400a <=( a851a ) or ( a852a );
 a9403a <=( a849a ) or ( a850a );
 a9404a <=( a9403a ) or ( a9400a );
 a9405a <=( a9404a ) or ( a9397a );
 a9408a <=( a847a ) or ( a848a );
 a9411a <=( a845a ) or ( a846a );
 a9412a <=( a9411a ) or ( a9408a );
 a9415a <=( a843a ) or ( a844a );
 a9418a <=( a841a ) or ( a842a );
 a9419a <=( a9418a ) or ( a9415a );
 a9420a <=( a9419a ) or ( a9412a );
 a9421a <=( a9420a ) or ( a9405a );
 a9422a <=( a9421a ) or ( a9392a );
 a9426a <=( a838a ) or ( a839a );
 a9427a <=( a840a ) or ( a9426a );
 a9430a <=( a836a ) or ( a837a );
 a9433a <=( a834a ) or ( a835a );
 a9434a <=( a9433a ) or ( a9430a );
 a9435a <=( a9434a ) or ( a9427a );
 a9439a <=( a831a ) or ( a832a );
 a9440a <=( a833a ) or ( a9439a );
 a9443a <=( a829a ) or ( a830a );
 a9446a <=( a827a ) or ( a828a );
 a9447a <=( a9446a ) or ( a9443a );
 a9448a <=( a9447a ) or ( a9440a );
 a9449a <=( a9448a ) or ( a9435a );
 a9453a <=( a824a ) or ( a825a );
 a9454a <=( a826a ) or ( a9453a );
 a9457a <=( a822a ) or ( a823a );
 a9460a <=( a820a ) or ( a821a );
 a9461a <=( a9460a ) or ( a9457a );
 a9462a <=( a9461a ) or ( a9454a );
 a9465a <=( a818a ) or ( a819a );
 a9468a <=( a816a ) or ( a817a );
 a9469a <=( a9468a ) or ( a9465a );
 a9472a <=( a814a ) or ( a815a );
 a9475a <=( a812a ) or ( a813a );
 a9476a <=( a9475a ) or ( a9472a );
 a9477a <=( a9476a ) or ( a9469a );
 a9478a <=( a9477a ) or ( a9462a );
 a9479a <=( a9478a ) or ( a9449a );
 a9480a <=( a9479a ) or ( a9422a );
 a9481a <=( a9480a ) or ( a9365a );
 a9485a <=( a809a ) or ( a810a );
 a9486a <=( a811a ) or ( a9485a );
 a9489a <=( a807a ) or ( a808a );
 a9492a <=( a805a ) or ( a806a );
 a9493a <=( a9492a ) or ( a9489a );
 a9494a <=( a9493a ) or ( a9486a );
 a9498a <=( a802a ) or ( a803a );
 a9499a <=( a804a ) or ( a9498a );
 a9502a <=( a800a ) or ( a801a );
 a9505a <=( a798a ) or ( a799a );
 a9506a <=( a9505a ) or ( a9502a );
 a9507a <=( a9506a ) or ( a9499a );
 a9508a <=( a9507a ) or ( a9494a );
 a9512a <=( a795a ) or ( a796a );
 a9513a <=( a797a ) or ( a9512a );
 a9516a <=( a793a ) or ( a794a );
 a9519a <=( a791a ) or ( a792a );
 a9520a <=( a9519a ) or ( a9516a );
 a9521a <=( a9520a ) or ( a9513a );
 a9524a <=( a789a ) or ( a790a );
 a9527a <=( a787a ) or ( a788a );
 a9528a <=( a9527a ) or ( a9524a );
 a9531a <=( a785a ) or ( a786a );
 a9534a <=( a783a ) or ( a784a );
 a9535a <=( a9534a ) or ( a9531a );
 a9536a <=( a9535a ) or ( a9528a );
 a9537a <=( a9536a ) or ( a9521a );
 a9538a <=( a9537a ) or ( a9508a );
 a9542a <=( a780a ) or ( a781a );
 a9543a <=( a782a ) or ( a9542a );
 a9546a <=( a778a ) or ( a779a );
 a9549a <=( a776a ) or ( a777a );
 a9550a <=( a9549a ) or ( a9546a );
 a9551a <=( a9550a ) or ( a9543a );
 a9555a <=( a773a ) or ( a774a );
 a9556a <=( a775a ) or ( a9555a );
 a9559a <=( a771a ) or ( a772a );
 a9562a <=( a769a ) or ( a770a );
 a9563a <=( a9562a ) or ( a9559a );
 a9564a <=( a9563a ) or ( a9556a );
 a9565a <=( a9564a ) or ( a9551a );
 a9569a <=( a766a ) or ( a767a );
 a9570a <=( a768a ) or ( a9569a );
 a9573a <=( a764a ) or ( a765a );
 a9576a <=( a762a ) or ( a763a );
 a9577a <=( a9576a ) or ( a9573a );
 a9578a <=( a9577a ) or ( a9570a );
 a9581a <=( a760a ) or ( a761a );
 a9584a <=( a758a ) or ( a759a );
 a9585a <=( a9584a ) or ( a9581a );
 a9588a <=( a756a ) or ( a757a );
 a9591a <=( a754a ) or ( a755a );
 a9592a <=( a9591a ) or ( a9588a );
 a9593a <=( a9592a ) or ( a9585a );
 a9594a <=( a9593a ) or ( a9578a );
 a9595a <=( a9594a ) or ( a9565a );
 a9596a <=( a9595a ) or ( a9538a );
 a9600a <=( a751a ) or ( a752a );
 a9601a <=( a753a ) or ( a9600a );
 a9604a <=( a749a ) or ( a750a );
 a9607a <=( a747a ) or ( a748a );
 a9608a <=( a9607a ) or ( a9604a );
 a9609a <=( a9608a ) or ( a9601a );
 a9613a <=( a744a ) or ( a745a );
 a9614a <=( a746a ) or ( a9613a );
 a9617a <=( a742a ) or ( a743a );
 a9620a <=( a740a ) or ( a741a );
 a9621a <=( a9620a ) or ( a9617a );
 a9622a <=( a9621a ) or ( a9614a );
 a9623a <=( a9622a ) or ( a9609a );
 a9627a <=( a737a ) or ( a738a );
 a9628a <=( a739a ) or ( a9627a );
 a9631a <=( a735a ) or ( a736a );
 a9634a <=( a733a ) or ( a734a );
 a9635a <=( a9634a ) or ( a9631a );
 a9636a <=( a9635a ) or ( a9628a );
 a9639a <=( a731a ) or ( a732a );
 a9642a <=( a729a ) or ( a730a );
 a9643a <=( a9642a ) or ( a9639a );
 a9646a <=( a727a ) or ( a728a );
 a9649a <=( a725a ) or ( a726a );
 a9650a <=( a9649a ) or ( a9646a );
 a9651a <=( a9650a ) or ( a9643a );
 a9652a <=( a9651a ) or ( a9636a );
 a9653a <=( a9652a ) or ( a9623a );
 a9657a <=( a722a ) or ( a723a );
 a9658a <=( a724a ) or ( a9657a );
 a9661a <=( a720a ) or ( a721a );
 a9664a <=( a718a ) or ( a719a );
 a9665a <=( a9664a ) or ( a9661a );
 a9666a <=( a9665a ) or ( a9658a );
 a9670a <=( a715a ) or ( a716a );
 a9671a <=( a717a ) or ( a9670a );
 a9674a <=( a713a ) or ( a714a );
 a9677a <=( a711a ) or ( a712a );
 a9678a <=( a9677a ) or ( a9674a );
 a9679a <=( a9678a ) or ( a9671a );
 a9680a <=( a9679a ) or ( a9666a );
 a9684a <=( a708a ) or ( a709a );
 a9685a <=( a710a ) or ( a9684a );
 a9688a <=( a706a ) or ( a707a );
 a9691a <=( a704a ) or ( a705a );
 a9692a <=( a9691a ) or ( a9688a );
 a9693a <=( a9692a ) or ( a9685a );
 a9696a <=( a702a ) or ( a703a );
 a9699a <=( a700a ) or ( a701a );
 a9700a <=( a9699a ) or ( a9696a );
 a9703a <=( a698a ) or ( a699a );
 a9706a <=( a696a ) or ( a697a );
 a9707a <=( a9706a ) or ( a9703a );
 a9708a <=( a9707a ) or ( a9700a );
 a9709a <=( a9708a ) or ( a9693a );
 a9710a <=( a9709a ) or ( a9680a );
 a9711a <=( a9710a ) or ( a9653a );
 a9712a <=( a9711a ) or ( a9596a );
 a9713a <=( a9712a ) or ( a9481a );
 a9717a <=( a693a ) or ( a694a );
 a9718a <=( a695a ) or ( a9717a );
 a9721a <=( a691a ) or ( a692a );
 a9724a <=( a689a ) or ( a690a );
 a9725a <=( a9724a ) or ( a9721a );
 a9726a <=( a9725a ) or ( a9718a );
 a9730a <=( a686a ) or ( a687a );
 a9731a <=( a688a ) or ( a9730a );
 a9734a <=( a684a ) or ( a685a );
 a9737a <=( a682a ) or ( a683a );
 a9738a <=( a9737a ) or ( a9734a );
 a9739a <=( a9738a ) or ( a9731a );
 a9740a <=( a9739a ) or ( a9726a );
 a9744a <=( a679a ) or ( a680a );
 a9745a <=( a681a ) or ( a9744a );
 a9748a <=( a677a ) or ( a678a );
 a9751a <=( a675a ) or ( a676a );
 a9752a <=( a9751a ) or ( a9748a );
 a9753a <=( a9752a ) or ( a9745a );
 a9756a <=( a673a ) or ( a674a );
 a9759a <=( a671a ) or ( a672a );
 a9760a <=( a9759a ) or ( a9756a );
 a9763a <=( a669a ) or ( a670a );
 a9766a <=( a667a ) or ( a668a );
 a9767a <=( a9766a ) or ( a9763a );
 a9768a <=( a9767a ) or ( a9760a );
 a9769a <=( a9768a ) or ( a9753a );
 a9770a <=( a9769a ) or ( a9740a );
 a9774a <=( a664a ) or ( a665a );
 a9775a <=( a666a ) or ( a9774a );
 a9778a <=( a662a ) or ( a663a );
 a9781a <=( a660a ) or ( a661a );
 a9782a <=( a9781a ) or ( a9778a );
 a9783a <=( a9782a ) or ( a9775a );
 a9787a <=( a657a ) or ( a658a );
 a9788a <=( a659a ) or ( a9787a );
 a9791a <=( a655a ) or ( a656a );
 a9794a <=( a653a ) or ( a654a );
 a9795a <=( a9794a ) or ( a9791a );
 a9796a <=( a9795a ) or ( a9788a );
 a9797a <=( a9796a ) or ( a9783a );
 a9801a <=( a650a ) or ( a651a );
 a9802a <=( a652a ) or ( a9801a );
 a9805a <=( a648a ) or ( a649a );
 a9808a <=( a646a ) or ( a647a );
 a9809a <=( a9808a ) or ( a9805a );
 a9810a <=( a9809a ) or ( a9802a );
 a9813a <=( a644a ) or ( a645a );
 a9816a <=( a642a ) or ( a643a );
 a9817a <=( a9816a ) or ( a9813a );
 a9820a <=( a640a ) or ( a641a );
 a9823a <=( a638a ) or ( a639a );
 a9824a <=( a9823a ) or ( a9820a );
 a9825a <=( a9824a ) or ( a9817a );
 a9826a <=( a9825a ) or ( a9810a );
 a9827a <=( a9826a ) or ( a9797a );
 a9828a <=( a9827a ) or ( a9770a );
 a9832a <=( a635a ) or ( a636a );
 a9833a <=( a637a ) or ( a9832a );
 a9836a <=( a633a ) or ( a634a );
 a9839a <=( a631a ) or ( a632a );
 a9840a <=( a9839a ) or ( a9836a );
 a9841a <=( a9840a ) or ( a9833a );
 a9845a <=( a628a ) or ( a629a );
 a9846a <=( a630a ) or ( a9845a );
 a9849a <=( a626a ) or ( a627a );
 a9852a <=( a624a ) or ( a625a );
 a9853a <=( a9852a ) or ( a9849a );
 a9854a <=( a9853a ) or ( a9846a );
 a9855a <=( a9854a ) or ( a9841a );
 a9859a <=( a621a ) or ( a622a );
 a9860a <=( a623a ) or ( a9859a );
 a9863a <=( a619a ) or ( a620a );
 a9866a <=( a617a ) or ( a618a );
 a9867a <=( a9866a ) or ( a9863a );
 a9868a <=( a9867a ) or ( a9860a );
 a9871a <=( a615a ) or ( a616a );
 a9874a <=( a613a ) or ( a614a );
 a9875a <=( a9874a ) or ( a9871a );
 a9878a <=( a611a ) or ( a612a );
 a9881a <=( a609a ) or ( a610a );
 a9882a <=( a9881a ) or ( a9878a );
 a9883a <=( a9882a ) or ( a9875a );
 a9884a <=( a9883a ) or ( a9868a );
 a9885a <=( a9884a ) or ( a9855a );
 a9889a <=( a606a ) or ( a607a );
 a9890a <=( a608a ) or ( a9889a );
 a9893a <=( a604a ) or ( a605a );
 a9896a <=( a602a ) or ( a603a );
 a9897a <=( a9896a ) or ( a9893a );
 a9898a <=( a9897a ) or ( a9890a );
 a9902a <=( a599a ) or ( a600a );
 a9903a <=( a601a ) or ( a9902a );
 a9906a <=( a597a ) or ( a598a );
 a9909a <=( a595a ) or ( a596a );
 a9910a <=( a9909a ) or ( a9906a );
 a9911a <=( a9910a ) or ( a9903a );
 a9912a <=( a9911a ) or ( a9898a );
 a9916a <=( a592a ) or ( a593a );
 a9917a <=( a594a ) or ( a9916a );
 a9920a <=( a590a ) or ( a591a );
 a9923a <=( a588a ) or ( a589a );
 a9924a <=( a9923a ) or ( a9920a );
 a9925a <=( a9924a ) or ( a9917a );
 a9928a <=( a586a ) or ( a587a );
 a9931a <=( a584a ) or ( a585a );
 a9932a <=( a9931a ) or ( a9928a );
 a9935a <=( a582a ) or ( a583a );
 a9938a <=( a580a ) or ( a581a );
 a9939a <=( a9938a ) or ( a9935a );
 a9940a <=( a9939a ) or ( a9932a );
 a9941a <=( a9940a ) or ( a9925a );
 a9942a <=( a9941a ) or ( a9912a );
 a9943a <=( a9942a ) or ( a9885a );
 a9944a <=( a9943a ) or ( a9828a );
 a9948a <=( a577a ) or ( a578a );
 a9949a <=( a579a ) or ( a9948a );
 a9952a <=( a575a ) or ( a576a );
 a9955a <=( a573a ) or ( a574a );
 a9956a <=( a9955a ) or ( a9952a );
 a9957a <=( a9956a ) or ( a9949a );
 a9961a <=( a570a ) or ( a571a );
 a9962a <=( a572a ) or ( a9961a );
 a9965a <=( a568a ) or ( a569a );
 a9968a <=( a566a ) or ( a567a );
 a9969a <=( a9968a ) or ( a9965a );
 a9970a <=( a9969a ) or ( a9962a );
 a9971a <=( a9970a ) or ( a9957a );
 a9975a <=( a563a ) or ( a564a );
 a9976a <=( a565a ) or ( a9975a );
 a9979a <=( a561a ) or ( a562a );
 a9982a <=( a559a ) or ( a560a );
 a9983a <=( a9982a ) or ( a9979a );
 a9984a <=( a9983a ) or ( a9976a );
 a9987a <=( a557a ) or ( a558a );
 a9990a <=( a555a ) or ( a556a );
 a9991a <=( a9990a ) or ( a9987a );
 a9994a <=( a553a ) or ( a554a );
 a9997a <=( a551a ) or ( a552a );
 a9998a <=( a9997a ) or ( a9994a );
 a9999a <=( a9998a ) or ( a9991a );
 a10000a <=( a9999a ) or ( a9984a );
 a10001a <=( a10000a ) or ( a9971a );
 a10005a <=( a548a ) or ( a549a );
 a10006a <=( a550a ) or ( a10005a );
 a10009a <=( a546a ) or ( a547a );
 a10012a <=( a544a ) or ( a545a );
 a10013a <=( a10012a ) or ( a10009a );
 a10014a <=( a10013a ) or ( a10006a );
 a10018a <=( a541a ) or ( a542a );
 a10019a <=( a543a ) or ( a10018a );
 a10022a <=( a539a ) or ( a540a );
 a10025a <=( a537a ) or ( a538a );
 a10026a <=( a10025a ) or ( a10022a );
 a10027a <=( a10026a ) or ( a10019a );
 a10028a <=( a10027a ) or ( a10014a );
 a10032a <=( a534a ) or ( a535a );
 a10033a <=( a536a ) or ( a10032a );
 a10036a <=( a532a ) or ( a533a );
 a10039a <=( a530a ) or ( a531a );
 a10040a <=( a10039a ) or ( a10036a );
 a10041a <=( a10040a ) or ( a10033a );
 a10044a <=( a528a ) or ( a529a );
 a10047a <=( a526a ) or ( a527a );
 a10048a <=( a10047a ) or ( a10044a );
 a10051a <=( a524a ) or ( a525a );
 a10054a <=( a522a ) or ( a523a );
 a10055a <=( a10054a ) or ( a10051a );
 a10056a <=( a10055a ) or ( a10048a );
 a10057a <=( a10056a ) or ( a10041a );
 a10058a <=( a10057a ) or ( a10028a );
 a10059a <=( a10058a ) or ( a10001a );
 a10063a <=( a519a ) or ( a520a );
 a10064a <=( a521a ) or ( a10063a );
 a10067a <=( a517a ) or ( a518a );
 a10070a <=( a515a ) or ( a516a );
 a10071a <=( a10070a ) or ( a10067a );
 a10072a <=( a10071a ) or ( a10064a );
 a10076a <=( a512a ) or ( a513a );
 a10077a <=( a514a ) or ( a10076a );
 a10080a <=( a510a ) or ( a511a );
 a10083a <=( a508a ) or ( a509a );
 a10084a <=( a10083a ) or ( a10080a );
 a10085a <=( a10084a ) or ( a10077a );
 a10086a <=( a10085a ) or ( a10072a );
 a10090a <=( a505a ) or ( a506a );
 a10091a <=( a507a ) or ( a10090a );
 a10094a <=( a503a ) or ( a504a );
 a10097a <=( a501a ) or ( a502a );
 a10098a <=( a10097a ) or ( a10094a );
 a10099a <=( a10098a ) or ( a10091a );
 a10102a <=( a499a ) or ( a500a );
 a10105a <=( a497a ) or ( a498a );
 a10106a <=( a10105a ) or ( a10102a );
 a10109a <=( a495a ) or ( a496a );
 a10112a <=( a493a ) or ( a494a );
 a10113a <=( a10112a ) or ( a10109a );
 a10114a <=( a10113a ) or ( a10106a );
 a10115a <=( a10114a ) or ( a10099a );
 a10116a <=( a10115a ) or ( a10086a );
 a10120a <=( a490a ) or ( a491a );
 a10121a <=( a492a ) or ( a10120a );
 a10124a <=( a488a ) or ( a489a );
 a10127a <=( a486a ) or ( a487a );
 a10128a <=( a10127a ) or ( a10124a );
 a10129a <=( a10128a ) or ( a10121a );
 a10133a <=( a483a ) or ( a484a );
 a10134a <=( a485a ) or ( a10133a );
 a10137a <=( a481a ) or ( a482a );
 a10140a <=( a479a ) or ( a480a );
 a10141a <=( a10140a ) or ( a10137a );
 a10142a <=( a10141a ) or ( a10134a );
 a10143a <=( a10142a ) or ( a10129a );
 a10147a <=( a476a ) or ( a477a );
 a10148a <=( a478a ) or ( a10147a );
 a10151a <=( a474a ) or ( a475a );
 a10154a <=( a472a ) or ( a473a );
 a10155a <=( a10154a ) or ( a10151a );
 a10156a <=( a10155a ) or ( a10148a );
 a10159a <=( a470a ) or ( a471a );
 a10162a <=( a468a ) or ( a469a );
 a10163a <=( a10162a ) or ( a10159a );
 a10166a <=( a466a ) or ( a467a );
 a10169a <=( a464a ) or ( a465a );
 a10170a <=( a10169a ) or ( a10166a );
 a10171a <=( a10170a ) or ( a10163a );
 a10172a <=( a10171a ) or ( a10156a );
 a10173a <=( a10172a ) or ( a10143a );
 a10174a <=( a10173a ) or ( a10116a );
 a10175a <=( a10174a ) or ( a10059a );
 a10176a <=( a10175a ) or ( a9944a );
 a10177a <=( a10176a ) or ( a9713a );
 a10181a <=( a461a ) or ( a462a );
 a10182a <=( a463a ) or ( a10181a );
 a10185a <=( a459a ) or ( a460a );
 a10188a <=( a457a ) or ( a458a );
 a10189a <=( a10188a ) or ( a10185a );
 a10190a <=( a10189a ) or ( a10182a );
 a10194a <=( a454a ) or ( a455a );
 a10195a <=( a456a ) or ( a10194a );
 a10198a <=( a452a ) or ( a453a );
 a10201a <=( a450a ) or ( a451a );
 a10202a <=( a10201a ) or ( a10198a );
 a10203a <=( a10202a ) or ( a10195a );
 a10204a <=( a10203a ) or ( a10190a );
 a10208a <=( a447a ) or ( a448a );
 a10209a <=( a449a ) or ( a10208a );
 a10212a <=( a445a ) or ( a446a );
 a10215a <=( a443a ) or ( a444a );
 a10216a <=( a10215a ) or ( a10212a );
 a10217a <=( a10216a ) or ( a10209a );
 a10221a <=( a440a ) or ( a441a );
 a10222a <=( a442a ) or ( a10221a );
 a10225a <=( a438a ) or ( a439a );
 a10228a <=( a436a ) or ( a437a );
 a10229a <=( a10228a ) or ( a10225a );
 a10230a <=( a10229a ) or ( a10222a );
 a10231a <=( a10230a ) or ( a10217a );
 a10232a <=( a10231a ) or ( a10204a );
 a10236a <=( a433a ) or ( a434a );
 a10237a <=( a435a ) or ( a10236a );
 a10240a <=( a431a ) or ( a432a );
 a10243a <=( a429a ) or ( a430a );
 a10244a <=( a10243a ) or ( a10240a );
 a10245a <=( a10244a ) or ( a10237a );
 a10249a <=( a426a ) or ( a427a );
 a10250a <=( a428a ) or ( a10249a );
 a10253a <=( a424a ) or ( a425a );
 a10256a <=( a422a ) or ( a423a );
 a10257a <=( a10256a ) or ( a10253a );
 a10258a <=( a10257a ) or ( a10250a );
 a10259a <=( a10258a ) or ( a10245a );
 a10263a <=( a419a ) or ( a420a );
 a10264a <=( a421a ) or ( a10263a );
 a10267a <=( a417a ) or ( a418a );
 a10270a <=( a415a ) or ( a416a );
 a10271a <=( a10270a ) or ( a10267a );
 a10272a <=( a10271a ) or ( a10264a );
 a10275a <=( a413a ) or ( a414a );
 a10278a <=( a411a ) or ( a412a );
 a10279a <=( a10278a ) or ( a10275a );
 a10282a <=( a409a ) or ( a410a );
 a10285a <=( a407a ) or ( a408a );
 a10286a <=( a10285a ) or ( a10282a );
 a10287a <=( a10286a ) or ( a10279a );
 a10288a <=( a10287a ) or ( a10272a );
 a10289a <=( a10288a ) or ( a10259a );
 a10290a <=( a10289a ) or ( a10232a );
 a10294a <=( a404a ) or ( a405a );
 a10295a <=( a406a ) or ( a10294a );
 a10298a <=( a402a ) or ( a403a );
 a10301a <=( a400a ) or ( a401a );
 a10302a <=( a10301a ) or ( a10298a );
 a10303a <=( a10302a ) or ( a10295a );
 a10307a <=( a397a ) or ( a398a );
 a10308a <=( a399a ) or ( a10307a );
 a10311a <=( a395a ) or ( a396a );
 a10314a <=( a393a ) or ( a394a );
 a10315a <=( a10314a ) or ( a10311a );
 a10316a <=( a10315a ) or ( a10308a );
 a10317a <=( a10316a ) or ( a10303a );
 a10321a <=( a390a ) or ( a391a );
 a10322a <=( a392a ) or ( a10321a );
 a10325a <=( a388a ) or ( a389a );
 a10328a <=( a386a ) or ( a387a );
 a10329a <=( a10328a ) or ( a10325a );
 a10330a <=( a10329a ) or ( a10322a );
 a10333a <=( a384a ) or ( a385a );
 a10336a <=( a382a ) or ( a383a );
 a10337a <=( a10336a ) or ( a10333a );
 a10340a <=( a380a ) or ( a381a );
 a10343a <=( a378a ) or ( a379a );
 a10344a <=( a10343a ) or ( a10340a );
 a10345a <=( a10344a ) or ( a10337a );
 a10346a <=( a10345a ) or ( a10330a );
 a10347a <=( a10346a ) or ( a10317a );
 a10351a <=( a375a ) or ( a376a );
 a10352a <=( a377a ) or ( a10351a );
 a10355a <=( a373a ) or ( a374a );
 a10358a <=( a371a ) or ( a372a );
 a10359a <=( a10358a ) or ( a10355a );
 a10360a <=( a10359a ) or ( a10352a );
 a10364a <=( a368a ) or ( a369a );
 a10365a <=( a370a ) or ( a10364a );
 a10368a <=( a366a ) or ( a367a );
 a10371a <=( a364a ) or ( a365a );
 a10372a <=( a10371a ) or ( a10368a );
 a10373a <=( a10372a ) or ( a10365a );
 a10374a <=( a10373a ) or ( a10360a );
 a10378a <=( a361a ) or ( a362a );
 a10379a <=( a363a ) or ( a10378a );
 a10382a <=( a359a ) or ( a360a );
 a10385a <=( a357a ) or ( a358a );
 a10386a <=( a10385a ) or ( a10382a );
 a10387a <=( a10386a ) or ( a10379a );
 a10390a <=( a355a ) or ( a356a );
 a10393a <=( a353a ) or ( a354a );
 a10394a <=( a10393a ) or ( a10390a );
 a10397a <=( a351a ) or ( a352a );
 a10400a <=( a349a ) or ( a350a );
 a10401a <=( a10400a ) or ( a10397a );
 a10402a <=( a10401a ) or ( a10394a );
 a10403a <=( a10402a ) or ( a10387a );
 a10404a <=( a10403a ) or ( a10374a );
 a10405a <=( a10404a ) or ( a10347a );
 a10406a <=( a10405a ) or ( a10290a );
 a10410a <=( a346a ) or ( a347a );
 a10411a <=( a348a ) or ( a10410a );
 a10414a <=( a344a ) or ( a345a );
 a10417a <=( a342a ) or ( a343a );
 a10418a <=( a10417a ) or ( a10414a );
 a10419a <=( a10418a ) or ( a10411a );
 a10423a <=( a339a ) or ( a340a );
 a10424a <=( a341a ) or ( a10423a );
 a10427a <=( a337a ) or ( a338a );
 a10430a <=( a335a ) or ( a336a );
 a10431a <=( a10430a ) or ( a10427a );
 a10432a <=( a10431a ) or ( a10424a );
 a10433a <=( a10432a ) or ( a10419a );
 a10437a <=( a332a ) or ( a333a );
 a10438a <=( a334a ) or ( a10437a );
 a10441a <=( a330a ) or ( a331a );
 a10444a <=( a328a ) or ( a329a );
 a10445a <=( a10444a ) or ( a10441a );
 a10446a <=( a10445a ) or ( a10438a );
 a10449a <=( a326a ) or ( a327a );
 a10452a <=( a324a ) or ( a325a );
 a10453a <=( a10452a ) or ( a10449a );
 a10456a <=( a322a ) or ( a323a );
 a10459a <=( a320a ) or ( a321a );
 a10460a <=( a10459a ) or ( a10456a );
 a10461a <=( a10460a ) or ( a10453a );
 a10462a <=( a10461a ) or ( a10446a );
 a10463a <=( a10462a ) or ( a10433a );
 a10467a <=( a317a ) or ( a318a );
 a10468a <=( a319a ) or ( a10467a );
 a10471a <=( a315a ) or ( a316a );
 a10474a <=( a313a ) or ( a314a );
 a10475a <=( a10474a ) or ( a10471a );
 a10476a <=( a10475a ) or ( a10468a );
 a10480a <=( a310a ) or ( a311a );
 a10481a <=( a312a ) or ( a10480a );
 a10484a <=( a308a ) or ( a309a );
 a10487a <=( a306a ) or ( a307a );
 a10488a <=( a10487a ) or ( a10484a );
 a10489a <=( a10488a ) or ( a10481a );
 a10490a <=( a10489a ) or ( a10476a );
 a10494a <=( a303a ) or ( a304a );
 a10495a <=( a305a ) or ( a10494a );
 a10498a <=( a301a ) or ( a302a );
 a10501a <=( a299a ) or ( a300a );
 a10502a <=( a10501a ) or ( a10498a );
 a10503a <=( a10502a ) or ( a10495a );
 a10506a <=( a297a ) or ( a298a );
 a10509a <=( a295a ) or ( a296a );
 a10510a <=( a10509a ) or ( a10506a );
 a10513a <=( a293a ) or ( a294a );
 a10516a <=( a291a ) or ( a292a );
 a10517a <=( a10516a ) or ( a10513a );
 a10518a <=( a10517a ) or ( a10510a );
 a10519a <=( a10518a ) or ( a10503a );
 a10520a <=( a10519a ) or ( a10490a );
 a10521a <=( a10520a ) or ( a10463a );
 a10525a <=( a288a ) or ( a289a );
 a10526a <=( a290a ) or ( a10525a );
 a10529a <=( a286a ) or ( a287a );
 a10532a <=( a284a ) or ( a285a );
 a10533a <=( a10532a ) or ( a10529a );
 a10534a <=( a10533a ) or ( a10526a );
 a10538a <=( a281a ) or ( a282a );
 a10539a <=( a283a ) or ( a10538a );
 a10542a <=( a279a ) or ( a280a );
 a10545a <=( a277a ) or ( a278a );
 a10546a <=( a10545a ) or ( a10542a );
 a10547a <=( a10546a ) or ( a10539a );
 a10548a <=( a10547a ) or ( a10534a );
 a10552a <=( a274a ) or ( a275a );
 a10553a <=( a276a ) or ( a10552a );
 a10556a <=( a272a ) or ( a273a );
 a10559a <=( a270a ) or ( a271a );
 a10560a <=( a10559a ) or ( a10556a );
 a10561a <=( a10560a ) or ( a10553a );
 a10564a <=( a268a ) or ( a269a );
 a10567a <=( a266a ) or ( a267a );
 a10568a <=( a10567a ) or ( a10564a );
 a10571a <=( a264a ) or ( a265a );
 a10574a <=( a262a ) or ( a263a );
 a10575a <=( a10574a ) or ( a10571a );
 a10576a <=( a10575a ) or ( a10568a );
 a10577a <=( a10576a ) or ( a10561a );
 a10578a <=( a10577a ) or ( a10548a );
 a10582a <=( a259a ) or ( a260a );
 a10583a <=( a261a ) or ( a10582a );
 a10586a <=( a257a ) or ( a258a );
 a10589a <=( a255a ) or ( a256a );
 a10590a <=( a10589a ) or ( a10586a );
 a10591a <=( a10590a ) or ( a10583a );
 a10595a <=( a252a ) or ( a253a );
 a10596a <=( a254a ) or ( a10595a );
 a10599a <=( a250a ) or ( a251a );
 a10602a <=( a248a ) or ( a249a );
 a10603a <=( a10602a ) or ( a10599a );
 a10604a <=( a10603a ) or ( a10596a );
 a10605a <=( a10604a ) or ( a10591a );
 a10609a <=( a245a ) or ( a246a );
 a10610a <=( a247a ) or ( a10609a );
 a10613a <=( a243a ) or ( a244a );
 a10616a <=( a241a ) or ( a242a );
 a10617a <=( a10616a ) or ( a10613a );
 a10618a <=( a10617a ) or ( a10610a );
 a10621a <=( a239a ) or ( a240a );
 a10624a <=( a237a ) or ( a238a );
 a10625a <=( a10624a ) or ( a10621a );
 a10628a <=( a235a ) or ( a236a );
 a10631a <=( a233a ) or ( a234a );
 a10632a <=( a10631a ) or ( a10628a );
 a10633a <=( a10632a ) or ( a10625a );
 a10634a <=( a10633a ) or ( a10618a );
 a10635a <=( a10634a ) or ( a10605a );
 a10636a <=( a10635a ) or ( a10578a );
 a10637a <=( a10636a ) or ( a10521a );
 a10638a <=( a10637a ) or ( a10406a );
 a10642a <=( a230a ) or ( a231a );
 a10643a <=( a232a ) or ( a10642a );
 a10646a <=( a228a ) or ( a229a );
 a10649a <=( a226a ) or ( a227a );
 a10650a <=( a10649a ) or ( a10646a );
 a10651a <=( a10650a ) or ( a10643a );
 a10655a <=( a223a ) or ( a224a );
 a10656a <=( a225a ) or ( a10655a );
 a10659a <=( a221a ) or ( a222a );
 a10662a <=( a219a ) or ( a220a );
 a10663a <=( a10662a ) or ( a10659a );
 a10664a <=( a10663a ) or ( a10656a );
 a10665a <=( a10664a ) or ( a10651a );
 a10669a <=( a216a ) or ( a217a );
 a10670a <=( a218a ) or ( a10669a );
 a10673a <=( a214a ) or ( a215a );
 a10676a <=( a212a ) or ( a213a );
 a10677a <=( a10676a ) or ( a10673a );
 a10678a <=( a10677a ) or ( a10670a );
 a10681a <=( a210a ) or ( a211a );
 a10684a <=( a208a ) or ( a209a );
 a10685a <=( a10684a ) or ( a10681a );
 a10688a <=( a206a ) or ( a207a );
 a10691a <=( a204a ) or ( a205a );
 a10692a <=( a10691a ) or ( a10688a );
 a10693a <=( a10692a ) or ( a10685a );
 a10694a <=( a10693a ) or ( a10678a );
 a10695a <=( a10694a ) or ( a10665a );
 a10699a <=( a201a ) or ( a202a );
 a10700a <=( a203a ) or ( a10699a );
 a10703a <=( a199a ) or ( a200a );
 a10706a <=( a197a ) or ( a198a );
 a10707a <=( a10706a ) or ( a10703a );
 a10708a <=( a10707a ) or ( a10700a );
 a10712a <=( a194a ) or ( a195a );
 a10713a <=( a196a ) or ( a10712a );
 a10716a <=( a192a ) or ( a193a );
 a10719a <=( a190a ) or ( a191a );
 a10720a <=( a10719a ) or ( a10716a );
 a10721a <=( a10720a ) or ( a10713a );
 a10722a <=( a10721a ) or ( a10708a );
 a10726a <=( a187a ) or ( a188a );
 a10727a <=( a189a ) or ( a10726a );
 a10730a <=( a185a ) or ( a186a );
 a10733a <=( a183a ) or ( a184a );
 a10734a <=( a10733a ) or ( a10730a );
 a10735a <=( a10734a ) or ( a10727a );
 a10738a <=( a181a ) or ( a182a );
 a10741a <=( a179a ) or ( a180a );
 a10742a <=( a10741a ) or ( a10738a );
 a10745a <=( a177a ) or ( a178a );
 a10748a <=( a175a ) or ( a176a );
 a10749a <=( a10748a ) or ( a10745a );
 a10750a <=( a10749a ) or ( a10742a );
 a10751a <=( a10750a ) or ( a10735a );
 a10752a <=( a10751a ) or ( a10722a );
 a10753a <=( a10752a ) or ( a10695a );
 a10757a <=( a172a ) or ( a173a );
 a10758a <=( a174a ) or ( a10757a );
 a10761a <=( a170a ) or ( a171a );
 a10764a <=( a168a ) or ( a169a );
 a10765a <=( a10764a ) or ( a10761a );
 a10766a <=( a10765a ) or ( a10758a );
 a10770a <=( a165a ) or ( a166a );
 a10771a <=( a167a ) or ( a10770a );
 a10774a <=( a163a ) or ( a164a );
 a10777a <=( a161a ) or ( a162a );
 a10778a <=( a10777a ) or ( a10774a );
 a10779a <=( a10778a ) or ( a10771a );
 a10780a <=( a10779a ) or ( a10766a );
 a10784a <=( a158a ) or ( a159a );
 a10785a <=( a160a ) or ( a10784a );
 a10788a <=( a156a ) or ( a157a );
 a10791a <=( a154a ) or ( a155a );
 a10792a <=( a10791a ) or ( a10788a );
 a10793a <=( a10792a ) or ( a10785a );
 a10796a <=( a152a ) or ( a153a );
 a10799a <=( a150a ) or ( a151a );
 a10800a <=( a10799a ) or ( a10796a );
 a10803a <=( a148a ) or ( a149a );
 a10806a <=( a146a ) or ( a147a );
 a10807a <=( a10806a ) or ( a10803a );
 a10808a <=( a10807a ) or ( a10800a );
 a10809a <=( a10808a ) or ( a10793a );
 a10810a <=( a10809a ) or ( a10780a );
 a10814a <=( a143a ) or ( a144a );
 a10815a <=( a145a ) or ( a10814a );
 a10818a <=( a141a ) or ( a142a );
 a10821a <=( a139a ) or ( a140a );
 a10822a <=( a10821a ) or ( a10818a );
 a10823a <=( a10822a ) or ( a10815a );
 a10827a <=( a136a ) or ( a137a );
 a10828a <=( a138a ) or ( a10827a );
 a10831a <=( a134a ) or ( a135a );
 a10834a <=( a132a ) or ( a133a );
 a10835a <=( a10834a ) or ( a10831a );
 a10836a <=( a10835a ) or ( a10828a );
 a10837a <=( a10836a ) or ( a10823a );
 a10841a <=( a129a ) or ( a130a );
 a10842a <=( a131a ) or ( a10841a );
 a10845a <=( a127a ) or ( a128a );
 a10848a <=( a125a ) or ( a126a );
 a10849a <=( a10848a ) or ( a10845a );
 a10850a <=( a10849a ) or ( a10842a );
 a10853a <=( a123a ) or ( a124a );
 a10856a <=( a121a ) or ( a122a );
 a10857a <=( a10856a ) or ( a10853a );
 a10860a <=( a119a ) or ( a120a );
 a10863a <=( a117a ) or ( a118a );
 a10864a <=( a10863a ) or ( a10860a );
 a10865a <=( a10864a ) or ( a10857a );
 a10866a <=( a10865a ) or ( a10850a );
 a10867a <=( a10866a ) or ( a10837a );
 a10868a <=( a10867a ) or ( a10810a );
 a10869a <=( a10868a ) or ( a10753a );
 a10873a <=( a114a ) or ( a115a );
 a10874a <=( a116a ) or ( a10873a );
 a10877a <=( a112a ) or ( a113a );
 a10880a <=( a110a ) or ( a111a );
 a10881a <=( a10880a ) or ( a10877a );
 a10882a <=( a10881a ) or ( a10874a );
 a10886a <=( a107a ) or ( a108a );
 a10887a <=( a109a ) or ( a10886a );
 a10890a <=( a105a ) or ( a106a );
 a10893a <=( a103a ) or ( a104a );
 a10894a <=( a10893a ) or ( a10890a );
 a10895a <=( a10894a ) or ( a10887a );
 a10896a <=( a10895a ) or ( a10882a );
 a10900a <=( a100a ) or ( a101a );
 a10901a <=( a102a ) or ( a10900a );
 a10904a <=( a98a ) or ( a99a );
 a10907a <=( a96a ) or ( a97a );
 a10908a <=( a10907a ) or ( a10904a );
 a10909a <=( a10908a ) or ( a10901a );
 a10912a <=( a94a ) or ( a95a );
 a10915a <=( a92a ) or ( a93a );
 a10916a <=( a10915a ) or ( a10912a );
 a10919a <=( a90a ) or ( a91a );
 a10922a <=( a88a ) or ( a89a );
 a10923a <=( a10922a ) or ( a10919a );
 a10924a <=( a10923a ) or ( a10916a );
 a10925a <=( a10924a ) or ( a10909a );
 a10926a <=( a10925a ) or ( a10896a );
 a10930a <=( a85a ) or ( a86a );
 a10931a <=( a87a ) or ( a10930a );
 a10934a <=( a83a ) or ( a84a );
 a10937a <=( a81a ) or ( a82a );
 a10938a <=( a10937a ) or ( a10934a );
 a10939a <=( a10938a ) or ( a10931a );
 a10943a <=( a78a ) or ( a79a );
 a10944a <=( a80a ) or ( a10943a );
 a10947a <=( a76a ) or ( a77a );
 a10950a <=( a74a ) or ( a75a );
 a10951a <=( a10950a ) or ( a10947a );
 a10952a <=( a10951a ) or ( a10944a );
 a10953a <=( a10952a ) or ( a10939a );
 a10957a <=( a71a ) or ( a72a );
 a10958a <=( a73a ) or ( a10957a );
 a10961a <=( a69a ) or ( a70a );
 a10964a <=( a67a ) or ( a68a );
 a10965a <=( a10964a ) or ( a10961a );
 a10966a <=( a10965a ) or ( a10958a );
 a10969a <=( a65a ) or ( a66a );
 a10972a <=( a63a ) or ( a64a );
 a10973a <=( a10972a ) or ( a10969a );
 a10976a <=( a61a ) or ( a62a );
 a10979a <=( a59a ) or ( a60a );
 a10980a <=( a10979a ) or ( a10976a );
 a10981a <=( a10980a ) or ( a10973a );
 a10982a <=( a10981a ) or ( a10966a );
 a10983a <=( a10982a ) or ( a10953a );
 a10984a <=( a10983a ) or ( a10926a );
 a10988a <=( a56a ) or ( a57a );
 a10989a <=( a58a ) or ( a10988a );
 a10992a <=( a54a ) or ( a55a );
 a10995a <=( a52a ) or ( a53a );
 a10996a <=( a10995a ) or ( a10992a );
 a10997a <=( a10996a ) or ( a10989a );
 a11001a <=( a49a ) or ( a50a );
 a11002a <=( a51a ) or ( a11001a );
 a11005a <=( a47a ) or ( a48a );
 a11008a <=( a45a ) or ( a46a );
 a11009a <=( a11008a ) or ( a11005a );
 a11010a <=( a11009a ) or ( a11002a );
 a11011a <=( a11010a ) or ( a10997a );
 a11015a <=( a42a ) or ( a43a );
 a11016a <=( a44a ) or ( a11015a );
 a11019a <=( a40a ) or ( a41a );
 a11022a <=( a38a ) or ( a39a );
 a11023a <=( a11022a ) or ( a11019a );
 a11024a <=( a11023a ) or ( a11016a );
 a11027a <=( a36a ) or ( a37a );
 a11030a <=( a34a ) or ( a35a );
 a11031a <=( a11030a ) or ( a11027a );
 a11034a <=( a32a ) or ( a33a );
 a11037a <=( a30a ) or ( a31a );
 a11038a <=( a11037a ) or ( a11034a );
 a11039a <=( a11038a ) or ( a11031a );
 a11040a <=( a11039a ) or ( a11024a );
 a11041a <=( a11040a ) or ( a11011a );
 a11045a <=( a27a ) or ( a28a );
 a11046a <=( a29a ) or ( a11045a );
 a11049a <=( a25a ) or ( a26a );
 a11052a <=( a23a ) or ( a24a );
 a11053a <=( a11052a ) or ( a11049a );
 a11054a <=( a11053a ) or ( a11046a );
 a11058a <=( a20a ) or ( a21a );
 a11059a <=( a22a ) or ( a11058a );
 a11062a <=( a18a ) or ( a19a );
 a11065a <=( a16a ) or ( a17a );
 a11066a <=( a11065a ) or ( a11062a );
 a11067a <=( a11066a ) or ( a11059a );
 a11068a <=( a11067a ) or ( a11054a );
 a11072a <=( a13a ) or ( a14a );
 a11073a <=( a15a ) or ( a11072a );
 a11076a <=( a11a ) or ( a12a );
 a11079a <=( a9a ) or ( a10a );
 a11080a <=( a11079a ) or ( a11076a );
 a11081a <=( a11080a ) or ( a11073a );
 a11084a <=( a7a ) or ( a8a );
 a11087a <=( a5a ) or ( a6a );
 a11088a <=( a11087a ) or ( a11084a );
 a11091a <=( a3a ) or ( a4a );
 a11094a <=( a1a ) or ( a2a );
 a11095a <=( a11094a ) or ( a11091a );
 a11096a <=( a11095a ) or ( a11088a );
 a11097a <=( a11096a ) or ( a11081a );
 a11098a <=( a11097a ) or ( a11068a );
 a11099a <=( a11098a ) or ( a11041a );
 a11100a <=( a11099a ) or ( a10984a );
 a11101a <=( a11100a ) or ( a10869a );
 a11102a <=( a11101a ) or ( a10638a );
 a11103a <=( a11102a ) or ( a10177a );
 a11104a <=( a11103a ) or ( a9252a );
 a11107a <=( A200  and  (not A199) );
 a11110a <=( A202  and  A201 );
 a11111a <=( a11110a  and  a11107a );
 a11114a <=( A233  and  (not A232) );
 a11117a <=( A235  and  A234 );
 a11118a <=( a11117a  and  a11114a );
 a11121a <=( A200  and  (not A199) );
 a11124a <=( A202  and  A201 );
 a11125a <=( a11124a  and  a11121a );
 a11128a <=( A233  and  (not A232) );
 a11131a <=( A236  and  A234 );
 a11132a <=( a11131a  and  a11128a );
 a11135a <=( A200  and  (not A199) );
 a11138a <=( A202  and  A201 );
 a11139a <=( a11138a  and  a11135a );
 a11142a <=( (not A233)  and  A232 );
 a11145a <=( A235  and  A234 );
 a11146a <=( a11145a  and  a11142a );
 a11149a <=( A200  and  (not A199) );
 a11152a <=( A202  and  A201 );
 a11153a <=( a11152a  and  a11149a );
 a11156a <=( (not A233)  and  A232 );
 a11159a <=( A236  and  A234 );
 a11160a <=( a11159a  and  a11156a );
 a11163a <=( A200  and  (not A199) );
 a11166a <=( A203  and  A201 );
 a11167a <=( a11166a  and  a11163a );
 a11170a <=( A233  and  (not A232) );
 a11173a <=( A235  and  A234 );
 a11174a <=( a11173a  and  a11170a );
 a11177a <=( A200  and  (not A199) );
 a11180a <=( A203  and  A201 );
 a11181a <=( a11180a  and  a11177a );
 a11184a <=( A233  and  (not A232) );
 a11187a <=( A236  and  A234 );
 a11188a <=( a11187a  and  a11184a );
 a11191a <=( A200  and  (not A199) );
 a11194a <=( A203  and  A201 );
 a11195a <=( a11194a  and  a11191a );
 a11198a <=( (not A233)  and  A232 );
 a11201a <=( A235  and  A234 );
 a11202a <=( a11201a  and  a11198a );
 a11205a <=( A200  and  (not A199) );
 a11208a <=( A203  and  A201 );
 a11209a <=( a11208a  and  a11205a );
 a11212a <=( (not A233)  and  A232 );
 a11215a <=( A236  and  A234 );
 a11216a <=( a11215a  and  a11212a );
 a11219a <=( (not A200)  and  A199 );
 a11222a <=( A202  and  A201 );
 a11223a <=( a11222a  and  a11219a );
 a11226a <=( A233  and  (not A232) );
 a11229a <=( A235  and  A234 );
 a11230a <=( a11229a  and  a11226a );
 a11233a <=( (not A200)  and  A199 );
 a11236a <=( A202  and  A201 );
 a11237a <=( a11236a  and  a11233a );
 a11240a <=( A233  and  (not A232) );
 a11243a <=( A236  and  A234 );
 a11244a <=( a11243a  and  a11240a );
 a11247a <=( (not A200)  and  A199 );
 a11250a <=( A202  and  A201 );
 a11251a <=( a11250a  and  a11247a );
 a11254a <=( (not A233)  and  A232 );
 a11257a <=( A235  and  A234 );
 a11258a <=( a11257a  and  a11254a );
 a11261a <=( (not A200)  and  A199 );
 a11264a <=( A202  and  A201 );
 a11265a <=( a11264a  and  a11261a );
 a11268a <=( (not A233)  and  A232 );
 a11271a <=( A236  and  A234 );
 a11272a <=( a11271a  and  a11268a );
 a11275a <=( (not A200)  and  A199 );
 a11278a <=( A203  and  A201 );
 a11279a <=( a11278a  and  a11275a );
 a11282a <=( A233  and  (not A232) );
 a11285a <=( A235  and  A234 );
 a11286a <=( a11285a  and  a11282a );
 a11289a <=( (not A200)  and  A199 );
 a11292a <=( A203  and  A201 );
 a11293a <=( a11292a  and  a11289a );
 a11296a <=( A233  and  (not A232) );
 a11299a <=( A236  and  A234 );
 a11300a <=( a11299a  and  a11296a );
 a11303a <=( (not A200)  and  A199 );
 a11306a <=( A203  and  A201 );
 a11307a <=( a11306a  and  a11303a );
 a11310a <=( (not A233)  and  A232 );
 a11313a <=( A235  and  A234 );
 a11314a <=( a11313a  and  a11310a );
 a11317a <=( (not A200)  and  A199 );
 a11320a <=( A203  and  A201 );
 a11321a <=( a11320a  and  a11317a );
 a11324a <=( (not A233)  and  A232 );
 a11327a <=( A236  and  A234 );
 a11328a <=( a11327a  and  a11324a );
 a11331a <=( A168  and  (not A170) );
 a11334a <=( (not A166)  and  A167 );
 a11335a <=( a11334a  and  a11331a );
 a11338a <=( A233  and  (not A232) );
 a11341a <=( A235  and  A234 );
 a11342a <=( a11341a  and  a11338a );
 a11345a <=( A168  and  (not A170) );
 a11348a <=( (not A166)  and  A167 );
 a11349a <=( a11348a  and  a11345a );
 a11352a <=( A233  and  (not A232) );
 a11355a <=( A236  and  A234 );
 a11356a <=( a11355a  and  a11352a );
 a11359a <=( A168  and  (not A170) );
 a11362a <=( (not A166)  and  A167 );
 a11363a <=( a11362a  and  a11359a );
 a11366a <=( (not A233)  and  A232 );
 a11369a <=( A235  and  A234 );
 a11370a <=( a11369a  and  a11366a );
 a11373a <=( A168  and  (not A170) );
 a11376a <=( (not A166)  and  A167 );
 a11377a <=( a11376a  and  a11373a );
 a11380a <=( (not A233)  and  A232 );
 a11383a <=( A236  and  A234 );
 a11384a <=( a11383a  and  a11380a );
 a11387a <=( A168  and  (not A170) );
 a11390a <=( A166  and  (not A167) );
 a11391a <=( a11390a  and  a11387a );
 a11394a <=( A233  and  (not A232) );
 a11397a <=( A235  and  A234 );
 a11398a <=( a11397a  and  a11394a );
 a11401a <=( A168  and  (not A170) );
 a11404a <=( A166  and  (not A167) );
 a11405a <=( a11404a  and  a11401a );
 a11408a <=( A233  and  (not A232) );
 a11411a <=( A236  and  A234 );
 a11412a <=( a11411a  and  a11408a );
 a11415a <=( A168  and  (not A170) );
 a11418a <=( A166  and  (not A167) );
 a11419a <=( a11418a  and  a11415a );
 a11422a <=( (not A233)  and  A232 );
 a11425a <=( A235  and  A234 );
 a11426a <=( a11425a  and  a11422a );
 a11429a <=( A168  and  (not A170) );
 a11432a <=( A166  and  (not A167) );
 a11433a <=( a11432a  and  a11429a );
 a11436a <=( (not A233)  and  A232 );
 a11439a <=( A236  and  A234 );
 a11440a <=( a11439a  and  a11436a );
 a11443a <=( A168  and  A169 );
 a11446a <=( (not A166)  and  A167 );
 a11447a <=( a11446a  and  a11443a );
 a11450a <=( A233  and  (not A232) );
 a11453a <=( A235  and  A234 );
 a11454a <=( a11453a  and  a11450a );
 a11457a <=( A168  and  A169 );
 a11460a <=( (not A166)  and  A167 );
 a11461a <=( a11460a  and  a11457a );
 a11464a <=( A233  and  (not A232) );
 a11467a <=( A236  and  A234 );
 a11468a <=( a11467a  and  a11464a );
 a11471a <=( A168  and  A169 );
 a11474a <=( (not A166)  and  A167 );
 a11475a <=( a11474a  and  a11471a );
 a11478a <=( (not A233)  and  A232 );
 a11481a <=( A235  and  A234 );
 a11482a <=( a11481a  and  a11478a );
 a11485a <=( A168  and  A169 );
 a11488a <=( (not A166)  and  A167 );
 a11489a <=( a11488a  and  a11485a );
 a11492a <=( (not A233)  and  A232 );
 a11495a <=( A236  and  A234 );
 a11496a <=( a11495a  and  a11492a );
 a11499a <=( A168  and  A169 );
 a11502a <=( A166  and  (not A167) );
 a11503a <=( a11502a  and  a11499a );
 a11506a <=( A233  and  (not A232) );
 a11509a <=( A235  and  A234 );
 a11510a <=( a11509a  and  a11506a );
 a11513a <=( A168  and  A169 );
 a11516a <=( A166  and  (not A167) );
 a11517a <=( a11516a  and  a11513a );
 a11520a <=( A233  and  (not A232) );
 a11523a <=( A236  and  A234 );
 a11524a <=( a11523a  and  a11520a );
 a11527a <=( A168  and  A169 );
 a11530a <=( A166  and  (not A167) );
 a11531a <=( a11530a  and  a11527a );
 a11534a <=( (not A233)  and  A232 );
 a11537a <=( A235  and  A234 );
 a11538a <=( a11537a  and  a11534a );
 a11541a <=( A168  and  A169 );
 a11544a <=( A166  and  (not A167) );
 a11545a <=( a11544a  and  a11541a );
 a11548a <=( (not A233)  and  A232 );
 a11551a <=( A236  and  A234 );
 a11552a <=( a11551a  and  a11548a );
 a11555a <=( A200  and  (not A199) );
 a11558a <=( A202  and  A201 );
 a11559a <=( a11558a  and  a11555a );
 a11562a <=( A233  and  (not A232) );
 a11566a <=( (not A236)  and  (not A235) );
 a11567a <=( (not A234)  and  a11566a );
 a11568a <=( a11567a  and  a11562a );
 a11571a <=( A200  and  (not A199) );
 a11574a <=( A202  and  A201 );
 a11575a <=( a11574a  and  a11571a );
 a11578a <=( (not A233)  and  A232 );
 a11582a <=( (not A236)  and  (not A235) );
 a11583a <=( (not A234)  and  a11582a );
 a11584a <=( a11583a  and  a11578a );
 a11587a <=( A200  and  (not A199) );
 a11590a <=( A203  and  A201 );
 a11591a <=( a11590a  and  a11587a );
 a11594a <=( A233  and  (not A232) );
 a11598a <=( (not A236)  and  (not A235) );
 a11599a <=( (not A234)  and  a11598a );
 a11600a <=( a11599a  and  a11594a );
 a11603a <=( A200  and  (not A199) );
 a11606a <=( A203  and  A201 );
 a11607a <=( a11606a  and  a11603a );
 a11610a <=( (not A233)  and  A232 );
 a11614a <=( (not A236)  and  (not A235) );
 a11615a <=( (not A234)  and  a11614a );
 a11616a <=( a11615a  and  a11610a );
 a11619a <=( A200  and  (not A199) );
 a11622a <=( (not A202)  and  (not A201) );
 a11623a <=( a11622a  and  a11619a );
 a11626a <=( (not A232)  and  (not A203) );
 a11630a <=( A235  and  A234 );
 a11631a <=( A233  and  a11630a );
 a11632a <=( a11631a  and  a11626a );
 a11635a <=( A200  and  (not A199) );
 a11638a <=( (not A202)  and  (not A201) );
 a11639a <=( a11638a  and  a11635a );
 a11642a <=( (not A232)  and  (not A203) );
 a11646a <=( A236  and  A234 );
 a11647a <=( A233  and  a11646a );
 a11648a <=( a11647a  and  a11642a );
 a11651a <=( A200  and  (not A199) );
 a11654a <=( (not A202)  and  (not A201) );
 a11655a <=( a11654a  and  a11651a );
 a11658a <=( A232  and  (not A203) );
 a11662a <=( A235  and  A234 );
 a11663a <=( (not A233)  and  a11662a );
 a11664a <=( a11663a  and  a11658a );
 a11667a <=( A200  and  (not A199) );
 a11670a <=( (not A202)  and  (not A201) );
 a11671a <=( a11670a  and  a11667a );
 a11674a <=( A232  and  (not A203) );
 a11678a <=( A236  and  A234 );
 a11679a <=( (not A233)  and  a11678a );
 a11680a <=( a11679a  and  a11674a );
 a11683a <=( (not A200)  and  A199 );
 a11686a <=( A202  and  A201 );
 a11687a <=( a11686a  and  a11683a );
 a11690a <=( A233  and  (not A232) );
 a11694a <=( (not A236)  and  (not A235) );
 a11695a <=( (not A234)  and  a11694a );
 a11696a <=( a11695a  and  a11690a );
 a11699a <=( (not A200)  and  A199 );
 a11702a <=( A202  and  A201 );
 a11703a <=( a11702a  and  a11699a );
 a11706a <=( (not A233)  and  A232 );
 a11710a <=( (not A236)  and  (not A235) );
 a11711a <=( (not A234)  and  a11710a );
 a11712a <=( a11711a  and  a11706a );
 a11715a <=( (not A200)  and  A199 );
 a11718a <=( A203  and  A201 );
 a11719a <=( a11718a  and  a11715a );
 a11722a <=( A233  and  (not A232) );
 a11726a <=( (not A236)  and  (not A235) );
 a11727a <=( (not A234)  and  a11726a );
 a11728a <=( a11727a  and  a11722a );
 a11731a <=( (not A200)  and  A199 );
 a11734a <=( A203  and  A201 );
 a11735a <=( a11734a  and  a11731a );
 a11738a <=( (not A233)  and  A232 );
 a11742a <=( (not A236)  and  (not A235) );
 a11743a <=( (not A234)  and  a11742a );
 a11744a <=( a11743a  and  a11738a );
 a11747a <=( (not A200)  and  A199 );
 a11750a <=( (not A202)  and  (not A201) );
 a11751a <=( a11750a  and  a11747a );
 a11754a <=( (not A232)  and  (not A203) );
 a11758a <=( A235  and  A234 );
 a11759a <=( A233  and  a11758a );
 a11760a <=( a11759a  and  a11754a );
 a11763a <=( (not A200)  and  A199 );
 a11766a <=( (not A202)  and  (not A201) );
 a11767a <=( a11766a  and  a11763a );
 a11770a <=( (not A232)  and  (not A203) );
 a11774a <=( A236  and  A234 );
 a11775a <=( A233  and  a11774a );
 a11776a <=( a11775a  and  a11770a );
 a11779a <=( (not A200)  and  A199 );
 a11782a <=( (not A202)  and  (not A201) );
 a11783a <=( a11782a  and  a11779a );
 a11786a <=( A232  and  (not A203) );
 a11790a <=( A235  and  A234 );
 a11791a <=( (not A233)  and  a11790a );
 a11792a <=( a11791a  and  a11786a );
 a11795a <=( (not A200)  and  A199 );
 a11798a <=( (not A202)  and  (not A201) );
 a11799a <=( a11798a  and  a11795a );
 a11802a <=( A232  and  (not A203) );
 a11806a <=( A236  and  A234 );
 a11807a <=( (not A233)  and  a11806a );
 a11808a <=( a11807a  and  a11802a );
 a11811a <=( A168  and  (not A170) );
 a11814a <=( (not A166)  and  A167 );
 a11815a <=( a11814a  and  a11811a );
 a11818a <=( A233  and  (not A232) );
 a11822a <=( (not A236)  and  (not A235) );
 a11823a <=( (not A234)  and  a11822a );
 a11824a <=( a11823a  and  a11818a );
 a11827a <=( A168  and  (not A170) );
 a11830a <=( (not A166)  and  A167 );
 a11831a <=( a11830a  and  a11827a );
 a11834a <=( (not A233)  and  A232 );
 a11838a <=( (not A236)  and  (not A235) );
 a11839a <=( (not A234)  and  a11838a );
 a11840a <=( a11839a  and  a11834a );
 a11843a <=( A168  and  (not A170) );
 a11846a <=( A166  and  (not A167) );
 a11847a <=( a11846a  and  a11843a );
 a11850a <=( A233  and  (not A232) );
 a11854a <=( (not A236)  and  (not A235) );
 a11855a <=( (not A234)  and  a11854a );
 a11856a <=( a11855a  and  a11850a );
 a11859a <=( A168  and  (not A170) );
 a11862a <=( A166  and  (not A167) );
 a11863a <=( a11862a  and  a11859a );
 a11866a <=( (not A233)  and  A232 );
 a11870a <=( (not A236)  and  (not A235) );
 a11871a <=( (not A234)  and  a11870a );
 a11872a <=( a11871a  and  a11866a );
 a11875a <=( A168  and  A169 );
 a11878a <=( (not A166)  and  A167 );
 a11879a <=( a11878a  and  a11875a );
 a11882a <=( A233  and  (not A232) );
 a11886a <=( (not A236)  and  (not A235) );
 a11887a <=( (not A234)  and  a11886a );
 a11888a <=( a11887a  and  a11882a );
 a11891a <=( A168  and  A169 );
 a11894a <=( (not A166)  and  A167 );
 a11895a <=( a11894a  and  a11891a );
 a11898a <=( (not A233)  and  A232 );
 a11902a <=( (not A236)  and  (not A235) );
 a11903a <=( (not A234)  and  a11902a );
 a11904a <=( a11903a  and  a11898a );
 a11907a <=( A168  and  A169 );
 a11910a <=( A166  and  (not A167) );
 a11911a <=( a11910a  and  a11907a );
 a11914a <=( A233  and  (not A232) );
 a11918a <=( (not A236)  and  (not A235) );
 a11919a <=( (not A234)  and  a11918a );
 a11920a <=( a11919a  and  a11914a );
 a11923a <=( A168  and  A169 );
 a11926a <=( A166  and  (not A167) );
 a11927a <=( a11926a  and  a11923a );
 a11930a <=( (not A233)  and  A232 );
 a11934a <=( (not A236)  and  (not A235) );
 a11935a <=( (not A234)  and  a11934a );
 a11936a <=( a11935a  and  a11930a );
 a11939a <=( (not A169)  and  A170 );
 a11942a <=( A167  and  (not A168) );
 a11943a <=( a11942a  and  a11939a );
 a11946a <=( (not A232)  and  (not A166) );
 a11950a <=( A235  and  A234 );
 a11951a <=( A233  and  a11950a );
 a11952a <=( a11951a  and  a11946a );
 a11955a <=( (not A169)  and  A170 );
 a11958a <=( A167  and  (not A168) );
 a11959a <=( a11958a  and  a11955a );
 a11962a <=( (not A232)  and  (not A166) );
 a11966a <=( A236  and  A234 );
 a11967a <=( A233  and  a11966a );
 a11968a <=( a11967a  and  a11962a );
 a11971a <=( (not A169)  and  A170 );
 a11974a <=( A167  and  (not A168) );
 a11975a <=( a11974a  and  a11971a );
 a11978a <=( A232  and  (not A166) );
 a11982a <=( A235  and  A234 );
 a11983a <=( (not A233)  and  a11982a );
 a11984a <=( a11983a  and  a11978a );
 a11987a <=( (not A169)  and  A170 );
 a11990a <=( A167  and  (not A168) );
 a11991a <=( a11990a  and  a11987a );
 a11994a <=( A232  and  (not A166) );
 a11998a <=( A236  and  A234 );
 a11999a <=( (not A233)  and  a11998a );
 a12000a <=( a11999a  and  a11994a );
 a12003a <=( (not A169)  and  A170 );
 a12006a <=( (not A167)  and  (not A168) );
 a12007a <=( a12006a  and  a12003a );
 a12010a <=( (not A232)  and  A166 );
 a12014a <=( A235  and  A234 );
 a12015a <=( A233  and  a12014a );
 a12016a <=( a12015a  and  a12010a );
 a12019a <=( (not A169)  and  A170 );
 a12022a <=( (not A167)  and  (not A168) );
 a12023a <=( a12022a  and  a12019a );
 a12026a <=( (not A232)  and  A166 );
 a12030a <=( A236  and  A234 );
 a12031a <=( A233  and  a12030a );
 a12032a <=( a12031a  and  a12026a );
 a12035a <=( (not A169)  and  A170 );
 a12038a <=( (not A167)  and  (not A168) );
 a12039a <=( a12038a  and  a12035a );
 a12042a <=( A232  and  A166 );
 a12046a <=( A235  and  A234 );
 a12047a <=( (not A233)  and  a12046a );
 a12048a <=( a12047a  and  a12042a );
 a12051a <=( (not A169)  and  A170 );
 a12054a <=( (not A167)  and  (not A168) );
 a12055a <=( a12054a  and  a12051a );
 a12058a <=( A232  and  A166 );
 a12062a <=( A236  and  A234 );
 a12063a <=( (not A233)  and  a12062a );
 a12064a <=( a12063a  and  a12058a );
 a12067a <=( A200  and  (not A199) );
 a12071a <=( (not A203)  and  (not A202) );
 a12072a <=( (not A201)  and  a12071a );
 a12073a <=( a12072a  and  a12067a );
 a12076a <=( A233  and  (not A232) );
 a12080a <=( (not A236)  and  (not A235) );
 a12081a <=( (not A234)  and  a12080a );
 a12082a <=( a12081a  and  a12076a );
 a12085a <=( A200  and  (not A199) );
 a12089a <=( (not A203)  and  (not A202) );
 a12090a <=( (not A201)  and  a12089a );
 a12091a <=( a12090a  and  a12085a );
 a12094a <=( (not A233)  and  A232 );
 a12098a <=( (not A236)  and  (not A235) );
 a12099a <=( (not A234)  and  a12098a );
 a12100a <=( a12099a  and  a12094a );
 a12103a <=( (not A200)  and  A199 );
 a12107a <=( (not A203)  and  (not A202) );
 a12108a <=( (not A201)  and  a12107a );
 a12109a <=( a12108a  and  a12103a );
 a12112a <=( A233  and  (not A232) );
 a12116a <=( (not A236)  and  (not A235) );
 a12117a <=( (not A234)  and  a12116a );
 a12118a <=( a12117a  and  a12112a );
 a12121a <=( (not A200)  and  A199 );
 a12125a <=( (not A203)  and  (not A202) );
 a12126a <=( (not A201)  and  a12125a );
 a12127a <=( a12126a  and  a12121a );
 a12130a <=( (not A233)  and  A232 );
 a12134a <=( (not A236)  and  (not A235) );
 a12135a <=( (not A234)  and  a12134a );
 a12136a <=( a12135a  and  a12130a );
 a12139a <=( A166  and  A167 );
 a12143a <=( (not A265)  and  A202 );
 a12144a <=( (not A201)  and  a12143a );
 a12145a <=( a12144a  and  a12139a );
 a12148a <=( A267  and  A266 );
 a12152a <=( A301  and  (not A300) );
 a12153a <=( A268  and  a12152a );
 a12154a <=( a12153a  and  a12148a );
 a12157a <=( A166  and  A167 );
 a12161a <=( (not A265)  and  A202 );
 a12162a <=( (not A201)  and  a12161a );
 a12163a <=( a12162a  and  a12157a );
 a12166a <=( A267  and  A266 );
 a12170a <=( A302  and  (not A300) );
 a12171a <=( A268  and  a12170a );
 a12172a <=( a12171a  and  a12166a );
 a12175a <=( A166  and  A167 );
 a12179a <=( (not A265)  and  A202 );
 a12180a <=( (not A201)  and  a12179a );
 a12181a <=( a12180a  and  a12175a );
 a12184a <=( A267  and  A266 );
 a12188a <=( A299  and  A298 );
 a12189a <=( A268  and  a12188a );
 a12190a <=( a12189a  and  a12184a );
 a12193a <=( A166  and  A167 );
 a12197a <=( (not A265)  and  A202 );
 a12198a <=( (not A201)  and  a12197a );
 a12199a <=( a12198a  and  a12193a );
 a12202a <=( A267  and  A266 );
 a12206a <=( (not A299)  and  (not A298) );
 a12207a <=( A268  and  a12206a );
 a12208a <=( a12207a  and  a12202a );
 a12211a <=( A166  and  A167 );
 a12215a <=( (not A265)  and  A202 );
 a12216a <=( (not A201)  and  a12215a );
 a12217a <=( a12216a  and  a12211a );
 a12220a <=( A267  and  A266 );
 a12224a <=( A301  and  (not A300) );
 a12225a <=( A269  and  a12224a );
 a12226a <=( a12225a  and  a12220a );
 a12229a <=( A166  and  A167 );
 a12233a <=( (not A265)  and  A202 );
 a12234a <=( (not A201)  and  a12233a );
 a12235a <=( a12234a  and  a12229a );
 a12238a <=( A267  and  A266 );
 a12242a <=( A302  and  (not A300) );
 a12243a <=( A269  and  a12242a );
 a12244a <=( a12243a  and  a12238a );
 a12247a <=( A166  and  A167 );
 a12251a <=( (not A265)  and  A202 );
 a12252a <=( (not A201)  and  a12251a );
 a12253a <=( a12252a  and  a12247a );
 a12256a <=( A267  and  A266 );
 a12260a <=( A299  and  A298 );
 a12261a <=( A269  and  a12260a );
 a12262a <=( a12261a  and  a12256a );
 a12265a <=( A166  and  A167 );
 a12269a <=( (not A265)  and  A202 );
 a12270a <=( (not A201)  and  a12269a );
 a12271a <=( a12270a  and  a12265a );
 a12274a <=( A267  and  A266 );
 a12278a <=( (not A299)  and  (not A298) );
 a12279a <=( A269  and  a12278a );
 a12280a <=( a12279a  and  a12274a );
 a12283a <=( A166  and  A167 );
 a12287a <=( A265  and  A202 );
 a12288a <=( (not A201)  and  a12287a );
 a12289a <=( a12288a  and  a12283a );
 a12292a <=( A267  and  (not A266) );
 a12296a <=( A301  and  (not A300) );
 a12297a <=( A268  and  a12296a );
 a12298a <=( a12297a  and  a12292a );
 a12301a <=( A166  and  A167 );
 a12305a <=( A265  and  A202 );
 a12306a <=( (not A201)  and  a12305a );
 a12307a <=( a12306a  and  a12301a );
 a12310a <=( A267  and  (not A266) );
 a12314a <=( A302  and  (not A300) );
 a12315a <=( A268  and  a12314a );
 a12316a <=( a12315a  and  a12310a );
 a12319a <=( A166  and  A167 );
 a12323a <=( A265  and  A202 );
 a12324a <=( (not A201)  and  a12323a );
 a12325a <=( a12324a  and  a12319a );
 a12328a <=( A267  and  (not A266) );
 a12332a <=( A299  and  A298 );
 a12333a <=( A268  and  a12332a );
 a12334a <=( a12333a  and  a12328a );
 a12337a <=( A166  and  A167 );
 a12341a <=( A265  and  A202 );
 a12342a <=( (not A201)  and  a12341a );
 a12343a <=( a12342a  and  a12337a );
 a12346a <=( A267  and  (not A266) );
 a12350a <=( (not A299)  and  (not A298) );
 a12351a <=( A268  and  a12350a );
 a12352a <=( a12351a  and  a12346a );
 a12355a <=( A166  and  A167 );
 a12359a <=( A265  and  A202 );
 a12360a <=( (not A201)  and  a12359a );
 a12361a <=( a12360a  and  a12355a );
 a12364a <=( A267  and  (not A266) );
 a12368a <=( A301  and  (not A300) );
 a12369a <=( A269  and  a12368a );
 a12370a <=( a12369a  and  a12364a );
 a12373a <=( A166  and  A167 );
 a12377a <=( A265  and  A202 );
 a12378a <=( (not A201)  and  a12377a );
 a12379a <=( a12378a  and  a12373a );
 a12382a <=( A267  and  (not A266) );
 a12386a <=( A302  and  (not A300) );
 a12387a <=( A269  and  a12386a );
 a12388a <=( a12387a  and  a12382a );
 a12391a <=( A166  and  A167 );
 a12395a <=( A265  and  A202 );
 a12396a <=( (not A201)  and  a12395a );
 a12397a <=( a12396a  and  a12391a );
 a12400a <=( A267  and  (not A266) );
 a12404a <=( A299  and  A298 );
 a12405a <=( A269  and  a12404a );
 a12406a <=( a12405a  and  a12400a );
 a12409a <=( A166  and  A167 );
 a12413a <=( A265  and  A202 );
 a12414a <=( (not A201)  and  a12413a );
 a12415a <=( a12414a  and  a12409a );
 a12418a <=( A267  and  (not A266) );
 a12422a <=( (not A299)  and  (not A298) );
 a12423a <=( A269  and  a12422a );
 a12424a <=( a12423a  and  a12418a );
 a12427a <=( A166  and  A167 );
 a12431a <=( (not A265)  and  A203 );
 a12432a <=( (not A201)  and  a12431a );
 a12433a <=( a12432a  and  a12427a );
 a12436a <=( A267  and  A266 );
 a12440a <=( A301  and  (not A300) );
 a12441a <=( A268  and  a12440a );
 a12442a <=( a12441a  and  a12436a );
 a12445a <=( A166  and  A167 );
 a12449a <=( (not A265)  and  A203 );
 a12450a <=( (not A201)  and  a12449a );
 a12451a <=( a12450a  and  a12445a );
 a12454a <=( A267  and  A266 );
 a12458a <=( A302  and  (not A300) );
 a12459a <=( A268  and  a12458a );
 a12460a <=( a12459a  and  a12454a );
 a12463a <=( A166  and  A167 );
 a12467a <=( (not A265)  and  A203 );
 a12468a <=( (not A201)  and  a12467a );
 a12469a <=( a12468a  and  a12463a );
 a12472a <=( A267  and  A266 );
 a12476a <=( A299  and  A298 );
 a12477a <=( A268  and  a12476a );
 a12478a <=( a12477a  and  a12472a );
 a12481a <=( A166  and  A167 );
 a12485a <=( (not A265)  and  A203 );
 a12486a <=( (not A201)  and  a12485a );
 a12487a <=( a12486a  and  a12481a );
 a12490a <=( A267  and  A266 );
 a12494a <=( (not A299)  and  (not A298) );
 a12495a <=( A268  and  a12494a );
 a12496a <=( a12495a  and  a12490a );
 a12499a <=( A166  and  A167 );
 a12503a <=( (not A265)  and  A203 );
 a12504a <=( (not A201)  and  a12503a );
 a12505a <=( a12504a  and  a12499a );
 a12508a <=( A267  and  A266 );
 a12512a <=( A301  and  (not A300) );
 a12513a <=( A269  and  a12512a );
 a12514a <=( a12513a  and  a12508a );
 a12517a <=( A166  and  A167 );
 a12521a <=( (not A265)  and  A203 );
 a12522a <=( (not A201)  and  a12521a );
 a12523a <=( a12522a  and  a12517a );
 a12526a <=( A267  and  A266 );
 a12530a <=( A302  and  (not A300) );
 a12531a <=( A269  and  a12530a );
 a12532a <=( a12531a  and  a12526a );
 a12535a <=( A166  and  A167 );
 a12539a <=( (not A265)  and  A203 );
 a12540a <=( (not A201)  and  a12539a );
 a12541a <=( a12540a  and  a12535a );
 a12544a <=( A267  and  A266 );
 a12548a <=( A299  and  A298 );
 a12549a <=( A269  and  a12548a );
 a12550a <=( a12549a  and  a12544a );
 a12553a <=( A166  and  A167 );
 a12557a <=( (not A265)  and  A203 );
 a12558a <=( (not A201)  and  a12557a );
 a12559a <=( a12558a  and  a12553a );
 a12562a <=( A267  and  A266 );
 a12566a <=( (not A299)  and  (not A298) );
 a12567a <=( A269  and  a12566a );
 a12568a <=( a12567a  and  a12562a );
 a12571a <=( A166  and  A167 );
 a12575a <=( A265  and  A203 );
 a12576a <=( (not A201)  and  a12575a );
 a12577a <=( a12576a  and  a12571a );
 a12580a <=( A267  and  (not A266) );
 a12584a <=( A301  and  (not A300) );
 a12585a <=( A268  and  a12584a );
 a12586a <=( a12585a  and  a12580a );
 a12589a <=( A166  and  A167 );
 a12593a <=( A265  and  A203 );
 a12594a <=( (not A201)  and  a12593a );
 a12595a <=( a12594a  and  a12589a );
 a12598a <=( A267  and  (not A266) );
 a12602a <=( A302  and  (not A300) );
 a12603a <=( A268  and  a12602a );
 a12604a <=( a12603a  and  a12598a );
 a12607a <=( A166  and  A167 );
 a12611a <=( A265  and  A203 );
 a12612a <=( (not A201)  and  a12611a );
 a12613a <=( a12612a  and  a12607a );
 a12616a <=( A267  and  (not A266) );
 a12620a <=( A299  and  A298 );
 a12621a <=( A268  and  a12620a );
 a12622a <=( a12621a  and  a12616a );
 a12625a <=( A166  and  A167 );
 a12629a <=( A265  and  A203 );
 a12630a <=( (not A201)  and  a12629a );
 a12631a <=( a12630a  and  a12625a );
 a12634a <=( A267  and  (not A266) );
 a12638a <=( (not A299)  and  (not A298) );
 a12639a <=( A268  and  a12638a );
 a12640a <=( a12639a  and  a12634a );
 a12643a <=( A166  and  A167 );
 a12647a <=( A265  and  A203 );
 a12648a <=( (not A201)  and  a12647a );
 a12649a <=( a12648a  and  a12643a );
 a12652a <=( A267  and  (not A266) );
 a12656a <=( A301  and  (not A300) );
 a12657a <=( A269  and  a12656a );
 a12658a <=( a12657a  and  a12652a );
 a12661a <=( A166  and  A167 );
 a12665a <=( A265  and  A203 );
 a12666a <=( (not A201)  and  a12665a );
 a12667a <=( a12666a  and  a12661a );
 a12670a <=( A267  and  (not A266) );
 a12674a <=( A302  and  (not A300) );
 a12675a <=( A269  and  a12674a );
 a12676a <=( a12675a  and  a12670a );
 a12679a <=( A166  and  A167 );
 a12683a <=( A265  and  A203 );
 a12684a <=( (not A201)  and  a12683a );
 a12685a <=( a12684a  and  a12679a );
 a12688a <=( A267  and  (not A266) );
 a12692a <=( A299  and  A298 );
 a12693a <=( A269  and  a12692a );
 a12694a <=( a12693a  and  a12688a );
 a12697a <=( A166  and  A167 );
 a12701a <=( A265  and  A203 );
 a12702a <=( (not A201)  and  a12701a );
 a12703a <=( a12702a  and  a12697a );
 a12706a <=( A267  and  (not A266) );
 a12710a <=( (not A299)  and  (not A298) );
 a12711a <=( A269  and  a12710a );
 a12712a <=( a12711a  and  a12706a );
 a12715a <=( A166  and  A167 );
 a12719a <=( (not A265)  and  A200 );
 a12720a <=( A199  and  a12719a );
 a12721a <=( a12720a  and  a12715a );
 a12724a <=( A267  and  A266 );
 a12728a <=( A301  and  (not A300) );
 a12729a <=( A268  and  a12728a );
 a12730a <=( a12729a  and  a12724a );
 a12733a <=( A166  and  A167 );
 a12737a <=( (not A265)  and  A200 );
 a12738a <=( A199  and  a12737a );
 a12739a <=( a12738a  and  a12733a );
 a12742a <=( A267  and  A266 );
 a12746a <=( A302  and  (not A300) );
 a12747a <=( A268  and  a12746a );
 a12748a <=( a12747a  and  a12742a );
 a12751a <=( A166  and  A167 );
 a12755a <=( (not A265)  and  A200 );
 a12756a <=( A199  and  a12755a );
 a12757a <=( a12756a  and  a12751a );
 a12760a <=( A267  and  A266 );
 a12764a <=( A299  and  A298 );
 a12765a <=( A268  and  a12764a );
 a12766a <=( a12765a  and  a12760a );
 a12769a <=( A166  and  A167 );
 a12773a <=( (not A265)  and  A200 );
 a12774a <=( A199  and  a12773a );
 a12775a <=( a12774a  and  a12769a );
 a12778a <=( A267  and  A266 );
 a12782a <=( (not A299)  and  (not A298) );
 a12783a <=( A268  and  a12782a );
 a12784a <=( a12783a  and  a12778a );
 a12787a <=( A166  and  A167 );
 a12791a <=( (not A265)  and  A200 );
 a12792a <=( A199  and  a12791a );
 a12793a <=( a12792a  and  a12787a );
 a12796a <=( A267  and  A266 );
 a12800a <=( A301  and  (not A300) );
 a12801a <=( A269  and  a12800a );
 a12802a <=( a12801a  and  a12796a );
 a12805a <=( A166  and  A167 );
 a12809a <=( (not A265)  and  A200 );
 a12810a <=( A199  and  a12809a );
 a12811a <=( a12810a  and  a12805a );
 a12814a <=( A267  and  A266 );
 a12818a <=( A302  and  (not A300) );
 a12819a <=( A269  and  a12818a );
 a12820a <=( a12819a  and  a12814a );
 a12823a <=( A166  and  A167 );
 a12827a <=( (not A265)  and  A200 );
 a12828a <=( A199  and  a12827a );
 a12829a <=( a12828a  and  a12823a );
 a12832a <=( A267  and  A266 );
 a12836a <=( A299  and  A298 );
 a12837a <=( A269  and  a12836a );
 a12838a <=( a12837a  and  a12832a );
 a12841a <=( A166  and  A167 );
 a12845a <=( (not A265)  and  A200 );
 a12846a <=( A199  and  a12845a );
 a12847a <=( a12846a  and  a12841a );
 a12850a <=( A267  and  A266 );
 a12854a <=( (not A299)  and  (not A298) );
 a12855a <=( A269  and  a12854a );
 a12856a <=( a12855a  and  a12850a );
 a12859a <=( A166  and  A167 );
 a12863a <=( A265  and  A200 );
 a12864a <=( A199  and  a12863a );
 a12865a <=( a12864a  and  a12859a );
 a12868a <=( A267  and  (not A266) );
 a12872a <=( A301  and  (not A300) );
 a12873a <=( A268  and  a12872a );
 a12874a <=( a12873a  and  a12868a );
 a12877a <=( A166  and  A167 );
 a12881a <=( A265  and  A200 );
 a12882a <=( A199  and  a12881a );
 a12883a <=( a12882a  and  a12877a );
 a12886a <=( A267  and  (not A266) );
 a12890a <=( A302  and  (not A300) );
 a12891a <=( A268  and  a12890a );
 a12892a <=( a12891a  and  a12886a );
 a12895a <=( A166  and  A167 );
 a12899a <=( A265  and  A200 );
 a12900a <=( A199  and  a12899a );
 a12901a <=( a12900a  and  a12895a );
 a12904a <=( A267  and  (not A266) );
 a12908a <=( A299  and  A298 );
 a12909a <=( A268  and  a12908a );
 a12910a <=( a12909a  and  a12904a );
 a12913a <=( A166  and  A167 );
 a12917a <=( A265  and  A200 );
 a12918a <=( A199  and  a12917a );
 a12919a <=( a12918a  and  a12913a );
 a12922a <=( A267  and  (not A266) );
 a12926a <=( (not A299)  and  (not A298) );
 a12927a <=( A268  and  a12926a );
 a12928a <=( a12927a  and  a12922a );
 a12931a <=( A166  and  A167 );
 a12935a <=( A265  and  A200 );
 a12936a <=( A199  and  a12935a );
 a12937a <=( a12936a  and  a12931a );
 a12940a <=( A267  and  (not A266) );
 a12944a <=( A301  and  (not A300) );
 a12945a <=( A269  and  a12944a );
 a12946a <=( a12945a  and  a12940a );
 a12949a <=( A166  and  A167 );
 a12953a <=( A265  and  A200 );
 a12954a <=( A199  and  a12953a );
 a12955a <=( a12954a  and  a12949a );
 a12958a <=( A267  and  (not A266) );
 a12962a <=( A302  and  (not A300) );
 a12963a <=( A269  and  a12962a );
 a12964a <=( a12963a  and  a12958a );
 a12967a <=( A166  and  A167 );
 a12971a <=( A265  and  A200 );
 a12972a <=( A199  and  a12971a );
 a12973a <=( a12972a  and  a12967a );
 a12976a <=( A267  and  (not A266) );
 a12980a <=( A299  and  A298 );
 a12981a <=( A269  and  a12980a );
 a12982a <=( a12981a  and  a12976a );
 a12985a <=( A166  and  A167 );
 a12989a <=( A265  and  A200 );
 a12990a <=( A199  and  a12989a );
 a12991a <=( a12990a  and  a12985a );
 a12994a <=( A267  and  (not A266) );
 a12998a <=( (not A299)  and  (not A298) );
 a12999a <=( A269  and  a12998a );
 a13000a <=( a12999a  and  a12994a );
 a13003a <=( A166  and  A167 );
 a13007a <=( (not A265)  and  (not A200) );
 a13008a <=( (not A199)  and  a13007a );
 a13009a <=( a13008a  and  a13003a );
 a13012a <=( A267  and  A266 );
 a13016a <=( A301  and  (not A300) );
 a13017a <=( A268  and  a13016a );
 a13018a <=( a13017a  and  a13012a );
 a13021a <=( A166  and  A167 );
 a13025a <=( (not A265)  and  (not A200) );
 a13026a <=( (not A199)  and  a13025a );
 a13027a <=( a13026a  and  a13021a );
 a13030a <=( A267  and  A266 );
 a13034a <=( A302  and  (not A300) );
 a13035a <=( A268  and  a13034a );
 a13036a <=( a13035a  and  a13030a );
 a13039a <=( A166  and  A167 );
 a13043a <=( (not A265)  and  (not A200) );
 a13044a <=( (not A199)  and  a13043a );
 a13045a <=( a13044a  and  a13039a );
 a13048a <=( A267  and  A266 );
 a13052a <=( A299  and  A298 );
 a13053a <=( A268  and  a13052a );
 a13054a <=( a13053a  and  a13048a );
 a13057a <=( A166  and  A167 );
 a13061a <=( (not A265)  and  (not A200) );
 a13062a <=( (not A199)  and  a13061a );
 a13063a <=( a13062a  and  a13057a );
 a13066a <=( A267  and  A266 );
 a13070a <=( (not A299)  and  (not A298) );
 a13071a <=( A268  and  a13070a );
 a13072a <=( a13071a  and  a13066a );
 a13075a <=( A166  and  A167 );
 a13079a <=( (not A265)  and  (not A200) );
 a13080a <=( (not A199)  and  a13079a );
 a13081a <=( a13080a  and  a13075a );
 a13084a <=( A267  and  A266 );
 a13088a <=( A301  and  (not A300) );
 a13089a <=( A269  and  a13088a );
 a13090a <=( a13089a  and  a13084a );
 a13093a <=( A166  and  A167 );
 a13097a <=( (not A265)  and  (not A200) );
 a13098a <=( (not A199)  and  a13097a );
 a13099a <=( a13098a  and  a13093a );
 a13102a <=( A267  and  A266 );
 a13106a <=( A302  and  (not A300) );
 a13107a <=( A269  and  a13106a );
 a13108a <=( a13107a  and  a13102a );
 a13111a <=( A166  and  A167 );
 a13115a <=( (not A265)  and  (not A200) );
 a13116a <=( (not A199)  and  a13115a );
 a13117a <=( a13116a  and  a13111a );
 a13120a <=( A267  and  A266 );
 a13124a <=( A299  and  A298 );
 a13125a <=( A269  and  a13124a );
 a13126a <=( a13125a  and  a13120a );
 a13129a <=( A166  and  A167 );
 a13133a <=( (not A265)  and  (not A200) );
 a13134a <=( (not A199)  and  a13133a );
 a13135a <=( a13134a  and  a13129a );
 a13138a <=( A267  and  A266 );
 a13142a <=( (not A299)  and  (not A298) );
 a13143a <=( A269  and  a13142a );
 a13144a <=( a13143a  and  a13138a );
 a13147a <=( A166  and  A167 );
 a13151a <=( A265  and  (not A200) );
 a13152a <=( (not A199)  and  a13151a );
 a13153a <=( a13152a  and  a13147a );
 a13156a <=( A267  and  (not A266) );
 a13160a <=( A301  and  (not A300) );
 a13161a <=( A268  and  a13160a );
 a13162a <=( a13161a  and  a13156a );
 a13165a <=( A166  and  A167 );
 a13169a <=( A265  and  (not A200) );
 a13170a <=( (not A199)  and  a13169a );
 a13171a <=( a13170a  and  a13165a );
 a13174a <=( A267  and  (not A266) );
 a13178a <=( A302  and  (not A300) );
 a13179a <=( A268  and  a13178a );
 a13180a <=( a13179a  and  a13174a );
 a13183a <=( A166  and  A167 );
 a13187a <=( A265  and  (not A200) );
 a13188a <=( (not A199)  and  a13187a );
 a13189a <=( a13188a  and  a13183a );
 a13192a <=( A267  and  (not A266) );
 a13196a <=( A299  and  A298 );
 a13197a <=( A268  and  a13196a );
 a13198a <=( a13197a  and  a13192a );
 a13201a <=( A166  and  A167 );
 a13205a <=( A265  and  (not A200) );
 a13206a <=( (not A199)  and  a13205a );
 a13207a <=( a13206a  and  a13201a );
 a13210a <=( A267  and  (not A266) );
 a13214a <=( (not A299)  and  (not A298) );
 a13215a <=( A268  and  a13214a );
 a13216a <=( a13215a  and  a13210a );
 a13219a <=( A166  and  A167 );
 a13223a <=( A265  and  (not A200) );
 a13224a <=( (not A199)  and  a13223a );
 a13225a <=( a13224a  and  a13219a );
 a13228a <=( A267  and  (not A266) );
 a13232a <=( A301  and  (not A300) );
 a13233a <=( A269  and  a13232a );
 a13234a <=( a13233a  and  a13228a );
 a13237a <=( A166  and  A167 );
 a13241a <=( A265  and  (not A200) );
 a13242a <=( (not A199)  and  a13241a );
 a13243a <=( a13242a  and  a13237a );
 a13246a <=( A267  and  (not A266) );
 a13250a <=( A302  and  (not A300) );
 a13251a <=( A269  and  a13250a );
 a13252a <=( a13251a  and  a13246a );
 a13255a <=( A166  and  A167 );
 a13259a <=( A265  and  (not A200) );
 a13260a <=( (not A199)  and  a13259a );
 a13261a <=( a13260a  and  a13255a );
 a13264a <=( A267  and  (not A266) );
 a13268a <=( A299  and  A298 );
 a13269a <=( A269  and  a13268a );
 a13270a <=( a13269a  and  a13264a );
 a13273a <=( A166  and  A167 );
 a13277a <=( A265  and  (not A200) );
 a13278a <=( (not A199)  and  a13277a );
 a13279a <=( a13278a  and  a13273a );
 a13282a <=( A267  and  (not A266) );
 a13286a <=( (not A299)  and  (not A298) );
 a13287a <=( A269  and  a13286a );
 a13288a <=( a13287a  and  a13282a );
 a13291a <=( (not A166)  and  (not A167) );
 a13295a <=( (not A265)  and  A202 );
 a13296a <=( (not A201)  and  a13295a );
 a13297a <=( a13296a  and  a13291a );
 a13300a <=( A267  and  A266 );
 a13304a <=( A301  and  (not A300) );
 a13305a <=( A268  and  a13304a );
 a13306a <=( a13305a  and  a13300a );
 a13309a <=( (not A166)  and  (not A167) );
 a13313a <=( (not A265)  and  A202 );
 a13314a <=( (not A201)  and  a13313a );
 a13315a <=( a13314a  and  a13309a );
 a13318a <=( A267  and  A266 );
 a13322a <=( A302  and  (not A300) );
 a13323a <=( A268  and  a13322a );
 a13324a <=( a13323a  and  a13318a );
 a13327a <=( (not A166)  and  (not A167) );
 a13331a <=( (not A265)  and  A202 );
 a13332a <=( (not A201)  and  a13331a );
 a13333a <=( a13332a  and  a13327a );
 a13336a <=( A267  and  A266 );
 a13340a <=( A299  and  A298 );
 a13341a <=( A268  and  a13340a );
 a13342a <=( a13341a  and  a13336a );
 a13345a <=( (not A166)  and  (not A167) );
 a13349a <=( (not A265)  and  A202 );
 a13350a <=( (not A201)  and  a13349a );
 a13351a <=( a13350a  and  a13345a );
 a13354a <=( A267  and  A266 );
 a13358a <=( (not A299)  and  (not A298) );
 a13359a <=( A268  and  a13358a );
 a13360a <=( a13359a  and  a13354a );
 a13363a <=( (not A166)  and  (not A167) );
 a13367a <=( (not A265)  and  A202 );
 a13368a <=( (not A201)  and  a13367a );
 a13369a <=( a13368a  and  a13363a );
 a13372a <=( A267  and  A266 );
 a13376a <=( A301  and  (not A300) );
 a13377a <=( A269  and  a13376a );
 a13378a <=( a13377a  and  a13372a );
 a13381a <=( (not A166)  and  (not A167) );
 a13385a <=( (not A265)  and  A202 );
 a13386a <=( (not A201)  and  a13385a );
 a13387a <=( a13386a  and  a13381a );
 a13390a <=( A267  and  A266 );
 a13394a <=( A302  and  (not A300) );
 a13395a <=( A269  and  a13394a );
 a13396a <=( a13395a  and  a13390a );
 a13399a <=( (not A166)  and  (not A167) );
 a13403a <=( (not A265)  and  A202 );
 a13404a <=( (not A201)  and  a13403a );
 a13405a <=( a13404a  and  a13399a );
 a13408a <=( A267  and  A266 );
 a13412a <=( A299  and  A298 );
 a13413a <=( A269  and  a13412a );
 a13414a <=( a13413a  and  a13408a );
 a13417a <=( (not A166)  and  (not A167) );
 a13421a <=( (not A265)  and  A202 );
 a13422a <=( (not A201)  and  a13421a );
 a13423a <=( a13422a  and  a13417a );
 a13426a <=( A267  and  A266 );
 a13430a <=( (not A299)  and  (not A298) );
 a13431a <=( A269  and  a13430a );
 a13432a <=( a13431a  and  a13426a );
 a13435a <=( (not A166)  and  (not A167) );
 a13439a <=( A265  and  A202 );
 a13440a <=( (not A201)  and  a13439a );
 a13441a <=( a13440a  and  a13435a );
 a13444a <=( A267  and  (not A266) );
 a13448a <=( A301  and  (not A300) );
 a13449a <=( A268  and  a13448a );
 a13450a <=( a13449a  and  a13444a );
 a13453a <=( (not A166)  and  (not A167) );
 a13457a <=( A265  and  A202 );
 a13458a <=( (not A201)  and  a13457a );
 a13459a <=( a13458a  and  a13453a );
 a13462a <=( A267  and  (not A266) );
 a13466a <=( A302  and  (not A300) );
 a13467a <=( A268  and  a13466a );
 a13468a <=( a13467a  and  a13462a );
 a13471a <=( (not A166)  and  (not A167) );
 a13475a <=( A265  and  A202 );
 a13476a <=( (not A201)  and  a13475a );
 a13477a <=( a13476a  and  a13471a );
 a13480a <=( A267  and  (not A266) );
 a13484a <=( A299  and  A298 );
 a13485a <=( A268  and  a13484a );
 a13486a <=( a13485a  and  a13480a );
 a13489a <=( (not A166)  and  (not A167) );
 a13493a <=( A265  and  A202 );
 a13494a <=( (not A201)  and  a13493a );
 a13495a <=( a13494a  and  a13489a );
 a13498a <=( A267  and  (not A266) );
 a13502a <=( (not A299)  and  (not A298) );
 a13503a <=( A268  and  a13502a );
 a13504a <=( a13503a  and  a13498a );
 a13507a <=( (not A166)  and  (not A167) );
 a13511a <=( A265  and  A202 );
 a13512a <=( (not A201)  and  a13511a );
 a13513a <=( a13512a  and  a13507a );
 a13516a <=( A267  and  (not A266) );
 a13520a <=( A301  and  (not A300) );
 a13521a <=( A269  and  a13520a );
 a13522a <=( a13521a  and  a13516a );
 a13525a <=( (not A166)  and  (not A167) );
 a13529a <=( A265  and  A202 );
 a13530a <=( (not A201)  and  a13529a );
 a13531a <=( a13530a  and  a13525a );
 a13534a <=( A267  and  (not A266) );
 a13538a <=( A302  and  (not A300) );
 a13539a <=( A269  and  a13538a );
 a13540a <=( a13539a  and  a13534a );
 a13543a <=( (not A166)  and  (not A167) );
 a13547a <=( A265  and  A202 );
 a13548a <=( (not A201)  and  a13547a );
 a13549a <=( a13548a  and  a13543a );
 a13552a <=( A267  and  (not A266) );
 a13556a <=( A299  and  A298 );
 a13557a <=( A269  and  a13556a );
 a13558a <=( a13557a  and  a13552a );
 a13561a <=( (not A166)  and  (not A167) );
 a13565a <=( A265  and  A202 );
 a13566a <=( (not A201)  and  a13565a );
 a13567a <=( a13566a  and  a13561a );
 a13570a <=( A267  and  (not A266) );
 a13574a <=( (not A299)  and  (not A298) );
 a13575a <=( A269  and  a13574a );
 a13576a <=( a13575a  and  a13570a );
 a13579a <=( (not A166)  and  (not A167) );
 a13583a <=( (not A265)  and  A203 );
 a13584a <=( (not A201)  and  a13583a );
 a13585a <=( a13584a  and  a13579a );
 a13588a <=( A267  and  A266 );
 a13592a <=( A301  and  (not A300) );
 a13593a <=( A268  and  a13592a );
 a13594a <=( a13593a  and  a13588a );
 a13597a <=( (not A166)  and  (not A167) );
 a13601a <=( (not A265)  and  A203 );
 a13602a <=( (not A201)  and  a13601a );
 a13603a <=( a13602a  and  a13597a );
 a13606a <=( A267  and  A266 );
 a13610a <=( A302  and  (not A300) );
 a13611a <=( A268  and  a13610a );
 a13612a <=( a13611a  and  a13606a );
 a13615a <=( (not A166)  and  (not A167) );
 a13619a <=( (not A265)  and  A203 );
 a13620a <=( (not A201)  and  a13619a );
 a13621a <=( a13620a  and  a13615a );
 a13624a <=( A267  and  A266 );
 a13628a <=( A299  and  A298 );
 a13629a <=( A268  and  a13628a );
 a13630a <=( a13629a  and  a13624a );
 a13633a <=( (not A166)  and  (not A167) );
 a13637a <=( (not A265)  and  A203 );
 a13638a <=( (not A201)  and  a13637a );
 a13639a <=( a13638a  and  a13633a );
 a13642a <=( A267  and  A266 );
 a13646a <=( (not A299)  and  (not A298) );
 a13647a <=( A268  and  a13646a );
 a13648a <=( a13647a  and  a13642a );
 a13651a <=( (not A166)  and  (not A167) );
 a13655a <=( (not A265)  and  A203 );
 a13656a <=( (not A201)  and  a13655a );
 a13657a <=( a13656a  and  a13651a );
 a13660a <=( A267  and  A266 );
 a13664a <=( A301  and  (not A300) );
 a13665a <=( A269  and  a13664a );
 a13666a <=( a13665a  and  a13660a );
 a13669a <=( (not A166)  and  (not A167) );
 a13673a <=( (not A265)  and  A203 );
 a13674a <=( (not A201)  and  a13673a );
 a13675a <=( a13674a  and  a13669a );
 a13678a <=( A267  and  A266 );
 a13682a <=( A302  and  (not A300) );
 a13683a <=( A269  and  a13682a );
 a13684a <=( a13683a  and  a13678a );
 a13687a <=( (not A166)  and  (not A167) );
 a13691a <=( (not A265)  and  A203 );
 a13692a <=( (not A201)  and  a13691a );
 a13693a <=( a13692a  and  a13687a );
 a13696a <=( A267  and  A266 );
 a13700a <=( A299  and  A298 );
 a13701a <=( A269  and  a13700a );
 a13702a <=( a13701a  and  a13696a );
 a13705a <=( (not A166)  and  (not A167) );
 a13709a <=( (not A265)  and  A203 );
 a13710a <=( (not A201)  and  a13709a );
 a13711a <=( a13710a  and  a13705a );
 a13714a <=( A267  and  A266 );
 a13718a <=( (not A299)  and  (not A298) );
 a13719a <=( A269  and  a13718a );
 a13720a <=( a13719a  and  a13714a );
 a13723a <=( (not A166)  and  (not A167) );
 a13727a <=( A265  and  A203 );
 a13728a <=( (not A201)  and  a13727a );
 a13729a <=( a13728a  and  a13723a );
 a13732a <=( A267  and  (not A266) );
 a13736a <=( A301  and  (not A300) );
 a13737a <=( A268  and  a13736a );
 a13738a <=( a13737a  and  a13732a );
 a13741a <=( (not A166)  and  (not A167) );
 a13745a <=( A265  and  A203 );
 a13746a <=( (not A201)  and  a13745a );
 a13747a <=( a13746a  and  a13741a );
 a13750a <=( A267  and  (not A266) );
 a13754a <=( A302  and  (not A300) );
 a13755a <=( A268  and  a13754a );
 a13756a <=( a13755a  and  a13750a );
 a13759a <=( (not A166)  and  (not A167) );
 a13763a <=( A265  and  A203 );
 a13764a <=( (not A201)  and  a13763a );
 a13765a <=( a13764a  and  a13759a );
 a13768a <=( A267  and  (not A266) );
 a13772a <=( A299  and  A298 );
 a13773a <=( A268  and  a13772a );
 a13774a <=( a13773a  and  a13768a );
 a13777a <=( (not A166)  and  (not A167) );
 a13781a <=( A265  and  A203 );
 a13782a <=( (not A201)  and  a13781a );
 a13783a <=( a13782a  and  a13777a );
 a13786a <=( A267  and  (not A266) );
 a13790a <=( (not A299)  and  (not A298) );
 a13791a <=( A268  and  a13790a );
 a13792a <=( a13791a  and  a13786a );
 a13795a <=( (not A166)  and  (not A167) );
 a13799a <=( A265  and  A203 );
 a13800a <=( (not A201)  and  a13799a );
 a13801a <=( a13800a  and  a13795a );
 a13804a <=( A267  and  (not A266) );
 a13808a <=( A301  and  (not A300) );
 a13809a <=( A269  and  a13808a );
 a13810a <=( a13809a  and  a13804a );
 a13813a <=( (not A166)  and  (not A167) );
 a13817a <=( A265  and  A203 );
 a13818a <=( (not A201)  and  a13817a );
 a13819a <=( a13818a  and  a13813a );
 a13822a <=( A267  and  (not A266) );
 a13826a <=( A302  and  (not A300) );
 a13827a <=( A269  and  a13826a );
 a13828a <=( a13827a  and  a13822a );
 a13831a <=( (not A166)  and  (not A167) );
 a13835a <=( A265  and  A203 );
 a13836a <=( (not A201)  and  a13835a );
 a13837a <=( a13836a  and  a13831a );
 a13840a <=( A267  and  (not A266) );
 a13844a <=( A299  and  A298 );
 a13845a <=( A269  and  a13844a );
 a13846a <=( a13845a  and  a13840a );
 a13849a <=( (not A166)  and  (not A167) );
 a13853a <=( A265  and  A203 );
 a13854a <=( (not A201)  and  a13853a );
 a13855a <=( a13854a  and  a13849a );
 a13858a <=( A267  and  (not A266) );
 a13862a <=( (not A299)  and  (not A298) );
 a13863a <=( A269  and  a13862a );
 a13864a <=( a13863a  and  a13858a );
 a13867a <=( (not A166)  and  (not A167) );
 a13871a <=( (not A265)  and  A200 );
 a13872a <=( A199  and  a13871a );
 a13873a <=( a13872a  and  a13867a );
 a13876a <=( A267  and  A266 );
 a13880a <=( A301  and  (not A300) );
 a13881a <=( A268  and  a13880a );
 a13882a <=( a13881a  and  a13876a );
 a13885a <=( (not A166)  and  (not A167) );
 a13889a <=( (not A265)  and  A200 );
 a13890a <=( A199  and  a13889a );
 a13891a <=( a13890a  and  a13885a );
 a13894a <=( A267  and  A266 );
 a13898a <=( A302  and  (not A300) );
 a13899a <=( A268  and  a13898a );
 a13900a <=( a13899a  and  a13894a );
 a13903a <=( (not A166)  and  (not A167) );
 a13907a <=( (not A265)  and  A200 );
 a13908a <=( A199  and  a13907a );
 a13909a <=( a13908a  and  a13903a );
 a13912a <=( A267  and  A266 );
 a13916a <=( A299  and  A298 );
 a13917a <=( A268  and  a13916a );
 a13918a <=( a13917a  and  a13912a );
 a13921a <=( (not A166)  and  (not A167) );
 a13925a <=( (not A265)  and  A200 );
 a13926a <=( A199  and  a13925a );
 a13927a <=( a13926a  and  a13921a );
 a13930a <=( A267  and  A266 );
 a13934a <=( (not A299)  and  (not A298) );
 a13935a <=( A268  and  a13934a );
 a13936a <=( a13935a  and  a13930a );
 a13939a <=( (not A166)  and  (not A167) );
 a13943a <=( (not A265)  and  A200 );
 a13944a <=( A199  and  a13943a );
 a13945a <=( a13944a  and  a13939a );
 a13948a <=( A267  and  A266 );
 a13952a <=( A301  and  (not A300) );
 a13953a <=( A269  and  a13952a );
 a13954a <=( a13953a  and  a13948a );
 a13957a <=( (not A166)  and  (not A167) );
 a13961a <=( (not A265)  and  A200 );
 a13962a <=( A199  and  a13961a );
 a13963a <=( a13962a  and  a13957a );
 a13966a <=( A267  and  A266 );
 a13970a <=( A302  and  (not A300) );
 a13971a <=( A269  and  a13970a );
 a13972a <=( a13971a  and  a13966a );
 a13975a <=( (not A166)  and  (not A167) );
 a13979a <=( (not A265)  and  A200 );
 a13980a <=( A199  and  a13979a );
 a13981a <=( a13980a  and  a13975a );
 a13984a <=( A267  and  A266 );
 a13988a <=( A299  and  A298 );
 a13989a <=( A269  and  a13988a );
 a13990a <=( a13989a  and  a13984a );
 a13993a <=( (not A166)  and  (not A167) );
 a13997a <=( (not A265)  and  A200 );
 a13998a <=( A199  and  a13997a );
 a13999a <=( a13998a  and  a13993a );
 a14002a <=( A267  and  A266 );
 a14006a <=( (not A299)  and  (not A298) );
 a14007a <=( A269  and  a14006a );
 a14008a <=( a14007a  and  a14002a );
 a14011a <=( (not A166)  and  (not A167) );
 a14015a <=( A265  and  A200 );
 a14016a <=( A199  and  a14015a );
 a14017a <=( a14016a  and  a14011a );
 a14020a <=( A267  and  (not A266) );
 a14024a <=( A301  and  (not A300) );
 a14025a <=( A268  and  a14024a );
 a14026a <=( a14025a  and  a14020a );
 a14029a <=( (not A166)  and  (not A167) );
 a14033a <=( A265  and  A200 );
 a14034a <=( A199  and  a14033a );
 a14035a <=( a14034a  and  a14029a );
 a14038a <=( A267  and  (not A266) );
 a14042a <=( A302  and  (not A300) );
 a14043a <=( A268  and  a14042a );
 a14044a <=( a14043a  and  a14038a );
 a14047a <=( (not A166)  and  (not A167) );
 a14051a <=( A265  and  A200 );
 a14052a <=( A199  and  a14051a );
 a14053a <=( a14052a  and  a14047a );
 a14056a <=( A267  and  (not A266) );
 a14060a <=( A299  and  A298 );
 a14061a <=( A268  and  a14060a );
 a14062a <=( a14061a  and  a14056a );
 a14065a <=( (not A166)  and  (not A167) );
 a14069a <=( A265  and  A200 );
 a14070a <=( A199  and  a14069a );
 a14071a <=( a14070a  and  a14065a );
 a14074a <=( A267  and  (not A266) );
 a14078a <=( (not A299)  and  (not A298) );
 a14079a <=( A268  and  a14078a );
 a14080a <=( a14079a  and  a14074a );
 a14083a <=( (not A166)  and  (not A167) );
 a14087a <=( A265  and  A200 );
 a14088a <=( A199  and  a14087a );
 a14089a <=( a14088a  and  a14083a );
 a14092a <=( A267  and  (not A266) );
 a14096a <=( A301  and  (not A300) );
 a14097a <=( A269  and  a14096a );
 a14098a <=( a14097a  and  a14092a );
 a14101a <=( (not A166)  and  (not A167) );
 a14105a <=( A265  and  A200 );
 a14106a <=( A199  and  a14105a );
 a14107a <=( a14106a  and  a14101a );
 a14110a <=( A267  and  (not A266) );
 a14114a <=( A302  and  (not A300) );
 a14115a <=( A269  and  a14114a );
 a14116a <=( a14115a  and  a14110a );
 a14119a <=( (not A166)  and  (not A167) );
 a14123a <=( A265  and  A200 );
 a14124a <=( A199  and  a14123a );
 a14125a <=( a14124a  and  a14119a );
 a14128a <=( A267  and  (not A266) );
 a14132a <=( A299  and  A298 );
 a14133a <=( A269  and  a14132a );
 a14134a <=( a14133a  and  a14128a );
 a14137a <=( (not A166)  and  (not A167) );
 a14141a <=( A265  and  A200 );
 a14142a <=( A199  and  a14141a );
 a14143a <=( a14142a  and  a14137a );
 a14146a <=( A267  and  (not A266) );
 a14150a <=( (not A299)  and  (not A298) );
 a14151a <=( A269  and  a14150a );
 a14152a <=( a14151a  and  a14146a );
 a14155a <=( (not A166)  and  (not A167) );
 a14159a <=( (not A265)  and  (not A200) );
 a14160a <=( (not A199)  and  a14159a );
 a14161a <=( a14160a  and  a14155a );
 a14164a <=( A267  and  A266 );
 a14168a <=( A301  and  (not A300) );
 a14169a <=( A268  and  a14168a );
 a14170a <=( a14169a  and  a14164a );
 a14173a <=( (not A166)  and  (not A167) );
 a14177a <=( (not A265)  and  (not A200) );
 a14178a <=( (not A199)  and  a14177a );
 a14179a <=( a14178a  and  a14173a );
 a14182a <=( A267  and  A266 );
 a14186a <=( A302  and  (not A300) );
 a14187a <=( A268  and  a14186a );
 a14188a <=( a14187a  and  a14182a );
 a14191a <=( (not A166)  and  (not A167) );
 a14195a <=( (not A265)  and  (not A200) );
 a14196a <=( (not A199)  and  a14195a );
 a14197a <=( a14196a  and  a14191a );
 a14200a <=( A267  and  A266 );
 a14204a <=( A299  and  A298 );
 a14205a <=( A268  and  a14204a );
 a14206a <=( a14205a  and  a14200a );
 a14209a <=( (not A166)  and  (not A167) );
 a14213a <=( (not A265)  and  (not A200) );
 a14214a <=( (not A199)  and  a14213a );
 a14215a <=( a14214a  and  a14209a );
 a14218a <=( A267  and  A266 );
 a14222a <=( (not A299)  and  (not A298) );
 a14223a <=( A268  and  a14222a );
 a14224a <=( a14223a  and  a14218a );
 a14227a <=( (not A166)  and  (not A167) );
 a14231a <=( (not A265)  and  (not A200) );
 a14232a <=( (not A199)  and  a14231a );
 a14233a <=( a14232a  and  a14227a );
 a14236a <=( A267  and  A266 );
 a14240a <=( A301  and  (not A300) );
 a14241a <=( A269  and  a14240a );
 a14242a <=( a14241a  and  a14236a );
 a14245a <=( (not A166)  and  (not A167) );
 a14249a <=( (not A265)  and  (not A200) );
 a14250a <=( (not A199)  and  a14249a );
 a14251a <=( a14250a  and  a14245a );
 a14254a <=( A267  and  A266 );
 a14258a <=( A302  and  (not A300) );
 a14259a <=( A269  and  a14258a );
 a14260a <=( a14259a  and  a14254a );
 a14263a <=( (not A166)  and  (not A167) );
 a14267a <=( (not A265)  and  (not A200) );
 a14268a <=( (not A199)  and  a14267a );
 a14269a <=( a14268a  and  a14263a );
 a14272a <=( A267  and  A266 );
 a14276a <=( A299  and  A298 );
 a14277a <=( A269  and  a14276a );
 a14278a <=( a14277a  and  a14272a );
 a14281a <=( (not A166)  and  (not A167) );
 a14285a <=( (not A265)  and  (not A200) );
 a14286a <=( (not A199)  and  a14285a );
 a14287a <=( a14286a  and  a14281a );
 a14290a <=( A267  and  A266 );
 a14294a <=( (not A299)  and  (not A298) );
 a14295a <=( A269  and  a14294a );
 a14296a <=( a14295a  and  a14290a );
 a14299a <=( (not A166)  and  (not A167) );
 a14303a <=( A265  and  (not A200) );
 a14304a <=( (not A199)  and  a14303a );
 a14305a <=( a14304a  and  a14299a );
 a14308a <=( A267  and  (not A266) );
 a14312a <=( A301  and  (not A300) );
 a14313a <=( A268  and  a14312a );
 a14314a <=( a14313a  and  a14308a );
 a14317a <=( (not A166)  and  (not A167) );
 a14321a <=( A265  and  (not A200) );
 a14322a <=( (not A199)  and  a14321a );
 a14323a <=( a14322a  and  a14317a );
 a14326a <=( A267  and  (not A266) );
 a14330a <=( A302  and  (not A300) );
 a14331a <=( A268  and  a14330a );
 a14332a <=( a14331a  and  a14326a );
 a14335a <=( (not A166)  and  (not A167) );
 a14339a <=( A265  and  (not A200) );
 a14340a <=( (not A199)  and  a14339a );
 a14341a <=( a14340a  and  a14335a );
 a14344a <=( A267  and  (not A266) );
 a14348a <=( A299  and  A298 );
 a14349a <=( A268  and  a14348a );
 a14350a <=( a14349a  and  a14344a );
 a14353a <=( (not A166)  and  (not A167) );
 a14357a <=( A265  and  (not A200) );
 a14358a <=( (not A199)  and  a14357a );
 a14359a <=( a14358a  and  a14353a );
 a14362a <=( A267  and  (not A266) );
 a14366a <=( (not A299)  and  (not A298) );
 a14367a <=( A268  and  a14366a );
 a14368a <=( a14367a  and  a14362a );
 a14371a <=( (not A166)  and  (not A167) );
 a14375a <=( A265  and  (not A200) );
 a14376a <=( (not A199)  and  a14375a );
 a14377a <=( a14376a  and  a14371a );
 a14380a <=( A267  and  (not A266) );
 a14384a <=( A301  and  (not A300) );
 a14385a <=( A269  and  a14384a );
 a14386a <=( a14385a  and  a14380a );
 a14389a <=( (not A166)  and  (not A167) );
 a14393a <=( A265  and  (not A200) );
 a14394a <=( (not A199)  and  a14393a );
 a14395a <=( a14394a  and  a14389a );
 a14398a <=( A267  and  (not A266) );
 a14402a <=( A302  and  (not A300) );
 a14403a <=( A269  and  a14402a );
 a14404a <=( a14403a  and  a14398a );
 a14407a <=( (not A166)  and  (not A167) );
 a14411a <=( A265  and  (not A200) );
 a14412a <=( (not A199)  and  a14411a );
 a14413a <=( a14412a  and  a14407a );
 a14416a <=( A267  and  (not A266) );
 a14420a <=( A299  and  A298 );
 a14421a <=( A269  and  a14420a );
 a14422a <=( a14421a  and  a14416a );
 a14425a <=( (not A166)  and  (not A167) );
 a14429a <=( A265  and  (not A200) );
 a14430a <=( (not A199)  and  a14429a );
 a14431a <=( a14430a  and  a14425a );
 a14434a <=( A267  and  (not A266) );
 a14438a <=( (not A299)  and  (not A298) );
 a14439a <=( A269  and  a14438a );
 a14440a <=( a14439a  and  a14434a );
 a14443a <=( (not A168)  and  (not A170) );
 a14447a <=( (not A265)  and  A202 );
 a14448a <=( (not A201)  and  a14447a );
 a14449a <=( a14448a  and  a14443a );
 a14452a <=( A267  and  A266 );
 a14456a <=( A301  and  (not A300) );
 a14457a <=( A268  and  a14456a );
 a14458a <=( a14457a  and  a14452a );
 a14461a <=( (not A168)  and  (not A170) );
 a14465a <=( (not A265)  and  A202 );
 a14466a <=( (not A201)  and  a14465a );
 a14467a <=( a14466a  and  a14461a );
 a14470a <=( A267  and  A266 );
 a14474a <=( A302  and  (not A300) );
 a14475a <=( A268  and  a14474a );
 a14476a <=( a14475a  and  a14470a );
 a14479a <=( (not A168)  and  (not A170) );
 a14483a <=( (not A265)  and  A202 );
 a14484a <=( (not A201)  and  a14483a );
 a14485a <=( a14484a  and  a14479a );
 a14488a <=( A267  and  A266 );
 a14492a <=( A299  and  A298 );
 a14493a <=( A268  and  a14492a );
 a14494a <=( a14493a  and  a14488a );
 a14497a <=( (not A168)  and  (not A170) );
 a14501a <=( (not A265)  and  A202 );
 a14502a <=( (not A201)  and  a14501a );
 a14503a <=( a14502a  and  a14497a );
 a14506a <=( A267  and  A266 );
 a14510a <=( (not A299)  and  (not A298) );
 a14511a <=( A268  and  a14510a );
 a14512a <=( a14511a  and  a14506a );
 a14515a <=( (not A168)  and  (not A170) );
 a14519a <=( (not A265)  and  A202 );
 a14520a <=( (not A201)  and  a14519a );
 a14521a <=( a14520a  and  a14515a );
 a14524a <=( A267  and  A266 );
 a14528a <=( A301  and  (not A300) );
 a14529a <=( A269  and  a14528a );
 a14530a <=( a14529a  and  a14524a );
 a14533a <=( (not A168)  and  (not A170) );
 a14537a <=( (not A265)  and  A202 );
 a14538a <=( (not A201)  and  a14537a );
 a14539a <=( a14538a  and  a14533a );
 a14542a <=( A267  and  A266 );
 a14546a <=( A302  and  (not A300) );
 a14547a <=( A269  and  a14546a );
 a14548a <=( a14547a  and  a14542a );
 a14551a <=( (not A168)  and  (not A170) );
 a14555a <=( (not A265)  and  A202 );
 a14556a <=( (not A201)  and  a14555a );
 a14557a <=( a14556a  and  a14551a );
 a14560a <=( A267  and  A266 );
 a14564a <=( A299  and  A298 );
 a14565a <=( A269  and  a14564a );
 a14566a <=( a14565a  and  a14560a );
 a14569a <=( (not A168)  and  (not A170) );
 a14573a <=( (not A265)  and  A202 );
 a14574a <=( (not A201)  and  a14573a );
 a14575a <=( a14574a  and  a14569a );
 a14578a <=( A267  and  A266 );
 a14582a <=( (not A299)  and  (not A298) );
 a14583a <=( A269  and  a14582a );
 a14584a <=( a14583a  and  a14578a );
 a14587a <=( (not A168)  and  (not A170) );
 a14591a <=( A265  and  A202 );
 a14592a <=( (not A201)  and  a14591a );
 a14593a <=( a14592a  and  a14587a );
 a14596a <=( A267  and  (not A266) );
 a14600a <=( A301  and  (not A300) );
 a14601a <=( A268  and  a14600a );
 a14602a <=( a14601a  and  a14596a );
 a14605a <=( (not A168)  and  (not A170) );
 a14609a <=( A265  and  A202 );
 a14610a <=( (not A201)  and  a14609a );
 a14611a <=( a14610a  and  a14605a );
 a14614a <=( A267  and  (not A266) );
 a14618a <=( A302  and  (not A300) );
 a14619a <=( A268  and  a14618a );
 a14620a <=( a14619a  and  a14614a );
 a14623a <=( (not A168)  and  (not A170) );
 a14627a <=( A265  and  A202 );
 a14628a <=( (not A201)  and  a14627a );
 a14629a <=( a14628a  and  a14623a );
 a14632a <=( A267  and  (not A266) );
 a14636a <=( A299  and  A298 );
 a14637a <=( A268  and  a14636a );
 a14638a <=( a14637a  and  a14632a );
 a14641a <=( (not A168)  and  (not A170) );
 a14645a <=( A265  and  A202 );
 a14646a <=( (not A201)  and  a14645a );
 a14647a <=( a14646a  and  a14641a );
 a14650a <=( A267  and  (not A266) );
 a14654a <=( (not A299)  and  (not A298) );
 a14655a <=( A268  and  a14654a );
 a14656a <=( a14655a  and  a14650a );
 a14659a <=( (not A168)  and  (not A170) );
 a14663a <=( A265  and  A202 );
 a14664a <=( (not A201)  and  a14663a );
 a14665a <=( a14664a  and  a14659a );
 a14668a <=( A267  and  (not A266) );
 a14672a <=( A301  and  (not A300) );
 a14673a <=( A269  and  a14672a );
 a14674a <=( a14673a  and  a14668a );
 a14677a <=( (not A168)  and  (not A170) );
 a14681a <=( A265  and  A202 );
 a14682a <=( (not A201)  and  a14681a );
 a14683a <=( a14682a  and  a14677a );
 a14686a <=( A267  and  (not A266) );
 a14690a <=( A302  and  (not A300) );
 a14691a <=( A269  and  a14690a );
 a14692a <=( a14691a  and  a14686a );
 a14695a <=( (not A168)  and  (not A170) );
 a14699a <=( A265  and  A202 );
 a14700a <=( (not A201)  and  a14699a );
 a14701a <=( a14700a  and  a14695a );
 a14704a <=( A267  and  (not A266) );
 a14708a <=( A299  and  A298 );
 a14709a <=( A269  and  a14708a );
 a14710a <=( a14709a  and  a14704a );
 a14713a <=( (not A168)  and  (not A170) );
 a14717a <=( A265  and  A202 );
 a14718a <=( (not A201)  and  a14717a );
 a14719a <=( a14718a  and  a14713a );
 a14722a <=( A267  and  (not A266) );
 a14726a <=( (not A299)  and  (not A298) );
 a14727a <=( A269  and  a14726a );
 a14728a <=( a14727a  and  a14722a );
 a14731a <=( (not A168)  and  (not A170) );
 a14735a <=( (not A265)  and  A203 );
 a14736a <=( (not A201)  and  a14735a );
 a14737a <=( a14736a  and  a14731a );
 a14740a <=( A267  and  A266 );
 a14744a <=( A301  and  (not A300) );
 a14745a <=( A268  and  a14744a );
 a14746a <=( a14745a  and  a14740a );
 a14749a <=( (not A168)  and  (not A170) );
 a14753a <=( (not A265)  and  A203 );
 a14754a <=( (not A201)  and  a14753a );
 a14755a <=( a14754a  and  a14749a );
 a14758a <=( A267  and  A266 );
 a14762a <=( A302  and  (not A300) );
 a14763a <=( A268  and  a14762a );
 a14764a <=( a14763a  and  a14758a );
 a14767a <=( (not A168)  and  (not A170) );
 a14771a <=( (not A265)  and  A203 );
 a14772a <=( (not A201)  and  a14771a );
 a14773a <=( a14772a  and  a14767a );
 a14776a <=( A267  and  A266 );
 a14780a <=( A299  and  A298 );
 a14781a <=( A268  and  a14780a );
 a14782a <=( a14781a  and  a14776a );
 a14785a <=( (not A168)  and  (not A170) );
 a14789a <=( (not A265)  and  A203 );
 a14790a <=( (not A201)  and  a14789a );
 a14791a <=( a14790a  and  a14785a );
 a14794a <=( A267  and  A266 );
 a14798a <=( (not A299)  and  (not A298) );
 a14799a <=( A268  and  a14798a );
 a14800a <=( a14799a  and  a14794a );
 a14803a <=( (not A168)  and  (not A170) );
 a14807a <=( (not A265)  and  A203 );
 a14808a <=( (not A201)  and  a14807a );
 a14809a <=( a14808a  and  a14803a );
 a14812a <=( A267  and  A266 );
 a14816a <=( A301  and  (not A300) );
 a14817a <=( A269  and  a14816a );
 a14818a <=( a14817a  and  a14812a );
 a14821a <=( (not A168)  and  (not A170) );
 a14825a <=( (not A265)  and  A203 );
 a14826a <=( (not A201)  and  a14825a );
 a14827a <=( a14826a  and  a14821a );
 a14830a <=( A267  and  A266 );
 a14834a <=( A302  and  (not A300) );
 a14835a <=( A269  and  a14834a );
 a14836a <=( a14835a  and  a14830a );
 a14839a <=( (not A168)  and  (not A170) );
 a14843a <=( (not A265)  and  A203 );
 a14844a <=( (not A201)  and  a14843a );
 a14845a <=( a14844a  and  a14839a );
 a14848a <=( A267  and  A266 );
 a14852a <=( A299  and  A298 );
 a14853a <=( A269  and  a14852a );
 a14854a <=( a14853a  and  a14848a );
 a14857a <=( (not A168)  and  (not A170) );
 a14861a <=( (not A265)  and  A203 );
 a14862a <=( (not A201)  and  a14861a );
 a14863a <=( a14862a  and  a14857a );
 a14866a <=( A267  and  A266 );
 a14870a <=( (not A299)  and  (not A298) );
 a14871a <=( A269  and  a14870a );
 a14872a <=( a14871a  and  a14866a );
 a14875a <=( (not A168)  and  (not A170) );
 a14879a <=( A265  and  A203 );
 a14880a <=( (not A201)  and  a14879a );
 a14881a <=( a14880a  and  a14875a );
 a14884a <=( A267  and  (not A266) );
 a14888a <=( A301  and  (not A300) );
 a14889a <=( A268  and  a14888a );
 a14890a <=( a14889a  and  a14884a );
 a14893a <=( (not A168)  and  (not A170) );
 a14897a <=( A265  and  A203 );
 a14898a <=( (not A201)  and  a14897a );
 a14899a <=( a14898a  and  a14893a );
 a14902a <=( A267  and  (not A266) );
 a14906a <=( A302  and  (not A300) );
 a14907a <=( A268  and  a14906a );
 a14908a <=( a14907a  and  a14902a );
 a14911a <=( (not A168)  and  (not A170) );
 a14915a <=( A265  and  A203 );
 a14916a <=( (not A201)  and  a14915a );
 a14917a <=( a14916a  and  a14911a );
 a14920a <=( A267  and  (not A266) );
 a14924a <=( A299  and  A298 );
 a14925a <=( A268  and  a14924a );
 a14926a <=( a14925a  and  a14920a );
 a14929a <=( (not A168)  and  (not A170) );
 a14933a <=( A265  and  A203 );
 a14934a <=( (not A201)  and  a14933a );
 a14935a <=( a14934a  and  a14929a );
 a14938a <=( A267  and  (not A266) );
 a14942a <=( (not A299)  and  (not A298) );
 a14943a <=( A268  and  a14942a );
 a14944a <=( a14943a  and  a14938a );
 a14947a <=( (not A168)  and  (not A170) );
 a14951a <=( A265  and  A203 );
 a14952a <=( (not A201)  and  a14951a );
 a14953a <=( a14952a  and  a14947a );
 a14956a <=( A267  and  (not A266) );
 a14960a <=( A301  and  (not A300) );
 a14961a <=( A269  and  a14960a );
 a14962a <=( a14961a  and  a14956a );
 a14965a <=( (not A168)  and  (not A170) );
 a14969a <=( A265  and  A203 );
 a14970a <=( (not A201)  and  a14969a );
 a14971a <=( a14970a  and  a14965a );
 a14974a <=( A267  and  (not A266) );
 a14978a <=( A302  and  (not A300) );
 a14979a <=( A269  and  a14978a );
 a14980a <=( a14979a  and  a14974a );
 a14983a <=( (not A168)  and  (not A170) );
 a14987a <=( A265  and  A203 );
 a14988a <=( (not A201)  and  a14987a );
 a14989a <=( a14988a  and  a14983a );
 a14992a <=( A267  and  (not A266) );
 a14996a <=( A299  and  A298 );
 a14997a <=( A269  and  a14996a );
 a14998a <=( a14997a  and  a14992a );
 a15001a <=( (not A168)  and  (not A170) );
 a15005a <=( A265  and  A203 );
 a15006a <=( (not A201)  and  a15005a );
 a15007a <=( a15006a  and  a15001a );
 a15010a <=( A267  and  (not A266) );
 a15014a <=( (not A299)  and  (not A298) );
 a15015a <=( A269  and  a15014a );
 a15016a <=( a15015a  and  a15010a );
 a15019a <=( (not A168)  and  (not A170) );
 a15023a <=( (not A265)  and  A200 );
 a15024a <=( A199  and  a15023a );
 a15025a <=( a15024a  and  a15019a );
 a15028a <=( A267  and  A266 );
 a15032a <=( A301  and  (not A300) );
 a15033a <=( A268  and  a15032a );
 a15034a <=( a15033a  and  a15028a );
 a15037a <=( (not A168)  and  (not A170) );
 a15041a <=( (not A265)  and  A200 );
 a15042a <=( A199  and  a15041a );
 a15043a <=( a15042a  and  a15037a );
 a15046a <=( A267  and  A266 );
 a15050a <=( A302  and  (not A300) );
 a15051a <=( A268  and  a15050a );
 a15052a <=( a15051a  and  a15046a );
 a15055a <=( (not A168)  and  (not A170) );
 a15059a <=( (not A265)  and  A200 );
 a15060a <=( A199  and  a15059a );
 a15061a <=( a15060a  and  a15055a );
 a15064a <=( A267  and  A266 );
 a15068a <=( A299  and  A298 );
 a15069a <=( A268  and  a15068a );
 a15070a <=( a15069a  and  a15064a );
 a15073a <=( (not A168)  and  (not A170) );
 a15077a <=( (not A265)  and  A200 );
 a15078a <=( A199  and  a15077a );
 a15079a <=( a15078a  and  a15073a );
 a15082a <=( A267  and  A266 );
 a15086a <=( (not A299)  and  (not A298) );
 a15087a <=( A268  and  a15086a );
 a15088a <=( a15087a  and  a15082a );
 a15091a <=( (not A168)  and  (not A170) );
 a15095a <=( (not A265)  and  A200 );
 a15096a <=( A199  and  a15095a );
 a15097a <=( a15096a  and  a15091a );
 a15100a <=( A267  and  A266 );
 a15104a <=( A301  and  (not A300) );
 a15105a <=( A269  and  a15104a );
 a15106a <=( a15105a  and  a15100a );
 a15109a <=( (not A168)  and  (not A170) );
 a15113a <=( (not A265)  and  A200 );
 a15114a <=( A199  and  a15113a );
 a15115a <=( a15114a  and  a15109a );
 a15118a <=( A267  and  A266 );
 a15122a <=( A302  and  (not A300) );
 a15123a <=( A269  and  a15122a );
 a15124a <=( a15123a  and  a15118a );
 a15127a <=( (not A168)  and  (not A170) );
 a15131a <=( (not A265)  and  A200 );
 a15132a <=( A199  and  a15131a );
 a15133a <=( a15132a  and  a15127a );
 a15136a <=( A267  and  A266 );
 a15140a <=( A299  and  A298 );
 a15141a <=( A269  and  a15140a );
 a15142a <=( a15141a  and  a15136a );
 a15145a <=( (not A168)  and  (not A170) );
 a15149a <=( (not A265)  and  A200 );
 a15150a <=( A199  and  a15149a );
 a15151a <=( a15150a  and  a15145a );
 a15154a <=( A267  and  A266 );
 a15158a <=( (not A299)  and  (not A298) );
 a15159a <=( A269  and  a15158a );
 a15160a <=( a15159a  and  a15154a );
 a15163a <=( (not A168)  and  (not A170) );
 a15167a <=( A265  and  A200 );
 a15168a <=( A199  and  a15167a );
 a15169a <=( a15168a  and  a15163a );
 a15172a <=( A267  and  (not A266) );
 a15176a <=( A301  and  (not A300) );
 a15177a <=( A268  and  a15176a );
 a15178a <=( a15177a  and  a15172a );
 a15181a <=( (not A168)  and  (not A170) );
 a15185a <=( A265  and  A200 );
 a15186a <=( A199  and  a15185a );
 a15187a <=( a15186a  and  a15181a );
 a15190a <=( A267  and  (not A266) );
 a15194a <=( A302  and  (not A300) );
 a15195a <=( A268  and  a15194a );
 a15196a <=( a15195a  and  a15190a );
 a15199a <=( (not A168)  and  (not A170) );
 a15203a <=( A265  and  A200 );
 a15204a <=( A199  and  a15203a );
 a15205a <=( a15204a  and  a15199a );
 a15208a <=( A267  and  (not A266) );
 a15212a <=( A299  and  A298 );
 a15213a <=( A268  and  a15212a );
 a15214a <=( a15213a  and  a15208a );
 a15217a <=( (not A168)  and  (not A170) );
 a15221a <=( A265  and  A200 );
 a15222a <=( A199  and  a15221a );
 a15223a <=( a15222a  and  a15217a );
 a15226a <=( A267  and  (not A266) );
 a15230a <=( (not A299)  and  (not A298) );
 a15231a <=( A268  and  a15230a );
 a15232a <=( a15231a  and  a15226a );
 a15235a <=( (not A168)  and  (not A170) );
 a15239a <=( A265  and  A200 );
 a15240a <=( A199  and  a15239a );
 a15241a <=( a15240a  and  a15235a );
 a15244a <=( A267  and  (not A266) );
 a15248a <=( A301  and  (not A300) );
 a15249a <=( A269  and  a15248a );
 a15250a <=( a15249a  and  a15244a );
 a15253a <=( (not A168)  and  (not A170) );
 a15257a <=( A265  and  A200 );
 a15258a <=( A199  and  a15257a );
 a15259a <=( a15258a  and  a15253a );
 a15262a <=( A267  and  (not A266) );
 a15266a <=( A302  and  (not A300) );
 a15267a <=( A269  and  a15266a );
 a15268a <=( a15267a  and  a15262a );
 a15271a <=( (not A168)  and  (not A170) );
 a15275a <=( A265  and  A200 );
 a15276a <=( A199  and  a15275a );
 a15277a <=( a15276a  and  a15271a );
 a15280a <=( A267  and  (not A266) );
 a15284a <=( A299  and  A298 );
 a15285a <=( A269  and  a15284a );
 a15286a <=( a15285a  and  a15280a );
 a15289a <=( (not A168)  and  (not A170) );
 a15293a <=( A265  and  A200 );
 a15294a <=( A199  and  a15293a );
 a15295a <=( a15294a  and  a15289a );
 a15298a <=( A267  and  (not A266) );
 a15302a <=( (not A299)  and  (not A298) );
 a15303a <=( A269  and  a15302a );
 a15304a <=( a15303a  and  a15298a );
 a15307a <=( (not A168)  and  (not A170) );
 a15311a <=( (not A265)  and  (not A200) );
 a15312a <=( (not A199)  and  a15311a );
 a15313a <=( a15312a  and  a15307a );
 a15316a <=( A267  and  A266 );
 a15320a <=( A301  and  (not A300) );
 a15321a <=( A268  and  a15320a );
 a15322a <=( a15321a  and  a15316a );
 a15325a <=( (not A168)  and  (not A170) );
 a15329a <=( (not A265)  and  (not A200) );
 a15330a <=( (not A199)  and  a15329a );
 a15331a <=( a15330a  and  a15325a );
 a15334a <=( A267  and  A266 );
 a15338a <=( A302  and  (not A300) );
 a15339a <=( A268  and  a15338a );
 a15340a <=( a15339a  and  a15334a );
 a15343a <=( (not A168)  and  (not A170) );
 a15347a <=( (not A265)  and  (not A200) );
 a15348a <=( (not A199)  and  a15347a );
 a15349a <=( a15348a  and  a15343a );
 a15352a <=( A267  and  A266 );
 a15356a <=( A299  and  A298 );
 a15357a <=( A268  and  a15356a );
 a15358a <=( a15357a  and  a15352a );
 a15361a <=( (not A168)  and  (not A170) );
 a15365a <=( (not A265)  and  (not A200) );
 a15366a <=( (not A199)  and  a15365a );
 a15367a <=( a15366a  and  a15361a );
 a15370a <=( A267  and  A266 );
 a15374a <=( (not A299)  and  (not A298) );
 a15375a <=( A268  and  a15374a );
 a15376a <=( a15375a  and  a15370a );
 a15379a <=( (not A168)  and  (not A170) );
 a15383a <=( (not A265)  and  (not A200) );
 a15384a <=( (not A199)  and  a15383a );
 a15385a <=( a15384a  and  a15379a );
 a15388a <=( A267  and  A266 );
 a15392a <=( A301  and  (not A300) );
 a15393a <=( A269  and  a15392a );
 a15394a <=( a15393a  and  a15388a );
 a15397a <=( (not A168)  and  (not A170) );
 a15401a <=( (not A265)  and  (not A200) );
 a15402a <=( (not A199)  and  a15401a );
 a15403a <=( a15402a  and  a15397a );
 a15406a <=( A267  and  A266 );
 a15410a <=( A302  and  (not A300) );
 a15411a <=( A269  and  a15410a );
 a15412a <=( a15411a  and  a15406a );
 a15415a <=( (not A168)  and  (not A170) );
 a15419a <=( (not A265)  and  (not A200) );
 a15420a <=( (not A199)  and  a15419a );
 a15421a <=( a15420a  and  a15415a );
 a15424a <=( A267  and  A266 );
 a15428a <=( A299  and  A298 );
 a15429a <=( A269  and  a15428a );
 a15430a <=( a15429a  and  a15424a );
 a15433a <=( (not A168)  and  (not A170) );
 a15437a <=( (not A265)  and  (not A200) );
 a15438a <=( (not A199)  and  a15437a );
 a15439a <=( a15438a  and  a15433a );
 a15442a <=( A267  and  A266 );
 a15446a <=( (not A299)  and  (not A298) );
 a15447a <=( A269  and  a15446a );
 a15448a <=( a15447a  and  a15442a );
 a15451a <=( (not A168)  and  (not A170) );
 a15455a <=( A265  and  (not A200) );
 a15456a <=( (not A199)  and  a15455a );
 a15457a <=( a15456a  and  a15451a );
 a15460a <=( A267  and  (not A266) );
 a15464a <=( A301  and  (not A300) );
 a15465a <=( A268  and  a15464a );
 a15466a <=( a15465a  and  a15460a );
 a15469a <=( (not A168)  and  (not A170) );
 a15473a <=( A265  and  (not A200) );
 a15474a <=( (not A199)  and  a15473a );
 a15475a <=( a15474a  and  a15469a );
 a15478a <=( A267  and  (not A266) );
 a15482a <=( A302  and  (not A300) );
 a15483a <=( A268  and  a15482a );
 a15484a <=( a15483a  and  a15478a );
 a15487a <=( (not A168)  and  (not A170) );
 a15491a <=( A265  and  (not A200) );
 a15492a <=( (not A199)  and  a15491a );
 a15493a <=( a15492a  and  a15487a );
 a15496a <=( A267  and  (not A266) );
 a15500a <=( A299  and  A298 );
 a15501a <=( A268  and  a15500a );
 a15502a <=( a15501a  and  a15496a );
 a15505a <=( (not A168)  and  (not A170) );
 a15509a <=( A265  and  (not A200) );
 a15510a <=( (not A199)  and  a15509a );
 a15511a <=( a15510a  and  a15505a );
 a15514a <=( A267  and  (not A266) );
 a15518a <=( (not A299)  and  (not A298) );
 a15519a <=( A268  and  a15518a );
 a15520a <=( a15519a  and  a15514a );
 a15523a <=( (not A168)  and  (not A170) );
 a15527a <=( A265  and  (not A200) );
 a15528a <=( (not A199)  and  a15527a );
 a15529a <=( a15528a  and  a15523a );
 a15532a <=( A267  and  (not A266) );
 a15536a <=( A301  and  (not A300) );
 a15537a <=( A269  and  a15536a );
 a15538a <=( a15537a  and  a15532a );
 a15541a <=( (not A168)  and  (not A170) );
 a15545a <=( A265  and  (not A200) );
 a15546a <=( (not A199)  and  a15545a );
 a15547a <=( a15546a  and  a15541a );
 a15550a <=( A267  and  (not A266) );
 a15554a <=( A302  and  (not A300) );
 a15555a <=( A269  and  a15554a );
 a15556a <=( a15555a  and  a15550a );
 a15559a <=( (not A168)  and  (not A170) );
 a15563a <=( A265  and  (not A200) );
 a15564a <=( (not A199)  and  a15563a );
 a15565a <=( a15564a  and  a15559a );
 a15568a <=( A267  and  (not A266) );
 a15572a <=( A299  and  A298 );
 a15573a <=( A269  and  a15572a );
 a15574a <=( a15573a  and  a15568a );
 a15577a <=( (not A168)  and  (not A170) );
 a15581a <=( A265  and  (not A200) );
 a15582a <=( (not A199)  and  a15581a );
 a15583a <=( a15582a  and  a15577a );
 a15586a <=( A267  and  (not A266) );
 a15590a <=( (not A299)  and  (not A298) );
 a15591a <=( A269  and  a15590a );
 a15592a <=( a15591a  and  a15586a );
 a15595a <=( (not A168)  and  A169 );
 a15599a <=( (not A265)  and  A202 );
 a15600a <=( (not A201)  and  a15599a );
 a15601a <=( a15600a  and  a15595a );
 a15604a <=( A267  and  A266 );
 a15608a <=( A301  and  (not A300) );
 a15609a <=( A268  and  a15608a );
 a15610a <=( a15609a  and  a15604a );
 a15613a <=( (not A168)  and  A169 );
 a15617a <=( (not A265)  and  A202 );
 a15618a <=( (not A201)  and  a15617a );
 a15619a <=( a15618a  and  a15613a );
 a15622a <=( A267  and  A266 );
 a15626a <=( A302  and  (not A300) );
 a15627a <=( A268  and  a15626a );
 a15628a <=( a15627a  and  a15622a );
 a15631a <=( (not A168)  and  A169 );
 a15635a <=( (not A265)  and  A202 );
 a15636a <=( (not A201)  and  a15635a );
 a15637a <=( a15636a  and  a15631a );
 a15640a <=( A267  and  A266 );
 a15644a <=( A299  and  A298 );
 a15645a <=( A268  and  a15644a );
 a15646a <=( a15645a  and  a15640a );
 a15649a <=( (not A168)  and  A169 );
 a15653a <=( (not A265)  and  A202 );
 a15654a <=( (not A201)  and  a15653a );
 a15655a <=( a15654a  and  a15649a );
 a15658a <=( A267  and  A266 );
 a15662a <=( (not A299)  and  (not A298) );
 a15663a <=( A268  and  a15662a );
 a15664a <=( a15663a  and  a15658a );
 a15667a <=( (not A168)  and  A169 );
 a15671a <=( (not A265)  and  A202 );
 a15672a <=( (not A201)  and  a15671a );
 a15673a <=( a15672a  and  a15667a );
 a15676a <=( A267  and  A266 );
 a15680a <=( A301  and  (not A300) );
 a15681a <=( A269  and  a15680a );
 a15682a <=( a15681a  and  a15676a );
 a15685a <=( (not A168)  and  A169 );
 a15689a <=( (not A265)  and  A202 );
 a15690a <=( (not A201)  and  a15689a );
 a15691a <=( a15690a  and  a15685a );
 a15694a <=( A267  and  A266 );
 a15698a <=( A302  and  (not A300) );
 a15699a <=( A269  and  a15698a );
 a15700a <=( a15699a  and  a15694a );
 a15703a <=( (not A168)  and  A169 );
 a15707a <=( (not A265)  and  A202 );
 a15708a <=( (not A201)  and  a15707a );
 a15709a <=( a15708a  and  a15703a );
 a15712a <=( A267  and  A266 );
 a15716a <=( A299  and  A298 );
 a15717a <=( A269  and  a15716a );
 a15718a <=( a15717a  and  a15712a );
 a15721a <=( (not A168)  and  A169 );
 a15725a <=( (not A265)  and  A202 );
 a15726a <=( (not A201)  and  a15725a );
 a15727a <=( a15726a  and  a15721a );
 a15730a <=( A267  and  A266 );
 a15734a <=( (not A299)  and  (not A298) );
 a15735a <=( A269  and  a15734a );
 a15736a <=( a15735a  and  a15730a );
 a15739a <=( (not A168)  and  A169 );
 a15743a <=( A265  and  A202 );
 a15744a <=( (not A201)  and  a15743a );
 a15745a <=( a15744a  and  a15739a );
 a15748a <=( A267  and  (not A266) );
 a15752a <=( A301  and  (not A300) );
 a15753a <=( A268  and  a15752a );
 a15754a <=( a15753a  and  a15748a );
 a15757a <=( (not A168)  and  A169 );
 a15761a <=( A265  and  A202 );
 a15762a <=( (not A201)  and  a15761a );
 a15763a <=( a15762a  and  a15757a );
 a15766a <=( A267  and  (not A266) );
 a15770a <=( A302  and  (not A300) );
 a15771a <=( A268  and  a15770a );
 a15772a <=( a15771a  and  a15766a );
 a15775a <=( (not A168)  and  A169 );
 a15779a <=( A265  and  A202 );
 a15780a <=( (not A201)  and  a15779a );
 a15781a <=( a15780a  and  a15775a );
 a15784a <=( A267  and  (not A266) );
 a15788a <=( A299  and  A298 );
 a15789a <=( A268  and  a15788a );
 a15790a <=( a15789a  and  a15784a );
 a15793a <=( (not A168)  and  A169 );
 a15797a <=( A265  and  A202 );
 a15798a <=( (not A201)  and  a15797a );
 a15799a <=( a15798a  and  a15793a );
 a15802a <=( A267  and  (not A266) );
 a15806a <=( (not A299)  and  (not A298) );
 a15807a <=( A268  and  a15806a );
 a15808a <=( a15807a  and  a15802a );
 a15811a <=( (not A168)  and  A169 );
 a15815a <=( A265  and  A202 );
 a15816a <=( (not A201)  and  a15815a );
 a15817a <=( a15816a  and  a15811a );
 a15820a <=( A267  and  (not A266) );
 a15824a <=( A301  and  (not A300) );
 a15825a <=( A269  and  a15824a );
 a15826a <=( a15825a  and  a15820a );
 a15829a <=( (not A168)  and  A169 );
 a15833a <=( A265  and  A202 );
 a15834a <=( (not A201)  and  a15833a );
 a15835a <=( a15834a  and  a15829a );
 a15838a <=( A267  and  (not A266) );
 a15842a <=( A302  and  (not A300) );
 a15843a <=( A269  and  a15842a );
 a15844a <=( a15843a  and  a15838a );
 a15847a <=( (not A168)  and  A169 );
 a15851a <=( A265  and  A202 );
 a15852a <=( (not A201)  and  a15851a );
 a15853a <=( a15852a  and  a15847a );
 a15856a <=( A267  and  (not A266) );
 a15860a <=( A299  and  A298 );
 a15861a <=( A269  and  a15860a );
 a15862a <=( a15861a  and  a15856a );
 a15865a <=( (not A168)  and  A169 );
 a15869a <=( A265  and  A202 );
 a15870a <=( (not A201)  and  a15869a );
 a15871a <=( a15870a  and  a15865a );
 a15874a <=( A267  and  (not A266) );
 a15878a <=( (not A299)  and  (not A298) );
 a15879a <=( A269  and  a15878a );
 a15880a <=( a15879a  and  a15874a );
 a15883a <=( (not A168)  and  A169 );
 a15887a <=( (not A265)  and  A203 );
 a15888a <=( (not A201)  and  a15887a );
 a15889a <=( a15888a  and  a15883a );
 a15892a <=( A267  and  A266 );
 a15896a <=( A301  and  (not A300) );
 a15897a <=( A268  and  a15896a );
 a15898a <=( a15897a  and  a15892a );
 a15901a <=( (not A168)  and  A169 );
 a15905a <=( (not A265)  and  A203 );
 a15906a <=( (not A201)  and  a15905a );
 a15907a <=( a15906a  and  a15901a );
 a15910a <=( A267  and  A266 );
 a15914a <=( A302  and  (not A300) );
 a15915a <=( A268  and  a15914a );
 a15916a <=( a15915a  and  a15910a );
 a15919a <=( (not A168)  and  A169 );
 a15923a <=( (not A265)  and  A203 );
 a15924a <=( (not A201)  and  a15923a );
 a15925a <=( a15924a  and  a15919a );
 a15928a <=( A267  and  A266 );
 a15932a <=( A299  and  A298 );
 a15933a <=( A268  and  a15932a );
 a15934a <=( a15933a  and  a15928a );
 a15937a <=( (not A168)  and  A169 );
 a15941a <=( (not A265)  and  A203 );
 a15942a <=( (not A201)  and  a15941a );
 a15943a <=( a15942a  and  a15937a );
 a15946a <=( A267  and  A266 );
 a15950a <=( (not A299)  and  (not A298) );
 a15951a <=( A268  and  a15950a );
 a15952a <=( a15951a  and  a15946a );
 a15955a <=( (not A168)  and  A169 );
 a15959a <=( (not A265)  and  A203 );
 a15960a <=( (not A201)  and  a15959a );
 a15961a <=( a15960a  and  a15955a );
 a15964a <=( A267  and  A266 );
 a15968a <=( A301  and  (not A300) );
 a15969a <=( A269  and  a15968a );
 a15970a <=( a15969a  and  a15964a );
 a15973a <=( (not A168)  and  A169 );
 a15977a <=( (not A265)  and  A203 );
 a15978a <=( (not A201)  and  a15977a );
 a15979a <=( a15978a  and  a15973a );
 a15982a <=( A267  and  A266 );
 a15986a <=( A302  and  (not A300) );
 a15987a <=( A269  and  a15986a );
 a15988a <=( a15987a  and  a15982a );
 a15991a <=( (not A168)  and  A169 );
 a15995a <=( (not A265)  and  A203 );
 a15996a <=( (not A201)  and  a15995a );
 a15997a <=( a15996a  and  a15991a );
 a16000a <=( A267  and  A266 );
 a16004a <=( A299  and  A298 );
 a16005a <=( A269  and  a16004a );
 a16006a <=( a16005a  and  a16000a );
 a16009a <=( (not A168)  and  A169 );
 a16013a <=( (not A265)  and  A203 );
 a16014a <=( (not A201)  and  a16013a );
 a16015a <=( a16014a  and  a16009a );
 a16018a <=( A267  and  A266 );
 a16022a <=( (not A299)  and  (not A298) );
 a16023a <=( A269  and  a16022a );
 a16024a <=( a16023a  and  a16018a );
 a16027a <=( (not A168)  and  A169 );
 a16031a <=( A265  and  A203 );
 a16032a <=( (not A201)  and  a16031a );
 a16033a <=( a16032a  and  a16027a );
 a16036a <=( A267  and  (not A266) );
 a16040a <=( A301  and  (not A300) );
 a16041a <=( A268  and  a16040a );
 a16042a <=( a16041a  and  a16036a );
 a16045a <=( (not A168)  and  A169 );
 a16049a <=( A265  and  A203 );
 a16050a <=( (not A201)  and  a16049a );
 a16051a <=( a16050a  and  a16045a );
 a16054a <=( A267  and  (not A266) );
 a16058a <=( A302  and  (not A300) );
 a16059a <=( A268  and  a16058a );
 a16060a <=( a16059a  and  a16054a );
 a16063a <=( (not A168)  and  A169 );
 a16067a <=( A265  and  A203 );
 a16068a <=( (not A201)  and  a16067a );
 a16069a <=( a16068a  and  a16063a );
 a16072a <=( A267  and  (not A266) );
 a16076a <=( A299  and  A298 );
 a16077a <=( A268  and  a16076a );
 a16078a <=( a16077a  and  a16072a );
 a16081a <=( (not A168)  and  A169 );
 a16085a <=( A265  and  A203 );
 a16086a <=( (not A201)  and  a16085a );
 a16087a <=( a16086a  and  a16081a );
 a16090a <=( A267  and  (not A266) );
 a16094a <=( (not A299)  and  (not A298) );
 a16095a <=( A268  and  a16094a );
 a16096a <=( a16095a  and  a16090a );
 a16099a <=( (not A168)  and  A169 );
 a16103a <=( A265  and  A203 );
 a16104a <=( (not A201)  and  a16103a );
 a16105a <=( a16104a  and  a16099a );
 a16108a <=( A267  and  (not A266) );
 a16112a <=( A301  and  (not A300) );
 a16113a <=( A269  and  a16112a );
 a16114a <=( a16113a  and  a16108a );
 a16117a <=( (not A168)  and  A169 );
 a16121a <=( A265  and  A203 );
 a16122a <=( (not A201)  and  a16121a );
 a16123a <=( a16122a  and  a16117a );
 a16126a <=( A267  and  (not A266) );
 a16130a <=( A302  and  (not A300) );
 a16131a <=( A269  and  a16130a );
 a16132a <=( a16131a  and  a16126a );
 a16135a <=( (not A168)  and  A169 );
 a16139a <=( A265  and  A203 );
 a16140a <=( (not A201)  and  a16139a );
 a16141a <=( a16140a  and  a16135a );
 a16144a <=( A267  and  (not A266) );
 a16148a <=( A299  and  A298 );
 a16149a <=( A269  and  a16148a );
 a16150a <=( a16149a  and  a16144a );
 a16153a <=( (not A168)  and  A169 );
 a16157a <=( A265  and  A203 );
 a16158a <=( (not A201)  and  a16157a );
 a16159a <=( a16158a  and  a16153a );
 a16162a <=( A267  and  (not A266) );
 a16166a <=( (not A299)  and  (not A298) );
 a16167a <=( A269  and  a16166a );
 a16168a <=( a16167a  and  a16162a );
 a16171a <=( (not A168)  and  A169 );
 a16175a <=( (not A265)  and  A200 );
 a16176a <=( A199  and  a16175a );
 a16177a <=( a16176a  and  a16171a );
 a16180a <=( A267  and  A266 );
 a16184a <=( A301  and  (not A300) );
 a16185a <=( A268  and  a16184a );
 a16186a <=( a16185a  and  a16180a );
 a16189a <=( (not A168)  and  A169 );
 a16193a <=( (not A265)  and  A200 );
 a16194a <=( A199  and  a16193a );
 a16195a <=( a16194a  and  a16189a );
 a16198a <=( A267  and  A266 );
 a16202a <=( A302  and  (not A300) );
 a16203a <=( A268  and  a16202a );
 a16204a <=( a16203a  and  a16198a );
 a16207a <=( (not A168)  and  A169 );
 a16211a <=( (not A265)  and  A200 );
 a16212a <=( A199  and  a16211a );
 a16213a <=( a16212a  and  a16207a );
 a16216a <=( A267  and  A266 );
 a16220a <=( A299  and  A298 );
 a16221a <=( A268  and  a16220a );
 a16222a <=( a16221a  and  a16216a );
 a16225a <=( (not A168)  and  A169 );
 a16229a <=( (not A265)  and  A200 );
 a16230a <=( A199  and  a16229a );
 a16231a <=( a16230a  and  a16225a );
 a16234a <=( A267  and  A266 );
 a16238a <=( (not A299)  and  (not A298) );
 a16239a <=( A268  and  a16238a );
 a16240a <=( a16239a  and  a16234a );
 a16243a <=( (not A168)  and  A169 );
 a16247a <=( (not A265)  and  A200 );
 a16248a <=( A199  and  a16247a );
 a16249a <=( a16248a  and  a16243a );
 a16252a <=( A267  and  A266 );
 a16256a <=( A301  and  (not A300) );
 a16257a <=( A269  and  a16256a );
 a16258a <=( a16257a  and  a16252a );
 a16261a <=( (not A168)  and  A169 );
 a16265a <=( (not A265)  and  A200 );
 a16266a <=( A199  and  a16265a );
 a16267a <=( a16266a  and  a16261a );
 a16270a <=( A267  and  A266 );
 a16274a <=( A302  and  (not A300) );
 a16275a <=( A269  and  a16274a );
 a16276a <=( a16275a  and  a16270a );
 a16279a <=( (not A168)  and  A169 );
 a16283a <=( (not A265)  and  A200 );
 a16284a <=( A199  and  a16283a );
 a16285a <=( a16284a  and  a16279a );
 a16288a <=( A267  and  A266 );
 a16292a <=( A299  and  A298 );
 a16293a <=( A269  and  a16292a );
 a16294a <=( a16293a  and  a16288a );
 a16297a <=( (not A168)  and  A169 );
 a16301a <=( (not A265)  and  A200 );
 a16302a <=( A199  and  a16301a );
 a16303a <=( a16302a  and  a16297a );
 a16306a <=( A267  and  A266 );
 a16310a <=( (not A299)  and  (not A298) );
 a16311a <=( A269  and  a16310a );
 a16312a <=( a16311a  and  a16306a );
 a16315a <=( (not A168)  and  A169 );
 a16319a <=( A265  and  A200 );
 a16320a <=( A199  and  a16319a );
 a16321a <=( a16320a  and  a16315a );
 a16324a <=( A267  and  (not A266) );
 a16328a <=( A301  and  (not A300) );
 a16329a <=( A268  and  a16328a );
 a16330a <=( a16329a  and  a16324a );
 a16333a <=( (not A168)  and  A169 );
 a16337a <=( A265  and  A200 );
 a16338a <=( A199  and  a16337a );
 a16339a <=( a16338a  and  a16333a );
 a16342a <=( A267  and  (not A266) );
 a16346a <=( A302  and  (not A300) );
 a16347a <=( A268  and  a16346a );
 a16348a <=( a16347a  and  a16342a );
 a16351a <=( (not A168)  and  A169 );
 a16355a <=( A265  and  A200 );
 a16356a <=( A199  and  a16355a );
 a16357a <=( a16356a  and  a16351a );
 a16360a <=( A267  and  (not A266) );
 a16364a <=( A299  and  A298 );
 a16365a <=( A268  and  a16364a );
 a16366a <=( a16365a  and  a16360a );
 a16369a <=( (not A168)  and  A169 );
 a16373a <=( A265  and  A200 );
 a16374a <=( A199  and  a16373a );
 a16375a <=( a16374a  and  a16369a );
 a16378a <=( A267  and  (not A266) );
 a16382a <=( (not A299)  and  (not A298) );
 a16383a <=( A268  and  a16382a );
 a16384a <=( a16383a  and  a16378a );
 a16387a <=( (not A168)  and  A169 );
 a16391a <=( A265  and  A200 );
 a16392a <=( A199  and  a16391a );
 a16393a <=( a16392a  and  a16387a );
 a16396a <=( A267  and  (not A266) );
 a16400a <=( A301  and  (not A300) );
 a16401a <=( A269  and  a16400a );
 a16402a <=( a16401a  and  a16396a );
 a16405a <=( (not A168)  and  A169 );
 a16409a <=( A265  and  A200 );
 a16410a <=( A199  and  a16409a );
 a16411a <=( a16410a  and  a16405a );
 a16414a <=( A267  and  (not A266) );
 a16418a <=( A302  and  (not A300) );
 a16419a <=( A269  and  a16418a );
 a16420a <=( a16419a  and  a16414a );
 a16423a <=( (not A168)  and  A169 );
 a16427a <=( A265  and  A200 );
 a16428a <=( A199  and  a16427a );
 a16429a <=( a16428a  and  a16423a );
 a16432a <=( A267  and  (not A266) );
 a16436a <=( A299  and  A298 );
 a16437a <=( A269  and  a16436a );
 a16438a <=( a16437a  and  a16432a );
 a16441a <=( (not A168)  and  A169 );
 a16445a <=( A265  and  A200 );
 a16446a <=( A199  and  a16445a );
 a16447a <=( a16446a  and  a16441a );
 a16450a <=( A267  and  (not A266) );
 a16454a <=( (not A299)  and  (not A298) );
 a16455a <=( A269  and  a16454a );
 a16456a <=( a16455a  and  a16450a );
 a16459a <=( (not A168)  and  A169 );
 a16463a <=( (not A265)  and  (not A200) );
 a16464a <=( (not A199)  and  a16463a );
 a16465a <=( a16464a  and  a16459a );
 a16468a <=( A267  and  A266 );
 a16472a <=( A301  and  (not A300) );
 a16473a <=( A268  and  a16472a );
 a16474a <=( a16473a  and  a16468a );
 a16477a <=( (not A168)  and  A169 );
 a16481a <=( (not A265)  and  (not A200) );
 a16482a <=( (not A199)  and  a16481a );
 a16483a <=( a16482a  and  a16477a );
 a16486a <=( A267  and  A266 );
 a16490a <=( A302  and  (not A300) );
 a16491a <=( A268  and  a16490a );
 a16492a <=( a16491a  and  a16486a );
 a16495a <=( (not A168)  and  A169 );
 a16499a <=( (not A265)  and  (not A200) );
 a16500a <=( (not A199)  and  a16499a );
 a16501a <=( a16500a  and  a16495a );
 a16504a <=( A267  and  A266 );
 a16508a <=( A299  and  A298 );
 a16509a <=( A268  and  a16508a );
 a16510a <=( a16509a  and  a16504a );
 a16513a <=( (not A168)  and  A169 );
 a16517a <=( (not A265)  and  (not A200) );
 a16518a <=( (not A199)  and  a16517a );
 a16519a <=( a16518a  and  a16513a );
 a16522a <=( A267  and  A266 );
 a16526a <=( (not A299)  and  (not A298) );
 a16527a <=( A268  and  a16526a );
 a16528a <=( a16527a  and  a16522a );
 a16531a <=( (not A168)  and  A169 );
 a16535a <=( (not A265)  and  (not A200) );
 a16536a <=( (not A199)  and  a16535a );
 a16537a <=( a16536a  and  a16531a );
 a16540a <=( A267  and  A266 );
 a16544a <=( A301  and  (not A300) );
 a16545a <=( A269  and  a16544a );
 a16546a <=( a16545a  and  a16540a );
 a16549a <=( (not A168)  and  A169 );
 a16553a <=( (not A265)  and  (not A200) );
 a16554a <=( (not A199)  and  a16553a );
 a16555a <=( a16554a  and  a16549a );
 a16558a <=( A267  and  A266 );
 a16562a <=( A302  and  (not A300) );
 a16563a <=( A269  and  a16562a );
 a16564a <=( a16563a  and  a16558a );
 a16567a <=( (not A168)  and  A169 );
 a16571a <=( (not A265)  and  (not A200) );
 a16572a <=( (not A199)  and  a16571a );
 a16573a <=( a16572a  and  a16567a );
 a16576a <=( A267  and  A266 );
 a16580a <=( A299  and  A298 );
 a16581a <=( A269  and  a16580a );
 a16582a <=( a16581a  and  a16576a );
 a16585a <=( (not A168)  and  A169 );
 a16589a <=( (not A265)  and  (not A200) );
 a16590a <=( (not A199)  and  a16589a );
 a16591a <=( a16590a  and  a16585a );
 a16594a <=( A267  and  A266 );
 a16598a <=( (not A299)  and  (not A298) );
 a16599a <=( A269  and  a16598a );
 a16600a <=( a16599a  and  a16594a );
 a16603a <=( (not A168)  and  A169 );
 a16607a <=( A265  and  (not A200) );
 a16608a <=( (not A199)  and  a16607a );
 a16609a <=( a16608a  and  a16603a );
 a16612a <=( A267  and  (not A266) );
 a16616a <=( A301  and  (not A300) );
 a16617a <=( A268  and  a16616a );
 a16618a <=( a16617a  and  a16612a );
 a16621a <=( (not A168)  and  A169 );
 a16625a <=( A265  and  (not A200) );
 a16626a <=( (not A199)  and  a16625a );
 a16627a <=( a16626a  and  a16621a );
 a16630a <=( A267  and  (not A266) );
 a16634a <=( A302  and  (not A300) );
 a16635a <=( A268  and  a16634a );
 a16636a <=( a16635a  and  a16630a );
 a16639a <=( (not A168)  and  A169 );
 a16643a <=( A265  and  (not A200) );
 a16644a <=( (not A199)  and  a16643a );
 a16645a <=( a16644a  and  a16639a );
 a16648a <=( A267  and  (not A266) );
 a16652a <=( A299  and  A298 );
 a16653a <=( A268  and  a16652a );
 a16654a <=( a16653a  and  a16648a );
 a16657a <=( (not A168)  and  A169 );
 a16661a <=( A265  and  (not A200) );
 a16662a <=( (not A199)  and  a16661a );
 a16663a <=( a16662a  and  a16657a );
 a16666a <=( A267  and  (not A266) );
 a16670a <=( (not A299)  and  (not A298) );
 a16671a <=( A268  and  a16670a );
 a16672a <=( a16671a  and  a16666a );
 a16675a <=( (not A168)  and  A169 );
 a16679a <=( A265  and  (not A200) );
 a16680a <=( (not A199)  and  a16679a );
 a16681a <=( a16680a  and  a16675a );
 a16684a <=( A267  and  (not A266) );
 a16688a <=( A301  and  (not A300) );
 a16689a <=( A269  and  a16688a );
 a16690a <=( a16689a  and  a16684a );
 a16693a <=( (not A168)  and  A169 );
 a16697a <=( A265  and  (not A200) );
 a16698a <=( (not A199)  and  a16697a );
 a16699a <=( a16698a  and  a16693a );
 a16702a <=( A267  and  (not A266) );
 a16706a <=( A302  and  (not A300) );
 a16707a <=( A269  and  a16706a );
 a16708a <=( a16707a  and  a16702a );
 a16711a <=( (not A168)  and  A169 );
 a16715a <=( A265  and  (not A200) );
 a16716a <=( (not A199)  and  a16715a );
 a16717a <=( a16716a  and  a16711a );
 a16720a <=( A267  and  (not A266) );
 a16724a <=( A299  and  A298 );
 a16725a <=( A269  and  a16724a );
 a16726a <=( a16725a  and  a16720a );
 a16729a <=( (not A168)  and  A169 );
 a16733a <=( A265  and  (not A200) );
 a16734a <=( (not A199)  and  a16733a );
 a16735a <=( a16734a  and  a16729a );
 a16738a <=( A267  and  (not A266) );
 a16742a <=( (not A299)  and  (not A298) );
 a16743a <=( A269  and  a16742a );
 a16744a <=( a16743a  and  a16738a );
 a16747a <=( (not A169)  and  A170 );
 a16751a <=( (not A166)  and  A167 );
 a16752a <=( (not A168)  and  a16751a );
 a16753a <=( a16752a  and  a16747a );
 a16756a <=( A233  and  (not A232) );
 a16760a <=( (not A236)  and  (not A235) );
 a16761a <=( (not A234)  and  a16760a );
 a16762a <=( a16761a  and  a16756a );
 a16765a <=( (not A169)  and  A170 );
 a16769a <=( (not A166)  and  A167 );
 a16770a <=( (not A168)  and  a16769a );
 a16771a <=( a16770a  and  a16765a );
 a16774a <=( (not A233)  and  A232 );
 a16778a <=( (not A236)  and  (not A235) );
 a16779a <=( (not A234)  and  a16778a );
 a16780a <=( a16779a  and  a16774a );
 a16783a <=( (not A169)  and  A170 );
 a16787a <=( A166  and  (not A167) );
 a16788a <=( (not A168)  and  a16787a );
 a16789a <=( a16788a  and  a16783a );
 a16792a <=( A233  and  (not A232) );
 a16796a <=( (not A236)  and  (not A235) );
 a16797a <=( (not A234)  and  a16796a );
 a16798a <=( a16797a  and  a16792a );
 a16801a <=( (not A169)  and  A170 );
 a16805a <=( A166  and  (not A167) );
 a16806a <=( (not A168)  and  a16805a );
 a16807a <=( a16806a  and  a16801a );
 a16810a <=( (not A233)  and  A232 );
 a16814a <=( (not A236)  and  (not A235) );
 a16815a <=( (not A234)  and  a16814a );
 a16816a <=( a16815a  and  a16810a );
 a16819a <=( A166  and  A167 );
 a16823a <=( (not A203)  and  (not A202) );
 a16824a <=( A201  and  a16823a );
 a16825a <=( a16824a  and  a16819a );
 a16829a <=( A267  and  A266 );
 a16830a <=( (not A265)  and  a16829a );
 a16834a <=( A301  and  (not A300) );
 a16835a <=( A268  and  a16834a );
 a16836a <=( a16835a  and  a16830a );
 a16839a <=( A166  and  A167 );
 a16843a <=( (not A203)  and  (not A202) );
 a16844a <=( A201  and  a16843a );
 a16845a <=( a16844a  and  a16839a );
 a16849a <=( A267  and  A266 );
 a16850a <=( (not A265)  and  a16849a );
 a16854a <=( A302  and  (not A300) );
 a16855a <=( A268  and  a16854a );
 a16856a <=( a16855a  and  a16850a );
 a16859a <=( A166  and  A167 );
 a16863a <=( (not A203)  and  (not A202) );
 a16864a <=( A201  and  a16863a );
 a16865a <=( a16864a  and  a16859a );
 a16869a <=( A267  and  A266 );
 a16870a <=( (not A265)  and  a16869a );
 a16874a <=( A299  and  A298 );
 a16875a <=( A268  and  a16874a );
 a16876a <=( a16875a  and  a16870a );
 a16879a <=( A166  and  A167 );
 a16883a <=( (not A203)  and  (not A202) );
 a16884a <=( A201  and  a16883a );
 a16885a <=( a16884a  and  a16879a );
 a16889a <=( A267  and  A266 );
 a16890a <=( (not A265)  and  a16889a );
 a16894a <=( (not A299)  and  (not A298) );
 a16895a <=( A268  and  a16894a );
 a16896a <=( a16895a  and  a16890a );
 a16899a <=( A166  and  A167 );
 a16903a <=( (not A203)  and  (not A202) );
 a16904a <=( A201  and  a16903a );
 a16905a <=( a16904a  and  a16899a );
 a16909a <=( A267  and  A266 );
 a16910a <=( (not A265)  and  a16909a );
 a16914a <=( A301  and  (not A300) );
 a16915a <=( A269  and  a16914a );
 a16916a <=( a16915a  and  a16910a );
 a16919a <=( A166  and  A167 );
 a16923a <=( (not A203)  and  (not A202) );
 a16924a <=( A201  and  a16923a );
 a16925a <=( a16924a  and  a16919a );
 a16929a <=( A267  and  A266 );
 a16930a <=( (not A265)  and  a16929a );
 a16934a <=( A302  and  (not A300) );
 a16935a <=( A269  and  a16934a );
 a16936a <=( a16935a  and  a16930a );
 a16939a <=( A166  and  A167 );
 a16943a <=( (not A203)  and  (not A202) );
 a16944a <=( A201  and  a16943a );
 a16945a <=( a16944a  and  a16939a );
 a16949a <=( A267  and  A266 );
 a16950a <=( (not A265)  and  a16949a );
 a16954a <=( A299  and  A298 );
 a16955a <=( A269  and  a16954a );
 a16956a <=( a16955a  and  a16950a );
 a16959a <=( A166  and  A167 );
 a16963a <=( (not A203)  and  (not A202) );
 a16964a <=( A201  and  a16963a );
 a16965a <=( a16964a  and  a16959a );
 a16969a <=( A267  and  A266 );
 a16970a <=( (not A265)  and  a16969a );
 a16974a <=( (not A299)  and  (not A298) );
 a16975a <=( A269  and  a16974a );
 a16976a <=( a16975a  and  a16970a );
 a16979a <=( A166  and  A167 );
 a16983a <=( (not A203)  and  (not A202) );
 a16984a <=( A201  and  a16983a );
 a16985a <=( a16984a  and  a16979a );
 a16989a <=( A267  and  (not A266) );
 a16990a <=( A265  and  a16989a );
 a16994a <=( A301  and  (not A300) );
 a16995a <=( A268  and  a16994a );
 a16996a <=( a16995a  and  a16990a );
 a16999a <=( A166  and  A167 );
 a17003a <=( (not A203)  and  (not A202) );
 a17004a <=( A201  and  a17003a );
 a17005a <=( a17004a  and  a16999a );
 a17009a <=( A267  and  (not A266) );
 a17010a <=( A265  and  a17009a );
 a17014a <=( A302  and  (not A300) );
 a17015a <=( A268  and  a17014a );
 a17016a <=( a17015a  and  a17010a );
 a17019a <=( A166  and  A167 );
 a17023a <=( (not A203)  and  (not A202) );
 a17024a <=( A201  and  a17023a );
 a17025a <=( a17024a  and  a17019a );
 a17029a <=( A267  and  (not A266) );
 a17030a <=( A265  and  a17029a );
 a17034a <=( A299  and  A298 );
 a17035a <=( A268  and  a17034a );
 a17036a <=( a17035a  and  a17030a );
 a17039a <=( A166  and  A167 );
 a17043a <=( (not A203)  and  (not A202) );
 a17044a <=( A201  and  a17043a );
 a17045a <=( a17044a  and  a17039a );
 a17049a <=( A267  and  (not A266) );
 a17050a <=( A265  and  a17049a );
 a17054a <=( (not A299)  and  (not A298) );
 a17055a <=( A268  and  a17054a );
 a17056a <=( a17055a  and  a17050a );
 a17059a <=( A166  and  A167 );
 a17063a <=( (not A203)  and  (not A202) );
 a17064a <=( A201  and  a17063a );
 a17065a <=( a17064a  and  a17059a );
 a17069a <=( A267  and  (not A266) );
 a17070a <=( A265  and  a17069a );
 a17074a <=( A301  and  (not A300) );
 a17075a <=( A269  and  a17074a );
 a17076a <=( a17075a  and  a17070a );
 a17079a <=( A166  and  A167 );
 a17083a <=( (not A203)  and  (not A202) );
 a17084a <=( A201  and  a17083a );
 a17085a <=( a17084a  and  a17079a );
 a17089a <=( A267  and  (not A266) );
 a17090a <=( A265  and  a17089a );
 a17094a <=( A302  and  (not A300) );
 a17095a <=( A269  and  a17094a );
 a17096a <=( a17095a  and  a17090a );
 a17099a <=( A166  and  A167 );
 a17103a <=( (not A203)  and  (not A202) );
 a17104a <=( A201  and  a17103a );
 a17105a <=( a17104a  and  a17099a );
 a17109a <=( A267  and  (not A266) );
 a17110a <=( A265  and  a17109a );
 a17114a <=( A299  and  A298 );
 a17115a <=( A269  and  a17114a );
 a17116a <=( a17115a  and  a17110a );
 a17119a <=( A166  and  A167 );
 a17123a <=( (not A203)  and  (not A202) );
 a17124a <=( A201  and  a17123a );
 a17125a <=( a17124a  and  a17119a );
 a17129a <=( A267  and  (not A266) );
 a17130a <=( A265  and  a17129a );
 a17134a <=( (not A299)  and  (not A298) );
 a17135a <=( A269  and  a17134a );
 a17136a <=( a17135a  and  a17130a );
 a17139a <=( A166  and  A167 );
 a17143a <=( (not A265)  and  A202 );
 a17144a <=( (not A201)  and  a17143a );
 a17145a <=( a17144a  and  a17139a );
 a17149a <=( A268  and  A267 );
 a17150a <=( A266  and  a17149a );
 a17154a <=( (not A302)  and  (not A301) );
 a17155a <=( A300  and  a17154a );
 a17156a <=( a17155a  and  a17150a );
 a17159a <=( A166  and  A167 );
 a17163a <=( (not A265)  and  A202 );
 a17164a <=( (not A201)  and  a17163a );
 a17165a <=( a17164a  and  a17159a );
 a17169a <=( A269  and  A267 );
 a17170a <=( A266  and  a17169a );
 a17174a <=( (not A302)  and  (not A301) );
 a17175a <=( A300  and  a17174a );
 a17176a <=( a17175a  and  a17170a );
 a17179a <=( A166  and  A167 );
 a17183a <=( (not A265)  and  A202 );
 a17184a <=( (not A201)  and  a17183a );
 a17185a <=( a17184a  and  a17179a );
 a17189a <=( (not A268)  and  (not A267) );
 a17190a <=( A266  and  a17189a );
 a17194a <=( A301  and  (not A300) );
 a17195a <=( (not A269)  and  a17194a );
 a17196a <=( a17195a  and  a17190a );
 a17199a <=( A166  and  A167 );
 a17203a <=( (not A265)  and  A202 );
 a17204a <=( (not A201)  and  a17203a );
 a17205a <=( a17204a  and  a17199a );
 a17209a <=( (not A268)  and  (not A267) );
 a17210a <=( A266  and  a17209a );
 a17214a <=( A302  and  (not A300) );
 a17215a <=( (not A269)  and  a17214a );
 a17216a <=( a17215a  and  a17210a );
 a17219a <=( A166  and  A167 );
 a17223a <=( (not A265)  and  A202 );
 a17224a <=( (not A201)  and  a17223a );
 a17225a <=( a17224a  and  a17219a );
 a17229a <=( (not A268)  and  (not A267) );
 a17230a <=( A266  and  a17229a );
 a17234a <=( A299  and  A298 );
 a17235a <=( (not A269)  and  a17234a );
 a17236a <=( a17235a  and  a17230a );
 a17239a <=( A166  and  A167 );
 a17243a <=( (not A265)  and  A202 );
 a17244a <=( (not A201)  and  a17243a );
 a17245a <=( a17244a  and  a17239a );
 a17249a <=( (not A268)  and  (not A267) );
 a17250a <=( A266  and  a17249a );
 a17254a <=( (not A299)  and  (not A298) );
 a17255a <=( (not A269)  and  a17254a );
 a17256a <=( a17255a  and  a17250a );
 a17259a <=( A166  and  A167 );
 a17263a <=( A265  and  A202 );
 a17264a <=( (not A201)  and  a17263a );
 a17265a <=( a17264a  and  a17259a );
 a17269a <=( A268  and  A267 );
 a17270a <=( (not A266)  and  a17269a );
 a17274a <=( (not A302)  and  (not A301) );
 a17275a <=( A300  and  a17274a );
 a17276a <=( a17275a  and  a17270a );
 a17279a <=( A166  and  A167 );
 a17283a <=( A265  and  A202 );
 a17284a <=( (not A201)  and  a17283a );
 a17285a <=( a17284a  and  a17279a );
 a17289a <=( A269  and  A267 );
 a17290a <=( (not A266)  and  a17289a );
 a17294a <=( (not A302)  and  (not A301) );
 a17295a <=( A300  and  a17294a );
 a17296a <=( a17295a  and  a17290a );
 a17299a <=( A166  and  A167 );
 a17303a <=( A265  and  A202 );
 a17304a <=( (not A201)  and  a17303a );
 a17305a <=( a17304a  and  a17299a );
 a17309a <=( (not A268)  and  (not A267) );
 a17310a <=( (not A266)  and  a17309a );
 a17314a <=( A301  and  (not A300) );
 a17315a <=( (not A269)  and  a17314a );
 a17316a <=( a17315a  and  a17310a );
 a17319a <=( A166  and  A167 );
 a17323a <=( A265  and  A202 );
 a17324a <=( (not A201)  and  a17323a );
 a17325a <=( a17324a  and  a17319a );
 a17329a <=( (not A268)  and  (not A267) );
 a17330a <=( (not A266)  and  a17329a );
 a17334a <=( A302  and  (not A300) );
 a17335a <=( (not A269)  and  a17334a );
 a17336a <=( a17335a  and  a17330a );
 a17339a <=( A166  and  A167 );
 a17343a <=( A265  and  A202 );
 a17344a <=( (not A201)  and  a17343a );
 a17345a <=( a17344a  and  a17339a );
 a17349a <=( (not A268)  and  (not A267) );
 a17350a <=( (not A266)  and  a17349a );
 a17354a <=( A299  and  A298 );
 a17355a <=( (not A269)  and  a17354a );
 a17356a <=( a17355a  and  a17350a );
 a17359a <=( A166  and  A167 );
 a17363a <=( A265  and  A202 );
 a17364a <=( (not A201)  and  a17363a );
 a17365a <=( a17364a  and  a17359a );
 a17369a <=( (not A268)  and  (not A267) );
 a17370a <=( (not A266)  and  a17369a );
 a17374a <=( (not A299)  and  (not A298) );
 a17375a <=( (not A269)  and  a17374a );
 a17376a <=( a17375a  and  a17370a );
 a17379a <=( A166  and  A167 );
 a17383a <=( (not A265)  and  A203 );
 a17384a <=( (not A201)  and  a17383a );
 a17385a <=( a17384a  and  a17379a );
 a17389a <=( A268  and  A267 );
 a17390a <=( A266  and  a17389a );
 a17394a <=( (not A302)  and  (not A301) );
 a17395a <=( A300  and  a17394a );
 a17396a <=( a17395a  and  a17390a );
 a17399a <=( A166  and  A167 );
 a17403a <=( (not A265)  and  A203 );
 a17404a <=( (not A201)  and  a17403a );
 a17405a <=( a17404a  and  a17399a );
 a17409a <=( A269  and  A267 );
 a17410a <=( A266  and  a17409a );
 a17414a <=( (not A302)  and  (not A301) );
 a17415a <=( A300  and  a17414a );
 a17416a <=( a17415a  and  a17410a );
 a17419a <=( A166  and  A167 );
 a17423a <=( (not A265)  and  A203 );
 a17424a <=( (not A201)  and  a17423a );
 a17425a <=( a17424a  and  a17419a );
 a17429a <=( (not A268)  and  (not A267) );
 a17430a <=( A266  and  a17429a );
 a17434a <=( A301  and  (not A300) );
 a17435a <=( (not A269)  and  a17434a );
 a17436a <=( a17435a  and  a17430a );
 a17439a <=( A166  and  A167 );
 a17443a <=( (not A265)  and  A203 );
 a17444a <=( (not A201)  and  a17443a );
 a17445a <=( a17444a  and  a17439a );
 a17449a <=( (not A268)  and  (not A267) );
 a17450a <=( A266  and  a17449a );
 a17454a <=( A302  and  (not A300) );
 a17455a <=( (not A269)  and  a17454a );
 a17456a <=( a17455a  and  a17450a );
 a17459a <=( A166  and  A167 );
 a17463a <=( (not A265)  and  A203 );
 a17464a <=( (not A201)  and  a17463a );
 a17465a <=( a17464a  and  a17459a );
 a17469a <=( (not A268)  and  (not A267) );
 a17470a <=( A266  and  a17469a );
 a17474a <=( A299  and  A298 );
 a17475a <=( (not A269)  and  a17474a );
 a17476a <=( a17475a  and  a17470a );
 a17479a <=( A166  and  A167 );
 a17483a <=( (not A265)  and  A203 );
 a17484a <=( (not A201)  and  a17483a );
 a17485a <=( a17484a  and  a17479a );
 a17489a <=( (not A268)  and  (not A267) );
 a17490a <=( A266  and  a17489a );
 a17494a <=( (not A299)  and  (not A298) );
 a17495a <=( (not A269)  and  a17494a );
 a17496a <=( a17495a  and  a17490a );
 a17499a <=( A166  and  A167 );
 a17503a <=( A265  and  A203 );
 a17504a <=( (not A201)  and  a17503a );
 a17505a <=( a17504a  and  a17499a );
 a17509a <=( A268  and  A267 );
 a17510a <=( (not A266)  and  a17509a );
 a17514a <=( (not A302)  and  (not A301) );
 a17515a <=( A300  and  a17514a );
 a17516a <=( a17515a  and  a17510a );
 a17519a <=( A166  and  A167 );
 a17523a <=( A265  and  A203 );
 a17524a <=( (not A201)  and  a17523a );
 a17525a <=( a17524a  and  a17519a );
 a17529a <=( A269  and  A267 );
 a17530a <=( (not A266)  and  a17529a );
 a17534a <=( (not A302)  and  (not A301) );
 a17535a <=( A300  and  a17534a );
 a17536a <=( a17535a  and  a17530a );
 a17539a <=( A166  and  A167 );
 a17543a <=( A265  and  A203 );
 a17544a <=( (not A201)  and  a17543a );
 a17545a <=( a17544a  and  a17539a );
 a17549a <=( (not A268)  and  (not A267) );
 a17550a <=( (not A266)  and  a17549a );
 a17554a <=( A301  and  (not A300) );
 a17555a <=( (not A269)  and  a17554a );
 a17556a <=( a17555a  and  a17550a );
 a17559a <=( A166  and  A167 );
 a17563a <=( A265  and  A203 );
 a17564a <=( (not A201)  and  a17563a );
 a17565a <=( a17564a  and  a17559a );
 a17569a <=( (not A268)  and  (not A267) );
 a17570a <=( (not A266)  and  a17569a );
 a17574a <=( A302  and  (not A300) );
 a17575a <=( (not A269)  and  a17574a );
 a17576a <=( a17575a  and  a17570a );
 a17579a <=( A166  and  A167 );
 a17583a <=( A265  and  A203 );
 a17584a <=( (not A201)  and  a17583a );
 a17585a <=( a17584a  and  a17579a );
 a17589a <=( (not A268)  and  (not A267) );
 a17590a <=( (not A266)  and  a17589a );
 a17594a <=( A299  and  A298 );
 a17595a <=( (not A269)  and  a17594a );
 a17596a <=( a17595a  and  a17590a );
 a17599a <=( A166  and  A167 );
 a17603a <=( A265  and  A203 );
 a17604a <=( (not A201)  and  a17603a );
 a17605a <=( a17604a  and  a17599a );
 a17609a <=( (not A268)  and  (not A267) );
 a17610a <=( (not A266)  and  a17609a );
 a17614a <=( (not A299)  and  (not A298) );
 a17615a <=( (not A269)  and  a17614a );
 a17616a <=( a17615a  and  a17610a );
 a17619a <=( A166  and  A167 );
 a17623a <=( (not A265)  and  A200 );
 a17624a <=( A199  and  a17623a );
 a17625a <=( a17624a  and  a17619a );
 a17629a <=( A268  and  A267 );
 a17630a <=( A266  and  a17629a );
 a17634a <=( (not A302)  and  (not A301) );
 a17635a <=( A300  and  a17634a );
 a17636a <=( a17635a  and  a17630a );
 a17639a <=( A166  and  A167 );
 a17643a <=( (not A265)  and  A200 );
 a17644a <=( A199  and  a17643a );
 a17645a <=( a17644a  and  a17639a );
 a17649a <=( A269  and  A267 );
 a17650a <=( A266  and  a17649a );
 a17654a <=( (not A302)  and  (not A301) );
 a17655a <=( A300  and  a17654a );
 a17656a <=( a17655a  and  a17650a );
 a17659a <=( A166  and  A167 );
 a17663a <=( (not A265)  and  A200 );
 a17664a <=( A199  and  a17663a );
 a17665a <=( a17664a  and  a17659a );
 a17669a <=( (not A268)  and  (not A267) );
 a17670a <=( A266  and  a17669a );
 a17674a <=( A301  and  (not A300) );
 a17675a <=( (not A269)  and  a17674a );
 a17676a <=( a17675a  and  a17670a );
 a17679a <=( A166  and  A167 );
 a17683a <=( (not A265)  and  A200 );
 a17684a <=( A199  and  a17683a );
 a17685a <=( a17684a  and  a17679a );
 a17689a <=( (not A268)  and  (not A267) );
 a17690a <=( A266  and  a17689a );
 a17694a <=( A302  and  (not A300) );
 a17695a <=( (not A269)  and  a17694a );
 a17696a <=( a17695a  and  a17690a );
 a17699a <=( A166  and  A167 );
 a17703a <=( (not A265)  and  A200 );
 a17704a <=( A199  and  a17703a );
 a17705a <=( a17704a  and  a17699a );
 a17709a <=( (not A268)  and  (not A267) );
 a17710a <=( A266  and  a17709a );
 a17714a <=( A299  and  A298 );
 a17715a <=( (not A269)  and  a17714a );
 a17716a <=( a17715a  and  a17710a );
 a17719a <=( A166  and  A167 );
 a17723a <=( (not A265)  and  A200 );
 a17724a <=( A199  and  a17723a );
 a17725a <=( a17724a  and  a17719a );
 a17729a <=( (not A268)  and  (not A267) );
 a17730a <=( A266  and  a17729a );
 a17734a <=( (not A299)  and  (not A298) );
 a17735a <=( (not A269)  and  a17734a );
 a17736a <=( a17735a  and  a17730a );
 a17739a <=( A166  and  A167 );
 a17743a <=( A265  and  A200 );
 a17744a <=( A199  and  a17743a );
 a17745a <=( a17744a  and  a17739a );
 a17749a <=( A268  and  A267 );
 a17750a <=( (not A266)  and  a17749a );
 a17754a <=( (not A302)  and  (not A301) );
 a17755a <=( A300  and  a17754a );
 a17756a <=( a17755a  and  a17750a );
 a17759a <=( A166  and  A167 );
 a17763a <=( A265  and  A200 );
 a17764a <=( A199  and  a17763a );
 a17765a <=( a17764a  and  a17759a );
 a17769a <=( A269  and  A267 );
 a17770a <=( (not A266)  and  a17769a );
 a17774a <=( (not A302)  and  (not A301) );
 a17775a <=( A300  and  a17774a );
 a17776a <=( a17775a  and  a17770a );
 a17779a <=( A166  and  A167 );
 a17783a <=( A265  and  A200 );
 a17784a <=( A199  and  a17783a );
 a17785a <=( a17784a  and  a17779a );
 a17789a <=( (not A268)  and  (not A267) );
 a17790a <=( (not A266)  and  a17789a );
 a17794a <=( A301  and  (not A300) );
 a17795a <=( (not A269)  and  a17794a );
 a17796a <=( a17795a  and  a17790a );
 a17799a <=( A166  and  A167 );
 a17803a <=( A265  and  A200 );
 a17804a <=( A199  and  a17803a );
 a17805a <=( a17804a  and  a17799a );
 a17809a <=( (not A268)  and  (not A267) );
 a17810a <=( (not A266)  and  a17809a );
 a17814a <=( A302  and  (not A300) );
 a17815a <=( (not A269)  and  a17814a );
 a17816a <=( a17815a  and  a17810a );
 a17819a <=( A166  and  A167 );
 a17823a <=( A265  and  A200 );
 a17824a <=( A199  and  a17823a );
 a17825a <=( a17824a  and  a17819a );
 a17829a <=( (not A268)  and  (not A267) );
 a17830a <=( (not A266)  and  a17829a );
 a17834a <=( A299  and  A298 );
 a17835a <=( (not A269)  and  a17834a );
 a17836a <=( a17835a  and  a17830a );
 a17839a <=( A166  and  A167 );
 a17843a <=( A265  and  A200 );
 a17844a <=( A199  and  a17843a );
 a17845a <=( a17844a  and  a17839a );
 a17849a <=( (not A268)  and  (not A267) );
 a17850a <=( (not A266)  and  a17849a );
 a17854a <=( (not A299)  and  (not A298) );
 a17855a <=( (not A269)  and  a17854a );
 a17856a <=( a17855a  and  a17850a );
 a17859a <=( A166  and  A167 );
 a17863a <=( (not A265)  and  (not A200) );
 a17864a <=( (not A199)  and  a17863a );
 a17865a <=( a17864a  and  a17859a );
 a17869a <=( A268  and  A267 );
 a17870a <=( A266  and  a17869a );
 a17874a <=( (not A302)  and  (not A301) );
 a17875a <=( A300  and  a17874a );
 a17876a <=( a17875a  and  a17870a );
 a17879a <=( A166  and  A167 );
 a17883a <=( (not A265)  and  (not A200) );
 a17884a <=( (not A199)  and  a17883a );
 a17885a <=( a17884a  and  a17879a );
 a17889a <=( A269  and  A267 );
 a17890a <=( A266  and  a17889a );
 a17894a <=( (not A302)  and  (not A301) );
 a17895a <=( A300  and  a17894a );
 a17896a <=( a17895a  and  a17890a );
 a17899a <=( A166  and  A167 );
 a17903a <=( (not A265)  and  (not A200) );
 a17904a <=( (not A199)  and  a17903a );
 a17905a <=( a17904a  and  a17899a );
 a17909a <=( (not A268)  and  (not A267) );
 a17910a <=( A266  and  a17909a );
 a17914a <=( A301  and  (not A300) );
 a17915a <=( (not A269)  and  a17914a );
 a17916a <=( a17915a  and  a17910a );
 a17919a <=( A166  and  A167 );
 a17923a <=( (not A265)  and  (not A200) );
 a17924a <=( (not A199)  and  a17923a );
 a17925a <=( a17924a  and  a17919a );
 a17929a <=( (not A268)  and  (not A267) );
 a17930a <=( A266  and  a17929a );
 a17934a <=( A302  and  (not A300) );
 a17935a <=( (not A269)  and  a17934a );
 a17936a <=( a17935a  and  a17930a );
 a17939a <=( A166  and  A167 );
 a17943a <=( (not A265)  and  (not A200) );
 a17944a <=( (not A199)  and  a17943a );
 a17945a <=( a17944a  and  a17939a );
 a17949a <=( (not A268)  and  (not A267) );
 a17950a <=( A266  and  a17949a );
 a17954a <=( A299  and  A298 );
 a17955a <=( (not A269)  and  a17954a );
 a17956a <=( a17955a  and  a17950a );
 a17959a <=( A166  and  A167 );
 a17963a <=( (not A265)  and  (not A200) );
 a17964a <=( (not A199)  and  a17963a );
 a17965a <=( a17964a  and  a17959a );
 a17969a <=( (not A268)  and  (not A267) );
 a17970a <=( A266  and  a17969a );
 a17974a <=( (not A299)  and  (not A298) );
 a17975a <=( (not A269)  and  a17974a );
 a17976a <=( a17975a  and  a17970a );
 a17979a <=( A166  and  A167 );
 a17983a <=( A265  and  (not A200) );
 a17984a <=( (not A199)  and  a17983a );
 a17985a <=( a17984a  and  a17979a );
 a17989a <=( A268  and  A267 );
 a17990a <=( (not A266)  and  a17989a );
 a17994a <=( (not A302)  and  (not A301) );
 a17995a <=( A300  and  a17994a );
 a17996a <=( a17995a  and  a17990a );
 a17999a <=( A166  and  A167 );
 a18003a <=( A265  and  (not A200) );
 a18004a <=( (not A199)  and  a18003a );
 a18005a <=( a18004a  and  a17999a );
 a18009a <=( A269  and  A267 );
 a18010a <=( (not A266)  and  a18009a );
 a18014a <=( (not A302)  and  (not A301) );
 a18015a <=( A300  and  a18014a );
 a18016a <=( a18015a  and  a18010a );
 a18019a <=( A166  and  A167 );
 a18023a <=( A265  and  (not A200) );
 a18024a <=( (not A199)  and  a18023a );
 a18025a <=( a18024a  and  a18019a );
 a18029a <=( (not A268)  and  (not A267) );
 a18030a <=( (not A266)  and  a18029a );
 a18034a <=( A301  and  (not A300) );
 a18035a <=( (not A269)  and  a18034a );
 a18036a <=( a18035a  and  a18030a );
 a18039a <=( A166  and  A167 );
 a18043a <=( A265  and  (not A200) );
 a18044a <=( (not A199)  and  a18043a );
 a18045a <=( a18044a  and  a18039a );
 a18049a <=( (not A268)  and  (not A267) );
 a18050a <=( (not A266)  and  a18049a );
 a18054a <=( A302  and  (not A300) );
 a18055a <=( (not A269)  and  a18054a );
 a18056a <=( a18055a  and  a18050a );
 a18059a <=( A166  and  A167 );
 a18063a <=( A265  and  (not A200) );
 a18064a <=( (not A199)  and  a18063a );
 a18065a <=( a18064a  and  a18059a );
 a18069a <=( (not A268)  and  (not A267) );
 a18070a <=( (not A266)  and  a18069a );
 a18074a <=( A299  and  A298 );
 a18075a <=( (not A269)  and  a18074a );
 a18076a <=( a18075a  and  a18070a );
 a18079a <=( A166  and  A167 );
 a18083a <=( A265  and  (not A200) );
 a18084a <=( (not A199)  and  a18083a );
 a18085a <=( a18084a  and  a18079a );
 a18089a <=( (not A268)  and  (not A267) );
 a18090a <=( (not A266)  and  a18089a );
 a18094a <=( (not A299)  and  (not A298) );
 a18095a <=( (not A269)  and  a18094a );
 a18096a <=( a18095a  and  a18090a );
 a18099a <=( (not A166)  and  (not A167) );
 a18103a <=( (not A203)  and  (not A202) );
 a18104a <=( A201  and  a18103a );
 a18105a <=( a18104a  and  a18099a );
 a18109a <=( A267  and  A266 );
 a18110a <=( (not A265)  and  a18109a );
 a18114a <=( A301  and  (not A300) );
 a18115a <=( A268  and  a18114a );
 a18116a <=( a18115a  and  a18110a );
 a18119a <=( (not A166)  and  (not A167) );
 a18123a <=( (not A203)  and  (not A202) );
 a18124a <=( A201  and  a18123a );
 a18125a <=( a18124a  and  a18119a );
 a18129a <=( A267  and  A266 );
 a18130a <=( (not A265)  and  a18129a );
 a18134a <=( A302  and  (not A300) );
 a18135a <=( A268  and  a18134a );
 a18136a <=( a18135a  and  a18130a );
 a18139a <=( (not A166)  and  (not A167) );
 a18143a <=( (not A203)  and  (not A202) );
 a18144a <=( A201  and  a18143a );
 a18145a <=( a18144a  and  a18139a );
 a18149a <=( A267  and  A266 );
 a18150a <=( (not A265)  and  a18149a );
 a18154a <=( A299  and  A298 );
 a18155a <=( A268  and  a18154a );
 a18156a <=( a18155a  and  a18150a );
 a18159a <=( (not A166)  and  (not A167) );
 a18163a <=( (not A203)  and  (not A202) );
 a18164a <=( A201  and  a18163a );
 a18165a <=( a18164a  and  a18159a );
 a18169a <=( A267  and  A266 );
 a18170a <=( (not A265)  and  a18169a );
 a18174a <=( (not A299)  and  (not A298) );
 a18175a <=( A268  and  a18174a );
 a18176a <=( a18175a  and  a18170a );
 a18179a <=( (not A166)  and  (not A167) );
 a18183a <=( (not A203)  and  (not A202) );
 a18184a <=( A201  and  a18183a );
 a18185a <=( a18184a  and  a18179a );
 a18189a <=( A267  and  A266 );
 a18190a <=( (not A265)  and  a18189a );
 a18194a <=( A301  and  (not A300) );
 a18195a <=( A269  and  a18194a );
 a18196a <=( a18195a  and  a18190a );
 a18199a <=( (not A166)  and  (not A167) );
 a18203a <=( (not A203)  and  (not A202) );
 a18204a <=( A201  and  a18203a );
 a18205a <=( a18204a  and  a18199a );
 a18209a <=( A267  and  A266 );
 a18210a <=( (not A265)  and  a18209a );
 a18214a <=( A302  and  (not A300) );
 a18215a <=( A269  and  a18214a );
 a18216a <=( a18215a  and  a18210a );
 a18219a <=( (not A166)  and  (not A167) );
 a18223a <=( (not A203)  and  (not A202) );
 a18224a <=( A201  and  a18223a );
 a18225a <=( a18224a  and  a18219a );
 a18229a <=( A267  and  A266 );
 a18230a <=( (not A265)  and  a18229a );
 a18234a <=( A299  and  A298 );
 a18235a <=( A269  and  a18234a );
 a18236a <=( a18235a  and  a18230a );
 a18239a <=( (not A166)  and  (not A167) );
 a18243a <=( (not A203)  and  (not A202) );
 a18244a <=( A201  and  a18243a );
 a18245a <=( a18244a  and  a18239a );
 a18249a <=( A267  and  A266 );
 a18250a <=( (not A265)  and  a18249a );
 a18254a <=( (not A299)  and  (not A298) );
 a18255a <=( A269  and  a18254a );
 a18256a <=( a18255a  and  a18250a );
 a18259a <=( (not A166)  and  (not A167) );
 a18263a <=( (not A203)  and  (not A202) );
 a18264a <=( A201  and  a18263a );
 a18265a <=( a18264a  and  a18259a );
 a18269a <=( A267  and  (not A266) );
 a18270a <=( A265  and  a18269a );
 a18274a <=( A301  and  (not A300) );
 a18275a <=( A268  and  a18274a );
 a18276a <=( a18275a  and  a18270a );
 a18279a <=( (not A166)  and  (not A167) );
 a18283a <=( (not A203)  and  (not A202) );
 a18284a <=( A201  and  a18283a );
 a18285a <=( a18284a  and  a18279a );
 a18289a <=( A267  and  (not A266) );
 a18290a <=( A265  and  a18289a );
 a18294a <=( A302  and  (not A300) );
 a18295a <=( A268  and  a18294a );
 a18296a <=( a18295a  and  a18290a );
 a18299a <=( (not A166)  and  (not A167) );
 a18303a <=( (not A203)  and  (not A202) );
 a18304a <=( A201  and  a18303a );
 a18305a <=( a18304a  and  a18299a );
 a18309a <=( A267  and  (not A266) );
 a18310a <=( A265  and  a18309a );
 a18314a <=( A299  and  A298 );
 a18315a <=( A268  and  a18314a );
 a18316a <=( a18315a  and  a18310a );
 a18319a <=( (not A166)  and  (not A167) );
 a18323a <=( (not A203)  and  (not A202) );
 a18324a <=( A201  and  a18323a );
 a18325a <=( a18324a  and  a18319a );
 a18329a <=( A267  and  (not A266) );
 a18330a <=( A265  and  a18329a );
 a18334a <=( (not A299)  and  (not A298) );
 a18335a <=( A268  and  a18334a );
 a18336a <=( a18335a  and  a18330a );
 a18339a <=( (not A166)  and  (not A167) );
 a18343a <=( (not A203)  and  (not A202) );
 a18344a <=( A201  and  a18343a );
 a18345a <=( a18344a  and  a18339a );
 a18349a <=( A267  and  (not A266) );
 a18350a <=( A265  and  a18349a );
 a18354a <=( A301  and  (not A300) );
 a18355a <=( A269  and  a18354a );
 a18356a <=( a18355a  and  a18350a );
 a18359a <=( (not A166)  and  (not A167) );
 a18363a <=( (not A203)  and  (not A202) );
 a18364a <=( A201  and  a18363a );
 a18365a <=( a18364a  and  a18359a );
 a18369a <=( A267  and  (not A266) );
 a18370a <=( A265  and  a18369a );
 a18374a <=( A302  and  (not A300) );
 a18375a <=( A269  and  a18374a );
 a18376a <=( a18375a  and  a18370a );
 a18379a <=( (not A166)  and  (not A167) );
 a18383a <=( (not A203)  and  (not A202) );
 a18384a <=( A201  and  a18383a );
 a18385a <=( a18384a  and  a18379a );
 a18389a <=( A267  and  (not A266) );
 a18390a <=( A265  and  a18389a );
 a18394a <=( A299  and  A298 );
 a18395a <=( A269  and  a18394a );
 a18396a <=( a18395a  and  a18390a );
 a18399a <=( (not A166)  and  (not A167) );
 a18403a <=( (not A203)  and  (not A202) );
 a18404a <=( A201  and  a18403a );
 a18405a <=( a18404a  and  a18399a );
 a18409a <=( A267  and  (not A266) );
 a18410a <=( A265  and  a18409a );
 a18414a <=( (not A299)  and  (not A298) );
 a18415a <=( A269  and  a18414a );
 a18416a <=( a18415a  and  a18410a );
 a18419a <=( (not A166)  and  (not A167) );
 a18423a <=( (not A265)  and  A202 );
 a18424a <=( (not A201)  and  a18423a );
 a18425a <=( a18424a  and  a18419a );
 a18429a <=( A268  and  A267 );
 a18430a <=( A266  and  a18429a );
 a18434a <=( (not A302)  and  (not A301) );
 a18435a <=( A300  and  a18434a );
 a18436a <=( a18435a  and  a18430a );
 a18439a <=( (not A166)  and  (not A167) );
 a18443a <=( (not A265)  and  A202 );
 a18444a <=( (not A201)  and  a18443a );
 a18445a <=( a18444a  and  a18439a );
 a18449a <=( A269  and  A267 );
 a18450a <=( A266  and  a18449a );
 a18454a <=( (not A302)  and  (not A301) );
 a18455a <=( A300  and  a18454a );
 a18456a <=( a18455a  and  a18450a );
 a18459a <=( (not A166)  and  (not A167) );
 a18463a <=( (not A265)  and  A202 );
 a18464a <=( (not A201)  and  a18463a );
 a18465a <=( a18464a  and  a18459a );
 a18469a <=( (not A268)  and  (not A267) );
 a18470a <=( A266  and  a18469a );
 a18474a <=( A301  and  (not A300) );
 a18475a <=( (not A269)  and  a18474a );
 a18476a <=( a18475a  and  a18470a );
 a18479a <=( (not A166)  and  (not A167) );
 a18483a <=( (not A265)  and  A202 );
 a18484a <=( (not A201)  and  a18483a );
 a18485a <=( a18484a  and  a18479a );
 a18489a <=( (not A268)  and  (not A267) );
 a18490a <=( A266  and  a18489a );
 a18494a <=( A302  and  (not A300) );
 a18495a <=( (not A269)  and  a18494a );
 a18496a <=( a18495a  and  a18490a );
 a18499a <=( (not A166)  and  (not A167) );
 a18503a <=( (not A265)  and  A202 );
 a18504a <=( (not A201)  and  a18503a );
 a18505a <=( a18504a  and  a18499a );
 a18509a <=( (not A268)  and  (not A267) );
 a18510a <=( A266  and  a18509a );
 a18514a <=( A299  and  A298 );
 a18515a <=( (not A269)  and  a18514a );
 a18516a <=( a18515a  and  a18510a );
 a18519a <=( (not A166)  and  (not A167) );
 a18523a <=( (not A265)  and  A202 );
 a18524a <=( (not A201)  and  a18523a );
 a18525a <=( a18524a  and  a18519a );
 a18529a <=( (not A268)  and  (not A267) );
 a18530a <=( A266  and  a18529a );
 a18534a <=( (not A299)  and  (not A298) );
 a18535a <=( (not A269)  and  a18534a );
 a18536a <=( a18535a  and  a18530a );
 a18539a <=( (not A166)  and  (not A167) );
 a18543a <=( A265  and  A202 );
 a18544a <=( (not A201)  and  a18543a );
 a18545a <=( a18544a  and  a18539a );
 a18549a <=( A268  and  A267 );
 a18550a <=( (not A266)  and  a18549a );
 a18554a <=( (not A302)  and  (not A301) );
 a18555a <=( A300  and  a18554a );
 a18556a <=( a18555a  and  a18550a );
 a18559a <=( (not A166)  and  (not A167) );
 a18563a <=( A265  and  A202 );
 a18564a <=( (not A201)  and  a18563a );
 a18565a <=( a18564a  and  a18559a );
 a18569a <=( A269  and  A267 );
 a18570a <=( (not A266)  and  a18569a );
 a18574a <=( (not A302)  and  (not A301) );
 a18575a <=( A300  and  a18574a );
 a18576a <=( a18575a  and  a18570a );
 a18579a <=( (not A166)  and  (not A167) );
 a18583a <=( A265  and  A202 );
 a18584a <=( (not A201)  and  a18583a );
 a18585a <=( a18584a  and  a18579a );
 a18589a <=( (not A268)  and  (not A267) );
 a18590a <=( (not A266)  and  a18589a );
 a18594a <=( A301  and  (not A300) );
 a18595a <=( (not A269)  and  a18594a );
 a18596a <=( a18595a  and  a18590a );
 a18599a <=( (not A166)  and  (not A167) );
 a18603a <=( A265  and  A202 );
 a18604a <=( (not A201)  and  a18603a );
 a18605a <=( a18604a  and  a18599a );
 a18609a <=( (not A268)  and  (not A267) );
 a18610a <=( (not A266)  and  a18609a );
 a18614a <=( A302  and  (not A300) );
 a18615a <=( (not A269)  and  a18614a );
 a18616a <=( a18615a  and  a18610a );
 a18619a <=( (not A166)  and  (not A167) );
 a18623a <=( A265  and  A202 );
 a18624a <=( (not A201)  and  a18623a );
 a18625a <=( a18624a  and  a18619a );
 a18629a <=( (not A268)  and  (not A267) );
 a18630a <=( (not A266)  and  a18629a );
 a18634a <=( A299  and  A298 );
 a18635a <=( (not A269)  and  a18634a );
 a18636a <=( a18635a  and  a18630a );
 a18639a <=( (not A166)  and  (not A167) );
 a18643a <=( A265  and  A202 );
 a18644a <=( (not A201)  and  a18643a );
 a18645a <=( a18644a  and  a18639a );
 a18649a <=( (not A268)  and  (not A267) );
 a18650a <=( (not A266)  and  a18649a );
 a18654a <=( (not A299)  and  (not A298) );
 a18655a <=( (not A269)  and  a18654a );
 a18656a <=( a18655a  and  a18650a );
 a18659a <=( (not A166)  and  (not A167) );
 a18663a <=( (not A265)  and  A203 );
 a18664a <=( (not A201)  and  a18663a );
 a18665a <=( a18664a  and  a18659a );
 a18669a <=( A268  and  A267 );
 a18670a <=( A266  and  a18669a );
 a18674a <=( (not A302)  and  (not A301) );
 a18675a <=( A300  and  a18674a );
 a18676a <=( a18675a  and  a18670a );
 a18679a <=( (not A166)  and  (not A167) );
 a18683a <=( (not A265)  and  A203 );
 a18684a <=( (not A201)  and  a18683a );
 a18685a <=( a18684a  and  a18679a );
 a18689a <=( A269  and  A267 );
 a18690a <=( A266  and  a18689a );
 a18694a <=( (not A302)  and  (not A301) );
 a18695a <=( A300  and  a18694a );
 a18696a <=( a18695a  and  a18690a );
 a18699a <=( (not A166)  and  (not A167) );
 a18703a <=( (not A265)  and  A203 );
 a18704a <=( (not A201)  and  a18703a );
 a18705a <=( a18704a  and  a18699a );
 a18709a <=( (not A268)  and  (not A267) );
 a18710a <=( A266  and  a18709a );
 a18714a <=( A301  and  (not A300) );
 a18715a <=( (not A269)  and  a18714a );
 a18716a <=( a18715a  and  a18710a );
 a18719a <=( (not A166)  and  (not A167) );
 a18723a <=( (not A265)  and  A203 );
 a18724a <=( (not A201)  and  a18723a );
 a18725a <=( a18724a  and  a18719a );
 a18729a <=( (not A268)  and  (not A267) );
 a18730a <=( A266  and  a18729a );
 a18734a <=( A302  and  (not A300) );
 a18735a <=( (not A269)  and  a18734a );
 a18736a <=( a18735a  and  a18730a );
 a18739a <=( (not A166)  and  (not A167) );
 a18743a <=( (not A265)  and  A203 );
 a18744a <=( (not A201)  and  a18743a );
 a18745a <=( a18744a  and  a18739a );
 a18749a <=( (not A268)  and  (not A267) );
 a18750a <=( A266  and  a18749a );
 a18754a <=( A299  and  A298 );
 a18755a <=( (not A269)  and  a18754a );
 a18756a <=( a18755a  and  a18750a );
 a18759a <=( (not A166)  and  (not A167) );
 a18763a <=( (not A265)  and  A203 );
 a18764a <=( (not A201)  and  a18763a );
 a18765a <=( a18764a  and  a18759a );
 a18769a <=( (not A268)  and  (not A267) );
 a18770a <=( A266  and  a18769a );
 a18774a <=( (not A299)  and  (not A298) );
 a18775a <=( (not A269)  and  a18774a );
 a18776a <=( a18775a  and  a18770a );
 a18779a <=( (not A166)  and  (not A167) );
 a18783a <=( A265  and  A203 );
 a18784a <=( (not A201)  and  a18783a );
 a18785a <=( a18784a  and  a18779a );
 a18789a <=( A268  and  A267 );
 a18790a <=( (not A266)  and  a18789a );
 a18794a <=( (not A302)  and  (not A301) );
 a18795a <=( A300  and  a18794a );
 a18796a <=( a18795a  and  a18790a );
 a18799a <=( (not A166)  and  (not A167) );
 a18803a <=( A265  and  A203 );
 a18804a <=( (not A201)  and  a18803a );
 a18805a <=( a18804a  and  a18799a );
 a18809a <=( A269  and  A267 );
 a18810a <=( (not A266)  and  a18809a );
 a18814a <=( (not A302)  and  (not A301) );
 a18815a <=( A300  and  a18814a );
 a18816a <=( a18815a  and  a18810a );
 a18819a <=( (not A166)  and  (not A167) );
 a18823a <=( A265  and  A203 );
 a18824a <=( (not A201)  and  a18823a );
 a18825a <=( a18824a  and  a18819a );
 a18829a <=( (not A268)  and  (not A267) );
 a18830a <=( (not A266)  and  a18829a );
 a18834a <=( A301  and  (not A300) );
 a18835a <=( (not A269)  and  a18834a );
 a18836a <=( a18835a  and  a18830a );
 a18839a <=( (not A166)  and  (not A167) );
 a18843a <=( A265  and  A203 );
 a18844a <=( (not A201)  and  a18843a );
 a18845a <=( a18844a  and  a18839a );
 a18849a <=( (not A268)  and  (not A267) );
 a18850a <=( (not A266)  and  a18849a );
 a18854a <=( A302  and  (not A300) );
 a18855a <=( (not A269)  and  a18854a );
 a18856a <=( a18855a  and  a18850a );
 a18859a <=( (not A166)  and  (not A167) );
 a18863a <=( A265  and  A203 );
 a18864a <=( (not A201)  and  a18863a );
 a18865a <=( a18864a  and  a18859a );
 a18869a <=( (not A268)  and  (not A267) );
 a18870a <=( (not A266)  and  a18869a );
 a18874a <=( A299  and  A298 );
 a18875a <=( (not A269)  and  a18874a );
 a18876a <=( a18875a  and  a18870a );
 a18879a <=( (not A166)  and  (not A167) );
 a18883a <=( A265  and  A203 );
 a18884a <=( (not A201)  and  a18883a );
 a18885a <=( a18884a  and  a18879a );
 a18889a <=( (not A268)  and  (not A267) );
 a18890a <=( (not A266)  and  a18889a );
 a18894a <=( (not A299)  and  (not A298) );
 a18895a <=( (not A269)  and  a18894a );
 a18896a <=( a18895a  and  a18890a );
 a18899a <=( (not A166)  and  (not A167) );
 a18903a <=( (not A265)  and  A200 );
 a18904a <=( A199  and  a18903a );
 a18905a <=( a18904a  and  a18899a );
 a18909a <=( A268  and  A267 );
 a18910a <=( A266  and  a18909a );
 a18914a <=( (not A302)  and  (not A301) );
 a18915a <=( A300  and  a18914a );
 a18916a <=( a18915a  and  a18910a );
 a18919a <=( (not A166)  and  (not A167) );
 a18923a <=( (not A265)  and  A200 );
 a18924a <=( A199  and  a18923a );
 a18925a <=( a18924a  and  a18919a );
 a18929a <=( A269  and  A267 );
 a18930a <=( A266  and  a18929a );
 a18934a <=( (not A302)  and  (not A301) );
 a18935a <=( A300  and  a18934a );
 a18936a <=( a18935a  and  a18930a );
 a18939a <=( (not A166)  and  (not A167) );
 a18943a <=( (not A265)  and  A200 );
 a18944a <=( A199  and  a18943a );
 a18945a <=( a18944a  and  a18939a );
 a18949a <=( (not A268)  and  (not A267) );
 a18950a <=( A266  and  a18949a );
 a18954a <=( A301  and  (not A300) );
 a18955a <=( (not A269)  and  a18954a );
 a18956a <=( a18955a  and  a18950a );
 a18959a <=( (not A166)  and  (not A167) );
 a18963a <=( (not A265)  and  A200 );
 a18964a <=( A199  and  a18963a );
 a18965a <=( a18964a  and  a18959a );
 a18969a <=( (not A268)  and  (not A267) );
 a18970a <=( A266  and  a18969a );
 a18974a <=( A302  and  (not A300) );
 a18975a <=( (not A269)  and  a18974a );
 a18976a <=( a18975a  and  a18970a );
 a18979a <=( (not A166)  and  (not A167) );
 a18983a <=( (not A265)  and  A200 );
 a18984a <=( A199  and  a18983a );
 a18985a <=( a18984a  and  a18979a );
 a18989a <=( (not A268)  and  (not A267) );
 a18990a <=( A266  and  a18989a );
 a18994a <=( A299  and  A298 );
 a18995a <=( (not A269)  and  a18994a );
 a18996a <=( a18995a  and  a18990a );
 a18999a <=( (not A166)  and  (not A167) );
 a19003a <=( (not A265)  and  A200 );
 a19004a <=( A199  and  a19003a );
 a19005a <=( a19004a  and  a18999a );
 a19009a <=( (not A268)  and  (not A267) );
 a19010a <=( A266  and  a19009a );
 a19014a <=( (not A299)  and  (not A298) );
 a19015a <=( (not A269)  and  a19014a );
 a19016a <=( a19015a  and  a19010a );
 a19019a <=( (not A166)  and  (not A167) );
 a19023a <=( A265  and  A200 );
 a19024a <=( A199  and  a19023a );
 a19025a <=( a19024a  and  a19019a );
 a19029a <=( A268  and  A267 );
 a19030a <=( (not A266)  and  a19029a );
 a19034a <=( (not A302)  and  (not A301) );
 a19035a <=( A300  and  a19034a );
 a19036a <=( a19035a  and  a19030a );
 a19039a <=( (not A166)  and  (not A167) );
 a19043a <=( A265  and  A200 );
 a19044a <=( A199  and  a19043a );
 a19045a <=( a19044a  and  a19039a );
 a19049a <=( A269  and  A267 );
 a19050a <=( (not A266)  and  a19049a );
 a19054a <=( (not A302)  and  (not A301) );
 a19055a <=( A300  and  a19054a );
 a19056a <=( a19055a  and  a19050a );
 a19059a <=( (not A166)  and  (not A167) );
 a19063a <=( A265  and  A200 );
 a19064a <=( A199  and  a19063a );
 a19065a <=( a19064a  and  a19059a );
 a19069a <=( (not A268)  and  (not A267) );
 a19070a <=( (not A266)  and  a19069a );
 a19074a <=( A301  and  (not A300) );
 a19075a <=( (not A269)  and  a19074a );
 a19076a <=( a19075a  and  a19070a );
 a19079a <=( (not A166)  and  (not A167) );
 a19083a <=( A265  and  A200 );
 a19084a <=( A199  and  a19083a );
 a19085a <=( a19084a  and  a19079a );
 a19089a <=( (not A268)  and  (not A267) );
 a19090a <=( (not A266)  and  a19089a );
 a19094a <=( A302  and  (not A300) );
 a19095a <=( (not A269)  and  a19094a );
 a19096a <=( a19095a  and  a19090a );
 a19099a <=( (not A166)  and  (not A167) );
 a19103a <=( A265  and  A200 );
 a19104a <=( A199  and  a19103a );
 a19105a <=( a19104a  and  a19099a );
 a19109a <=( (not A268)  and  (not A267) );
 a19110a <=( (not A266)  and  a19109a );
 a19114a <=( A299  and  A298 );
 a19115a <=( (not A269)  and  a19114a );
 a19116a <=( a19115a  and  a19110a );
 a19119a <=( (not A166)  and  (not A167) );
 a19123a <=( A265  and  A200 );
 a19124a <=( A199  and  a19123a );
 a19125a <=( a19124a  and  a19119a );
 a19129a <=( (not A268)  and  (not A267) );
 a19130a <=( (not A266)  and  a19129a );
 a19134a <=( (not A299)  and  (not A298) );
 a19135a <=( (not A269)  and  a19134a );
 a19136a <=( a19135a  and  a19130a );
 a19139a <=( (not A166)  and  (not A167) );
 a19143a <=( (not A265)  and  (not A200) );
 a19144a <=( (not A199)  and  a19143a );
 a19145a <=( a19144a  and  a19139a );
 a19149a <=( A268  and  A267 );
 a19150a <=( A266  and  a19149a );
 a19154a <=( (not A302)  and  (not A301) );
 a19155a <=( A300  and  a19154a );
 a19156a <=( a19155a  and  a19150a );
 a19159a <=( (not A166)  and  (not A167) );
 a19163a <=( (not A265)  and  (not A200) );
 a19164a <=( (not A199)  and  a19163a );
 a19165a <=( a19164a  and  a19159a );
 a19169a <=( A269  and  A267 );
 a19170a <=( A266  and  a19169a );
 a19174a <=( (not A302)  and  (not A301) );
 a19175a <=( A300  and  a19174a );
 a19176a <=( a19175a  and  a19170a );
 a19179a <=( (not A166)  and  (not A167) );
 a19183a <=( (not A265)  and  (not A200) );
 a19184a <=( (not A199)  and  a19183a );
 a19185a <=( a19184a  and  a19179a );
 a19189a <=( (not A268)  and  (not A267) );
 a19190a <=( A266  and  a19189a );
 a19194a <=( A301  and  (not A300) );
 a19195a <=( (not A269)  and  a19194a );
 a19196a <=( a19195a  and  a19190a );
 a19199a <=( (not A166)  and  (not A167) );
 a19203a <=( (not A265)  and  (not A200) );
 a19204a <=( (not A199)  and  a19203a );
 a19205a <=( a19204a  and  a19199a );
 a19209a <=( (not A268)  and  (not A267) );
 a19210a <=( A266  and  a19209a );
 a19214a <=( A302  and  (not A300) );
 a19215a <=( (not A269)  and  a19214a );
 a19216a <=( a19215a  and  a19210a );
 a19219a <=( (not A166)  and  (not A167) );
 a19223a <=( (not A265)  and  (not A200) );
 a19224a <=( (not A199)  and  a19223a );
 a19225a <=( a19224a  and  a19219a );
 a19229a <=( (not A268)  and  (not A267) );
 a19230a <=( A266  and  a19229a );
 a19234a <=( A299  and  A298 );
 a19235a <=( (not A269)  and  a19234a );
 a19236a <=( a19235a  and  a19230a );
 a19239a <=( (not A166)  and  (not A167) );
 a19243a <=( (not A265)  and  (not A200) );
 a19244a <=( (not A199)  and  a19243a );
 a19245a <=( a19244a  and  a19239a );
 a19249a <=( (not A268)  and  (not A267) );
 a19250a <=( A266  and  a19249a );
 a19254a <=( (not A299)  and  (not A298) );
 a19255a <=( (not A269)  and  a19254a );
 a19256a <=( a19255a  and  a19250a );
 a19259a <=( (not A166)  and  (not A167) );
 a19263a <=( A265  and  (not A200) );
 a19264a <=( (not A199)  and  a19263a );
 a19265a <=( a19264a  and  a19259a );
 a19269a <=( A268  and  A267 );
 a19270a <=( (not A266)  and  a19269a );
 a19274a <=( (not A302)  and  (not A301) );
 a19275a <=( A300  and  a19274a );
 a19276a <=( a19275a  and  a19270a );
 a19279a <=( (not A166)  and  (not A167) );
 a19283a <=( A265  and  (not A200) );
 a19284a <=( (not A199)  and  a19283a );
 a19285a <=( a19284a  and  a19279a );
 a19289a <=( A269  and  A267 );
 a19290a <=( (not A266)  and  a19289a );
 a19294a <=( (not A302)  and  (not A301) );
 a19295a <=( A300  and  a19294a );
 a19296a <=( a19295a  and  a19290a );
 a19299a <=( (not A166)  and  (not A167) );
 a19303a <=( A265  and  (not A200) );
 a19304a <=( (not A199)  and  a19303a );
 a19305a <=( a19304a  and  a19299a );
 a19309a <=( (not A268)  and  (not A267) );
 a19310a <=( (not A266)  and  a19309a );
 a19314a <=( A301  and  (not A300) );
 a19315a <=( (not A269)  and  a19314a );
 a19316a <=( a19315a  and  a19310a );
 a19319a <=( (not A166)  and  (not A167) );
 a19323a <=( A265  and  (not A200) );
 a19324a <=( (not A199)  and  a19323a );
 a19325a <=( a19324a  and  a19319a );
 a19329a <=( (not A268)  and  (not A267) );
 a19330a <=( (not A266)  and  a19329a );
 a19334a <=( A302  and  (not A300) );
 a19335a <=( (not A269)  and  a19334a );
 a19336a <=( a19335a  and  a19330a );
 a19339a <=( (not A166)  and  (not A167) );
 a19343a <=( A265  and  (not A200) );
 a19344a <=( (not A199)  and  a19343a );
 a19345a <=( a19344a  and  a19339a );
 a19349a <=( (not A268)  and  (not A267) );
 a19350a <=( (not A266)  and  a19349a );
 a19354a <=( A299  and  A298 );
 a19355a <=( (not A269)  and  a19354a );
 a19356a <=( a19355a  and  a19350a );
 a19359a <=( (not A166)  and  (not A167) );
 a19363a <=( A265  and  (not A200) );
 a19364a <=( (not A199)  and  a19363a );
 a19365a <=( a19364a  and  a19359a );
 a19369a <=( (not A268)  and  (not A267) );
 a19370a <=( (not A266)  and  a19369a );
 a19374a <=( (not A299)  and  (not A298) );
 a19375a <=( (not A269)  and  a19374a );
 a19376a <=( a19375a  and  a19370a );
 a19379a <=( (not A168)  and  (not A170) );
 a19383a <=( (not A203)  and  (not A202) );
 a19384a <=( A201  and  a19383a );
 a19385a <=( a19384a  and  a19379a );
 a19389a <=( A267  and  A266 );
 a19390a <=( (not A265)  and  a19389a );
 a19394a <=( A301  and  (not A300) );
 a19395a <=( A268  and  a19394a );
 a19396a <=( a19395a  and  a19390a );
 a19399a <=( (not A168)  and  (not A170) );
 a19403a <=( (not A203)  and  (not A202) );
 a19404a <=( A201  and  a19403a );
 a19405a <=( a19404a  and  a19399a );
 a19409a <=( A267  and  A266 );
 a19410a <=( (not A265)  and  a19409a );
 a19414a <=( A302  and  (not A300) );
 a19415a <=( A268  and  a19414a );
 a19416a <=( a19415a  and  a19410a );
 a19419a <=( (not A168)  and  (not A170) );
 a19423a <=( (not A203)  and  (not A202) );
 a19424a <=( A201  and  a19423a );
 a19425a <=( a19424a  and  a19419a );
 a19429a <=( A267  and  A266 );
 a19430a <=( (not A265)  and  a19429a );
 a19434a <=( A299  and  A298 );
 a19435a <=( A268  and  a19434a );
 a19436a <=( a19435a  and  a19430a );
 a19439a <=( (not A168)  and  (not A170) );
 a19443a <=( (not A203)  and  (not A202) );
 a19444a <=( A201  and  a19443a );
 a19445a <=( a19444a  and  a19439a );
 a19449a <=( A267  and  A266 );
 a19450a <=( (not A265)  and  a19449a );
 a19454a <=( (not A299)  and  (not A298) );
 a19455a <=( A268  and  a19454a );
 a19456a <=( a19455a  and  a19450a );
 a19459a <=( (not A168)  and  (not A170) );
 a19463a <=( (not A203)  and  (not A202) );
 a19464a <=( A201  and  a19463a );
 a19465a <=( a19464a  and  a19459a );
 a19469a <=( A267  and  A266 );
 a19470a <=( (not A265)  and  a19469a );
 a19474a <=( A301  and  (not A300) );
 a19475a <=( A269  and  a19474a );
 a19476a <=( a19475a  and  a19470a );
 a19479a <=( (not A168)  and  (not A170) );
 a19483a <=( (not A203)  and  (not A202) );
 a19484a <=( A201  and  a19483a );
 a19485a <=( a19484a  and  a19479a );
 a19489a <=( A267  and  A266 );
 a19490a <=( (not A265)  and  a19489a );
 a19494a <=( A302  and  (not A300) );
 a19495a <=( A269  and  a19494a );
 a19496a <=( a19495a  and  a19490a );
 a19499a <=( (not A168)  and  (not A170) );
 a19503a <=( (not A203)  and  (not A202) );
 a19504a <=( A201  and  a19503a );
 a19505a <=( a19504a  and  a19499a );
 a19509a <=( A267  and  A266 );
 a19510a <=( (not A265)  and  a19509a );
 a19514a <=( A299  and  A298 );
 a19515a <=( A269  and  a19514a );
 a19516a <=( a19515a  and  a19510a );
 a19519a <=( (not A168)  and  (not A170) );
 a19523a <=( (not A203)  and  (not A202) );
 a19524a <=( A201  and  a19523a );
 a19525a <=( a19524a  and  a19519a );
 a19529a <=( A267  and  A266 );
 a19530a <=( (not A265)  and  a19529a );
 a19534a <=( (not A299)  and  (not A298) );
 a19535a <=( A269  and  a19534a );
 a19536a <=( a19535a  and  a19530a );
 a19539a <=( (not A168)  and  (not A170) );
 a19543a <=( (not A203)  and  (not A202) );
 a19544a <=( A201  and  a19543a );
 a19545a <=( a19544a  and  a19539a );
 a19549a <=( A267  and  (not A266) );
 a19550a <=( A265  and  a19549a );
 a19554a <=( A301  and  (not A300) );
 a19555a <=( A268  and  a19554a );
 a19556a <=( a19555a  and  a19550a );
 a19559a <=( (not A168)  and  (not A170) );
 a19563a <=( (not A203)  and  (not A202) );
 a19564a <=( A201  and  a19563a );
 a19565a <=( a19564a  and  a19559a );
 a19569a <=( A267  and  (not A266) );
 a19570a <=( A265  and  a19569a );
 a19574a <=( A302  and  (not A300) );
 a19575a <=( A268  and  a19574a );
 a19576a <=( a19575a  and  a19570a );
 a19579a <=( (not A168)  and  (not A170) );
 a19583a <=( (not A203)  and  (not A202) );
 a19584a <=( A201  and  a19583a );
 a19585a <=( a19584a  and  a19579a );
 a19589a <=( A267  and  (not A266) );
 a19590a <=( A265  and  a19589a );
 a19594a <=( A299  and  A298 );
 a19595a <=( A268  and  a19594a );
 a19596a <=( a19595a  and  a19590a );
 a19599a <=( (not A168)  and  (not A170) );
 a19603a <=( (not A203)  and  (not A202) );
 a19604a <=( A201  and  a19603a );
 a19605a <=( a19604a  and  a19599a );
 a19609a <=( A267  and  (not A266) );
 a19610a <=( A265  and  a19609a );
 a19614a <=( (not A299)  and  (not A298) );
 a19615a <=( A268  and  a19614a );
 a19616a <=( a19615a  and  a19610a );
 a19619a <=( (not A168)  and  (not A170) );
 a19623a <=( (not A203)  and  (not A202) );
 a19624a <=( A201  and  a19623a );
 a19625a <=( a19624a  and  a19619a );
 a19629a <=( A267  and  (not A266) );
 a19630a <=( A265  and  a19629a );
 a19634a <=( A301  and  (not A300) );
 a19635a <=( A269  and  a19634a );
 a19636a <=( a19635a  and  a19630a );
 a19639a <=( (not A168)  and  (not A170) );
 a19643a <=( (not A203)  and  (not A202) );
 a19644a <=( A201  and  a19643a );
 a19645a <=( a19644a  and  a19639a );
 a19649a <=( A267  and  (not A266) );
 a19650a <=( A265  and  a19649a );
 a19654a <=( A302  and  (not A300) );
 a19655a <=( A269  and  a19654a );
 a19656a <=( a19655a  and  a19650a );
 a19659a <=( (not A168)  and  (not A170) );
 a19663a <=( (not A203)  and  (not A202) );
 a19664a <=( A201  and  a19663a );
 a19665a <=( a19664a  and  a19659a );
 a19669a <=( A267  and  (not A266) );
 a19670a <=( A265  and  a19669a );
 a19674a <=( A299  and  A298 );
 a19675a <=( A269  and  a19674a );
 a19676a <=( a19675a  and  a19670a );
 a19679a <=( (not A168)  and  (not A170) );
 a19683a <=( (not A203)  and  (not A202) );
 a19684a <=( A201  and  a19683a );
 a19685a <=( a19684a  and  a19679a );
 a19689a <=( A267  and  (not A266) );
 a19690a <=( A265  and  a19689a );
 a19694a <=( (not A299)  and  (not A298) );
 a19695a <=( A269  and  a19694a );
 a19696a <=( a19695a  and  a19690a );
 a19699a <=( (not A168)  and  (not A170) );
 a19703a <=( (not A265)  and  A202 );
 a19704a <=( (not A201)  and  a19703a );
 a19705a <=( a19704a  and  a19699a );
 a19709a <=( A268  and  A267 );
 a19710a <=( A266  and  a19709a );
 a19714a <=( (not A302)  and  (not A301) );
 a19715a <=( A300  and  a19714a );
 a19716a <=( a19715a  and  a19710a );
 a19719a <=( (not A168)  and  (not A170) );
 a19723a <=( (not A265)  and  A202 );
 a19724a <=( (not A201)  and  a19723a );
 a19725a <=( a19724a  and  a19719a );
 a19729a <=( A269  and  A267 );
 a19730a <=( A266  and  a19729a );
 a19734a <=( (not A302)  and  (not A301) );
 a19735a <=( A300  and  a19734a );
 a19736a <=( a19735a  and  a19730a );
 a19739a <=( (not A168)  and  (not A170) );
 a19743a <=( (not A265)  and  A202 );
 a19744a <=( (not A201)  and  a19743a );
 a19745a <=( a19744a  and  a19739a );
 a19749a <=( (not A268)  and  (not A267) );
 a19750a <=( A266  and  a19749a );
 a19754a <=( A301  and  (not A300) );
 a19755a <=( (not A269)  and  a19754a );
 a19756a <=( a19755a  and  a19750a );
 a19759a <=( (not A168)  and  (not A170) );
 a19763a <=( (not A265)  and  A202 );
 a19764a <=( (not A201)  and  a19763a );
 a19765a <=( a19764a  and  a19759a );
 a19769a <=( (not A268)  and  (not A267) );
 a19770a <=( A266  and  a19769a );
 a19774a <=( A302  and  (not A300) );
 a19775a <=( (not A269)  and  a19774a );
 a19776a <=( a19775a  and  a19770a );
 a19779a <=( (not A168)  and  (not A170) );
 a19783a <=( (not A265)  and  A202 );
 a19784a <=( (not A201)  and  a19783a );
 a19785a <=( a19784a  and  a19779a );
 a19789a <=( (not A268)  and  (not A267) );
 a19790a <=( A266  and  a19789a );
 a19794a <=( A299  and  A298 );
 a19795a <=( (not A269)  and  a19794a );
 a19796a <=( a19795a  and  a19790a );
 a19799a <=( (not A168)  and  (not A170) );
 a19803a <=( (not A265)  and  A202 );
 a19804a <=( (not A201)  and  a19803a );
 a19805a <=( a19804a  and  a19799a );
 a19809a <=( (not A268)  and  (not A267) );
 a19810a <=( A266  and  a19809a );
 a19814a <=( (not A299)  and  (not A298) );
 a19815a <=( (not A269)  and  a19814a );
 a19816a <=( a19815a  and  a19810a );
 a19819a <=( (not A168)  and  (not A170) );
 a19823a <=( A265  and  A202 );
 a19824a <=( (not A201)  and  a19823a );
 a19825a <=( a19824a  and  a19819a );
 a19829a <=( A268  and  A267 );
 a19830a <=( (not A266)  and  a19829a );
 a19834a <=( (not A302)  and  (not A301) );
 a19835a <=( A300  and  a19834a );
 a19836a <=( a19835a  and  a19830a );
 a19839a <=( (not A168)  and  (not A170) );
 a19843a <=( A265  and  A202 );
 a19844a <=( (not A201)  and  a19843a );
 a19845a <=( a19844a  and  a19839a );
 a19849a <=( A269  and  A267 );
 a19850a <=( (not A266)  and  a19849a );
 a19854a <=( (not A302)  and  (not A301) );
 a19855a <=( A300  and  a19854a );
 a19856a <=( a19855a  and  a19850a );
 a19859a <=( (not A168)  and  (not A170) );
 a19863a <=( A265  and  A202 );
 a19864a <=( (not A201)  and  a19863a );
 a19865a <=( a19864a  and  a19859a );
 a19869a <=( (not A268)  and  (not A267) );
 a19870a <=( (not A266)  and  a19869a );
 a19874a <=( A301  and  (not A300) );
 a19875a <=( (not A269)  and  a19874a );
 a19876a <=( a19875a  and  a19870a );
 a19879a <=( (not A168)  and  (not A170) );
 a19883a <=( A265  and  A202 );
 a19884a <=( (not A201)  and  a19883a );
 a19885a <=( a19884a  and  a19879a );
 a19889a <=( (not A268)  and  (not A267) );
 a19890a <=( (not A266)  and  a19889a );
 a19894a <=( A302  and  (not A300) );
 a19895a <=( (not A269)  and  a19894a );
 a19896a <=( a19895a  and  a19890a );
 a19899a <=( (not A168)  and  (not A170) );
 a19903a <=( A265  and  A202 );
 a19904a <=( (not A201)  and  a19903a );
 a19905a <=( a19904a  and  a19899a );
 a19909a <=( (not A268)  and  (not A267) );
 a19910a <=( (not A266)  and  a19909a );
 a19914a <=( A299  and  A298 );
 a19915a <=( (not A269)  and  a19914a );
 a19916a <=( a19915a  and  a19910a );
 a19919a <=( (not A168)  and  (not A170) );
 a19923a <=( A265  and  A202 );
 a19924a <=( (not A201)  and  a19923a );
 a19925a <=( a19924a  and  a19919a );
 a19929a <=( (not A268)  and  (not A267) );
 a19930a <=( (not A266)  and  a19929a );
 a19934a <=( (not A299)  and  (not A298) );
 a19935a <=( (not A269)  and  a19934a );
 a19936a <=( a19935a  and  a19930a );
 a19939a <=( (not A168)  and  (not A170) );
 a19943a <=( (not A265)  and  A203 );
 a19944a <=( (not A201)  and  a19943a );
 a19945a <=( a19944a  and  a19939a );
 a19949a <=( A268  and  A267 );
 a19950a <=( A266  and  a19949a );
 a19954a <=( (not A302)  and  (not A301) );
 a19955a <=( A300  and  a19954a );
 a19956a <=( a19955a  and  a19950a );
 a19959a <=( (not A168)  and  (not A170) );
 a19963a <=( (not A265)  and  A203 );
 a19964a <=( (not A201)  and  a19963a );
 a19965a <=( a19964a  and  a19959a );
 a19969a <=( A269  and  A267 );
 a19970a <=( A266  and  a19969a );
 a19974a <=( (not A302)  and  (not A301) );
 a19975a <=( A300  and  a19974a );
 a19976a <=( a19975a  and  a19970a );
 a19979a <=( (not A168)  and  (not A170) );
 a19983a <=( (not A265)  and  A203 );
 a19984a <=( (not A201)  and  a19983a );
 a19985a <=( a19984a  and  a19979a );
 a19989a <=( (not A268)  and  (not A267) );
 a19990a <=( A266  and  a19989a );
 a19994a <=( A301  and  (not A300) );
 a19995a <=( (not A269)  and  a19994a );
 a19996a <=( a19995a  and  a19990a );
 a19999a <=( (not A168)  and  (not A170) );
 a20003a <=( (not A265)  and  A203 );
 a20004a <=( (not A201)  and  a20003a );
 a20005a <=( a20004a  and  a19999a );
 a20009a <=( (not A268)  and  (not A267) );
 a20010a <=( A266  and  a20009a );
 a20014a <=( A302  and  (not A300) );
 a20015a <=( (not A269)  and  a20014a );
 a20016a <=( a20015a  and  a20010a );
 a20019a <=( (not A168)  and  (not A170) );
 a20023a <=( (not A265)  and  A203 );
 a20024a <=( (not A201)  and  a20023a );
 a20025a <=( a20024a  and  a20019a );
 a20029a <=( (not A268)  and  (not A267) );
 a20030a <=( A266  and  a20029a );
 a20034a <=( A299  and  A298 );
 a20035a <=( (not A269)  and  a20034a );
 a20036a <=( a20035a  and  a20030a );
 a20039a <=( (not A168)  and  (not A170) );
 a20043a <=( (not A265)  and  A203 );
 a20044a <=( (not A201)  and  a20043a );
 a20045a <=( a20044a  and  a20039a );
 a20049a <=( (not A268)  and  (not A267) );
 a20050a <=( A266  and  a20049a );
 a20054a <=( (not A299)  and  (not A298) );
 a20055a <=( (not A269)  and  a20054a );
 a20056a <=( a20055a  and  a20050a );
 a20059a <=( (not A168)  and  (not A170) );
 a20063a <=( A265  and  A203 );
 a20064a <=( (not A201)  and  a20063a );
 a20065a <=( a20064a  and  a20059a );
 a20069a <=( A268  and  A267 );
 a20070a <=( (not A266)  and  a20069a );
 a20074a <=( (not A302)  and  (not A301) );
 a20075a <=( A300  and  a20074a );
 a20076a <=( a20075a  and  a20070a );
 a20079a <=( (not A168)  and  (not A170) );
 a20083a <=( A265  and  A203 );
 a20084a <=( (not A201)  and  a20083a );
 a20085a <=( a20084a  and  a20079a );
 a20089a <=( A269  and  A267 );
 a20090a <=( (not A266)  and  a20089a );
 a20094a <=( (not A302)  and  (not A301) );
 a20095a <=( A300  and  a20094a );
 a20096a <=( a20095a  and  a20090a );
 a20099a <=( (not A168)  and  (not A170) );
 a20103a <=( A265  and  A203 );
 a20104a <=( (not A201)  and  a20103a );
 a20105a <=( a20104a  and  a20099a );
 a20109a <=( (not A268)  and  (not A267) );
 a20110a <=( (not A266)  and  a20109a );
 a20114a <=( A301  and  (not A300) );
 a20115a <=( (not A269)  and  a20114a );
 a20116a <=( a20115a  and  a20110a );
 a20119a <=( (not A168)  and  (not A170) );
 a20123a <=( A265  and  A203 );
 a20124a <=( (not A201)  and  a20123a );
 a20125a <=( a20124a  and  a20119a );
 a20129a <=( (not A268)  and  (not A267) );
 a20130a <=( (not A266)  and  a20129a );
 a20134a <=( A302  and  (not A300) );
 a20135a <=( (not A269)  and  a20134a );
 a20136a <=( a20135a  and  a20130a );
 a20139a <=( (not A168)  and  (not A170) );
 a20143a <=( A265  and  A203 );
 a20144a <=( (not A201)  and  a20143a );
 a20145a <=( a20144a  and  a20139a );
 a20149a <=( (not A268)  and  (not A267) );
 a20150a <=( (not A266)  and  a20149a );
 a20154a <=( A299  and  A298 );
 a20155a <=( (not A269)  and  a20154a );
 a20156a <=( a20155a  and  a20150a );
 a20159a <=( (not A168)  and  (not A170) );
 a20163a <=( A265  and  A203 );
 a20164a <=( (not A201)  and  a20163a );
 a20165a <=( a20164a  and  a20159a );
 a20169a <=( (not A268)  and  (not A267) );
 a20170a <=( (not A266)  and  a20169a );
 a20174a <=( (not A299)  and  (not A298) );
 a20175a <=( (not A269)  and  a20174a );
 a20176a <=( a20175a  and  a20170a );
 a20179a <=( (not A168)  and  (not A170) );
 a20183a <=( (not A265)  and  A200 );
 a20184a <=( A199  and  a20183a );
 a20185a <=( a20184a  and  a20179a );
 a20189a <=( A268  and  A267 );
 a20190a <=( A266  and  a20189a );
 a20194a <=( (not A302)  and  (not A301) );
 a20195a <=( A300  and  a20194a );
 a20196a <=( a20195a  and  a20190a );
 a20199a <=( (not A168)  and  (not A170) );
 a20203a <=( (not A265)  and  A200 );
 a20204a <=( A199  and  a20203a );
 a20205a <=( a20204a  and  a20199a );
 a20209a <=( A269  and  A267 );
 a20210a <=( A266  and  a20209a );
 a20214a <=( (not A302)  and  (not A301) );
 a20215a <=( A300  and  a20214a );
 a20216a <=( a20215a  and  a20210a );
 a20219a <=( (not A168)  and  (not A170) );
 a20223a <=( (not A265)  and  A200 );
 a20224a <=( A199  and  a20223a );
 a20225a <=( a20224a  and  a20219a );
 a20229a <=( (not A268)  and  (not A267) );
 a20230a <=( A266  and  a20229a );
 a20234a <=( A301  and  (not A300) );
 a20235a <=( (not A269)  and  a20234a );
 a20236a <=( a20235a  and  a20230a );
 a20239a <=( (not A168)  and  (not A170) );
 a20243a <=( (not A265)  and  A200 );
 a20244a <=( A199  and  a20243a );
 a20245a <=( a20244a  and  a20239a );
 a20249a <=( (not A268)  and  (not A267) );
 a20250a <=( A266  and  a20249a );
 a20254a <=( A302  and  (not A300) );
 a20255a <=( (not A269)  and  a20254a );
 a20256a <=( a20255a  and  a20250a );
 a20259a <=( (not A168)  and  (not A170) );
 a20263a <=( (not A265)  and  A200 );
 a20264a <=( A199  and  a20263a );
 a20265a <=( a20264a  and  a20259a );
 a20269a <=( (not A268)  and  (not A267) );
 a20270a <=( A266  and  a20269a );
 a20274a <=( A299  and  A298 );
 a20275a <=( (not A269)  and  a20274a );
 a20276a <=( a20275a  and  a20270a );
 a20279a <=( (not A168)  and  (not A170) );
 a20283a <=( (not A265)  and  A200 );
 a20284a <=( A199  and  a20283a );
 a20285a <=( a20284a  and  a20279a );
 a20289a <=( (not A268)  and  (not A267) );
 a20290a <=( A266  and  a20289a );
 a20294a <=( (not A299)  and  (not A298) );
 a20295a <=( (not A269)  and  a20294a );
 a20296a <=( a20295a  and  a20290a );
 a20299a <=( (not A168)  and  (not A170) );
 a20303a <=( A265  and  A200 );
 a20304a <=( A199  and  a20303a );
 a20305a <=( a20304a  and  a20299a );
 a20309a <=( A268  and  A267 );
 a20310a <=( (not A266)  and  a20309a );
 a20314a <=( (not A302)  and  (not A301) );
 a20315a <=( A300  and  a20314a );
 a20316a <=( a20315a  and  a20310a );
 a20319a <=( (not A168)  and  (not A170) );
 a20323a <=( A265  and  A200 );
 a20324a <=( A199  and  a20323a );
 a20325a <=( a20324a  and  a20319a );
 a20329a <=( A269  and  A267 );
 a20330a <=( (not A266)  and  a20329a );
 a20334a <=( (not A302)  and  (not A301) );
 a20335a <=( A300  and  a20334a );
 a20336a <=( a20335a  and  a20330a );
 a20339a <=( (not A168)  and  (not A170) );
 a20343a <=( A265  and  A200 );
 a20344a <=( A199  and  a20343a );
 a20345a <=( a20344a  and  a20339a );
 a20349a <=( (not A268)  and  (not A267) );
 a20350a <=( (not A266)  and  a20349a );
 a20354a <=( A301  and  (not A300) );
 a20355a <=( (not A269)  and  a20354a );
 a20356a <=( a20355a  and  a20350a );
 a20359a <=( (not A168)  and  (not A170) );
 a20363a <=( A265  and  A200 );
 a20364a <=( A199  and  a20363a );
 a20365a <=( a20364a  and  a20359a );
 a20369a <=( (not A268)  and  (not A267) );
 a20370a <=( (not A266)  and  a20369a );
 a20374a <=( A302  and  (not A300) );
 a20375a <=( (not A269)  and  a20374a );
 a20376a <=( a20375a  and  a20370a );
 a20379a <=( (not A168)  and  (not A170) );
 a20383a <=( A265  and  A200 );
 a20384a <=( A199  and  a20383a );
 a20385a <=( a20384a  and  a20379a );
 a20389a <=( (not A268)  and  (not A267) );
 a20390a <=( (not A266)  and  a20389a );
 a20394a <=( A299  and  A298 );
 a20395a <=( (not A269)  and  a20394a );
 a20396a <=( a20395a  and  a20390a );
 a20399a <=( (not A168)  and  (not A170) );
 a20403a <=( A265  and  A200 );
 a20404a <=( A199  and  a20403a );
 a20405a <=( a20404a  and  a20399a );
 a20409a <=( (not A268)  and  (not A267) );
 a20410a <=( (not A266)  and  a20409a );
 a20414a <=( (not A299)  and  (not A298) );
 a20415a <=( (not A269)  and  a20414a );
 a20416a <=( a20415a  and  a20410a );
 a20419a <=( (not A168)  and  (not A170) );
 a20423a <=( (not A265)  and  (not A200) );
 a20424a <=( (not A199)  and  a20423a );
 a20425a <=( a20424a  and  a20419a );
 a20429a <=( A268  and  A267 );
 a20430a <=( A266  and  a20429a );
 a20434a <=( (not A302)  and  (not A301) );
 a20435a <=( A300  and  a20434a );
 a20436a <=( a20435a  and  a20430a );
 a20439a <=( (not A168)  and  (not A170) );
 a20443a <=( (not A265)  and  (not A200) );
 a20444a <=( (not A199)  and  a20443a );
 a20445a <=( a20444a  and  a20439a );
 a20449a <=( A269  and  A267 );
 a20450a <=( A266  and  a20449a );
 a20454a <=( (not A302)  and  (not A301) );
 a20455a <=( A300  and  a20454a );
 a20456a <=( a20455a  and  a20450a );
 a20459a <=( (not A168)  and  (not A170) );
 a20463a <=( (not A265)  and  (not A200) );
 a20464a <=( (not A199)  and  a20463a );
 a20465a <=( a20464a  and  a20459a );
 a20469a <=( (not A268)  and  (not A267) );
 a20470a <=( A266  and  a20469a );
 a20474a <=( A301  and  (not A300) );
 a20475a <=( (not A269)  and  a20474a );
 a20476a <=( a20475a  and  a20470a );
 a20479a <=( (not A168)  and  (not A170) );
 a20483a <=( (not A265)  and  (not A200) );
 a20484a <=( (not A199)  and  a20483a );
 a20485a <=( a20484a  and  a20479a );
 a20489a <=( (not A268)  and  (not A267) );
 a20490a <=( A266  and  a20489a );
 a20494a <=( A302  and  (not A300) );
 a20495a <=( (not A269)  and  a20494a );
 a20496a <=( a20495a  and  a20490a );
 a20499a <=( (not A168)  and  (not A170) );
 a20503a <=( (not A265)  and  (not A200) );
 a20504a <=( (not A199)  and  a20503a );
 a20505a <=( a20504a  and  a20499a );
 a20509a <=( (not A268)  and  (not A267) );
 a20510a <=( A266  and  a20509a );
 a20514a <=( A299  and  A298 );
 a20515a <=( (not A269)  and  a20514a );
 a20516a <=( a20515a  and  a20510a );
 a20519a <=( (not A168)  and  (not A170) );
 a20523a <=( (not A265)  and  (not A200) );
 a20524a <=( (not A199)  and  a20523a );
 a20525a <=( a20524a  and  a20519a );
 a20529a <=( (not A268)  and  (not A267) );
 a20530a <=( A266  and  a20529a );
 a20534a <=( (not A299)  and  (not A298) );
 a20535a <=( (not A269)  and  a20534a );
 a20536a <=( a20535a  and  a20530a );
 a20539a <=( (not A168)  and  (not A170) );
 a20543a <=( A265  and  (not A200) );
 a20544a <=( (not A199)  and  a20543a );
 a20545a <=( a20544a  and  a20539a );
 a20549a <=( A268  and  A267 );
 a20550a <=( (not A266)  and  a20549a );
 a20554a <=( (not A302)  and  (not A301) );
 a20555a <=( A300  and  a20554a );
 a20556a <=( a20555a  and  a20550a );
 a20559a <=( (not A168)  and  (not A170) );
 a20563a <=( A265  and  (not A200) );
 a20564a <=( (not A199)  and  a20563a );
 a20565a <=( a20564a  and  a20559a );
 a20569a <=( A269  and  A267 );
 a20570a <=( (not A266)  and  a20569a );
 a20574a <=( (not A302)  and  (not A301) );
 a20575a <=( A300  and  a20574a );
 a20576a <=( a20575a  and  a20570a );
 a20579a <=( (not A168)  and  (not A170) );
 a20583a <=( A265  and  (not A200) );
 a20584a <=( (not A199)  and  a20583a );
 a20585a <=( a20584a  and  a20579a );
 a20589a <=( (not A268)  and  (not A267) );
 a20590a <=( (not A266)  and  a20589a );
 a20594a <=( A301  and  (not A300) );
 a20595a <=( (not A269)  and  a20594a );
 a20596a <=( a20595a  and  a20590a );
 a20599a <=( (not A168)  and  (not A170) );
 a20603a <=( A265  and  (not A200) );
 a20604a <=( (not A199)  and  a20603a );
 a20605a <=( a20604a  and  a20599a );
 a20609a <=( (not A268)  and  (not A267) );
 a20610a <=( (not A266)  and  a20609a );
 a20614a <=( A302  and  (not A300) );
 a20615a <=( (not A269)  and  a20614a );
 a20616a <=( a20615a  and  a20610a );
 a20619a <=( (not A168)  and  (not A170) );
 a20623a <=( A265  and  (not A200) );
 a20624a <=( (not A199)  and  a20623a );
 a20625a <=( a20624a  and  a20619a );
 a20629a <=( (not A268)  and  (not A267) );
 a20630a <=( (not A266)  and  a20629a );
 a20634a <=( A299  and  A298 );
 a20635a <=( (not A269)  and  a20634a );
 a20636a <=( a20635a  and  a20630a );
 a20639a <=( (not A168)  and  (not A170) );
 a20643a <=( A265  and  (not A200) );
 a20644a <=( (not A199)  and  a20643a );
 a20645a <=( a20644a  and  a20639a );
 a20649a <=( (not A268)  and  (not A267) );
 a20650a <=( (not A266)  and  a20649a );
 a20654a <=( (not A299)  and  (not A298) );
 a20655a <=( (not A269)  and  a20654a );
 a20656a <=( a20655a  and  a20650a );
 a20659a <=( (not A168)  and  A169 );
 a20663a <=( (not A203)  and  (not A202) );
 a20664a <=( A201  and  a20663a );
 a20665a <=( a20664a  and  a20659a );
 a20669a <=( A267  and  A266 );
 a20670a <=( (not A265)  and  a20669a );
 a20674a <=( A301  and  (not A300) );
 a20675a <=( A268  and  a20674a );
 a20676a <=( a20675a  and  a20670a );
 a20679a <=( (not A168)  and  A169 );
 a20683a <=( (not A203)  and  (not A202) );
 a20684a <=( A201  and  a20683a );
 a20685a <=( a20684a  and  a20679a );
 a20689a <=( A267  and  A266 );
 a20690a <=( (not A265)  and  a20689a );
 a20694a <=( A302  and  (not A300) );
 a20695a <=( A268  and  a20694a );
 a20696a <=( a20695a  and  a20690a );
 a20699a <=( (not A168)  and  A169 );
 a20703a <=( (not A203)  and  (not A202) );
 a20704a <=( A201  and  a20703a );
 a20705a <=( a20704a  and  a20699a );
 a20709a <=( A267  and  A266 );
 a20710a <=( (not A265)  and  a20709a );
 a20714a <=( A299  and  A298 );
 a20715a <=( A268  and  a20714a );
 a20716a <=( a20715a  and  a20710a );
 a20719a <=( (not A168)  and  A169 );
 a20723a <=( (not A203)  and  (not A202) );
 a20724a <=( A201  and  a20723a );
 a20725a <=( a20724a  and  a20719a );
 a20729a <=( A267  and  A266 );
 a20730a <=( (not A265)  and  a20729a );
 a20734a <=( (not A299)  and  (not A298) );
 a20735a <=( A268  and  a20734a );
 a20736a <=( a20735a  and  a20730a );
 a20739a <=( (not A168)  and  A169 );
 a20743a <=( (not A203)  and  (not A202) );
 a20744a <=( A201  and  a20743a );
 a20745a <=( a20744a  and  a20739a );
 a20749a <=( A267  and  A266 );
 a20750a <=( (not A265)  and  a20749a );
 a20754a <=( A301  and  (not A300) );
 a20755a <=( A269  and  a20754a );
 a20756a <=( a20755a  and  a20750a );
 a20759a <=( (not A168)  and  A169 );
 a20763a <=( (not A203)  and  (not A202) );
 a20764a <=( A201  and  a20763a );
 a20765a <=( a20764a  and  a20759a );
 a20769a <=( A267  and  A266 );
 a20770a <=( (not A265)  and  a20769a );
 a20774a <=( A302  and  (not A300) );
 a20775a <=( A269  and  a20774a );
 a20776a <=( a20775a  and  a20770a );
 a20779a <=( (not A168)  and  A169 );
 a20783a <=( (not A203)  and  (not A202) );
 a20784a <=( A201  and  a20783a );
 a20785a <=( a20784a  and  a20779a );
 a20789a <=( A267  and  A266 );
 a20790a <=( (not A265)  and  a20789a );
 a20794a <=( A299  and  A298 );
 a20795a <=( A269  and  a20794a );
 a20796a <=( a20795a  and  a20790a );
 a20799a <=( (not A168)  and  A169 );
 a20803a <=( (not A203)  and  (not A202) );
 a20804a <=( A201  and  a20803a );
 a20805a <=( a20804a  and  a20799a );
 a20809a <=( A267  and  A266 );
 a20810a <=( (not A265)  and  a20809a );
 a20814a <=( (not A299)  and  (not A298) );
 a20815a <=( A269  and  a20814a );
 a20816a <=( a20815a  and  a20810a );
 a20819a <=( (not A168)  and  A169 );
 a20823a <=( (not A203)  and  (not A202) );
 a20824a <=( A201  and  a20823a );
 a20825a <=( a20824a  and  a20819a );
 a20829a <=( A267  and  (not A266) );
 a20830a <=( A265  and  a20829a );
 a20834a <=( A301  and  (not A300) );
 a20835a <=( A268  and  a20834a );
 a20836a <=( a20835a  and  a20830a );
 a20839a <=( (not A168)  and  A169 );
 a20843a <=( (not A203)  and  (not A202) );
 a20844a <=( A201  and  a20843a );
 a20845a <=( a20844a  and  a20839a );
 a20849a <=( A267  and  (not A266) );
 a20850a <=( A265  and  a20849a );
 a20854a <=( A302  and  (not A300) );
 a20855a <=( A268  and  a20854a );
 a20856a <=( a20855a  and  a20850a );
 a20859a <=( (not A168)  and  A169 );
 a20863a <=( (not A203)  and  (not A202) );
 a20864a <=( A201  and  a20863a );
 a20865a <=( a20864a  and  a20859a );
 a20869a <=( A267  and  (not A266) );
 a20870a <=( A265  and  a20869a );
 a20874a <=( A299  and  A298 );
 a20875a <=( A268  and  a20874a );
 a20876a <=( a20875a  and  a20870a );
 a20879a <=( (not A168)  and  A169 );
 a20883a <=( (not A203)  and  (not A202) );
 a20884a <=( A201  and  a20883a );
 a20885a <=( a20884a  and  a20879a );
 a20889a <=( A267  and  (not A266) );
 a20890a <=( A265  and  a20889a );
 a20894a <=( (not A299)  and  (not A298) );
 a20895a <=( A268  and  a20894a );
 a20896a <=( a20895a  and  a20890a );
 a20899a <=( (not A168)  and  A169 );
 a20903a <=( (not A203)  and  (not A202) );
 a20904a <=( A201  and  a20903a );
 a20905a <=( a20904a  and  a20899a );
 a20909a <=( A267  and  (not A266) );
 a20910a <=( A265  and  a20909a );
 a20914a <=( A301  and  (not A300) );
 a20915a <=( A269  and  a20914a );
 a20916a <=( a20915a  and  a20910a );
 a20919a <=( (not A168)  and  A169 );
 a20923a <=( (not A203)  and  (not A202) );
 a20924a <=( A201  and  a20923a );
 a20925a <=( a20924a  and  a20919a );
 a20929a <=( A267  and  (not A266) );
 a20930a <=( A265  and  a20929a );
 a20934a <=( A302  and  (not A300) );
 a20935a <=( A269  and  a20934a );
 a20936a <=( a20935a  and  a20930a );
 a20939a <=( (not A168)  and  A169 );
 a20943a <=( (not A203)  and  (not A202) );
 a20944a <=( A201  and  a20943a );
 a20945a <=( a20944a  and  a20939a );
 a20949a <=( A267  and  (not A266) );
 a20950a <=( A265  and  a20949a );
 a20954a <=( A299  and  A298 );
 a20955a <=( A269  and  a20954a );
 a20956a <=( a20955a  and  a20950a );
 a20959a <=( (not A168)  and  A169 );
 a20963a <=( (not A203)  and  (not A202) );
 a20964a <=( A201  and  a20963a );
 a20965a <=( a20964a  and  a20959a );
 a20969a <=( A267  and  (not A266) );
 a20970a <=( A265  and  a20969a );
 a20974a <=( (not A299)  and  (not A298) );
 a20975a <=( A269  and  a20974a );
 a20976a <=( a20975a  and  a20970a );
 a20979a <=( (not A168)  and  A169 );
 a20983a <=( (not A265)  and  A202 );
 a20984a <=( (not A201)  and  a20983a );
 a20985a <=( a20984a  and  a20979a );
 a20989a <=( A268  and  A267 );
 a20990a <=( A266  and  a20989a );
 a20994a <=( (not A302)  and  (not A301) );
 a20995a <=( A300  and  a20994a );
 a20996a <=( a20995a  and  a20990a );
 a20999a <=( (not A168)  and  A169 );
 a21003a <=( (not A265)  and  A202 );
 a21004a <=( (not A201)  and  a21003a );
 a21005a <=( a21004a  and  a20999a );
 a21009a <=( A269  and  A267 );
 a21010a <=( A266  and  a21009a );
 a21014a <=( (not A302)  and  (not A301) );
 a21015a <=( A300  and  a21014a );
 a21016a <=( a21015a  and  a21010a );
 a21019a <=( (not A168)  and  A169 );
 a21023a <=( (not A265)  and  A202 );
 a21024a <=( (not A201)  and  a21023a );
 a21025a <=( a21024a  and  a21019a );
 a21029a <=( (not A268)  and  (not A267) );
 a21030a <=( A266  and  a21029a );
 a21034a <=( A301  and  (not A300) );
 a21035a <=( (not A269)  and  a21034a );
 a21036a <=( a21035a  and  a21030a );
 a21039a <=( (not A168)  and  A169 );
 a21043a <=( (not A265)  and  A202 );
 a21044a <=( (not A201)  and  a21043a );
 a21045a <=( a21044a  and  a21039a );
 a21049a <=( (not A268)  and  (not A267) );
 a21050a <=( A266  and  a21049a );
 a21054a <=( A302  and  (not A300) );
 a21055a <=( (not A269)  and  a21054a );
 a21056a <=( a21055a  and  a21050a );
 a21059a <=( (not A168)  and  A169 );
 a21063a <=( (not A265)  and  A202 );
 a21064a <=( (not A201)  and  a21063a );
 a21065a <=( a21064a  and  a21059a );
 a21069a <=( (not A268)  and  (not A267) );
 a21070a <=( A266  and  a21069a );
 a21074a <=( A299  and  A298 );
 a21075a <=( (not A269)  and  a21074a );
 a21076a <=( a21075a  and  a21070a );
 a21079a <=( (not A168)  and  A169 );
 a21083a <=( (not A265)  and  A202 );
 a21084a <=( (not A201)  and  a21083a );
 a21085a <=( a21084a  and  a21079a );
 a21089a <=( (not A268)  and  (not A267) );
 a21090a <=( A266  and  a21089a );
 a21094a <=( (not A299)  and  (not A298) );
 a21095a <=( (not A269)  and  a21094a );
 a21096a <=( a21095a  and  a21090a );
 a21099a <=( (not A168)  and  A169 );
 a21103a <=( A265  and  A202 );
 a21104a <=( (not A201)  and  a21103a );
 a21105a <=( a21104a  and  a21099a );
 a21109a <=( A268  and  A267 );
 a21110a <=( (not A266)  and  a21109a );
 a21114a <=( (not A302)  and  (not A301) );
 a21115a <=( A300  and  a21114a );
 a21116a <=( a21115a  and  a21110a );
 a21119a <=( (not A168)  and  A169 );
 a21123a <=( A265  and  A202 );
 a21124a <=( (not A201)  and  a21123a );
 a21125a <=( a21124a  and  a21119a );
 a21129a <=( A269  and  A267 );
 a21130a <=( (not A266)  and  a21129a );
 a21134a <=( (not A302)  and  (not A301) );
 a21135a <=( A300  and  a21134a );
 a21136a <=( a21135a  and  a21130a );
 a21139a <=( (not A168)  and  A169 );
 a21143a <=( A265  and  A202 );
 a21144a <=( (not A201)  and  a21143a );
 a21145a <=( a21144a  and  a21139a );
 a21149a <=( (not A268)  and  (not A267) );
 a21150a <=( (not A266)  and  a21149a );
 a21154a <=( A301  and  (not A300) );
 a21155a <=( (not A269)  and  a21154a );
 a21156a <=( a21155a  and  a21150a );
 a21159a <=( (not A168)  and  A169 );
 a21163a <=( A265  and  A202 );
 a21164a <=( (not A201)  and  a21163a );
 a21165a <=( a21164a  and  a21159a );
 a21169a <=( (not A268)  and  (not A267) );
 a21170a <=( (not A266)  and  a21169a );
 a21174a <=( A302  and  (not A300) );
 a21175a <=( (not A269)  and  a21174a );
 a21176a <=( a21175a  and  a21170a );
 a21179a <=( (not A168)  and  A169 );
 a21183a <=( A265  and  A202 );
 a21184a <=( (not A201)  and  a21183a );
 a21185a <=( a21184a  and  a21179a );
 a21189a <=( (not A268)  and  (not A267) );
 a21190a <=( (not A266)  and  a21189a );
 a21194a <=( A299  and  A298 );
 a21195a <=( (not A269)  and  a21194a );
 a21196a <=( a21195a  and  a21190a );
 a21199a <=( (not A168)  and  A169 );
 a21203a <=( A265  and  A202 );
 a21204a <=( (not A201)  and  a21203a );
 a21205a <=( a21204a  and  a21199a );
 a21209a <=( (not A268)  and  (not A267) );
 a21210a <=( (not A266)  and  a21209a );
 a21214a <=( (not A299)  and  (not A298) );
 a21215a <=( (not A269)  and  a21214a );
 a21216a <=( a21215a  and  a21210a );
 a21219a <=( (not A168)  and  A169 );
 a21223a <=( (not A265)  and  A203 );
 a21224a <=( (not A201)  and  a21223a );
 a21225a <=( a21224a  and  a21219a );
 a21229a <=( A268  and  A267 );
 a21230a <=( A266  and  a21229a );
 a21234a <=( (not A302)  and  (not A301) );
 a21235a <=( A300  and  a21234a );
 a21236a <=( a21235a  and  a21230a );
 a21239a <=( (not A168)  and  A169 );
 a21243a <=( (not A265)  and  A203 );
 a21244a <=( (not A201)  and  a21243a );
 a21245a <=( a21244a  and  a21239a );
 a21249a <=( A269  and  A267 );
 a21250a <=( A266  and  a21249a );
 a21254a <=( (not A302)  and  (not A301) );
 a21255a <=( A300  and  a21254a );
 a21256a <=( a21255a  and  a21250a );
 a21259a <=( (not A168)  and  A169 );
 a21263a <=( (not A265)  and  A203 );
 a21264a <=( (not A201)  and  a21263a );
 a21265a <=( a21264a  and  a21259a );
 a21269a <=( (not A268)  and  (not A267) );
 a21270a <=( A266  and  a21269a );
 a21274a <=( A301  and  (not A300) );
 a21275a <=( (not A269)  and  a21274a );
 a21276a <=( a21275a  and  a21270a );
 a21279a <=( (not A168)  and  A169 );
 a21283a <=( (not A265)  and  A203 );
 a21284a <=( (not A201)  and  a21283a );
 a21285a <=( a21284a  and  a21279a );
 a21289a <=( (not A268)  and  (not A267) );
 a21290a <=( A266  and  a21289a );
 a21294a <=( A302  and  (not A300) );
 a21295a <=( (not A269)  and  a21294a );
 a21296a <=( a21295a  and  a21290a );
 a21299a <=( (not A168)  and  A169 );
 a21303a <=( (not A265)  and  A203 );
 a21304a <=( (not A201)  and  a21303a );
 a21305a <=( a21304a  and  a21299a );
 a21309a <=( (not A268)  and  (not A267) );
 a21310a <=( A266  and  a21309a );
 a21314a <=( A299  and  A298 );
 a21315a <=( (not A269)  and  a21314a );
 a21316a <=( a21315a  and  a21310a );
 a21319a <=( (not A168)  and  A169 );
 a21323a <=( (not A265)  and  A203 );
 a21324a <=( (not A201)  and  a21323a );
 a21325a <=( a21324a  and  a21319a );
 a21329a <=( (not A268)  and  (not A267) );
 a21330a <=( A266  and  a21329a );
 a21334a <=( (not A299)  and  (not A298) );
 a21335a <=( (not A269)  and  a21334a );
 a21336a <=( a21335a  and  a21330a );
 a21339a <=( (not A168)  and  A169 );
 a21343a <=( A265  and  A203 );
 a21344a <=( (not A201)  and  a21343a );
 a21345a <=( a21344a  and  a21339a );
 a21349a <=( A268  and  A267 );
 a21350a <=( (not A266)  and  a21349a );
 a21354a <=( (not A302)  and  (not A301) );
 a21355a <=( A300  and  a21354a );
 a21356a <=( a21355a  and  a21350a );
 a21359a <=( (not A168)  and  A169 );
 a21363a <=( A265  and  A203 );
 a21364a <=( (not A201)  and  a21363a );
 a21365a <=( a21364a  and  a21359a );
 a21369a <=( A269  and  A267 );
 a21370a <=( (not A266)  and  a21369a );
 a21374a <=( (not A302)  and  (not A301) );
 a21375a <=( A300  and  a21374a );
 a21376a <=( a21375a  and  a21370a );
 a21379a <=( (not A168)  and  A169 );
 a21383a <=( A265  and  A203 );
 a21384a <=( (not A201)  and  a21383a );
 a21385a <=( a21384a  and  a21379a );
 a21389a <=( (not A268)  and  (not A267) );
 a21390a <=( (not A266)  and  a21389a );
 a21394a <=( A301  and  (not A300) );
 a21395a <=( (not A269)  and  a21394a );
 a21396a <=( a21395a  and  a21390a );
 a21399a <=( (not A168)  and  A169 );
 a21403a <=( A265  and  A203 );
 a21404a <=( (not A201)  and  a21403a );
 a21405a <=( a21404a  and  a21399a );
 a21409a <=( (not A268)  and  (not A267) );
 a21410a <=( (not A266)  and  a21409a );
 a21414a <=( A302  and  (not A300) );
 a21415a <=( (not A269)  and  a21414a );
 a21416a <=( a21415a  and  a21410a );
 a21419a <=( (not A168)  and  A169 );
 a21423a <=( A265  and  A203 );
 a21424a <=( (not A201)  and  a21423a );
 a21425a <=( a21424a  and  a21419a );
 a21429a <=( (not A268)  and  (not A267) );
 a21430a <=( (not A266)  and  a21429a );
 a21434a <=( A299  and  A298 );
 a21435a <=( (not A269)  and  a21434a );
 a21436a <=( a21435a  and  a21430a );
 a21439a <=( (not A168)  and  A169 );
 a21443a <=( A265  and  A203 );
 a21444a <=( (not A201)  and  a21443a );
 a21445a <=( a21444a  and  a21439a );
 a21449a <=( (not A268)  and  (not A267) );
 a21450a <=( (not A266)  and  a21449a );
 a21454a <=( (not A299)  and  (not A298) );
 a21455a <=( (not A269)  and  a21454a );
 a21456a <=( a21455a  and  a21450a );
 a21459a <=( (not A168)  and  A169 );
 a21463a <=( (not A265)  and  A200 );
 a21464a <=( A199  and  a21463a );
 a21465a <=( a21464a  and  a21459a );
 a21469a <=( A268  and  A267 );
 a21470a <=( A266  and  a21469a );
 a21474a <=( (not A302)  and  (not A301) );
 a21475a <=( A300  and  a21474a );
 a21476a <=( a21475a  and  a21470a );
 a21479a <=( (not A168)  and  A169 );
 a21483a <=( (not A265)  and  A200 );
 a21484a <=( A199  and  a21483a );
 a21485a <=( a21484a  and  a21479a );
 a21489a <=( A269  and  A267 );
 a21490a <=( A266  and  a21489a );
 a21494a <=( (not A302)  and  (not A301) );
 a21495a <=( A300  and  a21494a );
 a21496a <=( a21495a  and  a21490a );
 a21499a <=( (not A168)  and  A169 );
 a21503a <=( (not A265)  and  A200 );
 a21504a <=( A199  and  a21503a );
 a21505a <=( a21504a  and  a21499a );
 a21509a <=( (not A268)  and  (not A267) );
 a21510a <=( A266  and  a21509a );
 a21514a <=( A301  and  (not A300) );
 a21515a <=( (not A269)  and  a21514a );
 a21516a <=( a21515a  and  a21510a );
 a21519a <=( (not A168)  and  A169 );
 a21523a <=( (not A265)  and  A200 );
 a21524a <=( A199  and  a21523a );
 a21525a <=( a21524a  and  a21519a );
 a21529a <=( (not A268)  and  (not A267) );
 a21530a <=( A266  and  a21529a );
 a21534a <=( A302  and  (not A300) );
 a21535a <=( (not A269)  and  a21534a );
 a21536a <=( a21535a  and  a21530a );
 a21539a <=( (not A168)  and  A169 );
 a21543a <=( (not A265)  and  A200 );
 a21544a <=( A199  and  a21543a );
 a21545a <=( a21544a  and  a21539a );
 a21549a <=( (not A268)  and  (not A267) );
 a21550a <=( A266  and  a21549a );
 a21554a <=( A299  and  A298 );
 a21555a <=( (not A269)  and  a21554a );
 a21556a <=( a21555a  and  a21550a );
 a21559a <=( (not A168)  and  A169 );
 a21563a <=( (not A265)  and  A200 );
 a21564a <=( A199  and  a21563a );
 a21565a <=( a21564a  and  a21559a );
 a21569a <=( (not A268)  and  (not A267) );
 a21570a <=( A266  and  a21569a );
 a21574a <=( (not A299)  and  (not A298) );
 a21575a <=( (not A269)  and  a21574a );
 a21576a <=( a21575a  and  a21570a );
 a21579a <=( (not A168)  and  A169 );
 a21583a <=( A265  and  A200 );
 a21584a <=( A199  and  a21583a );
 a21585a <=( a21584a  and  a21579a );
 a21589a <=( A268  and  A267 );
 a21590a <=( (not A266)  and  a21589a );
 a21594a <=( (not A302)  and  (not A301) );
 a21595a <=( A300  and  a21594a );
 a21596a <=( a21595a  and  a21590a );
 a21599a <=( (not A168)  and  A169 );
 a21603a <=( A265  and  A200 );
 a21604a <=( A199  and  a21603a );
 a21605a <=( a21604a  and  a21599a );
 a21609a <=( A269  and  A267 );
 a21610a <=( (not A266)  and  a21609a );
 a21614a <=( (not A302)  and  (not A301) );
 a21615a <=( A300  and  a21614a );
 a21616a <=( a21615a  and  a21610a );
 a21619a <=( (not A168)  and  A169 );
 a21623a <=( A265  and  A200 );
 a21624a <=( A199  and  a21623a );
 a21625a <=( a21624a  and  a21619a );
 a21629a <=( (not A268)  and  (not A267) );
 a21630a <=( (not A266)  and  a21629a );
 a21634a <=( A301  and  (not A300) );
 a21635a <=( (not A269)  and  a21634a );
 a21636a <=( a21635a  and  a21630a );
 a21639a <=( (not A168)  and  A169 );
 a21643a <=( A265  and  A200 );
 a21644a <=( A199  and  a21643a );
 a21645a <=( a21644a  and  a21639a );
 a21649a <=( (not A268)  and  (not A267) );
 a21650a <=( (not A266)  and  a21649a );
 a21654a <=( A302  and  (not A300) );
 a21655a <=( (not A269)  and  a21654a );
 a21656a <=( a21655a  and  a21650a );
 a21659a <=( (not A168)  and  A169 );
 a21663a <=( A265  and  A200 );
 a21664a <=( A199  and  a21663a );
 a21665a <=( a21664a  and  a21659a );
 a21669a <=( (not A268)  and  (not A267) );
 a21670a <=( (not A266)  and  a21669a );
 a21674a <=( A299  and  A298 );
 a21675a <=( (not A269)  and  a21674a );
 a21676a <=( a21675a  and  a21670a );
 a21679a <=( (not A168)  and  A169 );
 a21683a <=( A265  and  A200 );
 a21684a <=( A199  and  a21683a );
 a21685a <=( a21684a  and  a21679a );
 a21689a <=( (not A268)  and  (not A267) );
 a21690a <=( (not A266)  and  a21689a );
 a21694a <=( (not A299)  and  (not A298) );
 a21695a <=( (not A269)  and  a21694a );
 a21696a <=( a21695a  and  a21690a );
 a21699a <=( (not A168)  and  A169 );
 a21703a <=( (not A265)  and  (not A200) );
 a21704a <=( (not A199)  and  a21703a );
 a21705a <=( a21704a  and  a21699a );
 a21709a <=( A268  and  A267 );
 a21710a <=( A266  and  a21709a );
 a21714a <=( (not A302)  and  (not A301) );
 a21715a <=( A300  and  a21714a );
 a21716a <=( a21715a  and  a21710a );
 a21719a <=( (not A168)  and  A169 );
 a21723a <=( (not A265)  and  (not A200) );
 a21724a <=( (not A199)  and  a21723a );
 a21725a <=( a21724a  and  a21719a );
 a21729a <=( A269  and  A267 );
 a21730a <=( A266  and  a21729a );
 a21734a <=( (not A302)  and  (not A301) );
 a21735a <=( A300  and  a21734a );
 a21736a <=( a21735a  and  a21730a );
 a21739a <=( (not A168)  and  A169 );
 a21743a <=( (not A265)  and  (not A200) );
 a21744a <=( (not A199)  and  a21743a );
 a21745a <=( a21744a  and  a21739a );
 a21749a <=( (not A268)  and  (not A267) );
 a21750a <=( A266  and  a21749a );
 a21754a <=( A301  and  (not A300) );
 a21755a <=( (not A269)  and  a21754a );
 a21756a <=( a21755a  and  a21750a );
 a21759a <=( (not A168)  and  A169 );
 a21763a <=( (not A265)  and  (not A200) );
 a21764a <=( (not A199)  and  a21763a );
 a21765a <=( a21764a  and  a21759a );
 a21769a <=( (not A268)  and  (not A267) );
 a21770a <=( A266  and  a21769a );
 a21774a <=( A302  and  (not A300) );
 a21775a <=( (not A269)  and  a21774a );
 a21776a <=( a21775a  and  a21770a );
 a21779a <=( (not A168)  and  A169 );
 a21783a <=( (not A265)  and  (not A200) );
 a21784a <=( (not A199)  and  a21783a );
 a21785a <=( a21784a  and  a21779a );
 a21789a <=( (not A268)  and  (not A267) );
 a21790a <=( A266  and  a21789a );
 a21794a <=( A299  and  A298 );
 a21795a <=( (not A269)  and  a21794a );
 a21796a <=( a21795a  and  a21790a );
 a21799a <=( (not A168)  and  A169 );
 a21803a <=( (not A265)  and  (not A200) );
 a21804a <=( (not A199)  and  a21803a );
 a21805a <=( a21804a  and  a21799a );
 a21809a <=( (not A268)  and  (not A267) );
 a21810a <=( A266  and  a21809a );
 a21814a <=( (not A299)  and  (not A298) );
 a21815a <=( (not A269)  and  a21814a );
 a21816a <=( a21815a  and  a21810a );
 a21819a <=( (not A168)  and  A169 );
 a21823a <=( A265  and  (not A200) );
 a21824a <=( (not A199)  and  a21823a );
 a21825a <=( a21824a  and  a21819a );
 a21829a <=( A268  and  A267 );
 a21830a <=( (not A266)  and  a21829a );
 a21834a <=( (not A302)  and  (not A301) );
 a21835a <=( A300  and  a21834a );
 a21836a <=( a21835a  and  a21830a );
 a21839a <=( (not A168)  and  A169 );
 a21843a <=( A265  and  (not A200) );
 a21844a <=( (not A199)  and  a21843a );
 a21845a <=( a21844a  and  a21839a );
 a21849a <=( A269  and  A267 );
 a21850a <=( (not A266)  and  a21849a );
 a21854a <=( (not A302)  and  (not A301) );
 a21855a <=( A300  and  a21854a );
 a21856a <=( a21855a  and  a21850a );
 a21859a <=( (not A168)  and  A169 );
 a21863a <=( A265  and  (not A200) );
 a21864a <=( (not A199)  and  a21863a );
 a21865a <=( a21864a  and  a21859a );
 a21869a <=( (not A268)  and  (not A267) );
 a21870a <=( (not A266)  and  a21869a );
 a21874a <=( A301  and  (not A300) );
 a21875a <=( (not A269)  and  a21874a );
 a21876a <=( a21875a  and  a21870a );
 a21879a <=( (not A168)  and  A169 );
 a21883a <=( A265  and  (not A200) );
 a21884a <=( (not A199)  and  a21883a );
 a21885a <=( a21884a  and  a21879a );
 a21889a <=( (not A268)  and  (not A267) );
 a21890a <=( (not A266)  and  a21889a );
 a21894a <=( A302  and  (not A300) );
 a21895a <=( (not A269)  and  a21894a );
 a21896a <=( a21895a  and  a21890a );
 a21899a <=( (not A168)  and  A169 );
 a21903a <=( A265  and  (not A200) );
 a21904a <=( (not A199)  and  a21903a );
 a21905a <=( a21904a  and  a21899a );
 a21909a <=( (not A268)  and  (not A267) );
 a21910a <=( (not A266)  and  a21909a );
 a21914a <=( A299  and  A298 );
 a21915a <=( (not A269)  and  a21914a );
 a21916a <=( a21915a  and  a21910a );
 a21919a <=( (not A168)  and  A169 );
 a21923a <=( A265  and  (not A200) );
 a21924a <=( (not A199)  and  a21923a );
 a21925a <=( a21924a  and  a21919a );
 a21929a <=( (not A268)  and  (not A267) );
 a21930a <=( (not A266)  and  a21929a );
 a21934a <=( (not A299)  and  (not A298) );
 a21935a <=( (not A269)  and  a21934a );
 a21936a <=( a21935a  and  a21930a );
 a21939a <=( (not A169)  and  A170 );
 a21943a <=( A202  and  (not A201) );
 a21944a <=( A168  and  a21943a );
 a21945a <=( a21944a  and  a21939a );
 a21949a <=( A267  and  A266 );
 a21950a <=( (not A265)  and  a21949a );
 a21954a <=( A301  and  (not A300) );
 a21955a <=( A268  and  a21954a );
 a21956a <=( a21955a  and  a21950a );
 a21959a <=( (not A169)  and  A170 );
 a21963a <=( A202  and  (not A201) );
 a21964a <=( A168  and  a21963a );
 a21965a <=( a21964a  and  a21959a );
 a21969a <=( A267  and  A266 );
 a21970a <=( (not A265)  and  a21969a );
 a21974a <=( A302  and  (not A300) );
 a21975a <=( A268  and  a21974a );
 a21976a <=( a21975a  and  a21970a );
 a21979a <=( (not A169)  and  A170 );
 a21983a <=( A202  and  (not A201) );
 a21984a <=( A168  and  a21983a );
 a21985a <=( a21984a  and  a21979a );
 a21989a <=( A267  and  A266 );
 a21990a <=( (not A265)  and  a21989a );
 a21994a <=( A299  and  A298 );
 a21995a <=( A268  and  a21994a );
 a21996a <=( a21995a  and  a21990a );
 a21999a <=( (not A169)  and  A170 );
 a22003a <=( A202  and  (not A201) );
 a22004a <=( A168  and  a22003a );
 a22005a <=( a22004a  and  a21999a );
 a22009a <=( A267  and  A266 );
 a22010a <=( (not A265)  and  a22009a );
 a22014a <=( (not A299)  and  (not A298) );
 a22015a <=( A268  and  a22014a );
 a22016a <=( a22015a  and  a22010a );
 a22019a <=( (not A169)  and  A170 );
 a22023a <=( A202  and  (not A201) );
 a22024a <=( A168  and  a22023a );
 a22025a <=( a22024a  and  a22019a );
 a22029a <=( A267  and  A266 );
 a22030a <=( (not A265)  and  a22029a );
 a22034a <=( A301  and  (not A300) );
 a22035a <=( A269  and  a22034a );
 a22036a <=( a22035a  and  a22030a );
 a22039a <=( (not A169)  and  A170 );
 a22043a <=( A202  and  (not A201) );
 a22044a <=( A168  and  a22043a );
 a22045a <=( a22044a  and  a22039a );
 a22049a <=( A267  and  A266 );
 a22050a <=( (not A265)  and  a22049a );
 a22054a <=( A302  and  (not A300) );
 a22055a <=( A269  and  a22054a );
 a22056a <=( a22055a  and  a22050a );
 a22059a <=( (not A169)  and  A170 );
 a22063a <=( A202  and  (not A201) );
 a22064a <=( A168  and  a22063a );
 a22065a <=( a22064a  and  a22059a );
 a22069a <=( A267  and  A266 );
 a22070a <=( (not A265)  and  a22069a );
 a22074a <=( A299  and  A298 );
 a22075a <=( A269  and  a22074a );
 a22076a <=( a22075a  and  a22070a );
 a22079a <=( (not A169)  and  A170 );
 a22083a <=( A202  and  (not A201) );
 a22084a <=( A168  and  a22083a );
 a22085a <=( a22084a  and  a22079a );
 a22089a <=( A267  and  A266 );
 a22090a <=( (not A265)  and  a22089a );
 a22094a <=( (not A299)  and  (not A298) );
 a22095a <=( A269  and  a22094a );
 a22096a <=( a22095a  and  a22090a );
 a22099a <=( (not A169)  and  A170 );
 a22103a <=( A202  and  (not A201) );
 a22104a <=( A168  and  a22103a );
 a22105a <=( a22104a  and  a22099a );
 a22109a <=( A267  and  (not A266) );
 a22110a <=( A265  and  a22109a );
 a22114a <=( A301  and  (not A300) );
 a22115a <=( A268  and  a22114a );
 a22116a <=( a22115a  and  a22110a );
 a22119a <=( (not A169)  and  A170 );
 a22123a <=( A202  and  (not A201) );
 a22124a <=( A168  and  a22123a );
 a22125a <=( a22124a  and  a22119a );
 a22129a <=( A267  and  (not A266) );
 a22130a <=( A265  and  a22129a );
 a22134a <=( A302  and  (not A300) );
 a22135a <=( A268  and  a22134a );
 a22136a <=( a22135a  and  a22130a );
 a22139a <=( (not A169)  and  A170 );
 a22143a <=( A202  and  (not A201) );
 a22144a <=( A168  and  a22143a );
 a22145a <=( a22144a  and  a22139a );
 a22149a <=( A267  and  (not A266) );
 a22150a <=( A265  and  a22149a );
 a22154a <=( A299  and  A298 );
 a22155a <=( A268  and  a22154a );
 a22156a <=( a22155a  and  a22150a );
 a22159a <=( (not A169)  and  A170 );
 a22163a <=( A202  and  (not A201) );
 a22164a <=( A168  and  a22163a );
 a22165a <=( a22164a  and  a22159a );
 a22169a <=( A267  and  (not A266) );
 a22170a <=( A265  and  a22169a );
 a22174a <=( (not A299)  and  (not A298) );
 a22175a <=( A268  and  a22174a );
 a22176a <=( a22175a  and  a22170a );
 a22179a <=( (not A169)  and  A170 );
 a22183a <=( A202  and  (not A201) );
 a22184a <=( A168  and  a22183a );
 a22185a <=( a22184a  and  a22179a );
 a22189a <=( A267  and  (not A266) );
 a22190a <=( A265  and  a22189a );
 a22194a <=( A301  and  (not A300) );
 a22195a <=( A269  and  a22194a );
 a22196a <=( a22195a  and  a22190a );
 a22199a <=( (not A169)  and  A170 );
 a22203a <=( A202  and  (not A201) );
 a22204a <=( A168  and  a22203a );
 a22205a <=( a22204a  and  a22199a );
 a22209a <=( A267  and  (not A266) );
 a22210a <=( A265  and  a22209a );
 a22214a <=( A302  and  (not A300) );
 a22215a <=( A269  and  a22214a );
 a22216a <=( a22215a  and  a22210a );
 a22219a <=( (not A169)  and  A170 );
 a22223a <=( A202  and  (not A201) );
 a22224a <=( A168  and  a22223a );
 a22225a <=( a22224a  and  a22219a );
 a22229a <=( A267  and  (not A266) );
 a22230a <=( A265  and  a22229a );
 a22234a <=( A299  and  A298 );
 a22235a <=( A269  and  a22234a );
 a22236a <=( a22235a  and  a22230a );
 a22239a <=( (not A169)  and  A170 );
 a22243a <=( A202  and  (not A201) );
 a22244a <=( A168  and  a22243a );
 a22245a <=( a22244a  and  a22239a );
 a22249a <=( A267  and  (not A266) );
 a22250a <=( A265  and  a22249a );
 a22254a <=( (not A299)  and  (not A298) );
 a22255a <=( A269  and  a22254a );
 a22256a <=( a22255a  and  a22250a );
 a22259a <=( (not A169)  and  A170 );
 a22263a <=( A203  and  (not A201) );
 a22264a <=( A168  and  a22263a );
 a22265a <=( a22264a  and  a22259a );
 a22269a <=( A267  and  A266 );
 a22270a <=( (not A265)  and  a22269a );
 a22274a <=( A301  and  (not A300) );
 a22275a <=( A268  and  a22274a );
 a22276a <=( a22275a  and  a22270a );
 a22279a <=( (not A169)  and  A170 );
 a22283a <=( A203  and  (not A201) );
 a22284a <=( A168  and  a22283a );
 a22285a <=( a22284a  and  a22279a );
 a22289a <=( A267  and  A266 );
 a22290a <=( (not A265)  and  a22289a );
 a22294a <=( A302  and  (not A300) );
 a22295a <=( A268  and  a22294a );
 a22296a <=( a22295a  and  a22290a );
 a22299a <=( (not A169)  and  A170 );
 a22303a <=( A203  and  (not A201) );
 a22304a <=( A168  and  a22303a );
 a22305a <=( a22304a  and  a22299a );
 a22309a <=( A267  and  A266 );
 a22310a <=( (not A265)  and  a22309a );
 a22314a <=( A299  and  A298 );
 a22315a <=( A268  and  a22314a );
 a22316a <=( a22315a  and  a22310a );
 a22319a <=( (not A169)  and  A170 );
 a22323a <=( A203  and  (not A201) );
 a22324a <=( A168  and  a22323a );
 a22325a <=( a22324a  and  a22319a );
 a22329a <=( A267  and  A266 );
 a22330a <=( (not A265)  and  a22329a );
 a22334a <=( (not A299)  and  (not A298) );
 a22335a <=( A268  and  a22334a );
 a22336a <=( a22335a  and  a22330a );
 a22339a <=( (not A169)  and  A170 );
 a22343a <=( A203  and  (not A201) );
 a22344a <=( A168  and  a22343a );
 a22345a <=( a22344a  and  a22339a );
 a22349a <=( A267  and  A266 );
 a22350a <=( (not A265)  and  a22349a );
 a22354a <=( A301  and  (not A300) );
 a22355a <=( A269  and  a22354a );
 a22356a <=( a22355a  and  a22350a );
 a22359a <=( (not A169)  and  A170 );
 a22363a <=( A203  and  (not A201) );
 a22364a <=( A168  and  a22363a );
 a22365a <=( a22364a  and  a22359a );
 a22369a <=( A267  and  A266 );
 a22370a <=( (not A265)  and  a22369a );
 a22374a <=( A302  and  (not A300) );
 a22375a <=( A269  and  a22374a );
 a22376a <=( a22375a  and  a22370a );
 a22379a <=( (not A169)  and  A170 );
 a22383a <=( A203  and  (not A201) );
 a22384a <=( A168  and  a22383a );
 a22385a <=( a22384a  and  a22379a );
 a22389a <=( A267  and  A266 );
 a22390a <=( (not A265)  and  a22389a );
 a22394a <=( A299  and  A298 );
 a22395a <=( A269  and  a22394a );
 a22396a <=( a22395a  and  a22390a );
 a22399a <=( (not A169)  and  A170 );
 a22403a <=( A203  and  (not A201) );
 a22404a <=( A168  and  a22403a );
 a22405a <=( a22404a  and  a22399a );
 a22409a <=( A267  and  A266 );
 a22410a <=( (not A265)  and  a22409a );
 a22414a <=( (not A299)  and  (not A298) );
 a22415a <=( A269  and  a22414a );
 a22416a <=( a22415a  and  a22410a );
 a22419a <=( (not A169)  and  A170 );
 a22423a <=( A203  and  (not A201) );
 a22424a <=( A168  and  a22423a );
 a22425a <=( a22424a  and  a22419a );
 a22429a <=( A267  and  (not A266) );
 a22430a <=( A265  and  a22429a );
 a22434a <=( A301  and  (not A300) );
 a22435a <=( A268  and  a22434a );
 a22436a <=( a22435a  and  a22430a );
 a22439a <=( (not A169)  and  A170 );
 a22443a <=( A203  and  (not A201) );
 a22444a <=( A168  and  a22443a );
 a22445a <=( a22444a  and  a22439a );
 a22449a <=( A267  and  (not A266) );
 a22450a <=( A265  and  a22449a );
 a22454a <=( A302  and  (not A300) );
 a22455a <=( A268  and  a22454a );
 a22456a <=( a22455a  and  a22450a );
 a22459a <=( (not A169)  and  A170 );
 a22463a <=( A203  and  (not A201) );
 a22464a <=( A168  and  a22463a );
 a22465a <=( a22464a  and  a22459a );
 a22469a <=( A267  and  (not A266) );
 a22470a <=( A265  and  a22469a );
 a22474a <=( A299  and  A298 );
 a22475a <=( A268  and  a22474a );
 a22476a <=( a22475a  and  a22470a );
 a22479a <=( (not A169)  and  A170 );
 a22483a <=( A203  and  (not A201) );
 a22484a <=( A168  and  a22483a );
 a22485a <=( a22484a  and  a22479a );
 a22489a <=( A267  and  (not A266) );
 a22490a <=( A265  and  a22489a );
 a22494a <=( (not A299)  and  (not A298) );
 a22495a <=( A268  and  a22494a );
 a22496a <=( a22495a  and  a22490a );
 a22499a <=( (not A169)  and  A170 );
 a22503a <=( A203  and  (not A201) );
 a22504a <=( A168  and  a22503a );
 a22505a <=( a22504a  and  a22499a );
 a22509a <=( A267  and  (not A266) );
 a22510a <=( A265  and  a22509a );
 a22514a <=( A301  and  (not A300) );
 a22515a <=( A269  and  a22514a );
 a22516a <=( a22515a  and  a22510a );
 a22519a <=( (not A169)  and  A170 );
 a22523a <=( A203  and  (not A201) );
 a22524a <=( A168  and  a22523a );
 a22525a <=( a22524a  and  a22519a );
 a22529a <=( A267  and  (not A266) );
 a22530a <=( A265  and  a22529a );
 a22534a <=( A302  and  (not A300) );
 a22535a <=( A269  and  a22534a );
 a22536a <=( a22535a  and  a22530a );
 a22539a <=( (not A169)  and  A170 );
 a22543a <=( A203  and  (not A201) );
 a22544a <=( A168  and  a22543a );
 a22545a <=( a22544a  and  a22539a );
 a22549a <=( A267  and  (not A266) );
 a22550a <=( A265  and  a22549a );
 a22554a <=( A299  and  A298 );
 a22555a <=( A269  and  a22554a );
 a22556a <=( a22555a  and  a22550a );
 a22559a <=( (not A169)  and  A170 );
 a22563a <=( A203  and  (not A201) );
 a22564a <=( A168  and  a22563a );
 a22565a <=( a22564a  and  a22559a );
 a22569a <=( A267  and  (not A266) );
 a22570a <=( A265  and  a22569a );
 a22574a <=( (not A299)  and  (not A298) );
 a22575a <=( A269  and  a22574a );
 a22576a <=( a22575a  and  a22570a );
 a22579a <=( (not A169)  and  A170 );
 a22583a <=( A200  and  A199 );
 a22584a <=( A168  and  a22583a );
 a22585a <=( a22584a  and  a22579a );
 a22589a <=( A267  and  A266 );
 a22590a <=( (not A265)  and  a22589a );
 a22594a <=( A301  and  (not A300) );
 a22595a <=( A268  and  a22594a );
 a22596a <=( a22595a  and  a22590a );
 a22599a <=( (not A169)  and  A170 );
 a22603a <=( A200  and  A199 );
 a22604a <=( A168  and  a22603a );
 a22605a <=( a22604a  and  a22599a );
 a22609a <=( A267  and  A266 );
 a22610a <=( (not A265)  and  a22609a );
 a22614a <=( A302  and  (not A300) );
 a22615a <=( A268  and  a22614a );
 a22616a <=( a22615a  and  a22610a );
 a22619a <=( (not A169)  and  A170 );
 a22623a <=( A200  and  A199 );
 a22624a <=( A168  and  a22623a );
 a22625a <=( a22624a  and  a22619a );
 a22629a <=( A267  and  A266 );
 a22630a <=( (not A265)  and  a22629a );
 a22634a <=( A299  and  A298 );
 a22635a <=( A268  and  a22634a );
 a22636a <=( a22635a  and  a22630a );
 a22639a <=( (not A169)  and  A170 );
 a22643a <=( A200  and  A199 );
 a22644a <=( A168  and  a22643a );
 a22645a <=( a22644a  and  a22639a );
 a22649a <=( A267  and  A266 );
 a22650a <=( (not A265)  and  a22649a );
 a22654a <=( (not A299)  and  (not A298) );
 a22655a <=( A268  and  a22654a );
 a22656a <=( a22655a  and  a22650a );
 a22659a <=( (not A169)  and  A170 );
 a22663a <=( A200  and  A199 );
 a22664a <=( A168  and  a22663a );
 a22665a <=( a22664a  and  a22659a );
 a22669a <=( A267  and  A266 );
 a22670a <=( (not A265)  and  a22669a );
 a22674a <=( A301  and  (not A300) );
 a22675a <=( A269  and  a22674a );
 a22676a <=( a22675a  and  a22670a );
 a22679a <=( (not A169)  and  A170 );
 a22683a <=( A200  and  A199 );
 a22684a <=( A168  and  a22683a );
 a22685a <=( a22684a  and  a22679a );
 a22689a <=( A267  and  A266 );
 a22690a <=( (not A265)  and  a22689a );
 a22694a <=( A302  and  (not A300) );
 a22695a <=( A269  and  a22694a );
 a22696a <=( a22695a  and  a22690a );
 a22699a <=( (not A169)  and  A170 );
 a22703a <=( A200  and  A199 );
 a22704a <=( A168  and  a22703a );
 a22705a <=( a22704a  and  a22699a );
 a22709a <=( A267  and  A266 );
 a22710a <=( (not A265)  and  a22709a );
 a22714a <=( A299  and  A298 );
 a22715a <=( A269  and  a22714a );
 a22716a <=( a22715a  and  a22710a );
 a22719a <=( (not A169)  and  A170 );
 a22723a <=( A200  and  A199 );
 a22724a <=( A168  and  a22723a );
 a22725a <=( a22724a  and  a22719a );
 a22729a <=( A267  and  A266 );
 a22730a <=( (not A265)  and  a22729a );
 a22734a <=( (not A299)  and  (not A298) );
 a22735a <=( A269  and  a22734a );
 a22736a <=( a22735a  and  a22730a );
 a22739a <=( (not A169)  and  A170 );
 a22743a <=( A200  and  A199 );
 a22744a <=( A168  and  a22743a );
 a22745a <=( a22744a  and  a22739a );
 a22749a <=( A267  and  (not A266) );
 a22750a <=( A265  and  a22749a );
 a22754a <=( A301  and  (not A300) );
 a22755a <=( A268  and  a22754a );
 a22756a <=( a22755a  and  a22750a );
 a22759a <=( (not A169)  and  A170 );
 a22763a <=( A200  and  A199 );
 a22764a <=( A168  and  a22763a );
 a22765a <=( a22764a  and  a22759a );
 a22769a <=( A267  and  (not A266) );
 a22770a <=( A265  and  a22769a );
 a22774a <=( A302  and  (not A300) );
 a22775a <=( A268  and  a22774a );
 a22776a <=( a22775a  and  a22770a );
 a22779a <=( (not A169)  and  A170 );
 a22783a <=( A200  and  A199 );
 a22784a <=( A168  and  a22783a );
 a22785a <=( a22784a  and  a22779a );
 a22789a <=( A267  and  (not A266) );
 a22790a <=( A265  and  a22789a );
 a22794a <=( A299  and  A298 );
 a22795a <=( A268  and  a22794a );
 a22796a <=( a22795a  and  a22790a );
 a22799a <=( (not A169)  and  A170 );
 a22803a <=( A200  and  A199 );
 a22804a <=( A168  and  a22803a );
 a22805a <=( a22804a  and  a22799a );
 a22809a <=( A267  and  (not A266) );
 a22810a <=( A265  and  a22809a );
 a22814a <=( (not A299)  and  (not A298) );
 a22815a <=( A268  and  a22814a );
 a22816a <=( a22815a  and  a22810a );
 a22819a <=( (not A169)  and  A170 );
 a22823a <=( A200  and  A199 );
 a22824a <=( A168  and  a22823a );
 a22825a <=( a22824a  and  a22819a );
 a22829a <=( A267  and  (not A266) );
 a22830a <=( A265  and  a22829a );
 a22834a <=( A301  and  (not A300) );
 a22835a <=( A269  and  a22834a );
 a22836a <=( a22835a  and  a22830a );
 a22839a <=( (not A169)  and  A170 );
 a22843a <=( A200  and  A199 );
 a22844a <=( A168  and  a22843a );
 a22845a <=( a22844a  and  a22839a );
 a22849a <=( A267  and  (not A266) );
 a22850a <=( A265  and  a22849a );
 a22854a <=( A302  and  (not A300) );
 a22855a <=( A269  and  a22854a );
 a22856a <=( a22855a  and  a22850a );
 a22859a <=( (not A169)  and  A170 );
 a22863a <=( A200  and  A199 );
 a22864a <=( A168  and  a22863a );
 a22865a <=( a22864a  and  a22859a );
 a22869a <=( A267  and  (not A266) );
 a22870a <=( A265  and  a22869a );
 a22874a <=( A299  and  A298 );
 a22875a <=( A269  and  a22874a );
 a22876a <=( a22875a  and  a22870a );
 a22879a <=( (not A169)  and  A170 );
 a22883a <=( A200  and  A199 );
 a22884a <=( A168  and  a22883a );
 a22885a <=( a22884a  and  a22879a );
 a22889a <=( A267  and  (not A266) );
 a22890a <=( A265  and  a22889a );
 a22894a <=( (not A299)  and  (not A298) );
 a22895a <=( A269  and  a22894a );
 a22896a <=( a22895a  and  a22890a );
 a22899a <=( (not A169)  and  A170 );
 a22903a <=( (not A200)  and  (not A199) );
 a22904a <=( A168  and  a22903a );
 a22905a <=( a22904a  and  a22899a );
 a22909a <=( A267  and  A266 );
 a22910a <=( (not A265)  and  a22909a );
 a22914a <=( A301  and  (not A300) );
 a22915a <=( A268  and  a22914a );
 a22916a <=( a22915a  and  a22910a );
 a22919a <=( (not A169)  and  A170 );
 a22923a <=( (not A200)  and  (not A199) );
 a22924a <=( A168  and  a22923a );
 a22925a <=( a22924a  and  a22919a );
 a22929a <=( A267  and  A266 );
 a22930a <=( (not A265)  and  a22929a );
 a22934a <=( A302  and  (not A300) );
 a22935a <=( A268  and  a22934a );
 a22936a <=( a22935a  and  a22930a );
 a22939a <=( (not A169)  and  A170 );
 a22943a <=( (not A200)  and  (not A199) );
 a22944a <=( A168  and  a22943a );
 a22945a <=( a22944a  and  a22939a );
 a22949a <=( A267  and  A266 );
 a22950a <=( (not A265)  and  a22949a );
 a22954a <=( A299  and  A298 );
 a22955a <=( A268  and  a22954a );
 a22956a <=( a22955a  and  a22950a );
 a22959a <=( (not A169)  and  A170 );
 a22963a <=( (not A200)  and  (not A199) );
 a22964a <=( A168  and  a22963a );
 a22965a <=( a22964a  and  a22959a );
 a22969a <=( A267  and  A266 );
 a22970a <=( (not A265)  and  a22969a );
 a22974a <=( (not A299)  and  (not A298) );
 a22975a <=( A268  and  a22974a );
 a22976a <=( a22975a  and  a22970a );
 a22979a <=( (not A169)  and  A170 );
 a22983a <=( (not A200)  and  (not A199) );
 a22984a <=( A168  and  a22983a );
 a22985a <=( a22984a  and  a22979a );
 a22989a <=( A267  and  A266 );
 a22990a <=( (not A265)  and  a22989a );
 a22994a <=( A301  and  (not A300) );
 a22995a <=( A269  and  a22994a );
 a22996a <=( a22995a  and  a22990a );
 a22999a <=( (not A169)  and  A170 );
 a23003a <=( (not A200)  and  (not A199) );
 a23004a <=( A168  and  a23003a );
 a23005a <=( a23004a  and  a22999a );
 a23009a <=( A267  and  A266 );
 a23010a <=( (not A265)  and  a23009a );
 a23014a <=( A302  and  (not A300) );
 a23015a <=( A269  and  a23014a );
 a23016a <=( a23015a  and  a23010a );
 a23019a <=( (not A169)  and  A170 );
 a23023a <=( (not A200)  and  (not A199) );
 a23024a <=( A168  and  a23023a );
 a23025a <=( a23024a  and  a23019a );
 a23029a <=( A267  and  A266 );
 a23030a <=( (not A265)  and  a23029a );
 a23034a <=( A299  and  A298 );
 a23035a <=( A269  and  a23034a );
 a23036a <=( a23035a  and  a23030a );
 a23039a <=( (not A169)  and  A170 );
 a23043a <=( (not A200)  and  (not A199) );
 a23044a <=( A168  and  a23043a );
 a23045a <=( a23044a  and  a23039a );
 a23049a <=( A267  and  A266 );
 a23050a <=( (not A265)  and  a23049a );
 a23054a <=( (not A299)  and  (not A298) );
 a23055a <=( A269  and  a23054a );
 a23056a <=( a23055a  and  a23050a );
 a23059a <=( (not A169)  and  A170 );
 a23063a <=( (not A200)  and  (not A199) );
 a23064a <=( A168  and  a23063a );
 a23065a <=( a23064a  and  a23059a );
 a23069a <=( A267  and  (not A266) );
 a23070a <=( A265  and  a23069a );
 a23074a <=( A301  and  (not A300) );
 a23075a <=( A268  and  a23074a );
 a23076a <=( a23075a  and  a23070a );
 a23079a <=( (not A169)  and  A170 );
 a23083a <=( (not A200)  and  (not A199) );
 a23084a <=( A168  and  a23083a );
 a23085a <=( a23084a  and  a23079a );
 a23089a <=( A267  and  (not A266) );
 a23090a <=( A265  and  a23089a );
 a23094a <=( A302  and  (not A300) );
 a23095a <=( A268  and  a23094a );
 a23096a <=( a23095a  and  a23090a );
 a23099a <=( (not A169)  and  A170 );
 a23103a <=( (not A200)  and  (not A199) );
 a23104a <=( A168  and  a23103a );
 a23105a <=( a23104a  and  a23099a );
 a23109a <=( A267  and  (not A266) );
 a23110a <=( A265  and  a23109a );
 a23114a <=( A299  and  A298 );
 a23115a <=( A268  and  a23114a );
 a23116a <=( a23115a  and  a23110a );
 a23119a <=( (not A169)  and  A170 );
 a23123a <=( (not A200)  and  (not A199) );
 a23124a <=( A168  and  a23123a );
 a23125a <=( a23124a  and  a23119a );
 a23129a <=( A267  and  (not A266) );
 a23130a <=( A265  and  a23129a );
 a23134a <=( (not A299)  and  (not A298) );
 a23135a <=( A268  and  a23134a );
 a23136a <=( a23135a  and  a23130a );
 a23139a <=( (not A169)  and  A170 );
 a23143a <=( (not A200)  and  (not A199) );
 a23144a <=( A168  and  a23143a );
 a23145a <=( a23144a  and  a23139a );
 a23149a <=( A267  and  (not A266) );
 a23150a <=( A265  and  a23149a );
 a23154a <=( A301  and  (not A300) );
 a23155a <=( A269  and  a23154a );
 a23156a <=( a23155a  and  a23150a );
 a23159a <=( (not A169)  and  A170 );
 a23163a <=( (not A200)  and  (not A199) );
 a23164a <=( A168  and  a23163a );
 a23165a <=( a23164a  and  a23159a );
 a23169a <=( A267  and  (not A266) );
 a23170a <=( A265  and  a23169a );
 a23174a <=( A302  and  (not A300) );
 a23175a <=( A269  and  a23174a );
 a23176a <=( a23175a  and  a23170a );
 a23179a <=( (not A169)  and  A170 );
 a23183a <=( (not A200)  and  (not A199) );
 a23184a <=( A168  and  a23183a );
 a23185a <=( a23184a  and  a23179a );
 a23189a <=( A267  and  (not A266) );
 a23190a <=( A265  and  a23189a );
 a23194a <=( A299  and  A298 );
 a23195a <=( A269  and  a23194a );
 a23196a <=( a23195a  and  a23190a );
 a23199a <=( (not A169)  and  A170 );
 a23203a <=( (not A200)  and  (not A199) );
 a23204a <=( A168  and  a23203a );
 a23205a <=( a23204a  and  a23199a );
 a23209a <=( A267  and  (not A266) );
 a23210a <=( A265  and  a23209a );
 a23214a <=( (not A299)  and  (not A298) );
 a23215a <=( A269  and  a23214a );
 a23216a <=( a23215a  and  a23210a );
 a23220a <=( A201  and  A166 );
 a23221a <=( A167  and  a23220a );
 a23225a <=( (not A265)  and  (not A203) );
 a23226a <=( (not A202)  and  a23225a );
 a23227a <=( a23226a  and  a23221a );
 a23231a <=( A268  and  A267 );
 a23232a <=( A266  and  a23231a );
 a23236a <=( (not A302)  and  (not A301) );
 a23237a <=( A300  and  a23236a );
 a23238a <=( a23237a  and  a23232a );
 a23242a <=( A201  and  A166 );
 a23243a <=( A167  and  a23242a );
 a23247a <=( (not A265)  and  (not A203) );
 a23248a <=( (not A202)  and  a23247a );
 a23249a <=( a23248a  and  a23243a );
 a23253a <=( A269  and  A267 );
 a23254a <=( A266  and  a23253a );
 a23258a <=( (not A302)  and  (not A301) );
 a23259a <=( A300  and  a23258a );
 a23260a <=( a23259a  and  a23254a );
 a23264a <=( A201  and  A166 );
 a23265a <=( A167  and  a23264a );
 a23269a <=( (not A265)  and  (not A203) );
 a23270a <=( (not A202)  and  a23269a );
 a23271a <=( a23270a  and  a23265a );
 a23275a <=( (not A268)  and  (not A267) );
 a23276a <=( A266  and  a23275a );
 a23280a <=( A301  and  (not A300) );
 a23281a <=( (not A269)  and  a23280a );
 a23282a <=( a23281a  and  a23276a );
 a23286a <=( A201  and  A166 );
 a23287a <=( A167  and  a23286a );
 a23291a <=( (not A265)  and  (not A203) );
 a23292a <=( (not A202)  and  a23291a );
 a23293a <=( a23292a  and  a23287a );
 a23297a <=( (not A268)  and  (not A267) );
 a23298a <=( A266  and  a23297a );
 a23302a <=( A302  and  (not A300) );
 a23303a <=( (not A269)  and  a23302a );
 a23304a <=( a23303a  and  a23298a );
 a23308a <=( A201  and  A166 );
 a23309a <=( A167  and  a23308a );
 a23313a <=( (not A265)  and  (not A203) );
 a23314a <=( (not A202)  and  a23313a );
 a23315a <=( a23314a  and  a23309a );
 a23319a <=( (not A268)  and  (not A267) );
 a23320a <=( A266  and  a23319a );
 a23324a <=( A299  and  A298 );
 a23325a <=( (not A269)  and  a23324a );
 a23326a <=( a23325a  and  a23320a );
 a23330a <=( A201  and  A166 );
 a23331a <=( A167  and  a23330a );
 a23335a <=( (not A265)  and  (not A203) );
 a23336a <=( (not A202)  and  a23335a );
 a23337a <=( a23336a  and  a23331a );
 a23341a <=( (not A268)  and  (not A267) );
 a23342a <=( A266  and  a23341a );
 a23346a <=( (not A299)  and  (not A298) );
 a23347a <=( (not A269)  and  a23346a );
 a23348a <=( a23347a  and  a23342a );
 a23352a <=( A201  and  A166 );
 a23353a <=( A167  and  a23352a );
 a23357a <=( A265  and  (not A203) );
 a23358a <=( (not A202)  and  a23357a );
 a23359a <=( a23358a  and  a23353a );
 a23363a <=( A268  and  A267 );
 a23364a <=( (not A266)  and  a23363a );
 a23368a <=( (not A302)  and  (not A301) );
 a23369a <=( A300  and  a23368a );
 a23370a <=( a23369a  and  a23364a );
 a23374a <=( A201  and  A166 );
 a23375a <=( A167  and  a23374a );
 a23379a <=( A265  and  (not A203) );
 a23380a <=( (not A202)  and  a23379a );
 a23381a <=( a23380a  and  a23375a );
 a23385a <=( A269  and  A267 );
 a23386a <=( (not A266)  and  a23385a );
 a23390a <=( (not A302)  and  (not A301) );
 a23391a <=( A300  and  a23390a );
 a23392a <=( a23391a  and  a23386a );
 a23396a <=( A201  and  A166 );
 a23397a <=( A167  and  a23396a );
 a23401a <=( A265  and  (not A203) );
 a23402a <=( (not A202)  and  a23401a );
 a23403a <=( a23402a  and  a23397a );
 a23407a <=( (not A268)  and  (not A267) );
 a23408a <=( (not A266)  and  a23407a );
 a23412a <=( A301  and  (not A300) );
 a23413a <=( (not A269)  and  a23412a );
 a23414a <=( a23413a  and  a23408a );
 a23418a <=( A201  and  A166 );
 a23419a <=( A167  and  a23418a );
 a23423a <=( A265  and  (not A203) );
 a23424a <=( (not A202)  and  a23423a );
 a23425a <=( a23424a  and  a23419a );
 a23429a <=( (not A268)  and  (not A267) );
 a23430a <=( (not A266)  and  a23429a );
 a23434a <=( A302  and  (not A300) );
 a23435a <=( (not A269)  and  a23434a );
 a23436a <=( a23435a  and  a23430a );
 a23440a <=( A201  and  A166 );
 a23441a <=( A167  and  a23440a );
 a23445a <=( A265  and  (not A203) );
 a23446a <=( (not A202)  and  a23445a );
 a23447a <=( a23446a  and  a23441a );
 a23451a <=( (not A268)  and  (not A267) );
 a23452a <=( (not A266)  and  a23451a );
 a23456a <=( A299  and  A298 );
 a23457a <=( (not A269)  and  a23456a );
 a23458a <=( a23457a  and  a23452a );
 a23462a <=( A201  and  A166 );
 a23463a <=( A167  and  a23462a );
 a23467a <=( A265  and  (not A203) );
 a23468a <=( (not A202)  and  a23467a );
 a23469a <=( a23468a  and  a23463a );
 a23473a <=( (not A268)  and  (not A267) );
 a23474a <=( (not A266)  and  a23473a );
 a23478a <=( (not A299)  and  (not A298) );
 a23479a <=( (not A269)  and  a23478a );
 a23480a <=( a23479a  and  a23474a );
 a23484a <=( (not A201)  and  A166 );
 a23485a <=( A167  and  a23484a );
 a23489a <=( A266  and  (not A265) );
 a23490a <=( A202  and  a23489a );
 a23491a <=( a23490a  and  a23485a );
 a23495a <=( (not A269)  and  (not A268) );
 a23496a <=( (not A267)  and  a23495a );
 a23500a <=( (not A302)  and  (not A301) );
 a23501a <=( A300  and  a23500a );
 a23502a <=( a23501a  and  a23496a );
 a23506a <=( (not A201)  and  A166 );
 a23507a <=( A167  and  a23506a );
 a23511a <=( (not A266)  and  A265 );
 a23512a <=( A202  and  a23511a );
 a23513a <=( a23512a  and  a23507a );
 a23517a <=( (not A269)  and  (not A268) );
 a23518a <=( (not A267)  and  a23517a );
 a23522a <=( (not A302)  and  (not A301) );
 a23523a <=( A300  and  a23522a );
 a23524a <=( a23523a  and  a23518a );
 a23528a <=( (not A201)  and  A166 );
 a23529a <=( A167  and  a23528a );
 a23533a <=( A266  and  (not A265) );
 a23534a <=( A203  and  a23533a );
 a23535a <=( a23534a  and  a23529a );
 a23539a <=( (not A269)  and  (not A268) );
 a23540a <=( (not A267)  and  a23539a );
 a23544a <=( (not A302)  and  (not A301) );
 a23545a <=( A300  and  a23544a );
 a23546a <=( a23545a  and  a23540a );
 a23550a <=( (not A201)  and  A166 );
 a23551a <=( A167  and  a23550a );
 a23555a <=( (not A266)  and  A265 );
 a23556a <=( A203  and  a23555a );
 a23557a <=( a23556a  and  a23551a );
 a23561a <=( (not A269)  and  (not A268) );
 a23562a <=( (not A267)  and  a23561a );
 a23566a <=( (not A302)  and  (not A301) );
 a23567a <=( A300  and  a23566a );
 a23568a <=( a23567a  and  a23562a );
 a23572a <=( A199  and  A166 );
 a23573a <=( A167  and  a23572a );
 a23577a <=( A266  and  (not A265) );
 a23578a <=( A200  and  a23577a );
 a23579a <=( a23578a  and  a23573a );
 a23583a <=( (not A269)  and  (not A268) );
 a23584a <=( (not A267)  and  a23583a );
 a23588a <=( (not A302)  and  (not A301) );
 a23589a <=( A300  and  a23588a );
 a23590a <=( a23589a  and  a23584a );
 a23594a <=( A199  and  A166 );
 a23595a <=( A167  and  a23594a );
 a23599a <=( (not A266)  and  A265 );
 a23600a <=( A200  and  a23599a );
 a23601a <=( a23600a  and  a23595a );
 a23605a <=( (not A269)  and  (not A268) );
 a23606a <=( (not A267)  and  a23605a );
 a23610a <=( (not A302)  and  (not A301) );
 a23611a <=( A300  and  a23610a );
 a23612a <=( a23611a  and  a23606a );
 a23616a <=( (not A199)  and  A166 );
 a23617a <=( A167  and  a23616a );
 a23621a <=( A202  and  A201 );
 a23622a <=( A200  and  a23621a );
 a23623a <=( a23622a  and  a23617a );
 a23627a <=( A298  and  A268 );
 a23628a <=( (not A267)  and  a23627a );
 a23632a <=( A301  and  A300 );
 a23633a <=( (not A299)  and  a23632a );
 a23634a <=( a23633a  and  a23628a );
 a23638a <=( (not A199)  and  A166 );
 a23639a <=( A167  and  a23638a );
 a23643a <=( A202  and  A201 );
 a23644a <=( A200  and  a23643a );
 a23645a <=( a23644a  and  a23639a );
 a23649a <=( A298  and  A268 );
 a23650a <=( (not A267)  and  a23649a );
 a23654a <=( A302  and  A300 );
 a23655a <=( (not A299)  and  a23654a );
 a23656a <=( a23655a  and  a23650a );
 a23660a <=( (not A199)  and  A166 );
 a23661a <=( A167  and  a23660a );
 a23665a <=( A202  and  A201 );
 a23666a <=( A200  and  a23665a );
 a23667a <=( a23666a  and  a23661a );
 a23671a <=( (not A298)  and  A268 );
 a23672a <=( (not A267)  and  a23671a );
 a23676a <=( A301  and  A300 );
 a23677a <=( A299  and  a23676a );
 a23678a <=( a23677a  and  a23672a );
 a23682a <=( (not A199)  and  A166 );
 a23683a <=( A167  and  a23682a );
 a23687a <=( A202  and  A201 );
 a23688a <=( A200  and  a23687a );
 a23689a <=( a23688a  and  a23683a );
 a23693a <=( (not A298)  and  A268 );
 a23694a <=( (not A267)  and  a23693a );
 a23698a <=( A302  and  A300 );
 a23699a <=( A299  and  a23698a );
 a23700a <=( a23699a  and  a23694a );
 a23704a <=( (not A199)  and  A166 );
 a23705a <=( A167  and  a23704a );
 a23709a <=( A202  and  A201 );
 a23710a <=( A200  and  a23709a );
 a23711a <=( a23710a  and  a23705a );
 a23715a <=( A298  and  A269 );
 a23716a <=( (not A267)  and  a23715a );
 a23720a <=( A301  and  A300 );
 a23721a <=( (not A299)  and  a23720a );
 a23722a <=( a23721a  and  a23716a );
 a23726a <=( (not A199)  and  A166 );
 a23727a <=( A167  and  a23726a );
 a23731a <=( A202  and  A201 );
 a23732a <=( A200  and  a23731a );
 a23733a <=( a23732a  and  a23727a );
 a23737a <=( A298  and  A269 );
 a23738a <=( (not A267)  and  a23737a );
 a23742a <=( A302  and  A300 );
 a23743a <=( (not A299)  and  a23742a );
 a23744a <=( a23743a  and  a23738a );
 a23748a <=( (not A199)  and  A166 );
 a23749a <=( A167  and  a23748a );
 a23753a <=( A202  and  A201 );
 a23754a <=( A200  and  a23753a );
 a23755a <=( a23754a  and  a23749a );
 a23759a <=( (not A298)  and  A269 );
 a23760a <=( (not A267)  and  a23759a );
 a23764a <=( A301  and  A300 );
 a23765a <=( A299  and  a23764a );
 a23766a <=( a23765a  and  a23760a );
 a23770a <=( (not A199)  and  A166 );
 a23771a <=( A167  and  a23770a );
 a23775a <=( A202  and  A201 );
 a23776a <=( A200  and  a23775a );
 a23777a <=( a23776a  and  a23771a );
 a23781a <=( (not A298)  and  A269 );
 a23782a <=( (not A267)  and  a23781a );
 a23786a <=( A302  and  A300 );
 a23787a <=( A299  and  a23786a );
 a23788a <=( a23787a  and  a23782a );
 a23792a <=( (not A199)  and  A166 );
 a23793a <=( A167  and  a23792a );
 a23797a <=( A202  and  A201 );
 a23798a <=( A200  and  a23797a );
 a23799a <=( a23798a  and  a23793a );
 a23803a <=( A298  and  A266 );
 a23804a <=( A265  and  a23803a );
 a23808a <=( A301  and  A300 );
 a23809a <=( (not A299)  and  a23808a );
 a23810a <=( a23809a  and  a23804a );
 a23814a <=( (not A199)  and  A166 );
 a23815a <=( A167  and  a23814a );
 a23819a <=( A202  and  A201 );
 a23820a <=( A200  and  a23819a );
 a23821a <=( a23820a  and  a23815a );
 a23825a <=( A298  and  A266 );
 a23826a <=( A265  and  a23825a );
 a23830a <=( A302  and  A300 );
 a23831a <=( (not A299)  and  a23830a );
 a23832a <=( a23831a  and  a23826a );
 a23836a <=( (not A199)  and  A166 );
 a23837a <=( A167  and  a23836a );
 a23841a <=( A202  and  A201 );
 a23842a <=( A200  and  a23841a );
 a23843a <=( a23842a  and  a23837a );
 a23847a <=( (not A298)  and  A266 );
 a23848a <=( A265  and  a23847a );
 a23852a <=( A301  and  A300 );
 a23853a <=( A299  and  a23852a );
 a23854a <=( a23853a  and  a23848a );
 a23858a <=( (not A199)  and  A166 );
 a23859a <=( A167  and  a23858a );
 a23863a <=( A202  and  A201 );
 a23864a <=( A200  and  a23863a );
 a23865a <=( a23864a  and  a23859a );
 a23869a <=( (not A298)  and  A266 );
 a23870a <=( A265  and  a23869a );
 a23874a <=( A302  and  A300 );
 a23875a <=( A299  and  a23874a );
 a23876a <=( a23875a  and  a23870a );
 a23880a <=( (not A199)  and  A166 );
 a23881a <=( A167  and  a23880a );
 a23885a <=( A202  and  A201 );
 a23886a <=( A200  and  a23885a );
 a23887a <=( a23886a  and  a23881a );
 a23891a <=( A298  and  (not A266) );
 a23892a <=( (not A265)  and  a23891a );
 a23896a <=( A301  and  A300 );
 a23897a <=( (not A299)  and  a23896a );
 a23898a <=( a23897a  and  a23892a );
 a23902a <=( (not A199)  and  A166 );
 a23903a <=( A167  and  a23902a );
 a23907a <=( A202  and  A201 );
 a23908a <=( A200  and  a23907a );
 a23909a <=( a23908a  and  a23903a );
 a23913a <=( A298  and  (not A266) );
 a23914a <=( (not A265)  and  a23913a );
 a23918a <=( A302  and  A300 );
 a23919a <=( (not A299)  and  a23918a );
 a23920a <=( a23919a  and  a23914a );
 a23924a <=( (not A199)  and  A166 );
 a23925a <=( A167  and  a23924a );
 a23929a <=( A202  and  A201 );
 a23930a <=( A200  and  a23929a );
 a23931a <=( a23930a  and  a23925a );
 a23935a <=( (not A298)  and  (not A266) );
 a23936a <=( (not A265)  and  a23935a );
 a23940a <=( A301  and  A300 );
 a23941a <=( A299  and  a23940a );
 a23942a <=( a23941a  and  a23936a );
 a23946a <=( (not A199)  and  A166 );
 a23947a <=( A167  and  a23946a );
 a23951a <=( A202  and  A201 );
 a23952a <=( A200  and  a23951a );
 a23953a <=( a23952a  and  a23947a );
 a23957a <=( (not A298)  and  (not A266) );
 a23958a <=( (not A265)  and  a23957a );
 a23962a <=( A302  and  A300 );
 a23963a <=( A299  and  a23962a );
 a23964a <=( a23963a  and  a23958a );
 a23968a <=( (not A199)  and  A166 );
 a23969a <=( A167  and  a23968a );
 a23973a <=( A203  and  A201 );
 a23974a <=( A200  and  a23973a );
 a23975a <=( a23974a  and  a23969a );
 a23979a <=( A298  and  A268 );
 a23980a <=( (not A267)  and  a23979a );
 a23984a <=( A301  and  A300 );
 a23985a <=( (not A299)  and  a23984a );
 a23986a <=( a23985a  and  a23980a );
 a23990a <=( (not A199)  and  A166 );
 a23991a <=( A167  and  a23990a );
 a23995a <=( A203  and  A201 );
 a23996a <=( A200  and  a23995a );
 a23997a <=( a23996a  and  a23991a );
 a24001a <=( A298  and  A268 );
 a24002a <=( (not A267)  and  a24001a );
 a24006a <=( A302  and  A300 );
 a24007a <=( (not A299)  and  a24006a );
 a24008a <=( a24007a  and  a24002a );
 a24012a <=( (not A199)  and  A166 );
 a24013a <=( A167  and  a24012a );
 a24017a <=( A203  and  A201 );
 a24018a <=( A200  and  a24017a );
 a24019a <=( a24018a  and  a24013a );
 a24023a <=( (not A298)  and  A268 );
 a24024a <=( (not A267)  and  a24023a );
 a24028a <=( A301  and  A300 );
 a24029a <=( A299  and  a24028a );
 a24030a <=( a24029a  and  a24024a );
 a24034a <=( (not A199)  and  A166 );
 a24035a <=( A167  and  a24034a );
 a24039a <=( A203  and  A201 );
 a24040a <=( A200  and  a24039a );
 a24041a <=( a24040a  and  a24035a );
 a24045a <=( (not A298)  and  A268 );
 a24046a <=( (not A267)  and  a24045a );
 a24050a <=( A302  and  A300 );
 a24051a <=( A299  and  a24050a );
 a24052a <=( a24051a  and  a24046a );
 a24056a <=( (not A199)  and  A166 );
 a24057a <=( A167  and  a24056a );
 a24061a <=( A203  and  A201 );
 a24062a <=( A200  and  a24061a );
 a24063a <=( a24062a  and  a24057a );
 a24067a <=( A298  and  A269 );
 a24068a <=( (not A267)  and  a24067a );
 a24072a <=( A301  and  A300 );
 a24073a <=( (not A299)  and  a24072a );
 a24074a <=( a24073a  and  a24068a );
 a24078a <=( (not A199)  and  A166 );
 a24079a <=( A167  and  a24078a );
 a24083a <=( A203  and  A201 );
 a24084a <=( A200  and  a24083a );
 a24085a <=( a24084a  and  a24079a );
 a24089a <=( A298  and  A269 );
 a24090a <=( (not A267)  and  a24089a );
 a24094a <=( A302  and  A300 );
 a24095a <=( (not A299)  and  a24094a );
 a24096a <=( a24095a  and  a24090a );
 a24100a <=( (not A199)  and  A166 );
 a24101a <=( A167  and  a24100a );
 a24105a <=( A203  and  A201 );
 a24106a <=( A200  and  a24105a );
 a24107a <=( a24106a  and  a24101a );
 a24111a <=( (not A298)  and  A269 );
 a24112a <=( (not A267)  and  a24111a );
 a24116a <=( A301  and  A300 );
 a24117a <=( A299  and  a24116a );
 a24118a <=( a24117a  and  a24112a );
 a24122a <=( (not A199)  and  A166 );
 a24123a <=( A167  and  a24122a );
 a24127a <=( A203  and  A201 );
 a24128a <=( A200  and  a24127a );
 a24129a <=( a24128a  and  a24123a );
 a24133a <=( (not A298)  and  A269 );
 a24134a <=( (not A267)  and  a24133a );
 a24138a <=( A302  and  A300 );
 a24139a <=( A299  and  a24138a );
 a24140a <=( a24139a  and  a24134a );
 a24144a <=( (not A199)  and  A166 );
 a24145a <=( A167  and  a24144a );
 a24149a <=( A203  and  A201 );
 a24150a <=( A200  and  a24149a );
 a24151a <=( a24150a  and  a24145a );
 a24155a <=( A298  and  A266 );
 a24156a <=( A265  and  a24155a );
 a24160a <=( A301  and  A300 );
 a24161a <=( (not A299)  and  a24160a );
 a24162a <=( a24161a  and  a24156a );
 a24166a <=( (not A199)  and  A166 );
 a24167a <=( A167  and  a24166a );
 a24171a <=( A203  and  A201 );
 a24172a <=( A200  and  a24171a );
 a24173a <=( a24172a  and  a24167a );
 a24177a <=( A298  and  A266 );
 a24178a <=( A265  and  a24177a );
 a24182a <=( A302  and  A300 );
 a24183a <=( (not A299)  and  a24182a );
 a24184a <=( a24183a  and  a24178a );
 a24188a <=( (not A199)  and  A166 );
 a24189a <=( A167  and  a24188a );
 a24193a <=( A203  and  A201 );
 a24194a <=( A200  and  a24193a );
 a24195a <=( a24194a  and  a24189a );
 a24199a <=( (not A298)  and  A266 );
 a24200a <=( A265  and  a24199a );
 a24204a <=( A301  and  A300 );
 a24205a <=( A299  and  a24204a );
 a24206a <=( a24205a  and  a24200a );
 a24210a <=( (not A199)  and  A166 );
 a24211a <=( A167  and  a24210a );
 a24215a <=( A203  and  A201 );
 a24216a <=( A200  and  a24215a );
 a24217a <=( a24216a  and  a24211a );
 a24221a <=( (not A298)  and  A266 );
 a24222a <=( A265  and  a24221a );
 a24226a <=( A302  and  A300 );
 a24227a <=( A299  and  a24226a );
 a24228a <=( a24227a  and  a24222a );
 a24232a <=( (not A199)  and  A166 );
 a24233a <=( A167  and  a24232a );
 a24237a <=( A203  and  A201 );
 a24238a <=( A200  and  a24237a );
 a24239a <=( a24238a  and  a24233a );
 a24243a <=( A298  and  (not A266) );
 a24244a <=( (not A265)  and  a24243a );
 a24248a <=( A301  and  A300 );
 a24249a <=( (not A299)  and  a24248a );
 a24250a <=( a24249a  and  a24244a );
 a24254a <=( (not A199)  and  A166 );
 a24255a <=( A167  and  a24254a );
 a24259a <=( A203  and  A201 );
 a24260a <=( A200  and  a24259a );
 a24261a <=( a24260a  and  a24255a );
 a24265a <=( A298  and  (not A266) );
 a24266a <=( (not A265)  and  a24265a );
 a24270a <=( A302  and  A300 );
 a24271a <=( (not A299)  and  a24270a );
 a24272a <=( a24271a  and  a24266a );
 a24276a <=( (not A199)  and  A166 );
 a24277a <=( A167  and  a24276a );
 a24281a <=( A203  and  A201 );
 a24282a <=( A200  and  a24281a );
 a24283a <=( a24282a  and  a24277a );
 a24287a <=( (not A298)  and  (not A266) );
 a24288a <=( (not A265)  and  a24287a );
 a24292a <=( A301  and  A300 );
 a24293a <=( A299  and  a24292a );
 a24294a <=( a24293a  and  a24288a );
 a24298a <=( (not A199)  and  A166 );
 a24299a <=( A167  and  a24298a );
 a24303a <=( A203  and  A201 );
 a24304a <=( A200  and  a24303a );
 a24305a <=( a24304a  and  a24299a );
 a24309a <=( (not A298)  and  (not A266) );
 a24310a <=( (not A265)  and  a24309a );
 a24314a <=( A302  and  A300 );
 a24315a <=( A299  and  a24314a );
 a24316a <=( a24315a  and  a24310a );
 a24320a <=( A199  and  A166 );
 a24321a <=( A167  and  a24320a );
 a24325a <=( A202  and  A201 );
 a24326a <=( (not A200)  and  a24325a );
 a24327a <=( a24326a  and  a24321a );
 a24331a <=( A298  and  A268 );
 a24332a <=( (not A267)  and  a24331a );
 a24336a <=( A301  and  A300 );
 a24337a <=( (not A299)  and  a24336a );
 a24338a <=( a24337a  and  a24332a );
 a24342a <=( A199  and  A166 );
 a24343a <=( A167  and  a24342a );
 a24347a <=( A202  and  A201 );
 a24348a <=( (not A200)  and  a24347a );
 a24349a <=( a24348a  and  a24343a );
 a24353a <=( A298  and  A268 );
 a24354a <=( (not A267)  and  a24353a );
 a24358a <=( A302  and  A300 );
 a24359a <=( (not A299)  and  a24358a );
 a24360a <=( a24359a  and  a24354a );
 a24364a <=( A199  and  A166 );
 a24365a <=( A167  and  a24364a );
 a24369a <=( A202  and  A201 );
 a24370a <=( (not A200)  and  a24369a );
 a24371a <=( a24370a  and  a24365a );
 a24375a <=( (not A298)  and  A268 );
 a24376a <=( (not A267)  and  a24375a );
 a24380a <=( A301  and  A300 );
 a24381a <=( A299  and  a24380a );
 a24382a <=( a24381a  and  a24376a );
 a24386a <=( A199  and  A166 );
 a24387a <=( A167  and  a24386a );
 a24391a <=( A202  and  A201 );
 a24392a <=( (not A200)  and  a24391a );
 a24393a <=( a24392a  and  a24387a );
 a24397a <=( (not A298)  and  A268 );
 a24398a <=( (not A267)  and  a24397a );
 a24402a <=( A302  and  A300 );
 a24403a <=( A299  and  a24402a );
 a24404a <=( a24403a  and  a24398a );
 a24408a <=( A199  and  A166 );
 a24409a <=( A167  and  a24408a );
 a24413a <=( A202  and  A201 );
 a24414a <=( (not A200)  and  a24413a );
 a24415a <=( a24414a  and  a24409a );
 a24419a <=( A298  and  A269 );
 a24420a <=( (not A267)  and  a24419a );
 a24424a <=( A301  and  A300 );
 a24425a <=( (not A299)  and  a24424a );
 a24426a <=( a24425a  and  a24420a );
 a24430a <=( A199  and  A166 );
 a24431a <=( A167  and  a24430a );
 a24435a <=( A202  and  A201 );
 a24436a <=( (not A200)  and  a24435a );
 a24437a <=( a24436a  and  a24431a );
 a24441a <=( A298  and  A269 );
 a24442a <=( (not A267)  and  a24441a );
 a24446a <=( A302  and  A300 );
 a24447a <=( (not A299)  and  a24446a );
 a24448a <=( a24447a  and  a24442a );
 a24452a <=( A199  and  A166 );
 a24453a <=( A167  and  a24452a );
 a24457a <=( A202  and  A201 );
 a24458a <=( (not A200)  and  a24457a );
 a24459a <=( a24458a  and  a24453a );
 a24463a <=( (not A298)  and  A269 );
 a24464a <=( (not A267)  and  a24463a );
 a24468a <=( A301  and  A300 );
 a24469a <=( A299  and  a24468a );
 a24470a <=( a24469a  and  a24464a );
 a24474a <=( A199  and  A166 );
 a24475a <=( A167  and  a24474a );
 a24479a <=( A202  and  A201 );
 a24480a <=( (not A200)  and  a24479a );
 a24481a <=( a24480a  and  a24475a );
 a24485a <=( (not A298)  and  A269 );
 a24486a <=( (not A267)  and  a24485a );
 a24490a <=( A302  and  A300 );
 a24491a <=( A299  and  a24490a );
 a24492a <=( a24491a  and  a24486a );
 a24496a <=( A199  and  A166 );
 a24497a <=( A167  and  a24496a );
 a24501a <=( A202  and  A201 );
 a24502a <=( (not A200)  and  a24501a );
 a24503a <=( a24502a  and  a24497a );
 a24507a <=( A298  and  A266 );
 a24508a <=( A265  and  a24507a );
 a24512a <=( A301  and  A300 );
 a24513a <=( (not A299)  and  a24512a );
 a24514a <=( a24513a  and  a24508a );
 a24518a <=( A199  and  A166 );
 a24519a <=( A167  and  a24518a );
 a24523a <=( A202  and  A201 );
 a24524a <=( (not A200)  and  a24523a );
 a24525a <=( a24524a  and  a24519a );
 a24529a <=( A298  and  A266 );
 a24530a <=( A265  and  a24529a );
 a24534a <=( A302  and  A300 );
 a24535a <=( (not A299)  and  a24534a );
 a24536a <=( a24535a  and  a24530a );
 a24540a <=( A199  and  A166 );
 a24541a <=( A167  and  a24540a );
 a24545a <=( A202  and  A201 );
 a24546a <=( (not A200)  and  a24545a );
 a24547a <=( a24546a  and  a24541a );
 a24551a <=( (not A298)  and  A266 );
 a24552a <=( A265  and  a24551a );
 a24556a <=( A301  and  A300 );
 a24557a <=( A299  and  a24556a );
 a24558a <=( a24557a  and  a24552a );
 a24562a <=( A199  and  A166 );
 a24563a <=( A167  and  a24562a );
 a24567a <=( A202  and  A201 );
 a24568a <=( (not A200)  and  a24567a );
 a24569a <=( a24568a  and  a24563a );
 a24573a <=( (not A298)  and  A266 );
 a24574a <=( A265  and  a24573a );
 a24578a <=( A302  and  A300 );
 a24579a <=( A299  and  a24578a );
 a24580a <=( a24579a  and  a24574a );
 a24584a <=( A199  and  A166 );
 a24585a <=( A167  and  a24584a );
 a24589a <=( A202  and  A201 );
 a24590a <=( (not A200)  and  a24589a );
 a24591a <=( a24590a  and  a24585a );
 a24595a <=( A298  and  (not A266) );
 a24596a <=( (not A265)  and  a24595a );
 a24600a <=( A301  and  A300 );
 a24601a <=( (not A299)  and  a24600a );
 a24602a <=( a24601a  and  a24596a );
 a24606a <=( A199  and  A166 );
 a24607a <=( A167  and  a24606a );
 a24611a <=( A202  and  A201 );
 a24612a <=( (not A200)  and  a24611a );
 a24613a <=( a24612a  and  a24607a );
 a24617a <=( A298  and  (not A266) );
 a24618a <=( (not A265)  and  a24617a );
 a24622a <=( A302  and  A300 );
 a24623a <=( (not A299)  and  a24622a );
 a24624a <=( a24623a  and  a24618a );
 a24628a <=( A199  and  A166 );
 a24629a <=( A167  and  a24628a );
 a24633a <=( A202  and  A201 );
 a24634a <=( (not A200)  and  a24633a );
 a24635a <=( a24634a  and  a24629a );
 a24639a <=( (not A298)  and  (not A266) );
 a24640a <=( (not A265)  and  a24639a );
 a24644a <=( A301  and  A300 );
 a24645a <=( A299  and  a24644a );
 a24646a <=( a24645a  and  a24640a );
 a24650a <=( A199  and  A166 );
 a24651a <=( A167  and  a24650a );
 a24655a <=( A202  and  A201 );
 a24656a <=( (not A200)  and  a24655a );
 a24657a <=( a24656a  and  a24651a );
 a24661a <=( (not A298)  and  (not A266) );
 a24662a <=( (not A265)  and  a24661a );
 a24666a <=( A302  and  A300 );
 a24667a <=( A299  and  a24666a );
 a24668a <=( a24667a  and  a24662a );
 a24672a <=( A199  and  A166 );
 a24673a <=( A167  and  a24672a );
 a24677a <=( A203  and  A201 );
 a24678a <=( (not A200)  and  a24677a );
 a24679a <=( a24678a  and  a24673a );
 a24683a <=( A298  and  A268 );
 a24684a <=( (not A267)  and  a24683a );
 a24688a <=( A301  and  A300 );
 a24689a <=( (not A299)  and  a24688a );
 a24690a <=( a24689a  and  a24684a );
 a24694a <=( A199  and  A166 );
 a24695a <=( A167  and  a24694a );
 a24699a <=( A203  and  A201 );
 a24700a <=( (not A200)  and  a24699a );
 a24701a <=( a24700a  and  a24695a );
 a24705a <=( A298  and  A268 );
 a24706a <=( (not A267)  and  a24705a );
 a24710a <=( A302  and  A300 );
 a24711a <=( (not A299)  and  a24710a );
 a24712a <=( a24711a  and  a24706a );
 a24716a <=( A199  and  A166 );
 a24717a <=( A167  and  a24716a );
 a24721a <=( A203  and  A201 );
 a24722a <=( (not A200)  and  a24721a );
 a24723a <=( a24722a  and  a24717a );
 a24727a <=( (not A298)  and  A268 );
 a24728a <=( (not A267)  and  a24727a );
 a24732a <=( A301  and  A300 );
 a24733a <=( A299  and  a24732a );
 a24734a <=( a24733a  and  a24728a );
 a24738a <=( A199  and  A166 );
 a24739a <=( A167  and  a24738a );
 a24743a <=( A203  and  A201 );
 a24744a <=( (not A200)  and  a24743a );
 a24745a <=( a24744a  and  a24739a );
 a24749a <=( (not A298)  and  A268 );
 a24750a <=( (not A267)  and  a24749a );
 a24754a <=( A302  and  A300 );
 a24755a <=( A299  and  a24754a );
 a24756a <=( a24755a  and  a24750a );
 a24760a <=( A199  and  A166 );
 a24761a <=( A167  and  a24760a );
 a24765a <=( A203  and  A201 );
 a24766a <=( (not A200)  and  a24765a );
 a24767a <=( a24766a  and  a24761a );
 a24771a <=( A298  and  A269 );
 a24772a <=( (not A267)  and  a24771a );
 a24776a <=( A301  and  A300 );
 a24777a <=( (not A299)  and  a24776a );
 a24778a <=( a24777a  and  a24772a );
 a24782a <=( A199  and  A166 );
 a24783a <=( A167  and  a24782a );
 a24787a <=( A203  and  A201 );
 a24788a <=( (not A200)  and  a24787a );
 a24789a <=( a24788a  and  a24783a );
 a24793a <=( A298  and  A269 );
 a24794a <=( (not A267)  and  a24793a );
 a24798a <=( A302  and  A300 );
 a24799a <=( (not A299)  and  a24798a );
 a24800a <=( a24799a  and  a24794a );
 a24804a <=( A199  and  A166 );
 a24805a <=( A167  and  a24804a );
 a24809a <=( A203  and  A201 );
 a24810a <=( (not A200)  and  a24809a );
 a24811a <=( a24810a  and  a24805a );
 a24815a <=( (not A298)  and  A269 );
 a24816a <=( (not A267)  and  a24815a );
 a24820a <=( A301  and  A300 );
 a24821a <=( A299  and  a24820a );
 a24822a <=( a24821a  and  a24816a );
 a24826a <=( A199  and  A166 );
 a24827a <=( A167  and  a24826a );
 a24831a <=( A203  and  A201 );
 a24832a <=( (not A200)  and  a24831a );
 a24833a <=( a24832a  and  a24827a );
 a24837a <=( (not A298)  and  A269 );
 a24838a <=( (not A267)  and  a24837a );
 a24842a <=( A302  and  A300 );
 a24843a <=( A299  and  a24842a );
 a24844a <=( a24843a  and  a24838a );
 a24848a <=( A199  and  A166 );
 a24849a <=( A167  and  a24848a );
 a24853a <=( A203  and  A201 );
 a24854a <=( (not A200)  and  a24853a );
 a24855a <=( a24854a  and  a24849a );
 a24859a <=( A298  and  A266 );
 a24860a <=( A265  and  a24859a );
 a24864a <=( A301  and  A300 );
 a24865a <=( (not A299)  and  a24864a );
 a24866a <=( a24865a  and  a24860a );
 a24870a <=( A199  and  A166 );
 a24871a <=( A167  and  a24870a );
 a24875a <=( A203  and  A201 );
 a24876a <=( (not A200)  and  a24875a );
 a24877a <=( a24876a  and  a24871a );
 a24881a <=( A298  and  A266 );
 a24882a <=( A265  and  a24881a );
 a24886a <=( A302  and  A300 );
 a24887a <=( (not A299)  and  a24886a );
 a24888a <=( a24887a  and  a24882a );
 a24892a <=( A199  and  A166 );
 a24893a <=( A167  and  a24892a );
 a24897a <=( A203  and  A201 );
 a24898a <=( (not A200)  and  a24897a );
 a24899a <=( a24898a  and  a24893a );
 a24903a <=( (not A298)  and  A266 );
 a24904a <=( A265  and  a24903a );
 a24908a <=( A301  and  A300 );
 a24909a <=( A299  and  a24908a );
 a24910a <=( a24909a  and  a24904a );
 a24914a <=( A199  and  A166 );
 a24915a <=( A167  and  a24914a );
 a24919a <=( A203  and  A201 );
 a24920a <=( (not A200)  and  a24919a );
 a24921a <=( a24920a  and  a24915a );
 a24925a <=( (not A298)  and  A266 );
 a24926a <=( A265  and  a24925a );
 a24930a <=( A302  and  A300 );
 a24931a <=( A299  and  a24930a );
 a24932a <=( a24931a  and  a24926a );
 a24936a <=( A199  and  A166 );
 a24937a <=( A167  and  a24936a );
 a24941a <=( A203  and  A201 );
 a24942a <=( (not A200)  and  a24941a );
 a24943a <=( a24942a  and  a24937a );
 a24947a <=( A298  and  (not A266) );
 a24948a <=( (not A265)  and  a24947a );
 a24952a <=( A301  and  A300 );
 a24953a <=( (not A299)  and  a24952a );
 a24954a <=( a24953a  and  a24948a );
 a24958a <=( A199  and  A166 );
 a24959a <=( A167  and  a24958a );
 a24963a <=( A203  and  A201 );
 a24964a <=( (not A200)  and  a24963a );
 a24965a <=( a24964a  and  a24959a );
 a24969a <=( A298  and  (not A266) );
 a24970a <=( (not A265)  and  a24969a );
 a24974a <=( A302  and  A300 );
 a24975a <=( (not A299)  and  a24974a );
 a24976a <=( a24975a  and  a24970a );
 a24980a <=( A199  and  A166 );
 a24981a <=( A167  and  a24980a );
 a24985a <=( A203  and  A201 );
 a24986a <=( (not A200)  and  a24985a );
 a24987a <=( a24986a  and  a24981a );
 a24991a <=( (not A298)  and  (not A266) );
 a24992a <=( (not A265)  and  a24991a );
 a24996a <=( A301  and  A300 );
 a24997a <=( A299  and  a24996a );
 a24998a <=( a24997a  and  a24992a );
 a25002a <=( A199  and  A166 );
 a25003a <=( A167  and  a25002a );
 a25007a <=( A203  and  A201 );
 a25008a <=( (not A200)  and  a25007a );
 a25009a <=( a25008a  and  a25003a );
 a25013a <=( (not A298)  and  (not A266) );
 a25014a <=( (not A265)  and  a25013a );
 a25018a <=( A302  and  A300 );
 a25019a <=( A299  and  a25018a );
 a25020a <=( a25019a  and  a25014a );
 a25024a <=( (not A199)  and  A166 );
 a25025a <=( A167  and  a25024a );
 a25029a <=( A266  and  (not A265) );
 a25030a <=( (not A200)  and  a25029a );
 a25031a <=( a25030a  and  a25025a );
 a25035a <=( (not A269)  and  (not A268) );
 a25036a <=( (not A267)  and  a25035a );
 a25040a <=( (not A302)  and  (not A301) );
 a25041a <=( A300  and  a25040a );
 a25042a <=( a25041a  and  a25036a );
 a25046a <=( (not A199)  and  A166 );
 a25047a <=( A167  and  a25046a );
 a25051a <=( (not A266)  and  A265 );
 a25052a <=( (not A200)  and  a25051a );
 a25053a <=( a25052a  and  a25047a );
 a25057a <=( (not A269)  and  (not A268) );
 a25058a <=( (not A267)  and  a25057a );
 a25062a <=( (not A302)  and  (not A301) );
 a25063a <=( A300  and  a25062a );
 a25064a <=( a25063a  and  a25058a );
 a25068a <=( A201  and  (not A166) );
 a25069a <=( (not A167)  and  a25068a );
 a25073a <=( (not A265)  and  (not A203) );
 a25074a <=( (not A202)  and  a25073a );
 a25075a <=( a25074a  and  a25069a );
 a25079a <=( A268  and  A267 );
 a25080a <=( A266  and  a25079a );
 a25084a <=( (not A302)  and  (not A301) );
 a25085a <=( A300  and  a25084a );
 a25086a <=( a25085a  and  a25080a );
 a25090a <=( A201  and  (not A166) );
 a25091a <=( (not A167)  and  a25090a );
 a25095a <=( (not A265)  and  (not A203) );
 a25096a <=( (not A202)  and  a25095a );
 a25097a <=( a25096a  and  a25091a );
 a25101a <=( A269  and  A267 );
 a25102a <=( A266  and  a25101a );
 a25106a <=( (not A302)  and  (not A301) );
 a25107a <=( A300  and  a25106a );
 a25108a <=( a25107a  and  a25102a );
 a25112a <=( A201  and  (not A166) );
 a25113a <=( (not A167)  and  a25112a );
 a25117a <=( (not A265)  and  (not A203) );
 a25118a <=( (not A202)  and  a25117a );
 a25119a <=( a25118a  and  a25113a );
 a25123a <=( (not A268)  and  (not A267) );
 a25124a <=( A266  and  a25123a );
 a25128a <=( A301  and  (not A300) );
 a25129a <=( (not A269)  and  a25128a );
 a25130a <=( a25129a  and  a25124a );
 a25134a <=( A201  and  (not A166) );
 a25135a <=( (not A167)  and  a25134a );
 a25139a <=( (not A265)  and  (not A203) );
 a25140a <=( (not A202)  and  a25139a );
 a25141a <=( a25140a  and  a25135a );
 a25145a <=( (not A268)  and  (not A267) );
 a25146a <=( A266  and  a25145a );
 a25150a <=( A302  and  (not A300) );
 a25151a <=( (not A269)  and  a25150a );
 a25152a <=( a25151a  and  a25146a );
 a25156a <=( A201  and  (not A166) );
 a25157a <=( (not A167)  and  a25156a );
 a25161a <=( (not A265)  and  (not A203) );
 a25162a <=( (not A202)  and  a25161a );
 a25163a <=( a25162a  and  a25157a );
 a25167a <=( (not A268)  and  (not A267) );
 a25168a <=( A266  and  a25167a );
 a25172a <=( A299  and  A298 );
 a25173a <=( (not A269)  and  a25172a );
 a25174a <=( a25173a  and  a25168a );
 a25178a <=( A201  and  (not A166) );
 a25179a <=( (not A167)  and  a25178a );
 a25183a <=( (not A265)  and  (not A203) );
 a25184a <=( (not A202)  and  a25183a );
 a25185a <=( a25184a  and  a25179a );
 a25189a <=( (not A268)  and  (not A267) );
 a25190a <=( A266  and  a25189a );
 a25194a <=( (not A299)  and  (not A298) );
 a25195a <=( (not A269)  and  a25194a );
 a25196a <=( a25195a  and  a25190a );
 a25200a <=( A201  and  (not A166) );
 a25201a <=( (not A167)  and  a25200a );
 a25205a <=( A265  and  (not A203) );
 a25206a <=( (not A202)  and  a25205a );
 a25207a <=( a25206a  and  a25201a );
 a25211a <=( A268  and  A267 );
 a25212a <=( (not A266)  and  a25211a );
 a25216a <=( (not A302)  and  (not A301) );
 a25217a <=( A300  and  a25216a );
 a25218a <=( a25217a  and  a25212a );
 a25222a <=( A201  and  (not A166) );
 a25223a <=( (not A167)  and  a25222a );
 a25227a <=( A265  and  (not A203) );
 a25228a <=( (not A202)  and  a25227a );
 a25229a <=( a25228a  and  a25223a );
 a25233a <=( A269  and  A267 );
 a25234a <=( (not A266)  and  a25233a );
 a25238a <=( (not A302)  and  (not A301) );
 a25239a <=( A300  and  a25238a );
 a25240a <=( a25239a  and  a25234a );
 a25244a <=( A201  and  (not A166) );
 a25245a <=( (not A167)  and  a25244a );
 a25249a <=( A265  and  (not A203) );
 a25250a <=( (not A202)  and  a25249a );
 a25251a <=( a25250a  and  a25245a );
 a25255a <=( (not A268)  and  (not A267) );
 a25256a <=( (not A266)  and  a25255a );
 a25260a <=( A301  and  (not A300) );
 a25261a <=( (not A269)  and  a25260a );
 a25262a <=( a25261a  and  a25256a );
 a25266a <=( A201  and  (not A166) );
 a25267a <=( (not A167)  and  a25266a );
 a25271a <=( A265  and  (not A203) );
 a25272a <=( (not A202)  and  a25271a );
 a25273a <=( a25272a  and  a25267a );
 a25277a <=( (not A268)  and  (not A267) );
 a25278a <=( (not A266)  and  a25277a );
 a25282a <=( A302  and  (not A300) );
 a25283a <=( (not A269)  and  a25282a );
 a25284a <=( a25283a  and  a25278a );
 a25288a <=( A201  and  (not A166) );
 a25289a <=( (not A167)  and  a25288a );
 a25293a <=( A265  and  (not A203) );
 a25294a <=( (not A202)  and  a25293a );
 a25295a <=( a25294a  and  a25289a );
 a25299a <=( (not A268)  and  (not A267) );
 a25300a <=( (not A266)  and  a25299a );
 a25304a <=( A299  and  A298 );
 a25305a <=( (not A269)  and  a25304a );
 a25306a <=( a25305a  and  a25300a );
 a25310a <=( A201  and  (not A166) );
 a25311a <=( (not A167)  and  a25310a );
 a25315a <=( A265  and  (not A203) );
 a25316a <=( (not A202)  and  a25315a );
 a25317a <=( a25316a  and  a25311a );
 a25321a <=( (not A268)  and  (not A267) );
 a25322a <=( (not A266)  and  a25321a );
 a25326a <=( (not A299)  and  (not A298) );
 a25327a <=( (not A269)  and  a25326a );
 a25328a <=( a25327a  and  a25322a );
 a25332a <=( (not A201)  and  (not A166) );
 a25333a <=( (not A167)  and  a25332a );
 a25337a <=( A266  and  (not A265) );
 a25338a <=( A202  and  a25337a );
 a25339a <=( a25338a  and  a25333a );
 a25343a <=( (not A269)  and  (not A268) );
 a25344a <=( (not A267)  and  a25343a );
 a25348a <=( (not A302)  and  (not A301) );
 a25349a <=( A300  and  a25348a );
 a25350a <=( a25349a  and  a25344a );
 a25354a <=( (not A201)  and  (not A166) );
 a25355a <=( (not A167)  and  a25354a );
 a25359a <=( (not A266)  and  A265 );
 a25360a <=( A202  and  a25359a );
 a25361a <=( a25360a  and  a25355a );
 a25365a <=( (not A269)  and  (not A268) );
 a25366a <=( (not A267)  and  a25365a );
 a25370a <=( (not A302)  and  (not A301) );
 a25371a <=( A300  and  a25370a );
 a25372a <=( a25371a  and  a25366a );
 a25376a <=( (not A201)  and  (not A166) );
 a25377a <=( (not A167)  and  a25376a );
 a25381a <=( A266  and  (not A265) );
 a25382a <=( A203  and  a25381a );
 a25383a <=( a25382a  and  a25377a );
 a25387a <=( (not A269)  and  (not A268) );
 a25388a <=( (not A267)  and  a25387a );
 a25392a <=( (not A302)  and  (not A301) );
 a25393a <=( A300  and  a25392a );
 a25394a <=( a25393a  and  a25388a );
 a25398a <=( (not A201)  and  (not A166) );
 a25399a <=( (not A167)  and  a25398a );
 a25403a <=( (not A266)  and  A265 );
 a25404a <=( A203  and  a25403a );
 a25405a <=( a25404a  and  a25399a );
 a25409a <=( (not A269)  and  (not A268) );
 a25410a <=( (not A267)  and  a25409a );
 a25414a <=( (not A302)  and  (not A301) );
 a25415a <=( A300  and  a25414a );
 a25416a <=( a25415a  and  a25410a );
 a25420a <=( A199  and  (not A166) );
 a25421a <=( (not A167)  and  a25420a );
 a25425a <=( A266  and  (not A265) );
 a25426a <=( A200  and  a25425a );
 a25427a <=( a25426a  and  a25421a );
 a25431a <=( (not A269)  and  (not A268) );
 a25432a <=( (not A267)  and  a25431a );
 a25436a <=( (not A302)  and  (not A301) );
 a25437a <=( A300  and  a25436a );
 a25438a <=( a25437a  and  a25432a );
 a25442a <=( A199  and  (not A166) );
 a25443a <=( (not A167)  and  a25442a );
 a25447a <=( (not A266)  and  A265 );
 a25448a <=( A200  and  a25447a );
 a25449a <=( a25448a  and  a25443a );
 a25453a <=( (not A269)  and  (not A268) );
 a25454a <=( (not A267)  and  a25453a );
 a25458a <=( (not A302)  and  (not A301) );
 a25459a <=( A300  and  a25458a );
 a25460a <=( a25459a  and  a25454a );
 a25464a <=( (not A199)  and  (not A166) );
 a25465a <=( (not A167)  and  a25464a );
 a25469a <=( A202  and  A201 );
 a25470a <=( A200  and  a25469a );
 a25471a <=( a25470a  and  a25465a );
 a25475a <=( A298  and  A268 );
 a25476a <=( (not A267)  and  a25475a );
 a25480a <=( A301  and  A300 );
 a25481a <=( (not A299)  and  a25480a );
 a25482a <=( a25481a  and  a25476a );
 a25486a <=( (not A199)  and  (not A166) );
 a25487a <=( (not A167)  and  a25486a );
 a25491a <=( A202  and  A201 );
 a25492a <=( A200  and  a25491a );
 a25493a <=( a25492a  and  a25487a );
 a25497a <=( A298  and  A268 );
 a25498a <=( (not A267)  and  a25497a );
 a25502a <=( A302  and  A300 );
 a25503a <=( (not A299)  and  a25502a );
 a25504a <=( a25503a  and  a25498a );
 a25508a <=( (not A199)  and  (not A166) );
 a25509a <=( (not A167)  and  a25508a );
 a25513a <=( A202  and  A201 );
 a25514a <=( A200  and  a25513a );
 a25515a <=( a25514a  and  a25509a );
 a25519a <=( (not A298)  and  A268 );
 a25520a <=( (not A267)  and  a25519a );
 a25524a <=( A301  and  A300 );
 a25525a <=( A299  and  a25524a );
 a25526a <=( a25525a  and  a25520a );
 a25530a <=( (not A199)  and  (not A166) );
 a25531a <=( (not A167)  and  a25530a );
 a25535a <=( A202  and  A201 );
 a25536a <=( A200  and  a25535a );
 a25537a <=( a25536a  and  a25531a );
 a25541a <=( (not A298)  and  A268 );
 a25542a <=( (not A267)  and  a25541a );
 a25546a <=( A302  and  A300 );
 a25547a <=( A299  and  a25546a );
 a25548a <=( a25547a  and  a25542a );
 a25552a <=( (not A199)  and  (not A166) );
 a25553a <=( (not A167)  and  a25552a );
 a25557a <=( A202  and  A201 );
 a25558a <=( A200  and  a25557a );
 a25559a <=( a25558a  and  a25553a );
 a25563a <=( A298  and  A269 );
 a25564a <=( (not A267)  and  a25563a );
 a25568a <=( A301  and  A300 );
 a25569a <=( (not A299)  and  a25568a );
 a25570a <=( a25569a  and  a25564a );
 a25574a <=( (not A199)  and  (not A166) );
 a25575a <=( (not A167)  and  a25574a );
 a25579a <=( A202  and  A201 );
 a25580a <=( A200  and  a25579a );
 a25581a <=( a25580a  and  a25575a );
 a25585a <=( A298  and  A269 );
 a25586a <=( (not A267)  and  a25585a );
 a25590a <=( A302  and  A300 );
 a25591a <=( (not A299)  and  a25590a );
 a25592a <=( a25591a  and  a25586a );
 a25596a <=( (not A199)  and  (not A166) );
 a25597a <=( (not A167)  and  a25596a );
 a25601a <=( A202  and  A201 );
 a25602a <=( A200  and  a25601a );
 a25603a <=( a25602a  and  a25597a );
 a25607a <=( (not A298)  and  A269 );
 a25608a <=( (not A267)  and  a25607a );
 a25612a <=( A301  and  A300 );
 a25613a <=( A299  and  a25612a );
 a25614a <=( a25613a  and  a25608a );
 a25618a <=( (not A199)  and  (not A166) );
 a25619a <=( (not A167)  and  a25618a );
 a25623a <=( A202  and  A201 );
 a25624a <=( A200  and  a25623a );
 a25625a <=( a25624a  and  a25619a );
 a25629a <=( (not A298)  and  A269 );
 a25630a <=( (not A267)  and  a25629a );
 a25634a <=( A302  and  A300 );
 a25635a <=( A299  and  a25634a );
 a25636a <=( a25635a  and  a25630a );
 a25640a <=( (not A199)  and  (not A166) );
 a25641a <=( (not A167)  and  a25640a );
 a25645a <=( A202  and  A201 );
 a25646a <=( A200  and  a25645a );
 a25647a <=( a25646a  and  a25641a );
 a25651a <=( A298  and  A266 );
 a25652a <=( A265  and  a25651a );
 a25656a <=( A301  and  A300 );
 a25657a <=( (not A299)  and  a25656a );
 a25658a <=( a25657a  and  a25652a );
 a25662a <=( (not A199)  and  (not A166) );
 a25663a <=( (not A167)  and  a25662a );
 a25667a <=( A202  and  A201 );
 a25668a <=( A200  and  a25667a );
 a25669a <=( a25668a  and  a25663a );
 a25673a <=( A298  and  A266 );
 a25674a <=( A265  and  a25673a );
 a25678a <=( A302  and  A300 );
 a25679a <=( (not A299)  and  a25678a );
 a25680a <=( a25679a  and  a25674a );
 a25684a <=( (not A199)  and  (not A166) );
 a25685a <=( (not A167)  and  a25684a );
 a25689a <=( A202  and  A201 );
 a25690a <=( A200  and  a25689a );
 a25691a <=( a25690a  and  a25685a );
 a25695a <=( (not A298)  and  A266 );
 a25696a <=( A265  and  a25695a );
 a25700a <=( A301  and  A300 );
 a25701a <=( A299  and  a25700a );
 a25702a <=( a25701a  and  a25696a );
 a25706a <=( (not A199)  and  (not A166) );
 a25707a <=( (not A167)  and  a25706a );
 a25711a <=( A202  and  A201 );
 a25712a <=( A200  and  a25711a );
 a25713a <=( a25712a  and  a25707a );
 a25717a <=( (not A298)  and  A266 );
 a25718a <=( A265  and  a25717a );
 a25722a <=( A302  and  A300 );
 a25723a <=( A299  and  a25722a );
 a25724a <=( a25723a  and  a25718a );
 a25728a <=( (not A199)  and  (not A166) );
 a25729a <=( (not A167)  and  a25728a );
 a25733a <=( A202  and  A201 );
 a25734a <=( A200  and  a25733a );
 a25735a <=( a25734a  and  a25729a );
 a25739a <=( A298  and  (not A266) );
 a25740a <=( (not A265)  and  a25739a );
 a25744a <=( A301  and  A300 );
 a25745a <=( (not A299)  and  a25744a );
 a25746a <=( a25745a  and  a25740a );
 a25750a <=( (not A199)  and  (not A166) );
 a25751a <=( (not A167)  and  a25750a );
 a25755a <=( A202  and  A201 );
 a25756a <=( A200  and  a25755a );
 a25757a <=( a25756a  and  a25751a );
 a25761a <=( A298  and  (not A266) );
 a25762a <=( (not A265)  and  a25761a );
 a25766a <=( A302  and  A300 );
 a25767a <=( (not A299)  and  a25766a );
 a25768a <=( a25767a  and  a25762a );
 a25772a <=( (not A199)  and  (not A166) );
 a25773a <=( (not A167)  and  a25772a );
 a25777a <=( A202  and  A201 );
 a25778a <=( A200  and  a25777a );
 a25779a <=( a25778a  and  a25773a );
 a25783a <=( (not A298)  and  (not A266) );
 a25784a <=( (not A265)  and  a25783a );
 a25788a <=( A301  and  A300 );
 a25789a <=( A299  and  a25788a );
 a25790a <=( a25789a  and  a25784a );
 a25794a <=( (not A199)  and  (not A166) );
 a25795a <=( (not A167)  and  a25794a );
 a25799a <=( A202  and  A201 );
 a25800a <=( A200  and  a25799a );
 a25801a <=( a25800a  and  a25795a );
 a25805a <=( (not A298)  and  (not A266) );
 a25806a <=( (not A265)  and  a25805a );
 a25810a <=( A302  and  A300 );
 a25811a <=( A299  and  a25810a );
 a25812a <=( a25811a  and  a25806a );
 a25816a <=( (not A199)  and  (not A166) );
 a25817a <=( (not A167)  and  a25816a );
 a25821a <=( A203  and  A201 );
 a25822a <=( A200  and  a25821a );
 a25823a <=( a25822a  and  a25817a );
 a25827a <=( A298  and  A268 );
 a25828a <=( (not A267)  and  a25827a );
 a25832a <=( A301  and  A300 );
 a25833a <=( (not A299)  and  a25832a );
 a25834a <=( a25833a  and  a25828a );
 a25838a <=( (not A199)  and  (not A166) );
 a25839a <=( (not A167)  and  a25838a );
 a25843a <=( A203  and  A201 );
 a25844a <=( A200  and  a25843a );
 a25845a <=( a25844a  and  a25839a );
 a25849a <=( A298  and  A268 );
 a25850a <=( (not A267)  and  a25849a );
 a25854a <=( A302  and  A300 );
 a25855a <=( (not A299)  and  a25854a );
 a25856a <=( a25855a  and  a25850a );
 a25860a <=( (not A199)  and  (not A166) );
 a25861a <=( (not A167)  and  a25860a );
 a25865a <=( A203  and  A201 );
 a25866a <=( A200  and  a25865a );
 a25867a <=( a25866a  and  a25861a );
 a25871a <=( (not A298)  and  A268 );
 a25872a <=( (not A267)  and  a25871a );
 a25876a <=( A301  and  A300 );
 a25877a <=( A299  and  a25876a );
 a25878a <=( a25877a  and  a25872a );
 a25882a <=( (not A199)  and  (not A166) );
 a25883a <=( (not A167)  and  a25882a );
 a25887a <=( A203  and  A201 );
 a25888a <=( A200  and  a25887a );
 a25889a <=( a25888a  and  a25883a );
 a25893a <=( (not A298)  and  A268 );
 a25894a <=( (not A267)  and  a25893a );
 a25898a <=( A302  and  A300 );
 a25899a <=( A299  and  a25898a );
 a25900a <=( a25899a  and  a25894a );
 a25904a <=( (not A199)  and  (not A166) );
 a25905a <=( (not A167)  and  a25904a );
 a25909a <=( A203  and  A201 );
 a25910a <=( A200  and  a25909a );
 a25911a <=( a25910a  and  a25905a );
 a25915a <=( A298  and  A269 );
 a25916a <=( (not A267)  and  a25915a );
 a25920a <=( A301  and  A300 );
 a25921a <=( (not A299)  and  a25920a );
 a25922a <=( a25921a  and  a25916a );
 a25926a <=( (not A199)  and  (not A166) );
 a25927a <=( (not A167)  and  a25926a );
 a25931a <=( A203  and  A201 );
 a25932a <=( A200  and  a25931a );
 a25933a <=( a25932a  and  a25927a );
 a25937a <=( A298  and  A269 );
 a25938a <=( (not A267)  and  a25937a );
 a25942a <=( A302  and  A300 );
 a25943a <=( (not A299)  and  a25942a );
 a25944a <=( a25943a  and  a25938a );
 a25948a <=( (not A199)  and  (not A166) );
 a25949a <=( (not A167)  and  a25948a );
 a25953a <=( A203  and  A201 );
 a25954a <=( A200  and  a25953a );
 a25955a <=( a25954a  and  a25949a );
 a25959a <=( (not A298)  and  A269 );
 a25960a <=( (not A267)  and  a25959a );
 a25964a <=( A301  and  A300 );
 a25965a <=( A299  and  a25964a );
 a25966a <=( a25965a  and  a25960a );
 a25970a <=( (not A199)  and  (not A166) );
 a25971a <=( (not A167)  and  a25970a );
 a25975a <=( A203  and  A201 );
 a25976a <=( A200  and  a25975a );
 a25977a <=( a25976a  and  a25971a );
 a25981a <=( (not A298)  and  A269 );
 a25982a <=( (not A267)  and  a25981a );
 a25986a <=( A302  and  A300 );
 a25987a <=( A299  and  a25986a );
 a25988a <=( a25987a  and  a25982a );
 a25992a <=( (not A199)  and  (not A166) );
 a25993a <=( (not A167)  and  a25992a );
 a25997a <=( A203  and  A201 );
 a25998a <=( A200  and  a25997a );
 a25999a <=( a25998a  and  a25993a );
 a26003a <=( A298  and  A266 );
 a26004a <=( A265  and  a26003a );
 a26008a <=( A301  and  A300 );
 a26009a <=( (not A299)  and  a26008a );
 a26010a <=( a26009a  and  a26004a );
 a26014a <=( (not A199)  and  (not A166) );
 a26015a <=( (not A167)  and  a26014a );
 a26019a <=( A203  and  A201 );
 a26020a <=( A200  and  a26019a );
 a26021a <=( a26020a  and  a26015a );
 a26025a <=( A298  and  A266 );
 a26026a <=( A265  and  a26025a );
 a26030a <=( A302  and  A300 );
 a26031a <=( (not A299)  and  a26030a );
 a26032a <=( a26031a  and  a26026a );
 a26036a <=( (not A199)  and  (not A166) );
 a26037a <=( (not A167)  and  a26036a );
 a26041a <=( A203  and  A201 );
 a26042a <=( A200  and  a26041a );
 a26043a <=( a26042a  and  a26037a );
 a26047a <=( (not A298)  and  A266 );
 a26048a <=( A265  and  a26047a );
 a26052a <=( A301  and  A300 );
 a26053a <=( A299  and  a26052a );
 a26054a <=( a26053a  and  a26048a );
 a26058a <=( (not A199)  and  (not A166) );
 a26059a <=( (not A167)  and  a26058a );
 a26063a <=( A203  and  A201 );
 a26064a <=( A200  and  a26063a );
 a26065a <=( a26064a  and  a26059a );
 a26069a <=( (not A298)  and  A266 );
 a26070a <=( A265  and  a26069a );
 a26074a <=( A302  and  A300 );
 a26075a <=( A299  and  a26074a );
 a26076a <=( a26075a  and  a26070a );
 a26080a <=( (not A199)  and  (not A166) );
 a26081a <=( (not A167)  and  a26080a );
 a26085a <=( A203  and  A201 );
 a26086a <=( A200  and  a26085a );
 a26087a <=( a26086a  and  a26081a );
 a26091a <=( A298  and  (not A266) );
 a26092a <=( (not A265)  and  a26091a );
 a26096a <=( A301  and  A300 );
 a26097a <=( (not A299)  and  a26096a );
 a26098a <=( a26097a  and  a26092a );
 a26102a <=( (not A199)  and  (not A166) );
 a26103a <=( (not A167)  and  a26102a );
 a26107a <=( A203  and  A201 );
 a26108a <=( A200  and  a26107a );
 a26109a <=( a26108a  and  a26103a );
 a26113a <=( A298  and  (not A266) );
 a26114a <=( (not A265)  and  a26113a );
 a26118a <=( A302  and  A300 );
 a26119a <=( (not A299)  and  a26118a );
 a26120a <=( a26119a  and  a26114a );
 a26124a <=( (not A199)  and  (not A166) );
 a26125a <=( (not A167)  and  a26124a );
 a26129a <=( A203  and  A201 );
 a26130a <=( A200  and  a26129a );
 a26131a <=( a26130a  and  a26125a );
 a26135a <=( (not A298)  and  (not A266) );
 a26136a <=( (not A265)  and  a26135a );
 a26140a <=( A301  and  A300 );
 a26141a <=( A299  and  a26140a );
 a26142a <=( a26141a  and  a26136a );
 a26146a <=( (not A199)  and  (not A166) );
 a26147a <=( (not A167)  and  a26146a );
 a26151a <=( A203  and  A201 );
 a26152a <=( A200  and  a26151a );
 a26153a <=( a26152a  and  a26147a );
 a26157a <=( (not A298)  and  (not A266) );
 a26158a <=( (not A265)  and  a26157a );
 a26162a <=( A302  and  A300 );
 a26163a <=( A299  and  a26162a );
 a26164a <=( a26163a  and  a26158a );
 a26168a <=( A199  and  (not A166) );
 a26169a <=( (not A167)  and  a26168a );
 a26173a <=( A202  and  A201 );
 a26174a <=( (not A200)  and  a26173a );
 a26175a <=( a26174a  and  a26169a );
 a26179a <=( A298  and  A268 );
 a26180a <=( (not A267)  and  a26179a );
 a26184a <=( A301  and  A300 );
 a26185a <=( (not A299)  and  a26184a );
 a26186a <=( a26185a  and  a26180a );
 a26190a <=( A199  and  (not A166) );
 a26191a <=( (not A167)  and  a26190a );
 a26195a <=( A202  and  A201 );
 a26196a <=( (not A200)  and  a26195a );
 a26197a <=( a26196a  and  a26191a );
 a26201a <=( A298  and  A268 );
 a26202a <=( (not A267)  and  a26201a );
 a26206a <=( A302  and  A300 );
 a26207a <=( (not A299)  and  a26206a );
 a26208a <=( a26207a  and  a26202a );
 a26212a <=( A199  and  (not A166) );
 a26213a <=( (not A167)  and  a26212a );
 a26217a <=( A202  and  A201 );
 a26218a <=( (not A200)  and  a26217a );
 a26219a <=( a26218a  and  a26213a );
 a26223a <=( (not A298)  and  A268 );
 a26224a <=( (not A267)  and  a26223a );
 a26228a <=( A301  and  A300 );
 a26229a <=( A299  and  a26228a );
 a26230a <=( a26229a  and  a26224a );
 a26234a <=( A199  and  (not A166) );
 a26235a <=( (not A167)  and  a26234a );
 a26239a <=( A202  and  A201 );
 a26240a <=( (not A200)  and  a26239a );
 a26241a <=( a26240a  and  a26235a );
 a26245a <=( (not A298)  and  A268 );
 a26246a <=( (not A267)  and  a26245a );
 a26250a <=( A302  and  A300 );
 a26251a <=( A299  and  a26250a );
 a26252a <=( a26251a  and  a26246a );
 a26256a <=( A199  and  (not A166) );
 a26257a <=( (not A167)  and  a26256a );
 a26261a <=( A202  and  A201 );
 a26262a <=( (not A200)  and  a26261a );
 a26263a <=( a26262a  and  a26257a );
 a26267a <=( A298  and  A269 );
 a26268a <=( (not A267)  and  a26267a );
 a26272a <=( A301  and  A300 );
 a26273a <=( (not A299)  and  a26272a );
 a26274a <=( a26273a  and  a26268a );
 a26278a <=( A199  and  (not A166) );
 a26279a <=( (not A167)  and  a26278a );
 a26283a <=( A202  and  A201 );
 a26284a <=( (not A200)  and  a26283a );
 a26285a <=( a26284a  and  a26279a );
 a26289a <=( A298  and  A269 );
 a26290a <=( (not A267)  and  a26289a );
 a26294a <=( A302  and  A300 );
 a26295a <=( (not A299)  and  a26294a );
 a26296a <=( a26295a  and  a26290a );
 a26300a <=( A199  and  (not A166) );
 a26301a <=( (not A167)  and  a26300a );
 a26305a <=( A202  and  A201 );
 a26306a <=( (not A200)  and  a26305a );
 a26307a <=( a26306a  and  a26301a );
 a26311a <=( (not A298)  and  A269 );
 a26312a <=( (not A267)  and  a26311a );
 a26316a <=( A301  and  A300 );
 a26317a <=( A299  and  a26316a );
 a26318a <=( a26317a  and  a26312a );
 a26322a <=( A199  and  (not A166) );
 a26323a <=( (not A167)  and  a26322a );
 a26327a <=( A202  and  A201 );
 a26328a <=( (not A200)  and  a26327a );
 a26329a <=( a26328a  and  a26323a );
 a26333a <=( (not A298)  and  A269 );
 a26334a <=( (not A267)  and  a26333a );
 a26338a <=( A302  and  A300 );
 a26339a <=( A299  and  a26338a );
 a26340a <=( a26339a  and  a26334a );
 a26344a <=( A199  and  (not A166) );
 a26345a <=( (not A167)  and  a26344a );
 a26349a <=( A202  and  A201 );
 a26350a <=( (not A200)  and  a26349a );
 a26351a <=( a26350a  and  a26345a );
 a26355a <=( A298  and  A266 );
 a26356a <=( A265  and  a26355a );
 a26360a <=( A301  and  A300 );
 a26361a <=( (not A299)  and  a26360a );
 a26362a <=( a26361a  and  a26356a );
 a26366a <=( A199  and  (not A166) );
 a26367a <=( (not A167)  and  a26366a );
 a26371a <=( A202  and  A201 );
 a26372a <=( (not A200)  and  a26371a );
 a26373a <=( a26372a  and  a26367a );
 a26377a <=( A298  and  A266 );
 a26378a <=( A265  and  a26377a );
 a26382a <=( A302  and  A300 );
 a26383a <=( (not A299)  and  a26382a );
 a26384a <=( a26383a  and  a26378a );
 a26388a <=( A199  and  (not A166) );
 a26389a <=( (not A167)  and  a26388a );
 a26393a <=( A202  and  A201 );
 a26394a <=( (not A200)  and  a26393a );
 a26395a <=( a26394a  and  a26389a );
 a26399a <=( (not A298)  and  A266 );
 a26400a <=( A265  and  a26399a );
 a26404a <=( A301  and  A300 );
 a26405a <=( A299  and  a26404a );
 a26406a <=( a26405a  and  a26400a );
 a26410a <=( A199  and  (not A166) );
 a26411a <=( (not A167)  and  a26410a );
 a26415a <=( A202  and  A201 );
 a26416a <=( (not A200)  and  a26415a );
 a26417a <=( a26416a  and  a26411a );
 a26421a <=( (not A298)  and  A266 );
 a26422a <=( A265  and  a26421a );
 a26426a <=( A302  and  A300 );
 a26427a <=( A299  and  a26426a );
 a26428a <=( a26427a  and  a26422a );
 a26432a <=( A199  and  (not A166) );
 a26433a <=( (not A167)  and  a26432a );
 a26437a <=( A202  and  A201 );
 a26438a <=( (not A200)  and  a26437a );
 a26439a <=( a26438a  and  a26433a );
 a26443a <=( A298  and  (not A266) );
 a26444a <=( (not A265)  and  a26443a );
 a26448a <=( A301  and  A300 );
 a26449a <=( (not A299)  and  a26448a );
 a26450a <=( a26449a  and  a26444a );
 a26454a <=( A199  and  (not A166) );
 a26455a <=( (not A167)  and  a26454a );
 a26459a <=( A202  and  A201 );
 a26460a <=( (not A200)  and  a26459a );
 a26461a <=( a26460a  and  a26455a );
 a26465a <=( A298  and  (not A266) );
 a26466a <=( (not A265)  and  a26465a );
 a26470a <=( A302  and  A300 );
 a26471a <=( (not A299)  and  a26470a );
 a26472a <=( a26471a  and  a26466a );
 a26476a <=( A199  and  (not A166) );
 a26477a <=( (not A167)  and  a26476a );
 a26481a <=( A202  and  A201 );
 a26482a <=( (not A200)  and  a26481a );
 a26483a <=( a26482a  and  a26477a );
 a26487a <=( (not A298)  and  (not A266) );
 a26488a <=( (not A265)  and  a26487a );
 a26492a <=( A301  and  A300 );
 a26493a <=( A299  and  a26492a );
 a26494a <=( a26493a  and  a26488a );
 a26498a <=( A199  and  (not A166) );
 a26499a <=( (not A167)  and  a26498a );
 a26503a <=( A202  and  A201 );
 a26504a <=( (not A200)  and  a26503a );
 a26505a <=( a26504a  and  a26499a );
 a26509a <=( (not A298)  and  (not A266) );
 a26510a <=( (not A265)  and  a26509a );
 a26514a <=( A302  and  A300 );
 a26515a <=( A299  and  a26514a );
 a26516a <=( a26515a  and  a26510a );
 a26520a <=( A199  and  (not A166) );
 a26521a <=( (not A167)  and  a26520a );
 a26525a <=( A203  and  A201 );
 a26526a <=( (not A200)  and  a26525a );
 a26527a <=( a26526a  and  a26521a );
 a26531a <=( A298  and  A268 );
 a26532a <=( (not A267)  and  a26531a );
 a26536a <=( A301  and  A300 );
 a26537a <=( (not A299)  and  a26536a );
 a26538a <=( a26537a  and  a26532a );
 a26542a <=( A199  and  (not A166) );
 a26543a <=( (not A167)  and  a26542a );
 a26547a <=( A203  and  A201 );
 a26548a <=( (not A200)  and  a26547a );
 a26549a <=( a26548a  and  a26543a );
 a26553a <=( A298  and  A268 );
 a26554a <=( (not A267)  and  a26553a );
 a26558a <=( A302  and  A300 );
 a26559a <=( (not A299)  and  a26558a );
 a26560a <=( a26559a  and  a26554a );
 a26564a <=( A199  and  (not A166) );
 a26565a <=( (not A167)  and  a26564a );
 a26569a <=( A203  and  A201 );
 a26570a <=( (not A200)  and  a26569a );
 a26571a <=( a26570a  and  a26565a );
 a26575a <=( (not A298)  and  A268 );
 a26576a <=( (not A267)  and  a26575a );
 a26580a <=( A301  and  A300 );
 a26581a <=( A299  and  a26580a );
 a26582a <=( a26581a  and  a26576a );
 a26586a <=( A199  and  (not A166) );
 a26587a <=( (not A167)  and  a26586a );
 a26591a <=( A203  and  A201 );
 a26592a <=( (not A200)  and  a26591a );
 a26593a <=( a26592a  and  a26587a );
 a26597a <=( (not A298)  and  A268 );
 a26598a <=( (not A267)  and  a26597a );
 a26602a <=( A302  and  A300 );
 a26603a <=( A299  and  a26602a );
 a26604a <=( a26603a  and  a26598a );
 a26608a <=( A199  and  (not A166) );
 a26609a <=( (not A167)  and  a26608a );
 a26613a <=( A203  and  A201 );
 a26614a <=( (not A200)  and  a26613a );
 a26615a <=( a26614a  and  a26609a );
 a26619a <=( A298  and  A269 );
 a26620a <=( (not A267)  and  a26619a );
 a26624a <=( A301  and  A300 );
 a26625a <=( (not A299)  and  a26624a );
 a26626a <=( a26625a  and  a26620a );
 a26630a <=( A199  and  (not A166) );
 a26631a <=( (not A167)  and  a26630a );
 a26635a <=( A203  and  A201 );
 a26636a <=( (not A200)  and  a26635a );
 a26637a <=( a26636a  and  a26631a );
 a26641a <=( A298  and  A269 );
 a26642a <=( (not A267)  and  a26641a );
 a26646a <=( A302  and  A300 );
 a26647a <=( (not A299)  and  a26646a );
 a26648a <=( a26647a  and  a26642a );
 a26652a <=( A199  and  (not A166) );
 a26653a <=( (not A167)  and  a26652a );
 a26657a <=( A203  and  A201 );
 a26658a <=( (not A200)  and  a26657a );
 a26659a <=( a26658a  and  a26653a );
 a26663a <=( (not A298)  and  A269 );
 a26664a <=( (not A267)  and  a26663a );
 a26668a <=( A301  and  A300 );
 a26669a <=( A299  and  a26668a );
 a26670a <=( a26669a  and  a26664a );
 a26674a <=( A199  and  (not A166) );
 a26675a <=( (not A167)  and  a26674a );
 a26679a <=( A203  and  A201 );
 a26680a <=( (not A200)  and  a26679a );
 a26681a <=( a26680a  and  a26675a );
 a26685a <=( (not A298)  and  A269 );
 a26686a <=( (not A267)  and  a26685a );
 a26690a <=( A302  and  A300 );
 a26691a <=( A299  and  a26690a );
 a26692a <=( a26691a  and  a26686a );
 a26696a <=( A199  and  (not A166) );
 a26697a <=( (not A167)  and  a26696a );
 a26701a <=( A203  and  A201 );
 a26702a <=( (not A200)  and  a26701a );
 a26703a <=( a26702a  and  a26697a );
 a26707a <=( A298  and  A266 );
 a26708a <=( A265  and  a26707a );
 a26712a <=( A301  and  A300 );
 a26713a <=( (not A299)  and  a26712a );
 a26714a <=( a26713a  and  a26708a );
 a26718a <=( A199  and  (not A166) );
 a26719a <=( (not A167)  and  a26718a );
 a26723a <=( A203  and  A201 );
 a26724a <=( (not A200)  and  a26723a );
 a26725a <=( a26724a  and  a26719a );
 a26729a <=( A298  and  A266 );
 a26730a <=( A265  and  a26729a );
 a26734a <=( A302  and  A300 );
 a26735a <=( (not A299)  and  a26734a );
 a26736a <=( a26735a  and  a26730a );
 a26740a <=( A199  and  (not A166) );
 a26741a <=( (not A167)  and  a26740a );
 a26745a <=( A203  and  A201 );
 a26746a <=( (not A200)  and  a26745a );
 a26747a <=( a26746a  and  a26741a );
 a26751a <=( (not A298)  and  A266 );
 a26752a <=( A265  and  a26751a );
 a26756a <=( A301  and  A300 );
 a26757a <=( A299  and  a26756a );
 a26758a <=( a26757a  and  a26752a );
 a26762a <=( A199  and  (not A166) );
 a26763a <=( (not A167)  and  a26762a );
 a26767a <=( A203  and  A201 );
 a26768a <=( (not A200)  and  a26767a );
 a26769a <=( a26768a  and  a26763a );
 a26773a <=( (not A298)  and  A266 );
 a26774a <=( A265  and  a26773a );
 a26778a <=( A302  and  A300 );
 a26779a <=( A299  and  a26778a );
 a26780a <=( a26779a  and  a26774a );
 a26784a <=( A199  and  (not A166) );
 a26785a <=( (not A167)  and  a26784a );
 a26789a <=( A203  and  A201 );
 a26790a <=( (not A200)  and  a26789a );
 a26791a <=( a26790a  and  a26785a );
 a26795a <=( A298  and  (not A266) );
 a26796a <=( (not A265)  and  a26795a );
 a26800a <=( A301  and  A300 );
 a26801a <=( (not A299)  and  a26800a );
 a26802a <=( a26801a  and  a26796a );
 a26806a <=( A199  and  (not A166) );
 a26807a <=( (not A167)  and  a26806a );
 a26811a <=( A203  and  A201 );
 a26812a <=( (not A200)  and  a26811a );
 a26813a <=( a26812a  and  a26807a );
 a26817a <=( A298  and  (not A266) );
 a26818a <=( (not A265)  and  a26817a );
 a26822a <=( A302  and  A300 );
 a26823a <=( (not A299)  and  a26822a );
 a26824a <=( a26823a  and  a26818a );
 a26828a <=( A199  and  (not A166) );
 a26829a <=( (not A167)  and  a26828a );
 a26833a <=( A203  and  A201 );
 a26834a <=( (not A200)  and  a26833a );
 a26835a <=( a26834a  and  a26829a );
 a26839a <=( (not A298)  and  (not A266) );
 a26840a <=( (not A265)  and  a26839a );
 a26844a <=( A301  and  A300 );
 a26845a <=( A299  and  a26844a );
 a26846a <=( a26845a  and  a26840a );
 a26850a <=( A199  and  (not A166) );
 a26851a <=( (not A167)  and  a26850a );
 a26855a <=( A203  and  A201 );
 a26856a <=( (not A200)  and  a26855a );
 a26857a <=( a26856a  and  a26851a );
 a26861a <=( (not A298)  and  (not A266) );
 a26862a <=( (not A265)  and  a26861a );
 a26866a <=( A302  and  A300 );
 a26867a <=( A299  and  a26866a );
 a26868a <=( a26867a  and  a26862a );
 a26872a <=( (not A199)  and  (not A166) );
 a26873a <=( (not A167)  and  a26872a );
 a26877a <=( A266  and  (not A265) );
 a26878a <=( (not A200)  and  a26877a );
 a26879a <=( a26878a  and  a26873a );
 a26883a <=( (not A269)  and  (not A268) );
 a26884a <=( (not A267)  and  a26883a );
 a26888a <=( (not A302)  and  (not A301) );
 a26889a <=( A300  and  a26888a );
 a26890a <=( a26889a  and  a26884a );
 a26894a <=( (not A199)  and  (not A166) );
 a26895a <=( (not A167)  and  a26894a );
 a26899a <=( (not A266)  and  A265 );
 a26900a <=( (not A200)  and  a26899a );
 a26901a <=( a26900a  and  a26895a );
 a26905a <=( (not A269)  and  (not A268) );
 a26906a <=( (not A267)  and  a26905a );
 a26910a <=( (not A302)  and  (not A301) );
 a26911a <=( A300  and  a26910a );
 a26912a <=( a26911a  and  a26906a );
 a26916a <=( A167  and  A168 );
 a26917a <=( (not A170)  and  a26916a );
 a26921a <=( A202  and  (not A201) );
 a26922a <=( (not A166)  and  a26921a );
 a26923a <=( a26922a  and  a26917a );
 a26927a <=( A298  and  A268 );
 a26928a <=( (not A267)  and  a26927a );
 a26932a <=( A301  and  A300 );
 a26933a <=( (not A299)  and  a26932a );
 a26934a <=( a26933a  and  a26928a );
 a26938a <=( A167  and  A168 );
 a26939a <=( (not A170)  and  a26938a );
 a26943a <=( A202  and  (not A201) );
 a26944a <=( (not A166)  and  a26943a );
 a26945a <=( a26944a  and  a26939a );
 a26949a <=( A298  and  A268 );
 a26950a <=( (not A267)  and  a26949a );
 a26954a <=( A302  and  A300 );
 a26955a <=( (not A299)  and  a26954a );
 a26956a <=( a26955a  and  a26950a );
 a26960a <=( A167  and  A168 );
 a26961a <=( (not A170)  and  a26960a );
 a26965a <=( A202  and  (not A201) );
 a26966a <=( (not A166)  and  a26965a );
 a26967a <=( a26966a  and  a26961a );
 a26971a <=( (not A298)  and  A268 );
 a26972a <=( (not A267)  and  a26971a );
 a26976a <=( A301  and  A300 );
 a26977a <=( A299  and  a26976a );
 a26978a <=( a26977a  and  a26972a );
 a26982a <=( A167  and  A168 );
 a26983a <=( (not A170)  and  a26982a );
 a26987a <=( A202  and  (not A201) );
 a26988a <=( (not A166)  and  a26987a );
 a26989a <=( a26988a  and  a26983a );
 a26993a <=( (not A298)  and  A268 );
 a26994a <=( (not A267)  and  a26993a );
 a26998a <=( A302  and  A300 );
 a26999a <=( A299  and  a26998a );
 a27000a <=( a26999a  and  a26994a );
 a27004a <=( A167  and  A168 );
 a27005a <=( (not A170)  and  a27004a );
 a27009a <=( A202  and  (not A201) );
 a27010a <=( (not A166)  and  a27009a );
 a27011a <=( a27010a  and  a27005a );
 a27015a <=( A298  and  A269 );
 a27016a <=( (not A267)  and  a27015a );
 a27020a <=( A301  and  A300 );
 a27021a <=( (not A299)  and  a27020a );
 a27022a <=( a27021a  and  a27016a );
 a27026a <=( A167  and  A168 );
 a27027a <=( (not A170)  and  a27026a );
 a27031a <=( A202  and  (not A201) );
 a27032a <=( (not A166)  and  a27031a );
 a27033a <=( a27032a  and  a27027a );
 a27037a <=( A298  and  A269 );
 a27038a <=( (not A267)  and  a27037a );
 a27042a <=( A302  and  A300 );
 a27043a <=( (not A299)  and  a27042a );
 a27044a <=( a27043a  and  a27038a );
 a27048a <=( A167  and  A168 );
 a27049a <=( (not A170)  and  a27048a );
 a27053a <=( A202  and  (not A201) );
 a27054a <=( (not A166)  and  a27053a );
 a27055a <=( a27054a  and  a27049a );
 a27059a <=( (not A298)  and  A269 );
 a27060a <=( (not A267)  and  a27059a );
 a27064a <=( A301  and  A300 );
 a27065a <=( A299  and  a27064a );
 a27066a <=( a27065a  and  a27060a );
 a27070a <=( A167  and  A168 );
 a27071a <=( (not A170)  and  a27070a );
 a27075a <=( A202  and  (not A201) );
 a27076a <=( (not A166)  and  a27075a );
 a27077a <=( a27076a  and  a27071a );
 a27081a <=( (not A298)  and  A269 );
 a27082a <=( (not A267)  and  a27081a );
 a27086a <=( A302  and  A300 );
 a27087a <=( A299  and  a27086a );
 a27088a <=( a27087a  and  a27082a );
 a27092a <=( A167  and  A168 );
 a27093a <=( (not A170)  and  a27092a );
 a27097a <=( A202  and  (not A201) );
 a27098a <=( (not A166)  and  a27097a );
 a27099a <=( a27098a  and  a27093a );
 a27103a <=( A298  and  A266 );
 a27104a <=( A265  and  a27103a );
 a27108a <=( A301  and  A300 );
 a27109a <=( (not A299)  and  a27108a );
 a27110a <=( a27109a  and  a27104a );
 a27114a <=( A167  and  A168 );
 a27115a <=( (not A170)  and  a27114a );
 a27119a <=( A202  and  (not A201) );
 a27120a <=( (not A166)  and  a27119a );
 a27121a <=( a27120a  and  a27115a );
 a27125a <=( A298  and  A266 );
 a27126a <=( A265  and  a27125a );
 a27130a <=( A302  and  A300 );
 a27131a <=( (not A299)  and  a27130a );
 a27132a <=( a27131a  and  a27126a );
 a27136a <=( A167  and  A168 );
 a27137a <=( (not A170)  and  a27136a );
 a27141a <=( A202  and  (not A201) );
 a27142a <=( (not A166)  and  a27141a );
 a27143a <=( a27142a  and  a27137a );
 a27147a <=( (not A298)  and  A266 );
 a27148a <=( A265  and  a27147a );
 a27152a <=( A301  and  A300 );
 a27153a <=( A299  and  a27152a );
 a27154a <=( a27153a  and  a27148a );
 a27158a <=( A167  and  A168 );
 a27159a <=( (not A170)  and  a27158a );
 a27163a <=( A202  and  (not A201) );
 a27164a <=( (not A166)  and  a27163a );
 a27165a <=( a27164a  and  a27159a );
 a27169a <=( (not A298)  and  A266 );
 a27170a <=( A265  and  a27169a );
 a27174a <=( A302  and  A300 );
 a27175a <=( A299  and  a27174a );
 a27176a <=( a27175a  and  a27170a );
 a27180a <=( A167  and  A168 );
 a27181a <=( (not A170)  and  a27180a );
 a27185a <=( A202  and  (not A201) );
 a27186a <=( (not A166)  and  a27185a );
 a27187a <=( a27186a  and  a27181a );
 a27191a <=( A298  and  (not A266) );
 a27192a <=( (not A265)  and  a27191a );
 a27196a <=( A301  and  A300 );
 a27197a <=( (not A299)  and  a27196a );
 a27198a <=( a27197a  and  a27192a );
 a27202a <=( A167  and  A168 );
 a27203a <=( (not A170)  and  a27202a );
 a27207a <=( A202  and  (not A201) );
 a27208a <=( (not A166)  and  a27207a );
 a27209a <=( a27208a  and  a27203a );
 a27213a <=( A298  and  (not A266) );
 a27214a <=( (not A265)  and  a27213a );
 a27218a <=( A302  and  A300 );
 a27219a <=( (not A299)  and  a27218a );
 a27220a <=( a27219a  and  a27214a );
 a27224a <=( A167  and  A168 );
 a27225a <=( (not A170)  and  a27224a );
 a27229a <=( A202  and  (not A201) );
 a27230a <=( (not A166)  and  a27229a );
 a27231a <=( a27230a  and  a27225a );
 a27235a <=( (not A298)  and  (not A266) );
 a27236a <=( (not A265)  and  a27235a );
 a27240a <=( A301  and  A300 );
 a27241a <=( A299  and  a27240a );
 a27242a <=( a27241a  and  a27236a );
 a27246a <=( A167  and  A168 );
 a27247a <=( (not A170)  and  a27246a );
 a27251a <=( A202  and  (not A201) );
 a27252a <=( (not A166)  and  a27251a );
 a27253a <=( a27252a  and  a27247a );
 a27257a <=( (not A298)  and  (not A266) );
 a27258a <=( (not A265)  and  a27257a );
 a27262a <=( A302  and  A300 );
 a27263a <=( A299  and  a27262a );
 a27264a <=( a27263a  and  a27258a );
 a27268a <=( A167  and  A168 );
 a27269a <=( (not A170)  and  a27268a );
 a27273a <=( A203  and  (not A201) );
 a27274a <=( (not A166)  and  a27273a );
 a27275a <=( a27274a  and  a27269a );
 a27279a <=( A298  and  A268 );
 a27280a <=( (not A267)  and  a27279a );
 a27284a <=( A301  and  A300 );
 a27285a <=( (not A299)  and  a27284a );
 a27286a <=( a27285a  and  a27280a );
 a27290a <=( A167  and  A168 );
 a27291a <=( (not A170)  and  a27290a );
 a27295a <=( A203  and  (not A201) );
 a27296a <=( (not A166)  and  a27295a );
 a27297a <=( a27296a  and  a27291a );
 a27301a <=( A298  and  A268 );
 a27302a <=( (not A267)  and  a27301a );
 a27306a <=( A302  and  A300 );
 a27307a <=( (not A299)  and  a27306a );
 a27308a <=( a27307a  and  a27302a );
 a27312a <=( A167  and  A168 );
 a27313a <=( (not A170)  and  a27312a );
 a27317a <=( A203  and  (not A201) );
 a27318a <=( (not A166)  and  a27317a );
 a27319a <=( a27318a  and  a27313a );
 a27323a <=( (not A298)  and  A268 );
 a27324a <=( (not A267)  and  a27323a );
 a27328a <=( A301  and  A300 );
 a27329a <=( A299  and  a27328a );
 a27330a <=( a27329a  and  a27324a );
 a27334a <=( A167  and  A168 );
 a27335a <=( (not A170)  and  a27334a );
 a27339a <=( A203  and  (not A201) );
 a27340a <=( (not A166)  and  a27339a );
 a27341a <=( a27340a  and  a27335a );
 a27345a <=( (not A298)  and  A268 );
 a27346a <=( (not A267)  and  a27345a );
 a27350a <=( A302  and  A300 );
 a27351a <=( A299  and  a27350a );
 a27352a <=( a27351a  and  a27346a );
 a27356a <=( A167  and  A168 );
 a27357a <=( (not A170)  and  a27356a );
 a27361a <=( A203  and  (not A201) );
 a27362a <=( (not A166)  and  a27361a );
 a27363a <=( a27362a  and  a27357a );
 a27367a <=( A298  and  A269 );
 a27368a <=( (not A267)  and  a27367a );
 a27372a <=( A301  and  A300 );
 a27373a <=( (not A299)  and  a27372a );
 a27374a <=( a27373a  and  a27368a );
 a27378a <=( A167  and  A168 );
 a27379a <=( (not A170)  and  a27378a );
 a27383a <=( A203  and  (not A201) );
 a27384a <=( (not A166)  and  a27383a );
 a27385a <=( a27384a  and  a27379a );
 a27389a <=( A298  and  A269 );
 a27390a <=( (not A267)  and  a27389a );
 a27394a <=( A302  and  A300 );
 a27395a <=( (not A299)  and  a27394a );
 a27396a <=( a27395a  and  a27390a );
 a27400a <=( A167  and  A168 );
 a27401a <=( (not A170)  and  a27400a );
 a27405a <=( A203  and  (not A201) );
 a27406a <=( (not A166)  and  a27405a );
 a27407a <=( a27406a  and  a27401a );
 a27411a <=( (not A298)  and  A269 );
 a27412a <=( (not A267)  and  a27411a );
 a27416a <=( A301  and  A300 );
 a27417a <=( A299  and  a27416a );
 a27418a <=( a27417a  and  a27412a );
 a27422a <=( A167  and  A168 );
 a27423a <=( (not A170)  and  a27422a );
 a27427a <=( A203  and  (not A201) );
 a27428a <=( (not A166)  and  a27427a );
 a27429a <=( a27428a  and  a27423a );
 a27433a <=( (not A298)  and  A269 );
 a27434a <=( (not A267)  and  a27433a );
 a27438a <=( A302  and  A300 );
 a27439a <=( A299  and  a27438a );
 a27440a <=( a27439a  and  a27434a );
 a27444a <=( A167  and  A168 );
 a27445a <=( (not A170)  and  a27444a );
 a27449a <=( A203  and  (not A201) );
 a27450a <=( (not A166)  and  a27449a );
 a27451a <=( a27450a  and  a27445a );
 a27455a <=( A298  and  A266 );
 a27456a <=( A265  and  a27455a );
 a27460a <=( A301  and  A300 );
 a27461a <=( (not A299)  and  a27460a );
 a27462a <=( a27461a  and  a27456a );
 a27466a <=( A167  and  A168 );
 a27467a <=( (not A170)  and  a27466a );
 a27471a <=( A203  and  (not A201) );
 a27472a <=( (not A166)  and  a27471a );
 a27473a <=( a27472a  and  a27467a );
 a27477a <=( A298  and  A266 );
 a27478a <=( A265  and  a27477a );
 a27482a <=( A302  and  A300 );
 a27483a <=( (not A299)  and  a27482a );
 a27484a <=( a27483a  and  a27478a );
 a27488a <=( A167  and  A168 );
 a27489a <=( (not A170)  and  a27488a );
 a27493a <=( A203  and  (not A201) );
 a27494a <=( (not A166)  and  a27493a );
 a27495a <=( a27494a  and  a27489a );
 a27499a <=( (not A298)  and  A266 );
 a27500a <=( A265  and  a27499a );
 a27504a <=( A301  and  A300 );
 a27505a <=( A299  and  a27504a );
 a27506a <=( a27505a  and  a27500a );
 a27510a <=( A167  and  A168 );
 a27511a <=( (not A170)  and  a27510a );
 a27515a <=( A203  and  (not A201) );
 a27516a <=( (not A166)  and  a27515a );
 a27517a <=( a27516a  and  a27511a );
 a27521a <=( (not A298)  and  A266 );
 a27522a <=( A265  and  a27521a );
 a27526a <=( A302  and  A300 );
 a27527a <=( A299  and  a27526a );
 a27528a <=( a27527a  and  a27522a );
 a27532a <=( A167  and  A168 );
 a27533a <=( (not A170)  and  a27532a );
 a27537a <=( A203  and  (not A201) );
 a27538a <=( (not A166)  and  a27537a );
 a27539a <=( a27538a  and  a27533a );
 a27543a <=( A298  and  (not A266) );
 a27544a <=( (not A265)  and  a27543a );
 a27548a <=( A301  and  A300 );
 a27549a <=( (not A299)  and  a27548a );
 a27550a <=( a27549a  and  a27544a );
 a27554a <=( A167  and  A168 );
 a27555a <=( (not A170)  and  a27554a );
 a27559a <=( A203  and  (not A201) );
 a27560a <=( (not A166)  and  a27559a );
 a27561a <=( a27560a  and  a27555a );
 a27565a <=( A298  and  (not A266) );
 a27566a <=( (not A265)  and  a27565a );
 a27570a <=( A302  and  A300 );
 a27571a <=( (not A299)  and  a27570a );
 a27572a <=( a27571a  and  a27566a );
 a27576a <=( A167  and  A168 );
 a27577a <=( (not A170)  and  a27576a );
 a27581a <=( A203  and  (not A201) );
 a27582a <=( (not A166)  and  a27581a );
 a27583a <=( a27582a  and  a27577a );
 a27587a <=( (not A298)  and  (not A266) );
 a27588a <=( (not A265)  and  a27587a );
 a27592a <=( A301  and  A300 );
 a27593a <=( A299  and  a27592a );
 a27594a <=( a27593a  and  a27588a );
 a27598a <=( A167  and  A168 );
 a27599a <=( (not A170)  and  a27598a );
 a27603a <=( A203  and  (not A201) );
 a27604a <=( (not A166)  and  a27603a );
 a27605a <=( a27604a  and  a27599a );
 a27609a <=( (not A298)  and  (not A266) );
 a27610a <=( (not A265)  and  a27609a );
 a27614a <=( A302  and  A300 );
 a27615a <=( A299  and  a27614a );
 a27616a <=( a27615a  and  a27610a );
 a27620a <=( A167  and  A168 );
 a27621a <=( (not A170)  and  a27620a );
 a27625a <=( A200  and  A199 );
 a27626a <=( (not A166)  and  a27625a );
 a27627a <=( a27626a  and  a27621a );
 a27631a <=( A298  and  A268 );
 a27632a <=( (not A267)  and  a27631a );
 a27636a <=( A301  and  A300 );
 a27637a <=( (not A299)  and  a27636a );
 a27638a <=( a27637a  and  a27632a );
 a27642a <=( A167  and  A168 );
 a27643a <=( (not A170)  and  a27642a );
 a27647a <=( A200  and  A199 );
 a27648a <=( (not A166)  and  a27647a );
 a27649a <=( a27648a  and  a27643a );
 a27653a <=( A298  and  A268 );
 a27654a <=( (not A267)  and  a27653a );
 a27658a <=( A302  and  A300 );
 a27659a <=( (not A299)  and  a27658a );
 a27660a <=( a27659a  and  a27654a );
 a27664a <=( A167  and  A168 );
 a27665a <=( (not A170)  and  a27664a );
 a27669a <=( A200  and  A199 );
 a27670a <=( (not A166)  and  a27669a );
 a27671a <=( a27670a  and  a27665a );
 a27675a <=( (not A298)  and  A268 );
 a27676a <=( (not A267)  and  a27675a );
 a27680a <=( A301  and  A300 );
 a27681a <=( A299  and  a27680a );
 a27682a <=( a27681a  and  a27676a );
 a27686a <=( A167  and  A168 );
 a27687a <=( (not A170)  and  a27686a );
 a27691a <=( A200  and  A199 );
 a27692a <=( (not A166)  and  a27691a );
 a27693a <=( a27692a  and  a27687a );
 a27697a <=( (not A298)  and  A268 );
 a27698a <=( (not A267)  and  a27697a );
 a27702a <=( A302  and  A300 );
 a27703a <=( A299  and  a27702a );
 a27704a <=( a27703a  and  a27698a );
 a27708a <=( A167  and  A168 );
 a27709a <=( (not A170)  and  a27708a );
 a27713a <=( A200  and  A199 );
 a27714a <=( (not A166)  and  a27713a );
 a27715a <=( a27714a  and  a27709a );
 a27719a <=( A298  and  A269 );
 a27720a <=( (not A267)  and  a27719a );
 a27724a <=( A301  and  A300 );
 a27725a <=( (not A299)  and  a27724a );
 a27726a <=( a27725a  and  a27720a );
 a27730a <=( A167  and  A168 );
 a27731a <=( (not A170)  and  a27730a );
 a27735a <=( A200  and  A199 );
 a27736a <=( (not A166)  and  a27735a );
 a27737a <=( a27736a  and  a27731a );
 a27741a <=( A298  and  A269 );
 a27742a <=( (not A267)  and  a27741a );
 a27746a <=( A302  and  A300 );
 a27747a <=( (not A299)  and  a27746a );
 a27748a <=( a27747a  and  a27742a );
 a27752a <=( A167  and  A168 );
 a27753a <=( (not A170)  and  a27752a );
 a27757a <=( A200  and  A199 );
 a27758a <=( (not A166)  and  a27757a );
 a27759a <=( a27758a  and  a27753a );
 a27763a <=( (not A298)  and  A269 );
 a27764a <=( (not A267)  and  a27763a );
 a27768a <=( A301  and  A300 );
 a27769a <=( A299  and  a27768a );
 a27770a <=( a27769a  and  a27764a );
 a27774a <=( A167  and  A168 );
 a27775a <=( (not A170)  and  a27774a );
 a27779a <=( A200  and  A199 );
 a27780a <=( (not A166)  and  a27779a );
 a27781a <=( a27780a  and  a27775a );
 a27785a <=( (not A298)  and  A269 );
 a27786a <=( (not A267)  and  a27785a );
 a27790a <=( A302  and  A300 );
 a27791a <=( A299  and  a27790a );
 a27792a <=( a27791a  and  a27786a );
 a27796a <=( A167  and  A168 );
 a27797a <=( (not A170)  and  a27796a );
 a27801a <=( A200  and  A199 );
 a27802a <=( (not A166)  and  a27801a );
 a27803a <=( a27802a  and  a27797a );
 a27807a <=( A298  and  A266 );
 a27808a <=( A265  and  a27807a );
 a27812a <=( A301  and  A300 );
 a27813a <=( (not A299)  and  a27812a );
 a27814a <=( a27813a  and  a27808a );
 a27818a <=( A167  and  A168 );
 a27819a <=( (not A170)  and  a27818a );
 a27823a <=( A200  and  A199 );
 a27824a <=( (not A166)  and  a27823a );
 a27825a <=( a27824a  and  a27819a );
 a27829a <=( A298  and  A266 );
 a27830a <=( A265  and  a27829a );
 a27834a <=( A302  and  A300 );
 a27835a <=( (not A299)  and  a27834a );
 a27836a <=( a27835a  and  a27830a );
 a27840a <=( A167  and  A168 );
 a27841a <=( (not A170)  and  a27840a );
 a27845a <=( A200  and  A199 );
 a27846a <=( (not A166)  and  a27845a );
 a27847a <=( a27846a  and  a27841a );
 a27851a <=( (not A298)  and  A266 );
 a27852a <=( A265  and  a27851a );
 a27856a <=( A301  and  A300 );
 a27857a <=( A299  and  a27856a );
 a27858a <=( a27857a  and  a27852a );
 a27862a <=( A167  and  A168 );
 a27863a <=( (not A170)  and  a27862a );
 a27867a <=( A200  and  A199 );
 a27868a <=( (not A166)  and  a27867a );
 a27869a <=( a27868a  and  a27863a );
 a27873a <=( (not A298)  and  A266 );
 a27874a <=( A265  and  a27873a );
 a27878a <=( A302  and  A300 );
 a27879a <=( A299  and  a27878a );
 a27880a <=( a27879a  and  a27874a );
 a27884a <=( A167  and  A168 );
 a27885a <=( (not A170)  and  a27884a );
 a27889a <=( A200  and  A199 );
 a27890a <=( (not A166)  and  a27889a );
 a27891a <=( a27890a  and  a27885a );
 a27895a <=( A298  and  (not A266) );
 a27896a <=( (not A265)  and  a27895a );
 a27900a <=( A301  and  A300 );
 a27901a <=( (not A299)  and  a27900a );
 a27902a <=( a27901a  and  a27896a );
 a27906a <=( A167  and  A168 );
 a27907a <=( (not A170)  and  a27906a );
 a27911a <=( A200  and  A199 );
 a27912a <=( (not A166)  and  a27911a );
 a27913a <=( a27912a  and  a27907a );
 a27917a <=( A298  and  (not A266) );
 a27918a <=( (not A265)  and  a27917a );
 a27922a <=( A302  and  A300 );
 a27923a <=( (not A299)  and  a27922a );
 a27924a <=( a27923a  and  a27918a );
 a27928a <=( A167  and  A168 );
 a27929a <=( (not A170)  and  a27928a );
 a27933a <=( A200  and  A199 );
 a27934a <=( (not A166)  and  a27933a );
 a27935a <=( a27934a  and  a27929a );
 a27939a <=( (not A298)  and  (not A266) );
 a27940a <=( (not A265)  and  a27939a );
 a27944a <=( A301  and  A300 );
 a27945a <=( A299  and  a27944a );
 a27946a <=( a27945a  and  a27940a );
 a27950a <=( A167  and  A168 );
 a27951a <=( (not A170)  and  a27950a );
 a27955a <=( A200  and  A199 );
 a27956a <=( (not A166)  and  a27955a );
 a27957a <=( a27956a  and  a27951a );
 a27961a <=( (not A298)  and  (not A266) );
 a27962a <=( (not A265)  and  a27961a );
 a27966a <=( A302  and  A300 );
 a27967a <=( A299  and  a27966a );
 a27968a <=( a27967a  and  a27962a );
 a27972a <=( A167  and  A168 );
 a27973a <=( (not A170)  and  a27972a );
 a27977a <=( (not A200)  and  (not A199) );
 a27978a <=( (not A166)  and  a27977a );
 a27979a <=( a27978a  and  a27973a );
 a27983a <=( A298  and  A268 );
 a27984a <=( (not A267)  and  a27983a );
 a27988a <=( A301  and  A300 );
 a27989a <=( (not A299)  and  a27988a );
 a27990a <=( a27989a  and  a27984a );
 a27994a <=( A167  and  A168 );
 a27995a <=( (not A170)  and  a27994a );
 a27999a <=( (not A200)  and  (not A199) );
 a28000a <=( (not A166)  and  a27999a );
 a28001a <=( a28000a  and  a27995a );
 a28005a <=( A298  and  A268 );
 a28006a <=( (not A267)  and  a28005a );
 a28010a <=( A302  and  A300 );
 a28011a <=( (not A299)  and  a28010a );
 a28012a <=( a28011a  and  a28006a );
 a28016a <=( A167  and  A168 );
 a28017a <=( (not A170)  and  a28016a );
 a28021a <=( (not A200)  and  (not A199) );
 a28022a <=( (not A166)  and  a28021a );
 a28023a <=( a28022a  and  a28017a );
 a28027a <=( (not A298)  and  A268 );
 a28028a <=( (not A267)  and  a28027a );
 a28032a <=( A301  and  A300 );
 a28033a <=( A299  and  a28032a );
 a28034a <=( a28033a  and  a28028a );
 a28038a <=( A167  and  A168 );
 a28039a <=( (not A170)  and  a28038a );
 a28043a <=( (not A200)  and  (not A199) );
 a28044a <=( (not A166)  and  a28043a );
 a28045a <=( a28044a  and  a28039a );
 a28049a <=( (not A298)  and  A268 );
 a28050a <=( (not A267)  and  a28049a );
 a28054a <=( A302  and  A300 );
 a28055a <=( A299  and  a28054a );
 a28056a <=( a28055a  and  a28050a );
 a28060a <=( A167  and  A168 );
 a28061a <=( (not A170)  and  a28060a );
 a28065a <=( (not A200)  and  (not A199) );
 a28066a <=( (not A166)  and  a28065a );
 a28067a <=( a28066a  and  a28061a );
 a28071a <=( A298  and  A269 );
 a28072a <=( (not A267)  and  a28071a );
 a28076a <=( A301  and  A300 );
 a28077a <=( (not A299)  and  a28076a );
 a28078a <=( a28077a  and  a28072a );
 a28082a <=( A167  and  A168 );
 a28083a <=( (not A170)  and  a28082a );
 a28087a <=( (not A200)  and  (not A199) );
 a28088a <=( (not A166)  and  a28087a );
 a28089a <=( a28088a  and  a28083a );
 a28093a <=( A298  and  A269 );
 a28094a <=( (not A267)  and  a28093a );
 a28098a <=( A302  and  A300 );
 a28099a <=( (not A299)  and  a28098a );
 a28100a <=( a28099a  and  a28094a );
 a28104a <=( A167  and  A168 );
 a28105a <=( (not A170)  and  a28104a );
 a28109a <=( (not A200)  and  (not A199) );
 a28110a <=( (not A166)  and  a28109a );
 a28111a <=( a28110a  and  a28105a );
 a28115a <=( (not A298)  and  A269 );
 a28116a <=( (not A267)  and  a28115a );
 a28120a <=( A301  and  A300 );
 a28121a <=( A299  and  a28120a );
 a28122a <=( a28121a  and  a28116a );
 a28126a <=( A167  and  A168 );
 a28127a <=( (not A170)  and  a28126a );
 a28131a <=( (not A200)  and  (not A199) );
 a28132a <=( (not A166)  and  a28131a );
 a28133a <=( a28132a  and  a28127a );
 a28137a <=( (not A298)  and  A269 );
 a28138a <=( (not A267)  and  a28137a );
 a28142a <=( A302  and  A300 );
 a28143a <=( A299  and  a28142a );
 a28144a <=( a28143a  and  a28138a );
 a28148a <=( A167  and  A168 );
 a28149a <=( (not A170)  and  a28148a );
 a28153a <=( (not A200)  and  (not A199) );
 a28154a <=( (not A166)  and  a28153a );
 a28155a <=( a28154a  and  a28149a );
 a28159a <=( A298  and  A266 );
 a28160a <=( A265  and  a28159a );
 a28164a <=( A301  and  A300 );
 a28165a <=( (not A299)  and  a28164a );
 a28166a <=( a28165a  and  a28160a );
 a28170a <=( A167  and  A168 );
 a28171a <=( (not A170)  and  a28170a );
 a28175a <=( (not A200)  and  (not A199) );
 a28176a <=( (not A166)  and  a28175a );
 a28177a <=( a28176a  and  a28171a );
 a28181a <=( A298  and  A266 );
 a28182a <=( A265  and  a28181a );
 a28186a <=( A302  and  A300 );
 a28187a <=( (not A299)  and  a28186a );
 a28188a <=( a28187a  and  a28182a );
 a28192a <=( A167  and  A168 );
 a28193a <=( (not A170)  and  a28192a );
 a28197a <=( (not A200)  and  (not A199) );
 a28198a <=( (not A166)  and  a28197a );
 a28199a <=( a28198a  and  a28193a );
 a28203a <=( (not A298)  and  A266 );
 a28204a <=( A265  and  a28203a );
 a28208a <=( A301  and  A300 );
 a28209a <=( A299  and  a28208a );
 a28210a <=( a28209a  and  a28204a );
 a28214a <=( A167  and  A168 );
 a28215a <=( (not A170)  and  a28214a );
 a28219a <=( (not A200)  and  (not A199) );
 a28220a <=( (not A166)  and  a28219a );
 a28221a <=( a28220a  and  a28215a );
 a28225a <=( (not A298)  and  A266 );
 a28226a <=( A265  and  a28225a );
 a28230a <=( A302  and  A300 );
 a28231a <=( A299  and  a28230a );
 a28232a <=( a28231a  and  a28226a );
 a28236a <=( A167  and  A168 );
 a28237a <=( (not A170)  and  a28236a );
 a28241a <=( (not A200)  and  (not A199) );
 a28242a <=( (not A166)  and  a28241a );
 a28243a <=( a28242a  and  a28237a );
 a28247a <=( A298  and  (not A266) );
 a28248a <=( (not A265)  and  a28247a );
 a28252a <=( A301  and  A300 );
 a28253a <=( (not A299)  and  a28252a );
 a28254a <=( a28253a  and  a28248a );
 a28258a <=( A167  and  A168 );
 a28259a <=( (not A170)  and  a28258a );
 a28263a <=( (not A200)  and  (not A199) );
 a28264a <=( (not A166)  and  a28263a );
 a28265a <=( a28264a  and  a28259a );
 a28269a <=( A298  and  (not A266) );
 a28270a <=( (not A265)  and  a28269a );
 a28274a <=( A302  and  A300 );
 a28275a <=( (not A299)  and  a28274a );
 a28276a <=( a28275a  and  a28270a );
 a28280a <=( A167  and  A168 );
 a28281a <=( (not A170)  and  a28280a );
 a28285a <=( (not A200)  and  (not A199) );
 a28286a <=( (not A166)  and  a28285a );
 a28287a <=( a28286a  and  a28281a );
 a28291a <=( (not A298)  and  (not A266) );
 a28292a <=( (not A265)  and  a28291a );
 a28296a <=( A301  and  A300 );
 a28297a <=( A299  and  a28296a );
 a28298a <=( a28297a  and  a28292a );
 a28302a <=( A167  and  A168 );
 a28303a <=( (not A170)  and  a28302a );
 a28307a <=( (not A200)  and  (not A199) );
 a28308a <=( (not A166)  and  a28307a );
 a28309a <=( a28308a  and  a28303a );
 a28313a <=( (not A298)  and  (not A266) );
 a28314a <=( (not A265)  and  a28313a );
 a28318a <=( A302  and  A300 );
 a28319a <=( A299  and  a28318a );
 a28320a <=( a28319a  and  a28314a );
 a28324a <=( (not A167)  and  A168 );
 a28325a <=( (not A170)  and  a28324a );
 a28329a <=( A202  and  (not A201) );
 a28330a <=( A166  and  a28329a );
 a28331a <=( a28330a  and  a28325a );
 a28335a <=( A298  and  A268 );
 a28336a <=( (not A267)  and  a28335a );
 a28340a <=( A301  and  A300 );
 a28341a <=( (not A299)  and  a28340a );
 a28342a <=( a28341a  and  a28336a );
 a28346a <=( (not A167)  and  A168 );
 a28347a <=( (not A170)  and  a28346a );
 a28351a <=( A202  and  (not A201) );
 a28352a <=( A166  and  a28351a );
 a28353a <=( a28352a  and  a28347a );
 a28357a <=( A298  and  A268 );
 a28358a <=( (not A267)  and  a28357a );
 a28362a <=( A302  and  A300 );
 a28363a <=( (not A299)  and  a28362a );
 a28364a <=( a28363a  and  a28358a );
 a28368a <=( (not A167)  and  A168 );
 a28369a <=( (not A170)  and  a28368a );
 a28373a <=( A202  and  (not A201) );
 a28374a <=( A166  and  a28373a );
 a28375a <=( a28374a  and  a28369a );
 a28379a <=( (not A298)  and  A268 );
 a28380a <=( (not A267)  and  a28379a );
 a28384a <=( A301  and  A300 );
 a28385a <=( A299  and  a28384a );
 a28386a <=( a28385a  and  a28380a );
 a28390a <=( (not A167)  and  A168 );
 a28391a <=( (not A170)  and  a28390a );
 a28395a <=( A202  and  (not A201) );
 a28396a <=( A166  and  a28395a );
 a28397a <=( a28396a  and  a28391a );
 a28401a <=( (not A298)  and  A268 );
 a28402a <=( (not A267)  and  a28401a );
 a28406a <=( A302  and  A300 );
 a28407a <=( A299  and  a28406a );
 a28408a <=( a28407a  and  a28402a );
 a28412a <=( (not A167)  and  A168 );
 a28413a <=( (not A170)  and  a28412a );
 a28417a <=( A202  and  (not A201) );
 a28418a <=( A166  and  a28417a );
 a28419a <=( a28418a  and  a28413a );
 a28423a <=( A298  and  A269 );
 a28424a <=( (not A267)  and  a28423a );
 a28428a <=( A301  and  A300 );
 a28429a <=( (not A299)  and  a28428a );
 a28430a <=( a28429a  and  a28424a );
 a28434a <=( (not A167)  and  A168 );
 a28435a <=( (not A170)  and  a28434a );
 a28439a <=( A202  and  (not A201) );
 a28440a <=( A166  and  a28439a );
 a28441a <=( a28440a  and  a28435a );
 a28445a <=( A298  and  A269 );
 a28446a <=( (not A267)  and  a28445a );
 a28450a <=( A302  and  A300 );
 a28451a <=( (not A299)  and  a28450a );
 a28452a <=( a28451a  and  a28446a );
 a28456a <=( (not A167)  and  A168 );
 a28457a <=( (not A170)  and  a28456a );
 a28461a <=( A202  and  (not A201) );
 a28462a <=( A166  and  a28461a );
 a28463a <=( a28462a  and  a28457a );
 a28467a <=( (not A298)  and  A269 );
 a28468a <=( (not A267)  and  a28467a );
 a28472a <=( A301  and  A300 );
 a28473a <=( A299  and  a28472a );
 a28474a <=( a28473a  and  a28468a );
 a28478a <=( (not A167)  and  A168 );
 a28479a <=( (not A170)  and  a28478a );
 a28483a <=( A202  and  (not A201) );
 a28484a <=( A166  and  a28483a );
 a28485a <=( a28484a  and  a28479a );
 a28489a <=( (not A298)  and  A269 );
 a28490a <=( (not A267)  and  a28489a );
 a28494a <=( A302  and  A300 );
 a28495a <=( A299  and  a28494a );
 a28496a <=( a28495a  and  a28490a );
 a28500a <=( (not A167)  and  A168 );
 a28501a <=( (not A170)  and  a28500a );
 a28505a <=( A202  and  (not A201) );
 a28506a <=( A166  and  a28505a );
 a28507a <=( a28506a  and  a28501a );
 a28511a <=( A298  and  A266 );
 a28512a <=( A265  and  a28511a );
 a28516a <=( A301  and  A300 );
 a28517a <=( (not A299)  and  a28516a );
 a28518a <=( a28517a  and  a28512a );
 a28522a <=( (not A167)  and  A168 );
 a28523a <=( (not A170)  and  a28522a );
 a28527a <=( A202  and  (not A201) );
 a28528a <=( A166  and  a28527a );
 a28529a <=( a28528a  and  a28523a );
 a28533a <=( A298  and  A266 );
 a28534a <=( A265  and  a28533a );
 a28538a <=( A302  and  A300 );
 a28539a <=( (not A299)  and  a28538a );
 a28540a <=( a28539a  and  a28534a );
 a28544a <=( (not A167)  and  A168 );
 a28545a <=( (not A170)  and  a28544a );
 a28549a <=( A202  and  (not A201) );
 a28550a <=( A166  and  a28549a );
 a28551a <=( a28550a  and  a28545a );
 a28555a <=( (not A298)  and  A266 );
 a28556a <=( A265  and  a28555a );
 a28560a <=( A301  and  A300 );
 a28561a <=( A299  and  a28560a );
 a28562a <=( a28561a  and  a28556a );
 a28566a <=( (not A167)  and  A168 );
 a28567a <=( (not A170)  and  a28566a );
 a28571a <=( A202  and  (not A201) );
 a28572a <=( A166  and  a28571a );
 a28573a <=( a28572a  and  a28567a );
 a28577a <=( (not A298)  and  A266 );
 a28578a <=( A265  and  a28577a );
 a28582a <=( A302  and  A300 );
 a28583a <=( A299  and  a28582a );
 a28584a <=( a28583a  and  a28578a );
 a28588a <=( (not A167)  and  A168 );
 a28589a <=( (not A170)  and  a28588a );
 a28593a <=( A202  and  (not A201) );
 a28594a <=( A166  and  a28593a );
 a28595a <=( a28594a  and  a28589a );
 a28599a <=( A298  and  (not A266) );
 a28600a <=( (not A265)  and  a28599a );
 a28604a <=( A301  and  A300 );
 a28605a <=( (not A299)  and  a28604a );
 a28606a <=( a28605a  and  a28600a );
 a28610a <=( (not A167)  and  A168 );
 a28611a <=( (not A170)  and  a28610a );
 a28615a <=( A202  and  (not A201) );
 a28616a <=( A166  and  a28615a );
 a28617a <=( a28616a  and  a28611a );
 a28621a <=( A298  and  (not A266) );
 a28622a <=( (not A265)  and  a28621a );
 a28626a <=( A302  and  A300 );
 a28627a <=( (not A299)  and  a28626a );
 a28628a <=( a28627a  and  a28622a );
 a28632a <=( (not A167)  and  A168 );
 a28633a <=( (not A170)  and  a28632a );
 a28637a <=( A202  and  (not A201) );
 a28638a <=( A166  and  a28637a );
 a28639a <=( a28638a  and  a28633a );
 a28643a <=( (not A298)  and  (not A266) );
 a28644a <=( (not A265)  and  a28643a );
 a28648a <=( A301  and  A300 );
 a28649a <=( A299  and  a28648a );
 a28650a <=( a28649a  and  a28644a );
 a28654a <=( (not A167)  and  A168 );
 a28655a <=( (not A170)  and  a28654a );
 a28659a <=( A202  and  (not A201) );
 a28660a <=( A166  and  a28659a );
 a28661a <=( a28660a  and  a28655a );
 a28665a <=( (not A298)  and  (not A266) );
 a28666a <=( (not A265)  and  a28665a );
 a28670a <=( A302  and  A300 );
 a28671a <=( A299  and  a28670a );
 a28672a <=( a28671a  and  a28666a );
 a28676a <=( (not A167)  and  A168 );
 a28677a <=( (not A170)  and  a28676a );
 a28681a <=( A203  and  (not A201) );
 a28682a <=( A166  and  a28681a );
 a28683a <=( a28682a  and  a28677a );
 a28687a <=( A298  and  A268 );
 a28688a <=( (not A267)  and  a28687a );
 a28692a <=( A301  and  A300 );
 a28693a <=( (not A299)  and  a28692a );
 a28694a <=( a28693a  and  a28688a );
 a28698a <=( (not A167)  and  A168 );
 a28699a <=( (not A170)  and  a28698a );
 a28703a <=( A203  and  (not A201) );
 a28704a <=( A166  and  a28703a );
 a28705a <=( a28704a  and  a28699a );
 a28709a <=( A298  and  A268 );
 a28710a <=( (not A267)  and  a28709a );
 a28714a <=( A302  and  A300 );
 a28715a <=( (not A299)  and  a28714a );
 a28716a <=( a28715a  and  a28710a );
 a28720a <=( (not A167)  and  A168 );
 a28721a <=( (not A170)  and  a28720a );
 a28725a <=( A203  and  (not A201) );
 a28726a <=( A166  and  a28725a );
 a28727a <=( a28726a  and  a28721a );
 a28731a <=( (not A298)  and  A268 );
 a28732a <=( (not A267)  and  a28731a );
 a28736a <=( A301  and  A300 );
 a28737a <=( A299  and  a28736a );
 a28738a <=( a28737a  and  a28732a );
 a28742a <=( (not A167)  and  A168 );
 a28743a <=( (not A170)  and  a28742a );
 a28747a <=( A203  and  (not A201) );
 a28748a <=( A166  and  a28747a );
 a28749a <=( a28748a  and  a28743a );
 a28753a <=( (not A298)  and  A268 );
 a28754a <=( (not A267)  and  a28753a );
 a28758a <=( A302  and  A300 );
 a28759a <=( A299  and  a28758a );
 a28760a <=( a28759a  and  a28754a );
 a28764a <=( (not A167)  and  A168 );
 a28765a <=( (not A170)  and  a28764a );
 a28769a <=( A203  and  (not A201) );
 a28770a <=( A166  and  a28769a );
 a28771a <=( a28770a  and  a28765a );
 a28775a <=( A298  and  A269 );
 a28776a <=( (not A267)  and  a28775a );
 a28780a <=( A301  and  A300 );
 a28781a <=( (not A299)  and  a28780a );
 a28782a <=( a28781a  and  a28776a );
 a28786a <=( (not A167)  and  A168 );
 a28787a <=( (not A170)  and  a28786a );
 a28791a <=( A203  and  (not A201) );
 a28792a <=( A166  and  a28791a );
 a28793a <=( a28792a  and  a28787a );
 a28797a <=( A298  and  A269 );
 a28798a <=( (not A267)  and  a28797a );
 a28802a <=( A302  and  A300 );
 a28803a <=( (not A299)  and  a28802a );
 a28804a <=( a28803a  and  a28798a );
 a28808a <=( (not A167)  and  A168 );
 a28809a <=( (not A170)  and  a28808a );
 a28813a <=( A203  and  (not A201) );
 a28814a <=( A166  and  a28813a );
 a28815a <=( a28814a  and  a28809a );
 a28819a <=( (not A298)  and  A269 );
 a28820a <=( (not A267)  and  a28819a );
 a28824a <=( A301  and  A300 );
 a28825a <=( A299  and  a28824a );
 a28826a <=( a28825a  and  a28820a );
 a28830a <=( (not A167)  and  A168 );
 a28831a <=( (not A170)  and  a28830a );
 a28835a <=( A203  and  (not A201) );
 a28836a <=( A166  and  a28835a );
 a28837a <=( a28836a  and  a28831a );
 a28841a <=( (not A298)  and  A269 );
 a28842a <=( (not A267)  and  a28841a );
 a28846a <=( A302  and  A300 );
 a28847a <=( A299  and  a28846a );
 a28848a <=( a28847a  and  a28842a );
 a28852a <=( (not A167)  and  A168 );
 a28853a <=( (not A170)  and  a28852a );
 a28857a <=( A203  and  (not A201) );
 a28858a <=( A166  and  a28857a );
 a28859a <=( a28858a  and  a28853a );
 a28863a <=( A298  and  A266 );
 a28864a <=( A265  and  a28863a );
 a28868a <=( A301  and  A300 );
 a28869a <=( (not A299)  and  a28868a );
 a28870a <=( a28869a  and  a28864a );
 a28874a <=( (not A167)  and  A168 );
 a28875a <=( (not A170)  and  a28874a );
 a28879a <=( A203  and  (not A201) );
 a28880a <=( A166  and  a28879a );
 a28881a <=( a28880a  and  a28875a );
 a28885a <=( A298  and  A266 );
 a28886a <=( A265  and  a28885a );
 a28890a <=( A302  and  A300 );
 a28891a <=( (not A299)  and  a28890a );
 a28892a <=( a28891a  and  a28886a );
 a28896a <=( (not A167)  and  A168 );
 a28897a <=( (not A170)  and  a28896a );
 a28901a <=( A203  and  (not A201) );
 a28902a <=( A166  and  a28901a );
 a28903a <=( a28902a  and  a28897a );
 a28907a <=( (not A298)  and  A266 );
 a28908a <=( A265  and  a28907a );
 a28912a <=( A301  and  A300 );
 a28913a <=( A299  and  a28912a );
 a28914a <=( a28913a  and  a28908a );
 a28918a <=( (not A167)  and  A168 );
 a28919a <=( (not A170)  and  a28918a );
 a28923a <=( A203  and  (not A201) );
 a28924a <=( A166  and  a28923a );
 a28925a <=( a28924a  and  a28919a );
 a28929a <=( (not A298)  and  A266 );
 a28930a <=( A265  and  a28929a );
 a28934a <=( A302  and  A300 );
 a28935a <=( A299  and  a28934a );
 a28936a <=( a28935a  and  a28930a );
 a28940a <=( (not A167)  and  A168 );
 a28941a <=( (not A170)  and  a28940a );
 a28945a <=( A203  and  (not A201) );
 a28946a <=( A166  and  a28945a );
 a28947a <=( a28946a  and  a28941a );
 a28951a <=( A298  and  (not A266) );
 a28952a <=( (not A265)  and  a28951a );
 a28956a <=( A301  and  A300 );
 a28957a <=( (not A299)  and  a28956a );
 a28958a <=( a28957a  and  a28952a );
 a28962a <=( (not A167)  and  A168 );
 a28963a <=( (not A170)  and  a28962a );
 a28967a <=( A203  and  (not A201) );
 a28968a <=( A166  and  a28967a );
 a28969a <=( a28968a  and  a28963a );
 a28973a <=( A298  and  (not A266) );
 a28974a <=( (not A265)  and  a28973a );
 a28978a <=( A302  and  A300 );
 a28979a <=( (not A299)  and  a28978a );
 a28980a <=( a28979a  and  a28974a );
 a28984a <=( (not A167)  and  A168 );
 a28985a <=( (not A170)  and  a28984a );
 a28989a <=( A203  and  (not A201) );
 a28990a <=( A166  and  a28989a );
 a28991a <=( a28990a  and  a28985a );
 a28995a <=( (not A298)  and  (not A266) );
 a28996a <=( (not A265)  and  a28995a );
 a29000a <=( A301  and  A300 );
 a29001a <=( A299  and  a29000a );
 a29002a <=( a29001a  and  a28996a );
 a29006a <=( (not A167)  and  A168 );
 a29007a <=( (not A170)  and  a29006a );
 a29011a <=( A203  and  (not A201) );
 a29012a <=( A166  and  a29011a );
 a29013a <=( a29012a  and  a29007a );
 a29017a <=( (not A298)  and  (not A266) );
 a29018a <=( (not A265)  and  a29017a );
 a29022a <=( A302  and  A300 );
 a29023a <=( A299  and  a29022a );
 a29024a <=( a29023a  and  a29018a );
 a29028a <=( (not A167)  and  A168 );
 a29029a <=( (not A170)  and  a29028a );
 a29033a <=( A200  and  A199 );
 a29034a <=( A166  and  a29033a );
 a29035a <=( a29034a  and  a29029a );
 a29039a <=( A298  and  A268 );
 a29040a <=( (not A267)  and  a29039a );
 a29044a <=( A301  and  A300 );
 a29045a <=( (not A299)  and  a29044a );
 a29046a <=( a29045a  and  a29040a );
 a29050a <=( (not A167)  and  A168 );
 a29051a <=( (not A170)  and  a29050a );
 a29055a <=( A200  and  A199 );
 a29056a <=( A166  and  a29055a );
 a29057a <=( a29056a  and  a29051a );
 a29061a <=( A298  and  A268 );
 a29062a <=( (not A267)  and  a29061a );
 a29066a <=( A302  and  A300 );
 a29067a <=( (not A299)  and  a29066a );
 a29068a <=( a29067a  and  a29062a );
 a29072a <=( (not A167)  and  A168 );
 a29073a <=( (not A170)  and  a29072a );
 a29077a <=( A200  and  A199 );
 a29078a <=( A166  and  a29077a );
 a29079a <=( a29078a  and  a29073a );
 a29083a <=( (not A298)  and  A268 );
 a29084a <=( (not A267)  and  a29083a );
 a29088a <=( A301  and  A300 );
 a29089a <=( A299  and  a29088a );
 a29090a <=( a29089a  and  a29084a );
 a29094a <=( (not A167)  and  A168 );
 a29095a <=( (not A170)  and  a29094a );
 a29099a <=( A200  and  A199 );
 a29100a <=( A166  and  a29099a );
 a29101a <=( a29100a  and  a29095a );
 a29105a <=( (not A298)  and  A268 );
 a29106a <=( (not A267)  and  a29105a );
 a29110a <=( A302  and  A300 );
 a29111a <=( A299  and  a29110a );
 a29112a <=( a29111a  and  a29106a );
 a29116a <=( (not A167)  and  A168 );
 a29117a <=( (not A170)  and  a29116a );
 a29121a <=( A200  and  A199 );
 a29122a <=( A166  and  a29121a );
 a29123a <=( a29122a  and  a29117a );
 a29127a <=( A298  and  A269 );
 a29128a <=( (not A267)  and  a29127a );
 a29132a <=( A301  and  A300 );
 a29133a <=( (not A299)  and  a29132a );
 a29134a <=( a29133a  and  a29128a );
 a29138a <=( (not A167)  and  A168 );
 a29139a <=( (not A170)  and  a29138a );
 a29143a <=( A200  and  A199 );
 a29144a <=( A166  and  a29143a );
 a29145a <=( a29144a  and  a29139a );
 a29149a <=( A298  and  A269 );
 a29150a <=( (not A267)  and  a29149a );
 a29154a <=( A302  and  A300 );
 a29155a <=( (not A299)  and  a29154a );
 a29156a <=( a29155a  and  a29150a );
 a29160a <=( (not A167)  and  A168 );
 a29161a <=( (not A170)  and  a29160a );
 a29165a <=( A200  and  A199 );
 a29166a <=( A166  and  a29165a );
 a29167a <=( a29166a  and  a29161a );
 a29171a <=( (not A298)  and  A269 );
 a29172a <=( (not A267)  and  a29171a );
 a29176a <=( A301  and  A300 );
 a29177a <=( A299  and  a29176a );
 a29178a <=( a29177a  and  a29172a );
 a29182a <=( (not A167)  and  A168 );
 a29183a <=( (not A170)  and  a29182a );
 a29187a <=( A200  and  A199 );
 a29188a <=( A166  and  a29187a );
 a29189a <=( a29188a  and  a29183a );
 a29193a <=( (not A298)  and  A269 );
 a29194a <=( (not A267)  and  a29193a );
 a29198a <=( A302  and  A300 );
 a29199a <=( A299  and  a29198a );
 a29200a <=( a29199a  and  a29194a );
 a29204a <=( (not A167)  and  A168 );
 a29205a <=( (not A170)  and  a29204a );
 a29209a <=( A200  and  A199 );
 a29210a <=( A166  and  a29209a );
 a29211a <=( a29210a  and  a29205a );
 a29215a <=( A298  and  A266 );
 a29216a <=( A265  and  a29215a );
 a29220a <=( A301  and  A300 );
 a29221a <=( (not A299)  and  a29220a );
 a29222a <=( a29221a  and  a29216a );
 a29226a <=( (not A167)  and  A168 );
 a29227a <=( (not A170)  and  a29226a );
 a29231a <=( A200  and  A199 );
 a29232a <=( A166  and  a29231a );
 a29233a <=( a29232a  and  a29227a );
 a29237a <=( A298  and  A266 );
 a29238a <=( A265  and  a29237a );
 a29242a <=( A302  and  A300 );
 a29243a <=( (not A299)  and  a29242a );
 a29244a <=( a29243a  and  a29238a );
 a29248a <=( (not A167)  and  A168 );
 a29249a <=( (not A170)  and  a29248a );
 a29253a <=( A200  and  A199 );
 a29254a <=( A166  and  a29253a );
 a29255a <=( a29254a  and  a29249a );
 a29259a <=( (not A298)  and  A266 );
 a29260a <=( A265  and  a29259a );
 a29264a <=( A301  and  A300 );
 a29265a <=( A299  and  a29264a );
 a29266a <=( a29265a  and  a29260a );
 a29270a <=( (not A167)  and  A168 );
 a29271a <=( (not A170)  and  a29270a );
 a29275a <=( A200  and  A199 );
 a29276a <=( A166  and  a29275a );
 a29277a <=( a29276a  and  a29271a );
 a29281a <=( (not A298)  and  A266 );
 a29282a <=( A265  and  a29281a );
 a29286a <=( A302  and  A300 );
 a29287a <=( A299  and  a29286a );
 a29288a <=( a29287a  and  a29282a );
 a29292a <=( (not A167)  and  A168 );
 a29293a <=( (not A170)  and  a29292a );
 a29297a <=( A200  and  A199 );
 a29298a <=( A166  and  a29297a );
 a29299a <=( a29298a  and  a29293a );
 a29303a <=( A298  and  (not A266) );
 a29304a <=( (not A265)  and  a29303a );
 a29308a <=( A301  and  A300 );
 a29309a <=( (not A299)  and  a29308a );
 a29310a <=( a29309a  and  a29304a );
 a29314a <=( (not A167)  and  A168 );
 a29315a <=( (not A170)  and  a29314a );
 a29319a <=( A200  and  A199 );
 a29320a <=( A166  and  a29319a );
 a29321a <=( a29320a  and  a29315a );
 a29325a <=( A298  and  (not A266) );
 a29326a <=( (not A265)  and  a29325a );
 a29330a <=( A302  and  A300 );
 a29331a <=( (not A299)  and  a29330a );
 a29332a <=( a29331a  and  a29326a );
 a29336a <=( (not A167)  and  A168 );
 a29337a <=( (not A170)  and  a29336a );
 a29341a <=( A200  and  A199 );
 a29342a <=( A166  and  a29341a );
 a29343a <=( a29342a  and  a29337a );
 a29347a <=( (not A298)  and  (not A266) );
 a29348a <=( (not A265)  and  a29347a );
 a29352a <=( A301  and  A300 );
 a29353a <=( A299  and  a29352a );
 a29354a <=( a29353a  and  a29348a );
 a29358a <=( (not A167)  and  A168 );
 a29359a <=( (not A170)  and  a29358a );
 a29363a <=( A200  and  A199 );
 a29364a <=( A166  and  a29363a );
 a29365a <=( a29364a  and  a29359a );
 a29369a <=( (not A298)  and  (not A266) );
 a29370a <=( (not A265)  and  a29369a );
 a29374a <=( A302  and  A300 );
 a29375a <=( A299  and  a29374a );
 a29376a <=( a29375a  and  a29370a );
 a29380a <=( (not A167)  and  A168 );
 a29381a <=( (not A170)  and  a29380a );
 a29385a <=( (not A200)  and  (not A199) );
 a29386a <=( A166  and  a29385a );
 a29387a <=( a29386a  and  a29381a );
 a29391a <=( A298  and  A268 );
 a29392a <=( (not A267)  and  a29391a );
 a29396a <=( A301  and  A300 );
 a29397a <=( (not A299)  and  a29396a );
 a29398a <=( a29397a  and  a29392a );
 a29402a <=( (not A167)  and  A168 );
 a29403a <=( (not A170)  and  a29402a );
 a29407a <=( (not A200)  and  (not A199) );
 a29408a <=( A166  and  a29407a );
 a29409a <=( a29408a  and  a29403a );
 a29413a <=( A298  and  A268 );
 a29414a <=( (not A267)  and  a29413a );
 a29418a <=( A302  and  A300 );
 a29419a <=( (not A299)  and  a29418a );
 a29420a <=( a29419a  and  a29414a );
 a29424a <=( (not A167)  and  A168 );
 a29425a <=( (not A170)  and  a29424a );
 a29429a <=( (not A200)  and  (not A199) );
 a29430a <=( A166  and  a29429a );
 a29431a <=( a29430a  and  a29425a );
 a29435a <=( (not A298)  and  A268 );
 a29436a <=( (not A267)  and  a29435a );
 a29440a <=( A301  and  A300 );
 a29441a <=( A299  and  a29440a );
 a29442a <=( a29441a  and  a29436a );
 a29446a <=( (not A167)  and  A168 );
 a29447a <=( (not A170)  and  a29446a );
 a29451a <=( (not A200)  and  (not A199) );
 a29452a <=( A166  and  a29451a );
 a29453a <=( a29452a  and  a29447a );
 a29457a <=( (not A298)  and  A268 );
 a29458a <=( (not A267)  and  a29457a );
 a29462a <=( A302  and  A300 );
 a29463a <=( A299  and  a29462a );
 a29464a <=( a29463a  and  a29458a );
 a29468a <=( (not A167)  and  A168 );
 a29469a <=( (not A170)  and  a29468a );
 a29473a <=( (not A200)  and  (not A199) );
 a29474a <=( A166  and  a29473a );
 a29475a <=( a29474a  and  a29469a );
 a29479a <=( A298  and  A269 );
 a29480a <=( (not A267)  and  a29479a );
 a29484a <=( A301  and  A300 );
 a29485a <=( (not A299)  and  a29484a );
 a29486a <=( a29485a  and  a29480a );
 a29490a <=( (not A167)  and  A168 );
 a29491a <=( (not A170)  and  a29490a );
 a29495a <=( (not A200)  and  (not A199) );
 a29496a <=( A166  and  a29495a );
 a29497a <=( a29496a  and  a29491a );
 a29501a <=( A298  and  A269 );
 a29502a <=( (not A267)  and  a29501a );
 a29506a <=( A302  and  A300 );
 a29507a <=( (not A299)  and  a29506a );
 a29508a <=( a29507a  and  a29502a );
 a29512a <=( (not A167)  and  A168 );
 a29513a <=( (not A170)  and  a29512a );
 a29517a <=( (not A200)  and  (not A199) );
 a29518a <=( A166  and  a29517a );
 a29519a <=( a29518a  and  a29513a );
 a29523a <=( (not A298)  and  A269 );
 a29524a <=( (not A267)  and  a29523a );
 a29528a <=( A301  and  A300 );
 a29529a <=( A299  and  a29528a );
 a29530a <=( a29529a  and  a29524a );
 a29534a <=( (not A167)  and  A168 );
 a29535a <=( (not A170)  and  a29534a );
 a29539a <=( (not A200)  and  (not A199) );
 a29540a <=( A166  and  a29539a );
 a29541a <=( a29540a  and  a29535a );
 a29545a <=( (not A298)  and  A269 );
 a29546a <=( (not A267)  and  a29545a );
 a29550a <=( A302  and  A300 );
 a29551a <=( A299  and  a29550a );
 a29552a <=( a29551a  and  a29546a );
 a29556a <=( (not A167)  and  A168 );
 a29557a <=( (not A170)  and  a29556a );
 a29561a <=( (not A200)  and  (not A199) );
 a29562a <=( A166  and  a29561a );
 a29563a <=( a29562a  and  a29557a );
 a29567a <=( A298  and  A266 );
 a29568a <=( A265  and  a29567a );
 a29572a <=( A301  and  A300 );
 a29573a <=( (not A299)  and  a29572a );
 a29574a <=( a29573a  and  a29568a );
 a29578a <=( (not A167)  and  A168 );
 a29579a <=( (not A170)  and  a29578a );
 a29583a <=( (not A200)  and  (not A199) );
 a29584a <=( A166  and  a29583a );
 a29585a <=( a29584a  and  a29579a );
 a29589a <=( A298  and  A266 );
 a29590a <=( A265  and  a29589a );
 a29594a <=( A302  and  A300 );
 a29595a <=( (not A299)  and  a29594a );
 a29596a <=( a29595a  and  a29590a );
 a29600a <=( (not A167)  and  A168 );
 a29601a <=( (not A170)  and  a29600a );
 a29605a <=( (not A200)  and  (not A199) );
 a29606a <=( A166  and  a29605a );
 a29607a <=( a29606a  and  a29601a );
 a29611a <=( (not A298)  and  A266 );
 a29612a <=( A265  and  a29611a );
 a29616a <=( A301  and  A300 );
 a29617a <=( A299  and  a29616a );
 a29618a <=( a29617a  and  a29612a );
 a29622a <=( (not A167)  and  A168 );
 a29623a <=( (not A170)  and  a29622a );
 a29627a <=( (not A200)  and  (not A199) );
 a29628a <=( A166  and  a29627a );
 a29629a <=( a29628a  and  a29623a );
 a29633a <=( (not A298)  and  A266 );
 a29634a <=( A265  and  a29633a );
 a29638a <=( A302  and  A300 );
 a29639a <=( A299  and  a29638a );
 a29640a <=( a29639a  and  a29634a );
 a29644a <=( (not A167)  and  A168 );
 a29645a <=( (not A170)  and  a29644a );
 a29649a <=( (not A200)  and  (not A199) );
 a29650a <=( A166  and  a29649a );
 a29651a <=( a29650a  and  a29645a );
 a29655a <=( A298  and  (not A266) );
 a29656a <=( (not A265)  and  a29655a );
 a29660a <=( A301  and  A300 );
 a29661a <=( (not A299)  and  a29660a );
 a29662a <=( a29661a  and  a29656a );
 a29666a <=( (not A167)  and  A168 );
 a29667a <=( (not A170)  and  a29666a );
 a29671a <=( (not A200)  and  (not A199) );
 a29672a <=( A166  and  a29671a );
 a29673a <=( a29672a  and  a29667a );
 a29677a <=( A298  and  (not A266) );
 a29678a <=( (not A265)  and  a29677a );
 a29682a <=( A302  and  A300 );
 a29683a <=( (not A299)  and  a29682a );
 a29684a <=( a29683a  and  a29678a );
 a29688a <=( (not A167)  and  A168 );
 a29689a <=( (not A170)  and  a29688a );
 a29693a <=( (not A200)  and  (not A199) );
 a29694a <=( A166  and  a29693a );
 a29695a <=( a29694a  and  a29689a );
 a29699a <=( (not A298)  and  (not A266) );
 a29700a <=( (not A265)  and  a29699a );
 a29704a <=( A301  and  A300 );
 a29705a <=( A299  and  a29704a );
 a29706a <=( a29705a  and  a29700a );
 a29710a <=( (not A167)  and  A168 );
 a29711a <=( (not A170)  and  a29710a );
 a29715a <=( (not A200)  and  (not A199) );
 a29716a <=( A166  and  a29715a );
 a29717a <=( a29716a  and  a29711a );
 a29721a <=( (not A298)  and  (not A266) );
 a29722a <=( (not A265)  and  a29721a );
 a29726a <=( A302  and  A300 );
 a29727a <=( A299  and  a29726a );
 a29728a <=( a29727a  and  a29722a );
 a29732a <=( A201  and  (not A168) );
 a29733a <=( (not A170)  and  a29732a );
 a29737a <=( (not A265)  and  (not A203) );
 a29738a <=( (not A202)  and  a29737a );
 a29739a <=( a29738a  and  a29733a );
 a29743a <=( A268  and  A267 );
 a29744a <=( A266  and  a29743a );
 a29748a <=( (not A302)  and  (not A301) );
 a29749a <=( A300  and  a29748a );
 a29750a <=( a29749a  and  a29744a );
 a29754a <=( A201  and  (not A168) );
 a29755a <=( (not A170)  and  a29754a );
 a29759a <=( (not A265)  and  (not A203) );
 a29760a <=( (not A202)  and  a29759a );
 a29761a <=( a29760a  and  a29755a );
 a29765a <=( A269  and  A267 );
 a29766a <=( A266  and  a29765a );
 a29770a <=( (not A302)  and  (not A301) );
 a29771a <=( A300  and  a29770a );
 a29772a <=( a29771a  and  a29766a );
 a29776a <=( A201  and  (not A168) );
 a29777a <=( (not A170)  and  a29776a );
 a29781a <=( (not A265)  and  (not A203) );
 a29782a <=( (not A202)  and  a29781a );
 a29783a <=( a29782a  and  a29777a );
 a29787a <=( (not A268)  and  (not A267) );
 a29788a <=( A266  and  a29787a );
 a29792a <=( A301  and  (not A300) );
 a29793a <=( (not A269)  and  a29792a );
 a29794a <=( a29793a  and  a29788a );
 a29798a <=( A201  and  (not A168) );
 a29799a <=( (not A170)  and  a29798a );
 a29803a <=( (not A265)  and  (not A203) );
 a29804a <=( (not A202)  and  a29803a );
 a29805a <=( a29804a  and  a29799a );
 a29809a <=( (not A268)  and  (not A267) );
 a29810a <=( A266  and  a29809a );
 a29814a <=( A302  and  (not A300) );
 a29815a <=( (not A269)  and  a29814a );
 a29816a <=( a29815a  and  a29810a );
 a29820a <=( A201  and  (not A168) );
 a29821a <=( (not A170)  and  a29820a );
 a29825a <=( (not A265)  and  (not A203) );
 a29826a <=( (not A202)  and  a29825a );
 a29827a <=( a29826a  and  a29821a );
 a29831a <=( (not A268)  and  (not A267) );
 a29832a <=( A266  and  a29831a );
 a29836a <=( A299  and  A298 );
 a29837a <=( (not A269)  and  a29836a );
 a29838a <=( a29837a  and  a29832a );
 a29842a <=( A201  and  (not A168) );
 a29843a <=( (not A170)  and  a29842a );
 a29847a <=( (not A265)  and  (not A203) );
 a29848a <=( (not A202)  and  a29847a );
 a29849a <=( a29848a  and  a29843a );
 a29853a <=( (not A268)  and  (not A267) );
 a29854a <=( A266  and  a29853a );
 a29858a <=( (not A299)  and  (not A298) );
 a29859a <=( (not A269)  and  a29858a );
 a29860a <=( a29859a  and  a29854a );
 a29864a <=( A201  and  (not A168) );
 a29865a <=( (not A170)  and  a29864a );
 a29869a <=( A265  and  (not A203) );
 a29870a <=( (not A202)  and  a29869a );
 a29871a <=( a29870a  and  a29865a );
 a29875a <=( A268  and  A267 );
 a29876a <=( (not A266)  and  a29875a );
 a29880a <=( (not A302)  and  (not A301) );
 a29881a <=( A300  and  a29880a );
 a29882a <=( a29881a  and  a29876a );
 a29886a <=( A201  and  (not A168) );
 a29887a <=( (not A170)  and  a29886a );
 a29891a <=( A265  and  (not A203) );
 a29892a <=( (not A202)  and  a29891a );
 a29893a <=( a29892a  and  a29887a );
 a29897a <=( A269  and  A267 );
 a29898a <=( (not A266)  and  a29897a );
 a29902a <=( (not A302)  and  (not A301) );
 a29903a <=( A300  and  a29902a );
 a29904a <=( a29903a  and  a29898a );
 a29908a <=( A201  and  (not A168) );
 a29909a <=( (not A170)  and  a29908a );
 a29913a <=( A265  and  (not A203) );
 a29914a <=( (not A202)  and  a29913a );
 a29915a <=( a29914a  and  a29909a );
 a29919a <=( (not A268)  and  (not A267) );
 a29920a <=( (not A266)  and  a29919a );
 a29924a <=( A301  and  (not A300) );
 a29925a <=( (not A269)  and  a29924a );
 a29926a <=( a29925a  and  a29920a );
 a29930a <=( A201  and  (not A168) );
 a29931a <=( (not A170)  and  a29930a );
 a29935a <=( A265  and  (not A203) );
 a29936a <=( (not A202)  and  a29935a );
 a29937a <=( a29936a  and  a29931a );
 a29941a <=( (not A268)  and  (not A267) );
 a29942a <=( (not A266)  and  a29941a );
 a29946a <=( A302  and  (not A300) );
 a29947a <=( (not A269)  and  a29946a );
 a29948a <=( a29947a  and  a29942a );
 a29952a <=( A201  and  (not A168) );
 a29953a <=( (not A170)  and  a29952a );
 a29957a <=( A265  and  (not A203) );
 a29958a <=( (not A202)  and  a29957a );
 a29959a <=( a29958a  and  a29953a );
 a29963a <=( (not A268)  and  (not A267) );
 a29964a <=( (not A266)  and  a29963a );
 a29968a <=( A299  and  A298 );
 a29969a <=( (not A269)  and  a29968a );
 a29970a <=( a29969a  and  a29964a );
 a29974a <=( A201  and  (not A168) );
 a29975a <=( (not A170)  and  a29974a );
 a29979a <=( A265  and  (not A203) );
 a29980a <=( (not A202)  and  a29979a );
 a29981a <=( a29980a  and  a29975a );
 a29985a <=( (not A268)  and  (not A267) );
 a29986a <=( (not A266)  and  a29985a );
 a29990a <=( (not A299)  and  (not A298) );
 a29991a <=( (not A269)  and  a29990a );
 a29992a <=( a29991a  and  a29986a );
 a29996a <=( (not A201)  and  (not A168) );
 a29997a <=( (not A170)  and  a29996a );
 a30001a <=( A266  and  (not A265) );
 a30002a <=( A202  and  a30001a );
 a30003a <=( a30002a  and  a29997a );
 a30007a <=( (not A269)  and  (not A268) );
 a30008a <=( (not A267)  and  a30007a );
 a30012a <=( (not A302)  and  (not A301) );
 a30013a <=( A300  and  a30012a );
 a30014a <=( a30013a  and  a30008a );
 a30018a <=( (not A201)  and  (not A168) );
 a30019a <=( (not A170)  and  a30018a );
 a30023a <=( (not A266)  and  A265 );
 a30024a <=( A202  and  a30023a );
 a30025a <=( a30024a  and  a30019a );
 a30029a <=( (not A269)  and  (not A268) );
 a30030a <=( (not A267)  and  a30029a );
 a30034a <=( (not A302)  and  (not A301) );
 a30035a <=( A300  and  a30034a );
 a30036a <=( a30035a  and  a30030a );
 a30040a <=( (not A201)  and  (not A168) );
 a30041a <=( (not A170)  and  a30040a );
 a30045a <=( A266  and  (not A265) );
 a30046a <=( A203  and  a30045a );
 a30047a <=( a30046a  and  a30041a );
 a30051a <=( (not A269)  and  (not A268) );
 a30052a <=( (not A267)  and  a30051a );
 a30056a <=( (not A302)  and  (not A301) );
 a30057a <=( A300  and  a30056a );
 a30058a <=( a30057a  and  a30052a );
 a30062a <=( (not A201)  and  (not A168) );
 a30063a <=( (not A170)  and  a30062a );
 a30067a <=( (not A266)  and  A265 );
 a30068a <=( A203  and  a30067a );
 a30069a <=( a30068a  and  a30063a );
 a30073a <=( (not A269)  and  (not A268) );
 a30074a <=( (not A267)  and  a30073a );
 a30078a <=( (not A302)  and  (not A301) );
 a30079a <=( A300  and  a30078a );
 a30080a <=( a30079a  and  a30074a );
 a30084a <=( A199  and  (not A168) );
 a30085a <=( (not A170)  and  a30084a );
 a30089a <=( A266  and  (not A265) );
 a30090a <=( A200  and  a30089a );
 a30091a <=( a30090a  and  a30085a );
 a30095a <=( (not A269)  and  (not A268) );
 a30096a <=( (not A267)  and  a30095a );
 a30100a <=( (not A302)  and  (not A301) );
 a30101a <=( A300  and  a30100a );
 a30102a <=( a30101a  and  a30096a );
 a30106a <=( A199  and  (not A168) );
 a30107a <=( (not A170)  and  a30106a );
 a30111a <=( (not A266)  and  A265 );
 a30112a <=( A200  and  a30111a );
 a30113a <=( a30112a  and  a30107a );
 a30117a <=( (not A269)  and  (not A268) );
 a30118a <=( (not A267)  and  a30117a );
 a30122a <=( (not A302)  and  (not A301) );
 a30123a <=( A300  and  a30122a );
 a30124a <=( a30123a  and  a30118a );
 a30128a <=( (not A199)  and  (not A168) );
 a30129a <=( (not A170)  and  a30128a );
 a30133a <=( A202  and  A201 );
 a30134a <=( A200  and  a30133a );
 a30135a <=( a30134a  and  a30129a );
 a30139a <=( A298  and  A268 );
 a30140a <=( (not A267)  and  a30139a );
 a30144a <=( A301  and  A300 );
 a30145a <=( (not A299)  and  a30144a );
 a30146a <=( a30145a  and  a30140a );
 a30150a <=( (not A199)  and  (not A168) );
 a30151a <=( (not A170)  and  a30150a );
 a30155a <=( A202  and  A201 );
 a30156a <=( A200  and  a30155a );
 a30157a <=( a30156a  and  a30151a );
 a30161a <=( A298  and  A268 );
 a30162a <=( (not A267)  and  a30161a );
 a30166a <=( A302  and  A300 );
 a30167a <=( (not A299)  and  a30166a );
 a30168a <=( a30167a  and  a30162a );
 a30172a <=( (not A199)  and  (not A168) );
 a30173a <=( (not A170)  and  a30172a );
 a30177a <=( A202  and  A201 );
 a30178a <=( A200  and  a30177a );
 a30179a <=( a30178a  and  a30173a );
 a30183a <=( (not A298)  and  A268 );
 a30184a <=( (not A267)  and  a30183a );
 a30188a <=( A301  and  A300 );
 a30189a <=( A299  and  a30188a );
 a30190a <=( a30189a  and  a30184a );
 a30194a <=( (not A199)  and  (not A168) );
 a30195a <=( (not A170)  and  a30194a );
 a30199a <=( A202  and  A201 );
 a30200a <=( A200  and  a30199a );
 a30201a <=( a30200a  and  a30195a );
 a30205a <=( (not A298)  and  A268 );
 a30206a <=( (not A267)  and  a30205a );
 a30210a <=( A302  and  A300 );
 a30211a <=( A299  and  a30210a );
 a30212a <=( a30211a  and  a30206a );
 a30216a <=( (not A199)  and  (not A168) );
 a30217a <=( (not A170)  and  a30216a );
 a30221a <=( A202  and  A201 );
 a30222a <=( A200  and  a30221a );
 a30223a <=( a30222a  and  a30217a );
 a30227a <=( A298  and  A269 );
 a30228a <=( (not A267)  and  a30227a );
 a30232a <=( A301  and  A300 );
 a30233a <=( (not A299)  and  a30232a );
 a30234a <=( a30233a  and  a30228a );
 a30238a <=( (not A199)  and  (not A168) );
 a30239a <=( (not A170)  and  a30238a );
 a30243a <=( A202  and  A201 );
 a30244a <=( A200  and  a30243a );
 a30245a <=( a30244a  and  a30239a );
 a30249a <=( A298  and  A269 );
 a30250a <=( (not A267)  and  a30249a );
 a30254a <=( A302  and  A300 );
 a30255a <=( (not A299)  and  a30254a );
 a30256a <=( a30255a  and  a30250a );
 a30260a <=( (not A199)  and  (not A168) );
 a30261a <=( (not A170)  and  a30260a );
 a30265a <=( A202  and  A201 );
 a30266a <=( A200  and  a30265a );
 a30267a <=( a30266a  and  a30261a );
 a30271a <=( (not A298)  and  A269 );
 a30272a <=( (not A267)  and  a30271a );
 a30276a <=( A301  and  A300 );
 a30277a <=( A299  and  a30276a );
 a30278a <=( a30277a  and  a30272a );
 a30282a <=( (not A199)  and  (not A168) );
 a30283a <=( (not A170)  and  a30282a );
 a30287a <=( A202  and  A201 );
 a30288a <=( A200  and  a30287a );
 a30289a <=( a30288a  and  a30283a );
 a30293a <=( (not A298)  and  A269 );
 a30294a <=( (not A267)  and  a30293a );
 a30298a <=( A302  and  A300 );
 a30299a <=( A299  and  a30298a );
 a30300a <=( a30299a  and  a30294a );
 a30304a <=( (not A199)  and  (not A168) );
 a30305a <=( (not A170)  and  a30304a );
 a30309a <=( A202  and  A201 );
 a30310a <=( A200  and  a30309a );
 a30311a <=( a30310a  and  a30305a );
 a30315a <=( A298  and  A266 );
 a30316a <=( A265  and  a30315a );
 a30320a <=( A301  and  A300 );
 a30321a <=( (not A299)  and  a30320a );
 a30322a <=( a30321a  and  a30316a );
 a30326a <=( (not A199)  and  (not A168) );
 a30327a <=( (not A170)  and  a30326a );
 a30331a <=( A202  and  A201 );
 a30332a <=( A200  and  a30331a );
 a30333a <=( a30332a  and  a30327a );
 a30337a <=( A298  and  A266 );
 a30338a <=( A265  and  a30337a );
 a30342a <=( A302  and  A300 );
 a30343a <=( (not A299)  and  a30342a );
 a30344a <=( a30343a  and  a30338a );
 a30348a <=( (not A199)  and  (not A168) );
 a30349a <=( (not A170)  and  a30348a );
 a30353a <=( A202  and  A201 );
 a30354a <=( A200  and  a30353a );
 a30355a <=( a30354a  and  a30349a );
 a30359a <=( (not A298)  and  A266 );
 a30360a <=( A265  and  a30359a );
 a30364a <=( A301  and  A300 );
 a30365a <=( A299  and  a30364a );
 a30366a <=( a30365a  and  a30360a );
 a30370a <=( (not A199)  and  (not A168) );
 a30371a <=( (not A170)  and  a30370a );
 a30375a <=( A202  and  A201 );
 a30376a <=( A200  and  a30375a );
 a30377a <=( a30376a  and  a30371a );
 a30381a <=( (not A298)  and  A266 );
 a30382a <=( A265  and  a30381a );
 a30386a <=( A302  and  A300 );
 a30387a <=( A299  and  a30386a );
 a30388a <=( a30387a  and  a30382a );
 a30392a <=( (not A199)  and  (not A168) );
 a30393a <=( (not A170)  and  a30392a );
 a30397a <=( A202  and  A201 );
 a30398a <=( A200  and  a30397a );
 a30399a <=( a30398a  and  a30393a );
 a30403a <=( A298  and  (not A266) );
 a30404a <=( (not A265)  and  a30403a );
 a30408a <=( A301  and  A300 );
 a30409a <=( (not A299)  and  a30408a );
 a30410a <=( a30409a  and  a30404a );
 a30414a <=( (not A199)  and  (not A168) );
 a30415a <=( (not A170)  and  a30414a );
 a30419a <=( A202  and  A201 );
 a30420a <=( A200  and  a30419a );
 a30421a <=( a30420a  and  a30415a );
 a30425a <=( A298  and  (not A266) );
 a30426a <=( (not A265)  and  a30425a );
 a30430a <=( A302  and  A300 );
 a30431a <=( (not A299)  and  a30430a );
 a30432a <=( a30431a  and  a30426a );
 a30436a <=( (not A199)  and  (not A168) );
 a30437a <=( (not A170)  and  a30436a );
 a30441a <=( A202  and  A201 );
 a30442a <=( A200  and  a30441a );
 a30443a <=( a30442a  and  a30437a );
 a30447a <=( (not A298)  and  (not A266) );
 a30448a <=( (not A265)  and  a30447a );
 a30452a <=( A301  and  A300 );
 a30453a <=( A299  and  a30452a );
 a30454a <=( a30453a  and  a30448a );
 a30458a <=( (not A199)  and  (not A168) );
 a30459a <=( (not A170)  and  a30458a );
 a30463a <=( A202  and  A201 );
 a30464a <=( A200  and  a30463a );
 a30465a <=( a30464a  and  a30459a );
 a30469a <=( (not A298)  and  (not A266) );
 a30470a <=( (not A265)  and  a30469a );
 a30474a <=( A302  and  A300 );
 a30475a <=( A299  and  a30474a );
 a30476a <=( a30475a  and  a30470a );
 a30480a <=( (not A199)  and  (not A168) );
 a30481a <=( (not A170)  and  a30480a );
 a30485a <=( A203  and  A201 );
 a30486a <=( A200  and  a30485a );
 a30487a <=( a30486a  and  a30481a );
 a30491a <=( A298  and  A268 );
 a30492a <=( (not A267)  and  a30491a );
 a30496a <=( A301  and  A300 );
 a30497a <=( (not A299)  and  a30496a );
 a30498a <=( a30497a  and  a30492a );
 a30502a <=( (not A199)  and  (not A168) );
 a30503a <=( (not A170)  and  a30502a );
 a30507a <=( A203  and  A201 );
 a30508a <=( A200  and  a30507a );
 a30509a <=( a30508a  and  a30503a );
 a30513a <=( A298  and  A268 );
 a30514a <=( (not A267)  and  a30513a );
 a30518a <=( A302  and  A300 );
 a30519a <=( (not A299)  and  a30518a );
 a30520a <=( a30519a  and  a30514a );
 a30524a <=( (not A199)  and  (not A168) );
 a30525a <=( (not A170)  and  a30524a );
 a30529a <=( A203  and  A201 );
 a30530a <=( A200  and  a30529a );
 a30531a <=( a30530a  and  a30525a );
 a30535a <=( (not A298)  and  A268 );
 a30536a <=( (not A267)  and  a30535a );
 a30540a <=( A301  and  A300 );
 a30541a <=( A299  and  a30540a );
 a30542a <=( a30541a  and  a30536a );
 a30546a <=( (not A199)  and  (not A168) );
 a30547a <=( (not A170)  and  a30546a );
 a30551a <=( A203  and  A201 );
 a30552a <=( A200  and  a30551a );
 a30553a <=( a30552a  and  a30547a );
 a30557a <=( (not A298)  and  A268 );
 a30558a <=( (not A267)  and  a30557a );
 a30562a <=( A302  and  A300 );
 a30563a <=( A299  and  a30562a );
 a30564a <=( a30563a  and  a30558a );
 a30568a <=( (not A199)  and  (not A168) );
 a30569a <=( (not A170)  and  a30568a );
 a30573a <=( A203  and  A201 );
 a30574a <=( A200  and  a30573a );
 a30575a <=( a30574a  and  a30569a );
 a30579a <=( A298  and  A269 );
 a30580a <=( (not A267)  and  a30579a );
 a30584a <=( A301  and  A300 );
 a30585a <=( (not A299)  and  a30584a );
 a30586a <=( a30585a  and  a30580a );
 a30590a <=( (not A199)  and  (not A168) );
 a30591a <=( (not A170)  and  a30590a );
 a30595a <=( A203  and  A201 );
 a30596a <=( A200  and  a30595a );
 a30597a <=( a30596a  and  a30591a );
 a30601a <=( A298  and  A269 );
 a30602a <=( (not A267)  and  a30601a );
 a30606a <=( A302  and  A300 );
 a30607a <=( (not A299)  and  a30606a );
 a30608a <=( a30607a  and  a30602a );
 a30612a <=( (not A199)  and  (not A168) );
 a30613a <=( (not A170)  and  a30612a );
 a30617a <=( A203  and  A201 );
 a30618a <=( A200  and  a30617a );
 a30619a <=( a30618a  and  a30613a );
 a30623a <=( (not A298)  and  A269 );
 a30624a <=( (not A267)  and  a30623a );
 a30628a <=( A301  and  A300 );
 a30629a <=( A299  and  a30628a );
 a30630a <=( a30629a  and  a30624a );
 a30634a <=( (not A199)  and  (not A168) );
 a30635a <=( (not A170)  and  a30634a );
 a30639a <=( A203  and  A201 );
 a30640a <=( A200  and  a30639a );
 a30641a <=( a30640a  and  a30635a );
 a30645a <=( (not A298)  and  A269 );
 a30646a <=( (not A267)  and  a30645a );
 a30650a <=( A302  and  A300 );
 a30651a <=( A299  and  a30650a );
 a30652a <=( a30651a  and  a30646a );
 a30656a <=( (not A199)  and  (not A168) );
 a30657a <=( (not A170)  and  a30656a );
 a30661a <=( A203  and  A201 );
 a30662a <=( A200  and  a30661a );
 a30663a <=( a30662a  and  a30657a );
 a30667a <=( A298  and  A266 );
 a30668a <=( A265  and  a30667a );
 a30672a <=( A301  and  A300 );
 a30673a <=( (not A299)  and  a30672a );
 a30674a <=( a30673a  and  a30668a );
 a30678a <=( (not A199)  and  (not A168) );
 a30679a <=( (not A170)  and  a30678a );
 a30683a <=( A203  and  A201 );
 a30684a <=( A200  and  a30683a );
 a30685a <=( a30684a  and  a30679a );
 a30689a <=( A298  and  A266 );
 a30690a <=( A265  and  a30689a );
 a30694a <=( A302  and  A300 );
 a30695a <=( (not A299)  and  a30694a );
 a30696a <=( a30695a  and  a30690a );
 a30700a <=( (not A199)  and  (not A168) );
 a30701a <=( (not A170)  and  a30700a );
 a30705a <=( A203  and  A201 );
 a30706a <=( A200  and  a30705a );
 a30707a <=( a30706a  and  a30701a );
 a30711a <=( (not A298)  and  A266 );
 a30712a <=( A265  and  a30711a );
 a30716a <=( A301  and  A300 );
 a30717a <=( A299  and  a30716a );
 a30718a <=( a30717a  and  a30712a );
 a30722a <=( (not A199)  and  (not A168) );
 a30723a <=( (not A170)  and  a30722a );
 a30727a <=( A203  and  A201 );
 a30728a <=( A200  and  a30727a );
 a30729a <=( a30728a  and  a30723a );
 a30733a <=( (not A298)  and  A266 );
 a30734a <=( A265  and  a30733a );
 a30738a <=( A302  and  A300 );
 a30739a <=( A299  and  a30738a );
 a30740a <=( a30739a  and  a30734a );
 a30744a <=( (not A199)  and  (not A168) );
 a30745a <=( (not A170)  and  a30744a );
 a30749a <=( A203  and  A201 );
 a30750a <=( A200  and  a30749a );
 a30751a <=( a30750a  and  a30745a );
 a30755a <=( A298  and  (not A266) );
 a30756a <=( (not A265)  and  a30755a );
 a30760a <=( A301  and  A300 );
 a30761a <=( (not A299)  and  a30760a );
 a30762a <=( a30761a  and  a30756a );
 a30766a <=( (not A199)  and  (not A168) );
 a30767a <=( (not A170)  and  a30766a );
 a30771a <=( A203  and  A201 );
 a30772a <=( A200  and  a30771a );
 a30773a <=( a30772a  and  a30767a );
 a30777a <=( A298  and  (not A266) );
 a30778a <=( (not A265)  and  a30777a );
 a30782a <=( A302  and  A300 );
 a30783a <=( (not A299)  and  a30782a );
 a30784a <=( a30783a  and  a30778a );
 a30788a <=( (not A199)  and  (not A168) );
 a30789a <=( (not A170)  and  a30788a );
 a30793a <=( A203  and  A201 );
 a30794a <=( A200  and  a30793a );
 a30795a <=( a30794a  and  a30789a );
 a30799a <=( (not A298)  and  (not A266) );
 a30800a <=( (not A265)  and  a30799a );
 a30804a <=( A301  and  A300 );
 a30805a <=( A299  and  a30804a );
 a30806a <=( a30805a  and  a30800a );
 a30810a <=( (not A199)  and  (not A168) );
 a30811a <=( (not A170)  and  a30810a );
 a30815a <=( A203  and  A201 );
 a30816a <=( A200  and  a30815a );
 a30817a <=( a30816a  and  a30811a );
 a30821a <=( (not A298)  and  (not A266) );
 a30822a <=( (not A265)  and  a30821a );
 a30826a <=( A302  and  A300 );
 a30827a <=( A299  and  a30826a );
 a30828a <=( a30827a  and  a30822a );
 a30832a <=( A199  and  (not A168) );
 a30833a <=( (not A170)  and  a30832a );
 a30837a <=( A202  and  A201 );
 a30838a <=( (not A200)  and  a30837a );
 a30839a <=( a30838a  and  a30833a );
 a30843a <=( A298  and  A268 );
 a30844a <=( (not A267)  and  a30843a );
 a30848a <=( A301  and  A300 );
 a30849a <=( (not A299)  and  a30848a );
 a30850a <=( a30849a  and  a30844a );
 a30854a <=( A199  and  (not A168) );
 a30855a <=( (not A170)  and  a30854a );
 a30859a <=( A202  and  A201 );
 a30860a <=( (not A200)  and  a30859a );
 a30861a <=( a30860a  and  a30855a );
 a30865a <=( A298  and  A268 );
 a30866a <=( (not A267)  and  a30865a );
 a30870a <=( A302  and  A300 );
 a30871a <=( (not A299)  and  a30870a );
 a30872a <=( a30871a  and  a30866a );
 a30876a <=( A199  and  (not A168) );
 a30877a <=( (not A170)  and  a30876a );
 a30881a <=( A202  and  A201 );
 a30882a <=( (not A200)  and  a30881a );
 a30883a <=( a30882a  and  a30877a );
 a30887a <=( (not A298)  and  A268 );
 a30888a <=( (not A267)  and  a30887a );
 a30892a <=( A301  and  A300 );
 a30893a <=( A299  and  a30892a );
 a30894a <=( a30893a  and  a30888a );
 a30898a <=( A199  and  (not A168) );
 a30899a <=( (not A170)  and  a30898a );
 a30903a <=( A202  and  A201 );
 a30904a <=( (not A200)  and  a30903a );
 a30905a <=( a30904a  and  a30899a );
 a30909a <=( (not A298)  and  A268 );
 a30910a <=( (not A267)  and  a30909a );
 a30914a <=( A302  and  A300 );
 a30915a <=( A299  and  a30914a );
 a30916a <=( a30915a  and  a30910a );
 a30920a <=( A199  and  (not A168) );
 a30921a <=( (not A170)  and  a30920a );
 a30925a <=( A202  and  A201 );
 a30926a <=( (not A200)  and  a30925a );
 a30927a <=( a30926a  and  a30921a );
 a30931a <=( A298  and  A269 );
 a30932a <=( (not A267)  and  a30931a );
 a30936a <=( A301  and  A300 );
 a30937a <=( (not A299)  and  a30936a );
 a30938a <=( a30937a  and  a30932a );
 a30942a <=( A199  and  (not A168) );
 a30943a <=( (not A170)  and  a30942a );
 a30947a <=( A202  and  A201 );
 a30948a <=( (not A200)  and  a30947a );
 a30949a <=( a30948a  and  a30943a );
 a30953a <=( A298  and  A269 );
 a30954a <=( (not A267)  and  a30953a );
 a30958a <=( A302  and  A300 );
 a30959a <=( (not A299)  and  a30958a );
 a30960a <=( a30959a  and  a30954a );
 a30964a <=( A199  and  (not A168) );
 a30965a <=( (not A170)  and  a30964a );
 a30969a <=( A202  and  A201 );
 a30970a <=( (not A200)  and  a30969a );
 a30971a <=( a30970a  and  a30965a );
 a30975a <=( (not A298)  and  A269 );
 a30976a <=( (not A267)  and  a30975a );
 a30980a <=( A301  and  A300 );
 a30981a <=( A299  and  a30980a );
 a30982a <=( a30981a  and  a30976a );
 a30986a <=( A199  and  (not A168) );
 a30987a <=( (not A170)  and  a30986a );
 a30991a <=( A202  and  A201 );
 a30992a <=( (not A200)  and  a30991a );
 a30993a <=( a30992a  and  a30987a );
 a30997a <=( (not A298)  and  A269 );
 a30998a <=( (not A267)  and  a30997a );
 a31002a <=( A302  and  A300 );
 a31003a <=( A299  and  a31002a );
 a31004a <=( a31003a  and  a30998a );
 a31008a <=( A199  and  (not A168) );
 a31009a <=( (not A170)  and  a31008a );
 a31013a <=( A202  and  A201 );
 a31014a <=( (not A200)  and  a31013a );
 a31015a <=( a31014a  and  a31009a );
 a31019a <=( A298  and  A266 );
 a31020a <=( A265  and  a31019a );
 a31024a <=( A301  and  A300 );
 a31025a <=( (not A299)  and  a31024a );
 a31026a <=( a31025a  and  a31020a );
 a31030a <=( A199  and  (not A168) );
 a31031a <=( (not A170)  and  a31030a );
 a31035a <=( A202  and  A201 );
 a31036a <=( (not A200)  and  a31035a );
 a31037a <=( a31036a  and  a31031a );
 a31041a <=( A298  and  A266 );
 a31042a <=( A265  and  a31041a );
 a31046a <=( A302  and  A300 );
 a31047a <=( (not A299)  and  a31046a );
 a31048a <=( a31047a  and  a31042a );
 a31052a <=( A199  and  (not A168) );
 a31053a <=( (not A170)  and  a31052a );
 a31057a <=( A202  and  A201 );
 a31058a <=( (not A200)  and  a31057a );
 a31059a <=( a31058a  and  a31053a );
 a31063a <=( (not A298)  and  A266 );
 a31064a <=( A265  and  a31063a );
 a31068a <=( A301  and  A300 );
 a31069a <=( A299  and  a31068a );
 a31070a <=( a31069a  and  a31064a );
 a31074a <=( A199  and  (not A168) );
 a31075a <=( (not A170)  and  a31074a );
 a31079a <=( A202  and  A201 );
 a31080a <=( (not A200)  and  a31079a );
 a31081a <=( a31080a  and  a31075a );
 a31085a <=( (not A298)  and  A266 );
 a31086a <=( A265  and  a31085a );
 a31090a <=( A302  and  A300 );
 a31091a <=( A299  and  a31090a );
 a31092a <=( a31091a  and  a31086a );
 a31096a <=( A199  and  (not A168) );
 a31097a <=( (not A170)  and  a31096a );
 a31101a <=( A202  and  A201 );
 a31102a <=( (not A200)  and  a31101a );
 a31103a <=( a31102a  and  a31097a );
 a31107a <=( A298  and  (not A266) );
 a31108a <=( (not A265)  and  a31107a );
 a31112a <=( A301  and  A300 );
 a31113a <=( (not A299)  and  a31112a );
 a31114a <=( a31113a  and  a31108a );
 a31118a <=( A199  and  (not A168) );
 a31119a <=( (not A170)  and  a31118a );
 a31123a <=( A202  and  A201 );
 a31124a <=( (not A200)  and  a31123a );
 a31125a <=( a31124a  and  a31119a );
 a31129a <=( A298  and  (not A266) );
 a31130a <=( (not A265)  and  a31129a );
 a31134a <=( A302  and  A300 );
 a31135a <=( (not A299)  and  a31134a );
 a31136a <=( a31135a  and  a31130a );
 a31140a <=( A199  and  (not A168) );
 a31141a <=( (not A170)  and  a31140a );
 a31145a <=( A202  and  A201 );
 a31146a <=( (not A200)  and  a31145a );
 a31147a <=( a31146a  and  a31141a );
 a31151a <=( (not A298)  and  (not A266) );
 a31152a <=( (not A265)  and  a31151a );
 a31156a <=( A301  and  A300 );
 a31157a <=( A299  and  a31156a );
 a31158a <=( a31157a  and  a31152a );
 a31162a <=( A199  and  (not A168) );
 a31163a <=( (not A170)  and  a31162a );
 a31167a <=( A202  and  A201 );
 a31168a <=( (not A200)  and  a31167a );
 a31169a <=( a31168a  and  a31163a );
 a31173a <=( (not A298)  and  (not A266) );
 a31174a <=( (not A265)  and  a31173a );
 a31178a <=( A302  and  A300 );
 a31179a <=( A299  and  a31178a );
 a31180a <=( a31179a  and  a31174a );
 a31184a <=( A199  and  (not A168) );
 a31185a <=( (not A170)  and  a31184a );
 a31189a <=( A203  and  A201 );
 a31190a <=( (not A200)  and  a31189a );
 a31191a <=( a31190a  and  a31185a );
 a31195a <=( A298  and  A268 );
 a31196a <=( (not A267)  and  a31195a );
 a31200a <=( A301  and  A300 );
 a31201a <=( (not A299)  and  a31200a );
 a31202a <=( a31201a  and  a31196a );
 a31206a <=( A199  and  (not A168) );
 a31207a <=( (not A170)  and  a31206a );
 a31211a <=( A203  and  A201 );
 a31212a <=( (not A200)  and  a31211a );
 a31213a <=( a31212a  and  a31207a );
 a31217a <=( A298  and  A268 );
 a31218a <=( (not A267)  and  a31217a );
 a31222a <=( A302  and  A300 );
 a31223a <=( (not A299)  and  a31222a );
 a31224a <=( a31223a  and  a31218a );
 a31228a <=( A199  and  (not A168) );
 a31229a <=( (not A170)  and  a31228a );
 a31233a <=( A203  and  A201 );
 a31234a <=( (not A200)  and  a31233a );
 a31235a <=( a31234a  and  a31229a );
 a31239a <=( (not A298)  and  A268 );
 a31240a <=( (not A267)  and  a31239a );
 a31244a <=( A301  and  A300 );
 a31245a <=( A299  and  a31244a );
 a31246a <=( a31245a  and  a31240a );
 a31250a <=( A199  and  (not A168) );
 a31251a <=( (not A170)  and  a31250a );
 a31255a <=( A203  and  A201 );
 a31256a <=( (not A200)  and  a31255a );
 a31257a <=( a31256a  and  a31251a );
 a31261a <=( (not A298)  and  A268 );
 a31262a <=( (not A267)  and  a31261a );
 a31266a <=( A302  and  A300 );
 a31267a <=( A299  and  a31266a );
 a31268a <=( a31267a  and  a31262a );
 a31272a <=( A199  and  (not A168) );
 a31273a <=( (not A170)  and  a31272a );
 a31277a <=( A203  and  A201 );
 a31278a <=( (not A200)  and  a31277a );
 a31279a <=( a31278a  and  a31273a );
 a31283a <=( A298  and  A269 );
 a31284a <=( (not A267)  and  a31283a );
 a31288a <=( A301  and  A300 );
 a31289a <=( (not A299)  and  a31288a );
 a31290a <=( a31289a  and  a31284a );
 a31294a <=( A199  and  (not A168) );
 a31295a <=( (not A170)  and  a31294a );
 a31299a <=( A203  and  A201 );
 a31300a <=( (not A200)  and  a31299a );
 a31301a <=( a31300a  and  a31295a );
 a31305a <=( A298  and  A269 );
 a31306a <=( (not A267)  and  a31305a );
 a31310a <=( A302  and  A300 );
 a31311a <=( (not A299)  and  a31310a );
 a31312a <=( a31311a  and  a31306a );
 a31316a <=( A199  and  (not A168) );
 a31317a <=( (not A170)  and  a31316a );
 a31321a <=( A203  and  A201 );
 a31322a <=( (not A200)  and  a31321a );
 a31323a <=( a31322a  and  a31317a );
 a31327a <=( (not A298)  and  A269 );
 a31328a <=( (not A267)  and  a31327a );
 a31332a <=( A301  and  A300 );
 a31333a <=( A299  and  a31332a );
 a31334a <=( a31333a  and  a31328a );
 a31338a <=( A199  and  (not A168) );
 a31339a <=( (not A170)  and  a31338a );
 a31343a <=( A203  and  A201 );
 a31344a <=( (not A200)  and  a31343a );
 a31345a <=( a31344a  and  a31339a );
 a31349a <=( (not A298)  and  A269 );
 a31350a <=( (not A267)  and  a31349a );
 a31354a <=( A302  and  A300 );
 a31355a <=( A299  and  a31354a );
 a31356a <=( a31355a  and  a31350a );
 a31360a <=( A199  and  (not A168) );
 a31361a <=( (not A170)  and  a31360a );
 a31365a <=( A203  and  A201 );
 a31366a <=( (not A200)  and  a31365a );
 a31367a <=( a31366a  and  a31361a );
 a31371a <=( A298  and  A266 );
 a31372a <=( A265  and  a31371a );
 a31376a <=( A301  and  A300 );
 a31377a <=( (not A299)  and  a31376a );
 a31378a <=( a31377a  and  a31372a );
 a31382a <=( A199  and  (not A168) );
 a31383a <=( (not A170)  and  a31382a );
 a31387a <=( A203  and  A201 );
 a31388a <=( (not A200)  and  a31387a );
 a31389a <=( a31388a  and  a31383a );
 a31393a <=( A298  and  A266 );
 a31394a <=( A265  and  a31393a );
 a31398a <=( A302  and  A300 );
 a31399a <=( (not A299)  and  a31398a );
 a31400a <=( a31399a  and  a31394a );
 a31404a <=( A199  and  (not A168) );
 a31405a <=( (not A170)  and  a31404a );
 a31409a <=( A203  and  A201 );
 a31410a <=( (not A200)  and  a31409a );
 a31411a <=( a31410a  and  a31405a );
 a31415a <=( (not A298)  and  A266 );
 a31416a <=( A265  and  a31415a );
 a31420a <=( A301  and  A300 );
 a31421a <=( A299  and  a31420a );
 a31422a <=( a31421a  and  a31416a );
 a31426a <=( A199  and  (not A168) );
 a31427a <=( (not A170)  and  a31426a );
 a31431a <=( A203  and  A201 );
 a31432a <=( (not A200)  and  a31431a );
 a31433a <=( a31432a  and  a31427a );
 a31437a <=( (not A298)  and  A266 );
 a31438a <=( A265  and  a31437a );
 a31442a <=( A302  and  A300 );
 a31443a <=( A299  and  a31442a );
 a31444a <=( a31443a  and  a31438a );
 a31448a <=( A199  and  (not A168) );
 a31449a <=( (not A170)  and  a31448a );
 a31453a <=( A203  and  A201 );
 a31454a <=( (not A200)  and  a31453a );
 a31455a <=( a31454a  and  a31449a );
 a31459a <=( A298  and  (not A266) );
 a31460a <=( (not A265)  and  a31459a );
 a31464a <=( A301  and  A300 );
 a31465a <=( (not A299)  and  a31464a );
 a31466a <=( a31465a  and  a31460a );
 a31470a <=( A199  and  (not A168) );
 a31471a <=( (not A170)  and  a31470a );
 a31475a <=( A203  and  A201 );
 a31476a <=( (not A200)  and  a31475a );
 a31477a <=( a31476a  and  a31471a );
 a31481a <=( A298  and  (not A266) );
 a31482a <=( (not A265)  and  a31481a );
 a31486a <=( A302  and  A300 );
 a31487a <=( (not A299)  and  a31486a );
 a31488a <=( a31487a  and  a31482a );
 a31492a <=( A199  and  (not A168) );
 a31493a <=( (not A170)  and  a31492a );
 a31497a <=( A203  and  A201 );
 a31498a <=( (not A200)  and  a31497a );
 a31499a <=( a31498a  and  a31493a );
 a31503a <=( (not A298)  and  (not A266) );
 a31504a <=( (not A265)  and  a31503a );
 a31508a <=( A301  and  A300 );
 a31509a <=( A299  and  a31508a );
 a31510a <=( a31509a  and  a31504a );
 a31514a <=( A199  and  (not A168) );
 a31515a <=( (not A170)  and  a31514a );
 a31519a <=( A203  and  A201 );
 a31520a <=( (not A200)  and  a31519a );
 a31521a <=( a31520a  and  a31515a );
 a31525a <=( (not A298)  and  (not A266) );
 a31526a <=( (not A265)  and  a31525a );
 a31530a <=( A302  and  A300 );
 a31531a <=( A299  and  a31530a );
 a31532a <=( a31531a  and  a31526a );
 a31536a <=( (not A199)  and  (not A168) );
 a31537a <=( (not A170)  and  a31536a );
 a31541a <=( A266  and  (not A265) );
 a31542a <=( (not A200)  and  a31541a );
 a31543a <=( a31542a  and  a31537a );
 a31547a <=( (not A269)  and  (not A268) );
 a31548a <=( (not A267)  and  a31547a );
 a31552a <=( (not A302)  and  (not A301) );
 a31553a <=( A300  and  a31552a );
 a31554a <=( a31553a  and  a31548a );
 a31558a <=( (not A199)  and  (not A168) );
 a31559a <=( (not A170)  and  a31558a );
 a31563a <=( (not A266)  and  A265 );
 a31564a <=( (not A200)  and  a31563a );
 a31565a <=( a31564a  and  a31559a );
 a31569a <=( (not A269)  and  (not A268) );
 a31570a <=( (not A267)  and  a31569a );
 a31574a <=( (not A302)  and  (not A301) );
 a31575a <=( A300  and  a31574a );
 a31576a <=( a31575a  and  a31570a );
 a31580a <=( A167  and  A168 );
 a31581a <=( A169  and  a31580a );
 a31585a <=( A202  and  (not A201) );
 a31586a <=( (not A166)  and  a31585a );
 a31587a <=( a31586a  and  a31581a );
 a31591a <=( A298  and  A268 );
 a31592a <=( (not A267)  and  a31591a );
 a31596a <=( A301  and  A300 );
 a31597a <=( (not A299)  and  a31596a );
 a31598a <=( a31597a  and  a31592a );
 a31602a <=( A167  and  A168 );
 a31603a <=( A169  and  a31602a );
 a31607a <=( A202  and  (not A201) );
 a31608a <=( (not A166)  and  a31607a );
 a31609a <=( a31608a  and  a31603a );
 a31613a <=( A298  and  A268 );
 a31614a <=( (not A267)  and  a31613a );
 a31618a <=( A302  and  A300 );
 a31619a <=( (not A299)  and  a31618a );
 a31620a <=( a31619a  and  a31614a );
 a31624a <=( A167  and  A168 );
 a31625a <=( A169  and  a31624a );
 a31629a <=( A202  and  (not A201) );
 a31630a <=( (not A166)  and  a31629a );
 a31631a <=( a31630a  and  a31625a );
 a31635a <=( (not A298)  and  A268 );
 a31636a <=( (not A267)  and  a31635a );
 a31640a <=( A301  and  A300 );
 a31641a <=( A299  and  a31640a );
 a31642a <=( a31641a  and  a31636a );
 a31646a <=( A167  and  A168 );
 a31647a <=( A169  and  a31646a );
 a31651a <=( A202  and  (not A201) );
 a31652a <=( (not A166)  and  a31651a );
 a31653a <=( a31652a  and  a31647a );
 a31657a <=( (not A298)  and  A268 );
 a31658a <=( (not A267)  and  a31657a );
 a31662a <=( A302  and  A300 );
 a31663a <=( A299  and  a31662a );
 a31664a <=( a31663a  and  a31658a );
 a31668a <=( A167  and  A168 );
 a31669a <=( A169  and  a31668a );
 a31673a <=( A202  and  (not A201) );
 a31674a <=( (not A166)  and  a31673a );
 a31675a <=( a31674a  and  a31669a );
 a31679a <=( A298  and  A269 );
 a31680a <=( (not A267)  and  a31679a );
 a31684a <=( A301  and  A300 );
 a31685a <=( (not A299)  and  a31684a );
 a31686a <=( a31685a  and  a31680a );
 a31690a <=( A167  and  A168 );
 a31691a <=( A169  and  a31690a );
 a31695a <=( A202  and  (not A201) );
 a31696a <=( (not A166)  and  a31695a );
 a31697a <=( a31696a  and  a31691a );
 a31701a <=( A298  and  A269 );
 a31702a <=( (not A267)  and  a31701a );
 a31706a <=( A302  and  A300 );
 a31707a <=( (not A299)  and  a31706a );
 a31708a <=( a31707a  and  a31702a );
 a31712a <=( A167  and  A168 );
 a31713a <=( A169  and  a31712a );
 a31717a <=( A202  and  (not A201) );
 a31718a <=( (not A166)  and  a31717a );
 a31719a <=( a31718a  and  a31713a );
 a31723a <=( (not A298)  and  A269 );
 a31724a <=( (not A267)  and  a31723a );
 a31728a <=( A301  and  A300 );
 a31729a <=( A299  and  a31728a );
 a31730a <=( a31729a  and  a31724a );
 a31734a <=( A167  and  A168 );
 a31735a <=( A169  and  a31734a );
 a31739a <=( A202  and  (not A201) );
 a31740a <=( (not A166)  and  a31739a );
 a31741a <=( a31740a  and  a31735a );
 a31745a <=( (not A298)  and  A269 );
 a31746a <=( (not A267)  and  a31745a );
 a31750a <=( A302  and  A300 );
 a31751a <=( A299  and  a31750a );
 a31752a <=( a31751a  and  a31746a );
 a31756a <=( A167  and  A168 );
 a31757a <=( A169  and  a31756a );
 a31761a <=( A202  and  (not A201) );
 a31762a <=( (not A166)  and  a31761a );
 a31763a <=( a31762a  and  a31757a );
 a31767a <=( A298  and  A266 );
 a31768a <=( A265  and  a31767a );
 a31772a <=( A301  and  A300 );
 a31773a <=( (not A299)  and  a31772a );
 a31774a <=( a31773a  and  a31768a );
 a31778a <=( A167  and  A168 );
 a31779a <=( A169  and  a31778a );
 a31783a <=( A202  and  (not A201) );
 a31784a <=( (not A166)  and  a31783a );
 a31785a <=( a31784a  and  a31779a );
 a31789a <=( A298  and  A266 );
 a31790a <=( A265  and  a31789a );
 a31794a <=( A302  and  A300 );
 a31795a <=( (not A299)  and  a31794a );
 a31796a <=( a31795a  and  a31790a );
 a31800a <=( A167  and  A168 );
 a31801a <=( A169  and  a31800a );
 a31805a <=( A202  and  (not A201) );
 a31806a <=( (not A166)  and  a31805a );
 a31807a <=( a31806a  and  a31801a );
 a31811a <=( (not A298)  and  A266 );
 a31812a <=( A265  and  a31811a );
 a31816a <=( A301  and  A300 );
 a31817a <=( A299  and  a31816a );
 a31818a <=( a31817a  and  a31812a );
 a31822a <=( A167  and  A168 );
 a31823a <=( A169  and  a31822a );
 a31827a <=( A202  and  (not A201) );
 a31828a <=( (not A166)  and  a31827a );
 a31829a <=( a31828a  and  a31823a );
 a31833a <=( (not A298)  and  A266 );
 a31834a <=( A265  and  a31833a );
 a31838a <=( A302  and  A300 );
 a31839a <=( A299  and  a31838a );
 a31840a <=( a31839a  and  a31834a );
 a31844a <=( A167  and  A168 );
 a31845a <=( A169  and  a31844a );
 a31849a <=( A202  and  (not A201) );
 a31850a <=( (not A166)  and  a31849a );
 a31851a <=( a31850a  and  a31845a );
 a31855a <=( A298  and  (not A266) );
 a31856a <=( (not A265)  and  a31855a );
 a31860a <=( A301  and  A300 );
 a31861a <=( (not A299)  and  a31860a );
 a31862a <=( a31861a  and  a31856a );
 a31866a <=( A167  and  A168 );
 a31867a <=( A169  and  a31866a );
 a31871a <=( A202  and  (not A201) );
 a31872a <=( (not A166)  and  a31871a );
 a31873a <=( a31872a  and  a31867a );
 a31877a <=( A298  and  (not A266) );
 a31878a <=( (not A265)  and  a31877a );
 a31882a <=( A302  and  A300 );
 a31883a <=( (not A299)  and  a31882a );
 a31884a <=( a31883a  and  a31878a );
 a31888a <=( A167  and  A168 );
 a31889a <=( A169  and  a31888a );
 a31893a <=( A202  and  (not A201) );
 a31894a <=( (not A166)  and  a31893a );
 a31895a <=( a31894a  and  a31889a );
 a31899a <=( (not A298)  and  (not A266) );
 a31900a <=( (not A265)  and  a31899a );
 a31904a <=( A301  and  A300 );
 a31905a <=( A299  and  a31904a );
 a31906a <=( a31905a  and  a31900a );
 a31910a <=( A167  and  A168 );
 a31911a <=( A169  and  a31910a );
 a31915a <=( A202  and  (not A201) );
 a31916a <=( (not A166)  and  a31915a );
 a31917a <=( a31916a  and  a31911a );
 a31921a <=( (not A298)  and  (not A266) );
 a31922a <=( (not A265)  and  a31921a );
 a31926a <=( A302  and  A300 );
 a31927a <=( A299  and  a31926a );
 a31928a <=( a31927a  and  a31922a );
 a31932a <=( A167  and  A168 );
 a31933a <=( A169  and  a31932a );
 a31937a <=( A203  and  (not A201) );
 a31938a <=( (not A166)  and  a31937a );
 a31939a <=( a31938a  and  a31933a );
 a31943a <=( A298  and  A268 );
 a31944a <=( (not A267)  and  a31943a );
 a31948a <=( A301  and  A300 );
 a31949a <=( (not A299)  and  a31948a );
 a31950a <=( a31949a  and  a31944a );
 a31954a <=( A167  and  A168 );
 a31955a <=( A169  and  a31954a );
 a31959a <=( A203  and  (not A201) );
 a31960a <=( (not A166)  and  a31959a );
 a31961a <=( a31960a  and  a31955a );
 a31965a <=( A298  and  A268 );
 a31966a <=( (not A267)  and  a31965a );
 a31970a <=( A302  and  A300 );
 a31971a <=( (not A299)  and  a31970a );
 a31972a <=( a31971a  and  a31966a );
 a31976a <=( A167  and  A168 );
 a31977a <=( A169  and  a31976a );
 a31981a <=( A203  and  (not A201) );
 a31982a <=( (not A166)  and  a31981a );
 a31983a <=( a31982a  and  a31977a );
 a31987a <=( (not A298)  and  A268 );
 a31988a <=( (not A267)  and  a31987a );
 a31992a <=( A301  and  A300 );
 a31993a <=( A299  and  a31992a );
 a31994a <=( a31993a  and  a31988a );
 a31998a <=( A167  and  A168 );
 a31999a <=( A169  and  a31998a );
 a32003a <=( A203  and  (not A201) );
 a32004a <=( (not A166)  and  a32003a );
 a32005a <=( a32004a  and  a31999a );
 a32009a <=( (not A298)  and  A268 );
 a32010a <=( (not A267)  and  a32009a );
 a32014a <=( A302  and  A300 );
 a32015a <=( A299  and  a32014a );
 a32016a <=( a32015a  and  a32010a );
 a32020a <=( A167  and  A168 );
 a32021a <=( A169  and  a32020a );
 a32025a <=( A203  and  (not A201) );
 a32026a <=( (not A166)  and  a32025a );
 a32027a <=( a32026a  and  a32021a );
 a32031a <=( A298  and  A269 );
 a32032a <=( (not A267)  and  a32031a );
 a32036a <=( A301  and  A300 );
 a32037a <=( (not A299)  and  a32036a );
 a32038a <=( a32037a  and  a32032a );
 a32042a <=( A167  and  A168 );
 a32043a <=( A169  and  a32042a );
 a32047a <=( A203  and  (not A201) );
 a32048a <=( (not A166)  and  a32047a );
 a32049a <=( a32048a  and  a32043a );
 a32053a <=( A298  and  A269 );
 a32054a <=( (not A267)  and  a32053a );
 a32058a <=( A302  and  A300 );
 a32059a <=( (not A299)  and  a32058a );
 a32060a <=( a32059a  and  a32054a );
 a32064a <=( A167  and  A168 );
 a32065a <=( A169  and  a32064a );
 a32069a <=( A203  and  (not A201) );
 a32070a <=( (not A166)  and  a32069a );
 a32071a <=( a32070a  and  a32065a );
 a32075a <=( (not A298)  and  A269 );
 a32076a <=( (not A267)  and  a32075a );
 a32080a <=( A301  and  A300 );
 a32081a <=( A299  and  a32080a );
 a32082a <=( a32081a  and  a32076a );
 a32086a <=( A167  and  A168 );
 a32087a <=( A169  and  a32086a );
 a32091a <=( A203  and  (not A201) );
 a32092a <=( (not A166)  and  a32091a );
 a32093a <=( a32092a  and  a32087a );
 a32097a <=( (not A298)  and  A269 );
 a32098a <=( (not A267)  and  a32097a );
 a32102a <=( A302  and  A300 );
 a32103a <=( A299  and  a32102a );
 a32104a <=( a32103a  and  a32098a );
 a32108a <=( A167  and  A168 );
 a32109a <=( A169  and  a32108a );
 a32113a <=( A203  and  (not A201) );
 a32114a <=( (not A166)  and  a32113a );
 a32115a <=( a32114a  and  a32109a );
 a32119a <=( A298  and  A266 );
 a32120a <=( A265  and  a32119a );
 a32124a <=( A301  and  A300 );
 a32125a <=( (not A299)  and  a32124a );
 a32126a <=( a32125a  and  a32120a );
 a32130a <=( A167  and  A168 );
 a32131a <=( A169  and  a32130a );
 a32135a <=( A203  and  (not A201) );
 a32136a <=( (not A166)  and  a32135a );
 a32137a <=( a32136a  and  a32131a );
 a32141a <=( A298  and  A266 );
 a32142a <=( A265  and  a32141a );
 a32146a <=( A302  and  A300 );
 a32147a <=( (not A299)  and  a32146a );
 a32148a <=( a32147a  and  a32142a );
 a32152a <=( A167  and  A168 );
 a32153a <=( A169  and  a32152a );
 a32157a <=( A203  and  (not A201) );
 a32158a <=( (not A166)  and  a32157a );
 a32159a <=( a32158a  and  a32153a );
 a32163a <=( (not A298)  and  A266 );
 a32164a <=( A265  and  a32163a );
 a32168a <=( A301  and  A300 );
 a32169a <=( A299  and  a32168a );
 a32170a <=( a32169a  and  a32164a );
 a32174a <=( A167  and  A168 );
 a32175a <=( A169  and  a32174a );
 a32179a <=( A203  and  (not A201) );
 a32180a <=( (not A166)  and  a32179a );
 a32181a <=( a32180a  and  a32175a );
 a32185a <=( (not A298)  and  A266 );
 a32186a <=( A265  and  a32185a );
 a32190a <=( A302  and  A300 );
 a32191a <=( A299  and  a32190a );
 a32192a <=( a32191a  and  a32186a );
 a32196a <=( A167  and  A168 );
 a32197a <=( A169  and  a32196a );
 a32201a <=( A203  and  (not A201) );
 a32202a <=( (not A166)  and  a32201a );
 a32203a <=( a32202a  and  a32197a );
 a32207a <=( A298  and  (not A266) );
 a32208a <=( (not A265)  and  a32207a );
 a32212a <=( A301  and  A300 );
 a32213a <=( (not A299)  and  a32212a );
 a32214a <=( a32213a  and  a32208a );
 a32218a <=( A167  and  A168 );
 a32219a <=( A169  and  a32218a );
 a32223a <=( A203  and  (not A201) );
 a32224a <=( (not A166)  and  a32223a );
 a32225a <=( a32224a  and  a32219a );
 a32229a <=( A298  and  (not A266) );
 a32230a <=( (not A265)  and  a32229a );
 a32234a <=( A302  and  A300 );
 a32235a <=( (not A299)  and  a32234a );
 a32236a <=( a32235a  and  a32230a );
 a32240a <=( A167  and  A168 );
 a32241a <=( A169  and  a32240a );
 a32245a <=( A203  and  (not A201) );
 a32246a <=( (not A166)  and  a32245a );
 a32247a <=( a32246a  and  a32241a );
 a32251a <=( (not A298)  and  (not A266) );
 a32252a <=( (not A265)  and  a32251a );
 a32256a <=( A301  and  A300 );
 a32257a <=( A299  and  a32256a );
 a32258a <=( a32257a  and  a32252a );
 a32262a <=( A167  and  A168 );
 a32263a <=( A169  and  a32262a );
 a32267a <=( A203  and  (not A201) );
 a32268a <=( (not A166)  and  a32267a );
 a32269a <=( a32268a  and  a32263a );
 a32273a <=( (not A298)  and  (not A266) );
 a32274a <=( (not A265)  and  a32273a );
 a32278a <=( A302  and  A300 );
 a32279a <=( A299  and  a32278a );
 a32280a <=( a32279a  and  a32274a );
 a32284a <=( A167  and  A168 );
 a32285a <=( A169  and  a32284a );
 a32289a <=( A200  and  A199 );
 a32290a <=( (not A166)  and  a32289a );
 a32291a <=( a32290a  and  a32285a );
 a32295a <=( A298  and  A268 );
 a32296a <=( (not A267)  and  a32295a );
 a32300a <=( A301  and  A300 );
 a32301a <=( (not A299)  and  a32300a );
 a32302a <=( a32301a  and  a32296a );
 a32306a <=( A167  and  A168 );
 a32307a <=( A169  and  a32306a );
 a32311a <=( A200  and  A199 );
 a32312a <=( (not A166)  and  a32311a );
 a32313a <=( a32312a  and  a32307a );
 a32317a <=( A298  and  A268 );
 a32318a <=( (not A267)  and  a32317a );
 a32322a <=( A302  and  A300 );
 a32323a <=( (not A299)  and  a32322a );
 a32324a <=( a32323a  and  a32318a );
 a32328a <=( A167  and  A168 );
 a32329a <=( A169  and  a32328a );
 a32333a <=( A200  and  A199 );
 a32334a <=( (not A166)  and  a32333a );
 a32335a <=( a32334a  and  a32329a );
 a32339a <=( (not A298)  and  A268 );
 a32340a <=( (not A267)  and  a32339a );
 a32344a <=( A301  and  A300 );
 a32345a <=( A299  and  a32344a );
 a32346a <=( a32345a  and  a32340a );
 a32350a <=( A167  and  A168 );
 a32351a <=( A169  and  a32350a );
 a32355a <=( A200  and  A199 );
 a32356a <=( (not A166)  and  a32355a );
 a32357a <=( a32356a  and  a32351a );
 a32361a <=( (not A298)  and  A268 );
 a32362a <=( (not A267)  and  a32361a );
 a32366a <=( A302  and  A300 );
 a32367a <=( A299  and  a32366a );
 a32368a <=( a32367a  and  a32362a );
 a32372a <=( A167  and  A168 );
 a32373a <=( A169  and  a32372a );
 a32377a <=( A200  and  A199 );
 a32378a <=( (not A166)  and  a32377a );
 a32379a <=( a32378a  and  a32373a );
 a32383a <=( A298  and  A269 );
 a32384a <=( (not A267)  and  a32383a );
 a32388a <=( A301  and  A300 );
 a32389a <=( (not A299)  and  a32388a );
 a32390a <=( a32389a  and  a32384a );
 a32394a <=( A167  and  A168 );
 a32395a <=( A169  and  a32394a );
 a32399a <=( A200  and  A199 );
 a32400a <=( (not A166)  and  a32399a );
 a32401a <=( a32400a  and  a32395a );
 a32405a <=( A298  and  A269 );
 a32406a <=( (not A267)  and  a32405a );
 a32410a <=( A302  and  A300 );
 a32411a <=( (not A299)  and  a32410a );
 a32412a <=( a32411a  and  a32406a );
 a32416a <=( A167  and  A168 );
 a32417a <=( A169  and  a32416a );
 a32421a <=( A200  and  A199 );
 a32422a <=( (not A166)  and  a32421a );
 a32423a <=( a32422a  and  a32417a );
 a32427a <=( (not A298)  and  A269 );
 a32428a <=( (not A267)  and  a32427a );
 a32432a <=( A301  and  A300 );
 a32433a <=( A299  and  a32432a );
 a32434a <=( a32433a  and  a32428a );
 a32438a <=( A167  and  A168 );
 a32439a <=( A169  and  a32438a );
 a32443a <=( A200  and  A199 );
 a32444a <=( (not A166)  and  a32443a );
 a32445a <=( a32444a  and  a32439a );
 a32449a <=( (not A298)  and  A269 );
 a32450a <=( (not A267)  and  a32449a );
 a32454a <=( A302  and  A300 );
 a32455a <=( A299  and  a32454a );
 a32456a <=( a32455a  and  a32450a );
 a32460a <=( A167  and  A168 );
 a32461a <=( A169  and  a32460a );
 a32465a <=( A200  and  A199 );
 a32466a <=( (not A166)  and  a32465a );
 a32467a <=( a32466a  and  a32461a );
 a32471a <=( A298  and  A266 );
 a32472a <=( A265  and  a32471a );
 a32476a <=( A301  and  A300 );
 a32477a <=( (not A299)  and  a32476a );
 a32478a <=( a32477a  and  a32472a );
 a32482a <=( A167  and  A168 );
 a32483a <=( A169  and  a32482a );
 a32487a <=( A200  and  A199 );
 a32488a <=( (not A166)  and  a32487a );
 a32489a <=( a32488a  and  a32483a );
 a32493a <=( A298  and  A266 );
 a32494a <=( A265  and  a32493a );
 a32498a <=( A302  and  A300 );
 a32499a <=( (not A299)  and  a32498a );
 a32500a <=( a32499a  and  a32494a );
 a32504a <=( A167  and  A168 );
 a32505a <=( A169  and  a32504a );
 a32509a <=( A200  and  A199 );
 a32510a <=( (not A166)  and  a32509a );
 a32511a <=( a32510a  and  a32505a );
 a32515a <=( (not A298)  and  A266 );
 a32516a <=( A265  and  a32515a );
 a32520a <=( A301  and  A300 );
 a32521a <=( A299  and  a32520a );
 a32522a <=( a32521a  and  a32516a );
 a32526a <=( A167  and  A168 );
 a32527a <=( A169  and  a32526a );
 a32531a <=( A200  and  A199 );
 a32532a <=( (not A166)  and  a32531a );
 a32533a <=( a32532a  and  a32527a );
 a32537a <=( (not A298)  and  A266 );
 a32538a <=( A265  and  a32537a );
 a32542a <=( A302  and  A300 );
 a32543a <=( A299  and  a32542a );
 a32544a <=( a32543a  and  a32538a );
 a32548a <=( A167  and  A168 );
 a32549a <=( A169  and  a32548a );
 a32553a <=( A200  and  A199 );
 a32554a <=( (not A166)  and  a32553a );
 a32555a <=( a32554a  and  a32549a );
 a32559a <=( A298  and  (not A266) );
 a32560a <=( (not A265)  and  a32559a );
 a32564a <=( A301  and  A300 );
 a32565a <=( (not A299)  and  a32564a );
 a32566a <=( a32565a  and  a32560a );
 a32570a <=( A167  and  A168 );
 a32571a <=( A169  and  a32570a );
 a32575a <=( A200  and  A199 );
 a32576a <=( (not A166)  and  a32575a );
 a32577a <=( a32576a  and  a32571a );
 a32581a <=( A298  and  (not A266) );
 a32582a <=( (not A265)  and  a32581a );
 a32586a <=( A302  and  A300 );
 a32587a <=( (not A299)  and  a32586a );
 a32588a <=( a32587a  and  a32582a );
 a32592a <=( A167  and  A168 );
 a32593a <=( A169  and  a32592a );
 a32597a <=( A200  and  A199 );
 a32598a <=( (not A166)  and  a32597a );
 a32599a <=( a32598a  and  a32593a );
 a32603a <=( (not A298)  and  (not A266) );
 a32604a <=( (not A265)  and  a32603a );
 a32608a <=( A301  and  A300 );
 a32609a <=( A299  and  a32608a );
 a32610a <=( a32609a  and  a32604a );
 a32614a <=( A167  and  A168 );
 a32615a <=( A169  and  a32614a );
 a32619a <=( A200  and  A199 );
 a32620a <=( (not A166)  and  a32619a );
 a32621a <=( a32620a  and  a32615a );
 a32625a <=( (not A298)  and  (not A266) );
 a32626a <=( (not A265)  and  a32625a );
 a32630a <=( A302  and  A300 );
 a32631a <=( A299  and  a32630a );
 a32632a <=( a32631a  and  a32626a );
 a32636a <=( A167  and  A168 );
 a32637a <=( A169  and  a32636a );
 a32641a <=( (not A200)  and  (not A199) );
 a32642a <=( (not A166)  and  a32641a );
 a32643a <=( a32642a  and  a32637a );
 a32647a <=( A298  and  A268 );
 a32648a <=( (not A267)  and  a32647a );
 a32652a <=( A301  and  A300 );
 a32653a <=( (not A299)  and  a32652a );
 a32654a <=( a32653a  and  a32648a );
 a32658a <=( A167  and  A168 );
 a32659a <=( A169  and  a32658a );
 a32663a <=( (not A200)  and  (not A199) );
 a32664a <=( (not A166)  and  a32663a );
 a32665a <=( a32664a  and  a32659a );
 a32669a <=( A298  and  A268 );
 a32670a <=( (not A267)  and  a32669a );
 a32674a <=( A302  and  A300 );
 a32675a <=( (not A299)  and  a32674a );
 a32676a <=( a32675a  and  a32670a );
 a32680a <=( A167  and  A168 );
 a32681a <=( A169  and  a32680a );
 a32685a <=( (not A200)  and  (not A199) );
 a32686a <=( (not A166)  and  a32685a );
 a32687a <=( a32686a  and  a32681a );
 a32691a <=( (not A298)  and  A268 );
 a32692a <=( (not A267)  and  a32691a );
 a32696a <=( A301  and  A300 );
 a32697a <=( A299  and  a32696a );
 a32698a <=( a32697a  and  a32692a );
 a32702a <=( A167  and  A168 );
 a32703a <=( A169  and  a32702a );
 a32707a <=( (not A200)  and  (not A199) );
 a32708a <=( (not A166)  and  a32707a );
 a32709a <=( a32708a  and  a32703a );
 a32713a <=( (not A298)  and  A268 );
 a32714a <=( (not A267)  and  a32713a );
 a32718a <=( A302  and  A300 );
 a32719a <=( A299  and  a32718a );
 a32720a <=( a32719a  and  a32714a );
 a32724a <=( A167  and  A168 );
 a32725a <=( A169  and  a32724a );
 a32729a <=( (not A200)  and  (not A199) );
 a32730a <=( (not A166)  and  a32729a );
 a32731a <=( a32730a  and  a32725a );
 a32735a <=( A298  and  A269 );
 a32736a <=( (not A267)  and  a32735a );
 a32740a <=( A301  and  A300 );
 a32741a <=( (not A299)  and  a32740a );
 a32742a <=( a32741a  and  a32736a );
 a32746a <=( A167  and  A168 );
 a32747a <=( A169  and  a32746a );
 a32751a <=( (not A200)  and  (not A199) );
 a32752a <=( (not A166)  and  a32751a );
 a32753a <=( a32752a  and  a32747a );
 a32757a <=( A298  and  A269 );
 a32758a <=( (not A267)  and  a32757a );
 a32762a <=( A302  and  A300 );
 a32763a <=( (not A299)  and  a32762a );
 a32764a <=( a32763a  and  a32758a );
 a32768a <=( A167  and  A168 );
 a32769a <=( A169  and  a32768a );
 a32773a <=( (not A200)  and  (not A199) );
 a32774a <=( (not A166)  and  a32773a );
 a32775a <=( a32774a  and  a32769a );
 a32779a <=( (not A298)  and  A269 );
 a32780a <=( (not A267)  and  a32779a );
 a32784a <=( A301  and  A300 );
 a32785a <=( A299  and  a32784a );
 a32786a <=( a32785a  and  a32780a );
 a32790a <=( A167  and  A168 );
 a32791a <=( A169  and  a32790a );
 a32795a <=( (not A200)  and  (not A199) );
 a32796a <=( (not A166)  and  a32795a );
 a32797a <=( a32796a  and  a32791a );
 a32801a <=( (not A298)  and  A269 );
 a32802a <=( (not A267)  and  a32801a );
 a32806a <=( A302  and  A300 );
 a32807a <=( A299  and  a32806a );
 a32808a <=( a32807a  and  a32802a );
 a32812a <=( A167  and  A168 );
 a32813a <=( A169  and  a32812a );
 a32817a <=( (not A200)  and  (not A199) );
 a32818a <=( (not A166)  and  a32817a );
 a32819a <=( a32818a  and  a32813a );
 a32823a <=( A298  and  A266 );
 a32824a <=( A265  and  a32823a );
 a32828a <=( A301  and  A300 );
 a32829a <=( (not A299)  and  a32828a );
 a32830a <=( a32829a  and  a32824a );
 a32834a <=( A167  and  A168 );
 a32835a <=( A169  and  a32834a );
 a32839a <=( (not A200)  and  (not A199) );
 a32840a <=( (not A166)  and  a32839a );
 a32841a <=( a32840a  and  a32835a );
 a32845a <=( A298  and  A266 );
 a32846a <=( A265  and  a32845a );
 a32850a <=( A302  and  A300 );
 a32851a <=( (not A299)  and  a32850a );
 a32852a <=( a32851a  and  a32846a );
 a32856a <=( A167  and  A168 );
 a32857a <=( A169  and  a32856a );
 a32861a <=( (not A200)  and  (not A199) );
 a32862a <=( (not A166)  and  a32861a );
 a32863a <=( a32862a  and  a32857a );
 a32867a <=( (not A298)  and  A266 );
 a32868a <=( A265  and  a32867a );
 a32872a <=( A301  and  A300 );
 a32873a <=( A299  and  a32872a );
 a32874a <=( a32873a  and  a32868a );
 a32878a <=( A167  and  A168 );
 a32879a <=( A169  and  a32878a );
 a32883a <=( (not A200)  and  (not A199) );
 a32884a <=( (not A166)  and  a32883a );
 a32885a <=( a32884a  and  a32879a );
 a32889a <=( (not A298)  and  A266 );
 a32890a <=( A265  and  a32889a );
 a32894a <=( A302  and  A300 );
 a32895a <=( A299  and  a32894a );
 a32896a <=( a32895a  and  a32890a );
 a32900a <=( A167  and  A168 );
 a32901a <=( A169  and  a32900a );
 a32905a <=( (not A200)  and  (not A199) );
 a32906a <=( (not A166)  and  a32905a );
 a32907a <=( a32906a  and  a32901a );
 a32911a <=( A298  and  (not A266) );
 a32912a <=( (not A265)  and  a32911a );
 a32916a <=( A301  and  A300 );
 a32917a <=( (not A299)  and  a32916a );
 a32918a <=( a32917a  and  a32912a );
 a32922a <=( A167  and  A168 );
 a32923a <=( A169  and  a32922a );
 a32927a <=( (not A200)  and  (not A199) );
 a32928a <=( (not A166)  and  a32927a );
 a32929a <=( a32928a  and  a32923a );
 a32933a <=( A298  and  (not A266) );
 a32934a <=( (not A265)  and  a32933a );
 a32938a <=( A302  and  A300 );
 a32939a <=( (not A299)  and  a32938a );
 a32940a <=( a32939a  and  a32934a );
 a32944a <=( A167  and  A168 );
 a32945a <=( A169  and  a32944a );
 a32949a <=( (not A200)  and  (not A199) );
 a32950a <=( (not A166)  and  a32949a );
 a32951a <=( a32950a  and  a32945a );
 a32955a <=( (not A298)  and  (not A266) );
 a32956a <=( (not A265)  and  a32955a );
 a32960a <=( A301  and  A300 );
 a32961a <=( A299  and  a32960a );
 a32962a <=( a32961a  and  a32956a );
 a32966a <=( A167  and  A168 );
 a32967a <=( A169  and  a32966a );
 a32971a <=( (not A200)  and  (not A199) );
 a32972a <=( (not A166)  and  a32971a );
 a32973a <=( a32972a  and  a32967a );
 a32977a <=( (not A298)  and  (not A266) );
 a32978a <=( (not A265)  and  a32977a );
 a32982a <=( A302  and  A300 );
 a32983a <=( A299  and  a32982a );
 a32984a <=( a32983a  and  a32978a );
 a32988a <=( (not A167)  and  A168 );
 a32989a <=( A169  and  a32988a );
 a32993a <=( A202  and  (not A201) );
 a32994a <=( A166  and  a32993a );
 a32995a <=( a32994a  and  a32989a );
 a32999a <=( A298  and  A268 );
 a33000a <=( (not A267)  and  a32999a );
 a33004a <=( A301  and  A300 );
 a33005a <=( (not A299)  and  a33004a );
 a33006a <=( a33005a  and  a33000a );
 a33010a <=( (not A167)  and  A168 );
 a33011a <=( A169  and  a33010a );
 a33015a <=( A202  and  (not A201) );
 a33016a <=( A166  and  a33015a );
 a33017a <=( a33016a  and  a33011a );
 a33021a <=( A298  and  A268 );
 a33022a <=( (not A267)  and  a33021a );
 a33026a <=( A302  and  A300 );
 a33027a <=( (not A299)  and  a33026a );
 a33028a <=( a33027a  and  a33022a );
 a33032a <=( (not A167)  and  A168 );
 a33033a <=( A169  and  a33032a );
 a33037a <=( A202  and  (not A201) );
 a33038a <=( A166  and  a33037a );
 a33039a <=( a33038a  and  a33033a );
 a33043a <=( (not A298)  and  A268 );
 a33044a <=( (not A267)  and  a33043a );
 a33048a <=( A301  and  A300 );
 a33049a <=( A299  and  a33048a );
 a33050a <=( a33049a  and  a33044a );
 a33054a <=( (not A167)  and  A168 );
 a33055a <=( A169  and  a33054a );
 a33059a <=( A202  and  (not A201) );
 a33060a <=( A166  and  a33059a );
 a33061a <=( a33060a  and  a33055a );
 a33065a <=( (not A298)  and  A268 );
 a33066a <=( (not A267)  and  a33065a );
 a33070a <=( A302  and  A300 );
 a33071a <=( A299  and  a33070a );
 a33072a <=( a33071a  and  a33066a );
 a33076a <=( (not A167)  and  A168 );
 a33077a <=( A169  and  a33076a );
 a33081a <=( A202  and  (not A201) );
 a33082a <=( A166  and  a33081a );
 a33083a <=( a33082a  and  a33077a );
 a33087a <=( A298  and  A269 );
 a33088a <=( (not A267)  and  a33087a );
 a33092a <=( A301  and  A300 );
 a33093a <=( (not A299)  and  a33092a );
 a33094a <=( a33093a  and  a33088a );
 a33098a <=( (not A167)  and  A168 );
 a33099a <=( A169  and  a33098a );
 a33103a <=( A202  and  (not A201) );
 a33104a <=( A166  and  a33103a );
 a33105a <=( a33104a  and  a33099a );
 a33109a <=( A298  and  A269 );
 a33110a <=( (not A267)  and  a33109a );
 a33114a <=( A302  and  A300 );
 a33115a <=( (not A299)  and  a33114a );
 a33116a <=( a33115a  and  a33110a );
 a33120a <=( (not A167)  and  A168 );
 a33121a <=( A169  and  a33120a );
 a33125a <=( A202  and  (not A201) );
 a33126a <=( A166  and  a33125a );
 a33127a <=( a33126a  and  a33121a );
 a33131a <=( (not A298)  and  A269 );
 a33132a <=( (not A267)  and  a33131a );
 a33136a <=( A301  and  A300 );
 a33137a <=( A299  and  a33136a );
 a33138a <=( a33137a  and  a33132a );
 a33142a <=( (not A167)  and  A168 );
 a33143a <=( A169  and  a33142a );
 a33147a <=( A202  and  (not A201) );
 a33148a <=( A166  and  a33147a );
 a33149a <=( a33148a  and  a33143a );
 a33153a <=( (not A298)  and  A269 );
 a33154a <=( (not A267)  and  a33153a );
 a33158a <=( A302  and  A300 );
 a33159a <=( A299  and  a33158a );
 a33160a <=( a33159a  and  a33154a );
 a33164a <=( (not A167)  and  A168 );
 a33165a <=( A169  and  a33164a );
 a33169a <=( A202  and  (not A201) );
 a33170a <=( A166  and  a33169a );
 a33171a <=( a33170a  and  a33165a );
 a33175a <=( A298  and  A266 );
 a33176a <=( A265  and  a33175a );
 a33180a <=( A301  and  A300 );
 a33181a <=( (not A299)  and  a33180a );
 a33182a <=( a33181a  and  a33176a );
 a33186a <=( (not A167)  and  A168 );
 a33187a <=( A169  and  a33186a );
 a33191a <=( A202  and  (not A201) );
 a33192a <=( A166  and  a33191a );
 a33193a <=( a33192a  and  a33187a );
 a33197a <=( A298  and  A266 );
 a33198a <=( A265  and  a33197a );
 a33202a <=( A302  and  A300 );
 a33203a <=( (not A299)  and  a33202a );
 a33204a <=( a33203a  and  a33198a );
 a33208a <=( (not A167)  and  A168 );
 a33209a <=( A169  and  a33208a );
 a33213a <=( A202  and  (not A201) );
 a33214a <=( A166  and  a33213a );
 a33215a <=( a33214a  and  a33209a );
 a33219a <=( (not A298)  and  A266 );
 a33220a <=( A265  and  a33219a );
 a33224a <=( A301  and  A300 );
 a33225a <=( A299  and  a33224a );
 a33226a <=( a33225a  and  a33220a );
 a33230a <=( (not A167)  and  A168 );
 a33231a <=( A169  and  a33230a );
 a33235a <=( A202  and  (not A201) );
 a33236a <=( A166  and  a33235a );
 a33237a <=( a33236a  and  a33231a );
 a33241a <=( (not A298)  and  A266 );
 a33242a <=( A265  and  a33241a );
 a33246a <=( A302  and  A300 );
 a33247a <=( A299  and  a33246a );
 a33248a <=( a33247a  and  a33242a );
 a33252a <=( (not A167)  and  A168 );
 a33253a <=( A169  and  a33252a );
 a33257a <=( A202  and  (not A201) );
 a33258a <=( A166  and  a33257a );
 a33259a <=( a33258a  and  a33253a );
 a33263a <=( A298  and  (not A266) );
 a33264a <=( (not A265)  and  a33263a );
 a33268a <=( A301  and  A300 );
 a33269a <=( (not A299)  and  a33268a );
 a33270a <=( a33269a  and  a33264a );
 a33274a <=( (not A167)  and  A168 );
 a33275a <=( A169  and  a33274a );
 a33279a <=( A202  and  (not A201) );
 a33280a <=( A166  and  a33279a );
 a33281a <=( a33280a  and  a33275a );
 a33285a <=( A298  and  (not A266) );
 a33286a <=( (not A265)  and  a33285a );
 a33290a <=( A302  and  A300 );
 a33291a <=( (not A299)  and  a33290a );
 a33292a <=( a33291a  and  a33286a );
 a33296a <=( (not A167)  and  A168 );
 a33297a <=( A169  and  a33296a );
 a33301a <=( A202  and  (not A201) );
 a33302a <=( A166  and  a33301a );
 a33303a <=( a33302a  and  a33297a );
 a33307a <=( (not A298)  and  (not A266) );
 a33308a <=( (not A265)  and  a33307a );
 a33312a <=( A301  and  A300 );
 a33313a <=( A299  and  a33312a );
 a33314a <=( a33313a  and  a33308a );
 a33318a <=( (not A167)  and  A168 );
 a33319a <=( A169  and  a33318a );
 a33323a <=( A202  and  (not A201) );
 a33324a <=( A166  and  a33323a );
 a33325a <=( a33324a  and  a33319a );
 a33329a <=( (not A298)  and  (not A266) );
 a33330a <=( (not A265)  and  a33329a );
 a33334a <=( A302  and  A300 );
 a33335a <=( A299  and  a33334a );
 a33336a <=( a33335a  and  a33330a );
 a33340a <=( (not A167)  and  A168 );
 a33341a <=( A169  and  a33340a );
 a33345a <=( A203  and  (not A201) );
 a33346a <=( A166  and  a33345a );
 a33347a <=( a33346a  and  a33341a );
 a33351a <=( A298  and  A268 );
 a33352a <=( (not A267)  and  a33351a );
 a33356a <=( A301  and  A300 );
 a33357a <=( (not A299)  and  a33356a );
 a33358a <=( a33357a  and  a33352a );
 a33362a <=( (not A167)  and  A168 );
 a33363a <=( A169  and  a33362a );
 a33367a <=( A203  and  (not A201) );
 a33368a <=( A166  and  a33367a );
 a33369a <=( a33368a  and  a33363a );
 a33373a <=( A298  and  A268 );
 a33374a <=( (not A267)  and  a33373a );
 a33378a <=( A302  and  A300 );
 a33379a <=( (not A299)  and  a33378a );
 a33380a <=( a33379a  and  a33374a );
 a33384a <=( (not A167)  and  A168 );
 a33385a <=( A169  and  a33384a );
 a33389a <=( A203  and  (not A201) );
 a33390a <=( A166  and  a33389a );
 a33391a <=( a33390a  and  a33385a );
 a33395a <=( (not A298)  and  A268 );
 a33396a <=( (not A267)  and  a33395a );
 a33400a <=( A301  and  A300 );
 a33401a <=( A299  and  a33400a );
 a33402a <=( a33401a  and  a33396a );
 a33406a <=( (not A167)  and  A168 );
 a33407a <=( A169  and  a33406a );
 a33411a <=( A203  and  (not A201) );
 a33412a <=( A166  and  a33411a );
 a33413a <=( a33412a  and  a33407a );
 a33417a <=( (not A298)  and  A268 );
 a33418a <=( (not A267)  and  a33417a );
 a33422a <=( A302  and  A300 );
 a33423a <=( A299  and  a33422a );
 a33424a <=( a33423a  and  a33418a );
 a33428a <=( (not A167)  and  A168 );
 a33429a <=( A169  and  a33428a );
 a33433a <=( A203  and  (not A201) );
 a33434a <=( A166  and  a33433a );
 a33435a <=( a33434a  and  a33429a );
 a33439a <=( A298  and  A269 );
 a33440a <=( (not A267)  and  a33439a );
 a33444a <=( A301  and  A300 );
 a33445a <=( (not A299)  and  a33444a );
 a33446a <=( a33445a  and  a33440a );
 a33450a <=( (not A167)  and  A168 );
 a33451a <=( A169  and  a33450a );
 a33455a <=( A203  and  (not A201) );
 a33456a <=( A166  and  a33455a );
 a33457a <=( a33456a  and  a33451a );
 a33461a <=( A298  and  A269 );
 a33462a <=( (not A267)  and  a33461a );
 a33466a <=( A302  and  A300 );
 a33467a <=( (not A299)  and  a33466a );
 a33468a <=( a33467a  and  a33462a );
 a33472a <=( (not A167)  and  A168 );
 a33473a <=( A169  and  a33472a );
 a33477a <=( A203  and  (not A201) );
 a33478a <=( A166  and  a33477a );
 a33479a <=( a33478a  and  a33473a );
 a33483a <=( (not A298)  and  A269 );
 a33484a <=( (not A267)  and  a33483a );
 a33488a <=( A301  and  A300 );
 a33489a <=( A299  and  a33488a );
 a33490a <=( a33489a  and  a33484a );
 a33494a <=( (not A167)  and  A168 );
 a33495a <=( A169  and  a33494a );
 a33499a <=( A203  and  (not A201) );
 a33500a <=( A166  and  a33499a );
 a33501a <=( a33500a  and  a33495a );
 a33505a <=( (not A298)  and  A269 );
 a33506a <=( (not A267)  and  a33505a );
 a33510a <=( A302  and  A300 );
 a33511a <=( A299  and  a33510a );
 a33512a <=( a33511a  and  a33506a );
 a33516a <=( (not A167)  and  A168 );
 a33517a <=( A169  and  a33516a );
 a33521a <=( A203  and  (not A201) );
 a33522a <=( A166  and  a33521a );
 a33523a <=( a33522a  and  a33517a );
 a33527a <=( A298  and  A266 );
 a33528a <=( A265  and  a33527a );
 a33532a <=( A301  and  A300 );
 a33533a <=( (not A299)  and  a33532a );
 a33534a <=( a33533a  and  a33528a );
 a33538a <=( (not A167)  and  A168 );
 a33539a <=( A169  and  a33538a );
 a33543a <=( A203  and  (not A201) );
 a33544a <=( A166  and  a33543a );
 a33545a <=( a33544a  and  a33539a );
 a33549a <=( A298  and  A266 );
 a33550a <=( A265  and  a33549a );
 a33554a <=( A302  and  A300 );
 a33555a <=( (not A299)  and  a33554a );
 a33556a <=( a33555a  and  a33550a );
 a33560a <=( (not A167)  and  A168 );
 a33561a <=( A169  and  a33560a );
 a33565a <=( A203  and  (not A201) );
 a33566a <=( A166  and  a33565a );
 a33567a <=( a33566a  and  a33561a );
 a33571a <=( (not A298)  and  A266 );
 a33572a <=( A265  and  a33571a );
 a33576a <=( A301  and  A300 );
 a33577a <=( A299  and  a33576a );
 a33578a <=( a33577a  and  a33572a );
 a33582a <=( (not A167)  and  A168 );
 a33583a <=( A169  and  a33582a );
 a33587a <=( A203  and  (not A201) );
 a33588a <=( A166  and  a33587a );
 a33589a <=( a33588a  and  a33583a );
 a33593a <=( (not A298)  and  A266 );
 a33594a <=( A265  and  a33593a );
 a33598a <=( A302  and  A300 );
 a33599a <=( A299  and  a33598a );
 a33600a <=( a33599a  and  a33594a );
 a33604a <=( (not A167)  and  A168 );
 a33605a <=( A169  and  a33604a );
 a33609a <=( A203  and  (not A201) );
 a33610a <=( A166  and  a33609a );
 a33611a <=( a33610a  and  a33605a );
 a33615a <=( A298  and  (not A266) );
 a33616a <=( (not A265)  and  a33615a );
 a33620a <=( A301  and  A300 );
 a33621a <=( (not A299)  and  a33620a );
 a33622a <=( a33621a  and  a33616a );
 a33626a <=( (not A167)  and  A168 );
 a33627a <=( A169  and  a33626a );
 a33631a <=( A203  and  (not A201) );
 a33632a <=( A166  and  a33631a );
 a33633a <=( a33632a  and  a33627a );
 a33637a <=( A298  and  (not A266) );
 a33638a <=( (not A265)  and  a33637a );
 a33642a <=( A302  and  A300 );
 a33643a <=( (not A299)  and  a33642a );
 a33644a <=( a33643a  and  a33638a );
 a33648a <=( (not A167)  and  A168 );
 a33649a <=( A169  and  a33648a );
 a33653a <=( A203  and  (not A201) );
 a33654a <=( A166  and  a33653a );
 a33655a <=( a33654a  and  a33649a );
 a33659a <=( (not A298)  and  (not A266) );
 a33660a <=( (not A265)  and  a33659a );
 a33664a <=( A301  and  A300 );
 a33665a <=( A299  and  a33664a );
 a33666a <=( a33665a  and  a33660a );
 a33670a <=( (not A167)  and  A168 );
 a33671a <=( A169  and  a33670a );
 a33675a <=( A203  and  (not A201) );
 a33676a <=( A166  and  a33675a );
 a33677a <=( a33676a  and  a33671a );
 a33681a <=( (not A298)  and  (not A266) );
 a33682a <=( (not A265)  and  a33681a );
 a33686a <=( A302  and  A300 );
 a33687a <=( A299  and  a33686a );
 a33688a <=( a33687a  and  a33682a );
 a33692a <=( (not A167)  and  A168 );
 a33693a <=( A169  and  a33692a );
 a33697a <=( A200  and  A199 );
 a33698a <=( A166  and  a33697a );
 a33699a <=( a33698a  and  a33693a );
 a33703a <=( A298  and  A268 );
 a33704a <=( (not A267)  and  a33703a );
 a33708a <=( A301  and  A300 );
 a33709a <=( (not A299)  and  a33708a );
 a33710a <=( a33709a  and  a33704a );
 a33714a <=( (not A167)  and  A168 );
 a33715a <=( A169  and  a33714a );
 a33719a <=( A200  and  A199 );
 a33720a <=( A166  and  a33719a );
 a33721a <=( a33720a  and  a33715a );
 a33725a <=( A298  and  A268 );
 a33726a <=( (not A267)  and  a33725a );
 a33730a <=( A302  and  A300 );
 a33731a <=( (not A299)  and  a33730a );
 a33732a <=( a33731a  and  a33726a );
 a33736a <=( (not A167)  and  A168 );
 a33737a <=( A169  and  a33736a );
 a33741a <=( A200  and  A199 );
 a33742a <=( A166  and  a33741a );
 a33743a <=( a33742a  and  a33737a );
 a33747a <=( (not A298)  and  A268 );
 a33748a <=( (not A267)  and  a33747a );
 a33752a <=( A301  and  A300 );
 a33753a <=( A299  and  a33752a );
 a33754a <=( a33753a  and  a33748a );
 a33758a <=( (not A167)  and  A168 );
 a33759a <=( A169  and  a33758a );
 a33763a <=( A200  and  A199 );
 a33764a <=( A166  and  a33763a );
 a33765a <=( a33764a  and  a33759a );
 a33769a <=( (not A298)  and  A268 );
 a33770a <=( (not A267)  and  a33769a );
 a33774a <=( A302  and  A300 );
 a33775a <=( A299  and  a33774a );
 a33776a <=( a33775a  and  a33770a );
 a33780a <=( (not A167)  and  A168 );
 a33781a <=( A169  and  a33780a );
 a33785a <=( A200  and  A199 );
 a33786a <=( A166  and  a33785a );
 a33787a <=( a33786a  and  a33781a );
 a33791a <=( A298  and  A269 );
 a33792a <=( (not A267)  and  a33791a );
 a33796a <=( A301  and  A300 );
 a33797a <=( (not A299)  and  a33796a );
 a33798a <=( a33797a  and  a33792a );
 a33802a <=( (not A167)  and  A168 );
 a33803a <=( A169  and  a33802a );
 a33807a <=( A200  and  A199 );
 a33808a <=( A166  and  a33807a );
 a33809a <=( a33808a  and  a33803a );
 a33813a <=( A298  and  A269 );
 a33814a <=( (not A267)  and  a33813a );
 a33818a <=( A302  and  A300 );
 a33819a <=( (not A299)  and  a33818a );
 a33820a <=( a33819a  and  a33814a );
 a33824a <=( (not A167)  and  A168 );
 a33825a <=( A169  and  a33824a );
 a33829a <=( A200  and  A199 );
 a33830a <=( A166  and  a33829a );
 a33831a <=( a33830a  and  a33825a );
 a33835a <=( (not A298)  and  A269 );
 a33836a <=( (not A267)  and  a33835a );
 a33840a <=( A301  and  A300 );
 a33841a <=( A299  and  a33840a );
 a33842a <=( a33841a  and  a33836a );
 a33846a <=( (not A167)  and  A168 );
 a33847a <=( A169  and  a33846a );
 a33851a <=( A200  and  A199 );
 a33852a <=( A166  and  a33851a );
 a33853a <=( a33852a  and  a33847a );
 a33857a <=( (not A298)  and  A269 );
 a33858a <=( (not A267)  and  a33857a );
 a33862a <=( A302  and  A300 );
 a33863a <=( A299  and  a33862a );
 a33864a <=( a33863a  and  a33858a );
 a33868a <=( (not A167)  and  A168 );
 a33869a <=( A169  and  a33868a );
 a33873a <=( A200  and  A199 );
 a33874a <=( A166  and  a33873a );
 a33875a <=( a33874a  and  a33869a );
 a33879a <=( A298  and  A266 );
 a33880a <=( A265  and  a33879a );
 a33884a <=( A301  and  A300 );
 a33885a <=( (not A299)  and  a33884a );
 a33886a <=( a33885a  and  a33880a );
 a33890a <=( (not A167)  and  A168 );
 a33891a <=( A169  and  a33890a );
 a33895a <=( A200  and  A199 );
 a33896a <=( A166  and  a33895a );
 a33897a <=( a33896a  and  a33891a );
 a33901a <=( A298  and  A266 );
 a33902a <=( A265  and  a33901a );
 a33906a <=( A302  and  A300 );
 a33907a <=( (not A299)  and  a33906a );
 a33908a <=( a33907a  and  a33902a );
 a33912a <=( (not A167)  and  A168 );
 a33913a <=( A169  and  a33912a );
 a33917a <=( A200  and  A199 );
 a33918a <=( A166  and  a33917a );
 a33919a <=( a33918a  and  a33913a );
 a33923a <=( (not A298)  and  A266 );
 a33924a <=( A265  and  a33923a );
 a33928a <=( A301  and  A300 );
 a33929a <=( A299  and  a33928a );
 a33930a <=( a33929a  and  a33924a );
 a33934a <=( (not A167)  and  A168 );
 a33935a <=( A169  and  a33934a );
 a33939a <=( A200  and  A199 );
 a33940a <=( A166  and  a33939a );
 a33941a <=( a33940a  and  a33935a );
 a33945a <=( (not A298)  and  A266 );
 a33946a <=( A265  and  a33945a );
 a33950a <=( A302  and  A300 );
 a33951a <=( A299  and  a33950a );
 a33952a <=( a33951a  and  a33946a );
 a33956a <=( (not A167)  and  A168 );
 a33957a <=( A169  and  a33956a );
 a33961a <=( A200  and  A199 );
 a33962a <=( A166  and  a33961a );
 a33963a <=( a33962a  and  a33957a );
 a33967a <=( A298  and  (not A266) );
 a33968a <=( (not A265)  and  a33967a );
 a33972a <=( A301  and  A300 );
 a33973a <=( (not A299)  and  a33972a );
 a33974a <=( a33973a  and  a33968a );
 a33978a <=( (not A167)  and  A168 );
 a33979a <=( A169  and  a33978a );
 a33983a <=( A200  and  A199 );
 a33984a <=( A166  and  a33983a );
 a33985a <=( a33984a  and  a33979a );
 a33989a <=( A298  and  (not A266) );
 a33990a <=( (not A265)  and  a33989a );
 a33994a <=( A302  and  A300 );
 a33995a <=( (not A299)  and  a33994a );
 a33996a <=( a33995a  and  a33990a );
 a34000a <=( (not A167)  and  A168 );
 a34001a <=( A169  and  a34000a );
 a34005a <=( A200  and  A199 );
 a34006a <=( A166  and  a34005a );
 a34007a <=( a34006a  and  a34001a );
 a34011a <=( (not A298)  and  (not A266) );
 a34012a <=( (not A265)  and  a34011a );
 a34016a <=( A301  and  A300 );
 a34017a <=( A299  and  a34016a );
 a34018a <=( a34017a  and  a34012a );
 a34022a <=( (not A167)  and  A168 );
 a34023a <=( A169  and  a34022a );
 a34027a <=( A200  and  A199 );
 a34028a <=( A166  and  a34027a );
 a34029a <=( a34028a  and  a34023a );
 a34033a <=( (not A298)  and  (not A266) );
 a34034a <=( (not A265)  and  a34033a );
 a34038a <=( A302  and  A300 );
 a34039a <=( A299  and  a34038a );
 a34040a <=( a34039a  and  a34034a );
 a34044a <=( (not A167)  and  A168 );
 a34045a <=( A169  and  a34044a );
 a34049a <=( (not A200)  and  (not A199) );
 a34050a <=( A166  and  a34049a );
 a34051a <=( a34050a  and  a34045a );
 a34055a <=( A298  and  A268 );
 a34056a <=( (not A267)  and  a34055a );
 a34060a <=( A301  and  A300 );
 a34061a <=( (not A299)  and  a34060a );
 a34062a <=( a34061a  and  a34056a );
 a34066a <=( (not A167)  and  A168 );
 a34067a <=( A169  and  a34066a );
 a34071a <=( (not A200)  and  (not A199) );
 a34072a <=( A166  and  a34071a );
 a34073a <=( a34072a  and  a34067a );
 a34077a <=( A298  and  A268 );
 a34078a <=( (not A267)  and  a34077a );
 a34082a <=( A302  and  A300 );
 a34083a <=( (not A299)  and  a34082a );
 a34084a <=( a34083a  and  a34078a );
 a34088a <=( (not A167)  and  A168 );
 a34089a <=( A169  and  a34088a );
 a34093a <=( (not A200)  and  (not A199) );
 a34094a <=( A166  and  a34093a );
 a34095a <=( a34094a  and  a34089a );
 a34099a <=( (not A298)  and  A268 );
 a34100a <=( (not A267)  and  a34099a );
 a34104a <=( A301  and  A300 );
 a34105a <=( A299  and  a34104a );
 a34106a <=( a34105a  and  a34100a );
 a34110a <=( (not A167)  and  A168 );
 a34111a <=( A169  and  a34110a );
 a34115a <=( (not A200)  and  (not A199) );
 a34116a <=( A166  and  a34115a );
 a34117a <=( a34116a  and  a34111a );
 a34121a <=( (not A298)  and  A268 );
 a34122a <=( (not A267)  and  a34121a );
 a34126a <=( A302  and  A300 );
 a34127a <=( A299  and  a34126a );
 a34128a <=( a34127a  and  a34122a );
 a34132a <=( (not A167)  and  A168 );
 a34133a <=( A169  and  a34132a );
 a34137a <=( (not A200)  and  (not A199) );
 a34138a <=( A166  and  a34137a );
 a34139a <=( a34138a  and  a34133a );
 a34143a <=( A298  and  A269 );
 a34144a <=( (not A267)  and  a34143a );
 a34148a <=( A301  and  A300 );
 a34149a <=( (not A299)  and  a34148a );
 a34150a <=( a34149a  and  a34144a );
 a34154a <=( (not A167)  and  A168 );
 a34155a <=( A169  and  a34154a );
 a34159a <=( (not A200)  and  (not A199) );
 a34160a <=( A166  and  a34159a );
 a34161a <=( a34160a  and  a34155a );
 a34165a <=( A298  and  A269 );
 a34166a <=( (not A267)  and  a34165a );
 a34170a <=( A302  and  A300 );
 a34171a <=( (not A299)  and  a34170a );
 a34172a <=( a34171a  and  a34166a );
 a34176a <=( (not A167)  and  A168 );
 a34177a <=( A169  and  a34176a );
 a34181a <=( (not A200)  and  (not A199) );
 a34182a <=( A166  and  a34181a );
 a34183a <=( a34182a  and  a34177a );
 a34187a <=( (not A298)  and  A269 );
 a34188a <=( (not A267)  and  a34187a );
 a34192a <=( A301  and  A300 );
 a34193a <=( A299  and  a34192a );
 a34194a <=( a34193a  and  a34188a );
 a34198a <=( (not A167)  and  A168 );
 a34199a <=( A169  and  a34198a );
 a34203a <=( (not A200)  and  (not A199) );
 a34204a <=( A166  and  a34203a );
 a34205a <=( a34204a  and  a34199a );
 a34209a <=( (not A298)  and  A269 );
 a34210a <=( (not A267)  and  a34209a );
 a34214a <=( A302  and  A300 );
 a34215a <=( A299  and  a34214a );
 a34216a <=( a34215a  and  a34210a );
 a34220a <=( (not A167)  and  A168 );
 a34221a <=( A169  and  a34220a );
 a34225a <=( (not A200)  and  (not A199) );
 a34226a <=( A166  and  a34225a );
 a34227a <=( a34226a  and  a34221a );
 a34231a <=( A298  and  A266 );
 a34232a <=( A265  and  a34231a );
 a34236a <=( A301  and  A300 );
 a34237a <=( (not A299)  and  a34236a );
 a34238a <=( a34237a  and  a34232a );
 a34242a <=( (not A167)  and  A168 );
 a34243a <=( A169  and  a34242a );
 a34247a <=( (not A200)  and  (not A199) );
 a34248a <=( A166  and  a34247a );
 a34249a <=( a34248a  and  a34243a );
 a34253a <=( A298  and  A266 );
 a34254a <=( A265  and  a34253a );
 a34258a <=( A302  and  A300 );
 a34259a <=( (not A299)  and  a34258a );
 a34260a <=( a34259a  and  a34254a );
 a34264a <=( (not A167)  and  A168 );
 a34265a <=( A169  and  a34264a );
 a34269a <=( (not A200)  and  (not A199) );
 a34270a <=( A166  and  a34269a );
 a34271a <=( a34270a  and  a34265a );
 a34275a <=( (not A298)  and  A266 );
 a34276a <=( A265  and  a34275a );
 a34280a <=( A301  and  A300 );
 a34281a <=( A299  and  a34280a );
 a34282a <=( a34281a  and  a34276a );
 a34286a <=( (not A167)  and  A168 );
 a34287a <=( A169  and  a34286a );
 a34291a <=( (not A200)  and  (not A199) );
 a34292a <=( A166  and  a34291a );
 a34293a <=( a34292a  and  a34287a );
 a34297a <=( (not A298)  and  A266 );
 a34298a <=( A265  and  a34297a );
 a34302a <=( A302  and  A300 );
 a34303a <=( A299  and  a34302a );
 a34304a <=( a34303a  and  a34298a );
 a34308a <=( (not A167)  and  A168 );
 a34309a <=( A169  and  a34308a );
 a34313a <=( (not A200)  and  (not A199) );
 a34314a <=( A166  and  a34313a );
 a34315a <=( a34314a  and  a34309a );
 a34319a <=( A298  and  (not A266) );
 a34320a <=( (not A265)  and  a34319a );
 a34324a <=( A301  and  A300 );
 a34325a <=( (not A299)  and  a34324a );
 a34326a <=( a34325a  and  a34320a );
 a34330a <=( (not A167)  and  A168 );
 a34331a <=( A169  and  a34330a );
 a34335a <=( (not A200)  and  (not A199) );
 a34336a <=( A166  and  a34335a );
 a34337a <=( a34336a  and  a34331a );
 a34341a <=( A298  and  (not A266) );
 a34342a <=( (not A265)  and  a34341a );
 a34346a <=( A302  and  A300 );
 a34347a <=( (not A299)  and  a34346a );
 a34348a <=( a34347a  and  a34342a );
 a34352a <=( (not A167)  and  A168 );
 a34353a <=( A169  and  a34352a );
 a34357a <=( (not A200)  and  (not A199) );
 a34358a <=( A166  and  a34357a );
 a34359a <=( a34358a  and  a34353a );
 a34363a <=( (not A298)  and  (not A266) );
 a34364a <=( (not A265)  and  a34363a );
 a34368a <=( A301  and  A300 );
 a34369a <=( A299  and  a34368a );
 a34370a <=( a34369a  and  a34364a );
 a34374a <=( (not A167)  and  A168 );
 a34375a <=( A169  and  a34374a );
 a34379a <=( (not A200)  and  (not A199) );
 a34380a <=( A166  and  a34379a );
 a34381a <=( a34380a  and  a34375a );
 a34385a <=( (not A298)  and  (not A266) );
 a34386a <=( (not A265)  and  a34385a );
 a34390a <=( A302  and  A300 );
 a34391a <=( A299  and  a34390a );
 a34392a <=( a34391a  and  a34386a );
 a34396a <=( A201  and  (not A168) );
 a34397a <=( A169  and  a34396a );
 a34401a <=( (not A265)  and  (not A203) );
 a34402a <=( (not A202)  and  a34401a );
 a34403a <=( a34402a  and  a34397a );
 a34407a <=( A268  and  A267 );
 a34408a <=( A266  and  a34407a );
 a34412a <=( (not A302)  and  (not A301) );
 a34413a <=( A300  and  a34412a );
 a34414a <=( a34413a  and  a34408a );
 a34418a <=( A201  and  (not A168) );
 a34419a <=( A169  and  a34418a );
 a34423a <=( (not A265)  and  (not A203) );
 a34424a <=( (not A202)  and  a34423a );
 a34425a <=( a34424a  and  a34419a );
 a34429a <=( A269  and  A267 );
 a34430a <=( A266  and  a34429a );
 a34434a <=( (not A302)  and  (not A301) );
 a34435a <=( A300  and  a34434a );
 a34436a <=( a34435a  and  a34430a );
 a34440a <=( A201  and  (not A168) );
 a34441a <=( A169  and  a34440a );
 a34445a <=( (not A265)  and  (not A203) );
 a34446a <=( (not A202)  and  a34445a );
 a34447a <=( a34446a  and  a34441a );
 a34451a <=( (not A268)  and  (not A267) );
 a34452a <=( A266  and  a34451a );
 a34456a <=( A301  and  (not A300) );
 a34457a <=( (not A269)  and  a34456a );
 a34458a <=( a34457a  and  a34452a );
 a34462a <=( A201  and  (not A168) );
 a34463a <=( A169  and  a34462a );
 a34467a <=( (not A265)  and  (not A203) );
 a34468a <=( (not A202)  and  a34467a );
 a34469a <=( a34468a  and  a34463a );
 a34473a <=( (not A268)  and  (not A267) );
 a34474a <=( A266  and  a34473a );
 a34478a <=( A302  and  (not A300) );
 a34479a <=( (not A269)  and  a34478a );
 a34480a <=( a34479a  and  a34474a );
 a34484a <=( A201  and  (not A168) );
 a34485a <=( A169  and  a34484a );
 a34489a <=( (not A265)  and  (not A203) );
 a34490a <=( (not A202)  and  a34489a );
 a34491a <=( a34490a  and  a34485a );
 a34495a <=( (not A268)  and  (not A267) );
 a34496a <=( A266  and  a34495a );
 a34500a <=( A299  and  A298 );
 a34501a <=( (not A269)  and  a34500a );
 a34502a <=( a34501a  and  a34496a );
 a34506a <=( A201  and  (not A168) );
 a34507a <=( A169  and  a34506a );
 a34511a <=( (not A265)  and  (not A203) );
 a34512a <=( (not A202)  and  a34511a );
 a34513a <=( a34512a  and  a34507a );
 a34517a <=( (not A268)  and  (not A267) );
 a34518a <=( A266  and  a34517a );
 a34522a <=( (not A299)  and  (not A298) );
 a34523a <=( (not A269)  and  a34522a );
 a34524a <=( a34523a  and  a34518a );
 a34528a <=( A201  and  (not A168) );
 a34529a <=( A169  and  a34528a );
 a34533a <=( A265  and  (not A203) );
 a34534a <=( (not A202)  and  a34533a );
 a34535a <=( a34534a  and  a34529a );
 a34539a <=( A268  and  A267 );
 a34540a <=( (not A266)  and  a34539a );
 a34544a <=( (not A302)  and  (not A301) );
 a34545a <=( A300  and  a34544a );
 a34546a <=( a34545a  and  a34540a );
 a34550a <=( A201  and  (not A168) );
 a34551a <=( A169  and  a34550a );
 a34555a <=( A265  and  (not A203) );
 a34556a <=( (not A202)  and  a34555a );
 a34557a <=( a34556a  and  a34551a );
 a34561a <=( A269  and  A267 );
 a34562a <=( (not A266)  and  a34561a );
 a34566a <=( (not A302)  and  (not A301) );
 a34567a <=( A300  and  a34566a );
 a34568a <=( a34567a  and  a34562a );
 a34572a <=( A201  and  (not A168) );
 a34573a <=( A169  and  a34572a );
 a34577a <=( A265  and  (not A203) );
 a34578a <=( (not A202)  and  a34577a );
 a34579a <=( a34578a  and  a34573a );
 a34583a <=( (not A268)  and  (not A267) );
 a34584a <=( (not A266)  and  a34583a );
 a34588a <=( A301  and  (not A300) );
 a34589a <=( (not A269)  and  a34588a );
 a34590a <=( a34589a  and  a34584a );
 a34594a <=( A201  and  (not A168) );
 a34595a <=( A169  and  a34594a );
 a34599a <=( A265  and  (not A203) );
 a34600a <=( (not A202)  and  a34599a );
 a34601a <=( a34600a  and  a34595a );
 a34605a <=( (not A268)  and  (not A267) );
 a34606a <=( (not A266)  and  a34605a );
 a34610a <=( A302  and  (not A300) );
 a34611a <=( (not A269)  and  a34610a );
 a34612a <=( a34611a  and  a34606a );
 a34616a <=( A201  and  (not A168) );
 a34617a <=( A169  and  a34616a );
 a34621a <=( A265  and  (not A203) );
 a34622a <=( (not A202)  and  a34621a );
 a34623a <=( a34622a  and  a34617a );
 a34627a <=( (not A268)  and  (not A267) );
 a34628a <=( (not A266)  and  a34627a );
 a34632a <=( A299  and  A298 );
 a34633a <=( (not A269)  and  a34632a );
 a34634a <=( a34633a  and  a34628a );
 a34638a <=( A201  and  (not A168) );
 a34639a <=( A169  and  a34638a );
 a34643a <=( A265  and  (not A203) );
 a34644a <=( (not A202)  and  a34643a );
 a34645a <=( a34644a  and  a34639a );
 a34649a <=( (not A268)  and  (not A267) );
 a34650a <=( (not A266)  and  a34649a );
 a34654a <=( (not A299)  and  (not A298) );
 a34655a <=( (not A269)  and  a34654a );
 a34656a <=( a34655a  and  a34650a );
 a34660a <=( (not A201)  and  (not A168) );
 a34661a <=( A169  and  a34660a );
 a34665a <=( A266  and  (not A265) );
 a34666a <=( A202  and  a34665a );
 a34667a <=( a34666a  and  a34661a );
 a34671a <=( (not A269)  and  (not A268) );
 a34672a <=( (not A267)  and  a34671a );
 a34676a <=( (not A302)  and  (not A301) );
 a34677a <=( A300  and  a34676a );
 a34678a <=( a34677a  and  a34672a );
 a34682a <=( (not A201)  and  (not A168) );
 a34683a <=( A169  and  a34682a );
 a34687a <=( (not A266)  and  A265 );
 a34688a <=( A202  and  a34687a );
 a34689a <=( a34688a  and  a34683a );
 a34693a <=( (not A269)  and  (not A268) );
 a34694a <=( (not A267)  and  a34693a );
 a34698a <=( (not A302)  and  (not A301) );
 a34699a <=( A300  and  a34698a );
 a34700a <=( a34699a  and  a34694a );
 a34704a <=( (not A201)  and  (not A168) );
 a34705a <=( A169  and  a34704a );
 a34709a <=( A266  and  (not A265) );
 a34710a <=( A203  and  a34709a );
 a34711a <=( a34710a  and  a34705a );
 a34715a <=( (not A269)  and  (not A268) );
 a34716a <=( (not A267)  and  a34715a );
 a34720a <=( (not A302)  and  (not A301) );
 a34721a <=( A300  and  a34720a );
 a34722a <=( a34721a  and  a34716a );
 a34726a <=( (not A201)  and  (not A168) );
 a34727a <=( A169  and  a34726a );
 a34731a <=( (not A266)  and  A265 );
 a34732a <=( A203  and  a34731a );
 a34733a <=( a34732a  and  a34727a );
 a34737a <=( (not A269)  and  (not A268) );
 a34738a <=( (not A267)  and  a34737a );
 a34742a <=( (not A302)  and  (not A301) );
 a34743a <=( A300  and  a34742a );
 a34744a <=( a34743a  and  a34738a );
 a34748a <=( A199  and  (not A168) );
 a34749a <=( A169  and  a34748a );
 a34753a <=( A266  and  (not A265) );
 a34754a <=( A200  and  a34753a );
 a34755a <=( a34754a  and  a34749a );
 a34759a <=( (not A269)  and  (not A268) );
 a34760a <=( (not A267)  and  a34759a );
 a34764a <=( (not A302)  and  (not A301) );
 a34765a <=( A300  and  a34764a );
 a34766a <=( a34765a  and  a34760a );
 a34770a <=( A199  and  (not A168) );
 a34771a <=( A169  and  a34770a );
 a34775a <=( (not A266)  and  A265 );
 a34776a <=( A200  and  a34775a );
 a34777a <=( a34776a  and  a34771a );
 a34781a <=( (not A269)  and  (not A268) );
 a34782a <=( (not A267)  and  a34781a );
 a34786a <=( (not A302)  and  (not A301) );
 a34787a <=( A300  and  a34786a );
 a34788a <=( a34787a  and  a34782a );
 a34792a <=( (not A199)  and  (not A168) );
 a34793a <=( A169  and  a34792a );
 a34797a <=( A202  and  A201 );
 a34798a <=( A200  and  a34797a );
 a34799a <=( a34798a  and  a34793a );
 a34803a <=( A298  and  A268 );
 a34804a <=( (not A267)  and  a34803a );
 a34808a <=( A301  and  A300 );
 a34809a <=( (not A299)  and  a34808a );
 a34810a <=( a34809a  and  a34804a );
 a34814a <=( (not A199)  and  (not A168) );
 a34815a <=( A169  and  a34814a );
 a34819a <=( A202  and  A201 );
 a34820a <=( A200  and  a34819a );
 a34821a <=( a34820a  and  a34815a );
 a34825a <=( A298  and  A268 );
 a34826a <=( (not A267)  and  a34825a );
 a34830a <=( A302  and  A300 );
 a34831a <=( (not A299)  and  a34830a );
 a34832a <=( a34831a  and  a34826a );
 a34836a <=( (not A199)  and  (not A168) );
 a34837a <=( A169  and  a34836a );
 a34841a <=( A202  and  A201 );
 a34842a <=( A200  and  a34841a );
 a34843a <=( a34842a  and  a34837a );
 a34847a <=( (not A298)  and  A268 );
 a34848a <=( (not A267)  and  a34847a );
 a34852a <=( A301  and  A300 );
 a34853a <=( A299  and  a34852a );
 a34854a <=( a34853a  and  a34848a );
 a34858a <=( (not A199)  and  (not A168) );
 a34859a <=( A169  and  a34858a );
 a34863a <=( A202  and  A201 );
 a34864a <=( A200  and  a34863a );
 a34865a <=( a34864a  and  a34859a );
 a34869a <=( (not A298)  and  A268 );
 a34870a <=( (not A267)  and  a34869a );
 a34874a <=( A302  and  A300 );
 a34875a <=( A299  and  a34874a );
 a34876a <=( a34875a  and  a34870a );
 a34880a <=( (not A199)  and  (not A168) );
 a34881a <=( A169  and  a34880a );
 a34885a <=( A202  and  A201 );
 a34886a <=( A200  and  a34885a );
 a34887a <=( a34886a  and  a34881a );
 a34891a <=( A298  and  A269 );
 a34892a <=( (not A267)  and  a34891a );
 a34896a <=( A301  and  A300 );
 a34897a <=( (not A299)  and  a34896a );
 a34898a <=( a34897a  and  a34892a );
 a34902a <=( (not A199)  and  (not A168) );
 a34903a <=( A169  and  a34902a );
 a34907a <=( A202  and  A201 );
 a34908a <=( A200  and  a34907a );
 a34909a <=( a34908a  and  a34903a );
 a34913a <=( A298  and  A269 );
 a34914a <=( (not A267)  and  a34913a );
 a34918a <=( A302  and  A300 );
 a34919a <=( (not A299)  and  a34918a );
 a34920a <=( a34919a  and  a34914a );
 a34924a <=( (not A199)  and  (not A168) );
 a34925a <=( A169  and  a34924a );
 a34929a <=( A202  and  A201 );
 a34930a <=( A200  and  a34929a );
 a34931a <=( a34930a  and  a34925a );
 a34935a <=( (not A298)  and  A269 );
 a34936a <=( (not A267)  and  a34935a );
 a34940a <=( A301  and  A300 );
 a34941a <=( A299  and  a34940a );
 a34942a <=( a34941a  and  a34936a );
 a34946a <=( (not A199)  and  (not A168) );
 a34947a <=( A169  and  a34946a );
 a34951a <=( A202  and  A201 );
 a34952a <=( A200  and  a34951a );
 a34953a <=( a34952a  and  a34947a );
 a34957a <=( (not A298)  and  A269 );
 a34958a <=( (not A267)  and  a34957a );
 a34962a <=( A302  and  A300 );
 a34963a <=( A299  and  a34962a );
 a34964a <=( a34963a  and  a34958a );
 a34968a <=( (not A199)  and  (not A168) );
 a34969a <=( A169  and  a34968a );
 a34973a <=( A202  and  A201 );
 a34974a <=( A200  and  a34973a );
 a34975a <=( a34974a  and  a34969a );
 a34979a <=( A298  and  A266 );
 a34980a <=( A265  and  a34979a );
 a34984a <=( A301  and  A300 );
 a34985a <=( (not A299)  and  a34984a );
 a34986a <=( a34985a  and  a34980a );
 a34990a <=( (not A199)  and  (not A168) );
 a34991a <=( A169  and  a34990a );
 a34995a <=( A202  and  A201 );
 a34996a <=( A200  and  a34995a );
 a34997a <=( a34996a  and  a34991a );
 a35001a <=( A298  and  A266 );
 a35002a <=( A265  and  a35001a );
 a35006a <=( A302  and  A300 );
 a35007a <=( (not A299)  and  a35006a );
 a35008a <=( a35007a  and  a35002a );
 a35012a <=( (not A199)  and  (not A168) );
 a35013a <=( A169  and  a35012a );
 a35017a <=( A202  and  A201 );
 a35018a <=( A200  and  a35017a );
 a35019a <=( a35018a  and  a35013a );
 a35023a <=( (not A298)  and  A266 );
 a35024a <=( A265  and  a35023a );
 a35028a <=( A301  and  A300 );
 a35029a <=( A299  and  a35028a );
 a35030a <=( a35029a  and  a35024a );
 a35034a <=( (not A199)  and  (not A168) );
 a35035a <=( A169  and  a35034a );
 a35039a <=( A202  and  A201 );
 a35040a <=( A200  and  a35039a );
 a35041a <=( a35040a  and  a35035a );
 a35045a <=( (not A298)  and  A266 );
 a35046a <=( A265  and  a35045a );
 a35050a <=( A302  and  A300 );
 a35051a <=( A299  and  a35050a );
 a35052a <=( a35051a  and  a35046a );
 a35056a <=( (not A199)  and  (not A168) );
 a35057a <=( A169  and  a35056a );
 a35061a <=( A202  and  A201 );
 a35062a <=( A200  and  a35061a );
 a35063a <=( a35062a  and  a35057a );
 a35067a <=( A298  and  (not A266) );
 a35068a <=( (not A265)  and  a35067a );
 a35072a <=( A301  and  A300 );
 a35073a <=( (not A299)  and  a35072a );
 a35074a <=( a35073a  and  a35068a );
 a35078a <=( (not A199)  and  (not A168) );
 a35079a <=( A169  and  a35078a );
 a35083a <=( A202  and  A201 );
 a35084a <=( A200  and  a35083a );
 a35085a <=( a35084a  and  a35079a );
 a35089a <=( A298  and  (not A266) );
 a35090a <=( (not A265)  and  a35089a );
 a35094a <=( A302  and  A300 );
 a35095a <=( (not A299)  and  a35094a );
 a35096a <=( a35095a  and  a35090a );
 a35100a <=( (not A199)  and  (not A168) );
 a35101a <=( A169  and  a35100a );
 a35105a <=( A202  and  A201 );
 a35106a <=( A200  and  a35105a );
 a35107a <=( a35106a  and  a35101a );
 a35111a <=( (not A298)  and  (not A266) );
 a35112a <=( (not A265)  and  a35111a );
 a35116a <=( A301  and  A300 );
 a35117a <=( A299  and  a35116a );
 a35118a <=( a35117a  and  a35112a );
 a35122a <=( (not A199)  and  (not A168) );
 a35123a <=( A169  and  a35122a );
 a35127a <=( A202  and  A201 );
 a35128a <=( A200  and  a35127a );
 a35129a <=( a35128a  and  a35123a );
 a35133a <=( (not A298)  and  (not A266) );
 a35134a <=( (not A265)  and  a35133a );
 a35138a <=( A302  and  A300 );
 a35139a <=( A299  and  a35138a );
 a35140a <=( a35139a  and  a35134a );
 a35144a <=( (not A199)  and  (not A168) );
 a35145a <=( A169  and  a35144a );
 a35149a <=( A203  and  A201 );
 a35150a <=( A200  and  a35149a );
 a35151a <=( a35150a  and  a35145a );
 a35155a <=( A298  and  A268 );
 a35156a <=( (not A267)  and  a35155a );
 a35160a <=( A301  and  A300 );
 a35161a <=( (not A299)  and  a35160a );
 a35162a <=( a35161a  and  a35156a );
 a35166a <=( (not A199)  and  (not A168) );
 a35167a <=( A169  and  a35166a );
 a35171a <=( A203  and  A201 );
 a35172a <=( A200  and  a35171a );
 a35173a <=( a35172a  and  a35167a );
 a35177a <=( A298  and  A268 );
 a35178a <=( (not A267)  and  a35177a );
 a35182a <=( A302  and  A300 );
 a35183a <=( (not A299)  and  a35182a );
 a35184a <=( a35183a  and  a35178a );
 a35188a <=( (not A199)  and  (not A168) );
 a35189a <=( A169  and  a35188a );
 a35193a <=( A203  and  A201 );
 a35194a <=( A200  and  a35193a );
 a35195a <=( a35194a  and  a35189a );
 a35199a <=( (not A298)  and  A268 );
 a35200a <=( (not A267)  and  a35199a );
 a35204a <=( A301  and  A300 );
 a35205a <=( A299  and  a35204a );
 a35206a <=( a35205a  and  a35200a );
 a35210a <=( (not A199)  and  (not A168) );
 a35211a <=( A169  and  a35210a );
 a35215a <=( A203  and  A201 );
 a35216a <=( A200  and  a35215a );
 a35217a <=( a35216a  and  a35211a );
 a35221a <=( (not A298)  and  A268 );
 a35222a <=( (not A267)  and  a35221a );
 a35226a <=( A302  and  A300 );
 a35227a <=( A299  and  a35226a );
 a35228a <=( a35227a  and  a35222a );
 a35232a <=( (not A199)  and  (not A168) );
 a35233a <=( A169  and  a35232a );
 a35237a <=( A203  and  A201 );
 a35238a <=( A200  and  a35237a );
 a35239a <=( a35238a  and  a35233a );
 a35243a <=( A298  and  A269 );
 a35244a <=( (not A267)  and  a35243a );
 a35248a <=( A301  and  A300 );
 a35249a <=( (not A299)  and  a35248a );
 a35250a <=( a35249a  and  a35244a );
 a35254a <=( (not A199)  and  (not A168) );
 a35255a <=( A169  and  a35254a );
 a35259a <=( A203  and  A201 );
 a35260a <=( A200  and  a35259a );
 a35261a <=( a35260a  and  a35255a );
 a35265a <=( A298  and  A269 );
 a35266a <=( (not A267)  and  a35265a );
 a35270a <=( A302  and  A300 );
 a35271a <=( (not A299)  and  a35270a );
 a35272a <=( a35271a  and  a35266a );
 a35276a <=( (not A199)  and  (not A168) );
 a35277a <=( A169  and  a35276a );
 a35281a <=( A203  and  A201 );
 a35282a <=( A200  and  a35281a );
 a35283a <=( a35282a  and  a35277a );
 a35287a <=( (not A298)  and  A269 );
 a35288a <=( (not A267)  and  a35287a );
 a35292a <=( A301  and  A300 );
 a35293a <=( A299  and  a35292a );
 a35294a <=( a35293a  and  a35288a );
 a35298a <=( (not A199)  and  (not A168) );
 a35299a <=( A169  and  a35298a );
 a35303a <=( A203  and  A201 );
 a35304a <=( A200  and  a35303a );
 a35305a <=( a35304a  and  a35299a );
 a35309a <=( (not A298)  and  A269 );
 a35310a <=( (not A267)  and  a35309a );
 a35314a <=( A302  and  A300 );
 a35315a <=( A299  and  a35314a );
 a35316a <=( a35315a  and  a35310a );
 a35320a <=( (not A199)  and  (not A168) );
 a35321a <=( A169  and  a35320a );
 a35325a <=( A203  and  A201 );
 a35326a <=( A200  and  a35325a );
 a35327a <=( a35326a  and  a35321a );
 a35331a <=( A298  and  A266 );
 a35332a <=( A265  and  a35331a );
 a35336a <=( A301  and  A300 );
 a35337a <=( (not A299)  and  a35336a );
 a35338a <=( a35337a  and  a35332a );
 a35342a <=( (not A199)  and  (not A168) );
 a35343a <=( A169  and  a35342a );
 a35347a <=( A203  and  A201 );
 a35348a <=( A200  and  a35347a );
 a35349a <=( a35348a  and  a35343a );
 a35353a <=( A298  and  A266 );
 a35354a <=( A265  and  a35353a );
 a35358a <=( A302  and  A300 );
 a35359a <=( (not A299)  and  a35358a );
 a35360a <=( a35359a  and  a35354a );
 a35364a <=( (not A199)  and  (not A168) );
 a35365a <=( A169  and  a35364a );
 a35369a <=( A203  and  A201 );
 a35370a <=( A200  and  a35369a );
 a35371a <=( a35370a  and  a35365a );
 a35375a <=( (not A298)  and  A266 );
 a35376a <=( A265  and  a35375a );
 a35380a <=( A301  and  A300 );
 a35381a <=( A299  and  a35380a );
 a35382a <=( a35381a  and  a35376a );
 a35386a <=( (not A199)  and  (not A168) );
 a35387a <=( A169  and  a35386a );
 a35391a <=( A203  and  A201 );
 a35392a <=( A200  and  a35391a );
 a35393a <=( a35392a  and  a35387a );
 a35397a <=( (not A298)  and  A266 );
 a35398a <=( A265  and  a35397a );
 a35402a <=( A302  and  A300 );
 a35403a <=( A299  and  a35402a );
 a35404a <=( a35403a  and  a35398a );
 a35408a <=( (not A199)  and  (not A168) );
 a35409a <=( A169  and  a35408a );
 a35413a <=( A203  and  A201 );
 a35414a <=( A200  and  a35413a );
 a35415a <=( a35414a  and  a35409a );
 a35419a <=( A298  and  (not A266) );
 a35420a <=( (not A265)  and  a35419a );
 a35424a <=( A301  and  A300 );
 a35425a <=( (not A299)  and  a35424a );
 a35426a <=( a35425a  and  a35420a );
 a35430a <=( (not A199)  and  (not A168) );
 a35431a <=( A169  and  a35430a );
 a35435a <=( A203  and  A201 );
 a35436a <=( A200  and  a35435a );
 a35437a <=( a35436a  and  a35431a );
 a35441a <=( A298  and  (not A266) );
 a35442a <=( (not A265)  and  a35441a );
 a35446a <=( A302  and  A300 );
 a35447a <=( (not A299)  and  a35446a );
 a35448a <=( a35447a  and  a35442a );
 a35452a <=( (not A199)  and  (not A168) );
 a35453a <=( A169  and  a35452a );
 a35457a <=( A203  and  A201 );
 a35458a <=( A200  and  a35457a );
 a35459a <=( a35458a  and  a35453a );
 a35463a <=( (not A298)  and  (not A266) );
 a35464a <=( (not A265)  and  a35463a );
 a35468a <=( A301  and  A300 );
 a35469a <=( A299  and  a35468a );
 a35470a <=( a35469a  and  a35464a );
 a35474a <=( (not A199)  and  (not A168) );
 a35475a <=( A169  and  a35474a );
 a35479a <=( A203  and  A201 );
 a35480a <=( A200  and  a35479a );
 a35481a <=( a35480a  and  a35475a );
 a35485a <=( (not A298)  and  (not A266) );
 a35486a <=( (not A265)  and  a35485a );
 a35490a <=( A302  and  A300 );
 a35491a <=( A299  and  a35490a );
 a35492a <=( a35491a  and  a35486a );
 a35496a <=( A199  and  (not A168) );
 a35497a <=( A169  and  a35496a );
 a35501a <=( A202  and  A201 );
 a35502a <=( (not A200)  and  a35501a );
 a35503a <=( a35502a  and  a35497a );
 a35507a <=( A298  and  A268 );
 a35508a <=( (not A267)  and  a35507a );
 a35512a <=( A301  and  A300 );
 a35513a <=( (not A299)  and  a35512a );
 a35514a <=( a35513a  and  a35508a );
 a35518a <=( A199  and  (not A168) );
 a35519a <=( A169  and  a35518a );
 a35523a <=( A202  and  A201 );
 a35524a <=( (not A200)  and  a35523a );
 a35525a <=( a35524a  and  a35519a );
 a35529a <=( A298  and  A268 );
 a35530a <=( (not A267)  and  a35529a );
 a35534a <=( A302  and  A300 );
 a35535a <=( (not A299)  and  a35534a );
 a35536a <=( a35535a  and  a35530a );
 a35540a <=( A199  and  (not A168) );
 a35541a <=( A169  and  a35540a );
 a35545a <=( A202  and  A201 );
 a35546a <=( (not A200)  and  a35545a );
 a35547a <=( a35546a  and  a35541a );
 a35551a <=( (not A298)  and  A268 );
 a35552a <=( (not A267)  and  a35551a );
 a35556a <=( A301  and  A300 );
 a35557a <=( A299  and  a35556a );
 a35558a <=( a35557a  and  a35552a );
 a35562a <=( A199  and  (not A168) );
 a35563a <=( A169  and  a35562a );
 a35567a <=( A202  and  A201 );
 a35568a <=( (not A200)  and  a35567a );
 a35569a <=( a35568a  and  a35563a );
 a35573a <=( (not A298)  and  A268 );
 a35574a <=( (not A267)  and  a35573a );
 a35578a <=( A302  and  A300 );
 a35579a <=( A299  and  a35578a );
 a35580a <=( a35579a  and  a35574a );
 a35584a <=( A199  and  (not A168) );
 a35585a <=( A169  and  a35584a );
 a35589a <=( A202  and  A201 );
 a35590a <=( (not A200)  and  a35589a );
 a35591a <=( a35590a  and  a35585a );
 a35595a <=( A298  and  A269 );
 a35596a <=( (not A267)  and  a35595a );
 a35600a <=( A301  and  A300 );
 a35601a <=( (not A299)  and  a35600a );
 a35602a <=( a35601a  and  a35596a );
 a35606a <=( A199  and  (not A168) );
 a35607a <=( A169  and  a35606a );
 a35611a <=( A202  and  A201 );
 a35612a <=( (not A200)  and  a35611a );
 a35613a <=( a35612a  and  a35607a );
 a35617a <=( A298  and  A269 );
 a35618a <=( (not A267)  and  a35617a );
 a35622a <=( A302  and  A300 );
 a35623a <=( (not A299)  and  a35622a );
 a35624a <=( a35623a  and  a35618a );
 a35628a <=( A199  and  (not A168) );
 a35629a <=( A169  and  a35628a );
 a35633a <=( A202  and  A201 );
 a35634a <=( (not A200)  and  a35633a );
 a35635a <=( a35634a  and  a35629a );
 a35639a <=( (not A298)  and  A269 );
 a35640a <=( (not A267)  and  a35639a );
 a35644a <=( A301  and  A300 );
 a35645a <=( A299  and  a35644a );
 a35646a <=( a35645a  and  a35640a );
 a35650a <=( A199  and  (not A168) );
 a35651a <=( A169  and  a35650a );
 a35655a <=( A202  and  A201 );
 a35656a <=( (not A200)  and  a35655a );
 a35657a <=( a35656a  and  a35651a );
 a35661a <=( (not A298)  and  A269 );
 a35662a <=( (not A267)  and  a35661a );
 a35666a <=( A302  and  A300 );
 a35667a <=( A299  and  a35666a );
 a35668a <=( a35667a  and  a35662a );
 a35672a <=( A199  and  (not A168) );
 a35673a <=( A169  and  a35672a );
 a35677a <=( A202  and  A201 );
 a35678a <=( (not A200)  and  a35677a );
 a35679a <=( a35678a  and  a35673a );
 a35683a <=( A298  and  A266 );
 a35684a <=( A265  and  a35683a );
 a35688a <=( A301  and  A300 );
 a35689a <=( (not A299)  and  a35688a );
 a35690a <=( a35689a  and  a35684a );
 a35694a <=( A199  and  (not A168) );
 a35695a <=( A169  and  a35694a );
 a35699a <=( A202  and  A201 );
 a35700a <=( (not A200)  and  a35699a );
 a35701a <=( a35700a  and  a35695a );
 a35705a <=( A298  and  A266 );
 a35706a <=( A265  and  a35705a );
 a35710a <=( A302  and  A300 );
 a35711a <=( (not A299)  and  a35710a );
 a35712a <=( a35711a  and  a35706a );
 a35716a <=( A199  and  (not A168) );
 a35717a <=( A169  and  a35716a );
 a35721a <=( A202  and  A201 );
 a35722a <=( (not A200)  and  a35721a );
 a35723a <=( a35722a  and  a35717a );
 a35727a <=( (not A298)  and  A266 );
 a35728a <=( A265  and  a35727a );
 a35732a <=( A301  and  A300 );
 a35733a <=( A299  and  a35732a );
 a35734a <=( a35733a  and  a35728a );
 a35738a <=( A199  and  (not A168) );
 a35739a <=( A169  and  a35738a );
 a35743a <=( A202  and  A201 );
 a35744a <=( (not A200)  and  a35743a );
 a35745a <=( a35744a  and  a35739a );
 a35749a <=( (not A298)  and  A266 );
 a35750a <=( A265  and  a35749a );
 a35754a <=( A302  and  A300 );
 a35755a <=( A299  and  a35754a );
 a35756a <=( a35755a  and  a35750a );
 a35760a <=( A199  and  (not A168) );
 a35761a <=( A169  and  a35760a );
 a35765a <=( A202  and  A201 );
 a35766a <=( (not A200)  and  a35765a );
 a35767a <=( a35766a  and  a35761a );
 a35771a <=( A298  and  (not A266) );
 a35772a <=( (not A265)  and  a35771a );
 a35776a <=( A301  and  A300 );
 a35777a <=( (not A299)  and  a35776a );
 a35778a <=( a35777a  and  a35772a );
 a35782a <=( A199  and  (not A168) );
 a35783a <=( A169  and  a35782a );
 a35787a <=( A202  and  A201 );
 a35788a <=( (not A200)  and  a35787a );
 a35789a <=( a35788a  and  a35783a );
 a35793a <=( A298  and  (not A266) );
 a35794a <=( (not A265)  and  a35793a );
 a35798a <=( A302  and  A300 );
 a35799a <=( (not A299)  and  a35798a );
 a35800a <=( a35799a  and  a35794a );
 a35804a <=( A199  and  (not A168) );
 a35805a <=( A169  and  a35804a );
 a35809a <=( A202  and  A201 );
 a35810a <=( (not A200)  and  a35809a );
 a35811a <=( a35810a  and  a35805a );
 a35815a <=( (not A298)  and  (not A266) );
 a35816a <=( (not A265)  and  a35815a );
 a35820a <=( A301  and  A300 );
 a35821a <=( A299  and  a35820a );
 a35822a <=( a35821a  and  a35816a );
 a35826a <=( A199  and  (not A168) );
 a35827a <=( A169  and  a35826a );
 a35831a <=( A202  and  A201 );
 a35832a <=( (not A200)  and  a35831a );
 a35833a <=( a35832a  and  a35827a );
 a35837a <=( (not A298)  and  (not A266) );
 a35838a <=( (not A265)  and  a35837a );
 a35842a <=( A302  and  A300 );
 a35843a <=( A299  and  a35842a );
 a35844a <=( a35843a  and  a35838a );
 a35848a <=( A199  and  (not A168) );
 a35849a <=( A169  and  a35848a );
 a35853a <=( A203  and  A201 );
 a35854a <=( (not A200)  and  a35853a );
 a35855a <=( a35854a  and  a35849a );
 a35859a <=( A298  and  A268 );
 a35860a <=( (not A267)  and  a35859a );
 a35864a <=( A301  and  A300 );
 a35865a <=( (not A299)  and  a35864a );
 a35866a <=( a35865a  and  a35860a );
 a35870a <=( A199  and  (not A168) );
 a35871a <=( A169  and  a35870a );
 a35875a <=( A203  and  A201 );
 a35876a <=( (not A200)  and  a35875a );
 a35877a <=( a35876a  and  a35871a );
 a35881a <=( A298  and  A268 );
 a35882a <=( (not A267)  and  a35881a );
 a35886a <=( A302  and  A300 );
 a35887a <=( (not A299)  and  a35886a );
 a35888a <=( a35887a  and  a35882a );
 a35892a <=( A199  and  (not A168) );
 a35893a <=( A169  and  a35892a );
 a35897a <=( A203  and  A201 );
 a35898a <=( (not A200)  and  a35897a );
 a35899a <=( a35898a  and  a35893a );
 a35903a <=( (not A298)  and  A268 );
 a35904a <=( (not A267)  and  a35903a );
 a35908a <=( A301  and  A300 );
 a35909a <=( A299  and  a35908a );
 a35910a <=( a35909a  and  a35904a );
 a35914a <=( A199  and  (not A168) );
 a35915a <=( A169  and  a35914a );
 a35919a <=( A203  and  A201 );
 a35920a <=( (not A200)  and  a35919a );
 a35921a <=( a35920a  and  a35915a );
 a35925a <=( (not A298)  and  A268 );
 a35926a <=( (not A267)  and  a35925a );
 a35930a <=( A302  and  A300 );
 a35931a <=( A299  and  a35930a );
 a35932a <=( a35931a  and  a35926a );
 a35936a <=( A199  and  (not A168) );
 a35937a <=( A169  and  a35936a );
 a35941a <=( A203  and  A201 );
 a35942a <=( (not A200)  and  a35941a );
 a35943a <=( a35942a  and  a35937a );
 a35947a <=( A298  and  A269 );
 a35948a <=( (not A267)  and  a35947a );
 a35952a <=( A301  and  A300 );
 a35953a <=( (not A299)  and  a35952a );
 a35954a <=( a35953a  and  a35948a );
 a35958a <=( A199  and  (not A168) );
 a35959a <=( A169  and  a35958a );
 a35963a <=( A203  and  A201 );
 a35964a <=( (not A200)  and  a35963a );
 a35965a <=( a35964a  and  a35959a );
 a35969a <=( A298  and  A269 );
 a35970a <=( (not A267)  and  a35969a );
 a35974a <=( A302  and  A300 );
 a35975a <=( (not A299)  and  a35974a );
 a35976a <=( a35975a  and  a35970a );
 a35980a <=( A199  and  (not A168) );
 a35981a <=( A169  and  a35980a );
 a35985a <=( A203  and  A201 );
 a35986a <=( (not A200)  and  a35985a );
 a35987a <=( a35986a  and  a35981a );
 a35991a <=( (not A298)  and  A269 );
 a35992a <=( (not A267)  and  a35991a );
 a35996a <=( A301  and  A300 );
 a35997a <=( A299  and  a35996a );
 a35998a <=( a35997a  and  a35992a );
 a36002a <=( A199  and  (not A168) );
 a36003a <=( A169  and  a36002a );
 a36007a <=( A203  and  A201 );
 a36008a <=( (not A200)  and  a36007a );
 a36009a <=( a36008a  and  a36003a );
 a36013a <=( (not A298)  and  A269 );
 a36014a <=( (not A267)  and  a36013a );
 a36018a <=( A302  and  A300 );
 a36019a <=( A299  and  a36018a );
 a36020a <=( a36019a  and  a36014a );
 a36024a <=( A199  and  (not A168) );
 a36025a <=( A169  and  a36024a );
 a36029a <=( A203  and  A201 );
 a36030a <=( (not A200)  and  a36029a );
 a36031a <=( a36030a  and  a36025a );
 a36035a <=( A298  and  A266 );
 a36036a <=( A265  and  a36035a );
 a36040a <=( A301  and  A300 );
 a36041a <=( (not A299)  and  a36040a );
 a36042a <=( a36041a  and  a36036a );
 a36046a <=( A199  and  (not A168) );
 a36047a <=( A169  and  a36046a );
 a36051a <=( A203  and  A201 );
 a36052a <=( (not A200)  and  a36051a );
 a36053a <=( a36052a  and  a36047a );
 a36057a <=( A298  and  A266 );
 a36058a <=( A265  and  a36057a );
 a36062a <=( A302  and  A300 );
 a36063a <=( (not A299)  and  a36062a );
 a36064a <=( a36063a  and  a36058a );
 a36068a <=( A199  and  (not A168) );
 a36069a <=( A169  and  a36068a );
 a36073a <=( A203  and  A201 );
 a36074a <=( (not A200)  and  a36073a );
 a36075a <=( a36074a  and  a36069a );
 a36079a <=( (not A298)  and  A266 );
 a36080a <=( A265  and  a36079a );
 a36084a <=( A301  and  A300 );
 a36085a <=( A299  and  a36084a );
 a36086a <=( a36085a  and  a36080a );
 a36090a <=( A199  and  (not A168) );
 a36091a <=( A169  and  a36090a );
 a36095a <=( A203  and  A201 );
 a36096a <=( (not A200)  and  a36095a );
 a36097a <=( a36096a  and  a36091a );
 a36101a <=( (not A298)  and  A266 );
 a36102a <=( A265  and  a36101a );
 a36106a <=( A302  and  A300 );
 a36107a <=( A299  and  a36106a );
 a36108a <=( a36107a  and  a36102a );
 a36112a <=( A199  and  (not A168) );
 a36113a <=( A169  and  a36112a );
 a36117a <=( A203  and  A201 );
 a36118a <=( (not A200)  and  a36117a );
 a36119a <=( a36118a  and  a36113a );
 a36123a <=( A298  and  (not A266) );
 a36124a <=( (not A265)  and  a36123a );
 a36128a <=( A301  and  A300 );
 a36129a <=( (not A299)  and  a36128a );
 a36130a <=( a36129a  and  a36124a );
 a36134a <=( A199  and  (not A168) );
 a36135a <=( A169  and  a36134a );
 a36139a <=( A203  and  A201 );
 a36140a <=( (not A200)  and  a36139a );
 a36141a <=( a36140a  and  a36135a );
 a36145a <=( A298  and  (not A266) );
 a36146a <=( (not A265)  and  a36145a );
 a36150a <=( A302  and  A300 );
 a36151a <=( (not A299)  and  a36150a );
 a36152a <=( a36151a  and  a36146a );
 a36156a <=( A199  and  (not A168) );
 a36157a <=( A169  and  a36156a );
 a36161a <=( A203  and  A201 );
 a36162a <=( (not A200)  and  a36161a );
 a36163a <=( a36162a  and  a36157a );
 a36167a <=( (not A298)  and  (not A266) );
 a36168a <=( (not A265)  and  a36167a );
 a36172a <=( A301  and  A300 );
 a36173a <=( A299  and  a36172a );
 a36174a <=( a36173a  and  a36168a );
 a36178a <=( A199  and  (not A168) );
 a36179a <=( A169  and  a36178a );
 a36183a <=( A203  and  A201 );
 a36184a <=( (not A200)  and  a36183a );
 a36185a <=( a36184a  and  a36179a );
 a36189a <=( (not A298)  and  (not A266) );
 a36190a <=( (not A265)  and  a36189a );
 a36194a <=( A302  and  A300 );
 a36195a <=( A299  and  a36194a );
 a36196a <=( a36195a  and  a36190a );
 a36200a <=( (not A199)  and  (not A168) );
 a36201a <=( A169  and  a36200a );
 a36205a <=( A266  and  (not A265) );
 a36206a <=( (not A200)  and  a36205a );
 a36207a <=( a36206a  and  a36201a );
 a36211a <=( (not A269)  and  (not A268) );
 a36212a <=( (not A267)  and  a36211a );
 a36216a <=( (not A302)  and  (not A301) );
 a36217a <=( A300  and  a36216a );
 a36218a <=( a36217a  and  a36212a );
 a36222a <=( (not A199)  and  (not A168) );
 a36223a <=( A169  and  a36222a );
 a36227a <=( (not A266)  and  A265 );
 a36228a <=( (not A200)  and  a36227a );
 a36229a <=( a36228a  and  a36223a );
 a36233a <=( (not A269)  and  (not A268) );
 a36234a <=( (not A267)  and  a36233a );
 a36238a <=( (not A302)  and  (not A301) );
 a36239a <=( A300  and  a36238a );
 a36240a <=( a36239a  and  a36234a );
 a36244a <=( A168  and  (not A169) );
 a36245a <=( A170  and  a36244a );
 a36249a <=( (not A203)  and  (not A202) );
 a36250a <=( A201  and  a36249a );
 a36251a <=( a36250a  and  a36245a );
 a36255a <=( A267  and  A266 );
 a36256a <=( (not A265)  and  a36255a );
 a36260a <=( A301  and  (not A300) );
 a36261a <=( A268  and  a36260a );
 a36262a <=( a36261a  and  a36256a );
 a36266a <=( A168  and  (not A169) );
 a36267a <=( A170  and  a36266a );
 a36271a <=( (not A203)  and  (not A202) );
 a36272a <=( A201  and  a36271a );
 a36273a <=( a36272a  and  a36267a );
 a36277a <=( A267  and  A266 );
 a36278a <=( (not A265)  and  a36277a );
 a36282a <=( A302  and  (not A300) );
 a36283a <=( A268  and  a36282a );
 a36284a <=( a36283a  and  a36278a );
 a36288a <=( A168  and  (not A169) );
 a36289a <=( A170  and  a36288a );
 a36293a <=( (not A203)  and  (not A202) );
 a36294a <=( A201  and  a36293a );
 a36295a <=( a36294a  and  a36289a );
 a36299a <=( A267  and  A266 );
 a36300a <=( (not A265)  and  a36299a );
 a36304a <=( A299  and  A298 );
 a36305a <=( A268  and  a36304a );
 a36306a <=( a36305a  and  a36300a );
 a36310a <=( A168  and  (not A169) );
 a36311a <=( A170  and  a36310a );
 a36315a <=( (not A203)  and  (not A202) );
 a36316a <=( A201  and  a36315a );
 a36317a <=( a36316a  and  a36311a );
 a36321a <=( A267  and  A266 );
 a36322a <=( (not A265)  and  a36321a );
 a36326a <=( (not A299)  and  (not A298) );
 a36327a <=( A268  and  a36326a );
 a36328a <=( a36327a  and  a36322a );
 a36332a <=( A168  and  (not A169) );
 a36333a <=( A170  and  a36332a );
 a36337a <=( (not A203)  and  (not A202) );
 a36338a <=( A201  and  a36337a );
 a36339a <=( a36338a  and  a36333a );
 a36343a <=( A267  and  A266 );
 a36344a <=( (not A265)  and  a36343a );
 a36348a <=( A301  and  (not A300) );
 a36349a <=( A269  and  a36348a );
 a36350a <=( a36349a  and  a36344a );
 a36354a <=( A168  and  (not A169) );
 a36355a <=( A170  and  a36354a );
 a36359a <=( (not A203)  and  (not A202) );
 a36360a <=( A201  and  a36359a );
 a36361a <=( a36360a  and  a36355a );
 a36365a <=( A267  and  A266 );
 a36366a <=( (not A265)  and  a36365a );
 a36370a <=( A302  and  (not A300) );
 a36371a <=( A269  and  a36370a );
 a36372a <=( a36371a  and  a36366a );
 a36376a <=( A168  and  (not A169) );
 a36377a <=( A170  and  a36376a );
 a36381a <=( (not A203)  and  (not A202) );
 a36382a <=( A201  and  a36381a );
 a36383a <=( a36382a  and  a36377a );
 a36387a <=( A267  and  A266 );
 a36388a <=( (not A265)  and  a36387a );
 a36392a <=( A299  and  A298 );
 a36393a <=( A269  and  a36392a );
 a36394a <=( a36393a  and  a36388a );
 a36398a <=( A168  and  (not A169) );
 a36399a <=( A170  and  a36398a );
 a36403a <=( (not A203)  and  (not A202) );
 a36404a <=( A201  and  a36403a );
 a36405a <=( a36404a  and  a36399a );
 a36409a <=( A267  and  A266 );
 a36410a <=( (not A265)  and  a36409a );
 a36414a <=( (not A299)  and  (not A298) );
 a36415a <=( A269  and  a36414a );
 a36416a <=( a36415a  and  a36410a );
 a36420a <=( A168  and  (not A169) );
 a36421a <=( A170  and  a36420a );
 a36425a <=( (not A203)  and  (not A202) );
 a36426a <=( A201  and  a36425a );
 a36427a <=( a36426a  and  a36421a );
 a36431a <=( A267  and  (not A266) );
 a36432a <=( A265  and  a36431a );
 a36436a <=( A301  and  (not A300) );
 a36437a <=( A268  and  a36436a );
 a36438a <=( a36437a  and  a36432a );
 a36442a <=( A168  and  (not A169) );
 a36443a <=( A170  and  a36442a );
 a36447a <=( (not A203)  and  (not A202) );
 a36448a <=( A201  and  a36447a );
 a36449a <=( a36448a  and  a36443a );
 a36453a <=( A267  and  (not A266) );
 a36454a <=( A265  and  a36453a );
 a36458a <=( A302  and  (not A300) );
 a36459a <=( A268  and  a36458a );
 a36460a <=( a36459a  and  a36454a );
 a36464a <=( A168  and  (not A169) );
 a36465a <=( A170  and  a36464a );
 a36469a <=( (not A203)  and  (not A202) );
 a36470a <=( A201  and  a36469a );
 a36471a <=( a36470a  and  a36465a );
 a36475a <=( A267  and  (not A266) );
 a36476a <=( A265  and  a36475a );
 a36480a <=( A299  and  A298 );
 a36481a <=( A268  and  a36480a );
 a36482a <=( a36481a  and  a36476a );
 a36486a <=( A168  and  (not A169) );
 a36487a <=( A170  and  a36486a );
 a36491a <=( (not A203)  and  (not A202) );
 a36492a <=( A201  and  a36491a );
 a36493a <=( a36492a  and  a36487a );
 a36497a <=( A267  and  (not A266) );
 a36498a <=( A265  and  a36497a );
 a36502a <=( (not A299)  and  (not A298) );
 a36503a <=( A268  and  a36502a );
 a36504a <=( a36503a  and  a36498a );
 a36508a <=( A168  and  (not A169) );
 a36509a <=( A170  and  a36508a );
 a36513a <=( (not A203)  and  (not A202) );
 a36514a <=( A201  and  a36513a );
 a36515a <=( a36514a  and  a36509a );
 a36519a <=( A267  and  (not A266) );
 a36520a <=( A265  and  a36519a );
 a36524a <=( A301  and  (not A300) );
 a36525a <=( A269  and  a36524a );
 a36526a <=( a36525a  and  a36520a );
 a36530a <=( A168  and  (not A169) );
 a36531a <=( A170  and  a36530a );
 a36535a <=( (not A203)  and  (not A202) );
 a36536a <=( A201  and  a36535a );
 a36537a <=( a36536a  and  a36531a );
 a36541a <=( A267  and  (not A266) );
 a36542a <=( A265  and  a36541a );
 a36546a <=( A302  and  (not A300) );
 a36547a <=( A269  and  a36546a );
 a36548a <=( a36547a  and  a36542a );
 a36552a <=( A168  and  (not A169) );
 a36553a <=( A170  and  a36552a );
 a36557a <=( (not A203)  and  (not A202) );
 a36558a <=( A201  and  a36557a );
 a36559a <=( a36558a  and  a36553a );
 a36563a <=( A267  and  (not A266) );
 a36564a <=( A265  and  a36563a );
 a36568a <=( A299  and  A298 );
 a36569a <=( A269  and  a36568a );
 a36570a <=( a36569a  and  a36564a );
 a36574a <=( A168  and  (not A169) );
 a36575a <=( A170  and  a36574a );
 a36579a <=( (not A203)  and  (not A202) );
 a36580a <=( A201  and  a36579a );
 a36581a <=( a36580a  and  a36575a );
 a36585a <=( A267  and  (not A266) );
 a36586a <=( A265  and  a36585a );
 a36590a <=( (not A299)  and  (not A298) );
 a36591a <=( A269  and  a36590a );
 a36592a <=( a36591a  and  a36586a );
 a36596a <=( A168  and  (not A169) );
 a36597a <=( A170  and  a36596a );
 a36601a <=( (not A265)  and  A202 );
 a36602a <=( (not A201)  and  a36601a );
 a36603a <=( a36602a  and  a36597a );
 a36607a <=( A268  and  A267 );
 a36608a <=( A266  and  a36607a );
 a36612a <=( (not A302)  and  (not A301) );
 a36613a <=( A300  and  a36612a );
 a36614a <=( a36613a  and  a36608a );
 a36618a <=( A168  and  (not A169) );
 a36619a <=( A170  and  a36618a );
 a36623a <=( (not A265)  and  A202 );
 a36624a <=( (not A201)  and  a36623a );
 a36625a <=( a36624a  and  a36619a );
 a36629a <=( A269  and  A267 );
 a36630a <=( A266  and  a36629a );
 a36634a <=( (not A302)  and  (not A301) );
 a36635a <=( A300  and  a36634a );
 a36636a <=( a36635a  and  a36630a );
 a36640a <=( A168  and  (not A169) );
 a36641a <=( A170  and  a36640a );
 a36645a <=( (not A265)  and  A202 );
 a36646a <=( (not A201)  and  a36645a );
 a36647a <=( a36646a  and  a36641a );
 a36651a <=( (not A268)  and  (not A267) );
 a36652a <=( A266  and  a36651a );
 a36656a <=( A301  and  (not A300) );
 a36657a <=( (not A269)  and  a36656a );
 a36658a <=( a36657a  and  a36652a );
 a36662a <=( A168  and  (not A169) );
 a36663a <=( A170  and  a36662a );
 a36667a <=( (not A265)  and  A202 );
 a36668a <=( (not A201)  and  a36667a );
 a36669a <=( a36668a  and  a36663a );
 a36673a <=( (not A268)  and  (not A267) );
 a36674a <=( A266  and  a36673a );
 a36678a <=( A302  and  (not A300) );
 a36679a <=( (not A269)  and  a36678a );
 a36680a <=( a36679a  and  a36674a );
 a36684a <=( A168  and  (not A169) );
 a36685a <=( A170  and  a36684a );
 a36689a <=( (not A265)  and  A202 );
 a36690a <=( (not A201)  and  a36689a );
 a36691a <=( a36690a  and  a36685a );
 a36695a <=( (not A268)  and  (not A267) );
 a36696a <=( A266  and  a36695a );
 a36700a <=( A299  and  A298 );
 a36701a <=( (not A269)  and  a36700a );
 a36702a <=( a36701a  and  a36696a );
 a36706a <=( A168  and  (not A169) );
 a36707a <=( A170  and  a36706a );
 a36711a <=( (not A265)  and  A202 );
 a36712a <=( (not A201)  and  a36711a );
 a36713a <=( a36712a  and  a36707a );
 a36717a <=( (not A268)  and  (not A267) );
 a36718a <=( A266  and  a36717a );
 a36722a <=( (not A299)  and  (not A298) );
 a36723a <=( (not A269)  and  a36722a );
 a36724a <=( a36723a  and  a36718a );
 a36728a <=( A168  and  (not A169) );
 a36729a <=( A170  and  a36728a );
 a36733a <=( A265  and  A202 );
 a36734a <=( (not A201)  and  a36733a );
 a36735a <=( a36734a  and  a36729a );
 a36739a <=( A268  and  A267 );
 a36740a <=( (not A266)  and  a36739a );
 a36744a <=( (not A302)  and  (not A301) );
 a36745a <=( A300  and  a36744a );
 a36746a <=( a36745a  and  a36740a );
 a36750a <=( A168  and  (not A169) );
 a36751a <=( A170  and  a36750a );
 a36755a <=( A265  and  A202 );
 a36756a <=( (not A201)  and  a36755a );
 a36757a <=( a36756a  and  a36751a );
 a36761a <=( A269  and  A267 );
 a36762a <=( (not A266)  and  a36761a );
 a36766a <=( (not A302)  and  (not A301) );
 a36767a <=( A300  and  a36766a );
 a36768a <=( a36767a  and  a36762a );
 a36772a <=( A168  and  (not A169) );
 a36773a <=( A170  and  a36772a );
 a36777a <=( A265  and  A202 );
 a36778a <=( (not A201)  and  a36777a );
 a36779a <=( a36778a  and  a36773a );
 a36783a <=( (not A268)  and  (not A267) );
 a36784a <=( (not A266)  and  a36783a );
 a36788a <=( A301  and  (not A300) );
 a36789a <=( (not A269)  and  a36788a );
 a36790a <=( a36789a  and  a36784a );
 a36794a <=( A168  and  (not A169) );
 a36795a <=( A170  and  a36794a );
 a36799a <=( A265  and  A202 );
 a36800a <=( (not A201)  and  a36799a );
 a36801a <=( a36800a  and  a36795a );
 a36805a <=( (not A268)  and  (not A267) );
 a36806a <=( (not A266)  and  a36805a );
 a36810a <=( A302  and  (not A300) );
 a36811a <=( (not A269)  and  a36810a );
 a36812a <=( a36811a  and  a36806a );
 a36816a <=( A168  and  (not A169) );
 a36817a <=( A170  and  a36816a );
 a36821a <=( A265  and  A202 );
 a36822a <=( (not A201)  and  a36821a );
 a36823a <=( a36822a  and  a36817a );
 a36827a <=( (not A268)  and  (not A267) );
 a36828a <=( (not A266)  and  a36827a );
 a36832a <=( A299  and  A298 );
 a36833a <=( (not A269)  and  a36832a );
 a36834a <=( a36833a  and  a36828a );
 a36838a <=( A168  and  (not A169) );
 a36839a <=( A170  and  a36838a );
 a36843a <=( A265  and  A202 );
 a36844a <=( (not A201)  and  a36843a );
 a36845a <=( a36844a  and  a36839a );
 a36849a <=( (not A268)  and  (not A267) );
 a36850a <=( (not A266)  and  a36849a );
 a36854a <=( (not A299)  and  (not A298) );
 a36855a <=( (not A269)  and  a36854a );
 a36856a <=( a36855a  and  a36850a );
 a36860a <=( A168  and  (not A169) );
 a36861a <=( A170  and  a36860a );
 a36865a <=( (not A265)  and  A203 );
 a36866a <=( (not A201)  and  a36865a );
 a36867a <=( a36866a  and  a36861a );
 a36871a <=( A268  and  A267 );
 a36872a <=( A266  and  a36871a );
 a36876a <=( (not A302)  and  (not A301) );
 a36877a <=( A300  and  a36876a );
 a36878a <=( a36877a  and  a36872a );
 a36882a <=( A168  and  (not A169) );
 a36883a <=( A170  and  a36882a );
 a36887a <=( (not A265)  and  A203 );
 a36888a <=( (not A201)  and  a36887a );
 a36889a <=( a36888a  and  a36883a );
 a36893a <=( A269  and  A267 );
 a36894a <=( A266  and  a36893a );
 a36898a <=( (not A302)  and  (not A301) );
 a36899a <=( A300  and  a36898a );
 a36900a <=( a36899a  and  a36894a );
 a36904a <=( A168  and  (not A169) );
 a36905a <=( A170  and  a36904a );
 a36909a <=( (not A265)  and  A203 );
 a36910a <=( (not A201)  and  a36909a );
 a36911a <=( a36910a  and  a36905a );
 a36915a <=( (not A268)  and  (not A267) );
 a36916a <=( A266  and  a36915a );
 a36920a <=( A301  and  (not A300) );
 a36921a <=( (not A269)  and  a36920a );
 a36922a <=( a36921a  and  a36916a );
 a36926a <=( A168  and  (not A169) );
 a36927a <=( A170  and  a36926a );
 a36931a <=( (not A265)  and  A203 );
 a36932a <=( (not A201)  and  a36931a );
 a36933a <=( a36932a  and  a36927a );
 a36937a <=( (not A268)  and  (not A267) );
 a36938a <=( A266  and  a36937a );
 a36942a <=( A302  and  (not A300) );
 a36943a <=( (not A269)  and  a36942a );
 a36944a <=( a36943a  and  a36938a );
 a36948a <=( A168  and  (not A169) );
 a36949a <=( A170  and  a36948a );
 a36953a <=( (not A265)  and  A203 );
 a36954a <=( (not A201)  and  a36953a );
 a36955a <=( a36954a  and  a36949a );
 a36959a <=( (not A268)  and  (not A267) );
 a36960a <=( A266  and  a36959a );
 a36964a <=( A299  and  A298 );
 a36965a <=( (not A269)  and  a36964a );
 a36966a <=( a36965a  and  a36960a );
 a36970a <=( A168  and  (not A169) );
 a36971a <=( A170  and  a36970a );
 a36975a <=( (not A265)  and  A203 );
 a36976a <=( (not A201)  and  a36975a );
 a36977a <=( a36976a  and  a36971a );
 a36981a <=( (not A268)  and  (not A267) );
 a36982a <=( A266  and  a36981a );
 a36986a <=( (not A299)  and  (not A298) );
 a36987a <=( (not A269)  and  a36986a );
 a36988a <=( a36987a  and  a36982a );
 a36992a <=( A168  and  (not A169) );
 a36993a <=( A170  and  a36992a );
 a36997a <=( A265  and  A203 );
 a36998a <=( (not A201)  and  a36997a );
 a36999a <=( a36998a  and  a36993a );
 a37003a <=( A268  and  A267 );
 a37004a <=( (not A266)  and  a37003a );
 a37008a <=( (not A302)  and  (not A301) );
 a37009a <=( A300  and  a37008a );
 a37010a <=( a37009a  and  a37004a );
 a37014a <=( A168  and  (not A169) );
 a37015a <=( A170  and  a37014a );
 a37019a <=( A265  and  A203 );
 a37020a <=( (not A201)  and  a37019a );
 a37021a <=( a37020a  and  a37015a );
 a37025a <=( A269  and  A267 );
 a37026a <=( (not A266)  and  a37025a );
 a37030a <=( (not A302)  and  (not A301) );
 a37031a <=( A300  and  a37030a );
 a37032a <=( a37031a  and  a37026a );
 a37036a <=( A168  and  (not A169) );
 a37037a <=( A170  and  a37036a );
 a37041a <=( A265  and  A203 );
 a37042a <=( (not A201)  and  a37041a );
 a37043a <=( a37042a  and  a37037a );
 a37047a <=( (not A268)  and  (not A267) );
 a37048a <=( (not A266)  and  a37047a );
 a37052a <=( A301  and  (not A300) );
 a37053a <=( (not A269)  and  a37052a );
 a37054a <=( a37053a  and  a37048a );
 a37058a <=( A168  and  (not A169) );
 a37059a <=( A170  and  a37058a );
 a37063a <=( A265  and  A203 );
 a37064a <=( (not A201)  and  a37063a );
 a37065a <=( a37064a  and  a37059a );
 a37069a <=( (not A268)  and  (not A267) );
 a37070a <=( (not A266)  and  a37069a );
 a37074a <=( A302  and  (not A300) );
 a37075a <=( (not A269)  and  a37074a );
 a37076a <=( a37075a  and  a37070a );
 a37080a <=( A168  and  (not A169) );
 a37081a <=( A170  and  a37080a );
 a37085a <=( A265  and  A203 );
 a37086a <=( (not A201)  and  a37085a );
 a37087a <=( a37086a  and  a37081a );
 a37091a <=( (not A268)  and  (not A267) );
 a37092a <=( (not A266)  and  a37091a );
 a37096a <=( A299  and  A298 );
 a37097a <=( (not A269)  and  a37096a );
 a37098a <=( a37097a  and  a37092a );
 a37102a <=( A168  and  (not A169) );
 a37103a <=( A170  and  a37102a );
 a37107a <=( A265  and  A203 );
 a37108a <=( (not A201)  and  a37107a );
 a37109a <=( a37108a  and  a37103a );
 a37113a <=( (not A268)  and  (not A267) );
 a37114a <=( (not A266)  and  a37113a );
 a37118a <=( (not A299)  and  (not A298) );
 a37119a <=( (not A269)  and  a37118a );
 a37120a <=( a37119a  and  a37114a );
 a37124a <=( A168  and  (not A169) );
 a37125a <=( A170  and  a37124a );
 a37129a <=( (not A265)  and  A200 );
 a37130a <=( A199  and  a37129a );
 a37131a <=( a37130a  and  a37125a );
 a37135a <=( A268  and  A267 );
 a37136a <=( A266  and  a37135a );
 a37140a <=( (not A302)  and  (not A301) );
 a37141a <=( A300  and  a37140a );
 a37142a <=( a37141a  and  a37136a );
 a37146a <=( A168  and  (not A169) );
 a37147a <=( A170  and  a37146a );
 a37151a <=( (not A265)  and  A200 );
 a37152a <=( A199  and  a37151a );
 a37153a <=( a37152a  and  a37147a );
 a37157a <=( A269  and  A267 );
 a37158a <=( A266  and  a37157a );
 a37162a <=( (not A302)  and  (not A301) );
 a37163a <=( A300  and  a37162a );
 a37164a <=( a37163a  and  a37158a );
 a37168a <=( A168  and  (not A169) );
 a37169a <=( A170  and  a37168a );
 a37173a <=( (not A265)  and  A200 );
 a37174a <=( A199  and  a37173a );
 a37175a <=( a37174a  and  a37169a );
 a37179a <=( (not A268)  and  (not A267) );
 a37180a <=( A266  and  a37179a );
 a37184a <=( A301  and  (not A300) );
 a37185a <=( (not A269)  and  a37184a );
 a37186a <=( a37185a  and  a37180a );
 a37190a <=( A168  and  (not A169) );
 a37191a <=( A170  and  a37190a );
 a37195a <=( (not A265)  and  A200 );
 a37196a <=( A199  and  a37195a );
 a37197a <=( a37196a  and  a37191a );
 a37201a <=( (not A268)  and  (not A267) );
 a37202a <=( A266  and  a37201a );
 a37206a <=( A302  and  (not A300) );
 a37207a <=( (not A269)  and  a37206a );
 a37208a <=( a37207a  and  a37202a );
 a37212a <=( A168  and  (not A169) );
 a37213a <=( A170  and  a37212a );
 a37217a <=( (not A265)  and  A200 );
 a37218a <=( A199  and  a37217a );
 a37219a <=( a37218a  and  a37213a );
 a37223a <=( (not A268)  and  (not A267) );
 a37224a <=( A266  and  a37223a );
 a37228a <=( A299  and  A298 );
 a37229a <=( (not A269)  and  a37228a );
 a37230a <=( a37229a  and  a37224a );
 a37234a <=( A168  and  (not A169) );
 a37235a <=( A170  and  a37234a );
 a37239a <=( (not A265)  and  A200 );
 a37240a <=( A199  and  a37239a );
 a37241a <=( a37240a  and  a37235a );
 a37245a <=( (not A268)  and  (not A267) );
 a37246a <=( A266  and  a37245a );
 a37250a <=( (not A299)  and  (not A298) );
 a37251a <=( (not A269)  and  a37250a );
 a37252a <=( a37251a  and  a37246a );
 a37256a <=( A168  and  (not A169) );
 a37257a <=( A170  and  a37256a );
 a37261a <=( A265  and  A200 );
 a37262a <=( A199  and  a37261a );
 a37263a <=( a37262a  and  a37257a );
 a37267a <=( A268  and  A267 );
 a37268a <=( (not A266)  and  a37267a );
 a37272a <=( (not A302)  and  (not A301) );
 a37273a <=( A300  and  a37272a );
 a37274a <=( a37273a  and  a37268a );
 a37278a <=( A168  and  (not A169) );
 a37279a <=( A170  and  a37278a );
 a37283a <=( A265  and  A200 );
 a37284a <=( A199  and  a37283a );
 a37285a <=( a37284a  and  a37279a );
 a37289a <=( A269  and  A267 );
 a37290a <=( (not A266)  and  a37289a );
 a37294a <=( (not A302)  and  (not A301) );
 a37295a <=( A300  and  a37294a );
 a37296a <=( a37295a  and  a37290a );
 a37300a <=( A168  and  (not A169) );
 a37301a <=( A170  and  a37300a );
 a37305a <=( A265  and  A200 );
 a37306a <=( A199  and  a37305a );
 a37307a <=( a37306a  and  a37301a );
 a37311a <=( (not A268)  and  (not A267) );
 a37312a <=( (not A266)  and  a37311a );
 a37316a <=( A301  and  (not A300) );
 a37317a <=( (not A269)  and  a37316a );
 a37318a <=( a37317a  and  a37312a );
 a37322a <=( A168  and  (not A169) );
 a37323a <=( A170  and  a37322a );
 a37327a <=( A265  and  A200 );
 a37328a <=( A199  and  a37327a );
 a37329a <=( a37328a  and  a37323a );
 a37333a <=( (not A268)  and  (not A267) );
 a37334a <=( (not A266)  and  a37333a );
 a37338a <=( A302  and  (not A300) );
 a37339a <=( (not A269)  and  a37338a );
 a37340a <=( a37339a  and  a37334a );
 a37344a <=( A168  and  (not A169) );
 a37345a <=( A170  and  a37344a );
 a37349a <=( A265  and  A200 );
 a37350a <=( A199  and  a37349a );
 a37351a <=( a37350a  and  a37345a );
 a37355a <=( (not A268)  and  (not A267) );
 a37356a <=( (not A266)  and  a37355a );
 a37360a <=( A299  and  A298 );
 a37361a <=( (not A269)  and  a37360a );
 a37362a <=( a37361a  and  a37356a );
 a37366a <=( A168  and  (not A169) );
 a37367a <=( A170  and  a37366a );
 a37371a <=( A265  and  A200 );
 a37372a <=( A199  and  a37371a );
 a37373a <=( a37372a  and  a37367a );
 a37377a <=( (not A268)  and  (not A267) );
 a37378a <=( (not A266)  and  a37377a );
 a37382a <=( (not A299)  and  (not A298) );
 a37383a <=( (not A269)  and  a37382a );
 a37384a <=( a37383a  and  a37378a );
 a37388a <=( A168  and  (not A169) );
 a37389a <=( A170  and  a37388a );
 a37393a <=( (not A265)  and  (not A200) );
 a37394a <=( (not A199)  and  a37393a );
 a37395a <=( a37394a  and  a37389a );
 a37399a <=( A268  and  A267 );
 a37400a <=( A266  and  a37399a );
 a37404a <=( (not A302)  and  (not A301) );
 a37405a <=( A300  and  a37404a );
 a37406a <=( a37405a  and  a37400a );
 a37410a <=( A168  and  (not A169) );
 a37411a <=( A170  and  a37410a );
 a37415a <=( (not A265)  and  (not A200) );
 a37416a <=( (not A199)  and  a37415a );
 a37417a <=( a37416a  and  a37411a );
 a37421a <=( A269  and  A267 );
 a37422a <=( A266  and  a37421a );
 a37426a <=( (not A302)  and  (not A301) );
 a37427a <=( A300  and  a37426a );
 a37428a <=( a37427a  and  a37422a );
 a37432a <=( A168  and  (not A169) );
 a37433a <=( A170  and  a37432a );
 a37437a <=( (not A265)  and  (not A200) );
 a37438a <=( (not A199)  and  a37437a );
 a37439a <=( a37438a  and  a37433a );
 a37443a <=( (not A268)  and  (not A267) );
 a37444a <=( A266  and  a37443a );
 a37448a <=( A301  and  (not A300) );
 a37449a <=( (not A269)  and  a37448a );
 a37450a <=( a37449a  and  a37444a );
 a37454a <=( A168  and  (not A169) );
 a37455a <=( A170  and  a37454a );
 a37459a <=( (not A265)  and  (not A200) );
 a37460a <=( (not A199)  and  a37459a );
 a37461a <=( a37460a  and  a37455a );
 a37465a <=( (not A268)  and  (not A267) );
 a37466a <=( A266  and  a37465a );
 a37470a <=( A302  and  (not A300) );
 a37471a <=( (not A269)  and  a37470a );
 a37472a <=( a37471a  and  a37466a );
 a37476a <=( A168  and  (not A169) );
 a37477a <=( A170  and  a37476a );
 a37481a <=( (not A265)  and  (not A200) );
 a37482a <=( (not A199)  and  a37481a );
 a37483a <=( a37482a  and  a37477a );
 a37487a <=( (not A268)  and  (not A267) );
 a37488a <=( A266  and  a37487a );
 a37492a <=( A299  and  A298 );
 a37493a <=( (not A269)  and  a37492a );
 a37494a <=( a37493a  and  a37488a );
 a37498a <=( A168  and  (not A169) );
 a37499a <=( A170  and  a37498a );
 a37503a <=( (not A265)  and  (not A200) );
 a37504a <=( (not A199)  and  a37503a );
 a37505a <=( a37504a  and  a37499a );
 a37509a <=( (not A268)  and  (not A267) );
 a37510a <=( A266  and  a37509a );
 a37514a <=( (not A299)  and  (not A298) );
 a37515a <=( (not A269)  and  a37514a );
 a37516a <=( a37515a  and  a37510a );
 a37520a <=( A168  and  (not A169) );
 a37521a <=( A170  and  a37520a );
 a37525a <=( A265  and  (not A200) );
 a37526a <=( (not A199)  and  a37525a );
 a37527a <=( a37526a  and  a37521a );
 a37531a <=( A268  and  A267 );
 a37532a <=( (not A266)  and  a37531a );
 a37536a <=( (not A302)  and  (not A301) );
 a37537a <=( A300  and  a37536a );
 a37538a <=( a37537a  and  a37532a );
 a37542a <=( A168  and  (not A169) );
 a37543a <=( A170  and  a37542a );
 a37547a <=( A265  and  (not A200) );
 a37548a <=( (not A199)  and  a37547a );
 a37549a <=( a37548a  and  a37543a );
 a37553a <=( A269  and  A267 );
 a37554a <=( (not A266)  and  a37553a );
 a37558a <=( (not A302)  and  (not A301) );
 a37559a <=( A300  and  a37558a );
 a37560a <=( a37559a  and  a37554a );
 a37564a <=( A168  and  (not A169) );
 a37565a <=( A170  and  a37564a );
 a37569a <=( A265  and  (not A200) );
 a37570a <=( (not A199)  and  a37569a );
 a37571a <=( a37570a  and  a37565a );
 a37575a <=( (not A268)  and  (not A267) );
 a37576a <=( (not A266)  and  a37575a );
 a37580a <=( A301  and  (not A300) );
 a37581a <=( (not A269)  and  a37580a );
 a37582a <=( a37581a  and  a37576a );
 a37586a <=( A168  and  (not A169) );
 a37587a <=( A170  and  a37586a );
 a37591a <=( A265  and  (not A200) );
 a37592a <=( (not A199)  and  a37591a );
 a37593a <=( a37592a  and  a37587a );
 a37597a <=( (not A268)  and  (not A267) );
 a37598a <=( (not A266)  and  a37597a );
 a37602a <=( A302  and  (not A300) );
 a37603a <=( (not A269)  and  a37602a );
 a37604a <=( a37603a  and  a37598a );
 a37608a <=( A168  and  (not A169) );
 a37609a <=( A170  and  a37608a );
 a37613a <=( A265  and  (not A200) );
 a37614a <=( (not A199)  and  a37613a );
 a37615a <=( a37614a  and  a37609a );
 a37619a <=( (not A268)  and  (not A267) );
 a37620a <=( (not A266)  and  a37619a );
 a37624a <=( A299  and  A298 );
 a37625a <=( (not A269)  and  a37624a );
 a37626a <=( a37625a  and  a37620a );
 a37630a <=( A168  and  (not A169) );
 a37631a <=( A170  and  a37630a );
 a37635a <=( A265  and  (not A200) );
 a37636a <=( (not A199)  and  a37635a );
 a37637a <=( a37636a  and  a37631a );
 a37641a <=( (not A268)  and  (not A267) );
 a37642a <=( (not A266)  and  a37641a );
 a37646a <=( (not A299)  and  (not A298) );
 a37647a <=( (not A269)  and  a37646a );
 a37648a <=( a37647a  and  a37642a );
 a37652a <=( A201  and  A166 );
 a37653a <=( A167  and  a37652a );
 a37657a <=( (not A265)  and  (not A203) );
 a37658a <=( (not A202)  and  a37657a );
 a37659a <=( a37658a  and  a37653a );
 a37663a <=( (not A268)  and  (not A267) );
 a37664a <=( A266  and  a37663a );
 a37667a <=( A300  and  (not A269) );
 a37670a <=( (not A302)  and  (not A301) );
 a37671a <=( a37670a  and  a37667a );
 a37672a <=( a37671a  and  a37664a );
 a37676a <=( A201  and  A166 );
 a37677a <=( A167  and  a37676a );
 a37681a <=( A265  and  (not A203) );
 a37682a <=( (not A202)  and  a37681a );
 a37683a <=( a37682a  and  a37677a );
 a37687a <=( (not A268)  and  (not A267) );
 a37688a <=( (not A266)  and  a37687a );
 a37691a <=( A300  and  (not A269) );
 a37694a <=( (not A302)  and  (not A301) );
 a37695a <=( a37694a  and  a37691a );
 a37696a <=( a37695a  and  a37688a );
 a37700a <=( (not A199)  and  A166 );
 a37701a <=( A167  and  a37700a );
 a37705a <=( A202  and  A201 );
 a37706a <=( A200  and  a37705a );
 a37707a <=( a37706a  and  a37701a );
 a37711a <=( (not A269)  and  (not A268) );
 a37712a <=( A267  and  a37711a );
 a37715a <=( (not A299)  and  A298 );
 a37718a <=( A301  and  A300 );
 a37719a <=( a37718a  and  a37715a );
 a37720a <=( a37719a  and  a37712a );
 a37724a <=( (not A199)  and  A166 );
 a37725a <=( A167  and  a37724a );
 a37729a <=( A202  and  A201 );
 a37730a <=( A200  and  a37729a );
 a37731a <=( a37730a  and  a37725a );
 a37735a <=( (not A269)  and  (not A268) );
 a37736a <=( A267  and  a37735a );
 a37739a <=( (not A299)  and  A298 );
 a37742a <=( A302  and  A300 );
 a37743a <=( a37742a  and  a37739a );
 a37744a <=( a37743a  and  a37736a );
 a37748a <=( (not A199)  and  A166 );
 a37749a <=( A167  and  a37748a );
 a37753a <=( A202  and  A201 );
 a37754a <=( A200  and  a37753a );
 a37755a <=( a37754a  and  a37749a );
 a37759a <=( (not A269)  and  (not A268) );
 a37760a <=( A267  and  a37759a );
 a37763a <=( A299  and  (not A298) );
 a37766a <=( A301  and  A300 );
 a37767a <=( a37766a  and  a37763a );
 a37768a <=( a37767a  and  a37760a );
 a37772a <=( (not A199)  and  A166 );
 a37773a <=( A167  and  a37772a );
 a37777a <=( A202  and  A201 );
 a37778a <=( A200  and  a37777a );
 a37779a <=( a37778a  and  a37773a );
 a37783a <=( (not A269)  and  (not A268) );
 a37784a <=( A267  and  a37783a );
 a37787a <=( A299  and  (not A298) );
 a37790a <=( A302  and  A300 );
 a37791a <=( a37790a  and  a37787a );
 a37792a <=( a37791a  and  a37784a );
 a37796a <=( (not A199)  and  A166 );
 a37797a <=( A167  and  a37796a );
 a37801a <=( A202  and  A201 );
 a37802a <=( A200  and  a37801a );
 a37803a <=( a37802a  and  a37797a );
 a37807a <=( A298  and  A268 );
 a37808a <=( (not A267)  and  a37807a );
 a37811a <=( (not A300)  and  (not A299) );
 a37814a <=( (not A302)  and  (not A301) );
 a37815a <=( a37814a  and  a37811a );
 a37816a <=( a37815a  and  a37808a );
 a37820a <=( (not A199)  and  A166 );
 a37821a <=( A167  and  a37820a );
 a37825a <=( A202  and  A201 );
 a37826a <=( A200  and  a37825a );
 a37827a <=( a37826a  and  a37821a );
 a37831a <=( (not A298)  and  A268 );
 a37832a <=( (not A267)  and  a37831a );
 a37835a <=( (not A300)  and  A299 );
 a37838a <=( (not A302)  and  (not A301) );
 a37839a <=( a37838a  and  a37835a );
 a37840a <=( a37839a  and  a37832a );
 a37844a <=( (not A199)  and  A166 );
 a37845a <=( A167  and  a37844a );
 a37849a <=( A202  and  A201 );
 a37850a <=( A200  and  a37849a );
 a37851a <=( a37850a  and  a37845a );
 a37855a <=( A298  and  A269 );
 a37856a <=( (not A267)  and  a37855a );
 a37859a <=( (not A300)  and  (not A299) );
 a37862a <=( (not A302)  and  (not A301) );
 a37863a <=( a37862a  and  a37859a );
 a37864a <=( a37863a  and  a37856a );
 a37868a <=( (not A199)  and  A166 );
 a37869a <=( A167  and  a37868a );
 a37873a <=( A202  and  A201 );
 a37874a <=( A200  and  a37873a );
 a37875a <=( a37874a  and  a37869a );
 a37879a <=( (not A298)  and  A269 );
 a37880a <=( (not A267)  and  a37879a );
 a37883a <=( (not A300)  and  A299 );
 a37886a <=( (not A302)  and  (not A301) );
 a37887a <=( a37886a  and  a37883a );
 a37888a <=( a37887a  and  a37880a );
 a37892a <=( (not A199)  and  A166 );
 a37893a <=( A167  and  a37892a );
 a37897a <=( A202  and  A201 );
 a37898a <=( A200  and  a37897a );
 a37899a <=( a37898a  and  a37893a );
 a37903a <=( A298  and  A266 );
 a37904a <=( A265  and  a37903a );
 a37907a <=( (not A300)  and  (not A299) );
 a37910a <=( (not A302)  and  (not A301) );
 a37911a <=( a37910a  and  a37907a );
 a37912a <=( a37911a  and  a37904a );
 a37916a <=( (not A199)  and  A166 );
 a37917a <=( A167  and  a37916a );
 a37921a <=( A202  and  A201 );
 a37922a <=( A200  and  a37921a );
 a37923a <=( a37922a  and  a37917a );
 a37927a <=( (not A298)  and  A266 );
 a37928a <=( A265  and  a37927a );
 a37931a <=( (not A300)  and  A299 );
 a37934a <=( (not A302)  and  (not A301) );
 a37935a <=( a37934a  and  a37931a );
 a37936a <=( a37935a  and  a37928a );
 a37940a <=( (not A199)  and  A166 );
 a37941a <=( A167  and  a37940a );
 a37945a <=( A202  and  A201 );
 a37946a <=( A200  and  a37945a );
 a37947a <=( a37946a  and  a37941a );
 a37951a <=( A298  and  (not A266) );
 a37952a <=( (not A265)  and  a37951a );
 a37955a <=( (not A300)  and  (not A299) );
 a37958a <=( (not A302)  and  (not A301) );
 a37959a <=( a37958a  and  a37955a );
 a37960a <=( a37959a  and  a37952a );
 a37964a <=( (not A199)  and  A166 );
 a37965a <=( A167  and  a37964a );
 a37969a <=( A202  and  A201 );
 a37970a <=( A200  and  a37969a );
 a37971a <=( a37970a  and  a37965a );
 a37975a <=( (not A298)  and  (not A266) );
 a37976a <=( (not A265)  and  a37975a );
 a37979a <=( (not A300)  and  A299 );
 a37982a <=( (not A302)  and  (not A301) );
 a37983a <=( a37982a  and  a37979a );
 a37984a <=( a37983a  and  a37976a );
 a37988a <=( (not A199)  and  A166 );
 a37989a <=( A167  and  a37988a );
 a37993a <=( A203  and  A201 );
 a37994a <=( A200  and  a37993a );
 a37995a <=( a37994a  and  a37989a );
 a37999a <=( (not A269)  and  (not A268) );
 a38000a <=( A267  and  a37999a );
 a38003a <=( (not A299)  and  A298 );
 a38006a <=( A301  and  A300 );
 a38007a <=( a38006a  and  a38003a );
 a38008a <=( a38007a  and  a38000a );
 a38012a <=( (not A199)  and  A166 );
 a38013a <=( A167  and  a38012a );
 a38017a <=( A203  and  A201 );
 a38018a <=( A200  and  a38017a );
 a38019a <=( a38018a  and  a38013a );
 a38023a <=( (not A269)  and  (not A268) );
 a38024a <=( A267  and  a38023a );
 a38027a <=( (not A299)  and  A298 );
 a38030a <=( A302  and  A300 );
 a38031a <=( a38030a  and  a38027a );
 a38032a <=( a38031a  and  a38024a );
 a38036a <=( (not A199)  and  A166 );
 a38037a <=( A167  and  a38036a );
 a38041a <=( A203  and  A201 );
 a38042a <=( A200  and  a38041a );
 a38043a <=( a38042a  and  a38037a );
 a38047a <=( (not A269)  and  (not A268) );
 a38048a <=( A267  and  a38047a );
 a38051a <=( A299  and  (not A298) );
 a38054a <=( A301  and  A300 );
 a38055a <=( a38054a  and  a38051a );
 a38056a <=( a38055a  and  a38048a );
 a38060a <=( (not A199)  and  A166 );
 a38061a <=( A167  and  a38060a );
 a38065a <=( A203  and  A201 );
 a38066a <=( A200  and  a38065a );
 a38067a <=( a38066a  and  a38061a );
 a38071a <=( (not A269)  and  (not A268) );
 a38072a <=( A267  and  a38071a );
 a38075a <=( A299  and  (not A298) );
 a38078a <=( A302  and  A300 );
 a38079a <=( a38078a  and  a38075a );
 a38080a <=( a38079a  and  a38072a );
 a38084a <=( (not A199)  and  A166 );
 a38085a <=( A167  and  a38084a );
 a38089a <=( A203  and  A201 );
 a38090a <=( A200  and  a38089a );
 a38091a <=( a38090a  and  a38085a );
 a38095a <=( A298  and  A268 );
 a38096a <=( (not A267)  and  a38095a );
 a38099a <=( (not A300)  and  (not A299) );
 a38102a <=( (not A302)  and  (not A301) );
 a38103a <=( a38102a  and  a38099a );
 a38104a <=( a38103a  and  a38096a );
 a38108a <=( (not A199)  and  A166 );
 a38109a <=( A167  and  a38108a );
 a38113a <=( A203  and  A201 );
 a38114a <=( A200  and  a38113a );
 a38115a <=( a38114a  and  a38109a );
 a38119a <=( (not A298)  and  A268 );
 a38120a <=( (not A267)  and  a38119a );
 a38123a <=( (not A300)  and  A299 );
 a38126a <=( (not A302)  and  (not A301) );
 a38127a <=( a38126a  and  a38123a );
 a38128a <=( a38127a  and  a38120a );
 a38132a <=( (not A199)  and  A166 );
 a38133a <=( A167  and  a38132a );
 a38137a <=( A203  and  A201 );
 a38138a <=( A200  and  a38137a );
 a38139a <=( a38138a  and  a38133a );
 a38143a <=( A298  and  A269 );
 a38144a <=( (not A267)  and  a38143a );
 a38147a <=( (not A300)  and  (not A299) );
 a38150a <=( (not A302)  and  (not A301) );
 a38151a <=( a38150a  and  a38147a );
 a38152a <=( a38151a  and  a38144a );
 a38156a <=( (not A199)  and  A166 );
 a38157a <=( A167  and  a38156a );
 a38161a <=( A203  and  A201 );
 a38162a <=( A200  and  a38161a );
 a38163a <=( a38162a  and  a38157a );
 a38167a <=( (not A298)  and  A269 );
 a38168a <=( (not A267)  and  a38167a );
 a38171a <=( (not A300)  and  A299 );
 a38174a <=( (not A302)  and  (not A301) );
 a38175a <=( a38174a  and  a38171a );
 a38176a <=( a38175a  and  a38168a );
 a38180a <=( (not A199)  and  A166 );
 a38181a <=( A167  and  a38180a );
 a38185a <=( A203  and  A201 );
 a38186a <=( A200  and  a38185a );
 a38187a <=( a38186a  and  a38181a );
 a38191a <=( A298  and  A266 );
 a38192a <=( A265  and  a38191a );
 a38195a <=( (not A300)  and  (not A299) );
 a38198a <=( (not A302)  and  (not A301) );
 a38199a <=( a38198a  and  a38195a );
 a38200a <=( a38199a  and  a38192a );
 a38204a <=( (not A199)  and  A166 );
 a38205a <=( A167  and  a38204a );
 a38209a <=( A203  and  A201 );
 a38210a <=( A200  and  a38209a );
 a38211a <=( a38210a  and  a38205a );
 a38215a <=( (not A298)  and  A266 );
 a38216a <=( A265  and  a38215a );
 a38219a <=( (not A300)  and  A299 );
 a38222a <=( (not A302)  and  (not A301) );
 a38223a <=( a38222a  and  a38219a );
 a38224a <=( a38223a  and  a38216a );
 a38228a <=( (not A199)  and  A166 );
 a38229a <=( A167  and  a38228a );
 a38233a <=( A203  and  A201 );
 a38234a <=( A200  and  a38233a );
 a38235a <=( a38234a  and  a38229a );
 a38239a <=( A298  and  (not A266) );
 a38240a <=( (not A265)  and  a38239a );
 a38243a <=( (not A300)  and  (not A299) );
 a38246a <=( (not A302)  and  (not A301) );
 a38247a <=( a38246a  and  a38243a );
 a38248a <=( a38247a  and  a38240a );
 a38252a <=( (not A199)  and  A166 );
 a38253a <=( A167  and  a38252a );
 a38257a <=( A203  and  A201 );
 a38258a <=( A200  and  a38257a );
 a38259a <=( a38258a  and  a38253a );
 a38263a <=( (not A298)  and  (not A266) );
 a38264a <=( (not A265)  and  a38263a );
 a38267a <=( (not A300)  and  A299 );
 a38270a <=( (not A302)  and  (not A301) );
 a38271a <=( a38270a  and  a38267a );
 a38272a <=( a38271a  and  a38264a );
 a38276a <=( (not A199)  and  A166 );
 a38277a <=( A167  and  a38276a );
 a38281a <=( (not A202)  and  (not A201) );
 a38282a <=( A200  and  a38281a );
 a38283a <=( a38282a  and  a38277a );
 a38287a <=( A268  and  (not A267) );
 a38288a <=( (not A203)  and  a38287a );
 a38291a <=( (not A299)  and  A298 );
 a38294a <=( A301  and  A300 );
 a38295a <=( a38294a  and  a38291a );
 a38296a <=( a38295a  and  a38288a );
 a38300a <=( (not A199)  and  A166 );
 a38301a <=( A167  and  a38300a );
 a38305a <=( (not A202)  and  (not A201) );
 a38306a <=( A200  and  a38305a );
 a38307a <=( a38306a  and  a38301a );
 a38311a <=( A268  and  (not A267) );
 a38312a <=( (not A203)  and  a38311a );
 a38315a <=( (not A299)  and  A298 );
 a38318a <=( A302  and  A300 );
 a38319a <=( a38318a  and  a38315a );
 a38320a <=( a38319a  and  a38312a );
 a38324a <=( (not A199)  and  A166 );
 a38325a <=( A167  and  a38324a );
 a38329a <=( (not A202)  and  (not A201) );
 a38330a <=( A200  and  a38329a );
 a38331a <=( a38330a  and  a38325a );
 a38335a <=( A268  and  (not A267) );
 a38336a <=( (not A203)  and  a38335a );
 a38339a <=( A299  and  (not A298) );
 a38342a <=( A301  and  A300 );
 a38343a <=( a38342a  and  a38339a );
 a38344a <=( a38343a  and  a38336a );
 a38348a <=( (not A199)  and  A166 );
 a38349a <=( A167  and  a38348a );
 a38353a <=( (not A202)  and  (not A201) );
 a38354a <=( A200  and  a38353a );
 a38355a <=( a38354a  and  a38349a );
 a38359a <=( A268  and  (not A267) );
 a38360a <=( (not A203)  and  a38359a );
 a38363a <=( A299  and  (not A298) );
 a38366a <=( A302  and  A300 );
 a38367a <=( a38366a  and  a38363a );
 a38368a <=( a38367a  and  a38360a );
 a38372a <=( (not A199)  and  A166 );
 a38373a <=( A167  and  a38372a );
 a38377a <=( (not A202)  and  (not A201) );
 a38378a <=( A200  and  a38377a );
 a38379a <=( a38378a  and  a38373a );
 a38383a <=( A269  and  (not A267) );
 a38384a <=( (not A203)  and  a38383a );
 a38387a <=( (not A299)  and  A298 );
 a38390a <=( A301  and  A300 );
 a38391a <=( a38390a  and  a38387a );
 a38392a <=( a38391a  and  a38384a );
 a38396a <=( (not A199)  and  A166 );
 a38397a <=( A167  and  a38396a );
 a38401a <=( (not A202)  and  (not A201) );
 a38402a <=( A200  and  a38401a );
 a38403a <=( a38402a  and  a38397a );
 a38407a <=( A269  and  (not A267) );
 a38408a <=( (not A203)  and  a38407a );
 a38411a <=( (not A299)  and  A298 );
 a38414a <=( A302  and  A300 );
 a38415a <=( a38414a  and  a38411a );
 a38416a <=( a38415a  and  a38408a );
 a38420a <=( (not A199)  and  A166 );
 a38421a <=( A167  and  a38420a );
 a38425a <=( (not A202)  and  (not A201) );
 a38426a <=( A200  and  a38425a );
 a38427a <=( a38426a  and  a38421a );
 a38431a <=( A269  and  (not A267) );
 a38432a <=( (not A203)  and  a38431a );
 a38435a <=( A299  and  (not A298) );
 a38438a <=( A301  and  A300 );
 a38439a <=( a38438a  and  a38435a );
 a38440a <=( a38439a  and  a38432a );
 a38444a <=( (not A199)  and  A166 );
 a38445a <=( A167  and  a38444a );
 a38449a <=( (not A202)  and  (not A201) );
 a38450a <=( A200  and  a38449a );
 a38451a <=( a38450a  and  a38445a );
 a38455a <=( A269  and  (not A267) );
 a38456a <=( (not A203)  and  a38455a );
 a38459a <=( A299  and  (not A298) );
 a38462a <=( A302  and  A300 );
 a38463a <=( a38462a  and  a38459a );
 a38464a <=( a38463a  and  a38456a );
 a38468a <=( (not A199)  and  A166 );
 a38469a <=( A167  and  a38468a );
 a38473a <=( (not A202)  and  (not A201) );
 a38474a <=( A200  and  a38473a );
 a38475a <=( a38474a  and  a38469a );
 a38479a <=( A266  and  A265 );
 a38480a <=( (not A203)  and  a38479a );
 a38483a <=( (not A299)  and  A298 );
 a38486a <=( A301  and  A300 );
 a38487a <=( a38486a  and  a38483a );
 a38488a <=( a38487a  and  a38480a );
 a38492a <=( (not A199)  and  A166 );
 a38493a <=( A167  and  a38492a );
 a38497a <=( (not A202)  and  (not A201) );
 a38498a <=( A200  and  a38497a );
 a38499a <=( a38498a  and  a38493a );
 a38503a <=( A266  and  A265 );
 a38504a <=( (not A203)  and  a38503a );
 a38507a <=( (not A299)  and  A298 );
 a38510a <=( A302  and  A300 );
 a38511a <=( a38510a  and  a38507a );
 a38512a <=( a38511a  and  a38504a );
 a38516a <=( (not A199)  and  A166 );
 a38517a <=( A167  and  a38516a );
 a38521a <=( (not A202)  and  (not A201) );
 a38522a <=( A200  and  a38521a );
 a38523a <=( a38522a  and  a38517a );
 a38527a <=( A266  and  A265 );
 a38528a <=( (not A203)  and  a38527a );
 a38531a <=( A299  and  (not A298) );
 a38534a <=( A301  and  A300 );
 a38535a <=( a38534a  and  a38531a );
 a38536a <=( a38535a  and  a38528a );
 a38540a <=( (not A199)  and  A166 );
 a38541a <=( A167  and  a38540a );
 a38545a <=( (not A202)  and  (not A201) );
 a38546a <=( A200  and  a38545a );
 a38547a <=( a38546a  and  a38541a );
 a38551a <=( A266  and  A265 );
 a38552a <=( (not A203)  and  a38551a );
 a38555a <=( A299  and  (not A298) );
 a38558a <=( A302  and  A300 );
 a38559a <=( a38558a  and  a38555a );
 a38560a <=( a38559a  and  a38552a );
 a38564a <=( (not A199)  and  A166 );
 a38565a <=( A167  and  a38564a );
 a38569a <=( (not A202)  and  (not A201) );
 a38570a <=( A200  and  a38569a );
 a38571a <=( a38570a  and  a38565a );
 a38575a <=( (not A266)  and  (not A265) );
 a38576a <=( (not A203)  and  a38575a );
 a38579a <=( (not A299)  and  A298 );
 a38582a <=( A301  and  A300 );
 a38583a <=( a38582a  and  a38579a );
 a38584a <=( a38583a  and  a38576a );
 a38588a <=( (not A199)  and  A166 );
 a38589a <=( A167  and  a38588a );
 a38593a <=( (not A202)  and  (not A201) );
 a38594a <=( A200  and  a38593a );
 a38595a <=( a38594a  and  a38589a );
 a38599a <=( (not A266)  and  (not A265) );
 a38600a <=( (not A203)  and  a38599a );
 a38603a <=( (not A299)  and  A298 );
 a38606a <=( A302  and  A300 );
 a38607a <=( a38606a  and  a38603a );
 a38608a <=( a38607a  and  a38600a );
 a38612a <=( (not A199)  and  A166 );
 a38613a <=( A167  and  a38612a );
 a38617a <=( (not A202)  and  (not A201) );
 a38618a <=( A200  and  a38617a );
 a38619a <=( a38618a  and  a38613a );
 a38623a <=( (not A266)  and  (not A265) );
 a38624a <=( (not A203)  and  a38623a );
 a38627a <=( A299  and  (not A298) );
 a38630a <=( A301  and  A300 );
 a38631a <=( a38630a  and  a38627a );
 a38632a <=( a38631a  and  a38624a );
 a38636a <=( (not A199)  and  A166 );
 a38637a <=( A167  and  a38636a );
 a38641a <=( (not A202)  and  (not A201) );
 a38642a <=( A200  and  a38641a );
 a38643a <=( a38642a  and  a38637a );
 a38647a <=( (not A266)  and  (not A265) );
 a38648a <=( (not A203)  and  a38647a );
 a38651a <=( A299  and  (not A298) );
 a38654a <=( A302  and  A300 );
 a38655a <=( a38654a  and  a38651a );
 a38656a <=( a38655a  and  a38648a );
 a38660a <=( A199  and  A166 );
 a38661a <=( A167  and  a38660a );
 a38665a <=( A202  and  A201 );
 a38666a <=( (not A200)  and  a38665a );
 a38667a <=( a38666a  and  a38661a );
 a38671a <=( (not A269)  and  (not A268) );
 a38672a <=( A267  and  a38671a );
 a38675a <=( (not A299)  and  A298 );
 a38678a <=( A301  and  A300 );
 a38679a <=( a38678a  and  a38675a );
 a38680a <=( a38679a  and  a38672a );
 a38684a <=( A199  and  A166 );
 a38685a <=( A167  and  a38684a );
 a38689a <=( A202  and  A201 );
 a38690a <=( (not A200)  and  a38689a );
 a38691a <=( a38690a  and  a38685a );
 a38695a <=( (not A269)  and  (not A268) );
 a38696a <=( A267  and  a38695a );
 a38699a <=( (not A299)  and  A298 );
 a38702a <=( A302  and  A300 );
 a38703a <=( a38702a  and  a38699a );
 a38704a <=( a38703a  and  a38696a );
 a38708a <=( A199  and  A166 );
 a38709a <=( A167  and  a38708a );
 a38713a <=( A202  and  A201 );
 a38714a <=( (not A200)  and  a38713a );
 a38715a <=( a38714a  and  a38709a );
 a38719a <=( (not A269)  and  (not A268) );
 a38720a <=( A267  and  a38719a );
 a38723a <=( A299  and  (not A298) );
 a38726a <=( A301  and  A300 );
 a38727a <=( a38726a  and  a38723a );
 a38728a <=( a38727a  and  a38720a );
 a38732a <=( A199  and  A166 );
 a38733a <=( A167  and  a38732a );
 a38737a <=( A202  and  A201 );
 a38738a <=( (not A200)  and  a38737a );
 a38739a <=( a38738a  and  a38733a );
 a38743a <=( (not A269)  and  (not A268) );
 a38744a <=( A267  and  a38743a );
 a38747a <=( A299  and  (not A298) );
 a38750a <=( A302  and  A300 );
 a38751a <=( a38750a  and  a38747a );
 a38752a <=( a38751a  and  a38744a );
 a38756a <=( A199  and  A166 );
 a38757a <=( A167  and  a38756a );
 a38761a <=( A202  and  A201 );
 a38762a <=( (not A200)  and  a38761a );
 a38763a <=( a38762a  and  a38757a );
 a38767a <=( A298  and  A268 );
 a38768a <=( (not A267)  and  a38767a );
 a38771a <=( (not A300)  and  (not A299) );
 a38774a <=( (not A302)  and  (not A301) );
 a38775a <=( a38774a  and  a38771a );
 a38776a <=( a38775a  and  a38768a );
 a38780a <=( A199  and  A166 );
 a38781a <=( A167  and  a38780a );
 a38785a <=( A202  and  A201 );
 a38786a <=( (not A200)  and  a38785a );
 a38787a <=( a38786a  and  a38781a );
 a38791a <=( (not A298)  and  A268 );
 a38792a <=( (not A267)  and  a38791a );
 a38795a <=( (not A300)  and  A299 );
 a38798a <=( (not A302)  and  (not A301) );
 a38799a <=( a38798a  and  a38795a );
 a38800a <=( a38799a  and  a38792a );
 a38804a <=( A199  and  A166 );
 a38805a <=( A167  and  a38804a );
 a38809a <=( A202  and  A201 );
 a38810a <=( (not A200)  and  a38809a );
 a38811a <=( a38810a  and  a38805a );
 a38815a <=( A298  and  A269 );
 a38816a <=( (not A267)  and  a38815a );
 a38819a <=( (not A300)  and  (not A299) );
 a38822a <=( (not A302)  and  (not A301) );
 a38823a <=( a38822a  and  a38819a );
 a38824a <=( a38823a  and  a38816a );
 a38828a <=( A199  and  A166 );
 a38829a <=( A167  and  a38828a );
 a38833a <=( A202  and  A201 );
 a38834a <=( (not A200)  and  a38833a );
 a38835a <=( a38834a  and  a38829a );
 a38839a <=( (not A298)  and  A269 );
 a38840a <=( (not A267)  and  a38839a );
 a38843a <=( (not A300)  and  A299 );
 a38846a <=( (not A302)  and  (not A301) );
 a38847a <=( a38846a  and  a38843a );
 a38848a <=( a38847a  and  a38840a );
 a38852a <=( A199  and  A166 );
 a38853a <=( A167  and  a38852a );
 a38857a <=( A202  and  A201 );
 a38858a <=( (not A200)  and  a38857a );
 a38859a <=( a38858a  and  a38853a );
 a38863a <=( A298  and  A266 );
 a38864a <=( A265  and  a38863a );
 a38867a <=( (not A300)  and  (not A299) );
 a38870a <=( (not A302)  and  (not A301) );
 a38871a <=( a38870a  and  a38867a );
 a38872a <=( a38871a  and  a38864a );
 a38876a <=( A199  and  A166 );
 a38877a <=( A167  and  a38876a );
 a38881a <=( A202  and  A201 );
 a38882a <=( (not A200)  and  a38881a );
 a38883a <=( a38882a  and  a38877a );
 a38887a <=( (not A298)  and  A266 );
 a38888a <=( A265  and  a38887a );
 a38891a <=( (not A300)  and  A299 );
 a38894a <=( (not A302)  and  (not A301) );
 a38895a <=( a38894a  and  a38891a );
 a38896a <=( a38895a  and  a38888a );
 a38900a <=( A199  and  A166 );
 a38901a <=( A167  and  a38900a );
 a38905a <=( A202  and  A201 );
 a38906a <=( (not A200)  and  a38905a );
 a38907a <=( a38906a  and  a38901a );
 a38911a <=( A298  and  (not A266) );
 a38912a <=( (not A265)  and  a38911a );
 a38915a <=( (not A300)  and  (not A299) );
 a38918a <=( (not A302)  and  (not A301) );
 a38919a <=( a38918a  and  a38915a );
 a38920a <=( a38919a  and  a38912a );
 a38924a <=( A199  and  A166 );
 a38925a <=( A167  and  a38924a );
 a38929a <=( A202  and  A201 );
 a38930a <=( (not A200)  and  a38929a );
 a38931a <=( a38930a  and  a38925a );
 a38935a <=( (not A298)  and  (not A266) );
 a38936a <=( (not A265)  and  a38935a );
 a38939a <=( (not A300)  and  A299 );
 a38942a <=( (not A302)  and  (not A301) );
 a38943a <=( a38942a  and  a38939a );
 a38944a <=( a38943a  and  a38936a );
 a38948a <=( A199  and  A166 );
 a38949a <=( A167  and  a38948a );
 a38953a <=( A203  and  A201 );
 a38954a <=( (not A200)  and  a38953a );
 a38955a <=( a38954a  and  a38949a );
 a38959a <=( (not A269)  and  (not A268) );
 a38960a <=( A267  and  a38959a );
 a38963a <=( (not A299)  and  A298 );
 a38966a <=( A301  and  A300 );
 a38967a <=( a38966a  and  a38963a );
 a38968a <=( a38967a  and  a38960a );
 a38972a <=( A199  and  A166 );
 a38973a <=( A167  and  a38972a );
 a38977a <=( A203  and  A201 );
 a38978a <=( (not A200)  and  a38977a );
 a38979a <=( a38978a  and  a38973a );
 a38983a <=( (not A269)  and  (not A268) );
 a38984a <=( A267  and  a38983a );
 a38987a <=( (not A299)  and  A298 );
 a38990a <=( A302  and  A300 );
 a38991a <=( a38990a  and  a38987a );
 a38992a <=( a38991a  and  a38984a );
 a38996a <=( A199  and  A166 );
 a38997a <=( A167  and  a38996a );
 a39001a <=( A203  and  A201 );
 a39002a <=( (not A200)  and  a39001a );
 a39003a <=( a39002a  and  a38997a );
 a39007a <=( (not A269)  and  (not A268) );
 a39008a <=( A267  and  a39007a );
 a39011a <=( A299  and  (not A298) );
 a39014a <=( A301  and  A300 );
 a39015a <=( a39014a  and  a39011a );
 a39016a <=( a39015a  and  a39008a );
 a39020a <=( A199  and  A166 );
 a39021a <=( A167  and  a39020a );
 a39025a <=( A203  and  A201 );
 a39026a <=( (not A200)  and  a39025a );
 a39027a <=( a39026a  and  a39021a );
 a39031a <=( (not A269)  and  (not A268) );
 a39032a <=( A267  and  a39031a );
 a39035a <=( A299  and  (not A298) );
 a39038a <=( A302  and  A300 );
 a39039a <=( a39038a  and  a39035a );
 a39040a <=( a39039a  and  a39032a );
 a39044a <=( A199  and  A166 );
 a39045a <=( A167  and  a39044a );
 a39049a <=( A203  and  A201 );
 a39050a <=( (not A200)  and  a39049a );
 a39051a <=( a39050a  and  a39045a );
 a39055a <=( A298  and  A268 );
 a39056a <=( (not A267)  and  a39055a );
 a39059a <=( (not A300)  and  (not A299) );
 a39062a <=( (not A302)  and  (not A301) );
 a39063a <=( a39062a  and  a39059a );
 a39064a <=( a39063a  and  a39056a );
 a39068a <=( A199  and  A166 );
 a39069a <=( A167  and  a39068a );
 a39073a <=( A203  and  A201 );
 a39074a <=( (not A200)  and  a39073a );
 a39075a <=( a39074a  and  a39069a );
 a39079a <=( (not A298)  and  A268 );
 a39080a <=( (not A267)  and  a39079a );
 a39083a <=( (not A300)  and  A299 );
 a39086a <=( (not A302)  and  (not A301) );
 a39087a <=( a39086a  and  a39083a );
 a39088a <=( a39087a  and  a39080a );
 a39092a <=( A199  and  A166 );
 a39093a <=( A167  and  a39092a );
 a39097a <=( A203  and  A201 );
 a39098a <=( (not A200)  and  a39097a );
 a39099a <=( a39098a  and  a39093a );
 a39103a <=( A298  and  A269 );
 a39104a <=( (not A267)  and  a39103a );
 a39107a <=( (not A300)  and  (not A299) );
 a39110a <=( (not A302)  and  (not A301) );
 a39111a <=( a39110a  and  a39107a );
 a39112a <=( a39111a  and  a39104a );
 a39116a <=( A199  and  A166 );
 a39117a <=( A167  and  a39116a );
 a39121a <=( A203  and  A201 );
 a39122a <=( (not A200)  and  a39121a );
 a39123a <=( a39122a  and  a39117a );
 a39127a <=( (not A298)  and  A269 );
 a39128a <=( (not A267)  and  a39127a );
 a39131a <=( (not A300)  and  A299 );
 a39134a <=( (not A302)  and  (not A301) );
 a39135a <=( a39134a  and  a39131a );
 a39136a <=( a39135a  and  a39128a );
 a39140a <=( A199  and  A166 );
 a39141a <=( A167  and  a39140a );
 a39145a <=( A203  and  A201 );
 a39146a <=( (not A200)  and  a39145a );
 a39147a <=( a39146a  and  a39141a );
 a39151a <=( A298  and  A266 );
 a39152a <=( A265  and  a39151a );
 a39155a <=( (not A300)  and  (not A299) );
 a39158a <=( (not A302)  and  (not A301) );
 a39159a <=( a39158a  and  a39155a );
 a39160a <=( a39159a  and  a39152a );
 a39164a <=( A199  and  A166 );
 a39165a <=( A167  and  a39164a );
 a39169a <=( A203  and  A201 );
 a39170a <=( (not A200)  and  a39169a );
 a39171a <=( a39170a  and  a39165a );
 a39175a <=( (not A298)  and  A266 );
 a39176a <=( A265  and  a39175a );
 a39179a <=( (not A300)  and  A299 );
 a39182a <=( (not A302)  and  (not A301) );
 a39183a <=( a39182a  and  a39179a );
 a39184a <=( a39183a  and  a39176a );
 a39188a <=( A199  and  A166 );
 a39189a <=( A167  and  a39188a );
 a39193a <=( A203  and  A201 );
 a39194a <=( (not A200)  and  a39193a );
 a39195a <=( a39194a  and  a39189a );
 a39199a <=( A298  and  (not A266) );
 a39200a <=( (not A265)  and  a39199a );
 a39203a <=( (not A300)  and  (not A299) );
 a39206a <=( (not A302)  and  (not A301) );
 a39207a <=( a39206a  and  a39203a );
 a39208a <=( a39207a  and  a39200a );
 a39212a <=( A199  and  A166 );
 a39213a <=( A167  and  a39212a );
 a39217a <=( A203  and  A201 );
 a39218a <=( (not A200)  and  a39217a );
 a39219a <=( a39218a  and  a39213a );
 a39223a <=( (not A298)  and  (not A266) );
 a39224a <=( (not A265)  and  a39223a );
 a39227a <=( (not A300)  and  A299 );
 a39230a <=( (not A302)  and  (not A301) );
 a39231a <=( a39230a  and  a39227a );
 a39232a <=( a39231a  and  a39224a );
 a39236a <=( A199  and  A166 );
 a39237a <=( A167  and  a39236a );
 a39241a <=( (not A202)  and  (not A201) );
 a39242a <=( (not A200)  and  a39241a );
 a39243a <=( a39242a  and  a39237a );
 a39247a <=( A268  and  (not A267) );
 a39248a <=( (not A203)  and  a39247a );
 a39251a <=( (not A299)  and  A298 );
 a39254a <=( A301  and  A300 );
 a39255a <=( a39254a  and  a39251a );
 a39256a <=( a39255a  and  a39248a );
 a39260a <=( A199  and  A166 );
 a39261a <=( A167  and  a39260a );
 a39265a <=( (not A202)  and  (not A201) );
 a39266a <=( (not A200)  and  a39265a );
 a39267a <=( a39266a  and  a39261a );
 a39271a <=( A268  and  (not A267) );
 a39272a <=( (not A203)  and  a39271a );
 a39275a <=( (not A299)  and  A298 );
 a39278a <=( A302  and  A300 );
 a39279a <=( a39278a  and  a39275a );
 a39280a <=( a39279a  and  a39272a );
 a39284a <=( A199  and  A166 );
 a39285a <=( A167  and  a39284a );
 a39289a <=( (not A202)  and  (not A201) );
 a39290a <=( (not A200)  and  a39289a );
 a39291a <=( a39290a  and  a39285a );
 a39295a <=( A268  and  (not A267) );
 a39296a <=( (not A203)  and  a39295a );
 a39299a <=( A299  and  (not A298) );
 a39302a <=( A301  and  A300 );
 a39303a <=( a39302a  and  a39299a );
 a39304a <=( a39303a  and  a39296a );
 a39308a <=( A199  and  A166 );
 a39309a <=( A167  and  a39308a );
 a39313a <=( (not A202)  and  (not A201) );
 a39314a <=( (not A200)  and  a39313a );
 a39315a <=( a39314a  and  a39309a );
 a39319a <=( A268  and  (not A267) );
 a39320a <=( (not A203)  and  a39319a );
 a39323a <=( A299  and  (not A298) );
 a39326a <=( A302  and  A300 );
 a39327a <=( a39326a  and  a39323a );
 a39328a <=( a39327a  and  a39320a );
 a39332a <=( A199  and  A166 );
 a39333a <=( A167  and  a39332a );
 a39337a <=( (not A202)  and  (not A201) );
 a39338a <=( (not A200)  and  a39337a );
 a39339a <=( a39338a  and  a39333a );
 a39343a <=( A269  and  (not A267) );
 a39344a <=( (not A203)  and  a39343a );
 a39347a <=( (not A299)  and  A298 );
 a39350a <=( A301  and  A300 );
 a39351a <=( a39350a  and  a39347a );
 a39352a <=( a39351a  and  a39344a );
 a39356a <=( A199  and  A166 );
 a39357a <=( A167  and  a39356a );
 a39361a <=( (not A202)  and  (not A201) );
 a39362a <=( (not A200)  and  a39361a );
 a39363a <=( a39362a  and  a39357a );
 a39367a <=( A269  and  (not A267) );
 a39368a <=( (not A203)  and  a39367a );
 a39371a <=( (not A299)  and  A298 );
 a39374a <=( A302  and  A300 );
 a39375a <=( a39374a  and  a39371a );
 a39376a <=( a39375a  and  a39368a );
 a39380a <=( A199  and  A166 );
 a39381a <=( A167  and  a39380a );
 a39385a <=( (not A202)  and  (not A201) );
 a39386a <=( (not A200)  and  a39385a );
 a39387a <=( a39386a  and  a39381a );
 a39391a <=( A269  and  (not A267) );
 a39392a <=( (not A203)  and  a39391a );
 a39395a <=( A299  and  (not A298) );
 a39398a <=( A301  and  A300 );
 a39399a <=( a39398a  and  a39395a );
 a39400a <=( a39399a  and  a39392a );
 a39404a <=( A199  and  A166 );
 a39405a <=( A167  and  a39404a );
 a39409a <=( (not A202)  and  (not A201) );
 a39410a <=( (not A200)  and  a39409a );
 a39411a <=( a39410a  and  a39405a );
 a39415a <=( A269  and  (not A267) );
 a39416a <=( (not A203)  and  a39415a );
 a39419a <=( A299  and  (not A298) );
 a39422a <=( A302  and  A300 );
 a39423a <=( a39422a  and  a39419a );
 a39424a <=( a39423a  and  a39416a );
 a39428a <=( A199  and  A166 );
 a39429a <=( A167  and  a39428a );
 a39433a <=( (not A202)  and  (not A201) );
 a39434a <=( (not A200)  and  a39433a );
 a39435a <=( a39434a  and  a39429a );
 a39439a <=( A266  and  A265 );
 a39440a <=( (not A203)  and  a39439a );
 a39443a <=( (not A299)  and  A298 );
 a39446a <=( A301  and  A300 );
 a39447a <=( a39446a  and  a39443a );
 a39448a <=( a39447a  and  a39440a );
 a39452a <=( A199  and  A166 );
 a39453a <=( A167  and  a39452a );
 a39457a <=( (not A202)  and  (not A201) );
 a39458a <=( (not A200)  and  a39457a );
 a39459a <=( a39458a  and  a39453a );
 a39463a <=( A266  and  A265 );
 a39464a <=( (not A203)  and  a39463a );
 a39467a <=( (not A299)  and  A298 );
 a39470a <=( A302  and  A300 );
 a39471a <=( a39470a  and  a39467a );
 a39472a <=( a39471a  and  a39464a );
 a39476a <=( A199  and  A166 );
 a39477a <=( A167  and  a39476a );
 a39481a <=( (not A202)  and  (not A201) );
 a39482a <=( (not A200)  and  a39481a );
 a39483a <=( a39482a  and  a39477a );
 a39487a <=( A266  and  A265 );
 a39488a <=( (not A203)  and  a39487a );
 a39491a <=( A299  and  (not A298) );
 a39494a <=( A301  and  A300 );
 a39495a <=( a39494a  and  a39491a );
 a39496a <=( a39495a  and  a39488a );
 a39500a <=( A199  and  A166 );
 a39501a <=( A167  and  a39500a );
 a39505a <=( (not A202)  and  (not A201) );
 a39506a <=( (not A200)  and  a39505a );
 a39507a <=( a39506a  and  a39501a );
 a39511a <=( A266  and  A265 );
 a39512a <=( (not A203)  and  a39511a );
 a39515a <=( A299  and  (not A298) );
 a39518a <=( A302  and  A300 );
 a39519a <=( a39518a  and  a39515a );
 a39520a <=( a39519a  and  a39512a );
 a39524a <=( A199  and  A166 );
 a39525a <=( A167  and  a39524a );
 a39529a <=( (not A202)  and  (not A201) );
 a39530a <=( (not A200)  and  a39529a );
 a39531a <=( a39530a  and  a39525a );
 a39535a <=( (not A266)  and  (not A265) );
 a39536a <=( (not A203)  and  a39535a );
 a39539a <=( (not A299)  and  A298 );
 a39542a <=( A301  and  A300 );
 a39543a <=( a39542a  and  a39539a );
 a39544a <=( a39543a  and  a39536a );
 a39548a <=( A199  and  A166 );
 a39549a <=( A167  and  a39548a );
 a39553a <=( (not A202)  and  (not A201) );
 a39554a <=( (not A200)  and  a39553a );
 a39555a <=( a39554a  and  a39549a );
 a39559a <=( (not A266)  and  (not A265) );
 a39560a <=( (not A203)  and  a39559a );
 a39563a <=( (not A299)  and  A298 );
 a39566a <=( A302  and  A300 );
 a39567a <=( a39566a  and  a39563a );
 a39568a <=( a39567a  and  a39560a );
 a39572a <=( A199  and  A166 );
 a39573a <=( A167  and  a39572a );
 a39577a <=( (not A202)  and  (not A201) );
 a39578a <=( (not A200)  and  a39577a );
 a39579a <=( a39578a  and  a39573a );
 a39583a <=( (not A266)  and  (not A265) );
 a39584a <=( (not A203)  and  a39583a );
 a39587a <=( A299  and  (not A298) );
 a39590a <=( A301  and  A300 );
 a39591a <=( a39590a  and  a39587a );
 a39592a <=( a39591a  and  a39584a );
 a39596a <=( A199  and  A166 );
 a39597a <=( A167  and  a39596a );
 a39601a <=( (not A202)  and  (not A201) );
 a39602a <=( (not A200)  and  a39601a );
 a39603a <=( a39602a  and  a39597a );
 a39607a <=( (not A266)  and  (not A265) );
 a39608a <=( (not A203)  and  a39607a );
 a39611a <=( A299  and  (not A298) );
 a39614a <=( A302  and  A300 );
 a39615a <=( a39614a  and  a39611a );
 a39616a <=( a39615a  and  a39608a );
 a39620a <=( A201  and  (not A166) );
 a39621a <=( (not A167)  and  a39620a );
 a39625a <=( (not A265)  and  (not A203) );
 a39626a <=( (not A202)  and  a39625a );
 a39627a <=( a39626a  and  a39621a );
 a39631a <=( (not A268)  and  (not A267) );
 a39632a <=( A266  and  a39631a );
 a39635a <=( A300  and  (not A269) );
 a39638a <=( (not A302)  and  (not A301) );
 a39639a <=( a39638a  and  a39635a );
 a39640a <=( a39639a  and  a39632a );
 a39644a <=( A201  and  (not A166) );
 a39645a <=( (not A167)  and  a39644a );
 a39649a <=( A265  and  (not A203) );
 a39650a <=( (not A202)  and  a39649a );
 a39651a <=( a39650a  and  a39645a );
 a39655a <=( (not A268)  and  (not A267) );
 a39656a <=( (not A266)  and  a39655a );
 a39659a <=( A300  and  (not A269) );
 a39662a <=( (not A302)  and  (not A301) );
 a39663a <=( a39662a  and  a39659a );
 a39664a <=( a39663a  and  a39656a );
 a39668a <=( (not A199)  and  (not A166) );
 a39669a <=( (not A167)  and  a39668a );
 a39673a <=( A202  and  A201 );
 a39674a <=( A200  and  a39673a );
 a39675a <=( a39674a  and  a39669a );
 a39679a <=( (not A269)  and  (not A268) );
 a39680a <=( A267  and  a39679a );
 a39683a <=( (not A299)  and  A298 );
 a39686a <=( A301  and  A300 );
 a39687a <=( a39686a  and  a39683a );
 a39688a <=( a39687a  and  a39680a );
 a39692a <=( (not A199)  and  (not A166) );
 a39693a <=( (not A167)  and  a39692a );
 a39697a <=( A202  and  A201 );
 a39698a <=( A200  and  a39697a );
 a39699a <=( a39698a  and  a39693a );
 a39703a <=( (not A269)  and  (not A268) );
 a39704a <=( A267  and  a39703a );
 a39707a <=( (not A299)  and  A298 );
 a39710a <=( A302  and  A300 );
 a39711a <=( a39710a  and  a39707a );
 a39712a <=( a39711a  and  a39704a );
 a39716a <=( (not A199)  and  (not A166) );
 a39717a <=( (not A167)  and  a39716a );
 a39721a <=( A202  and  A201 );
 a39722a <=( A200  and  a39721a );
 a39723a <=( a39722a  and  a39717a );
 a39727a <=( (not A269)  and  (not A268) );
 a39728a <=( A267  and  a39727a );
 a39731a <=( A299  and  (not A298) );
 a39734a <=( A301  and  A300 );
 a39735a <=( a39734a  and  a39731a );
 a39736a <=( a39735a  and  a39728a );
 a39740a <=( (not A199)  and  (not A166) );
 a39741a <=( (not A167)  and  a39740a );
 a39745a <=( A202  and  A201 );
 a39746a <=( A200  and  a39745a );
 a39747a <=( a39746a  and  a39741a );
 a39751a <=( (not A269)  and  (not A268) );
 a39752a <=( A267  and  a39751a );
 a39755a <=( A299  and  (not A298) );
 a39758a <=( A302  and  A300 );
 a39759a <=( a39758a  and  a39755a );
 a39760a <=( a39759a  and  a39752a );
 a39764a <=( (not A199)  and  (not A166) );
 a39765a <=( (not A167)  and  a39764a );
 a39769a <=( A202  and  A201 );
 a39770a <=( A200  and  a39769a );
 a39771a <=( a39770a  and  a39765a );
 a39775a <=( A298  and  A268 );
 a39776a <=( (not A267)  and  a39775a );
 a39779a <=( (not A300)  and  (not A299) );
 a39782a <=( (not A302)  and  (not A301) );
 a39783a <=( a39782a  and  a39779a );
 a39784a <=( a39783a  and  a39776a );
 a39788a <=( (not A199)  and  (not A166) );
 a39789a <=( (not A167)  and  a39788a );
 a39793a <=( A202  and  A201 );
 a39794a <=( A200  and  a39793a );
 a39795a <=( a39794a  and  a39789a );
 a39799a <=( (not A298)  and  A268 );
 a39800a <=( (not A267)  and  a39799a );
 a39803a <=( (not A300)  and  A299 );
 a39806a <=( (not A302)  and  (not A301) );
 a39807a <=( a39806a  and  a39803a );
 a39808a <=( a39807a  and  a39800a );
 a39812a <=( (not A199)  and  (not A166) );
 a39813a <=( (not A167)  and  a39812a );
 a39817a <=( A202  and  A201 );
 a39818a <=( A200  and  a39817a );
 a39819a <=( a39818a  and  a39813a );
 a39823a <=( A298  and  A269 );
 a39824a <=( (not A267)  and  a39823a );
 a39827a <=( (not A300)  and  (not A299) );
 a39830a <=( (not A302)  and  (not A301) );
 a39831a <=( a39830a  and  a39827a );
 a39832a <=( a39831a  and  a39824a );
 a39836a <=( (not A199)  and  (not A166) );
 a39837a <=( (not A167)  and  a39836a );
 a39841a <=( A202  and  A201 );
 a39842a <=( A200  and  a39841a );
 a39843a <=( a39842a  and  a39837a );
 a39847a <=( (not A298)  and  A269 );
 a39848a <=( (not A267)  and  a39847a );
 a39851a <=( (not A300)  and  A299 );
 a39854a <=( (not A302)  and  (not A301) );
 a39855a <=( a39854a  and  a39851a );
 a39856a <=( a39855a  and  a39848a );
 a39860a <=( (not A199)  and  (not A166) );
 a39861a <=( (not A167)  and  a39860a );
 a39865a <=( A202  and  A201 );
 a39866a <=( A200  and  a39865a );
 a39867a <=( a39866a  and  a39861a );
 a39871a <=( A298  and  A266 );
 a39872a <=( A265  and  a39871a );
 a39875a <=( (not A300)  and  (not A299) );
 a39878a <=( (not A302)  and  (not A301) );
 a39879a <=( a39878a  and  a39875a );
 a39880a <=( a39879a  and  a39872a );
 a39884a <=( (not A199)  and  (not A166) );
 a39885a <=( (not A167)  and  a39884a );
 a39889a <=( A202  and  A201 );
 a39890a <=( A200  and  a39889a );
 a39891a <=( a39890a  and  a39885a );
 a39895a <=( (not A298)  and  A266 );
 a39896a <=( A265  and  a39895a );
 a39899a <=( (not A300)  and  A299 );
 a39902a <=( (not A302)  and  (not A301) );
 a39903a <=( a39902a  and  a39899a );
 a39904a <=( a39903a  and  a39896a );
 a39908a <=( (not A199)  and  (not A166) );
 a39909a <=( (not A167)  and  a39908a );
 a39913a <=( A202  and  A201 );
 a39914a <=( A200  and  a39913a );
 a39915a <=( a39914a  and  a39909a );
 a39919a <=( A298  and  (not A266) );
 a39920a <=( (not A265)  and  a39919a );
 a39923a <=( (not A300)  and  (not A299) );
 a39926a <=( (not A302)  and  (not A301) );
 a39927a <=( a39926a  and  a39923a );
 a39928a <=( a39927a  and  a39920a );
 a39932a <=( (not A199)  and  (not A166) );
 a39933a <=( (not A167)  and  a39932a );
 a39937a <=( A202  and  A201 );
 a39938a <=( A200  and  a39937a );
 a39939a <=( a39938a  and  a39933a );
 a39943a <=( (not A298)  and  (not A266) );
 a39944a <=( (not A265)  and  a39943a );
 a39947a <=( (not A300)  and  A299 );
 a39950a <=( (not A302)  and  (not A301) );
 a39951a <=( a39950a  and  a39947a );
 a39952a <=( a39951a  and  a39944a );
 a39956a <=( (not A199)  and  (not A166) );
 a39957a <=( (not A167)  and  a39956a );
 a39961a <=( A203  and  A201 );
 a39962a <=( A200  and  a39961a );
 a39963a <=( a39962a  and  a39957a );
 a39967a <=( (not A269)  and  (not A268) );
 a39968a <=( A267  and  a39967a );
 a39971a <=( (not A299)  and  A298 );
 a39974a <=( A301  and  A300 );
 a39975a <=( a39974a  and  a39971a );
 a39976a <=( a39975a  and  a39968a );
 a39980a <=( (not A199)  and  (not A166) );
 a39981a <=( (not A167)  and  a39980a );
 a39985a <=( A203  and  A201 );
 a39986a <=( A200  and  a39985a );
 a39987a <=( a39986a  and  a39981a );
 a39991a <=( (not A269)  and  (not A268) );
 a39992a <=( A267  and  a39991a );
 a39995a <=( (not A299)  and  A298 );
 a39998a <=( A302  and  A300 );
 a39999a <=( a39998a  and  a39995a );
 a40000a <=( a39999a  and  a39992a );
 a40004a <=( (not A199)  and  (not A166) );
 a40005a <=( (not A167)  and  a40004a );
 a40009a <=( A203  and  A201 );
 a40010a <=( A200  and  a40009a );
 a40011a <=( a40010a  and  a40005a );
 a40015a <=( (not A269)  and  (not A268) );
 a40016a <=( A267  and  a40015a );
 a40019a <=( A299  and  (not A298) );
 a40022a <=( A301  and  A300 );
 a40023a <=( a40022a  and  a40019a );
 a40024a <=( a40023a  and  a40016a );
 a40028a <=( (not A199)  and  (not A166) );
 a40029a <=( (not A167)  and  a40028a );
 a40033a <=( A203  and  A201 );
 a40034a <=( A200  and  a40033a );
 a40035a <=( a40034a  and  a40029a );
 a40039a <=( (not A269)  and  (not A268) );
 a40040a <=( A267  and  a40039a );
 a40043a <=( A299  and  (not A298) );
 a40046a <=( A302  and  A300 );
 a40047a <=( a40046a  and  a40043a );
 a40048a <=( a40047a  and  a40040a );
 a40052a <=( (not A199)  and  (not A166) );
 a40053a <=( (not A167)  and  a40052a );
 a40057a <=( A203  and  A201 );
 a40058a <=( A200  and  a40057a );
 a40059a <=( a40058a  and  a40053a );
 a40063a <=( A298  and  A268 );
 a40064a <=( (not A267)  and  a40063a );
 a40067a <=( (not A300)  and  (not A299) );
 a40070a <=( (not A302)  and  (not A301) );
 a40071a <=( a40070a  and  a40067a );
 a40072a <=( a40071a  and  a40064a );
 a40076a <=( (not A199)  and  (not A166) );
 a40077a <=( (not A167)  and  a40076a );
 a40081a <=( A203  and  A201 );
 a40082a <=( A200  and  a40081a );
 a40083a <=( a40082a  and  a40077a );
 a40087a <=( (not A298)  and  A268 );
 a40088a <=( (not A267)  and  a40087a );
 a40091a <=( (not A300)  and  A299 );
 a40094a <=( (not A302)  and  (not A301) );
 a40095a <=( a40094a  and  a40091a );
 a40096a <=( a40095a  and  a40088a );
 a40100a <=( (not A199)  and  (not A166) );
 a40101a <=( (not A167)  and  a40100a );
 a40105a <=( A203  and  A201 );
 a40106a <=( A200  and  a40105a );
 a40107a <=( a40106a  and  a40101a );
 a40111a <=( A298  and  A269 );
 a40112a <=( (not A267)  and  a40111a );
 a40115a <=( (not A300)  and  (not A299) );
 a40118a <=( (not A302)  and  (not A301) );
 a40119a <=( a40118a  and  a40115a );
 a40120a <=( a40119a  and  a40112a );
 a40124a <=( (not A199)  and  (not A166) );
 a40125a <=( (not A167)  and  a40124a );
 a40129a <=( A203  and  A201 );
 a40130a <=( A200  and  a40129a );
 a40131a <=( a40130a  and  a40125a );
 a40135a <=( (not A298)  and  A269 );
 a40136a <=( (not A267)  and  a40135a );
 a40139a <=( (not A300)  and  A299 );
 a40142a <=( (not A302)  and  (not A301) );
 a40143a <=( a40142a  and  a40139a );
 a40144a <=( a40143a  and  a40136a );
 a40148a <=( (not A199)  and  (not A166) );
 a40149a <=( (not A167)  and  a40148a );
 a40153a <=( A203  and  A201 );
 a40154a <=( A200  and  a40153a );
 a40155a <=( a40154a  and  a40149a );
 a40159a <=( A298  and  A266 );
 a40160a <=( A265  and  a40159a );
 a40163a <=( (not A300)  and  (not A299) );
 a40166a <=( (not A302)  and  (not A301) );
 a40167a <=( a40166a  and  a40163a );
 a40168a <=( a40167a  and  a40160a );
 a40172a <=( (not A199)  and  (not A166) );
 a40173a <=( (not A167)  and  a40172a );
 a40177a <=( A203  and  A201 );
 a40178a <=( A200  and  a40177a );
 a40179a <=( a40178a  and  a40173a );
 a40183a <=( (not A298)  and  A266 );
 a40184a <=( A265  and  a40183a );
 a40187a <=( (not A300)  and  A299 );
 a40190a <=( (not A302)  and  (not A301) );
 a40191a <=( a40190a  and  a40187a );
 a40192a <=( a40191a  and  a40184a );
 a40196a <=( (not A199)  and  (not A166) );
 a40197a <=( (not A167)  and  a40196a );
 a40201a <=( A203  and  A201 );
 a40202a <=( A200  and  a40201a );
 a40203a <=( a40202a  and  a40197a );
 a40207a <=( A298  and  (not A266) );
 a40208a <=( (not A265)  and  a40207a );
 a40211a <=( (not A300)  and  (not A299) );
 a40214a <=( (not A302)  and  (not A301) );
 a40215a <=( a40214a  and  a40211a );
 a40216a <=( a40215a  and  a40208a );
 a40220a <=( (not A199)  and  (not A166) );
 a40221a <=( (not A167)  and  a40220a );
 a40225a <=( A203  and  A201 );
 a40226a <=( A200  and  a40225a );
 a40227a <=( a40226a  and  a40221a );
 a40231a <=( (not A298)  and  (not A266) );
 a40232a <=( (not A265)  and  a40231a );
 a40235a <=( (not A300)  and  A299 );
 a40238a <=( (not A302)  and  (not A301) );
 a40239a <=( a40238a  and  a40235a );
 a40240a <=( a40239a  and  a40232a );
 a40244a <=( (not A199)  and  (not A166) );
 a40245a <=( (not A167)  and  a40244a );
 a40249a <=( (not A202)  and  (not A201) );
 a40250a <=( A200  and  a40249a );
 a40251a <=( a40250a  and  a40245a );
 a40255a <=( A268  and  (not A267) );
 a40256a <=( (not A203)  and  a40255a );
 a40259a <=( (not A299)  and  A298 );
 a40262a <=( A301  and  A300 );
 a40263a <=( a40262a  and  a40259a );
 a40264a <=( a40263a  and  a40256a );
 a40268a <=( (not A199)  and  (not A166) );
 a40269a <=( (not A167)  and  a40268a );
 a40273a <=( (not A202)  and  (not A201) );
 a40274a <=( A200  and  a40273a );
 a40275a <=( a40274a  and  a40269a );
 a40279a <=( A268  and  (not A267) );
 a40280a <=( (not A203)  and  a40279a );
 a40283a <=( (not A299)  and  A298 );
 a40286a <=( A302  and  A300 );
 a40287a <=( a40286a  and  a40283a );
 a40288a <=( a40287a  and  a40280a );
 a40292a <=( (not A199)  and  (not A166) );
 a40293a <=( (not A167)  and  a40292a );
 a40297a <=( (not A202)  and  (not A201) );
 a40298a <=( A200  and  a40297a );
 a40299a <=( a40298a  and  a40293a );
 a40303a <=( A268  and  (not A267) );
 a40304a <=( (not A203)  and  a40303a );
 a40307a <=( A299  and  (not A298) );
 a40310a <=( A301  and  A300 );
 a40311a <=( a40310a  and  a40307a );
 a40312a <=( a40311a  and  a40304a );
 a40316a <=( (not A199)  and  (not A166) );
 a40317a <=( (not A167)  and  a40316a );
 a40321a <=( (not A202)  and  (not A201) );
 a40322a <=( A200  and  a40321a );
 a40323a <=( a40322a  and  a40317a );
 a40327a <=( A268  and  (not A267) );
 a40328a <=( (not A203)  and  a40327a );
 a40331a <=( A299  and  (not A298) );
 a40334a <=( A302  and  A300 );
 a40335a <=( a40334a  and  a40331a );
 a40336a <=( a40335a  and  a40328a );
 a40340a <=( (not A199)  and  (not A166) );
 a40341a <=( (not A167)  and  a40340a );
 a40345a <=( (not A202)  and  (not A201) );
 a40346a <=( A200  and  a40345a );
 a40347a <=( a40346a  and  a40341a );
 a40351a <=( A269  and  (not A267) );
 a40352a <=( (not A203)  and  a40351a );
 a40355a <=( (not A299)  and  A298 );
 a40358a <=( A301  and  A300 );
 a40359a <=( a40358a  and  a40355a );
 a40360a <=( a40359a  and  a40352a );
 a40364a <=( (not A199)  and  (not A166) );
 a40365a <=( (not A167)  and  a40364a );
 a40369a <=( (not A202)  and  (not A201) );
 a40370a <=( A200  and  a40369a );
 a40371a <=( a40370a  and  a40365a );
 a40375a <=( A269  and  (not A267) );
 a40376a <=( (not A203)  and  a40375a );
 a40379a <=( (not A299)  and  A298 );
 a40382a <=( A302  and  A300 );
 a40383a <=( a40382a  and  a40379a );
 a40384a <=( a40383a  and  a40376a );
 a40388a <=( (not A199)  and  (not A166) );
 a40389a <=( (not A167)  and  a40388a );
 a40393a <=( (not A202)  and  (not A201) );
 a40394a <=( A200  and  a40393a );
 a40395a <=( a40394a  and  a40389a );
 a40399a <=( A269  and  (not A267) );
 a40400a <=( (not A203)  and  a40399a );
 a40403a <=( A299  and  (not A298) );
 a40406a <=( A301  and  A300 );
 a40407a <=( a40406a  and  a40403a );
 a40408a <=( a40407a  and  a40400a );
 a40412a <=( (not A199)  and  (not A166) );
 a40413a <=( (not A167)  and  a40412a );
 a40417a <=( (not A202)  and  (not A201) );
 a40418a <=( A200  and  a40417a );
 a40419a <=( a40418a  and  a40413a );
 a40423a <=( A269  and  (not A267) );
 a40424a <=( (not A203)  and  a40423a );
 a40427a <=( A299  and  (not A298) );
 a40430a <=( A302  and  A300 );
 a40431a <=( a40430a  and  a40427a );
 a40432a <=( a40431a  and  a40424a );
 a40436a <=( (not A199)  and  (not A166) );
 a40437a <=( (not A167)  and  a40436a );
 a40441a <=( (not A202)  and  (not A201) );
 a40442a <=( A200  and  a40441a );
 a40443a <=( a40442a  and  a40437a );
 a40447a <=( A266  and  A265 );
 a40448a <=( (not A203)  and  a40447a );
 a40451a <=( (not A299)  and  A298 );
 a40454a <=( A301  and  A300 );
 a40455a <=( a40454a  and  a40451a );
 a40456a <=( a40455a  and  a40448a );
 a40460a <=( (not A199)  and  (not A166) );
 a40461a <=( (not A167)  and  a40460a );
 a40465a <=( (not A202)  and  (not A201) );
 a40466a <=( A200  and  a40465a );
 a40467a <=( a40466a  and  a40461a );
 a40471a <=( A266  and  A265 );
 a40472a <=( (not A203)  and  a40471a );
 a40475a <=( (not A299)  and  A298 );
 a40478a <=( A302  and  A300 );
 a40479a <=( a40478a  and  a40475a );
 a40480a <=( a40479a  and  a40472a );
 a40484a <=( (not A199)  and  (not A166) );
 a40485a <=( (not A167)  and  a40484a );
 a40489a <=( (not A202)  and  (not A201) );
 a40490a <=( A200  and  a40489a );
 a40491a <=( a40490a  and  a40485a );
 a40495a <=( A266  and  A265 );
 a40496a <=( (not A203)  and  a40495a );
 a40499a <=( A299  and  (not A298) );
 a40502a <=( A301  and  A300 );
 a40503a <=( a40502a  and  a40499a );
 a40504a <=( a40503a  and  a40496a );
 a40508a <=( (not A199)  and  (not A166) );
 a40509a <=( (not A167)  and  a40508a );
 a40513a <=( (not A202)  and  (not A201) );
 a40514a <=( A200  and  a40513a );
 a40515a <=( a40514a  and  a40509a );
 a40519a <=( A266  and  A265 );
 a40520a <=( (not A203)  and  a40519a );
 a40523a <=( A299  and  (not A298) );
 a40526a <=( A302  and  A300 );
 a40527a <=( a40526a  and  a40523a );
 a40528a <=( a40527a  and  a40520a );
 a40532a <=( (not A199)  and  (not A166) );
 a40533a <=( (not A167)  and  a40532a );
 a40537a <=( (not A202)  and  (not A201) );
 a40538a <=( A200  and  a40537a );
 a40539a <=( a40538a  and  a40533a );
 a40543a <=( (not A266)  and  (not A265) );
 a40544a <=( (not A203)  and  a40543a );
 a40547a <=( (not A299)  and  A298 );
 a40550a <=( A301  and  A300 );
 a40551a <=( a40550a  and  a40547a );
 a40552a <=( a40551a  and  a40544a );
 a40556a <=( (not A199)  and  (not A166) );
 a40557a <=( (not A167)  and  a40556a );
 a40561a <=( (not A202)  and  (not A201) );
 a40562a <=( A200  and  a40561a );
 a40563a <=( a40562a  and  a40557a );
 a40567a <=( (not A266)  and  (not A265) );
 a40568a <=( (not A203)  and  a40567a );
 a40571a <=( (not A299)  and  A298 );
 a40574a <=( A302  and  A300 );
 a40575a <=( a40574a  and  a40571a );
 a40576a <=( a40575a  and  a40568a );
 a40580a <=( (not A199)  and  (not A166) );
 a40581a <=( (not A167)  and  a40580a );
 a40585a <=( (not A202)  and  (not A201) );
 a40586a <=( A200  and  a40585a );
 a40587a <=( a40586a  and  a40581a );
 a40591a <=( (not A266)  and  (not A265) );
 a40592a <=( (not A203)  and  a40591a );
 a40595a <=( A299  and  (not A298) );
 a40598a <=( A301  and  A300 );
 a40599a <=( a40598a  and  a40595a );
 a40600a <=( a40599a  and  a40592a );
 a40604a <=( (not A199)  and  (not A166) );
 a40605a <=( (not A167)  and  a40604a );
 a40609a <=( (not A202)  and  (not A201) );
 a40610a <=( A200  and  a40609a );
 a40611a <=( a40610a  and  a40605a );
 a40615a <=( (not A266)  and  (not A265) );
 a40616a <=( (not A203)  and  a40615a );
 a40619a <=( A299  and  (not A298) );
 a40622a <=( A302  and  A300 );
 a40623a <=( a40622a  and  a40619a );
 a40624a <=( a40623a  and  a40616a );
 a40628a <=( A199  and  (not A166) );
 a40629a <=( (not A167)  and  a40628a );
 a40633a <=( A202  and  A201 );
 a40634a <=( (not A200)  and  a40633a );
 a40635a <=( a40634a  and  a40629a );
 a40639a <=( (not A269)  and  (not A268) );
 a40640a <=( A267  and  a40639a );
 a40643a <=( (not A299)  and  A298 );
 a40646a <=( A301  and  A300 );
 a40647a <=( a40646a  and  a40643a );
 a40648a <=( a40647a  and  a40640a );
 a40652a <=( A199  and  (not A166) );
 a40653a <=( (not A167)  and  a40652a );
 a40657a <=( A202  and  A201 );
 a40658a <=( (not A200)  and  a40657a );
 a40659a <=( a40658a  and  a40653a );
 a40663a <=( (not A269)  and  (not A268) );
 a40664a <=( A267  and  a40663a );
 a40667a <=( (not A299)  and  A298 );
 a40670a <=( A302  and  A300 );
 a40671a <=( a40670a  and  a40667a );
 a40672a <=( a40671a  and  a40664a );
 a40676a <=( A199  and  (not A166) );
 a40677a <=( (not A167)  and  a40676a );
 a40681a <=( A202  and  A201 );
 a40682a <=( (not A200)  and  a40681a );
 a40683a <=( a40682a  and  a40677a );
 a40687a <=( (not A269)  and  (not A268) );
 a40688a <=( A267  and  a40687a );
 a40691a <=( A299  and  (not A298) );
 a40694a <=( A301  and  A300 );
 a40695a <=( a40694a  and  a40691a );
 a40696a <=( a40695a  and  a40688a );
 a40700a <=( A199  and  (not A166) );
 a40701a <=( (not A167)  and  a40700a );
 a40705a <=( A202  and  A201 );
 a40706a <=( (not A200)  and  a40705a );
 a40707a <=( a40706a  and  a40701a );
 a40711a <=( (not A269)  and  (not A268) );
 a40712a <=( A267  and  a40711a );
 a40715a <=( A299  and  (not A298) );
 a40718a <=( A302  and  A300 );
 a40719a <=( a40718a  and  a40715a );
 a40720a <=( a40719a  and  a40712a );
 a40724a <=( A199  and  (not A166) );
 a40725a <=( (not A167)  and  a40724a );
 a40729a <=( A202  and  A201 );
 a40730a <=( (not A200)  and  a40729a );
 a40731a <=( a40730a  and  a40725a );
 a40735a <=( A298  and  A268 );
 a40736a <=( (not A267)  and  a40735a );
 a40739a <=( (not A300)  and  (not A299) );
 a40742a <=( (not A302)  and  (not A301) );
 a40743a <=( a40742a  and  a40739a );
 a40744a <=( a40743a  and  a40736a );
 a40748a <=( A199  and  (not A166) );
 a40749a <=( (not A167)  and  a40748a );
 a40753a <=( A202  and  A201 );
 a40754a <=( (not A200)  and  a40753a );
 a40755a <=( a40754a  and  a40749a );
 a40759a <=( (not A298)  and  A268 );
 a40760a <=( (not A267)  and  a40759a );
 a40763a <=( (not A300)  and  A299 );
 a40766a <=( (not A302)  and  (not A301) );
 a40767a <=( a40766a  and  a40763a );
 a40768a <=( a40767a  and  a40760a );
 a40772a <=( A199  and  (not A166) );
 a40773a <=( (not A167)  and  a40772a );
 a40777a <=( A202  and  A201 );
 a40778a <=( (not A200)  and  a40777a );
 a40779a <=( a40778a  and  a40773a );
 a40783a <=( A298  and  A269 );
 a40784a <=( (not A267)  and  a40783a );
 a40787a <=( (not A300)  and  (not A299) );
 a40790a <=( (not A302)  and  (not A301) );
 a40791a <=( a40790a  and  a40787a );
 a40792a <=( a40791a  and  a40784a );
 a40796a <=( A199  and  (not A166) );
 a40797a <=( (not A167)  and  a40796a );
 a40801a <=( A202  and  A201 );
 a40802a <=( (not A200)  and  a40801a );
 a40803a <=( a40802a  and  a40797a );
 a40807a <=( (not A298)  and  A269 );
 a40808a <=( (not A267)  and  a40807a );
 a40811a <=( (not A300)  and  A299 );
 a40814a <=( (not A302)  and  (not A301) );
 a40815a <=( a40814a  and  a40811a );
 a40816a <=( a40815a  and  a40808a );
 a40820a <=( A199  and  (not A166) );
 a40821a <=( (not A167)  and  a40820a );
 a40825a <=( A202  and  A201 );
 a40826a <=( (not A200)  and  a40825a );
 a40827a <=( a40826a  and  a40821a );
 a40831a <=( A298  and  A266 );
 a40832a <=( A265  and  a40831a );
 a40835a <=( (not A300)  and  (not A299) );
 a40838a <=( (not A302)  and  (not A301) );
 a40839a <=( a40838a  and  a40835a );
 a40840a <=( a40839a  and  a40832a );
 a40844a <=( A199  and  (not A166) );
 a40845a <=( (not A167)  and  a40844a );
 a40849a <=( A202  and  A201 );
 a40850a <=( (not A200)  and  a40849a );
 a40851a <=( a40850a  and  a40845a );
 a40855a <=( (not A298)  and  A266 );
 a40856a <=( A265  and  a40855a );
 a40859a <=( (not A300)  and  A299 );
 a40862a <=( (not A302)  and  (not A301) );
 a40863a <=( a40862a  and  a40859a );
 a40864a <=( a40863a  and  a40856a );
 a40868a <=( A199  and  (not A166) );
 a40869a <=( (not A167)  and  a40868a );
 a40873a <=( A202  and  A201 );
 a40874a <=( (not A200)  and  a40873a );
 a40875a <=( a40874a  and  a40869a );
 a40879a <=( A298  and  (not A266) );
 a40880a <=( (not A265)  and  a40879a );
 a40883a <=( (not A300)  and  (not A299) );
 a40886a <=( (not A302)  and  (not A301) );
 a40887a <=( a40886a  and  a40883a );
 a40888a <=( a40887a  and  a40880a );
 a40892a <=( A199  and  (not A166) );
 a40893a <=( (not A167)  and  a40892a );
 a40897a <=( A202  and  A201 );
 a40898a <=( (not A200)  and  a40897a );
 a40899a <=( a40898a  and  a40893a );
 a40903a <=( (not A298)  and  (not A266) );
 a40904a <=( (not A265)  and  a40903a );
 a40907a <=( (not A300)  and  A299 );
 a40910a <=( (not A302)  and  (not A301) );
 a40911a <=( a40910a  and  a40907a );
 a40912a <=( a40911a  and  a40904a );
 a40916a <=( A199  and  (not A166) );
 a40917a <=( (not A167)  and  a40916a );
 a40921a <=( A203  and  A201 );
 a40922a <=( (not A200)  and  a40921a );
 a40923a <=( a40922a  and  a40917a );
 a40927a <=( (not A269)  and  (not A268) );
 a40928a <=( A267  and  a40927a );
 a40931a <=( (not A299)  and  A298 );
 a40934a <=( A301  and  A300 );
 a40935a <=( a40934a  and  a40931a );
 a40936a <=( a40935a  and  a40928a );
 a40940a <=( A199  and  (not A166) );
 a40941a <=( (not A167)  and  a40940a );
 a40945a <=( A203  and  A201 );
 a40946a <=( (not A200)  and  a40945a );
 a40947a <=( a40946a  and  a40941a );
 a40951a <=( (not A269)  and  (not A268) );
 a40952a <=( A267  and  a40951a );
 a40955a <=( (not A299)  and  A298 );
 a40958a <=( A302  and  A300 );
 a40959a <=( a40958a  and  a40955a );
 a40960a <=( a40959a  and  a40952a );
 a40964a <=( A199  and  (not A166) );
 a40965a <=( (not A167)  and  a40964a );
 a40969a <=( A203  and  A201 );
 a40970a <=( (not A200)  and  a40969a );
 a40971a <=( a40970a  and  a40965a );
 a40975a <=( (not A269)  and  (not A268) );
 a40976a <=( A267  and  a40975a );
 a40979a <=( A299  and  (not A298) );
 a40982a <=( A301  and  A300 );
 a40983a <=( a40982a  and  a40979a );
 a40984a <=( a40983a  and  a40976a );
 a40988a <=( A199  and  (not A166) );
 a40989a <=( (not A167)  and  a40988a );
 a40993a <=( A203  and  A201 );
 a40994a <=( (not A200)  and  a40993a );
 a40995a <=( a40994a  and  a40989a );
 a40999a <=( (not A269)  and  (not A268) );
 a41000a <=( A267  and  a40999a );
 a41003a <=( A299  and  (not A298) );
 a41006a <=( A302  and  A300 );
 a41007a <=( a41006a  and  a41003a );
 a41008a <=( a41007a  and  a41000a );
 a41012a <=( A199  and  (not A166) );
 a41013a <=( (not A167)  and  a41012a );
 a41017a <=( A203  and  A201 );
 a41018a <=( (not A200)  and  a41017a );
 a41019a <=( a41018a  and  a41013a );
 a41023a <=( A298  and  A268 );
 a41024a <=( (not A267)  and  a41023a );
 a41027a <=( (not A300)  and  (not A299) );
 a41030a <=( (not A302)  and  (not A301) );
 a41031a <=( a41030a  and  a41027a );
 a41032a <=( a41031a  and  a41024a );
 a41036a <=( A199  and  (not A166) );
 a41037a <=( (not A167)  and  a41036a );
 a41041a <=( A203  and  A201 );
 a41042a <=( (not A200)  and  a41041a );
 a41043a <=( a41042a  and  a41037a );
 a41047a <=( (not A298)  and  A268 );
 a41048a <=( (not A267)  and  a41047a );
 a41051a <=( (not A300)  and  A299 );
 a41054a <=( (not A302)  and  (not A301) );
 a41055a <=( a41054a  and  a41051a );
 a41056a <=( a41055a  and  a41048a );
 a41060a <=( A199  and  (not A166) );
 a41061a <=( (not A167)  and  a41060a );
 a41065a <=( A203  and  A201 );
 a41066a <=( (not A200)  and  a41065a );
 a41067a <=( a41066a  and  a41061a );
 a41071a <=( A298  and  A269 );
 a41072a <=( (not A267)  and  a41071a );
 a41075a <=( (not A300)  and  (not A299) );
 a41078a <=( (not A302)  and  (not A301) );
 a41079a <=( a41078a  and  a41075a );
 a41080a <=( a41079a  and  a41072a );
 a41084a <=( A199  and  (not A166) );
 a41085a <=( (not A167)  and  a41084a );
 a41089a <=( A203  and  A201 );
 a41090a <=( (not A200)  and  a41089a );
 a41091a <=( a41090a  and  a41085a );
 a41095a <=( (not A298)  and  A269 );
 a41096a <=( (not A267)  and  a41095a );
 a41099a <=( (not A300)  and  A299 );
 a41102a <=( (not A302)  and  (not A301) );
 a41103a <=( a41102a  and  a41099a );
 a41104a <=( a41103a  and  a41096a );
 a41108a <=( A199  and  (not A166) );
 a41109a <=( (not A167)  and  a41108a );
 a41113a <=( A203  and  A201 );
 a41114a <=( (not A200)  and  a41113a );
 a41115a <=( a41114a  and  a41109a );
 a41119a <=( A298  and  A266 );
 a41120a <=( A265  and  a41119a );
 a41123a <=( (not A300)  and  (not A299) );
 a41126a <=( (not A302)  and  (not A301) );
 a41127a <=( a41126a  and  a41123a );
 a41128a <=( a41127a  and  a41120a );
 a41132a <=( A199  and  (not A166) );
 a41133a <=( (not A167)  and  a41132a );
 a41137a <=( A203  and  A201 );
 a41138a <=( (not A200)  and  a41137a );
 a41139a <=( a41138a  and  a41133a );
 a41143a <=( (not A298)  and  A266 );
 a41144a <=( A265  and  a41143a );
 a41147a <=( (not A300)  and  A299 );
 a41150a <=( (not A302)  and  (not A301) );
 a41151a <=( a41150a  and  a41147a );
 a41152a <=( a41151a  and  a41144a );
 a41156a <=( A199  and  (not A166) );
 a41157a <=( (not A167)  and  a41156a );
 a41161a <=( A203  and  A201 );
 a41162a <=( (not A200)  and  a41161a );
 a41163a <=( a41162a  and  a41157a );
 a41167a <=( A298  and  (not A266) );
 a41168a <=( (not A265)  and  a41167a );
 a41171a <=( (not A300)  and  (not A299) );
 a41174a <=( (not A302)  and  (not A301) );
 a41175a <=( a41174a  and  a41171a );
 a41176a <=( a41175a  and  a41168a );
 a41180a <=( A199  and  (not A166) );
 a41181a <=( (not A167)  and  a41180a );
 a41185a <=( A203  and  A201 );
 a41186a <=( (not A200)  and  a41185a );
 a41187a <=( a41186a  and  a41181a );
 a41191a <=( (not A298)  and  (not A266) );
 a41192a <=( (not A265)  and  a41191a );
 a41195a <=( (not A300)  and  A299 );
 a41198a <=( (not A302)  and  (not A301) );
 a41199a <=( a41198a  and  a41195a );
 a41200a <=( a41199a  and  a41192a );
 a41204a <=( A199  and  (not A166) );
 a41205a <=( (not A167)  and  a41204a );
 a41209a <=( (not A202)  and  (not A201) );
 a41210a <=( (not A200)  and  a41209a );
 a41211a <=( a41210a  and  a41205a );
 a41215a <=( A268  and  (not A267) );
 a41216a <=( (not A203)  and  a41215a );
 a41219a <=( (not A299)  and  A298 );
 a41222a <=( A301  and  A300 );
 a41223a <=( a41222a  and  a41219a );
 a41224a <=( a41223a  and  a41216a );
 a41228a <=( A199  and  (not A166) );
 a41229a <=( (not A167)  and  a41228a );
 a41233a <=( (not A202)  and  (not A201) );
 a41234a <=( (not A200)  and  a41233a );
 a41235a <=( a41234a  and  a41229a );
 a41239a <=( A268  and  (not A267) );
 a41240a <=( (not A203)  and  a41239a );
 a41243a <=( (not A299)  and  A298 );
 a41246a <=( A302  and  A300 );
 a41247a <=( a41246a  and  a41243a );
 a41248a <=( a41247a  and  a41240a );
 a41252a <=( A199  and  (not A166) );
 a41253a <=( (not A167)  and  a41252a );
 a41257a <=( (not A202)  and  (not A201) );
 a41258a <=( (not A200)  and  a41257a );
 a41259a <=( a41258a  and  a41253a );
 a41263a <=( A268  and  (not A267) );
 a41264a <=( (not A203)  and  a41263a );
 a41267a <=( A299  and  (not A298) );
 a41270a <=( A301  and  A300 );
 a41271a <=( a41270a  and  a41267a );
 a41272a <=( a41271a  and  a41264a );
 a41276a <=( A199  and  (not A166) );
 a41277a <=( (not A167)  and  a41276a );
 a41281a <=( (not A202)  and  (not A201) );
 a41282a <=( (not A200)  and  a41281a );
 a41283a <=( a41282a  and  a41277a );
 a41287a <=( A268  and  (not A267) );
 a41288a <=( (not A203)  and  a41287a );
 a41291a <=( A299  and  (not A298) );
 a41294a <=( A302  and  A300 );
 a41295a <=( a41294a  and  a41291a );
 a41296a <=( a41295a  and  a41288a );
 a41300a <=( A199  and  (not A166) );
 a41301a <=( (not A167)  and  a41300a );
 a41305a <=( (not A202)  and  (not A201) );
 a41306a <=( (not A200)  and  a41305a );
 a41307a <=( a41306a  and  a41301a );
 a41311a <=( A269  and  (not A267) );
 a41312a <=( (not A203)  and  a41311a );
 a41315a <=( (not A299)  and  A298 );
 a41318a <=( A301  and  A300 );
 a41319a <=( a41318a  and  a41315a );
 a41320a <=( a41319a  and  a41312a );
 a41324a <=( A199  and  (not A166) );
 a41325a <=( (not A167)  and  a41324a );
 a41329a <=( (not A202)  and  (not A201) );
 a41330a <=( (not A200)  and  a41329a );
 a41331a <=( a41330a  and  a41325a );
 a41335a <=( A269  and  (not A267) );
 a41336a <=( (not A203)  and  a41335a );
 a41339a <=( (not A299)  and  A298 );
 a41342a <=( A302  and  A300 );
 a41343a <=( a41342a  and  a41339a );
 a41344a <=( a41343a  and  a41336a );
 a41348a <=( A199  and  (not A166) );
 a41349a <=( (not A167)  and  a41348a );
 a41353a <=( (not A202)  and  (not A201) );
 a41354a <=( (not A200)  and  a41353a );
 a41355a <=( a41354a  and  a41349a );
 a41359a <=( A269  and  (not A267) );
 a41360a <=( (not A203)  and  a41359a );
 a41363a <=( A299  and  (not A298) );
 a41366a <=( A301  and  A300 );
 a41367a <=( a41366a  and  a41363a );
 a41368a <=( a41367a  and  a41360a );
 a41372a <=( A199  and  (not A166) );
 a41373a <=( (not A167)  and  a41372a );
 a41377a <=( (not A202)  and  (not A201) );
 a41378a <=( (not A200)  and  a41377a );
 a41379a <=( a41378a  and  a41373a );
 a41383a <=( A269  and  (not A267) );
 a41384a <=( (not A203)  and  a41383a );
 a41387a <=( A299  and  (not A298) );
 a41390a <=( A302  and  A300 );
 a41391a <=( a41390a  and  a41387a );
 a41392a <=( a41391a  and  a41384a );
 a41396a <=( A199  and  (not A166) );
 a41397a <=( (not A167)  and  a41396a );
 a41401a <=( (not A202)  and  (not A201) );
 a41402a <=( (not A200)  and  a41401a );
 a41403a <=( a41402a  and  a41397a );
 a41407a <=( A266  and  A265 );
 a41408a <=( (not A203)  and  a41407a );
 a41411a <=( (not A299)  and  A298 );
 a41414a <=( A301  and  A300 );
 a41415a <=( a41414a  and  a41411a );
 a41416a <=( a41415a  and  a41408a );
 a41420a <=( A199  and  (not A166) );
 a41421a <=( (not A167)  and  a41420a );
 a41425a <=( (not A202)  and  (not A201) );
 a41426a <=( (not A200)  and  a41425a );
 a41427a <=( a41426a  and  a41421a );
 a41431a <=( A266  and  A265 );
 a41432a <=( (not A203)  and  a41431a );
 a41435a <=( (not A299)  and  A298 );
 a41438a <=( A302  and  A300 );
 a41439a <=( a41438a  and  a41435a );
 a41440a <=( a41439a  and  a41432a );
 a41444a <=( A199  and  (not A166) );
 a41445a <=( (not A167)  and  a41444a );
 a41449a <=( (not A202)  and  (not A201) );
 a41450a <=( (not A200)  and  a41449a );
 a41451a <=( a41450a  and  a41445a );
 a41455a <=( A266  and  A265 );
 a41456a <=( (not A203)  and  a41455a );
 a41459a <=( A299  and  (not A298) );
 a41462a <=( A301  and  A300 );
 a41463a <=( a41462a  and  a41459a );
 a41464a <=( a41463a  and  a41456a );
 a41468a <=( A199  and  (not A166) );
 a41469a <=( (not A167)  and  a41468a );
 a41473a <=( (not A202)  and  (not A201) );
 a41474a <=( (not A200)  and  a41473a );
 a41475a <=( a41474a  and  a41469a );
 a41479a <=( A266  and  A265 );
 a41480a <=( (not A203)  and  a41479a );
 a41483a <=( A299  and  (not A298) );
 a41486a <=( A302  and  A300 );
 a41487a <=( a41486a  and  a41483a );
 a41488a <=( a41487a  and  a41480a );
 a41492a <=( A199  and  (not A166) );
 a41493a <=( (not A167)  and  a41492a );
 a41497a <=( (not A202)  and  (not A201) );
 a41498a <=( (not A200)  and  a41497a );
 a41499a <=( a41498a  and  a41493a );
 a41503a <=( (not A266)  and  (not A265) );
 a41504a <=( (not A203)  and  a41503a );
 a41507a <=( (not A299)  and  A298 );
 a41510a <=( A301  and  A300 );
 a41511a <=( a41510a  and  a41507a );
 a41512a <=( a41511a  and  a41504a );
 a41516a <=( A199  and  (not A166) );
 a41517a <=( (not A167)  and  a41516a );
 a41521a <=( (not A202)  and  (not A201) );
 a41522a <=( (not A200)  and  a41521a );
 a41523a <=( a41522a  and  a41517a );
 a41527a <=( (not A266)  and  (not A265) );
 a41528a <=( (not A203)  and  a41527a );
 a41531a <=( (not A299)  and  A298 );
 a41534a <=( A302  and  A300 );
 a41535a <=( a41534a  and  a41531a );
 a41536a <=( a41535a  and  a41528a );
 a41540a <=( A199  and  (not A166) );
 a41541a <=( (not A167)  and  a41540a );
 a41545a <=( (not A202)  and  (not A201) );
 a41546a <=( (not A200)  and  a41545a );
 a41547a <=( a41546a  and  a41541a );
 a41551a <=( (not A266)  and  (not A265) );
 a41552a <=( (not A203)  and  a41551a );
 a41555a <=( A299  and  (not A298) );
 a41558a <=( A301  and  A300 );
 a41559a <=( a41558a  and  a41555a );
 a41560a <=( a41559a  and  a41552a );
 a41564a <=( A199  and  (not A166) );
 a41565a <=( (not A167)  and  a41564a );
 a41569a <=( (not A202)  and  (not A201) );
 a41570a <=( (not A200)  and  a41569a );
 a41571a <=( a41570a  and  a41565a );
 a41575a <=( (not A266)  and  (not A265) );
 a41576a <=( (not A203)  and  a41575a );
 a41579a <=( A299  and  (not A298) );
 a41582a <=( A302  and  A300 );
 a41583a <=( a41582a  and  a41579a );
 a41584a <=( a41583a  and  a41576a );
 a41588a <=( A167  and  A168 );
 a41589a <=( (not A170)  and  a41588a );
 a41593a <=( (not A202)  and  A201 );
 a41594a <=( (not A166)  and  a41593a );
 a41595a <=( a41594a  and  a41589a );
 a41599a <=( A268  and  (not A267) );
 a41600a <=( (not A203)  and  a41599a );
 a41603a <=( (not A299)  and  A298 );
 a41606a <=( A301  and  A300 );
 a41607a <=( a41606a  and  a41603a );
 a41608a <=( a41607a  and  a41600a );
 a41612a <=( A167  and  A168 );
 a41613a <=( (not A170)  and  a41612a );
 a41617a <=( (not A202)  and  A201 );
 a41618a <=( (not A166)  and  a41617a );
 a41619a <=( a41618a  and  a41613a );
 a41623a <=( A268  and  (not A267) );
 a41624a <=( (not A203)  and  a41623a );
 a41627a <=( (not A299)  and  A298 );
 a41630a <=( A302  and  A300 );
 a41631a <=( a41630a  and  a41627a );
 a41632a <=( a41631a  and  a41624a );
 a41636a <=( A167  and  A168 );
 a41637a <=( (not A170)  and  a41636a );
 a41641a <=( (not A202)  and  A201 );
 a41642a <=( (not A166)  and  a41641a );
 a41643a <=( a41642a  and  a41637a );
 a41647a <=( A268  and  (not A267) );
 a41648a <=( (not A203)  and  a41647a );
 a41651a <=( A299  and  (not A298) );
 a41654a <=( A301  and  A300 );
 a41655a <=( a41654a  and  a41651a );
 a41656a <=( a41655a  and  a41648a );
 a41660a <=( A167  and  A168 );
 a41661a <=( (not A170)  and  a41660a );
 a41665a <=( (not A202)  and  A201 );
 a41666a <=( (not A166)  and  a41665a );
 a41667a <=( a41666a  and  a41661a );
 a41671a <=( A268  and  (not A267) );
 a41672a <=( (not A203)  and  a41671a );
 a41675a <=( A299  and  (not A298) );
 a41678a <=( A302  and  A300 );
 a41679a <=( a41678a  and  a41675a );
 a41680a <=( a41679a  and  a41672a );
 a41684a <=( A167  and  A168 );
 a41685a <=( (not A170)  and  a41684a );
 a41689a <=( (not A202)  and  A201 );
 a41690a <=( (not A166)  and  a41689a );
 a41691a <=( a41690a  and  a41685a );
 a41695a <=( A269  and  (not A267) );
 a41696a <=( (not A203)  and  a41695a );
 a41699a <=( (not A299)  and  A298 );
 a41702a <=( A301  and  A300 );
 a41703a <=( a41702a  and  a41699a );
 a41704a <=( a41703a  and  a41696a );
 a41708a <=( A167  and  A168 );
 a41709a <=( (not A170)  and  a41708a );
 a41713a <=( (not A202)  and  A201 );
 a41714a <=( (not A166)  and  a41713a );
 a41715a <=( a41714a  and  a41709a );
 a41719a <=( A269  and  (not A267) );
 a41720a <=( (not A203)  and  a41719a );
 a41723a <=( (not A299)  and  A298 );
 a41726a <=( A302  and  A300 );
 a41727a <=( a41726a  and  a41723a );
 a41728a <=( a41727a  and  a41720a );
 a41732a <=( A167  and  A168 );
 a41733a <=( (not A170)  and  a41732a );
 a41737a <=( (not A202)  and  A201 );
 a41738a <=( (not A166)  and  a41737a );
 a41739a <=( a41738a  and  a41733a );
 a41743a <=( A269  and  (not A267) );
 a41744a <=( (not A203)  and  a41743a );
 a41747a <=( A299  and  (not A298) );
 a41750a <=( A301  and  A300 );
 a41751a <=( a41750a  and  a41747a );
 a41752a <=( a41751a  and  a41744a );
 a41756a <=( A167  and  A168 );
 a41757a <=( (not A170)  and  a41756a );
 a41761a <=( (not A202)  and  A201 );
 a41762a <=( (not A166)  and  a41761a );
 a41763a <=( a41762a  and  a41757a );
 a41767a <=( A269  and  (not A267) );
 a41768a <=( (not A203)  and  a41767a );
 a41771a <=( A299  and  (not A298) );
 a41774a <=( A302  and  A300 );
 a41775a <=( a41774a  and  a41771a );
 a41776a <=( a41775a  and  a41768a );
 a41780a <=( A167  and  A168 );
 a41781a <=( (not A170)  and  a41780a );
 a41785a <=( (not A202)  and  A201 );
 a41786a <=( (not A166)  and  a41785a );
 a41787a <=( a41786a  and  a41781a );
 a41791a <=( A266  and  A265 );
 a41792a <=( (not A203)  and  a41791a );
 a41795a <=( (not A299)  and  A298 );
 a41798a <=( A301  and  A300 );
 a41799a <=( a41798a  and  a41795a );
 a41800a <=( a41799a  and  a41792a );
 a41804a <=( A167  and  A168 );
 a41805a <=( (not A170)  and  a41804a );
 a41809a <=( (not A202)  and  A201 );
 a41810a <=( (not A166)  and  a41809a );
 a41811a <=( a41810a  and  a41805a );
 a41815a <=( A266  and  A265 );
 a41816a <=( (not A203)  and  a41815a );
 a41819a <=( (not A299)  and  A298 );
 a41822a <=( A302  and  A300 );
 a41823a <=( a41822a  and  a41819a );
 a41824a <=( a41823a  and  a41816a );
 a41828a <=( A167  and  A168 );
 a41829a <=( (not A170)  and  a41828a );
 a41833a <=( (not A202)  and  A201 );
 a41834a <=( (not A166)  and  a41833a );
 a41835a <=( a41834a  and  a41829a );
 a41839a <=( A266  and  A265 );
 a41840a <=( (not A203)  and  a41839a );
 a41843a <=( A299  and  (not A298) );
 a41846a <=( A301  and  A300 );
 a41847a <=( a41846a  and  a41843a );
 a41848a <=( a41847a  and  a41840a );
 a41852a <=( A167  and  A168 );
 a41853a <=( (not A170)  and  a41852a );
 a41857a <=( (not A202)  and  A201 );
 a41858a <=( (not A166)  and  a41857a );
 a41859a <=( a41858a  and  a41853a );
 a41863a <=( A266  and  A265 );
 a41864a <=( (not A203)  and  a41863a );
 a41867a <=( A299  and  (not A298) );
 a41870a <=( A302  and  A300 );
 a41871a <=( a41870a  and  a41867a );
 a41872a <=( a41871a  and  a41864a );
 a41876a <=( A167  and  A168 );
 a41877a <=( (not A170)  and  a41876a );
 a41881a <=( (not A202)  and  A201 );
 a41882a <=( (not A166)  and  a41881a );
 a41883a <=( a41882a  and  a41877a );
 a41887a <=( (not A266)  and  (not A265) );
 a41888a <=( (not A203)  and  a41887a );
 a41891a <=( (not A299)  and  A298 );
 a41894a <=( A301  and  A300 );
 a41895a <=( a41894a  and  a41891a );
 a41896a <=( a41895a  and  a41888a );
 a41900a <=( A167  and  A168 );
 a41901a <=( (not A170)  and  a41900a );
 a41905a <=( (not A202)  and  A201 );
 a41906a <=( (not A166)  and  a41905a );
 a41907a <=( a41906a  and  a41901a );
 a41911a <=( (not A266)  and  (not A265) );
 a41912a <=( (not A203)  and  a41911a );
 a41915a <=( (not A299)  and  A298 );
 a41918a <=( A302  and  A300 );
 a41919a <=( a41918a  and  a41915a );
 a41920a <=( a41919a  and  a41912a );
 a41924a <=( A167  and  A168 );
 a41925a <=( (not A170)  and  a41924a );
 a41929a <=( (not A202)  and  A201 );
 a41930a <=( (not A166)  and  a41929a );
 a41931a <=( a41930a  and  a41925a );
 a41935a <=( (not A266)  and  (not A265) );
 a41936a <=( (not A203)  and  a41935a );
 a41939a <=( A299  and  (not A298) );
 a41942a <=( A301  and  A300 );
 a41943a <=( a41942a  and  a41939a );
 a41944a <=( a41943a  and  a41936a );
 a41948a <=( A167  and  A168 );
 a41949a <=( (not A170)  and  a41948a );
 a41953a <=( (not A202)  and  A201 );
 a41954a <=( (not A166)  and  a41953a );
 a41955a <=( a41954a  and  a41949a );
 a41959a <=( (not A266)  and  (not A265) );
 a41960a <=( (not A203)  and  a41959a );
 a41963a <=( A299  and  (not A298) );
 a41966a <=( A302  and  A300 );
 a41967a <=( a41966a  and  a41963a );
 a41968a <=( a41967a  and  a41960a );
 a41972a <=( A167  and  A168 );
 a41973a <=( (not A170)  and  a41972a );
 a41977a <=( A202  and  (not A201) );
 a41978a <=( (not A166)  and  a41977a );
 a41979a <=( a41978a  and  a41973a );
 a41983a <=( (not A269)  and  (not A268) );
 a41984a <=( A267  and  a41983a );
 a41987a <=( (not A299)  and  A298 );
 a41990a <=( A301  and  A300 );
 a41991a <=( a41990a  and  a41987a );
 a41992a <=( a41991a  and  a41984a );
 a41996a <=( A167  and  A168 );
 a41997a <=( (not A170)  and  a41996a );
 a42001a <=( A202  and  (not A201) );
 a42002a <=( (not A166)  and  a42001a );
 a42003a <=( a42002a  and  a41997a );
 a42007a <=( (not A269)  and  (not A268) );
 a42008a <=( A267  and  a42007a );
 a42011a <=( (not A299)  and  A298 );
 a42014a <=( A302  and  A300 );
 a42015a <=( a42014a  and  a42011a );
 a42016a <=( a42015a  and  a42008a );
 a42020a <=( A167  and  A168 );
 a42021a <=( (not A170)  and  a42020a );
 a42025a <=( A202  and  (not A201) );
 a42026a <=( (not A166)  and  a42025a );
 a42027a <=( a42026a  and  a42021a );
 a42031a <=( (not A269)  and  (not A268) );
 a42032a <=( A267  and  a42031a );
 a42035a <=( A299  and  (not A298) );
 a42038a <=( A301  and  A300 );
 a42039a <=( a42038a  and  a42035a );
 a42040a <=( a42039a  and  a42032a );
 a42044a <=( A167  and  A168 );
 a42045a <=( (not A170)  and  a42044a );
 a42049a <=( A202  and  (not A201) );
 a42050a <=( (not A166)  and  a42049a );
 a42051a <=( a42050a  and  a42045a );
 a42055a <=( (not A269)  and  (not A268) );
 a42056a <=( A267  and  a42055a );
 a42059a <=( A299  and  (not A298) );
 a42062a <=( A302  and  A300 );
 a42063a <=( a42062a  and  a42059a );
 a42064a <=( a42063a  and  a42056a );
 a42068a <=( A167  and  A168 );
 a42069a <=( (not A170)  and  a42068a );
 a42073a <=( A202  and  (not A201) );
 a42074a <=( (not A166)  and  a42073a );
 a42075a <=( a42074a  and  a42069a );
 a42079a <=( A298  and  A268 );
 a42080a <=( (not A267)  and  a42079a );
 a42083a <=( (not A300)  and  (not A299) );
 a42086a <=( (not A302)  and  (not A301) );
 a42087a <=( a42086a  and  a42083a );
 a42088a <=( a42087a  and  a42080a );
 a42092a <=( A167  and  A168 );
 a42093a <=( (not A170)  and  a42092a );
 a42097a <=( A202  and  (not A201) );
 a42098a <=( (not A166)  and  a42097a );
 a42099a <=( a42098a  and  a42093a );
 a42103a <=( (not A298)  and  A268 );
 a42104a <=( (not A267)  and  a42103a );
 a42107a <=( (not A300)  and  A299 );
 a42110a <=( (not A302)  and  (not A301) );
 a42111a <=( a42110a  and  a42107a );
 a42112a <=( a42111a  and  a42104a );
 a42116a <=( A167  and  A168 );
 a42117a <=( (not A170)  and  a42116a );
 a42121a <=( A202  and  (not A201) );
 a42122a <=( (not A166)  and  a42121a );
 a42123a <=( a42122a  and  a42117a );
 a42127a <=( A298  and  A269 );
 a42128a <=( (not A267)  and  a42127a );
 a42131a <=( (not A300)  and  (not A299) );
 a42134a <=( (not A302)  and  (not A301) );
 a42135a <=( a42134a  and  a42131a );
 a42136a <=( a42135a  and  a42128a );
 a42140a <=( A167  and  A168 );
 a42141a <=( (not A170)  and  a42140a );
 a42145a <=( A202  and  (not A201) );
 a42146a <=( (not A166)  and  a42145a );
 a42147a <=( a42146a  and  a42141a );
 a42151a <=( (not A298)  and  A269 );
 a42152a <=( (not A267)  and  a42151a );
 a42155a <=( (not A300)  and  A299 );
 a42158a <=( (not A302)  and  (not A301) );
 a42159a <=( a42158a  and  a42155a );
 a42160a <=( a42159a  and  a42152a );
 a42164a <=( A167  and  A168 );
 a42165a <=( (not A170)  and  a42164a );
 a42169a <=( A202  and  (not A201) );
 a42170a <=( (not A166)  and  a42169a );
 a42171a <=( a42170a  and  a42165a );
 a42175a <=( A298  and  A266 );
 a42176a <=( A265  and  a42175a );
 a42179a <=( (not A300)  and  (not A299) );
 a42182a <=( (not A302)  and  (not A301) );
 a42183a <=( a42182a  and  a42179a );
 a42184a <=( a42183a  and  a42176a );
 a42188a <=( A167  and  A168 );
 a42189a <=( (not A170)  and  a42188a );
 a42193a <=( A202  and  (not A201) );
 a42194a <=( (not A166)  and  a42193a );
 a42195a <=( a42194a  and  a42189a );
 a42199a <=( (not A298)  and  A266 );
 a42200a <=( A265  and  a42199a );
 a42203a <=( (not A300)  and  A299 );
 a42206a <=( (not A302)  and  (not A301) );
 a42207a <=( a42206a  and  a42203a );
 a42208a <=( a42207a  and  a42200a );
 a42212a <=( A167  and  A168 );
 a42213a <=( (not A170)  and  a42212a );
 a42217a <=( A202  and  (not A201) );
 a42218a <=( (not A166)  and  a42217a );
 a42219a <=( a42218a  and  a42213a );
 a42223a <=( A298  and  (not A266) );
 a42224a <=( (not A265)  and  a42223a );
 a42227a <=( (not A300)  and  (not A299) );
 a42230a <=( (not A302)  and  (not A301) );
 a42231a <=( a42230a  and  a42227a );
 a42232a <=( a42231a  and  a42224a );
 a42236a <=( A167  and  A168 );
 a42237a <=( (not A170)  and  a42236a );
 a42241a <=( A202  and  (not A201) );
 a42242a <=( (not A166)  and  a42241a );
 a42243a <=( a42242a  and  a42237a );
 a42247a <=( (not A298)  and  (not A266) );
 a42248a <=( (not A265)  and  a42247a );
 a42251a <=( (not A300)  and  A299 );
 a42254a <=( (not A302)  and  (not A301) );
 a42255a <=( a42254a  and  a42251a );
 a42256a <=( a42255a  and  a42248a );
 a42260a <=( A167  and  A168 );
 a42261a <=( (not A170)  and  a42260a );
 a42265a <=( A203  and  (not A201) );
 a42266a <=( (not A166)  and  a42265a );
 a42267a <=( a42266a  and  a42261a );
 a42271a <=( (not A269)  and  (not A268) );
 a42272a <=( A267  and  a42271a );
 a42275a <=( (not A299)  and  A298 );
 a42278a <=( A301  and  A300 );
 a42279a <=( a42278a  and  a42275a );
 a42280a <=( a42279a  and  a42272a );
 a42284a <=( A167  and  A168 );
 a42285a <=( (not A170)  and  a42284a );
 a42289a <=( A203  and  (not A201) );
 a42290a <=( (not A166)  and  a42289a );
 a42291a <=( a42290a  and  a42285a );
 a42295a <=( (not A269)  and  (not A268) );
 a42296a <=( A267  and  a42295a );
 a42299a <=( (not A299)  and  A298 );
 a42302a <=( A302  and  A300 );
 a42303a <=( a42302a  and  a42299a );
 a42304a <=( a42303a  and  a42296a );
 a42308a <=( A167  and  A168 );
 a42309a <=( (not A170)  and  a42308a );
 a42313a <=( A203  and  (not A201) );
 a42314a <=( (not A166)  and  a42313a );
 a42315a <=( a42314a  and  a42309a );
 a42319a <=( (not A269)  and  (not A268) );
 a42320a <=( A267  and  a42319a );
 a42323a <=( A299  and  (not A298) );
 a42326a <=( A301  and  A300 );
 a42327a <=( a42326a  and  a42323a );
 a42328a <=( a42327a  and  a42320a );
 a42332a <=( A167  and  A168 );
 a42333a <=( (not A170)  and  a42332a );
 a42337a <=( A203  and  (not A201) );
 a42338a <=( (not A166)  and  a42337a );
 a42339a <=( a42338a  and  a42333a );
 a42343a <=( (not A269)  and  (not A268) );
 a42344a <=( A267  and  a42343a );
 a42347a <=( A299  and  (not A298) );
 a42350a <=( A302  and  A300 );
 a42351a <=( a42350a  and  a42347a );
 a42352a <=( a42351a  and  a42344a );
 a42356a <=( A167  and  A168 );
 a42357a <=( (not A170)  and  a42356a );
 a42361a <=( A203  and  (not A201) );
 a42362a <=( (not A166)  and  a42361a );
 a42363a <=( a42362a  and  a42357a );
 a42367a <=( A298  and  A268 );
 a42368a <=( (not A267)  and  a42367a );
 a42371a <=( (not A300)  and  (not A299) );
 a42374a <=( (not A302)  and  (not A301) );
 a42375a <=( a42374a  and  a42371a );
 a42376a <=( a42375a  and  a42368a );
 a42380a <=( A167  and  A168 );
 a42381a <=( (not A170)  and  a42380a );
 a42385a <=( A203  and  (not A201) );
 a42386a <=( (not A166)  and  a42385a );
 a42387a <=( a42386a  and  a42381a );
 a42391a <=( (not A298)  and  A268 );
 a42392a <=( (not A267)  and  a42391a );
 a42395a <=( (not A300)  and  A299 );
 a42398a <=( (not A302)  and  (not A301) );
 a42399a <=( a42398a  and  a42395a );
 a42400a <=( a42399a  and  a42392a );
 a42404a <=( A167  and  A168 );
 a42405a <=( (not A170)  and  a42404a );
 a42409a <=( A203  and  (not A201) );
 a42410a <=( (not A166)  and  a42409a );
 a42411a <=( a42410a  and  a42405a );
 a42415a <=( A298  and  A269 );
 a42416a <=( (not A267)  and  a42415a );
 a42419a <=( (not A300)  and  (not A299) );
 a42422a <=( (not A302)  and  (not A301) );
 a42423a <=( a42422a  and  a42419a );
 a42424a <=( a42423a  and  a42416a );
 a42428a <=( A167  and  A168 );
 a42429a <=( (not A170)  and  a42428a );
 a42433a <=( A203  and  (not A201) );
 a42434a <=( (not A166)  and  a42433a );
 a42435a <=( a42434a  and  a42429a );
 a42439a <=( (not A298)  and  A269 );
 a42440a <=( (not A267)  and  a42439a );
 a42443a <=( (not A300)  and  A299 );
 a42446a <=( (not A302)  and  (not A301) );
 a42447a <=( a42446a  and  a42443a );
 a42448a <=( a42447a  and  a42440a );
 a42452a <=( A167  and  A168 );
 a42453a <=( (not A170)  and  a42452a );
 a42457a <=( A203  and  (not A201) );
 a42458a <=( (not A166)  and  a42457a );
 a42459a <=( a42458a  and  a42453a );
 a42463a <=( A298  and  A266 );
 a42464a <=( A265  and  a42463a );
 a42467a <=( (not A300)  and  (not A299) );
 a42470a <=( (not A302)  and  (not A301) );
 a42471a <=( a42470a  and  a42467a );
 a42472a <=( a42471a  and  a42464a );
 a42476a <=( A167  and  A168 );
 a42477a <=( (not A170)  and  a42476a );
 a42481a <=( A203  and  (not A201) );
 a42482a <=( (not A166)  and  a42481a );
 a42483a <=( a42482a  and  a42477a );
 a42487a <=( (not A298)  and  A266 );
 a42488a <=( A265  and  a42487a );
 a42491a <=( (not A300)  and  A299 );
 a42494a <=( (not A302)  and  (not A301) );
 a42495a <=( a42494a  and  a42491a );
 a42496a <=( a42495a  and  a42488a );
 a42500a <=( A167  and  A168 );
 a42501a <=( (not A170)  and  a42500a );
 a42505a <=( A203  and  (not A201) );
 a42506a <=( (not A166)  and  a42505a );
 a42507a <=( a42506a  and  a42501a );
 a42511a <=( A298  and  (not A266) );
 a42512a <=( (not A265)  and  a42511a );
 a42515a <=( (not A300)  and  (not A299) );
 a42518a <=( (not A302)  and  (not A301) );
 a42519a <=( a42518a  and  a42515a );
 a42520a <=( a42519a  and  a42512a );
 a42524a <=( A167  and  A168 );
 a42525a <=( (not A170)  and  a42524a );
 a42529a <=( A203  and  (not A201) );
 a42530a <=( (not A166)  and  a42529a );
 a42531a <=( a42530a  and  a42525a );
 a42535a <=( (not A298)  and  (not A266) );
 a42536a <=( (not A265)  and  a42535a );
 a42539a <=( (not A300)  and  A299 );
 a42542a <=( (not A302)  and  (not A301) );
 a42543a <=( a42542a  and  a42539a );
 a42544a <=( a42543a  and  a42536a );
 a42548a <=( A167  and  A168 );
 a42549a <=( (not A170)  and  a42548a );
 a42553a <=( A200  and  A199 );
 a42554a <=( (not A166)  and  a42553a );
 a42555a <=( a42554a  and  a42549a );
 a42559a <=( (not A269)  and  (not A268) );
 a42560a <=( A267  and  a42559a );
 a42563a <=( (not A299)  and  A298 );
 a42566a <=( A301  and  A300 );
 a42567a <=( a42566a  and  a42563a );
 a42568a <=( a42567a  and  a42560a );
 a42572a <=( A167  and  A168 );
 a42573a <=( (not A170)  and  a42572a );
 a42577a <=( A200  and  A199 );
 a42578a <=( (not A166)  and  a42577a );
 a42579a <=( a42578a  and  a42573a );
 a42583a <=( (not A269)  and  (not A268) );
 a42584a <=( A267  and  a42583a );
 a42587a <=( (not A299)  and  A298 );
 a42590a <=( A302  and  A300 );
 a42591a <=( a42590a  and  a42587a );
 a42592a <=( a42591a  and  a42584a );
 a42596a <=( A167  and  A168 );
 a42597a <=( (not A170)  and  a42596a );
 a42601a <=( A200  and  A199 );
 a42602a <=( (not A166)  and  a42601a );
 a42603a <=( a42602a  and  a42597a );
 a42607a <=( (not A269)  and  (not A268) );
 a42608a <=( A267  and  a42607a );
 a42611a <=( A299  and  (not A298) );
 a42614a <=( A301  and  A300 );
 a42615a <=( a42614a  and  a42611a );
 a42616a <=( a42615a  and  a42608a );
 a42620a <=( A167  and  A168 );
 a42621a <=( (not A170)  and  a42620a );
 a42625a <=( A200  and  A199 );
 a42626a <=( (not A166)  and  a42625a );
 a42627a <=( a42626a  and  a42621a );
 a42631a <=( (not A269)  and  (not A268) );
 a42632a <=( A267  and  a42631a );
 a42635a <=( A299  and  (not A298) );
 a42638a <=( A302  and  A300 );
 a42639a <=( a42638a  and  a42635a );
 a42640a <=( a42639a  and  a42632a );
 a42644a <=( A167  and  A168 );
 a42645a <=( (not A170)  and  a42644a );
 a42649a <=( A200  and  A199 );
 a42650a <=( (not A166)  and  a42649a );
 a42651a <=( a42650a  and  a42645a );
 a42655a <=( A298  and  A268 );
 a42656a <=( (not A267)  and  a42655a );
 a42659a <=( (not A300)  and  (not A299) );
 a42662a <=( (not A302)  and  (not A301) );
 a42663a <=( a42662a  and  a42659a );
 a42664a <=( a42663a  and  a42656a );
 a42668a <=( A167  and  A168 );
 a42669a <=( (not A170)  and  a42668a );
 a42673a <=( A200  and  A199 );
 a42674a <=( (not A166)  and  a42673a );
 a42675a <=( a42674a  and  a42669a );
 a42679a <=( (not A298)  and  A268 );
 a42680a <=( (not A267)  and  a42679a );
 a42683a <=( (not A300)  and  A299 );
 a42686a <=( (not A302)  and  (not A301) );
 a42687a <=( a42686a  and  a42683a );
 a42688a <=( a42687a  and  a42680a );
 a42692a <=( A167  and  A168 );
 a42693a <=( (not A170)  and  a42692a );
 a42697a <=( A200  and  A199 );
 a42698a <=( (not A166)  and  a42697a );
 a42699a <=( a42698a  and  a42693a );
 a42703a <=( A298  and  A269 );
 a42704a <=( (not A267)  and  a42703a );
 a42707a <=( (not A300)  and  (not A299) );
 a42710a <=( (not A302)  and  (not A301) );
 a42711a <=( a42710a  and  a42707a );
 a42712a <=( a42711a  and  a42704a );
 a42716a <=( A167  and  A168 );
 a42717a <=( (not A170)  and  a42716a );
 a42721a <=( A200  and  A199 );
 a42722a <=( (not A166)  and  a42721a );
 a42723a <=( a42722a  and  a42717a );
 a42727a <=( (not A298)  and  A269 );
 a42728a <=( (not A267)  and  a42727a );
 a42731a <=( (not A300)  and  A299 );
 a42734a <=( (not A302)  and  (not A301) );
 a42735a <=( a42734a  and  a42731a );
 a42736a <=( a42735a  and  a42728a );
 a42740a <=( A167  and  A168 );
 a42741a <=( (not A170)  and  a42740a );
 a42745a <=( A200  and  A199 );
 a42746a <=( (not A166)  and  a42745a );
 a42747a <=( a42746a  and  a42741a );
 a42751a <=( A298  and  A266 );
 a42752a <=( A265  and  a42751a );
 a42755a <=( (not A300)  and  (not A299) );
 a42758a <=( (not A302)  and  (not A301) );
 a42759a <=( a42758a  and  a42755a );
 a42760a <=( a42759a  and  a42752a );
 a42764a <=( A167  and  A168 );
 a42765a <=( (not A170)  and  a42764a );
 a42769a <=( A200  and  A199 );
 a42770a <=( (not A166)  and  a42769a );
 a42771a <=( a42770a  and  a42765a );
 a42775a <=( (not A298)  and  A266 );
 a42776a <=( A265  and  a42775a );
 a42779a <=( (not A300)  and  A299 );
 a42782a <=( (not A302)  and  (not A301) );
 a42783a <=( a42782a  and  a42779a );
 a42784a <=( a42783a  and  a42776a );
 a42788a <=( A167  and  A168 );
 a42789a <=( (not A170)  and  a42788a );
 a42793a <=( A200  and  A199 );
 a42794a <=( (not A166)  and  a42793a );
 a42795a <=( a42794a  and  a42789a );
 a42799a <=( A298  and  (not A266) );
 a42800a <=( (not A265)  and  a42799a );
 a42803a <=( (not A300)  and  (not A299) );
 a42806a <=( (not A302)  and  (not A301) );
 a42807a <=( a42806a  and  a42803a );
 a42808a <=( a42807a  and  a42800a );
 a42812a <=( A167  and  A168 );
 a42813a <=( (not A170)  and  a42812a );
 a42817a <=( A200  and  A199 );
 a42818a <=( (not A166)  and  a42817a );
 a42819a <=( a42818a  and  a42813a );
 a42823a <=( (not A298)  and  (not A266) );
 a42824a <=( (not A265)  and  a42823a );
 a42827a <=( (not A300)  and  A299 );
 a42830a <=( (not A302)  and  (not A301) );
 a42831a <=( a42830a  and  a42827a );
 a42832a <=( a42831a  and  a42824a );
 a42836a <=( A167  and  A168 );
 a42837a <=( (not A170)  and  a42836a );
 a42841a <=( (not A200)  and  (not A199) );
 a42842a <=( (not A166)  and  a42841a );
 a42843a <=( a42842a  and  a42837a );
 a42847a <=( (not A269)  and  (not A268) );
 a42848a <=( A267  and  a42847a );
 a42851a <=( (not A299)  and  A298 );
 a42854a <=( A301  and  A300 );
 a42855a <=( a42854a  and  a42851a );
 a42856a <=( a42855a  and  a42848a );
 a42860a <=( A167  and  A168 );
 a42861a <=( (not A170)  and  a42860a );
 a42865a <=( (not A200)  and  (not A199) );
 a42866a <=( (not A166)  and  a42865a );
 a42867a <=( a42866a  and  a42861a );
 a42871a <=( (not A269)  and  (not A268) );
 a42872a <=( A267  and  a42871a );
 a42875a <=( (not A299)  and  A298 );
 a42878a <=( A302  and  A300 );
 a42879a <=( a42878a  and  a42875a );
 a42880a <=( a42879a  and  a42872a );
 a42884a <=( A167  and  A168 );
 a42885a <=( (not A170)  and  a42884a );
 a42889a <=( (not A200)  and  (not A199) );
 a42890a <=( (not A166)  and  a42889a );
 a42891a <=( a42890a  and  a42885a );
 a42895a <=( (not A269)  and  (not A268) );
 a42896a <=( A267  and  a42895a );
 a42899a <=( A299  and  (not A298) );
 a42902a <=( A301  and  A300 );
 a42903a <=( a42902a  and  a42899a );
 a42904a <=( a42903a  and  a42896a );
 a42908a <=( A167  and  A168 );
 a42909a <=( (not A170)  and  a42908a );
 a42913a <=( (not A200)  and  (not A199) );
 a42914a <=( (not A166)  and  a42913a );
 a42915a <=( a42914a  and  a42909a );
 a42919a <=( (not A269)  and  (not A268) );
 a42920a <=( A267  and  a42919a );
 a42923a <=( A299  and  (not A298) );
 a42926a <=( A302  and  A300 );
 a42927a <=( a42926a  and  a42923a );
 a42928a <=( a42927a  and  a42920a );
 a42932a <=( A167  and  A168 );
 a42933a <=( (not A170)  and  a42932a );
 a42937a <=( (not A200)  and  (not A199) );
 a42938a <=( (not A166)  and  a42937a );
 a42939a <=( a42938a  and  a42933a );
 a42943a <=( A298  and  A268 );
 a42944a <=( (not A267)  and  a42943a );
 a42947a <=( (not A300)  and  (not A299) );
 a42950a <=( (not A302)  and  (not A301) );
 a42951a <=( a42950a  and  a42947a );
 a42952a <=( a42951a  and  a42944a );
 a42956a <=( A167  and  A168 );
 a42957a <=( (not A170)  and  a42956a );
 a42961a <=( (not A200)  and  (not A199) );
 a42962a <=( (not A166)  and  a42961a );
 a42963a <=( a42962a  and  a42957a );
 a42967a <=( (not A298)  and  A268 );
 a42968a <=( (not A267)  and  a42967a );
 a42971a <=( (not A300)  and  A299 );
 a42974a <=( (not A302)  and  (not A301) );
 a42975a <=( a42974a  and  a42971a );
 a42976a <=( a42975a  and  a42968a );
 a42980a <=( A167  and  A168 );
 a42981a <=( (not A170)  and  a42980a );
 a42985a <=( (not A200)  and  (not A199) );
 a42986a <=( (not A166)  and  a42985a );
 a42987a <=( a42986a  and  a42981a );
 a42991a <=( A298  and  A269 );
 a42992a <=( (not A267)  and  a42991a );
 a42995a <=( (not A300)  and  (not A299) );
 a42998a <=( (not A302)  and  (not A301) );
 a42999a <=( a42998a  and  a42995a );
 a43000a <=( a42999a  and  a42992a );
 a43004a <=( A167  and  A168 );
 a43005a <=( (not A170)  and  a43004a );
 a43009a <=( (not A200)  and  (not A199) );
 a43010a <=( (not A166)  and  a43009a );
 a43011a <=( a43010a  and  a43005a );
 a43015a <=( (not A298)  and  A269 );
 a43016a <=( (not A267)  and  a43015a );
 a43019a <=( (not A300)  and  A299 );
 a43022a <=( (not A302)  and  (not A301) );
 a43023a <=( a43022a  and  a43019a );
 a43024a <=( a43023a  and  a43016a );
 a43028a <=( A167  and  A168 );
 a43029a <=( (not A170)  and  a43028a );
 a43033a <=( (not A200)  and  (not A199) );
 a43034a <=( (not A166)  and  a43033a );
 a43035a <=( a43034a  and  a43029a );
 a43039a <=( A298  and  A266 );
 a43040a <=( A265  and  a43039a );
 a43043a <=( (not A300)  and  (not A299) );
 a43046a <=( (not A302)  and  (not A301) );
 a43047a <=( a43046a  and  a43043a );
 a43048a <=( a43047a  and  a43040a );
 a43052a <=( A167  and  A168 );
 a43053a <=( (not A170)  and  a43052a );
 a43057a <=( (not A200)  and  (not A199) );
 a43058a <=( (not A166)  and  a43057a );
 a43059a <=( a43058a  and  a43053a );
 a43063a <=( (not A298)  and  A266 );
 a43064a <=( A265  and  a43063a );
 a43067a <=( (not A300)  and  A299 );
 a43070a <=( (not A302)  and  (not A301) );
 a43071a <=( a43070a  and  a43067a );
 a43072a <=( a43071a  and  a43064a );
 a43076a <=( A167  and  A168 );
 a43077a <=( (not A170)  and  a43076a );
 a43081a <=( (not A200)  and  (not A199) );
 a43082a <=( (not A166)  and  a43081a );
 a43083a <=( a43082a  and  a43077a );
 a43087a <=( A298  and  (not A266) );
 a43088a <=( (not A265)  and  a43087a );
 a43091a <=( (not A300)  and  (not A299) );
 a43094a <=( (not A302)  and  (not A301) );
 a43095a <=( a43094a  and  a43091a );
 a43096a <=( a43095a  and  a43088a );
 a43100a <=( A167  and  A168 );
 a43101a <=( (not A170)  and  a43100a );
 a43105a <=( (not A200)  and  (not A199) );
 a43106a <=( (not A166)  and  a43105a );
 a43107a <=( a43106a  and  a43101a );
 a43111a <=( (not A298)  and  (not A266) );
 a43112a <=( (not A265)  and  a43111a );
 a43115a <=( (not A300)  and  A299 );
 a43118a <=( (not A302)  and  (not A301) );
 a43119a <=( a43118a  and  a43115a );
 a43120a <=( a43119a  and  a43112a );
 a43124a <=( (not A167)  and  A168 );
 a43125a <=( (not A170)  and  a43124a );
 a43129a <=( (not A202)  and  A201 );
 a43130a <=( A166  and  a43129a );
 a43131a <=( a43130a  and  a43125a );
 a43135a <=( A268  and  (not A267) );
 a43136a <=( (not A203)  and  a43135a );
 a43139a <=( (not A299)  and  A298 );
 a43142a <=( A301  and  A300 );
 a43143a <=( a43142a  and  a43139a );
 a43144a <=( a43143a  and  a43136a );
 a43148a <=( (not A167)  and  A168 );
 a43149a <=( (not A170)  and  a43148a );
 a43153a <=( (not A202)  and  A201 );
 a43154a <=( A166  and  a43153a );
 a43155a <=( a43154a  and  a43149a );
 a43159a <=( A268  and  (not A267) );
 a43160a <=( (not A203)  and  a43159a );
 a43163a <=( (not A299)  and  A298 );
 a43166a <=( A302  and  A300 );
 a43167a <=( a43166a  and  a43163a );
 a43168a <=( a43167a  and  a43160a );
 a43172a <=( (not A167)  and  A168 );
 a43173a <=( (not A170)  and  a43172a );
 a43177a <=( (not A202)  and  A201 );
 a43178a <=( A166  and  a43177a );
 a43179a <=( a43178a  and  a43173a );
 a43183a <=( A268  and  (not A267) );
 a43184a <=( (not A203)  and  a43183a );
 a43187a <=( A299  and  (not A298) );
 a43190a <=( A301  and  A300 );
 a43191a <=( a43190a  and  a43187a );
 a43192a <=( a43191a  and  a43184a );
 a43196a <=( (not A167)  and  A168 );
 a43197a <=( (not A170)  and  a43196a );
 a43201a <=( (not A202)  and  A201 );
 a43202a <=( A166  and  a43201a );
 a43203a <=( a43202a  and  a43197a );
 a43207a <=( A268  and  (not A267) );
 a43208a <=( (not A203)  and  a43207a );
 a43211a <=( A299  and  (not A298) );
 a43214a <=( A302  and  A300 );
 a43215a <=( a43214a  and  a43211a );
 a43216a <=( a43215a  and  a43208a );
 a43220a <=( (not A167)  and  A168 );
 a43221a <=( (not A170)  and  a43220a );
 a43225a <=( (not A202)  and  A201 );
 a43226a <=( A166  and  a43225a );
 a43227a <=( a43226a  and  a43221a );
 a43231a <=( A269  and  (not A267) );
 a43232a <=( (not A203)  and  a43231a );
 a43235a <=( (not A299)  and  A298 );
 a43238a <=( A301  and  A300 );
 a43239a <=( a43238a  and  a43235a );
 a43240a <=( a43239a  and  a43232a );
 a43244a <=( (not A167)  and  A168 );
 a43245a <=( (not A170)  and  a43244a );
 a43249a <=( (not A202)  and  A201 );
 a43250a <=( A166  and  a43249a );
 a43251a <=( a43250a  and  a43245a );
 a43255a <=( A269  and  (not A267) );
 a43256a <=( (not A203)  and  a43255a );
 a43259a <=( (not A299)  and  A298 );
 a43262a <=( A302  and  A300 );
 a43263a <=( a43262a  and  a43259a );
 a43264a <=( a43263a  and  a43256a );
 a43268a <=( (not A167)  and  A168 );
 a43269a <=( (not A170)  and  a43268a );
 a43273a <=( (not A202)  and  A201 );
 a43274a <=( A166  and  a43273a );
 a43275a <=( a43274a  and  a43269a );
 a43279a <=( A269  and  (not A267) );
 a43280a <=( (not A203)  and  a43279a );
 a43283a <=( A299  and  (not A298) );
 a43286a <=( A301  and  A300 );
 a43287a <=( a43286a  and  a43283a );
 a43288a <=( a43287a  and  a43280a );
 a43292a <=( (not A167)  and  A168 );
 a43293a <=( (not A170)  and  a43292a );
 a43297a <=( (not A202)  and  A201 );
 a43298a <=( A166  and  a43297a );
 a43299a <=( a43298a  and  a43293a );
 a43303a <=( A269  and  (not A267) );
 a43304a <=( (not A203)  and  a43303a );
 a43307a <=( A299  and  (not A298) );
 a43310a <=( A302  and  A300 );
 a43311a <=( a43310a  and  a43307a );
 a43312a <=( a43311a  and  a43304a );
 a43316a <=( (not A167)  and  A168 );
 a43317a <=( (not A170)  and  a43316a );
 a43321a <=( (not A202)  and  A201 );
 a43322a <=( A166  and  a43321a );
 a43323a <=( a43322a  and  a43317a );
 a43327a <=( A266  and  A265 );
 a43328a <=( (not A203)  and  a43327a );
 a43331a <=( (not A299)  and  A298 );
 a43334a <=( A301  and  A300 );
 a43335a <=( a43334a  and  a43331a );
 a43336a <=( a43335a  and  a43328a );
 a43340a <=( (not A167)  and  A168 );
 a43341a <=( (not A170)  and  a43340a );
 a43345a <=( (not A202)  and  A201 );
 a43346a <=( A166  and  a43345a );
 a43347a <=( a43346a  and  a43341a );
 a43351a <=( A266  and  A265 );
 a43352a <=( (not A203)  and  a43351a );
 a43355a <=( (not A299)  and  A298 );
 a43358a <=( A302  and  A300 );
 a43359a <=( a43358a  and  a43355a );
 a43360a <=( a43359a  and  a43352a );
 a43364a <=( (not A167)  and  A168 );
 a43365a <=( (not A170)  and  a43364a );
 a43369a <=( (not A202)  and  A201 );
 a43370a <=( A166  and  a43369a );
 a43371a <=( a43370a  and  a43365a );
 a43375a <=( A266  and  A265 );
 a43376a <=( (not A203)  and  a43375a );
 a43379a <=( A299  and  (not A298) );
 a43382a <=( A301  and  A300 );
 a43383a <=( a43382a  and  a43379a );
 a43384a <=( a43383a  and  a43376a );
 a43388a <=( (not A167)  and  A168 );
 a43389a <=( (not A170)  and  a43388a );
 a43393a <=( (not A202)  and  A201 );
 a43394a <=( A166  and  a43393a );
 a43395a <=( a43394a  and  a43389a );
 a43399a <=( A266  and  A265 );
 a43400a <=( (not A203)  and  a43399a );
 a43403a <=( A299  and  (not A298) );
 a43406a <=( A302  and  A300 );
 a43407a <=( a43406a  and  a43403a );
 a43408a <=( a43407a  and  a43400a );
 a43412a <=( (not A167)  and  A168 );
 a43413a <=( (not A170)  and  a43412a );
 a43417a <=( (not A202)  and  A201 );
 a43418a <=( A166  and  a43417a );
 a43419a <=( a43418a  and  a43413a );
 a43423a <=( (not A266)  and  (not A265) );
 a43424a <=( (not A203)  and  a43423a );
 a43427a <=( (not A299)  and  A298 );
 a43430a <=( A301  and  A300 );
 a43431a <=( a43430a  and  a43427a );
 a43432a <=( a43431a  and  a43424a );
 a43436a <=( (not A167)  and  A168 );
 a43437a <=( (not A170)  and  a43436a );
 a43441a <=( (not A202)  and  A201 );
 a43442a <=( A166  and  a43441a );
 a43443a <=( a43442a  and  a43437a );
 a43447a <=( (not A266)  and  (not A265) );
 a43448a <=( (not A203)  and  a43447a );
 a43451a <=( (not A299)  and  A298 );
 a43454a <=( A302  and  A300 );
 a43455a <=( a43454a  and  a43451a );
 a43456a <=( a43455a  and  a43448a );
 a43460a <=( (not A167)  and  A168 );
 a43461a <=( (not A170)  and  a43460a );
 a43465a <=( (not A202)  and  A201 );
 a43466a <=( A166  and  a43465a );
 a43467a <=( a43466a  and  a43461a );
 a43471a <=( (not A266)  and  (not A265) );
 a43472a <=( (not A203)  and  a43471a );
 a43475a <=( A299  and  (not A298) );
 a43478a <=( A301  and  A300 );
 a43479a <=( a43478a  and  a43475a );
 a43480a <=( a43479a  and  a43472a );
 a43484a <=( (not A167)  and  A168 );
 a43485a <=( (not A170)  and  a43484a );
 a43489a <=( (not A202)  and  A201 );
 a43490a <=( A166  and  a43489a );
 a43491a <=( a43490a  and  a43485a );
 a43495a <=( (not A266)  and  (not A265) );
 a43496a <=( (not A203)  and  a43495a );
 a43499a <=( A299  and  (not A298) );
 a43502a <=( A302  and  A300 );
 a43503a <=( a43502a  and  a43499a );
 a43504a <=( a43503a  and  a43496a );
 a43508a <=( (not A167)  and  A168 );
 a43509a <=( (not A170)  and  a43508a );
 a43513a <=( A202  and  (not A201) );
 a43514a <=( A166  and  a43513a );
 a43515a <=( a43514a  and  a43509a );
 a43519a <=( (not A269)  and  (not A268) );
 a43520a <=( A267  and  a43519a );
 a43523a <=( (not A299)  and  A298 );
 a43526a <=( A301  and  A300 );
 a43527a <=( a43526a  and  a43523a );
 a43528a <=( a43527a  and  a43520a );
 a43532a <=( (not A167)  and  A168 );
 a43533a <=( (not A170)  and  a43532a );
 a43537a <=( A202  and  (not A201) );
 a43538a <=( A166  and  a43537a );
 a43539a <=( a43538a  and  a43533a );
 a43543a <=( (not A269)  and  (not A268) );
 a43544a <=( A267  and  a43543a );
 a43547a <=( (not A299)  and  A298 );
 a43550a <=( A302  and  A300 );
 a43551a <=( a43550a  and  a43547a );
 a43552a <=( a43551a  and  a43544a );
 a43556a <=( (not A167)  and  A168 );
 a43557a <=( (not A170)  and  a43556a );
 a43561a <=( A202  and  (not A201) );
 a43562a <=( A166  and  a43561a );
 a43563a <=( a43562a  and  a43557a );
 a43567a <=( (not A269)  and  (not A268) );
 a43568a <=( A267  and  a43567a );
 a43571a <=( A299  and  (not A298) );
 a43574a <=( A301  and  A300 );
 a43575a <=( a43574a  and  a43571a );
 a43576a <=( a43575a  and  a43568a );
 a43580a <=( (not A167)  and  A168 );
 a43581a <=( (not A170)  and  a43580a );
 a43585a <=( A202  and  (not A201) );
 a43586a <=( A166  and  a43585a );
 a43587a <=( a43586a  and  a43581a );
 a43591a <=( (not A269)  and  (not A268) );
 a43592a <=( A267  and  a43591a );
 a43595a <=( A299  and  (not A298) );
 a43598a <=( A302  and  A300 );
 a43599a <=( a43598a  and  a43595a );
 a43600a <=( a43599a  and  a43592a );
 a43604a <=( (not A167)  and  A168 );
 a43605a <=( (not A170)  and  a43604a );
 a43609a <=( A202  and  (not A201) );
 a43610a <=( A166  and  a43609a );
 a43611a <=( a43610a  and  a43605a );
 a43615a <=( A298  and  A268 );
 a43616a <=( (not A267)  and  a43615a );
 a43619a <=( (not A300)  and  (not A299) );
 a43622a <=( (not A302)  and  (not A301) );
 a43623a <=( a43622a  and  a43619a );
 a43624a <=( a43623a  and  a43616a );
 a43628a <=( (not A167)  and  A168 );
 a43629a <=( (not A170)  and  a43628a );
 a43633a <=( A202  and  (not A201) );
 a43634a <=( A166  and  a43633a );
 a43635a <=( a43634a  and  a43629a );
 a43639a <=( (not A298)  and  A268 );
 a43640a <=( (not A267)  and  a43639a );
 a43643a <=( (not A300)  and  A299 );
 a43646a <=( (not A302)  and  (not A301) );
 a43647a <=( a43646a  and  a43643a );
 a43648a <=( a43647a  and  a43640a );
 a43652a <=( (not A167)  and  A168 );
 a43653a <=( (not A170)  and  a43652a );
 a43657a <=( A202  and  (not A201) );
 a43658a <=( A166  and  a43657a );
 a43659a <=( a43658a  and  a43653a );
 a43663a <=( A298  and  A269 );
 a43664a <=( (not A267)  and  a43663a );
 a43667a <=( (not A300)  and  (not A299) );
 a43670a <=( (not A302)  and  (not A301) );
 a43671a <=( a43670a  and  a43667a );
 a43672a <=( a43671a  and  a43664a );
 a43676a <=( (not A167)  and  A168 );
 a43677a <=( (not A170)  and  a43676a );
 a43681a <=( A202  and  (not A201) );
 a43682a <=( A166  and  a43681a );
 a43683a <=( a43682a  and  a43677a );
 a43687a <=( (not A298)  and  A269 );
 a43688a <=( (not A267)  and  a43687a );
 a43691a <=( (not A300)  and  A299 );
 a43694a <=( (not A302)  and  (not A301) );
 a43695a <=( a43694a  and  a43691a );
 a43696a <=( a43695a  and  a43688a );
 a43700a <=( (not A167)  and  A168 );
 a43701a <=( (not A170)  and  a43700a );
 a43705a <=( A202  and  (not A201) );
 a43706a <=( A166  and  a43705a );
 a43707a <=( a43706a  and  a43701a );
 a43711a <=( A298  and  A266 );
 a43712a <=( A265  and  a43711a );
 a43715a <=( (not A300)  and  (not A299) );
 a43718a <=( (not A302)  and  (not A301) );
 a43719a <=( a43718a  and  a43715a );
 a43720a <=( a43719a  and  a43712a );
 a43724a <=( (not A167)  and  A168 );
 a43725a <=( (not A170)  and  a43724a );
 a43729a <=( A202  and  (not A201) );
 a43730a <=( A166  and  a43729a );
 a43731a <=( a43730a  and  a43725a );
 a43735a <=( (not A298)  and  A266 );
 a43736a <=( A265  and  a43735a );
 a43739a <=( (not A300)  and  A299 );
 a43742a <=( (not A302)  and  (not A301) );
 a43743a <=( a43742a  and  a43739a );
 a43744a <=( a43743a  and  a43736a );
 a43748a <=( (not A167)  and  A168 );
 a43749a <=( (not A170)  and  a43748a );
 a43753a <=( A202  and  (not A201) );
 a43754a <=( A166  and  a43753a );
 a43755a <=( a43754a  and  a43749a );
 a43759a <=( A298  and  (not A266) );
 a43760a <=( (not A265)  and  a43759a );
 a43763a <=( (not A300)  and  (not A299) );
 a43766a <=( (not A302)  and  (not A301) );
 a43767a <=( a43766a  and  a43763a );
 a43768a <=( a43767a  and  a43760a );
 a43772a <=( (not A167)  and  A168 );
 a43773a <=( (not A170)  and  a43772a );
 a43777a <=( A202  and  (not A201) );
 a43778a <=( A166  and  a43777a );
 a43779a <=( a43778a  and  a43773a );
 a43783a <=( (not A298)  and  (not A266) );
 a43784a <=( (not A265)  and  a43783a );
 a43787a <=( (not A300)  and  A299 );
 a43790a <=( (not A302)  and  (not A301) );
 a43791a <=( a43790a  and  a43787a );
 a43792a <=( a43791a  and  a43784a );
 a43796a <=( (not A167)  and  A168 );
 a43797a <=( (not A170)  and  a43796a );
 a43801a <=( A203  and  (not A201) );
 a43802a <=( A166  and  a43801a );
 a43803a <=( a43802a  and  a43797a );
 a43807a <=( (not A269)  and  (not A268) );
 a43808a <=( A267  and  a43807a );
 a43811a <=( (not A299)  and  A298 );
 a43814a <=( A301  and  A300 );
 a43815a <=( a43814a  and  a43811a );
 a43816a <=( a43815a  and  a43808a );
 a43820a <=( (not A167)  and  A168 );
 a43821a <=( (not A170)  and  a43820a );
 a43825a <=( A203  and  (not A201) );
 a43826a <=( A166  and  a43825a );
 a43827a <=( a43826a  and  a43821a );
 a43831a <=( (not A269)  and  (not A268) );
 a43832a <=( A267  and  a43831a );
 a43835a <=( (not A299)  and  A298 );
 a43838a <=( A302  and  A300 );
 a43839a <=( a43838a  and  a43835a );
 a43840a <=( a43839a  and  a43832a );
 a43844a <=( (not A167)  and  A168 );
 a43845a <=( (not A170)  and  a43844a );
 a43849a <=( A203  and  (not A201) );
 a43850a <=( A166  and  a43849a );
 a43851a <=( a43850a  and  a43845a );
 a43855a <=( (not A269)  and  (not A268) );
 a43856a <=( A267  and  a43855a );
 a43859a <=( A299  and  (not A298) );
 a43862a <=( A301  and  A300 );
 a43863a <=( a43862a  and  a43859a );
 a43864a <=( a43863a  and  a43856a );
 a43868a <=( (not A167)  and  A168 );
 a43869a <=( (not A170)  and  a43868a );
 a43873a <=( A203  and  (not A201) );
 a43874a <=( A166  and  a43873a );
 a43875a <=( a43874a  and  a43869a );
 a43879a <=( (not A269)  and  (not A268) );
 a43880a <=( A267  and  a43879a );
 a43883a <=( A299  and  (not A298) );
 a43886a <=( A302  and  A300 );
 a43887a <=( a43886a  and  a43883a );
 a43888a <=( a43887a  and  a43880a );
 a43892a <=( (not A167)  and  A168 );
 a43893a <=( (not A170)  and  a43892a );
 a43897a <=( A203  and  (not A201) );
 a43898a <=( A166  and  a43897a );
 a43899a <=( a43898a  and  a43893a );
 a43903a <=( A298  and  A268 );
 a43904a <=( (not A267)  and  a43903a );
 a43907a <=( (not A300)  and  (not A299) );
 a43910a <=( (not A302)  and  (not A301) );
 a43911a <=( a43910a  and  a43907a );
 a43912a <=( a43911a  and  a43904a );
 a43916a <=( (not A167)  and  A168 );
 a43917a <=( (not A170)  and  a43916a );
 a43921a <=( A203  and  (not A201) );
 a43922a <=( A166  and  a43921a );
 a43923a <=( a43922a  and  a43917a );
 a43927a <=( (not A298)  and  A268 );
 a43928a <=( (not A267)  and  a43927a );
 a43931a <=( (not A300)  and  A299 );
 a43934a <=( (not A302)  and  (not A301) );
 a43935a <=( a43934a  and  a43931a );
 a43936a <=( a43935a  and  a43928a );
 a43940a <=( (not A167)  and  A168 );
 a43941a <=( (not A170)  and  a43940a );
 a43945a <=( A203  and  (not A201) );
 a43946a <=( A166  and  a43945a );
 a43947a <=( a43946a  and  a43941a );
 a43951a <=( A298  and  A269 );
 a43952a <=( (not A267)  and  a43951a );
 a43955a <=( (not A300)  and  (not A299) );
 a43958a <=( (not A302)  and  (not A301) );
 a43959a <=( a43958a  and  a43955a );
 a43960a <=( a43959a  and  a43952a );
 a43964a <=( (not A167)  and  A168 );
 a43965a <=( (not A170)  and  a43964a );
 a43969a <=( A203  and  (not A201) );
 a43970a <=( A166  and  a43969a );
 a43971a <=( a43970a  and  a43965a );
 a43975a <=( (not A298)  and  A269 );
 a43976a <=( (not A267)  and  a43975a );
 a43979a <=( (not A300)  and  A299 );
 a43982a <=( (not A302)  and  (not A301) );
 a43983a <=( a43982a  and  a43979a );
 a43984a <=( a43983a  and  a43976a );
 a43988a <=( (not A167)  and  A168 );
 a43989a <=( (not A170)  and  a43988a );
 a43993a <=( A203  and  (not A201) );
 a43994a <=( A166  and  a43993a );
 a43995a <=( a43994a  and  a43989a );
 a43999a <=( A298  and  A266 );
 a44000a <=( A265  and  a43999a );
 a44003a <=( (not A300)  and  (not A299) );
 a44006a <=( (not A302)  and  (not A301) );
 a44007a <=( a44006a  and  a44003a );
 a44008a <=( a44007a  and  a44000a );
 a44012a <=( (not A167)  and  A168 );
 a44013a <=( (not A170)  and  a44012a );
 a44017a <=( A203  and  (not A201) );
 a44018a <=( A166  and  a44017a );
 a44019a <=( a44018a  and  a44013a );
 a44023a <=( (not A298)  and  A266 );
 a44024a <=( A265  and  a44023a );
 a44027a <=( (not A300)  and  A299 );
 a44030a <=( (not A302)  and  (not A301) );
 a44031a <=( a44030a  and  a44027a );
 a44032a <=( a44031a  and  a44024a );
 a44036a <=( (not A167)  and  A168 );
 a44037a <=( (not A170)  and  a44036a );
 a44041a <=( A203  and  (not A201) );
 a44042a <=( A166  and  a44041a );
 a44043a <=( a44042a  and  a44037a );
 a44047a <=( A298  and  (not A266) );
 a44048a <=( (not A265)  and  a44047a );
 a44051a <=( (not A300)  and  (not A299) );
 a44054a <=( (not A302)  and  (not A301) );
 a44055a <=( a44054a  and  a44051a );
 a44056a <=( a44055a  and  a44048a );
 a44060a <=( (not A167)  and  A168 );
 a44061a <=( (not A170)  and  a44060a );
 a44065a <=( A203  and  (not A201) );
 a44066a <=( A166  and  a44065a );
 a44067a <=( a44066a  and  a44061a );
 a44071a <=( (not A298)  and  (not A266) );
 a44072a <=( (not A265)  and  a44071a );
 a44075a <=( (not A300)  and  A299 );
 a44078a <=( (not A302)  and  (not A301) );
 a44079a <=( a44078a  and  a44075a );
 a44080a <=( a44079a  and  a44072a );
 a44084a <=( (not A167)  and  A168 );
 a44085a <=( (not A170)  and  a44084a );
 a44089a <=( A200  and  A199 );
 a44090a <=( A166  and  a44089a );
 a44091a <=( a44090a  and  a44085a );
 a44095a <=( (not A269)  and  (not A268) );
 a44096a <=( A267  and  a44095a );
 a44099a <=( (not A299)  and  A298 );
 a44102a <=( A301  and  A300 );
 a44103a <=( a44102a  and  a44099a );
 a44104a <=( a44103a  and  a44096a );
 a44108a <=( (not A167)  and  A168 );
 a44109a <=( (not A170)  and  a44108a );
 a44113a <=( A200  and  A199 );
 a44114a <=( A166  and  a44113a );
 a44115a <=( a44114a  and  a44109a );
 a44119a <=( (not A269)  and  (not A268) );
 a44120a <=( A267  and  a44119a );
 a44123a <=( (not A299)  and  A298 );
 a44126a <=( A302  and  A300 );
 a44127a <=( a44126a  and  a44123a );
 a44128a <=( a44127a  and  a44120a );
 a44132a <=( (not A167)  and  A168 );
 a44133a <=( (not A170)  and  a44132a );
 a44137a <=( A200  and  A199 );
 a44138a <=( A166  and  a44137a );
 a44139a <=( a44138a  and  a44133a );
 a44143a <=( (not A269)  and  (not A268) );
 a44144a <=( A267  and  a44143a );
 a44147a <=( A299  and  (not A298) );
 a44150a <=( A301  and  A300 );
 a44151a <=( a44150a  and  a44147a );
 a44152a <=( a44151a  and  a44144a );
 a44156a <=( (not A167)  and  A168 );
 a44157a <=( (not A170)  and  a44156a );
 a44161a <=( A200  and  A199 );
 a44162a <=( A166  and  a44161a );
 a44163a <=( a44162a  and  a44157a );
 a44167a <=( (not A269)  and  (not A268) );
 a44168a <=( A267  and  a44167a );
 a44171a <=( A299  and  (not A298) );
 a44174a <=( A302  and  A300 );
 a44175a <=( a44174a  and  a44171a );
 a44176a <=( a44175a  and  a44168a );
 a44180a <=( (not A167)  and  A168 );
 a44181a <=( (not A170)  and  a44180a );
 a44185a <=( A200  and  A199 );
 a44186a <=( A166  and  a44185a );
 a44187a <=( a44186a  and  a44181a );
 a44191a <=( A298  and  A268 );
 a44192a <=( (not A267)  and  a44191a );
 a44195a <=( (not A300)  and  (not A299) );
 a44198a <=( (not A302)  and  (not A301) );
 a44199a <=( a44198a  and  a44195a );
 a44200a <=( a44199a  and  a44192a );
 a44204a <=( (not A167)  and  A168 );
 a44205a <=( (not A170)  and  a44204a );
 a44209a <=( A200  and  A199 );
 a44210a <=( A166  and  a44209a );
 a44211a <=( a44210a  and  a44205a );
 a44215a <=( (not A298)  and  A268 );
 a44216a <=( (not A267)  and  a44215a );
 a44219a <=( (not A300)  and  A299 );
 a44222a <=( (not A302)  and  (not A301) );
 a44223a <=( a44222a  and  a44219a );
 a44224a <=( a44223a  and  a44216a );
 a44228a <=( (not A167)  and  A168 );
 a44229a <=( (not A170)  and  a44228a );
 a44233a <=( A200  and  A199 );
 a44234a <=( A166  and  a44233a );
 a44235a <=( a44234a  and  a44229a );
 a44239a <=( A298  and  A269 );
 a44240a <=( (not A267)  and  a44239a );
 a44243a <=( (not A300)  and  (not A299) );
 a44246a <=( (not A302)  and  (not A301) );
 a44247a <=( a44246a  and  a44243a );
 a44248a <=( a44247a  and  a44240a );
 a44252a <=( (not A167)  and  A168 );
 a44253a <=( (not A170)  and  a44252a );
 a44257a <=( A200  and  A199 );
 a44258a <=( A166  and  a44257a );
 a44259a <=( a44258a  and  a44253a );
 a44263a <=( (not A298)  and  A269 );
 a44264a <=( (not A267)  and  a44263a );
 a44267a <=( (not A300)  and  A299 );
 a44270a <=( (not A302)  and  (not A301) );
 a44271a <=( a44270a  and  a44267a );
 a44272a <=( a44271a  and  a44264a );
 a44276a <=( (not A167)  and  A168 );
 a44277a <=( (not A170)  and  a44276a );
 a44281a <=( A200  and  A199 );
 a44282a <=( A166  and  a44281a );
 a44283a <=( a44282a  and  a44277a );
 a44287a <=( A298  and  A266 );
 a44288a <=( A265  and  a44287a );
 a44291a <=( (not A300)  and  (not A299) );
 a44294a <=( (not A302)  and  (not A301) );
 a44295a <=( a44294a  and  a44291a );
 a44296a <=( a44295a  and  a44288a );
 a44300a <=( (not A167)  and  A168 );
 a44301a <=( (not A170)  and  a44300a );
 a44305a <=( A200  and  A199 );
 a44306a <=( A166  and  a44305a );
 a44307a <=( a44306a  and  a44301a );
 a44311a <=( (not A298)  and  A266 );
 a44312a <=( A265  and  a44311a );
 a44315a <=( (not A300)  and  A299 );
 a44318a <=( (not A302)  and  (not A301) );
 a44319a <=( a44318a  and  a44315a );
 a44320a <=( a44319a  and  a44312a );
 a44324a <=( (not A167)  and  A168 );
 a44325a <=( (not A170)  and  a44324a );
 a44329a <=( A200  and  A199 );
 a44330a <=( A166  and  a44329a );
 a44331a <=( a44330a  and  a44325a );
 a44335a <=( A298  and  (not A266) );
 a44336a <=( (not A265)  and  a44335a );
 a44339a <=( (not A300)  and  (not A299) );
 a44342a <=( (not A302)  and  (not A301) );
 a44343a <=( a44342a  and  a44339a );
 a44344a <=( a44343a  and  a44336a );
 a44348a <=( (not A167)  and  A168 );
 a44349a <=( (not A170)  and  a44348a );
 a44353a <=( A200  and  A199 );
 a44354a <=( A166  and  a44353a );
 a44355a <=( a44354a  and  a44349a );
 a44359a <=( (not A298)  and  (not A266) );
 a44360a <=( (not A265)  and  a44359a );
 a44363a <=( (not A300)  and  A299 );
 a44366a <=( (not A302)  and  (not A301) );
 a44367a <=( a44366a  and  a44363a );
 a44368a <=( a44367a  and  a44360a );
 a44372a <=( (not A167)  and  A168 );
 a44373a <=( (not A170)  and  a44372a );
 a44377a <=( (not A200)  and  (not A199) );
 a44378a <=( A166  and  a44377a );
 a44379a <=( a44378a  and  a44373a );
 a44383a <=( (not A269)  and  (not A268) );
 a44384a <=( A267  and  a44383a );
 a44387a <=( (not A299)  and  A298 );
 a44390a <=( A301  and  A300 );
 a44391a <=( a44390a  and  a44387a );
 a44392a <=( a44391a  and  a44384a );
 a44396a <=( (not A167)  and  A168 );
 a44397a <=( (not A170)  and  a44396a );
 a44401a <=( (not A200)  and  (not A199) );
 a44402a <=( A166  and  a44401a );
 a44403a <=( a44402a  and  a44397a );
 a44407a <=( (not A269)  and  (not A268) );
 a44408a <=( A267  and  a44407a );
 a44411a <=( (not A299)  and  A298 );
 a44414a <=( A302  and  A300 );
 a44415a <=( a44414a  and  a44411a );
 a44416a <=( a44415a  and  a44408a );
 a44420a <=( (not A167)  and  A168 );
 a44421a <=( (not A170)  and  a44420a );
 a44425a <=( (not A200)  and  (not A199) );
 a44426a <=( A166  and  a44425a );
 a44427a <=( a44426a  and  a44421a );
 a44431a <=( (not A269)  and  (not A268) );
 a44432a <=( A267  and  a44431a );
 a44435a <=( A299  and  (not A298) );
 a44438a <=( A301  and  A300 );
 a44439a <=( a44438a  and  a44435a );
 a44440a <=( a44439a  and  a44432a );
 a44444a <=( (not A167)  and  A168 );
 a44445a <=( (not A170)  and  a44444a );
 a44449a <=( (not A200)  and  (not A199) );
 a44450a <=( A166  and  a44449a );
 a44451a <=( a44450a  and  a44445a );
 a44455a <=( (not A269)  and  (not A268) );
 a44456a <=( A267  and  a44455a );
 a44459a <=( A299  and  (not A298) );
 a44462a <=( A302  and  A300 );
 a44463a <=( a44462a  and  a44459a );
 a44464a <=( a44463a  and  a44456a );
 a44468a <=( (not A167)  and  A168 );
 a44469a <=( (not A170)  and  a44468a );
 a44473a <=( (not A200)  and  (not A199) );
 a44474a <=( A166  and  a44473a );
 a44475a <=( a44474a  and  a44469a );
 a44479a <=( A298  and  A268 );
 a44480a <=( (not A267)  and  a44479a );
 a44483a <=( (not A300)  and  (not A299) );
 a44486a <=( (not A302)  and  (not A301) );
 a44487a <=( a44486a  and  a44483a );
 a44488a <=( a44487a  and  a44480a );
 a44492a <=( (not A167)  and  A168 );
 a44493a <=( (not A170)  and  a44492a );
 a44497a <=( (not A200)  and  (not A199) );
 a44498a <=( A166  and  a44497a );
 a44499a <=( a44498a  and  a44493a );
 a44503a <=( (not A298)  and  A268 );
 a44504a <=( (not A267)  and  a44503a );
 a44507a <=( (not A300)  and  A299 );
 a44510a <=( (not A302)  and  (not A301) );
 a44511a <=( a44510a  and  a44507a );
 a44512a <=( a44511a  and  a44504a );
 a44516a <=( (not A167)  and  A168 );
 a44517a <=( (not A170)  and  a44516a );
 a44521a <=( (not A200)  and  (not A199) );
 a44522a <=( A166  and  a44521a );
 a44523a <=( a44522a  and  a44517a );
 a44527a <=( A298  and  A269 );
 a44528a <=( (not A267)  and  a44527a );
 a44531a <=( (not A300)  and  (not A299) );
 a44534a <=( (not A302)  and  (not A301) );
 a44535a <=( a44534a  and  a44531a );
 a44536a <=( a44535a  and  a44528a );
 a44540a <=( (not A167)  and  A168 );
 a44541a <=( (not A170)  and  a44540a );
 a44545a <=( (not A200)  and  (not A199) );
 a44546a <=( A166  and  a44545a );
 a44547a <=( a44546a  and  a44541a );
 a44551a <=( (not A298)  and  A269 );
 a44552a <=( (not A267)  and  a44551a );
 a44555a <=( (not A300)  and  A299 );
 a44558a <=( (not A302)  and  (not A301) );
 a44559a <=( a44558a  and  a44555a );
 a44560a <=( a44559a  and  a44552a );
 a44564a <=( (not A167)  and  A168 );
 a44565a <=( (not A170)  and  a44564a );
 a44569a <=( (not A200)  and  (not A199) );
 a44570a <=( A166  and  a44569a );
 a44571a <=( a44570a  and  a44565a );
 a44575a <=( A298  and  A266 );
 a44576a <=( A265  and  a44575a );
 a44579a <=( (not A300)  and  (not A299) );
 a44582a <=( (not A302)  and  (not A301) );
 a44583a <=( a44582a  and  a44579a );
 a44584a <=( a44583a  and  a44576a );
 a44588a <=( (not A167)  and  A168 );
 a44589a <=( (not A170)  and  a44588a );
 a44593a <=( (not A200)  and  (not A199) );
 a44594a <=( A166  and  a44593a );
 a44595a <=( a44594a  and  a44589a );
 a44599a <=( (not A298)  and  A266 );
 a44600a <=( A265  and  a44599a );
 a44603a <=( (not A300)  and  A299 );
 a44606a <=( (not A302)  and  (not A301) );
 a44607a <=( a44606a  and  a44603a );
 a44608a <=( a44607a  and  a44600a );
 a44612a <=( (not A167)  and  A168 );
 a44613a <=( (not A170)  and  a44612a );
 a44617a <=( (not A200)  and  (not A199) );
 a44618a <=( A166  and  a44617a );
 a44619a <=( a44618a  and  a44613a );
 a44623a <=( A298  and  (not A266) );
 a44624a <=( (not A265)  and  a44623a );
 a44627a <=( (not A300)  and  (not A299) );
 a44630a <=( (not A302)  and  (not A301) );
 a44631a <=( a44630a  and  a44627a );
 a44632a <=( a44631a  and  a44624a );
 a44636a <=( (not A167)  and  A168 );
 a44637a <=( (not A170)  and  a44636a );
 a44641a <=( (not A200)  and  (not A199) );
 a44642a <=( A166  and  a44641a );
 a44643a <=( a44642a  and  a44637a );
 a44647a <=( (not A298)  and  (not A266) );
 a44648a <=( (not A265)  and  a44647a );
 a44651a <=( (not A300)  and  A299 );
 a44654a <=( (not A302)  and  (not A301) );
 a44655a <=( a44654a  and  a44651a );
 a44656a <=( a44655a  and  a44648a );
 a44660a <=( A201  and  (not A168) );
 a44661a <=( (not A170)  and  a44660a );
 a44665a <=( (not A265)  and  (not A203) );
 a44666a <=( (not A202)  and  a44665a );
 a44667a <=( a44666a  and  a44661a );
 a44671a <=( (not A268)  and  (not A267) );
 a44672a <=( A266  and  a44671a );
 a44675a <=( A300  and  (not A269) );
 a44678a <=( (not A302)  and  (not A301) );
 a44679a <=( a44678a  and  a44675a );
 a44680a <=( a44679a  and  a44672a );
 a44684a <=( A201  and  (not A168) );
 a44685a <=( (not A170)  and  a44684a );
 a44689a <=( A265  and  (not A203) );
 a44690a <=( (not A202)  and  a44689a );
 a44691a <=( a44690a  and  a44685a );
 a44695a <=( (not A268)  and  (not A267) );
 a44696a <=( (not A266)  and  a44695a );
 a44699a <=( A300  and  (not A269) );
 a44702a <=( (not A302)  and  (not A301) );
 a44703a <=( a44702a  and  a44699a );
 a44704a <=( a44703a  and  a44696a );
 a44708a <=( (not A199)  and  (not A168) );
 a44709a <=( (not A170)  and  a44708a );
 a44713a <=( A202  and  A201 );
 a44714a <=( A200  and  a44713a );
 a44715a <=( a44714a  and  a44709a );
 a44719a <=( (not A269)  and  (not A268) );
 a44720a <=( A267  and  a44719a );
 a44723a <=( (not A299)  and  A298 );
 a44726a <=( A301  and  A300 );
 a44727a <=( a44726a  and  a44723a );
 a44728a <=( a44727a  and  a44720a );
 a44732a <=( (not A199)  and  (not A168) );
 a44733a <=( (not A170)  and  a44732a );
 a44737a <=( A202  and  A201 );
 a44738a <=( A200  and  a44737a );
 a44739a <=( a44738a  and  a44733a );
 a44743a <=( (not A269)  and  (not A268) );
 a44744a <=( A267  and  a44743a );
 a44747a <=( (not A299)  and  A298 );
 a44750a <=( A302  and  A300 );
 a44751a <=( a44750a  and  a44747a );
 a44752a <=( a44751a  and  a44744a );
 a44756a <=( (not A199)  and  (not A168) );
 a44757a <=( (not A170)  and  a44756a );
 a44761a <=( A202  and  A201 );
 a44762a <=( A200  and  a44761a );
 a44763a <=( a44762a  and  a44757a );
 a44767a <=( (not A269)  and  (not A268) );
 a44768a <=( A267  and  a44767a );
 a44771a <=( A299  and  (not A298) );
 a44774a <=( A301  and  A300 );
 a44775a <=( a44774a  and  a44771a );
 a44776a <=( a44775a  and  a44768a );
 a44780a <=( (not A199)  and  (not A168) );
 a44781a <=( (not A170)  and  a44780a );
 a44785a <=( A202  and  A201 );
 a44786a <=( A200  and  a44785a );
 a44787a <=( a44786a  and  a44781a );
 a44791a <=( (not A269)  and  (not A268) );
 a44792a <=( A267  and  a44791a );
 a44795a <=( A299  and  (not A298) );
 a44798a <=( A302  and  A300 );
 a44799a <=( a44798a  and  a44795a );
 a44800a <=( a44799a  and  a44792a );
 a44804a <=( (not A199)  and  (not A168) );
 a44805a <=( (not A170)  and  a44804a );
 a44809a <=( A202  and  A201 );
 a44810a <=( A200  and  a44809a );
 a44811a <=( a44810a  and  a44805a );
 a44815a <=( A298  and  A268 );
 a44816a <=( (not A267)  and  a44815a );
 a44819a <=( (not A300)  and  (not A299) );
 a44822a <=( (not A302)  and  (not A301) );
 a44823a <=( a44822a  and  a44819a );
 a44824a <=( a44823a  and  a44816a );
 a44828a <=( (not A199)  and  (not A168) );
 a44829a <=( (not A170)  and  a44828a );
 a44833a <=( A202  and  A201 );
 a44834a <=( A200  and  a44833a );
 a44835a <=( a44834a  and  a44829a );
 a44839a <=( (not A298)  and  A268 );
 a44840a <=( (not A267)  and  a44839a );
 a44843a <=( (not A300)  and  A299 );
 a44846a <=( (not A302)  and  (not A301) );
 a44847a <=( a44846a  and  a44843a );
 a44848a <=( a44847a  and  a44840a );
 a44852a <=( (not A199)  and  (not A168) );
 a44853a <=( (not A170)  and  a44852a );
 a44857a <=( A202  and  A201 );
 a44858a <=( A200  and  a44857a );
 a44859a <=( a44858a  and  a44853a );
 a44863a <=( A298  and  A269 );
 a44864a <=( (not A267)  and  a44863a );
 a44867a <=( (not A300)  and  (not A299) );
 a44870a <=( (not A302)  and  (not A301) );
 a44871a <=( a44870a  and  a44867a );
 a44872a <=( a44871a  and  a44864a );
 a44876a <=( (not A199)  and  (not A168) );
 a44877a <=( (not A170)  and  a44876a );
 a44881a <=( A202  and  A201 );
 a44882a <=( A200  and  a44881a );
 a44883a <=( a44882a  and  a44877a );
 a44887a <=( (not A298)  and  A269 );
 a44888a <=( (not A267)  and  a44887a );
 a44891a <=( (not A300)  and  A299 );
 a44894a <=( (not A302)  and  (not A301) );
 a44895a <=( a44894a  and  a44891a );
 a44896a <=( a44895a  and  a44888a );
 a44900a <=( (not A199)  and  (not A168) );
 a44901a <=( (not A170)  and  a44900a );
 a44905a <=( A202  and  A201 );
 a44906a <=( A200  and  a44905a );
 a44907a <=( a44906a  and  a44901a );
 a44911a <=( A298  and  A266 );
 a44912a <=( A265  and  a44911a );
 a44915a <=( (not A300)  and  (not A299) );
 a44918a <=( (not A302)  and  (not A301) );
 a44919a <=( a44918a  and  a44915a );
 a44920a <=( a44919a  and  a44912a );
 a44924a <=( (not A199)  and  (not A168) );
 a44925a <=( (not A170)  and  a44924a );
 a44929a <=( A202  and  A201 );
 a44930a <=( A200  and  a44929a );
 a44931a <=( a44930a  and  a44925a );
 a44935a <=( (not A298)  and  A266 );
 a44936a <=( A265  and  a44935a );
 a44939a <=( (not A300)  and  A299 );
 a44942a <=( (not A302)  and  (not A301) );
 a44943a <=( a44942a  and  a44939a );
 a44944a <=( a44943a  and  a44936a );
 a44948a <=( (not A199)  and  (not A168) );
 a44949a <=( (not A170)  and  a44948a );
 a44953a <=( A202  and  A201 );
 a44954a <=( A200  and  a44953a );
 a44955a <=( a44954a  and  a44949a );
 a44959a <=( A298  and  (not A266) );
 a44960a <=( (not A265)  and  a44959a );
 a44963a <=( (not A300)  and  (not A299) );
 a44966a <=( (not A302)  and  (not A301) );
 a44967a <=( a44966a  and  a44963a );
 a44968a <=( a44967a  and  a44960a );
 a44972a <=( (not A199)  and  (not A168) );
 a44973a <=( (not A170)  and  a44972a );
 a44977a <=( A202  and  A201 );
 a44978a <=( A200  and  a44977a );
 a44979a <=( a44978a  and  a44973a );
 a44983a <=( (not A298)  and  (not A266) );
 a44984a <=( (not A265)  and  a44983a );
 a44987a <=( (not A300)  and  A299 );
 a44990a <=( (not A302)  and  (not A301) );
 a44991a <=( a44990a  and  a44987a );
 a44992a <=( a44991a  and  a44984a );
 a44996a <=( (not A199)  and  (not A168) );
 a44997a <=( (not A170)  and  a44996a );
 a45001a <=( A203  and  A201 );
 a45002a <=( A200  and  a45001a );
 a45003a <=( a45002a  and  a44997a );
 a45007a <=( (not A269)  and  (not A268) );
 a45008a <=( A267  and  a45007a );
 a45011a <=( (not A299)  and  A298 );
 a45014a <=( A301  and  A300 );
 a45015a <=( a45014a  and  a45011a );
 a45016a <=( a45015a  and  a45008a );
 a45020a <=( (not A199)  and  (not A168) );
 a45021a <=( (not A170)  and  a45020a );
 a45025a <=( A203  and  A201 );
 a45026a <=( A200  and  a45025a );
 a45027a <=( a45026a  and  a45021a );
 a45031a <=( (not A269)  and  (not A268) );
 a45032a <=( A267  and  a45031a );
 a45035a <=( (not A299)  and  A298 );
 a45038a <=( A302  and  A300 );
 a45039a <=( a45038a  and  a45035a );
 a45040a <=( a45039a  and  a45032a );
 a45044a <=( (not A199)  and  (not A168) );
 a45045a <=( (not A170)  and  a45044a );
 a45049a <=( A203  and  A201 );
 a45050a <=( A200  and  a45049a );
 a45051a <=( a45050a  and  a45045a );
 a45055a <=( (not A269)  and  (not A268) );
 a45056a <=( A267  and  a45055a );
 a45059a <=( A299  and  (not A298) );
 a45062a <=( A301  and  A300 );
 a45063a <=( a45062a  and  a45059a );
 a45064a <=( a45063a  and  a45056a );
 a45068a <=( (not A199)  and  (not A168) );
 a45069a <=( (not A170)  and  a45068a );
 a45073a <=( A203  and  A201 );
 a45074a <=( A200  and  a45073a );
 a45075a <=( a45074a  and  a45069a );
 a45079a <=( (not A269)  and  (not A268) );
 a45080a <=( A267  and  a45079a );
 a45083a <=( A299  and  (not A298) );
 a45086a <=( A302  and  A300 );
 a45087a <=( a45086a  and  a45083a );
 a45088a <=( a45087a  and  a45080a );
 a45092a <=( (not A199)  and  (not A168) );
 a45093a <=( (not A170)  and  a45092a );
 a45097a <=( A203  and  A201 );
 a45098a <=( A200  and  a45097a );
 a45099a <=( a45098a  and  a45093a );
 a45103a <=( A298  and  A268 );
 a45104a <=( (not A267)  and  a45103a );
 a45107a <=( (not A300)  and  (not A299) );
 a45110a <=( (not A302)  and  (not A301) );
 a45111a <=( a45110a  and  a45107a );
 a45112a <=( a45111a  and  a45104a );
 a45116a <=( (not A199)  and  (not A168) );
 a45117a <=( (not A170)  and  a45116a );
 a45121a <=( A203  and  A201 );
 a45122a <=( A200  and  a45121a );
 a45123a <=( a45122a  and  a45117a );
 a45127a <=( (not A298)  and  A268 );
 a45128a <=( (not A267)  and  a45127a );
 a45131a <=( (not A300)  and  A299 );
 a45134a <=( (not A302)  and  (not A301) );
 a45135a <=( a45134a  and  a45131a );
 a45136a <=( a45135a  and  a45128a );
 a45140a <=( (not A199)  and  (not A168) );
 a45141a <=( (not A170)  and  a45140a );
 a45145a <=( A203  and  A201 );
 a45146a <=( A200  and  a45145a );
 a45147a <=( a45146a  and  a45141a );
 a45151a <=( A298  and  A269 );
 a45152a <=( (not A267)  and  a45151a );
 a45155a <=( (not A300)  and  (not A299) );
 a45158a <=( (not A302)  and  (not A301) );
 a45159a <=( a45158a  and  a45155a );
 a45160a <=( a45159a  and  a45152a );
 a45164a <=( (not A199)  and  (not A168) );
 a45165a <=( (not A170)  and  a45164a );
 a45169a <=( A203  and  A201 );
 a45170a <=( A200  and  a45169a );
 a45171a <=( a45170a  and  a45165a );
 a45175a <=( (not A298)  and  A269 );
 a45176a <=( (not A267)  and  a45175a );
 a45179a <=( (not A300)  and  A299 );
 a45182a <=( (not A302)  and  (not A301) );
 a45183a <=( a45182a  and  a45179a );
 a45184a <=( a45183a  and  a45176a );
 a45188a <=( (not A199)  and  (not A168) );
 a45189a <=( (not A170)  and  a45188a );
 a45193a <=( A203  and  A201 );
 a45194a <=( A200  and  a45193a );
 a45195a <=( a45194a  and  a45189a );
 a45199a <=( A298  and  A266 );
 a45200a <=( A265  and  a45199a );
 a45203a <=( (not A300)  and  (not A299) );
 a45206a <=( (not A302)  and  (not A301) );
 a45207a <=( a45206a  and  a45203a );
 a45208a <=( a45207a  and  a45200a );
 a45212a <=( (not A199)  and  (not A168) );
 a45213a <=( (not A170)  and  a45212a );
 a45217a <=( A203  and  A201 );
 a45218a <=( A200  and  a45217a );
 a45219a <=( a45218a  and  a45213a );
 a45223a <=( (not A298)  and  A266 );
 a45224a <=( A265  and  a45223a );
 a45227a <=( (not A300)  and  A299 );
 a45230a <=( (not A302)  and  (not A301) );
 a45231a <=( a45230a  and  a45227a );
 a45232a <=( a45231a  and  a45224a );
 a45236a <=( (not A199)  and  (not A168) );
 a45237a <=( (not A170)  and  a45236a );
 a45241a <=( A203  and  A201 );
 a45242a <=( A200  and  a45241a );
 a45243a <=( a45242a  and  a45237a );
 a45247a <=( A298  and  (not A266) );
 a45248a <=( (not A265)  and  a45247a );
 a45251a <=( (not A300)  and  (not A299) );
 a45254a <=( (not A302)  and  (not A301) );
 a45255a <=( a45254a  and  a45251a );
 a45256a <=( a45255a  and  a45248a );
 a45260a <=( (not A199)  and  (not A168) );
 a45261a <=( (not A170)  and  a45260a );
 a45265a <=( A203  and  A201 );
 a45266a <=( A200  and  a45265a );
 a45267a <=( a45266a  and  a45261a );
 a45271a <=( (not A298)  and  (not A266) );
 a45272a <=( (not A265)  and  a45271a );
 a45275a <=( (not A300)  and  A299 );
 a45278a <=( (not A302)  and  (not A301) );
 a45279a <=( a45278a  and  a45275a );
 a45280a <=( a45279a  and  a45272a );
 a45284a <=( (not A199)  and  (not A168) );
 a45285a <=( (not A170)  and  a45284a );
 a45289a <=( (not A202)  and  (not A201) );
 a45290a <=( A200  and  a45289a );
 a45291a <=( a45290a  and  a45285a );
 a45295a <=( A268  and  (not A267) );
 a45296a <=( (not A203)  and  a45295a );
 a45299a <=( (not A299)  and  A298 );
 a45302a <=( A301  and  A300 );
 a45303a <=( a45302a  and  a45299a );
 a45304a <=( a45303a  and  a45296a );
 a45308a <=( (not A199)  and  (not A168) );
 a45309a <=( (not A170)  and  a45308a );
 a45313a <=( (not A202)  and  (not A201) );
 a45314a <=( A200  and  a45313a );
 a45315a <=( a45314a  and  a45309a );
 a45319a <=( A268  and  (not A267) );
 a45320a <=( (not A203)  and  a45319a );
 a45323a <=( (not A299)  and  A298 );
 a45326a <=( A302  and  A300 );
 a45327a <=( a45326a  and  a45323a );
 a45328a <=( a45327a  and  a45320a );
 a45332a <=( (not A199)  and  (not A168) );
 a45333a <=( (not A170)  and  a45332a );
 a45337a <=( (not A202)  and  (not A201) );
 a45338a <=( A200  and  a45337a );
 a45339a <=( a45338a  and  a45333a );
 a45343a <=( A268  and  (not A267) );
 a45344a <=( (not A203)  and  a45343a );
 a45347a <=( A299  and  (not A298) );
 a45350a <=( A301  and  A300 );
 a45351a <=( a45350a  and  a45347a );
 a45352a <=( a45351a  and  a45344a );
 a45356a <=( (not A199)  and  (not A168) );
 a45357a <=( (not A170)  and  a45356a );
 a45361a <=( (not A202)  and  (not A201) );
 a45362a <=( A200  and  a45361a );
 a45363a <=( a45362a  and  a45357a );
 a45367a <=( A268  and  (not A267) );
 a45368a <=( (not A203)  and  a45367a );
 a45371a <=( A299  and  (not A298) );
 a45374a <=( A302  and  A300 );
 a45375a <=( a45374a  and  a45371a );
 a45376a <=( a45375a  and  a45368a );
 a45380a <=( (not A199)  and  (not A168) );
 a45381a <=( (not A170)  and  a45380a );
 a45385a <=( (not A202)  and  (not A201) );
 a45386a <=( A200  and  a45385a );
 a45387a <=( a45386a  and  a45381a );
 a45391a <=( A269  and  (not A267) );
 a45392a <=( (not A203)  and  a45391a );
 a45395a <=( (not A299)  and  A298 );
 a45398a <=( A301  and  A300 );
 a45399a <=( a45398a  and  a45395a );
 a45400a <=( a45399a  and  a45392a );
 a45404a <=( (not A199)  and  (not A168) );
 a45405a <=( (not A170)  and  a45404a );
 a45409a <=( (not A202)  and  (not A201) );
 a45410a <=( A200  and  a45409a );
 a45411a <=( a45410a  and  a45405a );
 a45415a <=( A269  and  (not A267) );
 a45416a <=( (not A203)  and  a45415a );
 a45419a <=( (not A299)  and  A298 );
 a45422a <=( A302  and  A300 );
 a45423a <=( a45422a  and  a45419a );
 a45424a <=( a45423a  and  a45416a );
 a45428a <=( (not A199)  and  (not A168) );
 a45429a <=( (not A170)  and  a45428a );
 a45433a <=( (not A202)  and  (not A201) );
 a45434a <=( A200  and  a45433a );
 a45435a <=( a45434a  and  a45429a );
 a45439a <=( A269  and  (not A267) );
 a45440a <=( (not A203)  and  a45439a );
 a45443a <=( A299  and  (not A298) );
 a45446a <=( A301  and  A300 );
 a45447a <=( a45446a  and  a45443a );
 a45448a <=( a45447a  and  a45440a );
 a45452a <=( (not A199)  and  (not A168) );
 a45453a <=( (not A170)  and  a45452a );
 a45457a <=( (not A202)  and  (not A201) );
 a45458a <=( A200  and  a45457a );
 a45459a <=( a45458a  and  a45453a );
 a45463a <=( A269  and  (not A267) );
 a45464a <=( (not A203)  and  a45463a );
 a45467a <=( A299  and  (not A298) );
 a45470a <=( A302  and  A300 );
 a45471a <=( a45470a  and  a45467a );
 a45472a <=( a45471a  and  a45464a );
 a45476a <=( (not A199)  and  (not A168) );
 a45477a <=( (not A170)  and  a45476a );
 a45481a <=( (not A202)  and  (not A201) );
 a45482a <=( A200  and  a45481a );
 a45483a <=( a45482a  and  a45477a );
 a45487a <=( A266  and  A265 );
 a45488a <=( (not A203)  and  a45487a );
 a45491a <=( (not A299)  and  A298 );
 a45494a <=( A301  and  A300 );
 a45495a <=( a45494a  and  a45491a );
 a45496a <=( a45495a  and  a45488a );
 a45500a <=( (not A199)  and  (not A168) );
 a45501a <=( (not A170)  and  a45500a );
 a45505a <=( (not A202)  and  (not A201) );
 a45506a <=( A200  and  a45505a );
 a45507a <=( a45506a  and  a45501a );
 a45511a <=( A266  and  A265 );
 a45512a <=( (not A203)  and  a45511a );
 a45515a <=( (not A299)  and  A298 );
 a45518a <=( A302  and  A300 );
 a45519a <=( a45518a  and  a45515a );
 a45520a <=( a45519a  and  a45512a );
 a45524a <=( (not A199)  and  (not A168) );
 a45525a <=( (not A170)  and  a45524a );
 a45529a <=( (not A202)  and  (not A201) );
 a45530a <=( A200  and  a45529a );
 a45531a <=( a45530a  and  a45525a );
 a45535a <=( A266  and  A265 );
 a45536a <=( (not A203)  and  a45535a );
 a45539a <=( A299  and  (not A298) );
 a45542a <=( A301  and  A300 );
 a45543a <=( a45542a  and  a45539a );
 a45544a <=( a45543a  and  a45536a );
 a45548a <=( (not A199)  and  (not A168) );
 a45549a <=( (not A170)  and  a45548a );
 a45553a <=( (not A202)  and  (not A201) );
 a45554a <=( A200  and  a45553a );
 a45555a <=( a45554a  and  a45549a );
 a45559a <=( A266  and  A265 );
 a45560a <=( (not A203)  and  a45559a );
 a45563a <=( A299  and  (not A298) );
 a45566a <=( A302  and  A300 );
 a45567a <=( a45566a  and  a45563a );
 a45568a <=( a45567a  and  a45560a );
 a45572a <=( (not A199)  and  (not A168) );
 a45573a <=( (not A170)  and  a45572a );
 a45577a <=( (not A202)  and  (not A201) );
 a45578a <=( A200  and  a45577a );
 a45579a <=( a45578a  and  a45573a );
 a45583a <=( (not A266)  and  (not A265) );
 a45584a <=( (not A203)  and  a45583a );
 a45587a <=( (not A299)  and  A298 );
 a45590a <=( A301  and  A300 );
 a45591a <=( a45590a  and  a45587a );
 a45592a <=( a45591a  and  a45584a );
 a45596a <=( (not A199)  and  (not A168) );
 a45597a <=( (not A170)  and  a45596a );
 a45601a <=( (not A202)  and  (not A201) );
 a45602a <=( A200  and  a45601a );
 a45603a <=( a45602a  and  a45597a );
 a45607a <=( (not A266)  and  (not A265) );
 a45608a <=( (not A203)  and  a45607a );
 a45611a <=( (not A299)  and  A298 );
 a45614a <=( A302  and  A300 );
 a45615a <=( a45614a  and  a45611a );
 a45616a <=( a45615a  and  a45608a );
 a45620a <=( (not A199)  and  (not A168) );
 a45621a <=( (not A170)  and  a45620a );
 a45625a <=( (not A202)  and  (not A201) );
 a45626a <=( A200  and  a45625a );
 a45627a <=( a45626a  and  a45621a );
 a45631a <=( (not A266)  and  (not A265) );
 a45632a <=( (not A203)  and  a45631a );
 a45635a <=( A299  and  (not A298) );
 a45638a <=( A301  and  A300 );
 a45639a <=( a45638a  and  a45635a );
 a45640a <=( a45639a  and  a45632a );
 a45644a <=( (not A199)  and  (not A168) );
 a45645a <=( (not A170)  and  a45644a );
 a45649a <=( (not A202)  and  (not A201) );
 a45650a <=( A200  and  a45649a );
 a45651a <=( a45650a  and  a45645a );
 a45655a <=( (not A266)  and  (not A265) );
 a45656a <=( (not A203)  and  a45655a );
 a45659a <=( A299  and  (not A298) );
 a45662a <=( A302  and  A300 );
 a45663a <=( a45662a  and  a45659a );
 a45664a <=( a45663a  and  a45656a );
 a45668a <=( A199  and  (not A168) );
 a45669a <=( (not A170)  and  a45668a );
 a45673a <=( A202  and  A201 );
 a45674a <=( (not A200)  and  a45673a );
 a45675a <=( a45674a  and  a45669a );
 a45679a <=( (not A269)  and  (not A268) );
 a45680a <=( A267  and  a45679a );
 a45683a <=( (not A299)  and  A298 );
 a45686a <=( A301  and  A300 );
 a45687a <=( a45686a  and  a45683a );
 a45688a <=( a45687a  and  a45680a );
 a45692a <=( A199  and  (not A168) );
 a45693a <=( (not A170)  and  a45692a );
 a45697a <=( A202  and  A201 );
 a45698a <=( (not A200)  and  a45697a );
 a45699a <=( a45698a  and  a45693a );
 a45703a <=( (not A269)  and  (not A268) );
 a45704a <=( A267  and  a45703a );
 a45707a <=( (not A299)  and  A298 );
 a45710a <=( A302  and  A300 );
 a45711a <=( a45710a  and  a45707a );
 a45712a <=( a45711a  and  a45704a );
 a45716a <=( A199  and  (not A168) );
 a45717a <=( (not A170)  and  a45716a );
 a45721a <=( A202  and  A201 );
 a45722a <=( (not A200)  and  a45721a );
 a45723a <=( a45722a  and  a45717a );
 a45727a <=( (not A269)  and  (not A268) );
 a45728a <=( A267  and  a45727a );
 a45731a <=( A299  and  (not A298) );
 a45734a <=( A301  and  A300 );
 a45735a <=( a45734a  and  a45731a );
 a45736a <=( a45735a  and  a45728a );
 a45740a <=( A199  and  (not A168) );
 a45741a <=( (not A170)  and  a45740a );
 a45745a <=( A202  and  A201 );
 a45746a <=( (not A200)  and  a45745a );
 a45747a <=( a45746a  and  a45741a );
 a45751a <=( (not A269)  and  (not A268) );
 a45752a <=( A267  and  a45751a );
 a45755a <=( A299  and  (not A298) );
 a45758a <=( A302  and  A300 );
 a45759a <=( a45758a  and  a45755a );
 a45760a <=( a45759a  and  a45752a );
 a45764a <=( A199  and  (not A168) );
 a45765a <=( (not A170)  and  a45764a );
 a45769a <=( A202  and  A201 );
 a45770a <=( (not A200)  and  a45769a );
 a45771a <=( a45770a  and  a45765a );
 a45775a <=( A298  and  A268 );
 a45776a <=( (not A267)  and  a45775a );
 a45779a <=( (not A300)  and  (not A299) );
 a45782a <=( (not A302)  and  (not A301) );
 a45783a <=( a45782a  and  a45779a );
 a45784a <=( a45783a  and  a45776a );
 a45788a <=( A199  and  (not A168) );
 a45789a <=( (not A170)  and  a45788a );
 a45793a <=( A202  and  A201 );
 a45794a <=( (not A200)  and  a45793a );
 a45795a <=( a45794a  and  a45789a );
 a45799a <=( (not A298)  and  A268 );
 a45800a <=( (not A267)  and  a45799a );
 a45803a <=( (not A300)  and  A299 );
 a45806a <=( (not A302)  and  (not A301) );
 a45807a <=( a45806a  and  a45803a );
 a45808a <=( a45807a  and  a45800a );
 a45812a <=( A199  and  (not A168) );
 a45813a <=( (not A170)  and  a45812a );
 a45817a <=( A202  and  A201 );
 a45818a <=( (not A200)  and  a45817a );
 a45819a <=( a45818a  and  a45813a );
 a45823a <=( A298  and  A269 );
 a45824a <=( (not A267)  and  a45823a );
 a45827a <=( (not A300)  and  (not A299) );
 a45830a <=( (not A302)  and  (not A301) );
 a45831a <=( a45830a  and  a45827a );
 a45832a <=( a45831a  and  a45824a );
 a45836a <=( A199  and  (not A168) );
 a45837a <=( (not A170)  and  a45836a );
 a45841a <=( A202  and  A201 );
 a45842a <=( (not A200)  and  a45841a );
 a45843a <=( a45842a  and  a45837a );
 a45847a <=( (not A298)  and  A269 );
 a45848a <=( (not A267)  and  a45847a );
 a45851a <=( (not A300)  and  A299 );
 a45854a <=( (not A302)  and  (not A301) );
 a45855a <=( a45854a  and  a45851a );
 a45856a <=( a45855a  and  a45848a );
 a45860a <=( A199  and  (not A168) );
 a45861a <=( (not A170)  and  a45860a );
 a45865a <=( A202  and  A201 );
 a45866a <=( (not A200)  and  a45865a );
 a45867a <=( a45866a  and  a45861a );
 a45871a <=( A298  and  A266 );
 a45872a <=( A265  and  a45871a );
 a45875a <=( (not A300)  and  (not A299) );
 a45878a <=( (not A302)  and  (not A301) );
 a45879a <=( a45878a  and  a45875a );
 a45880a <=( a45879a  and  a45872a );
 a45884a <=( A199  and  (not A168) );
 a45885a <=( (not A170)  and  a45884a );
 a45889a <=( A202  and  A201 );
 a45890a <=( (not A200)  and  a45889a );
 a45891a <=( a45890a  and  a45885a );
 a45895a <=( (not A298)  and  A266 );
 a45896a <=( A265  and  a45895a );
 a45899a <=( (not A300)  and  A299 );
 a45902a <=( (not A302)  and  (not A301) );
 a45903a <=( a45902a  and  a45899a );
 a45904a <=( a45903a  and  a45896a );
 a45908a <=( A199  and  (not A168) );
 a45909a <=( (not A170)  and  a45908a );
 a45913a <=( A202  and  A201 );
 a45914a <=( (not A200)  and  a45913a );
 a45915a <=( a45914a  and  a45909a );
 a45919a <=( A298  and  (not A266) );
 a45920a <=( (not A265)  and  a45919a );
 a45923a <=( (not A300)  and  (not A299) );
 a45926a <=( (not A302)  and  (not A301) );
 a45927a <=( a45926a  and  a45923a );
 a45928a <=( a45927a  and  a45920a );
 a45932a <=( A199  and  (not A168) );
 a45933a <=( (not A170)  and  a45932a );
 a45937a <=( A202  and  A201 );
 a45938a <=( (not A200)  and  a45937a );
 a45939a <=( a45938a  and  a45933a );
 a45943a <=( (not A298)  and  (not A266) );
 a45944a <=( (not A265)  and  a45943a );
 a45947a <=( (not A300)  and  A299 );
 a45950a <=( (not A302)  and  (not A301) );
 a45951a <=( a45950a  and  a45947a );
 a45952a <=( a45951a  and  a45944a );
 a45956a <=( A199  and  (not A168) );
 a45957a <=( (not A170)  and  a45956a );
 a45961a <=( A203  and  A201 );
 a45962a <=( (not A200)  and  a45961a );
 a45963a <=( a45962a  and  a45957a );
 a45967a <=( (not A269)  and  (not A268) );
 a45968a <=( A267  and  a45967a );
 a45971a <=( (not A299)  and  A298 );
 a45974a <=( A301  and  A300 );
 a45975a <=( a45974a  and  a45971a );
 a45976a <=( a45975a  and  a45968a );
 a45980a <=( A199  and  (not A168) );
 a45981a <=( (not A170)  and  a45980a );
 a45985a <=( A203  and  A201 );
 a45986a <=( (not A200)  and  a45985a );
 a45987a <=( a45986a  and  a45981a );
 a45991a <=( (not A269)  and  (not A268) );
 a45992a <=( A267  and  a45991a );
 a45995a <=( (not A299)  and  A298 );
 a45998a <=( A302  and  A300 );
 a45999a <=( a45998a  and  a45995a );
 a46000a <=( a45999a  and  a45992a );
 a46004a <=( A199  and  (not A168) );
 a46005a <=( (not A170)  and  a46004a );
 a46009a <=( A203  and  A201 );
 a46010a <=( (not A200)  and  a46009a );
 a46011a <=( a46010a  and  a46005a );
 a46015a <=( (not A269)  and  (not A268) );
 a46016a <=( A267  and  a46015a );
 a46019a <=( A299  and  (not A298) );
 a46022a <=( A301  and  A300 );
 a46023a <=( a46022a  and  a46019a );
 a46024a <=( a46023a  and  a46016a );
 a46028a <=( A199  and  (not A168) );
 a46029a <=( (not A170)  and  a46028a );
 a46033a <=( A203  and  A201 );
 a46034a <=( (not A200)  and  a46033a );
 a46035a <=( a46034a  and  a46029a );
 a46039a <=( (not A269)  and  (not A268) );
 a46040a <=( A267  and  a46039a );
 a46043a <=( A299  and  (not A298) );
 a46046a <=( A302  and  A300 );
 a46047a <=( a46046a  and  a46043a );
 a46048a <=( a46047a  and  a46040a );
 a46052a <=( A199  and  (not A168) );
 a46053a <=( (not A170)  and  a46052a );
 a46057a <=( A203  and  A201 );
 a46058a <=( (not A200)  and  a46057a );
 a46059a <=( a46058a  and  a46053a );
 a46063a <=( A298  and  A268 );
 a46064a <=( (not A267)  and  a46063a );
 a46067a <=( (not A300)  and  (not A299) );
 a46070a <=( (not A302)  and  (not A301) );
 a46071a <=( a46070a  and  a46067a );
 a46072a <=( a46071a  and  a46064a );
 a46076a <=( A199  and  (not A168) );
 a46077a <=( (not A170)  and  a46076a );
 a46081a <=( A203  and  A201 );
 a46082a <=( (not A200)  and  a46081a );
 a46083a <=( a46082a  and  a46077a );
 a46087a <=( (not A298)  and  A268 );
 a46088a <=( (not A267)  and  a46087a );
 a46091a <=( (not A300)  and  A299 );
 a46094a <=( (not A302)  and  (not A301) );
 a46095a <=( a46094a  and  a46091a );
 a46096a <=( a46095a  and  a46088a );
 a46100a <=( A199  and  (not A168) );
 a46101a <=( (not A170)  and  a46100a );
 a46105a <=( A203  and  A201 );
 a46106a <=( (not A200)  and  a46105a );
 a46107a <=( a46106a  and  a46101a );
 a46111a <=( A298  and  A269 );
 a46112a <=( (not A267)  and  a46111a );
 a46115a <=( (not A300)  and  (not A299) );
 a46118a <=( (not A302)  and  (not A301) );
 a46119a <=( a46118a  and  a46115a );
 a46120a <=( a46119a  and  a46112a );
 a46124a <=( A199  and  (not A168) );
 a46125a <=( (not A170)  and  a46124a );
 a46129a <=( A203  and  A201 );
 a46130a <=( (not A200)  and  a46129a );
 a46131a <=( a46130a  and  a46125a );
 a46135a <=( (not A298)  and  A269 );
 a46136a <=( (not A267)  and  a46135a );
 a46139a <=( (not A300)  and  A299 );
 a46142a <=( (not A302)  and  (not A301) );
 a46143a <=( a46142a  and  a46139a );
 a46144a <=( a46143a  and  a46136a );
 a46148a <=( A199  and  (not A168) );
 a46149a <=( (not A170)  and  a46148a );
 a46153a <=( A203  and  A201 );
 a46154a <=( (not A200)  and  a46153a );
 a46155a <=( a46154a  and  a46149a );
 a46159a <=( A298  and  A266 );
 a46160a <=( A265  and  a46159a );
 a46163a <=( (not A300)  and  (not A299) );
 a46166a <=( (not A302)  and  (not A301) );
 a46167a <=( a46166a  and  a46163a );
 a46168a <=( a46167a  and  a46160a );
 a46172a <=( A199  and  (not A168) );
 a46173a <=( (not A170)  and  a46172a );
 a46177a <=( A203  and  A201 );
 a46178a <=( (not A200)  and  a46177a );
 a46179a <=( a46178a  and  a46173a );
 a46183a <=( (not A298)  and  A266 );
 a46184a <=( A265  and  a46183a );
 a46187a <=( (not A300)  and  A299 );
 a46190a <=( (not A302)  and  (not A301) );
 a46191a <=( a46190a  and  a46187a );
 a46192a <=( a46191a  and  a46184a );
 a46196a <=( A199  and  (not A168) );
 a46197a <=( (not A170)  and  a46196a );
 a46201a <=( A203  and  A201 );
 a46202a <=( (not A200)  and  a46201a );
 a46203a <=( a46202a  and  a46197a );
 a46207a <=( A298  and  (not A266) );
 a46208a <=( (not A265)  and  a46207a );
 a46211a <=( (not A300)  and  (not A299) );
 a46214a <=( (not A302)  and  (not A301) );
 a46215a <=( a46214a  and  a46211a );
 a46216a <=( a46215a  and  a46208a );
 a46220a <=( A199  and  (not A168) );
 a46221a <=( (not A170)  and  a46220a );
 a46225a <=( A203  and  A201 );
 a46226a <=( (not A200)  and  a46225a );
 a46227a <=( a46226a  and  a46221a );
 a46231a <=( (not A298)  and  (not A266) );
 a46232a <=( (not A265)  and  a46231a );
 a46235a <=( (not A300)  and  A299 );
 a46238a <=( (not A302)  and  (not A301) );
 a46239a <=( a46238a  and  a46235a );
 a46240a <=( a46239a  and  a46232a );
 a46244a <=( A199  and  (not A168) );
 a46245a <=( (not A170)  and  a46244a );
 a46249a <=( (not A202)  and  (not A201) );
 a46250a <=( (not A200)  and  a46249a );
 a46251a <=( a46250a  and  a46245a );
 a46255a <=( A268  and  (not A267) );
 a46256a <=( (not A203)  and  a46255a );
 a46259a <=( (not A299)  and  A298 );
 a46262a <=( A301  and  A300 );
 a46263a <=( a46262a  and  a46259a );
 a46264a <=( a46263a  and  a46256a );
 a46268a <=( A199  and  (not A168) );
 a46269a <=( (not A170)  and  a46268a );
 a46273a <=( (not A202)  and  (not A201) );
 a46274a <=( (not A200)  and  a46273a );
 a46275a <=( a46274a  and  a46269a );
 a46279a <=( A268  and  (not A267) );
 a46280a <=( (not A203)  and  a46279a );
 a46283a <=( (not A299)  and  A298 );
 a46286a <=( A302  and  A300 );
 a46287a <=( a46286a  and  a46283a );
 a46288a <=( a46287a  and  a46280a );
 a46292a <=( A199  and  (not A168) );
 a46293a <=( (not A170)  and  a46292a );
 a46297a <=( (not A202)  and  (not A201) );
 a46298a <=( (not A200)  and  a46297a );
 a46299a <=( a46298a  and  a46293a );
 a46303a <=( A268  and  (not A267) );
 a46304a <=( (not A203)  and  a46303a );
 a46307a <=( A299  and  (not A298) );
 a46310a <=( A301  and  A300 );
 a46311a <=( a46310a  and  a46307a );
 a46312a <=( a46311a  and  a46304a );
 a46316a <=( A199  and  (not A168) );
 a46317a <=( (not A170)  and  a46316a );
 a46321a <=( (not A202)  and  (not A201) );
 a46322a <=( (not A200)  and  a46321a );
 a46323a <=( a46322a  and  a46317a );
 a46327a <=( A268  and  (not A267) );
 a46328a <=( (not A203)  and  a46327a );
 a46331a <=( A299  and  (not A298) );
 a46334a <=( A302  and  A300 );
 a46335a <=( a46334a  and  a46331a );
 a46336a <=( a46335a  and  a46328a );
 a46340a <=( A199  and  (not A168) );
 a46341a <=( (not A170)  and  a46340a );
 a46345a <=( (not A202)  and  (not A201) );
 a46346a <=( (not A200)  and  a46345a );
 a46347a <=( a46346a  and  a46341a );
 a46351a <=( A269  and  (not A267) );
 a46352a <=( (not A203)  and  a46351a );
 a46355a <=( (not A299)  and  A298 );
 a46358a <=( A301  and  A300 );
 a46359a <=( a46358a  and  a46355a );
 a46360a <=( a46359a  and  a46352a );
 a46364a <=( A199  and  (not A168) );
 a46365a <=( (not A170)  and  a46364a );
 a46369a <=( (not A202)  and  (not A201) );
 a46370a <=( (not A200)  and  a46369a );
 a46371a <=( a46370a  and  a46365a );
 a46375a <=( A269  and  (not A267) );
 a46376a <=( (not A203)  and  a46375a );
 a46379a <=( (not A299)  and  A298 );
 a46382a <=( A302  and  A300 );
 a46383a <=( a46382a  and  a46379a );
 a46384a <=( a46383a  and  a46376a );
 a46388a <=( A199  and  (not A168) );
 a46389a <=( (not A170)  and  a46388a );
 a46393a <=( (not A202)  and  (not A201) );
 a46394a <=( (not A200)  and  a46393a );
 a46395a <=( a46394a  and  a46389a );
 a46399a <=( A269  and  (not A267) );
 a46400a <=( (not A203)  and  a46399a );
 a46403a <=( A299  and  (not A298) );
 a46406a <=( A301  and  A300 );
 a46407a <=( a46406a  and  a46403a );
 a46408a <=( a46407a  and  a46400a );
 a46412a <=( A199  and  (not A168) );
 a46413a <=( (not A170)  and  a46412a );
 a46417a <=( (not A202)  and  (not A201) );
 a46418a <=( (not A200)  and  a46417a );
 a46419a <=( a46418a  and  a46413a );
 a46423a <=( A269  and  (not A267) );
 a46424a <=( (not A203)  and  a46423a );
 a46427a <=( A299  and  (not A298) );
 a46430a <=( A302  and  A300 );
 a46431a <=( a46430a  and  a46427a );
 a46432a <=( a46431a  and  a46424a );
 a46436a <=( A199  and  (not A168) );
 a46437a <=( (not A170)  and  a46436a );
 a46441a <=( (not A202)  and  (not A201) );
 a46442a <=( (not A200)  and  a46441a );
 a46443a <=( a46442a  and  a46437a );
 a46447a <=( A266  and  A265 );
 a46448a <=( (not A203)  and  a46447a );
 a46451a <=( (not A299)  and  A298 );
 a46454a <=( A301  and  A300 );
 a46455a <=( a46454a  and  a46451a );
 a46456a <=( a46455a  and  a46448a );
 a46460a <=( A199  and  (not A168) );
 a46461a <=( (not A170)  and  a46460a );
 a46465a <=( (not A202)  and  (not A201) );
 a46466a <=( (not A200)  and  a46465a );
 a46467a <=( a46466a  and  a46461a );
 a46471a <=( A266  and  A265 );
 a46472a <=( (not A203)  and  a46471a );
 a46475a <=( (not A299)  and  A298 );
 a46478a <=( A302  and  A300 );
 a46479a <=( a46478a  and  a46475a );
 a46480a <=( a46479a  and  a46472a );
 a46484a <=( A199  and  (not A168) );
 a46485a <=( (not A170)  and  a46484a );
 a46489a <=( (not A202)  and  (not A201) );
 a46490a <=( (not A200)  and  a46489a );
 a46491a <=( a46490a  and  a46485a );
 a46495a <=( A266  and  A265 );
 a46496a <=( (not A203)  and  a46495a );
 a46499a <=( A299  and  (not A298) );
 a46502a <=( A301  and  A300 );
 a46503a <=( a46502a  and  a46499a );
 a46504a <=( a46503a  and  a46496a );
 a46508a <=( A199  and  (not A168) );
 a46509a <=( (not A170)  and  a46508a );
 a46513a <=( (not A202)  and  (not A201) );
 a46514a <=( (not A200)  and  a46513a );
 a46515a <=( a46514a  and  a46509a );
 a46519a <=( A266  and  A265 );
 a46520a <=( (not A203)  and  a46519a );
 a46523a <=( A299  and  (not A298) );
 a46526a <=( A302  and  A300 );
 a46527a <=( a46526a  and  a46523a );
 a46528a <=( a46527a  and  a46520a );
 a46532a <=( A199  and  (not A168) );
 a46533a <=( (not A170)  and  a46532a );
 a46537a <=( (not A202)  and  (not A201) );
 a46538a <=( (not A200)  and  a46537a );
 a46539a <=( a46538a  and  a46533a );
 a46543a <=( (not A266)  and  (not A265) );
 a46544a <=( (not A203)  and  a46543a );
 a46547a <=( (not A299)  and  A298 );
 a46550a <=( A301  and  A300 );
 a46551a <=( a46550a  and  a46547a );
 a46552a <=( a46551a  and  a46544a );
 a46556a <=( A199  and  (not A168) );
 a46557a <=( (not A170)  and  a46556a );
 a46561a <=( (not A202)  and  (not A201) );
 a46562a <=( (not A200)  and  a46561a );
 a46563a <=( a46562a  and  a46557a );
 a46567a <=( (not A266)  and  (not A265) );
 a46568a <=( (not A203)  and  a46567a );
 a46571a <=( (not A299)  and  A298 );
 a46574a <=( A302  and  A300 );
 a46575a <=( a46574a  and  a46571a );
 a46576a <=( a46575a  and  a46568a );
 a46580a <=( A199  and  (not A168) );
 a46581a <=( (not A170)  and  a46580a );
 a46585a <=( (not A202)  and  (not A201) );
 a46586a <=( (not A200)  and  a46585a );
 a46587a <=( a46586a  and  a46581a );
 a46591a <=( (not A266)  and  (not A265) );
 a46592a <=( (not A203)  and  a46591a );
 a46595a <=( A299  and  (not A298) );
 a46598a <=( A301  and  A300 );
 a46599a <=( a46598a  and  a46595a );
 a46600a <=( a46599a  and  a46592a );
 a46604a <=( A199  and  (not A168) );
 a46605a <=( (not A170)  and  a46604a );
 a46609a <=( (not A202)  and  (not A201) );
 a46610a <=( (not A200)  and  a46609a );
 a46611a <=( a46610a  and  a46605a );
 a46615a <=( (not A266)  and  (not A265) );
 a46616a <=( (not A203)  and  a46615a );
 a46619a <=( A299  and  (not A298) );
 a46622a <=( A302  and  A300 );
 a46623a <=( a46622a  and  a46619a );
 a46624a <=( a46623a  and  a46616a );
 a46628a <=( A167  and  A168 );
 a46629a <=( A169  and  a46628a );
 a46633a <=( (not A202)  and  A201 );
 a46634a <=( (not A166)  and  a46633a );
 a46635a <=( a46634a  and  a46629a );
 a46639a <=( A268  and  (not A267) );
 a46640a <=( (not A203)  and  a46639a );
 a46643a <=( (not A299)  and  A298 );
 a46646a <=( A301  and  A300 );
 a46647a <=( a46646a  and  a46643a );
 a46648a <=( a46647a  and  a46640a );
 a46652a <=( A167  and  A168 );
 a46653a <=( A169  and  a46652a );
 a46657a <=( (not A202)  and  A201 );
 a46658a <=( (not A166)  and  a46657a );
 a46659a <=( a46658a  and  a46653a );
 a46663a <=( A268  and  (not A267) );
 a46664a <=( (not A203)  and  a46663a );
 a46667a <=( (not A299)  and  A298 );
 a46670a <=( A302  and  A300 );
 a46671a <=( a46670a  and  a46667a );
 a46672a <=( a46671a  and  a46664a );
 a46676a <=( A167  and  A168 );
 a46677a <=( A169  and  a46676a );
 a46681a <=( (not A202)  and  A201 );
 a46682a <=( (not A166)  and  a46681a );
 a46683a <=( a46682a  and  a46677a );
 a46687a <=( A268  and  (not A267) );
 a46688a <=( (not A203)  and  a46687a );
 a46691a <=( A299  and  (not A298) );
 a46694a <=( A301  and  A300 );
 a46695a <=( a46694a  and  a46691a );
 a46696a <=( a46695a  and  a46688a );
 a46700a <=( A167  and  A168 );
 a46701a <=( A169  and  a46700a );
 a46705a <=( (not A202)  and  A201 );
 a46706a <=( (not A166)  and  a46705a );
 a46707a <=( a46706a  and  a46701a );
 a46711a <=( A268  and  (not A267) );
 a46712a <=( (not A203)  and  a46711a );
 a46715a <=( A299  and  (not A298) );
 a46718a <=( A302  and  A300 );
 a46719a <=( a46718a  and  a46715a );
 a46720a <=( a46719a  and  a46712a );
 a46724a <=( A167  and  A168 );
 a46725a <=( A169  and  a46724a );
 a46729a <=( (not A202)  and  A201 );
 a46730a <=( (not A166)  and  a46729a );
 a46731a <=( a46730a  and  a46725a );
 a46735a <=( A269  and  (not A267) );
 a46736a <=( (not A203)  and  a46735a );
 a46739a <=( (not A299)  and  A298 );
 a46742a <=( A301  and  A300 );
 a46743a <=( a46742a  and  a46739a );
 a46744a <=( a46743a  and  a46736a );
 a46748a <=( A167  and  A168 );
 a46749a <=( A169  and  a46748a );
 a46753a <=( (not A202)  and  A201 );
 a46754a <=( (not A166)  and  a46753a );
 a46755a <=( a46754a  and  a46749a );
 a46759a <=( A269  and  (not A267) );
 a46760a <=( (not A203)  and  a46759a );
 a46763a <=( (not A299)  and  A298 );
 a46766a <=( A302  and  A300 );
 a46767a <=( a46766a  and  a46763a );
 a46768a <=( a46767a  and  a46760a );
 a46772a <=( A167  and  A168 );
 a46773a <=( A169  and  a46772a );
 a46777a <=( (not A202)  and  A201 );
 a46778a <=( (not A166)  and  a46777a );
 a46779a <=( a46778a  and  a46773a );
 a46783a <=( A269  and  (not A267) );
 a46784a <=( (not A203)  and  a46783a );
 a46787a <=( A299  and  (not A298) );
 a46790a <=( A301  and  A300 );
 a46791a <=( a46790a  and  a46787a );
 a46792a <=( a46791a  and  a46784a );
 a46796a <=( A167  and  A168 );
 a46797a <=( A169  and  a46796a );
 a46801a <=( (not A202)  and  A201 );
 a46802a <=( (not A166)  and  a46801a );
 a46803a <=( a46802a  and  a46797a );
 a46807a <=( A269  and  (not A267) );
 a46808a <=( (not A203)  and  a46807a );
 a46811a <=( A299  and  (not A298) );
 a46814a <=( A302  and  A300 );
 a46815a <=( a46814a  and  a46811a );
 a46816a <=( a46815a  and  a46808a );
 a46820a <=( A167  and  A168 );
 a46821a <=( A169  and  a46820a );
 a46825a <=( (not A202)  and  A201 );
 a46826a <=( (not A166)  and  a46825a );
 a46827a <=( a46826a  and  a46821a );
 a46831a <=( A266  and  A265 );
 a46832a <=( (not A203)  and  a46831a );
 a46835a <=( (not A299)  and  A298 );
 a46838a <=( A301  and  A300 );
 a46839a <=( a46838a  and  a46835a );
 a46840a <=( a46839a  and  a46832a );
 a46844a <=( A167  and  A168 );
 a46845a <=( A169  and  a46844a );
 a46849a <=( (not A202)  and  A201 );
 a46850a <=( (not A166)  and  a46849a );
 a46851a <=( a46850a  and  a46845a );
 a46855a <=( A266  and  A265 );
 a46856a <=( (not A203)  and  a46855a );
 a46859a <=( (not A299)  and  A298 );
 a46862a <=( A302  and  A300 );
 a46863a <=( a46862a  and  a46859a );
 a46864a <=( a46863a  and  a46856a );
 a46868a <=( A167  and  A168 );
 a46869a <=( A169  and  a46868a );
 a46873a <=( (not A202)  and  A201 );
 a46874a <=( (not A166)  and  a46873a );
 a46875a <=( a46874a  and  a46869a );
 a46879a <=( A266  and  A265 );
 a46880a <=( (not A203)  and  a46879a );
 a46883a <=( A299  and  (not A298) );
 a46886a <=( A301  and  A300 );
 a46887a <=( a46886a  and  a46883a );
 a46888a <=( a46887a  and  a46880a );
 a46892a <=( A167  and  A168 );
 a46893a <=( A169  and  a46892a );
 a46897a <=( (not A202)  and  A201 );
 a46898a <=( (not A166)  and  a46897a );
 a46899a <=( a46898a  and  a46893a );
 a46903a <=( A266  and  A265 );
 a46904a <=( (not A203)  and  a46903a );
 a46907a <=( A299  and  (not A298) );
 a46910a <=( A302  and  A300 );
 a46911a <=( a46910a  and  a46907a );
 a46912a <=( a46911a  and  a46904a );
 a46916a <=( A167  and  A168 );
 a46917a <=( A169  and  a46916a );
 a46921a <=( (not A202)  and  A201 );
 a46922a <=( (not A166)  and  a46921a );
 a46923a <=( a46922a  and  a46917a );
 a46927a <=( (not A266)  and  (not A265) );
 a46928a <=( (not A203)  and  a46927a );
 a46931a <=( (not A299)  and  A298 );
 a46934a <=( A301  and  A300 );
 a46935a <=( a46934a  and  a46931a );
 a46936a <=( a46935a  and  a46928a );
 a46940a <=( A167  and  A168 );
 a46941a <=( A169  and  a46940a );
 a46945a <=( (not A202)  and  A201 );
 a46946a <=( (not A166)  and  a46945a );
 a46947a <=( a46946a  and  a46941a );
 a46951a <=( (not A266)  and  (not A265) );
 a46952a <=( (not A203)  and  a46951a );
 a46955a <=( (not A299)  and  A298 );
 a46958a <=( A302  and  A300 );
 a46959a <=( a46958a  and  a46955a );
 a46960a <=( a46959a  and  a46952a );
 a46964a <=( A167  and  A168 );
 a46965a <=( A169  and  a46964a );
 a46969a <=( (not A202)  and  A201 );
 a46970a <=( (not A166)  and  a46969a );
 a46971a <=( a46970a  and  a46965a );
 a46975a <=( (not A266)  and  (not A265) );
 a46976a <=( (not A203)  and  a46975a );
 a46979a <=( A299  and  (not A298) );
 a46982a <=( A301  and  A300 );
 a46983a <=( a46982a  and  a46979a );
 a46984a <=( a46983a  and  a46976a );
 a46988a <=( A167  and  A168 );
 a46989a <=( A169  and  a46988a );
 a46993a <=( (not A202)  and  A201 );
 a46994a <=( (not A166)  and  a46993a );
 a46995a <=( a46994a  and  a46989a );
 a46999a <=( (not A266)  and  (not A265) );
 a47000a <=( (not A203)  and  a46999a );
 a47003a <=( A299  and  (not A298) );
 a47006a <=( A302  and  A300 );
 a47007a <=( a47006a  and  a47003a );
 a47008a <=( a47007a  and  a47000a );
 a47012a <=( A167  and  A168 );
 a47013a <=( A169  and  a47012a );
 a47017a <=( A202  and  (not A201) );
 a47018a <=( (not A166)  and  a47017a );
 a47019a <=( a47018a  and  a47013a );
 a47023a <=( (not A269)  and  (not A268) );
 a47024a <=( A267  and  a47023a );
 a47027a <=( (not A299)  and  A298 );
 a47030a <=( A301  and  A300 );
 a47031a <=( a47030a  and  a47027a );
 a47032a <=( a47031a  and  a47024a );
 a47036a <=( A167  and  A168 );
 a47037a <=( A169  and  a47036a );
 a47041a <=( A202  and  (not A201) );
 a47042a <=( (not A166)  and  a47041a );
 a47043a <=( a47042a  and  a47037a );
 a47047a <=( (not A269)  and  (not A268) );
 a47048a <=( A267  and  a47047a );
 a47051a <=( (not A299)  and  A298 );
 a47054a <=( A302  and  A300 );
 a47055a <=( a47054a  and  a47051a );
 a47056a <=( a47055a  and  a47048a );
 a47060a <=( A167  and  A168 );
 a47061a <=( A169  and  a47060a );
 a47065a <=( A202  and  (not A201) );
 a47066a <=( (not A166)  and  a47065a );
 a47067a <=( a47066a  and  a47061a );
 a47071a <=( (not A269)  and  (not A268) );
 a47072a <=( A267  and  a47071a );
 a47075a <=( A299  and  (not A298) );
 a47078a <=( A301  and  A300 );
 a47079a <=( a47078a  and  a47075a );
 a47080a <=( a47079a  and  a47072a );
 a47084a <=( A167  and  A168 );
 a47085a <=( A169  and  a47084a );
 a47089a <=( A202  and  (not A201) );
 a47090a <=( (not A166)  and  a47089a );
 a47091a <=( a47090a  and  a47085a );
 a47095a <=( (not A269)  and  (not A268) );
 a47096a <=( A267  and  a47095a );
 a47099a <=( A299  and  (not A298) );
 a47102a <=( A302  and  A300 );
 a47103a <=( a47102a  and  a47099a );
 a47104a <=( a47103a  and  a47096a );
 a47108a <=( A167  and  A168 );
 a47109a <=( A169  and  a47108a );
 a47113a <=( A202  and  (not A201) );
 a47114a <=( (not A166)  and  a47113a );
 a47115a <=( a47114a  and  a47109a );
 a47119a <=( A298  and  A268 );
 a47120a <=( (not A267)  and  a47119a );
 a47123a <=( (not A300)  and  (not A299) );
 a47126a <=( (not A302)  and  (not A301) );
 a47127a <=( a47126a  and  a47123a );
 a47128a <=( a47127a  and  a47120a );
 a47132a <=( A167  and  A168 );
 a47133a <=( A169  and  a47132a );
 a47137a <=( A202  and  (not A201) );
 a47138a <=( (not A166)  and  a47137a );
 a47139a <=( a47138a  and  a47133a );
 a47143a <=( (not A298)  and  A268 );
 a47144a <=( (not A267)  and  a47143a );
 a47147a <=( (not A300)  and  A299 );
 a47150a <=( (not A302)  and  (not A301) );
 a47151a <=( a47150a  and  a47147a );
 a47152a <=( a47151a  and  a47144a );
 a47156a <=( A167  and  A168 );
 a47157a <=( A169  and  a47156a );
 a47161a <=( A202  and  (not A201) );
 a47162a <=( (not A166)  and  a47161a );
 a47163a <=( a47162a  and  a47157a );
 a47167a <=( A298  and  A269 );
 a47168a <=( (not A267)  and  a47167a );
 a47171a <=( (not A300)  and  (not A299) );
 a47174a <=( (not A302)  and  (not A301) );
 a47175a <=( a47174a  and  a47171a );
 a47176a <=( a47175a  and  a47168a );
 a47180a <=( A167  and  A168 );
 a47181a <=( A169  and  a47180a );
 a47185a <=( A202  and  (not A201) );
 a47186a <=( (not A166)  and  a47185a );
 a47187a <=( a47186a  and  a47181a );
 a47191a <=( (not A298)  and  A269 );
 a47192a <=( (not A267)  and  a47191a );
 a47195a <=( (not A300)  and  A299 );
 a47198a <=( (not A302)  and  (not A301) );
 a47199a <=( a47198a  and  a47195a );
 a47200a <=( a47199a  and  a47192a );
 a47204a <=( A167  and  A168 );
 a47205a <=( A169  and  a47204a );
 a47209a <=( A202  and  (not A201) );
 a47210a <=( (not A166)  and  a47209a );
 a47211a <=( a47210a  and  a47205a );
 a47215a <=( A298  and  A266 );
 a47216a <=( A265  and  a47215a );
 a47219a <=( (not A300)  and  (not A299) );
 a47222a <=( (not A302)  and  (not A301) );
 a47223a <=( a47222a  and  a47219a );
 a47224a <=( a47223a  and  a47216a );
 a47228a <=( A167  and  A168 );
 a47229a <=( A169  and  a47228a );
 a47233a <=( A202  and  (not A201) );
 a47234a <=( (not A166)  and  a47233a );
 a47235a <=( a47234a  and  a47229a );
 a47239a <=( (not A298)  and  A266 );
 a47240a <=( A265  and  a47239a );
 a47243a <=( (not A300)  and  A299 );
 a47246a <=( (not A302)  and  (not A301) );
 a47247a <=( a47246a  and  a47243a );
 a47248a <=( a47247a  and  a47240a );
 a47252a <=( A167  and  A168 );
 a47253a <=( A169  and  a47252a );
 a47257a <=( A202  and  (not A201) );
 a47258a <=( (not A166)  and  a47257a );
 a47259a <=( a47258a  and  a47253a );
 a47263a <=( A298  and  (not A266) );
 a47264a <=( (not A265)  and  a47263a );
 a47267a <=( (not A300)  and  (not A299) );
 a47270a <=( (not A302)  and  (not A301) );
 a47271a <=( a47270a  and  a47267a );
 a47272a <=( a47271a  and  a47264a );
 a47276a <=( A167  and  A168 );
 a47277a <=( A169  and  a47276a );
 a47281a <=( A202  and  (not A201) );
 a47282a <=( (not A166)  and  a47281a );
 a47283a <=( a47282a  and  a47277a );
 a47287a <=( (not A298)  and  (not A266) );
 a47288a <=( (not A265)  and  a47287a );
 a47291a <=( (not A300)  and  A299 );
 a47294a <=( (not A302)  and  (not A301) );
 a47295a <=( a47294a  and  a47291a );
 a47296a <=( a47295a  and  a47288a );
 a47300a <=( A167  and  A168 );
 a47301a <=( A169  and  a47300a );
 a47305a <=( A203  and  (not A201) );
 a47306a <=( (not A166)  and  a47305a );
 a47307a <=( a47306a  and  a47301a );
 a47311a <=( (not A269)  and  (not A268) );
 a47312a <=( A267  and  a47311a );
 a47315a <=( (not A299)  and  A298 );
 a47318a <=( A301  and  A300 );
 a47319a <=( a47318a  and  a47315a );
 a47320a <=( a47319a  and  a47312a );
 a47324a <=( A167  and  A168 );
 a47325a <=( A169  and  a47324a );
 a47329a <=( A203  and  (not A201) );
 a47330a <=( (not A166)  and  a47329a );
 a47331a <=( a47330a  and  a47325a );
 a47335a <=( (not A269)  and  (not A268) );
 a47336a <=( A267  and  a47335a );
 a47339a <=( (not A299)  and  A298 );
 a47342a <=( A302  and  A300 );
 a47343a <=( a47342a  and  a47339a );
 a47344a <=( a47343a  and  a47336a );
 a47348a <=( A167  and  A168 );
 a47349a <=( A169  and  a47348a );
 a47353a <=( A203  and  (not A201) );
 a47354a <=( (not A166)  and  a47353a );
 a47355a <=( a47354a  and  a47349a );
 a47359a <=( (not A269)  and  (not A268) );
 a47360a <=( A267  and  a47359a );
 a47363a <=( A299  and  (not A298) );
 a47366a <=( A301  and  A300 );
 a47367a <=( a47366a  and  a47363a );
 a47368a <=( a47367a  and  a47360a );
 a47372a <=( A167  and  A168 );
 a47373a <=( A169  and  a47372a );
 a47377a <=( A203  and  (not A201) );
 a47378a <=( (not A166)  and  a47377a );
 a47379a <=( a47378a  and  a47373a );
 a47383a <=( (not A269)  and  (not A268) );
 a47384a <=( A267  and  a47383a );
 a47387a <=( A299  and  (not A298) );
 a47390a <=( A302  and  A300 );
 a47391a <=( a47390a  and  a47387a );
 a47392a <=( a47391a  and  a47384a );
 a47396a <=( A167  and  A168 );
 a47397a <=( A169  and  a47396a );
 a47401a <=( A203  and  (not A201) );
 a47402a <=( (not A166)  and  a47401a );
 a47403a <=( a47402a  and  a47397a );
 a47407a <=( A298  and  A268 );
 a47408a <=( (not A267)  and  a47407a );
 a47411a <=( (not A300)  and  (not A299) );
 a47414a <=( (not A302)  and  (not A301) );
 a47415a <=( a47414a  and  a47411a );
 a47416a <=( a47415a  and  a47408a );
 a47420a <=( A167  and  A168 );
 a47421a <=( A169  and  a47420a );
 a47425a <=( A203  and  (not A201) );
 a47426a <=( (not A166)  and  a47425a );
 a47427a <=( a47426a  and  a47421a );
 a47431a <=( (not A298)  and  A268 );
 a47432a <=( (not A267)  and  a47431a );
 a47435a <=( (not A300)  and  A299 );
 a47438a <=( (not A302)  and  (not A301) );
 a47439a <=( a47438a  and  a47435a );
 a47440a <=( a47439a  and  a47432a );
 a47444a <=( A167  and  A168 );
 a47445a <=( A169  and  a47444a );
 a47449a <=( A203  and  (not A201) );
 a47450a <=( (not A166)  and  a47449a );
 a47451a <=( a47450a  and  a47445a );
 a47455a <=( A298  and  A269 );
 a47456a <=( (not A267)  and  a47455a );
 a47459a <=( (not A300)  and  (not A299) );
 a47462a <=( (not A302)  and  (not A301) );
 a47463a <=( a47462a  and  a47459a );
 a47464a <=( a47463a  and  a47456a );
 a47468a <=( A167  and  A168 );
 a47469a <=( A169  and  a47468a );
 a47473a <=( A203  and  (not A201) );
 a47474a <=( (not A166)  and  a47473a );
 a47475a <=( a47474a  and  a47469a );
 a47479a <=( (not A298)  and  A269 );
 a47480a <=( (not A267)  and  a47479a );
 a47483a <=( (not A300)  and  A299 );
 a47486a <=( (not A302)  and  (not A301) );
 a47487a <=( a47486a  and  a47483a );
 a47488a <=( a47487a  and  a47480a );
 a47492a <=( A167  and  A168 );
 a47493a <=( A169  and  a47492a );
 a47497a <=( A203  and  (not A201) );
 a47498a <=( (not A166)  and  a47497a );
 a47499a <=( a47498a  and  a47493a );
 a47503a <=( A298  and  A266 );
 a47504a <=( A265  and  a47503a );
 a47507a <=( (not A300)  and  (not A299) );
 a47510a <=( (not A302)  and  (not A301) );
 a47511a <=( a47510a  and  a47507a );
 a47512a <=( a47511a  and  a47504a );
 a47516a <=( A167  and  A168 );
 a47517a <=( A169  and  a47516a );
 a47521a <=( A203  and  (not A201) );
 a47522a <=( (not A166)  and  a47521a );
 a47523a <=( a47522a  and  a47517a );
 a47527a <=( (not A298)  and  A266 );
 a47528a <=( A265  and  a47527a );
 a47531a <=( (not A300)  and  A299 );
 a47534a <=( (not A302)  and  (not A301) );
 a47535a <=( a47534a  and  a47531a );
 a47536a <=( a47535a  and  a47528a );
 a47540a <=( A167  and  A168 );
 a47541a <=( A169  and  a47540a );
 a47545a <=( A203  and  (not A201) );
 a47546a <=( (not A166)  and  a47545a );
 a47547a <=( a47546a  and  a47541a );
 a47551a <=( A298  and  (not A266) );
 a47552a <=( (not A265)  and  a47551a );
 a47555a <=( (not A300)  and  (not A299) );
 a47558a <=( (not A302)  and  (not A301) );
 a47559a <=( a47558a  and  a47555a );
 a47560a <=( a47559a  and  a47552a );
 a47564a <=( A167  and  A168 );
 a47565a <=( A169  and  a47564a );
 a47569a <=( A203  and  (not A201) );
 a47570a <=( (not A166)  and  a47569a );
 a47571a <=( a47570a  and  a47565a );
 a47575a <=( (not A298)  and  (not A266) );
 a47576a <=( (not A265)  and  a47575a );
 a47579a <=( (not A300)  and  A299 );
 a47582a <=( (not A302)  and  (not A301) );
 a47583a <=( a47582a  and  a47579a );
 a47584a <=( a47583a  and  a47576a );
 a47588a <=( A167  and  A168 );
 a47589a <=( A169  and  a47588a );
 a47593a <=( A200  and  A199 );
 a47594a <=( (not A166)  and  a47593a );
 a47595a <=( a47594a  and  a47589a );
 a47599a <=( (not A269)  and  (not A268) );
 a47600a <=( A267  and  a47599a );
 a47603a <=( (not A299)  and  A298 );
 a47606a <=( A301  and  A300 );
 a47607a <=( a47606a  and  a47603a );
 a47608a <=( a47607a  and  a47600a );
 a47612a <=( A167  and  A168 );
 a47613a <=( A169  and  a47612a );
 a47617a <=( A200  and  A199 );
 a47618a <=( (not A166)  and  a47617a );
 a47619a <=( a47618a  and  a47613a );
 a47623a <=( (not A269)  and  (not A268) );
 a47624a <=( A267  and  a47623a );
 a47627a <=( (not A299)  and  A298 );
 a47630a <=( A302  and  A300 );
 a47631a <=( a47630a  and  a47627a );
 a47632a <=( a47631a  and  a47624a );
 a47636a <=( A167  and  A168 );
 a47637a <=( A169  and  a47636a );
 a47641a <=( A200  and  A199 );
 a47642a <=( (not A166)  and  a47641a );
 a47643a <=( a47642a  and  a47637a );
 a47647a <=( (not A269)  and  (not A268) );
 a47648a <=( A267  and  a47647a );
 a47651a <=( A299  and  (not A298) );
 a47654a <=( A301  and  A300 );
 a47655a <=( a47654a  and  a47651a );
 a47656a <=( a47655a  and  a47648a );
 a47660a <=( A167  and  A168 );
 a47661a <=( A169  and  a47660a );
 a47665a <=( A200  and  A199 );
 a47666a <=( (not A166)  and  a47665a );
 a47667a <=( a47666a  and  a47661a );
 a47671a <=( (not A269)  and  (not A268) );
 a47672a <=( A267  and  a47671a );
 a47675a <=( A299  and  (not A298) );
 a47678a <=( A302  and  A300 );
 a47679a <=( a47678a  and  a47675a );
 a47680a <=( a47679a  and  a47672a );
 a47684a <=( A167  and  A168 );
 a47685a <=( A169  and  a47684a );
 a47689a <=( A200  and  A199 );
 a47690a <=( (not A166)  and  a47689a );
 a47691a <=( a47690a  and  a47685a );
 a47695a <=( A298  and  A268 );
 a47696a <=( (not A267)  and  a47695a );
 a47699a <=( (not A300)  and  (not A299) );
 a47702a <=( (not A302)  and  (not A301) );
 a47703a <=( a47702a  and  a47699a );
 a47704a <=( a47703a  and  a47696a );
 a47708a <=( A167  and  A168 );
 a47709a <=( A169  and  a47708a );
 a47713a <=( A200  and  A199 );
 a47714a <=( (not A166)  and  a47713a );
 a47715a <=( a47714a  and  a47709a );
 a47719a <=( (not A298)  and  A268 );
 a47720a <=( (not A267)  and  a47719a );
 a47723a <=( (not A300)  and  A299 );
 a47726a <=( (not A302)  and  (not A301) );
 a47727a <=( a47726a  and  a47723a );
 a47728a <=( a47727a  and  a47720a );
 a47732a <=( A167  and  A168 );
 a47733a <=( A169  and  a47732a );
 a47737a <=( A200  and  A199 );
 a47738a <=( (not A166)  and  a47737a );
 a47739a <=( a47738a  and  a47733a );
 a47743a <=( A298  and  A269 );
 a47744a <=( (not A267)  and  a47743a );
 a47747a <=( (not A300)  and  (not A299) );
 a47750a <=( (not A302)  and  (not A301) );
 a47751a <=( a47750a  and  a47747a );
 a47752a <=( a47751a  and  a47744a );
 a47756a <=( A167  and  A168 );
 a47757a <=( A169  and  a47756a );
 a47761a <=( A200  and  A199 );
 a47762a <=( (not A166)  and  a47761a );
 a47763a <=( a47762a  and  a47757a );
 a47767a <=( (not A298)  and  A269 );
 a47768a <=( (not A267)  and  a47767a );
 a47771a <=( (not A300)  and  A299 );
 a47774a <=( (not A302)  and  (not A301) );
 a47775a <=( a47774a  and  a47771a );
 a47776a <=( a47775a  and  a47768a );
 a47780a <=( A167  and  A168 );
 a47781a <=( A169  and  a47780a );
 a47785a <=( A200  and  A199 );
 a47786a <=( (not A166)  and  a47785a );
 a47787a <=( a47786a  and  a47781a );
 a47791a <=( A298  and  A266 );
 a47792a <=( A265  and  a47791a );
 a47795a <=( (not A300)  and  (not A299) );
 a47798a <=( (not A302)  and  (not A301) );
 a47799a <=( a47798a  and  a47795a );
 a47800a <=( a47799a  and  a47792a );
 a47804a <=( A167  and  A168 );
 a47805a <=( A169  and  a47804a );
 a47809a <=( A200  and  A199 );
 a47810a <=( (not A166)  and  a47809a );
 a47811a <=( a47810a  and  a47805a );
 a47815a <=( (not A298)  and  A266 );
 a47816a <=( A265  and  a47815a );
 a47819a <=( (not A300)  and  A299 );
 a47822a <=( (not A302)  and  (not A301) );
 a47823a <=( a47822a  and  a47819a );
 a47824a <=( a47823a  and  a47816a );
 a47828a <=( A167  and  A168 );
 a47829a <=( A169  and  a47828a );
 a47833a <=( A200  and  A199 );
 a47834a <=( (not A166)  and  a47833a );
 a47835a <=( a47834a  and  a47829a );
 a47839a <=( A298  and  (not A266) );
 a47840a <=( (not A265)  and  a47839a );
 a47843a <=( (not A300)  and  (not A299) );
 a47846a <=( (not A302)  and  (not A301) );
 a47847a <=( a47846a  and  a47843a );
 a47848a <=( a47847a  and  a47840a );
 a47852a <=( A167  and  A168 );
 a47853a <=( A169  and  a47852a );
 a47857a <=( A200  and  A199 );
 a47858a <=( (not A166)  and  a47857a );
 a47859a <=( a47858a  and  a47853a );
 a47863a <=( (not A298)  and  (not A266) );
 a47864a <=( (not A265)  and  a47863a );
 a47867a <=( (not A300)  and  A299 );
 a47870a <=( (not A302)  and  (not A301) );
 a47871a <=( a47870a  and  a47867a );
 a47872a <=( a47871a  and  a47864a );
 a47876a <=( A167  and  A168 );
 a47877a <=( A169  and  a47876a );
 a47881a <=( (not A200)  and  (not A199) );
 a47882a <=( (not A166)  and  a47881a );
 a47883a <=( a47882a  and  a47877a );
 a47887a <=( (not A269)  and  (not A268) );
 a47888a <=( A267  and  a47887a );
 a47891a <=( (not A299)  and  A298 );
 a47894a <=( A301  and  A300 );
 a47895a <=( a47894a  and  a47891a );
 a47896a <=( a47895a  and  a47888a );
 a47900a <=( A167  and  A168 );
 a47901a <=( A169  and  a47900a );
 a47905a <=( (not A200)  and  (not A199) );
 a47906a <=( (not A166)  and  a47905a );
 a47907a <=( a47906a  and  a47901a );
 a47911a <=( (not A269)  and  (not A268) );
 a47912a <=( A267  and  a47911a );
 a47915a <=( (not A299)  and  A298 );
 a47918a <=( A302  and  A300 );
 a47919a <=( a47918a  and  a47915a );
 a47920a <=( a47919a  and  a47912a );
 a47924a <=( A167  and  A168 );
 a47925a <=( A169  and  a47924a );
 a47929a <=( (not A200)  and  (not A199) );
 a47930a <=( (not A166)  and  a47929a );
 a47931a <=( a47930a  and  a47925a );
 a47935a <=( (not A269)  and  (not A268) );
 a47936a <=( A267  and  a47935a );
 a47939a <=( A299  and  (not A298) );
 a47942a <=( A301  and  A300 );
 a47943a <=( a47942a  and  a47939a );
 a47944a <=( a47943a  and  a47936a );
 a47948a <=( A167  and  A168 );
 a47949a <=( A169  and  a47948a );
 a47953a <=( (not A200)  and  (not A199) );
 a47954a <=( (not A166)  and  a47953a );
 a47955a <=( a47954a  and  a47949a );
 a47959a <=( (not A269)  and  (not A268) );
 a47960a <=( A267  and  a47959a );
 a47963a <=( A299  and  (not A298) );
 a47966a <=( A302  and  A300 );
 a47967a <=( a47966a  and  a47963a );
 a47968a <=( a47967a  and  a47960a );
 a47972a <=( A167  and  A168 );
 a47973a <=( A169  and  a47972a );
 a47977a <=( (not A200)  and  (not A199) );
 a47978a <=( (not A166)  and  a47977a );
 a47979a <=( a47978a  and  a47973a );
 a47983a <=( A298  and  A268 );
 a47984a <=( (not A267)  and  a47983a );
 a47987a <=( (not A300)  and  (not A299) );
 a47990a <=( (not A302)  and  (not A301) );
 a47991a <=( a47990a  and  a47987a );
 a47992a <=( a47991a  and  a47984a );
 a47996a <=( A167  and  A168 );
 a47997a <=( A169  and  a47996a );
 a48001a <=( (not A200)  and  (not A199) );
 a48002a <=( (not A166)  and  a48001a );
 a48003a <=( a48002a  and  a47997a );
 a48007a <=( (not A298)  and  A268 );
 a48008a <=( (not A267)  and  a48007a );
 a48011a <=( (not A300)  and  A299 );
 a48014a <=( (not A302)  and  (not A301) );
 a48015a <=( a48014a  and  a48011a );
 a48016a <=( a48015a  and  a48008a );
 a48020a <=( A167  and  A168 );
 a48021a <=( A169  and  a48020a );
 a48025a <=( (not A200)  and  (not A199) );
 a48026a <=( (not A166)  and  a48025a );
 a48027a <=( a48026a  and  a48021a );
 a48031a <=( A298  and  A269 );
 a48032a <=( (not A267)  and  a48031a );
 a48035a <=( (not A300)  and  (not A299) );
 a48038a <=( (not A302)  and  (not A301) );
 a48039a <=( a48038a  and  a48035a );
 a48040a <=( a48039a  and  a48032a );
 a48044a <=( A167  and  A168 );
 a48045a <=( A169  and  a48044a );
 a48049a <=( (not A200)  and  (not A199) );
 a48050a <=( (not A166)  and  a48049a );
 a48051a <=( a48050a  and  a48045a );
 a48055a <=( (not A298)  and  A269 );
 a48056a <=( (not A267)  and  a48055a );
 a48059a <=( (not A300)  and  A299 );
 a48062a <=( (not A302)  and  (not A301) );
 a48063a <=( a48062a  and  a48059a );
 a48064a <=( a48063a  and  a48056a );
 a48068a <=( A167  and  A168 );
 a48069a <=( A169  and  a48068a );
 a48073a <=( (not A200)  and  (not A199) );
 a48074a <=( (not A166)  and  a48073a );
 a48075a <=( a48074a  and  a48069a );
 a48079a <=( A298  and  A266 );
 a48080a <=( A265  and  a48079a );
 a48083a <=( (not A300)  and  (not A299) );
 a48086a <=( (not A302)  and  (not A301) );
 a48087a <=( a48086a  and  a48083a );
 a48088a <=( a48087a  and  a48080a );
 a48092a <=( A167  and  A168 );
 a48093a <=( A169  and  a48092a );
 a48097a <=( (not A200)  and  (not A199) );
 a48098a <=( (not A166)  and  a48097a );
 a48099a <=( a48098a  and  a48093a );
 a48103a <=( (not A298)  and  A266 );
 a48104a <=( A265  and  a48103a );
 a48107a <=( (not A300)  and  A299 );
 a48110a <=( (not A302)  and  (not A301) );
 a48111a <=( a48110a  and  a48107a );
 a48112a <=( a48111a  and  a48104a );
 a48116a <=( A167  and  A168 );
 a48117a <=( A169  and  a48116a );
 a48121a <=( (not A200)  and  (not A199) );
 a48122a <=( (not A166)  and  a48121a );
 a48123a <=( a48122a  and  a48117a );
 a48127a <=( A298  and  (not A266) );
 a48128a <=( (not A265)  and  a48127a );
 a48131a <=( (not A300)  and  (not A299) );
 a48134a <=( (not A302)  and  (not A301) );
 a48135a <=( a48134a  and  a48131a );
 a48136a <=( a48135a  and  a48128a );
 a48140a <=( A167  and  A168 );
 a48141a <=( A169  and  a48140a );
 a48145a <=( (not A200)  and  (not A199) );
 a48146a <=( (not A166)  and  a48145a );
 a48147a <=( a48146a  and  a48141a );
 a48151a <=( (not A298)  and  (not A266) );
 a48152a <=( (not A265)  and  a48151a );
 a48155a <=( (not A300)  and  A299 );
 a48158a <=( (not A302)  and  (not A301) );
 a48159a <=( a48158a  and  a48155a );
 a48160a <=( a48159a  and  a48152a );
 a48164a <=( (not A167)  and  A168 );
 a48165a <=( A169  and  a48164a );
 a48169a <=( (not A202)  and  A201 );
 a48170a <=( A166  and  a48169a );
 a48171a <=( a48170a  and  a48165a );
 a48175a <=( A268  and  (not A267) );
 a48176a <=( (not A203)  and  a48175a );
 a48179a <=( (not A299)  and  A298 );
 a48182a <=( A301  and  A300 );
 a48183a <=( a48182a  and  a48179a );
 a48184a <=( a48183a  and  a48176a );
 a48188a <=( (not A167)  and  A168 );
 a48189a <=( A169  and  a48188a );
 a48193a <=( (not A202)  and  A201 );
 a48194a <=( A166  and  a48193a );
 a48195a <=( a48194a  and  a48189a );
 a48199a <=( A268  and  (not A267) );
 a48200a <=( (not A203)  and  a48199a );
 a48203a <=( (not A299)  and  A298 );
 a48206a <=( A302  and  A300 );
 a48207a <=( a48206a  and  a48203a );
 a48208a <=( a48207a  and  a48200a );
 a48212a <=( (not A167)  and  A168 );
 a48213a <=( A169  and  a48212a );
 a48217a <=( (not A202)  and  A201 );
 a48218a <=( A166  and  a48217a );
 a48219a <=( a48218a  and  a48213a );
 a48223a <=( A268  and  (not A267) );
 a48224a <=( (not A203)  and  a48223a );
 a48227a <=( A299  and  (not A298) );
 a48230a <=( A301  and  A300 );
 a48231a <=( a48230a  and  a48227a );
 a48232a <=( a48231a  and  a48224a );
 a48236a <=( (not A167)  and  A168 );
 a48237a <=( A169  and  a48236a );
 a48241a <=( (not A202)  and  A201 );
 a48242a <=( A166  and  a48241a );
 a48243a <=( a48242a  and  a48237a );
 a48247a <=( A268  and  (not A267) );
 a48248a <=( (not A203)  and  a48247a );
 a48251a <=( A299  and  (not A298) );
 a48254a <=( A302  and  A300 );
 a48255a <=( a48254a  and  a48251a );
 a48256a <=( a48255a  and  a48248a );
 a48260a <=( (not A167)  and  A168 );
 a48261a <=( A169  and  a48260a );
 a48265a <=( (not A202)  and  A201 );
 a48266a <=( A166  and  a48265a );
 a48267a <=( a48266a  and  a48261a );
 a48271a <=( A269  and  (not A267) );
 a48272a <=( (not A203)  and  a48271a );
 a48275a <=( (not A299)  and  A298 );
 a48278a <=( A301  and  A300 );
 a48279a <=( a48278a  and  a48275a );
 a48280a <=( a48279a  and  a48272a );
 a48284a <=( (not A167)  and  A168 );
 a48285a <=( A169  and  a48284a );
 a48289a <=( (not A202)  and  A201 );
 a48290a <=( A166  and  a48289a );
 a48291a <=( a48290a  and  a48285a );
 a48295a <=( A269  and  (not A267) );
 a48296a <=( (not A203)  and  a48295a );
 a48299a <=( (not A299)  and  A298 );
 a48302a <=( A302  and  A300 );
 a48303a <=( a48302a  and  a48299a );
 a48304a <=( a48303a  and  a48296a );
 a48308a <=( (not A167)  and  A168 );
 a48309a <=( A169  and  a48308a );
 a48313a <=( (not A202)  and  A201 );
 a48314a <=( A166  and  a48313a );
 a48315a <=( a48314a  and  a48309a );
 a48319a <=( A269  and  (not A267) );
 a48320a <=( (not A203)  and  a48319a );
 a48323a <=( A299  and  (not A298) );
 a48326a <=( A301  and  A300 );
 a48327a <=( a48326a  and  a48323a );
 a48328a <=( a48327a  and  a48320a );
 a48332a <=( (not A167)  and  A168 );
 a48333a <=( A169  and  a48332a );
 a48337a <=( (not A202)  and  A201 );
 a48338a <=( A166  and  a48337a );
 a48339a <=( a48338a  and  a48333a );
 a48343a <=( A269  and  (not A267) );
 a48344a <=( (not A203)  and  a48343a );
 a48347a <=( A299  and  (not A298) );
 a48350a <=( A302  and  A300 );
 a48351a <=( a48350a  and  a48347a );
 a48352a <=( a48351a  and  a48344a );
 a48356a <=( (not A167)  and  A168 );
 a48357a <=( A169  and  a48356a );
 a48361a <=( (not A202)  and  A201 );
 a48362a <=( A166  and  a48361a );
 a48363a <=( a48362a  and  a48357a );
 a48367a <=( A266  and  A265 );
 a48368a <=( (not A203)  and  a48367a );
 a48371a <=( (not A299)  and  A298 );
 a48374a <=( A301  and  A300 );
 a48375a <=( a48374a  and  a48371a );
 a48376a <=( a48375a  and  a48368a );
 a48380a <=( (not A167)  and  A168 );
 a48381a <=( A169  and  a48380a );
 a48385a <=( (not A202)  and  A201 );
 a48386a <=( A166  and  a48385a );
 a48387a <=( a48386a  and  a48381a );
 a48391a <=( A266  and  A265 );
 a48392a <=( (not A203)  and  a48391a );
 a48395a <=( (not A299)  and  A298 );
 a48398a <=( A302  and  A300 );
 a48399a <=( a48398a  and  a48395a );
 a48400a <=( a48399a  and  a48392a );
 a48404a <=( (not A167)  and  A168 );
 a48405a <=( A169  and  a48404a );
 a48409a <=( (not A202)  and  A201 );
 a48410a <=( A166  and  a48409a );
 a48411a <=( a48410a  and  a48405a );
 a48415a <=( A266  and  A265 );
 a48416a <=( (not A203)  and  a48415a );
 a48419a <=( A299  and  (not A298) );
 a48422a <=( A301  and  A300 );
 a48423a <=( a48422a  and  a48419a );
 a48424a <=( a48423a  and  a48416a );
 a48428a <=( (not A167)  and  A168 );
 a48429a <=( A169  and  a48428a );
 a48433a <=( (not A202)  and  A201 );
 a48434a <=( A166  and  a48433a );
 a48435a <=( a48434a  and  a48429a );
 a48439a <=( A266  and  A265 );
 a48440a <=( (not A203)  and  a48439a );
 a48443a <=( A299  and  (not A298) );
 a48446a <=( A302  and  A300 );
 a48447a <=( a48446a  and  a48443a );
 a48448a <=( a48447a  and  a48440a );
 a48452a <=( (not A167)  and  A168 );
 a48453a <=( A169  and  a48452a );
 a48457a <=( (not A202)  and  A201 );
 a48458a <=( A166  and  a48457a );
 a48459a <=( a48458a  and  a48453a );
 a48463a <=( (not A266)  and  (not A265) );
 a48464a <=( (not A203)  and  a48463a );
 a48467a <=( (not A299)  and  A298 );
 a48470a <=( A301  and  A300 );
 a48471a <=( a48470a  and  a48467a );
 a48472a <=( a48471a  and  a48464a );
 a48476a <=( (not A167)  and  A168 );
 a48477a <=( A169  and  a48476a );
 a48481a <=( (not A202)  and  A201 );
 a48482a <=( A166  and  a48481a );
 a48483a <=( a48482a  and  a48477a );
 a48487a <=( (not A266)  and  (not A265) );
 a48488a <=( (not A203)  and  a48487a );
 a48491a <=( (not A299)  and  A298 );
 a48494a <=( A302  and  A300 );
 a48495a <=( a48494a  and  a48491a );
 a48496a <=( a48495a  and  a48488a );
 a48500a <=( (not A167)  and  A168 );
 a48501a <=( A169  and  a48500a );
 a48505a <=( (not A202)  and  A201 );
 a48506a <=( A166  and  a48505a );
 a48507a <=( a48506a  and  a48501a );
 a48511a <=( (not A266)  and  (not A265) );
 a48512a <=( (not A203)  and  a48511a );
 a48515a <=( A299  and  (not A298) );
 a48518a <=( A301  and  A300 );
 a48519a <=( a48518a  and  a48515a );
 a48520a <=( a48519a  and  a48512a );
 a48524a <=( (not A167)  and  A168 );
 a48525a <=( A169  and  a48524a );
 a48529a <=( (not A202)  and  A201 );
 a48530a <=( A166  and  a48529a );
 a48531a <=( a48530a  and  a48525a );
 a48535a <=( (not A266)  and  (not A265) );
 a48536a <=( (not A203)  and  a48535a );
 a48539a <=( A299  and  (not A298) );
 a48542a <=( A302  and  A300 );
 a48543a <=( a48542a  and  a48539a );
 a48544a <=( a48543a  and  a48536a );
 a48548a <=( (not A167)  and  A168 );
 a48549a <=( A169  and  a48548a );
 a48553a <=( A202  and  (not A201) );
 a48554a <=( A166  and  a48553a );
 a48555a <=( a48554a  and  a48549a );
 a48559a <=( (not A269)  and  (not A268) );
 a48560a <=( A267  and  a48559a );
 a48563a <=( (not A299)  and  A298 );
 a48566a <=( A301  and  A300 );
 a48567a <=( a48566a  and  a48563a );
 a48568a <=( a48567a  and  a48560a );
 a48572a <=( (not A167)  and  A168 );
 a48573a <=( A169  and  a48572a );
 a48577a <=( A202  and  (not A201) );
 a48578a <=( A166  and  a48577a );
 a48579a <=( a48578a  and  a48573a );
 a48583a <=( (not A269)  and  (not A268) );
 a48584a <=( A267  and  a48583a );
 a48587a <=( (not A299)  and  A298 );
 a48590a <=( A302  and  A300 );
 a48591a <=( a48590a  and  a48587a );
 a48592a <=( a48591a  and  a48584a );
 a48596a <=( (not A167)  and  A168 );
 a48597a <=( A169  and  a48596a );
 a48601a <=( A202  and  (not A201) );
 a48602a <=( A166  and  a48601a );
 a48603a <=( a48602a  and  a48597a );
 a48607a <=( (not A269)  and  (not A268) );
 a48608a <=( A267  and  a48607a );
 a48611a <=( A299  and  (not A298) );
 a48614a <=( A301  and  A300 );
 a48615a <=( a48614a  and  a48611a );
 a48616a <=( a48615a  and  a48608a );
 a48620a <=( (not A167)  and  A168 );
 a48621a <=( A169  and  a48620a );
 a48625a <=( A202  and  (not A201) );
 a48626a <=( A166  and  a48625a );
 a48627a <=( a48626a  and  a48621a );
 a48631a <=( (not A269)  and  (not A268) );
 a48632a <=( A267  and  a48631a );
 a48635a <=( A299  and  (not A298) );
 a48638a <=( A302  and  A300 );
 a48639a <=( a48638a  and  a48635a );
 a48640a <=( a48639a  and  a48632a );
 a48644a <=( (not A167)  and  A168 );
 a48645a <=( A169  and  a48644a );
 a48649a <=( A202  and  (not A201) );
 a48650a <=( A166  and  a48649a );
 a48651a <=( a48650a  and  a48645a );
 a48655a <=( A298  and  A268 );
 a48656a <=( (not A267)  and  a48655a );
 a48659a <=( (not A300)  and  (not A299) );
 a48662a <=( (not A302)  and  (not A301) );
 a48663a <=( a48662a  and  a48659a );
 a48664a <=( a48663a  and  a48656a );
 a48668a <=( (not A167)  and  A168 );
 a48669a <=( A169  and  a48668a );
 a48673a <=( A202  and  (not A201) );
 a48674a <=( A166  and  a48673a );
 a48675a <=( a48674a  and  a48669a );
 a48679a <=( (not A298)  and  A268 );
 a48680a <=( (not A267)  and  a48679a );
 a48683a <=( (not A300)  and  A299 );
 a48686a <=( (not A302)  and  (not A301) );
 a48687a <=( a48686a  and  a48683a );
 a48688a <=( a48687a  and  a48680a );
 a48692a <=( (not A167)  and  A168 );
 a48693a <=( A169  and  a48692a );
 a48697a <=( A202  and  (not A201) );
 a48698a <=( A166  and  a48697a );
 a48699a <=( a48698a  and  a48693a );
 a48703a <=( A298  and  A269 );
 a48704a <=( (not A267)  and  a48703a );
 a48707a <=( (not A300)  and  (not A299) );
 a48710a <=( (not A302)  and  (not A301) );
 a48711a <=( a48710a  and  a48707a );
 a48712a <=( a48711a  and  a48704a );
 a48716a <=( (not A167)  and  A168 );
 a48717a <=( A169  and  a48716a );
 a48721a <=( A202  and  (not A201) );
 a48722a <=( A166  and  a48721a );
 a48723a <=( a48722a  and  a48717a );
 a48727a <=( (not A298)  and  A269 );
 a48728a <=( (not A267)  and  a48727a );
 a48731a <=( (not A300)  and  A299 );
 a48734a <=( (not A302)  and  (not A301) );
 a48735a <=( a48734a  and  a48731a );
 a48736a <=( a48735a  and  a48728a );
 a48740a <=( (not A167)  and  A168 );
 a48741a <=( A169  and  a48740a );
 a48745a <=( A202  and  (not A201) );
 a48746a <=( A166  and  a48745a );
 a48747a <=( a48746a  and  a48741a );
 a48751a <=( A298  and  A266 );
 a48752a <=( A265  and  a48751a );
 a48755a <=( (not A300)  and  (not A299) );
 a48758a <=( (not A302)  and  (not A301) );
 a48759a <=( a48758a  and  a48755a );
 a48760a <=( a48759a  and  a48752a );
 a48764a <=( (not A167)  and  A168 );
 a48765a <=( A169  and  a48764a );
 a48769a <=( A202  and  (not A201) );
 a48770a <=( A166  and  a48769a );
 a48771a <=( a48770a  and  a48765a );
 a48775a <=( (not A298)  and  A266 );
 a48776a <=( A265  and  a48775a );
 a48779a <=( (not A300)  and  A299 );
 a48782a <=( (not A302)  and  (not A301) );
 a48783a <=( a48782a  and  a48779a );
 a48784a <=( a48783a  and  a48776a );
 a48788a <=( (not A167)  and  A168 );
 a48789a <=( A169  and  a48788a );
 a48793a <=( A202  and  (not A201) );
 a48794a <=( A166  and  a48793a );
 a48795a <=( a48794a  and  a48789a );
 a48799a <=( A298  and  (not A266) );
 a48800a <=( (not A265)  and  a48799a );
 a48803a <=( (not A300)  and  (not A299) );
 a48806a <=( (not A302)  and  (not A301) );
 a48807a <=( a48806a  and  a48803a );
 a48808a <=( a48807a  and  a48800a );
 a48812a <=( (not A167)  and  A168 );
 a48813a <=( A169  and  a48812a );
 a48817a <=( A202  and  (not A201) );
 a48818a <=( A166  and  a48817a );
 a48819a <=( a48818a  and  a48813a );
 a48823a <=( (not A298)  and  (not A266) );
 a48824a <=( (not A265)  and  a48823a );
 a48827a <=( (not A300)  and  A299 );
 a48830a <=( (not A302)  and  (not A301) );
 a48831a <=( a48830a  and  a48827a );
 a48832a <=( a48831a  and  a48824a );
 a48836a <=( (not A167)  and  A168 );
 a48837a <=( A169  and  a48836a );
 a48841a <=( A203  and  (not A201) );
 a48842a <=( A166  and  a48841a );
 a48843a <=( a48842a  and  a48837a );
 a48847a <=( (not A269)  and  (not A268) );
 a48848a <=( A267  and  a48847a );
 a48851a <=( (not A299)  and  A298 );
 a48854a <=( A301  and  A300 );
 a48855a <=( a48854a  and  a48851a );
 a48856a <=( a48855a  and  a48848a );
 a48860a <=( (not A167)  and  A168 );
 a48861a <=( A169  and  a48860a );
 a48865a <=( A203  and  (not A201) );
 a48866a <=( A166  and  a48865a );
 a48867a <=( a48866a  and  a48861a );
 a48871a <=( (not A269)  and  (not A268) );
 a48872a <=( A267  and  a48871a );
 a48875a <=( (not A299)  and  A298 );
 a48878a <=( A302  and  A300 );
 a48879a <=( a48878a  and  a48875a );
 a48880a <=( a48879a  and  a48872a );
 a48884a <=( (not A167)  and  A168 );
 a48885a <=( A169  and  a48884a );
 a48889a <=( A203  and  (not A201) );
 a48890a <=( A166  and  a48889a );
 a48891a <=( a48890a  and  a48885a );
 a48895a <=( (not A269)  and  (not A268) );
 a48896a <=( A267  and  a48895a );
 a48899a <=( A299  and  (not A298) );
 a48902a <=( A301  and  A300 );
 a48903a <=( a48902a  and  a48899a );
 a48904a <=( a48903a  and  a48896a );
 a48908a <=( (not A167)  and  A168 );
 a48909a <=( A169  and  a48908a );
 a48913a <=( A203  and  (not A201) );
 a48914a <=( A166  and  a48913a );
 a48915a <=( a48914a  and  a48909a );
 a48919a <=( (not A269)  and  (not A268) );
 a48920a <=( A267  and  a48919a );
 a48923a <=( A299  and  (not A298) );
 a48926a <=( A302  and  A300 );
 a48927a <=( a48926a  and  a48923a );
 a48928a <=( a48927a  and  a48920a );
 a48932a <=( (not A167)  and  A168 );
 a48933a <=( A169  and  a48932a );
 a48937a <=( A203  and  (not A201) );
 a48938a <=( A166  and  a48937a );
 a48939a <=( a48938a  and  a48933a );
 a48943a <=( A298  and  A268 );
 a48944a <=( (not A267)  and  a48943a );
 a48947a <=( (not A300)  and  (not A299) );
 a48950a <=( (not A302)  and  (not A301) );
 a48951a <=( a48950a  and  a48947a );
 a48952a <=( a48951a  and  a48944a );
 a48956a <=( (not A167)  and  A168 );
 a48957a <=( A169  and  a48956a );
 a48961a <=( A203  and  (not A201) );
 a48962a <=( A166  and  a48961a );
 a48963a <=( a48962a  and  a48957a );
 a48967a <=( (not A298)  and  A268 );
 a48968a <=( (not A267)  and  a48967a );
 a48971a <=( (not A300)  and  A299 );
 a48974a <=( (not A302)  and  (not A301) );
 a48975a <=( a48974a  and  a48971a );
 a48976a <=( a48975a  and  a48968a );
 a48980a <=( (not A167)  and  A168 );
 a48981a <=( A169  and  a48980a );
 a48985a <=( A203  and  (not A201) );
 a48986a <=( A166  and  a48985a );
 a48987a <=( a48986a  and  a48981a );
 a48991a <=( A298  and  A269 );
 a48992a <=( (not A267)  and  a48991a );
 a48995a <=( (not A300)  and  (not A299) );
 a48998a <=( (not A302)  and  (not A301) );
 a48999a <=( a48998a  and  a48995a );
 a49000a <=( a48999a  and  a48992a );
 a49004a <=( (not A167)  and  A168 );
 a49005a <=( A169  and  a49004a );
 a49009a <=( A203  and  (not A201) );
 a49010a <=( A166  and  a49009a );
 a49011a <=( a49010a  and  a49005a );
 a49015a <=( (not A298)  and  A269 );
 a49016a <=( (not A267)  and  a49015a );
 a49019a <=( (not A300)  and  A299 );
 a49022a <=( (not A302)  and  (not A301) );
 a49023a <=( a49022a  and  a49019a );
 a49024a <=( a49023a  and  a49016a );
 a49028a <=( (not A167)  and  A168 );
 a49029a <=( A169  and  a49028a );
 a49033a <=( A203  and  (not A201) );
 a49034a <=( A166  and  a49033a );
 a49035a <=( a49034a  and  a49029a );
 a49039a <=( A298  and  A266 );
 a49040a <=( A265  and  a49039a );
 a49043a <=( (not A300)  and  (not A299) );
 a49046a <=( (not A302)  and  (not A301) );
 a49047a <=( a49046a  and  a49043a );
 a49048a <=( a49047a  and  a49040a );
 a49052a <=( (not A167)  and  A168 );
 a49053a <=( A169  and  a49052a );
 a49057a <=( A203  and  (not A201) );
 a49058a <=( A166  and  a49057a );
 a49059a <=( a49058a  and  a49053a );
 a49063a <=( (not A298)  and  A266 );
 a49064a <=( A265  and  a49063a );
 a49067a <=( (not A300)  and  A299 );
 a49070a <=( (not A302)  and  (not A301) );
 a49071a <=( a49070a  and  a49067a );
 a49072a <=( a49071a  and  a49064a );
 a49076a <=( (not A167)  and  A168 );
 a49077a <=( A169  and  a49076a );
 a49081a <=( A203  and  (not A201) );
 a49082a <=( A166  and  a49081a );
 a49083a <=( a49082a  and  a49077a );
 a49087a <=( A298  and  (not A266) );
 a49088a <=( (not A265)  and  a49087a );
 a49091a <=( (not A300)  and  (not A299) );
 a49094a <=( (not A302)  and  (not A301) );
 a49095a <=( a49094a  and  a49091a );
 a49096a <=( a49095a  and  a49088a );
 a49100a <=( (not A167)  and  A168 );
 a49101a <=( A169  and  a49100a );
 a49105a <=( A203  and  (not A201) );
 a49106a <=( A166  and  a49105a );
 a49107a <=( a49106a  and  a49101a );
 a49111a <=( (not A298)  and  (not A266) );
 a49112a <=( (not A265)  and  a49111a );
 a49115a <=( (not A300)  and  A299 );
 a49118a <=( (not A302)  and  (not A301) );
 a49119a <=( a49118a  and  a49115a );
 a49120a <=( a49119a  and  a49112a );
 a49124a <=( (not A167)  and  A168 );
 a49125a <=( A169  and  a49124a );
 a49129a <=( A200  and  A199 );
 a49130a <=( A166  and  a49129a );
 a49131a <=( a49130a  and  a49125a );
 a49135a <=( (not A269)  and  (not A268) );
 a49136a <=( A267  and  a49135a );
 a49139a <=( (not A299)  and  A298 );
 a49142a <=( A301  and  A300 );
 a49143a <=( a49142a  and  a49139a );
 a49144a <=( a49143a  and  a49136a );
 a49148a <=( (not A167)  and  A168 );
 a49149a <=( A169  and  a49148a );
 a49153a <=( A200  and  A199 );
 a49154a <=( A166  and  a49153a );
 a49155a <=( a49154a  and  a49149a );
 a49159a <=( (not A269)  and  (not A268) );
 a49160a <=( A267  and  a49159a );
 a49163a <=( (not A299)  and  A298 );
 a49166a <=( A302  and  A300 );
 a49167a <=( a49166a  and  a49163a );
 a49168a <=( a49167a  and  a49160a );
 a49172a <=( (not A167)  and  A168 );
 a49173a <=( A169  and  a49172a );
 a49177a <=( A200  and  A199 );
 a49178a <=( A166  and  a49177a );
 a49179a <=( a49178a  and  a49173a );
 a49183a <=( (not A269)  and  (not A268) );
 a49184a <=( A267  and  a49183a );
 a49187a <=( A299  and  (not A298) );
 a49190a <=( A301  and  A300 );
 a49191a <=( a49190a  and  a49187a );
 a49192a <=( a49191a  and  a49184a );
 a49196a <=( (not A167)  and  A168 );
 a49197a <=( A169  and  a49196a );
 a49201a <=( A200  and  A199 );
 a49202a <=( A166  and  a49201a );
 a49203a <=( a49202a  and  a49197a );
 a49207a <=( (not A269)  and  (not A268) );
 a49208a <=( A267  and  a49207a );
 a49211a <=( A299  and  (not A298) );
 a49214a <=( A302  and  A300 );
 a49215a <=( a49214a  and  a49211a );
 a49216a <=( a49215a  and  a49208a );
 a49220a <=( (not A167)  and  A168 );
 a49221a <=( A169  and  a49220a );
 a49225a <=( A200  and  A199 );
 a49226a <=( A166  and  a49225a );
 a49227a <=( a49226a  and  a49221a );
 a49231a <=( A298  and  A268 );
 a49232a <=( (not A267)  and  a49231a );
 a49235a <=( (not A300)  and  (not A299) );
 a49238a <=( (not A302)  and  (not A301) );
 a49239a <=( a49238a  and  a49235a );
 a49240a <=( a49239a  and  a49232a );
 a49244a <=( (not A167)  and  A168 );
 a49245a <=( A169  and  a49244a );
 a49249a <=( A200  and  A199 );
 a49250a <=( A166  and  a49249a );
 a49251a <=( a49250a  and  a49245a );
 a49255a <=( (not A298)  and  A268 );
 a49256a <=( (not A267)  and  a49255a );
 a49259a <=( (not A300)  and  A299 );
 a49262a <=( (not A302)  and  (not A301) );
 a49263a <=( a49262a  and  a49259a );
 a49264a <=( a49263a  and  a49256a );
 a49268a <=( (not A167)  and  A168 );
 a49269a <=( A169  and  a49268a );
 a49273a <=( A200  and  A199 );
 a49274a <=( A166  and  a49273a );
 a49275a <=( a49274a  and  a49269a );
 a49279a <=( A298  and  A269 );
 a49280a <=( (not A267)  and  a49279a );
 a49283a <=( (not A300)  and  (not A299) );
 a49286a <=( (not A302)  and  (not A301) );
 a49287a <=( a49286a  and  a49283a );
 a49288a <=( a49287a  and  a49280a );
 a49292a <=( (not A167)  and  A168 );
 a49293a <=( A169  and  a49292a );
 a49297a <=( A200  and  A199 );
 a49298a <=( A166  and  a49297a );
 a49299a <=( a49298a  and  a49293a );
 a49303a <=( (not A298)  and  A269 );
 a49304a <=( (not A267)  and  a49303a );
 a49307a <=( (not A300)  and  A299 );
 a49310a <=( (not A302)  and  (not A301) );
 a49311a <=( a49310a  and  a49307a );
 a49312a <=( a49311a  and  a49304a );
 a49316a <=( (not A167)  and  A168 );
 a49317a <=( A169  and  a49316a );
 a49321a <=( A200  and  A199 );
 a49322a <=( A166  and  a49321a );
 a49323a <=( a49322a  and  a49317a );
 a49327a <=( A298  and  A266 );
 a49328a <=( A265  and  a49327a );
 a49331a <=( (not A300)  and  (not A299) );
 a49334a <=( (not A302)  and  (not A301) );
 a49335a <=( a49334a  and  a49331a );
 a49336a <=( a49335a  and  a49328a );
 a49340a <=( (not A167)  and  A168 );
 a49341a <=( A169  and  a49340a );
 a49345a <=( A200  and  A199 );
 a49346a <=( A166  and  a49345a );
 a49347a <=( a49346a  and  a49341a );
 a49351a <=( (not A298)  and  A266 );
 a49352a <=( A265  and  a49351a );
 a49355a <=( (not A300)  and  A299 );
 a49358a <=( (not A302)  and  (not A301) );
 a49359a <=( a49358a  and  a49355a );
 a49360a <=( a49359a  and  a49352a );
 a49364a <=( (not A167)  and  A168 );
 a49365a <=( A169  and  a49364a );
 a49369a <=( A200  and  A199 );
 a49370a <=( A166  and  a49369a );
 a49371a <=( a49370a  and  a49365a );
 a49375a <=( A298  and  (not A266) );
 a49376a <=( (not A265)  and  a49375a );
 a49379a <=( (not A300)  and  (not A299) );
 a49382a <=( (not A302)  and  (not A301) );
 a49383a <=( a49382a  and  a49379a );
 a49384a <=( a49383a  and  a49376a );
 a49388a <=( (not A167)  and  A168 );
 a49389a <=( A169  and  a49388a );
 a49393a <=( A200  and  A199 );
 a49394a <=( A166  and  a49393a );
 a49395a <=( a49394a  and  a49389a );
 a49399a <=( (not A298)  and  (not A266) );
 a49400a <=( (not A265)  and  a49399a );
 a49403a <=( (not A300)  and  A299 );
 a49406a <=( (not A302)  and  (not A301) );
 a49407a <=( a49406a  and  a49403a );
 a49408a <=( a49407a  and  a49400a );
 a49412a <=( (not A167)  and  A168 );
 a49413a <=( A169  and  a49412a );
 a49417a <=( (not A200)  and  (not A199) );
 a49418a <=( A166  and  a49417a );
 a49419a <=( a49418a  and  a49413a );
 a49423a <=( (not A269)  and  (not A268) );
 a49424a <=( A267  and  a49423a );
 a49427a <=( (not A299)  and  A298 );
 a49430a <=( A301  and  A300 );
 a49431a <=( a49430a  and  a49427a );
 a49432a <=( a49431a  and  a49424a );
 a49436a <=( (not A167)  and  A168 );
 a49437a <=( A169  and  a49436a );
 a49441a <=( (not A200)  and  (not A199) );
 a49442a <=( A166  and  a49441a );
 a49443a <=( a49442a  and  a49437a );
 a49447a <=( (not A269)  and  (not A268) );
 a49448a <=( A267  and  a49447a );
 a49451a <=( (not A299)  and  A298 );
 a49454a <=( A302  and  A300 );
 a49455a <=( a49454a  and  a49451a );
 a49456a <=( a49455a  and  a49448a );
 a49460a <=( (not A167)  and  A168 );
 a49461a <=( A169  and  a49460a );
 a49465a <=( (not A200)  and  (not A199) );
 a49466a <=( A166  and  a49465a );
 a49467a <=( a49466a  and  a49461a );
 a49471a <=( (not A269)  and  (not A268) );
 a49472a <=( A267  and  a49471a );
 a49475a <=( A299  and  (not A298) );
 a49478a <=( A301  and  A300 );
 a49479a <=( a49478a  and  a49475a );
 a49480a <=( a49479a  and  a49472a );
 a49484a <=( (not A167)  and  A168 );
 a49485a <=( A169  and  a49484a );
 a49489a <=( (not A200)  and  (not A199) );
 a49490a <=( A166  and  a49489a );
 a49491a <=( a49490a  and  a49485a );
 a49495a <=( (not A269)  and  (not A268) );
 a49496a <=( A267  and  a49495a );
 a49499a <=( A299  and  (not A298) );
 a49502a <=( A302  and  A300 );
 a49503a <=( a49502a  and  a49499a );
 a49504a <=( a49503a  and  a49496a );
 a49508a <=( (not A167)  and  A168 );
 a49509a <=( A169  and  a49508a );
 a49513a <=( (not A200)  and  (not A199) );
 a49514a <=( A166  and  a49513a );
 a49515a <=( a49514a  and  a49509a );
 a49519a <=( A298  and  A268 );
 a49520a <=( (not A267)  and  a49519a );
 a49523a <=( (not A300)  and  (not A299) );
 a49526a <=( (not A302)  and  (not A301) );
 a49527a <=( a49526a  and  a49523a );
 a49528a <=( a49527a  and  a49520a );
 a49532a <=( (not A167)  and  A168 );
 a49533a <=( A169  and  a49532a );
 a49537a <=( (not A200)  and  (not A199) );
 a49538a <=( A166  and  a49537a );
 a49539a <=( a49538a  and  a49533a );
 a49543a <=( (not A298)  and  A268 );
 a49544a <=( (not A267)  and  a49543a );
 a49547a <=( (not A300)  and  A299 );
 a49550a <=( (not A302)  and  (not A301) );
 a49551a <=( a49550a  and  a49547a );
 a49552a <=( a49551a  and  a49544a );
 a49556a <=( (not A167)  and  A168 );
 a49557a <=( A169  and  a49556a );
 a49561a <=( (not A200)  and  (not A199) );
 a49562a <=( A166  and  a49561a );
 a49563a <=( a49562a  and  a49557a );
 a49567a <=( A298  and  A269 );
 a49568a <=( (not A267)  and  a49567a );
 a49571a <=( (not A300)  and  (not A299) );
 a49574a <=( (not A302)  and  (not A301) );
 a49575a <=( a49574a  and  a49571a );
 a49576a <=( a49575a  and  a49568a );
 a49580a <=( (not A167)  and  A168 );
 a49581a <=( A169  and  a49580a );
 a49585a <=( (not A200)  and  (not A199) );
 a49586a <=( A166  and  a49585a );
 a49587a <=( a49586a  and  a49581a );
 a49591a <=( (not A298)  and  A269 );
 a49592a <=( (not A267)  and  a49591a );
 a49595a <=( (not A300)  and  A299 );
 a49598a <=( (not A302)  and  (not A301) );
 a49599a <=( a49598a  and  a49595a );
 a49600a <=( a49599a  and  a49592a );
 a49604a <=( (not A167)  and  A168 );
 a49605a <=( A169  and  a49604a );
 a49609a <=( (not A200)  and  (not A199) );
 a49610a <=( A166  and  a49609a );
 a49611a <=( a49610a  and  a49605a );
 a49615a <=( A298  and  A266 );
 a49616a <=( A265  and  a49615a );
 a49619a <=( (not A300)  and  (not A299) );
 a49622a <=( (not A302)  and  (not A301) );
 a49623a <=( a49622a  and  a49619a );
 a49624a <=( a49623a  and  a49616a );
 a49628a <=( (not A167)  and  A168 );
 a49629a <=( A169  and  a49628a );
 a49633a <=( (not A200)  and  (not A199) );
 a49634a <=( A166  and  a49633a );
 a49635a <=( a49634a  and  a49629a );
 a49639a <=( (not A298)  and  A266 );
 a49640a <=( A265  and  a49639a );
 a49643a <=( (not A300)  and  A299 );
 a49646a <=( (not A302)  and  (not A301) );
 a49647a <=( a49646a  and  a49643a );
 a49648a <=( a49647a  and  a49640a );
 a49652a <=( (not A167)  and  A168 );
 a49653a <=( A169  and  a49652a );
 a49657a <=( (not A200)  and  (not A199) );
 a49658a <=( A166  and  a49657a );
 a49659a <=( a49658a  and  a49653a );
 a49663a <=( A298  and  (not A266) );
 a49664a <=( (not A265)  and  a49663a );
 a49667a <=( (not A300)  and  (not A299) );
 a49670a <=( (not A302)  and  (not A301) );
 a49671a <=( a49670a  and  a49667a );
 a49672a <=( a49671a  and  a49664a );
 a49676a <=( (not A167)  and  A168 );
 a49677a <=( A169  and  a49676a );
 a49681a <=( (not A200)  and  (not A199) );
 a49682a <=( A166  and  a49681a );
 a49683a <=( a49682a  and  a49677a );
 a49687a <=( (not A298)  and  (not A266) );
 a49688a <=( (not A265)  and  a49687a );
 a49691a <=( (not A300)  and  A299 );
 a49694a <=( (not A302)  and  (not A301) );
 a49695a <=( a49694a  and  a49691a );
 a49696a <=( a49695a  and  a49688a );
 a49700a <=( A201  and  (not A168) );
 a49701a <=( A169  and  a49700a );
 a49705a <=( (not A265)  and  (not A203) );
 a49706a <=( (not A202)  and  a49705a );
 a49707a <=( a49706a  and  a49701a );
 a49711a <=( (not A268)  and  (not A267) );
 a49712a <=( A266  and  a49711a );
 a49715a <=( A300  and  (not A269) );
 a49718a <=( (not A302)  and  (not A301) );
 a49719a <=( a49718a  and  a49715a );
 a49720a <=( a49719a  and  a49712a );
 a49724a <=( A201  and  (not A168) );
 a49725a <=( A169  and  a49724a );
 a49729a <=( A265  and  (not A203) );
 a49730a <=( (not A202)  and  a49729a );
 a49731a <=( a49730a  and  a49725a );
 a49735a <=( (not A268)  and  (not A267) );
 a49736a <=( (not A266)  and  a49735a );
 a49739a <=( A300  and  (not A269) );
 a49742a <=( (not A302)  and  (not A301) );
 a49743a <=( a49742a  and  a49739a );
 a49744a <=( a49743a  and  a49736a );
 a49748a <=( (not A199)  and  (not A168) );
 a49749a <=( A169  and  a49748a );
 a49753a <=( A202  and  A201 );
 a49754a <=( A200  and  a49753a );
 a49755a <=( a49754a  and  a49749a );
 a49759a <=( (not A269)  and  (not A268) );
 a49760a <=( A267  and  a49759a );
 a49763a <=( (not A299)  and  A298 );
 a49766a <=( A301  and  A300 );
 a49767a <=( a49766a  and  a49763a );
 a49768a <=( a49767a  and  a49760a );
 a49772a <=( (not A199)  and  (not A168) );
 a49773a <=( A169  and  a49772a );
 a49777a <=( A202  and  A201 );
 a49778a <=( A200  and  a49777a );
 a49779a <=( a49778a  and  a49773a );
 a49783a <=( (not A269)  and  (not A268) );
 a49784a <=( A267  and  a49783a );
 a49787a <=( (not A299)  and  A298 );
 a49790a <=( A302  and  A300 );
 a49791a <=( a49790a  and  a49787a );
 a49792a <=( a49791a  and  a49784a );
 a49796a <=( (not A199)  and  (not A168) );
 a49797a <=( A169  and  a49796a );
 a49801a <=( A202  and  A201 );
 a49802a <=( A200  and  a49801a );
 a49803a <=( a49802a  and  a49797a );
 a49807a <=( (not A269)  and  (not A268) );
 a49808a <=( A267  and  a49807a );
 a49811a <=( A299  and  (not A298) );
 a49814a <=( A301  and  A300 );
 a49815a <=( a49814a  and  a49811a );
 a49816a <=( a49815a  and  a49808a );
 a49820a <=( (not A199)  and  (not A168) );
 a49821a <=( A169  and  a49820a );
 a49825a <=( A202  and  A201 );
 a49826a <=( A200  and  a49825a );
 a49827a <=( a49826a  and  a49821a );
 a49831a <=( (not A269)  and  (not A268) );
 a49832a <=( A267  and  a49831a );
 a49835a <=( A299  and  (not A298) );
 a49838a <=( A302  and  A300 );
 a49839a <=( a49838a  and  a49835a );
 a49840a <=( a49839a  and  a49832a );
 a49844a <=( (not A199)  and  (not A168) );
 a49845a <=( A169  and  a49844a );
 a49849a <=( A202  and  A201 );
 a49850a <=( A200  and  a49849a );
 a49851a <=( a49850a  and  a49845a );
 a49855a <=( A298  and  A268 );
 a49856a <=( (not A267)  and  a49855a );
 a49859a <=( (not A300)  and  (not A299) );
 a49862a <=( (not A302)  and  (not A301) );
 a49863a <=( a49862a  and  a49859a );
 a49864a <=( a49863a  and  a49856a );
 a49868a <=( (not A199)  and  (not A168) );
 a49869a <=( A169  and  a49868a );
 a49873a <=( A202  and  A201 );
 a49874a <=( A200  and  a49873a );
 a49875a <=( a49874a  and  a49869a );
 a49879a <=( (not A298)  and  A268 );
 a49880a <=( (not A267)  and  a49879a );
 a49883a <=( (not A300)  and  A299 );
 a49886a <=( (not A302)  and  (not A301) );
 a49887a <=( a49886a  and  a49883a );
 a49888a <=( a49887a  and  a49880a );
 a49892a <=( (not A199)  and  (not A168) );
 a49893a <=( A169  and  a49892a );
 a49897a <=( A202  and  A201 );
 a49898a <=( A200  and  a49897a );
 a49899a <=( a49898a  and  a49893a );
 a49903a <=( A298  and  A269 );
 a49904a <=( (not A267)  and  a49903a );
 a49907a <=( (not A300)  and  (not A299) );
 a49910a <=( (not A302)  and  (not A301) );
 a49911a <=( a49910a  and  a49907a );
 a49912a <=( a49911a  and  a49904a );
 a49916a <=( (not A199)  and  (not A168) );
 a49917a <=( A169  and  a49916a );
 a49921a <=( A202  and  A201 );
 a49922a <=( A200  and  a49921a );
 a49923a <=( a49922a  and  a49917a );
 a49927a <=( (not A298)  and  A269 );
 a49928a <=( (not A267)  and  a49927a );
 a49931a <=( (not A300)  and  A299 );
 a49934a <=( (not A302)  and  (not A301) );
 a49935a <=( a49934a  and  a49931a );
 a49936a <=( a49935a  and  a49928a );
 a49940a <=( (not A199)  and  (not A168) );
 a49941a <=( A169  and  a49940a );
 a49945a <=( A202  and  A201 );
 a49946a <=( A200  and  a49945a );
 a49947a <=( a49946a  and  a49941a );
 a49951a <=( A298  and  A266 );
 a49952a <=( A265  and  a49951a );
 a49955a <=( (not A300)  and  (not A299) );
 a49958a <=( (not A302)  and  (not A301) );
 a49959a <=( a49958a  and  a49955a );
 a49960a <=( a49959a  and  a49952a );
 a49964a <=( (not A199)  and  (not A168) );
 a49965a <=( A169  and  a49964a );
 a49969a <=( A202  and  A201 );
 a49970a <=( A200  and  a49969a );
 a49971a <=( a49970a  and  a49965a );
 a49975a <=( (not A298)  and  A266 );
 a49976a <=( A265  and  a49975a );
 a49979a <=( (not A300)  and  A299 );
 a49982a <=( (not A302)  and  (not A301) );
 a49983a <=( a49982a  and  a49979a );
 a49984a <=( a49983a  and  a49976a );
 a49988a <=( (not A199)  and  (not A168) );
 a49989a <=( A169  and  a49988a );
 a49993a <=( A202  and  A201 );
 a49994a <=( A200  and  a49993a );
 a49995a <=( a49994a  and  a49989a );
 a49999a <=( A298  and  (not A266) );
 a50000a <=( (not A265)  and  a49999a );
 a50003a <=( (not A300)  and  (not A299) );
 a50006a <=( (not A302)  and  (not A301) );
 a50007a <=( a50006a  and  a50003a );
 a50008a <=( a50007a  and  a50000a );
 a50012a <=( (not A199)  and  (not A168) );
 a50013a <=( A169  and  a50012a );
 a50017a <=( A202  and  A201 );
 a50018a <=( A200  and  a50017a );
 a50019a <=( a50018a  and  a50013a );
 a50023a <=( (not A298)  and  (not A266) );
 a50024a <=( (not A265)  and  a50023a );
 a50027a <=( (not A300)  and  A299 );
 a50030a <=( (not A302)  and  (not A301) );
 a50031a <=( a50030a  and  a50027a );
 a50032a <=( a50031a  and  a50024a );
 a50036a <=( (not A199)  and  (not A168) );
 a50037a <=( A169  and  a50036a );
 a50041a <=( A203  and  A201 );
 a50042a <=( A200  and  a50041a );
 a50043a <=( a50042a  and  a50037a );
 a50047a <=( (not A269)  and  (not A268) );
 a50048a <=( A267  and  a50047a );
 a50051a <=( (not A299)  and  A298 );
 a50054a <=( A301  and  A300 );
 a50055a <=( a50054a  and  a50051a );
 a50056a <=( a50055a  and  a50048a );
 a50060a <=( (not A199)  and  (not A168) );
 a50061a <=( A169  and  a50060a );
 a50065a <=( A203  and  A201 );
 a50066a <=( A200  and  a50065a );
 a50067a <=( a50066a  and  a50061a );
 a50071a <=( (not A269)  and  (not A268) );
 a50072a <=( A267  and  a50071a );
 a50075a <=( (not A299)  and  A298 );
 a50078a <=( A302  and  A300 );
 a50079a <=( a50078a  and  a50075a );
 a50080a <=( a50079a  and  a50072a );
 a50084a <=( (not A199)  and  (not A168) );
 a50085a <=( A169  and  a50084a );
 a50089a <=( A203  and  A201 );
 a50090a <=( A200  and  a50089a );
 a50091a <=( a50090a  and  a50085a );
 a50095a <=( (not A269)  and  (not A268) );
 a50096a <=( A267  and  a50095a );
 a50099a <=( A299  and  (not A298) );
 a50102a <=( A301  and  A300 );
 a50103a <=( a50102a  and  a50099a );
 a50104a <=( a50103a  and  a50096a );
 a50108a <=( (not A199)  and  (not A168) );
 a50109a <=( A169  and  a50108a );
 a50113a <=( A203  and  A201 );
 a50114a <=( A200  and  a50113a );
 a50115a <=( a50114a  and  a50109a );
 a50119a <=( (not A269)  and  (not A268) );
 a50120a <=( A267  and  a50119a );
 a50123a <=( A299  and  (not A298) );
 a50126a <=( A302  and  A300 );
 a50127a <=( a50126a  and  a50123a );
 a50128a <=( a50127a  and  a50120a );
 a50132a <=( (not A199)  and  (not A168) );
 a50133a <=( A169  and  a50132a );
 a50137a <=( A203  and  A201 );
 a50138a <=( A200  and  a50137a );
 a50139a <=( a50138a  and  a50133a );
 a50143a <=( A298  and  A268 );
 a50144a <=( (not A267)  and  a50143a );
 a50147a <=( (not A300)  and  (not A299) );
 a50150a <=( (not A302)  and  (not A301) );
 a50151a <=( a50150a  and  a50147a );
 a50152a <=( a50151a  and  a50144a );
 a50156a <=( (not A199)  and  (not A168) );
 a50157a <=( A169  and  a50156a );
 a50161a <=( A203  and  A201 );
 a50162a <=( A200  and  a50161a );
 a50163a <=( a50162a  and  a50157a );
 a50167a <=( (not A298)  and  A268 );
 a50168a <=( (not A267)  and  a50167a );
 a50171a <=( (not A300)  and  A299 );
 a50174a <=( (not A302)  and  (not A301) );
 a50175a <=( a50174a  and  a50171a );
 a50176a <=( a50175a  and  a50168a );
 a50180a <=( (not A199)  and  (not A168) );
 a50181a <=( A169  and  a50180a );
 a50185a <=( A203  and  A201 );
 a50186a <=( A200  and  a50185a );
 a50187a <=( a50186a  and  a50181a );
 a50191a <=( A298  and  A269 );
 a50192a <=( (not A267)  and  a50191a );
 a50195a <=( (not A300)  and  (not A299) );
 a50198a <=( (not A302)  and  (not A301) );
 a50199a <=( a50198a  and  a50195a );
 a50200a <=( a50199a  and  a50192a );
 a50204a <=( (not A199)  and  (not A168) );
 a50205a <=( A169  and  a50204a );
 a50209a <=( A203  and  A201 );
 a50210a <=( A200  and  a50209a );
 a50211a <=( a50210a  and  a50205a );
 a50215a <=( (not A298)  and  A269 );
 a50216a <=( (not A267)  and  a50215a );
 a50219a <=( (not A300)  and  A299 );
 a50222a <=( (not A302)  and  (not A301) );
 a50223a <=( a50222a  and  a50219a );
 a50224a <=( a50223a  and  a50216a );
 a50228a <=( (not A199)  and  (not A168) );
 a50229a <=( A169  and  a50228a );
 a50233a <=( A203  and  A201 );
 a50234a <=( A200  and  a50233a );
 a50235a <=( a50234a  and  a50229a );
 a50239a <=( A298  and  A266 );
 a50240a <=( A265  and  a50239a );
 a50243a <=( (not A300)  and  (not A299) );
 a50246a <=( (not A302)  and  (not A301) );
 a50247a <=( a50246a  and  a50243a );
 a50248a <=( a50247a  and  a50240a );
 a50252a <=( (not A199)  and  (not A168) );
 a50253a <=( A169  and  a50252a );
 a50257a <=( A203  and  A201 );
 a50258a <=( A200  and  a50257a );
 a50259a <=( a50258a  and  a50253a );
 a50263a <=( (not A298)  and  A266 );
 a50264a <=( A265  and  a50263a );
 a50267a <=( (not A300)  and  A299 );
 a50270a <=( (not A302)  and  (not A301) );
 a50271a <=( a50270a  and  a50267a );
 a50272a <=( a50271a  and  a50264a );
 a50276a <=( (not A199)  and  (not A168) );
 a50277a <=( A169  and  a50276a );
 a50281a <=( A203  and  A201 );
 a50282a <=( A200  and  a50281a );
 a50283a <=( a50282a  and  a50277a );
 a50287a <=( A298  and  (not A266) );
 a50288a <=( (not A265)  and  a50287a );
 a50291a <=( (not A300)  and  (not A299) );
 a50294a <=( (not A302)  and  (not A301) );
 a50295a <=( a50294a  and  a50291a );
 a50296a <=( a50295a  and  a50288a );
 a50300a <=( (not A199)  and  (not A168) );
 a50301a <=( A169  and  a50300a );
 a50305a <=( A203  and  A201 );
 a50306a <=( A200  and  a50305a );
 a50307a <=( a50306a  and  a50301a );
 a50311a <=( (not A298)  and  (not A266) );
 a50312a <=( (not A265)  and  a50311a );
 a50315a <=( (not A300)  and  A299 );
 a50318a <=( (not A302)  and  (not A301) );
 a50319a <=( a50318a  and  a50315a );
 a50320a <=( a50319a  and  a50312a );
 a50324a <=( (not A199)  and  (not A168) );
 a50325a <=( A169  and  a50324a );
 a50329a <=( (not A202)  and  (not A201) );
 a50330a <=( A200  and  a50329a );
 a50331a <=( a50330a  and  a50325a );
 a50335a <=( A268  and  (not A267) );
 a50336a <=( (not A203)  and  a50335a );
 a50339a <=( (not A299)  and  A298 );
 a50342a <=( A301  and  A300 );
 a50343a <=( a50342a  and  a50339a );
 a50344a <=( a50343a  and  a50336a );
 a50348a <=( (not A199)  and  (not A168) );
 a50349a <=( A169  and  a50348a );
 a50353a <=( (not A202)  and  (not A201) );
 a50354a <=( A200  and  a50353a );
 a50355a <=( a50354a  and  a50349a );
 a50359a <=( A268  and  (not A267) );
 a50360a <=( (not A203)  and  a50359a );
 a50363a <=( (not A299)  and  A298 );
 a50366a <=( A302  and  A300 );
 a50367a <=( a50366a  and  a50363a );
 a50368a <=( a50367a  and  a50360a );
 a50372a <=( (not A199)  and  (not A168) );
 a50373a <=( A169  and  a50372a );
 a50377a <=( (not A202)  and  (not A201) );
 a50378a <=( A200  and  a50377a );
 a50379a <=( a50378a  and  a50373a );
 a50383a <=( A268  and  (not A267) );
 a50384a <=( (not A203)  and  a50383a );
 a50387a <=( A299  and  (not A298) );
 a50390a <=( A301  and  A300 );
 a50391a <=( a50390a  and  a50387a );
 a50392a <=( a50391a  and  a50384a );
 a50396a <=( (not A199)  and  (not A168) );
 a50397a <=( A169  and  a50396a );
 a50401a <=( (not A202)  and  (not A201) );
 a50402a <=( A200  and  a50401a );
 a50403a <=( a50402a  and  a50397a );
 a50407a <=( A268  and  (not A267) );
 a50408a <=( (not A203)  and  a50407a );
 a50411a <=( A299  and  (not A298) );
 a50414a <=( A302  and  A300 );
 a50415a <=( a50414a  and  a50411a );
 a50416a <=( a50415a  and  a50408a );
 a50420a <=( (not A199)  and  (not A168) );
 a50421a <=( A169  and  a50420a );
 a50425a <=( (not A202)  and  (not A201) );
 a50426a <=( A200  and  a50425a );
 a50427a <=( a50426a  and  a50421a );
 a50431a <=( A269  and  (not A267) );
 a50432a <=( (not A203)  and  a50431a );
 a50435a <=( (not A299)  and  A298 );
 a50438a <=( A301  and  A300 );
 a50439a <=( a50438a  and  a50435a );
 a50440a <=( a50439a  and  a50432a );
 a50444a <=( (not A199)  and  (not A168) );
 a50445a <=( A169  and  a50444a );
 a50449a <=( (not A202)  and  (not A201) );
 a50450a <=( A200  and  a50449a );
 a50451a <=( a50450a  and  a50445a );
 a50455a <=( A269  and  (not A267) );
 a50456a <=( (not A203)  and  a50455a );
 a50459a <=( (not A299)  and  A298 );
 a50462a <=( A302  and  A300 );
 a50463a <=( a50462a  and  a50459a );
 a50464a <=( a50463a  and  a50456a );
 a50468a <=( (not A199)  and  (not A168) );
 a50469a <=( A169  and  a50468a );
 a50473a <=( (not A202)  and  (not A201) );
 a50474a <=( A200  and  a50473a );
 a50475a <=( a50474a  and  a50469a );
 a50479a <=( A269  and  (not A267) );
 a50480a <=( (not A203)  and  a50479a );
 a50483a <=( A299  and  (not A298) );
 a50486a <=( A301  and  A300 );
 a50487a <=( a50486a  and  a50483a );
 a50488a <=( a50487a  and  a50480a );
 a50492a <=( (not A199)  and  (not A168) );
 a50493a <=( A169  and  a50492a );
 a50497a <=( (not A202)  and  (not A201) );
 a50498a <=( A200  and  a50497a );
 a50499a <=( a50498a  and  a50493a );
 a50503a <=( A269  and  (not A267) );
 a50504a <=( (not A203)  and  a50503a );
 a50507a <=( A299  and  (not A298) );
 a50510a <=( A302  and  A300 );
 a50511a <=( a50510a  and  a50507a );
 a50512a <=( a50511a  and  a50504a );
 a50516a <=( (not A199)  and  (not A168) );
 a50517a <=( A169  and  a50516a );
 a50521a <=( (not A202)  and  (not A201) );
 a50522a <=( A200  and  a50521a );
 a50523a <=( a50522a  and  a50517a );
 a50527a <=( A266  and  A265 );
 a50528a <=( (not A203)  and  a50527a );
 a50531a <=( (not A299)  and  A298 );
 a50534a <=( A301  and  A300 );
 a50535a <=( a50534a  and  a50531a );
 a50536a <=( a50535a  and  a50528a );
 a50540a <=( (not A199)  and  (not A168) );
 a50541a <=( A169  and  a50540a );
 a50545a <=( (not A202)  and  (not A201) );
 a50546a <=( A200  and  a50545a );
 a50547a <=( a50546a  and  a50541a );
 a50551a <=( A266  and  A265 );
 a50552a <=( (not A203)  and  a50551a );
 a50555a <=( (not A299)  and  A298 );
 a50558a <=( A302  and  A300 );
 a50559a <=( a50558a  and  a50555a );
 a50560a <=( a50559a  and  a50552a );
 a50564a <=( (not A199)  and  (not A168) );
 a50565a <=( A169  and  a50564a );
 a50569a <=( (not A202)  and  (not A201) );
 a50570a <=( A200  and  a50569a );
 a50571a <=( a50570a  and  a50565a );
 a50575a <=( A266  and  A265 );
 a50576a <=( (not A203)  and  a50575a );
 a50579a <=( A299  and  (not A298) );
 a50582a <=( A301  and  A300 );
 a50583a <=( a50582a  and  a50579a );
 a50584a <=( a50583a  and  a50576a );
 a50588a <=( (not A199)  and  (not A168) );
 a50589a <=( A169  and  a50588a );
 a50593a <=( (not A202)  and  (not A201) );
 a50594a <=( A200  and  a50593a );
 a50595a <=( a50594a  and  a50589a );
 a50599a <=( A266  and  A265 );
 a50600a <=( (not A203)  and  a50599a );
 a50603a <=( A299  and  (not A298) );
 a50606a <=( A302  and  A300 );
 a50607a <=( a50606a  and  a50603a );
 a50608a <=( a50607a  and  a50600a );
 a50612a <=( (not A199)  and  (not A168) );
 a50613a <=( A169  and  a50612a );
 a50617a <=( (not A202)  and  (not A201) );
 a50618a <=( A200  and  a50617a );
 a50619a <=( a50618a  and  a50613a );
 a50623a <=( (not A266)  and  (not A265) );
 a50624a <=( (not A203)  and  a50623a );
 a50627a <=( (not A299)  and  A298 );
 a50630a <=( A301  and  A300 );
 a50631a <=( a50630a  and  a50627a );
 a50632a <=( a50631a  and  a50624a );
 a50636a <=( (not A199)  and  (not A168) );
 a50637a <=( A169  and  a50636a );
 a50641a <=( (not A202)  and  (not A201) );
 a50642a <=( A200  and  a50641a );
 a50643a <=( a50642a  and  a50637a );
 a50647a <=( (not A266)  and  (not A265) );
 a50648a <=( (not A203)  and  a50647a );
 a50651a <=( (not A299)  and  A298 );
 a50654a <=( A302  and  A300 );
 a50655a <=( a50654a  and  a50651a );
 a50656a <=( a50655a  and  a50648a );
 a50660a <=( (not A199)  and  (not A168) );
 a50661a <=( A169  and  a50660a );
 a50665a <=( (not A202)  and  (not A201) );
 a50666a <=( A200  and  a50665a );
 a50667a <=( a50666a  and  a50661a );
 a50671a <=( (not A266)  and  (not A265) );
 a50672a <=( (not A203)  and  a50671a );
 a50675a <=( A299  and  (not A298) );
 a50678a <=( A301  and  A300 );
 a50679a <=( a50678a  and  a50675a );
 a50680a <=( a50679a  and  a50672a );
 a50684a <=( (not A199)  and  (not A168) );
 a50685a <=( A169  and  a50684a );
 a50689a <=( (not A202)  and  (not A201) );
 a50690a <=( A200  and  a50689a );
 a50691a <=( a50690a  and  a50685a );
 a50695a <=( (not A266)  and  (not A265) );
 a50696a <=( (not A203)  and  a50695a );
 a50699a <=( A299  and  (not A298) );
 a50702a <=( A302  and  A300 );
 a50703a <=( a50702a  and  a50699a );
 a50704a <=( a50703a  and  a50696a );
 a50708a <=( A199  and  (not A168) );
 a50709a <=( A169  and  a50708a );
 a50713a <=( A202  and  A201 );
 a50714a <=( (not A200)  and  a50713a );
 a50715a <=( a50714a  and  a50709a );
 a50719a <=( (not A269)  and  (not A268) );
 a50720a <=( A267  and  a50719a );
 a50723a <=( (not A299)  and  A298 );
 a50726a <=( A301  and  A300 );
 a50727a <=( a50726a  and  a50723a );
 a50728a <=( a50727a  and  a50720a );
 a50732a <=( A199  and  (not A168) );
 a50733a <=( A169  and  a50732a );
 a50737a <=( A202  and  A201 );
 a50738a <=( (not A200)  and  a50737a );
 a50739a <=( a50738a  and  a50733a );
 a50743a <=( (not A269)  and  (not A268) );
 a50744a <=( A267  and  a50743a );
 a50747a <=( (not A299)  and  A298 );
 a50750a <=( A302  and  A300 );
 a50751a <=( a50750a  and  a50747a );
 a50752a <=( a50751a  and  a50744a );
 a50756a <=( A199  and  (not A168) );
 a50757a <=( A169  and  a50756a );
 a50761a <=( A202  and  A201 );
 a50762a <=( (not A200)  and  a50761a );
 a50763a <=( a50762a  and  a50757a );
 a50767a <=( (not A269)  and  (not A268) );
 a50768a <=( A267  and  a50767a );
 a50771a <=( A299  and  (not A298) );
 a50774a <=( A301  and  A300 );
 a50775a <=( a50774a  and  a50771a );
 a50776a <=( a50775a  and  a50768a );
 a50780a <=( A199  and  (not A168) );
 a50781a <=( A169  and  a50780a );
 a50785a <=( A202  and  A201 );
 a50786a <=( (not A200)  and  a50785a );
 a50787a <=( a50786a  and  a50781a );
 a50791a <=( (not A269)  and  (not A268) );
 a50792a <=( A267  and  a50791a );
 a50795a <=( A299  and  (not A298) );
 a50798a <=( A302  and  A300 );
 a50799a <=( a50798a  and  a50795a );
 a50800a <=( a50799a  and  a50792a );
 a50804a <=( A199  and  (not A168) );
 a50805a <=( A169  and  a50804a );
 a50809a <=( A202  and  A201 );
 a50810a <=( (not A200)  and  a50809a );
 a50811a <=( a50810a  and  a50805a );
 a50815a <=( A298  and  A268 );
 a50816a <=( (not A267)  and  a50815a );
 a50819a <=( (not A300)  and  (not A299) );
 a50822a <=( (not A302)  and  (not A301) );
 a50823a <=( a50822a  and  a50819a );
 a50824a <=( a50823a  and  a50816a );
 a50828a <=( A199  and  (not A168) );
 a50829a <=( A169  and  a50828a );
 a50833a <=( A202  and  A201 );
 a50834a <=( (not A200)  and  a50833a );
 a50835a <=( a50834a  and  a50829a );
 a50839a <=( (not A298)  and  A268 );
 a50840a <=( (not A267)  and  a50839a );
 a50843a <=( (not A300)  and  A299 );
 a50846a <=( (not A302)  and  (not A301) );
 a50847a <=( a50846a  and  a50843a );
 a50848a <=( a50847a  and  a50840a );
 a50852a <=( A199  and  (not A168) );
 a50853a <=( A169  and  a50852a );
 a50857a <=( A202  and  A201 );
 a50858a <=( (not A200)  and  a50857a );
 a50859a <=( a50858a  and  a50853a );
 a50863a <=( A298  and  A269 );
 a50864a <=( (not A267)  and  a50863a );
 a50867a <=( (not A300)  and  (not A299) );
 a50870a <=( (not A302)  and  (not A301) );
 a50871a <=( a50870a  and  a50867a );
 a50872a <=( a50871a  and  a50864a );
 a50876a <=( A199  and  (not A168) );
 a50877a <=( A169  and  a50876a );
 a50881a <=( A202  and  A201 );
 a50882a <=( (not A200)  and  a50881a );
 a50883a <=( a50882a  and  a50877a );
 a50887a <=( (not A298)  and  A269 );
 a50888a <=( (not A267)  and  a50887a );
 a50891a <=( (not A300)  and  A299 );
 a50894a <=( (not A302)  and  (not A301) );
 a50895a <=( a50894a  and  a50891a );
 a50896a <=( a50895a  and  a50888a );
 a50900a <=( A199  and  (not A168) );
 a50901a <=( A169  and  a50900a );
 a50905a <=( A202  and  A201 );
 a50906a <=( (not A200)  and  a50905a );
 a50907a <=( a50906a  and  a50901a );
 a50911a <=( A298  and  A266 );
 a50912a <=( A265  and  a50911a );
 a50915a <=( (not A300)  and  (not A299) );
 a50918a <=( (not A302)  and  (not A301) );
 a50919a <=( a50918a  and  a50915a );
 a50920a <=( a50919a  and  a50912a );
 a50924a <=( A199  and  (not A168) );
 a50925a <=( A169  and  a50924a );
 a50929a <=( A202  and  A201 );
 a50930a <=( (not A200)  and  a50929a );
 a50931a <=( a50930a  and  a50925a );
 a50935a <=( (not A298)  and  A266 );
 a50936a <=( A265  and  a50935a );
 a50939a <=( (not A300)  and  A299 );
 a50942a <=( (not A302)  and  (not A301) );
 a50943a <=( a50942a  and  a50939a );
 a50944a <=( a50943a  and  a50936a );
 a50948a <=( A199  and  (not A168) );
 a50949a <=( A169  and  a50948a );
 a50953a <=( A202  and  A201 );
 a50954a <=( (not A200)  and  a50953a );
 a50955a <=( a50954a  and  a50949a );
 a50959a <=( A298  and  (not A266) );
 a50960a <=( (not A265)  and  a50959a );
 a50963a <=( (not A300)  and  (not A299) );
 a50966a <=( (not A302)  and  (not A301) );
 a50967a <=( a50966a  and  a50963a );
 a50968a <=( a50967a  and  a50960a );
 a50972a <=( A199  and  (not A168) );
 a50973a <=( A169  and  a50972a );
 a50977a <=( A202  and  A201 );
 a50978a <=( (not A200)  and  a50977a );
 a50979a <=( a50978a  and  a50973a );
 a50983a <=( (not A298)  and  (not A266) );
 a50984a <=( (not A265)  and  a50983a );
 a50987a <=( (not A300)  and  A299 );
 a50990a <=( (not A302)  and  (not A301) );
 a50991a <=( a50990a  and  a50987a );
 a50992a <=( a50991a  and  a50984a );
 a50996a <=( A199  and  (not A168) );
 a50997a <=( A169  and  a50996a );
 a51001a <=( A203  and  A201 );
 a51002a <=( (not A200)  and  a51001a );
 a51003a <=( a51002a  and  a50997a );
 a51007a <=( (not A269)  and  (not A268) );
 a51008a <=( A267  and  a51007a );
 a51011a <=( (not A299)  and  A298 );
 a51014a <=( A301  and  A300 );
 a51015a <=( a51014a  and  a51011a );
 a51016a <=( a51015a  and  a51008a );
 a51020a <=( A199  and  (not A168) );
 a51021a <=( A169  and  a51020a );
 a51025a <=( A203  and  A201 );
 a51026a <=( (not A200)  and  a51025a );
 a51027a <=( a51026a  and  a51021a );
 a51031a <=( (not A269)  and  (not A268) );
 a51032a <=( A267  and  a51031a );
 a51035a <=( (not A299)  and  A298 );
 a51038a <=( A302  and  A300 );
 a51039a <=( a51038a  and  a51035a );
 a51040a <=( a51039a  and  a51032a );
 a51044a <=( A199  and  (not A168) );
 a51045a <=( A169  and  a51044a );
 a51049a <=( A203  and  A201 );
 a51050a <=( (not A200)  and  a51049a );
 a51051a <=( a51050a  and  a51045a );
 a51055a <=( (not A269)  and  (not A268) );
 a51056a <=( A267  and  a51055a );
 a51059a <=( A299  and  (not A298) );
 a51062a <=( A301  and  A300 );
 a51063a <=( a51062a  and  a51059a );
 a51064a <=( a51063a  and  a51056a );
 a51068a <=( A199  and  (not A168) );
 a51069a <=( A169  and  a51068a );
 a51073a <=( A203  and  A201 );
 a51074a <=( (not A200)  and  a51073a );
 a51075a <=( a51074a  and  a51069a );
 a51079a <=( (not A269)  and  (not A268) );
 a51080a <=( A267  and  a51079a );
 a51083a <=( A299  and  (not A298) );
 a51086a <=( A302  and  A300 );
 a51087a <=( a51086a  and  a51083a );
 a51088a <=( a51087a  and  a51080a );
 a51092a <=( A199  and  (not A168) );
 a51093a <=( A169  and  a51092a );
 a51097a <=( A203  and  A201 );
 a51098a <=( (not A200)  and  a51097a );
 a51099a <=( a51098a  and  a51093a );
 a51103a <=( A298  and  A268 );
 a51104a <=( (not A267)  and  a51103a );
 a51107a <=( (not A300)  and  (not A299) );
 a51110a <=( (not A302)  and  (not A301) );
 a51111a <=( a51110a  and  a51107a );
 a51112a <=( a51111a  and  a51104a );
 a51116a <=( A199  and  (not A168) );
 a51117a <=( A169  and  a51116a );
 a51121a <=( A203  and  A201 );
 a51122a <=( (not A200)  and  a51121a );
 a51123a <=( a51122a  and  a51117a );
 a51127a <=( (not A298)  and  A268 );
 a51128a <=( (not A267)  and  a51127a );
 a51131a <=( (not A300)  and  A299 );
 a51134a <=( (not A302)  and  (not A301) );
 a51135a <=( a51134a  and  a51131a );
 a51136a <=( a51135a  and  a51128a );
 a51140a <=( A199  and  (not A168) );
 a51141a <=( A169  and  a51140a );
 a51145a <=( A203  and  A201 );
 a51146a <=( (not A200)  and  a51145a );
 a51147a <=( a51146a  and  a51141a );
 a51151a <=( A298  and  A269 );
 a51152a <=( (not A267)  and  a51151a );
 a51155a <=( (not A300)  and  (not A299) );
 a51158a <=( (not A302)  and  (not A301) );
 a51159a <=( a51158a  and  a51155a );
 a51160a <=( a51159a  and  a51152a );
 a51164a <=( A199  and  (not A168) );
 a51165a <=( A169  and  a51164a );
 a51169a <=( A203  and  A201 );
 a51170a <=( (not A200)  and  a51169a );
 a51171a <=( a51170a  and  a51165a );
 a51175a <=( (not A298)  and  A269 );
 a51176a <=( (not A267)  and  a51175a );
 a51179a <=( (not A300)  and  A299 );
 a51182a <=( (not A302)  and  (not A301) );
 a51183a <=( a51182a  and  a51179a );
 a51184a <=( a51183a  and  a51176a );
 a51188a <=( A199  and  (not A168) );
 a51189a <=( A169  and  a51188a );
 a51193a <=( A203  and  A201 );
 a51194a <=( (not A200)  and  a51193a );
 a51195a <=( a51194a  and  a51189a );
 a51199a <=( A298  and  A266 );
 a51200a <=( A265  and  a51199a );
 a51203a <=( (not A300)  and  (not A299) );
 a51206a <=( (not A302)  and  (not A301) );
 a51207a <=( a51206a  and  a51203a );
 a51208a <=( a51207a  and  a51200a );
 a51212a <=( A199  and  (not A168) );
 a51213a <=( A169  and  a51212a );
 a51217a <=( A203  and  A201 );
 a51218a <=( (not A200)  and  a51217a );
 a51219a <=( a51218a  and  a51213a );
 a51223a <=( (not A298)  and  A266 );
 a51224a <=( A265  and  a51223a );
 a51227a <=( (not A300)  and  A299 );
 a51230a <=( (not A302)  and  (not A301) );
 a51231a <=( a51230a  and  a51227a );
 a51232a <=( a51231a  and  a51224a );
 a51236a <=( A199  and  (not A168) );
 a51237a <=( A169  and  a51236a );
 a51241a <=( A203  and  A201 );
 a51242a <=( (not A200)  and  a51241a );
 a51243a <=( a51242a  and  a51237a );
 a51247a <=( A298  and  (not A266) );
 a51248a <=( (not A265)  and  a51247a );
 a51251a <=( (not A300)  and  (not A299) );
 a51254a <=( (not A302)  and  (not A301) );
 a51255a <=( a51254a  and  a51251a );
 a51256a <=( a51255a  and  a51248a );
 a51260a <=( A199  and  (not A168) );
 a51261a <=( A169  and  a51260a );
 a51265a <=( A203  and  A201 );
 a51266a <=( (not A200)  and  a51265a );
 a51267a <=( a51266a  and  a51261a );
 a51271a <=( (not A298)  and  (not A266) );
 a51272a <=( (not A265)  and  a51271a );
 a51275a <=( (not A300)  and  A299 );
 a51278a <=( (not A302)  and  (not A301) );
 a51279a <=( a51278a  and  a51275a );
 a51280a <=( a51279a  and  a51272a );
 a51284a <=( A199  and  (not A168) );
 a51285a <=( A169  and  a51284a );
 a51289a <=( (not A202)  and  (not A201) );
 a51290a <=( (not A200)  and  a51289a );
 a51291a <=( a51290a  and  a51285a );
 a51295a <=( A268  and  (not A267) );
 a51296a <=( (not A203)  and  a51295a );
 a51299a <=( (not A299)  and  A298 );
 a51302a <=( A301  and  A300 );
 a51303a <=( a51302a  and  a51299a );
 a51304a <=( a51303a  and  a51296a );
 a51308a <=( A199  and  (not A168) );
 a51309a <=( A169  and  a51308a );
 a51313a <=( (not A202)  and  (not A201) );
 a51314a <=( (not A200)  and  a51313a );
 a51315a <=( a51314a  and  a51309a );
 a51319a <=( A268  and  (not A267) );
 a51320a <=( (not A203)  and  a51319a );
 a51323a <=( (not A299)  and  A298 );
 a51326a <=( A302  and  A300 );
 a51327a <=( a51326a  and  a51323a );
 a51328a <=( a51327a  and  a51320a );
 a51332a <=( A199  and  (not A168) );
 a51333a <=( A169  and  a51332a );
 a51337a <=( (not A202)  and  (not A201) );
 a51338a <=( (not A200)  and  a51337a );
 a51339a <=( a51338a  and  a51333a );
 a51343a <=( A268  and  (not A267) );
 a51344a <=( (not A203)  and  a51343a );
 a51347a <=( A299  and  (not A298) );
 a51350a <=( A301  and  A300 );
 a51351a <=( a51350a  and  a51347a );
 a51352a <=( a51351a  and  a51344a );
 a51356a <=( A199  and  (not A168) );
 a51357a <=( A169  and  a51356a );
 a51361a <=( (not A202)  and  (not A201) );
 a51362a <=( (not A200)  and  a51361a );
 a51363a <=( a51362a  and  a51357a );
 a51367a <=( A268  and  (not A267) );
 a51368a <=( (not A203)  and  a51367a );
 a51371a <=( A299  and  (not A298) );
 a51374a <=( A302  and  A300 );
 a51375a <=( a51374a  and  a51371a );
 a51376a <=( a51375a  and  a51368a );
 a51380a <=( A199  and  (not A168) );
 a51381a <=( A169  and  a51380a );
 a51385a <=( (not A202)  and  (not A201) );
 a51386a <=( (not A200)  and  a51385a );
 a51387a <=( a51386a  and  a51381a );
 a51391a <=( A269  and  (not A267) );
 a51392a <=( (not A203)  and  a51391a );
 a51395a <=( (not A299)  and  A298 );
 a51398a <=( A301  and  A300 );
 a51399a <=( a51398a  and  a51395a );
 a51400a <=( a51399a  and  a51392a );
 a51404a <=( A199  and  (not A168) );
 a51405a <=( A169  and  a51404a );
 a51409a <=( (not A202)  and  (not A201) );
 a51410a <=( (not A200)  and  a51409a );
 a51411a <=( a51410a  and  a51405a );
 a51415a <=( A269  and  (not A267) );
 a51416a <=( (not A203)  and  a51415a );
 a51419a <=( (not A299)  and  A298 );
 a51422a <=( A302  and  A300 );
 a51423a <=( a51422a  and  a51419a );
 a51424a <=( a51423a  and  a51416a );
 a51428a <=( A199  and  (not A168) );
 a51429a <=( A169  and  a51428a );
 a51433a <=( (not A202)  and  (not A201) );
 a51434a <=( (not A200)  and  a51433a );
 a51435a <=( a51434a  and  a51429a );
 a51439a <=( A269  and  (not A267) );
 a51440a <=( (not A203)  and  a51439a );
 a51443a <=( A299  and  (not A298) );
 a51446a <=( A301  and  A300 );
 a51447a <=( a51446a  and  a51443a );
 a51448a <=( a51447a  and  a51440a );
 a51452a <=( A199  and  (not A168) );
 a51453a <=( A169  and  a51452a );
 a51457a <=( (not A202)  and  (not A201) );
 a51458a <=( (not A200)  and  a51457a );
 a51459a <=( a51458a  and  a51453a );
 a51463a <=( A269  and  (not A267) );
 a51464a <=( (not A203)  and  a51463a );
 a51467a <=( A299  and  (not A298) );
 a51470a <=( A302  and  A300 );
 a51471a <=( a51470a  and  a51467a );
 a51472a <=( a51471a  and  a51464a );
 a51476a <=( A199  and  (not A168) );
 a51477a <=( A169  and  a51476a );
 a51481a <=( (not A202)  and  (not A201) );
 a51482a <=( (not A200)  and  a51481a );
 a51483a <=( a51482a  and  a51477a );
 a51487a <=( A266  and  A265 );
 a51488a <=( (not A203)  and  a51487a );
 a51491a <=( (not A299)  and  A298 );
 a51494a <=( A301  and  A300 );
 a51495a <=( a51494a  and  a51491a );
 a51496a <=( a51495a  and  a51488a );
 a51500a <=( A199  and  (not A168) );
 a51501a <=( A169  and  a51500a );
 a51505a <=( (not A202)  and  (not A201) );
 a51506a <=( (not A200)  and  a51505a );
 a51507a <=( a51506a  and  a51501a );
 a51511a <=( A266  and  A265 );
 a51512a <=( (not A203)  and  a51511a );
 a51515a <=( (not A299)  and  A298 );
 a51518a <=( A302  and  A300 );
 a51519a <=( a51518a  and  a51515a );
 a51520a <=( a51519a  and  a51512a );
 a51524a <=( A199  and  (not A168) );
 a51525a <=( A169  and  a51524a );
 a51529a <=( (not A202)  and  (not A201) );
 a51530a <=( (not A200)  and  a51529a );
 a51531a <=( a51530a  and  a51525a );
 a51535a <=( A266  and  A265 );
 a51536a <=( (not A203)  and  a51535a );
 a51539a <=( A299  and  (not A298) );
 a51542a <=( A301  and  A300 );
 a51543a <=( a51542a  and  a51539a );
 a51544a <=( a51543a  and  a51536a );
 a51548a <=( A199  and  (not A168) );
 a51549a <=( A169  and  a51548a );
 a51553a <=( (not A202)  and  (not A201) );
 a51554a <=( (not A200)  and  a51553a );
 a51555a <=( a51554a  and  a51549a );
 a51559a <=( A266  and  A265 );
 a51560a <=( (not A203)  and  a51559a );
 a51563a <=( A299  and  (not A298) );
 a51566a <=( A302  and  A300 );
 a51567a <=( a51566a  and  a51563a );
 a51568a <=( a51567a  and  a51560a );
 a51572a <=( A199  and  (not A168) );
 a51573a <=( A169  and  a51572a );
 a51577a <=( (not A202)  and  (not A201) );
 a51578a <=( (not A200)  and  a51577a );
 a51579a <=( a51578a  and  a51573a );
 a51583a <=( (not A266)  and  (not A265) );
 a51584a <=( (not A203)  and  a51583a );
 a51587a <=( (not A299)  and  A298 );
 a51590a <=( A301  and  A300 );
 a51591a <=( a51590a  and  a51587a );
 a51592a <=( a51591a  and  a51584a );
 a51596a <=( A199  and  (not A168) );
 a51597a <=( A169  and  a51596a );
 a51601a <=( (not A202)  and  (not A201) );
 a51602a <=( (not A200)  and  a51601a );
 a51603a <=( a51602a  and  a51597a );
 a51607a <=( (not A266)  and  (not A265) );
 a51608a <=( (not A203)  and  a51607a );
 a51611a <=( (not A299)  and  A298 );
 a51614a <=( A302  and  A300 );
 a51615a <=( a51614a  and  a51611a );
 a51616a <=( a51615a  and  a51608a );
 a51620a <=( A199  and  (not A168) );
 a51621a <=( A169  and  a51620a );
 a51625a <=( (not A202)  and  (not A201) );
 a51626a <=( (not A200)  and  a51625a );
 a51627a <=( a51626a  and  a51621a );
 a51631a <=( (not A266)  and  (not A265) );
 a51632a <=( (not A203)  and  a51631a );
 a51635a <=( A299  and  (not A298) );
 a51638a <=( A301  and  A300 );
 a51639a <=( a51638a  and  a51635a );
 a51640a <=( a51639a  and  a51632a );
 a51644a <=( A199  and  (not A168) );
 a51645a <=( A169  and  a51644a );
 a51649a <=( (not A202)  and  (not A201) );
 a51650a <=( (not A200)  and  a51649a );
 a51651a <=( a51650a  and  a51645a );
 a51655a <=( (not A266)  and  (not A265) );
 a51656a <=( (not A203)  and  a51655a );
 a51659a <=( A299  and  (not A298) );
 a51662a <=( A302  and  A300 );
 a51663a <=( a51662a  and  a51659a );
 a51664a <=( a51663a  and  a51656a );
 a51668a <=( A168  and  (not A169) );
 a51669a <=( A170  and  a51668a );
 a51673a <=( (not A203)  and  (not A202) );
 a51674a <=( A201  and  a51673a );
 a51675a <=( a51674a  and  a51669a );
 a51679a <=( A267  and  A266 );
 a51680a <=( (not A265)  and  a51679a );
 a51683a <=( A300  and  A268 );
 a51686a <=( (not A302)  and  (not A301) );
 a51687a <=( a51686a  and  a51683a );
 a51688a <=( a51687a  and  a51680a );
 a51692a <=( A168  and  (not A169) );
 a51693a <=( A170  and  a51692a );
 a51697a <=( (not A203)  and  (not A202) );
 a51698a <=( A201  and  a51697a );
 a51699a <=( a51698a  and  a51693a );
 a51703a <=( A267  and  A266 );
 a51704a <=( (not A265)  and  a51703a );
 a51707a <=( A300  and  A269 );
 a51710a <=( (not A302)  and  (not A301) );
 a51711a <=( a51710a  and  a51707a );
 a51712a <=( a51711a  and  a51704a );
 a51716a <=( A168  and  (not A169) );
 a51717a <=( A170  and  a51716a );
 a51721a <=( (not A203)  and  (not A202) );
 a51722a <=( A201  and  a51721a );
 a51723a <=( a51722a  and  a51717a );
 a51727a <=( (not A267)  and  A266 );
 a51728a <=( (not A265)  and  a51727a );
 a51731a <=( (not A269)  and  (not A268) );
 a51734a <=( A301  and  (not A300) );
 a51735a <=( a51734a  and  a51731a );
 a51736a <=( a51735a  and  a51728a );
 a51740a <=( A168  and  (not A169) );
 a51741a <=( A170  and  a51740a );
 a51745a <=( (not A203)  and  (not A202) );
 a51746a <=( A201  and  a51745a );
 a51747a <=( a51746a  and  a51741a );
 a51751a <=( (not A267)  and  A266 );
 a51752a <=( (not A265)  and  a51751a );
 a51755a <=( (not A269)  and  (not A268) );
 a51758a <=( A302  and  (not A300) );
 a51759a <=( a51758a  and  a51755a );
 a51760a <=( a51759a  and  a51752a );
 a51764a <=( A168  and  (not A169) );
 a51765a <=( A170  and  a51764a );
 a51769a <=( (not A203)  and  (not A202) );
 a51770a <=( A201  and  a51769a );
 a51771a <=( a51770a  and  a51765a );
 a51775a <=( (not A267)  and  A266 );
 a51776a <=( (not A265)  and  a51775a );
 a51779a <=( (not A269)  and  (not A268) );
 a51782a <=( A299  and  A298 );
 a51783a <=( a51782a  and  a51779a );
 a51784a <=( a51783a  and  a51776a );
 a51788a <=( A168  and  (not A169) );
 a51789a <=( A170  and  a51788a );
 a51793a <=( (not A203)  and  (not A202) );
 a51794a <=( A201  and  a51793a );
 a51795a <=( a51794a  and  a51789a );
 a51799a <=( (not A267)  and  A266 );
 a51800a <=( (not A265)  and  a51799a );
 a51803a <=( (not A269)  and  (not A268) );
 a51806a <=( (not A299)  and  (not A298) );
 a51807a <=( a51806a  and  a51803a );
 a51808a <=( a51807a  and  a51800a );
 a51812a <=( A168  and  (not A169) );
 a51813a <=( A170  and  a51812a );
 a51817a <=( (not A203)  and  (not A202) );
 a51818a <=( A201  and  a51817a );
 a51819a <=( a51818a  and  a51813a );
 a51823a <=( A267  and  (not A266) );
 a51824a <=( A265  and  a51823a );
 a51827a <=( A300  and  A268 );
 a51830a <=( (not A302)  and  (not A301) );
 a51831a <=( a51830a  and  a51827a );
 a51832a <=( a51831a  and  a51824a );
 a51836a <=( A168  and  (not A169) );
 a51837a <=( A170  and  a51836a );
 a51841a <=( (not A203)  and  (not A202) );
 a51842a <=( A201  and  a51841a );
 a51843a <=( a51842a  and  a51837a );
 a51847a <=( A267  and  (not A266) );
 a51848a <=( A265  and  a51847a );
 a51851a <=( A300  and  A269 );
 a51854a <=( (not A302)  and  (not A301) );
 a51855a <=( a51854a  and  a51851a );
 a51856a <=( a51855a  and  a51848a );
 a51860a <=( A168  and  (not A169) );
 a51861a <=( A170  and  a51860a );
 a51865a <=( (not A203)  and  (not A202) );
 a51866a <=( A201  and  a51865a );
 a51867a <=( a51866a  and  a51861a );
 a51871a <=( (not A267)  and  (not A266) );
 a51872a <=( A265  and  a51871a );
 a51875a <=( (not A269)  and  (not A268) );
 a51878a <=( A301  and  (not A300) );
 a51879a <=( a51878a  and  a51875a );
 a51880a <=( a51879a  and  a51872a );
 a51884a <=( A168  and  (not A169) );
 a51885a <=( A170  and  a51884a );
 a51889a <=( (not A203)  and  (not A202) );
 a51890a <=( A201  and  a51889a );
 a51891a <=( a51890a  and  a51885a );
 a51895a <=( (not A267)  and  (not A266) );
 a51896a <=( A265  and  a51895a );
 a51899a <=( (not A269)  and  (not A268) );
 a51902a <=( A302  and  (not A300) );
 a51903a <=( a51902a  and  a51899a );
 a51904a <=( a51903a  and  a51896a );
 a51908a <=( A168  and  (not A169) );
 a51909a <=( A170  and  a51908a );
 a51913a <=( (not A203)  and  (not A202) );
 a51914a <=( A201  and  a51913a );
 a51915a <=( a51914a  and  a51909a );
 a51919a <=( (not A267)  and  (not A266) );
 a51920a <=( A265  and  a51919a );
 a51923a <=( (not A269)  and  (not A268) );
 a51926a <=( A299  and  A298 );
 a51927a <=( a51926a  and  a51923a );
 a51928a <=( a51927a  and  a51920a );
 a51932a <=( A168  and  (not A169) );
 a51933a <=( A170  and  a51932a );
 a51937a <=( (not A203)  and  (not A202) );
 a51938a <=( A201  and  a51937a );
 a51939a <=( a51938a  and  a51933a );
 a51943a <=( (not A267)  and  (not A266) );
 a51944a <=( A265  and  a51943a );
 a51947a <=( (not A269)  and  (not A268) );
 a51950a <=( (not A299)  and  (not A298) );
 a51951a <=( a51950a  and  a51947a );
 a51952a <=( a51951a  and  a51944a );
 a51956a <=( A168  and  (not A169) );
 a51957a <=( A170  and  a51956a );
 a51961a <=( (not A265)  and  A202 );
 a51962a <=( (not A201)  and  a51961a );
 a51963a <=( a51962a  and  a51957a );
 a51967a <=( (not A268)  and  (not A267) );
 a51968a <=( A266  and  a51967a );
 a51971a <=( A300  and  (not A269) );
 a51974a <=( (not A302)  and  (not A301) );
 a51975a <=( a51974a  and  a51971a );
 a51976a <=( a51975a  and  a51968a );
 a51980a <=( A168  and  (not A169) );
 a51981a <=( A170  and  a51980a );
 a51985a <=( A265  and  A202 );
 a51986a <=( (not A201)  and  a51985a );
 a51987a <=( a51986a  and  a51981a );
 a51991a <=( (not A268)  and  (not A267) );
 a51992a <=( (not A266)  and  a51991a );
 a51995a <=( A300  and  (not A269) );
 a51998a <=( (not A302)  and  (not A301) );
 a51999a <=( a51998a  and  a51995a );
 a52000a <=( a51999a  and  a51992a );
 a52004a <=( A168  and  (not A169) );
 a52005a <=( A170  and  a52004a );
 a52009a <=( (not A265)  and  A203 );
 a52010a <=( (not A201)  and  a52009a );
 a52011a <=( a52010a  and  a52005a );
 a52015a <=( (not A268)  and  (not A267) );
 a52016a <=( A266  and  a52015a );
 a52019a <=( A300  and  (not A269) );
 a52022a <=( (not A302)  and  (not A301) );
 a52023a <=( a52022a  and  a52019a );
 a52024a <=( a52023a  and  a52016a );
 a52028a <=( A168  and  (not A169) );
 a52029a <=( A170  and  a52028a );
 a52033a <=( A265  and  A203 );
 a52034a <=( (not A201)  and  a52033a );
 a52035a <=( a52034a  and  a52029a );
 a52039a <=( (not A268)  and  (not A267) );
 a52040a <=( (not A266)  and  a52039a );
 a52043a <=( A300  and  (not A269) );
 a52046a <=( (not A302)  and  (not A301) );
 a52047a <=( a52046a  and  a52043a );
 a52048a <=( a52047a  and  a52040a );
 a52052a <=( A168  and  (not A169) );
 a52053a <=( A170  and  a52052a );
 a52057a <=( (not A265)  and  A200 );
 a52058a <=( A199  and  a52057a );
 a52059a <=( a52058a  and  a52053a );
 a52063a <=( (not A268)  and  (not A267) );
 a52064a <=( A266  and  a52063a );
 a52067a <=( A300  and  (not A269) );
 a52070a <=( (not A302)  and  (not A301) );
 a52071a <=( a52070a  and  a52067a );
 a52072a <=( a52071a  and  a52064a );
 a52076a <=( A168  and  (not A169) );
 a52077a <=( A170  and  a52076a );
 a52081a <=( A265  and  A200 );
 a52082a <=( A199  and  a52081a );
 a52083a <=( a52082a  and  a52077a );
 a52087a <=( (not A268)  and  (not A267) );
 a52088a <=( (not A266)  and  a52087a );
 a52091a <=( A300  and  (not A269) );
 a52094a <=( (not A302)  and  (not A301) );
 a52095a <=( a52094a  and  a52091a );
 a52096a <=( a52095a  and  a52088a );
 a52100a <=( A168  and  (not A169) );
 a52101a <=( A170  and  a52100a );
 a52105a <=( A201  and  A200 );
 a52106a <=( (not A199)  and  a52105a );
 a52107a <=( a52106a  and  a52101a );
 a52111a <=( A268  and  (not A267) );
 a52112a <=( A202  and  a52111a );
 a52115a <=( (not A299)  and  A298 );
 a52118a <=( A301  and  A300 );
 a52119a <=( a52118a  and  a52115a );
 a52120a <=( a52119a  and  a52112a );
 a52124a <=( A168  and  (not A169) );
 a52125a <=( A170  and  a52124a );
 a52129a <=( A201  and  A200 );
 a52130a <=( (not A199)  and  a52129a );
 a52131a <=( a52130a  and  a52125a );
 a52135a <=( A268  and  (not A267) );
 a52136a <=( A202  and  a52135a );
 a52139a <=( (not A299)  and  A298 );
 a52142a <=( A302  and  A300 );
 a52143a <=( a52142a  and  a52139a );
 a52144a <=( a52143a  and  a52136a );
 a52148a <=( A168  and  (not A169) );
 a52149a <=( A170  and  a52148a );
 a52153a <=( A201  and  A200 );
 a52154a <=( (not A199)  and  a52153a );
 a52155a <=( a52154a  and  a52149a );
 a52159a <=( A268  and  (not A267) );
 a52160a <=( A202  and  a52159a );
 a52163a <=( A299  and  (not A298) );
 a52166a <=( A301  and  A300 );
 a52167a <=( a52166a  and  a52163a );
 a52168a <=( a52167a  and  a52160a );
 a52172a <=( A168  and  (not A169) );
 a52173a <=( A170  and  a52172a );
 a52177a <=( A201  and  A200 );
 a52178a <=( (not A199)  and  a52177a );
 a52179a <=( a52178a  and  a52173a );
 a52183a <=( A268  and  (not A267) );
 a52184a <=( A202  and  a52183a );
 a52187a <=( A299  and  (not A298) );
 a52190a <=( A302  and  A300 );
 a52191a <=( a52190a  and  a52187a );
 a52192a <=( a52191a  and  a52184a );
 a52196a <=( A168  and  (not A169) );
 a52197a <=( A170  and  a52196a );
 a52201a <=( A201  and  A200 );
 a52202a <=( (not A199)  and  a52201a );
 a52203a <=( a52202a  and  a52197a );
 a52207a <=( A269  and  (not A267) );
 a52208a <=( A202  and  a52207a );
 a52211a <=( (not A299)  and  A298 );
 a52214a <=( A301  and  A300 );
 a52215a <=( a52214a  and  a52211a );
 a52216a <=( a52215a  and  a52208a );
 a52220a <=( A168  and  (not A169) );
 a52221a <=( A170  and  a52220a );
 a52225a <=( A201  and  A200 );
 a52226a <=( (not A199)  and  a52225a );
 a52227a <=( a52226a  and  a52221a );
 a52231a <=( A269  and  (not A267) );
 a52232a <=( A202  and  a52231a );
 a52235a <=( (not A299)  and  A298 );
 a52238a <=( A302  and  A300 );
 a52239a <=( a52238a  and  a52235a );
 a52240a <=( a52239a  and  a52232a );
 a52244a <=( A168  and  (not A169) );
 a52245a <=( A170  and  a52244a );
 a52249a <=( A201  and  A200 );
 a52250a <=( (not A199)  and  a52249a );
 a52251a <=( a52250a  and  a52245a );
 a52255a <=( A269  and  (not A267) );
 a52256a <=( A202  and  a52255a );
 a52259a <=( A299  and  (not A298) );
 a52262a <=( A301  and  A300 );
 a52263a <=( a52262a  and  a52259a );
 a52264a <=( a52263a  and  a52256a );
 a52268a <=( A168  and  (not A169) );
 a52269a <=( A170  and  a52268a );
 a52273a <=( A201  and  A200 );
 a52274a <=( (not A199)  and  a52273a );
 a52275a <=( a52274a  and  a52269a );
 a52279a <=( A269  and  (not A267) );
 a52280a <=( A202  and  a52279a );
 a52283a <=( A299  and  (not A298) );
 a52286a <=( A302  and  A300 );
 a52287a <=( a52286a  and  a52283a );
 a52288a <=( a52287a  and  a52280a );
 a52292a <=( A168  and  (not A169) );
 a52293a <=( A170  and  a52292a );
 a52297a <=( A201  and  A200 );
 a52298a <=( (not A199)  and  a52297a );
 a52299a <=( a52298a  and  a52293a );
 a52303a <=( A266  and  A265 );
 a52304a <=( A202  and  a52303a );
 a52307a <=( (not A299)  and  A298 );
 a52310a <=( A301  and  A300 );
 a52311a <=( a52310a  and  a52307a );
 a52312a <=( a52311a  and  a52304a );
 a52316a <=( A168  and  (not A169) );
 a52317a <=( A170  and  a52316a );
 a52321a <=( A201  and  A200 );
 a52322a <=( (not A199)  and  a52321a );
 a52323a <=( a52322a  and  a52317a );
 a52327a <=( A266  and  A265 );
 a52328a <=( A202  and  a52327a );
 a52331a <=( (not A299)  and  A298 );
 a52334a <=( A302  and  A300 );
 a52335a <=( a52334a  and  a52331a );
 a52336a <=( a52335a  and  a52328a );
 a52340a <=( A168  and  (not A169) );
 a52341a <=( A170  and  a52340a );
 a52345a <=( A201  and  A200 );
 a52346a <=( (not A199)  and  a52345a );
 a52347a <=( a52346a  and  a52341a );
 a52351a <=( A266  and  A265 );
 a52352a <=( A202  and  a52351a );
 a52355a <=( A299  and  (not A298) );
 a52358a <=( A301  and  A300 );
 a52359a <=( a52358a  and  a52355a );
 a52360a <=( a52359a  and  a52352a );
 a52364a <=( A168  and  (not A169) );
 a52365a <=( A170  and  a52364a );
 a52369a <=( A201  and  A200 );
 a52370a <=( (not A199)  and  a52369a );
 a52371a <=( a52370a  and  a52365a );
 a52375a <=( A266  and  A265 );
 a52376a <=( A202  and  a52375a );
 a52379a <=( A299  and  (not A298) );
 a52382a <=( A302  and  A300 );
 a52383a <=( a52382a  and  a52379a );
 a52384a <=( a52383a  and  a52376a );
 a52388a <=( A168  and  (not A169) );
 a52389a <=( A170  and  a52388a );
 a52393a <=( A201  and  A200 );
 a52394a <=( (not A199)  and  a52393a );
 a52395a <=( a52394a  and  a52389a );
 a52399a <=( (not A266)  and  (not A265) );
 a52400a <=( A202  and  a52399a );
 a52403a <=( (not A299)  and  A298 );
 a52406a <=( A301  and  A300 );
 a52407a <=( a52406a  and  a52403a );
 a52408a <=( a52407a  and  a52400a );
 a52412a <=( A168  and  (not A169) );
 a52413a <=( A170  and  a52412a );
 a52417a <=( A201  and  A200 );
 a52418a <=( (not A199)  and  a52417a );
 a52419a <=( a52418a  and  a52413a );
 a52423a <=( (not A266)  and  (not A265) );
 a52424a <=( A202  and  a52423a );
 a52427a <=( (not A299)  and  A298 );
 a52430a <=( A302  and  A300 );
 a52431a <=( a52430a  and  a52427a );
 a52432a <=( a52431a  and  a52424a );
 a52436a <=( A168  and  (not A169) );
 a52437a <=( A170  and  a52436a );
 a52441a <=( A201  and  A200 );
 a52442a <=( (not A199)  and  a52441a );
 a52443a <=( a52442a  and  a52437a );
 a52447a <=( (not A266)  and  (not A265) );
 a52448a <=( A202  and  a52447a );
 a52451a <=( A299  and  (not A298) );
 a52454a <=( A301  and  A300 );
 a52455a <=( a52454a  and  a52451a );
 a52456a <=( a52455a  and  a52448a );
 a52460a <=( A168  and  (not A169) );
 a52461a <=( A170  and  a52460a );
 a52465a <=( A201  and  A200 );
 a52466a <=( (not A199)  and  a52465a );
 a52467a <=( a52466a  and  a52461a );
 a52471a <=( (not A266)  and  (not A265) );
 a52472a <=( A202  and  a52471a );
 a52475a <=( A299  and  (not A298) );
 a52478a <=( A302  and  A300 );
 a52479a <=( a52478a  and  a52475a );
 a52480a <=( a52479a  and  a52472a );
 a52484a <=( A168  and  (not A169) );
 a52485a <=( A170  and  a52484a );
 a52489a <=( A201  and  A200 );
 a52490a <=( (not A199)  and  a52489a );
 a52491a <=( a52490a  and  a52485a );
 a52495a <=( A268  and  (not A267) );
 a52496a <=( A203  and  a52495a );
 a52499a <=( (not A299)  and  A298 );
 a52502a <=( A301  and  A300 );
 a52503a <=( a52502a  and  a52499a );
 a52504a <=( a52503a  and  a52496a );
 a52508a <=( A168  and  (not A169) );
 a52509a <=( A170  and  a52508a );
 a52513a <=( A201  and  A200 );
 a52514a <=( (not A199)  and  a52513a );
 a52515a <=( a52514a  and  a52509a );
 a52519a <=( A268  and  (not A267) );
 a52520a <=( A203  and  a52519a );
 a52523a <=( (not A299)  and  A298 );
 a52526a <=( A302  and  A300 );
 a52527a <=( a52526a  and  a52523a );
 a52528a <=( a52527a  and  a52520a );
 a52532a <=( A168  and  (not A169) );
 a52533a <=( A170  and  a52532a );
 a52537a <=( A201  and  A200 );
 a52538a <=( (not A199)  and  a52537a );
 a52539a <=( a52538a  and  a52533a );
 a52543a <=( A268  and  (not A267) );
 a52544a <=( A203  and  a52543a );
 a52547a <=( A299  and  (not A298) );
 a52550a <=( A301  and  A300 );
 a52551a <=( a52550a  and  a52547a );
 a52552a <=( a52551a  and  a52544a );
 a52556a <=( A168  and  (not A169) );
 a52557a <=( A170  and  a52556a );
 a52561a <=( A201  and  A200 );
 a52562a <=( (not A199)  and  a52561a );
 a52563a <=( a52562a  and  a52557a );
 a52567a <=( A268  and  (not A267) );
 a52568a <=( A203  and  a52567a );
 a52571a <=( A299  and  (not A298) );
 a52574a <=( A302  and  A300 );
 a52575a <=( a52574a  and  a52571a );
 a52576a <=( a52575a  and  a52568a );
 a52580a <=( A168  and  (not A169) );
 a52581a <=( A170  and  a52580a );
 a52585a <=( A201  and  A200 );
 a52586a <=( (not A199)  and  a52585a );
 a52587a <=( a52586a  and  a52581a );
 a52591a <=( A269  and  (not A267) );
 a52592a <=( A203  and  a52591a );
 a52595a <=( (not A299)  and  A298 );
 a52598a <=( A301  and  A300 );
 a52599a <=( a52598a  and  a52595a );
 a52600a <=( a52599a  and  a52592a );
 a52604a <=( A168  and  (not A169) );
 a52605a <=( A170  and  a52604a );
 a52609a <=( A201  and  A200 );
 a52610a <=( (not A199)  and  a52609a );
 a52611a <=( a52610a  and  a52605a );
 a52615a <=( A269  and  (not A267) );
 a52616a <=( A203  and  a52615a );
 a52619a <=( (not A299)  and  A298 );
 a52622a <=( A302  and  A300 );
 a52623a <=( a52622a  and  a52619a );
 a52624a <=( a52623a  and  a52616a );
 a52628a <=( A168  and  (not A169) );
 a52629a <=( A170  and  a52628a );
 a52633a <=( A201  and  A200 );
 a52634a <=( (not A199)  and  a52633a );
 a52635a <=( a52634a  and  a52629a );
 a52639a <=( A269  and  (not A267) );
 a52640a <=( A203  and  a52639a );
 a52643a <=( A299  and  (not A298) );
 a52646a <=( A301  and  A300 );
 a52647a <=( a52646a  and  a52643a );
 a52648a <=( a52647a  and  a52640a );
 a52652a <=( A168  and  (not A169) );
 a52653a <=( A170  and  a52652a );
 a52657a <=( A201  and  A200 );
 a52658a <=( (not A199)  and  a52657a );
 a52659a <=( a52658a  and  a52653a );
 a52663a <=( A269  and  (not A267) );
 a52664a <=( A203  and  a52663a );
 a52667a <=( A299  and  (not A298) );
 a52670a <=( A302  and  A300 );
 a52671a <=( a52670a  and  a52667a );
 a52672a <=( a52671a  and  a52664a );
 a52676a <=( A168  and  (not A169) );
 a52677a <=( A170  and  a52676a );
 a52681a <=( A201  and  A200 );
 a52682a <=( (not A199)  and  a52681a );
 a52683a <=( a52682a  and  a52677a );
 a52687a <=( A266  and  A265 );
 a52688a <=( A203  and  a52687a );
 a52691a <=( (not A299)  and  A298 );
 a52694a <=( A301  and  A300 );
 a52695a <=( a52694a  and  a52691a );
 a52696a <=( a52695a  and  a52688a );
 a52700a <=( A168  and  (not A169) );
 a52701a <=( A170  and  a52700a );
 a52705a <=( A201  and  A200 );
 a52706a <=( (not A199)  and  a52705a );
 a52707a <=( a52706a  and  a52701a );
 a52711a <=( A266  and  A265 );
 a52712a <=( A203  and  a52711a );
 a52715a <=( (not A299)  and  A298 );
 a52718a <=( A302  and  A300 );
 a52719a <=( a52718a  and  a52715a );
 a52720a <=( a52719a  and  a52712a );
 a52724a <=( A168  and  (not A169) );
 a52725a <=( A170  and  a52724a );
 a52729a <=( A201  and  A200 );
 a52730a <=( (not A199)  and  a52729a );
 a52731a <=( a52730a  and  a52725a );
 a52735a <=( A266  and  A265 );
 a52736a <=( A203  and  a52735a );
 a52739a <=( A299  and  (not A298) );
 a52742a <=( A301  and  A300 );
 a52743a <=( a52742a  and  a52739a );
 a52744a <=( a52743a  and  a52736a );
 a52748a <=( A168  and  (not A169) );
 a52749a <=( A170  and  a52748a );
 a52753a <=( A201  and  A200 );
 a52754a <=( (not A199)  and  a52753a );
 a52755a <=( a52754a  and  a52749a );
 a52759a <=( A266  and  A265 );
 a52760a <=( A203  and  a52759a );
 a52763a <=( A299  and  (not A298) );
 a52766a <=( A302  and  A300 );
 a52767a <=( a52766a  and  a52763a );
 a52768a <=( a52767a  and  a52760a );
 a52772a <=( A168  and  (not A169) );
 a52773a <=( A170  and  a52772a );
 a52777a <=( A201  and  A200 );
 a52778a <=( (not A199)  and  a52777a );
 a52779a <=( a52778a  and  a52773a );
 a52783a <=( (not A266)  and  (not A265) );
 a52784a <=( A203  and  a52783a );
 a52787a <=( (not A299)  and  A298 );
 a52790a <=( A301  and  A300 );
 a52791a <=( a52790a  and  a52787a );
 a52792a <=( a52791a  and  a52784a );
 a52796a <=( A168  and  (not A169) );
 a52797a <=( A170  and  a52796a );
 a52801a <=( A201  and  A200 );
 a52802a <=( (not A199)  and  a52801a );
 a52803a <=( a52802a  and  a52797a );
 a52807a <=( (not A266)  and  (not A265) );
 a52808a <=( A203  and  a52807a );
 a52811a <=( (not A299)  and  A298 );
 a52814a <=( A302  and  A300 );
 a52815a <=( a52814a  and  a52811a );
 a52816a <=( a52815a  and  a52808a );
 a52820a <=( A168  and  (not A169) );
 a52821a <=( A170  and  a52820a );
 a52825a <=( A201  and  A200 );
 a52826a <=( (not A199)  and  a52825a );
 a52827a <=( a52826a  and  a52821a );
 a52831a <=( (not A266)  and  (not A265) );
 a52832a <=( A203  and  a52831a );
 a52835a <=( A299  and  (not A298) );
 a52838a <=( A301  and  A300 );
 a52839a <=( a52838a  and  a52835a );
 a52840a <=( a52839a  and  a52832a );
 a52844a <=( A168  and  (not A169) );
 a52845a <=( A170  and  a52844a );
 a52849a <=( A201  and  A200 );
 a52850a <=( (not A199)  and  a52849a );
 a52851a <=( a52850a  and  a52845a );
 a52855a <=( (not A266)  and  (not A265) );
 a52856a <=( A203  and  a52855a );
 a52859a <=( A299  and  (not A298) );
 a52862a <=( A302  and  A300 );
 a52863a <=( a52862a  and  a52859a );
 a52864a <=( a52863a  and  a52856a );
 a52868a <=( A168  and  (not A169) );
 a52869a <=( A170  and  a52868a );
 a52873a <=( A201  and  (not A200) );
 a52874a <=( A199  and  a52873a );
 a52875a <=( a52874a  and  a52869a );
 a52879a <=( A268  and  (not A267) );
 a52880a <=( A202  and  a52879a );
 a52883a <=( (not A299)  and  A298 );
 a52886a <=( A301  and  A300 );
 a52887a <=( a52886a  and  a52883a );
 a52888a <=( a52887a  and  a52880a );
 a52892a <=( A168  and  (not A169) );
 a52893a <=( A170  and  a52892a );
 a52897a <=( A201  and  (not A200) );
 a52898a <=( A199  and  a52897a );
 a52899a <=( a52898a  and  a52893a );
 a52903a <=( A268  and  (not A267) );
 a52904a <=( A202  and  a52903a );
 a52907a <=( (not A299)  and  A298 );
 a52910a <=( A302  and  A300 );
 a52911a <=( a52910a  and  a52907a );
 a52912a <=( a52911a  and  a52904a );
 a52916a <=( A168  and  (not A169) );
 a52917a <=( A170  and  a52916a );
 a52921a <=( A201  and  (not A200) );
 a52922a <=( A199  and  a52921a );
 a52923a <=( a52922a  and  a52917a );
 a52927a <=( A268  and  (not A267) );
 a52928a <=( A202  and  a52927a );
 a52931a <=( A299  and  (not A298) );
 a52934a <=( A301  and  A300 );
 a52935a <=( a52934a  and  a52931a );
 a52936a <=( a52935a  and  a52928a );
 a52940a <=( A168  and  (not A169) );
 a52941a <=( A170  and  a52940a );
 a52945a <=( A201  and  (not A200) );
 a52946a <=( A199  and  a52945a );
 a52947a <=( a52946a  and  a52941a );
 a52951a <=( A268  and  (not A267) );
 a52952a <=( A202  and  a52951a );
 a52955a <=( A299  and  (not A298) );
 a52958a <=( A302  and  A300 );
 a52959a <=( a52958a  and  a52955a );
 a52960a <=( a52959a  and  a52952a );
 a52964a <=( A168  and  (not A169) );
 a52965a <=( A170  and  a52964a );
 a52969a <=( A201  and  (not A200) );
 a52970a <=( A199  and  a52969a );
 a52971a <=( a52970a  and  a52965a );
 a52975a <=( A269  and  (not A267) );
 a52976a <=( A202  and  a52975a );
 a52979a <=( (not A299)  and  A298 );
 a52982a <=( A301  and  A300 );
 a52983a <=( a52982a  and  a52979a );
 a52984a <=( a52983a  and  a52976a );
 a52988a <=( A168  and  (not A169) );
 a52989a <=( A170  and  a52988a );
 a52993a <=( A201  and  (not A200) );
 a52994a <=( A199  and  a52993a );
 a52995a <=( a52994a  and  a52989a );
 a52999a <=( A269  and  (not A267) );
 a53000a <=( A202  and  a52999a );
 a53003a <=( (not A299)  and  A298 );
 a53006a <=( A302  and  A300 );
 a53007a <=( a53006a  and  a53003a );
 a53008a <=( a53007a  and  a53000a );
 a53012a <=( A168  and  (not A169) );
 a53013a <=( A170  and  a53012a );
 a53017a <=( A201  and  (not A200) );
 a53018a <=( A199  and  a53017a );
 a53019a <=( a53018a  and  a53013a );
 a53023a <=( A269  and  (not A267) );
 a53024a <=( A202  and  a53023a );
 a53027a <=( A299  and  (not A298) );
 a53030a <=( A301  and  A300 );
 a53031a <=( a53030a  and  a53027a );
 a53032a <=( a53031a  and  a53024a );
 a53036a <=( A168  and  (not A169) );
 a53037a <=( A170  and  a53036a );
 a53041a <=( A201  and  (not A200) );
 a53042a <=( A199  and  a53041a );
 a53043a <=( a53042a  and  a53037a );
 a53047a <=( A269  and  (not A267) );
 a53048a <=( A202  and  a53047a );
 a53051a <=( A299  and  (not A298) );
 a53054a <=( A302  and  A300 );
 a53055a <=( a53054a  and  a53051a );
 a53056a <=( a53055a  and  a53048a );
 a53060a <=( A168  and  (not A169) );
 a53061a <=( A170  and  a53060a );
 a53065a <=( A201  and  (not A200) );
 a53066a <=( A199  and  a53065a );
 a53067a <=( a53066a  and  a53061a );
 a53071a <=( A266  and  A265 );
 a53072a <=( A202  and  a53071a );
 a53075a <=( (not A299)  and  A298 );
 a53078a <=( A301  and  A300 );
 a53079a <=( a53078a  and  a53075a );
 a53080a <=( a53079a  and  a53072a );
 a53084a <=( A168  and  (not A169) );
 a53085a <=( A170  and  a53084a );
 a53089a <=( A201  and  (not A200) );
 a53090a <=( A199  and  a53089a );
 a53091a <=( a53090a  and  a53085a );
 a53095a <=( A266  and  A265 );
 a53096a <=( A202  and  a53095a );
 a53099a <=( (not A299)  and  A298 );
 a53102a <=( A302  and  A300 );
 a53103a <=( a53102a  and  a53099a );
 a53104a <=( a53103a  and  a53096a );
 a53108a <=( A168  and  (not A169) );
 a53109a <=( A170  and  a53108a );
 a53113a <=( A201  and  (not A200) );
 a53114a <=( A199  and  a53113a );
 a53115a <=( a53114a  and  a53109a );
 a53119a <=( A266  and  A265 );
 a53120a <=( A202  and  a53119a );
 a53123a <=( A299  and  (not A298) );
 a53126a <=( A301  and  A300 );
 a53127a <=( a53126a  and  a53123a );
 a53128a <=( a53127a  and  a53120a );
 a53132a <=( A168  and  (not A169) );
 a53133a <=( A170  and  a53132a );
 a53137a <=( A201  and  (not A200) );
 a53138a <=( A199  and  a53137a );
 a53139a <=( a53138a  and  a53133a );
 a53143a <=( A266  and  A265 );
 a53144a <=( A202  and  a53143a );
 a53147a <=( A299  and  (not A298) );
 a53150a <=( A302  and  A300 );
 a53151a <=( a53150a  and  a53147a );
 a53152a <=( a53151a  and  a53144a );
 a53156a <=( A168  and  (not A169) );
 a53157a <=( A170  and  a53156a );
 a53161a <=( A201  and  (not A200) );
 a53162a <=( A199  and  a53161a );
 a53163a <=( a53162a  and  a53157a );
 a53167a <=( (not A266)  and  (not A265) );
 a53168a <=( A202  and  a53167a );
 a53171a <=( (not A299)  and  A298 );
 a53174a <=( A301  and  A300 );
 a53175a <=( a53174a  and  a53171a );
 a53176a <=( a53175a  and  a53168a );
 a53180a <=( A168  and  (not A169) );
 a53181a <=( A170  and  a53180a );
 a53185a <=( A201  and  (not A200) );
 a53186a <=( A199  and  a53185a );
 a53187a <=( a53186a  and  a53181a );
 a53191a <=( (not A266)  and  (not A265) );
 a53192a <=( A202  and  a53191a );
 a53195a <=( (not A299)  and  A298 );
 a53198a <=( A302  and  A300 );
 a53199a <=( a53198a  and  a53195a );
 a53200a <=( a53199a  and  a53192a );
 a53204a <=( A168  and  (not A169) );
 a53205a <=( A170  and  a53204a );
 a53209a <=( A201  and  (not A200) );
 a53210a <=( A199  and  a53209a );
 a53211a <=( a53210a  and  a53205a );
 a53215a <=( (not A266)  and  (not A265) );
 a53216a <=( A202  and  a53215a );
 a53219a <=( A299  and  (not A298) );
 a53222a <=( A301  and  A300 );
 a53223a <=( a53222a  and  a53219a );
 a53224a <=( a53223a  and  a53216a );
 a53228a <=( A168  and  (not A169) );
 a53229a <=( A170  and  a53228a );
 a53233a <=( A201  and  (not A200) );
 a53234a <=( A199  and  a53233a );
 a53235a <=( a53234a  and  a53229a );
 a53239a <=( (not A266)  and  (not A265) );
 a53240a <=( A202  and  a53239a );
 a53243a <=( A299  and  (not A298) );
 a53246a <=( A302  and  A300 );
 a53247a <=( a53246a  and  a53243a );
 a53248a <=( a53247a  and  a53240a );
 a53252a <=( A168  and  (not A169) );
 a53253a <=( A170  and  a53252a );
 a53257a <=( A201  and  (not A200) );
 a53258a <=( A199  and  a53257a );
 a53259a <=( a53258a  and  a53253a );
 a53263a <=( A268  and  (not A267) );
 a53264a <=( A203  and  a53263a );
 a53267a <=( (not A299)  and  A298 );
 a53270a <=( A301  and  A300 );
 a53271a <=( a53270a  and  a53267a );
 a53272a <=( a53271a  and  a53264a );
 a53276a <=( A168  and  (not A169) );
 a53277a <=( A170  and  a53276a );
 a53281a <=( A201  and  (not A200) );
 a53282a <=( A199  and  a53281a );
 a53283a <=( a53282a  and  a53277a );
 a53287a <=( A268  and  (not A267) );
 a53288a <=( A203  and  a53287a );
 a53291a <=( (not A299)  and  A298 );
 a53294a <=( A302  and  A300 );
 a53295a <=( a53294a  and  a53291a );
 a53296a <=( a53295a  and  a53288a );
 a53300a <=( A168  and  (not A169) );
 a53301a <=( A170  and  a53300a );
 a53305a <=( A201  and  (not A200) );
 a53306a <=( A199  and  a53305a );
 a53307a <=( a53306a  and  a53301a );
 a53311a <=( A268  and  (not A267) );
 a53312a <=( A203  and  a53311a );
 a53315a <=( A299  and  (not A298) );
 a53318a <=( A301  and  A300 );
 a53319a <=( a53318a  and  a53315a );
 a53320a <=( a53319a  and  a53312a );
 a53324a <=( A168  and  (not A169) );
 a53325a <=( A170  and  a53324a );
 a53329a <=( A201  and  (not A200) );
 a53330a <=( A199  and  a53329a );
 a53331a <=( a53330a  and  a53325a );
 a53335a <=( A268  and  (not A267) );
 a53336a <=( A203  and  a53335a );
 a53339a <=( A299  and  (not A298) );
 a53342a <=( A302  and  A300 );
 a53343a <=( a53342a  and  a53339a );
 a53344a <=( a53343a  and  a53336a );
 a53348a <=( A168  and  (not A169) );
 a53349a <=( A170  and  a53348a );
 a53353a <=( A201  and  (not A200) );
 a53354a <=( A199  and  a53353a );
 a53355a <=( a53354a  and  a53349a );
 a53359a <=( A269  and  (not A267) );
 a53360a <=( A203  and  a53359a );
 a53363a <=( (not A299)  and  A298 );
 a53366a <=( A301  and  A300 );
 a53367a <=( a53366a  and  a53363a );
 a53368a <=( a53367a  and  a53360a );
 a53372a <=( A168  and  (not A169) );
 a53373a <=( A170  and  a53372a );
 a53377a <=( A201  and  (not A200) );
 a53378a <=( A199  and  a53377a );
 a53379a <=( a53378a  and  a53373a );
 a53383a <=( A269  and  (not A267) );
 a53384a <=( A203  and  a53383a );
 a53387a <=( (not A299)  and  A298 );
 a53390a <=( A302  and  A300 );
 a53391a <=( a53390a  and  a53387a );
 a53392a <=( a53391a  and  a53384a );
 a53396a <=( A168  and  (not A169) );
 a53397a <=( A170  and  a53396a );
 a53401a <=( A201  and  (not A200) );
 a53402a <=( A199  and  a53401a );
 a53403a <=( a53402a  and  a53397a );
 a53407a <=( A269  and  (not A267) );
 a53408a <=( A203  and  a53407a );
 a53411a <=( A299  and  (not A298) );
 a53414a <=( A301  and  A300 );
 a53415a <=( a53414a  and  a53411a );
 a53416a <=( a53415a  and  a53408a );
 a53420a <=( A168  and  (not A169) );
 a53421a <=( A170  and  a53420a );
 a53425a <=( A201  and  (not A200) );
 a53426a <=( A199  and  a53425a );
 a53427a <=( a53426a  and  a53421a );
 a53431a <=( A269  and  (not A267) );
 a53432a <=( A203  and  a53431a );
 a53435a <=( A299  and  (not A298) );
 a53438a <=( A302  and  A300 );
 a53439a <=( a53438a  and  a53435a );
 a53440a <=( a53439a  and  a53432a );
 a53444a <=( A168  and  (not A169) );
 a53445a <=( A170  and  a53444a );
 a53449a <=( A201  and  (not A200) );
 a53450a <=( A199  and  a53449a );
 a53451a <=( a53450a  and  a53445a );
 a53455a <=( A266  and  A265 );
 a53456a <=( A203  and  a53455a );
 a53459a <=( (not A299)  and  A298 );
 a53462a <=( A301  and  A300 );
 a53463a <=( a53462a  and  a53459a );
 a53464a <=( a53463a  and  a53456a );
 a53468a <=( A168  and  (not A169) );
 a53469a <=( A170  and  a53468a );
 a53473a <=( A201  and  (not A200) );
 a53474a <=( A199  and  a53473a );
 a53475a <=( a53474a  and  a53469a );
 a53479a <=( A266  and  A265 );
 a53480a <=( A203  and  a53479a );
 a53483a <=( (not A299)  and  A298 );
 a53486a <=( A302  and  A300 );
 a53487a <=( a53486a  and  a53483a );
 a53488a <=( a53487a  and  a53480a );
 a53492a <=( A168  and  (not A169) );
 a53493a <=( A170  and  a53492a );
 a53497a <=( A201  and  (not A200) );
 a53498a <=( A199  and  a53497a );
 a53499a <=( a53498a  and  a53493a );
 a53503a <=( A266  and  A265 );
 a53504a <=( A203  and  a53503a );
 a53507a <=( A299  and  (not A298) );
 a53510a <=( A301  and  A300 );
 a53511a <=( a53510a  and  a53507a );
 a53512a <=( a53511a  and  a53504a );
 a53516a <=( A168  and  (not A169) );
 a53517a <=( A170  and  a53516a );
 a53521a <=( A201  and  (not A200) );
 a53522a <=( A199  and  a53521a );
 a53523a <=( a53522a  and  a53517a );
 a53527a <=( A266  and  A265 );
 a53528a <=( A203  and  a53527a );
 a53531a <=( A299  and  (not A298) );
 a53534a <=( A302  and  A300 );
 a53535a <=( a53534a  and  a53531a );
 a53536a <=( a53535a  and  a53528a );
 a53540a <=( A168  and  (not A169) );
 a53541a <=( A170  and  a53540a );
 a53545a <=( A201  and  (not A200) );
 a53546a <=( A199  and  a53545a );
 a53547a <=( a53546a  and  a53541a );
 a53551a <=( (not A266)  and  (not A265) );
 a53552a <=( A203  and  a53551a );
 a53555a <=( (not A299)  and  A298 );
 a53558a <=( A301  and  A300 );
 a53559a <=( a53558a  and  a53555a );
 a53560a <=( a53559a  and  a53552a );
 a53564a <=( A168  and  (not A169) );
 a53565a <=( A170  and  a53564a );
 a53569a <=( A201  and  (not A200) );
 a53570a <=( A199  and  a53569a );
 a53571a <=( a53570a  and  a53565a );
 a53575a <=( (not A266)  and  (not A265) );
 a53576a <=( A203  and  a53575a );
 a53579a <=( (not A299)  and  A298 );
 a53582a <=( A302  and  A300 );
 a53583a <=( a53582a  and  a53579a );
 a53584a <=( a53583a  and  a53576a );
 a53588a <=( A168  and  (not A169) );
 a53589a <=( A170  and  a53588a );
 a53593a <=( A201  and  (not A200) );
 a53594a <=( A199  and  a53593a );
 a53595a <=( a53594a  and  a53589a );
 a53599a <=( (not A266)  and  (not A265) );
 a53600a <=( A203  and  a53599a );
 a53603a <=( A299  and  (not A298) );
 a53606a <=( A301  and  A300 );
 a53607a <=( a53606a  and  a53603a );
 a53608a <=( a53607a  and  a53600a );
 a53612a <=( A168  and  (not A169) );
 a53613a <=( A170  and  a53612a );
 a53617a <=( A201  and  (not A200) );
 a53618a <=( A199  and  a53617a );
 a53619a <=( a53618a  and  a53613a );
 a53623a <=( (not A266)  and  (not A265) );
 a53624a <=( A203  and  a53623a );
 a53627a <=( A299  and  (not A298) );
 a53630a <=( A302  and  A300 );
 a53631a <=( a53630a  and  a53627a );
 a53632a <=( a53631a  and  a53624a );
 a53636a <=( A168  and  (not A169) );
 a53637a <=( A170  and  a53636a );
 a53641a <=( (not A265)  and  (not A200) );
 a53642a <=( (not A199)  and  a53641a );
 a53643a <=( a53642a  and  a53637a );
 a53647a <=( (not A268)  and  (not A267) );
 a53648a <=( A266  and  a53647a );
 a53651a <=( A300  and  (not A269) );
 a53654a <=( (not A302)  and  (not A301) );
 a53655a <=( a53654a  and  a53651a );
 a53656a <=( a53655a  and  a53648a );
 a53660a <=( A168  and  (not A169) );
 a53661a <=( A170  and  a53660a );
 a53665a <=( A265  and  (not A200) );
 a53666a <=( (not A199)  and  a53665a );
 a53667a <=( a53666a  and  a53661a );
 a53671a <=( (not A268)  and  (not A267) );
 a53672a <=( (not A266)  and  a53671a );
 a53675a <=( A300  and  (not A269) );
 a53678a <=( (not A302)  and  (not A301) );
 a53679a <=( a53678a  and  a53675a );
 a53680a <=( a53679a  and  a53672a );
 a53684a <=( (not A168)  and  (not A169) );
 a53685a <=( A170  and  a53684a );
 a53689a <=( (not A201)  and  (not A166) );
 a53690a <=( A167  and  a53689a );
 a53691a <=( a53690a  and  a53685a );
 a53695a <=( A268  and  (not A267) );
 a53696a <=( A202  and  a53695a );
 a53699a <=( (not A299)  and  A298 );
 a53702a <=( A301  and  A300 );
 a53703a <=( a53702a  and  a53699a );
 a53704a <=( a53703a  and  a53696a );
 a53708a <=( (not A168)  and  (not A169) );
 a53709a <=( A170  and  a53708a );
 a53713a <=( (not A201)  and  (not A166) );
 a53714a <=( A167  and  a53713a );
 a53715a <=( a53714a  and  a53709a );
 a53719a <=( A268  and  (not A267) );
 a53720a <=( A202  and  a53719a );
 a53723a <=( (not A299)  and  A298 );
 a53726a <=( A302  and  A300 );
 a53727a <=( a53726a  and  a53723a );
 a53728a <=( a53727a  and  a53720a );
 a53732a <=( (not A168)  and  (not A169) );
 a53733a <=( A170  and  a53732a );
 a53737a <=( (not A201)  and  (not A166) );
 a53738a <=( A167  and  a53737a );
 a53739a <=( a53738a  and  a53733a );
 a53743a <=( A268  and  (not A267) );
 a53744a <=( A202  and  a53743a );
 a53747a <=( A299  and  (not A298) );
 a53750a <=( A301  and  A300 );
 a53751a <=( a53750a  and  a53747a );
 a53752a <=( a53751a  and  a53744a );
 a53756a <=( (not A168)  and  (not A169) );
 a53757a <=( A170  and  a53756a );
 a53761a <=( (not A201)  and  (not A166) );
 a53762a <=( A167  and  a53761a );
 a53763a <=( a53762a  and  a53757a );
 a53767a <=( A268  and  (not A267) );
 a53768a <=( A202  and  a53767a );
 a53771a <=( A299  and  (not A298) );
 a53774a <=( A302  and  A300 );
 a53775a <=( a53774a  and  a53771a );
 a53776a <=( a53775a  and  a53768a );
 a53780a <=( (not A168)  and  (not A169) );
 a53781a <=( A170  and  a53780a );
 a53785a <=( (not A201)  and  (not A166) );
 a53786a <=( A167  and  a53785a );
 a53787a <=( a53786a  and  a53781a );
 a53791a <=( A269  and  (not A267) );
 a53792a <=( A202  and  a53791a );
 a53795a <=( (not A299)  and  A298 );
 a53798a <=( A301  and  A300 );
 a53799a <=( a53798a  and  a53795a );
 a53800a <=( a53799a  and  a53792a );
 a53804a <=( (not A168)  and  (not A169) );
 a53805a <=( A170  and  a53804a );
 a53809a <=( (not A201)  and  (not A166) );
 a53810a <=( A167  and  a53809a );
 a53811a <=( a53810a  and  a53805a );
 a53815a <=( A269  and  (not A267) );
 a53816a <=( A202  and  a53815a );
 a53819a <=( (not A299)  and  A298 );
 a53822a <=( A302  and  A300 );
 a53823a <=( a53822a  and  a53819a );
 a53824a <=( a53823a  and  a53816a );
 a53828a <=( (not A168)  and  (not A169) );
 a53829a <=( A170  and  a53828a );
 a53833a <=( (not A201)  and  (not A166) );
 a53834a <=( A167  and  a53833a );
 a53835a <=( a53834a  and  a53829a );
 a53839a <=( A269  and  (not A267) );
 a53840a <=( A202  and  a53839a );
 a53843a <=( A299  and  (not A298) );
 a53846a <=( A301  and  A300 );
 a53847a <=( a53846a  and  a53843a );
 a53848a <=( a53847a  and  a53840a );
 a53852a <=( (not A168)  and  (not A169) );
 a53853a <=( A170  and  a53852a );
 a53857a <=( (not A201)  and  (not A166) );
 a53858a <=( A167  and  a53857a );
 a53859a <=( a53858a  and  a53853a );
 a53863a <=( A269  and  (not A267) );
 a53864a <=( A202  and  a53863a );
 a53867a <=( A299  and  (not A298) );
 a53870a <=( A302  and  A300 );
 a53871a <=( a53870a  and  a53867a );
 a53872a <=( a53871a  and  a53864a );
 a53876a <=( (not A168)  and  (not A169) );
 a53877a <=( A170  and  a53876a );
 a53881a <=( (not A201)  and  (not A166) );
 a53882a <=( A167  and  a53881a );
 a53883a <=( a53882a  and  a53877a );
 a53887a <=( A266  and  A265 );
 a53888a <=( A202  and  a53887a );
 a53891a <=( (not A299)  and  A298 );
 a53894a <=( A301  and  A300 );
 a53895a <=( a53894a  and  a53891a );
 a53896a <=( a53895a  and  a53888a );
 a53900a <=( (not A168)  and  (not A169) );
 a53901a <=( A170  and  a53900a );
 a53905a <=( (not A201)  and  (not A166) );
 a53906a <=( A167  and  a53905a );
 a53907a <=( a53906a  and  a53901a );
 a53911a <=( A266  and  A265 );
 a53912a <=( A202  and  a53911a );
 a53915a <=( (not A299)  and  A298 );
 a53918a <=( A302  and  A300 );
 a53919a <=( a53918a  and  a53915a );
 a53920a <=( a53919a  and  a53912a );
 a53924a <=( (not A168)  and  (not A169) );
 a53925a <=( A170  and  a53924a );
 a53929a <=( (not A201)  and  (not A166) );
 a53930a <=( A167  and  a53929a );
 a53931a <=( a53930a  and  a53925a );
 a53935a <=( A266  and  A265 );
 a53936a <=( A202  and  a53935a );
 a53939a <=( A299  and  (not A298) );
 a53942a <=( A301  and  A300 );
 a53943a <=( a53942a  and  a53939a );
 a53944a <=( a53943a  and  a53936a );
 a53948a <=( (not A168)  and  (not A169) );
 a53949a <=( A170  and  a53948a );
 a53953a <=( (not A201)  and  (not A166) );
 a53954a <=( A167  and  a53953a );
 a53955a <=( a53954a  and  a53949a );
 a53959a <=( A266  and  A265 );
 a53960a <=( A202  and  a53959a );
 a53963a <=( A299  and  (not A298) );
 a53966a <=( A302  and  A300 );
 a53967a <=( a53966a  and  a53963a );
 a53968a <=( a53967a  and  a53960a );
 a53972a <=( (not A168)  and  (not A169) );
 a53973a <=( A170  and  a53972a );
 a53977a <=( (not A201)  and  (not A166) );
 a53978a <=( A167  and  a53977a );
 a53979a <=( a53978a  and  a53973a );
 a53983a <=( (not A266)  and  (not A265) );
 a53984a <=( A202  and  a53983a );
 a53987a <=( (not A299)  and  A298 );
 a53990a <=( A301  and  A300 );
 a53991a <=( a53990a  and  a53987a );
 a53992a <=( a53991a  and  a53984a );
 a53996a <=( (not A168)  and  (not A169) );
 a53997a <=( A170  and  a53996a );
 a54001a <=( (not A201)  and  (not A166) );
 a54002a <=( A167  and  a54001a );
 a54003a <=( a54002a  and  a53997a );
 a54007a <=( (not A266)  and  (not A265) );
 a54008a <=( A202  and  a54007a );
 a54011a <=( (not A299)  and  A298 );
 a54014a <=( A302  and  A300 );
 a54015a <=( a54014a  and  a54011a );
 a54016a <=( a54015a  and  a54008a );
 a54020a <=( (not A168)  and  (not A169) );
 a54021a <=( A170  and  a54020a );
 a54025a <=( (not A201)  and  (not A166) );
 a54026a <=( A167  and  a54025a );
 a54027a <=( a54026a  and  a54021a );
 a54031a <=( (not A266)  and  (not A265) );
 a54032a <=( A202  and  a54031a );
 a54035a <=( A299  and  (not A298) );
 a54038a <=( A301  and  A300 );
 a54039a <=( a54038a  and  a54035a );
 a54040a <=( a54039a  and  a54032a );
 a54044a <=( (not A168)  and  (not A169) );
 a54045a <=( A170  and  a54044a );
 a54049a <=( (not A201)  and  (not A166) );
 a54050a <=( A167  and  a54049a );
 a54051a <=( a54050a  and  a54045a );
 a54055a <=( (not A266)  and  (not A265) );
 a54056a <=( A202  and  a54055a );
 a54059a <=( A299  and  (not A298) );
 a54062a <=( A302  and  A300 );
 a54063a <=( a54062a  and  a54059a );
 a54064a <=( a54063a  and  a54056a );
 a54068a <=( (not A168)  and  (not A169) );
 a54069a <=( A170  and  a54068a );
 a54073a <=( (not A201)  and  (not A166) );
 a54074a <=( A167  and  a54073a );
 a54075a <=( a54074a  and  a54069a );
 a54079a <=( A268  and  (not A267) );
 a54080a <=( A203  and  a54079a );
 a54083a <=( (not A299)  and  A298 );
 a54086a <=( A301  and  A300 );
 a54087a <=( a54086a  and  a54083a );
 a54088a <=( a54087a  and  a54080a );
 a54092a <=( (not A168)  and  (not A169) );
 a54093a <=( A170  and  a54092a );
 a54097a <=( (not A201)  and  (not A166) );
 a54098a <=( A167  and  a54097a );
 a54099a <=( a54098a  and  a54093a );
 a54103a <=( A268  and  (not A267) );
 a54104a <=( A203  and  a54103a );
 a54107a <=( (not A299)  and  A298 );
 a54110a <=( A302  and  A300 );
 a54111a <=( a54110a  and  a54107a );
 a54112a <=( a54111a  and  a54104a );
 a54116a <=( (not A168)  and  (not A169) );
 a54117a <=( A170  and  a54116a );
 a54121a <=( (not A201)  and  (not A166) );
 a54122a <=( A167  and  a54121a );
 a54123a <=( a54122a  and  a54117a );
 a54127a <=( A268  and  (not A267) );
 a54128a <=( A203  and  a54127a );
 a54131a <=( A299  and  (not A298) );
 a54134a <=( A301  and  A300 );
 a54135a <=( a54134a  and  a54131a );
 a54136a <=( a54135a  and  a54128a );
 a54140a <=( (not A168)  and  (not A169) );
 a54141a <=( A170  and  a54140a );
 a54145a <=( (not A201)  and  (not A166) );
 a54146a <=( A167  and  a54145a );
 a54147a <=( a54146a  and  a54141a );
 a54151a <=( A268  and  (not A267) );
 a54152a <=( A203  and  a54151a );
 a54155a <=( A299  and  (not A298) );
 a54158a <=( A302  and  A300 );
 a54159a <=( a54158a  and  a54155a );
 a54160a <=( a54159a  and  a54152a );
 a54164a <=( (not A168)  and  (not A169) );
 a54165a <=( A170  and  a54164a );
 a54169a <=( (not A201)  and  (not A166) );
 a54170a <=( A167  and  a54169a );
 a54171a <=( a54170a  and  a54165a );
 a54175a <=( A269  and  (not A267) );
 a54176a <=( A203  and  a54175a );
 a54179a <=( (not A299)  and  A298 );
 a54182a <=( A301  and  A300 );
 a54183a <=( a54182a  and  a54179a );
 a54184a <=( a54183a  and  a54176a );
 a54188a <=( (not A168)  and  (not A169) );
 a54189a <=( A170  and  a54188a );
 a54193a <=( (not A201)  and  (not A166) );
 a54194a <=( A167  and  a54193a );
 a54195a <=( a54194a  and  a54189a );
 a54199a <=( A269  and  (not A267) );
 a54200a <=( A203  and  a54199a );
 a54203a <=( (not A299)  and  A298 );
 a54206a <=( A302  and  A300 );
 a54207a <=( a54206a  and  a54203a );
 a54208a <=( a54207a  and  a54200a );
 a54212a <=( (not A168)  and  (not A169) );
 a54213a <=( A170  and  a54212a );
 a54217a <=( (not A201)  and  (not A166) );
 a54218a <=( A167  and  a54217a );
 a54219a <=( a54218a  and  a54213a );
 a54223a <=( A269  and  (not A267) );
 a54224a <=( A203  and  a54223a );
 a54227a <=( A299  and  (not A298) );
 a54230a <=( A301  and  A300 );
 a54231a <=( a54230a  and  a54227a );
 a54232a <=( a54231a  and  a54224a );
 a54236a <=( (not A168)  and  (not A169) );
 a54237a <=( A170  and  a54236a );
 a54241a <=( (not A201)  and  (not A166) );
 a54242a <=( A167  and  a54241a );
 a54243a <=( a54242a  and  a54237a );
 a54247a <=( A269  and  (not A267) );
 a54248a <=( A203  and  a54247a );
 a54251a <=( A299  and  (not A298) );
 a54254a <=( A302  and  A300 );
 a54255a <=( a54254a  and  a54251a );
 a54256a <=( a54255a  and  a54248a );
 a54260a <=( (not A168)  and  (not A169) );
 a54261a <=( A170  and  a54260a );
 a54265a <=( (not A201)  and  (not A166) );
 a54266a <=( A167  and  a54265a );
 a54267a <=( a54266a  and  a54261a );
 a54271a <=( A266  and  A265 );
 a54272a <=( A203  and  a54271a );
 a54275a <=( (not A299)  and  A298 );
 a54278a <=( A301  and  A300 );
 a54279a <=( a54278a  and  a54275a );
 a54280a <=( a54279a  and  a54272a );
 a54284a <=( (not A168)  and  (not A169) );
 a54285a <=( A170  and  a54284a );
 a54289a <=( (not A201)  and  (not A166) );
 a54290a <=( A167  and  a54289a );
 a54291a <=( a54290a  and  a54285a );
 a54295a <=( A266  and  A265 );
 a54296a <=( A203  and  a54295a );
 a54299a <=( (not A299)  and  A298 );
 a54302a <=( A302  and  A300 );
 a54303a <=( a54302a  and  a54299a );
 a54304a <=( a54303a  and  a54296a );
 a54308a <=( (not A168)  and  (not A169) );
 a54309a <=( A170  and  a54308a );
 a54313a <=( (not A201)  and  (not A166) );
 a54314a <=( A167  and  a54313a );
 a54315a <=( a54314a  and  a54309a );
 a54319a <=( A266  and  A265 );
 a54320a <=( A203  and  a54319a );
 a54323a <=( A299  and  (not A298) );
 a54326a <=( A301  and  A300 );
 a54327a <=( a54326a  and  a54323a );
 a54328a <=( a54327a  and  a54320a );
 a54332a <=( (not A168)  and  (not A169) );
 a54333a <=( A170  and  a54332a );
 a54337a <=( (not A201)  and  (not A166) );
 a54338a <=( A167  and  a54337a );
 a54339a <=( a54338a  and  a54333a );
 a54343a <=( A266  and  A265 );
 a54344a <=( A203  and  a54343a );
 a54347a <=( A299  and  (not A298) );
 a54350a <=( A302  and  A300 );
 a54351a <=( a54350a  and  a54347a );
 a54352a <=( a54351a  and  a54344a );
 a54356a <=( (not A168)  and  (not A169) );
 a54357a <=( A170  and  a54356a );
 a54361a <=( (not A201)  and  (not A166) );
 a54362a <=( A167  and  a54361a );
 a54363a <=( a54362a  and  a54357a );
 a54367a <=( (not A266)  and  (not A265) );
 a54368a <=( A203  and  a54367a );
 a54371a <=( (not A299)  and  A298 );
 a54374a <=( A301  and  A300 );
 a54375a <=( a54374a  and  a54371a );
 a54376a <=( a54375a  and  a54368a );
 a54380a <=( (not A168)  and  (not A169) );
 a54381a <=( A170  and  a54380a );
 a54385a <=( (not A201)  and  (not A166) );
 a54386a <=( A167  and  a54385a );
 a54387a <=( a54386a  and  a54381a );
 a54391a <=( (not A266)  and  (not A265) );
 a54392a <=( A203  and  a54391a );
 a54395a <=( (not A299)  and  A298 );
 a54398a <=( A302  and  A300 );
 a54399a <=( a54398a  and  a54395a );
 a54400a <=( a54399a  and  a54392a );
 a54404a <=( (not A168)  and  (not A169) );
 a54405a <=( A170  and  a54404a );
 a54409a <=( (not A201)  and  (not A166) );
 a54410a <=( A167  and  a54409a );
 a54411a <=( a54410a  and  a54405a );
 a54415a <=( (not A266)  and  (not A265) );
 a54416a <=( A203  and  a54415a );
 a54419a <=( A299  and  (not A298) );
 a54422a <=( A301  and  A300 );
 a54423a <=( a54422a  and  a54419a );
 a54424a <=( a54423a  and  a54416a );
 a54428a <=( (not A168)  and  (not A169) );
 a54429a <=( A170  and  a54428a );
 a54433a <=( (not A201)  and  (not A166) );
 a54434a <=( A167  and  a54433a );
 a54435a <=( a54434a  and  a54429a );
 a54439a <=( (not A266)  and  (not A265) );
 a54440a <=( A203  and  a54439a );
 a54443a <=( A299  and  (not A298) );
 a54446a <=( A302  and  A300 );
 a54447a <=( a54446a  and  a54443a );
 a54448a <=( a54447a  and  a54440a );
 a54452a <=( (not A168)  and  (not A169) );
 a54453a <=( A170  and  a54452a );
 a54457a <=( A199  and  (not A166) );
 a54458a <=( A167  and  a54457a );
 a54459a <=( a54458a  and  a54453a );
 a54463a <=( A268  and  (not A267) );
 a54464a <=( A200  and  a54463a );
 a54467a <=( (not A299)  and  A298 );
 a54470a <=( A301  and  A300 );
 a54471a <=( a54470a  and  a54467a );
 a54472a <=( a54471a  and  a54464a );
 a54476a <=( (not A168)  and  (not A169) );
 a54477a <=( A170  and  a54476a );
 a54481a <=( A199  and  (not A166) );
 a54482a <=( A167  and  a54481a );
 a54483a <=( a54482a  and  a54477a );
 a54487a <=( A268  and  (not A267) );
 a54488a <=( A200  and  a54487a );
 a54491a <=( (not A299)  and  A298 );
 a54494a <=( A302  and  A300 );
 a54495a <=( a54494a  and  a54491a );
 a54496a <=( a54495a  and  a54488a );
 a54500a <=( (not A168)  and  (not A169) );
 a54501a <=( A170  and  a54500a );
 a54505a <=( A199  and  (not A166) );
 a54506a <=( A167  and  a54505a );
 a54507a <=( a54506a  and  a54501a );
 a54511a <=( A268  and  (not A267) );
 a54512a <=( A200  and  a54511a );
 a54515a <=( A299  and  (not A298) );
 a54518a <=( A301  and  A300 );
 a54519a <=( a54518a  and  a54515a );
 a54520a <=( a54519a  and  a54512a );
 a54524a <=( (not A168)  and  (not A169) );
 a54525a <=( A170  and  a54524a );
 a54529a <=( A199  and  (not A166) );
 a54530a <=( A167  and  a54529a );
 a54531a <=( a54530a  and  a54525a );
 a54535a <=( A268  and  (not A267) );
 a54536a <=( A200  and  a54535a );
 a54539a <=( A299  and  (not A298) );
 a54542a <=( A302  and  A300 );
 a54543a <=( a54542a  and  a54539a );
 a54544a <=( a54543a  and  a54536a );
 a54548a <=( (not A168)  and  (not A169) );
 a54549a <=( A170  and  a54548a );
 a54553a <=( A199  and  (not A166) );
 a54554a <=( A167  and  a54553a );
 a54555a <=( a54554a  and  a54549a );
 a54559a <=( A269  and  (not A267) );
 a54560a <=( A200  and  a54559a );
 a54563a <=( (not A299)  and  A298 );
 a54566a <=( A301  and  A300 );
 a54567a <=( a54566a  and  a54563a );
 a54568a <=( a54567a  and  a54560a );
 a54572a <=( (not A168)  and  (not A169) );
 a54573a <=( A170  and  a54572a );
 a54577a <=( A199  and  (not A166) );
 a54578a <=( A167  and  a54577a );
 a54579a <=( a54578a  and  a54573a );
 a54583a <=( A269  and  (not A267) );
 a54584a <=( A200  and  a54583a );
 a54587a <=( (not A299)  and  A298 );
 a54590a <=( A302  and  A300 );
 a54591a <=( a54590a  and  a54587a );
 a54592a <=( a54591a  and  a54584a );
 a54596a <=( (not A168)  and  (not A169) );
 a54597a <=( A170  and  a54596a );
 a54601a <=( A199  and  (not A166) );
 a54602a <=( A167  and  a54601a );
 a54603a <=( a54602a  and  a54597a );
 a54607a <=( A269  and  (not A267) );
 a54608a <=( A200  and  a54607a );
 a54611a <=( A299  and  (not A298) );
 a54614a <=( A301  and  A300 );
 a54615a <=( a54614a  and  a54611a );
 a54616a <=( a54615a  and  a54608a );
 a54620a <=( (not A168)  and  (not A169) );
 a54621a <=( A170  and  a54620a );
 a54625a <=( A199  and  (not A166) );
 a54626a <=( A167  and  a54625a );
 a54627a <=( a54626a  and  a54621a );
 a54631a <=( A269  and  (not A267) );
 a54632a <=( A200  and  a54631a );
 a54635a <=( A299  and  (not A298) );
 a54638a <=( A302  and  A300 );
 a54639a <=( a54638a  and  a54635a );
 a54640a <=( a54639a  and  a54632a );
 a54644a <=( (not A168)  and  (not A169) );
 a54645a <=( A170  and  a54644a );
 a54649a <=( A199  and  (not A166) );
 a54650a <=( A167  and  a54649a );
 a54651a <=( a54650a  and  a54645a );
 a54655a <=( A266  and  A265 );
 a54656a <=( A200  and  a54655a );
 a54659a <=( (not A299)  and  A298 );
 a54662a <=( A301  and  A300 );
 a54663a <=( a54662a  and  a54659a );
 a54664a <=( a54663a  and  a54656a );
 a54668a <=( (not A168)  and  (not A169) );
 a54669a <=( A170  and  a54668a );
 a54673a <=( A199  and  (not A166) );
 a54674a <=( A167  and  a54673a );
 a54675a <=( a54674a  and  a54669a );
 a54679a <=( A266  and  A265 );
 a54680a <=( A200  and  a54679a );
 a54683a <=( (not A299)  and  A298 );
 a54686a <=( A302  and  A300 );
 a54687a <=( a54686a  and  a54683a );
 a54688a <=( a54687a  and  a54680a );
 a54692a <=( (not A168)  and  (not A169) );
 a54693a <=( A170  and  a54692a );
 a54697a <=( A199  and  (not A166) );
 a54698a <=( A167  and  a54697a );
 a54699a <=( a54698a  and  a54693a );
 a54703a <=( A266  and  A265 );
 a54704a <=( A200  and  a54703a );
 a54707a <=( A299  and  (not A298) );
 a54710a <=( A301  and  A300 );
 a54711a <=( a54710a  and  a54707a );
 a54712a <=( a54711a  and  a54704a );
 a54716a <=( (not A168)  and  (not A169) );
 a54717a <=( A170  and  a54716a );
 a54721a <=( A199  and  (not A166) );
 a54722a <=( A167  and  a54721a );
 a54723a <=( a54722a  and  a54717a );
 a54727a <=( A266  and  A265 );
 a54728a <=( A200  and  a54727a );
 a54731a <=( A299  and  (not A298) );
 a54734a <=( A302  and  A300 );
 a54735a <=( a54734a  and  a54731a );
 a54736a <=( a54735a  and  a54728a );
 a54740a <=( (not A168)  and  (not A169) );
 a54741a <=( A170  and  a54740a );
 a54745a <=( A199  and  (not A166) );
 a54746a <=( A167  and  a54745a );
 a54747a <=( a54746a  and  a54741a );
 a54751a <=( (not A266)  and  (not A265) );
 a54752a <=( A200  and  a54751a );
 a54755a <=( (not A299)  and  A298 );
 a54758a <=( A301  and  A300 );
 a54759a <=( a54758a  and  a54755a );
 a54760a <=( a54759a  and  a54752a );
 a54764a <=( (not A168)  and  (not A169) );
 a54765a <=( A170  and  a54764a );
 a54769a <=( A199  and  (not A166) );
 a54770a <=( A167  and  a54769a );
 a54771a <=( a54770a  and  a54765a );
 a54775a <=( (not A266)  and  (not A265) );
 a54776a <=( A200  and  a54775a );
 a54779a <=( (not A299)  and  A298 );
 a54782a <=( A302  and  A300 );
 a54783a <=( a54782a  and  a54779a );
 a54784a <=( a54783a  and  a54776a );
 a54788a <=( (not A168)  and  (not A169) );
 a54789a <=( A170  and  a54788a );
 a54793a <=( A199  and  (not A166) );
 a54794a <=( A167  and  a54793a );
 a54795a <=( a54794a  and  a54789a );
 a54799a <=( (not A266)  and  (not A265) );
 a54800a <=( A200  and  a54799a );
 a54803a <=( A299  and  (not A298) );
 a54806a <=( A301  and  A300 );
 a54807a <=( a54806a  and  a54803a );
 a54808a <=( a54807a  and  a54800a );
 a54812a <=( (not A168)  and  (not A169) );
 a54813a <=( A170  and  a54812a );
 a54817a <=( A199  and  (not A166) );
 a54818a <=( A167  and  a54817a );
 a54819a <=( a54818a  and  a54813a );
 a54823a <=( (not A266)  and  (not A265) );
 a54824a <=( A200  and  a54823a );
 a54827a <=( A299  and  (not A298) );
 a54830a <=( A302  and  A300 );
 a54831a <=( a54830a  and  a54827a );
 a54832a <=( a54831a  and  a54824a );
 a54836a <=( (not A168)  and  (not A169) );
 a54837a <=( A170  and  a54836a );
 a54841a <=( (not A199)  and  (not A166) );
 a54842a <=( A167  and  a54841a );
 a54843a <=( a54842a  and  a54837a );
 a54847a <=( A268  and  (not A267) );
 a54848a <=( (not A200)  and  a54847a );
 a54851a <=( (not A299)  and  A298 );
 a54854a <=( A301  and  A300 );
 a54855a <=( a54854a  and  a54851a );
 a54856a <=( a54855a  and  a54848a );
 a54860a <=( (not A168)  and  (not A169) );
 a54861a <=( A170  and  a54860a );
 a54865a <=( (not A199)  and  (not A166) );
 a54866a <=( A167  and  a54865a );
 a54867a <=( a54866a  and  a54861a );
 a54871a <=( A268  and  (not A267) );
 a54872a <=( (not A200)  and  a54871a );
 a54875a <=( (not A299)  and  A298 );
 a54878a <=( A302  and  A300 );
 a54879a <=( a54878a  and  a54875a );
 a54880a <=( a54879a  and  a54872a );
 a54884a <=( (not A168)  and  (not A169) );
 a54885a <=( A170  and  a54884a );
 a54889a <=( (not A199)  and  (not A166) );
 a54890a <=( A167  and  a54889a );
 a54891a <=( a54890a  and  a54885a );
 a54895a <=( A268  and  (not A267) );
 a54896a <=( (not A200)  and  a54895a );
 a54899a <=( A299  and  (not A298) );
 a54902a <=( A301  and  A300 );
 a54903a <=( a54902a  and  a54899a );
 a54904a <=( a54903a  and  a54896a );
 a54908a <=( (not A168)  and  (not A169) );
 a54909a <=( A170  and  a54908a );
 a54913a <=( (not A199)  and  (not A166) );
 a54914a <=( A167  and  a54913a );
 a54915a <=( a54914a  and  a54909a );
 a54919a <=( A268  and  (not A267) );
 a54920a <=( (not A200)  and  a54919a );
 a54923a <=( A299  and  (not A298) );
 a54926a <=( A302  and  A300 );
 a54927a <=( a54926a  and  a54923a );
 a54928a <=( a54927a  and  a54920a );
 a54932a <=( (not A168)  and  (not A169) );
 a54933a <=( A170  and  a54932a );
 a54937a <=( (not A199)  and  (not A166) );
 a54938a <=( A167  and  a54937a );
 a54939a <=( a54938a  and  a54933a );
 a54943a <=( A269  and  (not A267) );
 a54944a <=( (not A200)  and  a54943a );
 a54947a <=( (not A299)  and  A298 );
 a54950a <=( A301  and  A300 );
 a54951a <=( a54950a  and  a54947a );
 a54952a <=( a54951a  and  a54944a );
 a54956a <=( (not A168)  and  (not A169) );
 a54957a <=( A170  and  a54956a );
 a54961a <=( (not A199)  and  (not A166) );
 a54962a <=( A167  and  a54961a );
 a54963a <=( a54962a  and  a54957a );
 a54967a <=( A269  and  (not A267) );
 a54968a <=( (not A200)  and  a54967a );
 a54971a <=( (not A299)  and  A298 );
 a54974a <=( A302  and  A300 );
 a54975a <=( a54974a  and  a54971a );
 a54976a <=( a54975a  and  a54968a );
 a54980a <=( (not A168)  and  (not A169) );
 a54981a <=( A170  and  a54980a );
 a54985a <=( (not A199)  and  (not A166) );
 a54986a <=( A167  and  a54985a );
 a54987a <=( a54986a  and  a54981a );
 a54991a <=( A269  and  (not A267) );
 a54992a <=( (not A200)  and  a54991a );
 a54995a <=( A299  and  (not A298) );
 a54998a <=( A301  and  A300 );
 a54999a <=( a54998a  and  a54995a );
 a55000a <=( a54999a  and  a54992a );
 a55004a <=( (not A168)  and  (not A169) );
 a55005a <=( A170  and  a55004a );
 a55009a <=( (not A199)  and  (not A166) );
 a55010a <=( A167  and  a55009a );
 a55011a <=( a55010a  and  a55005a );
 a55015a <=( A269  and  (not A267) );
 a55016a <=( (not A200)  and  a55015a );
 a55019a <=( A299  and  (not A298) );
 a55022a <=( A302  and  A300 );
 a55023a <=( a55022a  and  a55019a );
 a55024a <=( a55023a  and  a55016a );
 a55028a <=( (not A168)  and  (not A169) );
 a55029a <=( A170  and  a55028a );
 a55033a <=( (not A199)  and  (not A166) );
 a55034a <=( A167  and  a55033a );
 a55035a <=( a55034a  and  a55029a );
 a55039a <=( A266  and  A265 );
 a55040a <=( (not A200)  and  a55039a );
 a55043a <=( (not A299)  and  A298 );
 a55046a <=( A301  and  A300 );
 a55047a <=( a55046a  and  a55043a );
 a55048a <=( a55047a  and  a55040a );
 a55052a <=( (not A168)  and  (not A169) );
 a55053a <=( A170  and  a55052a );
 a55057a <=( (not A199)  and  (not A166) );
 a55058a <=( A167  and  a55057a );
 a55059a <=( a55058a  and  a55053a );
 a55063a <=( A266  and  A265 );
 a55064a <=( (not A200)  and  a55063a );
 a55067a <=( (not A299)  and  A298 );
 a55070a <=( A302  and  A300 );
 a55071a <=( a55070a  and  a55067a );
 a55072a <=( a55071a  and  a55064a );
 a55076a <=( (not A168)  and  (not A169) );
 a55077a <=( A170  and  a55076a );
 a55081a <=( (not A199)  and  (not A166) );
 a55082a <=( A167  and  a55081a );
 a55083a <=( a55082a  and  a55077a );
 a55087a <=( A266  and  A265 );
 a55088a <=( (not A200)  and  a55087a );
 a55091a <=( A299  and  (not A298) );
 a55094a <=( A301  and  A300 );
 a55095a <=( a55094a  and  a55091a );
 a55096a <=( a55095a  and  a55088a );
 a55100a <=( (not A168)  and  (not A169) );
 a55101a <=( A170  and  a55100a );
 a55105a <=( (not A199)  and  (not A166) );
 a55106a <=( A167  and  a55105a );
 a55107a <=( a55106a  and  a55101a );
 a55111a <=( A266  and  A265 );
 a55112a <=( (not A200)  and  a55111a );
 a55115a <=( A299  and  (not A298) );
 a55118a <=( A302  and  A300 );
 a55119a <=( a55118a  and  a55115a );
 a55120a <=( a55119a  and  a55112a );
 a55124a <=( (not A168)  and  (not A169) );
 a55125a <=( A170  and  a55124a );
 a55129a <=( (not A199)  and  (not A166) );
 a55130a <=( A167  and  a55129a );
 a55131a <=( a55130a  and  a55125a );
 a55135a <=( (not A266)  and  (not A265) );
 a55136a <=( (not A200)  and  a55135a );
 a55139a <=( (not A299)  and  A298 );
 a55142a <=( A301  and  A300 );
 a55143a <=( a55142a  and  a55139a );
 a55144a <=( a55143a  and  a55136a );
 a55148a <=( (not A168)  and  (not A169) );
 a55149a <=( A170  and  a55148a );
 a55153a <=( (not A199)  and  (not A166) );
 a55154a <=( A167  and  a55153a );
 a55155a <=( a55154a  and  a55149a );
 a55159a <=( (not A266)  and  (not A265) );
 a55160a <=( (not A200)  and  a55159a );
 a55163a <=( (not A299)  and  A298 );
 a55166a <=( A302  and  A300 );
 a55167a <=( a55166a  and  a55163a );
 a55168a <=( a55167a  and  a55160a );
 a55172a <=( (not A168)  and  (not A169) );
 a55173a <=( A170  and  a55172a );
 a55177a <=( (not A199)  and  (not A166) );
 a55178a <=( A167  and  a55177a );
 a55179a <=( a55178a  and  a55173a );
 a55183a <=( (not A266)  and  (not A265) );
 a55184a <=( (not A200)  and  a55183a );
 a55187a <=( A299  and  (not A298) );
 a55190a <=( A301  and  A300 );
 a55191a <=( a55190a  and  a55187a );
 a55192a <=( a55191a  and  a55184a );
 a55196a <=( (not A168)  and  (not A169) );
 a55197a <=( A170  and  a55196a );
 a55201a <=( (not A199)  and  (not A166) );
 a55202a <=( A167  and  a55201a );
 a55203a <=( a55202a  and  a55197a );
 a55207a <=( (not A266)  and  (not A265) );
 a55208a <=( (not A200)  and  a55207a );
 a55211a <=( A299  and  (not A298) );
 a55214a <=( A302  and  A300 );
 a55215a <=( a55214a  and  a55211a );
 a55216a <=( a55215a  and  a55208a );
 a55220a <=( (not A168)  and  (not A169) );
 a55221a <=( A170  and  a55220a );
 a55225a <=( (not A201)  and  A166 );
 a55226a <=( (not A167)  and  a55225a );
 a55227a <=( a55226a  and  a55221a );
 a55231a <=( A268  and  (not A267) );
 a55232a <=( A202  and  a55231a );
 a55235a <=( (not A299)  and  A298 );
 a55238a <=( A301  and  A300 );
 a55239a <=( a55238a  and  a55235a );
 a55240a <=( a55239a  and  a55232a );
 a55244a <=( (not A168)  and  (not A169) );
 a55245a <=( A170  and  a55244a );
 a55249a <=( (not A201)  and  A166 );
 a55250a <=( (not A167)  and  a55249a );
 a55251a <=( a55250a  and  a55245a );
 a55255a <=( A268  and  (not A267) );
 a55256a <=( A202  and  a55255a );
 a55259a <=( (not A299)  and  A298 );
 a55262a <=( A302  and  A300 );
 a55263a <=( a55262a  and  a55259a );
 a55264a <=( a55263a  and  a55256a );
 a55268a <=( (not A168)  and  (not A169) );
 a55269a <=( A170  and  a55268a );
 a55273a <=( (not A201)  and  A166 );
 a55274a <=( (not A167)  and  a55273a );
 a55275a <=( a55274a  and  a55269a );
 a55279a <=( A268  and  (not A267) );
 a55280a <=( A202  and  a55279a );
 a55283a <=( A299  and  (not A298) );
 a55286a <=( A301  and  A300 );
 a55287a <=( a55286a  and  a55283a );
 a55288a <=( a55287a  and  a55280a );
 a55292a <=( (not A168)  and  (not A169) );
 a55293a <=( A170  and  a55292a );
 a55297a <=( (not A201)  and  A166 );
 a55298a <=( (not A167)  and  a55297a );
 a55299a <=( a55298a  and  a55293a );
 a55303a <=( A268  and  (not A267) );
 a55304a <=( A202  and  a55303a );
 a55307a <=( A299  and  (not A298) );
 a55310a <=( A302  and  A300 );
 a55311a <=( a55310a  and  a55307a );
 a55312a <=( a55311a  and  a55304a );
 a55316a <=( (not A168)  and  (not A169) );
 a55317a <=( A170  and  a55316a );
 a55321a <=( (not A201)  and  A166 );
 a55322a <=( (not A167)  and  a55321a );
 a55323a <=( a55322a  and  a55317a );
 a55327a <=( A269  and  (not A267) );
 a55328a <=( A202  and  a55327a );
 a55331a <=( (not A299)  and  A298 );
 a55334a <=( A301  and  A300 );
 a55335a <=( a55334a  and  a55331a );
 a55336a <=( a55335a  and  a55328a );
 a55340a <=( (not A168)  and  (not A169) );
 a55341a <=( A170  and  a55340a );
 a55345a <=( (not A201)  and  A166 );
 a55346a <=( (not A167)  and  a55345a );
 a55347a <=( a55346a  and  a55341a );
 a55351a <=( A269  and  (not A267) );
 a55352a <=( A202  and  a55351a );
 a55355a <=( (not A299)  and  A298 );
 a55358a <=( A302  and  A300 );
 a55359a <=( a55358a  and  a55355a );
 a55360a <=( a55359a  and  a55352a );
 a55364a <=( (not A168)  and  (not A169) );
 a55365a <=( A170  and  a55364a );
 a55369a <=( (not A201)  and  A166 );
 a55370a <=( (not A167)  and  a55369a );
 a55371a <=( a55370a  and  a55365a );
 a55375a <=( A269  and  (not A267) );
 a55376a <=( A202  and  a55375a );
 a55379a <=( A299  and  (not A298) );
 a55382a <=( A301  and  A300 );
 a55383a <=( a55382a  and  a55379a );
 a55384a <=( a55383a  and  a55376a );
 a55388a <=( (not A168)  and  (not A169) );
 a55389a <=( A170  and  a55388a );
 a55393a <=( (not A201)  and  A166 );
 a55394a <=( (not A167)  and  a55393a );
 a55395a <=( a55394a  and  a55389a );
 a55399a <=( A269  and  (not A267) );
 a55400a <=( A202  and  a55399a );
 a55403a <=( A299  and  (not A298) );
 a55406a <=( A302  and  A300 );
 a55407a <=( a55406a  and  a55403a );
 a55408a <=( a55407a  and  a55400a );
 a55412a <=( (not A168)  and  (not A169) );
 a55413a <=( A170  and  a55412a );
 a55417a <=( (not A201)  and  A166 );
 a55418a <=( (not A167)  and  a55417a );
 a55419a <=( a55418a  and  a55413a );
 a55423a <=( A266  and  A265 );
 a55424a <=( A202  and  a55423a );
 a55427a <=( (not A299)  and  A298 );
 a55430a <=( A301  and  A300 );
 a55431a <=( a55430a  and  a55427a );
 a55432a <=( a55431a  and  a55424a );
 a55436a <=( (not A168)  and  (not A169) );
 a55437a <=( A170  and  a55436a );
 a55441a <=( (not A201)  and  A166 );
 a55442a <=( (not A167)  and  a55441a );
 a55443a <=( a55442a  and  a55437a );
 a55447a <=( A266  and  A265 );
 a55448a <=( A202  and  a55447a );
 a55451a <=( (not A299)  and  A298 );
 a55454a <=( A302  and  A300 );
 a55455a <=( a55454a  and  a55451a );
 a55456a <=( a55455a  and  a55448a );
 a55460a <=( (not A168)  and  (not A169) );
 a55461a <=( A170  and  a55460a );
 a55465a <=( (not A201)  and  A166 );
 a55466a <=( (not A167)  and  a55465a );
 a55467a <=( a55466a  and  a55461a );
 a55471a <=( A266  and  A265 );
 a55472a <=( A202  and  a55471a );
 a55475a <=( A299  and  (not A298) );
 a55478a <=( A301  and  A300 );
 a55479a <=( a55478a  and  a55475a );
 a55480a <=( a55479a  and  a55472a );
 a55484a <=( (not A168)  and  (not A169) );
 a55485a <=( A170  and  a55484a );
 a55489a <=( (not A201)  and  A166 );
 a55490a <=( (not A167)  and  a55489a );
 a55491a <=( a55490a  and  a55485a );
 a55495a <=( A266  and  A265 );
 a55496a <=( A202  and  a55495a );
 a55499a <=( A299  and  (not A298) );
 a55502a <=( A302  and  A300 );
 a55503a <=( a55502a  and  a55499a );
 a55504a <=( a55503a  and  a55496a );
 a55508a <=( (not A168)  and  (not A169) );
 a55509a <=( A170  and  a55508a );
 a55513a <=( (not A201)  and  A166 );
 a55514a <=( (not A167)  and  a55513a );
 a55515a <=( a55514a  and  a55509a );
 a55519a <=( (not A266)  and  (not A265) );
 a55520a <=( A202  and  a55519a );
 a55523a <=( (not A299)  and  A298 );
 a55526a <=( A301  and  A300 );
 a55527a <=( a55526a  and  a55523a );
 a55528a <=( a55527a  and  a55520a );
 a55532a <=( (not A168)  and  (not A169) );
 a55533a <=( A170  and  a55532a );
 a55537a <=( (not A201)  and  A166 );
 a55538a <=( (not A167)  and  a55537a );
 a55539a <=( a55538a  and  a55533a );
 a55543a <=( (not A266)  and  (not A265) );
 a55544a <=( A202  and  a55543a );
 a55547a <=( (not A299)  and  A298 );
 a55550a <=( A302  and  A300 );
 a55551a <=( a55550a  and  a55547a );
 a55552a <=( a55551a  and  a55544a );
 a55556a <=( (not A168)  and  (not A169) );
 a55557a <=( A170  and  a55556a );
 a55561a <=( (not A201)  and  A166 );
 a55562a <=( (not A167)  and  a55561a );
 a55563a <=( a55562a  and  a55557a );
 a55567a <=( (not A266)  and  (not A265) );
 a55568a <=( A202  and  a55567a );
 a55571a <=( A299  and  (not A298) );
 a55574a <=( A301  and  A300 );
 a55575a <=( a55574a  and  a55571a );
 a55576a <=( a55575a  and  a55568a );
 a55580a <=( (not A168)  and  (not A169) );
 a55581a <=( A170  and  a55580a );
 a55585a <=( (not A201)  and  A166 );
 a55586a <=( (not A167)  and  a55585a );
 a55587a <=( a55586a  and  a55581a );
 a55591a <=( (not A266)  and  (not A265) );
 a55592a <=( A202  and  a55591a );
 a55595a <=( A299  and  (not A298) );
 a55598a <=( A302  and  A300 );
 a55599a <=( a55598a  and  a55595a );
 a55600a <=( a55599a  and  a55592a );
 a55604a <=( (not A168)  and  (not A169) );
 a55605a <=( A170  and  a55604a );
 a55609a <=( (not A201)  and  A166 );
 a55610a <=( (not A167)  and  a55609a );
 a55611a <=( a55610a  and  a55605a );
 a55615a <=( A268  and  (not A267) );
 a55616a <=( A203  and  a55615a );
 a55619a <=( (not A299)  and  A298 );
 a55622a <=( A301  and  A300 );
 a55623a <=( a55622a  and  a55619a );
 a55624a <=( a55623a  and  a55616a );
 a55628a <=( (not A168)  and  (not A169) );
 a55629a <=( A170  and  a55628a );
 a55633a <=( (not A201)  and  A166 );
 a55634a <=( (not A167)  and  a55633a );
 a55635a <=( a55634a  and  a55629a );
 a55639a <=( A268  and  (not A267) );
 a55640a <=( A203  and  a55639a );
 a55643a <=( (not A299)  and  A298 );
 a55646a <=( A302  and  A300 );
 a55647a <=( a55646a  and  a55643a );
 a55648a <=( a55647a  and  a55640a );
 a55652a <=( (not A168)  and  (not A169) );
 a55653a <=( A170  and  a55652a );
 a55657a <=( (not A201)  and  A166 );
 a55658a <=( (not A167)  and  a55657a );
 a55659a <=( a55658a  and  a55653a );
 a55663a <=( A268  and  (not A267) );
 a55664a <=( A203  and  a55663a );
 a55667a <=( A299  and  (not A298) );
 a55670a <=( A301  and  A300 );
 a55671a <=( a55670a  and  a55667a );
 a55672a <=( a55671a  and  a55664a );
 a55676a <=( (not A168)  and  (not A169) );
 a55677a <=( A170  and  a55676a );
 a55681a <=( (not A201)  and  A166 );
 a55682a <=( (not A167)  and  a55681a );
 a55683a <=( a55682a  and  a55677a );
 a55687a <=( A268  and  (not A267) );
 a55688a <=( A203  and  a55687a );
 a55691a <=( A299  and  (not A298) );
 a55694a <=( A302  and  A300 );
 a55695a <=( a55694a  and  a55691a );
 a55696a <=( a55695a  and  a55688a );
 a55700a <=( (not A168)  and  (not A169) );
 a55701a <=( A170  and  a55700a );
 a55705a <=( (not A201)  and  A166 );
 a55706a <=( (not A167)  and  a55705a );
 a55707a <=( a55706a  and  a55701a );
 a55711a <=( A269  and  (not A267) );
 a55712a <=( A203  and  a55711a );
 a55715a <=( (not A299)  and  A298 );
 a55718a <=( A301  and  A300 );
 a55719a <=( a55718a  and  a55715a );
 a55720a <=( a55719a  and  a55712a );
 a55724a <=( (not A168)  and  (not A169) );
 a55725a <=( A170  and  a55724a );
 a55729a <=( (not A201)  and  A166 );
 a55730a <=( (not A167)  and  a55729a );
 a55731a <=( a55730a  and  a55725a );
 a55735a <=( A269  and  (not A267) );
 a55736a <=( A203  and  a55735a );
 a55739a <=( (not A299)  and  A298 );
 a55742a <=( A302  and  A300 );
 a55743a <=( a55742a  and  a55739a );
 a55744a <=( a55743a  and  a55736a );
 a55748a <=( (not A168)  and  (not A169) );
 a55749a <=( A170  and  a55748a );
 a55753a <=( (not A201)  and  A166 );
 a55754a <=( (not A167)  and  a55753a );
 a55755a <=( a55754a  and  a55749a );
 a55759a <=( A269  and  (not A267) );
 a55760a <=( A203  and  a55759a );
 a55763a <=( A299  and  (not A298) );
 a55766a <=( A301  and  A300 );
 a55767a <=( a55766a  and  a55763a );
 a55768a <=( a55767a  and  a55760a );
 a55772a <=( (not A168)  and  (not A169) );
 a55773a <=( A170  and  a55772a );
 a55777a <=( (not A201)  and  A166 );
 a55778a <=( (not A167)  and  a55777a );
 a55779a <=( a55778a  and  a55773a );
 a55783a <=( A269  and  (not A267) );
 a55784a <=( A203  and  a55783a );
 a55787a <=( A299  and  (not A298) );
 a55790a <=( A302  and  A300 );
 a55791a <=( a55790a  and  a55787a );
 a55792a <=( a55791a  and  a55784a );
 a55796a <=( (not A168)  and  (not A169) );
 a55797a <=( A170  and  a55796a );
 a55801a <=( (not A201)  and  A166 );
 a55802a <=( (not A167)  and  a55801a );
 a55803a <=( a55802a  and  a55797a );
 a55807a <=( A266  and  A265 );
 a55808a <=( A203  and  a55807a );
 a55811a <=( (not A299)  and  A298 );
 a55814a <=( A301  and  A300 );
 a55815a <=( a55814a  and  a55811a );
 a55816a <=( a55815a  and  a55808a );
 a55820a <=( (not A168)  and  (not A169) );
 a55821a <=( A170  and  a55820a );
 a55825a <=( (not A201)  and  A166 );
 a55826a <=( (not A167)  and  a55825a );
 a55827a <=( a55826a  and  a55821a );
 a55831a <=( A266  and  A265 );
 a55832a <=( A203  and  a55831a );
 a55835a <=( (not A299)  and  A298 );
 a55838a <=( A302  and  A300 );
 a55839a <=( a55838a  and  a55835a );
 a55840a <=( a55839a  and  a55832a );
 a55844a <=( (not A168)  and  (not A169) );
 a55845a <=( A170  and  a55844a );
 a55849a <=( (not A201)  and  A166 );
 a55850a <=( (not A167)  and  a55849a );
 a55851a <=( a55850a  and  a55845a );
 a55855a <=( A266  and  A265 );
 a55856a <=( A203  and  a55855a );
 a55859a <=( A299  and  (not A298) );
 a55862a <=( A301  and  A300 );
 a55863a <=( a55862a  and  a55859a );
 a55864a <=( a55863a  and  a55856a );
 a55868a <=( (not A168)  and  (not A169) );
 a55869a <=( A170  and  a55868a );
 a55873a <=( (not A201)  and  A166 );
 a55874a <=( (not A167)  and  a55873a );
 a55875a <=( a55874a  and  a55869a );
 a55879a <=( A266  and  A265 );
 a55880a <=( A203  and  a55879a );
 a55883a <=( A299  and  (not A298) );
 a55886a <=( A302  and  A300 );
 a55887a <=( a55886a  and  a55883a );
 a55888a <=( a55887a  and  a55880a );
 a55892a <=( (not A168)  and  (not A169) );
 a55893a <=( A170  and  a55892a );
 a55897a <=( (not A201)  and  A166 );
 a55898a <=( (not A167)  and  a55897a );
 a55899a <=( a55898a  and  a55893a );
 a55903a <=( (not A266)  and  (not A265) );
 a55904a <=( A203  and  a55903a );
 a55907a <=( (not A299)  and  A298 );
 a55910a <=( A301  and  A300 );
 a55911a <=( a55910a  and  a55907a );
 a55912a <=( a55911a  and  a55904a );
 a55916a <=( (not A168)  and  (not A169) );
 a55917a <=( A170  and  a55916a );
 a55921a <=( (not A201)  and  A166 );
 a55922a <=( (not A167)  and  a55921a );
 a55923a <=( a55922a  and  a55917a );
 a55927a <=( (not A266)  and  (not A265) );
 a55928a <=( A203  and  a55927a );
 a55931a <=( (not A299)  and  A298 );
 a55934a <=( A302  and  A300 );
 a55935a <=( a55934a  and  a55931a );
 a55936a <=( a55935a  and  a55928a );
 a55940a <=( (not A168)  and  (not A169) );
 a55941a <=( A170  and  a55940a );
 a55945a <=( (not A201)  and  A166 );
 a55946a <=( (not A167)  and  a55945a );
 a55947a <=( a55946a  and  a55941a );
 a55951a <=( (not A266)  and  (not A265) );
 a55952a <=( A203  and  a55951a );
 a55955a <=( A299  and  (not A298) );
 a55958a <=( A301  and  A300 );
 a55959a <=( a55958a  and  a55955a );
 a55960a <=( a55959a  and  a55952a );
 a55964a <=( (not A168)  and  (not A169) );
 a55965a <=( A170  and  a55964a );
 a55969a <=( (not A201)  and  A166 );
 a55970a <=( (not A167)  and  a55969a );
 a55971a <=( a55970a  and  a55965a );
 a55975a <=( (not A266)  and  (not A265) );
 a55976a <=( A203  and  a55975a );
 a55979a <=( A299  and  (not A298) );
 a55982a <=( A302  and  A300 );
 a55983a <=( a55982a  and  a55979a );
 a55984a <=( a55983a  and  a55976a );
 a55988a <=( (not A168)  and  (not A169) );
 a55989a <=( A170  and  a55988a );
 a55993a <=( A199  and  A166 );
 a55994a <=( (not A167)  and  a55993a );
 a55995a <=( a55994a  and  a55989a );
 a55999a <=( A268  and  (not A267) );
 a56000a <=( A200  and  a55999a );
 a56003a <=( (not A299)  and  A298 );
 a56006a <=( A301  and  A300 );
 a56007a <=( a56006a  and  a56003a );
 a56008a <=( a56007a  and  a56000a );
 a56012a <=( (not A168)  and  (not A169) );
 a56013a <=( A170  and  a56012a );
 a56017a <=( A199  and  A166 );
 a56018a <=( (not A167)  and  a56017a );
 a56019a <=( a56018a  and  a56013a );
 a56023a <=( A268  and  (not A267) );
 a56024a <=( A200  and  a56023a );
 a56027a <=( (not A299)  and  A298 );
 a56030a <=( A302  and  A300 );
 a56031a <=( a56030a  and  a56027a );
 a56032a <=( a56031a  and  a56024a );
 a56036a <=( (not A168)  and  (not A169) );
 a56037a <=( A170  and  a56036a );
 a56041a <=( A199  and  A166 );
 a56042a <=( (not A167)  and  a56041a );
 a56043a <=( a56042a  and  a56037a );
 a56047a <=( A268  and  (not A267) );
 a56048a <=( A200  and  a56047a );
 a56051a <=( A299  and  (not A298) );
 a56054a <=( A301  and  A300 );
 a56055a <=( a56054a  and  a56051a );
 a56056a <=( a56055a  and  a56048a );
 a56060a <=( (not A168)  and  (not A169) );
 a56061a <=( A170  and  a56060a );
 a56065a <=( A199  and  A166 );
 a56066a <=( (not A167)  and  a56065a );
 a56067a <=( a56066a  and  a56061a );
 a56071a <=( A268  and  (not A267) );
 a56072a <=( A200  and  a56071a );
 a56075a <=( A299  and  (not A298) );
 a56078a <=( A302  and  A300 );
 a56079a <=( a56078a  and  a56075a );
 a56080a <=( a56079a  and  a56072a );
 a56084a <=( (not A168)  and  (not A169) );
 a56085a <=( A170  and  a56084a );
 a56089a <=( A199  and  A166 );
 a56090a <=( (not A167)  and  a56089a );
 a56091a <=( a56090a  and  a56085a );
 a56095a <=( A269  and  (not A267) );
 a56096a <=( A200  and  a56095a );
 a56099a <=( (not A299)  and  A298 );
 a56102a <=( A301  and  A300 );
 a56103a <=( a56102a  and  a56099a );
 a56104a <=( a56103a  and  a56096a );
 a56108a <=( (not A168)  and  (not A169) );
 a56109a <=( A170  and  a56108a );
 a56113a <=( A199  and  A166 );
 a56114a <=( (not A167)  and  a56113a );
 a56115a <=( a56114a  and  a56109a );
 a56119a <=( A269  and  (not A267) );
 a56120a <=( A200  and  a56119a );
 a56123a <=( (not A299)  and  A298 );
 a56126a <=( A302  and  A300 );
 a56127a <=( a56126a  and  a56123a );
 a56128a <=( a56127a  and  a56120a );
 a56132a <=( (not A168)  and  (not A169) );
 a56133a <=( A170  and  a56132a );
 a56137a <=( A199  and  A166 );
 a56138a <=( (not A167)  and  a56137a );
 a56139a <=( a56138a  and  a56133a );
 a56143a <=( A269  and  (not A267) );
 a56144a <=( A200  and  a56143a );
 a56147a <=( A299  and  (not A298) );
 a56150a <=( A301  and  A300 );
 a56151a <=( a56150a  and  a56147a );
 a56152a <=( a56151a  and  a56144a );
 a56156a <=( (not A168)  and  (not A169) );
 a56157a <=( A170  and  a56156a );
 a56161a <=( A199  and  A166 );
 a56162a <=( (not A167)  and  a56161a );
 a56163a <=( a56162a  and  a56157a );
 a56167a <=( A269  and  (not A267) );
 a56168a <=( A200  and  a56167a );
 a56171a <=( A299  and  (not A298) );
 a56174a <=( A302  and  A300 );
 a56175a <=( a56174a  and  a56171a );
 a56176a <=( a56175a  and  a56168a );
 a56180a <=( (not A168)  and  (not A169) );
 a56181a <=( A170  and  a56180a );
 a56185a <=( A199  and  A166 );
 a56186a <=( (not A167)  and  a56185a );
 a56187a <=( a56186a  and  a56181a );
 a56191a <=( A266  and  A265 );
 a56192a <=( A200  and  a56191a );
 a56195a <=( (not A299)  and  A298 );
 a56198a <=( A301  and  A300 );
 a56199a <=( a56198a  and  a56195a );
 a56200a <=( a56199a  and  a56192a );
 a56204a <=( (not A168)  and  (not A169) );
 a56205a <=( A170  and  a56204a );
 a56209a <=( A199  and  A166 );
 a56210a <=( (not A167)  and  a56209a );
 a56211a <=( a56210a  and  a56205a );
 a56215a <=( A266  and  A265 );
 a56216a <=( A200  and  a56215a );
 a56219a <=( (not A299)  and  A298 );
 a56222a <=( A302  and  A300 );
 a56223a <=( a56222a  and  a56219a );
 a56224a <=( a56223a  and  a56216a );
 a56228a <=( (not A168)  and  (not A169) );
 a56229a <=( A170  and  a56228a );
 a56233a <=( A199  and  A166 );
 a56234a <=( (not A167)  and  a56233a );
 a56235a <=( a56234a  and  a56229a );
 a56239a <=( A266  and  A265 );
 a56240a <=( A200  and  a56239a );
 a56243a <=( A299  and  (not A298) );
 a56246a <=( A301  and  A300 );
 a56247a <=( a56246a  and  a56243a );
 a56248a <=( a56247a  and  a56240a );
 a56252a <=( (not A168)  and  (not A169) );
 a56253a <=( A170  and  a56252a );
 a56257a <=( A199  and  A166 );
 a56258a <=( (not A167)  and  a56257a );
 a56259a <=( a56258a  and  a56253a );
 a56263a <=( A266  and  A265 );
 a56264a <=( A200  and  a56263a );
 a56267a <=( A299  and  (not A298) );
 a56270a <=( A302  and  A300 );
 a56271a <=( a56270a  and  a56267a );
 a56272a <=( a56271a  and  a56264a );
 a56276a <=( (not A168)  and  (not A169) );
 a56277a <=( A170  and  a56276a );
 a56281a <=( A199  and  A166 );
 a56282a <=( (not A167)  and  a56281a );
 a56283a <=( a56282a  and  a56277a );
 a56287a <=( (not A266)  and  (not A265) );
 a56288a <=( A200  and  a56287a );
 a56291a <=( (not A299)  and  A298 );
 a56294a <=( A301  and  A300 );
 a56295a <=( a56294a  and  a56291a );
 a56296a <=( a56295a  and  a56288a );
 a56300a <=( (not A168)  and  (not A169) );
 a56301a <=( A170  and  a56300a );
 a56305a <=( A199  and  A166 );
 a56306a <=( (not A167)  and  a56305a );
 a56307a <=( a56306a  and  a56301a );
 a56311a <=( (not A266)  and  (not A265) );
 a56312a <=( A200  and  a56311a );
 a56315a <=( (not A299)  and  A298 );
 a56318a <=( A302  and  A300 );
 a56319a <=( a56318a  and  a56315a );
 a56320a <=( a56319a  and  a56312a );
 a56324a <=( (not A168)  and  (not A169) );
 a56325a <=( A170  and  a56324a );
 a56329a <=( A199  and  A166 );
 a56330a <=( (not A167)  and  a56329a );
 a56331a <=( a56330a  and  a56325a );
 a56335a <=( (not A266)  and  (not A265) );
 a56336a <=( A200  and  a56335a );
 a56339a <=( A299  and  (not A298) );
 a56342a <=( A301  and  A300 );
 a56343a <=( a56342a  and  a56339a );
 a56344a <=( a56343a  and  a56336a );
 a56348a <=( (not A168)  and  (not A169) );
 a56349a <=( A170  and  a56348a );
 a56353a <=( A199  and  A166 );
 a56354a <=( (not A167)  and  a56353a );
 a56355a <=( a56354a  and  a56349a );
 a56359a <=( (not A266)  and  (not A265) );
 a56360a <=( A200  and  a56359a );
 a56363a <=( A299  and  (not A298) );
 a56366a <=( A302  and  A300 );
 a56367a <=( a56366a  and  a56363a );
 a56368a <=( a56367a  and  a56360a );
 a56372a <=( (not A168)  and  (not A169) );
 a56373a <=( A170  and  a56372a );
 a56377a <=( (not A199)  and  A166 );
 a56378a <=( (not A167)  and  a56377a );
 a56379a <=( a56378a  and  a56373a );
 a56383a <=( A268  and  (not A267) );
 a56384a <=( (not A200)  and  a56383a );
 a56387a <=( (not A299)  and  A298 );
 a56390a <=( A301  and  A300 );
 a56391a <=( a56390a  and  a56387a );
 a56392a <=( a56391a  and  a56384a );
 a56396a <=( (not A168)  and  (not A169) );
 a56397a <=( A170  and  a56396a );
 a56401a <=( (not A199)  and  A166 );
 a56402a <=( (not A167)  and  a56401a );
 a56403a <=( a56402a  and  a56397a );
 a56407a <=( A268  and  (not A267) );
 a56408a <=( (not A200)  and  a56407a );
 a56411a <=( (not A299)  and  A298 );
 a56414a <=( A302  and  A300 );
 a56415a <=( a56414a  and  a56411a );
 a56416a <=( a56415a  and  a56408a );
 a56420a <=( (not A168)  and  (not A169) );
 a56421a <=( A170  and  a56420a );
 a56425a <=( (not A199)  and  A166 );
 a56426a <=( (not A167)  and  a56425a );
 a56427a <=( a56426a  and  a56421a );
 a56431a <=( A268  and  (not A267) );
 a56432a <=( (not A200)  and  a56431a );
 a56435a <=( A299  and  (not A298) );
 a56438a <=( A301  and  A300 );
 a56439a <=( a56438a  and  a56435a );
 a56440a <=( a56439a  and  a56432a );
 a56444a <=( (not A168)  and  (not A169) );
 a56445a <=( A170  and  a56444a );
 a56449a <=( (not A199)  and  A166 );
 a56450a <=( (not A167)  and  a56449a );
 a56451a <=( a56450a  and  a56445a );
 a56455a <=( A268  and  (not A267) );
 a56456a <=( (not A200)  and  a56455a );
 a56459a <=( A299  and  (not A298) );
 a56462a <=( A302  and  A300 );
 a56463a <=( a56462a  and  a56459a );
 a56464a <=( a56463a  and  a56456a );
 a56468a <=( (not A168)  and  (not A169) );
 a56469a <=( A170  and  a56468a );
 a56473a <=( (not A199)  and  A166 );
 a56474a <=( (not A167)  and  a56473a );
 a56475a <=( a56474a  and  a56469a );
 a56479a <=( A269  and  (not A267) );
 a56480a <=( (not A200)  and  a56479a );
 a56483a <=( (not A299)  and  A298 );
 a56486a <=( A301  and  A300 );
 a56487a <=( a56486a  and  a56483a );
 a56488a <=( a56487a  and  a56480a );
 a56492a <=( (not A168)  and  (not A169) );
 a56493a <=( A170  and  a56492a );
 a56497a <=( (not A199)  and  A166 );
 a56498a <=( (not A167)  and  a56497a );
 a56499a <=( a56498a  and  a56493a );
 a56503a <=( A269  and  (not A267) );
 a56504a <=( (not A200)  and  a56503a );
 a56507a <=( (not A299)  and  A298 );
 a56510a <=( A302  and  A300 );
 a56511a <=( a56510a  and  a56507a );
 a56512a <=( a56511a  and  a56504a );
 a56516a <=( (not A168)  and  (not A169) );
 a56517a <=( A170  and  a56516a );
 a56521a <=( (not A199)  and  A166 );
 a56522a <=( (not A167)  and  a56521a );
 a56523a <=( a56522a  and  a56517a );
 a56527a <=( A269  and  (not A267) );
 a56528a <=( (not A200)  and  a56527a );
 a56531a <=( A299  and  (not A298) );
 a56534a <=( A301  and  A300 );
 a56535a <=( a56534a  and  a56531a );
 a56536a <=( a56535a  and  a56528a );
 a56540a <=( (not A168)  and  (not A169) );
 a56541a <=( A170  and  a56540a );
 a56545a <=( (not A199)  and  A166 );
 a56546a <=( (not A167)  and  a56545a );
 a56547a <=( a56546a  and  a56541a );
 a56551a <=( A269  and  (not A267) );
 a56552a <=( (not A200)  and  a56551a );
 a56555a <=( A299  and  (not A298) );
 a56558a <=( A302  and  A300 );
 a56559a <=( a56558a  and  a56555a );
 a56560a <=( a56559a  and  a56552a );
 a56564a <=( (not A168)  and  (not A169) );
 a56565a <=( A170  and  a56564a );
 a56569a <=( (not A199)  and  A166 );
 a56570a <=( (not A167)  and  a56569a );
 a56571a <=( a56570a  and  a56565a );
 a56575a <=( A266  and  A265 );
 a56576a <=( (not A200)  and  a56575a );
 a56579a <=( (not A299)  and  A298 );
 a56582a <=( A301  and  A300 );
 a56583a <=( a56582a  and  a56579a );
 a56584a <=( a56583a  and  a56576a );
 a56588a <=( (not A168)  and  (not A169) );
 a56589a <=( A170  and  a56588a );
 a56593a <=( (not A199)  and  A166 );
 a56594a <=( (not A167)  and  a56593a );
 a56595a <=( a56594a  and  a56589a );
 a56599a <=( A266  and  A265 );
 a56600a <=( (not A200)  and  a56599a );
 a56603a <=( (not A299)  and  A298 );
 a56606a <=( A302  and  A300 );
 a56607a <=( a56606a  and  a56603a );
 a56608a <=( a56607a  and  a56600a );
 a56612a <=( (not A168)  and  (not A169) );
 a56613a <=( A170  and  a56612a );
 a56617a <=( (not A199)  and  A166 );
 a56618a <=( (not A167)  and  a56617a );
 a56619a <=( a56618a  and  a56613a );
 a56623a <=( A266  and  A265 );
 a56624a <=( (not A200)  and  a56623a );
 a56627a <=( A299  and  (not A298) );
 a56630a <=( A301  and  A300 );
 a56631a <=( a56630a  and  a56627a );
 a56632a <=( a56631a  and  a56624a );
 a56636a <=( (not A168)  and  (not A169) );
 a56637a <=( A170  and  a56636a );
 a56641a <=( (not A199)  and  A166 );
 a56642a <=( (not A167)  and  a56641a );
 a56643a <=( a56642a  and  a56637a );
 a56647a <=( A266  and  A265 );
 a56648a <=( (not A200)  and  a56647a );
 a56651a <=( A299  and  (not A298) );
 a56654a <=( A302  and  A300 );
 a56655a <=( a56654a  and  a56651a );
 a56656a <=( a56655a  and  a56648a );
 a56660a <=( (not A168)  and  (not A169) );
 a56661a <=( A170  and  a56660a );
 a56665a <=( (not A199)  and  A166 );
 a56666a <=( (not A167)  and  a56665a );
 a56667a <=( a56666a  and  a56661a );
 a56671a <=( (not A266)  and  (not A265) );
 a56672a <=( (not A200)  and  a56671a );
 a56675a <=( (not A299)  and  A298 );
 a56678a <=( A301  and  A300 );
 a56679a <=( a56678a  and  a56675a );
 a56680a <=( a56679a  and  a56672a );
 a56684a <=( (not A168)  and  (not A169) );
 a56685a <=( A170  and  a56684a );
 a56689a <=( (not A199)  and  A166 );
 a56690a <=( (not A167)  and  a56689a );
 a56691a <=( a56690a  and  a56685a );
 a56695a <=( (not A266)  and  (not A265) );
 a56696a <=( (not A200)  and  a56695a );
 a56699a <=( (not A299)  and  A298 );
 a56702a <=( A302  and  A300 );
 a56703a <=( a56702a  and  a56699a );
 a56704a <=( a56703a  and  a56696a );
 a56708a <=( (not A168)  and  (not A169) );
 a56709a <=( A170  and  a56708a );
 a56713a <=( (not A199)  and  A166 );
 a56714a <=( (not A167)  and  a56713a );
 a56715a <=( a56714a  and  a56709a );
 a56719a <=( (not A266)  and  (not A265) );
 a56720a <=( (not A200)  and  a56719a );
 a56723a <=( A299  and  (not A298) );
 a56726a <=( A301  and  A300 );
 a56727a <=( a56726a  and  a56723a );
 a56728a <=( a56727a  and  a56720a );
 a56732a <=( (not A168)  and  (not A169) );
 a56733a <=( A170  and  a56732a );
 a56737a <=( (not A199)  and  A166 );
 a56738a <=( (not A167)  and  a56737a );
 a56739a <=( a56738a  and  a56733a );
 a56743a <=( (not A266)  and  (not A265) );
 a56744a <=( (not A200)  and  a56743a );
 a56747a <=( A299  and  (not A298) );
 a56750a <=( A302  and  A300 );
 a56751a <=( a56750a  and  a56747a );
 a56752a <=( a56751a  and  a56744a );
 a56756a <=( (not A199)  and  A166 );
 a56757a <=( A167  and  a56756a );
 a56760a <=( A201  and  A200 );
 a56763a <=( A267  and  A202 );
 a56764a <=( a56763a  and  a56760a );
 a56765a <=( a56764a  and  a56757a );
 a56769a <=( A298  and  (not A269) );
 a56770a <=( (not A268)  and  a56769a );
 a56773a <=( (not A300)  and  (not A299) );
 a56776a <=( (not A302)  and  (not A301) );
 a56777a <=( a56776a  and  a56773a );
 a56778a <=( a56777a  and  a56770a );
 a56782a <=( (not A199)  and  A166 );
 a56783a <=( A167  and  a56782a );
 a56786a <=( A201  and  A200 );
 a56789a <=( A267  and  A202 );
 a56790a <=( a56789a  and  a56786a );
 a56791a <=( a56790a  and  a56783a );
 a56795a <=( (not A298)  and  (not A269) );
 a56796a <=( (not A268)  and  a56795a );
 a56799a <=( (not A300)  and  A299 );
 a56802a <=( (not A302)  and  (not A301) );
 a56803a <=( a56802a  and  a56799a );
 a56804a <=( a56803a  and  a56796a );
 a56808a <=( (not A199)  and  A166 );
 a56809a <=( A167  and  a56808a );
 a56812a <=( A201  and  A200 );
 a56815a <=( A267  and  A203 );
 a56816a <=( a56815a  and  a56812a );
 a56817a <=( a56816a  and  a56809a );
 a56821a <=( A298  and  (not A269) );
 a56822a <=( (not A268)  and  a56821a );
 a56825a <=( (not A300)  and  (not A299) );
 a56828a <=( (not A302)  and  (not A301) );
 a56829a <=( a56828a  and  a56825a );
 a56830a <=( a56829a  and  a56822a );
 a56834a <=( (not A199)  and  A166 );
 a56835a <=( A167  and  a56834a );
 a56838a <=( A201  and  A200 );
 a56841a <=( A267  and  A203 );
 a56842a <=( a56841a  and  a56838a );
 a56843a <=( a56842a  and  a56835a );
 a56847a <=( (not A298)  and  (not A269) );
 a56848a <=( (not A268)  and  a56847a );
 a56851a <=( (not A300)  and  A299 );
 a56854a <=( (not A302)  and  (not A301) );
 a56855a <=( a56854a  and  a56851a );
 a56856a <=( a56855a  and  a56848a );
 a56860a <=( (not A199)  and  A166 );
 a56861a <=( A167  and  a56860a );
 a56864a <=( (not A201)  and  A200 );
 a56867a <=( (not A203)  and  (not A202) );
 a56868a <=( a56867a  and  a56864a );
 a56869a <=( a56868a  and  a56861a );
 a56873a <=( (not A269)  and  (not A268) );
 a56874a <=( A267  and  a56873a );
 a56877a <=( (not A299)  and  A298 );
 a56880a <=( A301  and  A300 );
 a56881a <=( a56880a  and  a56877a );
 a56882a <=( a56881a  and  a56874a );
 a56886a <=( (not A199)  and  A166 );
 a56887a <=( A167  and  a56886a );
 a56890a <=( (not A201)  and  A200 );
 a56893a <=( (not A203)  and  (not A202) );
 a56894a <=( a56893a  and  a56890a );
 a56895a <=( a56894a  and  a56887a );
 a56899a <=( (not A269)  and  (not A268) );
 a56900a <=( A267  and  a56899a );
 a56903a <=( (not A299)  and  A298 );
 a56906a <=( A302  and  A300 );
 a56907a <=( a56906a  and  a56903a );
 a56908a <=( a56907a  and  a56900a );
 a56912a <=( (not A199)  and  A166 );
 a56913a <=( A167  and  a56912a );
 a56916a <=( (not A201)  and  A200 );
 a56919a <=( (not A203)  and  (not A202) );
 a56920a <=( a56919a  and  a56916a );
 a56921a <=( a56920a  and  a56913a );
 a56925a <=( (not A269)  and  (not A268) );
 a56926a <=( A267  and  a56925a );
 a56929a <=( A299  and  (not A298) );
 a56932a <=( A301  and  A300 );
 a56933a <=( a56932a  and  a56929a );
 a56934a <=( a56933a  and  a56926a );
 a56938a <=( (not A199)  and  A166 );
 a56939a <=( A167  and  a56938a );
 a56942a <=( (not A201)  and  A200 );
 a56945a <=( (not A203)  and  (not A202) );
 a56946a <=( a56945a  and  a56942a );
 a56947a <=( a56946a  and  a56939a );
 a56951a <=( (not A269)  and  (not A268) );
 a56952a <=( A267  and  a56951a );
 a56955a <=( A299  and  (not A298) );
 a56958a <=( A302  and  A300 );
 a56959a <=( a56958a  and  a56955a );
 a56960a <=( a56959a  and  a56952a );
 a56964a <=( (not A199)  and  A166 );
 a56965a <=( A167  and  a56964a );
 a56968a <=( (not A201)  and  A200 );
 a56971a <=( (not A203)  and  (not A202) );
 a56972a <=( a56971a  and  a56968a );
 a56973a <=( a56972a  and  a56965a );
 a56977a <=( A298  and  A268 );
 a56978a <=( (not A267)  and  a56977a );
 a56981a <=( (not A300)  and  (not A299) );
 a56984a <=( (not A302)  and  (not A301) );
 a56985a <=( a56984a  and  a56981a );
 a56986a <=( a56985a  and  a56978a );
 a56990a <=( (not A199)  and  A166 );
 a56991a <=( A167  and  a56990a );
 a56994a <=( (not A201)  and  A200 );
 a56997a <=( (not A203)  and  (not A202) );
 a56998a <=( a56997a  and  a56994a );
 a56999a <=( a56998a  and  a56991a );
 a57003a <=( (not A298)  and  A268 );
 a57004a <=( (not A267)  and  a57003a );
 a57007a <=( (not A300)  and  A299 );
 a57010a <=( (not A302)  and  (not A301) );
 a57011a <=( a57010a  and  a57007a );
 a57012a <=( a57011a  and  a57004a );
 a57016a <=( (not A199)  and  A166 );
 a57017a <=( A167  and  a57016a );
 a57020a <=( (not A201)  and  A200 );
 a57023a <=( (not A203)  and  (not A202) );
 a57024a <=( a57023a  and  a57020a );
 a57025a <=( a57024a  and  a57017a );
 a57029a <=( A298  and  A269 );
 a57030a <=( (not A267)  and  a57029a );
 a57033a <=( (not A300)  and  (not A299) );
 a57036a <=( (not A302)  and  (not A301) );
 a57037a <=( a57036a  and  a57033a );
 a57038a <=( a57037a  and  a57030a );
 a57042a <=( (not A199)  and  A166 );
 a57043a <=( A167  and  a57042a );
 a57046a <=( (not A201)  and  A200 );
 a57049a <=( (not A203)  and  (not A202) );
 a57050a <=( a57049a  and  a57046a );
 a57051a <=( a57050a  and  a57043a );
 a57055a <=( (not A298)  and  A269 );
 a57056a <=( (not A267)  and  a57055a );
 a57059a <=( (not A300)  and  A299 );
 a57062a <=( (not A302)  and  (not A301) );
 a57063a <=( a57062a  and  a57059a );
 a57064a <=( a57063a  and  a57056a );
 a57068a <=( (not A199)  and  A166 );
 a57069a <=( A167  and  a57068a );
 a57072a <=( (not A201)  and  A200 );
 a57075a <=( (not A203)  and  (not A202) );
 a57076a <=( a57075a  and  a57072a );
 a57077a <=( a57076a  and  a57069a );
 a57081a <=( A298  and  A266 );
 a57082a <=( A265  and  a57081a );
 a57085a <=( (not A300)  and  (not A299) );
 a57088a <=( (not A302)  and  (not A301) );
 a57089a <=( a57088a  and  a57085a );
 a57090a <=( a57089a  and  a57082a );
 a57094a <=( (not A199)  and  A166 );
 a57095a <=( A167  and  a57094a );
 a57098a <=( (not A201)  and  A200 );
 a57101a <=( (not A203)  and  (not A202) );
 a57102a <=( a57101a  and  a57098a );
 a57103a <=( a57102a  and  a57095a );
 a57107a <=( (not A298)  and  A266 );
 a57108a <=( A265  and  a57107a );
 a57111a <=( (not A300)  and  A299 );
 a57114a <=( (not A302)  and  (not A301) );
 a57115a <=( a57114a  and  a57111a );
 a57116a <=( a57115a  and  a57108a );
 a57120a <=( (not A199)  and  A166 );
 a57121a <=( A167  and  a57120a );
 a57124a <=( (not A201)  and  A200 );
 a57127a <=( (not A203)  and  (not A202) );
 a57128a <=( a57127a  and  a57124a );
 a57129a <=( a57128a  and  a57121a );
 a57133a <=( A298  and  (not A266) );
 a57134a <=( (not A265)  and  a57133a );
 a57137a <=( (not A300)  and  (not A299) );
 a57140a <=( (not A302)  and  (not A301) );
 a57141a <=( a57140a  and  a57137a );
 a57142a <=( a57141a  and  a57134a );
 a57146a <=( (not A199)  and  A166 );
 a57147a <=( A167  and  a57146a );
 a57150a <=( (not A201)  and  A200 );
 a57153a <=( (not A203)  and  (not A202) );
 a57154a <=( a57153a  and  a57150a );
 a57155a <=( a57154a  and  a57147a );
 a57159a <=( (not A298)  and  (not A266) );
 a57160a <=( (not A265)  and  a57159a );
 a57163a <=( (not A300)  and  A299 );
 a57166a <=( (not A302)  and  (not A301) );
 a57167a <=( a57166a  and  a57163a );
 a57168a <=( a57167a  and  a57160a );
 a57172a <=( A199  and  A166 );
 a57173a <=( A167  and  a57172a );
 a57176a <=( A201  and  (not A200) );
 a57179a <=( A267  and  A202 );
 a57180a <=( a57179a  and  a57176a );
 a57181a <=( a57180a  and  a57173a );
 a57185a <=( A298  and  (not A269) );
 a57186a <=( (not A268)  and  a57185a );
 a57189a <=( (not A300)  and  (not A299) );
 a57192a <=( (not A302)  and  (not A301) );
 a57193a <=( a57192a  and  a57189a );
 a57194a <=( a57193a  and  a57186a );
 a57198a <=( A199  and  A166 );
 a57199a <=( A167  and  a57198a );
 a57202a <=( A201  and  (not A200) );
 a57205a <=( A267  and  A202 );
 a57206a <=( a57205a  and  a57202a );
 a57207a <=( a57206a  and  a57199a );
 a57211a <=( (not A298)  and  (not A269) );
 a57212a <=( (not A268)  and  a57211a );
 a57215a <=( (not A300)  and  A299 );
 a57218a <=( (not A302)  and  (not A301) );
 a57219a <=( a57218a  and  a57215a );
 a57220a <=( a57219a  and  a57212a );
 a57224a <=( A199  and  A166 );
 a57225a <=( A167  and  a57224a );
 a57228a <=( A201  and  (not A200) );
 a57231a <=( A267  and  A203 );
 a57232a <=( a57231a  and  a57228a );
 a57233a <=( a57232a  and  a57225a );
 a57237a <=( A298  and  (not A269) );
 a57238a <=( (not A268)  and  a57237a );
 a57241a <=( (not A300)  and  (not A299) );
 a57244a <=( (not A302)  and  (not A301) );
 a57245a <=( a57244a  and  a57241a );
 a57246a <=( a57245a  and  a57238a );
 a57250a <=( A199  and  A166 );
 a57251a <=( A167  and  a57250a );
 a57254a <=( A201  and  (not A200) );
 a57257a <=( A267  and  A203 );
 a57258a <=( a57257a  and  a57254a );
 a57259a <=( a57258a  and  a57251a );
 a57263a <=( (not A298)  and  (not A269) );
 a57264a <=( (not A268)  and  a57263a );
 a57267a <=( (not A300)  and  A299 );
 a57270a <=( (not A302)  and  (not A301) );
 a57271a <=( a57270a  and  a57267a );
 a57272a <=( a57271a  and  a57264a );
 a57276a <=( A199  and  A166 );
 a57277a <=( A167  and  a57276a );
 a57280a <=( (not A201)  and  (not A200) );
 a57283a <=( (not A203)  and  (not A202) );
 a57284a <=( a57283a  and  a57280a );
 a57285a <=( a57284a  and  a57277a );
 a57289a <=( (not A269)  and  (not A268) );
 a57290a <=( A267  and  a57289a );
 a57293a <=( (not A299)  and  A298 );
 a57296a <=( A301  and  A300 );
 a57297a <=( a57296a  and  a57293a );
 a57298a <=( a57297a  and  a57290a );
 a57302a <=( A199  and  A166 );
 a57303a <=( A167  and  a57302a );
 a57306a <=( (not A201)  and  (not A200) );
 a57309a <=( (not A203)  and  (not A202) );
 a57310a <=( a57309a  and  a57306a );
 a57311a <=( a57310a  and  a57303a );
 a57315a <=( (not A269)  and  (not A268) );
 a57316a <=( A267  and  a57315a );
 a57319a <=( (not A299)  and  A298 );
 a57322a <=( A302  and  A300 );
 a57323a <=( a57322a  and  a57319a );
 a57324a <=( a57323a  and  a57316a );
 a57328a <=( A199  and  A166 );
 a57329a <=( A167  and  a57328a );
 a57332a <=( (not A201)  and  (not A200) );
 a57335a <=( (not A203)  and  (not A202) );
 a57336a <=( a57335a  and  a57332a );
 a57337a <=( a57336a  and  a57329a );
 a57341a <=( (not A269)  and  (not A268) );
 a57342a <=( A267  and  a57341a );
 a57345a <=( A299  and  (not A298) );
 a57348a <=( A301  and  A300 );
 a57349a <=( a57348a  and  a57345a );
 a57350a <=( a57349a  and  a57342a );
 a57354a <=( A199  and  A166 );
 a57355a <=( A167  and  a57354a );
 a57358a <=( (not A201)  and  (not A200) );
 a57361a <=( (not A203)  and  (not A202) );
 a57362a <=( a57361a  and  a57358a );
 a57363a <=( a57362a  and  a57355a );
 a57367a <=( (not A269)  and  (not A268) );
 a57368a <=( A267  and  a57367a );
 a57371a <=( A299  and  (not A298) );
 a57374a <=( A302  and  A300 );
 a57375a <=( a57374a  and  a57371a );
 a57376a <=( a57375a  and  a57368a );
 a57380a <=( A199  and  A166 );
 a57381a <=( A167  and  a57380a );
 a57384a <=( (not A201)  and  (not A200) );
 a57387a <=( (not A203)  and  (not A202) );
 a57388a <=( a57387a  and  a57384a );
 a57389a <=( a57388a  and  a57381a );
 a57393a <=( A298  and  A268 );
 a57394a <=( (not A267)  and  a57393a );
 a57397a <=( (not A300)  and  (not A299) );
 a57400a <=( (not A302)  and  (not A301) );
 a57401a <=( a57400a  and  a57397a );
 a57402a <=( a57401a  and  a57394a );
 a57406a <=( A199  and  A166 );
 a57407a <=( A167  and  a57406a );
 a57410a <=( (not A201)  and  (not A200) );
 a57413a <=( (not A203)  and  (not A202) );
 a57414a <=( a57413a  and  a57410a );
 a57415a <=( a57414a  and  a57407a );
 a57419a <=( (not A298)  and  A268 );
 a57420a <=( (not A267)  and  a57419a );
 a57423a <=( (not A300)  and  A299 );
 a57426a <=( (not A302)  and  (not A301) );
 a57427a <=( a57426a  and  a57423a );
 a57428a <=( a57427a  and  a57420a );
 a57432a <=( A199  and  A166 );
 a57433a <=( A167  and  a57432a );
 a57436a <=( (not A201)  and  (not A200) );
 a57439a <=( (not A203)  and  (not A202) );
 a57440a <=( a57439a  and  a57436a );
 a57441a <=( a57440a  and  a57433a );
 a57445a <=( A298  and  A269 );
 a57446a <=( (not A267)  and  a57445a );
 a57449a <=( (not A300)  and  (not A299) );
 a57452a <=( (not A302)  and  (not A301) );
 a57453a <=( a57452a  and  a57449a );
 a57454a <=( a57453a  and  a57446a );
 a57458a <=( A199  and  A166 );
 a57459a <=( A167  and  a57458a );
 a57462a <=( (not A201)  and  (not A200) );
 a57465a <=( (not A203)  and  (not A202) );
 a57466a <=( a57465a  and  a57462a );
 a57467a <=( a57466a  and  a57459a );
 a57471a <=( (not A298)  and  A269 );
 a57472a <=( (not A267)  and  a57471a );
 a57475a <=( (not A300)  and  A299 );
 a57478a <=( (not A302)  and  (not A301) );
 a57479a <=( a57478a  and  a57475a );
 a57480a <=( a57479a  and  a57472a );
 a57484a <=( A199  and  A166 );
 a57485a <=( A167  and  a57484a );
 a57488a <=( (not A201)  and  (not A200) );
 a57491a <=( (not A203)  and  (not A202) );
 a57492a <=( a57491a  and  a57488a );
 a57493a <=( a57492a  and  a57485a );
 a57497a <=( A298  and  A266 );
 a57498a <=( A265  and  a57497a );
 a57501a <=( (not A300)  and  (not A299) );
 a57504a <=( (not A302)  and  (not A301) );
 a57505a <=( a57504a  and  a57501a );
 a57506a <=( a57505a  and  a57498a );
 a57510a <=( A199  and  A166 );
 a57511a <=( A167  and  a57510a );
 a57514a <=( (not A201)  and  (not A200) );
 a57517a <=( (not A203)  and  (not A202) );
 a57518a <=( a57517a  and  a57514a );
 a57519a <=( a57518a  and  a57511a );
 a57523a <=( (not A298)  and  A266 );
 a57524a <=( A265  and  a57523a );
 a57527a <=( (not A300)  and  A299 );
 a57530a <=( (not A302)  and  (not A301) );
 a57531a <=( a57530a  and  a57527a );
 a57532a <=( a57531a  and  a57524a );
 a57536a <=( A199  and  A166 );
 a57537a <=( A167  and  a57536a );
 a57540a <=( (not A201)  and  (not A200) );
 a57543a <=( (not A203)  and  (not A202) );
 a57544a <=( a57543a  and  a57540a );
 a57545a <=( a57544a  and  a57537a );
 a57549a <=( A298  and  (not A266) );
 a57550a <=( (not A265)  and  a57549a );
 a57553a <=( (not A300)  and  (not A299) );
 a57556a <=( (not A302)  and  (not A301) );
 a57557a <=( a57556a  and  a57553a );
 a57558a <=( a57557a  and  a57550a );
 a57562a <=( A199  and  A166 );
 a57563a <=( A167  and  a57562a );
 a57566a <=( (not A201)  and  (not A200) );
 a57569a <=( (not A203)  and  (not A202) );
 a57570a <=( a57569a  and  a57566a );
 a57571a <=( a57570a  and  a57563a );
 a57575a <=( (not A298)  and  (not A266) );
 a57576a <=( (not A265)  and  a57575a );
 a57579a <=( (not A300)  and  A299 );
 a57582a <=( (not A302)  and  (not A301) );
 a57583a <=( a57582a  and  a57579a );
 a57584a <=( a57583a  and  a57576a );
 a57588a <=( (not A199)  and  (not A166) );
 a57589a <=( (not A167)  and  a57588a );
 a57592a <=( A201  and  A200 );
 a57595a <=( A267  and  A202 );
 a57596a <=( a57595a  and  a57592a );
 a57597a <=( a57596a  and  a57589a );
 a57601a <=( A298  and  (not A269) );
 a57602a <=( (not A268)  and  a57601a );
 a57605a <=( (not A300)  and  (not A299) );
 a57608a <=( (not A302)  and  (not A301) );
 a57609a <=( a57608a  and  a57605a );
 a57610a <=( a57609a  and  a57602a );
 a57614a <=( (not A199)  and  (not A166) );
 a57615a <=( (not A167)  and  a57614a );
 a57618a <=( A201  and  A200 );
 a57621a <=( A267  and  A202 );
 a57622a <=( a57621a  and  a57618a );
 a57623a <=( a57622a  and  a57615a );
 a57627a <=( (not A298)  and  (not A269) );
 a57628a <=( (not A268)  and  a57627a );
 a57631a <=( (not A300)  and  A299 );
 a57634a <=( (not A302)  and  (not A301) );
 a57635a <=( a57634a  and  a57631a );
 a57636a <=( a57635a  and  a57628a );
 a57640a <=( (not A199)  and  (not A166) );
 a57641a <=( (not A167)  and  a57640a );
 a57644a <=( A201  and  A200 );
 a57647a <=( A267  and  A203 );
 a57648a <=( a57647a  and  a57644a );
 a57649a <=( a57648a  and  a57641a );
 a57653a <=( A298  and  (not A269) );
 a57654a <=( (not A268)  and  a57653a );
 a57657a <=( (not A300)  and  (not A299) );
 a57660a <=( (not A302)  and  (not A301) );
 a57661a <=( a57660a  and  a57657a );
 a57662a <=( a57661a  and  a57654a );
 a57666a <=( (not A199)  and  (not A166) );
 a57667a <=( (not A167)  and  a57666a );
 a57670a <=( A201  and  A200 );
 a57673a <=( A267  and  A203 );
 a57674a <=( a57673a  and  a57670a );
 a57675a <=( a57674a  and  a57667a );
 a57679a <=( (not A298)  and  (not A269) );
 a57680a <=( (not A268)  and  a57679a );
 a57683a <=( (not A300)  and  A299 );
 a57686a <=( (not A302)  and  (not A301) );
 a57687a <=( a57686a  and  a57683a );
 a57688a <=( a57687a  and  a57680a );
 a57692a <=( (not A199)  and  (not A166) );
 a57693a <=( (not A167)  and  a57692a );
 a57696a <=( (not A201)  and  A200 );
 a57699a <=( (not A203)  and  (not A202) );
 a57700a <=( a57699a  and  a57696a );
 a57701a <=( a57700a  and  a57693a );
 a57705a <=( (not A269)  and  (not A268) );
 a57706a <=( A267  and  a57705a );
 a57709a <=( (not A299)  and  A298 );
 a57712a <=( A301  and  A300 );
 a57713a <=( a57712a  and  a57709a );
 a57714a <=( a57713a  and  a57706a );
 a57718a <=( (not A199)  and  (not A166) );
 a57719a <=( (not A167)  and  a57718a );
 a57722a <=( (not A201)  and  A200 );
 a57725a <=( (not A203)  and  (not A202) );
 a57726a <=( a57725a  and  a57722a );
 a57727a <=( a57726a  and  a57719a );
 a57731a <=( (not A269)  and  (not A268) );
 a57732a <=( A267  and  a57731a );
 a57735a <=( (not A299)  and  A298 );
 a57738a <=( A302  and  A300 );
 a57739a <=( a57738a  and  a57735a );
 a57740a <=( a57739a  and  a57732a );
 a57744a <=( (not A199)  and  (not A166) );
 a57745a <=( (not A167)  and  a57744a );
 a57748a <=( (not A201)  and  A200 );
 a57751a <=( (not A203)  and  (not A202) );
 a57752a <=( a57751a  and  a57748a );
 a57753a <=( a57752a  and  a57745a );
 a57757a <=( (not A269)  and  (not A268) );
 a57758a <=( A267  and  a57757a );
 a57761a <=( A299  and  (not A298) );
 a57764a <=( A301  and  A300 );
 a57765a <=( a57764a  and  a57761a );
 a57766a <=( a57765a  and  a57758a );
 a57770a <=( (not A199)  and  (not A166) );
 a57771a <=( (not A167)  and  a57770a );
 a57774a <=( (not A201)  and  A200 );
 a57777a <=( (not A203)  and  (not A202) );
 a57778a <=( a57777a  and  a57774a );
 a57779a <=( a57778a  and  a57771a );
 a57783a <=( (not A269)  and  (not A268) );
 a57784a <=( A267  and  a57783a );
 a57787a <=( A299  and  (not A298) );
 a57790a <=( A302  and  A300 );
 a57791a <=( a57790a  and  a57787a );
 a57792a <=( a57791a  and  a57784a );
 a57796a <=( (not A199)  and  (not A166) );
 a57797a <=( (not A167)  and  a57796a );
 a57800a <=( (not A201)  and  A200 );
 a57803a <=( (not A203)  and  (not A202) );
 a57804a <=( a57803a  and  a57800a );
 a57805a <=( a57804a  and  a57797a );
 a57809a <=( A298  and  A268 );
 a57810a <=( (not A267)  and  a57809a );
 a57813a <=( (not A300)  and  (not A299) );
 a57816a <=( (not A302)  and  (not A301) );
 a57817a <=( a57816a  and  a57813a );
 a57818a <=( a57817a  and  a57810a );
 a57822a <=( (not A199)  and  (not A166) );
 a57823a <=( (not A167)  and  a57822a );
 a57826a <=( (not A201)  and  A200 );
 a57829a <=( (not A203)  and  (not A202) );
 a57830a <=( a57829a  and  a57826a );
 a57831a <=( a57830a  and  a57823a );
 a57835a <=( (not A298)  and  A268 );
 a57836a <=( (not A267)  and  a57835a );
 a57839a <=( (not A300)  and  A299 );
 a57842a <=( (not A302)  and  (not A301) );
 a57843a <=( a57842a  and  a57839a );
 a57844a <=( a57843a  and  a57836a );
 a57848a <=( (not A199)  and  (not A166) );
 a57849a <=( (not A167)  and  a57848a );
 a57852a <=( (not A201)  and  A200 );
 a57855a <=( (not A203)  and  (not A202) );
 a57856a <=( a57855a  and  a57852a );
 a57857a <=( a57856a  and  a57849a );
 a57861a <=( A298  and  A269 );
 a57862a <=( (not A267)  and  a57861a );
 a57865a <=( (not A300)  and  (not A299) );
 a57868a <=( (not A302)  and  (not A301) );
 a57869a <=( a57868a  and  a57865a );
 a57870a <=( a57869a  and  a57862a );
 a57874a <=( (not A199)  and  (not A166) );
 a57875a <=( (not A167)  and  a57874a );
 a57878a <=( (not A201)  and  A200 );
 a57881a <=( (not A203)  and  (not A202) );
 a57882a <=( a57881a  and  a57878a );
 a57883a <=( a57882a  and  a57875a );
 a57887a <=( (not A298)  and  A269 );
 a57888a <=( (not A267)  and  a57887a );
 a57891a <=( (not A300)  and  A299 );
 a57894a <=( (not A302)  and  (not A301) );
 a57895a <=( a57894a  and  a57891a );
 a57896a <=( a57895a  and  a57888a );
 a57900a <=( (not A199)  and  (not A166) );
 a57901a <=( (not A167)  and  a57900a );
 a57904a <=( (not A201)  and  A200 );
 a57907a <=( (not A203)  and  (not A202) );
 a57908a <=( a57907a  and  a57904a );
 a57909a <=( a57908a  and  a57901a );
 a57913a <=( A298  and  A266 );
 a57914a <=( A265  and  a57913a );
 a57917a <=( (not A300)  and  (not A299) );
 a57920a <=( (not A302)  and  (not A301) );
 a57921a <=( a57920a  and  a57917a );
 a57922a <=( a57921a  and  a57914a );
 a57926a <=( (not A199)  and  (not A166) );
 a57927a <=( (not A167)  and  a57926a );
 a57930a <=( (not A201)  and  A200 );
 a57933a <=( (not A203)  and  (not A202) );
 a57934a <=( a57933a  and  a57930a );
 a57935a <=( a57934a  and  a57927a );
 a57939a <=( (not A298)  and  A266 );
 a57940a <=( A265  and  a57939a );
 a57943a <=( (not A300)  and  A299 );
 a57946a <=( (not A302)  and  (not A301) );
 a57947a <=( a57946a  and  a57943a );
 a57948a <=( a57947a  and  a57940a );
 a57952a <=( (not A199)  and  (not A166) );
 a57953a <=( (not A167)  and  a57952a );
 a57956a <=( (not A201)  and  A200 );
 a57959a <=( (not A203)  and  (not A202) );
 a57960a <=( a57959a  and  a57956a );
 a57961a <=( a57960a  and  a57953a );
 a57965a <=( A298  and  (not A266) );
 a57966a <=( (not A265)  and  a57965a );
 a57969a <=( (not A300)  and  (not A299) );
 a57972a <=( (not A302)  and  (not A301) );
 a57973a <=( a57972a  and  a57969a );
 a57974a <=( a57973a  and  a57966a );
 a57978a <=( (not A199)  and  (not A166) );
 a57979a <=( (not A167)  and  a57978a );
 a57982a <=( (not A201)  and  A200 );
 a57985a <=( (not A203)  and  (not A202) );
 a57986a <=( a57985a  and  a57982a );
 a57987a <=( a57986a  and  a57979a );
 a57991a <=( (not A298)  and  (not A266) );
 a57992a <=( (not A265)  and  a57991a );
 a57995a <=( (not A300)  and  A299 );
 a57998a <=( (not A302)  and  (not A301) );
 a57999a <=( a57998a  and  a57995a );
 a58000a <=( a57999a  and  a57992a );
 a58004a <=( A199  and  (not A166) );
 a58005a <=( (not A167)  and  a58004a );
 a58008a <=( A201  and  (not A200) );
 a58011a <=( A267  and  A202 );
 a58012a <=( a58011a  and  a58008a );
 a58013a <=( a58012a  and  a58005a );
 a58017a <=( A298  and  (not A269) );
 a58018a <=( (not A268)  and  a58017a );
 a58021a <=( (not A300)  and  (not A299) );
 a58024a <=( (not A302)  and  (not A301) );
 a58025a <=( a58024a  and  a58021a );
 a58026a <=( a58025a  and  a58018a );
 a58030a <=( A199  and  (not A166) );
 a58031a <=( (not A167)  and  a58030a );
 a58034a <=( A201  and  (not A200) );
 a58037a <=( A267  and  A202 );
 a58038a <=( a58037a  and  a58034a );
 a58039a <=( a58038a  and  a58031a );
 a58043a <=( (not A298)  and  (not A269) );
 a58044a <=( (not A268)  and  a58043a );
 a58047a <=( (not A300)  and  A299 );
 a58050a <=( (not A302)  and  (not A301) );
 a58051a <=( a58050a  and  a58047a );
 a58052a <=( a58051a  and  a58044a );
 a58056a <=( A199  and  (not A166) );
 a58057a <=( (not A167)  and  a58056a );
 a58060a <=( A201  and  (not A200) );
 a58063a <=( A267  and  A203 );
 a58064a <=( a58063a  and  a58060a );
 a58065a <=( a58064a  and  a58057a );
 a58069a <=( A298  and  (not A269) );
 a58070a <=( (not A268)  and  a58069a );
 a58073a <=( (not A300)  and  (not A299) );
 a58076a <=( (not A302)  and  (not A301) );
 a58077a <=( a58076a  and  a58073a );
 a58078a <=( a58077a  and  a58070a );
 a58082a <=( A199  and  (not A166) );
 a58083a <=( (not A167)  and  a58082a );
 a58086a <=( A201  and  (not A200) );
 a58089a <=( A267  and  A203 );
 a58090a <=( a58089a  and  a58086a );
 a58091a <=( a58090a  and  a58083a );
 a58095a <=( (not A298)  and  (not A269) );
 a58096a <=( (not A268)  and  a58095a );
 a58099a <=( (not A300)  and  A299 );
 a58102a <=( (not A302)  and  (not A301) );
 a58103a <=( a58102a  and  a58099a );
 a58104a <=( a58103a  and  a58096a );
 a58108a <=( A199  and  (not A166) );
 a58109a <=( (not A167)  and  a58108a );
 a58112a <=( (not A201)  and  (not A200) );
 a58115a <=( (not A203)  and  (not A202) );
 a58116a <=( a58115a  and  a58112a );
 a58117a <=( a58116a  and  a58109a );
 a58121a <=( (not A269)  and  (not A268) );
 a58122a <=( A267  and  a58121a );
 a58125a <=( (not A299)  and  A298 );
 a58128a <=( A301  and  A300 );
 a58129a <=( a58128a  and  a58125a );
 a58130a <=( a58129a  and  a58122a );
 a58134a <=( A199  and  (not A166) );
 a58135a <=( (not A167)  and  a58134a );
 a58138a <=( (not A201)  and  (not A200) );
 a58141a <=( (not A203)  and  (not A202) );
 a58142a <=( a58141a  and  a58138a );
 a58143a <=( a58142a  and  a58135a );
 a58147a <=( (not A269)  and  (not A268) );
 a58148a <=( A267  and  a58147a );
 a58151a <=( (not A299)  and  A298 );
 a58154a <=( A302  and  A300 );
 a58155a <=( a58154a  and  a58151a );
 a58156a <=( a58155a  and  a58148a );
 a58160a <=( A199  and  (not A166) );
 a58161a <=( (not A167)  and  a58160a );
 a58164a <=( (not A201)  and  (not A200) );
 a58167a <=( (not A203)  and  (not A202) );
 a58168a <=( a58167a  and  a58164a );
 a58169a <=( a58168a  and  a58161a );
 a58173a <=( (not A269)  and  (not A268) );
 a58174a <=( A267  and  a58173a );
 a58177a <=( A299  and  (not A298) );
 a58180a <=( A301  and  A300 );
 a58181a <=( a58180a  and  a58177a );
 a58182a <=( a58181a  and  a58174a );
 a58186a <=( A199  and  (not A166) );
 a58187a <=( (not A167)  and  a58186a );
 a58190a <=( (not A201)  and  (not A200) );
 a58193a <=( (not A203)  and  (not A202) );
 a58194a <=( a58193a  and  a58190a );
 a58195a <=( a58194a  and  a58187a );
 a58199a <=( (not A269)  and  (not A268) );
 a58200a <=( A267  and  a58199a );
 a58203a <=( A299  and  (not A298) );
 a58206a <=( A302  and  A300 );
 a58207a <=( a58206a  and  a58203a );
 a58208a <=( a58207a  and  a58200a );
 a58212a <=( A199  and  (not A166) );
 a58213a <=( (not A167)  and  a58212a );
 a58216a <=( (not A201)  and  (not A200) );
 a58219a <=( (not A203)  and  (not A202) );
 a58220a <=( a58219a  and  a58216a );
 a58221a <=( a58220a  and  a58213a );
 a58225a <=( A298  and  A268 );
 a58226a <=( (not A267)  and  a58225a );
 a58229a <=( (not A300)  and  (not A299) );
 a58232a <=( (not A302)  and  (not A301) );
 a58233a <=( a58232a  and  a58229a );
 a58234a <=( a58233a  and  a58226a );
 a58238a <=( A199  and  (not A166) );
 a58239a <=( (not A167)  and  a58238a );
 a58242a <=( (not A201)  and  (not A200) );
 a58245a <=( (not A203)  and  (not A202) );
 a58246a <=( a58245a  and  a58242a );
 a58247a <=( a58246a  and  a58239a );
 a58251a <=( (not A298)  and  A268 );
 a58252a <=( (not A267)  and  a58251a );
 a58255a <=( (not A300)  and  A299 );
 a58258a <=( (not A302)  and  (not A301) );
 a58259a <=( a58258a  and  a58255a );
 a58260a <=( a58259a  and  a58252a );
 a58264a <=( A199  and  (not A166) );
 a58265a <=( (not A167)  and  a58264a );
 a58268a <=( (not A201)  and  (not A200) );
 a58271a <=( (not A203)  and  (not A202) );
 a58272a <=( a58271a  and  a58268a );
 a58273a <=( a58272a  and  a58265a );
 a58277a <=( A298  and  A269 );
 a58278a <=( (not A267)  and  a58277a );
 a58281a <=( (not A300)  and  (not A299) );
 a58284a <=( (not A302)  and  (not A301) );
 a58285a <=( a58284a  and  a58281a );
 a58286a <=( a58285a  and  a58278a );
 a58290a <=( A199  and  (not A166) );
 a58291a <=( (not A167)  and  a58290a );
 a58294a <=( (not A201)  and  (not A200) );
 a58297a <=( (not A203)  and  (not A202) );
 a58298a <=( a58297a  and  a58294a );
 a58299a <=( a58298a  and  a58291a );
 a58303a <=( (not A298)  and  A269 );
 a58304a <=( (not A267)  and  a58303a );
 a58307a <=( (not A300)  and  A299 );
 a58310a <=( (not A302)  and  (not A301) );
 a58311a <=( a58310a  and  a58307a );
 a58312a <=( a58311a  and  a58304a );
 a58316a <=( A199  and  (not A166) );
 a58317a <=( (not A167)  and  a58316a );
 a58320a <=( (not A201)  and  (not A200) );
 a58323a <=( (not A203)  and  (not A202) );
 a58324a <=( a58323a  and  a58320a );
 a58325a <=( a58324a  and  a58317a );
 a58329a <=( A298  and  A266 );
 a58330a <=( A265  and  a58329a );
 a58333a <=( (not A300)  and  (not A299) );
 a58336a <=( (not A302)  and  (not A301) );
 a58337a <=( a58336a  and  a58333a );
 a58338a <=( a58337a  and  a58330a );
 a58342a <=( A199  and  (not A166) );
 a58343a <=( (not A167)  and  a58342a );
 a58346a <=( (not A201)  and  (not A200) );
 a58349a <=( (not A203)  and  (not A202) );
 a58350a <=( a58349a  and  a58346a );
 a58351a <=( a58350a  and  a58343a );
 a58355a <=( (not A298)  and  A266 );
 a58356a <=( A265  and  a58355a );
 a58359a <=( (not A300)  and  A299 );
 a58362a <=( (not A302)  and  (not A301) );
 a58363a <=( a58362a  and  a58359a );
 a58364a <=( a58363a  and  a58356a );
 a58368a <=( A199  and  (not A166) );
 a58369a <=( (not A167)  and  a58368a );
 a58372a <=( (not A201)  and  (not A200) );
 a58375a <=( (not A203)  and  (not A202) );
 a58376a <=( a58375a  and  a58372a );
 a58377a <=( a58376a  and  a58369a );
 a58381a <=( A298  and  (not A266) );
 a58382a <=( (not A265)  and  a58381a );
 a58385a <=( (not A300)  and  (not A299) );
 a58388a <=( (not A302)  and  (not A301) );
 a58389a <=( a58388a  and  a58385a );
 a58390a <=( a58389a  and  a58382a );
 a58394a <=( A199  and  (not A166) );
 a58395a <=( (not A167)  and  a58394a );
 a58398a <=( (not A201)  and  (not A200) );
 a58401a <=( (not A203)  and  (not A202) );
 a58402a <=( a58401a  and  a58398a );
 a58403a <=( a58402a  and  a58395a );
 a58407a <=( (not A298)  and  (not A266) );
 a58408a <=( (not A265)  and  a58407a );
 a58411a <=( (not A300)  and  A299 );
 a58414a <=( (not A302)  and  (not A301) );
 a58415a <=( a58414a  and  a58411a );
 a58416a <=( a58415a  and  a58408a );
 a58420a <=( A167  and  A168 );
 a58421a <=( (not A170)  and  a58420a );
 a58424a <=( A201  and  (not A166) );
 a58427a <=( (not A203)  and  (not A202) );
 a58428a <=( a58427a  and  a58424a );
 a58429a <=( a58428a  and  a58421a );
 a58433a <=( (not A269)  and  (not A268) );
 a58434a <=( A267  and  a58433a );
 a58437a <=( (not A299)  and  A298 );
 a58440a <=( A301  and  A300 );
 a58441a <=( a58440a  and  a58437a );
 a58442a <=( a58441a  and  a58434a );
 a58446a <=( A167  and  A168 );
 a58447a <=( (not A170)  and  a58446a );
 a58450a <=( A201  and  (not A166) );
 a58453a <=( (not A203)  and  (not A202) );
 a58454a <=( a58453a  and  a58450a );
 a58455a <=( a58454a  and  a58447a );
 a58459a <=( (not A269)  and  (not A268) );
 a58460a <=( A267  and  a58459a );
 a58463a <=( (not A299)  and  A298 );
 a58466a <=( A302  and  A300 );
 a58467a <=( a58466a  and  a58463a );
 a58468a <=( a58467a  and  a58460a );
 a58472a <=( A167  and  A168 );
 a58473a <=( (not A170)  and  a58472a );
 a58476a <=( A201  and  (not A166) );
 a58479a <=( (not A203)  and  (not A202) );
 a58480a <=( a58479a  and  a58476a );
 a58481a <=( a58480a  and  a58473a );
 a58485a <=( (not A269)  and  (not A268) );
 a58486a <=( A267  and  a58485a );
 a58489a <=( A299  and  (not A298) );
 a58492a <=( A301  and  A300 );
 a58493a <=( a58492a  and  a58489a );
 a58494a <=( a58493a  and  a58486a );
 a58498a <=( A167  and  A168 );
 a58499a <=( (not A170)  and  a58498a );
 a58502a <=( A201  and  (not A166) );
 a58505a <=( (not A203)  and  (not A202) );
 a58506a <=( a58505a  and  a58502a );
 a58507a <=( a58506a  and  a58499a );
 a58511a <=( (not A269)  and  (not A268) );
 a58512a <=( A267  and  a58511a );
 a58515a <=( A299  and  (not A298) );
 a58518a <=( A302  and  A300 );
 a58519a <=( a58518a  and  a58515a );
 a58520a <=( a58519a  and  a58512a );
 a58524a <=( A167  and  A168 );
 a58525a <=( (not A170)  and  a58524a );
 a58528a <=( A201  and  (not A166) );
 a58531a <=( (not A203)  and  (not A202) );
 a58532a <=( a58531a  and  a58528a );
 a58533a <=( a58532a  and  a58525a );
 a58537a <=( A298  and  A268 );
 a58538a <=( (not A267)  and  a58537a );
 a58541a <=( (not A300)  and  (not A299) );
 a58544a <=( (not A302)  and  (not A301) );
 a58545a <=( a58544a  and  a58541a );
 a58546a <=( a58545a  and  a58538a );
 a58550a <=( A167  and  A168 );
 a58551a <=( (not A170)  and  a58550a );
 a58554a <=( A201  and  (not A166) );
 a58557a <=( (not A203)  and  (not A202) );
 a58558a <=( a58557a  and  a58554a );
 a58559a <=( a58558a  and  a58551a );
 a58563a <=( (not A298)  and  A268 );
 a58564a <=( (not A267)  and  a58563a );
 a58567a <=( (not A300)  and  A299 );
 a58570a <=( (not A302)  and  (not A301) );
 a58571a <=( a58570a  and  a58567a );
 a58572a <=( a58571a  and  a58564a );
 a58576a <=( A167  and  A168 );
 a58577a <=( (not A170)  and  a58576a );
 a58580a <=( A201  and  (not A166) );
 a58583a <=( (not A203)  and  (not A202) );
 a58584a <=( a58583a  and  a58580a );
 a58585a <=( a58584a  and  a58577a );
 a58589a <=( A298  and  A269 );
 a58590a <=( (not A267)  and  a58589a );
 a58593a <=( (not A300)  and  (not A299) );
 a58596a <=( (not A302)  and  (not A301) );
 a58597a <=( a58596a  and  a58593a );
 a58598a <=( a58597a  and  a58590a );
 a58602a <=( A167  and  A168 );
 a58603a <=( (not A170)  and  a58602a );
 a58606a <=( A201  and  (not A166) );
 a58609a <=( (not A203)  and  (not A202) );
 a58610a <=( a58609a  and  a58606a );
 a58611a <=( a58610a  and  a58603a );
 a58615a <=( (not A298)  and  A269 );
 a58616a <=( (not A267)  and  a58615a );
 a58619a <=( (not A300)  and  A299 );
 a58622a <=( (not A302)  and  (not A301) );
 a58623a <=( a58622a  and  a58619a );
 a58624a <=( a58623a  and  a58616a );
 a58628a <=( A167  and  A168 );
 a58629a <=( (not A170)  and  a58628a );
 a58632a <=( A201  and  (not A166) );
 a58635a <=( (not A203)  and  (not A202) );
 a58636a <=( a58635a  and  a58632a );
 a58637a <=( a58636a  and  a58629a );
 a58641a <=( A298  and  A266 );
 a58642a <=( A265  and  a58641a );
 a58645a <=( (not A300)  and  (not A299) );
 a58648a <=( (not A302)  and  (not A301) );
 a58649a <=( a58648a  and  a58645a );
 a58650a <=( a58649a  and  a58642a );
 a58654a <=( A167  and  A168 );
 a58655a <=( (not A170)  and  a58654a );
 a58658a <=( A201  and  (not A166) );
 a58661a <=( (not A203)  and  (not A202) );
 a58662a <=( a58661a  and  a58658a );
 a58663a <=( a58662a  and  a58655a );
 a58667a <=( (not A298)  and  A266 );
 a58668a <=( A265  and  a58667a );
 a58671a <=( (not A300)  and  A299 );
 a58674a <=( (not A302)  and  (not A301) );
 a58675a <=( a58674a  and  a58671a );
 a58676a <=( a58675a  and  a58668a );
 a58680a <=( A167  and  A168 );
 a58681a <=( (not A170)  and  a58680a );
 a58684a <=( A201  and  (not A166) );
 a58687a <=( (not A203)  and  (not A202) );
 a58688a <=( a58687a  and  a58684a );
 a58689a <=( a58688a  and  a58681a );
 a58693a <=( A298  and  (not A266) );
 a58694a <=( (not A265)  and  a58693a );
 a58697a <=( (not A300)  and  (not A299) );
 a58700a <=( (not A302)  and  (not A301) );
 a58701a <=( a58700a  and  a58697a );
 a58702a <=( a58701a  and  a58694a );
 a58706a <=( A167  and  A168 );
 a58707a <=( (not A170)  and  a58706a );
 a58710a <=( A201  and  (not A166) );
 a58713a <=( (not A203)  and  (not A202) );
 a58714a <=( a58713a  and  a58710a );
 a58715a <=( a58714a  and  a58707a );
 a58719a <=( (not A298)  and  (not A266) );
 a58720a <=( (not A265)  and  a58719a );
 a58723a <=( (not A300)  and  A299 );
 a58726a <=( (not A302)  and  (not A301) );
 a58727a <=( a58726a  and  a58723a );
 a58728a <=( a58727a  and  a58720a );
 a58732a <=( A167  and  A168 );
 a58733a <=( (not A170)  and  a58732a );
 a58736a <=( (not A201)  and  (not A166) );
 a58739a <=( A267  and  A202 );
 a58740a <=( a58739a  and  a58736a );
 a58741a <=( a58740a  and  a58733a );
 a58745a <=( A298  and  (not A269) );
 a58746a <=( (not A268)  and  a58745a );
 a58749a <=( (not A300)  and  (not A299) );
 a58752a <=( (not A302)  and  (not A301) );
 a58753a <=( a58752a  and  a58749a );
 a58754a <=( a58753a  and  a58746a );
 a58758a <=( A167  and  A168 );
 a58759a <=( (not A170)  and  a58758a );
 a58762a <=( (not A201)  and  (not A166) );
 a58765a <=( A267  and  A202 );
 a58766a <=( a58765a  and  a58762a );
 a58767a <=( a58766a  and  a58759a );
 a58771a <=( (not A298)  and  (not A269) );
 a58772a <=( (not A268)  and  a58771a );
 a58775a <=( (not A300)  and  A299 );
 a58778a <=( (not A302)  and  (not A301) );
 a58779a <=( a58778a  and  a58775a );
 a58780a <=( a58779a  and  a58772a );
 a58784a <=( A167  and  A168 );
 a58785a <=( (not A170)  and  a58784a );
 a58788a <=( (not A201)  and  (not A166) );
 a58791a <=( A267  and  A203 );
 a58792a <=( a58791a  and  a58788a );
 a58793a <=( a58792a  and  a58785a );
 a58797a <=( A298  and  (not A269) );
 a58798a <=( (not A268)  and  a58797a );
 a58801a <=( (not A300)  and  (not A299) );
 a58804a <=( (not A302)  and  (not A301) );
 a58805a <=( a58804a  and  a58801a );
 a58806a <=( a58805a  and  a58798a );
 a58810a <=( A167  and  A168 );
 a58811a <=( (not A170)  and  a58810a );
 a58814a <=( (not A201)  and  (not A166) );
 a58817a <=( A267  and  A203 );
 a58818a <=( a58817a  and  a58814a );
 a58819a <=( a58818a  and  a58811a );
 a58823a <=( (not A298)  and  (not A269) );
 a58824a <=( (not A268)  and  a58823a );
 a58827a <=( (not A300)  and  A299 );
 a58830a <=( (not A302)  and  (not A301) );
 a58831a <=( a58830a  and  a58827a );
 a58832a <=( a58831a  and  a58824a );
 a58836a <=( A167  and  A168 );
 a58837a <=( (not A170)  and  a58836a );
 a58840a <=( A199  and  (not A166) );
 a58843a <=( A267  and  A200 );
 a58844a <=( a58843a  and  a58840a );
 a58845a <=( a58844a  and  a58837a );
 a58849a <=( A298  and  (not A269) );
 a58850a <=( (not A268)  and  a58849a );
 a58853a <=( (not A300)  and  (not A299) );
 a58856a <=( (not A302)  and  (not A301) );
 a58857a <=( a58856a  and  a58853a );
 a58858a <=( a58857a  and  a58850a );
 a58862a <=( A167  and  A168 );
 a58863a <=( (not A170)  and  a58862a );
 a58866a <=( A199  and  (not A166) );
 a58869a <=( A267  and  A200 );
 a58870a <=( a58869a  and  a58866a );
 a58871a <=( a58870a  and  a58863a );
 a58875a <=( (not A298)  and  (not A269) );
 a58876a <=( (not A268)  and  a58875a );
 a58879a <=( (not A300)  and  A299 );
 a58882a <=( (not A302)  and  (not A301) );
 a58883a <=( a58882a  and  a58879a );
 a58884a <=( a58883a  and  a58876a );
 a58888a <=( A167  and  A168 );
 a58889a <=( (not A170)  and  a58888a );
 a58892a <=( (not A199)  and  (not A166) );
 a58895a <=( A201  and  A200 );
 a58896a <=( a58895a  and  a58892a );
 a58897a <=( a58896a  and  a58889a );
 a58901a <=( A266  and  (not A265) );
 a58902a <=( A202  and  a58901a );
 a58905a <=( A268  and  A267 );
 a58908a <=( A301  and  (not A300) );
 a58909a <=( a58908a  and  a58905a );
 a58910a <=( a58909a  and  a58902a );
 a58914a <=( A167  and  A168 );
 a58915a <=( (not A170)  and  a58914a );
 a58918a <=( (not A199)  and  (not A166) );
 a58921a <=( A201  and  A200 );
 a58922a <=( a58921a  and  a58918a );
 a58923a <=( a58922a  and  a58915a );
 a58927a <=( A266  and  (not A265) );
 a58928a <=( A202  and  a58927a );
 a58931a <=( A268  and  A267 );
 a58934a <=( A302  and  (not A300) );
 a58935a <=( a58934a  and  a58931a );
 a58936a <=( a58935a  and  a58928a );
 a58940a <=( A167  and  A168 );
 a58941a <=( (not A170)  and  a58940a );
 a58944a <=( (not A199)  and  (not A166) );
 a58947a <=( A201  and  A200 );
 a58948a <=( a58947a  and  a58944a );
 a58949a <=( a58948a  and  a58941a );
 a58953a <=( A266  and  (not A265) );
 a58954a <=( A202  and  a58953a );
 a58957a <=( A268  and  A267 );
 a58960a <=( A299  and  A298 );
 a58961a <=( a58960a  and  a58957a );
 a58962a <=( a58961a  and  a58954a );
 a58966a <=( A167  and  A168 );
 a58967a <=( (not A170)  and  a58966a );
 a58970a <=( (not A199)  and  (not A166) );
 a58973a <=( A201  and  A200 );
 a58974a <=( a58973a  and  a58970a );
 a58975a <=( a58974a  and  a58967a );
 a58979a <=( A266  and  (not A265) );
 a58980a <=( A202  and  a58979a );
 a58983a <=( A268  and  A267 );
 a58986a <=( (not A299)  and  (not A298) );
 a58987a <=( a58986a  and  a58983a );
 a58988a <=( a58987a  and  a58980a );
 a58992a <=( A167  and  A168 );
 a58993a <=( (not A170)  and  a58992a );
 a58996a <=( (not A199)  and  (not A166) );
 a58999a <=( A201  and  A200 );
 a59000a <=( a58999a  and  a58996a );
 a59001a <=( a59000a  and  a58993a );
 a59005a <=( A266  and  (not A265) );
 a59006a <=( A202  and  a59005a );
 a59009a <=( A269  and  A267 );
 a59012a <=( A301  and  (not A300) );
 a59013a <=( a59012a  and  a59009a );
 a59014a <=( a59013a  and  a59006a );
 a59018a <=( A167  and  A168 );
 a59019a <=( (not A170)  and  a59018a );
 a59022a <=( (not A199)  and  (not A166) );
 a59025a <=( A201  and  A200 );
 a59026a <=( a59025a  and  a59022a );
 a59027a <=( a59026a  and  a59019a );
 a59031a <=( A266  and  (not A265) );
 a59032a <=( A202  and  a59031a );
 a59035a <=( A269  and  A267 );
 a59038a <=( A302  and  (not A300) );
 a59039a <=( a59038a  and  a59035a );
 a59040a <=( a59039a  and  a59032a );
 a59044a <=( A167  and  A168 );
 a59045a <=( (not A170)  and  a59044a );
 a59048a <=( (not A199)  and  (not A166) );
 a59051a <=( A201  and  A200 );
 a59052a <=( a59051a  and  a59048a );
 a59053a <=( a59052a  and  a59045a );
 a59057a <=( A266  and  (not A265) );
 a59058a <=( A202  and  a59057a );
 a59061a <=( A269  and  A267 );
 a59064a <=( A299  and  A298 );
 a59065a <=( a59064a  and  a59061a );
 a59066a <=( a59065a  and  a59058a );
 a59070a <=( A167  and  A168 );
 a59071a <=( (not A170)  and  a59070a );
 a59074a <=( (not A199)  and  (not A166) );
 a59077a <=( A201  and  A200 );
 a59078a <=( a59077a  and  a59074a );
 a59079a <=( a59078a  and  a59071a );
 a59083a <=( A266  and  (not A265) );
 a59084a <=( A202  and  a59083a );
 a59087a <=( A269  and  A267 );
 a59090a <=( (not A299)  and  (not A298) );
 a59091a <=( a59090a  and  a59087a );
 a59092a <=( a59091a  and  a59084a );
 a59096a <=( A167  and  A168 );
 a59097a <=( (not A170)  and  a59096a );
 a59100a <=( (not A199)  and  (not A166) );
 a59103a <=( A201  and  A200 );
 a59104a <=( a59103a  and  a59100a );
 a59105a <=( a59104a  and  a59097a );
 a59109a <=( (not A266)  and  A265 );
 a59110a <=( A202  and  a59109a );
 a59113a <=( A268  and  A267 );
 a59116a <=( A301  and  (not A300) );
 a59117a <=( a59116a  and  a59113a );
 a59118a <=( a59117a  and  a59110a );
 a59122a <=( A167  and  A168 );
 a59123a <=( (not A170)  and  a59122a );
 a59126a <=( (not A199)  and  (not A166) );
 a59129a <=( A201  and  A200 );
 a59130a <=( a59129a  and  a59126a );
 a59131a <=( a59130a  and  a59123a );
 a59135a <=( (not A266)  and  A265 );
 a59136a <=( A202  and  a59135a );
 a59139a <=( A268  and  A267 );
 a59142a <=( A302  and  (not A300) );
 a59143a <=( a59142a  and  a59139a );
 a59144a <=( a59143a  and  a59136a );
 a59148a <=( A167  and  A168 );
 a59149a <=( (not A170)  and  a59148a );
 a59152a <=( (not A199)  and  (not A166) );
 a59155a <=( A201  and  A200 );
 a59156a <=( a59155a  and  a59152a );
 a59157a <=( a59156a  and  a59149a );
 a59161a <=( (not A266)  and  A265 );
 a59162a <=( A202  and  a59161a );
 a59165a <=( A268  and  A267 );
 a59168a <=( A299  and  A298 );
 a59169a <=( a59168a  and  a59165a );
 a59170a <=( a59169a  and  a59162a );
 a59174a <=( A167  and  A168 );
 a59175a <=( (not A170)  and  a59174a );
 a59178a <=( (not A199)  and  (not A166) );
 a59181a <=( A201  and  A200 );
 a59182a <=( a59181a  and  a59178a );
 a59183a <=( a59182a  and  a59175a );
 a59187a <=( (not A266)  and  A265 );
 a59188a <=( A202  and  a59187a );
 a59191a <=( A268  and  A267 );
 a59194a <=( (not A299)  and  (not A298) );
 a59195a <=( a59194a  and  a59191a );
 a59196a <=( a59195a  and  a59188a );
 a59200a <=( A167  and  A168 );
 a59201a <=( (not A170)  and  a59200a );
 a59204a <=( (not A199)  and  (not A166) );
 a59207a <=( A201  and  A200 );
 a59208a <=( a59207a  and  a59204a );
 a59209a <=( a59208a  and  a59201a );
 a59213a <=( (not A266)  and  A265 );
 a59214a <=( A202  and  a59213a );
 a59217a <=( A269  and  A267 );
 a59220a <=( A301  and  (not A300) );
 a59221a <=( a59220a  and  a59217a );
 a59222a <=( a59221a  and  a59214a );
 a59226a <=( A167  and  A168 );
 a59227a <=( (not A170)  and  a59226a );
 a59230a <=( (not A199)  and  (not A166) );
 a59233a <=( A201  and  A200 );
 a59234a <=( a59233a  and  a59230a );
 a59235a <=( a59234a  and  a59227a );
 a59239a <=( (not A266)  and  A265 );
 a59240a <=( A202  and  a59239a );
 a59243a <=( A269  and  A267 );
 a59246a <=( A302  and  (not A300) );
 a59247a <=( a59246a  and  a59243a );
 a59248a <=( a59247a  and  a59240a );
 a59252a <=( A167  and  A168 );
 a59253a <=( (not A170)  and  a59252a );
 a59256a <=( (not A199)  and  (not A166) );
 a59259a <=( A201  and  A200 );
 a59260a <=( a59259a  and  a59256a );
 a59261a <=( a59260a  and  a59253a );
 a59265a <=( (not A266)  and  A265 );
 a59266a <=( A202  and  a59265a );
 a59269a <=( A269  and  A267 );
 a59272a <=( A299  and  A298 );
 a59273a <=( a59272a  and  a59269a );
 a59274a <=( a59273a  and  a59266a );
 a59278a <=( A167  and  A168 );
 a59279a <=( (not A170)  and  a59278a );
 a59282a <=( (not A199)  and  (not A166) );
 a59285a <=( A201  and  A200 );
 a59286a <=( a59285a  and  a59282a );
 a59287a <=( a59286a  and  a59279a );
 a59291a <=( (not A266)  and  A265 );
 a59292a <=( A202  and  a59291a );
 a59295a <=( A269  and  A267 );
 a59298a <=( (not A299)  and  (not A298) );
 a59299a <=( a59298a  and  a59295a );
 a59300a <=( a59299a  and  a59292a );
 a59304a <=( A167  and  A168 );
 a59305a <=( (not A170)  and  a59304a );
 a59308a <=( (not A199)  and  (not A166) );
 a59311a <=( A201  and  A200 );
 a59312a <=( a59311a  and  a59308a );
 a59313a <=( a59312a  and  a59305a );
 a59317a <=( A266  and  (not A265) );
 a59318a <=( A203  and  a59317a );
 a59321a <=( A268  and  A267 );
 a59324a <=( A301  and  (not A300) );
 a59325a <=( a59324a  and  a59321a );
 a59326a <=( a59325a  and  a59318a );
 a59330a <=( A167  and  A168 );
 a59331a <=( (not A170)  and  a59330a );
 a59334a <=( (not A199)  and  (not A166) );
 a59337a <=( A201  and  A200 );
 a59338a <=( a59337a  and  a59334a );
 a59339a <=( a59338a  and  a59331a );
 a59343a <=( A266  and  (not A265) );
 a59344a <=( A203  and  a59343a );
 a59347a <=( A268  and  A267 );
 a59350a <=( A302  and  (not A300) );
 a59351a <=( a59350a  and  a59347a );
 a59352a <=( a59351a  and  a59344a );
 a59356a <=( A167  and  A168 );
 a59357a <=( (not A170)  and  a59356a );
 a59360a <=( (not A199)  and  (not A166) );
 a59363a <=( A201  and  A200 );
 a59364a <=( a59363a  and  a59360a );
 a59365a <=( a59364a  and  a59357a );
 a59369a <=( A266  and  (not A265) );
 a59370a <=( A203  and  a59369a );
 a59373a <=( A268  and  A267 );
 a59376a <=( A299  and  A298 );
 a59377a <=( a59376a  and  a59373a );
 a59378a <=( a59377a  and  a59370a );
 a59382a <=( A167  and  A168 );
 a59383a <=( (not A170)  and  a59382a );
 a59386a <=( (not A199)  and  (not A166) );
 a59389a <=( A201  and  A200 );
 a59390a <=( a59389a  and  a59386a );
 a59391a <=( a59390a  and  a59383a );
 a59395a <=( A266  and  (not A265) );
 a59396a <=( A203  and  a59395a );
 a59399a <=( A268  and  A267 );
 a59402a <=( (not A299)  and  (not A298) );
 a59403a <=( a59402a  and  a59399a );
 a59404a <=( a59403a  and  a59396a );
 a59408a <=( A167  and  A168 );
 a59409a <=( (not A170)  and  a59408a );
 a59412a <=( (not A199)  and  (not A166) );
 a59415a <=( A201  and  A200 );
 a59416a <=( a59415a  and  a59412a );
 a59417a <=( a59416a  and  a59409a );
 a59421a <=( A266  and  (not A265) );
 a59422a <=( A203  and  a59421a );
 a59425a <=( A269  and  A267 );
 a59428a <=( A301  and  (not A300) );
 a59429a <=( a59428a  and  a59425a );
 a59430a <=( a59429a  and  a59422a );
 a59434a <=( A167  and  A168 );
 a59435a <=( (not A170)  and  a59434a );
 a59438a <=( (not A199)  and  (not A166) );
 a59441a <=( A201  and  A200 );
 a59442a <=( a59441a  and  a59438a );
 a59443a <=( a59442a  and  a59435a );
 a59447a <=( A266  and  (not A265) );
 a59448a <=( A203  and  a59447a );
 a59451a <=( A269  and  A267 );
 a59454a <=( A302  and  (not A300) );
 a59455a <=( a59454a  and  a59451a );
 a59456a <=( a59455a  and  a59448a );
 a59460a <=( A167  and  A168 );
 a59461a <=( (not A170)  and  a59460a );
 a59464a <=( (not A199)  and  (not A166) );
 a59467a <=( A201  and  A200 );
 a59468a <=( a59467a  and  a59464a );
 a59469a <=( a59468a  and  a59461a );
 a59473a <=( A266  and  (not A265) );
 a59474a <=( A203  and  a59473a );
 a59477a <=( A269  and  A267 );
 a59480a <=( A299  and  A298 );
 a59481a <=( a59480a  and  a59477a );
 a59482a <=( a59481a  and  a59474a );
 a59486a <=( A167  and  A168 );
 a59487a <=( (not A170)  and  a59486a );
 a59490a <=( (not A199)  and  (not A166) );
 a59493a <=( A201  and  A200 );
 a59494a <=( a59493a  and  a59490a );
 a59495a <=( a59494a  and  a59487a );
 a59499a <=( A266  and  (not A265) );
 a59500a <=( A203  and  a59499a );
 a59503a <=( A269  and  A267 );
 a59506a <=( (not A299)  and  (not A298) );
 a59507a <=( a59506a  and  a59503a );
 a59508a <=( a59507a  and  a59500a );
 a59512a <=( A167  and  A168 );
 a59513a <=( (not A170)  and  a59512a );
 a59516a <=( (not A199)  and  (not A166) );
 a59519a <=( A201  and  A200 );
 a59520a <=( a59519a  and  a59516a );
 a59521a <=( a59520a  and  a59513a );
 a59525a <=( (not A266)  and  A265 );
 a59526a <=( A203  and  a59525a );
 a59529a <=( A268  and  A267 );
 a59532a <=( A301  and  (not A300) );
 a59533a <=( a59532a  and  a59529a );
 a59534a <=( a59533a  and  a59526a );
 a59538a <=( A167  and  A168 );
 a59539a <=( (not A170)  and  a59538a );
 a59542a <=( (not A199)  and  (not A166) );
 a59545a <=( A201  and  A200 );
 a59546a <=( a59545a  and  a59542a );
 a59547a <=( a59546a  and  a59539a );
 a59551a <=( (not A266)  and  A265 );
 a59552a <=( A203  and  a59551a );
 a59555a <=( A268  and  A267 );
 a59558a <=( A302  and  (not A300) );
 a59559a <=( a59558a  and  a59555a );
 a59560a <=( a59559a  and  a59552a );
 a59564a <=( A167  and  A168 );
 a59565a <=( (not A170)  and  a59564a );
 a59568a <=( (not A199)  and  (not A166) );
 a59571a <=( A201  and  A200 );
 a59572a <=( a59571a  and  a59568a );
 a59573a <=( a59572a  and  a59565a );
 a59577a <=( (not A266)  and  A265 );
 a59578a <=( A203  and  a59577a );
 a59581a <=( A268  and  A267 );
 a59584a <=( A299  and  A298 );
 a59585a <=( a59584a  and  a59581a );
 a59586a <=( a59585a  and  a59578a );
 a59590a <=( A167  and  A168 );
 a59591a <=( (not A170)  and  a59590a );
 a59594a <=( (not A199)  and  (not A166) );
 a59597a <=( A201  and  A200 );
 a59598a <=( a59597a  and  a59594a );
 a59599a <=( a59598a  and  a59591a );
 a59603a <=( (not A266)  and  A265 );
 a59604a <=( A203  and  a59603a );
 a59607a <=( A268  and  A267 );
 a59610a <=( (not A299)  and  (not A298) );
 a59611a <=( a59610a  and  a59607a );
 a59612a <=( a59611a  and  a59604a );
 a59616a <=( A167  and  A168 );
 a59617a <=( (not A170)  and  a59616a );
 a59620a <=( (not A199)  and  (not A166) );
 a59623a <=( A201  and  A200 );
 a59624a <=( a59623a  and  a59620a );
 a59625a <=( a59624a  and  a59617a );
 a59629a <=( (not A266)  and  A265 );
 a59630a <=( A203  and  a59629a );
 a59633a <=( A269  and  A267 );
 a59636a <=( A301  and  (not A300) );
 a59637a <=( a59636a  and  a59633a );
 a59638a <=( a59637a  and  a59630a );
 a59642a <=( A167  and  A168 );
 a59643a <=( (not A170)  and  a59642a );
 a59646a <=( (not A199)  and  (not A166) );
 a59649a <=( A201  and  A200 );
 a59650a <=( a59649a  and  a59646a );
 a59651a <=( a59650a  and  a59643a );
 a59655a <=( (not A266)  and  A265 );
 a59656a <=( A203  and  a59655a );
 a59659a <=( A269  and  A267 );
 a59662a <=( A302  and  (not A300) );
 a59663a <=( a59662a  and  a59659a );
 a59664a <=( a59663a  and  a59656a );
 a59668a <=( A167  and  A168 );
 a59669a <=( (not A170)  and  a59668a );
 a59672a <=( (not A199)  and  (not A166) );
 a59675a <=( A201  and  A200 );
 a59676a <=( a59675a  and  a59672a );
 a59677a <=( a59676a  and  a59669a );
 a59681a <=( (not A266)  and  A265 );
 a59682a <=( A203  and  a59681a );
 a59685a <=( A269  and  A267 );
 a59688a <=( A299  and  A298 );
 a59689a <=( a59688a  and  a59685a );
 a59690a <=( a59689a  and  a59682a );
 a59694a <=( A167  and  A168 );
 a59695a <=( (not A170)  and  a59694a );
 a59698a <=( (not A199)  and  (not A166) );
 a59701a <=( A201  and  A200 );
 a59702a <=( a59701a  and  a59698a );
 a59703a <=( a59702a  and  a59695a );
 a59707a <=( (not A266)  and  A265 );
 a59708a <=( A203  and  a59707a );
 a59711a <=( A269  and  A267 );
 a59714a <=( (not A299)  and  (not A298) );
 a59715a <=( a59714a  and  a59711a );
 a59716a <=( a59715a  and  a59708a );
 a59720a <=( A167  and  A168 );
 a59721a <=( (not A170)  and  a59720a );
 a59724a <=( A199  and  (not A166) );
 a59727a <=( A201  and  (not A200) );
 a59728a <=( a59727a  and  a59724a );
 a59729a <=( a59728a  and  a59721a );
 a59733a <=( A266  and  (not A265) );
 a59734a <=( A202  and  a59733a );
 a59737a <=( A268  and  A267 );
 a59740a <=( A301  and  (not A300) );
 a59741a <=( a59740a  and  a59737a );
 a59742a <=( a59741a  and  a59734a );
 a59746a <=( A167  and  A168 );
 a59747a <=( (not A170)  and  a59746a );
 a59750a <=( A199  and  (not A166) );
 a59753a <=( A201  and  (not A200) );
 a59754a <=( a59753a  and  a59750a );
 a59755a <=( a59754a  and  a59747a );
 a59759a <=( A266  and  (not A265) );
 a59760a <=( A202  and  a59759a );
 a59763a <=( A268  and  A267 );
 a59766a <=( A302  and  (not A300) );
 a59767a <=( a59766a  and  a59763a );
 a59768a <=( a59767a  and  a59760a );
 a59772a <=( A167  and  A168 );
 a59773a <=( (not A170)  and  a59772a );
 a59776a <=( A199  and  (not A166) );
 a59779a <=( A201  and  (not A200) );
 a59780a <=( a59779a  and  a59776a );
 a59781a <=( a59780a  and  a59773a );
 a59785a <=( A266  and  (not A265) );
 a59786a <=( A202  and  a59785a );
 a59789a <=( A268  and  A267 );
 a59792a <=( A299  and  A298 );
 a59793a <=( a59792a  and  a59789a );
 a59794a <=( a59793a  and  a59786a );
 a59798a <=( A167  and  A168 );
 a59799a <=( (not A170)  and  a59798a );
 a59802a <=( A199  and  (not A166) );
 a59805a <=( A201  and  (not A200) );
 a59806a <=( a59805a  and  a59802a );
 a59807a <=( a59806a  and  a59799a );
 a59811a <=( A266  and  (not A265) );
 a59812a <=( A202  and  a59811a );
 a59815a <=( A268  and  A267 );
 a59818a <=( (not A299)  and  (not A298) );
 a59819a <=( a59818a  and  a59815a );
 a59820a <=( a59819a  and  a59812a );
 a59824a <=( A167  and  A168 );
 a59825a <=( (not A170)  and  a59824a );
 a59828a <=( A199  and  (not A166) );
 a59831a <=( A201  and  (not A200) );
 a59832a <=( a59831a  and  a59828a );
 a59833a <=( a59832a  and  a59825a );
 a59837a <=( A266  and  (not A265) );
 a59838a <=( A202  and  a59837a );
 a59841a <=( A269  and  A267 );
 a59844a <=( A301  and  (not A300) );
 a59845a <=( a59844a  and  a59841a );
 a59846a <=( a59845a  and  a59838a );
 a59850a <=( A167  and  A168 );
 a59851a <=( (not A170)  and  a59850a );
 a59854a <=( A199  and  (not A166) );
 a59857a <=( A201  and  (not A200) );
 a59858a <=( a59857a  and  a59854a );
 a59859a <=( a59858a  and  a59851a );
 a59863a <=( A266  and  (not A265) );
 a59864a <=( A202  and  a59863a );
 a59867a <=( A269  and  A267 );
 a59870a <=( A302  and  (not A300) );
 a59871a <=( a59870a  and  a59867a );
 a59872a <=( a59871a  and  a59864a );
 a59876a <=( A167  and  A168 );
 a59877a <=( (not A170)  and  a59876a );
 a59880a <=( A199  and  (not A166) );
 a59883a <=( A201  and  (not A200) );
 a59884a <=( a59883a  and  a59880a );
 a59885a <=( a59884a  and  a59877a );
 a59889a <=( A266  and  (not A265) );
 a59890a <=( A202  and  a59889a );
 a59893a <=( A269  and  A267 );
 a59896a <=( A299  and  A298 );
 a59897a <=( a59896a  and  a59893a );
 a59898a <=( a59897a  and  a59890a );
 a59902a <=( A167  and  A168 );
 a59903a <=( (not A170)  and  a59902a );
 a59906a <=( A199  and  (not A166) );
 a59909a <=( A201  and  (not A200) );
 a59910a <=( a59909a  and  a59906a );
 a59911a <=( a59910a  and  a59903a );
 a59915a <=( A266  and  (not A265) );
 a59916a <=( A202  and  a59915a );
 a59919a <=( A269  and  A267 );
 a59922a <=( (not A299)  and  (not A298) );
 a59923a <=( a59922a  and  a59919a );
 a59924a <=( a59923a  and  a59916a );
 a59928a <=( A167  and  A168 );
 a59929a <=( (not A170)  and  a59928a );
 a59932a <=( A199  and  (not A166) );
 a59935a <=( A201  and  (not A200) );
 a59936a <=( a59935a  and  a59932a );
 a59937a <=( a59936a  and  a59929a );
 a59941a <=( (not A266)  and  A265 );
 a59942a <=( A202  and  a59941a );
 a59945a <=( A268  and  A267 );
 a59948a <=( A301  and  (not A300) );
 a59949a <=( a59948a  and  a59945a );
 a59950a <=( a59949a  and  a59942a );
 a59954a <=( A167  and  A168 );
 a59955a <=( (not A170)  and  a59954a );
 a59958a <=( A199  and  (not A166) );
 a59961a <=( A201  and  (not A200) );
 a59962a <=( a59961a  and  a59958a );
 a59963a <=( a59962a  and  a59955a );
 a59967a <=( (not A266)  and  A265 );
 a59968a <=( A202  and  a59967a );
 a59971a <=( A268  and  A267 );
 a59974a <=( A302  and  (not A300) );
 a59975a <=( a59974a  and  a59971a );
 a59976a <=( a59975a  and  a59968a );
 a59980a <=( A167  and  A168 );
 a59981a <=( (not A170)  and  a59980a );
 a59984a <=( A199  and  (not A166) );
 a59987a <=( A201  and  (not A200) );
 a59988a <=( a59987a  and  a59984a );
 a59989a <=( a59988a  and  a59981a );
 a59993a <=( (not A266)  and  A265 );
 a59994a <=( A202  and  a59993a );
 a59997a <=( A268  and  A267 );
 a60000a <=( A299  and  A298 );
 a60001a <=( a60000a  and  a59997a );
 a60002a <=( a60001a  and  a59994a );
 a60006a <=( A167  and  A168 );
 a60007a <=( (not A170)  and  a60006a );
 a60010a <=( A199  and  (not A166) );
 a60013a <=( A201  and  (not A200) );
 a60014a <=( a60013a  and  a60010a );
 a60015a <=( a60014a  and  a60007a );
 a60019a <=( (not A266)  and  A265 );
 a60020a <=( A202  and  a60019a );
 a60023a <=( A268  and  A267 );
 a60026a <=( (not A299)  and  (not A298) );
 a60027a <=( a60026a  and  a60023a );
 a60028a <=( a60027a  and  a60020a );
 a60032a <=( A167  and  A168 );
 a60033a <=( (not A170)  and  a60032a );
 a60036a <=( A199  and  (not A166) );
 a60039a <=( A201  and  (not A200) );
 a60040a <=( a60039a  and  a60036a );
 a60041a <=( a60040a  and  a60033a );
 a60045a <=( (not A266)  and  A265 );
 a60046a <=( A202  and  a60045a );
 a60049a <=( A269  and  A267 );
 a60052a <=( A301  and  (not A300) );
 a60053a <=( a60052a  and  a60049a );
 a60054a <=( a60053a  and  a60046a );
 a60058a <=( A167  and  A168 );
 a60059a <=( (not A170)  and  a60058a );
 a60062a <=( A199  and  (not A166) );
 a60065a <=( A201  and  (not A200) );
 a60066a <=( a60065a  and  a60062a );
 a60067a <=( a60066a  and  a60059a );
 a60071a <=( (not A266)  and  A265 );
 a60072a <=( A202  and  a60071a );
 a60075a <=( A269  and  A267 );
 a60078a <=( A302  and  (not A300) );
 a60079a <=( a60078a  and  a60075a );
 a60080a <=( a60079a  and  a60072a );
 a60084a <=( A167  and  A168 );
 a60085a <=( (not A170)  and  a60084a );
 a60088a <=( A199  and  (not A166) );
 a60091a <=( A201  and  (not A200) );
 a60092a <=( a60091a  and  a60088a );
 a60093a <=( a60092a  and  a60085a );
 a60097a <=( (not A266)  and  A265 );
 a60098a <=( A202  and  a60097a );
 a60101a <=( A269  and  A267 );
 a60104a <=( A299  and  A298 );
 a60105a <=( a60104a  and  a60101a );
 a60106a <=( a60105a  and  a60098a );
 a60110a <=( A167  and  A168 );
 a60111a <=( (not A170)  and  a60110a );
 a60114a <=( A199  and  (not A166) );
 a60117a <=( A201  and  (not A200) );
 a60118a <=( a60117a  and  a60114a );
 a60119a <=( a60118a  and  a60111a );
 a60123a <=( (not A266)  and  A265 );
 a60124a <=( A202  and  a60123a );
 a60127a <=( A269  and  A267 );
 a60130a <=( (not A299)  and  (not A298) );
 a60131a <=( a60130a  and  a60127a );
 a60132a <=( a60131a  and  a60124a );
 a60136a <=( A167  and  A168 );
 a60137a <=( (not A170)  and  a60136a );
 a60140a <=( A199  and  (not A166) );
 a60143a <=( A201  and  (not A200) );
 a60144a <=( a60143a  and  a60140a );
 a60145a <=( a60144a  and  a60137a );
 a60149a <=( A266  and  (not A265) );
 a60150a <=( A203  and  a60149a );
 a60153a <=( A268  and  A267 );
 a60156a <=( A301  and  (not A300) );
 a60157a <=( a60156a  and  a60153a );
 a60158a <=( a60157a  and  a60150a );
 a60162a <=( A167  and  A168 );
 a60163a <=( (not A170)  and  a60162a );
 a60166a <=( A199  and  (not A166) );
 a60169a <=( A201  and  (not A200) );
 a60170a <=( a60169a  and  a60166a );
 a60171a <=( a60170a  and  a60163a );
 a60175a <=( A266  and  (not A265) );
 a60176a <=( A203  and  a60175a );
 a60179a <=( A268  and  A267 );
 a60182a <=( A302  and  (not A300) );
 a60183a <=( a60182a  and  a60179a );
 a60184a <=( a60183a  and  a60176a );
 a60188a <=( A167  and  A168 );
 a60189a <=( (not A170)  and  a60188a );
 a60192a <=( A199  and  (not A166) );
 a60195a <=( A201  and  (not A200) );
 a60196a <=( a60195a  and  a60192a );
 a60197a <=( a60196a  and  a60189a );
 a60201a <=( A266  and  (not A265) );
 a60202a <=( A203  and  a60201a );
 a60205a <=( A268  and  A267 );
 a60208a <=( A299  and  A298 );
 a60209a <=( a60208a  and  a60205a );
 a60210a <=( a60209a  and  a60202a );
 a60214a <=( A167  and  A168 );
 a60215a <=( (not A170)  and  a60214a );
 a60218a <=( A199  and  (not A166) );
 a60221a <=( A201  and  (not A200) );
 a60222a <=( a60221a  and  a60218a );
 a60223a <=( a60222a  and  a60215a );
 a60227a <=( A266  and  (not A265) );
 a60228a <=( A203  and  a60227a );
 a60231a <=( A268  and  A267 );
 a60234a <=( (not A299)  and  (not A298) );
 a60235a <=( a60234a  and  a60231a );
 a60236a <=( a60235a  and  a60228a );
 a60240a <=( A167  and  A168 );
 a60241a <=( (not A170)  and  a60240a );
 a60244a <=( A199  and  (not A166) );
 a60247a <=( A201  and  (not A200) );
 a60248a <=( a60247a  and  a60244a );
 a60249a <=( a60248a  and  a60241a );
 a60253a <=( A266  and  (not A265) );
 a60254a <=( A203  and  a60253a );
 a60257a <=( A269  and  A267 );
 a60260a <=( A301  and  (not A300) );
 a60261a <=( a60260a  and  a60257a );
 a60262a <=( a60261a  and  a60254a );
 a60266a <=( A167  and  A168 );
 a60267a <=( (not A170)  and  a60266a );
 a60270a <=( A199  and  (not A166) );
 a60273a <=( A201  and  (not A200) );
 a60274a <=( a60273a  and  a60270a );
 a60275a <=( a60274a  and  a60267a );
 a60279a <=( A266  and  (not A265) );
 a60280a <=( A203  and  a60279a );
 a60283a <=( A269  and  A267 );
 a60286a <=( A302  and  (not A300) );
 a60287a <=( a60286a  and  a60283a );
 a60288a <=( a60287a  and  a60280a );
 a60292a <=( A167  and  A168 );
 a60293a <=( (not A170)  and  a60292a );
 a60296a <=( A199  and  (not A166) );
 a60299a <=( A201  and  (not A200) );
 a60300a <=( a60299a  and  a60296a );
 a60301a <=( a60300a  and  a60293a );
 a60305a <=( A266  and  (not A265) );
 a60306a <=( A203  and  a60305a );
 a60309a <=( A269  and  A267 );
 a60312a <=( A299  and  A298 );
 a60313a <=( a60312a  and  a60309a );
 a60314a <=( a60313a  and  a60306a );
 a60318a <=( A167  and  A168 );
 a60319a <=( (not A170)  and  a60318a );
 a60322a <=( A199  and  (not A166) );
 a60325a <=( A201  and  (not A200) );
 a60326a <=( a60325a  and  a60322a );
 a60327a <=( a60326a  and  a60319a );
 a60331a <=( A266  and  (not A265) );
 a60332a <=( A203  and  a60331a );
 a60335a <=( A269  and  A267 );
 a60338a <=( (not A299)  and  (not A298) );
 a60339a <=( a60338a  and  a60335a );
 a60340a <=( a60339a  and  a60332a );
 a60344a <=( A167  and  A168 );
 a60345a <=( (not A170)  and  a60344a );
 a60348a <=( A199  and  (not A166) );
 a60351a <=( A201  and  (not A200) );
 a60352a <=( a60351a  and  a60348a );
 a60353a <=( a60352a  and  a60345a );
 a60357a <=( (not A266)  and  A265 );
 a60358a <=( A203  and  a60357a );
 a60361a <=( A268  and  A267 );
 a60364a <=( A301  and  (not A300) );
 a60365a <=( a60364a  and  a60361a );
 a60366a <=( a60365a  and  a60358a );
 a60370a <=( A167  and  A168 );
 a60371a <=( (not A170)  and  a60370a );
 a60374a <=( A199  and  (not A166) );
 a60377a <=( A201  and  (not A200) );
 a60378a <=( a60377a  and  a60374a );
 a60379a <=( a60378a  and  a60371a );
 a60383a <=( (not A266)  and  A265 );
 a60384a <=( A203  and  a60383a );
 a60387a <=( A268  and  A267 );
 a60390a <=( A302  and  (not A300) );
 a60391a <=( a60390a  and  a60387a );
 a60392a <=( a60391a  and  a60384a );
 a60396a <=( A167  and  A168 );
 a60397a <=( (not A170)  and  a60396a );
 a60400a <=( A199  and  (not A166) );
 a60403a <=( A201  and  (not A200) );
 a60404a <=( a60403a  and  a60400a );
 a60405a <=( a60404a  and  a60397a );
 a60409a <=( (not A266)  and  A265 );
 a60410a <=( A203  and  a60409a );
 a60413a <=( A268  and  A267 );
 a60416a <=( A299  and  A298 );
 a60417a <=( a60416a  and  a60413a );
 a60418a <=( a60417a  and  a60410a );
 a60422a <=( A167  and  A168 );
 a60423a <=( (not A170)  and  a60422a );
 a60426a <=( A199  and  (not A166) );
 a60429a <=( A201  and  (not A200) );
 a60430a <=( a60429a  and  a60426a );
 a60431a <=( a60430a  and  a60423a );
 a60435a <=( (not A266)  and  A265 );
 a60436a <=( A203  and  a60435a );
 a60439a <=( A268  and  A267 );
 a60442a <=( (not A299)  and  (not A298) );
 a60443a <=( a60442a  and  a60439a );
 a60444a <=( a60443a  and  a60436a );
 a60448a <=( A167  and  A168 );
 a60449a <=( (not A170)  and  a60448a );
 a60452a <=( A199  and  (not A166) );
 a60455a <=( A201  and  (not A200) );
 a60456a <=( a60455a  and  a60452a );
 a60457a <=( a60456a  and  a60449a );
 a60461a <=( (not A266)  and  A265 );
 a60462a <=( A203  and  a60461a );
 a60465a <=( A269  and  A267 );
 a60468a <=( A301  and  (not A300) );
 a60469a <=( a60468a  and  a60465a );
 a60470a <=( a60469a  and  a60462a );
 a60474a <=( A167  and  A168 );
 a60475a <=( (not A170)  and  a60474a );
 a60478a <=( A199  and  (not A166) );
 a60481a <=( A201  and  (not A200) );
 a60482a <=( a60481a  and  a60478a );
 a60483a <=( a60482a  and  a60475a );
 a60487a <=( (not A266)  and  A265 );
 a60488a <=( A203  and  a60487a );
 a60491a <=( A269  and  A267 );
 a60494a <=( A302  and  (not A300) );
 a60495a <=( a60494a  and  a60491a );
 a60496a <=( a60495a  and  a60488a );
 a60500a <=( A167  and  A168 );
 a60501a <=( (not A170)  and  a60500a );
 a60504a <=( A199  and  (not A166) );
 a60507a <=( A201  and  (not A200) );
 a60508a <=( a60507a  and  a60504a );
 a60509a <=( a60508a  and  a60501a );
 a60513a <=( (not A266)  and  A265 );
 a60514a <=( A203  and  a60513a );
 a60517a <=( A269  and  A267 );
 a60520a <=( A299  and  A298 );
 a60521a <=( a60520a  and  a60517a );
 a60522a <=( a60521a  and  a60514a );
 a60526a <=( A167  and  A168 );
 a60527a <=( (not A170)  and  a60526a );
 a60530a <=( A199  and  (not A166) );
 a60533a <=( A201  and  (not A200) );
 a60534a <=( a60533a  and  a60530a );
 a60535a <=( a60534a  and  a60527a );
 a60539a <=( (not A266)  and  A265 );
 a60540a <=( A203  and  a60539a );
 a60543a <=( A269  and  A267 );
 a60546a <=( (not A299)  and  (not A298) );
 a60547a <=( a60546a  and  a60543a );
 a60548a <=( a60547a  and  a60540a );
 a60552a <=( A167  and  A168 );
 a60553a <=( (not A170)  and  a60552a );
 a60556a <=( (not A199)  and  (not A166) );
 a60559a <=( A267  and  (not A200) );
 a60560a <=( a60559a  and  a60556a );
 a60561a <=( a60560a  and  a60553a );
 a60565a <=( A298  and  (not A269) );
 a60566a <=( (not A268)  and  a60565a );
 a60569a <=( (not A300)  and  (not A299) );
 a60572a <=( (not A302)  and  (not A301) );
 a60573a <=( a60572a  and  a60569a );
 a60574a <=( a60573a  and  a60566a );
 a60578a <=( A167  and  A168 );
 a60579a <=( (not A170)  and  a60578a );
 a60582a <=( (not A199)  and  (not A166) );
 a60585a <=( A267  and  (not A200) );
 a60586a <=( a60585a  and  a60582a );
 a60587a <=( a60586a  and  a60579a );
 a60591a <=( (not A298)  and  (not A269) );
 a60592a <=( (not A268)  and  a60591a );
 a60595a <=( (not A300)  and  A299 );
 a60598a <=( (not A302)  and  (not A301) );
 a60599a <=( a60598a  and  a60595a );
 a60600a <=( a60599a  and  a60592a );
 a60604a <=( (not A167)  and  A168 );
 a60605a <=( (not A170)  and  a60604a );
 a60608a <=( A201  and  A166 );
 a60611a <=( (not A203)  and  (not A202) );
 a60612a <=( a60611a  and  a60608a );
 a60613a <=( a60612a  and  a60605a );
 a60617a <=( (not A269)  and  (not A268) );
 a60618a <=( A267  and  a60617a );
 a60621a <=( (not A299)  and  A298 );
 a60624a <=( A301  and  A300 );
 a60625a <=( a60624a  and  a60621a );
 a60626a <=( a60625a  and  a60618a );
 a60630a <=( (not A167)  and  A168 );
 a60631a <=( (not A170)  and  a60630a );
 a60634a <=( A201  and  A166 );
 a60637a <=( (not A203)  and  (not A202) );
 a60638a <=( a60637a  and  a60634a );
 a60639a <=( a60638a  and  a60631a );
 a60643a <=( (not A269)  and  (not A268) );
 a60644a <=( A267  and  a60643a );
 a60647a <=( (not A299)  and  A298 );
 a60650a <=( A302  and  A300 );
 a60651a <=( a60650a  and  a60647a );
 a60652a <=( a60651a  and  a60644a );
 a60656a <=( (not A167)  and  A168 );
 a60657a <=( (not A170)  and  a60656a );
 a60660a <=( A201  and  A166 );
 a60663a <=( (not A203)  and  (not A202) );
 a60664a <=( a60663a  and  a60660a );
 a60665a <=( a60664a  and  a60657a );
 a60669a <=( (not A269)  and  (not A268) );
 a60670a <=( A267  and  a60669a );
 a60673a <=( A299  and  (not A298) );
 a60676a <=( A301  and  A300 );
 a60677a <=( a60676a  and  a60673a );
 a60678a <=( a60677a  and  a60670a );
 a60682a <=( (not A167)  and  A168 );
 a60683a <=( (not A170)  and  a60682a );
 a60686a <=( A201  and  A166 );
 a60689a <=( (not A203)  and  (not A202) );
 a60690a <=( a60689a  and  a60686a );
 a60691a <=( a60690a  and  a60683a );
 a60695a <=( (not A269)  and  (not A268) );
 a60696a <=( A267  and  a60695a );
 a60699a <=( A299  and  (not A298) );
 a60702a <=( A302  and  A300 );
 a60703a <=( a60702a  and  a60699a );
 a60704a <=( a60703a  and  a60696a );
 a60708a <=( (not A167)  and  A168 );
 a60709a <=( (not A170)  and  a60708a );
 a60712a <=( A201  and  A166 );
 a60715a <=( (not A203)  and  (not A202) );
 a60716a <=( a60715a  and  a60712a );
 a60717a <=( a60716a  and  a60709a );
 a60721a <=( A298  and  A268 );
 a60722a <=( (not A267)  and  a60721a );
 a60725a <=( (not A300)  and  (not A299) );
 a60728a <=( (not A302)  and  (not A301) );
 a60729a <=( a60728a  and  a60725a );
 a60730a <=( a60729a  and  a60722a );
 a60734a <=( (not A167)  and  A168 );
 a60735a <=( (not A170)  and  a60734a );
 a60738a <=( A201  and  A166 );
 a60741a <=( (not A203)  and  (not A202) );
 a60742a <=( a60741a  and  a60738a );
 a60743a <=( a60742a  and  a60735a );
 a60747a <=( (not A298)  and  A268 );
 a60748a <=( (not A267)  and  a60747a );
 a60751a <=( (not A300)  and  A299 );
 a60754a <=( (not A302)  and  (not A301) );
 a60755a <=( a60754a  and  a60751a );
 a60756a <=( a60755a  and  a60748a );
 a60760a <=( (not A167)  and  A168 );
 a60761a <=( (not A170)  and  a60760a );
 a60764a <=( A201  and  A166 );
 a60767a <=( (not A203)  and  (not A202) );
 a60768a <=( a60767a  and  a60764a );
 a60769a <=( a60768a  and  a60761a );
 a60773a <=( A298  and  A269 );
 a60774a <=( (not A267)  and  a60773a );
 a60777a <=( (not A300)  and  (not A299) );
 a60780a <=( (not A302)  and  (not A301) );
 a60781a <=( a60780a  and  a60777a );
 a60782a <=( a60781a  and  a60774a );
 a60786a <=( (not A167)  and  A168 );
 a60787a <=( (not A170)  and  a60786a );
 a60790a <=( A201  and  A166 );
 a60793a <=( (not A203)  and  (not A202) );
 a60794a <=( a60793a  and  a60790a );
 a60795a <=( a60794a  and  a60787a );
 a60799a <=( (not A298)  and  A269 );
 a60800a <=( (not A267)  and  a60799a );
 a60803a <=( (not A300)  and  A299 );
 a60806a <=( (not A302)  and  (not A301) );
 a60807a <=( a60806a  and  a60803a );
 a60808a <=( a60807a  and  a60800a );
 a60812a <=( (not A167)  and  A168 );
 a60813a <=( (not A170)  and  a60812a );
 a60816a <=( A201  and  A166 );
 a60819a <=( (not A203)  and  (not A202) );
 a60820a <=( a60819a  and  a60816a );
 a60821a <=( a60820a  and  a60813a );
 a60825a <=( A298  and  A266 );
 a60826a <=( A265  and  a60825a );
 a60829a <=( (not A300)  and  (not A299) );
 a60832a <=( (not A302)  and  (not A301) );
 a60833a <=( a60832a  and  a60829a );
 a60834a <=( a60833a  and  a60826a );
 a60838a <=( (not A167)  and  A168 );
 a60839a <=( (not A170)  and  a60838a );
 a60842a <=( A201  and  A166 );
 a60845a <=( (not A203)  and  (not A202) );
 a60846a <=( a60845a  and  a60842a );
 a60847a <=( a60846a  and  a60839a );
 a60851a <=( (not A298)  and  A266 );
 a60852a <=( A265  and  a60851a );
 a60855a <=( (not A300)  and  A299 );
 a60858a <=( (not A302)  and  (not A301) );
 a60859a <=( a60858a  and  a60855a );
 a60860a <=( a60859a  and  a60852a );
 a60864a <=( (not A167)  and  A168 );
 a60865a <=( (not A170)  and  a60864a );
 a60868a <=( A201  and  A166 );
 a60871a <=( (not A203)  and  (not A202) );
 a60872a <=( a60871a  and  a60868a );
 a60873a <=( a60872a  and  a60865a );
 a60877a <=( A298  and  (not A266) );
 a60878a <=( (not A265)  and  a60877a );
 a60881a <=( (not A300)  and  (not A299) );
 a60884a <=( (not A302)  and  (not A301) );
 a60885a <=( a60884a  and  a60881a );
 a60886a <=( a60885a  and  a60878a );
 a60890a <=( (not A167)  and  A168 );
 a60891a <=( (not A170)  and  a60890a );
 a60894a <=( A201  and  A166 );
 a60897a <=( (not A203)  and  (not A202) );
 a60898a <=( a60897a  and  a60894a );
 a60899a <=( a60898a  and  a60891a );
 a60903a <=( (not A298)  and  (not A266) );
 a60904a <=( (not A265)  and  a60903a );
 a60907a <=( (not A300)  and  A299 );
 a60910a <=( (not A302)  and  (not A301) );
 a60911a <=( a60910a  and  a60907a );
 a60912a <=( a60911a  and  a60904a );
 a60916a <=( (not A167)  and  A168 );
 a60917a <=( (not A170)  and  a60916a );
 a60920a <=( (not A201)  and  A166 );
 a60923a <=( A267  and  A202 );
 a60924a <=( a60923a  and  a60920a );
 a60925a <=( a60924a  and  a60917a );
 a60929a <=( A298  and  (not A269) );
 a60930a <=( (not A268)  and  a60929a );
 a60933a <=( (not A300)  and  (not A299) );
 a60936a <=( (not A302)  and  (not A301) );
 a60937a <=( a60936a  and  a60933a );
 a60938a <=( a60937a  and  a60930a );
 a60942a <=( (not A167)  and  A168 );
 a60943a <=( (not A170)  and  a60942a );
 a60946a <=( (not A201)  and  A166 );
 a60949a <=( A267  and  A202 );
 a60950a <=( a60949a  and  a60946a );
 a60951a <=( a60950a  and  a60943a );
 a60955a <=( (not A298)  and  (not A269) );
 a60956a <=( (not A268)  and  a60955a );
 a60959a <=( (not A300)  and  A299 );
 a60962a <=( (not A302)  and  (not A301) );
 a60963a <=( a60962a  and  a60959a );
 a60964a <=( a60963a  and  a60956a );
 a60968a <=( (not A167)  and  A168 );
 a60969a <=( (not A170)  and  a60968a );
 a60972a <=( (not A201)  and  A166 );
 a60975a <=( A267  and  A203 );
 a60976a <=( a60975a  and  a60972a );
 a60977a <=( a60976a  and  a60969a );
 a60981a <=( A298  and  (not A269) );
 a60982a <=( (not A268)  and  a60981a );
 a60985a <=( (not A300)  and  (not A299) );
 a60988a <=( (not A302)  and  (not A301) );
 a60989a <=( a60988a  and  a60985a );
 a60990a <=( a60989a  and  a60982a );
 a60994a <=( (not A167)  and  A168 );
 a60995a <=( (not A170)  and  a60994a );
 a60998a <=( (not A201)  and  A166 );
 a61001a <=( A267  and  A203 );
 a61002a <=( a61001a  and  a60998a );
 a61003a <=( a61002a  and  a60995a );
 a61007a <=( (not A298)  and  (not A269) );
 a61008a <=( (not A268)  and  a61007a );
 a61011a <=( (not A300)  and  A299 );
 a61014a <=( (not A302)  and  (not A301) );
 a61015a <=( a61014a  and  a61011a );
 a61016a <=( a61015a  and  a61008a );
 a61020a <=( (not A167)  and  A168 );
 a61021a <=( (not A170)  and  a61020a );
 a61024a <=( A199  and  A166 );
 a61027a <=( A267  and  A200 );
 a61028a <=( a61027a  and  a61024a );
 a61029a <=( a61028a  and  a61021a );
 a61033a <=( A298  and  (not A269) );
 a61034a <=( (not A268)  and  a61033a );
 a61037a <=( (not A300)  and  (not A299) );
 a61040a <=( (not A302)  and  (not A301) );
 a61041a <=( a61040a  and  a61037a );
 a61042a <=( a61041a  and  a61034a );
 a61046a <=( (not A167)  and  A168 );
 a61047a <=( (not A170)  and  a61046a );
 a61050a <=( A199  and  A166 );
 a61053a <=( A267  and  A200 );
 a61054a <=( a61053a  and  a61050a );
 a61055a <=( a61054a  and  a61047a );
 a61059a <=( (not A298)  and  (not A269) );
 a61060a <=( (not A268)  and  a61059a );
 a61063a <=( (not A300)  and  A299 );
 a61066a <=( (not A302)  and  (not A301) );
 a61067a <=( a61066a  and  a61063a );
 a61068a <=( a61067a  and  a61060a );
 a61072a <=( (not A167)  and  A168 );
 a61073a <=( (not A170)  and  a61072a );
 a61076a <=( (not A199)  and  A166 );
 a61079a <=( A201  and  A200 );
 a61080a <=( a61079a  and  a61076a );
 a61081a <=( a61080a  and  a61073a );
 a61085a <=( A266  and  (not A265) );
 a61086a <=( A202  and  a61085a );
 a61089a <=( A268  and  A267 );
 a61092a <=( A301  and  (not A300) );
 a61093a <=( a61092a  and  a61089a );
 a61094a <=( a61093a  and  a61086a );
 a61098a <=( (not A167)  and  A168 );
 a61099a <=( (not A170)  and  a61098a );
 a61102a <=( (not A199)  and  A166 );
 a61105a <=( A201  and  A200 );
 a61106a <=( a61105a  and  a61102a );
 a61107a <=( a61106a  and  a61099a );
 a61111a <=( A266  and  (not A265) );
 a61112a <=( A202  and  a61111a );
 a61115a <=( A268  and  A267 );
 a61118a <=( A302  and  (not A300) );
 a61119a <=( a61118a  and  a61115a );
 a61120a <=( a61119a  and  a61112a );
 a61124a <=( (not A167)  and  A168 );
 a61125a <=( (not A170)  and  a61124a );
 a61128a <=( (not A199)  and  A166 );
 a61131a <=( A201  and  A200 );
 a61132a <=( a61131a  and  a61128a );
 a61133a <=( a61132a  and  a61125a );
 a61137a <=( A266  and  (not A265) );
 a61138a <=( A202  and  a61137a );
 a61141a <=( A268  and  A267 );
 a61144a <=( A299  and  A298 );
 a61145a <=( a61144a  and  a61141a );
 a61146a <=( a61145a  and  a61138a );
 a61150a <=( (not A167)  and  A168 );
 a61151a <=( (not A170)  and  a61150a );
 a61154a <=( (not A199)  and  A166 );
 a61157a <=( A201  and  A200 );
 a61158a <=( a61157a  and  a61154a );
 a61159a <=( a61158a  and  a61151a );
 a61163a <=( A266  and  (not A265) );
 a61164a <=( A202  and  a61163a );
 a61167a <=( A268  and  A267 );
 a61170a <=( (not A299)  and  (not A298) );
 a61171a <=( a61170a  and  a61167a );
 a61172a <=( a61171a  and  a61164a );
 a61176a <=( (not A167)  and  A168 );
 a61177a <=( (not A170)  and  a61176a );
 a61180a <=( (not A199)  and  A166 );
 a61183a <=( A201  and  A200 );
 a61184a <=( a61183a  and  a61180a );
 a61185a <=( a61184a  and  a61177a );
 a61189a <=( A266  and  (not A265) );
 a61190a <=( A202  and  a61189a );
 a61193a <=( A269  and  A267 );
 a61196a <=( A301  and  (not A300) );
 a61197a <=( a61196a  and  a61193a );
 a61198a <=( a61197a  and  a61190a );
 a61202a <=( (not A167)  and  A168 );
 a61203a <=( (not A170)  and  a61202a );
 a61206a <=( (not A199)  and  A166 );
 a61209a <=( A201  and  A200 );
 a61210a <=( a61209a  and  a61206a );
 a61211a <=( a61210a  and  a61203a );
 a61215a <=( A266  and  (not A265) );
 a61216a <=( A202  and  a61215a );
 a61219a <=( A269  and  A267 );
 a61222a <=( A302  and  (not A300) );
 a61223a <=( a61222a  and  a61219a );
 a61224a <=( a61223a  and  a61216a );
 a61228a <=( (not A167)  and  A168 );
 a61229a <=( (not A170)  and  a61228a );
 a61232a <=( (not A199)  and  A166 );
 a61235a <=( A201  and  A200 );
 a61236a <=( a61235a  and  a61232a );
 a61237a <=( a61236a  and  a61229a );
 a61241a <=( A266  and  (not A265) );
 a61242a <=( A202  and  a61241a );
 a61245a <=( A269  and  A267 );
 a61248a <=( A299  and  A298 );
 a61249a <=( a61248a  and  a61245a );
 a61250a <=( a61249a  and  a61242a );
 a61254a <=( (not A167)  and  A168 );
 a61255a <=( (not A170)  and  a61254a );
 a61258a <=( (not A199)  and  A166 );
 a61261a <=( A201  and  A200 );
 a61262a <=( a61261a  and  a61258a );
 a61263a <=( a61262a  and  a61255a );
 a61267a <=( A266  and  (not A265) );
 a61268a <=( A202  and  a61267a );
 a61271a <=( A269  and  A267 );
 a61274a <=( (not A299)  and  (not A298) );
 a61275a <=( a61274a  and  a61271a );
 a61276a <=( a61275a  and  a61268a );
 a61280a <=( (not A167)  and  A168 );
 a61281a <=( (not A170)  and  a61280a );
 a61284a <=( (not A199)  and  A166 );
 a61287a <=( A201  and  A200 );
 a61288a <=( a61287a  and  a61284a );
 a61289a <=( a61288a  and  a61281a );
 a61293a <=( (not A266)  and  A265 );
 a61294a <=( A202  and  a61293a );
 a61297a <=( A268  and  A267 );
 a61300a <=( A301  and  (not A300) );
 a61301a <=( a61300a  and  a61297a );
 a61302a <=( a61301a  and  a61294a );
 a61306a <=( (not A167)  and  A168 );
 a61307a <=( (not A170)  and  a61306a );
 a61310a <=( (not A199)  and  A166 );
 a61313a <=( A201  and  A200 );
 a61314a <=( a61313a  and  a61310a );
 a61315a <=( a61314a  and  a61307a );
 a61319a <=( (not A266)  and  A265 );
 a61320a <=( A202  and  a61319a );
 a61323a <=( A268  and  A267 );
 a61326a <=( A302  and  (not A300) );
 a61327a <=( a61326a  and  a61323a );
 a61328a <=( a61327a  and  a61320a );
 a61332a <=( (not A167)  and  A168 );
 a61333a <=( (not A170)  and  a61332a );
 a61336a <=( (not A199)  and  A166 );
 a61339a <=( A201  and  A200 );
 a61340a <=( a61339a  and  a61336a );
 a61341a <=( a61340a  and  a61333a );
 a61345a <=( (not A266)  and  A265 );
 a61346a <=( A202  and  a61345a );
 a61349a <=( A268  and  A267 );
 a61352a <=( A299  and  A298 );
 a61353a <=( a61352a  and  a61349a );
 a61354a <=( a61353a  and  a61346a );
 a61358a <=( (not A167)  and  A168 );
 a61359a <=( (not A170)  and  a61358a );
 a61362a <=( (not A199)  and  A166 );
 a61365a <=( A201  and  A200 );
 a61366a <=( a61365a  and  a61362a );
 a61367a <=( a61366a  and  a61359a );
 a61371a <=( (not A266)  and  A265 );
 a61372a <=( A202  and  a61371a );
 a61375a <=( A268  and  A267 );
 a61378a <=( (not A299)  and  (not A298) );
 a61379a <=( a61378a  and  a61375a );
 a61380a <=( a61379a  and  a61372a );
 a61384a <=( (not A167)  and  A168 );
 a61385a <=( (not A170)  and  a61384a );
 a61388a <=( (not A199)  and  A166 );
 a61391a <=( A201  and  A200 );
 a61392a <=( a61391a  and  a61388a );
 a61393a <=( a61392a  and  a61385a );
 a61397a <=( (not A266)  and  A265 );
 a61398a <=( A202  and  a61397a );
 a61401a <=( A269  and  A267 );
 a61404a <=( A301  and  (not A300) );
 a61405a <=( a61404a  and  a61401a );
 a61406a <=( a61405a  and  a61398a );
 a61410a <=( (not A167)  and  A168 );
 a61411a <=( (not A170)  and  a61410a );
 a61414a <=( (not A199)  and  A166 );
 a61417a <=( A201  and  A200 );
 a61418a <=( a61417a  and  a61414a );
 a61419a <=( a61418a  and  a61411a );
 a61423a <=( (not A266)  and  A265 );
 a61424a <=( A202  and  a61423a );
 a61427a <=( A269  and  A267 );
 a61430a <=( A302  and  (not A300) );
 a61431a <=( a61430a  and  a61427a );
 a61432a <=( a61431a  and  a61424a );
 a61436a <=( (not A167)  and  A168 );
 a61437a <=( (not A170)  and  a61436a );
 a61440a <=( (not A199)  and  A166 );
 a61443a <=( A201  and  A200 );
 a61444a <=( a61443a  and  a61440a );
 a61445a <=( a61444a  and  a61437a );
 a61449a <=( (not A266)  and  A265 );
 a61450a <=( A202  and  a61449a );
 a61453a <=( A269  and  A267 );
 a61456a <=( A299  and  A298 );
 a61457a <=( a61456a  and  a61453a );
 a61458a <=( a61457a  and  a61450a );
 a61462a <=( (not A167)  and  A168 );
 a61463a <=( (not A170)  and  a61462a );
 a61466a <=( (not A199)  and  A166 );
 a61469a <=( A201  and  A200 );
 a61470a <=( a61469a  and  a61466a );
 a61471a <=( a61470a  and  a61463a );
 a61475a <=( (not A266)  and  A265 );
 a61476a <=( A202  and  a61475a );
 a61479a <=( A269  and  A267 );
 a61482a <=( (not A299)  and  (not A298) );
 a61483a <=( a61482a  and  a61479a );
 a61484a <=( a61483a  and  a61476a );
 a61488a <=( (not A167)  and  A168 );
 a61489a <=( (not A170)  and  a61488a );
 a61492a <=( (not A199)  and  A166 );
 a61495a <=( A201  and  A200 );
 a61496a <=( a61495a  and  a61492a );
 a61497a <=( a61496a  and  a61489a );
 a61501a <=( A266  and  (not A265) );
 a61502a <=( A203  and  a61501a );
 a61505a <=( A268  and  A267 );
 a61508a <=( A301  and  (not A300) );
 a61509a <=( a61508a  and  a61505a );
 a61510a <=( a61509a  and  a61502a );
 a61514a <=( (not A167)  and  A168 );
 a61515a <=( (not A170)  and  a61514a );
 a61518a <=( (not A199)  and  A166 );
 a61521a <=( A201  and  A200 );
 a61522a <=( a61521a  and  a61518a );
 a61523a <=( a61522a  and  a61515a );
 a61527a <=( A266  and  (not A265) );
 a61528a <=( A203  and  a61527a );
 a61531a <=( A268  and  A267 );
 a61534a <=( A302  and  (not A300) );
 a61535a <=( a61534a  and  a61531a );
 a61536a <=( a61535a  and  a61528a );
 a61540a <=( (not A167)  and  A168 );
 a61541a <=( (not A170)  and  a61540a );
 a61544a <=( (not A199)  and  A166 );
 a61547a <=( A201  and  A200 );
 a61548a <=( a61547a  and  a61544a );
 a61549a <=( a61548a  and  a61541a );
 a61553a <=( A266  and  (not A265) );
 a61554a <=( A203  and  a61553a );
 a61557a <=( A268  and  A267 );
 a61560a <=( A299  and  A298 );
 a61561a <=( a61560a  and  a61557a );
 a61562a <=( a61561a  and  a61554a );
 a61566a <=( (not A167)  and  A168 );
 a61567a <=( (not A170)  and  a61566a );
 a61570a <=( (not A199)  and  A166 );
 a61573a <=( A201  and  A200 );
 a61574a <=( a61573a  and  a61570a );
 a61575a <=( a61574a  and  a61567a );
 a61579a <=( A266  and  (not A265) );
 a61580a <=( A203  and  a61579a );
 a61583a <=( A268  and  A267 );
 a61586a <=( (not A299)  and  (not A298) );
 a61587a <=( a61586a  and  a61583a );
 a61588a <=( a61587a  and  a61580a );
 a61592a <=( (not A167)  and  A168 );
 a61593a <=( (not A170)  and  a61592a );
 a61596a <=( (not A199)  and  A166 );
 a61599a <=( A201  and  A200 );
 a61600a <=( a61599a  and  a61596a );
 a61601a <=( a61600a  and  a61593a );
 a61605a <=( A266  and  (not A265) );
 a61606a <=( A203  and  a61605a );
 a61609a <=( A269  and  A267 );
 a61612a <=( A301  and  (not A300) );
 a61613a <=( a61612a  and  a61609a );
 a61614a <=( a61613a  and  a61606a );
 a61618a <=( (not A167)  and  A168 );
 a61619a <=( (not A170)  and  a61618a );
 a61622a <=( (not A199)  and  A166 );
 a61625a <=( A201  and  A200 );
 a61626a <=( a61625a  and  a61622a );
 a61627a <=( a61626a  and  a61619a );
 a61631a <=( A266  and  (not A265) );
 a61632a <=( A203  and  a61631a );
 a61635a <=( A269  and  A267 );
 a61638a <=( A302  and  (not A300) );
 a61639a <=( a61638a  and  a61635a );
 a61640a <=( a61639a  and  a61632a );
 a61644a <=( (not A167)  and  A168 );
 a61645a <=( (not A170)  and  a61644a );
 a61648a <=( (not A199)  and  A166 );
 a61651a <=( A201  and  A200 );
 a61652a <=( a61651a  and  a61648a );
 a61653a <=( a61652a  and  a61645a );
 a61657a <=( A266  and  (not A265) );
 a61658a <=( A203  and  a61657a );
 a61661a <=( A269  and  A267 );
 a61664a <=( A299  and  A298 );
 a61665a <=( a61664a  and  a61661a );
 a61666a <=( a61665a  and  a61658a );
 a61670a <=( (not A167)  and  A168 );
 a61671a <=( (not A170)  and  a61670a );
 a61674a <=( (not A199)  and  A166 );
 a61677a <=( A201  and  A200 );
 a61678a <=( a61677a  and  a61674a );
 a61679a <=( a61678a  and  a61671a );
 a61683a <=( A266  and  (not A265) );
 a61684a <=( A203  and  a61683a );
 a61687a <=( A269  and  A267 );
 a61690a <=( (not A299)  and  (not A298) );
 a61691a <=( a61690a  and  a61687a );
 a61692a <=( a61691a  and  a61684a );
 a61696a <=( (not A167)  and  A168 );
 a61697a <=( (not A170)  and  a61696a );
 a61700a <=( (not A199)  and  A166 );
 a61703a <=( A201  and  A200 );
 a61704a <=( a61703a  and  a61700a );
 a61705a <=( a61704a  and  a61697a );
 a61709a <=( (not A266)  and  A265 );
 a61710a <=( A203  and  a61709a );
 a61713a <=( A268  and  A267 );
 a61716a <=( A301  and  (not A300) );
 a61717a <=( a61716a  and  a61713a );
 a61718a <=( a61717a  and  a61710a );
 a61722a <=( (not A167)  and  A168 );
 a61723a <=( (not A170)  and  a61722a );
 a61726a <=( (not A199)  and  A166 );
 a61729a <=( A201  and  A200 );
 a61730a <=( a61729a  and  a61726a );
 a61731a <=( a61730a  and  a61723a );
 a61735a <=( (not A266)  and  A265 );
 a61736a <=( A203  and  a61735a );
 a61739a <=( A268  and  A267 );
 a61742a <=( A302  and  (not A300) );
 a61743a <=( a61742a  and  a61739a );
 a61744a <=( a61743a  and  a61736a );
 a61748a <=( (not A167)  and  A168 );
 a61749a <=( (not A170)  and  a61748a );
 a61752a <=( (not A199)  and  A166 );
 a61755a <=( A201  and  A200 );
 a61756a <=( a61755a  and  a61752a );
 a61757a <=( a61756a  and  a61749a );
 a61761a <=( (not A266)  and  A265 );
 a61762a <=( A203  and  a61761a );
 a61765a <=( A268  and  A267 );
 a61768a <=( A299  and  A298 );
 a61769a <=( a61768a  and  a61765a );
 a61770a <=( a61769a  and  a61762a );
 a61774a <=( (not A167)  and  A168 );
 a61775a <=( (not A170)  and  a61774a );
 a61778a <=( (not A199)  and  A166 );
 a61781a <=( A201  and  A200 );
 a61782a <=( a61781a  and  a61778a );
 a61783a <=( a61782a  and  a61775a );
 a61787a <=( (not A266)  and  A265 );
 a61788a <=( A203  and  a61787a );
 a61791a <=( A268  and  A267 );
 a61794a <=( (not A299)  and  (not A298) );
 a61795a <=( a61794a  and  a61791a );
 a61796a <=( a61795a  and  a61788a );
 a61800a <=( (not A167)  and  A168 );
 a61801a <=( (not A170)  and  a61800a );
 a61804a <=( (not A199)  and  A166 );
 a61807a <=( A201  and  A200 );
 a61808a <=( a61807a  and  a61804a );
 a61809a <=( a61808a  and  a61801a );
 a61813a <=( (not A266)  and  A265 );
 a61814a <=( A203  and  a61813a );
 a61817a <=( A269  and  A267 );
 a61820a <=( A301  and  (not A300) );
 a61821a <=( a61820a  and  a61817a );
 a61822a <=( a61821a  and  a61814a );
 a61826a <=( (not A167)  and  A168 );
 a61827a <=( (not A170)  and  a61826a );
 a61830a <=( (not A199)  and  A166 );
 a61833a <=( A201  and  A200 );
 a61834a <=( a61833a  and  a61830a );
 a61835a <=( a61834a  and  a61827a );
 a61839a <=( (not A266)  and  A265 );
 a61840a <=( A203  and  a61839a );
 a61843a <=( A269  and  A267 );
 a61846a <=( A302  and  (not A300) );
 a61847a <=( a61846a  and  a61843a );
 a61848a <=( a61847a  and  a61840a );
 a61852a <=( (not A167)  and  A168 );
 a61853a <=( (not A170)  and  a61852a );
 a61856a <=( (not A199)  and  A166 );
 a61859a <=( A201  and  A200 );
 a61860a <=( a61859a  and  a61856a );
 a61861a <=( a61860a  and  a61853a );
 a61865a <=( (not A266)  and  A265 );
 a61866a <=( A203  and  a61865a );
 a61869a <=( A269  and  A267 );
 a61872a <=( A299  and  A298 );
 a61873a <=( a61872a  and  a61869a );
 a61874a <=( a61873a  and  a61866a );
 a61878a <=( (not A167)  and  A168 );
 a61879a <=( (not A170)  and  a61878a );
 a61882a <=( (not A199)  and  A166 );
 a61885a <=( A201  and  A200 );
 a61886a <=( a61885a  and  a61882a );
 a61887a <=( a61886a  and  a61879a );
 a61891a <=( (not A266)  and  A265 );
 a61892a <=( A203  and  a61891a );
 a61895a <=( A269  and  A267 );
 a61898a <=( (not A299)  and  (not A298) );
 a61899a <=( a61898a  and  a61895a );
 a61900a <=( a61899a  and  a61892a );
 a61904a <=( (not A167)  and  A168 );
 a61905a <=( (not A170)  and  a61904a );
 a61908a <=( A199  and  A166 );
 a61911a <=( A201  and  (not A200) );
 a61912a <=( a61911a  and  a61908a );
 a61913a <=( a61912a  and  a61905a );
 a61917a <=( A266  and  (not A265) );
 a61918a <=( A202  and  a61917a );
 a61921a <=( A268  and  A267 );
 a61924a <=( A301  and  (not A300) );
 a61925a <=( a61924a  and  a61921a );
 a61926a <=( a61925a  and  a61918a );
 a61930a <=( (not A167)  and  A168 );
 a61931a <=( (not A170)  and  a61930a );
 a61934a <=( A199  and  A166 );
 a61937a <=( A201  and  (not A200) );
 a61938a <=( a61937a  and  a61934a );
 a61939a <=( a61938a  and  a61931a );
 a61943a <=( A266  and  (not A265) );
 a61944a <=( A202  and  a61943a );
 a61947a <=( A268  and  A267 );
 a61950a <=( A302  and  (not A300) );
 a61951a <=( a61950a  and  a61947a );
 a61952a <=( a61951a  and  a61944a );
 a61956a <=( (not A167)  and  A168 );
 a61957a <=( (not A170)  and  a61956a );
 a61960a <=( A199  and  A166 );
 a61963a <=( A201  and  (not A200) );
 a61964a <=( a61963a  and  a61960a );
 a61965a <=( a61964a  and  a61957a );
 a61969a <=( A266  and  (not A265) );
 a61970a <=( A202  and  a61969a );
 a61973a <=( A268  and  A267 );
 a61976a <=( A299  and  A298 );
 a61977a <=( a61976a  and  a61973a );
 a61978a <=( a61977a  and  a61970a );
 a61982a <=( (not A167)  and  A168 );
 a61983a <=( (not A170)  and  a61982a );
 a61986a <=( A199  and  A166 );
 a61989a <=( A201  and  (not A200) );
 a61990a <=( a61989a  and  a61986a );
 a61991a <=( a61990a  and  a61983a );
 a61995a <=( A266  and  (not A265) );
 a61996a <=( A202  and  a61995a );
 a61999a <=( A268  and  A267 );
 a62002a <=( (not A299)  and  (not A298) );
 a62003a <=( a62002a  and  a61999a );
 a62004a <=( a62003a  and  a61996a );
 a62008a <=( (not A167)  and  A168 );
 a62009a <=( (not A170)  and  a62008a );
 a62012a <=( A199  and  A166 );
 a62015a <=( A201  and  (not A200) );
 a62016a <=( a62015a  and  a62012a );
 a62017a <=( a62016a  and  a62009a );
 a62021a <=( A266  and  (not A265) );
 a62022a <=( A202  and  a62021a );
 a62025a <=( A269  and  A267 );
 a62028a <=( A301  and  (not A300) );
 a62029a <=( a62028a  and  a62025a );
 a62030a <=( a62029a  and  a62022a );
 a62034a <=( (not A167)  and  A168 );
 a62035a <=( (not A170)  and  a62034a );
 a62038a <=( A199  and  A166 );
 a62041a <=( A201  and  (not A200) );
 a62042a <=( a62041a  and  a62038a );
 a62043a <=( a62042a  and  a62035a );
 a62047a <=( A266  and  (not A265) );
 a62048a <=( A202  and  a62047a );
 a62051a <=( A269  and  A267 );
 a62054a <=( A302  and  (not A300) );
 a62055a <=( a62054a  and  a62051a );
 a62056a <=( a62055a  and  a62048a );
 a62060a <=( (not A167)  and  A168 );
 a62061a <=( (not A170)  and  a62060a );
 a62064a <=( A199  and  A166 );
 a62067a <=( A201  and  (not A200) );
 a62068a <=( a62067a  and  a62064a );
 a62069a <=( a62068a  and  a62061a );
 a62073a <=( A266  and  (not A265) );
 a62074a <=( A202  and  a62073a );
 a62077a <=( A269  and  A267 );
 a62080a <=( A299  and  A298 );
 a62081a <=( a62080a  and  a62077a );
 a62082a <=( a62081a  and  a62074a );
 a62086a <=( (not A167)  and  A168 );
 a62087a <=( (not A170)  and  a62086a );
 a62090a <=( A199  and  A166 );
 a62093a <=( A201  and  (not A200) );
 a62094a <=( a62093a  and  a62090a );
 a62095a <=( a62094a  and  a62087a );
 a62099a <=( A266  and  (not A265) );
 a62100a <=( A202  and  a62099a );
 a62103a <=( A269  and  A267 );
 a62106a <=( (not A299)  and  (not A298) );
 a62107a <=( a62106a  and  a62103a );
 a62108a <=( a62107a  and  a62100a );
 a62112a <=( (not A167)  and  A168 );
 a62113a <=( (not A170)  and  a62112a );
 a62116a <=( A199  and  A166 );
 a62119a <=( A201  and  (not A200) );
 a62120a <=( a62119a  and  a62116a );
 a62121a <=( a62120a  and  a62113a );
 a62125a <=( (not A266)  and  A265 );
 a62126a <=( A202  and  a62125a );
 a62129a <=( A268  and  A267 );
 a62132a <=( A301  and  (not A300) );
 a62133a <=( a62132a  and  a62129a );
 a62134a <=( a62133a  and  a62126a );
 a62138a <=( (not A167)  and  A168 );
 a62139a <=( (not A170)  and  a62138a );
 a62142a <=( A199  and  A166 );
 a62145a <=( A201  and  (not A200) );
 a62146a <=( a62145a  and  a62142a );
 a62147a <=( a62146a  and  a62139a );
 a62151a <=( (not A266)  and  A265 );
 a62152a <=( A202  and  a62151a );
 a62155a <=( A268  and  A267 );
 a62158a <=( A302  and  (not A300) );
 a62159a <=( a62158a  and  a62155a );
 a62160a <=( a62159a  and  a62152a );
 a62164a <=( (not A167)  and  A168 );
 a62165a <=( (not A170)  and  a62164a );
 a62168a <=( A199  and  A166 );
 a62171a <=( A201  and  (not A200) );
 a62172a <=( a62171a  and  a62168a );
 a62173a <=( a62172a  and  a62165a );
 a62177a <=( (not A266)  and  A265 );
 a62178a <=( A202  and  a62177a );
 a62181a <=( A268  and  A267 );
 a62184a <=( A299  and  A298 );
 a62185a <=( a62184a  and  a62181a );
 a62186a <=( a62185a  and  a62178a );
 a62190a <=( (not A167)  and  A168 );
 a62191a <=( (not A170)  and  a62190a );
 a62194a <=( A199  and  A166 );
 a62197a <=( A201  and  (not A200) );
 a62198a <=( a62197a  and  a62194a );
 a62199a <=( a62198a  and  a62191a );
 a62203a <=( (not A266)  and  A265 );
 a62204a <=( A202  and  a62203a );
 a62207a <=( A268  and  A267 );
 a62210a <=( (not A299)  and  (not A298) );
 a62211a <=( a62210a  and  a62207a );
 a62212a <=( a62211a  and  a62204a );
 a62216a <=( (not A167)  and  A168 );
 a62217a <=( (not A170)  and  a62216a );
 a62220a <=( A199  and  A166 );
 a62223a <=( A201  and  (not A200) );
 a62224a <=( a62223a  and  a62220a );
 a62225a <=( a62224a  and  a62217a );
 a62229a <=( (not A266)  and  A265 );
 a62230a <=( A202  and  a62229a );
 a62233a <=( A269  and  A267 );
 a62236a <=( A301  and  (not A300) );
 a62237a <=( a62236a  and  a62233a );
 a62238a <=( a62237a  and  a62230a );
 a62242a <=( (not A167)  and  A168 );
 a62243a <=( (not A170)  and  a62242a );
 a62246a <=( A199  and  A166 );
 a62249a <=( A201  and  (not A200) );
 a62250a <=( a62249a  and  a62246a );
 a62251a <=( a62250a  and  a62243a );
 a62255a <=( (not A266)  and  A265 );
 a62256a <=( A202  and  a62255a );
 a62259a <=( A269  and  A267 );
 a62262a <=( A302  and  (not A300) );
 a62263a <=( a62262a  and  a62259a );
 a62264a <=( a62263a  and  a62256a );
 a62268a <=( (not A167)  and  A168 );
 a62269a <=( (not A170)  and  a62268a );
 a62272a <=( A199  and  A166 );
 a62275a <=( A201  and  (not A200) );
 a62276a <=( a62275a  and  a62272a );
 a62277a <=( a62276a  and  a62269a );
 a62281a <=( (not A266)  and  A265 );
 a62282a <=( A202  and  a62281a );
 a62285a <=( A269  and  A267 );
 a62288a <=( A299  and  A298 );
 a62289a <=( a62288a  and  a62285a );
 a62290a <=( a62289a  and  a62282a );
 a62294a <=( (not A167)  and  A168 );
 a62295a <=( (not A170)  and  a62294a );
 a62298a <=( A199  and  A166 );
 a62301a <=( A201  and  (not A200) );
 a62302a <=( a62301a  and  a62298a );
 a62303a <=( a62302a  and  a62295a );
 a62307a <=( (not A266)  and  A265 );
 a62308a <=( A202  and  a62307a );
 a62311a <=( A269  and  A267 );
 a62314a <=( (not A299)  and  (not A298) );
 a62315a <=( a62314a  and  a62311a );
 a62316a <=( a62315a  and  a62308a );
 a62320a <=( (not A167)  and  A168 );
 a62321a <=( (not A170)  and  a62320a );
 a62324a <=( A199  and  A166 );
 a62327a <=( A201  and  (not A200) );
 a62328a <=( a62327a  and  a62324a );
 a62329a <=( a62328a  and  a62321a );
 a62333a <=( A266  and  (not A265) );
 a62334a <=( A203  and  a62333a );
 a62337a <=( A268  and  A267 );
 a62340a <=( A301  and  (not A300) );
 a62341a <=( a62340a  and  a62337a );
 a62342a <=( a62341a  and  a62334a );
 a62346a <=( (not A167)  and  A168 );
 a62347a <=( (not A170)  and  a62346a );
 a62350a <=( A199  and  A166 );
 a62353a <=( A201  and  (not A200) );
 a62354a <=( a62353a  and  a62350a );
 a62355a <=( a62354a  and  a62347a );
 a62359a <=( A266  and  (not A265) );
 a62360a <=( A203  and  a62359a );
 a62363a <=( A268  and  A267 );
 a62366a <=( A302  and  (not A300) );
 a62367a <=( a62366a  and  a62363a );
 a62368a <=( a62367a  and  a62360a );
 a62372a <=( (not A167)  and  A168 );
 a62373a <=( (not A170)  and  a62372a );
 a62376a <=( A199  and  A166 );
 a62379a <=( A201  and  (not A200) );
 a62380a <=( a62379a  and  a62376a );
 a62381a <=( a62380a  and  a62373a );
 a62385a <=( A266  and  (not A265) );
 a62386a <=( A203  and  a62385a );
 a62389a <=( A268  and  A267 );
 a62392a <=( A299  and  A298 );
 a62393a <=( a62392a  and  a62389a );
 a62394a <=( a62393a  and  a62386a );
 a62398a <=( (not A167)  and  A168 );
 a62399a <=( (not A170)  and  a62398a );
 a62402a <=( A199  and  A166 );
 a62405a <=( A201  and  (not A200) );
 a62406a <=( a62405a  and  a62402a );
 a62407a <=( a62406a  and  a62399a );
 a62411a <=( A266  and  (not A265) );
 a62412a <=( A203  and  a62411a );
 a62415a <=( A268  and  A267 );
 a62418a <=( (not A299)  and  (not A298) );
 a62419a <=( a62418a  and  a62415a );
 a62420a <=( a62419a  and  a62412a );
 a62424a <=( (not A167)  and  A168 );
 a62425a <=( (not A170)  and  a62424a );
 a62428a <=( A199  and  A166 );
 a62431a <=( A201  and  (not A200) );
 a62432a <=( a62431a  and  a62428a );
 a62433a <=( a62432a  and  a62425a );
 a62437a <=( A266  and  (not A265) );
 a62438a <=( A203  and  a62437a );
 a62441a <=( A269  and  A267 );
 a62444a <=( A301  and  (not A300) );
 a62445a <=( a62444a  and  a62441a );
 a62446a <=( a62445a  and  a62438a );
 a62450a <=( (not A167)  and  A168 );
 a62451a <=( (not A170)  and  a62450a );
 a62454a <=( A199  and  A166 );
 a62457a <=( A201  and  (not A200) );
 a62458a <=( a62457a  and  a62454a );
 a62459a <=( a62458a  and  a62451a );
 a62463a <=( A266  and  (not A265) );
 a62464a <=( A203  and  a62463a );
 a62467a <=( A269  and  A267 );
 a62470a <=( A302  and  (not A300) );
 a62471a <=( a62470a  and  a62467a );
 a62472a <=( a62471a  and  a62464a );
 a62476a <=( (not A167)  and  A168 );
 a62477a <=( (not A170)  and  a62476a );
 a62480a <=( A199  and  A166 );
 a62483a <=( A201  and  (not A200) );
 a62484a <=( a62483a  and  a62480a );
 a62485a <=( a62484a  and  a62477a );
 a62489a <=( A266  and  (not A265) );
 a62490a <=( A203  and  a62489a );
 a62493a <=( A269  and  A267 );
 a62496a <=( A299  and  A298 );
 a62497a <=( a62496a  and  a62493a );
 a62498a <=( a62497a  and  a62490a );
 a62502a <=( (not A167)  and  A168 );
 a62503a <=( (not A170)  and  a62502a );
 a62506a <=( A199  and  A166 );
 a62509a <=( A201  and  (not A200) );
 a62510a <=( a62509a  and  a62506a );
 a62511a <=( a62510a  and  a62503a );
 a62515a <=( A266  and  (not A265) );
 a62516a <=( A203  and  a62515a );
 a62519a <=( A269  and  A267 );
 a62522a <=( (not A299)  and  (not A298) );
 a62523a <=( a62522a  and  a62519a );
 a62524a <=( a62523a  and  a62516a );
 a62528a <=( (not A167)  and  A168 );
 a62529a <=( (not A170)  and  a62528a );
 a62532a <=( A199  and  A166 );
 a62535a <=( A201  and  (not A200) );
 a62536a <=( a62535a  and  a62532a );
 a62537a <=( a62536a  and  a62529a );
 a62541a <=( (not A266)  and  A265 );
 a62542a <=( A203  and  a62541a );
 a62545a <=( A268  and  A267 );
 a62548a <=( A301  and  (not A300) );
 a62549a <=( a62548a  and  a62545a );
 a62550a <=( a62549a  and  a62542a );
 a62554a <=( (not A167)  and  A168 );
 a62555a <=( (not A170)  and  a62554a );
 a62558a <=( A199  and  A166 );
 a62561a <=( A201  and  (not A200) );
 a62562a <=( a62561a  and  a62558a );
 a62563a <=( a62562a  and  a62555a );
 a62567a <=( (not A266)  and  A265 );
 a62568a <=( A203  and  a62567a );
 a62571a <=( A268  and  A267 );
 a62574a <=( A302  and  (not A300) );
 a62575a <=( a62574a  and  a62571a );
 a62576a <=( a62575a  and  a62568a );
 a62580a <=( (not A167)  and  A168 );
 a62581a <=( (not A170)  and  a62580a );
 a62584a <=( A199  and  A166 );
 a62587a <=( A201  and  (not A200) );
 a62588a <=( a62587a  and  a62584a );
 a62589a <=( a62588a  and  a62581a );
 a62593a <=( (not A266)  and  A265 );
 a62594a <=( A203  and  a62593a );
 a62597a <=( A268  and  A267 );
 a62600a <=( A299  and  A298 );
 a62601a <=( a62600a  and  a62597a );
 a62602a <=( a62601a  and  a62594a );
 a62606a <=( (not A167)  and  A168 );
 a62607a <=( (not A170)  and  a62606a );
 a62610a <=( A199  and  A166 );
 a62613a <=( A201  and  (not A200) );
 a62614a <=( a62613a  and  a62610a );
 a62615a <=( a62614a  and  a62607a );
 a62619a <=( (not A266)  and  A265 );
 a62620a <=( A203  and  a62619a );
 a62623a <=( A268  and  A267 );
 a62626a <=( (not A299)  and  (not A298) );
 a62627a <=( a62626a  and  a62623a );
 a62628a <=( a62627a  and  a62620a );
 a62632a <=( (not A167)  and  A168 );
 a62633a <=( (not A170)  and  a62632a );
 a62636a <=( A199  and  A166 );
 a62639a <=( A201  and  (not A200) );
 a62640a <=( a62639a  and  a62636a );
 a62641a <=( a62640a  and  a62633a );
 a62645a <=( (not A266)  and  A265 );
 a62646a <=( A203  and  a62645a );
 a62649a <=( A269  and  A267 );
 a62652a <=( A301  and  (not A300) );
 a62653a <=( a62652a  and  a62649a );
 a62654a <=( a62653a  and  a62646a );
 a62658a <=( (not A167)  and  A168 );
 a62659a <=( (not A170)  and  a62658a );
 a62662a <=( A199  and  A166 );
 a62665a <=( A201  and  (not A200) );
 a62666a <=( a62665a  and  a62662a );
 a62667a <=( a62666a  and  a62659a );
 a62671a <=( (not A266)  and  A265 );
 a62672a <=( A203  and  a62671a );
 a62675a <=( A269  and  A267 );
 a62678a <=( A302  and  (not A300) );
 a62679a <=( a62678a  and  a62675a );
 a62680a <=( a62679a  and  a62672a );
 a62684a <=( (not A167)  and  A168 );
 a62685a <=( (not A170)  and  a62684a );
 a62688a <=( A199  and  A166 );
 a62691a <=( A201  and  (not A200) );
 a62692a <=( a62691a  and  a62688a );
 a62693a <=( a62692a  and  a62685a );
 a62697a <=( (not A266)  and  A265 );
 a62698a <=( A203  and  a62697a );
 a62701a <=( A269  and  A267 );
 a62704a <=( A299  and  A298 );
 a62705a <=( a62704a  and  a62701a );
 a62706a <=( a62705a  and  a62698a );
 a62710a <=( (not A167)  and  A168 );
 a62711a <=( (not A170)  and  a62710a );
 a62714a <=( A199  and  A166 );
 a62717a <=( A201  and  (not A200) );
 a62718a <=( a62717a  and  a62714a );
 a62719a <=( a62718a  and  a62711a );
 a62723a <=( (not A266)  and  A265 );
 a62724a <=( A203  and  a62723a );
 a62727a <=( A269  and  A267 );
 a62730a <=( (not A299)  and  (not A298) );
 a62731a <=( a62730a  and  a62727a );
 a62732a <=( a62731a  and  a62724a );
 a62736a <=( (not A167)  and  A168 );
 a62737a <=( (not A170)  and  a62736a );
 a62740a <=( (not A199)  and  A166 );
 a62743a <=( A267  and  (not A200) );
 a62744a <=( a62743a  and  a62740a );
 a62745a <=( a62744a  and  a62737a );
 a62749a <=( A298  and  (not A269) );
 a62750a <=( (not A268)  and  a62749a );
 a62753a <=( (not A300)  and  (not A299) );
 a62756a <=( (not A302)  and  (not A301) );
 a62757a <=( a62756a  and  a62753a );
 a62758a <=( a62757a  and  a62750a );
 a62762a <=( (not A167)  and  A168 );
 a62763a <=( (not A170)  and  a62762a );
 a62766a <=( (not A199)  and  A166 );
 a62769a <=( A267  and  (not A200) );
 a62770a <=( a62769a  and  a62766a );
 a62771a <=( a62770a  and  a62763a );
 a62775a <=( (not A298)  and  (not A269) );
 a62776a <=( (not A268)  and  a62775a );
 a62779a <=( (not A300)  and  A299 );
 a62782a <=( (not A302)  and  (not A301) );
 a62783a <=( a62782a  and  a62779a );
 a62784a <=( a62783a  and  a62776a );
 a62788a <=( (not A199)  and  (not A168) );
 a62789a <=( (not A170)  and  a62788a );
 a62792a <=( A201  and  A200 );
 a62795a <=( A267  and  A202 );
 a62796a <=( a62795a  and  a62792a );
 a62797a <=( a62796a  and  a62789a );
 a62801a <=( A298  and  (not A269) );
 a62802a <=( (not A268)  and  a62801a );
 a62805a <=( (not A300)  and  (not A299) );
 a62808a <=( (not A302)  and  (not A301) );
 a62809a <=( a62808a  and  a62805a );
 a62810a <=( a62809a  and  a62802a );
 a62814a <=( (not A199)  and  (not A168) );
 a62815a <=( (not A170)  and  a62814a );
 a62818a <=( A201  and  A200 );
 a62821a <=( A267  and  A202 );
 a62822a <=( a62821a  and  a62818a );
 a62823a <=( a62822a  and  a62815a );
 a62827a <=( (not A298)  and  (not A269) );
 a62828a <=( (not A268)  and  a62827a );
 a62831a <=( (not A300)  and  A299 );
 a62834a <=( (not A302)  and  (not A301) );
 a62835a <=( a62834a  and  a62831a );
 a62836a <=( a62835a  and  a62828a );
 a62840a <=( (not A199)  and  (not A168) );
 a62841a <=( (not A170)  and  a62840a );
 a62844a <=( A201  and  A200 );
 a62847a <=( A267  and  A203 );
 a62848a <=( a62847a  and  a62844a );
 a62849a <=( a62848a  and  a62841a );
 a62853a <=( A298  and  (not A269) );
 a62854a <=( (not A268)  and  a62853a );
 a62857a <=( (not A300)  and  (not A299) );
 a62860a <=( (not A302)  and  (not A301) );
 a62861a <=( a62860a  and  a62857a );
 a62862a <=( a62861a  and  a62854a );
 a62866a <=( (not A199)  and  (not A168) );
 a62867a <=( (not A170)  and  a62866a );
 a62870a <=( A201  and  A200 );
 a62873a <=( A267  and  A203 );
 a62874a <=( a62873a  and  a62870a );
 a62875a <=( a62874a  and  a62867a );
 a62879a <=( (not A298)  and  (not A269) );
 a62880a <=( (not A268)  and  a62879a );
 a62883a <=( (not A300)  and  A299 );
 a62886a <=( (not A302)  and  (not A301) );
 a62887a <=( a62886a  and  a62883a );
 a62888a <=( a62887a  and  a62880a );
 a62892a <=( (not A199)  and  (not A168) );
 a62893a <=( (not A170)  and  a62892a );
 a62896a <=( (not A201)  and  A200 );
 a62899a <=( (not A203)  and  (not A202) );
 a62900a <=( a62899a  and  a62896a );
 a62901a <=( a62900a  and  a62893a );
 a62905a <=( (not A269)  and  (not A268) );
 a62906a <=( A267  and  a62905a );
 a62909a <=( (not A299)  and  A298 );
 a62912a <=( A301  and  A300 );
 a62913a <=( a62912a  and  a62909a );
 a62914a <=( a62913a  and  a62906a );
 a62918a <=( (not A199)  and  (not A168) );
 a62919a <=( (not A170)  and  a62918a );
 a62922a <=( (not A201)  and  A200 );
 a62925a <=( (not A203)  and  (not A202) );
 a62926a <=( a62925a  and  a62922a );
 a62927a <=( a62926a  and  a62919a );
 a62931a <=( (not A269)  and  (not A268) );
 a62932a <=( A267  and  a62931a );
 a62935a <=( (not A299)  and  A298 );
 a62938a <=( A302  and  A300 );
 a62939a <=( a62938a  and  a62935a );
 a62940a <=( a62939a  and  a62932a );
 a62944a <=( (not A199)  and  (not A168) );
 a62945a <=( (not A170)  and  a62944a );
 a62948a <=( (not A201)  and  A200 );
 a62951a <=( (not A203)  and  (not A202) );
 a62952a <=( a62951a  and  a62948a );
 a62953a <=( a62952a  and  a62945a );
 a62957a <=( (not A269)  and  (not A268) );
 a62958a <=( A267  and  a62957a );
 a62961a <=( A299  and  (not A298) );
 a62964a <=( A301  and  A300 );
 a62965a <=( a62964a  and  a62961a );
 a62966a <=( a62965a  and  a62958a );
 a62970a <=( (not A199)  and  (not A168) );
 a62971a <=( (not A170)  and  a62970a );
 a62974a <=( (not A201)  and  A200 );
 a62977a <=( (not A203)  and  (not A202) );
 a62978a <=( a62977a  and  a62974a );
 a62979a <=( a62978a  and  a62971a );
 a62983a <=( (not A269)  and  (not A268) );
 a62984a <=( A267  and  a62983a );
 a62987a <=( A299  and  (not A298) );
 a62990a <=( A302  and  A300 );
 a62991a <=( a62990a  and  a62987a );
 a62992a <=( a62991a  and  a62984a );
 a62996a <=( (not A199)  and  (not A168) );
 a62997a <=( (not A170)  and  a62996a );
 a63000a <=( (not A201)  and  A200 );
 a63003a <=( (not A203)  and  (not A202) );
 a63004a <=( a63003a  and  a63000a );
 a63005a <=( a63004a  and  a62997a );
 a63009a <=( A298  and  A268 );
 a63010a <=( (not A267)  and  a63009a );
 a63013a <=( (not A300)  and  (not A299) );
 a63016a <=( (not A302)  and  (not A301) );
 a63017a <=( a63016a  and  a63013a );
 a63018a <=( a63017a  and  a63010a );
 a63022a <=( (not A199)  and  (not A168) );
 a63023a <=( (not A170)  and  a63022a );
 a63026a <=( (not A201)  and  A200 );
 a63029a <=( (not A203)  and  (not A202) );
 a63030a <=( a63029a  and  a63026a );
 a63031a <=( a63030a  and  a63023a );
 a63035a <=( (not A298)  and  A268 );
 a63036a <=( (not A267)  and  a63035a );
 a63039a <=( (not A300)  and  A299 );
 a63042a <=( (not A302)  and  (not A301) );
 a63043a <=( a63042a  and  a63039a );
 a63044a <=( a63043a  and  a63036a );
 a63048a <=( (not A199)  and  (not A168) );
 a63049a <=( (not A170)  and  a63048a );
 a63052a <=( (not A201)  and  A200 );
 a63055a <=( (not A203)  and  (not A202) );
 a63056a <=( a63055a  and  a63052a );
 a63057a <=( a63056a  and  a63049a );
 a63061a <=( A298  and  A269 );
 a63062a <=( (not A267)  and  a63061a );
 a63065a <=( (not A300)  and  (not A299) );
 a63068a <=( (not A302)  and  (not A301) );
 a63069a <=( a63068a  and  a63065a );
 a63070a <=( a63069a  and  a63062a );
 a63074a <=( (not A199)  and  (not A168) );
 a63075a <=( (not A170)  and  a63074a );
 a63078a <=( (not A201)  and  A200 );
 a63081a <=( (not A203)  and  (not A202) );
 a63082a <=( a63081a  and  a63078a );
 a63083a <=( a63082a  and  a63075a );
 a63087a <=( (not A298)  and  A269 );
 a63088a <=( (not A267)  and  a63087a );
 a63091a <=( (not A300)  and  A299 );
 a63094a <=( (not A302)  and  (not A301) );
 a63095a <=( a63094a  and  a63091a );
 a63096a <=( a63095a  and  a63088a );
 a63100a <=( (not A199)  and  (not A168) );
 a63101a <=( (not A170)  and  a63100a );
 a63104a <=( (not A201)  and  A200 );
 a63107a <=( (not A203)  and  (not A202) );
 a63108a <=( a63107a  and  a63104a );
 a63109a <=( a63108a  and  a63101a );
 a63113a <=( A298  and  A266 );
 a63114a <=( A265  and  a63113a );
 a63117a <=( (not A300)  and  (not A299) );
 a63120a <=( (not A302)  and  (not A301) );
 a63121a <=( a63120a  and  a63117a );
 a63122a <=( a63121a  and  a63114a );
 a63126a <=( (not A199)  and  (not A168) );
 a63127a <=( (not A170)  and  a63126a );
 a63130a <=( (not A201)  and  A200 );
 a63133a <=( (not A203)  and  (not A202) );
 a63134a <=( a63133a  and  a63130a );
 a63135a <=( a63134a  and  a63127a );
 a63139a <=( (not A298)  and  A266 );
 a63140a <=( A265  and  a63139a );
 a63143a <=( (not A300)  and  A299 );
 a63146a <=( (not A302)  and  (not A301) );
 a63147a <=( a63146a  and  a63143a );
 a63148a <=( a63147a  and  a63140a );
 a63152a <=( (not A199)  and  (not A168) );
 a63153a <=( (not A170)  and  a63152a );
 a63156a <=( (not A201)  and  A200 );
 a63159a <=( (not A203)  and  (not A202) );
 a63160a <=( a63159a  and  a63156a );
 a63161a <=( a63160a  and  a63153a );
 a63165a <=( A298  and  (not A266) );
 a63166a <=( (not A265)  and  a63165a );
 a63169a <=( (not A300)  and  (not A299) );
 a63172a <=( (not A302)  and  (not A301) );
 a63173a <=( a63172a  and  a63169a );
 a63174a <=( a63173a  and  a63166a );
 a63178a <=( (not A199)  and  (not A168) );
 a63179a <=( (not A170)  and  a63178a );
 a63182a <=( (not A201)  and  A200 );
 a63185a <=( (not A203)  and  (not A202) );
 a63186a <=( a63185a  and  a63182a );
 a63187a <=( a63186a  and  a63179a );
 a63191a <=( (not A298)  and  (not A266) );
 a63192a <=( (not A265)  and  a63191a );
 a63195a <=( (not A300)  and  A299 );
 a63198a <=( (not A302)  and  (not A301) );
 a63199a <=( a63198a  and  a63195a );
 a63200a <=( a63199a  and  a63192a );
 a63204a <=( A199  and  (not A168) );
 a63205a <=( (not A170)  and  a63204a );
 a63208a <=( A201  and  (not A200) );
 a63211a <=( A267  and  A202 );
 a63212a <=( a63211a  and  a63208a );
 a63213a <=( a63212a  and  a63205a );
 a63217a <=( A298  and  (not A269) );
 a63218a <=( (not A268)  and  a63217a );
 a63221a <=( (not A300)  and  (not A299) );
 a63224a <=( (not A302)  and  (not A301) );
 a63225a <=( a63224a  and  a63221a );
 a63226a <=( a63225a  and  a63218a );
 a63230a <=( A199  and  (not A168) );
 a63231a <=( (not A170)  and  a63230a );
 a63234a <=( A201  and  (not A200) );
 a63237a <=( A267  and  A202 );
 a63238a <=( a63237a  and  a63234a );
 a63239a <=( a63238a  and  a63231a );
 a63243a <=( (not A298)  and  (not A269) );
 a63244a <=( (not A268)  and  a63243a );
 a63247a <=( (not A300)  and  A299 );
 a63250a <=( (not A302)  and  (not A301) );
 a63251a <=( a63250a  and  a63247a );
 a63252a <=( a63251a  and  a63244a );
 a63256a <=( A199  and  (not A168) );
 a63257a <=( (not A170)  and  a63256a );
 a63260a <=( A201  and  (not A200) );
 a63263a <=( A267  and  A203 );
 a63264a <=( a63263a  and  a63260a );
 a63265a <=( a63264a  and  a63257a );
 a63269a <=( A298  and  (not A269) );
 a63270a <=( (not A268)  and  a63269a );
 a63273a <=( (not A300)  and  (not A299) );
 a63276a <=( (not A302)  and  (not A301) );
 a63277a <=( a63276a  and  a63273a );
 a63278a <=( a63277a  and  a63270a );
 a63282a <=( A199  and  (not A168) );
 a63283a <=( (not A170)  and  a63282a );
 a63286a <=( A201  and  (not A200) );
 a63289a <=( A267  and  A203 );
 a63290a <=( a63289a  and  a63286a );
 a63291a <=( a63290a  and  a63283a );
 a63295a <=( (not A298)  and  (not A269) );
 a63296a <=( (not A268)  and  a63295a );
 a63299a <=( (not A300)  and  A299 );
 a63302a <=( (not A302)  and  (not A301) );
 a63303a <=( a63302a  and  a63299a );
 a63304a <=( a63303a  and  a63296a );
 a63308a <=( A199  and  (not A168) );
 a63309a <=( (not A170)  and  a63308a );
 a63312a <=( (not A201)  and  (not A200) );
 a63315a <=( (not A203)  and  (not A202) );
 a63316a <=( a63315a  and  a63312a );
 a63317a <=( a63316a  and  a63309a );
 a63321a <=( (not A269)  and  (not A268) );
 a63322a <=( A267  and  a63321a );
 a63325a <=( (not A299)  and  A298 );
 a63328a <=( A301  and  A300 );
 a63329a <=( a63328a  and  a63325a );
 a63330a <=( a63329a  and  a63322a );
 a63334a <=( A199  and  (not A168) );
 a63335a <=( (not A170)  and  a63334a );
 a63338a <=( (not A201)  and  (not A200) );
 a63341a <=( (not A203)  and  (not A202) );
 a63342a <=( a63341a  and  a63338a );
 a63343a <=( a63342a  and  a63335a );
 a63347a <=( (not A269)  and  (not A268) );
 a63348a <=( A267  and  a63347a );
 a63351a <=( (not A299)  and  A298 );
 a63354a <=( A302  and  A300 );
 a63355a <=( a63354a  and  a63351a );
 a63356a <=( a63355a  and  a63348a );
 a63360a <=( A199  and  (not A168) );
 a63361a <=( (not A170)  and  a63360a );
 a63364a <=( (not A201)  and  (not A200) );
 a63367a <=( (not A203)  and  (not A202) );
 a63368a <=( a63367a  and  a63364a );
 a63369a <=( a63368a  and  a63361a );
 a63373a <=( (not A269)  and  (not A268) );
 a63374a <=( A267  and  a63373a );
 a63377a <=( A299  and  (not A298) );
 a63380a <=( A301  and  A300 );
 a63381a <=( a63380a  and  a63377a );
 a63382a <=( a63381a  and  a63374a );
 a63386a <=( A199  and  (not A168) );
 a63387a <=( (not A170)  and  a63386a );
 a63390a <=( (not A201)  and  (not A200) );
 a63393a <=( (not A203)  and  (not A202) );
 a63394a <=( a63393a  and  a63390a );
 a63395a <=( a63394a  and  a63387a );
 a63399a <=( (not A269)  and  (not A268) );
 a63400a <=( A267  and  a63399a );
 a63403a <=( A299  and  (not A298) );
 a63406a <=( A302  and  A300 );
 a63407a <=( a63406a  and  a63403a );
 a63408a <=( a63407a  and  a63400a );
 a63412a <=( A199  and  (not A168) );
 a63413a <=( (not A170)  and  a63412a );
 a63416a <=( (not A201)  and  (not A200) );
 a63419a <=( (not A203)  and  (not A202) );
 a63420a <=( a63419a  and  a63416a );
 a63421a <=( a63420a  and  a63413a );
 a63425a <=( A298  and  A268 );
 a63426a <=( (not A267)  and  a63425a );
 a63429a <=( (not A300)  and  (not A299) );
 a63432a <=( (not A302)  and  (not A301) );
 a63433a <=( a63432a  and  a63429a );
 a63434a <=( a63433a  and  a63426a );
 a63438a <=( A199  and  (not A168) );
 a63439a <=( (not A170)  and  a63438a );
 a63442a <=( (not A201)  and  (not A200) );
 a63445a <=( (not A203)  and  (not A202) );
 a63446a <=( a63445a  and  a63442a );
 a63447a <=( a63446a  and  a63439a );
 a63451a <=( (not A298)  and  A268 );
 a63452a <=( (not A267)  and  a63451a );
 a63455a <=( (not A300)  and  A299 );
 a63458a <=( (not A302)  and  (not A301) );
 a63459a <=( a63458a  and  a63455a );
 a63460a <=( a63459a  and  a63452a );
 a63464a <=( A199  and  (not A168) );
 a63465a <=( (not A170)  and  a63464a );
 a63468a <=( (not A201)  and  (not A200) );
 a63471a <=( (not A203)  and  (not A202) );
 a63472a <=( a63471a  and  a63468a );
 a63473a <=( a63472a  and  a63465a );
 a63477a <=( A298  and  A269 );
 a63478a <=( (not A267)  and  a63477a );
 a63481a <=( (not A300)  and  (not A299) );
 a63484a <=( (not A302)  and  (not A301) );
 a63485a <=( a63484a  and  a63481a );
 a63486a <=( a63485a  and  a63478a );
 a63490a <=( A199  and  (not A168) );
 a63491a <=( (not A170)  and  a63490a );
 a63494a <=( (not A201)  and  (not A200) );
 a63497a <=( (not A203)  and  (not A202) );
 a63498a <=( a63497a  and  a63494a );
 a63499a <=( a63498a  and  a63491a );
 a63503a <=( (not A298)  and  A269 );
 a63504a <=( (not A267)  and  a63503a );
 a63507a <=( (not A300)  and  A299 );
 a63510a <=( (not A302)  and  (not A301) );
 a63511a <=( a63510a  and  a63507a );
 a63512a <=( a63511a  and  a63504a );
 a63516a <=( A199  and  (not A168) );
 a63517a <=( (not A170)  and  a63516a );
 a63520a <=( (not A201)  and  (not A200) );
 a63523a <=( (not A203)  and  (not A202) );
 a63524a <=( a63523a  and  a63520a );
 a63525a <=( a63524a  and  a63517a );
 a63529a <=( A298  and  A266 );
 a63530a <=( A265  and  a63529a );
 a63533a <=( (not A300)  and  (not A299) );
 a63536a <=( (not A302)  and  (not A301) );
 a63537a <=( a63536a  and  a63533a );
 a63538a <=( a63537a  and  a63530a );
 a63542a <=( A199  and  (not A168) );
 a63543a <=( (not A170)  and  a63542a );
 a63546a <=( (not A201)  and  (not A200) );
 a63549a <=( (not A203)  and  (not A202) );
 a63550a <=( a63549a  and  a63546a );
 a63551a <=( a63550a  and  a63543a );
 a63555a <=( (not A298)  and  A266 );
 a63556a <=( A265  and  a63555a );
 a63559a <=( (not A300)  and  A299 );
 a63562a <=( (not A302)  and  (not A301) );
 a63563a <=( a63562a  and  a63559a );
 a63564a <=( a63563a  and  a63556a );
 a63568a <=( A199  and  (not A168) );
 a63569a <=( (not A170)  and  a63568a );
 a63572a <=( (not A201)  and  (not A200) );
 a63575a <=( (not A203)  and  (not A202) );
 a63576a <=( a63575a  and  a63572a );
 a63577a <=( a63576a  and  a63569a );
 a63581a <=( A298  and  (not A266) );
 a63582a <=( (not A265)  and  a63581a );
 a63585a <=( (not A300)  and  (not A299) );
 a63588a <=( (not A302)  and  (not A301) );
 a63589a <=( a63588a  and  a63585a );
 a63590a <=( a63589a  and  a63582a );
 a63594a <=( A199  and  (not A168) );
 a63595a <=( (not A170)  and  a63594a );
 a63598a <=( (not A201)  and  (not A200) );
 a63601a <=( (not A203)  and  (not A202) );
 a63602a <=( a63601a  and  a63598a );
 a63603a <=( a63602a  and  a63595a );
 a63607a <=( (not A298)  and  (not A266) );
 a63608a <=( (not A265)  and  a63607a );
 a63611a <=( (not A300)  and  A299 );
 a63614a <=( (not A302)  and  (not A301) );
 a63615a <=( a63614a  and  a63611a );
 a63616a <=( a63615a  and  a63608a );
 a63620a <=( A167  and  A168 );
 a63621a <=( A169  and  a63620a );
 a63624a <=( A201  and  (not A166) );
 a63627a <=( (not A203)  and  (not A202) );
 a63628a <=( a63627a  and  a63624a );
 a63629a <=( a63628a  and  a63621a );
 a63633a <=( (not A269)  and  (not A268) );
 a63634a <=( A267  and  a63633a );
 a63637a <=( (not A299)  and  A298 );
 a63640a <=( A301  and  A300 );
 a63641a <=( a63640a  and  a63637a );
 a63642a <=( a63641a  and  a63634a );
 a63646a <=( A167  and  A168 );
 a63647a <=( A169  and  a63646a );
 a63650a <=( A201  and  (not A166) );
 a63653a <=( (not A203)  and  (not A202) );
 a63654a <=( a63653a  and  a63650a );
 a63655a <=( a63654a  and  a63647a );
 a63659a <=( (not A269)  and  (not A268) );
 a63660a <=( A267  and  a63659a );
 a63663a <=( (not A299)  and  A298 );
 a63666a <=( A302  and  A300 );
 a63667a <=( a63666a  and  a63663a );
 a63668a <=( a63667a  and  a63660a );
 a63672a <=( A167  and  A168 );
 a63673a <=( A169  and  a63672a );
 a63676a <=( A201  and  (not A166) );
 a63679a <=( (not A203)  and  (not A202) );
 a63680a <=( a63679a  and  a63676a );
 a63681a <=( a63680a  and  a63673a );
 a63685a <=( (not A269)  and  (not A268) );
 a63686a <=( A267  and  a63685a );
 a63689a <=( A299  and  (not A298) );
 a63692a <=( A301  and  A300 );
 a63693a <=( a63692a  and  a63689a );
 a63694a <=( a63693a  and  a63686a );
 a63698a <=( A167  and  A168 );
 a63699a <=( A169  and  a63698a );
 a63702a <=( A201  and  (not A166) );
 a63705a <=( (not A203)  and  (not A202) );
 a63706a <=( a63705a  and  a63702a );
 a63707a <=( a63706a  and  a63699a );
 a63711a <=( (not A269)  and  (not A268) );
 a63712a <=( A267  and  a63711a );
 a63715a <=( A299  and  (not A298) );
 a63718a <=( A302  and  A300 );
 a63719a <=( a63718a  and  a63715a );
 a63720a <=( a63719a  and  a63712a );
 a63724a <=( A167  and  A168 );
 a63725a <=( A169  and  a63724a );
 a63728a <=( A201  and  (not A166) );
 a63731a <=( (not A203)  and  (not A202) );
 a63732a <=( a63731a  and  a63728a );
 a63733a <=( a63732a  and  a63725a );
 a63737a <=( A298  and  A268 );
 a63738a <=( (not A267)  and  a63737a );
 a63741a <=( (not A300)  and  (not A299) );
 a63744a <=( (not A302)  and  (not A301) );
 a63745a <=( a63744a  and  a63741a );
 a63746a <=( a63745a  and  a63738a );
 a63750a <=( A167  and  A168 );
 a63751a <=( A169  and  a63750a );
 a63754a <=( A201  and  (not A166) );
 a63757a <=( (not A203)  and  (not A202) );
 a63758a <=( a63757a  and  a63754a );
 a63759a <=( a63758a  and  a63751a );
 a63763a <=( (not A298)  and  A268 );
 a63764a <=( (not A267)  and  a63763a );
 a63767a <=( (not A300)  and  A299 );
 a63770a <=( (not A302)  and  (not A301) );
 a63771a <=( a63770a  and  a63767a );
 a63772a <=( a63771a  and  a63764a );
 a63776a <=( A167  and  A168 );
 a63777a <=( A169  and  a63776a );
 a63780a <=( A201  and  (not A166) );
 a63783a <=( (not A203)  and  (not A202) );
 a63784a <=( a63783a  and  a63780a );
 a63785a <=( a63784a  and  a63777a );
 a63789a <=( A298  and  A269 );
 a63790a <=( (not A267)  and  a63789a );
 a63793a <=( (not A300)  and  (not A299) );
 a63796a <=( (not A302)  and  (not A301) );
 a63797a <=( a63796a  and  a63793a );
 a63798a <=( a63797a  and  a63790a );
 a63802a <=( A167  and  A168 );
 a63803a <=( A169  and  a63802a );
 a63806a <=( A201  and  (not A166) );
 a63809a <=( (not A203)  and  (not A202) );
 a63810a <=( a63809a  and  a63806a );
 a63811a <=( a63810a  and  a63803a );
 a63815a <=( (not A298)  and  A269 );
 a63816a <=( (not A267)  and  a63815a );
 a63819a <=( (not A300)  and  A299 );
 a63822a <=( (not A302)  and  (not A301) );
 a63823a <=( a63822a  and  a63819a );
 a63824a <=( a63823a  and  a63816a );
 a63828a <=( A167  and  A168 );
 a63829a <=( A169  and  a63828a );
 a63832a <=( A201  and  (not A166) );
 a63835a <=( (not A203)  and  (not A202) );
 a63836a <=( a63835a  and  a63832a );
 a63837a <=( a63836a  and  a63829a );
 a63841a <=( A298  and  A266 );
 a63842a <=( A265  and  a63841a );
 a63845a <=( (not A300)  and  (not A299) );
 a63848a <=( (not A302)  and  (not A301) );
 a63849a <=( a63848a  and  a63845a );
 a63850a <=( a63849a  and  a63842a );
 a63854a <=( A167  and  A168 );
 a63855a <=( A169  and  a63854a );
 a63858a <=( A201  and  (not A166) );
 a63861a <=( (not A203)  and  (not A202) );
 a63862a <=( a63861a  and  a63858a );
 a63863a <=( a63862a  and  a63855a );
 a63867a <=( (not A298)  and  A266 );
 a63868a <=( A265  and  a63867a );
 a63871a <=( (not A300)  and  A299 );
 a63874a <=( (not A302)  and  (not A301) );
 a63875a <=( a63874a  and  a63871a );
 a63876a <=( a63875a  and  a63868a );
 a63880a <=( A167  and  A168 );
 a63881a <=( A169  and  a63880a );
 a63884a <=( A201  and  (not A166) );
 a63887a <=( (not A203)  and  (not A202) );
 a63888a <=( a63887a  and  a63884a );
 a63889a <=( a63888a  and  a63881a );
 a63893a <=( A298  and  (not A266) );
 a63894a <=( (not A265)  and  a63893a );
 a63897a <=( (not A300)  and  (not A299) );
 a63900a <=( (not A302)  and  (not A301) );
 a63901a <=( a63900a  and  a63897a );
 a63902a <=( a63901a  and  a63894a );
 a63906a <=( A167  and  A168 );
 a63907a <=( A169  and  a63906a );
 a63910a <=( A201  and  (not A166) );
 a63913a <=( (not A203)  and  (not A202) );
 a63914a <=( a63913a  and  a63910a );
 a63915a <=( a63914a  and  a63907a );
 a63919a <=( (not A298)  and  (not A266) );
 a63920a <=( (not A265)  and  a63919a );
 a63923a <=( (not A300)  and  A299 );
 a63926a <=( (not A302)  and  (not A301) );
 a63927a <=( a63926a  and  a63923a );
 a63928a <=( a63927a  and  a63920a );
 a63932a <=( A167  and  A168 );
 a63933a <=( A169  and  a63932a );
 a63936a <=( (not A201)  and  (not A166) );
 a63939a <=( A267  and  A202 );
 a63940a <=( a63939a  and  a63936a );
 a63941a <=( a63940a  and  a63933a );
 a63945a <=( A298  and  (not A269) );
 a63946a <=( (not A268)  and  a63945a );
 a63949a <=( (not A300)  and  (not A299) );
 a63952a <=( (not A302)  and  (not A301) );
 a63953a <=( a63952a  and  a63949a );
 a63954a <=( a63953a  and  a63946a );
 a63958a <=( A167  and  A168 );
 a63959a <=( A169  and  a63958a );
 a63962a <=( (not A201)  and  (not A166) );
 a63965a <=( A267  and  A202 );
 a63966a <=( a63965a  and  a63962a );
 a63967a <=( a63966a  and  a63959a );
 a63971a <=( (not A298)  and  (not A269) );
 a63972a <=( (not A268)  and  a63971a );
 a63975a <=( (not A300)  and  A299 );
 a63978a <=( (not A302)  and  (not A301) );
 a63979a <=( a63978a  and  a63975a );
 a63980a <=( a63979a  and  a63972a );
 a63984a <=( A167  and  A168 );
 a63985a <=( A169  and  a63984a );
 a63988a <=( (not A201)  and  (not A166) );
 a63991a <=( A267  and  A203 );
 a63992a <=( a63991a  and  a63988a );
 a63993a <=( a63992a  and  a63985a );
 a63997a <=( A298  and  (not A269) );
 a63998a <=( (not A268)  and  a63997a );
 a64001a <=( (not A300)  and  (not A299) );
 a64004a <=( (not A302)  and  (not A301) );
 a64005a <=( a64004a  and  a64001a );
 a64006a <=( a64005a  and  a63998a );
 a64010a <=( A167  and  A168 );
 a64011a <=( A169  and  a64010a );
 a64014a <=( (not A201)  and  (not A166) );
 a64017a <=( A267  and  A203 );
 a64018a <=( a64017a  and  a64014a );
 a64019a <=( a64018a  and  a64011a );
 a64023a <=( (not A298)  and  (not A269) );
 a64024a <=( (not A268)  and  a64023a );
 a64027a <=( (not A300)  and  A299 );
 a64030a <=( (not A302)  and  (not A301) );
 a64031a <=( a64030a  and  a64027a );
 a64032a <=( a64031a  and  a64024a );
 a64036a <=( A167  and  A168 );
 a64037a <=( A169  and  a64036a );
 a64040a <=( A199  and  (not A166) );
 a64043a <=( A267  and  A200 );
 a64044a <=( a64043a  and  a64040a );
 a64045a <=( a64044a  and  a64037a );
 a64049a <=( A298  and  (not A269) );
 a64050a <=( (not A268)  and  a64049a );
 a64053a <=( (not A300)  and  (not A299) );
 a64056a <=( (not A302)  and  (not A301) );
 a64057a <=( a64056a  and  a64053a );
 a64058a <=( a64057a  and  a64050a );
 a64062a <=( A167  and  A168 );
 a64063a <=( A169  and  a64062a );
 a64066a <=( A199  and  (not A166) );
 a64069a <=( A267  and  A200 );
 a64070a <=( a64069a  and  a64066a );
 a64071a <=( a64070a  and  a64063a );
 a64075a <=( (not A298)  and  (not A269) );
 a64076a <=( (not A268)  and  a64075a );
 a64079a <=( (not A300)  and  A299 );
 a64082a <=( (not A302)  and  (not A301) );
 a64083a <=( a64082a  and  a64079a );
 a64084a <=( a64083a  and  a64076a );
 a64088a <=( A167  and  A168 );
 a64089a <=( A169  and  a64088a );
 a64092a <=( (not A199)  and  (not A166) );
 a64095a <=( A201  and  A200 );
 a64096a <=( a64095a  and  a64092a );
 a64097a <=( a64096a  and  a64089a );
 a64101a <=( A266  and  (not A265) );
 a64102a <=( A202  and  a64101a );
 a64105a <=( A268  and  A267 );
 a64108a <=( A301  and  (not A300) );
 a64109a <=( a64108a  and  a64105a );
 a64110a <=( a64109a  and  a64102a );
 a64114a <=( A167  and  A168 );
 a64115a <=( A169  and  a64114a );
 a64118a <=( (not A199)  and  (not A166) );
 a64121a <=( A201  and  A200 );
 a64122a <=( a64121a  and  a64118a );
 a64123a <=( a64122a  and  a64115a );
 a64127a <=( A266  and  (not A265) );
 a64128a <=( A202  and  a64127a );
 a64131a <=( A268  and  A267 );
 a64134a <=( A302  and  (not A300) );
 a64135a <=( a64134a  and  a64131a );
 a64136a <=( a64135a  and  a64128a );
 a64140a <=( A167  and  A168 );
 a64141a <=( A169  and  a64140a );
 a64144a <=( (not A199)  and  (not A166) );
 a64147a <=( A201  and  A200 );
 a64148a <=( a64147a  and  a64144a );
 a64149a <=( a64148a  and  a64141a );
 a64153a <=( A266  and  (not A265) );
 a64154a <=( A202  and  a64153a );
 a64157a <=( A268  and  A267 );
 a64160a <=( A299  and  A298 );
 a64161a <=( a64160a  and  a64157a );
 a64162a <=( a64161a  and  a64154a );
 a64166a <=( A167  and  A168 );
 a64167a <=( A169  and  a64166a );
 a64170a <=( (not A199)  and  (not A166) );
 a64173a <=( A201  and  A200 );
 a64174a <=( a64173a  and  a64170a );
 a64175a <=( a64174a  and  a64167a );
 a64179a <=( A266  and  (not A265) );
 a64180a <=( A202  and  a64179a );
 a64183a <=( A268  and  A267 );
 a64186a <=( (not A299)  and  (not A298) );
 a64187a <=( a64186a  and  a64183a );
 a64188a <=( a64187a  and  a64180a );
 a64192a <=( A167  and  A168 );
 a64193a <=( A169  and  a64192a );
 a64196a <=( (not A199)  and  (not A166) );
 a64199a <=( A201  and  A200 );
 a64200a <=( a64199a  and  a64196a );
 a64201a <=( a64200a  and  a64193a );
 a64205a <=( A266  and  (not A265) );
 a64206a <=( A202  and  a64205a );
 a64209a <=( A269  and  A267 );
 a64212a <=( A301  and  (not A300) );
 a64213a <=( a64212a  and  a64209a );
 a64214a <=( a64213a  and  a64206a );
 a64218a <=( A167  and  A168 );
 a64219a <=( A169  and  a64218a );
 a64222a <=( (not A199)  and  (not A166) );
 a64225a <=( A201  and  A200 );
 a64226a <=( a64225a  and  a64222a );
 a64227a <=( a64226a  and  a64219a );
 a64231a <=( A266  and  (not A265) );
 a64232a <=( A202  and  a64231a );
 a64235a <=( A269  and  A267 );
 a64238a <=( A302  and  (not A300) );
 a64239a <=( a64238a  and  a64235a );
 a64240a <=( a64239a  and  a64232a );
 a64244a <=( A167  and  A168 );
 a64245a <=( A169  and  a64244a );
 a64248a <=( (not A199)  and  (not A166) );
 a64251a <=( A201  and  A200 );
 a64252a <=( a64251a  and  a64248a );
 a64253a <=( a64252a  and  a64245a );
 a64257a <=( A266  and  (not A265) );
 a64258a <=( A202  and  a64257a );
 a64261a <=( A269  and  A267 );
 a64264a <=( A299  and  A298 );
 a64265a <=( a64264a  and  a64261a );
 a64266a <=( a64265a  and  a64258a );
 a64270a <=( A167  and  A168 );
 a64271a <=( A169  and  a64270a );
 a64274a <=( (not A199)  and  (not A166) );
 a64277a <=( A201  and  A200 );
 a64278a <=( a64277a  and  a64274a );
 a64279a <=( a64278a  and  a64271a );
 a64283a <=( A266  and  (not A265) );
 a64284a <=( A202  and  a64283a );
 a64287a <=( A269  and  A267 );
 a64290a <=( (not A299)  and  (not A298) );
 a64291a <=( a64290a  and  a64287a );
 a64292a <=( a64291a  and  a64284a );
 a64296a <=( A167  and  A168 );
 a64297a <=( A169  and  a64296a );
 a64300a <=( (not A199)  and  (not A166) );
 a64303a <=( A201  and  A200 );
 a64304a <=( a64303a  and  a64300a );
 a64305a <=( a64304a  and  a64297a );
 a64309a <=( (not A266)  and  A265 );
 a64310a <=( A202  and  a64309a );
 a64313a <=( A268  and  A267 );
 a64316a <=( A301  and  (not A300) );
 a64317a <=( a64316a  and  a64313a );
 a64318a <=( a64317a  and  a64310a );
 a64322a <=( A167  and  A168 );
 a64323a <=( A169  and  a64322a );
 a64326a <=( (not A199)  and  (not A166) );
 a64329a <=( A201  and  A200 );
 a64330a <=( a64329a  and  a64326a );
 a64331a <=( a64330a  and  a64323a );
 a64335a <=( (not A266)  and  A265 );
 a64336a <=( A202  and  a64335a );
 a64339a <=( A268  and  A267 );
 a64342a <=( A302  and  (not A300) );
 a64343a <=( a64342a  and  a64339a );
 a64344a <=( a64343a  and  a64336a );
 a64348a <=( A167  and  A168 );
 a64349a <=( A169  and  a64348a );
 a64352a <=( (not A199)  and  (not A166) );
 a64355a <=( A201  and  A200 );
 a64356a <=( a64355a  and  a64352a );
 a64357a <=( a64356a  and  a64349a );
 a64361a <=( (not A266)  and  A265 );
 a64362a <=( A202  and  a64361a );
 a64365a <=( A268  and  A267 );
 a64368a <=( A299  and  A298 );
 a64369a <=( a64368a  and  a64365a );
 a64370a <=( a64369a  and  a64362a );
 a64374a <=( A167  and  A168 );
 a64375a <=( A169  and  a64374a );
 a64378a <=( (not A199)  and  (not A166) );
 a64381a <=( A201  and  A200 );
 a64382a <=( a64381a  and  a64378a );
 a64383a <=( a64382a  and  a64375a );
 a64387a <=( (not A266)  and  A265 );
 a64388a <=( A202  and  a64387a );
 a64391a <=( A268  and  A267 );
 a64394a <=( (not A299)  and  (not A298) );
 a64395a <=( a64394a  and  a64391a );
 a64396a <=( a64395a  and  a64388a );
 a64400a <=( A167  and  A168 );
 a64401a <=( A169  and  a64400a );
 a64404a <=( (not A199)  and  (not A166) );
 a64407a <=( A201  and  A200 );
 a64408a <=( a64407a  and  a64404a );
 a64409a <=( a64408a  and  a64401a );
 a64413a <=( (not A266)  and  A265 );
 a64414a <=( A202  and  a64413a );
 a64417a <=( A269  and  A267 );
 a64420a <=( A301  and  (not A300) );
 a64421a <=( a64420a  and  a64417a );
 a64422a <=( a64421a  and  a64414a );
 a64426a <=( A167  and  A168 );
 a64427a <=( A169  and  a64426a );
 a64430a <=( (not A199)  and  (not A166) );
 a64433a <=( A201  and  A200 );
 a64434a <=( a64433a  and  a64430a );
 a64435a <=( a64434a  and  a64427a );
 a64439a <=( (not A266)  and  A265 );
 a64440a <=( A202  and  a64439a );
 a64443a <=( A269  and  A267 );
 a64446a <=( A302  and  (not A300) );
 a64447a <=( a64446a  and  a64443a );
 a64448a <=( a64447a  and  a64440a );
 a64452a <=( A167  and  A168 );
 a64453a <=( A169  and  a64452a );
 a64456a <=( (not A199)  and  (not A166) );
 a64459a <=( A201  and  A200 );
 a64460a <=( a64459a  and  a64456a );
 a64461a <=( a64460a  and  a64453a );
 a64465a <=( (not A266)  and  A265 );
 a64466a <=( A202  and  a64465a );
 a64469a <=( A269  and  A267 );
 a64472a <=( A299  and  A298 );
 a64473a <=( a64472a  and  a64469a );
 a64474a <=( a64473a  and  a64466a );
 a64478a <=( A167  and  A168 );
 a64479a <=( A169  and  a64478a );
 a64482a <=( (not A199)  and  (not A166) );
 a64485a <=( A201  and  A200 );
 a64486a <=( a64485a  and  a64482a );
 a64487a <=( a64486a  and  a64479a );
 a64491a <=( (not A266)  and  A265 );
 a64492a <=( A202  and  a64491a );
 a64495a <=( A269  and  A267 );
 a64498a <=( (not A299)  and  (not A298) );
 a64499a <=( a64498a  and  a64495a );
 a64500a <=( a64499a  and  a64492a );
 a64504a <=( A167  and  A168 );
 a64505a <=( A169  and  a64504a );
 a64508a <=( (not A199)  and  (not A166) );
 a64511a <=( A201  and  A200 );
 a64512a <=( a64511a  and  a64508a );
 a64513a <=( a64512a  and  a64505a );
 a64517a <=( A266  and  (not A265) );
 a64518a <=( A203  and  a64517a );
 a64521a <=( A268  and  A267 );
 a64524a <=( A301  and  (not A300) );
 a64525a <=( a64524a  and  a64521a );
 a64526a <=( a64525a  and  a64518a );
 a64530a <=( A167  and  A168 );
 a64531a <=( A169  and  a64530a );
 a64534a <=( (not A199)  and  (not A166) );
 a64537a <=( A201  and  A200 );
 a64538a <=( a64537a  and  a64534a );
 a64539a <=( a64538a  and  a64531a );
 a64543a <=( A266  and  (not A265) );
 a64544a <=( A203  and  a64543a );
 a64547a <=( A268  and  A267 );
 a64550a <=( A302  and  (not A300) );
 a64551a <=( a64550a  and  a64547a );
 a64552a <=( a64551a  and  a64544a );
 a64556a <=( A167  and  A168 );
 a64557a <=( A169  and  a64556a );
 a64560a <=( (not A199)  and  (not A166) );
 a64563a <=( A201  and  A200 );
 a64564a <=( a64563a  and  a64560a );
 a64565a <=( a64564a  and  a64557a );
 a64569a <=( A266  and  (not A265) );
 a64570a <=( A203  and  a64569a );
 a64573a <=( A268  and  A267 );
 a64576a <=( A299  and  A298 );
 a64577a <=( a64576a  and  a64573a );
 a64578a <=( a64577a  and  a64570a );
 a64582a <=( A167  and  A168 );
 a64583a <=( A169  and  a64582a );
 a64586a <=( (not A199)  and  (not A166) );
 a64589a <=( A201  and  A200 );
 a64590a <=( a64589a  and  a64586a );
 a64591a <=( a64590a  and  a64583a );
 a64595a <=( A266  and  (not A265) );
 a64596a <=( A203  and  a64595a );
 a64599a <=( A268  and  A267 );
 a64602a <=( (not A299)  and  (not A298) );
 a64603a <=( a64602a  and  a64599a );
 a64604a <=( a64603a  and  a64596a );
 a64608a <=( A167  and  A168 );
 a64609a <=( A169  and  a64608a );
 a64612a <=( (not A199)  and  (not A166) );
 a64615a <=( A201  and  A200 );
 a64616a <=( a64615a  and  a64612a );
 a64617a <=( a64616a  and  a64609a );
 a64621a <=( A266  and  (not A265) );
 a64622a <=( A203  and  a64621a );
 a64625a <=( A269  and  A267 );
 a64628a <=( A301  and  (not A300) );
 a64629a <=( a64628a  and  a64625a );
 a64630a <=( a64629a  and  a64622a );
 a64634a <=( A167  and  A168 );
 a64635a <=( A169  and  a64634a );
 a64638a <=( (not A199)  and  (not A166) );
 a64641a <=( A201  and  A200 );
 a64642a <=( a64641a  and  a64638a );
 a64643a <=( a64642a  and  a64635a );
 a64647a <=( A266  and  (not A265) );
 a64648a <=( A203  and  a64647a );
 a64651a <=( A269  and  A267 );
 a64654a <=( A302  and  (not A300) );
 a64655a <=( a64654a  and  a64651a );
 a64656a <=( a64655a  and  a64648a );
 a64660a <=( A167  and  A168 );
 a64661a <=( A169  and  a64660a );
 a64664a <=( (not A199)  and  (not A166) );
 a64667a <=( A201  and  A200 );
 a64668a <=( a64667a  and  a64664a );
 a64669a <=( a64668a  and  a64661a );
 a64673a <=( A266  and  (not A265) );
 a64674a <=( A203  and  a64673a );
 a64677a <=( A269  and  A267 );
 a64680a <=( A299  and  A298 );
 a64681a <=( a64680a  and  a64677a );
 a64682a <=( a64681a  and  a64674a );
 a64686a <=( A167  and  A168 );
 a64687a <=( A169  and  a64686a );
 a64690a <=( (not A199)  and  (not A166) );
 a64693a <=( A201  and  A200 );
 a64694a <=( a64693a  and  a64690a );
 a64695a <=( a64694a  and  a64687a );
 a64699a <=( A266  and  (not A265) );
 a64700a <=( A203  and  a64699a );
 a64703a <=( A269  and  A267 );
 a64706a <=( (not A299)  and  (not A298) );
 a64707a <=( a64706a  and  a64703a );
 a64708a <=( a64707a  and  a64700a );
 a64712a <=( A167  and  A168 );
 a64713a <=( A169  and  a64712a );
 a64716a <=( (not A199)  and  (not A166) );
 a64719a <=( A201  and  A200 );
 a64720a <=( a64719a  and  a64716a );
 a64721a <=( a64720a  and  a64713a );
 a64725a <=( (not A266)  and  A265 );
 a64726a <=( A203  and  a64725a );
 a64729a <=( A268  and  A267 );
 a64732a <=( A301  and  (not A300) );
 a64733a <=( a64732a  and  a64729a );
 a64734a <=( a64733a  and  a64726a );
 a64738a <=( A167  and  A168 );
 a64739a <=( A169  and  a64738a );
 a64742a <=( (not A199)  and  (not A166) );
 a64745a <=( A201  and  A200 );
 a64746a <=( a64745a  and  a64742a );
 a64747a <=( a64746a  and  a64739a );
 a64751a <=( (not A266)  and  A265 );
 a64752a <=( A203  and  a64751a );
 a64755a <=( A268  and  A267 );
 a64758a <=( A302  and  (not A300) );
 a64759a <=( a64758a  and  a64755a );
 a64760a <=( a64759a  and  a64752a );
 a64764a <=( A167  and  A168 );
 a64765a <=( A169  and  a64764a );
 a64768a <=( (not A199)  and  (not A166) );
 a64771a <=( A201  and  A200 );
 a64772a <=( a64771a  and  a64768a );
 a64773a <=( a64772a  and  a64765a );
 a64777a <=( (not A266)  and  A265 );
 a64778a <=( A203  and  a64777a );
 a64781a <=( A268  and  A267 );
 a64784a <=( A299  and  A298 );
 a64785a <=( a64784a  and  a64781a );
 a64786a <=( a64785a  and  a64778a );
 a64790a <=( A167  and  A168 );
 a64791a <=( A169  and  a64790a );
 a64794a <=( (not A199)  and  (not A166) );
 a64797a <=( A201  and  A200 );
 a64798a <=( a64797a  and  a64794a );
 a64799a <=( a64798a  and  a64791a );
 a64803a <=( (not A266)  and  A265 );
 a64804a <=( A203  and  a64803a );
 a64807a <=( A268  and  A267 );
 a64810a <=( (not A299)  and  (not A298) );
 a64811a <=( a64810a  and  a64807a );
 a64812a <=( a64811a  and  a64804a );
 a64816a <=( A167  and  A168 );
 a64817a <=( A169  and  a64816a );
 a64820a <=( (not A199)  and  (not A166) );
 a64823a <=( A201  and  A200 );
 a64824a <=( a64823a  and  a64820a );
 a64825a <=( a64824a  and  a64817a );
 a64829a <=( (not A266)  and  A265 );
 a64830a <=( A203  and  a64829a );
 a64833a <=( A269  and  A267 );
 a64836a <=( A301  and  (not A300) );
 a64837a <=( a64836a  and  a64833a );
 a64838a <=( a64837a  and  a64830a );
 a64842a <=( A167  and  A168 );
 a64843a <=( A169  and  a64842a );
 a64846a <=( (not A199)  and  (not A166) );
 a64849a <=( A201  and  A200 );
 a64850a <=( a64849a  and  a64846a );
 a64851a <=( a64850a  and  a64843a );
 a64855a <=( (not A266)  and  A265 );
 a64856a <=( A203  and  a64855a );
 a64859a <=( A269  and  A267 );
 a64862a <=( A302  and  (not A300) );
 a64863a <=( a64862a  and  a64859a );
 a64864a <=( a64863a  and  a64856a );
 a64868a <=( A167  and  A168 );
 a64869a <=( A169  and  a64868a );
 a64872a <=( (not A199)  and  (not A166) );
 a64875a <=( A201  and  A200 );
 a64876a <=( a64875a  and  a64872a );
 a64877a <=( a64876a  and  a64869a );
 a64881a <=( (not A266)  and  A265 );
 a64882a <=( A203  and  a64881a );
 a64885a <=( A269  and  A267 );
 a64888a <=( A299  and  A298 );
 a64889a <=( a64888a  and  a64885a );
 a64890a <=( a64889a  and  a64882a );
 a64894a <=( A167  and  A168 );
 a64895a <=( A169  and  a64894a );
 a64898a <=( (not A199)  and  (not A166) );
 a64901a <=( A201  and  A200 );
 a64902a <=( a64901a  and  a64898a );
 a64903a <=( a64902a  and  a64895a );
 a64907a <=( (not A266)  and  A265 );
 a64908a <=( A203  and  a64907a );
 a64911a <=( A269  and  A267 );
 a64914a <=( (not A299)  and  (not A298) );
 a64915a <=( a64914a  and  a64911a );
 a64916a <=( a64915a  and  a64908a );
 a64920a <=( A167  and  A168 );
 a64921a <=( A169  and  a64920a );
 a64924a <=( A199  and  (not A166) );
 a64927a <=( A201  and  (not A200) );
 a64928a <=( a64927a  and  a64924a );
 a64929a <=( a64928a  and  a64921a );
 a64933a <=( A266  and  (not A265) );
 a64934a <=( A202  and  a64933a );
 a64937a <=( A268  and  A267 );
 a64940a <=( A301  and  (not A300) );
 a64941a <=( a64940a  and  a64937a );
 a64942a <=( a64941a  and  a64934a );
 a64946a <=( A167  and  A168 );
 a64947a <=( A169  and  a64946a );
 a64950a <=( A199  and  (not A166) );
 a64953a <=( A201  and  (not A200) );
 a64954a <=( a64953a  and  a64950a );
 a64955a <=( a64954a  and  a64947a );
 a64959a <=( A266  and  (not A265) );
 a64960a <=( A202  and  a64959a );
 a64963a <=( A268  and  A267 );
 a64966a <=( A302  and  (not A300) );
 a64967a <=( a64966a  and  a64963a );
 a64968a <=( a64967a  and  a64960a );
 a64972a <=( A167  and  A168 );
 a64973a <=( A169  and  a64972a );
 a64976a <=( A199  and  (not A166) );
 a64979a <=( A201  and  (not A200) );
 a64980a <=( a64979a  and  a64976a );
 a64981a <=( a64980a  and  a64973a );
 a64985a <=( A266  and  (not A265) );
 a64986a <=( A202  and  a64985a );
 a64989a <=( A268  and  A267 );
 a64992a <=( A299  and  A298 );
 a64993a <=( a64992a  and  a64989a );
 a64994a <=( a64993a  and  a64986a );
 a64998a <=( A167  and  A168 );
 a64999a <=( A169  and  a64998a );
 a65002a <=( A199  and  (not A166) );
 a65005a <=( A201  and  (not A200) );
 a65006a <=( a65005a  and  a65002a );
 a65007a <=( a65006a  and  a64999a );
 a65011a <=( A266  and  (not A265) );
 a65012a <=( A202  and  a65011a );
 a65015a <=( A268  and  A267 );
 a65018a <=( (not A299)  and  (not A298) );
 a65019a <=( a65018a  and  a65015a );
 a65020a <=( a65019a  and  a65012a );
 a65024a <=( A167  and  A168 );
 a65025a <=( A169  and  a65024a );
 a65028a <=( A199  and  (not A166) );
 a65031a <=( A201  and  (not A200) );
 a65032a <=( a65031a  and  a65028a );
 a65033a <=( a65032a  and  a65025a );
 a65037a <=( A266  and  (not A265) );
 a65038a <=( A202  and  a65037a );
 a65041a <=( A269  and  A267 );
 a65044a <=( A301  and  (not A300) );
 a65045a <=( a65044a  and  a65041a );
 a65046a <=( a65045a  and  a65038a );
 a65050a <=( A167  and  A168 );
 a65051a <=( A169  and  a65050a );
 a65054a <=( A199  and  (not A166) );
 a65057a <=( A201  and  (not A200) );
 a65058a <=( a65057a  and  a65054a );
 a65059a <=( a65058a  and  a65051a );
 a65063a <=( A266  and  (not A265) );
 a65064a <=( A202  and  a65063a );
 a65067a <=( A269  and  A267 );
 a65070a <=( A302  and  (not A300) );
 a65071a <=( a65070a  and  a65067a );
 a65072a <=( a65071a  and  a65064a );
 a65076a <=( A167  and  A168 );
 a65077a <=( A169  and  a65076a );
 a65080a <=( A199  and  (not A166) );
 a65083a <=( A201  and  (not A200) );
 a65084a <=( a65083a  and  a65080a );
 a65085a <=( a65084a  and  a65077a );
 a65089a <=( A266  and  (not A265) );
 a65090a <=( A202  and  a65089a );
 a65093a <=( A269  and  A267 );
 a65096a <=( A299  and  A298 );
 a65097a <=( a65096a  and  a65093a );
 a65098a <=( a65097a  and  a65090a );
 a65102a <=( A167  and  A168 );
 a65103a <=( A169  and  a65102a );
 a65106a <=( A199  and  (not A166) );
 a65109a <=( A201  and  (not A200) );
 a65110a <=( a65109a  and  a65106a );
 a65111a <=( a65110a  and  a65103a );
 a65115a <=( A266  and  (not A265) );
 a65116a <=( A202  and  a65115a );
 a65119a <=( A269  and  A267 );
 a65122a <=( (not A299)  and  (not A298) );
 a65123a <=( a65122a  and  a65119a );
 a65124a <=( a65123a  and  a65116a );
 a65128a <=( A167  and  A168 );
 a65129a <=( A169  and  a65128a );
 a65132a <=( A199  and  (not A166) );
 a65135a <=( A201  and  (not A200) );
 a65136a <=( a65135a  and  a65132a );
 a65137a <=( a65136a  and  a65129a );
 a65141a <=( (not A266)  and  A265 );
 a65142a <=( A202  and  a65141a );
 a65145a <=( A268  and  A267 );
 a65148a <=( A301  and  (not A300) );
 a65149a <=( a65148a  and  a65145a );
 a65150a <=( a65149a  and  a65142a );
 a65154a <=( A167  and  A168 );
 a65155a <=( A169  and  a65154a );
 a65158a <=( A199  and  (not A166) );
 a65161a <=( A201  and  (not A200) );
 a65162a <=( a65161a  and  a65158a );
 a65163a <=( a65162a  and  a65155a );
 a65167a <=( (not A266)  and  A265 );
 a65168a <=( A202  and  a65167a );
 a65171a <=( A268  and  A267 );
 a65174a <=( A302  and  (not A300) );
 a65175a <=( a65174a  and  a65171a );
 a65176a <=( a65175a  and  a65168a );
 a65180a <=( A167  and  A168 );
 a65181a <=( A169  and  a65180a );
 a65184a <=( A199  and  (not A166) );
 a65187a <=( A201  and  (not A200) );
 a65188a <=( a65187a  and  a65184a );
 a65189a <=( a65188a  and  a65181a );
 a65193a <=( (not A266)  and  A265 );
 a65194a <=( A202  and  a65193a );
 a65197a <=( A268  and  A267 );
 a65200a <=( A299  and  A298 );
 a65201a <=( a65200a  and  a65197a );
 a65202a <=( a65201a  and  a65194a );
 a65206a <=( A167  and  A168 );
 a65207a <=( A169  and  a65206a );
 a65210a <=( A199  and  (not A166) );
 a65213a <=( A201  and  (not A200) );
 a65214a <=( a65213a  and  a65210a );
 a65215a <=( a65214a  and  a65207a );
 a65219a <=( (not A266)  and  A265 );
 a65220a <=( A202  and  a65219a );
 a65223a <=( A268  and  A267 );
 a65226a <=( (not A299)  and  (not A298) );
 a65227a <=( a65226a  and  a65223a );
 a65228a <=( a65227a  and  a65220a );
 a65232a <=( A167  and  A168 );
 a65233a <=( A169  and  a65232a );
 a65236a <=( A199  and  (not A166) );
 a65239a <=( A201  and  (not A200) );
 a65240a <=( a65239a  and  a65236a );
 a65241a <=( a65240a  and  a65233a );
 a65245a <=( (not A266)  and  A265 );
 a65246a <=( A202  and  a65245a );
 a65249a <=( A269  and  A267 );
 a65252a <=( A301  and  (not A300) );
 a65253a <=( a65252a  and  a65249a );
 a65254a <=( a65253a  and  a65246a );
 a65258a <=( A167  and  A168 );
 a65259a <=( A169  and  a65258a );
 a65262a <=( A199  and  (not A166) );
 a65265a <=( A201  and  (not A200) );
 a65266a <=( a65265a  and  a65262a );
 a65267a <=( a65266a  and  a65259a );
 a65271a <=( (not A266)  and  A265 );
 a65272a <=( A202  and  a65271a );
 a65275a <=( A269  and  A267 );
 a65278a <=( A302  and  (not A300) );
 a65279a <=( a65278a  and  a65275a );
 a65280a <=( a65279a  and  a65272a );
 a65284a <=( A167  and  A168 );
 a65285a <=( A169  and  a65284a );
 a65288a <=( A199  and  (not A166) );
 a65291a <=( A201  and  (not A200) );
 a65292a <=( a65291a  and  a65288a );
 a65293a <=( a65292a  and  a65285a );
 a65297a <=( (not A266)  and  A265 );
 a65298a <=( A202  and  a65297a );
 a65301a <=( A269  and  A267 );
 a65304a <=( A299  and  A298 );
 a65305a <=( a65304a  and  a65301a );
 a65306a <=( a65305a  and  a65298a );
 a65310a <=( A167  and  A168 );
 a65311a <=( A169  and  a65310a );
 a65314a <=( A199  and  (not A166) );
 a65317a <=( A201  and  (not A200) );
 a65318a <=( a65317a  and  a65314a );
 a65319a <=( a65318a  and  a65311a );
 a65323a <=( (not A266)  and  A265 );
 a65324a <=( A202  and  a65323a );
 a65327a <=( A269  and  A267 );
 a65330a <=( (not A299)  and  (not A298) );
 a65331a <=( a65330a  and  a65327a );
 a65332a <=( a65331a  and  a65324a );
 a65336a <=( A167  and  A168 );
 a65337a <=( A169  and  a65336a );
 a65340a <=( A199  and  (not A166) );
 a65343a <=( A201  and  (not A200) );
 a65344a <=( a65343a  and  a65340a );
 a65345a <=( a65344a  and  a65337a );
 a65349a <=( A266  and  (not A265) );
 a65350a <=( A203  and  a65349a );
 a65353a <=( A268  and  A267 );
 a65356a <=( A301  and  (not A300) );
 a65357a <=( a65356a  and  a65353a );
 a65358a <=( a65357a  and  a65350a );
 a65362a <=( A167  and  A168 );
 a65363a <=( A169  and  a65362a );
 a65366a <=( A199  and  (not A166) );
 a65369a <=( A201  and  (not A200) );
 a65370a <=( a65369a  and  a65366a );
 a65371a <=( a65370a  and  a65363a );
 a65375a <=( A266  and  (not A265) );
 a65376a <=( A203  and  a65375a );
 a65379a <=( A268  and  A267 );
 a65382a <=( A302  and  (not A300) );
 a65383a <=( a65382a  and  a65379a );
 a65384a <=( a65383a  and  a65376a );
 a65388a <=( A167  and  A168 );
 a65389a <=( A169  and  a65388a );
 a65392a <=( A199  and  (not A166) );
 a65395a <=( A201  and  (not A200) );
 a65396a <=( a65395a  and  a65392a );
 a65397a <=( a65396a  and  a65389a );
 a65401a <=( A266  and  (not A265) );
 a65402a <=( A203  and  a65401a );
 a65405a <=( A268  and  A267 );
 a65408a <=( A299  and  A298 );
 a65409a <=( a65408a  and  a65405a );
 a65410a <=( a65409a  and  a65402a );
 a65414a <=( A167  and  A168 );
 a65415a <=( A169  and  a65414a );
 a65418a <=( A199  and  (not A166) );
 a65421a <=( A201  and  (not A200) );
 a65422a <=( a65421a  and  a65418a );
 a65423a <=( a65422a  and  a65415a );
 a65427a <=( A266  and  (not A265) );
 a65428a <=( A203  and  a65427a );
 a65431a <=( A268  and  A267 );
 a65434a <=( (not A299)  and  (not A298) );
 a65435a <=( a65434a  and  a65431a );
 a65436a <=( a65435a  and  a65428a );
 a65440a <=( A167  and  A168 );
 a65441a <=( A169  and  a65440a );
 a65444a <=( A199  and  (not A166) );
 a65447a <=( A201  and  (not A200) );
 a65448a <=( a65447a  and  a65444a );
 a65449a <=( a65448a  and  a65441a );
 a65453a <=( A266  and  (not A265) );
 a65454a <=( A203  and  a65453a );
 a65457a <=( A269  and  A267 );
 a65460a <=( A301  and  (not A300) );
 a65461a <=( a65460a  and  a65457a );
 a65462a <=( a65461a  and  a65454a );
 a65466a <=( A167  and  A168 );
 a65467a <=( A169  and  a65466a );
 a65470a <=( A199  and  (not A166) );
 a65473a <=( A201  and  (not A200) );
 a65474a <=( a65473a  and  a65470a );
 a65475a <=( a65474a  and  a65467a );
 a65479a <=( A266  and  (not A265) );
 a65480a <=( A203  and  a65479a );
 a65483a <=( A269  and  A267 );
 a65486a <=( A302  and  (not A300) );
 a65487a <=( a65486a  and  a65483a );
 a65488a <=( a65487a  and  a65480a );
 a65492a <=( A167  and  A168 );
 a65493a <=( A169  and  a65492a );
 a65496a <=( A199  and  (not A166) );
 a65499a <=( A201  and  (not A200) );
 a65500a <=( a65499a  and  a65496a );
 a65501a <=( a65500a  and  a65493a );
 a65505a <=( A266  and  (not A265) );
 a65506a <=( A203  and  a65505a );
 a65509a <=( A269  and  A267 );
 a65512a <=( A299  and  A298 );
 a65513a <=( a65512a  and  a65509a );
 a65514a <=( a65513a  and  a65506a );
 a65518a <=( A167  and  A168 );
 a65519a <=( A169  and  a65518a );
 a65522a <=( A199  and  (not A166) );
 a65525a <=( A201  and  (not A200) );
 a65526a <=( a65525a  and  a65522a );
 a65527a <=( a65526a  and  a65519a );
 a65531a <=( A266  and  (not A265) );
 a65532a <=( A203  and  a65531a );
 a65535a <=( A269  and  A267 );
 a65538a <=( (not A299)  and  (not A298) );
 a65539a <=( a65538a  and  a65535a );
 a65540a <=( a65539a  and  a65532a );
 a65544a <=( A167  and  A168 );
 a65545a <=( A169  and  a65544a );
 a65548a <=( A199  and  (not A166) );
 a65551a <=( A201  and  (not A200) );
 a65552a <=( a65551a  and  a65548a );
 a65553a <=( a65552a  and  a65545a );
 a65557a <=( (not A266)  and  A265 );
 a65558a <=( A203  and  a65557a );
 a65561a <=( A268  and  A267 );
 a65564a <=( A301  and  (not A300) );
 a65565a <=( a65564a  and  a65561a );
 a65566a <=( a65565a  and  a65558a );
 a65570a <=( A167  and  A168 );
 a65571a <=( A169  and  a65570a );
 a65574a <=( A199  and  (not A166) );
 a65577a <=( A201  and  (not A200) );
 a65578a <=( a65577a  and  a65574a );
 a65579a <=( a65578a  and  a65571a );
 a65583a <=( (not A266)  and  A265 );
 a65584a <=( A203  and  a65583a );
 a65587a <=( A268  and  A267 );
 a65590a <=( A302  and  (not A300) );
 a65591a <=( a65590a  and  a65587a );
 a65592a <=( a65591a  and  a65584a );
 a65596a <=( A167  and  A168 );
 a65597a <=( A169  and  a65596a );
 a65600a <=( A199  and  (not A166) );
 a65603a <=( A201  and  (not A200) );
 a65604a <=( a65603a  and  a65600a );
 a65605a <=( a65604a  and  a65597a );
 a65609a <=( (not A266)  and  A265 );
 a65610a <=( A203  and  a65609a );
 a65613a <=( A268  and  A267 );
 a65616a <=( A299  and  A298 );
 a65617a <=( a65616a  and  a65613a );
 a65618a <=( a65617a  and  a65610a );
 a65622a <=( A167  and  A168 );
 a65623a <=( A169  and  a65622a );
 a65626a <=( A199  and  (not A166) );
 a65629a <=( A201  and  (not A200) );
 a65630a <=( a65629a  and  a65626a );
 a65631a <=( a65630a  and  a65623a );
 a65635a <=( (not A266)  and  A265 );
 a65636a <=( A203  and  a65635a );
 a65639a <=( A268  and  A267 );
 a65642a <=( (not A299)  and  (not A298) );
 a65643a <=( a65642a  and  a65639a );
 a65644a <=( a65643a  and  a65636a );
 a65648a <=( A167  and  A168 );
 a65649a <=( A169  and  a65648a );
 a65652a <=( A199  and  (not A166) );
 a65655a <=( A201  and  (not A200) );
 a65656a <=( a65655a  and  a65652a );
 a65657a <=( a65656a  and  a65649a );
 a65661a <=( (not A266)  and  A265 );
 a65662a <=( A203  and  a65661a );
 a65665a <=( A269  and  A267 );
 a65668a <=( A301  and  (not A300) );
 a65669a <=( a65668a  and  a65665a );
 a65670a <=( a65669a  and  a65662a );
 a65674a <=( A167  and  A168 );
 a65675a <=( A169  and  a65674a );
 a65678a <=( A199  and  (not A166) );
 a65681a <=( A201  and  (not A200) );
 a65682a <=( a65681a  and  a65678a );
 a65683a <=( a65682a  and  a65675a );
 a65687a <=( (not A266)  and  A265 );
 a65688a <=( A203  and  a65687a );
 a65691a <=( A269  and  A267 );
 a65694a <=( A302  and  (not A300) );
 a65695a <=( a65694a  and  a65691a );
 a65696a <=( a65695a  and  a65688a );
 a65700a <=( A167  and  A168 );
 a65701a <=( A169  and  a65700a );
 a65704a <=( A199  and  (not A166) );
 a65707a <=( A201  and  (not A200) );
 a65708a <=( a65707a  and  a65704a );
 a65709a <=( a65708a  and  a65701a );
 a65713a <=( (not A266)  and  A265 );
 a65714a <=( A203  and  a65713a );
 a65717a <=( A269  and  A267 );
 a65720a <=( A299  and  A298 );
 a65721a <=( a65720a  and  a65717a );
 a65722a <=( a65721a  and  a65714a );
 a65726a <=( A167  and  A168 );
 a65727a <=( A169  and  a65726a );
 a65730a <=( A199  and  (not A166) );
 a65733a <=( A201  and  (not A200) );
 a65734a <=( a65733a  and  a65730a );
 a65735a <=( a65734a  and  a65727a );
 a65739a <=( (not A266)  and  A265 );
 a65740a <=( A203  and  a65739a );
 a65743a <=( A269  and  A267 );
 a65746a <=( (not A299)  and  (not A298) );
 a65747a <=( a65746a  and  a65743a );
 a65748a <=( a65747a  and  a65740a );
 a65752a <=( A167  and  A168 );
 a65753a <=( A169  and  a65752a );
 a65756a <=( (not A199)  and  (not A166) );
 a65759a <=( A267  and  (not A200) );
 a65760a <=( a65759a  and  a65756a );
 a65761a <=( a65760a  and  a65753a );
 a65765a <=( A298  and  (not A269) );
 a65766a <=( (not A268)  and  a65765a );
 a65769a <=( (not A300)  and  (not A299) );
 a65772a <=( (not A302)  and  (not A301) );
 a65773a <=( a65772a  and  a65769a );
 a65774a <=( a65773a  and  a65766a );
 a65778a <=( A167  and  A168 );
 a65779a <=( A169  and  a65778a );
 a65782a <=( (not A199)  and  (not A166) );
 a65785a <=( A267  and  (not A200) );
 a65786a <=( a65785a  and  a65782a );
 a65787a <=( a65786a  and  a65779a );
 a65791a <=( (not A298)  and  (not A269) );
 a65792a <=( (not A268)  and  a65791a );
 a65795a <=( (not A300)  and  A299 );
 a65798a <=( (not A302)  and  (not A301) );
 a65799a <=( a65798a  and  a65795a );
 a65800a <=( a65799a  and  a65792a );
 a65804a <=( (not A167)  and  A168 );
 a65805a <=( A169  and  a65804a );
 a65808a <=( A201  and  A166 );
 a65811a <=( (not A203)  and  (not A202) );
 a65812a <=( a65811a  and  a65808a );
 a65813a <=( a65812a  and  a65805a );
 a65817a <=( (not A269)  and  (not A268) );
 a65818a <=( A267  and  a65817a );
 a65821a <=( (not A299)  and  A298 );
 a65824a <=( A301  and  A300 );
 a65825a <=( a65824a  and  a65821a );
 a65826a <=( a65825a  and  a65818a );
 a65830a <=( (not A167)  and  A168 );
 a65831a <=( A169  and  a65830a );
 a65834a <=( A201  and  A166 );
 a65837a <=( (not A203)  and  (not A202) );
 a65838a <=( a65837a  and  a65834a );
 a65839a <=( a65838a  and  a65831a );
 a65843a <=( (not A269)  and  (not A268) );
 a65844a <=( A267  and  a65843a );
 a65847a <=( (not A299)  and  A298 );
 a65850a <=( A302  and  A300 );
 a65851a <=( a65850a  and  a65847a );
 a65852a <=( a65851a  and  a65844a );
 a65856a <=( (not A167)  and  A168 );
 a65857a <=( A169  and  a65856a );
 a65860a <=( A201  and  A166 );
 a65863a <=( (not A203)  and  (not A202) );
 a65864a <=( a65863a  and  a65860a );
 a65865a <=( a65864a  and  a65857a );
 a65869a <=( (not A269)  and  (not A268) );
 a65870a <=( A267  and  a65869a );
 a65873a <=( A299  and  (not A298) );
 a65876a <=( A301  and  A300 );
 a65877a <=( a65876a  and  a65873a );
 a65878a <=( a65877a  and  a65870a );
 a65882a <=( (not A167)  and  A168 );
 a65883a <=( A169  and  a65882a );
 a65886a <=( A201  and  A166 );
 a65889a <=( (not A203)  and  (not A202) );
 a65890a <=( a65889a  and  a65886a );
 a65891a <=( a65890a  and  a65883a );
 a65895a <=( (not A269)  and  (not A268) );
 a65896a <=( A267  and  a65895a );
 a65899a <=( A299  and  (not A298) );
 a65902a <=( A302  and  A300 );
 a65903a <=( a65902a  and  a65899a );
 a65904a <=( a65903a  and  a65896a );
 a65908a <=( (not A167)  and  A168 );
 a65909a <=( A169  and  a65908a );
 a65912a <=( A201  and  A166 );
 a65915a <=( (not A203)  and  (not A202) );
 a65916a <=( a65915a  and  a65912a );
 a65917a <=( a65916a  and  a65909a );
 a65921a <=( A298  and  A268 );
 a65922a <=( (not A267)  and  a65921a );
 a65925a <=( (not A300)  and  (not A299) );
 a65928a <=( (not A302)  and  (not A301) );
 a65929a <=( a65928a  and  a65925a );
 a65930a <=( a65929a  and  a65922a );
 a65934a <=( (not A167)  and  A168 );
 a65935a <=( A169  and  a65934a );
 a65938a <=( A201  and  A166 );
 a65941a <=( (not A203)  and  (not A202) );
 a65942a <=( a65941a  and  a65938a );
 a65943a <=( a65942a  and  a65935a );
 a65947a <=( (not A298)  and  A268 );
 a65948a <=( (not A267)  and  a65947a );
 a65951a <=( (not A300)  and  A299 );
 a65954a <=( (not A302)  and  (not A301) );
 a65955a <=( a65954a  and  a65951a );
 a65956a <=( a65955a  and  a65948a );
 a65960a <=( (not A167)  and  A168 );
 a65961a <=( A169  and  a65960a );
 a65964a <=( A201  and  A166 );
 a65967a <=( (not A203)  and  (not A202) );
 a65968a <=( a65967a  and  a65964a );
 a65969a <=( a65968a  and  a65961a );
 a65973a <=( A298  and  A269 );
 a65974a <=( (not A267)  and  a65973a );
 a65977a <=( (not A300)  and  (not A299) );
 a65980a <=( (not A302)  and  (not A301) );
 a65981a <=( a65980a  and  a65977a );
 a65982a <=( a65981a  and  a65974a );
 a65986a <=( (not A167)  and  A168 );
 a65987a <=( A169  and  a65986a );
 a65990a <=( A201  and  A166 );
 a65993a <=( (not A203)  and  (not A202) );
 a65994a <=( a65993a  and  a65990a );
 a65995a <=( a65994a  and  a65987a );
 a65999a <=( (not A298)  and  A269 );
 a66000a <=( (not A267)  and  a65999a );
 a66003a <=( (not A300)  and  A299 );
 a66006a <=( (not A302)  and  (not A301) );
 a66007a <=( a66006a  and  a66003a );
 a66008a <=( a66007a  and  a66000a );
 a66012a <=( (not A167)  and  A168 );
 a66013a <=( A169  and  a66012a );
 a66016a <=( A201  and  A166 );
 a66019a <=( (not A203)  and  (not A202) );
 a66020a <=( a66019a  and  a66016a );
 a66021a <=( a66020a  and  a66013a );
 a66025a <=( A298  and  A266 );
 a66026a <=( A265  and  a66025a );
 a66029a <=( (not A300)  and  (not A299) );
 a66032a <=( (not A302)  and  (not A301) );
 a66033a <=( a66032a  and  a66029a );
 a66034a <=( a66033a  and  a66026a );
 a66038a <=( (not A167)  and  A168 );
 a66039a <=( A169  and  a66038a );
 a66042a <=( A201  and  A166 );
 a66045a <=( (not A203)  and  (not A202) );
 a66046a <=( a66045a  and  a66042a );
 a66047a <=( a66046a  and  a66039a );
 a66051a <=( (not A298)  and  A266 );
 a66052a <=( A265  and  a66051a );
 a66055a <=( (not A300)  and  A299 );
 a66058a <=( (not A302)  and  (not A301) );
 a66059a <=( a66058a  and  a66055a );
 a66060a <=( a66059a  and  a66052a );
 a66064a <=( (not A167)  and  A168 );
 a66065a <=( A169  and  a66064a );
 a66068a <=( A201  and  A166 );
 a66071a <=( (not A203)  and  (not A202) );
 a66072a <=( a66071a  and  a66068a );
 a66073a <=( a66072a  and  a66065a );
 a66077a <=( A298  and  (not A266) );
 a66078a <=( (not A265)  and  a66077a );
 a66081a <=( (not A300)  and  (not A299) );
 a66084a <=( (not A302)  and  (not A301) );
 a66085a <=( a66084a  and  a66081a );
 a66086a <=( a66085a  and  a66078a );
 a66090a <=( (not A167)  and  A168 );
 a66091a <=( A169  and  a66090a );
 a66094a <=( A201  and  A166 );
 a66097a <=( (not A203)  and  (not A202) );
 a66098a <=( a66097a  and  a66094a );
 a66099a <=( a66098a  and  a66091a );
 a66103a <=( (not A298)  and  (not A266) );
 a66104a <=( (not A265)  and  a66103a );
 a66107a <=( (not A300)  and  A299 );
 a66110a <=( (not A302)  and  (not A301) );
 a66111a <=( a66110a  and  a66107a );
 a66112a <=( a66111a  and  a66104a );
 a66116a <=( (not A167)  and  A168 );
 a66117a <=( A169  and  a66116a );
 a66120a <=( (not A201)  and  A166 );
 a66123a <=( A267  and  A202 );
 a66124a <=( a66123a  and  a66120a );
 a66125a <=( a66124a  and  a66117a );
 a66129a <=( A298  and  (not A269) );
 a66130a <=( (not A268)  and  a66129a );
 a66133a <=( (not A300)  and  (not A299) );
 a66136a <=( (not A302)  and  (not A301) );
 a66137a <=( a66136a  and  a66133a );
 a66138a <=( a66137a  and  a66130a );
 a66142a <=( (not A167)  and  A168 );
 a66143a <=( A169  and  a66142a );
 a66146a <=( (not A201)  and  A166 );
 a66149a <=( A267  and  A202 );
 a66150a <=( a66149a  and  a66146a );
 a66151a <=( a66150a  and  a66143a );
 a66155a <=( (not A298)  and  (not A269) );
 a66156a <=( (not A268)  and  a66155a );
 a66159a <=( (not A300)  and  A299 );
 a66162a <=( (not A302)  and  (not A301) );
 a66163a <=( a66162a  and  a66159a );
 a66164a <=( a66163a  and  a66156a );
 a66168a <=( (not A167)  and  A168 );
 a66169a <=( A169  and  a66168a );
 a66172a <=( (not A201)  and  A166 );
 a66175a <=( A267  and  A203 );
 a66176a <=( a66175a  and  a66172a );
 a66177a <=( a66176a  and  a66169a );
 a66181a <=( A298  and  (not A269) );
 a66182a <=( (not A268)  and  a66181a );
 a66185a <=( (not A300)  and  (not A299) );
 a66188a <=( (not A302)  and  (not A301) );
 a66189a <=( a66188a  and  a66185a );
 a66190a <=( a66189a  and  a66182a );
 a66194a <=( (not A167)  and  A168 );
 a66195a <=( A169  and  a66194a );
 a66198a <=( (not A201)  and  A166 );
 a66201a <=( A267  and  A203 );
 a66202a <=( a66201a  and  a66198a );
 a66203a <=( a66202a  and  a66195a );
 a66207a <=( (not A298)  and  (not A269) );
 a66208a <=( (not A268)  and  a66207a );
 a66211a <=( (not A300)  and  A299 );
 a66214a <=( (not A302)  and  (not A301) );
 a66215a <=( a66214a  and  a66211a );
 a66216a <=( a66215a  and  a66208a );
 a66220a <=( (not A167)  and  A168 );
 a66221a <=( A169  and  a66220a );
 a66224a <=( A199  and  A166 );
 a66227a <=( A267  and  A200 );
 a66228a <=( a66227a  and  a66224a );
 a66229a <=( a66228a  and  a66221a );
 a66233a <=( A298  and  (not A269) );
 a66234a <=( (not A268)  and  a66233a );
 a66237a <=( (not A300)  and  (not A299) );
 a66240a <=( (not A302)  and  (not A301) );
 a66241a <=( a66240a  and  a66237a );
 a66242a <=( a66241a  and  a66234a );
 a66246a <=( (not A167)  and  A168 );
 a66247a <=( A169  and  a66246a );
 a66250a <=( A199  and  A166 );
 a66253a <=( A267  and  A200 );
 a66254a <=( a66253a  and  a66250a );
 a66255a <=( a66254a  and  a66247a );
 a66259a <=( (not A298)  and  (not A269) );
 a66260a <=( (not A268)  and  a66259a );
 a66263a <=( (not A300)  and  A299 );
 a66266a <=( (not A302)  and  (not A301) );
 a66267a <=( a66266a  and  a66263a );
 a66268a <=( a66267a  and  a66260a );
 a66272a <=( (not A167)  and  A168 );
 a66273a <=( A169  and  a66272a );
 a66276a <=( (not A199)  and  A166 );
 a66279a <=( A201  and  A200 );
 a66280a <=( a66279a  and  a66276a );
 a66281a <=( a66280a  and  a66273a );
 a66285a <=( A266  and  (not A265) );
 a66286a <=( A202  and  a66285a );
 a66289a <=( A268  and  A267 );
 a66292a <=( A301  and  (not A300) );
 a66293a <=( a66292a  and  a66289a );
 a66294a <=( a66293a  and  a66286a );
 a66298a <=( (not A167)  and  A168 );
 a66299a <=( A169  and  a66298a );
 a66302a <=( (not A199)  and  A166 );
 a66305a <=( A201  and  A200 );
 a66306a <=( a66305a  and  a66302a );
 a66307a <=( a66306a  and  a66299a );
 a66311a <=( A266  and  (not A265) );
 a66312a <=( A202  and  a66311a );
 a66315a <=( A268  and  A267 );
 a66318a <=( A302  and  (not A300) );
 a66319a <=( a66318a  and  a66315a );
 a66320a <=( a66319a  and  a66312a );
 a66324a <=( (not A167)  and  A168 );
 a66325a <=( A169  and  a66324a );
 a66328a <=( (not A199)  and  A166 );
 a66331a <=( A201  and  A200 );
 a66332a <=( a66331a  and  a66328a );
 a66333a <=( a66332a  and  a66325a );
 a66337a <=( A266  and  (not A265) );
 a66338a <=( A202  and  a66337a );
 a66341a <=( A268  and  A267 );
 a66344a <=( A299  and  A298 );
 a66345a <=( a66344a  and  a66341a );
 a66346a <=( a66345a  and  a66338a );
 a66350a <=( (not A167)  and  A168 );
 a66351a <=( A169  and  a66350a );
 a66354a <=( (not A199)  and  A166 );
 a66357a <=( A201  and  A200 );
 a66358a <=( a66357a  and  a66354a );
 a66359a <=( a66358a  and  a66351a );
 a66363a <=( A266  and  (not A265) );
 a66364a <=( A202  and  a66363a );
 a66367a <=( A268  and  A267 );
 a66370a <=( (not A299)  and  (not A298) );
 a66371a <=( a66370a  and  a66367a );
 a66372a <=( a66371a  and  a66364a );
 a66376a <=( (not A167)  and  A168 );
 a66377a <=( A169  and  a66376a );
 a66380a <=( (not A199)  and  A166 );
 a66383a <=( A201  and  A200 );
 a66384a <=( a66383a  and  a66380a );
 a66385a <=( a66384a  and  a66377a );
 a66389a <=( A266  and  (not A265) );
 a66390a <=( A202  and  a66389a );
 a66393a <=( A269  and  A267 );
 a66396a <=( A301  and  (not A300) );
 a66397a <=( a66396a  and  a66393a );
 a66398a <=( a66397a  and  a66390a );
 a66402a <=( (not A167)  and  A168 );
 a66403a <=( A169  and  a66402a );
 a66406a <=( (not A199)  and  A166 );
 a66409a <=( A201  and  A200 );
 a66410a <=( a66409a  and  a66406a );
 a66411a <=( a66410a  and  a66403a );
 a66415a <=( A266  and  (not A265) );
 a66416a <=( A202  and  a66415a );
 a66419a <=( A269  and  A267 );
 a66422a <=( A302  and  (not A300) );
 a66423a <=( a66422a  and  a66419a );
 a66424a <=( a66423a  and  a66416a );
 a66428a <=( (not A167)  and  A168 );
 a66429a <=( A169  and  a66428a );
 a66432a <=( (not A199)  and  A166 );
 a66435a <=( A201  and  A200 );
 a66436a <=( a66435a  and  a66432a );
 a66437a <=( a66436a  and  a66429a );
 a66441a <=( A266  and  (not A265) );
 a66442a <=( A202  and  a66441a );
 a66445a <=( A269  and  A267 );
 a66448a <=( A299  and  A298 );
 a66449a <=( a66448a  and  a66445a );
 a66450a <=( a66449a  and  a66442a );
 a66454a <=( (not A167)  and  A168 );
 a66455a <=( A169  and  a66454a );
 a66458a <=( (not A199)  and  A166 );
 a66461a <=( A201  and  A200 );
 a66462a <=( a66461a  and  a66458a );
 a66463a <=( a66462a  and  a66455a );
 a66467a <=( A266  and  (not A265) );
 a66468a <=( A202  and  a66467a );
 a66471a <=( A269  and  A267 );
 a66474a <=( (not A299)  and  (not A298) );
 a66475a <=( a66474a  and  a66471a );
 a66476a <=( a66475a  and  a66468a );
 a66480a <=( (not A167)  and  A168 );
 a66481a <=( A169  and  a66480a );
 a66484a <=( (not A199)  and  A166 );
 a66487a <=( A201  and  A200 );
 a66488a <=( a66487a  and  a66484a );
 a66489a <=( a66488a  and  a66481a );
 a66493a <=( (not A266)  and  A265 );
 a66494a <=( A202  and  a66493a );
 a66497a <=( A268  and  A267 );
 a66500a <=( A301  and  (not A300) );
 a66501a <=( a66500a  and  a66497a );
 a66502a <=( a66501a  and  a66494a );
 a66506a <=( (not A167)  and  A168 );
 a66507a <=( A169  and  a66506a );
 a66510a <=( (not A199)  and  A166 );
 a66513a <=( A201  and  A200 );
 a66514a <=( a66513a  and  a66510a );
 a66515a <=( a66514a  and  a66507a );
 a66519a <=( (not A266)  and  A265 );
 a66520a <=( A202  and  a66519a );
 a66523a <=( A268  and  A267 );
 a66526a <=( A302  and  (not A300) );
 a66527a <=( a66526a  and  a66523a );
 a66528a <=( a66527a  and  a66520a );
 a66532a <=( (not A167)  and  A168 );
 a66533a <=( A169  and  a66532a );
 a66536a <=( (not A199)  and  A166 );
 a66539a <=( A201  and  A200 );
 a66540a <=( a66539a  and  a66536a );
 a66541a <=( a66540a  and  a66533a );
 a66545a <=( (not A266)  and  A265 );
 a66546a <=( A202  and  a66545a );
 a66549a <=( A268  and  A267 );
 a66552a <=( A299  and  A298 );
 a66553a <=( a66552a  and  a66549a );
 a66554a <=( a66553a  and  a66546a );
 a66558a <=( (not A167)  and  A168 );
 a66559a <=( A169  and  a66558a );
 a66562a <=( (not A199)  and  A166 );
 a66565a <=( A201  and  A200 );
 a66566a <=( a66565a  and  a66562a );
 a66567a <=( a66566a  and  a66559a );
 a66571a <=( (not A266)  and  A265 );
 a66572a <=( A202  and  a66571a );
 a66575a <=( A268  and  A267 );
 a66578a <=( (not A299)  and  (not A298) );
 a66579a <=( a66578a  and  a66575a );
 a66580a <=( a66579a  and  a66572a );
 a66584a <=( (not A167)  and  A168 );
 a66585a <=( A169  and  a66584a );
 a66588a <=( (not A199)  and  A166 );
 a66591a <=( A201  and  A200 );
 a66592a <=( a66591a  and  a66588a );
 a66593a <=( a66592a  and  a66585a );
 a66597a <=( (not A266)  and  A265 );
 a66598a <=( A202  and  a66597a );
 a66601a <=( A269  and  A267 );
 a66604a <=( A301  and  (not A300) );
 a66605a <=( a66604a  and  a66601a );
 a66606a <=( a66605a  and  a66598a );
 a66610a <=( (not A167)  and  A168 );
 a66611a <=( A169  and  a66610a );
 a66614a <=( (not A199)  and  A166 );
 a66617a <=( A201  and  A200 );
 a66618a <=( a66617a  and  a66614a );
 a66619a <=( a66618a  and  a66611a );
 a66623a <=( (not A266)  and  A265 );
 a66624a <=( A202  and  a66623a );
 a66627a <=( A269  and  A267 );
 a66630a <=( A302  and  (not A300) );
 a66631a <=( a66630a  and  a66627a );
 a66632a <=( a66631a  and  a66624a );
 a66636a <=( (not A167)  and  A168 );
 a66637a <=( A169  and  a66636a );
 a66640a <=( (not A199)  and  A166 );
 a66643a <=( A201  and  A200 );
 a66644a <=( a66643a  and  a66640a );
 a66645a <=( a66644a  and  a66637a );
 a66649a <=( (not A266)  and  A265 );
 a66650a <=( A202  and  a66649a );
 a66653a <=( A269  and  A267 );
 a66656a <=( A299  and  A298 );
 a66657a <=( a66656a  and  a66653a );
 a66658a <=( a66657a  and  a66650a );
 a66662a <=( (not A167)  and  A168 );
 a66663a <=( A169  and  a66662a );
 a66666a <=( (not A199)  and  A166 );
 a66669a <=( A201  and  A200 );
 a66670a <=( a66669a  and  a66666a );
 a66671a <=( a66670a  and  a66663a );
 a66675a <=( (not A266)  and  A265 );
 a66676a <=( A202  and  a66675a );
 a66679a <=( A269  and  A267 );
 a66682a <=( (not A299)  and  (not A298) );
 a66683a <=( a66682a  and  a66679a );
 a66684a <=( a66683a  and  a66676a );
 a66688a <=( (not A167)  and  A168 );
 a66689a <=( A169  and  a66688a );
 a66692a <=( (not A199)  and  A166 );
 a66695a <=( A201  and  A200 );
 a66696a <=( a66695a  and  a66692a );
 a66697a <=( a66696a  and  a66689a );
 a66701a <=( A266  and  (not A265) );
 a66702a <=( A203  and  a66701a );
 a66705a <=( A268  and  A267 );
 a66708a <=( A301  and  (not A300) );
 a66709a <=( a66708a  and  a66705a );
 a66710a <=( a66709a  and  a66702a );
 a66714a <=( (not A167)  and  A168 );
 a66715a <=( A169  and  a66714a );
 a66718a <=( (not A199)  and  A166 );
 a66721a <=( A201  and  A200 );
 a66722a <=( a66721a  and  a66718a );
 a66723a <=( a66722a  and  a66715a );
 a66727a <=( A266  and  (not A265) );
 a66728a <=( A203  and  a66727a );
 a66731a <=( A268  and  A267 );
 a66734a <=( A302  and  (not A300) );
 a66735a <=( a66734a  and  a66731a );
 a66736a <=( a66735a  and  a66728a );
 a66740a <=( (not A167)  and  A168 );
 a66741a <=( A169  and  a66740a );
 a66744a <=( (not A199)  and  A166 );
 a66747a <=( A201  and  A200 );
 a66748a <=( a66747a  and  a66744a );
 a66749a <=( a66748a  and  a66741a );
 a66753a <=( A266  and  (not A265) );
 a66754a <=( A203  and  a66753a );
 a66757a <=( A268  and  A267 );
 a66760a <=( A299  and  A298 );
 a66761a <=( a66760a  and  a66757a );
 a66762a <=( a66761a  and  a66754a );
 a66766a <=( (not A167)  and  A168 );
 a66767a <=( A169  and  a66766a );
 a66770a <=( (not A199)  and  A166 );
 a66773a <=( A201  and  A200 );
 a66774a <=( a66773a  and  a66770a );
 a66775a <=( a66774a  and  a66767a );
 a66779a <=( A266  and  (not A265) );
 a66780a <=( A203  and  a66779a );
 a66783a <=( A268  and  A267 );
 a66786a <=( (not A299)  and  (not A298) );
 a66787a <=( a66786a  and  a66783a );
 a66788a <=( a66787a  and  a66780a );
 a66792a <=( (not A167)  and  A168 );
 a66793a <=( A169  and  a66792a );
 a66796a <=( (not A199)  and  A166 );
 a66799a <=( A201  and  A200 );
 a66800a <=( a66799a  and  a66796a );
 a66801a <=( a66800a  and  a66793a );
 a66805a <=( A266  and  (not A265) );
 a66806a <=( A203  and  a66805a );
 a66809a <=( A269  and  A267 );
 a66812a <=( A301  and  (not A300) );
 a66813a <=( a66812a  and  a66809a );
 a66814a <=( a66813a  and  a66806a );
 a66818a <=( (not A167)  and  A168 );
 a66819a <=( A169  and  a66818a );
 a66822a <=( (not A199)  and  A166 );
 a66825a <=( A201  and  A200 );
 a66826a <=( a66825a  and  a66822a );
 a66827a <=( a66826a  and  a66819a );
 a66831a <=( A266  and  (not A265) );
 a66832a <=( A203  and  a66831a );
 a66835a <=( A269  and  A267 );
 a66838a <=( A302  and  (not A300) );
 a66839a <=( a66838a  and  a66835a );
 a66840a <=( a66839a  and  a66832a );
 a66844a <=( (not A167)  and  A168 );
 a66845a <=( A169  and  a66844a );
 a66848a <=( (not A199)  and  A166 );
 a66851a <=( A201  and  A200 );
 a66852a <=( a66851a  and  a66848a );
 a66853a <=( a66852a  and  a66845a );
 a66857a <=( A266  and  (not A265) );
 a66858a <=( A203  and  a66857a );
 a66861a <=( A269  and  A267 );
 a66864a <=( A299  and  A298 );
 a66865a <=( a66864a  and  a66861a );
 a66866a <=( a66865a  and  a66858a );
 a66870a <=( (not A167)  and  A168 );
 a66871a <=( A169  and  a66870a );
 a66874a <=( (not A199)  and  A166 );
 a66877a <=( A201  and  A200 );
 a66878a <=( a66877a  and  a66874a );
 a66879a <=( a66878a  and  a66871a );
 a66883a <=( A266  and  (not A265) );
 a66884a <=( A203  and  a66883a );
 a66887a <=( A269  and  A267 );
 a66890a <=( (not A299)  and  (not A298) );
 a66891a <=( a66890a  and  a66887a );
 a66892a <=( a66891a  and  a66884a );
 a66896a <=( (not A167)  and  A168 );
 a66897a <=( A169  and  a66896a );
 a66900a <=( (not A199)  and  A166 );
 a66903a <=( A201  and  A200 );
 a66904a <=( a66903a  and  a66900a );
 a66905a <=( a66904a  and  a66897a );
 a66909a <=( (not A266)  and  A265 );
 a66910a <=( A203  and  a66909a );
 a66913a <=( A268  and  A267 );
 a66916a <=( A301  and  (not A300) );
 a66917a <=( a66916a  and  a66913a );
 a66918a <=( a66917a  and  a66910a );
 a66922a <=( (not A167)  and  A168 );
 a66923a <=( A169  and  a66922a );
 a66926a <=( (not A199)  and  A166 );
 a66929a <=( A201  and  A200 );
 a66930a <=( a66929a  and  a66926a );
 a66931a <=( a66930a  and  a66923a );
 a66935a <=( (not A266)  and  A265 );
 a66936a <=( A203  and  a66935a );
 a66939a <=( A268  and  A267 );
 a66942a <=( A302  and  (not A300) );
 a66943a <=( a66942a  and  a66939a );
 a66944a <=( a66943a  and  a66936a );
 a66948a <=( (not A167)  and  A168 );
 a66949a <=( A169  and  a66948a );
 a66952a <=( (not A199)  and  A166 );
 a66955a <=( A201  and  A200 );
 a66956a <=( a66955a  and  a66952a );
 a66957a <=( a66956a  and  a66949a );
 a66961a <=( (not A266)  and  A265 );
 a66962a <=( A203  and  a66961a );
 a66965a <=( A268  and  A267 );
 a66968a <=( A299  and  A298 );
 a66969a <=( a66968a  and  a66965a );
 a66970a <=( a66969a  and  a66962a );
 a66974a <=( (not A167)  and  A168 );
 a66975a <=( A169  and  a66974a );
 a66978a <=( (not A199)  and  A166 );
 a66981a <=( A201  and  A200 );
 a66982a <=( a66981a  and  a66978a );
 a66983a <=( a66982a  and  a66975a );
 a66987a <=( (not A266)  and  A265 );
 a66988a <=( A203  and  a66987a );
 a66991a <=( A268  and  A267 );
 a66994a <=( (not A299)  and  (not A298) );
 a66995a <=( a66994a  and  a66991a );
 a66996a <=( a66995a  and  a66988a );
 a67000a <=( (not A167)  and  A168 );
 a67001a <=( A169  and  a67000a );
 a67004a <=( (not A199)  and  A166 );
 a67007a <=( A201  and  A200 );
 a67008a <=( a67007a  and  a67004a );
 a67009a <=( a67008a  and  a67001a );
 a67013a <=( (not A266)  and  A265 );
 a67014a <=( A203  and  a67013a );
 a67017a <=( A269  and  A267 );
 a67020a <=( A301  and  (not A300) );
 a67021a <=( a67020a  and  a67017a );
 a67022a <=( a67021a  and  a67014a );
 a67026a <=( (not A167)  and  A168 );
 a67027a <=( A169  and  a67026a );
 a67030a <=( (not A199)  and  A166 );
 a67033a <=( A201  and  A200 );
 a67034a <=( a67033a  and  a67030a );
 a67035a <=( a67034a  and  a67027a );
 a67039a <=( (not A266)  and  A265 );
 a67040a <=( A203  and  a67039a );
 a67043a <=( A269  and  A267 );
 a67046a <=( A302  and  (not A300) );
 a67047a <=( a67046a  and  a67043a );
 a67048a <=( a67047a  and  a67040a );
 a67052a <=( (not A167)  and  A168 );
 a67053a <=( A169  and  a67052a );
 a67056a <=( (not A199)  and  A166 );
 a67059a <=( A201  and  A200 );
 a67060a <=( a67059a  and  a67056a );
 a67061a <=( a67060a  and  a67053a );
 a67065a <=( (not A266)  and  A265 );
 a67066a <=( A203  and  a67065a );
 a67069a <=( A269  and  A267 );
 a67072a <=( A299  and  A298 );
 a67073a <=( a67072a  and  a67069a );
 a67074a <=( a67073a  and  a67066a );
 a67078a <=( (not A167)  and  A168 );
 a67079a <=( A169  and  a67078a );
 a67082a <=( (not A199)  and  A166 );
 a67085a <=( A201  and  A200 );
 a67086a <=( a67085a  and  a67082a );
 a67087a <=( a67086a  and  a67079a );
 a67091a <=( (not A266)  and  A265 );
 a67092a <=( A203  and  a67091a );
 a67095a <=( A269  and  A267 );
 a67098a <=( (not A299)  and  (not A298) );
 a67099a <=( a67098a  and  a67095a );
 a67100a <=( a67099a  and  a67092a );
 a67104a <=( (not A167)  and  A168 );
 a67105a <=( A169  and  a67104a );
 a67108a <=( A199  and  A166 );
 a67111a <=( A201  and  (not A200) );
 a67112a <=( a67111a  and  a67108a );
 a67113a <=( a67112a  and  a67105a );
 a67117a <=( A266  and  (not A265) );
 a67118a <=( A202  and  a67117a );
 a67121a <=( A268  and  A267 );
 a67124a <=( A301  and  (not A300) );
 a67125a <=( a67124a  and  a67121a );
 a67126a <=( a67125a  and  a67118a );
 a67130a <=( (not A167)  and  A168 );
 a67131a <=( A169  and  a67130a );
 a67134a <=( A199  and  A166 );
 a67137a <=( A201  and  (not A200) );
 a67138a <=( a67137a  and  a67134a );
 a67139a <=( a67138a  and  a67131a );
 a67143a <=( A266  and  (not A265) );
 a67144a <=( A202  and  a67143a );
 a67147a <=( A268  and  A267 );
 a67150a <=( A302  and  (not A300) );
 a67151a <=( a67150a  and  a67147a );
 a67152a <=( a67151a  and  a67144a );
 a67156a <=( (not A167)  and  A168 );
 a67157a <=( A169  and  a67156a );
 a67160a <=( A199  and  A166 );
 a67163a <=( A201  and  (not A200) );
 a67164a <=( a67163a  and  a67160a );
 a67165a <=( a67164a  and  a67157a );
 a67169a <=( A266  and  (not A265) );
 a67170a <=( A202  and  a67169a );
 a67173a <=( A268  and  A267 );
 a67176a <=( A299  and  A298 );
 a67177a <=( a67176a  and  a67173a );
 a67178a <=( a67177a  and  a67170a );
 a67182a <=( (not A167)  and  A168 );
 a67183a <=( A169  and  a67182a );
 a67186a <=( A199  and  A166 );
 a67189a <=( A201  and  (not A200) );
 a67190a <=( a67189a  and  a67186a );
 a67191a <=( a67190a  and  a67183a );
 a67195a <=( A266  and  (not A265) );
 a67196a <=( A202  and  a67195a );
 a67199a <=( A268  and  A267 );
 a67202a <=( (not A299)  and  (not A298) );
 a67203a <=( a67202a  and  a67199a );
 a67204a <=( a67203a  and  a67196a );
 a67208a <=( (not A167)  and  A168 );
 a67209a <=( A169  and  a67208a );
 a67212a <=( A199  and  A166 );
 a67215a <=( A201  and  (not A200) );
 a67216a <=( a67215a  and  a67212a );
 a67217a <=( a67216a  and  a67209a );
 a67221a <=( A266  and  (not A265) );
 a67222a <=( A202  and  a67221a );
 a67225a <=( A269  and  A267 );
 a67228a <=( A301  and  (not A300) );
 a67229a <=( a67228a  and  a67225a );
 a67230a <=( a67229a  and  a67222a );
 a67234a <=( (not A167)  and  A168 );
 a67235a <=( A169  and  a67234a );
 a67238a <=( A199  and  A166 );
 a67241a <=( A201  and  (not A200) );
 a67242a <=( a67241a  and  a67238a );
 a67243a <=( a67242a  and  a67235a );
 a67247a <=( A266  and  (not A265) );
 a67248a <=( A202  and  a67247a );
 a67251a <=( A269  and  A267 );
 a67254a <=( A302  and  (not A300) );
 a67255a <=( a67254a  and  a67251a );
 a67256a <=( a67255a  and  a67248a );
 a67260a <=( (not A167)  and  A168 );
 a67261a <=( A169  and  a67260a );
 a67264a <=( A199  and  A166 );
 a67267a <=( A201  and  (not A200) );
 a67268a <=( a67267a  and  a67264a );
 a67269a <=( a67268a  and  a67261a );
 a67273a <=( A266  and  (not A265) );
 a67274a <=( A202  and  a67273a );
 a67277a <=( A269  and  A267 );
 a67280a <=( A299  and  A298 );
 a67281a <=( a67280a  and  a67277a );
 a67282a <=( a67281a  and  a67274a );
 a67286a <=( (not A167)  and  A168 );
 a67287a <=( A169  and  a67286a );
 a67290a <=( A199  and  A166 );
 a67293a <=( A201  and  (not A200) );
 a67294a <=( a67293a  and  a67290a );
 a67295a <=( a67294a  and  a67287a );
 a67299a <=( A266  and  (not A265) );
 a67300a <=( A202  and  a67299a );
 a67303a <=( A269  and  A267 );
 a67306a <=( (not A299)  and  (not A298) );
 a67307a <=( a67306a  and  a67303a );
 a67308a <=( a67307a  and  a67300a );
 a67312a <=( (not A167)  and  A168 );
 a67313a <=( A169  and  a67312a );
 a67316a <=( A199  and  A166 );
 a67319a <=( A201  and  (not A200) );
 a67320a <=( a67319a  and  a67316a );
 a67321a <=( a67320a  and  a67313a );
 a67325a <=( (not A266)  and  A265 );
 a67326a <=( A202  and  a67325a );
 a67329a <=( A268  and  A267 );
 a67332a <=( A301  and  (not A300) );
 a67333a <=( a67332a  and  a67329a );
 a67334a <=( a67333a  and  a67326a );
 a67338a <=( (not A167)  and  A168 );
 a67339a <=( A169  and  a67338a );
 a67342a <=( A199  and  A166 );
 a67345a <=( A201  and  (not A200) );
 a67346a <=( a67345a  and  a67342a );
 a67347a <=( a67346a  and  a67339a );
 a67351a <=( (not A266)  and  A265 );
 a67352a <=( A202  and  a67351a );
 a67355a <=( A268  and  A267 );
 a67358a <=( A302  and  (not A300) );
 a67359a <=( a67358a  and  a67355a );
 a67360a <=( a67359a  and  a67352a );
 a67364a <=( (not A167)  and  A168 );
 a67365a <=( A169  and  a67364a );
 a67368a <=( A199  and  A166 );
 a67371a <=( A201  and  (not A200) );
 a67372a <=( a67371a  and  a67368a );
 a67373a <=( a67372a  and  a67365a );
 a67377a <=( (not A266)  and  A265 );
 a67378a <=( A202  and  a67377a );
 a67381a <=( A268  and  A267 );
 a67384a <=( A299  and  A298 );
 a67385a <=( a67384a  and  a67381a );
 a67386a <=( a67385a  and  a67378a );
 a67390a <=( (not A167)  and  A168 );
 a67391a <=( A169  and  a67390a );
 a67394a <=( A199  and  A166 );
 a67397a <=( A201  and  (not A200) );
 a67398a <=( a67397a  and  a67394a );
 a67399a <=( a67398a  and  a67391a );
 a67403a <=( (not A266)  and  A265 );
 a67404a <=( A202  and  a67403a );
 a67407a <=( A268  and  A267 );
 a67410a <=( (not A299)  and  (not A298) );
 a67411a <=( a67410a  and  a67407a );
 a67412a <=( a67411a  and  a67404a );
 a67416a <=( (not A167)  and  A168 );
 a67417a <=( A169  and  a67416a );
 a67420a <=( A199  and  A166 );
 a67423a <=( A201  and  (not A200) );
 a67424a <=( a67423a  and  a67420a );
 a67425a <=( a67424a  and  a67417a );
 a67429a <=( (not A266)  and  A265 );
 a67430a <=( A202  and  a67429a );
 a67433a <=( A269  and  A267 );
 a67436a <=( A301  and  (not A300) );
 a67437a <=( a67436a  and  a67433a );
 a67438a <=( a67437a  and  a67430a );
 a67442a <=( (not A167)  and  A168 );
 a67443a <=( A169  and  a67442a );
 a67446a <=( A199  and  A166 );
 a67449a <=( A201  and  (not A200) );
 a67450a <=( a67449a  and  a67446a );
 a67451a <=( a67450a  and  a67443a );
 a67455a <=( (not A266)  and  A265 );
 a67456a <=( A202  and  a67455a );
 a67459a <=( A269  and  A267 );
 a67462a <=( A302  and  (not A300) );
 a67463a <=( a67462a  and  a67459a );
 a67464a <=( a67463a  and  a67456a );
 a67468a <=( (not A167)  and  A168 );
 a67469a <=( A169  and  a67468a );
 a67472a <=( A199  and  A166 );
 a67475a <=( A201  and  (not A200) );
 a67476a <=( a67475a  and  a67472a );
 a67477a <=( a67476a  and  a67469a );
 a67481a <=( (not A266)  and  A265 );
 a67482a <=( A202  and  a67481a );
 a67485a <=( A269  and  A267 );
 a67488a <=( A299  and  A298 );
 a67489a <=( a67488a  and  a67485a );
 a67490a <=( a67489a  and  a67482a );
 a67494a <=( (not A167)  and  A168 );
 a67495a <=( A169  and  a67494a );
 a67498a <=( A199  and  A166 );
 a67501a <=( A201  and  (not A200) );
 a67502a <=( a67501a  and  a67498a );
 a67503a <=( a67502a  and  a67495a );
 a67507a <=( (not A266)  and  A265 );
 a67508a <=( A202  and  a67507a );
 a67511a <=( A269  and  A267 );
 a67514a <=( (not A299)  and  (not A298) );
 a67515a <=( a67514a  and  a67511a );
 a67516a <=( a67515a  and  a67508a );
 a67520a <=( (not A167)  and  A168 );
 a67521a <=( A169  and  a67520a );
 a67524a <=( A199  and  A166 );
 a67527a <=( A201  and  (not A200) );
 a67528a <=( a67527a  and  a67524a );
 a67529a <=( a67528a  and  a67521a );
 a67533a <=( A266  and  (not A265) );
 a67534a <=( A203  and  a67533a );
 a67537a <=( A268  and  A267 );
 a67540a <=( A301  and  (not A300) );
 a67541a <=( a67540a  and  a67537a );
 a67542a <=( a67541a  and  a67534a );
 a67546a <=( (not A167)  and  A168 );
 a67547a <=( A169  and  a67546a );
 a67550a <=( A199  and  A166 );
 a67553a <=( A201  and  (not A200) );
 a67554a <=( a67553a  and  a67550a );
 a67555a <=( a67554a  and  a67547a );
 a67559a <=( A266  and  (not A265) );
 a67560a <=( A203  and  a67559a );
 a67563a <=( A268  and  A267 );
 a67566a <=( A302  and  (not A300) );
 a67567a <=( a67566a  and  a67563a );
 a67568a <=( a67567a  and  a67560a );
 a67572a <=( (not A167)  and  A168 );
 a67573a <=( A169  and  a67572a );
 a67576a <=( A199  and  A166 );
 a67579a <=( A201  and  (not A200) );
 a67580a <=( a67579a  and  a67576a );
 a67581a <=( a67580a  and  a67573a );
 a67585a <=( A266  and  (not A265) );
 a67586a <=( A203  and  a67585a );
 a67589a <=( A268  and  A267 );
 a67592a <=( A299  and  A298 );
 a67593a <=( a67592a  and  a67589a );
 a67594a <=( a67593a  and  a67586a );
 a67598a <=( (not A167)  and  A168 );
 a67599a <=( A169  and  a67598a );
 a67602a <=( A199  and  A166 );
 a67605a <=( A201  and  (not A200) );
 a67606a <=( a67605a  and  a67602a );
 a67607a <=( a67606a  and  a67599a );
 a67611a <=( A266  and  (not A265) );
 a67612a <=( A203  and  a67611a );
 a67615a <=( A268  and  A267 );
 a67618a <=( (not A299)  and  (not A298) );
 a67619a <=( a67618a  and  a67615a );
 a67620a <=( a67619a  and  a67612a );
 a67624a <=( (not A167)  and  A168 );
 a67625a <=( A169  and  a67624a );
 a67628a <=( A199  and  A166 );
 a67631a <=( A201  and  (not A200) );
 a67632a <=( a67631a  and  a67628a );
 a67633a <=( a67632a  and  a67625a );
 a67637a <=( A266  and  (not A265) );
 a67638a <=( A203  and  a67637a );
 a67641a <=( A269  and  A267 );
 a67644a <=( A301  and  (not A300) );
 a67645a <=( a67644a  and  a67641a );
 a67646a <=( a67645a  and  a67638a );
 a67650a <=( (not A167)  and  A168 );
 a67651a <=( A169  and  a67650a );
 a67654a <=( A199  and  A166 );
 a67657a <=( A201  and  (not A200) );
 a67658a <=( a67657a  and  a67654a );
 a67659a <=( a67658a  and  a67651a );
 a67663a <=( A266  and  (not A265) );
 a67664a <=( A203  and  a67663a );
 a67667a <=( A269  and  A267 );
 a67670a <=( A302  and  (not A300) );
 a67671a <=( a67670a  and  a67667a );
 a67672a <=( a67671a  and  a67664a );
 a67676a <=( (not A167)  and  A168 );
 a67677a <=( A169  and  a67676a );
 a67680a <=( A199  and  A166 );
 a67683a <=( A201  and  (not A200) );
 a67684a <=( a67683a  and  a67680a );
 a67685a <=( a67684a  and  a67677a );
 a67689a <=( A266  and  (not A265) );
 a67690a <=( A203  and  a67689a );
 a67693a <=( A269  and  A267 );
 a67696a <=( A299  and  A298 );
 a67697a <=( a67696a  and  a67693a );
 a67698a <=( a67697a  and  a67690a );
 a67702a <=( (not A167)  and  A168 );
 a67703a <=( A169  and  a67702a );
 a67706a <=( A199  and  A166 );
 a67709a <=( A201  and  (not A200) );
 a67710a <=( a67709a  and  a67706a );
 a67711a <=( a67710a  and  a67703a );
 a67715a <=( A266  and  (not A265) );
 a67716a <=( A203  and  a67715a );
 a67719a <=( A269  and  A267 );
 a67722a <=( (not A299)  and  (not A298) );
 a67723a <=( a67722a  and  a67719a );
 a67724a <=( a67723a  and  a67716a );
 a67728a <=( (not A167)  and  A168 );
 a67729a <=( A169  and  a67728a );
 a67732a <=( A199  and  A166 );
 a67735a <=( A201  and  (not A200) );
 a67736a <=( a67735a  and  a67732a );
 a67737a <=( a67736a  and  a67729a );
 a67741a <=( (not A266)  and  A265 );
 a67742a <=( A203  and  a67741a );
 a67745a <=( A268  and  A267 );
 a67748a <=( A301  and  (not A300) );
 a67749a <=( a67748a  and  a67745a );
 a67750a <=( a67749a  and  a67742a );
 a67754a <=( (not A167)  and  A168 );
 a67755a <=( A169  and  a67754a );
 a67758a <=( A199  and  A166 );
 a67761a <=( A201  and  (not A200) );
 a67762a <=( a67761a  and  a67758a );
 a67763a <=( a67762a  and  a67755a );
 a67767a <=( (not A266)  and  A265 );
 a67768a <=( A203  and  a67767a );
 a67771a <=( A268  and  A267 );
 a67774a <=( A302  and  (not A300) );
 a67775a <=( a67774a  and  a67771a );
 a67776a <=( a67775a  and  a67768a );
 a67780a <=( (not A167)  and  A168 );
 a67781a <=( A169  and  a67780a );
 a67784a <=( A199  and  A166 );
 a67787a <=( A201  and  (not A200) );
 a67788a <=( a67787a  and  a67784a );
 a67789a <=( a67788a  and  a67781a );
 a67793a <=( (not A266)  and  A265 );
 a67794a <=( A203  and  a67793a );
 a67797a <=( A268  and  A267 );
 a67800a <=( A299  and  A298 );
 a67801a <=( a67800a  and  a67797a );
 a67802a <=( a67801a  and  a67794a );
 a67806a <=( (not A167)  and  A168 );
 a67807a <=( A169  and  a67806a );
 a67810a <=( A199  and  A166 );
 a67813a <=( A201  and  (not A200) );
 a67814a <=( a67813a  and  a67810a );
 a67815a <=( a67814a  and  a67807a );
 a67819a <=( (not A266)  and  A265 );
 a67820a <=( A203  and  a67819a );
 a67823a <=( A268  and  A267 );
 a67826a <=( (not A299)  and  (not A298) );
 a67827a <=( a67826a  and  a67823a );
 a67828a <=( a67827a  and  a67820a );
 a67832a <=( (not A167)  and  A168 );
 a67833a <=( A169  and  a67832a );
 a67836a <=( A199  and  A166 );
 a67839a <=( A201  and  (not A200) );
 a67840a <=( a67839a  and  a67836a );
 a67841a <=( a67840a  and  a67833a );
 a67845a <=( (not A266)  and  A265 );
 a67846a <=( A203  and  a67845a );
 a67849a <=( A269  and  A267 );
 a67852a <=( A301  and  (not A300) );
 a67853a <=( a67852a  and  a67849a );
 a67854a <=( a67853a  and  a67846a );
 a67858a <=( (not A167)  and  A168 );
 a67859a <=( A169  and  a67858a );
 a67862a <=( A199  and  A166 );
 a67865a <=( A201  and  (not A200) );
 a67866a <=( a67865a  and  a67862a );
 a67867a <=( a67866a  and  a67859a );
 a67871a <=( (not A266)  and  A265 );
 a67872a <=( A203  and  a67871a );
 a67875a <=( A269  and  A267 );
 a67878a <=( A302  and  (not A300) );
 a67879a <=( a67878a  and  a67875a );
 a67880a <=( a67879a  and  a67872a );
 a67884a <=( (not A167)  and  A168 );
 a67885a <=( A169  and  a67884a );
 a67888a <=( A199  and  A166 );
 a67891a <=( A201  and  (not A200) );
 a67892a <=( a67891a  and  a67888a );
 a67893a <=( a67892a  and  a67885a );
 a67897a <=( (not A266)  and  A265 );
 a67898a <=( A203  and  a67897a );
 a67901a <=( A269  and  A267 );
 a67904a <=( A299  and  A298 );
 a67905a <=( a67904a  and  a67901a );
 a67906a <=( a67905a  and  a67898a );
 a67910a <=( (not A167)  and  A168 );
 a67911a <=( A169  and  a67910a );
 a67914a <=( A199  and  A166 );
 a67917a <=( A201  and  (not A200) );
 a67918a <=( a67917a  and  a67914a );
 a67919a <=( a67918a  and  a67911a );
 a67923a <=( (not A266)  and  A265 );
 a67924a <=( A203  and  a67923a );
 a67927a <=( A269  and  A267 );
 a67930a <=( (not A299)  and  (not A298) );
 a67931a <=( a67930a  and  a67927a );
 a67932a <=( a67931a  and  a67924a );
 a67936a <=( (not A167)  and  A168 );
 a67937a <=( A169  and  a67936a );
 a67940a <=( (not A199)  and  A166 );
 a67943a <=( A267  and  (not A200) );
 a67944a <=( a67943a  and  a67940a );
 a67945a <=( a67944a  and  a67937a );
 a67949a <=( A298  and  (not A269) );
 a67950a <=( (not A268)  and  a67949a );
 a67953a <=( (not A300)  and  (not A299) );
 a67956a <=( (not A302)  and  (not A301) );
 a67957a <=( a67956a  and  a67953a );
 a67958a <=( a67957a  and  a67950a );
 a67962a <=( (not A167)  and  A168 );
 a67963a <=( A169  and  a67962a );
 a67966a <=( (not A199)  and  A166 );
 a67969a <=( A267  and  (not A200) );
 a67970a <=( a67969a  and  a67966a );
 a67971a <=( a67970a  and  a67963a );
 a67975a <=( (not A298)  and  (not A269) );
 a67976a <=( (not A268)  and  a67975a );
 a67979a <=( (not A300)  and  A299 );
 a67982a <=( (not A302)  and  (not A301) );
 a67983a <=( a67982a  and  a67979a );
 a67984a <=( a67983a  and  a67976a );
 a67988a <=( (not A199)  and  (not A168) );
 a67989a <=( A169  and  a67988a );
 a67992a <=( A201  and  A200 );
 a67995a <=( A267  and  A202 );
 a67996a <=( a67995a  and  a67992a );
 a67997a <=( a67996a  and  a67989a );
 a68001a <=( A298  and  (not A269) );
 a68002a <=( (not A268)  and  a68001a );
 a68005a <=( (not A300)  and  (not A299) );
 a68008a <=( (not A302)  and  (not A301) );
 a68009a <=( a68008a  and  a68005a );
 a68010a <=( a68009a  and  a68002a );
 a68014a <=( (not A199)  and  (not A168) );
 a68015a <=( A169  and  a68014a );
 a68018a <=( A201  and  A200 );
 a68021a <=( A267  and  A202 );
 a68022a <=( a68021a  and  a68018a );
 a68023a <=( a68022a  and  a68015a );
 a68027a <=( (not A298)  and  (not A269) );
 a68028a <=( (not A268)  and  a68027a );
 a68031a <=( (not A300)  and  A299 );
 a68034a <=( (not A302)  and  (not A301) );
 a68035a <=( a68034a  and  a68031a );
 a68036a <=( a68035a  and  a68028a );
 a68040a <=( (not A199)  and  (not A168) );
 a68041a <=( A169  and  a68040a );
 a68044a <=( A201  and  A200 );
 a68047a <=( A267  and  A203 );
 a68048a <=( a68047a  and  a68044a );
 a68049a <=( a68048a  and  a68041a );
 a68053a <=( A298  and  (not A269) );
 a68054a <=( (not A268)  and  a68053a );
 a68057a <=( (not A300)  and  (not A299) );
 a68060a <=( (not A302)  and  (not A301) );
 a68061a <=( a68060a  and  a68057a );
 a68062a <=( a68061a  and  a68054a );
 a68066a <=( (not A199)  and  (not A168) );
 a68067a <=( A169  and  a68066a );
 a68070a <=( A201  and  A200 );
 a68073a <=( A267  and  A203 );
 a68074a <=( a68073a  and  a68070a );
 a68075a <=( a68074a  and  a68067a );
 a68079a <=( (not A298)  and  (not A269) );
 a68080a <=( (not A268)  and  a68079a );
 a68083a <=( (not A300)  and  A299 );
 a68086a <=( (not A302)  and  (not A301) );
 a68087a <=( a68086a  and  a68083a );
 a68088a <=( a68087a  and  a68080a );
 a68092a <=( (not A199)  and  (not A168) );
 a68093a <=( A169  and  a68092a );
 a68096a <=( (not A201)  and  A200 );
 a68099a <=( (not A203)  and  (not A202) );
 a68100a <=( a68099a  and  a68096a );
 a68101a <=( a68100a  and  a68093a );
 a68105a <=( (not A269)  and  (not A268) );
 a68106a <=( A267  and  a68105a );
 a68109a <=( (not A299)  and  A298 );
 a68112a <=( A301  and  A300 );
 a68113a <=( a68112a  and  a68109a );
 a68114a <=( a68113a  and  a68106a );
 a68118a <=( (not A199)  and  (not A168) );
 a68119a <=( A169  and  a68118a );
 a68122a <=( (not A201)  and  A200 );
 a68125a <=( (not A203)  and  (not A202) );
 a68126a <=( a68125a  and  a68122a );
 a68127a <=( a68126a  and  a68119a );
 a68131a <=( (not A269)  and  (not A268) );
 a68132a <=( A267  and  a68131a );
 a68135a <=( (not A299)  and  A298 );
 a68138a <=( A302  and  A300 );
 a68139a <=( a68138a  and  a68135a );
 a68140a <=( a68139a  and  a68132a );
 a68144a <=( (not A199)  and  (not A168) );
 a68145a <=( A169  and  a68144a );
 a68148a <=( (not A201)  and  A200 );
 a68151a <=( (not A203)  and  (not A202) );
 a68152a <=( a68151a  and  a68148a );
 a68153a <=( a68152a  and  a68145a );
 a68157a <=( (not A269)  and  (not A268) );
 a68158a <=( A267  and  a68157a );
 a68161a <=( A299  and  (not A298) );
 a68164a <=( A301  and  A300 );
 a68165a <=( a68164a  and  a68161a );
 a68166a <=( a68165a  and  a68158a );
 a68170a <=( (not A199)  and  (not A168) );
 a68171a <=( A169  and  a68170a );
 a68174a <=( (not A201)  and  A200 );
 a68177a <=( (not A203)  and  (not A202) );
 a68178a <=( a68177a  and  a68174a );
 a68179a <=( a68178a  and  a68171a );
 a68183a <=( (not A269)  and  (not A268) );
 a68184a <=( A267  and  a68183a );
 a68187a <=( A299  and  (not A298) );
 a68190a <=( A302  and  A300 );
 a68191a <=( a68190a  and  a68187a );
 a68192a <=( a68191a  and  a68184a );
 a68196a <=( (not A199)  and  (not A168) );
 a68197a <=( A169  and  a68196a );
 a68200a <=( (not A201)  and  A200 );
 a68203a <=( (not A203)  and  (not A202) );
 a68204a <=( a68203a  and  a68200a );
 a68205a <=( a68204a  and  a68197a );
 a68209a <=( A298  and  A268 );
 a68210a <=( (not A267)  and  a68209a );
 a68213a <=( (not A300)  and  (not A299) );
 a68216a <=( (not A302)  and  (not A301) );
 a68217a <=( a68216a  and  a68213a );
 a68218a <=( a68217a  and  a68210a );
 a68222a <=( (not A199)  and  (not A168) );
 a68223a <=( A169  and  a68222a );
 a68226a <=( (not A201)  and  A200 );
 a68229a <=( (not A203)  and  (not A202) );
 a68230a <=( a68229a  and  a68226a );
 a68231a <=( a68230a  and  a68223a );
 a68235a <=( (not A298)  and  A268 );
 a68236a <=( (not A267)  and  a68235a );
 a68239a <=( (not A300)  and  A299 );
 a68242a <=( (not A302)  and  (not A301) );
 a68243a <=( a68242a  and  a68239a );
 a68244a <=( a68243a  and  a68236a );
 a68248a <=( (not A199)  and  (not A168) );
 a68249a <=( A169  and  a68248a );
 a68252a <=( (not A201)  and  A200 );
 a68255a <=( (not A203)  and  (not A202) );
 a68256a <=( a68255a  and  a68252a );
 a68257a <=( a68256a  and  a68249a );
 a68261a <=( A298  and  A269 );
 a68262a <=( (not A267)  and  a68261a );
 a68265a <=( (not A300)  and  (not A299) );
 a68268a <=( (not A302)  and  (not A301) );
 a68269a <=( a68268a  and  a68265a );
 a68270a <=( a68269a  and  a68262a );
 a68274a <=( (not A199)  and  (not A168) );
 a68275a <=( A169  and  a68274a );
 a68278a <=( (not A201)  and  A200 );
 a68281a <=( (not A203)  and  (not A202) );
 a68282a <=( a68281a  and  a68278a );
 a68283a <=( a68282a  and  a68275a );
 a68287a <=( (not A298)  and  A269 );
 a68288a <=( (not A267)  and  a68287a );
 a68291a <=( (not A300)  and  A299 );
 a68294a <=( (not A302)  and  (not A301) );
 a68295a <=( a68294a  and  a68291a );
 a68296a <=( a68295a  and  a68288a );
 a68300a <=( (not A199)  and  (not A168) );
 a68301a <=( A169  and  a68300a );
 a68304a <=( (not A201)  and  A200 );
 a68307a <=( (not A203)  and  (not A202) );
 a68308a <=( a68307a  and  a68304a );
 a68309a <=( a68308a  and  a68301a );
 a68313a <=( A298  and  A266 );
 a68314a <=( A265  and  a68313a );
 a68317a <=( (not A300)  and  (not A299) );
 a68320a <=( (not A302)  and  (not A301) );
 a68321a <=( a68320a  and  a68317a );
 a68322a <=( a68321a  and  a68314a );
 a68326a <=( (not A199)  and  (not A168) );
 a68327a <=( A169  and  a68326a );
 a68330a <=( (not A201)  and  A200 );
 a68333a <=( (not A203)  and  (not A202) );
 a68334a <=( a68333a  and  a68330a );
 a68335a <=( a68334a  and  a68327a );
 a68339a <=( (not A298)  and  A266 );
 a68340a <=( A265  and  a68339a );
 a68343a <=( (not A300)  and  A299 );
 a68346a <=( (not A302)  and  (not A301) );
 a68347a <=( a68346a  and  a68343a );
 a68348a <=( a68347a  and  a68340a );
 a68352a <=( (not A199)  and  (not A168) );
 a68353a <=( A169  and  a68352a );
 a68356a <=( (not A201)  and  A200 );
 a68359a <=( (not A203)  and  (not A202) );
 a68360a <=( a68359a  and  a68356a );
 a68361a <=( a68360a  and  a68353a );
 a68365a <=( A298  and  (not A266) );
 a68366a <=( (not A265)  and  a68365a );
 a68369a <=( (not A300)  and  (not A299) );
 a68372a <=( (not A302)  and  (not A301) );
 a68373a <=( a68372a  and  a68369a );
 a68374a <=( a68373a  and  a68366a );
 a68378a <=( (not A199)  and  (not A168) );
 a68379a <=( A169  and  a68378a );
 a68382a <=( (not A201)  and  A200 );
 a68385a <=( (not A203)  and  (not A202) );
 a68386a <=( a68385a  and  a68382a );
 a68387a <=( a68386a  and  a68379a );
 a68391a <=( (not A298)  and  (not A266) );
 a68392a <=( (not A265)  and  a68391a );
 a68395a <=( (not A300)  and  A299 );
 a68398a <=( (not A302)  and  (not A301) );
 a68399a <=( a68398a  and  a68395a );
 a68400a <=( a68399a  and  a68392a );
 a68404a <=( A199  and  (not A168) );
 a68405a <=( A169  and  a68404a );
 a68408a <=( A201  and  (not A200) );
 a68411a <=( A267  and  A202 );
 a68412a <=( a68411a  and  a68408a );
 a68413a <=( a68412a  and  a68405a );
 a68417a <=( A298  and  (not A269) );
 a68418a <=( (not A268)  and  a68417a );
 a68421a <=( (not A300)  and  (not A299) );
 a68424a <=( (not A302)  and  (not A301) );
 a68425a <=( a68424a  and  a68421a );
 a68426a <=( a68425a  and  a68418a );
 a68430a <=( A199  and  (not A168) );
 a68431a <=( A169  and  a68430a );
 a68434a <=( A201  and  (not A200) );
 a68437a <=( A267  and  A202 );
 a68438a <=( a68437a  and  a68434a );
 a68439a <=( a68438a  and  a68431a );
 a68443a <=( (not A298)  and  (not A269) );
 a68444a <=( (not A268)  and  a68443a );
 a68447a <=( (not A300)  and  A299 );
 a68450a <=( (not A302)  and  (not A301) );
 a68451a <=( a68450a  and  a68447a );
 a68452a <=( a68451a  and  a68444a );
 a68456a <=( A199  and  (not A168) );
 a68457a <=( A169  and  a68456a );
 a68460a <=( A201  and  (not A200) );
 a68463a <=( A267  and  A203 );
 a68464a <=( a68463a  and  a68460a );
 a68465a <=( a68464a  and  a68457a );
 a68469a <=( A298  and  (not A269) );
 a68470a <=( (not A268)  and  a68469a );
 a68473a <=( (not A300)  and  (not A299) );
 a68476a <=( (not A302)  and  (not A301) );
 a68477a <=( a68476a  and  a68473a );
 a68478a <=( a68477a  and  a68470a );
 a68482a <=( A199  and  (not A168) );
 a68483a <=( A169  and  a68482a );
 a68486a <=( A201  and  (not A200) );
 a68489a <=( A267  and  A203 );
 a68490a <=( a68489a  and  a68486a );
 a68491a <=( a68490a  and  a68483a );
 a68495a <=( (not A298)  and  (not A269) );
 a68496a <=( (not A268)  and  a68495a );
 a68499a <=( (not A300)  and  A299 );
 a68502a <=( (not A302)  and  (not A301) );
 a68503a <=( a68502a  and  a68499a );
 a68504a <=( a68503a  and  a68496a );
 a68508a <=( A199  and  (not A168) );
 a68509a <=( A169  and  a68508a );
 a68512a <=( (not A201)  and  (not A200) );
 a68515a <=( (not A203)  and  (not A202) );
 a68516a <=( a68515a  and  a68512a );
 a68517a <=( a68516a  and  a68509a );
 a68521a <=( (not A269)  and  (not A268) );
 a68522a <=( A267  and  a68521a );
 a68525a <=( (not A299)  and  A298 );
 a68528a <=( A301  and  A300 );
 a68529a <=( a68528a  and  a68525a );
 a68530a <=( a68529a  and  a68522a );
 a68534a <=( A199  and  (not A168) );
 a68535a <=( A169  and  a68534a );
 a68538a <=( (not A201)  and  (not A200) );
 a68541a <=( (not A203)  and  (not A202) );
 a68542a <=( a68541a  and  a68538a );
 a68543a <=( a68542a  and  a68535a );
 a68547a <=( (not A269)  and  (not A268) );
 a68548a <=( A267  and  a68547a );
 a68551a <=( (not A299)  and  A298 );
 a68554a <=( A302  and  A300 );
 a68555a <=( a68554a  and  a68551a );
 a68556a <=( a68555a  and  a68548a );
 a68560a <=( A199  and  (not A168) );
 a68561a <=( A169  and  a68560a );
 a68564a <=( (not A201)  and  (not A200) );
 a68567a <=( (not A203)  and  (not A202) );
 a68568a <=( a68567a  and  a68564a );
 a68569a <=( a68568a  and  a68561a );
 a68573a <=( (not A269)  and  (not A268) );
 a68574a <=( A267  and  a68573a );
 a68577a <=( A299  and  (not A298) );
 a68580a <=( A301  and  A300 );
 a68581a <=( a68580a  and  a68577a );
 a68582a <=( a68581a  and  a68574a );
 a68586a <=( A199  and  (not A168) );
 a68587a <=( A169  and  a68586a );
 a68590a <=( (not A201)  and  (not A200) );
 a68593a <=( (not A203)  and  (not A202) );
 a68594a <=( a68593a  and  a68590a );
 a68595a <=( a68594a  and  a68587a );
 a68599a <=( (not A269)  and  (not A268) );
 a68600a <=( A267  and  a68599a );
 a68603a <=( A299  and  (not A298) );
 a68606a <=( A302  and  A300 );
 a68607a <=( a68606a  and  a68603a );
 a68608a <=( a68607a  and  a68600a );
 a68612a <=( A199  and  (not A168) );
 a68613a <=( A169  and  a68612a );
 a68616a <=( (not A201)  and  (not A200) );
 a68619a <=( (not A203)  and  (not A202) );
 a68620a <=( a68619a  and  a68616a );
 a68621a <=( a68620a  and  a68613a );
 a68625a <=( A298  and  A268 );
 a68626a <=( (not A267)  and  a68625a );
 a68629a <=( (not A300)  and  (not A299) );
 a68632a <=( (not A302)  and  (not A301) );
 a68633a <=( a68632a  and  a68629a );
 a68634a <=( a68633a  and  a68626a );
 a68638a <=( A199  and  (not A168) );
 a68639a <=( A169  and  a68638a );
 a68642a <=( (not A201)  and  (not A200) );
 a68645a <=( (not A203)  and  (not A202) );
 a68646a <=( a68645a  and  a68642a );
 a68647a <=( a68646a  and  a68639a );
 a68651a <=( (not A298)  and  A268 );
 a68652a <=( (not A267)  and  a68651a );
 a68655a <=( (not A300)  and  A299 );
 a68658a <=( (not A302)  and  (not A301) );
 a68659a <=( a68658a  and  a68655a );
 a68660a <=( a68659a  and  a68652a );
 a68664a <=( A199  and  (not A168) );
 a68665a <=( A169  and  a68664a );
 a68668a <=( (not A201)  and  (not A200) );
 a68671a <=( (not A203)  and  (not A202) );
 a68672a <=( a68671a  and  a68668a );
 a68673a <=( a68672a  and  a68665a );
 a68677a <=( A298  and  A269 );
 a68678a <=( (not A267)  and  a68677a );
 a68681a <=( (not A300)  and  (not A299) );
 a68684a <=( (not A302)  and  (not A301) );
 a68685a <=( a68684a  and  a68681a );
 a68686a <=( a68685a  and  a68678a );
 a68690a <=( A199  and  (not A168) );
 a68691a <=( A169  and  a68690a );
 a68694a <=( (not A201)  and  (not A200) );
 a68697a <=( (not A203)  and  (not A202) );
 a68698a <=( a68697a  and  a68694a );
 a68699a <=( a68698a  and  a68691a );
 a68703a <=( (not A298)  and  A269 );
 a68704a <=( (not A267)  and  a68703a );
 a68707a <=( (not A300)  and  A299 );
 a68710a <=( (not A302)  and  (not A301) );
 a68711a <=( a68710a  and  a68707a );
 a68712a <=( a68711a  and  a68704a );
 a68716a <=( A199  and  (not A168) );
 a68717a <=( A169  and  a68716a );
 a68720a <=( (not A201)  and  (not A200) );
 a68723a <=( (not A203)  and  (not A202) );
 a68724a <=( a68723a  and  a68720a );
 a68725a <=( a68724a  and  a68717a );
 a68729a <=( A298  and  A266 );
 a68730a <=( A265  and  a68729a );
 a68733a <=( (not A300)  and  (not A299) );
 a68736a <=( (not A302)  and  (not A301) );
 a68737a <=( a68736a  and  a68733a );
 a68738a <=( a68737a  and  a68730a );
 a68742a <=( A199  and  (not A168) );
 a68743a <=( A169  and  a68742a );
 a68746a <=( (not A201)  and  (not A200) );
 a68749a <=( (not A203)  and  (not A202) );
 a68750a <=( a68749a  and  a68746a );
 a68751a <=( a68750a  and  a68743a );
 a68755a <=( (not A298)  and  A266 );
 a68756a <=( A265  and  a68755a );
 a68759a <=( (not A300)  and  A299 );
 a68762a <=( (not A302)  and  (not A301) );
 a68763a <=( a68762a  and  a68759a );
 a68764a <=( a68763a  and  a68756a );
 a68768a <=( A199  and  (not A168) );
 a68769a <=( A169  and  a68768a );
 a68772a <=( (not A201)  and  (not A200) );
 a68775a <=( (not A203)  and  (not A202) );
 a68776a <=( a68775a  and  a68772a );
 a68777a <=( a68776a  and  a68769a );
 a68781a <=( A298  and  (not A266) );
 a68782a <=( (not A265)  and  a68781a );
 a68785a <=( (not A300)  and  (not A299) );
 a68788a <=( (not A302)  and  (not A301) );
 a68789a <=( a68788a  and  a68785a );
 a68790a <=( a68789a  and  a68782a );
 a68794a <=( A199  and  (not A168) );
 a68795a <=( A169  and  a68794a );
 a68798a <=( (not A201)  and  (not A200) );
 a68801a <=( (not A203)  and  (not A202) );
 a68802a <=( a68801a  and  a68798a );
 a68803a <=( a68802a  and  a68795a );
 a68807a <=( (not A298)  and  (not A266) );
 a68808a <=( (not A265)  and  a68807a );
 a68811a <=( (not A300)  and  A299 );
 a68814a <=( (not A302)  and  (not A301) );
 a68815a <=( a68814a  and  a68811a );
 a68816a <=( a68815a  and  a68808a );
 a68820a <=( A168  and  (not A169) );
 a68821a <=( A170  and  a68820a );
 a68824a <=( (not A202)  and  A201 );
 a68827a <=( (not A265)  and  (not A203) );
 a68828a <=( a68827a  and  a68824a );
 a68829a <=( a68828a  and  a68821a );
 a68833a <=( (not A268)  and  (not A267) );
 a68834a <=( A266  and  a68833a );
 a68837a <=( A300  and  (not A269) );
 a68840a <=( (not A302)  and  (not A301) );
 a68841a <=( a68840a  and  a68837a );
 a68842a <=( a68841a  and  a68834a );
 a68846a <=( A168  and  (not A169) );
 a68847a <=( A170  and  a68846a );
 a68850a <=( (not A202)  and  A201 );
 a68853a <=( A265  and  (not A203) );
 a68854a <=( a68853a  and  a68850a );
 a68855a <=( a68854a  and  a68847a );
 a68859a <=( (not A268)  and  (not A267) );
 a68860a <=( (not A266)  and  a68859a );
 a68863a <=( A300  and  (not A269) );
 a68866a <=( (not A302)  and  (not A301) );
 a68867a <=( a68866a  and  a68863a );
 a68868a <=( a68867a  and  a68860a );
 a68872a <=( A168  and  (not A169) );
 a68873a <=( A170  and  a68872a );
 a68876a <=( A200  and  (not A199) );
 a68879a <=( A202  and  A201 );
 a68880a <=( a68879a  and  a68876a );
 a68881a <=( a68880a  and  a68873a );
 a68885a <=( (not A269)  and  (not A268) );
 a68886a <=( A267  and  a68885a );
 a68889a <=( (not A299)  and  A298 );
 a68892a <=( A301  and  A300 );
 a68893a <=( a68892a  and  a68889a );
 a68894a <=( a68893a  and  a68886a );
 a68898a <=( A168  and  (not A169) );
 a68899a <=( A170  and  a68898a );
 a68902a <=( A200  and  (not A199) );
 a68905a <=( A202  and  A201 );
 a68906a <=( a68905a  and  a68902a );
 a68907a <=( a68906a  and  a68899a );
 a68911a <=( (not A269)  and  (not A268) );
 a68912a <=( A267  and  a68911a );
 a68915a <=( (not A299)  and  A298 );
 a68918a <=( A302  and  A300 );
 a68919a <=( a68918a  and  a68915a );
 a68920a <=( a68919a  and  a68912a );
 a68924a <=( A168  and  (not A169) );
 a68925a <=( A170  and  a68924a );
 a68928a <=( A200  and  (not A199) );
 a68931a <=( A202  and  A201 );
 a68932a <=( a68931a  and  a68928a );
 a68933a <=( a68932a  and  a68925a );
 a68937a <=( (not A269)  and  (not A268) );
 a68938a <=( A267  and  a68937a );
 a68941a <=( A299  and  (not A298) );
 a68944a <=( A301  and  A300 );
 a68945a <=( a68944a  and  a68941a );
 a68946a <=( a68945a  and  a68938a );
 a68950a <=( A168  and  (not A169) );
 a68951a <=( A170  and  a68950a );
 a68954a <=( A200  and  (not A199) );
 a68957a <=( A202  and  A201 );
 a68958a <=( a68957a  and  a68954a );
 a68959a <=( a68958a  and  a68951a );
 a68963a <=( (not A269)  and  (not A268) );
 a68964a <=( A267  and  a68963a );
 a68967a <=( A299  and  (not A298) );
 a68970a <=( A302  and  A300 );
 a68971a <=( a68970a  and  a68967a );
 a68972a <=( a68971a  and  a68964a );
 a68976a <=( A168  and  (not A169) );
 a68977a <=( A170  and  a68976a );
 a68980a <=( A200  and  (not A199) );
 a68983a <=( A202  and  A201 );
 a68984a <=( a68983a  and  a68980a );
 a68985a <=( a68984a  and  a68977a );
 a68989a <=( A298  and  A268 );
 a68990a <=( (not A267)  and  a68989a );
 a68993a <=( (not A300)  and  (not A299) );
 a68996a <=( (not A302)  and  (not A301) );
 a68997a <=( a68996a  and  a68993a );
 a68998a <=( a68997a  and  a68990a );
 a69002a <=( A168  and  (not A169) );
 a69003a <=( A170  and  a69002a );
 a69006a <=( A200  and  (not A199) );
 a69009a <=( A202  and  A201 );
 a69010a <=( a69009a  and  a69006a );
 a69011a <=( a69010a  and  a69003a );
 a69015a <=( (not A298)  and  A268 );
 a69016a <=( (not A267)  and  a69015a );
 a69019a <=( (not A300)  and  A299 );
 a69022a <=( (not A302)  and  (not A301) );
 a69023a <=( a69022a  and  a69019a );
 a69024a <=( a69023a  and  a69016a );
 a69028a <=( A168  and  (not A169) );
 a69029a <=( A170  and  a69028a );
 a69032a <=( A200  and  (not A199) );
 a69035a <=( A202  and  A201 );
 a69036a <=( a69035a  and  a69032a );
 a69037a <=( a69036a  and  a69029a );
 a69041a <=( A298  and  A269 );
 a69042a <=( (not A267)  and  a69041a );
 a69045a <=( (not A300)  and  (not A299) );
 a69048a <=( (not A302)  and  (not A301) );
 a69049a <=( a69048a  and  a69045a );
 a69050a <=( a69049a  and  a69042a );
 a69054a <=( A168  and  (not A169) );
 a69055a <=( A170  and  a69054a );
 a69058a <=( A200  and  (not A199) );
 a69061a <=( A202  and  A201 );
 a69062a <=( a69061a  and  a69058a );
 a69063a <=( a69062a  and  a69055a );
 a69067a <=( (not A298)  and  A269 );
 a69068a <=( (not A267)  and  a69067a );
 a69071a <=( (not A300)  and  A299 );
 a69074a <=( (not A302)  and  (not A301) );
 a69075a <=( a69074a  and  a69071a );
 a69076a <=( a69075a  and  a69068a );
 a69080a <=( A168  and  (not A169) );
 a69081a <=( A170  and  a69080a );
 a69084a <=( A200  and  (not A199) );
 a69087a <=( A202  and  A201 );
 a69088a <=( a69087a  and  a69084a );
 a69089a <=( a69088a  and  a69081a );
 a69093a <=( A298  and  A266 );
 a69094a <=( A265  and  a69093a );
 a69097a <=( (not A300)  and  (not A299) );
 a69100a <=( (not A302)  and  (not A301) );
 a69101a <=( a69100a  and  a69097a );
 a69102a <=( a69101a  and  a69094a );
 a69106a <=( A168  and  (not A169) );
 a69107a <=( A170  and  a69106a );
 a69110a <=( A200  and  (not A199) );
 a69113a <=( A202  and  A201 );
 a69114a <=( a69113a  and  a69110a );
 a69115a <=( a69114a  and  a69107a );
 a69119a <=( (not A298)  and  A266 );
 a69120a <=( A265  and  a69119a );
 a69123a <=( (not A300)  and  A299 );
 a69126a <=( (not A302)  and  (not A301) );
 a69127a <=( a69126a  and  a69123a );
 a69128a <=( a69127a  and  a69120a );
 a69132a <=( A168  and  (not A169) );
 a69133a <=( A170  and  a69132a );
 a69136a <=( A200  and  (not A199) );
 a69139a <=( A202  and  A201 );
 a69140a <=( a69139a  and  a69136a );
 a69141a <=( a69140a  and  a69133a );
 a69145a <=( A298  and  (not A266) );
 a69146a <=( (not A265)  and  a69145a );
 a69149a <=( (not A300)  and  (not A299) );
 a69152a <=( (not A302)  and  (not A301) );
 a69153a <=( a69152a  and  a69149a );
 a69154a <=( a69153a  and  a69146a );
 a69158a <=( A168  and  (not A169) );
 a69159a <=( A170  and  a69158a );
 a69162a <=( A200  and  (not A199) );
 a69165a <=( A202  and  A201 );
 a69166a <=( a69165a  and  a69162a );
 a69167a <=( a69166a  and  a69159a );
 a69171a <=( (not A298)  and  (not A266) );
 a69172a <=( (not A265)  and  a69171a );
 a69175a <=( (not A300)  and  A299 );
 a69178a <=( (not A302)  and  (not A301) );
 a69179a <=( a69178a  and  a69175a );
 a69180a <=( a69179a  and  a69172a );
 a69184a <=( A168  and  (not A169) );
 a69185a <=( A170  and  a69184a );
 a69188a <=( A200  and  (not A199) );
 a69191a <=( A203  and  A201 );
 a69192a <=( a69191a  and  a69188a );
 a69193a <=( a69192a  and  a69185a );
 a69197a <=( (not A269)  and  (not A268) );
 a69198a <=( A267  and  a69197a );
 a69201a <=( (not A299)  and  A298 );
 a69204a <=( A301  and  A300 );
 a69205a <=( a69204a  and  a69201a );
 a69206a <=( a69205a  and  a69198a );
 a69210a <=( A168  and  (not A169) );
 a69211a <=( A170  and  a69210a );
 a69214a <=( A200  and  (not A199) );
 a69217a <=( A203  and  A201 );
 a69218a <=( a69217a  and  a69214a );
 a69219a <=( a69218a  and  a69211a );
 a69223a <=( (not A269)  and  (not A268) );
 a69224a <=( A267  and  a69223a );
 a69227a <=( (not A299)  and  A298 );
 a69230a <=( A302  and  A300 );
 a69231a <=( a69230a  and  a69227a );
 a69232a <=( a69231a  and  a69224a );
 a69236a <=( A168  and  (not A169) );
 a69237a <=( A170  and  a69236a );
 a69240a <=( A200  and  (not A199) );
 a69243a <=( A203  and  A201 );
 a69244a <=( a69243a  and  a69240a );
 a69245a <=( a69244a  and  a69237a );
 a69249a <=( (not A269)  and  (not A268) );
 a69250a <=( A267  and  a69249a );
 a69253a <=( A299  and  (not A298) );
 a69256a <=( A301  and  A300 );
 a69257a <=( a69256a  and  a69253a );
 a69258a <=( a69257a  and  a69250a );
 a69262a <=( A168  and  (not A169) );
 a69263a <=( A170  and  a69262a );
 a69266a <=( A200  and  (not A199) );
 a69269a <=( A203  and  A201 );
 a69270a <=( a69269a  and  a69266a );
 a69271a <=( a69270a  and  a69263a );
 a69275a <=( (not A269)  and  (not A268) );
 a69276a <=( A267  and  a69275a );
 a69279a <=( A299  and  (not A298) );
 a69282a <=( A302  and  A300 );
 a69283a <=( a69282a  and  a69279a );
 a69284a <=( a69283a  and  a69276a );
 a69288a <=( A168  and  (not A169) );
 a69289a <=( A170  and  a69288a );
 a69292a <=( A200  and  (not A199) );
 a69295a <=( A203  and  A201 );
 a69296a <=( a69295a  and  a69292a );
 a69297a <=( a69296a  and  a69289a );
 a69301a <=( A298  and  A268 );
 a69302a <=( (not A267)  and  a69301a );
 a69305a <=( (not A300)  and  (not A299) );
 a69308a <=( (not A302)  and  (not A301) );
 a69309a <=( a69308a  and  a69305a );
 a69310a <=( a69309a  and  a69302a );
 a69314a <=( A168  and  (not A169) );
 a69315a <=( A170  and  a69314a );
 a69318a <=( A200  and  (not A199) );
 a69321a <=( A203  and  A201 );
 a69322a <=( a69321a  and  a69318a );
 a69323a <=( a69322a  and  a69315a );
 a69327a <=( (not A298)  and  A268 );
 a69328a <=( (not A267)  and  a69327a );
 a69331a <=( (not A300)  and  A299 );
 a69334a <=( (not A302)  and  (not A301) );
 a69335a <=( a69334a  and  a69331a );
 a69336a <=( a69335a  and  a69328a );
 a69340a <=( A168  and  (not A169) );
 a69341a <=( A170  and  a69340a );
 a69344a <=( A200  and  (not A199) );
 a69347a <=( A203  and  A201 );
 a69348a <=( a69347a  and  a69344a );
 a69349a <=( a69348a  and  a69341a );
 a69353a <=( A298  and  A269 );
 a69354a <=( (not A267)  and  a69353a );
 a69357a <=( (not A300)  and  (not A299) );
 a69360a <=( (not A302)  and  (not A301) );
 a69361a <=( a69360a  and  a69357a );
 a69362a <=( a69361a  and  a69354a );
 a69366a <=( A168  and  (not A169) );
 a69367a <=( A170  and  a69366a );
 a69370a <=( A200  and  (not A199) );
 a69373a <=( A203  and  A201 );
 a69374a <=( a69373a  and  a69370a );
 a69375a <=( a69374a  and  a69367a );
 a69379a <=( (not A298)  and  A269 );
 a69380a <=( (not A267)  and  a69379a );
 a69383a <=( (not A300)  and  A299 );
 a69386a <=( (not A302)  and  (not A301) );
 a69387a <=( a69386a  and  a69383a );
 a69388a <=( a69387a  and  a69380a );
 a69392a <=( A168  and  (not A169) );
 a69393a <=( A170  and  a69392a );
 a69396a <=( A200  and  (not A199) );
 a69399a <=( A203  and  A201 );
 a69400a <=( a69399a  and  a69396a );
 a69401a <=( a69400a  and  a69393a );
 a69405a <=( A298  and  A266 );
 a69406a <=( A265  and  a69405a );
 a69409a <=( (not A300)  and  (not A299) );
 a69412a <=( (not A302)  and  (not A301) );
 a69413a <=( a69412a  and  a69409a );
 a69414a <=( a69413a  and  a69406a );
 a69418a <=( A168  and  (not A169) );
 a69419a <=( A170  and  a69418a );
 a69422a <=( A200  and  (not A199) );
 a69425a <=( A203  and  A201 );
 a69426a <=( a69425a  and  a69422a );
 a69427a <=( a69426a  and  a69419a );
 a69431a <=( (not A298)  and  A266 );
 a69432a <=( A265  and  a69431a );
 a69435a <=( (not A300)  and  A299 );
 a69438a <=( (not A302)  and  (not A301) );
 a69439a <=( a69438a  and  a69435a );
 a69440a <=( a69439a  and  a69432a );
 a69444a <=( A168  and  (not A169) );
 a69445a <=( A170  and  a69444a );
 a69448a <=( A200  and  (not A199) );
 a69451a <=( A203  and  A201 );
 a69452a <=( a69451a  and  a69448a );
 a69453a <=( a69452a  and  a69445a );
 a69457a <=( A298  and  (not A266) );
 a69458a <=( (not A265)  and  a69457a );
 a69461a <=( (not A300)  and  (not A299) );
 a69464a <=( (not A302)  and  (not A301) );
 a69465a <=( a69464a  and  a69461a );
 a69466a <=( a69465a  and  a69458a );
 a69470a <=( A168  and  (not A169) );
 a69471a <=( A170  and  a69470a );
 a69474a <=( A200  and  (not A199) );
 a69477a <=( A203  and  A201 );
 a69478a <=( a69477a  and  a69474a );
 a69479a <=( a69478a  and  a69471a );
 a69483a <=( (not A298)  and  (not A266) );
 a69484a <=( (not A265)  and  a69483a );
 a69487a <=( (not A300)  and  A299 );
 a69490a <=( (not A302)  and  (not A301) );
 a69491a <=( a69490a  and  a69487a );
 a69492a <=( a69491a  and  a69484a );
 a69496a <=( A168  and  (not A169) );
 a69497a <=( A170  and  a69496a );
 a69500a <=( A200  and  (not A199) );
 a69503a <=( (not A202)  and  (not A201) );
 a69504a <=( a69503a  and  a69500a );
 a69505a <=( a69504a  and  a69497a );
 a69509a <=( A268  and  (not A267) );
 a69510a <=( (not A203)  and  a69509a );
 a69513a <=( (not A299)  and  A298 );
 a69516a <=( A301  and  A300 );
 a69517a <=( a69516a  and  a69513a );
 a69518a <=( a69517a  and  a69510a );
 a69522a <=( A168  and  (not A169) );
 a69523a <=( A170  and  a69522a );
 a69526a <=( A200  and  (not A199) );
 a69529a <=( (not A202)  and  (not A201) );
 a69530a <=( a69529a  and  a69526a );
 a69531a <=( a69530a  and  a69523a );
 a69535a <=( A268  and  (not A267) );
 a69536a <=( (not A203)  and  a69535a );
 a69539a <=( (not A299)  and  A298 );
 a69542a <=( A302  and  A300 );
 a69543a <=( a69542a  and  a69539a );
 a69544a <=( a69543a  and  a69536a );
 a69548a <=( A168  and  (not A169) );
 a69549a <=( A170  and  a69548a );
 a69552a <=( A200  and  (not A199) );
 a69555a <=( (not A202)  and  (not A201) );
 a69556a <=( a69555a  and  a69552a );
 a69557a <=( a69556a  and  a69549a );
 a69561a <=( A268  and  (not A267) );
 a69562a <=( (not A203)  and  a69561a );
 a69565a <=( A299  and  (not A298) );
 a69568a <=( A301  and  A300 );
 a69569a <=( a69568a  and  a69565a );
 a69570a <=( a69569a  and  a69562a );
 a69574a <=( A168  and  (not A169) );
 a69575a <=( A170  and  a69574a );
 a69578a <=( A200  and  (not A199) );
 a69581a <=( (not A202)  and  (not A201) );
 a69582a <=( a69581a  and  a69578a );
 a69583a <=( a69582a  and  a69575a );
 a69587a <=( A268  and  (not A267) );
 a69588a <=( (not A203)  and  a69587a );
 a69591a <=( A299  and  (not A298) );
 a69594a <=( A302  and  A300 );
 a69595a <=( a69594a  and  a69591a );
 a69596a <=( a69595a  and  a69588a );
 a69600a <=( A168  and  (not A169) );
 a69601a <=( A170  and  a69600a );
 a69604a <=( A200  and  (not A199) );
 a69607a <=( (not A202)  and  (not A201) );
 a69608a <=( a69607a  and  a69604a );
 a69609a <=( a69608a  and  a69601a );
 a69613a <=( A269  and  (not A267) );
 a69614a <=( (not A203)  and  a69613a );
 a69617a <=( (not A299)  and  A298 );
 a69620a <=( A301  and  A300 );
 a69621a <=( a69620a  and  a69617a );
 a69622a <=( a69621a  and  a69614a );
 a69626a <=( A168  and  (not A169) );
 a69627a <=( A170  and  a69626a );
 a69630a <=( A200  and  (not A199) );
 a69633a <=( (not A202)  and  (not A201) );
 a69634a <=( a69633a  and  a69630a );
 a69635a <=( a69634a  and  a69627a );
 a69639a <=( A269  and  (not A267) );
 a69640a <=( (not A203)  and  a69639a );
 a69643a <=( (not A299)  and  A298 );
 a69646a <=( A302  and  A300 );
 a69647a <=( a69646a  and  a69643a );
 a69648a <=( a69647a  and  a69640a );
 a69652a <=( A168  and  (not A169) );
 a69653a <=( A170  and  a69652a );
 a69656a <=( A200  and  (not A199) );
 a69659a <=( (not A202)  and  (not A201) );
 a69660a <=( a69659a  and  a69656a );
 a69661a <=( a69660a  and  a69653a );
 a69665a <=( A269  and  (not A267) );
 a69666a <=( (not A203)  and  a69665a );
 a69669a <=( A299  and  (not A298) );
 a69672a <=( A301  and  A300 );
 a69673a <=( a69672a  and  a69669a );
 a69674a <=( a69673a  and  a69666a );
 a69678a <=( A168  and  (not A169) );
 a69679a <=( A170  and  a69678a );
 a69682a <=( A200  and  (not A199) );
 a69685a <=( (not A202)  and  (not A201) );
 a69686a <=( a69685a  and  a69682a );
 a69687a <=( a69686a  and  a69679a );
 a69691a <=( A269  and  (not A267) );
 a69692a <=( (not A203)  and  a69691a );
 a69695a <=( A299  and  (not A298) );
 a69698a <=( A302  and  A300 );
 a69699a <=( a69698a  and  a69695a );
 a69700a <=( a69699a  and  a69692a );
 a69704a <=( A168  and  (not A169) );
 a69705a <=( A170  and  a69704a );
 a69708a <=( A200  and  (not A199) );
 a69711a <=( (not A202)  and  (not A201) );
 a69712a <=( a69711a  and  a69708a );
 a69713a <=( a69712a  and  a69705a );
 a69717a <=( A266  and  A265 );
 a69718a <=( (not A203)  and  a69717a );
 a69721a <=( (not A299)  and  A298 );
 a69724a <=( A301  and  A300 );
 a69725a <=( a69724a  and  a69721a );
 a69726a <=( a69725a  and  a69718a );
 a69730a <=( A168  and  (not A169) );
 a69731a <=( A170  and  a69730a );
 a69734a <=( A200  and  (not A199) );
 a69737a <=( (not A202)  and  (not A201) );
 a69738a <=( a69737a  and  a69734a );
 a69739a <=( a69738a  and  a69731a );
 a69743a <=( A266  and  A265 );
 a69744a <=( (not A203)  and  a69743a );
 a69747a <=( (not A299)  and  A298 );
 a69750a <=( A302  and  A300 );
 a69751a <=( a69750a  and  a69747a );
 a69752a <=( a69751a  and  a69744a );
 a69756a <=( A168  and  (not A169) );
 a69757a <=( A170  and  a69756a );
 a69760a <=( A200  and  (not A199) );
 a69763a <=( (not A202)  and  (not A201) );
 a69764a <=( a69763a  and  a69760a );
 a69765a <=( a69764a  and  a69757a );
 a69769a <=( A266  and  A265 );
 a69770a <=( (not A203)  and  a69769a );
 a69773a <=( A299  and  (not A298) );
 a69776a <=( A301  and  A300 );
 a69777a <=( a69776a  and  a69773a );
 a69778a <=( a69777a  and  a69770a );
 a69782a <=( A168  and  (not A169) );
 a69783a <=( A170  and  a69782a );
 a69786a <=( A200  and  (not A199) );
 a69789a <=( (not A202)  and  (not A201) );
 a69790a <=( a69789a  and  a69786a );
 a69791a <=( a69790a  and  a69783a );
 a69795a <=( A266  and  A265 );
 a69796a <=( (not A203)  and  a69795a );
 a69799a <=( A299  and  (not A298) );
 a69802a <=( A302  and  A300 );
 a69803a <=( a69802a  and  a69799a );
 a69804a <=( a69803a  and  a69796a );
 a69808a <=( A168  and  (not A169) );
 a69809a <=( A170  and  a69808a );
 a69812a <=( A200  and  (not A199) );
 a69815a <=( (not A202)  and  (not A201) );
 a69816a <=( a69815a  and  a69812a );
 a69817a <=( a69816a  and  a69809a );
 a69821a <=( (not A266)  and  (not A265) );
 a69822a <=( (not A203)  and  a69821a );
 a69825a <=( (not A299)  and  A298 );
 a69828a <=( A301  and  A300 );
 a69829a <=( a69828a  and  a69825a );
 a69830a <=( a69829a  and  a69822a );
 a69834a <=( A168  and  (not A169) );
 a69835a <=( A170  and  a69834a );
 a69838a <=( A200  and  (not A199) );
 a69841a <=( (not A202)  and  (not A201) );
 a69842a <=( a69841a  and  a69838a );
 a69843a <=( a69842a  and  a69835a );
 a69847a <=( (not A266)  and  (not A265) );
 a69848a <=( (not A203)  and  a69847a );
 a69851a <=( (not A299)  and  A298 );
 a69854a <=( A302  and  A300 );
 a69855a <=( a69854a  and  a69851a );
 a69856a <=( a69855a  and  a69848a );
 a69860a <=( A168  and  (not A169) );
 a69861a <=( A170  and  a69860a );
 a69864a <=( A200  and  (not A199) );
 a69867a <=( (not A202)  and  (not A201) );
 a69868a <=( a69867a  and  a69864a );
 a69869a <=( a69868a  and  a69861a );
 a69873a <=( (not A266)  and  (not A265) );
 a69874a <=( (not A203)  and  a69873a );
 a69877a <=( A299  and  (not A298) );
 a69880a <=( A301  and  A300 );
 a69881a <=( a69880a  and  a69877a );
 a69882a <=( a69881a  and  a69874a );
 a69886a <=( A168  and  (not A169) );
 a69887a <=( A170  and  a69886a );
 a69890a <=( A200  and  (not A199) );
 a69893a <=( (not A202)  and  (not A201) );
 a69894a <=( a69893a  and  a69890a );
 a69895a <=( a69894a  and  a69887a );
 a69899a <=( (not A266)  and  (not A265) );
 a69900a <=( (not A203)  and  a69899a );
 a69903a <=( A299  and  (not A298) );
 a69906a <=( A302  and  A300 );
 a69907a <=( a69906a  and  a69903a );
 a69908a <=( a69907a  and  a69900a );
 a69912a <=( A168  and  (not A169) );
 a69913a <=( A170  and  a69912a );
 a69916a <=( (not A200)  and  A199 );
 a69919a <=( A202  and  A201 );
 a69920a <=( a69919a  and  a69916a );
 a69921a <=( a69920a  and  a69913a );
 a69925a <=( (not A269)  and  (not A268) );
 a69926a <=( A267  and  a69925a );
 a69929a <=( (not A299)  and  A298 );
 a69932a <=( A301  and  A300 );
 a69933a <=( a69932a  and  a69929a );
 a69934a <=( a69933a  and  a69926a );
 a69938a <=( A168  and  (not A169) );
 a69939a <=( A170  and  a69938a );
 a69942a <=( (not A200)  and  A199 );
 a69945a <=( A202  and  A201 );
 a69946a <=( a69945a  and  a69942a );
 a69947a <=( a69946a  and  a69939a );
 a69951a <=( (not A269)  and  (not A268) );
 a69952a <=( A267  and  a69951a );
 a69955a <=( (not A299)  and  A298 );
 a69958a <=( A302  and  A300 );
 a69959a <=( a69958a  and  a69955a );
 a69960a <=( a69959a  and  a69952a );
 a69964a <=( A168  and  (not A169) );
 a69965a <=( A170  and  a69964a );
 a69968a <=( (not A200)  and  A199 );
 a69971a <=( A202  and  A201 );
 a69972a <=( a69971a  and  a69968a );
 a69973a <=( a69972a  and  a69965a );
 a69977a <=( (not A269)  and  (not A268) );
 a69978a <=( A267  and  a69977a );
 a69981a <=( A299  and  (not A298) );
 a69984a <=( A301  and  A300 );
 a69985a <=( a69984a  and  a69981a );
 a69986a <=( a69985a  and  a69978a );
 a69990a <=( A168  and  (not A169) );
 a69991a <=( A170  and  a69990a );
 a69994a <=( (not A200)  and  A199 );
 a69997a <=( A202  and  A201 );
 a69998a <=( a69997a  and  a69994a );
 a69999a <=( a69998a  and  a69991a );
 a70003a <=( (not A269)  and  (not A268) );
 a70004a <=( A267  and  a70003a );
 a70007a <=( A299  and  (not A298) );
 a70010a <=( A302  and  A300 );
 a70011a <=( a70010a  and  a70007a );
 a70012a <=( a70011a  and  a70004a );
 a70016a <=( A168  and  (not A169) );
 a70017a <=( A170  and  a70016a );
 a70020a <=( (not A200)  and  A199 );
 a70023a <=( A202  and  A201 );
 a70024a <=( a70023a  and  a70020a );
 a70025a <=( a70024a  and  a70017a );
 a70029a <=( A298  and  A268 );
 a70030a <=( (not A267)  and  a70029a );
 a70033a <=( (not A300)  and  (not A299) );
 a70036a <=( (not A302)  and  (not A301) );
 a70037a <=( a70036a  and  a70033a );
 a70038a <=( a70037a  and  a70030a );
 a70042a <=( A168  and  (not A169) );
 a70043a <=( A170  and  a70042a );
 a70046a <=( (not A200)  and  A199 );
 a70049a <=( A202  and  A201 );
 a70050a <=( a70049a  and  a70046a );
 a70051a <=( a70050a  and  a70043a );
 a70055a <=( (not A298)  and  A268 );
 a70056a <=( (not A267)  and  a70055a );
 a70059a <=( (not A300)  and  A299 );
 a70062a <=( (not A302)  and  (not A301) );
 a70063a <=( a70062a  and  a70059a );
 a70064a <=( a70063a  and  a70056a );
 a70068a <=( A168  and  (not A169) );
 a70069a <=( A170  and  a70068a );
 a70072a <=( (not A200)  and  A199 );
 a70075a <=( A202  and  A201 );
 a70076a <=( a70075a  and  a70072a );
 a70077a <=( a70076a  and  a70069a );
 a70081a <=( A298  and  A269 );
 a70082a <=( (not A267)  and  a70081a );
 a70085a <=( (not A300)  and  (not A299) );
 a70088a <=( (not A302)  and  (not A301) );
 a70089a <=( a70088a  and  a70085a );
 a70090a <=( a70089a  and  a70082a );
 a70094a <=( A168  and  (not A169) );
 a70095a <=( A170  and  a70094a );
 a70098a <=( (not A200)  and  A199 );
 a70101a <=( A202  and  A201 );
 a70102a <=( a70101a  and  a70098a );
 a70103a <=( a70102a  and  a70095a );
 a70107a <=( (not A298)  and  A269 );
 a70108a <=( (not A267)  and  a70107a );
 a70111a <=( (not A300)  and  A299 );
 a70114a <=( (not A302)  and  (not A301) );
 a70115a <=( a70114a  and  a70111a );
 a70116a <=( a70115a  and  a70108a );
 a70120a <=( A168  and  (not A169) );
 a70121a <=( A170  and  a70120a );
 a70124a <=( (not A200)  and  A199 );
 a70127a <=( A202  and  A201 );
 a70128a <=( a70127a  and  a70124a );
 a70129a <=( a70128a  and  a70121a );
 a70133a <=( A298  and  A266 );
 a70134a <=( A265  and  a70133a );
 a70137a <=( (not A300)  and  (not A299) );
 a70140a <=( (not A302)  and  (not A301) );
 a70141a <=( a70140a  and  a70137a );
 a70142a <=( a70141a  and  a70134a );
 a70146a <=( A168  and  (not A169) );
 a70147a <=( A170  and  a70146a );
 a70150a <=( (not A200)  and  A199 );
 a70153a <=( A202  and  A201 );
 a70154a <=( a70153a  and  a70150a );
 a70155a <=( a70154a  and  a70147a );
 a70159a <=( (not A298)  and  A266 );
 a70160a <=( A265  and  a70159a );
 a70163a <=( (not A300)  and  A299 );
 a70166a <=( (not A302)  and  (not A301) );
 a70167a <=( a70166a  and  a70163a );
 a70168a <=( a70167a  and  a70160a );
 a70172a <=( A168  and  (not A169) );
 a70173a <=( A170  and  a70172a );
 a70176a <=( (not A200)  and  A199 );
 a70179a <=( A202  and  A201 );
 a70180a <=( a70179a  and  a70176a );
 a70181a <=( a70180a  and  a70173a );
 a70185a <=( A298  and  (not A266) );
 a70186a <=( (not A265)  and  a70185a );
 a70189a <=( (not A300)  and  (not A299) );
 a70192a <=( (not A302)  and  (not A301) );
 a70193a <=( a70192a  and  a70189a );
 a70194a <=( a70193a  and  a70186a );
 a70198a <=( A168  and  (not A169) );
 a70199a <=( A170  and  a70198a );
 a70202a <=( (not A200)  and  A199 );
 a70205a <=( A202  and  A201 );
 a70206a <=( a70205a  and  a70202a );
 a70207a <=( a70206a  and  a70199a );
 a70211a <=( (not A298)  and  (not A266) );
 a70212a <=( (not A265)  and  a70211a );
 a70215a <=( (not A300)  and  A299 );
 a70218a <=( (not A302)  and  (not A301) );
 a70219a <=( a70218a  and  a70215a );
 a70220a <=( a70219a  and  a70212a );
 a70224a <=( A168  and  (not A169) );
 a70225a <=( A170  and  a70224a );
 a70228a <=( (not A200)  and  A199 );
 a70231a <=( A203  and  A201 );
 a70232a <=( a70231a  and  a70228a );
 a70233a <=( a70232a  and  a70225a );
 a70237a <=( (not A269)  and  (not A268) );
 a70238a <=( A267  and  a70237a );
 a70241a <=( (not A299)  and  A298 );
 a70244a <=( A301  and  A300 );
 a70245a <=( a70244a  and  a70241a );
 a70246a <=( a70245a  and  a70238a );
 a70250a <=( A168  and  (not A169) );
 a70251a <=( A170  and  a70250a );
 a70254a <=( (not A200)  and  A199 );
 a70257a <=( A203  and  A201 );
 a70258a <=( a70257a  and  a70254a );
 a70259a <=( a70258a  and  a70251a );
 a70263a <=( (not A269)  and  (not A268) );
 a70264a <=( A267  and  a70263a );
 a70267a <=( (not A299)  and  A298 );
 a70270a <=( A302  and  A300 );
 a70271a <=( a70270a  and  a70267a );
 a70272a <=( a70271a  and  a70264a );
 a70276a <=( A168  and  (not A169) );
 a70277a <=( A170  and  a70276a );
 a70280a <=( (not A200)  and  A199 );
 a70283a <=( A203  and  A201 );
 a70284a <=( a70283a  and  a70280a );
 a70285a <=( a70284a  and  a70277a );
 a70289a <=( (not A269)  and  (not A268) );
 a70290a <=( A267  and  a70289a );
 a70293a <=( A299  and  (not A298) );
 a70296a <=( A301  and  A300 );
 a70297a <=( a70296a  and  a70293a );
 a70298a <=( a70297a  and  a70290a );
 a70302a <=( A168  and  (not A169) );
 a70303a <=( A170  and  a70302a );
 a70306a <=( (not A200)  and  A199 );
 a70309a <=( A203  and  A201 );
 a70310a <=( a70309a  and  a70306a );
 a70311a <=( a70310a  and  a70303a );
 a70315a <=( (not A269)  and  (not A268) );
 a70316a <=( A267  and  a70315a );
 a70319a <=( A299  and  (not A298) );
 a70322a <=( A302  and  A300 );
 a70323a <=( a70322a  and  a70319a );
 a70324a <=( a70323a  and  a70316a );
 a70328a <=( A168  and  (not A169) );
 a70329a <=( A170  and  a70328a );
 a70332a <=( (not A200)  and  A199 );
 a70335a <=( A203  and  A201 );
 a70336a <=( a70335a  and  a70332a );
 a70337a <=( a70336a  and  a70329a );
 a70341a <=( A298  and  A268 );
 a70342a <=( (not A267)  and  a70341a );
 a70345a <=( (not A300)  and  (not A299) );
 a70348a <=( (not A302)  and  (not A301) );
 a70349a <=( a70348a  and  a70345a );
 a70350a <=( a70349a  and  a70342a );
 a70354a <=( A168  and  (not A169) );
 a70355a <=( A170  and  a70354a );
 a70358a <=( (not A200)  and  A199 );
 a70361a <=( A203  and  A201 );
 a70362a <=( a70361a  and  a70358a );
 a70363a <=( a70362a  and  a70355a );
 a70367a <=( (not A298)  and  A268 );
 a70368a <=( (not A267)  and  a70367a );
 a70371a <=( (not A300)  and  A299 );
 a70374a <=( (not A302)  and  (not A301) );
 a70375a <=( a70374a  and  a70371a );
 a70376a <=( a70375a  and  a70368a );
 a70380a <=( A168  and  (not A169) );
 a70381a <=( A170  and  a70380a );
 a70384a <=( (not A200)  and  A199 );
 a70387a <=( A203  and  A201 );
 a70388a <=( a70387a  and  a70384a );
 a70389a <=( a70388a  and  a70381a );
 a70393a <=( A298  and  A269 );
 a70394a <=( (not A267)  and  a70393a );
 a70397a <=( (not A300)  and  (not A299) );
 a70400a <=( (not A302)  and  (not A301) );
 a70401a <=( a70400a  and  a70397a );
 a70402a <=( a70401a  and  a70394a );
 a70406a <=( A168  and  (not A169) );
 a70407a <=( A170  and  a70406a );
 a70410a <=( (not A200)  and  A199 );
 a70413a <=( A203  and  A201 );
 a70414a <=( a70413a  and  a70410a );
 a70415a <=( a70414a  and  a70407a );
 a70419a <=( (not A298)  and  A269 );
 a70420a <=( (not A267)  and  a70419a );
 a70423a <=( (not A300)  and  A299 );
 a70426a <=( (not A302)  and  (not A301) );
 a70427a <=( a70426a  and  a70423a );
 a70428a <=( a70427a  and  a70420a );
 a70432a <=( A168  and  (not A169) );
 a70433a <=( A170  and  a70432a );
 a70436a <=( (not A200)  and  A199 );
 a70439a <=( A203  and  A201 );
 a70440a <=( a70439a  and  a70436a );
 a70441a <=( a70440a  and  a70433a );
 a70445a <=( A298  and  A266 );
 a70446a <=( A265  and  a70445a );
 a70449a <=( (not A300)  and  (not A299) );
 a70452a <=( (not A302)  and  (not A301) );
 a70453a <=( a70452a  and  a70449a );
 a70454a <=( a70453a  and  a70446a );
 a70458a <=( A168  and  (not A169) );
 a70459a <=( A170  and  a70458a );
 a70462a <=( (not A200)  and  A199 );
 a70465a <=( A203  and  A201 );
 a70466a <=( a70465a  and  a70462a );
 a70467a <=( a70466a  and  a70459a );
 a70471a <=( (not A298)  and  A266 );
 a70472a <=( A265  and  a70471a );
 a70475a <=( (not A300)  and  A299 );
 a70478a <=( (not A302)  and  (not A301) );
 a70479a <=( a70478a  and  a70475a );
 a70480a <=( a70479a  and  a70472a );
 a70484a <=( A168  and  (not A169) );
 a70485a <=( A170  and  a70484a );
 a70488a <=( (not A200)  and  A199 );
 a70491a <=( A203  and  A201 );
 a70492a <=( a70491a  and  a70488a );
 a70493a <=( a70492a  and  a70485a );
 a70497a <=( A298  and  (not A266) );
 a70498a <=( (not A265)  and  a70497a );
 a70501a <=( (not A300)  and  (not A299) );
 a70504a <=( (not A302)  and  (not A301) );
 a70505a <=( a70504a  and  a70501a );
 a70506a <=( a70505a  and  a70498a );
 a70510a <=( A168  and  (not A169) );
 a70511a <=( A170  and  a70510a );
 a70514a <=( (not A200)  and  A199 );
 a70517a <=( A203  and  A201 );
 a70518a <=( a70517a  and  a70514a );
 a70519a <=( a70518a  and  a70511a );
 a70523a <=( (not A298)  and  (not A266) );
 a70524a <=( (not A265)  and  a70523a );
 a70527a <=( (not A300)  and  A299 );
 a70530a <=( (not A302)  and  (not A301) );
 a70531a <=( a70530a  and  a70527a );
 a70532a <=( a70531a  and  a70524a );
 a70536a <=( A168  and  (not A169) );
 a70537a <=( A170  and  a70536a );
 a70540a <=( (not A200)  and  A199 );
 a70543a <=( (not A202)  and  (not A201) );
 a70544a <=( a70543a  and  a70540a );
 a70545a <=( a70544a  and  a70537a );
 a70549a <=( A268  and  (not A267) );
 a70550a <=( (not A203)  and  a70549a );
 a70553a <=( (not A299)  and  A298 );
 a70556a <=( A301  and  A300 );
 a70557a <=( a70556a  and  a70553a );
 a70558a <=( a70557a  and  a70550a );
 a70562a <=( A168  and  (not A169) );
 a70563a <=( A170  and  a70562a );
 a70566a <=( (not A200)  and  A199 );
 a70569a <=( (not A202)  and  (not A201) );
 a70570a <=( a70569a  and  a70566a );
 a70571a <=( a70570a  and  a70563a );
 a70575a <=( A268  and  (not A267) );
 a70576a <=( (not A203)  and  a70575a );
 a70579a <=( (not A299)  and  A298 );
 a70582a <=( A302  and  A300 );
 a70583a <=( a70582a  and  a70579a );
 a70584a <=( a70583a  and  a70576a );
 a70588a <=( A168  and  (not A169) );
 a70589a <=( A170  and  a70588a );
 a70592a <=( (not A200)  and  A199 );
 a70595a <=( (not A202)  and  (not A201) );
 a70596a <=( a70595a  and  a70592a );
 a70597a <=( a70596a  and  a70589a );
 a70601a <=( A268  and  (not A267) );
 a70602a <=( (not A203)  and  a70601a );
 a70605a <=( A299  and  (not A298) );
 a70608a <=( A301  and  A300 );
 a70609a <=( a70608a  and  a70605a );
 a70610a <=( a70609a  and  a70602a );
 a70614a <=( A168  and  (not A169) );
 a70615a <=( A170  and  a70614a );
 a70618a <=( (not A200)  and  A199 );
 a70621a <=( (not A202)  and  (not A201) );
 a70622a <=( a70621a  and  a70618a );
 a70623a <=( a70622a  and  a70615a );
 a70627a <=( A268  and  (not A267) );
 a70628a <=( (not A203)  and  a70627a );
 a70631a <=( A299  and  (not A298) );
 a70634a <=( A302  and  A300 );
 a70635a <=( a70634a  and  a70631a );
 a70636a <=( a70635a  and  a70628a );
 a70640a <=( A168  and  (not A169) );
 a70641a <=( A170  and  a70640a );
 a70644a <=( (not A200)  and  A199 );
 a70647a <=( (not A202)  and  (not A201) );
 a70648a <=( a70647a  and  a70644a );
 a70649a <=( a70648a  and  a70641a );
 a70653a <=( A269  and  (not A267) );
 a70654a <=( (not A203)  and  a70653a );
 a70657a <=( (not A299)  and  A298 );
 a70660a <=( A301  and  A300 );
 a70661a <=( a70660a  and  a70657a );
 a70662a <=( a70661a  and  a70654a );
 a70666a <=( A168  and  (not A169) );
 a70667a <=( A170  and  a70666a );
 a70670a <=( (not A200)  and  A199 );
 a70673a <=( (not A202)  and  (not A201) );
 a70674a <=( a70673a  and  a70670a );
 a70675a <=( a70674a  and  a70667a );
 a70679a <=( A269  and  (not A267) );
 a70680a <=( (not A203)  and  a70679a );
 a70683a <=( (not A299)  and  A298 );
 a70686a <=( A302  and  A300 );
 a70687a <=( a70686a  and  a70683a );
 a70688a <=( a70687a  and  a70680a );
 a70692a <=( A168  and  (not A169) );
 a70693a <=( A170  and  a70692a );
 a70696a <=( (not A200)  and  A199 );
 a70699a <=( (not A202)  and  (not A201) );
 a70700a <=( a70699a  and  a70696a );
 a70701a <=( a70700a  and  a70693a );
 a70705a <=( A269  and  (not A267) );
 a70706a <=( (not A203)  and  a70705a );
 a70709a <=( A299  and  (not A298) );
 a70712a <=( A301  and  A300 );
 a70713a <=( a70712a  and  a70709a );
 a70714a <=( a70713a  and  a70706a );
 a70718a <=( A168  and  (not A169) );
 a70719a <=( A170  and  a70718a );
 a70722a <=( (not A200)  and  A199 );
 a70725a <=( (not A202)  and  (not A201) );
 a70726a <=( a70725a  and  a70722a );
 a70727a <=( a70726a  and  a70719a );
 a70731a <=( A269  and  (not A267) );
 a70732a <=( (not A203)  and  a70731a );
 a70735a <=( A299  and  (not A298) );
 a70738a <=( A302  and  A300 );
 a70739a <=( a70738a  and  a70735a );
 a70740a <=( a70739a  and  a70732a );
 a70744a <=( A168  and  (not A169) );
 a70745a <=( A170  and  a70744a );
 a70748a <=( (not A200)  and  A199 );
 a70751a <=( (not A202)  and  (not A201) );
 a70752a <=( a70751a  and  a70748a );
 a70753a <=( a70752a  and  a70745a );
 a70757a <=( A266  and  A265 );
 a70758a <=( (not A203)  and  a70757a );
 a70761a <=( (not A299)  and  A298 );
 a70764a <=( A301  and  A300 );
 a70765a <=( a70764a  and  a70761a );
 a70766a <=( a70765a  and  a70758a );
 a70770a <=( A168  and  (not A169) );
 a70771a <=( A170  and  a70770a );
 a70774a <=( (not A200)  and  A199 );
 a70777a <=( (not A202)  and  (not A201) );
 a70778a <=( a70777a  and  a70774a );
 a70779a <=( a70778a  and  a70771a );
 a70783a <=( A266  and  A265 );
 a70784a <=( (not A203)  and  a70783a );
 a70787a <=( (not A299)  and  A298 );
 a70790a <=( A302  and  A300 );
 a70791a <=( a70790a  and  a70787a );
 a70792a <=( a70791a  and  a70784a );
 a70796a <=( A168  and  (not A169) );
 a70797a <=( A170  and  a70796a );
 a70800a <=( (not A200)  and  A199 );
 a70803a <=( (not A202)  and  (not A201) );
 a70804a <=( a70803a  and  a70800a );
 a70805a <=( a70804a  and  a70797a );
 a70809a <=( A266  and  A265 );
 a70810a <=( (not A203)  and  a70809a );
 a70813a <=( A299  and  (not A298) );
 a70816a <=( A301  and  A300 );
 a70817a <=( a70816a  and  a70813a );
 a70818a <=( a70817a  and  a70810a );
 a70822a <=( A168  and  (not A169) );
 a70823a <=( A170  and  a70822a );
 a70826a <=( (not A200)  and  A199 );
 a70829a <=( (not A202)  and  (not A201) );
 a70830a <=( a70829a  and  a70826a );
 a70831a <=( a70830a  and  a70823a );
 a70835a <=( A266  and  A265 );
 a70836a <=( (not A203)  and  a70835a );
 a70839a <=( A299  and  (not A298) );
 a70842a <=( A302  and  A300 );
 a70843a <=( a70842a  and  a70839a );
 a70844a <=( a70843a  and  a70836a );
 a70848a <=( A168  and  (not A169) );
 a70849a <=( A170  and  a70848a );
 a70852a <=( (not A200)  and  A199 );
 a70855a <=( (not A202)  and  (not A201) );
 a70856a <=( a70855a  and  a70852a );
 a70857a <=( a70856a  and  a70849a );
 a70861a <=( (not A266)  and  (not A265) );
 a70862a <=( (not A203)  and  a70861a );
 a70865a <=( (not A299)  and  A298 );
 a70868a <=( A301  and  A300 );
 a70869a <=( a70868a  and  a70865a );
 a70870a <=( a70869a  and  a70862a );
 a70874a <=( A168  and  (not A169) );
 a70875a <=( A170  and  a70874a );
 a70878a <=( (not A200)  and  A199 );
 a70881a <=( (not A202)  and  (not A201) );
 a70882a <=( a70881a  and  a70878a );
 a70883a <=( a70882a  and  a70875a );
 a70887a <=( (not A266)  and  (not A265) );
 a70888a <=( (not A203)  and  a70887a );
 a70891a <=( (not A299)  and  A298 );
 a70894a <=( A302  and  A300 );
 a70895a <=( a70894a  and  a70891a );
 a70896a <=( a70895a  and  a70888a );
 a70900a <=( A168  and  (not A169) );
 a70901a <=( A170  and  a70900a );
 a70904a <=( (not A200)  and  A199 );
 a70907a <=( (not A202)  and  (not A201) );
 a70908a <=( a70907a  and  a70904a );
 a70909a <=( a70908a  and  a70901a );
 a70913a <=( (not A266)  and  (not A265) );
 a70914a <=( (not A203)  and  a70913a );
 a70917a <=( A299  and  (not A298) );
 a70920a <=( A301  and  A300 );
 a70921a <=( a70920a  and  a70917a );
 a70922a <=( a70921a  and  a70914a );
 a70926a <=( A168  and  (not A169) );
 a70927a <=( A170  and  a70926a );
 a70930a <=( (not A200)  and  A199 );
 a70933a <=( (not A202)  and  (not A201) );
 a70934a <=( a70933a  and  a70930a );
 a70935a <=( a70934a  and  a70927a );
 a70939a <=( (not A266)  and  (not A265) );
 a70940a <=( (not A203)  and  a70939a );
 a70943a <=( A299  and  (not A298) );
 a70946a <=( A302  and  A300 );
 a70947a <=( a70946a  and  a70943a );
 a70948a <=( a70947a  and  a70940a );
 a70952a <=( (not A168)  and  (not A169) );
 a70953a <=( A170  and  a70952a );
 a70956a <=( (not A166)  and  A167 );
 a70959a <=( (not A202)  and  A201 );
 a70960a <=( a70959a  and  a70956a );
 a70961a <=( a70960a  and  a70953a );
 a70965a <=( A268  and  (not A267) );
 a70966a <=( (not A203)  and  a70965a );
 a70969a <=( (not A299)  and  A298 );
 a70972a <=( A301  and  A300 );
 a70973a <=( a70972a  and  a70969a );
 a70974a <=( a70973a  and  a70966a );
 a70978a <=( (not A168)  and  (not A169) );
 a70979a <=( A170  and  a70978a );
 a70982a <=( (not A166)  and  A167 );
 a70985a <=( (not A202)  and  A201 );
 a70986a <=( a70985a  and  a70982a );
 a70987a <=( a70986a  and  a70979a );
 a70991a <=( A268  and  (not A267) );
 a70992a <=( (not A203)  and  a70991a );
 a70995a <=( (not A299)  and  A298 );
 a70998a <=( A302  and  A300 );
 a70999a <=( a70998a  and  a70995a );
 a71000a <=( a70999a  and  a70992a );
 a71004a <=( (not A168)  and  (not A169) );
 a71005a <=( A170  and  a71004a );
 a71008a <=( (not A166)  and  A167 );
 a71011a <=( (not A202)  and  A201 );
 a71012a <=( a71011a  and  a71008a );
 a71013a <=( a71012a  and  a71005a );
 a71017a <=( A268  and  (not A267) );
 a71018a <=( (not A203)  and  a71017a );
 a71021a <=( A299  and  (not A298) );
 a71024a <=( A301  and  A300 );
 a71025a <=( a71024a  and  a71021a );
 a71026a <=( a71025a  and  a71018a );
 a71030a <=( (not A168)  and  (not A169) );
 a71031a <=( A170  and  a71030a );
 a71034a <=( (not A166)  and  A167 );
 a71037a <=( (not A202)  and  A201 );
 a71038a <=( a71037a  and  a71034a );
 a71039a <=( a71038a  and  a71031a );
 a71043a <=( A268  and  (not A267) );
 a71044a <=( (not A203)  and  a71043a );
 a71047a <=( A299  and  (not A298) );
 a71050a <=( A302  and  A300 );
 a71051a <=( a71050a  and  a71047a );
 a71052a <=( a71051a  and  a71044a );
 a71056a <=( (not A168)  and  (not A169) );
 a71057a <=( A170  and  a71056a );
 a71060a <=( (not A166)  and  A167 );
 a71063a <=( (not A202)  and  A201 );
 a71064a <=( a71063a  and  a71060a );
 a71065a <=( a71064a  and  a71057a );
 a71069a <=( A269  and  (not A267) );
 a71070a <=( (not A203)  and  a71069a );
 a71073a <=( (not A299)  and  A298 );
 a71076a <=( A301  and  A300 );
 a71077a <=( a71076a  and  a71073a );
 a71078a <=( a71077a  and  a71070a );
 a71082a <=( (not A168)  and  (not A169) );
 a71083a <=( A170  and  a71082a );
 a71086a <=( (not A166)  and  A167 );
 a71089a <=( (not A202)  and  A201 );
 a71090a <=( a71089a  and  a71086a );
 a71091a <=( a71090a  and  a71083a );
 a71095a <=( A269  and  (not A267) );
 a71096a <=( (not A203)  and  a71095a );
 a71099a <=( (not A299)  and  A298 );
 a71102a <=( A302  and  A300 );
 a71103a <=( a71102a  and  a71099a );
 a71104a <=( a71103a  and  a71096a );
 a71108a <=( (not A168)  and  (not A169) );
 a71109a <=( A170  and  a71108a );
 a71112a <=( (not A166)  and  A167 );
 a71115a <=( (not A202)  and  A201 );
 a71116a <=( a71115a  and  a71112a );
 a71117a <=( a71116a  and  a71109a );
 a71121a <=( A269  and  (not A267) );
 a71122a <=( (not A203)  and  a71121a );
 a71125a <=( A299  and  (not A298) );
 a71128a <=( A301  and  A300 );
 a71129a <=( a71128a  and  a71125a );
 a71130a <=( a71129a  and  a71122a );
 a71134a <=( (not A168)  and  (not A169) );
 a71135a <=( A170  and  a71134a );
 a71138a <=( (not A166)  and  A167 );
 a71141a <=( (not A202)  and  A201 );
 a71142a <=( a71141a  and  a71138a );
 a71143a <=( a71142a  and  a71135a );
 a71147a <=( A269  and  (not A267) );
 a71148a <=( (not A203)  and  a71147a );
 a71151a <=( A299  and  (not A298) );
 a71154a <=( A302  and  A300 );
 a71155a <=( a71154a  and  a71151a );
 a71156a <=( a71155a  and  a71148a );
 a71160a <=( (not A168)  and  (not A169) );
 a71161a <=( A170  and  a71160a );
 a71164a <=( (not A166)  and  A167 );
 a71167a <=( (not A202)  and  A201 );
 a71168a <=( a71167a  and  a71164a );
 a71169a <=( a71168a  and  a71161a );
 a71173a <=( A266  and  A265 );
 a71174a <=( (not A203)  and  a71173a );
 a71177a <=( (not A299)  and  A298 );
 a71180a <=( A301  and  A300 );
 a71181a <=( a71180a  and  a71177a );
 a71182a <=( a71181a  and  a71174a );
 a71186a <=( (not A168)  and  (not A169) );
 a71187a <=( A170  and  a71186a );
 a71190a <=( (not A166)  and  A167 );
 a71193a <=( (not A202)  and  A201 );
 a71194a <=( a71193a  and  a71190a );
 a71195a <=( a71194a  and  a71187a );
 a71199a <=( A266  and  A265 );
 a71200a <=( (not A203)  and  a71199a );
 a71203a <=( (not A299)  and  A298 );
 a71206a <=( A302  and  A300 );
 a71207a <=( a71206a  and  a71203a );
 a71208a <=( a71207a  and  a71200a );
 a71212a <=( (not A168)  and  (not A169) );
 a71213a <=( A170  and  a71212a );
 a71216a <=( (not A166)  and  A167 );
 a71219a <=( (not A202)  and  A201 );
 a71220a <=( a71219a  and  a71216a );
 a71221a <=( a71220a  and  a71213a );
 a71225a <=( A266  and  A265 );
 a71226a <=( (not A203)  and  a71225a );
 a71229a <=( A299  and  (not A298) );
 a71232a <=( A301  and  A300 );
 a71233a <=( a71232a  and  a71229a );
 a71234a <=( a71233a  and  a71226a );
 a71238a <=( (not A168)  and  (not A169) );
 a71239a <=( A170  and  a71238a );
 a71242a <=( (not A166)  and  A167 );
 a71245a <=( (not A202)  and  A201 );
 a71246a <=( a71245a  and  a71242a );
 a71247a <=( a71246a  and  a71239a );
 a71251a <=( A266  and  A265 );
 a71252a <=( (not A203)  and  a71251a );
 a71255a <=( A299  and  (not A298) );
 a71258a <=( A302  and  A300 );
 a71259a <=( a71258a  and  a71255a );
 a71260a <=( a71259a  and  a71252a );
 a71264a <=( (not A168)  and  (not A169) );
 a71265a <=( A170  and  a71264a );
 a71268a <=( (not A166)  and  A167 );
 a71271a <=( (not A202)  and  A201 );
 a71272a <=( a71271a  and  a71268a );
 a71273a <=( a71272a  and  a71265a );
 a71277a <=( (not A266)  and  (not A265) );
 a71278a <=( (not A203)  and  a71277a );
 a71281a <=( (not A299)  and  A298 );
 a71284a <=( A301  and  A300 );
 a71285a <=( a71284a  and  a71281a );
 a71286a <=( a71285a  and  a71278a );
 a71290a <=( (not A168)  and  (not A169) );
 a71291a <=( A170  and  a71290a );
 a71294a <=( (not A166)  and  A167 );
 a71297a <=( (not A202)  and  A201 );
 a71298a <=( a71297a  and  a71294a );
 a71299a <=( a71298a  and  a71291a );
 a71303a <=( (not A266)  and  (not A265) );
 a71304a <=( (not A203)  and  a71303a );
 a71307a <=( (not A299)  and  A298 );
 a71310a <=( A302  and  A300 );
 a71311a <=( a71310a  and  a71307a );
 a71312a <=( a71311a  and  a71304a );
 a71316a <=( (not A168)  and  (not A169) );
 a71317a <=( A170  and  a71316a );
 a71320a <=( (not A166)  and  A167 );
 a71323a <=( (not A202)  and  A201 );
 a71324a <=( a71323a  and  a71320a );
 a71325a <=( a71324a  and  a71317a );
 a71329a <=( (not A266)  and  (not A265) );
 a71330a <=( (not A203)  and  a71329a );
 a71333a <=( A299  and  (not A298) );
 a71336a <=( A301  and  A300 );
 a71337a <=( a71336a  and  a71333a );
 a71338a <=( a71337a  and  a71330a );
 a71342a <=( (not A168)  and  (not A169) );
 a71343a <=( A170  and  a71342a );
 a71346a <=( (not A166)  and  A167 );
 a71349a <=( (not A202)  and  A201 );
 a71350a <=( a71349a  and  a71346a );
 a71351a <=( a71350a  and  a71343a );
 a71355a <=( (not A266)  and  (not A265) );
 a71356a <=( (not A203)  and  a71355a );
 a71359a <=( A299  and  (not A298) );
 a71362a <=( A302  and  A300 );
 a71363a <=( a71362a  and  a71359a );
 a71364a <=( a71363a  and  a71356a );
 a71368a <=( (not A168)  and  (not A169) );
 a71369a <=( A170  and  a71368a );
 a71372a <=( (not A166)  and  A167 );
 a71375a <=( A202  and  (not A201) );
 a71376a <=( a71375a  and  a71372a );
 a71377a <=( a71376a  and  a71369a );
 a71381a <=( (not A269)  and  (not A268) );
 a71382a <=( A267  and  a71381a );
 a71385a <=( (not A299)  and  A298 );
 a71388a <=( A301  and  A300 );
 a71389a <=( a71388a  and  a71385a );
 a71390a <=( a71389a  and  a71382a );
 a71394a <=( (not A168)  and  (not A169) );
 a71395a <=( A170  and  a71394a );
 a71398a <=( (not A166)  and  A167 );
 a71401a <=( A202  and  (not A201) );
 a71402a <=( a71401a  and  a71398a );
 a71403a <=( a71402a  and  a71395a );
 a71407a <=( (not A269)  and  (not A268) );
 a71408a <=( A267  and  a71407a );
 a71411a <=( (not A299)  and  A298 );
 a71414a <=( A302  and  A300 );
 a71415a <=( a71414a  and  a71411a );
 a71416a <=( a71415a  and  a71408a );
 a71420a <=( (not A168)  and  (not A169) );
 a71421a <=( A170  and  a71420a );
 a71424a <=( (not A166)  and  A167 );
 a71427a <=( A202  and  (not A201) );
 a71428a <=( a71427a  and  a71424a );
 a71429a <=( a71428a  and  a71421a );
 a71433a <=( (not A269)  and  (not A268) );
 a71434a <=( A267  and  a71433a );
 a71437a <=( A299  and  (not A298) );
 a71440a <=( A301  and  A300 );
 a71441a <=( a71440a  and  a71437a );
 a71442a <=( a71441a  and  a71434a );
 a71446a <=( (not A168)  and  (not A169) );
 a71447a <=( A170  and  a71446a );
 a71450a <=( (not A166)  and  A167 );
 a71453a <=( A202  and  (not A201) );
 a71454a <=( a71453a  and  a71450a );
 a71455a <=( a71454a  and  a71447a );
 a71459a <=( (not A269)  and  (not A268) );
 a71460a <=( A267  and  a71459a );
 a71463a <=( A299  and  (not A298) );
 a71466a <=( A302  and  A300 );
 a71467a <=( a71466a  and  a71463a );
 a71468a <=( a71467a  and  a71460a );
 a71472a <=( (not A168)  and  (not A169) );
 a71473a <=( A170  and  a71472a );
 a71476a <=( (not A166)  and  A167 );
 a71479a <=( A202  and  (not A201) );
 a71480a <=( a71479a  and  a71476a );
 a71481a <=( a71480a  and  a71473a );
 a71485a <=( A298  and  A268 );
 a71486a <=( (not A267)  and  a71485a );
 a71489a <=( (not A300)  and  (not A299) );
 a71492a <=( (not A302)  and  (not A301) );
 a71493a <=( a71492a  and  a71489a );
 a71494a <=( a71493a  and  a71486a );
 a71498a <=( (not A168)  and  (not A169) );
 a71499a <=( A170  and  a71498a );
 a71502a <=( (not A166)  and  A167 );
 a71505a <=( A202  and  (not A201) );
 a71506a <=( a71505a  and  a71502a );
 a71507a <=( a71506a  and  a71499a );
 a71511a <=( (not A298)  and  A268 );
 a71512a <=( (not A267)  and  a71511a );
 a71515a <=( (not A300)  and  A299 );
 a71518a <=( (not A302)  and  (not A301) );
 a71519a <=( a71518a  and  a71515a );
 a71520a <=( a71519a  and  a71512a );
 a71524a <=( (not A168)  and  (not A169) );
 a71525a <=( A170  and  a71524a );
 a71528a <=( (not A166)  and  A167 );
 a71531a <=( A202  and  (not A201) );
 a71532a <=( a71531a  and  a71528a );
 a71533a <=( a71532a  and  a71525a );
 a71537a <=( A298  and  A269 );
 a71538a <=( (not A267)  and  a71537a );
 a71541a <=( (not A300)  and  (not A299) );
 a71544a <=( (not A302)  and  (not A301) );
 a71545a <=( a71544a  and  a71541a );
 a71546a <=( a71545a  and  a71538a );
 a71550a <=( (not A168)  and  (not A169) );
 a71551a <=( A170  and  a71550a );
 a71554a <=( (not A166)  and  A167 );
 a71557a <=( A202  and  (not A201) );
 a71558a <=( a71557a  and  a71554a );
 a71559a <=( a71558a  and  a71551a );
 a71563a <=( (not A298)  and  A269 );
 a71564a <=( (not A267)  and  a71563a );
 a71567a <=( (not A300)  and  A299 );
 a71570a <=( (not A302)  and  (not A301) );
 a71571a <=( a71570a  and  a71567a );
 a71572a <=( a71571a  and  a71564a );
 a71576a <=( (not A168)  and  (not A169) );
 a71577a <=( A170  and  a71576a );
 a71580a <=( (not A166)  and  A167 );
 a71583a <=( A202  and  (not A201) );
 a71584a <=( a71583a  and  a71580a );
 a71585a <=( a71584a  and  a71577a );
 a71589a <=( A298  and  A266 );
 a71590a <=( A265  and  a71589a );
 a71593a <=( (not A300)  and  (not A299) );
 a71596a <=( (not A302)  and  (not A301) );
 a71597a <=( a71596a  and  a71593a );
 a71598a <=( a71597a  and  a71590a );
 a71602a <=( (not A168)  and  (not A169) );
 a71603a <=( A170  and  a71602a );
 a71606a <=( (not A166)  and  A167 );
 a71609a <=( A202  and  (not A201) );
 a71610a <=( a71609a  and  a71606a );
 a71611a <=( a71610a  and  a71603a );
 a71615a <=( (not A298)  and  A266 );
 a71616a <=( A265  and  a71615a );
 a71619a <=( (not A300)  and  A299 );
 a71622a <=( (not A302)  and  (not A301) );
 a71623a <=( a71622a  and  a71619a );
 a71624a <=( a71623a  and  a71616a );
 a71628a <=( (not A168)  and  (not A169) );
 a71629a <=( A170  and  a71628a );
 a71632a <=( (not A166)  and  A167 );
 a71635a <=( A202  and  (not A201) );
 a71636a <=( a71635a  and  a71632a );
 a71637a <=( a71636a  and  a71629a );
 a71641a <=( A298  and  (not A266) );
 a71642a <=( (not A265)  and  a71641a );
 a71645a <=( (not A300)  and  (not A299) );
 a71648a <=( (not A302)  and  (not A301) );
 a71649a <=( a71648a  and  a71645a );
 a71650a <=( a71649a  and  a71642a );
 a71654a <=( (not A168)  and  (not A169) );
 a71655a <=( A170  and  a71654a );
 a71658a <=( (not A166)  and  A167 );
 a71661a <=( A202  and  (not A201) );
 a71662a <=( a71661a  and  a71658a );
 a71663a <=( a71662a  and  a71655a );
 a71667a <=( (not A298)  and  (not A266) );
 a71668a <=( (not A265)  and  a71667a );
 a71671a <=( (not A300)  and  A299 );
 a71674a <=( (not A302)  and  (not A301) );
 a71675a <=( a71674a  and  a71671a );
 a71676a <=( a71675a  and  a71668a );
 a71680a <=( (not A168)  and  (not A169) );
 a71681a <=( A170  and  a71680a );
 a71684a <=( (not A166)  and  A167 );
 a71687a <=( A203  and  (not A201) );
 a71688a <=( a71687a  and  a71684a );
 a71689a <=( a71688a  and  a71681a );
 a71693a <=( (not A269)  and  (not A268) );
 a71694a <=( A267  and  a71693a );
 a71697a <=( (not A299)  and  A298 );
 a71700a <=( A301  and  A300 );
 a71701a <=( a71700a  and  a71697a );
 a71702a <=( a71701a  and  a71694a );
 a71706a <=( (not A168)  and  (not A169) );
 a71707a <=( A170  and  a71706a );
 a71710a <=( (not A166)  and  A167 );
 a71713a <=( A203  and  (not A201) );
 a71714a <=( a71713a  and  a71710a );
 a71715a <=( a71714a  and  a71707a );
 a71719a <=( (not A269)  and  (not A268) );
 a71720a <=( A267  and  a71719a );
 a71723a <=( (not A299)  and  A298 );
 a71726a <=( A302  and  A300 );
 a71727a <=( a71726a  and  a71723a );
 a71728a <=( a71727a  and  a71720a );
 a71732a <=( (not A168)  and  (not A169) );
 a71733a <=( A170  and  a71732a );
 a71736a <=( (not A166)  and  A167 );
 a71739a <=( A203  and  (not A201) );
 a71740a <=( a71739a  and  a71736a );
 a71741a <=( a71740a  and  a71733a );
 a71745a <=( (not A269)  and  (not A268) );
 a71746a <=( A267  and  a71745a );
 a71749a <=( A299  and  (not A298) );
 a71752a <=( A301  and  A300 );
 a71753a <=( a71752a  and  a71749a );
 a71754a <=( a71753a  and  a71746a );
 a71758a <=( (not A168)  and  (not A169) );
 a71759a <=( A170  and  a71758a );
 a71762a <=( (not A166)  and  A167 );
 a71765a <=( A203  and  (not A201) );
 a71766a <=( a71765a  and  a71762a );
 a71767a <=( a71766a  and  a71759a );
 a71771a <=( (not A269)  and  (not A268) );
 a71772a <=( A267  and  a71771a );
 a71775a <=( A299  and  (not A298) );
 a71778a <=( A302  and  A300 );
 a71779a <=( a71778a  and  a71775a );
 a71780a <=( a71779a  and  a71772a );
 a71784a <=( (not A168)  and  (not A169) );
 a71785a <=( A170  and  a71784a );
 a71788a <=( (not A166)  and  A167 );
 a71791a <=( A203  and  (not A201) );
 a71792a <=( a71791a  and  a71788a );
 a71793a <=( a71792a  and  a71785a );
 a71797a <=( A298  and  A268 );
 a71798a <=( (not A267)  and  a71797a );
 a71801a <=( (not A300)  and  (not A299) );
 a71804a <=( (not A302)  and  (not A301) );
 a71805a <=( a71804a  and  a71801a );
 a71806a <=( a71805a  and  a71798a );
 a71810a <=( (not A168)  and  (not A169) );
 a71811a <=( A170  and  a71810a );
 a71814a <=( (not A166)  and  A167 );
 a71817a <=( A203  and  (not A201) );
 a71818a <=( a71817a  and  a71814a );
 a71819a <=( a71818a  and  a71811a );
 a71823a <=( (not A298)  and  A268 );
 a71824a <=( (not A267)  and  a71823a );
 a71827a <=( (not A300)  and  A299 );
 a71830a <=( (not A302)  and  (not A301) );
 a71831a <=( a71830a  and  a71827a );
 a71832a <=( a71831a  and  a71824a );
 a71836a <=( (not A168)  and  (not A169) );
 a71837a <=( A170  and  a71836a );
 a71840a <=( (not A166)  and  A167 );
 a71843a <=( A203  and  (not A201) );
 a71844a <=( a71843a  and  a71840a );
 a71845a <=( a71844a  and  a71837a );
 a71849a <=( A298  and  A269 );
 a71850a <=( (not A267)  and  a71849a );
 a71853a <=( (not A300)  and  (not A299) );
 a71856a <=( (not A302)  and  (not A301) );
 a71857a <=( a71856a  and  a71853a );
 a71858a <=( a71857a  and  a71850a );
 a71862a <=( (not A168)  and  (not A169) );
 a71863a <=( A170  and  a71862a );
 a71866a <=( (not A166)  and  A167 );
 a71869a <=( A203  and  (not A201) );
 a71870a <=( a71869a  and  a71866a );
 a71871a <=( a71870a  and  a71863a );
 a71875a <=( (not A298)  and  A269 );
 a71876a <=( (not A267)  and  a71875a );
 a71879a <=( (not A300)  and  A299 );
 a71882a <=( (not A302)  and  (not A301) );
 a71883a <=( a71882a  and  a71879a );
 a71884a <=( a71883a  and  a71876a );
 a71888a <=( (not A168)  and  (not A169) );
 a71889a <=( A170  and  a71888a );
 a71892a <=( (not A166)  and  A167 );
 a71895a <=( A203  and  (not A201) );
 a71896a <=( a71895a  and  a71892a );
 a71897a <=( a71896a  and  a71889a );
 a71901a <=( A298  and  A266 );
 a71902a <=( A265  and  a71901a );
 a71905a <=( (not A300)  and  (not A299) );
 a71908a <=( (not A302)  and  (not A301) );
 a71909a <=( a71908a  and  a71905a );
 a71910a <=( a71909a  and  a71902a );
 a71914a <=( (not A168)  and  (not A169) );
 a71915a <=( A170  and  a71914a );
 a71918a <=( (not A166)  and  A167 );
 a71921a <=( A203  and  (not A201) );
 a71922a <=( a71921a  and  a71918a );
 a71923a <=( a71922a  and  a71915a );
 a71927a <=( (not A298)  and  A266 );
 a71928a <=( A265  and  a71927a );
 a71931a <=( (not A300)  and  A299 );
 a71934a <=( (not A302)  and  (not A301) );
 a71935a <=( a71934a  and  a71931a );
 a71936a <=( a71935a  and  a71928a );
 a71940a <=( (not A168)  and  (not A169) );
 a71941a <=( A170  and  a71940a );
 a71944a <=( (not A166)  and  A167 );
 a71947a <=( A203  and  (not A201) );
 a71948a <=( a71947a  and  a71944a );
 a71949a <=( a71948a  and  a71941a );
 a71953a <=( A298  and  (not A266) );
 a71954a <=( (not A265)  and  a71953a );
 a71957a <=( (not A300)  and  (not A299) );
 a71960a <=( (not A302)  and  (not A301) );
 a71961a <=( a71960a  and  a71957a );
 a71962a <=( a71961a  and  a71954a );
 a71966a <=( (not A168)  and  (not A169) );
 a71967a <=( A170  and  a71966a );
 a71970a <=( (not A166)  and  A167 );
 a71973a <=( A203  and  (not A201) );
 a71974a <=( a71973a  and  a71970a );
 a71975a <=( a71974a  and  a71967a );
 a71979a <=( (not A298)  and  (not A266) );
 a71980a <=( (not A265)  and  a71979a );
 a71983a <=( (not A300)  and  A299 );
 a71986a <=( (not A302)  and  (not A301) );
 a71987a <=( a71986a  and  a71983a );
 a71988a <=( a71987a  and  a71980a );
 a71992a <=( (not A168)  and  (not A169) );
 a71993a <=( A170  and  a71992a );
 a71996a <=( (not A166)  and  A167 );
 a71999a <=( A200  and  A199 );
 a72000a <=( a71999a  and  a71996a );
 a72001a <=( a72000a  and  a71993a );
 a72005a <=( (not A269)  and  (not A268) );
 a72006a <=( A267  and  a72005a );
 a72009a <=( (not A299)  and  A298 );
 a72012a <=( A301  and  A300 );
 a72013a <=( a72012a  and  a72009a );
 a72014a <=( a72013a  and  a72006a );
 a72018a <=( (not A168)  and  (not A169) );
 a72019a <=( A170  and  a72018a );
 a72022a <=( (not A166)  and  A167 );
 a72025a <=( A200  and  A199 );
 a72026a <=( a72025a  and  a72022a );
 a72027a <=( a72026a  and  a72019a );
 a72031a <=( (not A269)  and  (not A268) );
 a72032a <=( A267  and  a72031a );
 a72035a <=( (not A299)  and  A298 );
 a72038a <=( A302  and  A300 );
 a72039a <=( a72038a  and  a72035a );
 a72040a <=( a72039a  and  a72032a );
 a72044a <=( (not A168)  and  (not A169) );
 a72045a <=( A170  and  a72044a );
 a72048a <=( (not A166)  and  A167 );
 a72051a <=( A200  and  A199 );
 a72052a <=( a72051a  and  a72048a );
 a72053a <=( a72052a  and  a72045a );
 a72057a <=( (not A269)  and  (not A268) );
 a72058a <=( A267  and  a72057a );
 a72061a <=( A299  and  (not A298) );
 a72064a <=( A301  and  A300 );
 a72065a <=( a72064a  and  a72061a );
 a72066a <=( a72065a  and  a72058a );
 a72070a <=( (not A168)  and  (not A169) );
 a72071a <=( A170  and  a72070a );
 a72074a <=( (not A166)  and  A167 );
 a72077a <=( A200  and  A199 );
 a72078a <=( a72077a  and  a72074a );
 a72079a <=( a72078a  and  a72071a );
 a72083a <=( (not A269)  and  (not A268) );
 a72084a <=( A267  and  a72083a );
 a72087a <=( A299  and  (not A298) );
 a72090a <=( A302  and  A300 );
 a72091a <=( a72090a  and  a72087a );
 a72092a <=( a72091a  and  a72084a );
 a72096a <=( (not A168)  and  (not A169) );
 a72097a <=( A170  and  a72096a );
 a72100a <=( (not A166)  and  A167 );
 a72103a <=( A200  and  A199 );
 a72104a <=( a72103a  and  a72100a );
 a72105a <=( a72104a  and  a72097a );
 a72109a <=( A298  and  A268 );
 a72110a <=( (not A267)  and  a72109a );
 a72113a <=( (not A300)  and  (not A299) );
 a72116a <=( (not A302)  and  (not A301) );
 a72117a <=( a72116a  and  a72113a );
 a72118a <=( a72117a  and  a72110a );
 a72122a <=( (not A168)  and  (not A169) );
 a72123a <=( A170  and  a72122a );
 a72126a <=( (not A166)  and  A167 );
 a72129a <=( A200  and  A199 );
 a72130a <=( a72129a  and  a72126a );
 a72131a <=( a72130a  and  a72123a );
 a72135a <=( (not A298)  and  A268 );
 a72136a <=( (not A267)  and  a72135a );
 a72139a <=( (not A300)  and  A299 );
 a72142a <=( (not A302)  and  (not A301) );
 a72143a <=( a72142a  and  a72139a );
 a72144a <=( a72143a  and  a72136a );
 a72148a <=( (not A168)  and  (not A169) );
 a72149a <=( A170  and  a72148a );
 a72152a <=( (not A166)  and  A167 );
 a72155a <=( A200  and  A199 );
 a72156a <=( a72155a  and  a72152a );
 a72157a <=( a72156a  and  a72149a );
 a72161a <=( A298  and  A269 );
 a72162a <=( (not A267)  and  a72161a );
 a72165a <=( (not A300)  and  (not A299) );
 a72168a <=( (not A302)  and  (not A301) );
 a72169a <=( a72168a  and  a72165a );
 a72170a <=( a72169a  and  a72162a );
 a72174a <=( (not A168)  and  (not A169) );
 a72175a <=( A170  and  a72174a );
 a72178a <=( (not A166)  and  A167 );
 a72181a <=( A200  and  A199 );
 a72182a <=( a72181a  and  a72178a );
 a72183a <=( a72182a  and  a72175a );
 a72187a <=( (not A298)  and  A269 );
 a72188a <=( (not A267)  and  a72187a );
 a72191a <=( (not A300)  and  A299 );
 a72194a <=( (not A302)  and  (not A301) );
 a72195a <=( a72194a  and  a72191a );
 a72196a <=( a72195a  and  a72188a );
 a72200a <=( (not A168)  and  (not A169) );
 a72201a <=( A170  and  a72200a );
 a72204a <=( (not A166)  and  A167 );
 a72207a <=( A200  and  A199 );
 a72208a <=( a72207a  and  a72204a );
 a72209a <=( a72208a  and  a72201a );
 a72213a <=( A298  and  A266 );
 a72214a <=( A265  and  a72213a );
 a72217a <=( (not A300)  and  (not A299) );
 a72220a <=( (not A302)  and  (not A301) );
 a72221a <=( a72220a  and  a72217a );
 a72222a <=( a72221a  and  a72214a );
 a72226a <=( (not A168)  and  (not A169) );
 a72227a <=( A170  and  a72226a );
 a72230a <=( (not A166)  and  A167 );
 a72233a <=( A200  and  A199 );
 a72234a <=( a72233a  and  a72230a );
 a72235a <=( a72234a  and  a72227a );
 a72239a <=( (not A298)  and  A266 );
 a72240a <=( A265  and  a72239a );
 a72243a <=( (not A300)  and  A299 );
 a72246a <=( (not A302)  and  (not A301) );
 a72247a <=( a72246a  and  a72243a );
 a72248a <=( a72247a  and  a72240a );
 a72252a <=( (not A168)  and  (not A169) );
 a72253a <=( A170  and  a72252a );
 a72256a <=( (not A166)  and  A167 );
 a72259a <=( A200  and  A199 );
 a72260a <=( a72259a  and  a72256a );
 a72261a <=( a72260a  and  a72253a );
 a72265a <=( A298  and  (not A266) );
 a72266a <=( (not A265)  and  a72265a );
 a72269a <=( (not A300)  and  (not A299) );
 a72272a <=( (not A302)  and  (not A301) );
 a72273a <=( a72272a  and  a72269a );
 a72274a <=( a72273a  and  a72266a );
 a72278a <=( (not A168)  and  (not A169) );
 a72279a <=( A170  and  a72278a );
 a72282a <=( (not A166)  and  A167 );
 a72285a <=( A200  and  A199 );
 a72286a <=( a72285a  and  a72282a );
 a72287a <=( a72286a  and  a72279a );
 a72291a <=( (not A298)  and  (not A266) );
 a72292a <=( (not A265)  and  a72291a );
 a72295a <=( (not A300)  and  A299 );
 a72298a <=( (not A302)  and  (not A301) );
 a72299a <=( a72298a  and  a72295a );
 a72300a <=( a72299a  and  a72292a );
 a72304a <=( (not A168)  and  (not A169) );
 a72305a <=( A170  and  a72304a );
 a72308a <=( (not A166)  and  A167 );
 a72311a <=( (not A200)  and  (not A199) );
 a72312a <=( a72311a  and  a72308a );
 a72313a <=( a72312a  and  a72305a );
 a72317a <=( (not A269)  and  (not A268) );
 a72318a <=( A267  and  a72317a );
 a72321a <=( (not A299)  and  A298 );
 a72324a <=( A301  and  A300 );
 a72325a <=( a72324a  and  a72321a );
 a72326a <=( a72325a  and  a72318a );
 a72330a <=( (not A168)  and  (not A169) );
 a72331a <=( A170  and  a72330a );
 a72334a <=( (not A166)  and  A167 );
 a72337a <=( (not A200)  and  (not A199) );
 a72338a <=( a72337a  and  a72334a );
 a72339a <=( a72338a  and  a72331a );
 a72343a <=( (not A269)  and  (not A268) );
 a72344a <=( A267  and  a72343a );
 a72347a <=( (not A299)  and  A298 );
 a72350a <=( A302  and  A300 );
 a72351a <=( a72350a  and  a72347a );
 a72352a <=( a72351a  and  a72344a );
 a72356a <=( (not A168)  and  (not A169) );
 a72357a <=( A170  and  a72356a );
 a72360a <=( (not A166)  and  A167 );
 a72363a <=( (not A200)  and  (not A199) );
 a72364a <=( a72363a  and  a72360a );
 a72365a <=( a72364a  and  a72357a );
 a72369a <=( (not A269)  and  (not A268) );
 a72370a <=( A267  and  a72369a );
 a72373a <=( A299  and  (not A298) );
 a72376a <=( A301  and  A300 );
 a72377a <=( a72376a  and  a72373a );
 a72378a <=( a72377a  and  a72370a );
 a72382a <=( (not A168)  and  (not A169) );
 a72383a <=( A170  and  a72382a );
 a72386a <=( (not A166)  and  A167 );
 a72389a <=( (not A200)  and  (not A199) );
 a72390a <=( a72389a  and  a72386a );
 a72391a <=( a72390a  and  a72383a );
 a72395a <=( (not A269)  and  (not A268) );
 a72396a <=( A267  and  a72395a );
 a72399a <=( A299  and  (not A298) );
 a72402a <=( A302  and  A300 );
 a72403a <=( a72402a  and  a72399a );
 a72404a <=( a72403a  and  a72396a );
 a72408a <=( (not A168)  and  (not A169) );
 a72409a <=( A170  and  a72408a );
 a72412a <=( (not A166)  and  A167 );
 a72415a <=( (not A200)  and  (not A199) );
 a72416a <=( a72415a  and  a72412a );
 a72417a <=( a72416a  and  a72409a );
 a72421a <=( A298  and  A268 );
 a72422a <=( (not A267)  and  a72421a );
 a72425a <=( (not A300)  and  (not A299) );
 a72428a <=( (not A302)  and  (not A301) );
 a72429a <=( a72428a  and  a72425a );
 a72430a <=( a72429a  and  a72422a );
 a72434a <=( (not A168)  and  (not A169) );
 a72435a <=( A170  and  a72434a );
 a72438a <=( (not A166)  and  A167 );
 a72441a <=( (not A200)  and  (not A199) );
 a72442a <=( a72441a  and  a72438a );
 a72443a <=( a72442a  and  a72435a );
 a72447a <=( (not A298)  and  A268 );
 a72448a <=( (not A267)  and  a72447a );
 a72451a <=( (not A300)  and  A299 );
 a72454a <=( (not A302)  and  (not A301) );
 a72455a <=( a72454a  and  a72451a );
 a72456a <=( a72455a  and  a72448a );
 a72460a <=( (not A168)  and  (not A169) );
 a72461a <=( A170  and  a72460a );
 a72464a <=( (not A166)  and  A167 );
 a72467a <=( (not A200)  and  (not A199) );
 a72468a <=( a72467a  and  a72464a );
 a72469a <=( a72468a  and  a72461a );
 a72473a <=( A298  and  A269 );
 a72474a <=( (not A267)  and  a72473a );
 a72477a <=( (not A300)  and  (not A299) );
 a72480a <=( (not A302)  and  (not A301) );
 a72481a <=( a72480a  and  a72477a );
 a72482a <=( a72481a  and  a72474a );
 a72486a <=( (not A168)  and  (not A169) );
 a72487a <=( A170  and  a72486a );
 a72490a <=( (not A166)  and  A167 );
 a72493a <=( (not A200)  and  (not A199) );
 a72494a <=( a72493a  and  a72490a );
 a72495a <=( a72494a  and  a72487a );
 a72499a <=( (not A298)  and  A269 );
 a72500a <=( (not A267)  and  a72499a );
 a72503a <=( (not A300)  and  A299 );
 a72506a <=( (not A302)  and  (not A301) );
 a72507a <=( a72506a  and  a72503a );
 a72508a <=( a72507a  and  a72500a );
 a72512a <=( (not A168)  and  (not A169) );
 a72513a <=( A170  and  a72512a );
 a72516a <=( (not A166)  and  A167 );
 a72519a <=( (not A200)  and  (not A199) );
 a72520a <=( a72519a  and  a72516a );
 a72521a <=( a72520a  and  a72513a );
 a72525a <=( A298  and  A266 );
 a72526a <=( A265  and  a72525a );
 a72529a <=( (not A300)  and  (not A299) );
 a72532a <=( (not A302)  and  (not A301) );
 a72533a <=( a72532a  and  a72529a );
 a72534a <=( a72533a  and  a72526a );
 a72538a <=( (not A168)  and  (not A169) );
 a72539a <=( A170  and  a72538a );
 a72542a <=( (not A166)  and  A167 );
 a72545a <=( (not A200)  and  (not A199) );
 a72546a <=( a72545a  and  a72542a );
 a72547a <=( a72546a  and  a72539a );
 a72551a <=( (not A298)  and  A266 );
 a72552a <=( A265  and  a72551a );
 a72555a <=( (not A300)  and  A299 );
 a72558a <=( (not A302)  and  (not A301) );
 a72559a <=( a72558a  and  a72555a );
 a72560a <=( a72559a  and  a72552a );
 a72564a <=( (not A168)  and  (not A169) );
 a72565a <=( A170  and  a72564a );
 a72568a <=( (not A166)  and  A167 );
 a72571a <=( (not A200)  and  (not A199) );
 a72572a <=( a72571a  and  a72568a );
 a72573a <=( a72572a  and  a72565a );
 a72577a <=( A298  and  (not A266) );
 a72578a <=( (not A265)  and  a72577a );
 a72581a <=( (not A300)  and  (not A299) );
 a72584a <=( (not A302)  and  (not A301) );
 a72585a <=( a72584a  and  a72581a );
 a72586a <=( a72585a  and  a72578a );
 a72590a <=( (not A168)  and  (not A169) );
 a72591a <=( A170  and  a72590a );
 a72594a <=( (not A166)  and  A167 );
 a72597a <=( (not A200)  and  (not A199) );
 a72598a <=( a72597a  and  a72594a );
 a72599a <=( a72598a  and  a72591a );
 a72603a <=( (not A298)  and  (not A266) );
 a72604a <=( (not A265)  and  a72603a );
 a72607a <=( (not A300)  and  A299 );
 a72610a <=( (not A302)  and  (not A301) );
 a72611a <=( a72610a  and  a72607a );
 a72612a <=( a72611a  and  a72604a );
 a72616a <=( (not A168)  and  (not A169) );
 a72617a <=( A170  and  a72616a );
 a72620a <=( A166  and  (not A167) );
 a72623a <=( (not A202)  and  A201 );
 a72624a <=( a72623a  and  a72620a );
 a72625a <=( a72624a  and  a72617a );
 a72629a <=( A268  and  (not A267) );
 a72630a <=( (not A203)  and  a72629a );
 a72633a <=( (not A299)  and  A298 );
 a72636a <=( A301  and  A300 );
 a72637a <=( a72636a  and  a72633a );
 a72638a <=( a72637a  and  a72630a );
 a72642a <=( (not A168)  and  (not A169) );
 a72643a <=( A170  and  a72642a );
 a72646a <=( A166  and  (not A167) );
 a72649a <=( (not A202)  and  A201 );
 a72650a <=( a72649a  and  a72646a );
 a72651a <=( a72650a  and  a72643a );
 a72655a <=( A268  and  (not A267) );
 a72656a <=( (not A203)  and  a72655a );
 a72659a <=( (not A299)  and  A298 );
 a72662a <=( A302  and  A300 );
 a72663a <=( a72662a  and  a72659a );
 a72664a <=( a72663a  and  a72656a );
 a72668a <=( (not A168)  and  (not A169) );
 a72669a <=( A170  and  a72668a );
 a72672a <=( A166  and  (not A167) );
 a72675a <=( (not A202)  and  A201 );
 a72676a <=( a72675a  and  a72672a );
 a72677a <=( a72676a  and  a72669a );
 a72681a <=( A268  and  (not A267) );
 a72682a <=( (not A203)  and  a72681a );
 a72685a <=( A299  and  (not A298) );
 a72688a <=( A301  and  A300 );
 a72689a <=( a72688a  and  a72685a );
 a72690a <=( a72689a  and  a72682a );
 a72694a <=( (not A168)  and  (not A169) );
 a72695a <=( A170  and  a72694a );
 a72698a <=( A166  and  (not A167) );
 a72701a <=( (not A202)  and  A201 );
 a72702a <=( a72701a  and  a72698a );
 a72703a <=( a72702a  and  a72695a );
 a72707a <=( A268  and  (not A267) );
 a72708a <=( (not A203)  and  a72707a );
 a72711a <=( A299  and  (not A298) );
 a72714a <=( A302  and  A300 );
 a72715a <=( a72714a  and  a72711a );
 a72716a <=( a72715a  and  a72708a );
 a72720a <=( (not A168)  and  (not A169) );
 a72721a <=( A170  and  a72720a );
 a72724a <=( A166  and  (not A167) );
 a72727a <=( (not A202)  and  A201 );
 a72728a <=( a72727a  and  a72724a );
 a72729a <=( a72728a  and  a72721a );
 a72733a <=( A269  and  (not A267) );
 a72734a <=( (not A203)  and  a72733a );
 a72737a <=( (not A299)  and  A298 );
 a72740a <=( A301  and  A300 );
 a72741a <=( a72740a  and  a72737a );
 a72742a <=( a72741a  and  a72734a );
 a72746a <=( (not A168)  and  (not A169) );
 a72747a <=( A170  and  a72746a );
 a72750a <=( A166  and  (not A167) );
 a72753a <=( (not A202)  and  A201 );
 a72754a <=( a72753a  and  a72750a );
 a72755a <=( a72754a  and  a72747a );
 a72759a <=( A269  and  (not A267) );
 a72760a <=( (not A203)  and  a72759a );
 a72763a <=( (not A299)  and  A298 );
 a72766a <=( A302  and  A300 );
 a72767a <=( a72766a  and  a72763a );
 a72768a <=( a72767a  and  a72760a );
 a72772a <=( (not A168)  and  (not A169) );
 a72773a <=( A170  and  a72772a );
 a72776a <=( A166  and  (not A167) );
 a72779a <=( (not A202)  and  A201 );
 a72780a <=( a72779a  and  a72776a );
 a72781a <=( a72780a  and  a72773a );
 a72785a <=( A269  and  (not A267) );
 a72786a <=( (not A203)  and  a72785a );
 a72789a <=( A299  and  (not A298) );
 a72792a <=( A301  and  A300 );
 a72793a <=( a72792a  and  a72789a );
 a72794a <=( a72793a  and  a72786a );
 a72798a <=( (not A168)  and  (not A169) );
 a72799a <=( A170  and  a72798a );
 a72802a <=( A166  and  (not A167) );
 a72805a <=( (not A202)  and  A201 );
 a72806a <=( a72805a  and  a72802a );
 a72807a <=( a72806a  and  a72799a );
 a72811a <=( A269  and  (not A267) );
 a72812a <=( (not A203)  and  a72811a );
 a72815a <=( A299  and  (not A298) );
 a72818a <=( A302  and  A300 );
 a72819a <=( a72818a  and  a72815a );
 a72820a <=( a72819a  and  a72812a );
 a72824a <=( (not A168)  and  (not A169) );
 a72825a <=( A170  and  a72824a );
 a72828a <=( A166  and  (not A167) );
 a72831a <=( (not A202)  and  A201 );
 a72832a <=( a72831a  and  a72828a );
 a72833a <=( a72832a  and  a72825a );
 a72837a <=( A266  and  A265 );
 a72838a <=( (not A203)  and  a72837a );
 a72841a <=( (not A299)  and  A298 );
 a72844a <=( A301  and  A300 );
 a72845a <=( a72844a  and  a72841a );
 a72846a <=( a72845a  and  a72838a );
 a72850a <=( (not A168)  and  (not A169) );
 a72851a <=( A170  and  a72850a );
 a72854a <=( A166  and  (not A167) );
 a72857a <=( (not A202)  and  A201 );
 a72858a <=( a72857a  and  a72854a );
 a72859a <=( a72858a  and  a72851a );
 a72863a <=( A266  and  A265 );
 a72864a <=( (not A203)  and  a72863a );
 a72867a <=( (not A299)  and  A298 );
 a72870a <=( A302  and  A300 );
 a72871a <=( a72870a  and  a72867a );
 a72872a <=( a72871a  and  a72864a );
 a72876a <=( (not A168)  and  (not A169) );
 a72877a <=( A170  and  a72876a );
 a72880a <=( A166  and  (not A167) );
 a72883a <=( (not A202)  and  A201 );
 a72884a <=( a72883a  and  a72880a );
 a72885a <=( a72884a  and  a72877a );
 a72889a <=( A266  and  A265 );
 a72890a <=( (not A203)  and  a72889a );
 a72893a <=( A299  and  (not A298) );
 a72896a <=( A301  and  A300 );
 a72897a <=( a72896a  and  a72893a );
 a72898a <=( a72897a  and  a72890a );
 a72902a <=( (not A168)  and  (not A169) );
 a72903a <=( A170  and  a72902a );
 a72906a <=( A166  and  (not A167) );
 a72909a <=( (not A202)  and  A201 );
 a72910a <=( a72909a  and  a72906a );
 a72911a <=( a72910a  and  a72903a );
 a72915a <=( A266  and  A265 );
 a72916a <=( (not A203)  and  a72915a );
 a72919a <=( A299  and  (not A298) );
 a72922a <=( A302  and  A300 );
 a72923a <=( a72922a  and  a72919a );
 a72924a <=( a72923a  and  a72916a );
 a72928a <=( (not A168)  and  (not A169) );
 a72929a <=( A170  and  a72928a );
 a72932a <=( A166  and  (not A167) );
 a72935a <=( (not A202)  and  A201 );
 a72936a <=( a72935a  and  a72932a );
 a72937a <=( a72936a  and  a72929a );
 a72941a <=( (not A266)  and  (not A265) );
 a72942a <=( (not A203)  and  a72941a );
 a72945a <=( (not A299)  and  A298 );
 a72948a <=( A301  and  A300 );
 a72949a <=( a72948a  and  a72945a );
 a72950a <=( a72949a  and  a72942a );
 a72954a <=( (not A168)  and  (not A169) );
 a72955a <=( A170  and  a72954a );
 a72958a <=( A166  and  (not A167) );
 a72961a <=( (not A202)  and  A201 );
 a72962a <=( a72961a  and  a72958a );
 a72963a <=( a72962a  and  a72955a );
 a72967a <=( (not A266)  and  (not A265) );
 a72968a <=( (not A203)  and  a72967a );
 a72971a <=( (not A299)  and  A298 );
 a72974a <=( A302  and  A300 );
 a72975a <=( a72974a  and  a72971a );
 a72976a <=( a72975a  and  a72968a );
 a72980a <=( (not A168)  and  (not A169) );
 a72981a <=( A170  and  a72980a );
 a72984a <=( A166  and  (not A167) );
 a72987a <=( (not A202)  and  A201 );
 a72988a <=( a72987a  and  a72984a );
 a72989a <=( a72988a  and  a72981a );
 a72993a <=( (not A266)  and  (not A265) );
 a72994a <=( (not A203)  and  a72993a );
 a72997a <=( A299  and  (not A298) );
 a73000a <=( A301  and  A300 );
 a73001a <=( a73000a  and  a72997a );
 a73002a <=( a73001a  and  a72994a );
 a73006a <=( (not A168)  and  (not A169) );
 a73007a <=( A170  and  a73006a );
 a73010a <=( A166  and  (not A167) );
 a73013a <=( (not A202)  and  A201 );
 a73014a <=( a73013a  and  a73010a );
 a73015a <=( a73014a  and  a73007a );
 a73019a <=( (not A266)  and  (not A265) );
 a73020a <=( (not A203)  and  a73019a );
 a73023a <=( A299  and  (not A298) );
 a73026a <=( A302  and  A300 );
 a73027a <=( a73026a  and  a73023a );
 a73028a <=( a73027a  and  a73020a );
 a73032a <=( (not A168)  and  (not A169) );
 a73033a <=( A170  and  a73032a );
 a73036a <=( A166  and  (not A167) );
 a73039a <=( A202  and  (not A201) );
 a73040a <=( a73039a  and  a73036a );
 a73041a <=( a73040a  and  a73033a );
 a73045a <=( (not A269)  and  (not A268) );
 a73046a <=( A267  and  a73045a );
 a73049a <=( (not A299)  and  A298 );
 a73052a <=( A301  and  A300 );
 a73053a <=( a73052a  and  a73049a );
 a73054a <=( a73053a  and  a73046a );
 a73058a <=( (not A168)  and  (not A169) );
 a73059a <=( A170  and  a73058a );
 a73062a <=( A166  and  (not A167) );
 a73065a <=( A202  and  (not A201) );
 a73066a <=( a73065a  and  a73062a );
 a73067a <=( a73066a  and  a73059a );
 a73071a <=( (not A269)  and  (not A268) );
 a73072a <=( A267  and  a73071a );
 a73075a <=( (not A299)  and  A298 );
 a73078a <=( A302  and  A300 );
 a73079a <=( a73078a  and  a73075a );
 a73080a <=( a73079a  and  a73072a );
 a73084a <=( (not A168)  and  (not A169) );
 a73085a <=( A170  and  a73084a );
 a73088a <=( A166  and  (not A167) );
 a73091a <=( A202  and  (not A201) );
 a73092a <=( a73091a  and  a73088a );
 a73093a <=( a73092a  and  a73085a );
 a73097a <=( (not A269)  and  (not A268) );
 a73098a <=( A267  and  a73097a );
 a73101a <=( A299  and  (not A298) );
 a73104a <=( A301  and  A300 );
 a73105a <=( a73104a  and  a73101a );
 a73106a <=( a73105a  and  a73098a );
 a73110a <=( (not A168)  and  (not A169) );
 a73111a <=( A170  and  a73110a );
 a73114a <=( A166  and  (not A167) );
 a73117a <=( A202  and  (not A201) );
 a73118a <=( a73117a  and  a73114a );
 a73119a <=( a73118a  and  a73111a );
 a73123a <=( (not A269)  and  (not A268) );
 a73124a <=( A267  and  a73123a );
 a73127a <=( A299  and  (not A298) );
 a73130a <=( A302  and  A300 );
 a73131a <=( a73130a  and  a73127a );
 a73132a <=( a73131a  and  a73124a );
 a73136a <=( (not A168)  and  (not A169) );
 a73137a <=( A170  and  a73136a );
 a73140a <=( A166  and  (not A167) );
 a73143a <=( A202  and  (not A201) );
 a73144a <=( a73143a  and  a73140a );
 a73145a <=( a73144a  and  a73137a );
 a73149a <=( A298  and  A268 );
 a73150a <=( (not A267)  and  a73149a );
 a73153a <=( (not A300)  and  (not A299) );
 a73156a <=( (not A302)  and  (not A301) );
 a73157a <=( a73156a  and  a73153a );
 a73158a <=( a73157a  and  a73150a );
 a73162a <=( (not A168)  and  (not A169) );
 a73163a <=( A170  and  a73162a );
 a73166a <=( A166  and  (not A167) );
 a73169a <=( A202  and  (not A201) );
 a73170a <=( a73169a  and  a73166a );
 a73171a <=( a73170a  and  a73163a );
 a73175a <=( (not A298)  and  A268 );
 a73176a <=( (not A267)  and  a73175a );
 a73179a <=( (not A300)  and  A299 );
 a73182a <=( (not A302)  and  (not A301) );
 a73183a <=( a73182a  and  a73179a );
 a73184a <=( a73183a  and  a73176a );
 a73188a <=( (not A168)  and  (not A169) );
 a73189a <=( A170  and  a73188a );
 a73192a <=( A166  and  (not A167) );
 a73195a <=( A202  and  (not A201) );
 a73196a <=( a73195a  and  a73192a );
 a73197a <=( a73196a  and  a73189a );
 a73201a <=( A298  and  A269 );
 a73202a <=( (not A267)  and  a73201a );
 a73205a <=( (not A300)  and  (not A299) );
 a73208a <=( (not A302)  and  (not A301) );
 a73209a <=( a73208a  and  a73205a );
 a73210a <=( a73209a  and  a73202a );
 a73214a <=( (not A168)  and  (not A169) );
 a73215a <=( A170  and  a73214a );
 a73218a <=( A166  and  (not A167) );
 a73221a <=( A202  and  (not A201) );
 a73222a <=( a73221a  and  a73218a );
 a73223a <=( a73222a  and  a73215a );
 a73227a <=( (not A298)  and  A269 );
 a73228a <=( (not A267)  and  a73227a );
 a73231a <=( (not A300)  and  A299 );
 a73234a <=( (not A302)  and  (not A301) );
 a73235a <=( a73234a  and  a73231a );
 a73236a <=( a73235a  and  a73228a );
 a73240a <=( (not A168)  and  (not A169) );
 a73241a <=( A170  and  a73240a );
 a73244a <=( A166  and  (not A167) );
 a73247a <=( A202  and  (not A201) );
 a73248a <=( a73247a  and  a73244a );
 a73249a <=( a73248a  and  a73241a );
 a73253a <=( A298  and  A266 );
 a73254a <=( A265  and  a73253a );
 a73257a <=( (not A300)  and  (not A299) );
 a73260a <=( (not A302)  and  (not A301) );
 a73261a <=( a73260a  and  a73257a );
 a73262a <=( a73261a  and  a73254a );
 a73266a <=( (not A168)  and  (not A169) );
 a73267a <=( A170  and  a73266a );
 a73270a <=( A166  and  (not A167) );
 a73273a <=( A202  and  (not A201) );
 a73274a <=( a73273a  and  a73270a );
 a73275a <=( a73274a  and  a73267a );
 a73279a <=( (not A298)  and  A266 );
 a73280a <=( A265  and  a73279a );
 a73283a <=( (not A300)  and  A299 );
 a73286a <=( (not A302)  and  (not A301) );
 a73287a <=( a73286a  and  a73283a );
 a73288a <=( a73287a  and  a73280a );
 a73292a <=( (not A168)  and  (not A169) );
 a73293a <=( A170  and  a73292a );
 a73296a <=( A166  and  (not A167) );
 a73299a <=( A202  and  (not A201) );
 a73300a <=( a73299a  and  a73296a );
 a73301a <=( a73300a  and  a73293a );
 a73305a <=( A298  and  (not A266) );
 a73306a <=( (not A265)  and  a73305a );
 a73309a <=( (not A300)  and  (not A299) );
 a73312a <=( (not A302)  and  (not A301) );
 a73313a <=( a73312a  and  a73309a );
 a73314a <=( a73313a  and  a73306a );
 a73318a <=( (not A168)  and  (not A169) );
 a73319a <=( A170  and  a73318a );
 a73322a <=( A166  and  (not A167) );
 a73325a <=( A202  and  (not A201) );
 a73326a <=( a73325a  and  a73322a );
 a73327a <=( a73326a  and  a73319a );
 a73331a <=( (not A298)  and  (not A266) );
 a73332a <=( (not A265)  and  a73331a );
 a73335a <=( (not A300)  and  A299 );
 a73338a <=( (not A302)  and  (not A301) );
 a73339a <=( a73338a  and  a73335a );
 a73340a <=( a73339a  and  a73332a );
 a73344a <=( (not A168)  and  (not A169) );
 a73345a <=( A170  and  a73344a );
 a73348a <=( A166  and  (not A167) );
 a73351a <=( A203  and  (not A201) );
 a73352a <=( a73351a  and  a73348a );
 a73353a <=( a73352a  and  a73345a );
 a73357a <=( (not A269)  and  (not A268) );
 a73358a <=( A267  and  a73357a );
 a73361a <=( (not A299)  and  A298 );
 a73364a <=( A301  and  A300 );
 a73365a <=( a73364a  and  a73361a );
 a73366a <=( a73365a  and  a73358a );
 a73370a <=( (not A168)  and  (not A169) );
 a73371a <=( A170  and  a73370a );
 a73374a <=( A166  and  (not A167) );
 a73377a <=( A203  and  (not A201) );
 a73378a <=( a73377a  and  a73374a );
 a73379a <=( a73378a  and  a73371a );
 a73383a <=( (not A269)  and  (not A268) );
 a73384a <=( A267  and  a73383a );
 a73387a <=( (not A299)  and  A298 );
 a73390a <=( A302  and  A300 );
 a73391a <=( a73390a  and  a73387a );
 a73392a <=( a73391a  and  a73384a );
 a73396a <=( (not A168)  and  (not A169) );
 a73397a <=( A170  and  a73396a );
 a73400a <=( A166  and  (not A167) );
 a73403a <=( A203  and  (not A201) );
 a73404a <=( a73403a  and  a73400a );
 a73405a <=( a73404a  and  a73397a );
 a73409a <=( (not A269)  and  (not A268) );
 a73410a <=( A267  and  a73409a );
 a73413a <=( A299  and  (not A298) );
 a73416a <=( A301  and  A300 );
 a73417a <=( a73416a  and  a73413a );
 a73418a <=( a73417a  and  a73410a );
 a73422a <=( (not A168)  and  (not A169) );
 a73423a <=( A170  and  a73422a );
 a73426a <=( A166  and  (not A167) );
 a73429a <=( A203  and  (not A201) );
 a73430a <=( a73429a  and  a73426a );
 a73431a <=( a73430a  and  a73423a );
 a73435a <=( (not A269)  and  (not A268) );
 a73436a <=( A267  and  a73435a );
 a73439a <=( A299  and  (not A298) );
 a73442a <=( A302  and  A300 );
 a73443a <=( a73442a  and  a73439a );
 a73444a <=( a73443a  and  a73436a );
 a73448a <=( (not A168)  and  (not A169) );
 a73449a <=( A170  and  a73448a );
 a73452a <=( A166  and  (not A167) );
 a73455a <=( A203  and  (not A201) );
 a73456a <=( a73455a  and  a73452a );
 a73457a <=( a73456a  and  a73449a );
 a73461a <=( A298  and  A268 );
 a73462a <=( (not A267)  and  a73461a );
 a73465a <=( (not A300)  and  (not A299) );
 a73468a <=( (not A302)  and  (not A301) );
 a73469a <=( a73468a  and  a73465a );
 a73470a <=( a73469a  and  a73462a );
 a73474a <=( (not A168)  and  (not A169) );
 a73475a <=( A170  and  a73474a );
 a73478a <=( A166  and  (not A167) );
 a73481a <=( A203  and  (not A201) );
 a73482a <=( a73481a  and  a73478a );
 a73483a <=( a73482a  and  a73475a );
 a73487a <=( (not A298)  and  A268 );
 a73488a <=( (not A267)  and  a73487a );
 a73491a <=( (not A300)  and  A299 );
 a73494a <=( (not A302)  and  (not A301) );
 a73495a <=( a73494a  and  a73491a );
 a73496a <=( a73495a  and  a73488a );
 a73500a <=( (not A168)  and  (not A169) );
 a73501a <=( A170  and  a73500a );
 a73504a <=( A166  and  (not A167) );
 a73507a <=( A203  and  (not A201) );
 a73508a <=( a73507a  and  a73504a );
 a73509a <=( a73508a  and  a73501a );
 a73513a <=( A298  and  A269 );
 a73514a <=( (not A267)  and  a73513a );
 a73517a <=( (not A300)  and  (not A299) );
 a73520a <=( (not A302)  and  (not A301) );
 a73521a <=( a73520a  and  a73517a );
 a73522a <=( a73521a  and  a73514a );
 a73526a <=( (not A168)  and  (not A169) );
 a73527a <=( A170  and  a73526a );
 a73530a <=( A166  and  (not A167) );
 a73533a <=( A203  and  (not A201) );
 a73534a <=( a73533a  and  a73530a );
 a73535a <=( a73534a  and  a73527a );
 a73539a <=( (not A298)  and  A269 );
 a73540a <=( (not A267)  and  a73539a );
 a73543a <=( (not A300)  and  A299 );
 a73546a <=( (not A302)  and  (not A301) );
 a73547a <=( a73546a  and  a73543a );
 a73548a <=( a73547a  and  a73540a );
 a73552a <=( (not A168)  and  (not A169) );
 a73553a <=( A170  and  a73552a );
 a73556a <=( A166  and  (not A167) );
 a73559a <=( A203  and  (not A201) );
 a73560a <=( a73559a  and  a73556a );
 a73561a <=( a73560a  and  a73553a );
 a73565a <=( A298  and  A266 );
 a73566a <=( A265  and  a73565a );
 a73569a <=( (not A300)  and  (not A299) );
 a73572a <=( (not A302)  and  (not A301) );
 a73573a <=( a73572a  and  a73569a );
 a73574a <=( a73573a  and  a73566a );
 a73578a <=( (not A168)  and  (not A169) );
 a73579a <=( A170  and  a73578a );
 a73582a <=( A166  and  (not A167) );
 a73585a <=( A203  and  (not A201) );
 a73586a <=( a73585a  and  a73582a );
 a73587a <=( a73586a  and  a73579a );
 a73591a <=( (not A298)  and  A266 );
 a73592a <=( A265  and  a73591a );
 a73595a <=( (not A300)  and  A299 );
 a73598a <=( (not A302)  and  (not A301) );
 a73599a <=( a73598a  and  a73595a );
 a73600a <=( a73599a  and  a73592a );
 a73604a <=( (not A168)  and  (not A169) );
 a73605a <=( A170  and  a73604a );
 a73608a <=( A166  and  (not A167) );
 a73611a <=( A203  and  (not A201) );
 a73612a <=( a73611a  and  a73608a );
 a73613a <=( a73612a  and  a73605a );
 a73617a <=( A298  and  (not A266) );
 a73618a <=( (not A265)  and  a73617a );
 a73621a <=( (not A300)  and  (not A299) );
 a73624a <=( (not A302)  and  (not A301) );
 a73625a <=( a73624a  and  a73621a );
 a73626a <=( a73625a  and  a73618a );
 a73630a <=( (not A168)  and  (not A169) );
 a73631a <=( A170  and  a73630a );
 a73634a <=( A166  and  (not A167) );
 a73637a <=( A203  and  (not A201) );
 a73638a <=( a73637a  and  a73634a );
 a73639a <=( a73638a  and  a73631a );
 a73643a <=( (not A298)  and  (not A266) );
 a73644a <=( (not A265)  and  a73643a );
 a73647a <=( (not A300)  and  A299 );
 a73650a <=( (not A302)  and  (not A301) );
 a73651a <=( a73650a  and  a73647a );
 a73652a <=( a73651a  and  a73644a );
 a73656a <=( (not A168)  and  (not A169) );
 a73657a <=( A170  and  a73656a );
 a73660a <=( A166  and  (not A167) );
 a73663a <=( A200  and  A199 );
 a73664a <=( a73663a  and  a73660a );
 a73665a <=( a73664a  and  a73657a );
 a73669a <=( (not A269)  and  (not A268) );
 a73670a <=( A267  and  a73669a );
 a73673a <=( (not A299)  and  A298 );
 a73676a <=( A301  and  A300 );
 a73677a <=( a73676a  and  a73673a );
 a73678a <=( a73677a  and  a73670a );
 a73682a <=( (not A168)  and  (not A169) );
 a73683a <=( A170  and  a73682a );
 a73686a <=( A166  and  (not A167) );
 a73689a <=( A200  and  A199 );
 a73690a <=( a73689a  and  a73686a );
 a73691a <=( a73690a  and  a73683a );
 a73695a <=( (not A269)  and  (not A268) );
 a73696a <=( A267  and  a73695a );
 a73699a <=( (not A299)  and  A298 );
 a73702a <=( A302  and  A300 );
 a73703a <=( a73702a  and  a73699a );
 a73704a <=( a73703a  and  a73696a );
 a73708a <=( (not A168)  and  (not A169) );
 a73709a <=( A170  and  a73708a );
 a73712a <=( A166  and  (not A167) );
 a73715a <=( A200  and  A199 );
 a73716a <=( a73715a  and  a73712a );
 a73717a <=( a73716a  and  a73709a );
 a73721a <=( (not A269)  and  (not A268) );
 a73722a <=( A267  and  a73721a );
 a73725a <=( A299  and  (not A298) );
 a73728a <=( A301  and  A300 );
 a73729a <=( a73728a  and  a73725a );
 a73730a <=( a73729a  and  a73722a );
 a73734a <=( (not A168)  and  (not A169) );
 a73735a <=( A170  and  a73734a );
 a73738a <=( A166  and  (not A167) );
 a73741a <=( A200  and  A199 );
 a73742a <=( a73741a  and  a73738a );
 a73743a <=( a73742a  and  a73735a );
 a73747a <=( (not A269)  and  (not A268) );
 a73748a <=( A267  and  a73747a );
 a73751a <=( A299  and  (not A298) );
 a73754a <=( A302  and  A300 );
 a73755a <=( a73754a  and  a73751a );
 a73756a <=( a73755a  and  a73748a );
 a73760a <=( (not A168)  and  (not A169) );
 a73761a <=( A170  and  a73760a );
 a73764a <=( A166  and  (not A167) );
 a73767a <=( A200  and  A199 );
 a73768a <=( a73767a  and  a73764a );
 a73769a <=( a73768a  and  a73761a );
 a73773a <=( A298  and  A268 );
 a73774a <=( (not A267)  and  a73773a );
 a73777a <=( (not A300)  and  (not A299) );
 a73780a <=( (not A302)  and  (not A301) );
 a73781a <=( a73780a  and  a73777a );
 a73782a <=( a73781a  and  a73774a );
 a73786a <=( (not A168)  and  (not A169) );
 a73787a <=( A170  and  a73786a );
 a73790a <=( A166  and  (not A167) );
 a73793a <=( A200  and  A199 );
 a73794a <=( a73793a  and  a73790a );
 a73795a <=( a73794a  and  a73787a );
 a73799a <=( (not A298)  and  A268 );
 a73800a <=( (not A267)  and  a73799a );
 a73803a <=( (not A300)  and  A299 );
 a73806a <=( (not A302)  and  (not A301) );
 a73807a <=( a73806a  and  a73803a );
 a73808a <=( a73807a  and  a73800a );
 a73812a <=( (not A168)  and  (not A169) );
 a73813a <=( A170  and  a73812a );
 a73816a <=( A166  and  (not A167) );
 a73819a <=( A200  and  A199 );
 a73820a <=( a73819a  and  a73816a );
 a73821a <=( a73820a  and  a73813a );
 a73825a <=( A298  and  A269 );
 a73826a <=( (not A267)  and  a73825a );
 a73829a <=( (not A300)  and  (not A299) );
 a73832a <=( (not A302)  and  (not A301) );
 a73833a <=( a73832a  and  a73829a );
 a73834a <=( a73833a  and  a73826a );
 a73838a <=( (not A168)  and  (not A169) );
 a73839a <=( A170  and  a73838a );
 a73842a <=( A166  and  (not A167) );
 a73845a <=( A200  and  A199 );
 a73846a <=( a73845a  and  a73842a );
 a73847a <=( a73846a  and  a73839a );
 a73851a <=( (not A298)  and  A269 );
 a73852a <=( (not A267)  and  a73851a );
 a73855a <=( (not A300)  and  A299 );
 a73858a <=( (not A302)  and  (not A301) );
 a73859a <=( a73858a  and  a73855a );
 a73860a <=( a73859a  and  a73852a );
 a73864a <=( (not A168)  and  (not A169) );
 a73865a <=( A170  and  a73864a );
 a73868a <=( A166  and  (not A167) );
 a73871a <=( A200  and  A199 );
 a73872a <=( a73871a  and  a73868a );
 a73873a <=( a73872a  and  a73865a );
 a73877a <=( A298  and  A266 );
 a73878a <=( A265  and  a73877a );
 a73881a <=( (not A300)  and  (not A299) );
 a73884a <=( (not A302)  and  (not A301) );
 a73885a <=( a73884a  and  a73881a );
 a73886a <=( a73885a  and  a73878a );
 a73890a <=( (not A168)  and  (not A169) );
 a73891a <=( A170  and  a73890a );
 a73894a <=( A166  and  (not A167) );
 a73897a <=( A200  and  A199 );
 a73898a <=( a73897a  and  a73894a );
 a73899a <=( a73898a  and  a73891a );
 a73903a <=( (not A298)  and  A266 );
 a73904a <=( A265  and  a73903a );
 a73907a <=( (not A300)  and  A299 );
 a73910a <=( (not A302)  and  (not A301) );
 a73911a <=( a73910a  and  a73907a );
 a73912a <=( a73911a  and  a73904a );
 a73916a <=( (not A168)  and  (not A169) );
 a73917a <=( A170  and  a73916a );
 a73920a <=( A166  and  (not A167) );
 a73923a <=( A200  and  A199 );
 a73924a <=( a73923a  and  a73920a );
 a73925a <=( a73924a  and  a73917a );
 a73929a <=( A298  and  (not A266) );
 a73930a <=( (not A265)  and  a73929a );
 a73933a <=( (not A300)  and  (not A299) );
 a73936a <=( (not A302)  and  (not A301) );
 a73937a <=( a73936a  and  a73933a );
 a73938a <=( a73937a  and  a73930a );
 a73942a <=( (not A168)  and  (not A169) );
 a73943a <=( A170  and  a73942a );
 a73946a <=( A166  and  (not A167) );
 a73949a <=( A200  and  A199 );
 a73950a <=( a73949a  and  a73946a );
 a73951a <=( a73950a  and  a73943a );
 a73955a <=( (not A298)  and  (not A266) );
 a73956a <=( (not A265)  and  a73955a );
 a73959a <=( (not A300)  and  A299 );
 a73962a <=( (not A302)  and  (not A301) );
 a73963a <=( a73962a  and  a73959a );
 a73964a <=( a73963a  and  a73956a );
 a73968a <=( (not A168)  and  (not A169) );
 a73969a <=( A170  and  a73968a );
 a73972a <=( A166  and  (not A167) );
 a73975a <=( (not A200)  and  (not A199) );
 a73976a <=( a73975a  and  a73972a );
 a73977a <=( a73976a  and  a73969a );
 a73981a <=( (not A269)  and  (not A268) );
 a73982a <=( A267  and  a73981a );
 a73985a <=( (not A299)  and  A298 );
 a73988a <=( A301  and  A300 );
 a73989a <=( a73988a  and  a73985a );
 a73990a <=( a73989a  and  a73982a );
 a73994a <=( (not A168)  and  (not A169) );
 a73995a <=( A170  and  a73994a );
 a73998a <=( A166  and  (not A167) );
 a74001a <=( (not A200)  and  (not A199) );
 a74002a <=( a74001a  and  a73998a );
 a74003a <=( a74002a  and  a73995a );
 a74007a <=( (not A269)  and  (not A268) );
 a74008a <=( A267  and  a74007a );
 a74011a <=( (not A299)  and  A298 );
 a74014a <=( A302  and  A300 );
 a74015a <=( a74014a  and  a74011a );
 a74016a <=( a74015a  and  a74008a );
 a74020a <=( (not A168)  and  (not A169) );
 a74021a <=( A170  and  a74020a );
 a74024a <=( A166  and  (not A167) );
 a74027a <=( (not A200)  and  (not A199) );
 a74028a <=( a74027a  and  a74024a );
 a74029a <=( a74028a  and  a74021a );
 a74033a <=( (not A269)  and  (not A268) );
 a74034a <=( A267  and  a74033a );
 a74037a <=( A299  and  (not A298) );
 a74040a <=( A301  and  A300 );
 a74041a <=( a74040a  and  a74037a );
 a74042a <=( a74041a  and  a74034a );
 a74046a <=( (not A168)  and  (not A169) );
 a74047a <=( A170  and  a74046a );
 a74050a <=( A166  and  (not A167) );
 a74053a <=( (not A200)  and  (not A199) );
 a74054a <=( a74053a  and  a74050a );
 a74055a <=( a74054a  and  a74047a );
 a74059a <=( (not A269)  and  (not A268) );
 a74060a <=( A267  and  a74059a );
 a74063a <=( A299  and  (not A298) );
 a74066a <=( A302  and  A300 );
 a74067a <=( a74066a  and  a74063a );
 a74068a <=( a74067a  and  a74060a );
 a74072a <=( (not A168)  and  (not A169) );
 a74073a <=( A170  and  a74072a );
 a74076a <=( A166  and  (not A167) );
 a74079a <=( (not A200)  and  (not A199) );
 a74080a <=( a74079a  and  a74076a );
 a74081a <=( a74080a  and  a74073a );
 a74085a <=( A298  and  A268 );
 a74086a <=( (not A267)  and  a74085a );
 a74089a <=( (not A300)  and  (not A299) );
 a74092a <=( (not A302)  and  (not A301) );
 a74093a <=( a74092a  and  a74089a );
 a74094a <=( a74093a  and  a74086a );
 a74098a <=( (not A168)  and  (not A169) );
 a74099a <=( A170  and  a74098a );
 a74102a <=( A166  and  (not A167) );
 a74105a <=( (not A200)  and  (not A199) );
 a74106a <=( a74105a  and  a74102a );
 a74107a <=( a74106a  and  a74099a );
 a74111a <=( (not A298)  and  A268 );
 a74112a <=( (not A267)  and  a74111a );
 a74115a <=( (not A300)  and  A299 );
 a74118a <=( (not A302)  and  (not A301) );
 a74119a <=( a74118a  and  a74115a );
 a74120a <=( a74119a  and  a74112a );
 a74124a <=( (not A168)  and  (not A169) );
 a74125a <=( A170  and  a74124a );
 a74128a <=( A166  and  (not A167) );
 a74131a <=( (not A200)  and  (not A199) );
 a74132a <=( a74131a  and  a74128a );
 a74133a <=( a74132a  and  a74125a );
 a74137a <=( A298  and  A269 );
 a74138a <=( (not A267)  and  a74137a );
 a74141a <=( (not A300)  and  (not A299) );
 a74144a <=( (not A302)  and  (not A301) );
 a74145a <=( a74144a  and  a74141a );
 a74146a <=( a74145a  and  a74138a );
 a74150a <=( (not A168)  and  (not A169) );
 a74151a <=( A170  and  a74150a );
 a74154a <=( A166  and  (not A167) );
 a74157a <=( (not A200)  and  (not A199) );
 a74158a <=( a74157a  and  a74154a );
 a74159a <=( a74158a  and  a74151a );
 a74163a <=( (not A298)  and  A269 );
 a74164a <=( (not A267)  and  a74163a );
 a74167a <=( (not A300)  and  A299 );
 a74170a <=( (not A302)  and  (not A301) );
 a74171a <=( a74170a  and  a74167a );
 a74172a <=( a74171a  and  a74164a );
 a74176a <=( (not A168)  and  (not A169) );
 a74177a <=( A170  and  a74176a );
 a74180a <=( A166  and  (not A167) );
 a74183a <=( (not A200)  and  (not A199) );
 a74184a <=( a74183a  and  a74180a );
 a74185a <=( a74184a  and  a74177a );
 a74189a <=( A298  and  A266 );
 a74190a <=( A265  and  a74189a );
 a74193a <=( (not A300)  and  (not A299) );
 a74196a <=( (not A302)  and  (not A301) );
 a74197a <=( a74196a  and  a74193a );
 a74198a <=( a74197a  and  a74190a );
 a74202a <=( (not A168)  and  (not A169) );
 a74203a <=( A170  and  a74202a );
 a74206a <=( A166  and  (not A167) );
 a74209a <=( (not A200)  and  (not A199) );
 a74210a <=( a74209a  and  a74206a );
 a74211a <=( a74210a  and  a74203a );
 a74215a <=( (not A298)  and  A266 );
 a74216a <=( A265  and  a74215a );
 a74219a <=( (not A300)  and  A299 );
 a74222a <=( (not A302)  and  (not A301) );
 a74223a <=( a74222a  and  a74219a );
 a74224a <=( a74223a  and  a74216a );
 a74228a <=( (not A168)  and  (not A169) );
 a74229a <=( A170  and  a74228a );
 a74232a <=( A166  and  (not A167) );
 a74235a <=( (not A200)  and  (not A199) );
 a74236a <=( a74235a  and  a74232a );
 a74237a <=( a74236a  and  a74229a );
 a74241a <=( A298  and  (not A266) );
 a74242a <=( (not A265)  and  a74241a );
 a74245a <=( (not A300)  and  (not A299) );
 a74248a <=( (not A302)  and  (not A301) );
 a74249a <=( a74248a  and  a74245a );
 a74250a <=( a74249a  and  a74242a );
 a74254a <=( (not A168)  and  (not A169) );
 a74255a <=( A170  and  a74254a );
 a74258a <=( A166  and  (not A167) );
 a74261a <=( (not A200)  and  (not A199) );
 a74262a <=( a74261a  and  a74258a );
 a74263a <=( a74262a  and  a74255a );
 a74267a <=( (not A298)  and  (not A266) );
 a74268a <=( (not A265)  and  a74267a );
 a74271a <=( (not A300)  and  A299 );
 a74274a <=( (not A302)  and  (not A301) );
 a74275a <=( a74274a  and  a74271a );
 a74276a <=( a74275a  and  a74268a );
 a74280a <=( (not A199)  and  A166 );
 a74281a <=( A167  and  a74280a );
 a74284a <=( (not A201)  and  A200 );
 a74287a <=( (not A203)  and  (not A202) );
 a74288a <=( a74287a  and  a74284a );
 a74289a <=( a74288a  and  a74281a );
 a74292a <=( (not A268)  and  A267 );
 a74295a <=( A298  and  (not A269) );
 a74296a <=( a74295a  and  a74292a );
 a74299a <=( (not A300)  and  (not A299) );
 a74302a <=( (not A302)  and  (not A301) );
 a74303a <=( a74302a  and  a74299a );
 a74304a <=( a74303a  and  a74296a );
 a74308a <=( (not A199)  and  A166 );
 a74309a <=( A167  and  a74308a );
 a74312a <=( (not A201)  and  A200 );
 a74315a <=( (not A203)  and  (not A202) );
 a74316a <=( a74315a  and  a74312a );
 a74317a <=( a74316a  and  a74309a );
 a74320a <=( (not A268)  and  A267 );
 a74323a <=( (not A298)  and  (not A269) );
 a74324a <=( a74323a  and  a74320a );
 a74327a <=( (not A300)  and  A299 );
 a74330a <=( (not A302)  and  (not A301) );
 a74331a <=( a74330a  and  a74327a );
 a74332a <=( a74331a  and  a74324a );
 a74336a <=( A199  and  A166 );
 a74337a <=( A167  and  a74336a );
 a74340a <=( (not A201)  and  (not A200) );
 a74343a <=( (not A203)  and  (not A202) );
 a74344a <=( a74343a  and  a74340a );
 a74345a <=( a74344a  and  a74337a );
 a74348a <=( (not A268)  and  A267 );
 a74351a <=( A298  and  (not A269) );
 a74352a <=( a74351a  and  a74348a );
 a74355a <=( (not A300)  and  (not A299) );
 a74358a <=( (not A302)  and  (not A301) );
 a74359a <=( a74358a  and  a74355a );
 a74360a <=( a74359a  and  a74352a );
 a74364a <=( A199  and  A166 );
 a74365a <=( A167  and  a74364a );
 a74368a <=( (not A201)  and  (not A200) );
 a74371a <=( (not A203)  and  (not A202) );
 a74372a <=( a74371a  and  a74368a );
 a74373a <=( a74372a  and  a74365a );
 a74376a <=( (not A268)  and  A267 );
 a74379a <=( (not A298)  and  (not A269) );
 a74380a <=( a74379a  and  a74376a );
 a74383a <=( (not A300)  and  A299 );
 a74386a <=( (not A302)  and  (not A301) );
 a74387a <=( a74386a  and  a74383a );
 a74388a <=( a74387a  and  a74380a );
 a74392a <=( (not A199)  and  (not A166) );
 a74393a <=( (not A167)  and  a74392a );
 a74396a <=( (not A201)  and  A200 );
 a74399a <=( (not A203)  and  (not A202) );
 a74400a <=( a74399a  and  a74396a );
 a74401a <=( a74400a  and  a74393a );
 a74404a <=( (not A268)  and  A267 );
 a74407a <=( A298  and  (not A269) );
 a74408a <=( a74407a  and  a74404a );
 a74411a <=( (not A300)  and  (not A299) );
 a74414a <=( (not A302)  and  (not A301) );
 a74415a <=( a74414a  and  a74411a );
 a74416a <=( a74415a  and  a74408a );
 a74420a <=( (not A199)  and  (not A166) );
 a74421a <=( (not A167)  and  a74420a );
 a74424a <=( (not A201)  and  A200 );
 a74427a <=( (not A203)  and  (not A202) );
 a74428a <=( a74427a  and  a74424a );
 a74429a <=( a74428a  and  a74421a );
 a74432a <=( (not A268)  and  A267 );
 a74435a <=( (not A298)  and  (not A269) );
 a74436a <=( a74435a  and  a74432a );
 a74439a <=( (not A300)  and  A299 );
 a74442a <=( (not A302)  and  (not A301) );
 a74443a <=( a74442a  and  a74439a );
 a74444a <=( a74443a  and  a74436a );
 a74448a <=( A199  and  (not A166) );
 a74449a <=( (not A167)  and  a74448a );
 a74452a <=( (not A201)  and  (not A200) );
 a74455a <=( (not A203)  and  (not A202) );
 a74456a <=( a74455a  and  a74452a );
 a74457a <=( a74456a  and  a74449a );
 a74460a <=( (not A268)  and  A267 );
 a74463a <=( A298  and  (not A269) );
 a74464a <=( a74463a  and  a74460a );
 a74467a <=( (not A300)  and  (not A299) );
 a74470a <=( (not A302)  and  (not A301) );
 a74471a <=( a74470a  and  a74467a );
 a74472a <=( a74471a  and  a74464a );
 a74476a <=( A199  and  (not A166) );
 a74477a <=( (not A167)  and  a74476a );
 a74480a <=( (not A201)  and  (not A200) );
 a74483a <=( (not A203)  and  (not A202) );
 a74484a <=( a74483a  and  a74480a );
 a74485a <=( a74484a  and  a74477a );
 a74488a <=( (not A268)  and  A267 );
 a74491a <=( (not A298)  and  (not A269) );
 a74492a <=( a74491a  and  a74488a );
 a74495a <=( (not A300)  and  A299 );
 a74498a <=( (not A302)  and  (not A301) );
 a74499a <=( a74498a  and  a74495a );
 a74500a <=( a74499a  and  a74492a );
 a74504a <=( A167  and  A168 );
 a74505a <=( (not A170)  and  a74504a );
 a74508a <=( A201  and  (not A166) );
 a74511a <=( (not A203)  and  (not A202) );
 a74512a <=( a74511a  and  a74508a );
 a74513a <=( a74512a  and  a74505a );
 a74516a <=( (not A268)  and  A267 );
 a74519a <=( A298  and  (not A269) );
 a74520a <=( a74519a  and  a74516a );
 a74523a <=( (not A300)  and  (not A299) );
 a74526a <=( (not A302)  and  (not A301) );
 a74527a <=( a74526a  and  a74523a );
 a74528a <=( a74527a  and  a74520a );
 a74532a <=( A167  and  A168 );
 a74533a <=( (not A170)  and  a74532a );
 a74536a <=( A201  and  (not A166) );
 a74539a <=( (not A203)  and  (not A202) );
 a74540a <=( a74539a  and  a74536a );
 a74541a <=( a74540a  and  a74533a );
 a74544a <=( (not A268)  and  A267 );
 a74547a <=( (not A298)  and  (not A269) );
 a74548a <=( a74547a  and  a74544a );
 a74551a <=( (not A300)  and  A299 );
 a74554a <=( (not A302)  and  (not A301) );
 a74555a <=( a74554a  and  a74551a );
 a74556a <=( a74555a  and  a74548a );
 a74560a <=( A167  and  A168 );
 a74561a <=( (not A170)  and  a74560a );
 a74564a <=( (not A199)  and  (not A166) );
 a74567a <=( A201  and  A200 );
 a74568a <=( a74567a  and  a74564a );
 a74569a <=( a74568a  and  a74561a );
 a74572a <=( (not A265)  and  A202 );
 a74575a <=( A267  and  A266 );
 a74576a <=( a74575a  and  a74572a );
 a74579a <=( A300  and  A268 );
 a74582a <=( (not A302)  and  (not A301) );
 a74583a <=( a74582a  and  a74579a );
 a74584a <=( a74583a  and  a74576a );
 a74588a <=( A167  and  A168 );
 a74589a <=( (not A170)  and  a74588a );
 a74592a <=( (not A199)  and  (not A166) );
 a74595a <=( A201  and  A200 );
 a74596a <=( a74595a  and  a74592a );
 a74597a <=( a74596a  and  a74589a );
 a74600a <=( (not A265)  and  A202 );
 a74603a <=( A267  and  A266 );
 a74604a <=( a74603a  and  a74600a );
 a74607a <=( A300  and  A269 );
 a74610a <=( (not A302)  and  (not A301) );
 a74611a <=( a74610a  and  a74607a );
 a74612a <=( a74611a  and  a74604a );
 a74616a <=( A167  and  A168 );
 a74617a <=( (not A170)  and  a74616a );
 a74620a <=( (not A199)  and  (not A166) );
 a74623a <=( A201  and  A200 );
 a74624a <=( a74623a  and  a74620a );
 a74625a <=( a74624a  and  a74617a );
 a74628a <=( (not A265)  and  A202 );
 a74631a <=( (not A267)  and  A266 );
 a74632a <=( a74631a  and  a74628a );
 a74635a <=( (not A269)  and  (not A268) );
 a74638a <=( A301  and  (not A300) );
 a74639a <=( a74638a  and  a74635a );
 a74640a <=( a74639a  and  a74632a );
 a74644a <=( A167  and  A168 );
 a74645a <=( (not A170)  and  a74644a );
 a74648a <=( (not A199)  and  (not A166) );
 a74651a <=( A201  and  A200 );
 a74652a <=( a74651a  and  a74648a );
 a74653a <=( a74652a  and  a74645a );
 a74656a <=( (not A265)  and  A202 );
 a74659a <=( (not A267)  and  A266 );
 a74660a <=( a74659a  and  a74656a );
 a74663a <=( (not A269)  and  (not A268) );
 a74666a <=( A302  and  (not A300) );
 a74667a <=( a74666a  and  a74663a );
 a74668a <=( a74667a  and  a74660a );
 a74672a <=( A167  and  A168 );
 a74673a <=( (not A170)  and  a74672a );
 a74676a <=( (not A199)  and  (not A166) );
 a74679a <=( A201  and  A200 );
 a74680a <=( a74679a  and  a74676a );
 a74681a <=( a74680a  and  a74673a );
 a74684a <=( (not A265)  and  A202 );
 a74687a <=( (not A267)  and  A266 );
 a74688a <=( a74687a  and  a74684a );
 a74691a <=( (not A269)  and  (not A268) );
 a74694a <=( A299  and  A298 );
 a74695a <=( a74694a  and  a74691a );
 a74696a <=( a74695a  and  a74688a );
 a74700a <=( A167  and  A168 );
 a74701a <=( (not A170)  and  a74700a );
 a74704a <=( (not A199)  and  (not A166) );
 a74707a <=( A201  and  A200 );
 a74708a <=( a74707a  and  a74704a );
 a74709a <=( a74708a  and  a74701a );
 a74712a <=( (not A265)  and  A202 );
 a74715a <=( (not A267)  and  A266 );
 a74716a <=( a74715a  and  a74712a );
 a74719a <=( (not A269)  and  (not A268) );
 a74722a <=( (not A299)  and  (not A298) );
 a74723a <=( a74722a  and  a74719a );
 a74724a <=( a74723a  and  a74716a );
 a74728a <=( A167  and  A168 );
 a74729a <=( (not A170)  and  a74728a );
 a74732a <=( (not A199)  and  (not A166) );
 a74735a <=( A201  and  A200 );
 a74736a <=( a74735a  and  a74732a );
 a74737a <=( a74736a  and  a74729a );
 a74740a <=( A265  and  A202 );
 a74743a <=( A267  and  (not A266) );
 a74744a <=( a74743a  and  a74740a );
 a74747a <=( A300  and  A268 );
 a74750a <=( (not A302)  and  (not A301) );
 a74751a <=( a74750a  and  a74747a );
 a74752a <=( a74751a  and  a74744a );
 a74756a <=( A167  and  A168 );
 a74757a <=( (not A170)  and  a74756a );
 a74760a <=( (not A199)  and  (not A166) );
 a74763a <=( A201  and  A200 );
 a74764a <=( a74763a  and  a74760a );
 a74765a <=( a74764a  and  a74757a );
 a74768a <=( A265  and  A202 );
 a74771a <=( A267  and  (not A266) );
 a74772a <=( a74771a  and  a74768a );
 a74775a <=( A300  and  A269 );
 a74778a <=( (not A302)  and  (not A301) );
 a74779a <=( a74778a  and  a74775a );
 a74780a <=( a74779a  and  a74772a );
 a74784a <=( A167  and  A168 );
 a74785a <=( (not A170)  and  a74784a );
 a74788a <=( (not A199)  and  (not A166) );
 a74791a <=( A201  and  A200 );
 a74792a <=( a74791a  and  a74788a );
 a74793a <=( a74792a  and  a74785a );
 a74796a <=( A265  and  A202 );
 a74799a <=( (not A267)  and  (not A266) );
 a74800a <=( a74799a  and  a74796a );
 a74803a <=( (not A269)  and  (not A268) );
 a74806a <=( A301  and  (not A300) );
 a74807a <=( a74806a  and  a74803a );
 a74808a <=( a74807a  and  a74800a );
 a74812a <=( A167  and  A168 );
 a74813a <=( (not A170)  and  a74812a );
 a74816a <=( (not A199)  and  (not A166) );
 a74819a <=( A201  and  A200 );
 a74820a <=( a74819a  and  a74816a );
 a74821a <=( a74820a  and  a74813a );
 a74824a <=( A265  and  A202 );
 a74827a <=( (not A267)  and  (not A266) );
 a74828a <=( a74827a  and  a74824a );
 a74831a <=( (not A269)  and  (not A268) );
 a74834a <=( A302  and  (not A300) );
 a74835a <=( a74834a  and  a74831a );
 a74836a <=( a74835a  and  a74828a );
 a74840a <=( A167  and  A168 );
 a74841a <=( (not A170)  and  a74840a );
 a74844a <=( (not A199)  and  (not A166) );
 a74847a <=( A201  and  A200 );
 a74848a <=( a74847a  and  a74844a );
 a74849a <=( a74848a  and  a74841a );
 a74852a <=( A265  and  A202 );
 a74855a <=( (not A267)  and  (not A266) );
 a74856a <=( a74855a  and  a74852a );
 a74859a <=( (not A269)  and  (not A268) );
 a74862a <=( A299  and  A298 );
 a74863a <=( a74862a  and  a74859a );
 a74864a <=( a74863a  and  a74856a );
 a74868a <=( A167  and  A168 );
 a74869a <=( (not A170)  and  a74868a );
 a74872a <=( (not A199)  and  (not A166) );
 a74875a <=( A201  and  A200 );
 a74876a <=( a74875a  and  a74872a );
 a74877a <=( a74876a  and  a74869a );
 a74880a <=( A265  and  A202 );
 a74883a <=( (not A267)  and  (not A266) );
 a74884a <=( a74883a  and  a74880a );
 a74887a <=( (not A269)  and  (not A268) );
 a74890a <=( (not A299)  and  (not A298) );
 a74891a <=( a74890a  and  a74887a );
 a74892a <=( a74891a  and  a74884a );
 a74896a <=( A167  and  A168 );
 a74897a <=( (not A170)  and  a74896a );
 a74900a <=( (not A199)  and  (not A166) );
 a74903a <=( A201  and  A200 );
 a74904a <=( a74903a  and  a74900a );
 a74905a <=( a74904a  and  a74897a );
 a74908a <=( (not A265)  and  A203 );
 a74911a <=( A267  and  A266 );
 a74912a <=( a74911a  and  a74908a );
 a74915a <=( A300  and  A268 );
 a74918a <=( (not A302)  and  (not A301) );
 a74919a <=( a74918a  and  a74915a );
 a74920a <=( a74919a  and  a74912a );
 a74924a <=( A167  and  A168 );
 a74925a <=( (not A170)  and  a74924a );
 a74928a <=( (not A199)  and  (not A166) );
 a74931a <=( A201  and  A200 );
 a74932a <=( a74931a  and  a74928a );
 a74933a <=( a74932a  and  a74925a );
 a74936a <=( (not A265)  and  A203 );
 a74939a <=( A267  and  A266 );
 a74940a <=( a74939a  and  a74936a );
 a74943a <=( A300  and  A269 );
 a74946a <=( (not A302)  and  (not A301) );
 a74947a <=( a74946a  and  a74943a );
 a74948a <=( a74947a  and  a74940a );
 a74952a <=( A167  and  A168 );
 a74953a <=( (not A170)  and  a74952a );
 a74956a <=( (not A199)  and  (not A166) );
 a74959a <=( A201  and  A200 );
 a74960a <=( a74959a  and  a74956a );
 a74961a <=( a74960a  and  a74953a );
 a74964a <=( (not A265)  and  A203 );
 a74967a <=( (not A267)  and  A266 );
 a74968a <=( a74967a  and  a74964a );
 a74971a <=( (not A269)  and  (not A268) );
 a74974a <=( A301  and  (not A300) );
 a74975a <=( a74974a  and  a74971a );
 a74976a <=( a74975a  and  a74968a );
 a74980a <=( A167  and  A168 );
 a74981a <=( (not A170)  and  a74980a );
 a74984a <=( (not A199)  and  (not A166) );
 a74987a <=( A201  and  A200 );
 a74988a <=( a74987a  and  a74984a );
 a74989a <=( a74988a  and  a74981a );
 a74992a <=( (not A265)  and  A203 );
 a74995a <=( (not A267)  and  A266 );
 a74996a <=( a74995a  and  a74992a );
 a74999a <=( (not A269)  and  (not A268) );
 a75002a <=( A302  and  (not A300) );
 a75003a <=( a75002a  and  a74999a );
 a75004a <=( a75003a  and  a74996a );
 a75008a <=( A167  and  A168 );
 a75009a <=( (not A170)  and  a75008a );
 a75012a <=( (not A199)  and  (not A166) );
 a75015a <=( A201  and  A200 );
 a75016a <=( a75015a  and  a75012a );
 a75017a <=( a75016a  and  a75009a );
 a75020a <=( (not A265)  and  A203 );
 a75023a <=( (not A267)  and  A266 );
 a75024a <=( a75023a  and  a75020a );
 a75027a <=( (not A269)  and  (not A268) );
 a75030a <=( A299  and  A298 );
 a75031a <=( a75030a  and  a75027a );
 a75032a <=( a75031a  and  a75024a );
 a75036a <=( A167  and  A168 );
 a75037a <=( (not A170)  and  a75036a );
 a75040a <=( (not A199)  and  (not A166) );
 a75043a <=( A201  and  A200 );
 a75044a <=( a75043a  and  a75040a );
 a75045a <=( a75044a  and  a75037a );
 a75048a <=( (not A265)  and  A203 );
 a75051a <=( (not A267)  and  A266 );
 a75052a <=( a75051a  and  a75048a );
 a75055a <=( (not A269)  and  (not A268) );
 a75058a <=( (not A299)  and  (not A298) );
 a75059a <=( a75058a  and  a75055a );
 a75060a <=( a75059a  and  a75052a );
 a75064a <=( A167  and  A168 );
 a75065a <=( (not A170)  and  a75064a );
 a75068a <=( (not A199)  and  (not A166) );
 a75071a <=( A201  and  A200 );
 a75072a <=( a75071a  and  a75068a );
 a75073a <=( a75072a  and  a75065a );
 a75076a <=( A265  and  A203 );
 a75079a <=( A267  and  (not A266) );
 a75080a <=( a75079a  and  a75076a );
 a75083a <=( A300  and  A268 );
 a75086a <=( (not A302)  and  (not A301) );
 a75087a <=( a75086a  and  a75083a );
 a75088a <=( a75087a  and  a75080a );
 a75092a <=( A167  and  A168 );
 a75093a <=( (not A170)  and  a75092a );
 a75096a <=( (not A199)  and  (not A166) );
 a75099a <=( A201  and  A200 );
 a75100a <=( a75099a  and  a75096a );
 a75101a <=( a75100a  and  a75093a );
 a75104a <=( A265  and  A203 );
 a75107a <=( A267  and  (not A266) );
 a75108a <=( a75107a  and  a75104a );
 a75111a <=( A300  and  A269 );
 a75114a <=( (not A302)  and  (not A301) );
 a75115a <=( a75114a  and  a75111a );
 a75116a <=( a75115a  and  a75108a );
 a75120a <=( A167  and  A168 );
 a75121a <=( (not A170)  and  a75120a );
 a75124a <=( (not A199)  and  (not A166) );
 a75127a <=( A201  and  A200 );
 a75128a <=( a75127a  and  a75124a );
 a75129a <=( a75128a  and  a75121a );
 a75132a <=( A265  and  A203 );
 a75135a <=( (not A267)  and  (not A266) );
 a75136a <=( a75135a  and  a75132a );
 a75139a <=( (not A269)  and  (not A268) );
 a75142a <=( A301  and  (not A300) );
 a75143a <=( a75142a  and  a75139a );
 a75144a <=( a75143a  and  a75136a );
 a75148a <=( A167  and  A168 );
 a75149a <=( (not A170)  and  a75148a );
 a75152a <=( (not A199)  and  (not A166) );
 a75155a <=( A201  and  A200 );
 a75156a <=( a75155a  and  a75152a );
 a75157a <=( a75156a  and  a75149a );
 a75160a <=( A265  and  A203 );
 a75163a <=( (not A267)  and  (not A266) );
 a75164a <=( a75163a  and  a75160a );
 a75167a <=( (not A269)  and  (not A268) );
 a75170a <=( A302  and  (not A300) );
 a75171a <=( a75170a  and  a75167a );
 a75172a <=( a75171a  and  a75164a );
 a75176a <=( A167  and  A168 );
 a75177a <=( (not A170)  and  a75176a );
 a75180a <=( (not A199)  and  (not A166) );
 a75183a <=( A201  and  A200 );
 a75184a <=( a75183a  and  a75180a );
 a75185a <=( a75184a  and  a75177a );
 a75188a <=( A265  and  A203 );
 a75191a <=( (not A267)  and  (not A266) );
 a75192a <=( a75191a  and  a75188a );
 a75195a <=( (not A269)  and  (not A268) );
 a75198a <=( A299  and  A298 );
 a75199a <=( a75198a  and  a75195a );
 a75200a <=( a75199a  and  a75192a );
 a75204a <=( A167  and  A168 );
 a75205a <=( (not A170)  and  a75204a );
 a75208a <=( (not A199)  and  (not A166) );
 a75211a <=( A201  and  A200 );
 a75212a <=( a75211a  and  a75208a );
 a75213a <=( a75212a  and  a75205a );
 a75216a <=( A265  and  A203 );
 a75219a <=( (not A267)  and  (not A266) );
 a75220a <=( a75219a  and  a75216a );
 a75223a <=( (not A269)  and  (not A268) );
 a75226a <=( (not A299)  and  (not A298) );
 a75227a <=( a75226a  and  a75223a );
 a75228a <=( a75227a  and  a75220a );
 a75232a <=( A167  and  A168 );
 a75233a <=( (not A170)  and  a75232a );
 a75236a <=( (not A199)  and  (not A166) );
 a75239a <=( (not A201)  and  A200 );
 a75240a <=( a75239a  and  a75236a );
 a75241a <=( a75240a  and  a75233a );
 a75244a <=( (not A203)  and  (not A202) );
 a75247a <=( A266  and  (not A265) );
 a75248a <=( a75247a  and  a75244a );
 a75251a <=( A268  and  A267 );
 a75254a <=( A301  and  (not A300) );
 a75255a <=( a75254a  and  a75251a );
 a75256a <=( a75255a  and  a75248a );
 a75260a <=( A167  and  A168 );
 a75261a <=( (not A170)  and  a75260a );
 a75264a <=( (not A199)  and  (not A166) );
 a75267a <=( (not A201)  and  A200 );
 a75268a <=( a75267a  and  a75264a );
 a75269a <=( a75268a  and  a75261a );
 a75272a <=( (not A203)  and  (not A202) );
 a75275a <=( A266  and  (not A265) );
 a75276a <=( a75275a  and  a75272a );
 a75279a <=( A268  and  A267 );
 a75282a <=( A302  and  (not A300) );
 a75283a <=( a75282a  and  a75279a );
 a75284a <=( a75283a  and  a75276a );
 a75288a <=( A167  and  A168 );
 a75289a <=( (not A170)  and  a75288a );
 a75292a <=( (not A199)  and  (not A166) );
 a75295a <=( (not A201)  and  A200 );
 a75296a <=( a75295a  and  a75292a );
 a75297a <=( a75296a  and  a75289a );
 a75300a <=( (not A203)  and  (not A202) );
 a75303a <=( A266  and  (not A265) );
 a75304a <=( a75303a  and  a75300a );
 a75307a <=( A268  and  A267 );
 a75310a <=( A299  and  A298 );
 a75311a <=( a75310a  and  a75307a );
 a75312a <=( a75311a  and  a75304a );
 a75316a <=( A167  and  A168 );
 a75317a <=( (not A170)  and  a75316a );
 a75320a <=( (not A199)  and  (not A166) );
 a75323a <=( (not A201)  and  A200 );
 a75324a <=( a75323a  and  a75320a );
 a75325a <=( a75324a  and  a75317a );
 a75328a <=( (not A203)  and  (not A202) );
 a75331a <=( A266  and  (not A265) );
 a75332a <=( a75331a  and  a75328a );
 a75335a <=( A268  and  A267 );
 a75338a <=( (not A299)  and  (not A298) );
 a75339a <=( a75338a  and  a75335a );
 a75340a <=( a75339a  and  a75332a );
 a75344a <=( A167  and  A168 );
 a75345a <=( (not A170)  and  a75344a );
 a75348a <=( (not A199)  and  (not A166) );
 a75351a <=( (not A201)  and  A200 );
 a75352a <=( a75351a  and  a75348a );
 a75353a <=( a75352a  and  a75345a );
 a75356a <=( (not A203)  and  (not A202) );
 a75359a <=( A266  and  (not A265) );
 a75360a <=( a75359a  and  a75356a );
 a75363a <=( A269  and  A267 );
 a75366a <=( A301  and  (not A300) );
 a75367a <=( a75366a  and  a75363a );
 a75368a <=( a75367a  and  a75360a );
 a75372a <=( A167  and  A168 );
 a75373a <=( (not A170)  and  a75372a );
 a75376a <=( (not A199)  and  (not A166) );
 a75379a <=( (not A201)  and  A200 );
 a75380a <=( a75379a  and  a75376a );
 a75381a <=( a75380a  and  a75373a );
 a75384a <=( (not A203)  and  (not A202) );
 a75387a <=( A266  and  (not A265) );
 a75388a <=( a75387a  and  a75384a );
 a75391a <=( A269  and  A267 );
 a75394a <=( A302  and  (not A300) );
 a75395a <=( a75394a  and  a75391a );
 a75396a <=( a75395a  and  a75388a );
 a75400a <=( A167  and  A168 );
 a75401a <=( (not A170)  and  a75400a );
 a75404a <=( (not A199)  and  (not A166) );
 a75407a <=( (not A201)  and  A200 );
 a75408a <=( a75407a  and  a75404a );
 a75409a <=( a75408a  and  a75401a );
 a75412a <=( (not A203)  and  (not A202) );
 a75415a <=( A266  and  (not A265) );
 a75416a <=( a75415a  and  a75412a );
 a75419a <=( A269  and  A267 );
 a75422a <=( A299  and  A298 );
 a75423a <=( a75422a  and  a75419a );
 a75424a <=( a75423a  and  a75416a );
 a75428a <=( A167  and  A168 );
 a75429a <=( (not A170)  and  a75428a );
 a75432a <=( (not A199)  and  (not A166) );
 a75435a <=( (not A201)  and  A200 );
 a75436a <=( a75435a  and  a75432a );
 a75437a <=( a75436a  and  a75429a );
 a75440a <=( (not A203)  and  (not A202) );
 a75443a <=( A266  and  (not A265) );
 a75444a <=( a75443a  and  a75440a );
 a75447a <=( A269  and  A267 );
 a75450a <=( (not A299)  and  (not A298) );
 a75451a <=( a75450a  and  a75447a );
 a75452a <=( a75451a  and  a75444a );
 a75456a <=( A167  and  A168 );
 a75457a <=( (not A170)  and  a75456a );
 a75460a <=( (not A199)  and  (not A166) );
 a75463a <=( (not A201)  and  A200 );
 a75464a <=( a75463a  and  a75460a );
 a75465a <=( a75464a  and  a75457a );
 a75468a <=( (not A203)  and  (not A202) );
 a75471a <=( (not A266)  and  A265 );
 a75472a <=( a75471a  and  a75468a );
 a75475a <=( A268  and  A267 );
 a75478a <=( A301  and  (not A300) );
 a75479a <=( a75478a  and  a75475a );
 a75480a <=( a75479a  and  a75472a );
 a75484a <=( A167  and  A168 );
 a75485a <=( (not A170)  and  a75484a );
 a75488a <=( (not A199)  and  (not A166) );
 a75491a <=( (not A201)  and  A200 );
 a75492a <=( a75491a  and  a75488a );
 a75493a <=( a75492a  and  a75485a );
 a75496a <=( (not A203)  and  (not A202) );
 a75499a <=( (not A266)  and  A265 );
 a75500a <=( a75499a  and  a75496a );
 a75503a <=( A268  and  A267 );
 a75506a <=( A302  and  (not A300) );
 a75507a <=( a75506a  and  a75503a );
 a75508a <=( a75507a  and  a75500a );
 a75512a <=( A167  and  A168 );
 a75513a <=( (not A170)  and  a75512a );
 a75516a <=( (not A199)  and  (not A166) );
 a75519a <=( (not A201)  and  A200 );
 a75520a <=( a75519a  and  a75516a );
 a75521a <=( a75520a  and  a75513a );
 a75524a <=( (not A203)  and  (not A202) );
 a75527a <=( (not A266)  and  A265 );
 a75528a <=( a75527a  and  a75524a );
 a75531a <=( A268  and  A267 );
 a75534a <=( A299  and  A298 );
 a75535a <=( a75534a  and  a75531a );
 a75536a <=( a75535a  and  a75528a );
 a75540a <=( A167  and  A168 );
 a75541a <=( (not A170)  and  a75540a );
 a75544a <=( (not A199)  and  (not A166) );
 a75547a <=( (not A201)  and  A200 );
 a75548a <=( a75547a  and  a75544a );
 a75549a <=( a75548a  and  a75541a );
 a75552a <=( (not A203)  and  (not A202) );
 a75555a <=( (not A266)  and  A265 );
 a75556a <=( a75555a  and  a75552a );
 a75559a <=( A268  and  A267 );
 a75562a <=( (not A299)  and  (not A298) );
 a75563a <=( a75562a  and  a75559a );
 a75564a <=( a75563a  and  a75556a );
 a75568a <=( A167  and  A168 );
 a75569a <=( (not A170)  and  a75568a );
 a75572a <=( (not A199)  and  (not A166) );
 a75575a <=( (not A201)  and  A200 );
 a75576a <=( a75575a  and  a75572a );
 a75577a <=( a75576a  and  a75569a );
 a75580a <=( (not A203)  and  (not A202) );
 a75583a <=( (not A266)  and  A265 );
 a75584a <=( a75583a  and  a75580a );
 a75587a <=( A269  and  A267 );
 a75590a <=( A301  and  (not A300) );
 a75591a <=( a75590a  and  a75587a );
 a75592a <=( a75591a  and  a75584a );
 a75596a <=( A167  and  A168 );
 a75597a <=( (not A170)  and  a75596a );
 a75600a <=( (not A199)  and  (not A166) );
 a75603a <=( (not A201)  and  A200 );
 a75604a <=( a75603a  and  a75600a );
 a75605a <=( a75604a  and  a75597a );
 a75608a <=( (not A203)  and  (not A202) );
 a75611a <=( (not A266)  and  A265 );
 a75612a <=( a75611a  and  a75608a );
 a75615a <=( A269  and  A267 );
 a75618a <=( A302  and  (not A300) );
 a75619a <=( a75618a  and  a75615a );
 a75620a <=( a75619a  and  a75612a );
 a75624a <=( A167  and  A168 );
 a75625a <=( (not A170)  and  a75624a );
 a75628a <=( (not A199)  and  (not A166) );
 a75631a <=( (not A201)  and  A200 );
 a75632a <=( a75631a  and  a75628a );
 a75633a <=( a75632a  and  a75625a );
 a75636a <=( (not A203)  and  (not A202) );
 a75639a <=( (not A266)  and  A265 );
 a75640a <=( a75639a  and  a75636a );
 a75643a <=( A269  and  A267 );
 a75646a <=( A299  and  A298 );
 a75647a <=( a75646a  and  a75643a );
 a75648a <=( a75647a  and  a75640a );
 a75652a <=( A167  and  A168 );
 a75653a <=( (not A170)  and  a75652a );
 a75656a <=( (not A199)  and  (not A166) );
 a75659a <=( (not A201)  and  A200 );
 a75660a <=( a75659a  and  a75656a );
 a75661a <=( a75660a  and  a75653a );
 a75664a <=( (not A203)  and  (not A202) );
 a75667a <=( (not A266)  and  A265 );
 a75668a <=( a75667a  and  a75664a );
 a75671a <=( A269  and  A267 );
 a75674a <=( (not A299)  and  (not A298) );
 a75675a <=( a75674a  and  a75671a );
 a75676a <=( a75675a  and  a75668a );
 a75680a <=( A167  and  A168 );
 a75681a <=( (not A170)  and  a75680a );
 a75684a <=( A199  and  (not A166) );
 a75687a <=( A201  and  (not A200) );
 a75688a <=( a75687a  and  a75684a );
 a75689a <=( a75688a  and  a75681a );
 a75692a <=( (not A265)  and  A202 );
 a75695a <=( A267  and  A266 );
 a75696a <=( a75695a  and  a75692a );
 a75699a <=( A300  and  A268 );
 a75702a <=( (not A302)  and  (not A301) );
 a75703a <=( a75702a  and  a75699a );
 a75704a <=( a75703a  and  a75696a );
 a75708a <=( A167  and  A168 );
 a75709a <=( (not A170)  and  a75708a );
 a75712a <=( A199  and  (not A166) );
 a75715a <=( A201  and  (not A200) );
 a75716a <=( a75715a  and  a75712a );
 a75717a <=( a75716a  and  a75709a );
 a75720a <=( (not A265)  and  A202 );
 a75723a <=( A267  and  A266 );
 a75724a <=( a75723a  and  a75720a );
 a75727a <=( A300  and  A269 );
 a75730a <=( (not A302)  and  (not A301) );
 a75731a <=( a75730a  and  a75727a );
 a75732a <=( a75731a  and  a75724a );
 a75736a <=( A167  and  A168 );
 a75737a <=( (not A170)  and  a75736a );
 a75740a <=( A199  and  (not A166) );
 a75743a <=( A201  and  (not A200) );
 a75744a <=( a75743a  and  a75740a );
 a75745a <=( a75744a  and  a75737a );
 a75748a <=( (not A265)  and  A202 );
 a75751a <=( (not A267)  and  A266 );
 a75752a <=( a75751a  and  a75748a );
 a75755a <=( (not A269)  and  (not A268) );
 a75758a <=( A301  and  (not A300) );
 a75759a <=( a75758a  and  a75755a );
 a75760a <=( a75759a  and  a75752a );
 a75764a <=( A167  and  A168 );
 a75765a <=( (not A170)  and  a75764a );
 a75768a <=( A199  and  (not A166) );
 a75771a <=( A201  and  (not A200) );
 a75772a <=( a75771a  and  a75768a );
 a75773a <=( a75772a  and  a75765a );
 a75776a <=( (not A265)  and  A202 );
 a75779a <=( (not A267)  and  A266 );
 a75780a <=( a75779a  and  a75776a );
 a75783a <=( (not A269)  and  (not A268) );
 a75786a <=( A302  and  (not A300) );
 a75787a <=( a75786a  and  a75783a );
 a75788a <=( a75787a  and  a75780a );
 a75792a <=( A167  and  A168 );
 a75793a <=( (not A170)  and  a75792a );
 a75796a <=( A199  and  (not A166) );
 a75799a <=( A201  and  (not A200) );
 a75800a <=( a75799a  and  a75796a );
 a75801a <=( a75800a  and  a75793a );
 a75804a <=( (not A265)  and  A202 );
 a75807a <=( (not A267)  and  A266 );
 a75808a <=( a75807a  and  a75804a );
 a75811a <=( (not A269)  and  (not A268) );
 a75814a <=( A299  and  A298 );
 a75815a <=( a75814a  and  a75811a );
 a75816a <=( a75815a  and  a75808a );
 a75820a <=( A167  and  A168 );
 a75821a <=( (not A170)  and  a75820a );
 a75824a <=( A199  and  (not A166) );
 a75827a <=( A201  and  (not A200) );
 a75828a <=( a75827a  and  a75824a );
 a75829a <=( a75828a  and  a75821a );
 a75832a <=( (not A265)  and  A202 );
 a75835a <=( (not A267)  and  A266 );
 a75836a <=( a75835a  and  a75832a );
 a75839a <=( (not A269)  and  (not A268) );
 a75842a <=( (not A299)  and  (not A298) );
 a75843a <=( a75842a  and  a75839a );
 a75844a <=( a75843a  and  a75836a );
 a75848a <=( A167  and  A168 );
 a75849a <=( (not A170)  and  a75848a );
 a75852a <=( A199  and  (not A166) );
 a75855a <=( A201  and  (not A200) );
 a75856a <=( a75855a  and  a75852a );
 a75857a <=( a75856a  and  a75849a );
 a75860a <=( A265  and  A202 );
 a75863a <=( A267  and  (not A266) );
 a75864a <=( a75863a  and  a75860a );
 a75867a <=( A300  and  A268 );
 a75870a <=( (not A302)  and  (not A301) );
 a75871a <=( a75870a  and  a75867a );
 a75872a <=( a75871a  and  a75864a );
 a75876a <=( A167  and  A168 );
 a75877a <=( (not A170)  and  a75876a );
 a75880a <=( A199  and  (not A166) );
 a75883a <=( A201  and  (not A200) );
 a75884a <=( a75883a  and  a75880a );
 a75885a <=( a75884a  and  a75877a );
 a75888a <=( A265  and  A202 );
 a75891a <=( A267  and  (not A266) );
 a75892a <=( a75891a  and  a75888a );
 a75895a <=( A300  and  A269 );
 a75898a <=( (not A302)  and  (not A301) );
 a75899a <=( a75898a  and  a75895a );
 a75900a <=( a75899a  and  a75892a );
 a75904a <=( A167  and  A168 );
 a75905a <=( (not A170)  and  a75904a );
 a75908a <=( A199  and  (not A166) );
 a75911a <=( A201  and  (not A200) );
 a75912a <=( a75911a  and  a75908a );
 a75913a <=( a75912a  and  a75905a );
 a75916a <=( A265  and  A202 );
 a75919a <=( (not A267)  and  (not A266) );
 a75920a <=( a75919a  and  a75916a );
 a75923a <=( (not A269)  and  (not A268) );
 a75926a <=( A301  and  (not A300) );
 a75927a <=( a75926a  and  a75923a );
 a75928a <=( a75927a  and  a75920a );
 a75932a <=( A167  and  A168 );
 a75933a <=( (not A170)  and  a75932a );
 a75936a <=( A199  and  (not A166) );
 a75939a <=( A201  and  (not A200) );
 a75940a <=( a75939a  and  a75936a );
 a75941a <=( a75940a  and  a75933a );
 a75944a <=( A265  and  A202 );
 a75947a <=( (not A267)  and  (not A266) );
 a75948a <=( a75947a  and  a75944a );
 a75951a <=( (not A269)  and  (not A268) );
 a75954a <=( A302  and  (not A300) );
 a75955a <=( a75954a  and  a75951a );
 a75956a <=( a75955a  and  a75948a );
 a75960a <=( A167  and  A168 );
 a75961a <=( (not A170)  and  a75960a );
 a75964a <=( A199  and  (not A166) );
 a75967a <=( A201  and  (not A200) );
 a75968a <=( a75967a  and  a75964a );
 a75969a <=( a75968a  and  a75961a );
 a75972a <=( A265  and  A202 );
 a75975a <=( (not A267)  and  (not A266) );
 a75976a <=( a75975a  and  a75972a );
 a75979a <=( (not A269)  and  (not A268) );
 a75982a <=( A299  and  A298 );
 a75983a <=( a75982a  and  a75979a );
 a75984a <=( a75983a  and  a75976a );
 a75988a <=( A167  and  A168 );
 a75989a <=( (not A170)  and  a75988a );
 a75992a <=( A199  and  (not A166) );
 a75995a <=( A201  and  (not A200) );
 a75996a <=( a75995a  and  a75992a );
 a75997a <=( a75996a  and  a75989a );
 a76000a <=( A265  and  A202 );
 a76003a <=( (not A267)  and  (not A266) );
 a76004a <=( a76003a  and  a76000a );
 a76007a <=( (not A269)  and  (not A268) );
 a76010a <=( (not A299)  and  (not A298) );
 a76011a <=( a76010a  and  a76007a );
 a76012a <=( a76011a  and  a76004a );
 a76016a <=( A167  and  A168 );
 a76017a <=( (not A170)  and  a76016a );
 a76020a <=( A199  and  (not A166) );
 a76023a <=( A201  and  (not A200) );
 a76024a <=( a76023a  and  a76020a );
 a76025a <=( a76024a  and  a76017a );
 a76028a <=( (not A265)  and  A203 );
 a76031a <=( A267  and  A266 );
 a76032a <=( a76031a  and  a76028a );
 a76035a <=( A300  and  A268 );
 a76038a <=( (not A302)  and  (not A301) );
 a76039a <=( a76038a  and  a76035a );
 a76040a <=( a76039a  and  a76032a );
 a76044a <=( A167  and  A168 );
 a76045a <=( (not A170)  and  a76044a );
 a76048a <=( A199  and  (not A166) );
 a76051a <=( A201  and  (not A200) );
 a76052a <=( a76051a  and  a76048a );
 a76053a <=( a76052a  and  a76045a );
 a76056a <=( (not A265)  and  A203 );
 a76059a <=( A267  and  A266 );
 a76060a <=( a76059a  and  a76056a );
 a76063a <=( A300  and  A269 );
 a76066a <=( (not A302)  and  (not A301) );
 a76067a <=( a76066a  and  a76063a );
 a76068a <=( a76067a  and  a76060a );
 a76072a <=( A167  and  A168 );
 a76073a <=( (not A170)  and  a76072a );
 a76076a <=( A199  and  (not A166) );
 a76079a <=( A201  and  (not A200) );
 a76080a <=( a76079a  and  a76076a );
 a76081a <=( a76080a  and  a76073a );
 a76084a <=( (not A265)  and  A203 );
 a76087a <=( (not A267)  and  A266 );
 a76088a <=( a76087a  and  a76084a );
 a76091a <=( (not A269)  and  (not A268) );
 a76094a <=( A301  and  (not A300) );
 a76095a <=( a76094a  and  a76091a );
 a76096a <=( a76095a  and  a76088a );
 a76100a <=( A167  and  A168 );
 a76101a <=( (not A170)  and  a76100a );
 a76104a <=( A199  and  (not A166) );
 a76107a <=( A201  and  (not A200) );
 a76108a <=( a76107a  and  a76104a );
 a76109a <=( a76108a  and  a76101a );
 a76112a <=( (not A265)  and  A203 );
 a76115a <=( (not A267)  and  A266 );
 a76116a <=( a76115a  and  a76112a );
 a76119a <=( (not A269)  and  (not A268) );
 a76122a <=( A302  and  (not A300) );
 a76123a <=( a76122a  and  a76119a );
 a76124a <=( a76123a  and  a76116a );
 a76128a <=( A167  and  A168 );
 a76129a <=( (not A170)  and  a76128a );
 a76132a <=( A199  and  (not A166) );
 a76135a <=( A201  and  (not A200) );
 a76136a <=( a76135a  and  a76132a );
 a76137a <=( a76136a  and  a76129a );
 a76140a <=( (not A265)  and  A203 );
 a76143a <=( (not A267)  and  A266 );
 a76144a <=( a76143a  and  a76140a );
 a76147a <=( (not A269)  and  (not A268) );
 a76150a <=( A299  and  A298 );
 a76151a <=( a76150a  and  a76147a );
 a76152a <=( a76151a  and  a76144a );
 a76156a <=( A167  and  A168 );
 a76157a <=( (not A170)  and  a76156a );
 a76160a <=( A199  and  (not A166) );
 a76163a <=( A201  and  (not A200) );
 a76164a <=( a76163a  and  a76160a );
 a76165a <=( a76164a  and  a76157a );
 a76168a <=( (not A265)  and  A203 );
 a76171a <=( (not A267)  and  A266 );
 a76172a <=( a76171a  and  a76168a );
 a76175a <=( (not A269)  and  (not A268) );
 a76178a <=( (not A299)  and  (not A298) );
 a76179a <=( a76178a  and  a76175a );
 a76180a <=( a76179a  and  a76172a );
 a76184a <=( A167  and  A168 );
 a76185a <=( (not A170)  and  a76184a );
 a76188a <=( A199  and  (not A166) );
 a76191a <=( A201  and  (not A200) );
 a76192a <=( a76191a  and  a76188a );
 a76193a <=( a76192a  and  a76185a );
 a76196a <=( A265  and  A203 );
 a76199a <=( A267  and  (not A266) );
 a76200a <=( a76199a  and  a76196a );
 a76203a <=( A300  and  A268 );
 a76206a <=( (not A302)  and  (not A301) );
 a76207a <=( a76206a  and  a76203a );
 a76208a <=( a76207a  and  a76200a );
 a76212a <=( A167  and  A168 );
 a76213a <=( (not A170)  and  a76212a );
 a76216a <=( A199  and  (not A166) );
 a76219a <=( A201  and  (not A200) );
 a76220a <=( a76219a  and  a76216a );
 a76221a <=( a76220a  and  a76213a );
 a76224a <=( A265  and  A203 );
 a76227a <=( A267  and  (not A266) );
 a76228a <=( a76227a  and  a76224a );
 a76231a <=( A300  and  A269 );
 a76234a <=( (not A302)  and  (not A301) );
 a76235a <=( a76234a  and  a76231a );
 a76236a <=( a76235a  and  a76228a );
 a76240a <=( A167  and  A168 );
 a76241a <=( (not A170)  and  a76240a );
 a76244a <=( A199  and  (not A166) );
 a76247a <=( A201  and  (not A200) );
 a76248a <=( a76247a  and  a76244a );
 a76249a <=( a76248a  and  a76241a );
 a76252a <=( A265  and  A203 );
 a76255a <=( (not A267)  and  (not A266) );
 a76256a <=( a76255a  and  a76252a );
 a76259a <=( (not A269)  and  (not A268) );
 a76262a <=( A301  and  (not A300) );
 a76263a <=( a76262a  and  a76259a );
 a76264a <=( a76263a  and  a76256a );
 a76268a <=( A167  and  A168 );
 a76269a <=( (not A170)  and  a76268a );
 a76272a <=( A199  and  (not A166) );
 a76275a <=( A201  and  (not A200) );
 a76276a <=( a76275a  and  a76272a );
 a76277a <=( a76276a  and  a76269a );
 a76280a <=( A265  and  A203 );
 a76283a <=( (not A267)  and  (not A266) );
 a76284a <=( a76283a  and  a76280a );
 a76287a <=( (not A269)  and  (not A268) );
 a76290a <=( A302  and  (not A300) );
 a76291a <=( a76290a  and  a76287a );
 a76292a <=( a76291a  and  a76284a );
 a76296a <=( A167  and  A168 );
 a76297a <=( (not A170)  and  a76296a );
 a76300a <=( A199  and  (not A166) );
 a76303a <=( A201  and  (not A200) );
 a76304a <=( a76303a  and  a76300a );
 a76305a <=( a76304a  and  a76297a );
 a76308a <=( A265  and  A203 );
 a76311a <=( (not A267)  and  (not A266) );
 a76312a <=( a76311a  and  a76308a );
 a76315a <=( (not A269)  and  (not A268) );
 a76318a <=( A299  and  A298 );
 a76319a <=( a76318a  and  a76315a );
 a76320a <=( a76319a  and  a76312a );
 a76324a <=( A167  and  A168 );
 a76325a <=( (not A170)  and  a76324a );
 a76328a <=( A199  and  (not A166) );
 a76331a <=( A201  and  (not A200) );
 a76332a <=( a76331a  and  a76328a );
 a76333a <=( a76332a  and  a76325a );
 a76336a <=( A265  and  A203 );
 a76339a <=( (not A267)  and  (not A266) );
 a76340a <=( a76339a  and  a76336a );
 a76343a <=( (not A269)  and  (not A268) );
 a76346a <=( (not A299)  and  (not A298) );
 a76347a <=( a76346a  and  a76343a );
 a76348a <=( a76347a  and  a76340a );
 a76352a <=( A167  and  A168 );
 a76353a <=( (not A170)  and  a76352a );
 a76356a <=( A199  and  (not A166) );
 a76359a <=( (not A201)  and  (not A200) );
 a76360a <=( a76359a  and  a76356a );
 a76361a <=( a76360a  and  a76353a );
 a76364a <=( (not A203)  and  (not A202) );
 a76367a <=( A266  and  (not A265) );
 a76368a <=( a76367a  and  a76364a );
 a76371a <=( A268  and  A267 );
 a76374a <=( A301  and  (not A300) );
 a76375a <=( a76374a  and  a76371a );
 a76376a <=( a76375a  and  a76368a );
 a76380a <=( A167  and  A168 );
 a76381a <=( (not A170)  and  a76380a );
 a76384a <=( A199  and  (not A166) );
 a76387a <=( (not A201)  and  (not A200) );
 a76388a <=( a76387a  and  a76384a );
 a76389a <=( a76388a  and  a76381a );
 a76392a <=( (not A203)  and  (not A202) );
 a76395a <=( A266  and  (not A265) );
 a76396a <=( a76395a  and  a76392a );
 a76399a <=( A268  and  A267 );
 a76402a <=( A302  and  (not A300) );
 a76403a <=( a76402a  and  a76399a );
 a76404a <=( a76403a  and  a76396a );
 a76408a <=( A167  and  A168 );
 a76409a <=( (not A170)  and  a76408a );
 a76412a <=( A199  and  (not A166) );
 a76415a <=( (not A201)  and  (not A200) );
 a76416a <=( a76415a  and  a76412a );
 a76417a <=( a76416a  and  a76409a );
 a76420a <=( (not A203)  and  (not A202) );
 a76423a <=( A266  and  (not A265) );
 a76424a <=( a76423a  and  a76420a );
 a76427a <=( A268  and  A267 );
 a76430a <=( A299  and  A298 );
 a76431a <=( a76430a  and  a76427a );
 a76432a <=( a76431a  and  a76424a );
 a76436a <=( A167  and  A168 );
 a76437a <=( (not A170)  and  a76436a );
 a76440a <=( A199  and  (not A166) );
 a76443a <=( (not A201)  and  (not A200) );
 a76444a <=( a76443a  and  a76440a );
 a76445a <=( a76444a  and  a76437a );
 a76448a <=( (not A203)  and  (not A202) );
 a76451a <=( A266  and  (not A265) );
 a76452a <=( a76451a  and  a76448a );
 a76455a <=( A268  and  A267 );
 a76458a <=( (not A299)  and  (not A298) );
 a76459a <=( a76458a  and  a76455a );
 a76460a <=( a76459a  and  a76452a );
 a76464a <=( A167  and  A168 );
 a76465a <=( (not A170)  and  a76464a );
 a76468a <=( A199  and  (not A166) );
 a76471a <=( (not A201)  and  (not A200) );
 a76472a <=( a76471a  and  a76468a );
 a76473a <=( a76472a  and  a76465a );
 a76476a <=( (not A203)  and  (not A202) );
 a76479a <=( A266  and  (not A265) );
 a76480a <=( a76479a  and  a76476a );
 a76483a <=( A269  and  A267 );
 a76486a <=( A301  and  (not A300) );
 a76487a <=( a76486a  and  a76483a );
 a76488a <=( a76487a  and  a76480a );
 a76492a <=( A167  and  A168 );
 a76493a <=( (not A170)  and  a76492a );
 a76496a <=( A199  and  (not A166) );
 a76499a <=( (not A201)  and  (not A200) );
 a76500a <=( a76499a  and  a76496a );
 a76501a <=( a76500a  and  a76493a );
 a76504a <=( (not A203)  and  (not A202) );
 a76507a <=( A266  and  (not A265) );
 a76508a <=( a76507a  and  a76504a );
 a76511a <=( A269  and  A267 );
 a76514a <=( A302  and  (not A300) );
 a76515a <=( a76514a  and  a76511a );
 a76516a <=( a76515a  and  a76508a );
 a76520a <=( A167  and  A168 );
 a76521a <=( (not A170)  and  a76520a );
 a76524a <=( A199  and  (not A166) );
 a76527a <=( (not A201)  and  (not A200) );
 a76528a <=( a76527a  and  a76524a );
 a76529a <=( a76528a  and  a76521a );
 a76532a <=( (not A203)  and  (not A202) );
 a76535a <=( A266  and  (not A265) );
 a76536a <=( a76535a  and  a76532a );
 a76539a <=( A269  and  A267 );
 a76542a <=( A299  and  A298 );
 a76543a <=( a76542a  and  a76539a );
 a76544a <=( a76543a  and  a76536a );
 a76548a <=( A167  and  A168 );
 a76549a <=( (not A170)  and  a76548a );
 a76552a <=( A199  and  (not A166) );
 a76555a <=( (not A201)  and  (not A200) );
 a76556a <=( a76555a  and  a76552a );
 a76557a <=( a76556a  and  a76549a );
 a76560a <=( (not A203)  and  (not A202) );
 a76563a <=( A266  and  (not A265) );
 a76564a <=( a76563a  and  a76560a );
 a76567a <=( A269  and  A267 );
 a76570a <=( (not A299)  and  (not A298) );
 a76571a <=( a76570a  and  a76567a );
 a76572a <=( a76571a  and  a76564a );
 a76576a <=( A167  and  A168 );
 a76577a <=( (not A170)  and  a76576a );
 a76580a <=( A199  and  (not A166) );
 a76583a <=( (not A201)  and  (not A200) );
 a76584a <=( a76583a  and  a76580a );
 a76585a <=( a76584a  and  a76577a );
 a76588a <=( (not A203)  and  (not A202) );
 a76591a <=( (not A266)  and  A265 );
 a76592a <=( a76591a  and  a76588a );
 a76595a <=( A268  and  A267 );
 a76598a <=( A301  and  (not A300) );
 a76599a <=( a76598a  and  a76595a );
 a76600a <=( a76599a  and  a76592a );
 a76604a <=( A167  and  A168 );
 a76605a <=( (not A170)  and  a76604a );
 a76608a <=( A199  and  (not A166) );
 a76611a <=( (not A201)  and  (not A200) );
 a76612a <=( a76611a  and  a76608a );
 a76613a <=( a76612a  and  a76605a );
 a76616a <=( (not A203)  and  (not A202) );
 a76619a <=( (not A266)  and  A265 );
 a76620a <=( a76619a  and  a76616a );
 a76623a <=( A268  and  A267 );
 a76626a <=( A302  and  (not A300) );
 a76627a <=( a76626a  and  a76623a );
 a76628a <=( a76627a  and  a76620a );
 a76632a <=( A167  and  A168 );
 a76633a <=( (not A170)  and  a76632a );
 a76636a <=( A199  and  (not A166) );
 a76639a <=( (not A201)  and  (not A200) );
 a76640a <=( a76639a  and  a76636a );
 a76641a <=( a76640a  and  a76633a );
 a76644a <=( (not A203)  and  (not A202) );
 a76647a <=( (not A266)  and  A265 );
 a76648a <=( a76647a  and  a76644a );
 a76651a <=( A268  and  A267 );
 a76654a <=( A299  and  A298 );
 a76655a <=( a76654a  and  a76651a );
 a76656a <=( a76655a  and  a76648a );
 a76660a <=( A167  and  A168 );
 a76661a <=( (not A170)  and  a76660a );
 a76664a <=( A199  and  (not A166) );
 a76667a <=( (not A201)  and  (not A200) );
 a76668a <=( a76667a  and  a76664a );
 a76669a <=( a76668a  and  a76661a );
 a76672a <=( (not A203)  and  (not A202) );
 a76675a <=( (not A266)  and  A265 );
 a76676a <=( a76675a  and  a76672a );
 a76679a <=( A268  and  A267 );
 a76682a <=( (not A299)  and  (not A298) );
 a76683a <=( a76682a  and  a76679a );
 a76684a <=( a76683a  and  a76676a );
 a76688a <=( A167  and  A168 );
 a76689a <=( (not A170)  and  a76688a );
 a76692a <=( A199  and  (not A166) );
 a76695a <=( (not A201)  and  (not A200) );
 a76696a <=( a76695a  and  a76692a );
 a76697a <=( a76696a  and  a76689a );
 a76700a <=( (not A203)  and  (not A202) );
 a76703a <=( (not A266)  and  A265 );
 a76704a <=( a76703a  and  a76700a );
 a76707a <=( A269  and  A267 );
 a76710a <=( A301  and  (not A300) );
 a76711a <=( a76710a  and  a76707a );
 a76712a <=( a76711a  and  a76704a );
 a76716a <=( A167  and  A168 );
 a76717a <=( (not A170)  and  a76716a );
 a76720a <=( A199  and  (not A166) );
 a76723a <=( (not A201)  and  (not A200) );
 a76724a <=( a76723a  and  a76720a );
 a76725a <=( a76724a  and  a76717a );
 a76728a <=( (not A203)  and  (not A202) );
 a76731a <=( (not A266)  and  A265 );
 a76732a <=( a76731a  and  a76728a );
 a76735a <=( A269  and  A267 );
 a76738a <=( A302  and  (not A300) );
 a76739a <=( a76738a  and  a76735a );
 a76740a <=( a76739a  and  a76732a );
 a76744a <=( A167  and  A168 );
 a76745a <=( (not A170)  and  a76744a );
 a76748a <=( A199  and  (not A166) );
 a76751a <=( (not A201)  and  (not A200) );
 a76752a <=( a76751a  and  a76748a );
 a76753a <=( a76752a  and  a76745a );
 a76756a <=( (not A203)  and  (not A202) );
 a76759a <=( (not A266)  and  A265 );
 a76760a <=( a76759a  and  a76756a );
 a76763a <=( A269  and  A267 );
 a76766a <=( A299  and  A298 );
 a76767a <=( a76766a  and  a76763a );
 a76768a <=( a76767a  and  a76760a );
 a76772a <=( A167  and  A168 );
 a76773a <=( (not A170)  and  a76772a );
 a76776a <=( A199  and  (not A166) );
 a76779a <=( (not A201)  and  (not A200) );
 a76780a <=( a76779a  and  a76776a );
 a76781a <=( a76780a  and  a76773a );
 a76784a <=( (not A203)  and  (not A202) );
 a76787a <=( (not A266)  and  A265 );
 a76788a <=( a76787a  and  a76784a );
 a76791a <=( A269  and  A267 );
 a76794a <=( (not A299)  and  (not A298) );
 a76795a <=( a76794a  and  a76791a );
 a76796a <=( a76795a  and  a76788a );
 a76800a <=( (not A167)  and  A168 );
 a76801a <=( (not A170)  and  a76800a );
 a76804a <=( A201  and  A166 );
 a76807a <=( (not A203)  and  (not A202) );
 a76808a <=( a76807a  and  a76804a );
 a76809a <=( a76808a  and  a76801a );
 a76812a <=( (not A268)  and  A267 );
 a76815a <=( A298  and  (not A269) );
 a76816a <=( a76815a  and  a76812a );
 a76819a <=( (not A300)  and  (not A299) );
 a76822a <=( (not A302)  and  (not A301) );
 a76823a <=( a76822a  and  a76819a );
 a76824a <=( a76823a  and  a76816a );
 a76828a <=( (not A167)  and  A168 );
 a76829a <=( (not A170)  and  a76828a );
 a76832a <=( A201  and  A166 );
 a76835a <=( (not A203)  and  (not A202) );
 a76836a <=( a76835a  and  a76832a );
 a76837a <=( a76836a  and  a76829a );
 a76840a <=( (not A268)  and  A267 );
 a76843a <=( (not A298)  and  (not A269) );
 a76844a <=( a76843a  and  a76840a );
 a76847a <=( (not A300)  and  A299 );
 a76850a <=( (not A302)  and  (not A301) );
 a76851a <=( a76850a  and  a76847a );
 a76852a <=( a76851a  and  a76844a );
 a76856a <=( (not A167)  and  A168 );
 a76857a <=( (not A170)  and  a76856a );
 a76860a <=( (not A199)  and  A166 );
 a76863a <=( A201  and  A200 );
 a76864a <=( a76863a  and  a76860a );
 a76865a <=( a76864a  and  a76857a );
 a76868a <=( (not A265)  and  A202 );
 a76871a <=( A267  and  A266 );
 a76872a <=( a76871a  and  a76868a );
 a76875a <=( A300  and  A268 );
 a76878a <=( (not A302)  and  (not A301) );
 a76879a <=( a76878a  and  a76875a );
 a76880a <=( a76879a  and  a76872a );
 a76884a <=( (not A167)  and  A168 );
 a76885a <=( (not A170)  and  a76884a );
 a76888a <=( (not A199)  and  A166 );
 a76891a <=( A201  and  A200 );
 a76892a <=( a76891a  and  a76888a );
 a76893a <=( a76892a  and  a76885a );
 a76896a <=( (not A265)  and  A202 );
 a76899a <=( A267  and  A266 );
 a76900a <=( a76899a  and  a76896a );
 a76903a <=( A300  and  A269 );
 a76906a <=( (not A302)  and  (not A301) );
 a76907a <=( a76906a  and  a76903a );
 a76908a <=( a76907a  and  a76900a );
 a76912a <=( (not A167)  and  A168 );
 a76913a <=( (not A170)  and  a76912a );
 a76916a <=( (not A199)  and  A166 );
 a76919a <=( A201  and  A200 );
 a76920a <=( a76919a  and  a76916a );
 a76921a <=( a76920a  and  a76913a );
 a76924a <=( (not A265)  and  A202 );
 a76927a <=( (not A267)  and  A266 );
 a76928a <=( a76927a  and  a76924a );
 a76931a <=( (not A269)  and  (not A268) );
 a76934a <=( A301  and  (not A300) );
 a76935a <=( a76934a  and  a76931a );
 a76936a <=( a76935a  and  a76928a );
 a76940a <=( (not A167)  and  A168 );
 a76941a <=( (not A170)  and  a76940a );
 a76944a <=( (not A199)  and  A166 );
 a76947a <=( A201  and  A200 );
 a76948a <=( a76947a  and  a76944a );
 a76949a <=( a76948a  and  a76941a );
 a76952a <=( (not A265)  and  A202 );
 a76955a <=( (not A267)  and  A266 );
 a76956a <=( a76955a  and  a76952a );
 a76959a <=( (not A269)  and  (not A268) );
 a76962a <=( A302  and  (not A300) );
 a76963a <=( a76962a  and  a76959a );
 a76964a <=( a76963a  and  a76956a );
 a76968a <=( (not A167)  and  A168 );
 a76969a <=( (not A170)  and  a76968a );
 a76972a <=( (not A199)  and  A166 );
 a76975a <=( A201  and  A200 );
 a76976a <=( a76975a  and  a76972a );
 a76977a <=( a76976a  and  a76969a );
 a76980a <=( (not A265)  and  A202 );
 a76983a <=( (not A267)  and  A266 );
 a76984a <=( a76983a  and  a76980a );
 a76987a <=( (not A269)  and  (not A268) );
 a76990a <=( A299  and  A298 );
 a76991a <=( a76990a  and  a76987a );
 a76992a <=( a76991a  and  a76984a );
 a76996a <=( (not A167)  and  A168 );
 a76997a <=( (not A170)  and  a76996a );
 a77000a <=( (not A199)  and  A166 );
 a77003a <=( A201  and  A200 );
 a77004a <=( a77003a  and  a77000a );
 a77005a <=( a77004a  and  a76997a );
 a77008a <=( (not A265)  and  A202 );
 a77011a <=( (not A267)  and  A266 );
 a77012a <=( a77011a  and  a77008a );
 a77015a <=( (not A269)  and  (not A268) );
 a77018a <=( (not A299)  and  (not A298) );
 a77019a <=( a77018a  and  a77015a );
 a77020a <=( a77019a  and  a77012a );
 a77024a <=( (not A167)  and  A168 );
 a77025a <=( (not A170)  and  a77024a );
 a77028a <=( (not A199)  and  A166 );
 a77031a <=( A201  and  A200 );
 a77032a <=( a77031a  and  a77028a );
 a77033a <=( a77032a  and  a77025a );
 a77036a <=( A265  and  A202 );
 a77039a <=( A267  and  (not A266) );
 a77040a <=( a77039a  and  a77036a );
 a77043a <=( A300  and  A268 );
 a77046a <=( (not A302)  and  (not A301) );
 a77047a <=( a77046a  and  a77043a );
 a77048a <=( a77047a  and  a77040a );
 a77052a <=( (not A167)  and  A168 );
 a77053a <=( (not A170)  and  a77052a );
 a77056a <=( (not A199)  and  A166 );
 a77059a <=( A201  and  A200 );
 a77060a <=( a77059a  and  a77056a );
 a77061a <=( a77060a  and  a77053a );
 a77064a <=( A265  and  A202 );
 a77067a <=( A267  and  (not A266) );
 a77068a <=( a77067a  and  a77064a );
 a77071a <=( A300  and  A269 );
 a77074a <=( (not A302)  and  (not A301) );
 a77075a <=( a77074a  and  a77071a );
 a77076a <=( a77075a  and  a77068a );
 a77080a <=( (not A167)  and  A168 );
 a77081a <=( (not A170)  and  a77080a );
 a77084a <=( (not A199)  and  A166 );
 a77087a <=( A201  and  A200 );
 a77088a <=( a77087a  and  a77084a );
 a77089a <=( a77088a  and  a77081a );
 a77092a <=( A265  and  A202 );
 a77095a <=( (not A267)  and  (not A266) );
 a77096a <=( a77095a  and  a77092a );
 a77099a <=( (not A269)  and  (not A268) );
 a77102a <=( A301  and  (not A300) );
 a77103a <=( a77102a  and  a77099a );
 a77104a <=( a77103a  and  a77096a );
 a77108a <=( (not A167)  and  A168 );
 a77109a <=( (not A170)  and  a77108a );
 a77112a <=( (not A199)  and  A166 );
 a77115a <=( A201  and  A200 );
 a77116a <=( a77115a  and  a77112a );
 a77117a <=( a77116a  and  a77109a );
 a77120a <=( A265  and  A202 );
 a77123a <=( (not A267)  and  (not A266) );
 a77124a <=( a77123a  and  a77120a );
 a77127a <=( (not A269)  and  (not A268) );
 a77130a <=( A302  and  (not A300) );
 a77131a <=( a77130a  and  a77127a );
 a77132a <=( a77131a  and  a77124a );
 a77136a <=( (not A167)  and  A168 );
 a77137a <=( (not A170)  and  a77136a );
 a77140a <=( (not A199)  and  A166 );
 a77143a <=( A201  and  A200 );
 a77144a <=( a77143a  and  a77140a );
 a77145a <=( a77144a  and  a77137a );
 a77148a <=( A265  and  A202 );
 a77151a <=( (not A267)  and  (not A266) );
 a77152a <=( a77151a  and  a77148a );
 a77155a <=( (not A269)  and  (not A268) );
 a77158a <=( A299  and  A298 );
 a77159a <=( a77158a  and  a77155a );
 a77160a <=( a77159a  and  a77152a );
 a77164a <=( (not A167)  and  A168 );
 a77165a <=( (not A170)  and  a77164a );
 a77168a <=( (not A199)  and  A166 );
 a77171a <=( A201  and  A200 );
 a77172a <=( a77171a  and  a77168a );
 a77173a <=( a77172a  and  a77165a );
 a77176a <=( A265  and  A202 );
 a77179a <=( (not A267)  and  (not A266) );
 a77180a <=( a77179a  and  a77176a );
 a77183a <=( (not A269)  and  (not A268) );
 a77186a <=( (not A299)  and  (not A298) );
 a77187a <=( a77186a  and  a77183a );
 a77188a <=( a77187a  and  a77180a );
 a77192a <=( (not A167)  and  A168 );
 a77193a <=( (not A170)  and  a77192a );
 a77196a <=( (not A199)  and  A166 );
 a77199a <=( A201  and  A200 );
 a77200a <=( a77199a  and  a77196a );
 a77201a <=( a77200a  and  a77193a );
 a77204a <=( (not A265)  and  A203 );
 a77207a <=( A267  and  A266 );
 a77208a <=( a77207a  and  a77204a );
 a77211a <=( A300  and  A268 );
 a77214a <=( (not A302)  and  (not A301) );
 a77215a <=( a77214a  and  a77211a );
 a77216a <=( a77215a  and  a77208a );
 a77220a <=( (not A167)  and  A168 );
 a77221a <=( (not A170)  and  a77220a );
 a77224a <=( (not A199)  and  A166 );
 a77227a <=( A201  and  A200 );
 a77228a <=( a77227a  and  a77224a );
 a77229a <=( a77228a  and  a77221a );
 a77232a <=( (not A265)  and  A203 );
 a77235a <=( A267  and  A266 );
 a77236a <=( a77235a  and  a77232a );
 a77239a <=( A300  and  A269 );
 a77242a <=( (not A302)  and  (not A301) );
 a77243a <=( a77242a  and  a77239a );
 a77244a <=( a77243a  and  a77236a );
 a77248a <=( (not A167)  and  A168 );
 a77249a <=( (not A170)  and  a77248a );
 a77252a <=( (not A199)  and  A166 );
 a77255a <=( A201  and  A200 );
 a77256a <=( a77255a  and  a77252a );
 a77257a <=( a77256a  and  a77249a );
 a77260a <=( (not A265)  and  A203 );
 a77263a <=( (not A267)  and  A266 );
 a77264a <=( a77263a  and  a77260a );
 a77267a <=( (not A269)  and  (not A268) );
 a77270a <=( A301  and  (not A300) );
 a77271a <=( a77270a  and  a77267a );
 a77272a <=( a77271a  and  a77264a );
 a77276a <=( (not A167)  and  A168 );
 a77277a <=( (not A170)  and  a77276a );
 a77280a <=( (not A199)  and  A166 );
 a77283a <=( A201  and  A200 );
 a77284a <=( a77283a  and  a77280a );
 a77285a <=( a77284a  and  a77277a );
 a77288a <=( (not A265)  and  A203 );
 a77291a <=( (not A267)  and  A266 );
 a77292a <=( a77291a  and  a77288a );
 a77295a <=( (not A269)  and  (not A268) );
 a77298a <=( A302  and  (not A300) );
 a77299a <=( a77298a  and  a77295a );
 a77300a <=( a77299a  and  a77292a );
 a77304a <=( (not A167)  and  A168 );
 a77305a <=( (not A170)  and  a77304a );
 a77308a <=( (not A199)  and  A166 );
 a77311a <=( A201  and  A200 );
 a77312a <=( a77311a  and  a77308a );
 a77313a <=( a77312a  and  a77305a );
 a77316a <=( (not A265)  and  A203 );
 a77319a <=( (not A267)  and  A266 );
 a77320a <=( a77319a  and  a77316a );
 a77323a <=( (not A269)  and  (not A268) );
 a77326a <=( A299  and  A298 );
 a77327a <=( a77326a  and  a77323a );
 a77328a <=( a77327a  and  a77320a );
 a77332a <=( (not A167)  and  A168 );
 a77333a <=( (not A170)  and  a77332a );
 a77336a <=( (not A199)  and  A166 );
 a77339a <=( A201  and  A200 );
 a77340a <=( a77339a  and  a77336a );
 a77341a <=( a77340a  and  a77333a );
 a77344a <=( (not A265)  and  A203 );
 a77347a <=( (not A267)  and  A266 );
 a77348a <=( a77347a  and  a77344a );
 a77351a <=( (not A269)  and  (not A268) );
 a77354a <=( (not A299)  and  (not A298) );
 a77355a <=( a77354a  and  a77351a );
 a77356a <=( a77355a  and  a77348a );
 a77360a <=( (not A167)  and  A168 );
 a77361a <=( (not A170)  and  a77360a );
 a77364a <=( (not A199)  and  A166 );
 a77367a <=( A201  and  A200 );
 a77368a <=( a77367a  and  a77364a );
 a77369a <=( a77368a  and  a77361a );
 a77372a <=( A265  and  A203 );
 a77375a <=( A267  and  (not A266) );
 a77376a <=( a77375a  and  a77372a );
 a77379a <=( A300  and  A268 );
 a77382a <=( (not A302)  and  (not A301) );
 a77383a <=( a77382a  and  a77379a );
 a77384a <=( a77383a  and  a77376a );
 a77388a <=( (not A167)  and  A168 );
 a77389a <=( (not A170)  and  a77388a );
 a77392a <=( (not A199)  and  A166 );
 a77395a <=( A201  and  A200 );
 a77396a <=( a77395a  and  a77392a );
 a77397a <=( a77396a  and  a77389a );
 a77400a <=( A265  and  A203 );
 a77403a <=( A267  and  (not A266) );
 a77404a <=( a77403a  and  a77400a );
 a77407a <=( A300  and  A269 );
 a77410a <=( (not A302)  and  (not A301) );
 a77411a <=( a77410a  and  a77407a );
 a77412a <=( a77411a  and  a77404a );
 a77416a <=( (not A167)  and  A168 );
 a77417a <=( (not A170)  and  a77416a );
 a77420a <=( (not A199)  and  A166 );
 a77423a <=( A201  and  A200 );
 a77424a <=( a77423a  and  a77420a );
 a77425a <=( a77424a  and  a77417a );
 a77428a <=( A265  and  A203 );
 a77431a <=( (not A267)  and  (not A266) );
 a77432a <=( a77431a  and  a77428a );
 a77435a <=( (not A269)  and  (not A268) );
 a77438a <=( A301  and  (not A300) );
 a77439a <=( a77438a  and  a77435a );
 a77440a <=( a77439a  and  a77432a );
 a77444a <=( (not A167)  and  A168 );
 a77445a <=( (not A170)  and  a77444a );
 a77448a <=( (not A199)  and  A166 );
 a77451a <=( A201  and  A200 );
 a77452a <=( a77451a  and  a77448a );
 a77453a <=( a77452a  and  a77445a );
 a77456a <=( A265  and  A203 );
 a77459a <=( (not A267)  and  (not A266) );
 a77460a <=( a77459a  and  a77456a );
 a77463a <=( (not A269)  and  (not A268) );
 a77466a <=( A302  and  (not A300) );
 a77467a <=( a77466a  and  a77463a );
 a77468a <=( a77467a  and  a77460a );
 a77472a <=( (not A167)  and  A168 );
 a77473a <=( (not A170)  and  a77472a );
 a77476a <=( (not A199)  and  A166 );
 a77479a <=( A201  and  A200 );
 a77480a <=( a77479a  and  a77476a );
 a77481a <=( a77480a  and  a77473a );
 a77484a <=( A265  and  A203 );
 a77487a <=( (not A267)  and  (not A266) );
 a77488a <=( a77487a  and  a77484a );
 a77491a <=( (not A269)  and  (not A268) );
 a77494a <=( A299  and  A298 );
 a77495a <=( a77494a  and  a77491a );
 a77496a <=( a77495a  and  a77488a );
 a77500a <=( (not A167)  and  A168 );
 a77501a <=( (not A170)  and  a77500a );
 a77504a <=( (not A199)  and  A166 );
 a77507a <=( A201  and  A200 );
 a77508a <=( a77507a  and  a77504a );
 a77509a <=( a77508a  and  a77501a );
 a77512a <=( A265  and  A203 );
 a77515a <=( (not A267)  and  (not A266) );
 a77516a <=( a77515a  and  a77512a );
 a77519a <=( (not A269)  and  (not A268) );
 a77522a <=( (not A299)  and  (not A298) );
 a77523a <=( a77522a  and  a77519a );
 a77524a <=( a77523a  and  a77516a );
 a77528a <=( (not A167)  and  A168 );
 a77529a <=( (not A170)  and  a77528a );
 a77532a <=( (not A199)  and  A166 );
 a77535a <=( (not A201)  and  A200 );
 a77536a <=( a77535a  and  a77532a );
 a77537a <=( a77536a  and  a77529a );
 a77540a <=( (not A203)  and  (not A202) );
 a77543a <=( A266  and  (not A265) );
 a77544a <=( a77543a  and  a77540a );
 a77547a <=( A268  and  A267 );
 a77550a <=( A301  and  (not A300) );
 a77551a <=( a77550a  and  a77547a );
 a77552a <=( a77551a  and  a77544a );
 a77556a <=( (not A167)  and  A168 );
 a77557a <=( (not A170)  and  a77556a );
 a77560a <=( (not A199)  and  A166 );
 a77563a <=( (not A201)  and  A200 );
 a77564a <=( a77563a  and  a77560a );
 a77565a <=( a77564a  and  a77557a );
 a77568a <=( (not A203)  and  (not A202) );
 a77571a <=( A266  and  (not A265) );
 a77572a <=( a77571a  and  a77568a );
 a77575a <=( A268  and  A267 );
 a77578a <=( A302  and  (not A300) );
 a77579a <=( a77578a  and  a77575a );
 a77580a <=( a77579a  and  a77572a );
 a77584a <=( (not A167)  and  A168 );
 a77585a <=( (not A170)  and  a77584a );
 a77588a <=( (not A199)  and  A166 );
 a77591a <=( (not A201)  and  A200 );
 a77592a <=( a77591a  and  a77588a );
 a77593a <=( a77592a  and  a77585a );
 a77596a <=( (not A203)  and  (not A202) );
 a77599a <=( A266  and  (not A265) );
 a77600a <=( a77599a  and  a77596a );
 a77603a <=( A268  and  A267 );
 a77606a <=( A299  and  A298 );
 a77607a <=( a77606a  and  a77603a );
 a77608a <=( a77607a  and  a77600a );
 a77612a <=( (not A167)  and  A168 );
 a77613a <=( (not A170)  and  a77612a );
 a77616a <=( (not A199)  and  A166 );
 a77619a <=( (not A201)  and  A200 );
 a77620a <=( a77619a  and  a77616a );
 a77621a <=( a77620a  and  a77613a );
 a77624a <=( (not A203)  and  (not A202) );
 a77627a <=( A266  and  (not A265) );
 a77628a <=( a77627a  and  a77624a );
 a77631a <=( A268  and  A267 );
 a77634a <=( (not A299)  and  (not A298) );
 a77635a <=( a77634a  and  a77631a );
 a77636a <=( a77635a  and  a77628a );
 a77640a <=( (not A167)  and  A168 );
 a77641a <=( (not A170)  and  a77640a );
 a77644a <=( (not A199)  and  A166 );
 a77647a <=( (not A201)  and  A200 );
 a77648a <=( a77647a  and  a77644a );
 a77649a <=( a77648a  and  a77641a );
 a77652a <=( (not A203)  and  (not A202) );
 a77655a <=( A266  and  (not A265) );
 a77656a <=( a77655a  and  a77652a );
 a77659a <=( A269  and  A267 );
 a77662a <=( A301  and  (not A300) );
 a77663a <=( a77662a  and  a77659a );
 a77664a <=( a77663a  and  a77656a );
 a77668a <=( (not A167)  and  A168 );
 a77669a <=( (not A170)  and  a77668a );
 a77672a <=( (not A199)  and  A166 );
 a77675a <=( (not A201)  and  A200 );
 a77676a <=( a77675a  and  a77672a );
 a77677a <=( a77676a  and  a77669a );
 a77680a <=( (not A203)  and  (not A202) );
 a77683a <=( A266  and  (not A265) );
 a77684a <=( a77683a  and  a77680a );
 a77687a <=( A269  and  A267 );
 a77690a <=( A302  and  (not A300) );
 a77691a <=( a77690a  and  a77687a );
 a77692a <=( a77691a  and  a77684a );
 a77696a <=( (not A167)  and  A168 );
 a77697a <=( (not A170)  and  a77696a );
 a77700a <=( (not A199)  and  A166 );
 a77703a <=( (not A201)  and  A200 );
 a77704a <=( a77703a  and  a77700a );
 a77705a <=( a77704a  and  a77697a );
 a77708a <=( (not A203)  and  (not A202) );
 a77711a <=( A266  and  (not A265) );
 a77712a <=( a77711a  and  a77708a );
 a77715a <=( A269  and  A267 );
 a77718a <=( A299  and  A298 );
 a77719a <=( a77718a  and  a77715a );
 a77720a <=( a77719a  and  a77712a );
 a77724a <=( (not A167)  and  A168 );
 a77725a <=( (not A170)  and  a77724a );
 a77728a <=( (not A199)  and  A166 );
 a77731a <=( (not A201)  and  A200 );
 a77732a <=( a77731a  and  a77728a );
 a77733a <=( a77732a  and  a77725a );
 a77736a <=( (not A203)  and  (not A202) );
 a77739a <=( A266  and  (not A265) );
 a77740a <=( a77739a  and  a77736a );
 a77743a <=( A269  and  A267 );
 a77746a <=( (not A299)  and  (not A298) );
 a77747a <=( a77746a  and  a77743a );
 a77748a <=( a77747a  and  a77740a );
 a77752a <=( (not A167)  and  A168 );
 a77753a <=( (not A170)  and  a77752a );
 a77756a <=( (not A199)  and  A166 );
 a77759a <=( (not A201)  and  A200 );
 a77760a <=( a77759a  and  a77756a );
 a77761a <=( a77760a  and  a77753a );
 a77764a <=( (not A203)  and  (not A202) );
 a77767a <=( (not A266)  and  A265 );
 a77768a <=( a77767a  and  a77764a );
 a77771a <=( A268  and  A267 );
 a77774a <=( A301  and  (not A300) );
 a77775a <=( a77774a  and  a77771a );
 a77776a <=( a77775a  and  a77768a );
 a77780a <=( (not A167)  and  A168 );
 a77781a <=( (not A170)  and  a77780a );
 a77784a <=( (not A199)  and  A166 );
 a77787a <=( (not A201)  and  A200 );
 a77788a <=( a77787a  and  a77784a );
 a77789a <=( a77788a  and  a77781a );
 a77792a <=( (not A203)  and  (not A202) );
 a77795a <=( (not A266)  and  A265 );
 a77796a <=( a77795a  and  a77792a );
 a77799a <=( A268  and  A267 );
 a77802a <=( A302  and  (not A300) );
 a77803a <=( a77802a  and  a77799a );
 a77804a <=( a77803a  and  a77796a );
 a77808a <=( (not A167)  and  A168 );
 a77809a <=( (not A170)  and  a77808a );
 a77812a <=( (not A199)  and  A166 );
 a77815a <=( (not A201)  and  A200 );
 a77816a <=( a77815a  and  a77812a );
 a77817a <=( a77816a  and  a77809a );
 a77820a <=( (not A203)  and  (not A202) );
 a77823a <=( (not A266)  and  A265 );
 a77824a <=( a77823a  and  a77820a );
 a77827a <=( A268  and  A267 );
 a77830a <=( A299  and  A298 );
 a77831a <=( a77830a  and  a77827a );
 a77832a <=( a77831a  and  a77824a );
 a77836a <=( (not A167)  and  A168 );
 a77837a <=( (not A170)  and  a77836a );
 a77840a <=( (not A199)  and  A166 );
 a77843a <=( (not A201)  and  A200 );
 a77844a <=( a77843a  and  a77840a );
 a77845a <=( a77844a  and  a77837a );
 a77848a <=( (not A203)  and  (not A202) );
 a77851a <=( (not A266)  and  A265 );
 a77852a <=( a77851a  and  a77848a );
 a77855a <=( A268  and  A267 );
 a77858a <=( (not A299)  and  (not A298) );
 a77859a <=( a77858a  and  a77855a );
 a77860a <=( a77859a  and  a77852a );
 a77864a <=( (not A167)  and  A168 );
 a77865a <=( (not A170)  and  a77864a );
 a77868a <=( (not A199)  and  A166 );
 a77871a <=( (not A201)  and  A200 );
 a77872a <=( a77871a  and  a77868a );
 a77873a <=( a77872a  and  a77865a );
 a77876a <=( (not A203)  and  (not A202) );
 a77879a <=( (not A266)  and  A265 );
 a77880a <=( a77879a  and  a77876a );
 a77883a <=( A269  and  A267 );
 a77886a <=( A301  and  (not A300) );
 a77887a <=( a77886a  and  a77883a );
 a77888a <=( a77887a  and  a77880a );
 a77892a <=( (not A167)  and  A168 );
 a77893a <=( (not A170)  and  a77892a );
 a77896a <=( (not A199)  and  A166 );
 a77899a <=( (not A201)  and  A200 );
 a77900a <=( a77899a  and  a77896a );
 a77901a <=( a77900a  and  a77893a );
 a77904a <=( (not A203)  and  (not A202) );
 a77907a <=( (not A266)  and  A265 );
 a77908a <=( a77907a  and  a77904a );
 a77911a <=( A269  and  A267 );
 a77914a <=( A302  and  (not A300) );
 a77915a <=( a77914a  and  a77911a );
 a77916a <=( a77915a  and  a77908a );
 a77920a <=( (not A167)  and  A168 );
 a77921a <=( (not A170)  and  a77920a );
 a77924a <=( (not A199)  and  A166 );
 a77927a <=( (not A201)  and  A200 );
 a77928a <=( a77927a  and  a77924a );
 a77929a <=( a77928a  and  a77921a );
 a77932a <=( (not A203)  and  (not A202) );
 a77935a <=( (not A266)  and  A265 );
 a77936a <=( a77935a  and  a77932a );
 a77939a <=( A269  and  A267 );
 a77942a <=( A299  and  A298 );
 a77943a <=( a77942a  and  a77939a );
 a77944a <=( a77943a  and  a77936a );
 a77948a <=( (not A167)  and  A168 );
 a77949a <=( (not A170)  and  a77948a );
 a77952a <=( (not A199)  and  A166 );
 a77955a <=( (not A201)  and  A200 );
 a77956a <=( a77955a  and  a77952a );
 a77957a <=( a77956a  and  a77949a );
 a77960a <=( (not A203)  and  (not A202) );
 a77963a <=( (not A266)  and  A265 );
 a77964a <=( a77963a  and  a77960a );
 a77967a <=( A269  and  A267 );
 a77970a <=( (not A299)  and  (not A298) );
 a77971a <=( a77970a  and  a77967a );
 a77972a <=( a77971a  and  a77964a );
 a77976a <=( (not A167)  and  A168 );
 a77977a <=( (not A170)  and  a77976a );
 a77980a <=( A199  and  A166 );
 a77983a <=( A201  and  (not A200) );
 a77984a <=( a77983a  and  a77980a );
 a77985a <=( a77984a  and  a77977a );
 a77988a <=( (not A265)  and  A202 );
 a77991a <=( A267  and  A266 );
 a77992a <=( a77991a  and  a77988a );
 a77995a <=( A300  and  A268 );
 a77998a <=( (not A302)  and  (not A301) );
 a77999a <=( a77998a  and  a77995a );
 a78000a <=( a77999a  and  a77992a );
 a78004a <=( (not A167)  and  A168 );
 a78005a <=( (not A170)  and  a78004a );
 a78008a <=( A199  and  A166 );
 a78011a <=( A201  and  (not A200) );
 a78012a <=( a78011a  and  a78008a );
 a78013a <=( a78012a  and  a78005a );
 a78016a <=( (not A265)  and  A202 );
 a78019a <=( A267  and  A266 );
 a78020a <=( a78019a  and  a78016a );
 a78023a <=( A300  and  A269 );
 a78026a <=( (not A302)  and  (not A301) );
 a78027a <=( a78026a  and  a78023a );
 a78028a <=( a78027a  and  a78020a );
 a78032a <=( (not A167)  and  A168 );
 a78033a <=( (not A170)  and  a78032a );
 a78036a <=( A199  and  A166 );
 a78039a <=( A201  and  (not A200) );
 a78040a <=( a78039a  and  a78036a );
 a78041a <=( a78040a  and  a78033a );
 a78044a <=( (not A265)  and  A202 );
 a78047a <=( (not A267)  and  A266 );
 a78048a <=( a78047a  and  a78044a );
 a78051a <=( (not A269)  and  (not A268) );
 a78054a <=( A301  and  (not A300) );
 a78055a <=( a78054a  and  a78051a );
 a78056a <=( a78055a  and  a78048a );
 a78060a <=( (not A167)  and  A168 );
 a78061a <=( (not A170)  and  a78060a );
 a78064a <=( A199  and  A166 );
 a78067a <=( A201  and  (not A200) );
 a78068a <=( a78067a  and  a78064a );
 a78069a <=( a78068a  and  a78061a );
 a78072a <=( (not A265)  and  A202 );
 a78075a <=( (not A267)  and  A266 );
 a78076a <=( a78075a  and  a78072a );
 a78079a <=( (not A269)  and  (not A268) );
 a78082a <=( A302  and  (not A300) );
 a78083a <=( a78082a  and  a78079a );
 a78084a <=( a78083a  and  a78076a );
 a78088a <=( (not A167)  and  A168 );
 a78089a <=( (not A170)  and  a78088a );
 a78092a <=( A199  and  A166 );
 a78095a <=( A201  and  (not A200) );
 a78096a <=( a78095a  and  a78092a );
 a78097a <=( a78096a  and  a78089a );
 a78100a <=( (not A265)  and  A202 );
 a78103a <=( (not A267)  and  A266 );
 a78104a <=( a78103a  and  a78100a );
 a78107a <=( (not A269)  and  (not A268) );
 a78110a <=( A299  and  A298 );
 a78111a <=( a78110a  and  a78107a );
 a78112a <=( a78111a  and  a78104a );
 a78116a <=( (not A167)  and  A168 );
 a78117a <=( (not A170)  and  a78116a );
 a78120a <=( A199  and  A166 );
 a78123a <=( A201  and  (not A200) );
 a78124a <=( a78123a  and  a78120a );
 a78125a <=( a78124a  and  a78117a );
 a78128a <=( (not A265)  and  A202 );
 a78131a <=( (not A267)  and  A266 );
 a78132a <=( a78131a  and  a78128a );
 a78135a <=( (not A269)  and  (not A268) );
 a78138a <=( (not A299)  and  (not A298) );
 a78139a <=( a78138a  and  a78135a );
 a78140a <=( a78139a  and  a78132a );
 a78144a <=( (not A167)  and  A168 );
 a78145a <=( (not A170)  and  a78144a );
 a78148a <=( A199  and  A166 );
 a78151a <=( A201  and  (not A200) );
 a78152a <=( a78151a  and  a78148a );
 a78153a <=( a78152a  and  a78145a );
 a78156a <=( A265  and  A202 );
 a78159a <=( A267  and  (not A266) );
 a78160a <=( a78159a  and  a78156a );
 a78163a <=( A300  and  A268 );
 a78166a <=( (not A302)  and  (not A301) );
 a78167a <=( a78166a  and  a78163a );
 a78168a <=( a78167a  and  a78160a );
 a78172a <=( (not A167)  and  A168 );
 a78173a <=( (not A170)  and  a78172a );
 a78176a <=( A199  and  A166 );
 a78179a <=( A201  and  (not A200) );
 a78180a <=( a78179a  and  a78176a );
 a78181a <=( a78180a  and  a78173a );
 a78184a <=( A265  and  A202 );
 a78187a <=( A267  and  (not A266) );
 a78188a <=( a78187a  and  a78184a );
 a78191a <=( A300  and  A269 );
 a78194a <=( (not A302)  and  (not A301) );
 a78195a <=( a78194a  and  a78191a );
 a78196a <=( a78195a  and  a78188a );
 a78200a <=( (not A167)  and  A168 );
 a78201a <=( (not A170)  and  a78200a );
 a78204a <=( A199  and  A166 );
 a78207a <=( A201  and  (not A200) );
 a78208a <=( a78207a  and  a78204a );
 a78209a <=( a78208a  and  a78201a );
 a78212a <=( A265  and  A202 );
 a78215a <=( (not A267)  and  (not A266) );
 a78216a <=( a78215a  and  a78212a );
 a78219a <=( (not A269)  and  (not A268) );
 a78222a <=( A301  and  (not A300) );
 a78223a <=( a78222a  and  a78219a );
 a78224a <=( a78223a  and  a78216a );
 a78228a <=( (not A167)  and  A168 );
 a78229a <=( (not A170)  and  a78228a );
 a78232a <=( A199  and  A166 );
 a78235a <=( A201  and  (not A200) );
 a78236a <=( a78235a  and  a78232a );
 a78237a <=( a78236a  and  a78229a );
 a78240a <=( A265  and  A202 );
 a78243a <=( (not A267)  and  (not A266) );
 a78244a <=( a78243a  and  a78240a );
 a78247a <=( (not A269)  and  (not A268) );
 a78250a <=( A302  and  (not A300) );
 a78251a <=( a78250a  and  a78247a );
 a78252a <=( a78251a  and  a78244a );
 a78256a <=( (not A167)  and  A168 );
 a78257a <=( (not A170)  and  a78256a );
 a78260a <=( A199  and  A166 );
 a78263a <=( A201  and  (not A200) );
 a78264a <=( a78263a  and  a78260a );
 a78265a <=( a78264a  and  a78257a );
 a78268a <=( A265  and  A202 );
 a78271a <=( (not A267)  and  (not A266) );
 a78272a <=( a78271a  and  a78268a );
 a78275a <=( (not A269)  and  (not A268) );
 a78278a <=( A299  and  A298 );
 a78279a <=( a78278a  and  a78275a );
 a78280a <=( a78279a  and  a78272a );
 a78284a <=( (not A167)  and  A168 );
 a78285a <=( (not A170)  and  a78284a );
 a78288a <=( A199  and  A166 );
 a78291a <=( A201  and  (not A200) );
 a78292a <=( a78291a  and  a78288a );
 a78293a <=( a78292a  and  a78285a );
 a78296a <=( A265  and  A202 );
 a78299a <=( (not A267)  and  (not A266) );
 a78300a <=( a78299a  and  a78296a );
 a78303a <=( (not A269)  and  (not A268) );
 a78306a <=( (not A299)  and  (not A298) );
 a78307a <=( a78306a  and  a78303a );
 a78308a <=( a78307a  and  a78300a );
 a78312a <=( (not A167)  and  A168 );
 a78313a <=( (not A170)  and  a78312a );
 a78316a <=( A199  and  A166 );
 a78319a <=( A201  and  (not A200) );
 a78320a <=( a78319a  and  a78316a );
 a78321a <=( a78320a  and  a78313a );
 a78324a <=( (not A265)  and  A203 );
 a78327a <=( A267  and  A266 );
 a78328a <=( a78327a  and  a78324a );
 a78331a <=( A300  and  A268 );
 a78334a <=( (not A302)  and  (not A301) );
 a78335a <=( a78334a  and  a78331a );
 a78336a <=( a78335a  and  a78328a );
 a78340a <=( (not A167)  and  A168 );
 a78341a <=( (not A170)  and  a78340a );
 a78344a <=( A199  and  A166 );
 a78347a <=( A201  and  (not A200) );
 a78348a <=( a78347a  and  a78344a );
 a78349a <=( a78348a  and  a78341a );
 a78352a <=( (not A265)  and  A203 );
 a78355a <=( A267  and  A266 );
 a78356a <=( a78355a  and  a78352a );
 a78359a <=( A300  and  A269 );
 a78362a <=( (not A302)  and  (not A301) );
 a78363a <=( a78362a  and  a78359a );
 a78364a <=( a78363a  and  a78356a );
 a78368a <=( (not A167)  and  A168 );
 a78369a <=( (not A170)  and  a78368a );
 a78372a <=( A199  and  A166 );
 a78375a <=( A201  and  (not A200) );
 a78376a <=( a78375a  and  a78372a );
 a78377a <=( a78376a  and  a78369a );
 a78380a <=( (not A265)  and  A203 );
 a78383a <=( (not A267)  and  A266 );
 a78384a <=( a78383a  and  a78380a );
 a78387a <=( (not A269)  and  (not A268) );
 a78390a <=( A301  and  (not A300) );
 a78391a <=( a78390a  and  a78387a );
 a78392a <=( a78391a  and  a78384a );
 a78396a <=( (not A167)  and  A168 );
 a78397a <=( (not A170)  and  a78396a );
 a78400a <=( A199  and  A166 );
 a78403a <=( A201  and  (not A200) );
 a78404a <=( a78403a  and  a78400a );
 a78405a <=( a78404a  and  a78397a );
 a78408a <=( (not A265)  and  A203 );
 a78411a <=( (not A267)  and  A266 );
 a78412a <=( a78411a  and  a78408a );
 a78415a <=( (not A269)  and  (not A268) );
 a78418a <=( A302  and  (not A300) );
 a78419a <=( a78418a  and  a78415a );
 a78420a <=( a78419a  and  a78412a );
 a78424a <=( (not A167)  and  A168 );
 a78425a <=( (not A170)  and  a78424a );
 a78428a <=( A199  and  A166 );
 a78431a <=( A201  and  (not A200) );
 a78432a <=( a78431a  and  a78428a );
 a78433a <=( a78432a  and  a78425a );
 a78436a <=( (not A265)  and  A203 );
 a78439a <=( (not A267)  and  A266 );
 a78440a <=( a78439a  and  a78436a );
 a78443a <=( (not A269)  and  (not A268) );
 a78446a <=( A299  and  A298 );
 a78447a <=( a78446a  and  a78443a );
 a78448a <=( a78447a  and  a78440a );
 a78452a <=( (not A167)  and  A168 );
 a78453a <=( (not A170)  and  a78452a );
 a78456a <=( A199  and  A166 );
 a78459a <=( A201  and  (not A200) );
 a78460a <=( a78459a  and  a78456a );
 a78461a <=( a78460a  and  a78453a );
 a78464a <=( (not A265)  and  A203 );
 a78467a <=( (not A267)  and  A266 );
 a78468a <=( a78467a  and  a78464a );
 a78471a <=( (not A269)  and  (not A268) );
 a78474a <=( (not A299)  and  (not A298) );
 a78475a <=( a78474a  and  a78471a );
 a78476a <=( a78475a  and  a78468a );
 a78480a <=( (not A167)  and  A168 );
 a78481a <=( (not A170)  and  a78480a );
 a78484a <=( A199  and  A166 );
 a78487a <=( A201  and  (not A200) );
 a78488a <=( a78487a  and  a78484a );
 a78489a <=( a78488a  and  a78481a );
 a78492a <=( A265  and  A203 );
 a78495a <=( A267  and  (not A266) );
 a78496a <=( a78495a  and  a78492a );
 a78499a <=( A300  and  A268 );
 a78502a <=( (not A302)  and  (not A301) );
 a78503a <=( a78502a  and  a78499a );
 a78504a <=( a78503a  and  a78496a );
 a78508a <=( (not A167)  and  A168 );
 a78509a <=( (not A170)  and  a78508a );
 a78512a <=( A199  and  A166 );
 a78515a <=( A201  and  (not A200) );
 a78516a <=( a78515a  and  a78512a );
 a78517a <=( a78516a  and  a78509a );
 a78520a <=( A265  and  A203 );
 a78523a <=( A267  and  (not A266) );
 a78524a <=( a78523a  and  a78520a );
 a78527a <=( A300  and  A269 );
 a78530a <=( (not A302)  and  (not A301) );
 a78531a <=( a78530a  and  a78527a );
 a78532a <=( a78531a  and  a78524a );
 a78536a <=( (not A167)  and  A168 );
 a78537a <=( (not A170)  and  a78536a );
 a78540a <=( A199  and  A166 );
 a78543a <=( A201  and  (not A200) );
 a78544a <=( a78543a  and  a78540a );
 a78545a <=( a78544a  and  a78537a );
 a78548a <=( A265  and  A203 );
 a78551a <=( (not A267)  and  (not A266) );
 a78552a <=( a78551a  and  a78548a );
 a78555a <=( (not A269)  and  (not A268) );
 a78558a <=( A301  and  (not A300) );
 a78559a <=( a78558a  and  a78555a );
 a78560a <=( a78559a  and  a78552a );
 a78564a <=( (not A167)  and  A168 );
 a78565a <=( (not A170)  and  a78564a );
 a78568a <=( A199  and  A166 );
 a78571a <=( A201  and  (not A200) );
 a78572a <=( a78571a  and  a78568a );
 a78573a <=( a78572a  and  a78565a );
 a78576a <=( A265  and  A203 );
 a78579a <=( (not A267)  and  (not A266) );
 a78580a <=( a78579a  and  a78576a );
 a78583a <=( (not A269)  and  (not A268) );
 a78586a <=( A302  and  (not A300) );
 a78587a <=( a78586a  and  a78583a );
 a78588a <=( a78587a  and  a78580a );
 a78592a <=( (not A167)  and  A168 );
 a78593a <=( (not A170)  and  a78592a );
 a78596a <=( A199  and  A166 );
 a78599a <=( A201  and  (not A200) );
 a78600a <=( a78599a  and  a78596a );
 a78601a <=( a78600a  and  a78593a );
 a78604a <=( A265  and  A203 );
 a78607a <=( (not A267)  and  (not A266) );
 a78608a <=( a78607a  and  a78604a );
 a78611a <=( (not A269)  and  (not A268) );
 a78614a <=( A299  and  A298 );
 a78615a <=( a78614a  and  a78611a );
 a78616a <=( a78615a  and  a78608a );
 a78620a <=( (not A167)  and  A168 );
 a78621a <=( (not A170)  and  a78620a );
 a78624a <=( A199  and  A166 );
 a78627a <=( A201  and  (not A200) );
 a78628a <=( a78627a  and  a78624a );
 a78629a <=( a78628a  and  a78621a );
 a78632a <=( A265  and  A203 );
 a78635a <=( (not A267)  and  (not A266) );
 a78636a <=( a78635a  and  a78632a );
 a78639a <=( (not A269)  and  (not A268) );
 a78642a <=( (not A299)  and  (not A298) );
 a78643a <=( a78642a  and  a78639a );
 a78644a <=( a78643a  and  a78636a );
 a78648a <=( (not A167)  and  A168 );
 a78649a <=( (not A170)  and  a78648a );
 a78652a <=( A199  and  A166 );
 a78655a <=( (not A201)  and  (not A200) );
 a78656a <=( a78655a  and  a78652a );
 a78657a <=( a78656a  and  a78649a );
 a78660a <=( (not A203)  and  (not A202) );
 a78663a <=( A266  and  (not A265) );
 a78664a <=( a78663a  and  a78660a );
 a78667a <=( A268  and  A267 );
 a78670a <=( A301  and  (not A300) );
 a78671a <=( a78670a  and  a78667a );
 a78672a <=( a78671a  and  a78664a );
 a78676a <=( (not A167)  and  A168 );
 a78677a <=( (not A170)  and  a78676a );
 a78680a <=( A199  and  A166 );
 a78683a <=( (not A201)  and  (not A200) );
 a78684a <=( a78683a  and  a78680a );
 a78685a <=( a78684a  and  a78677a );
 a78688a <=( (not A203)  and  (not A202) );
 a78691a <=( A266  and  (not A265) );
 a78692a <=( a78691a  and  a78688a );
 a78695a <=( A268  and  A267 );
 a78698a <=( A302  and  (not A300) );
 a78699a <=( a78698a  and  a78695a );
 a78700a <=( a78699a  and  a78692a );
 a78704a <=( (not A167)  and  A168 );
 a78705a <=( (not A170)  and  a78704a );
 a78708a <=( A199  and  A166 );
 a78711a <=( (not A201)  and  (not A200) );
 a78712a <=( a78711a  and  a78708a );
 a78713a <=( a78712a  and  a78705a );
 a78716a <=( (not A203)  and  (not A202) );
 a78719a <=( A266  and  (not A265) );
 a78720a <=( a78719a  and  a78716a );
 a78723a <=( A268  and  A267 );
 a78726a <=( A299  and  A298 );
 a78727a <=( a78726a  and  a78723a );
 a78728a <=( a78727a  and  a78720a );
 a78732a <=( (not A167)  and  A168 );
 a78733a <=( (not A170)  and  a78732a );
 a78736a <=( A199  and  A166 );
 a78739a <=( (not A201)  and  (not A200) );
 a78740a <=( a78739a  and  a78736a );
 a78741a <=( a78740a  and  a78733a );
 a78744a <=( (not A203)  and  (not A202) );
 a78747a <=( A266  and  (not A265) );
 a78748a <=( a78747a  and  a78744a );
 a78751a <=( A268  and  A267 );
 a78754a <=( (not A299)  and  (not A298) );
 a78755a <=( a78754a  and  a78751a );
 a78756a <=( a78755a  and  a78748a );
 a78760a <=( (not A167)  and  A168 );
 a78761a <=( (not A170)  and  a78760a );
 a78764a <=( A199  and  A166 );
 a78767a <=( (not A201)  and  (not A200) );
 a78768a <=( a78767a  and  a78764a );
 a78769a <=( a78768a  and  a78761a );
 a78772a <=( (not A203)  and  (not A202) );
 a78775a <=( A266  and  (not A265) );
 a78776a <=( a78775a  and  a78772a );
 a78779a <=( A269  and  A267 );
 a78782a <=( A301  and  (not A300) );
 a78783a <=( a78782a  and  a78779a );
 a78784a <=( a78783a  and  a78776a );
 a78788a <=( (not A167)  and  A168 );
 a78789a <=( (not A170)  and  a78788a );
 a78792a <=( A199  and  A166 );
 a78795a <=( (not A201)  and  (not A200) );
 a78796a <=( a78795a  and  a78792a );
 a78797a <=( a78796a  and  a78789a );
 a78800a <=( (not A203)  and  (not A202) );
 a78803a <=( A266  and  (not A265) );
 a78804a <=( a78803a  and  a78800a );
 a78807a <=( A269  and  A267 );
 a78810a <=( A302  and  (not A300) );
 a78811a <=( a78810a  and  a78807a );
 a78812a <=( a78811a  and  a78804a );
 a78816a <=( (not A167)  and  A168 );
 a78817a <=( (not A170)  and  a78816a );
 a78820a <=( A199  and  A166 );
 a78823a <=( (not A201)  and  (not A200) );
 a78824a <=( a78823a  and  a78820a );
 a78825a <=( a78824a  and  a78817a );
 a78828a <=( (not A203)  and  (not A202) );
 a78831a <=( A266  and  (not A265) );
 a78832a <=( a78831a  and  a78828a );
 a78835a <=( A269  and  A267 );
 a78838a <=( A299  and  A298 );
 a78839a <=( a78838a  and  a78835a );
 a78840a <=( a78839a  and  a78832a );
 a78844a <=( (not A167)  and  A168 );
 a78845a <=( (not A170)  and  a78844a );
 a78848a <=( A199  and  A166 );
 a78851a <=( (not A201)  and  (not A200) );
 a78852a <=( a78851a  and  a78848a );
 a78853a <=( a78852a  and  a78845a );
 a78856a <=( (not A203)  and  (not A202) );
 a78859a <=( A266  and  (not A265) );
 a78860a <=( a78859a  and  a78856a );
 a78863a <=( A269  and  A267 );
 a78866a <=( (not A299)  and  (not A298) );
 a78867a <=( a78866a  and  a78863a );
 a78868a <=( a78867a  and  a78860a );
 a78872a <=( (not A167)  and  A168 );
 a78873a <=( (not A170)  and  a78872a );
 a78876a <=( A199  and  A166 );
 a78879a <=( (not A201)  and  (not A200) );
 a78880a <=( a78879a  and  a78876a );
 a78881a <=( a78880a  and  a78873a );
 a78884a <=( (not A203)  and  (not A202) );
 a78887a <=( (not A266)  and  A265 );
 a78888a <=( a78887a  and  a78884a );
 a78891a <=( A268  and  A267 );
 a78894a <=( A301  and  (not A300) );
 a78895a <=( a78894a  and  a78891a );
 a78896a <=( a78895a  and  a78888a );
 a78900a <=( (not A167)  and  A168 );
 a78901a <=( (not A170)  and  a78900a );
 a78904a <=( A199  and  A166 );
 a78907a <=( (not A201)  and  (not A200) );
 a78908a <=( a78907a  and  a78904a );
 a78909a <=( a78908a  and  a78901a );
 a78912a <=( (not A203)  and  (not A202) );
 a78915a <=( (not A266)  and  A265 );
 a78916a <=( a78915a  and  a78912a );
 a78919a <=( A268  and  A267 );
 a78922a <=( A302  and  (not A300) );
 a78923a <=( a78922a  and  a78919a );
 a78924a <=( a78923a  and  a78916a );
 a78928a <=( (not A167)  and  A168 );
 a78929a <=( (not A170)  and  a78928a );
 a78932a <=( A199  and  A166 );
 a78935a <=( (not A201)  and  (not A200) );
 a78936a <=( a78935a  and  a78932a );
 a78937a <=( a78936a  and  a78929a );
 a78940a <=( (not A203)  and  (not A202) );
 a78943a <=( (not A266)  and  A265 );
 a78944a <=( a78943a  and  a78940a );
 a78947a <=( A268  and  A267 );
 a78950a <=( A299  and  A298 );
 a78951a <=( a78950a  and  a78947a );
 a78952a <=( a78951a  and  a78944a );
 a78956a <=( (not A167)  and  A168 );
 a78957a <=( (not A170)  and  a78956a );
 a78960a <=( A199  and  A166 );
 a78963a <=( (not A201)  and  (not A200) );
 a78964a <=( a78963a  and  a78960a );
 a78965a <=( a78964a  and  a78957a );
 a78968a <=( (not A203)  and  (not A202) );
 a78971a <=( (not A266)  and  A265 );
 a78972a <=( a78971a  and  a78968a );
 a78975a <=( A268  and  A267 );
 a78978a <=( (not A299)  and  (not A298) );
 a78979a <=( a78978a  and  a78975a );
 a78980a <=( a78979a  and  a78972a );
 a78984a <=( (not A167)  and  A168 );
 a78985a <=( (not A170)  and  a78984a );
 a78988a <=( A199  and  A166 );
 a78991a <=( (not A201)  and  (not A200) );
 a78992a <=( a78991a  and  a78988a );
 a78993a <=( a78992a  and  a78985a );
 a78996a <=( (not A203)  and  (not A202) );
 a78999a <=( (not A266)  and  A265 );
 a79000a <=( a78999a  and  a78996a );
 a79003a <=( A269  and  A267 );
 a79006a <=( A301  and  (not A300) );
 a79007a <=( a79006a  and  a79003a );
 a79008a <=( a79007a  and  a79000a );
 a79012a <=( (not A167)  and  A168 );
 a79013a <=( (not A170)  and  a79012a );
 a79016a <=( A199  and  A166 );
 a79019a <=( (not A201)  and  (not A200) );
 a79020a <=( a79019a  and  a79016a );
 a79021a <=( a79020a  and  a79013a );
 a79024a <=( (not A203)  and  (not A202) );
 a79027a <=( (not A266)  and  A265 );
 a79028a <=( a79027a  and  a79024a );
 a79031a <=( A269  and  A267 );
 a79034a <=( A302  and  (not A300) );
 a79035a <=( a79034a  and  a79031a );
 a79036a <=( a79035a  and  a79028a );
 a79040a <=( (not A167)  and  A168 );
 a79041a <=( (not A170)  and  a79040a );
 a79044a <=( A199  and  A166 );
 a79047a <=( (not A201)  and  (not A200) );
 a79048a <=( a79047a  and  a79044a );
 a79049a <=( a79048a  and  a79041a );
 a79052a <=( (not A203)  and  (not A202) );
 a79055a <=( (not A266)  and  A265 );
 a79056a <=( a79055a  and  a79052a );
 a79059a <=( A269  and  A267 );
 a79062a <=( A299  and  A298 );
 a79063a <=( a79062a  and  a79059a );
 a79064a <=( a79063a  and  a79056a );
 a79068a <=( (not A167)  and  A168 );
 a79069a <=( (not A170)  and  a79068a );
 a79072a <=( A199  and  A166 );
 a79075a <=( (not A201)  and  (not A200) );
 a79076a <=( a79075a  and  a79072a );
 a79077a <=( a79076a  and  a79069a );
 a79080a <=( (not A203)  and  (not A202) );
 a79083a <=( (not A266)  and  A265 );
 a79084a <=( a79083a  and  a79080a );
 a79087a <=( A269  and  A267 );
 a79090a <=( (not A299)  and  (not A298) );
 a79091a <=( a79090a  and  a79087a );
 a79092a <=( a79091a  and  a79084a );
 a79096a <=( (not A199)  and  (not A168) );
 a79097a <=( (not A170)  and  a79096a );
 a79100a <=( (not A201)  and  A200 );
 a79103a <=( (not A203)  and  (not A202) );
 a79104a <=( a79103a  and  a79100a );
 a79105a <=( a79104a  and  a79097a );
 a79108a <=( (not A268)  and  A267 );
 a79111a <=( A298  and  (not A269) );
 a79112a <=( a79111a  and  a79108a );
 a79115a <=( (not A300)  and  (not A299) );
 a79118a <=( (not A302)  and  (not A301) );
 a79119a <=( a79118a  and  a79115a );
 a79120a <=( a79119a  and  a79112a );
 a79124a <=( (not A199)  and  (not A168) );
 a79125a <=( (not A170)  and  a79124a );
 a79128a <=( (not A201)  and  A200 );
 a79131a <=( (not A203)  and  (not A202) );
 a79132a <=( a79131a  and  a79128a );
 a79133a <=( a79132a  and  a79125a );
 a79136a <=( (not A268)  and  A267 );
 a79139a <=( (not A298)  and  (not A269) );
 a79140a <=( a79139a  and  a79136a );
 a79143a <=( (not A300)  and  A299 );
 a79146a <=( (not A302)  and  (not A301) );
 a79147a <=( a79146a  and  a79143a );
 a79148a <=( a79147a  and  a79140a );
 a79152a <=( A199  and  (not A168) );
 a79153a <=( (not A170)  and  a79152a );
 a79156a <=( (not A201)  and  (not A200) );
 a79159a <=( (not A203)  and  (not A202) );
 a79160a <=( a79159a  and  a79156a );
 a79161a <=( a79160a  and  a79153a );
 a79164a <=( (not A268)  and  A267 );
 a79167a <=( A298  and  (not A269) );
 a79168a <=( a79167a  and  a79164a );
 a79171a <=( (not A300)  and  (not A299) );
 a79174a <=( (not A302)  and  (not A301) );
 a79175a <=( a79174a  and  a79171a );
 a79176a <=( a79175a  and  a79168a );
 a79180a <=( A199  and  (not A168) );
 a79181a <=( (not A170)  and  a79180a );
 a79184a <=( (not A201)  and  (not A200) );
 a79187a <=( (not A203)  and  (not A202) );
 a79188a <=( a79187a  and  a79184a );
 a79189a <=( a79188a  and  a79181a );
 a79192a <=( (not A268)  and  A267 );
 a79195a <=( (not A298)  and  (not A269) );
 a79196a <=( a79195a  and  a79192a );
 a79199a <=( (not A300)  and  A299 );
 a79202a <=( (not A302)  and  (not A301) );
 a79203a <=( a79202a  and  a79199a );
 a79204a <=( a79203a  and  a79196a );
 a79208a <=( A167  and  A168 );
 a79209a <=( A169  and  a79208a );
 a79212a <=( A201  and  (not A166) );
 a79215a <=( (not A203)  and  (not A202) );
 a79216a <=( a79215a  and  a79212a );
 a79217a <=( a79216a  and  a79209a );
 a79220a <=( (not A268)  and  A267 );
 a79223a <=( A298  and  (not A269) );
 a79224a <=( a79223a  and  a79220a );
 a79227a <=( (not A300)  and  (not A299) );
 a79230a <=( (not A302)  and  (not A301) );
 a79231a <=( a79230a  and  a79227a );
 a79232a <=( a79231a  and  a79224a );
 a79236a <=( A167  and  A168 );
 a79237a <=( A169  and  a79236a );
 a79240a <=( A201  and  (not A166) );
 a79243a <=( (not A203)  and  (not A202) );
 a79244a <=( a79243a  and  a79240a );
 a79245a <=( a79244a  and  a79237a );
 a79248a <=( (not A268)  and  A267 );
 a79251a <=( (not A298)  and  (not A269) );
 a79252a <=( a79251a  and  a79248a );
 a79255a <=( (not A300)  and  A299 );
 a79258a <=( (not A302)  and  (not A301) );
 a79259a <=( a79258a  and  a79255a );
 a79260a <=( a79259a  and  a79252a );
 a79264a <=( A167  and  A168 );
 a79265a <=( A169  and  a79264a );
 a79268a <=( (not A199)  and  (not A166) );
 a79271a <=( A201  and  A200 );
 a79272a <=( a79271a  and  a79268a );
 a79273a <=( a79272a  and  a79265a );
 a79276a <=( (not A265)  and  A202 );
 a79279a <=( A267  and  A266 );
 a79280a <=( a79279a  and  a79276a );
 a79283a <=( A300  and  A268 );
 a79286a <=( (not A302)  and  (not A301) );
 a79287a <=( a79286a  and  a79283a );
 a79288a <=( a79287a  and  a79280a );
 a79292a <=( A167  and  A168 );
 a79293a <=( A169  and  a79292a );
 a79296a <=( (not A199)  and  (not A166) );
 a79299a <=( A201  and  A200 );
 a79300a <=( a79299a  and  a79296a );
 a79301a <=( a79300a  and  a79293a );
 a79304a <=( (not A265)  and  A202 );
 a79307a <=( A267  and  A266 );
 a79308a <=( a79307a  and  a79304a );
 a79311a <=( A300  and  A269 );
 a79314a <=( (not A302)  and  (not A301) );
 a79315a <=( a79314a  and  a79311a );
 a79316a <=( a79315a  and  a79308a );
 a79320a <=( A167  and  A168 );
 a79321a <=( A169  and  a79320a );
 a79324a <=( (not A199)  and  (not A166) );
 a79327a <=( A201  and  A200 );
 a79328a <=( a79327a  and  a79324a );
 a79329a <=( a79328a  and  a79321a );
 a79332a <=( (not A265)  and  A202 );
 a79335a <=( (not A267)  and  A266 );
 a79336a <=( a79335a  and  a79332a );
 a79339a <=( (not A269)  and  (not A268) );
 a79342a <=( A301  and  (not A300) );
 a79343a <=( a79342a  and  a79339a );
 a79344a <=( a79343a  and  a79336a );
 a79348a <=( A167  and  A168 );
 a79349a <=( A169  and  a79348a );
 a79352a <=( (not A199)  and  (not A166) );
 a79355a <=( A201  and  A200 );
 a79356a <=( a79355a  and  a79352a );
 a79357a <=( a79356a  and  a79349a );
 a79360a <=( (not A265)  and  A202 );
 a79363a <=( (not A267)  and  A266 );
 a79364a <=( a79363a  and  a79360a );
 a79367a <=( (not A269)  and  (not A268) );
 a79370a <=( A302  and  (not A300) );
 a79371a <=( a79370a  and  a79367a );
 a79372a <=( a79371a  and  a79364a );
 a79376a <=( A167  and  A168 );
 a79377a <=( A169  and  a79376a );
 a79380a <=( (not A199)  and  (not A166) );
 a79383a <=( A201  and  A200 );
 a79384a <=( a79383a  and  a79380a );
 a79385a <=( a79384a  and  a79377a );
 a79388a <=( (not A265)  and  A202 );
 a79391a <=( (not A267)  and  A266 );
 a79392a <=( a79391a  and  a79388a );
 a79395a <=( (not A269)  and  (not A268) );
 a79398a <=( A299  and  A298 );
 a79399a <=( a79398a  and  a79395a );
 a79400a <=( a79399a  and  a79392a );
 a79404a <=( A167  and  A168 );
 a79405a <=( A169  and  a79404a );
 a79408a <=( (not A199)  and  (not A166) );
 a79411a <=( A201  and  A200 );
 a79412a <=( a79411a  and  a79408a );
 a79413a <=( a79412a  and  a79405a );
 a79416a <=( (not A265)  and  A202 );
 a79419a <=( (not A267)  and  A266 );
 a79420a <=( a79419a  and  a79416a );
 a79423a <=( (not A269)  and  (not A268) );
 a79426a <=( (not A299)  and  (not A298) );
 a79427a <=( a79426a  and  a79423a );
 a79428a <=( a79427a  and  a79420a );
 a79432a <=( A167  and  A168 );
 a79433a <=( A169  and  a79432a );
 a79436a <=( (not A199)  and  (not A166) );
 a79439a <=( A201  and  A200 );
 a79440a <=( a79439a  and  a79436a );
 a79441a <=( a79440a  and  a79433a );
 a79444a <=( A265  and  A202 );
 a79447a <=( A267  and  (not A266) );
 a79448a <=( a79447a  and  a79444a );
 a79451a <=( A300  and  A268 );
 a79454a <=( (not A302)  and  (not A301) );
 a79455a <=( a79454a  and  a79451a );
 a79456a <=( a79455a  and  a79448a );
 a79460a <=( A167  and  A168 );
 a79461a <=( A169  and  a79460a );
 a79464a <=( (not A199)  and  (not A166) );
 a79467a <=( A201  and  A200 );
 a79468a <=( a79467a  and  a79464a );
 a79469a <=( a79468a  and  a79461a );
 a79472a <=( A265  and  A202 );
 a79475a <=( A267  and  (not A266) );
 a79476a <=( a79475a  and  a79472a );
 a79479a <=( A300  and  A269 );
 a79482a <=( (not A302)  and  (not A301) );
 a79483a <=( a79482a  and  a79479a );
 a79484a <=( a79483a  and  a79476a );
 a79488a <=( A167  and  A168 );
 a79489a <=( A169  and  a79488a );
 a79492a <=( (not A199)  and  (not A166) );
 a79495a <=( A201  and  A200 );
 a79496a <=( a79495a  and  a79492a );
 a79497a <=( a79496a  and  a79489a );
 a79500a <=( A265  and  A202 );
 a79503a <=( (not A267)  and  (not A266) );
 a79504a <=( a79503a  and  a79500a );
 a79507a <=( (not A269)  and  (not A268) );
 a79510a <=( A301  and  (not A300) );
 a79511a <=( a79510a  and  a79507a );
 a79512a <=( a79511a  and  a79504a );
 a79516a <=( A167  and  A168 );
 a79517a <=( A169  and  a79516a );
 a79520a <=( (not A199)  and  (not A166) );
 a79523a <=( A201  and  A200 );
 a79524a <=( a79523a  and  a79520a );
 a79525a <=( a79524a  and  a79517a );
 a79528a <=( A265  and  A202 );
 a79531a <=( (not A267)  and  (not A266) );
 a79532a <=( a79531a  and  a79528a );
 a79535a <=( (not A269)  and  (not A268) );
 a79538a <=( A302  and  (not A300) );
 a79539a <=( a79538a  and  a79535a );
 a79540a <=( a79539a  and  a79532a );
 a79544a <=( A167  and  A168 );
 a79545a <=( A169  and  a79544a );
 a79548a <=( (not A199)  and  (not A166) );
 a79551a <=( A201  and  A200 );
 a79552a <=( a79551a  and  a79548a );
 a79553a <=( a79552a  and  a79545a );
 a79556a <=( A265  and  A202 );
 a79559a <=( (not A267)  and  (not A266) );
 a79560a <=( a79559a  and  a79556a );
 a79563a <=( (not A269)  and  (not A268) );
 a79566a <=( A299  and  A298 );
 a79567a <=( a79566a  and  a79563a );
 a79568a <=( a79567a  and  a79560a );
 a79572a <=( A167  and  A168 );
 a79573a <=( A169  and  a79572a );
 a79576a <=( (not A199)  and  (not A166) );
 a79579a <=( A201  and  A200 );
 a79580a <=( a79579a  and  a79576a );
 a79581a <=( a79580a  and  a79573a );
 a79584a <=( A265  and  A202 );
 a79587a <=( (not A267)  and  (not A266) );
 a79588a <=( a79587a  and  a79584a );
 a79591a <=( (not A269)  and  (not A268) );
 a79594a <=( (not A299)  and  (not A298) );
 a79595a <=( a79594a  and  a79591a );
 a79596a <=( a79595a  and  a79588a );
 a79600a <=( A167  and  A168 );
 a79601a <=( A169  and  a79600a );
 a79604a <=( (not A199)  and  (not A166) );
 a79607a <=( A201  and  A200 );
 a79608a <=( a79607a  and  a79604a );
 a79609a <=( a79608a  and  a79601a );
 a79612a <=( (not A265)  and  A203 );
 a79615a <=( A267  and  A266 );
 a79616a <=( a79615a  and  a79612a );
 a79619a <=( A300  and  A268 );
 a79622a <=( (not A302)  and  (not A301) );
 a79623a <=( a79622a  and  a79619a );
 a79624a <=( a79623a  and  a79616a );
 a79628a <=( A167  and  A168 );
 a79629a <=( A169  and  a79628a );
 a79632a <=( (not A199)  and  (not A166) );
 a79635a <=( A201  and  A200 );
 a79636a <=( a79635a  and  a79632a );
 a79637a <=( a79636a  and  a79629a );
 a79640a <=( (not A265)  and  A203 );
 a79643a <=( A267  and  A266 );
 a79644a <=( a79643a  and  a79640a );
 a79647a <=( A300  and  A269 );
 a79650a <=( (not A302)  and  (not A301) );
 a79651a <=( a79650a  and  a79647a );
 a79652a <=( a79651a  and  a79644a );
 a79656a <=( A167  and  A168 );
 a79657a <=( A169  and  a79656a );
 a79660a <=( (not A199)  and  (not A166) );
 a79663a <=( A201  and  A200 );
 a79664a <=( a79663a  and  a79660a );
 a79665a <=( a79664a  and  a79657a );
 a79668a <=( (not A265)  and  A203 );
 a79671a <=( (not A267)  and  A266 );
 a79672a <=( a79671a  and  a79668a );
 a79675a <=( (not A269)  and  (not A268) );
 a79678a <=( A301  and  (not A300) );
 a79679a <=( a79678a  and  a79675a );
 a79680a <=( a79679a  and  a79672a );
 a79684a <=( A167  and  A168 );
 a79685a <=( A169  and  a79684a );
 a79688a <=( (not A199)  and  (not A166) );
 a79691a <=( A201  and  A200 );
 a79692a <=( a79691a  and  a79688a );
 a79693a <=( a79692a  and  a79685a );
 a79696a <=( (not A265)  and  A203 );
 a79699a <=( (not A267)  and  A266 );
 a79700a <=( a79699a  and  a79696a );
 a79703a <=( (not A269)  and  (not A268) );
 a79706a <=( A302  and  (not A300) );
 a79707a <=( a79706a  and  a79703a );
 a79708a <=( a79707a  and  a79700a );
 a79712a <=( A167  and  A168 );
 a79713a <=( A169  and  a79712a );
 a79716a <=( (not A199)  and  (not A166) );
 a79719a <=( A201  and  A200 );
 a79720a <=( a79719a  and  a79716a );
 a79721a <=( a79720a  and  a79713a );
 a79724a <=( (not A265)  and  A203 );
 a79727a <=( (not A267)  and  A266 );
 a79728a <=( a79727a  and  a79724a );
 a79731a <=( (not A269)  and  (not A268) );
 a79734a <=( A299  and  A298 );
 a79735a <=( a79734a  and  a79731a );
 a79736a <=( a79735a  and  a79728a );
 a79740a <=( A167  and  A168 );
 a79741a <=( A169  and  a79740a );
 a79744a <=( (not A199)  and  (not A166) );
 a79747a <=( A201  and  A200 );
 a79748a <=( a79747a  and  a79744a );
 a79749a <=( a79748a  and  a79741a );
 a79752a <=( (not A265)  and  A203 );
 a79755a <=( (not A267)  and  A266 );
 a79756a <=( a79755a  and  a79752a );
 a79759a <=( (not A269)  and  (not A268) );
 a79762a <=( (not A299)  and  (not A298) );
 a79763a <=( a79762a  and  a79759a );
 a79764a <=( a79763a  and  a79756a );
 a79768a <=( A167  and  A168 );
 a79769a <=( A169  and  a79768a );
 a79772a <=( (not A199)  and  (not A166) );
 a79775a <=( A201  and  A200 );
 a79776a <=( a79775a  and  a79772a );
 a79777a <=( a79776a  and  a79769a );
 a79780a <=( A265  and  A203 );
 a79783a <=( A267  and  (not A266) );
 a79784a <=( a79783a  and  a79780a );
 a79787a <=( A300  and  A268 );
 a79790a <=( (not A302)  and  (not A301) );
 a79791a <=( a79790a  and  a79787a );
 a79792a <=( a79791a  and  a79784a );
 a79796a <=( A167  and  A168 );
 a79797a <=( A169  and  a79796a );
 a79800a <=( (not A199)  and  (not A166) );
 a79803a <=( A201  and  A200 );
 a79804a <=( a79803a  and  a79800a );
 a79805a <=( a79804a  and  a79797a );
 a79808a <=( A265  and  A203 );
 a79811a <=( A267  and  (not A266) );
 a79812a <=( a79811a  and  a79808a );
 a79815a <=( A300  and  A269 );
 a79818a <=( (not A302)  and  (not A301) );
 a79819a <=( a79818a  and  a79815a );
 a79820a <=( a79819a  and  a79812a );
 a79824a <=( A167  and  A168 );
 a79825a <=( A169  and  a79824a );
 a79828a <=( (not A199)  and  (not A166) );
 a79831a <=( A201  and  A200 );
 a79832a <=( a79831a  and  a79828a );
 a79833a <=( a79832a  and  a79825a );
 a79836a <=( A265  and  A203 );
 a79839a <=( (not A267)  and  (not A266) );
 a79840a <=( a79839a  and  a79836a );
 a79843a <=( (not A269)  and  (not A268) );
 a79846a <=( A301  and  (not A300) );
 a79847a <=( a79846a  and  a79843a );
 a79848a <=( a79847a  and  a79840a );
 a79852a <=( A167  and  A168 );
 a79853a <=( A169  and  a79852a );
 a79856a <=( (not A199)  and  (not A166) );
 a79859a <=( A201  and  A200 );
 a79860a <=( a79859a  and  a79856a );
 a79861a <=( a79860a  and  a79853a );
 a79864a <=( A265  and  A203 );
 a79867a <=( (not A267)  and  (not A266) );
 a79868a <=( a79867a  and  a79864a );
 a79871a <=( (not A269)  and  (not A268) );
 a79874a <=( A302  and  (not A300) );
 a79875a <=( a79874a  and  a79871a );
 a79876a <=( a79875a  and  a79868a );
 a79880a <=( A167  and  A168 );
 a79881a <=( A169  and  a79880a );
 a79884a <=( (not A199)  and  (not A166) );
 a79887a <=( A201  and  A200 );
 a79888a <=( a79887a  and  a79884a );
 a79889a <=( a79888a  and  a79881a );
 a79892a <=( A265  and  A203 );
 a79895a <=( (not A267)  and  (not A266) );
 a79896a <=( a79895a  and  a79892a );
 a79899a <=( (not A269)  and  (not A268) );
 a79902a <=( A299  and  A298 );
 a79903a <=( a79902a  and  a79899a );
 a79904a <=( a79903a  and  a79896a );
 a79908a <=( A167  and  A168 );
 a79909a <=( A169  and  a79908a );
 a79912a <=( (not A199)  and  (not A166) );
 a79915a <=( A201  and  A200 );
 a79916a <=( a79915a  and  a79912a );
 a79917a <=( a79916a  and  a79909a );
 a79920a <=( A265  and  A203 );
 a79923a <=( (not A267)  and  (not A266) );
 a79924a <=( a79923a  and  a79920a );
 a79927a <=( (not A269)  and  (not A268) );
 a79930a <=( (not A299)  and  (not A298) );
 a79931a <=( a79930a  and  a79927a );
 a79932a <=( a79931a  and  a79924a );
 a79936a <=( A167  and  A168 );
 a79937a <=( A169  and  a79936a );
 a79940a <=( (not A199)  and  (not A166) );
 a79943a <=( (not A201)  and  A200 );
 a79944a <=( a79943a  and  a79940a );
 a79945a <=( a79944a  and  a79937a );
 a79948a <=( (not A203)  and  (not A202) );
 a79951a <=( A266  and  (not A265) );
 a79952a <=( a79951a  and  a79948a );
 a79955a <=( A268  and  A267 );
 a79958a <=( A301  and  (not A300) );
 a79959a <=( a79958a  and  a79955a );
 a79960a <=( a79959a  and  a79952a );
 a79964a <=( A167  and  A168 );
 a79965a <=( A169  and  a79964a );
 a79968a <=( (not A199)  and  (not A166) );
 a79971a <=( (not A201)  and  A200 );
 a79972a <=( a79971a  and  a79968a );
 a79973a <=( a79972a  and  a79965a );
 a79976a <=( (not A203)  and  (not A202) );
 a79979a <=( A266  and  (not A265) );
 a79980a <=( a79979a  and  a79976a );
 a79983a <=( A268  and  A267 );
 a79986a <=( A302  and  (not A300) );
 a79987a <=( a79986a  and  a79983a );
 a79988a <=( a79987a  and  a79980a );
 a79992a <=( A167  and  A168 );
 a79993a <=( A169  and  a79992a );
 a79996a <=( (not A199)  and  (not A166) );
 a79999a <=( (not A201)  and  A200 );
 a80000a <=( a79999a  and  a79996a );
 a80001a <=( a80000a  and  a79993a );
 a80004a <=( (not A203)  and  (not A202) );
 a80007a <=( A266  and  (not A265) );
 a80008a <=( a80007a  and  a80004a );
 a80011a <=( A268  and  A267 );
 a80014a <=( A299  and  A298 );
 a80015a <=( a80014a  and  a80011a );
 a80016a <=( a80015a  and  a80008a );
 a80020a <=( A167  and  A168 );
 a80021a <=( A169  and  a80020a );
 a80024a <=( (not A199)  and  (not A166) );
 a80027a <=( (not A201)  and  A200 );
 a80028a <=( a80027a  and  a80024a );
 a80029a <=( a80028a  and  a80021a );
 a80032a <=( (not A203)  and  (not A202) );
 a80035a <=( A266  and  (not A265) );
 a80036a <=( a80035a  and  a80032a );
 a80039a <=( A268  and  A267 );
 a80042a <=( (not A299)  and  (not A298) );
 a80043a <=( a80042a  and  a80039a );
 a80044a <=( a80043a  and  a80036a );
 a80048a <=( A167  and  A168 );
 a80049a <=( A169  and  a80048a );
 a80052a <=( (not A199)  and  (not A166) );
 a80055a <=( (not A201)  and  A200 );
 a80056a <=( a80055a  and  a80052a );
 a80057a <=( a80056a  and  a80049a );
 a80060a <=( (not A203)  and  (not A202) );
 a80063a <=( A266  and  (not A265) );
 a80064a <=( a80063a  and  a80060a );
 a80067a <=( A269  and  A267 );
 a80070a <=( A301  and  (not A300) );
 a80071a <=( a80070a  and  a80067a );
 a80072a <=( a80071a  and  a80064a );
 a80076a <=( A167  and  A168 );
 a80077a <=( A169  and  a80076a );
 a80080a <=( (not A199)  and  (not A166) );
 a80083a <=( (not A201)  and  A200 );
 a80084a <=( a80083a  and  a80080a );
 a80085a <=( a80084a  and  a80077a );
 a80088a <=( (not A203)  and  (not A202) );
 a80091a <=( A266  and  (not A265) );
 a80092a <=( a80091a  and  a80088a );
 a80095a <=( A269  and  A267 );
 a80098a <=( A302  and  (not A300) );
 a80099a <=( a80098a  and  a80095a );
 a80100a <=( a80099a  and  a80092a );
 a80104a <=( A167  and  A168 );
 a80105a <=( A169  and  a80104a );
 a80108a <=( (not A199)  and  (not A166) );
 a80111a <=( (not A201)  and  A200 );
 a80112a <=( a80111a  and  a80108a );
 a80113a <=( a80112a  and  a80105a );
 a80116a <=( (not A203)  and  (not A202) );
 a80119a <=( A266  and  (not A265) );
 a80120a <=( a80119a  and  a80116a );
 a80123a <=( A269  and  A267 );
 a80126a <=( A299  and  A298 );
 a80127a <=( a80126a  and  a80123a );
 a80128a <=( a80127a  and  a80120a );
 a80132a <=( A167  and  A168 );
 a80133a <=( A169  and  a80132a );
 a80136a <=( (not A199)  and  (not A166) );
 a80139a <=( (not A201)  and  A200 );
 a80140a <=( a80139a  and  a80136a );
 a80141a <=( a80140a  and  a80133a );
 a80144a <=( (not A203)  and  (not A202) );
 a80147a <=( A266  and  (not A265) );
 a80148a <=( a80147a  and  a80144a );
 a80151a <=( A269  and  A267 );
 a80154a <=( (not A299)  and  (not A298) );
 a80155a <=( a80154a  and  a80151a );
 a80156a <=( a80155a  and  a80148a );
 a80160a <=( A167  and  A168 );
 a80161a <=( A169  and  a80160a );
 a80164a <=( (not A199)  and  (not A166) );
 a80167a <=( (not A201)  and  A200 );
 a80168a <=( a80167a  and  a80164a );
 a80169a <=( a80168a  and  a80161a );
 a80172a <=( (not A203)  and  (not A202) );
 a80175a <=( (not A266)  and  A265 );
 a80176a <=( a80175a  and  a80172a );
 a80179a <=( A268  and  A267 );
 a80182a <=( A301  and  (not A300) );
 a80183a <=( a80182a  and  a80179a );
 a80184a <=( a80183a  and  a80176a );
 a80188a <=( A167  and  A168 );
 a80189a <=( A169  and  a80188a );
 a80192a <=( (not A199)  and  (not A166) );
 a80195a <=( (not A201)  and  A200 );
 a80196a <=( a80195a  and  a80192a );
 a80197a <=( a80196a  and  a80189a );
 a80200a <=( (not A203)  and  (not A202) );
 a80203a <=( (not A266)  and  A265 );
 a80204a <=( a80203a  and  a80200a );
 a80207a <=( A268  and  A267 );
 a80210a <=( A302  and  (not A300) );
 a80211a <=( a80210a  and  a80207a );
 a80212a <=( a80211a  and  a80204a );
 a80216a <=( A167  and  A168 );
 a80217a <=( A169  and  a80216a );
 a80220a <=( (not A199)  and  (not A166) );
 a80223a <=( (not A201)  and  A200 );
 a80224a <=( a80223a  and  a80220a );
 a80225a <=( a80224a  and  a80217a );
 a80228a <=( (not A203)  and  (not A202) );
 a80231a <=( (not A266)  and  A265 );
 a80232a <=( a80231a  and  a80228a );
 a80235a <=( A268  and  A267 );
 a80238a <=( A299  and  A298 );
 a80239a <=( a80238a  and  a80235a );
 a80240a <=( a80239a  and  a80232a );
 a80244a <=( A167  and  A168 );
 a80245a <=( A169  and  a80244a );
 a80248a <=( (not A199)  and  (not A166) );
 a80251a <=( (not A201)  and  A200 );
 a80252a <=( a80251a  and  a80248a );
 a80253a <=( a80252a  and  a80245a );
 a80256a <=( (not A203)  and  (not A202) );
 a80259a <=( (not A266)  and  A265 );
 a80260a <=( a80259a  and  a80256a );
 a80263a <=( A268  and  A267 );
 a80266a <=( (not A299)  and  (not A298) );
 a80267a <=( a80266a  and  a80263a );
 a80268a <=( a80267a  and  a80260a );
 a80272a <=( A167  and  A168 );
 a80273a <=( A169  and  a80272a );
 a80276a <=( (not A199)  and  (not A166) );
 a80279a <=( (not A201)  and  A200 );
 a80280a <=( a80279a  and  a80276a );
 a80281a <=( a80280a  and  a80273a );
 a80284a <=( (not A203)  and  (not A202) );
 a80287a <=( (not A266)  and  A265 );
 a80288a <=( a80287a  and  a80284a );
 a80291a <=( A269  and  A267 );
 a80294a <=( A301  and  (not A300) );
 a80295a <=( a80294a  and  a80291a );
 a80296a <=( a80295a  and  a80288a );
 a80300a <=( A167  and  A168 );
 a80301a <=( A169  and  a80300a );
 a80304a <=( (not A199)  and  (not A166) );
 a80307a <=( (not A201)  and  A200 );
 a80308a <=( a80307a  and  a80304a );
 a80309a <=( a80308a  and  a80301a );
 a80312a <=( (not A203)  and  (not A202) );
 a80315a <=( (not A266)  and  A265 );
 a80316a <=( a80315a  and  a80312a );
 a80319a <=( A269  and  A267 );
 a80322a <=( A302  and  (not A300) );
 a80323a <=( a80322a  and  a80319a );
 a80324a <=( a80323a  and  a80316a );
 a80328a <=( A167  and  A168 );
 a80329a <=( A169  and  a80328a );
 a80332a <=( (not A199)  and  (not A166) );
 a80335a <=( (not A201)  and  A200 );
 a80336a <=( a80335a  and  a80332a );
 a80337a <=( a80336a  and  a80329a );
 a80340a <=( (not A203)  and  (not A202) );
 a80343a <=( (not A266)  and  A265 );
 a80344a <=( a80343a  and  a80340a );
 a80347a <=( A269  and  A267 );
 a80350a <=( A299  and  A298 );
 a80351a <=( a80350a  and  a80347a );
 a80352a <=( a80351a  and  a80344a );
 a80356a <=( A167  and  A168 );
 a80357a <=( A169  and  a80356a );
 a80360a <=( (not A199)  and  (not A166) );
 a80363a <=( (not A201)  and  A200 );
 a80364a <=( a80363a  and  a80360a );
 a80365a <=( a80364a  and  a80357a );
 a80368a <=( (not A203)  and  (not A202) );
 a80371a <=( (not A266)  and  A265 );
 a80372a <=( a80371a  and  a80368a );
 a80375a <=( A269  and  A267 );
 a80378a <=( (not A299)  and  (not A298) );
 a80379a <=( a80378a  and  a80375a );
 a80380a <=( a80379a  and  a80372a );
 a80384a <=( A167  and  A168 );
 a80385a <=( A169  and  a80384a );
 a80388a <=( A199  and  (not A166) );
 a80391a <=( A201  and  (not A200) );
 a80392a <=( a80391a  and  a80388a );
 a80393a <=( a80392a  and  a80385a );
 a80396a <=( (not A265)  and  A202 );
 a80399a <=( A267  and  A266 );
 a80400a <=( a80399a  and  a80396a );
 a80403a <=( A300  and  A268 );
 a80406a <=( (not A302)  and  (not A301) );
 a80407a <=( a80406a  and  a80403a );
 a80408a <=( a80407a  and  a80400a );
 a80412a <=( A167  and  A168 );
 a80413a <=( A169  and  a80412a );
 a80416a <=( A199  and  (not A166) );
 a80419a <=( A201  and  (not A200) );
 a80420a <=( a80419a  and  a80416a );
 a80421a <=( a80420a  and  a80413a );
 a80424a <=( (not A265)  and  A202 );
 a80427a <=( A267  and  A266 );
 a80428a <=( a80427a  and  a80424a );
 a80431a <=( A300  and  A269 );
 a80434a <=( (not A302)  and  (not A301) );
 a80435a <=( a80434a  and  a80431a );
 a80436a <=( a80435a  and  a80428a );
 a80440a <=( A167  and  A168 );
 a80441a <=( A169  and  a80440a );
 a80444a <=( A199  and  (not A166) );
 a80447a <=( A201  and  (not A200) );
 a80448a <=( a80447a  and  a80444a );
 a80449a <=( a80448a  and  a80441a );
 a80452a <=( (not A265)  and  A202 );
 a80455a <=( (not A267)  and  A266 );
 a80456a <=( a80455a  and  a80452a );
 a80459a <=( (not A269)  and  (not A268) );
 a80462a <=( A301  and  (not A300) );
 a80463a <=( a80462a  and  a80459a );
 a80464a <=( a80463a  and  a80456a );
 a80468a <=( A167  and  A168 );
 a80469a <=( A169  and  a80468a );
 a80472a <=( A199  and  (not A166) );
 a80475a <=( A201  and  (not A200) );
 a80476a <=( a80475a  and  a80472a );
 a80477a <=( a80476a  and  a80469a );
 a80480a <=( (not A265)  and  A202 );
 a80483a <=( (not A267)  and  A266 );
 a80484a <=( a80483a  and  a80480a );
 a80487a <=( (not A269)  and  (not A268) );
 a80490a <=( A302  and  (not A300) );
 a80491a <=( a80490a  and  a80487a );
 a80492a <=( a80491a  and  a80484a );
 a80496a <=( A167  and  A168 );
 a80497a <=( A169  and  a80496a );
 a80500a <=( A199  and  (not A166) );
 a80503a <=( A201  and  (not A200) );
 a80504a <=( a80503a  and  a80500a );
 a80505a <=( a80504a  and  a80497a );
 a80508a <=( (not A265)  and  A202 );
 a80511a <=( (not A267)  and  A266 );
 a80512a <=( a80511a  and  a80508a );
 a80515a <=( (not A269)  and  (not A268) );
 a80518a <=( A299  and  A298 );
 a80519a <=( a80518a  and  a80515a );
 a80520a <=( a80519a  and  a80512a );
 a80524a <=( A167  and  A168 );
 a80525a <=( A169  and  a80524a );
 a80528a <=( A199  and  (not A166) );
 a80531a <=( A201  and  (not A200) );
 a80532a <=( a80531a  and  a80528a );
 a80533a <=( a80532a  and  a80525a );
 a80536a <=( (not A265)  and  A202 );
 a80539a <=( (not A267)  and  A266 );
 a80540a <=( a80539a  and  a80536a );
 a80543a <=( (not A269)  and  (not A268) );
 a80546a <=( (not A299)  and  (not A298) );
 a80547a <=( a80546a  and  a80543a );
 a80548a <=( a80547a  and  a80540a );
 a80552a <=( A167  and  A168 );
 a80553a <=( A169  and  a80552a );
 a80556a <=( A199  and  (not A166) );
 a80559a <=( A201  and  (not A200) );
 a80560a <=( a80559a  and  a80556a );
 a80561a <=( a80560a  and  a80553a );
 a80564a <=( A265  and  A202 );
 a80567a <=( A267  and  (not A266) );
 a80568a <=( a80567a  and  a80564a );
 a80571a <=( A300  and  A268 );
 a80574a <=( (not A302)  and  (not A301) );
 a80575a <=( a80574a  and  a80571a );
 a80576a <=( a80575a  and  a80568a );
 a80580a <=( A167  and  A168 );
 a80581a <=( A169  and  a80580a );
 a80584a <=( A199  and  (not A166) );
 a80587a <=( A201  and  (not A200) );
 a80588a <=( a80587a  and  a80584a );
 a80589a <=( a80588a  and  a80581a );
 a80592a <=( A265  and  A202 );
 a80595a <=( A267  and  (not A266) );
 a80596a <=( a80595a  and  a80592a );
 a80599a <=( A300  and  A269 );
 a80602a <=( (not A302)  and  (not A301) );
 a80603a <=( a80602a  and  a80599a );
 a80604a <=( a80603a  and  a80596a );
 a80608a <=( A167  and  A168 );
 a80609a <=( A169  and  a80608a );
 a80612a <=( A199  and  (not A166) );
 a80615a <=( A201  and  (not A200) );
 a80616a <=( a80615a  and  a80612a );
 a80617a <=( a80616a  and  a80609a );
 a80620a <=( A265  and  A202 );
 a80623a <=( (not A267)  and  (not A266) );
 a80624a <=( a80623a  and  a80620a );
 a80627a <=( (not A269)  and  (not A268) );
 a80630a <=( A301  and  (not A300) );
 a80631a <=( a80630a  and  a80627a );
 a80632a <=( a80631a  and  a80624a );
 a80636a <=( A167  and  A168 );
 a80637a <=( A169  and  a80636a );
 a80640a <=( A199  and  (not A166) );
 a80643a <=( A201  and  (not A200) );
 a80644a <=( a80643a  and  a80640a );
 a80645a <=( a80644a  and  a80637a );
 a80648a <=( A265  and  A202 );
 a80651a <=( (not A267)  and  (not A266) );
 a80652a <=( a80651a  and  a80648a );
 a80655a <=( (not A269)  and  (not A268) );
 a80658a <=( A302  and  (not A300) );
 a80659a <=( a80658a  and  a80655a );
 a80660a <=( a80659a  and  a80652a );
 a80664a <=( A167  and  A168 );
 a80665a <=( A169  and  a80664a );
 a80668a <=( A199  and  (not A166) );
 a80671a <=( A201  and  (not A200) );
 a80672a <=( a80671a  and  a80668a );
 a80673a <=( a80672a  and  a80665a );
 a80676a <=( A265  and  A202 );
 a80679a <=( (not A267)  and  (not A266) );
 a80680a <=( a80679a  and  a80676a );
 a80683a <=( (not A269)  and  (not A268) );
 a80686a <=( A299  and  A298 );
 a80687a <=( a80686a  and  a80683a );
 a80688a <=( a80687a  and  a80680a );
 a80692a <=( A167  and  A168 );
 a80693a <=( A169  and  a80692a );
 a80696a <=( A199  and  (not A166) );
 a80699a <=( A201  and  (not A200) );
 a80700a <=( a80699a  and  a80696a );
 a80701a <=( a80700a  and  a80693a );
 a80704a <=( A265  and  A202 );
 a80707a <=( (not A267)  and  (not A266) );
 a80708a <=( a80707a  and  a80704a );
 a80711a <=( (not A269)  and  (not A268) );
 a80714a <=( (not A299)  and  (not A298) );
 a80715a <=( a80714a  and  a80711a );
 a80716a <=( a80715a  and  a80708a );
 a80720a <=( A167  and  A168 );
 a80721a <=( A169  and  a80720a );
 a80724a <=( A199  and  (not A166) );
 a80727a <=( A201  and  (not A200) );
 a80728a <=( a80727a  and  a80724a );
 a80729a <=( a80728a  and  a80721a );
 a80732a <=( (not A265)  and  A203 );
 a80735a <=( A267  and  A266 );
 a80736a <=( a80735a  and  a80732a );
 a80739a <=( A300  and  A268 );
 a80742a <=( (not A302)  and  (not A301) );
 a80743a <=( a80742a  and  a80739a );
 a80744a <=( a80743a  and  a80736a );
 a80748a <=( A167  and  A168 );
 a80749a <=( A169  and  a80748a );
 a80752a <=( A199  and  (not A166) );
 a80755a <=( A201  and  (not A200) );
 a80756a <=( a80755a  and  a80752a );
 a80757a <=( a80756a  and  a80749a );
 a80760a <=( (not A265)  and  A203 );
 a80763a <=( A267  and  A266 );
 a80764a <=( a80763a  and  a80760a );
 a80767a <=( A300  and  A269 );
 a80770a <=( (not A302)  and  (not A301) );
 a80771a <=( a80770a  and  a80767a );
 a80772a <=( a80771a  and  a80764a );
 a80776a <=( A167  and  A168 );
 a80777a <=( A169  and  a80776a );
 a80780a <=( A199  and  (not A166) );
 a80783a <=( A201  and  (not A200) );
 a80784a <=( a80783a  and  a80780a );
 a80785a <=( a80784a  and  a80777a );
 a80788a <=( (not A265)  and  A203 );
 a80791a <=( (not A267)  and  A266 );
 a80792a <=( a80791a  and  a80788a );
 a80795a <=( (not A269)  and  (not A268) );
 a80798a <=( A301  and  (not A300) );
 a80799a <=( a80798a  and  a80795a );
 a80800a <=( a80799a  and  a80792a );
 a80804a <=( A167  and  A168 );
 a80805a <=( A169  and  a80804a );
 a80808a <=( A199  and  (not A166) );
 a80811a <=( A201  and  (not A200) );
 a80812a <=( a80811a  and  a80808a );
 a80813a <=( a80812a  and  a80805a );
 a80816a <=( (not A265)  and  A203 );
 a80819a <=( (not A267)  and  A266 );
 a80820a <=( a80819a  and  a80816a );
 a80823a <=( (not A269)  and  (not A268) );
 a80826a <=( A302  and  (not A300) );
 a80827a <=( a80826a  and  a80823a );
 a80828a <=( a80827a  and  a80820a );
 a80832a <=( A167  and  A168 );
 a80833a <=( A169  and  a80832a );
 a80836a <=( A199  and  (not A166) );
 a80839a <=( A201  and  (not A200) );
 a80840a <=( a80839a  and  a80836a );
 a80841a <=( a80840a  and  a80833a );
 a80844a <=( (not A265)  and  A203 );
 a80847a <=( (not A267)  and  A266 );
 a80848a <=( a80847a  and  a80844a );
 a80851a <=( (not A269)  and  (not A268) );
 a80854a <=( A299  and  A298 );
 a80855a <=( a80854a  and  a80851a );
 a80856a <=( a80855a  and  a80848a );
 a80860a <=( A167  and  A168 );
 a80861a <=( A169  and  a80860a );
 a80864a <=( A199  and  (not A166) );
 a80867a <=( A201  and  (not A200) );
 a80868a <=( a80867a  and  a80864a );
 a80869a <=( a80868a  and  a80861a );
 a80872a <=( (not A265)  and  A203 );
 a80875a <=( (not A267)  and  A266 );
 a80876a <=( a80875a  and  a80872a );
 a80879a <=( (not A269)  and  (not A268) );
 a80882a <=( (not A299)  and  (not A298) );
 a80883a <=( a80882a  and  a80879a );
 a80884a <=( a80883a  and  a80876a );
 a80888a <=( A167  and  A168 );
 a80889a <=( A169  and  a80888a );
 a80892a <=( A199  and  (not A166) );
 a80895a <=( A201  and  (not A200) );
 a80896a <=( a80895a  and  a80892a );
 a80897a <=( a80896a  and  a80889a );
 a80900a <=( A265  and  A203 );
 a80903a <=( A267  and  (not A266) );
 a80904a <=( a80903a  and  a80900a );
 a80907a <=( A300  and  A268 );
 a80910a <=( (not A302)  and  (not A301) );
 a80911a <=( a80910a  and  a80907a );
 a80912a <=( a80911a  and  a80904a );
 a80916a <=( A167  and  A168 );
 a80917a <=( A169  and  a80916a );
 a80920a <=( A199  and  (not A166) );
 a80923a <=( A201  and  (not A200) );
 a80924a <=( a80923a  and  a80920a );
 a80925a <=( a80924a  and  a80917a );
 a80928a <=( A265  and  A203 );
 a80931a <=( A267  and  (not A266) );
 a80932a <=( a80931a  and  a80928a );
 a80935a <=( A300  and  A269 );
 a80938a <=( (not A302)  and  (not A301) );
 a80939a <=( a80938a  and  a80935a );
 a80940a <=( a80939a  and  a80932a );
 a80944a <=( A167  and  A168 );
 a80945a <=( A169  and  a80944a );
 a80948a <=( A199  and  (not A166) );
 a80951a <=( A201  and  (not A200) );
 a80952a <=( a80951a  and  a80948a );
 a80953a <=( a80952a  and  a80945a );
 a80956a <=( A265  and  A203 );
 a80959a <=( (not A267)  and  (not A266) );
 a80960a <=( a80959a  and  a80956a );
 a80963a <=( (not A269)  and  (not A268) );
 a80966a <=( A301  and  (not A300) );
 a80967a <=( a80966a  and  a80963a );
 a80968a <=( a80967a  and  a80960a );
 a80972a <=( A167  and  A168 );
 a80973a <=( A169  and  a80972a );
 a80976a <=( A199  and  (not A166) );
 a80979a <=( A201  and  (not A200) );
 a80980a <=( a80979a  and  a80976a );
 a80981a <=( a80980a  and  a80973a );
 a80984a <=( A265  and  A203 );
 a80987a <=( (not A267)  and  (not A266) );
 a80988a <=( a80987a  and  a80984a );
 a80991a <=( (not A269)  and  (not A268) );
 a80994a <=( A302  and  (not A300) );
 a80995a <=( a80994a  and  a80991a );
 a80996a <=( a80995a  and  a80988a );
 a81000a <=( A167  and  A168 );
 a81001a <=( A169  and  a81000a );
 a81004a <=( A199  and  (not A166) );
 a81007a <=( A201  and  (not A200) );
 a81008a <=( a81007a  and  a81004a );
 a81009a <=( a81008a  and  a81001a );
 a81012a <=( A265  and  A203 );
 a81015a <=( (not A267)  and  (not A266) );
 a81016a <=( a81015a  and  a81012a );
 a81019a <=( (not A269)  and  (not A268) );
 a81022a <=( A299  and  A298 );
 a81023a <=( a81022a  and  a81019a );
 a81024a <=( a81023a  and  a81016a );
 a81028a <=( A167  and  A168 );
 a81029a <=( A169  and  a81028a );
 a81032a <=( A199  and  (not A166) );
 a81035a <=( A201  and  (not A200) );
 a81036a <=( a81035a  and  a81032a );
 a81037a <=( a81036a  and  a81029a );
 a81040a <=( A265  and  A203 );
 a81043a <=( (not A267)  and  (not A266) );
 a81044a <=( a81043a  and  a81040a );
 a81047a <=( (not A269)  and  (not A268) );
 a81050a <=( (not A299)  and  (not A298) );
 a81051a <=( a81050a  and  a81047a );
 a81052a <=( a81051a  and  a81044a );
 a81056a <=( A167  and  A168 );
 a81057a <=( A169  and  a81056a );
 a81060a <=( A199  and  (not A166) );
 a81063a <=( (not A201)  and  (not A200) );
 a81064a <=( a81063a  and  a81060a );
 a81065a <=( a81064a  and  a81057a );
 a81068a <=( (not A203)  and  (not A202) );
 a81071a <=( A266  and  (not A265) );
 a81072a <=( a81071a  and  a81068a );
 a81075a <=( A268  and  A267 );
 a81078a <=( A301  and  (not A300) );
 a81079a <=( a81078a  and  a81075a );
 a81080a <=( a81079a  and  a81072a );
 a81084a <=( A167  and  A168 );
 a81085a <=( A169  and  a81084a );
 a81088a <=( A199  and  (not A166) );
 a81091a <=( (not A201)  and  (not A200) );
 a81092a <=( a81091a  and  a81088a );
 a81093a <=( a81092a  and  a81085a );
 a81096a <=( (not A203)  and  (not A202) );
 a81099a <=( A266  and  (not A265) );
 a81100a <=( a81099a  and  a81096a );
 a81103a <=( A268  and  A267 );
 a81106a <=( A302  and  (not A300) );
 a81107a <=( a81106a  and  a81103a );
 a81108a <=( a81107a  and  a81100a );
 a81112a <=( A167  and  A168 );
 a81113a <=( A169  and  a81112a );
 a81116a <=( A199  and  (not A166) );
 a81119a <=( (not A201)  and  (not A200) );
 a81120a <=( a81119a  and  a81116a );
 a81121a <=( a81120a  and  a81113a );
 a81124a <=( (not A203)  and  (not A202) );
 a81127a <=( A266  and  (not A265) );
 a81128a <=( a81127a  and  a81124a );
 a81131a <=( A268  and  A267 );
 a81134a <=( A299  and  A298 );
 a81135a <=( a81134a  and  a81131a );
 a81136a <=( a81135a  and  a81128a );
 a81140a <=( A167  and  A168 );
 a81141a <=( A169  and  a81140a );
 a81144a <=( A199  and  (not A166) );
 a81147a <=( (not A201)  and  (not A200) );
 a81148a <=( a81147a  and  a81144a );
 a81149a <=( a81148a  and  a81141a );
 a81152a <=( (not A203)  and  (not A202) );
 a81155a <=( A266  and  (not A265) );
 a81156a <=( a81155a  and  a81152a );
 a81159a <=( A268  and  A267 );
 a81162a <=( (not A299)  and  (not A298) );
 a81163a <=( a81162a  and  a81159a );
 a81164a <=( a81163a  and  a81156a );
 a81168a <=( A167  and  A168 );
 a81169a <=( A169  and  a81168a );
 a81172a <=( A199  and  (not A166) );
 a81175a <=( (not A201)  and  (not A200) );
 a81176a <=( a81175a  and  a81172a );
 a81177a <=( a81176a  and  a81169a );
 a81180a <=( (not A203)  and  (not A202) );
 a81183a <=( A266  and  (not A265) );
 a81184a <=( a81183a  and  a81180a );
 a81187a <=( A269  and  A267 );
 a81190a <=( A301  and  (not A300) );
 a81191a <=( a81190a  and  a81187a );
 a81192a <=( a81191a  and  a81184a );
 a81196a <=( A167  and  A168 );
 a81197a <=( A169  and  a81196a );
 a81200a <=( A199  and  (not A166) );
 a81203a <=( (not A201)  and  (not A200) );
 a81204a <=( a81203a  and  a81200a );
 a81205a <=( a81204a  and  a81197a );
 a81208a <=( (not A203)  and  (not A202) );
 a81211a <=( A266  and  (not A265) );
 a81212a <=( a81211a  and  a81208a );
 a81215a <=( A269  and  A267 );
 a81218a <=( A302  and  (not A300) );
 a81219a <=( a81218a  and  a81215a );
 a81220a <=( a81219a  and  a81212a );
 a81224a <=( A167  and  A168 );
 a81225a <=( A169  and  a81224a );
 a81228a <=( A199  and  (not A166) );
 a81231a <=( (not A201)  and  (not A200) );
 a81232a <=( a81231a  and  a81228a );
 a81233a <=( a81232a  and  a81225a );
 a81236a <=( (not A203)  and  (not A202) );
 a81239a <=( A266  and  (not A265) );
 a81240a <=( a81239a  and  a81236a );
 a81243a <=( A269  and  A267 );
 a81246a <=( A299  and  A298 );
 a81247a <=( a81246a  and  a81243a );
 a81248a <=( a81247a  and  a81240a );
 a81252a <=( A167  and  A168 );
 a81253a <=( A169  and  a81252a );
 a81256a <=( A199  and  (not A166) );
 a81259a <=( (not A201)  and  (not A200) );
 a81260a <=( a81259a  and  a81256a );
 a81261a <=( a81260a  and  a81253a );
 a81264a <=( (not A203)  and  (not A202) );
 a81267a <=( A266  and  (not A265) );
 a81268a <=( a81267a  and  a81264a );
 a81271a <=( A269  and  A267 );
 a81274a <=( (not A299)  and  (not A298) );
 a81275a <=( a81274a  and  a81271a );
 a81276a <=( a81275a  and  a81268a );
 a81280a <=( A167  and  A168 );
 a81281a <=( A169  and  a81280a );
 a81284a <=( A199  and  (not A166) );
 a81287a <=( (not A201)  and  (not A200) );
 a81288a <=( a81287a  and  a81284a );
 a81289a <=( a81288a  and  a81281a );
 a81292a <=( (not A203)  and  (not A202) );
 a81295a <=( (not A266)  and  A265 );
 a81296a <=( a81295a  and  a81292a );
 a81299a <=( A268  and  A267 );
 a81302a <=( A301  and  (not A300) );
 a81303a <=( a81302a  and  a81299a );
 a81304a <=( a81303a  and  a81296a );
 a81308a <=( A167  and  A168 );
 a81309a <=( A169  and  a81308a );
 a81312a <=( A199  and  (not A166) );
 a81315a <=( (not A201)  and  (not A200) );
 a81316a <=( a81315a  and  a81312a );
 a81317a <=( a81316a  and  a81309a );
 a81320a <=( (not A203)  and  (not A202) );
 a81323a <=( (not A266)  and  A265 );
 a81324a <=( a81323a  and  a81320a );
 a81327a <=( A268  and  A267 );
 a81330a <=( A302  and  (not A300) );
 a81331a <=( a81330a  and  a81327a );
 a81332a <=( a81331a  and  a81324a );
 a81336a <=( A167  and  A168 );
 a81337a <=( A169  and  a81336a );
 a81340a <=( A199  and  (not A166) );
 a81343a <=( (not A201)  and  (not A200) );
 a81344a <=( a81343a  and  a81340a );
 a81345a <=( a81344a  and  a81337a );
 a81348a <=( (not A203)  and  (not A202) );
 a81351a <=( (not A266)  and  A265 );
 a81352a <=( a81351a  and  a81348a );
 a81355a <=( A268  and  A267 );
 a81358a <=( A299  and  A298 );
 a81359a <=( a81358a  and  a81355a );
 a81360a <=( a81359a  and  a81352a );
 a81364a <=( A167  and  A168 );
 a81365a <=( A169  and  a81364a );
 a81368a <=( A199  and  (not A166) );
 a81371a <=( (not A201)  and  (not A200) );
 a81372a <=( a81371a  and  a81368a );
 a81373a <=( a81372a  and  a81365a );
 a81376a <=( (not A203)  and  (not A202) );
 a81379a <=( (not A266)  and  A265 );
 a81380a <=( a81379a  and  a81376a );
 a81383a <=( A268  and  A267 );
 a81386a <=( (not A299)  and  (not A298) );
 a81387a <=( a81386a  and  a81383a );
 a81388a <=( a81387a  and  a81380a );
 a81392a <=( A167  and  A168 );
 a81393a <=( A169  and  a81392a );
 a81396a <=( A199  and  (not A166) );
 a81399a <=( (not A201)  and  (not A200) );
 a81400a <=( a81399a  and  a81396a );
 a81401a <=( a81400a  and  a81393a );
 a81404a <=( (not A203)  and  (not A202) );
 a81407a <=( (not A266)  and  A265 );
 a81408a <=( a81407a  and  a81404a );
 a81411a <=( A269  and  A267 );
 a81414a <=( A301  and  (not A300) );
 a81415a <=( a81414a  and  a81411a );
 a81416a <=( a81415a  and  a81408a );
 a81420a <=( A167  and  A168 );
 a81421a <=( A169  and  a81420a );
 a81424a <=( A199  and  (not A166) );
 a81427a <=( (not A201)  and  (not A200) );
 a81428a <=( a81427a  and  a81424a );
 a81429a <=( a81428a  and  a81421a );
 a81432a <=( (not A203)  and  (not A202) );
 a81435a <=( (not A266)  and  A265 );
 a81436a <=( a81435a  and  a81432a );
 a81439a <=( A269  and  A267 );
 a81442a <=( A302  and  (not A300) );
 a81443a <=( a81442a  and  a81439a );
 a81444a <=( a81443a  and  a81436a );
 a81448a <=( A167  and  A168 );
 a81449a <=( A169  and  a81448a );
 a81452a <=( A199  and  (not A166) );
 a81455a <=( (not A201)  and  (not A200) );
 a81456a <=( a81455a  and  a81452a );
 a81457a <=( a81456a  and  a81449a );
 a81460a <=( (not A203)  and  (not A202) );
 a81463a <=( (not A266)  and  A265 );
 a81464a <=( a81463a  and  a81460a );
 a81467a <=( A269  and  A267 );
 a81470a <=( A299  and  A298 );
 a81471a <=( a81470a  and  a81467a );
 a81472a <=( a81471a  and  a81464a );
 a81476a <=( A167  and  A168 );
 a81477a <=( A169  and  a81476a );
 a81480a <=( A199  and  (not A166) );
 a81483a <=( (not A201)  and  (not A200) );
 a81484a <=( a81483a  and  a81480a );
 a81485a <=( a81484a  and  a81477a );
 a81488a <=( (not A203)  and  (not A202) );
 a81491a <=( (not A266)  and  A265 );
 a81492a <=( a81491a  and  a81488a );
 a81495a <=( A269  and  A267 );
 a81498a <=( (not A299)  and  (not A298) );
 a81499a <=( a81498a  and  a81495a );
 a81500a <=( a81499a  and  a81492a );
 a81504a <=( (not A167)  and  A168 );
 a81505a <=( A169  and  a81504a );
 a81508a <=( A201  and  A166 );
 a81511a <=( (not A203)  and  (not A202) );
 a81512a <=( a81511a  and  a81508a );
 a81513a <=( a81512a  and  a81505a );
 a81516a <=( (not A268)  and  A267 );
 a81519a <=( A298  and  (not A269) );
 a81520a <=( a81519a  and  a81516a );
 a81523a <=( (not A300)  and  (not A299) );
 a81526a <=( (not A302)  and  (not A301) );
 a81527a <=( a81526a  and  a81523a );
 a81528a <=( a81527a  and  a81520a );
 a81532a <=( (not A167)  and  A168 );
 a81533a <=( A169  and  a81532a );
 a81536a <=( A201  and  A166 );
 a81539a <=( (not A203)  and  (not A202) );
 a81540a <=( a81539a  and  a81536a );
 a81541a <=( a81540a  and  a81533a );
 a81544a <=( (not A268)  and  A267 );
 a81547a <=( (not A298)  and  (not A269) );
 a81548a <=( a81547a  and  a81544a );
 a81551a <=( (not A300)  and  A299 );
 a81554a <=( (not A302)  and  (not A301) );
 a81555a <=( a81554a  and  a81551a );
 a81556a <=( a81555a  and  a81548a );
 a81560a <=( (not A167)  and  A168 );
 a81561a <=( A169  and  a81560a );
 a81564a <=( (not A199)  and  A166 );
 a81567a <=( A201  and  A200 );
 a81568a <=( a81567a  and  a81564a );
 a81569a <=( a81568a  and  a81561a );
 a81572a <=( (not A265)  and  A202 );
 a81575a <=( A267  and  A266 );
 a81576a <=( a81575a  and  a81572a );
 a81579a <=( A300  and  A268 );
 a81582a <=( (not A302)  and  (not A301) );
 a81583a <=( a81582a  and  a81579a );
 a81584a <=( a81583a  and  a81576a );
 a81588a <=( (not A167)  and  A168 );
 a81589a <=( A169  and  a81588a );
 a81592a <=( (not A199)  and  A166 );
 a81595a <=( A201  and  A200 );
 a81596a <=( a81595a  and  a81592a );
 a81597a <=( a81596a  and  a81589a );
 a81600a <=( (not A265)  and  A202 );
 a81603a <=( A267  and  A266 );
 a81604a <=( a81603a  and  a81600a );
 a81607a <=( A300  and  A269 );
 a81610a <=( (not A302)  and  (not A301) );
 a81611a <=( a81610a  and  a81607a );
 a81612a <=( a81611a  and  a81604a );
 a81616a <=( (not A167)  and  A168 );
 a81617a <=( A169  and  a81616a );
 a81620a <=( (not A199)  and  A166 );
 a81623a <=( A201  and  A200 );
 a81624a <=( a81623a  and  a81620a );
 a81625a <=( a81624a  and  a81617a );
 a81628a <=( (not A265)  and  A202 );
 a81631a <=( (not A267)  and  A266 );
 a81632a <=( a81631a  and  a81628a );
 a81635a <=( (not A269)  and  (not A268) );
 a81638a <=( A301  and  (not A300) );
 a81639a <=( a81638a  and  a81635a );
 a81640a <=( a81639a  and  a81632a );
 a81644a <=( (not A167)  and  A168 );
 a81645a <=( A169  and  a81644a );
 a81648a <=( (not A199)  and  A166 );
 a81651a <=( A201  and  A200 );
 a81652a <=( a81651a  and  a81648a );
 a81653a <=( a81652a  and  a81645a );
 a81656a <=( (not A265)  and  A202 );
 a81659a <=( (not A267)  and  A266 );
 a81660a <=( a81659a  and  a81656a );
 a81663a <=( (not A269)  and  (not A268) );
 a81666a <=( A302  and  (not A300) );
 a81667a <=( a81666a  and  a81663a );
 a81668a <=( a81667a  and  a81660a );
 a81672a <=( (not A167)  and  A168 );
 a81673a <=( A169  and  a81672a );
 a81676a <=( (not A199)  and  A166 );
 a81679a <=( A201  and  A200 );
 a81680a <=( a81679a  and  a81676a );
 a81681a <=( a81680a  and  a81673a );
 a81684a <=( (not A265)  and  A202 );
 a81687a <=( (not A267)  and  A266 );
 a81688a <=( a81687a  and  a81684a );
 a81691a <=( (not A269)  and  (not A268) );
 a81694a <=( A299  and  A298 );
 a81695a <=( a81694a  and  a81691a );
 a81696a <=( a81695a  and  a81688a );
 a81700a <=( (not A167)  and  A168 );
 a81701a <=( A169  and  a81700a );
 a81704a <=( (not A199)  and  A166 );
 a81707a <=( A201  and  A200 );
 a81708a <=( a81707a  and  a81704a );
 a81709a <=( a81708a  and  a81701a );
 a81712a <=( (not A265)  and  A202 );
 a81715a <=( (not A267)  and  A266 );
 a81716a <=( a81715a  and  a81712a );
 a81719a <=( (not A269)  and  (not A268) );
 a81722a <=( (not A299)  and  (not A298) );
 a81723a <=( a81722a  and  a81719a );
 a81724a <=( a81723a  and  a81716a );
 a81728a <=( (not A167)  and  A168 );
 a81729a <=( A169  and  a81728a );
 a81732a <=( (not A199)  and  A166 );
 a81735a <=( A201  and  A200 );
 a81736a <=( a81735a  and  a81732a );
 a81737a <=( a81736a  and  a81729a );
 a81740a <=( A265  and  A202 );
 a81743a <=( A267  and  (not A266) );
 a81744a <=( a81743a  and  a81740a );
 a81747a <=( A300  and  A268 );
 a81750a <=( (not A302)  and  (not A301) );
 a81751a <=( a81750a  and  a81747a );
 a81752a <=( a81751a  and  a81744a );
 a81756a <=( (not A167)  and  A168 );
 a81757a <=( A169  and  a81756a );
 a81760a <=( (not A199)  and  A166 );
 a81763a <=( A201  and  A200 );
 a81764a <=( a81763a  and  a81760a );
 a81765a <=( a81764a  and  a81757a );
 a81768a <=( A265  and  A202 );
 a81771a <=( A267  and  (not A266) );
 a81772a <=( a81771a  and  a81768a );
 a81775a <=( A300  and  A269 );
 a81778a <=( (not A302)  and  (not A301) );
 a81779a <=( a81778a  and  a81775a );
 a81780a <=( a81779a  and  a81772a );
 a81784a <=( (not A167)  and  A168 );
 a81785a <=( A169  and  a81784a );
 a81788a <=( (not A199)  and  A166 );
 a81791a <=( A201  and  A200 );
 a81792a <=( a81791a  and  a81788a );
 a81793a <=( a81792a  and  a81785a );
 a81796a <=( A265  and  A202 );
 a81799a <=( (not A267)  and  (not A266) );
 a81800a <=( a81799a  and  a81796a );
 a81803a <=( (not A269)  and  (not A268) );
 a81806a <=( A301  and  (not A300) );
 a81807a <=( a81806a  and  a81803a );
 a81808a <=( a81807a  and  a81800a );
 a81812a <=( (not A167)  and  A168 );
 a81813a <=( A169  and  a81812a );
 a81816a <=( (not A199)  and  A166 );
 a81819a <=( A201  and  A200 );
 a81820a <=( a81819a  and  a81816a );
 a81821a <=( a81820a  and  a81813a );
 a81824a <=( A265  and  A202 );
 a81827a <=( (not A267)  and  (not A266) );
 a81828a <=( a81827a  and  a81824a );
 a81831a <=( (not A269)  and  (not A268) );
 a81834a <=( A302  and  (not A300) );
 a81835a <=( a81834a  and  a81831a );
 a81836a <=( a81835a  and  a81828a );
 a81840a <=( (not A167)  and  A168 );
 a81841a <=( A169  and  a81840a );
 a81844a <=( (not A199)  and  A166 );
 a81847a <=( A201  and  A200 );
 a81848a <=( a81847a  and  a81844a );
 a81849a <=( a81848a  and  a81841a );
 a81852a <=( A265  and  A202 );
 a81855a <=( (not A267)  and  (not A266) );
 a81856a <=( a81855a  and  a81852a );
 a81859a <=( (not A269)  and  (not A268) );
 a81862a <=( A299  and  A298 );
 a81863a <=( a81862a  and  a81859a );
 a81864a <=( a81863a  and  a81856a );
 a81868a <=( (not A167)  and  A168 );
 a81869a <=( A169  and  a81868a );
 a81872a <=( (not A199)  and  A166 );
 a81875a <=( A201  and  A200 );
 a81876a <=( a81875a  and  a81872a );
 a81877a <=( a81876a  and  a81869a );
 a81880a <=( A265  and  A202 );
 a81883a <=( (not A267)  and  (not A266) );
 a81884a <=( a81883a  and  a81880a );
 a81887a <=( (not A269)  and  (not A268) );
 a81890a <=( (not A299)  and  (not A298) );
 a81891a <=( a81890a  and  a81887a );
 a81892a <=( a81891a  and  a81884a );
 a81896a <=( (not A167)  and  A168 );
 a81897a <=( A169  and  a81896a );
 a81900a <=( (not A199)  and  A166 );
 a81903a <=( A201  and  A200 );
 a81904a <=( a81903a  and  a81900a );
 a81905a <=( a81904a  and  a81897a );
 a81908a <=( (not A265)  and  A203 );
 a81911a <=( A267  and  A266 );
 a81912a <=( a81911a  and  a81908a );
 a81915a <=( A300  and  A268 );
 a81918a <=( (not A302)  and  (not A301) );
 a81919a <=( a81918a  and  a81915a );
 a81920a <=( a81919a  and  a81912a );
 a81924a <=( (not A167)  and  A168 );
 a81925a <=( A169  and  a81924a );
 a81928a <=( (not A199)  and  A166 );
 a81931a <=( A201  and  A200 );
 a81932a <=( a81931a  and  a81928a );
 a81933a <=( a81932a  and  a81925a );
 a81936a <=( (not A265)  and  A203 );
 a81939a <=( A267  and  A266 );
 a81940a <=( a81939a  and  a81936a );
 a81943a <=( A300  and  A269 );
 a81946a <=( (not A302)  and  (not A301) );
 a81947a <=( a81946a  and  a81943a );
 a81948a <=( a81947a  and  a81940a );
 a81952a <=( (not A167)  and  A168 );
 a81953a <=( A169  and  a81952a );
 a81956a <=( (not A199)  and  A166 );
 a81959a <=( A201  and  A200 );
 a81960a <=( a81959a  and  a81956a );
 a81961a <=( a81960a  and  a81953a );
 a81964a <=( (not A265)  and  A203 );
 a81967a <=( (not A267)  and  A266 );
 a81968a <=( a81967a  and  a81964a );
 a81971a <=( (not A269)  and  (not A268) );
 a81974a <=( A301  and  (not A300) );
 a81975a <=( a81974a  and  a81971a );
 a81976a <=( a81975a  and  a81968a );
 a81980a <=( (not A167)  and  A168 );
 a81981a <=( A169  and  a81980a );
 a81984a <=( (not A199)  and  A166 );
 a81987a <=( A201  and  A200 );
 a81988a <=( a81987a  and  a81984a );
 a81989a <=( a81988a  and  a81981a );
 a81992a <=( (not A265)  and  A203 );
 a81995a <=( (not A267)  and  A266 );
 a81996a <=( a81995a  and  a81992a );
 a81999a <=( (not A269)  and  (not A268) );
 a82002a <=( A302  and  (not A300) );
 a82003a <=( a82002a  and  a81999a );
 a82004a <=( a82003a  and  a81996a );
 a82008a <=( (not A167)  and  A168 );
 a82009a <=( A169  and  a82008a );
 a82012a <=( (not A199)  and  A166 );
 a82015a <=( A201  and  A200 );
 a82016a <=( a82015a  and  a82012a );
 a82017a <=( a82016a  and  a82009a );
 a82020a <=( (not A265)  and  A203 );
 a82023a <=( (not A267)  and  A266 );
 a82024a <=( a82023a  and  a82020a );
 a82027a <=( (not A269)  and  (not A268) );
 a82030a <=( A299  and  A298 );
 a82031a <=( a82030a  and  a82027a );
 a82032a <=( a82031a  and  a82024a );
 a82036a <=( (not A167)  and  A168 );
 a82037a <=( A169  and  a82036a );
 a82040a <=( (not A199)  and  A166 );
 a82043a <=( A201  and  A200 );
 a82044a <=( a82043a  and  a82040a );
 a82045a <=( a82044a  and  a82037a );
 a82048a <=( (not A265)  and  A203 );
 a82051a <=( (not A267)  and  A266 );
 a82052a <=( a82051a  and  a82048a );
 a82055a <=( (not A269)  and  (not A268) );
 a82058a <=( (not A299)  and  (not A298) );
 a82059a <=( a82058a  and  a82055a );
 a82060a <=( a82059a  and  a82052a );
 a82064a <=( (not A167)  and  A168 );
 a82065a <=( A169  and  a82064a );
 a82068a <=( (not A199)  and  A166 );
 a82071a <=( A201  and  A200 );
 a82072a <=( a82071a  and  a82068a );
 a82073a <=( a82072a  and  a82065a );
 a82076a <=( A265  and  A203 );
 a82079a <=( A267  and  (not A266) );
 a82080a <=( a82079a  and  a82076a );
 a82083a <=( A300  and  A268 );
 a82086a <=( (not A302)  and  (not A301) );
 a82087a <=( a82086a  and  a82083a );
 a82088a <=( a82087a  and  a82080a );
 a82092a <=( (not A167)  and  A168 );
 a82093a <=( A169  and  a82092a );
 a82096a <=( (not A199)  and  A166 );
 a82099a <=( A201  and  A200 );
 a82100a <=( a82099a  and  a82096a );
 a82101a <=( a82100a  and  a82093a );
 a82104a <=( A265  and  A203 );
 a82107a <=( A267  and  (not A266) );
 a82108a <=( a82107a  and  a82104a );
 a82111a <=( A300  and  A269 );
 a82114a <=( (not A302)  and  (not A301) );
 a82115a <=( a82114a  and  a82111a );
 a82116a <=( a82115a  and  a82108a );
 a82120a <=( (not A167)  and  A168 );
 a82121a <=( A169  and  a82120a );
 a82124a <=( (not A199)  and  A166 );
 a82127a <=( A201  and  A200 );
 a82128a <=( a82127a  and  a82124a );
 a82129a <=( a82128a  and  a82121a );
 a82132a <=( A265  and  A203 );
 a82135a <=( (not A267)  and  (not A266) );
 a82136a <=( a82135a  and  a82132a );
 a82139a <=( (not A269)  and  (not A268) );
 a82142a <=( A301  and  (not A300) );
 a82143a <=( a82142a  and  a82139a );
 a82144a <=( a82143a  and  a82136a );
 a82148a <=( (not A167)  and  A168 );
 a82149a <=( A169  and  a82148a );
 a82152a <=( (not A199)  and  A166 );
 a82155a <=( A201  and  A200 );
 a82156a <=( a82155a  and  a82152a );
 a82157a <=( a82156a  and  a82149a );
 a82160a <=( A265  and  A203 );
 a82163a <=( (not A267)  and  (not A266) );
 a82164a <=( a82163a  and  a82160a );
 a82167a <=( (not A269)  and  (not A268) );
 a82170a <=( A302  and  (not A300) );
 a82171a <=( a82170a  and  a82167a );
 a82172a <=( a82171a  and  a82164a );
 a82176a <=( (not A167)  and  A168 );
 a82177a <=( A169  and  a82176a );
 a82180a <=( (not A199)  and  A166 );
 a82183a <=( A201  and  A200 );
 a82184a <=( a82183a  and  a82180a );
 a82185a <=( a82184a  and  a82177a );
 a82188a <=( A265  and  A203 );
 a82191a <=( (not A267)  and  (not A266) );
 a82192a <=( a82191a  and  a82188a );
 a82195a <=( (not A269)  and  (not A268) );
 a82198a <=( A299  and  A298 );
 a82199a <=( a82198a  and  a82195a );
 a82200a <=( a82199a  and  a82192a );
 a82204a <=( (not A167)  and  A168 );
 a82205a <=( A169  and  a82204a );
 a82208a <=( (not A199)  and  A166 );
 a82211a <=( A201  and  A200 );
 a82212a <=( a82211a  and  a82208a );
 a82213a <=( a82212a  and  a82205a );
 a82216a <=( A265  and  A203 );
 a82219a <=( (not A267)  and  (not A266) );
 a82220a <=( a82219a  and  a82216a );
 a82223a <=( (not A269)  and  (not A268) );
 a82226a <=( (not A299)  and  (not A298) );
 a82227a <=( a82226a  and  a82223a );
 a82228a <=( a82227a  and  a82220a );
 a82232a <=( (not A167)  and  A168 );
 a82233a <=( A169  and  a82232a );
 a82236a <=( (not A199)  and  A166 );
 a82239a <=( (not A201)  and  A200 );
 a82240a <=( a82239a  and  a82236a );
 a82241a <=( a82240a  and  a82233a );
 a82244a <=( (not A203)  and  (not A202) );
 a82247a <=( A266  and  (not A265) );
 a82248a <=( a82247a  and  a82244a );
 a82251a <=( A268  and  A267 );
 a82254a <=( A301  and  (not A300) );
 a82255a <=( a82254a  and  a82251a );
 a82256a <=( a82255a  and  a82248a );
 a82260a <=( (not A167)  and  A168 );
 a82261a <=( A169  and  a82260a );
 a82264a <=( (not A199)  and  A166 );
 a82267a <=( (not A201)  and  A200 );
 a82268a <=( a82267a  and  a82264a );
 a82269a <=( a82268a  and  a82261a );
 a82272a <=( (not A203)  and  (not A202) );
 a82275a <=( A266  and  (not A265) );
 a82276a <=( a82275a  and  a82272a );
 a82279a <=( A268  and  A267 );
 a82282a <=( A302  and  (not A300) );
 a82283a <=( a82282a  and  a82279a );
 a82284a <=( a82283a  and  a82276a );
 a82288a <=( (not A167)  and  A168 );
 a82289a <=( A169  and  a82288a );
 a82292a <=( (not A199)  and  A166 );
 a82295a <=( (not A201)  and  A200 );
 a82296a <=( a82295a  and  a82292a );
 a82297a <=( a82296a  and  a82289a );
 a82300a <=( (not A203)  and  (not A202) );
 a82303a <=( A266  and  (not A265) );
 a82304a <=( a82303a  and  a82300a );
 a82307a <=( A268  and  A267 );
 a82310a <=( A299  and  A298 );
 a82311a <=( a82310a  and  a82307a );
 a82312a <=( a82311a  and  a82304a );
 a82316a <=( (not A167)  and  A168 );
 a82317a <=( A169  and  a82316a );
 a82320a <=( (not A199)  and  A166 );
 a82323a <=( (not A201)  and  A200 );
 a82324a <=( a82323a  and  a82320a );
 a82325a <=( a82324a  and  a82317a );
 a82328a <=( (not A203)  and  (not A202) );
 a82331a <=( A266  and  (not A265) );
 a82332a <=( a82331a  and  a82328a );
 a82335a <=( A268  and  A267 );
 a82338a <=( (not A299)  and  (not A298) );
 a82339a <=( a82338a  and  a82335a );
 a82340a <=( a82339a  and  a82332a );
 a82344a <=( (not A167)  and  A168 );
 a82345a <=( A169  and  a82344a );
 a82348a <=( (not A199)  and  A166 );
 a82351a <=( (not A201)  and  A200 );
 a82352a <=( a82351a  and  a82348a );
 a82353a <=( a82352a  and  a82345a );
 a82356a <=( (not A203)  and  (not A202) );
 a82359a <=( A266  and  (not A265) );
 a82360a <=( a82359a  and  a82356a );
 a82363a <=( A269  and  A267 );
 a82366a <=( A301  and  (not A300) );
 a82367a <=( a82366a  and  a82363a );
 a82368a <=( a82367a  and  a82360a );
 a82372a <=( (not A167)  and  A168 );
 a82373a <=( A169  and  a82372a );
 a82376a <=( (not A199)  and  A166 );
 a82379a <=( (not A201)  and  A200 );
 a82380a <=( a82379a  and  a82376a );
 a82381a <=( a82380a  and  a82373a );
 a82384a <=( (not A203)  and  (not A202) );
 a82387a <=( A266  and  (not A265) );
 a82388a <=( a82387a  and  a82384a );
 a82391a <=( A269  and  A267 );
 a82394a <=( A302  and  (not A300) );
 a82395a <=( a82394a  and  a82391a );
 a82396a <=( a82395a  and  a82388a );
 a82400a <=( (not A167)  and  A168 );
 a82401a <=( A169  and  a82400a );
 a82404a <=( (not A199)  and  A166 );
 a82407a <=( (not A201)  and  A200 );
 a82408a <=( a82407a  and  a82404a );
 a82409a <=( a82408a  and  a82401a );
 a82412a <=( (not A203)  and  (not A202) );
 a82415a <=( A266  and  (not A265) );
 a82416a <=( a82415a  and  a82412a );
 a82419a <=( A269  and  A267 );
 a82422a <=( A299  and  A298 );
 a82423a <=( a82422a  and  a82419a );
 a82424a <=( a82423a  and  a82416a );
 a82428a <=( (not A167)  and  A168 );
 a82429a <=( A169  and  a82428a );
 a82432a <=( (not A199)  and  A166 );
 a82435a <=( (not A201)  and  A200 );
 a82436a <=( a82435a  and  a82432a );
 a82437a <=( a82436a  and  a82429a );
 a82440a <=( (not A203)  and  (not A202) );
 a82443a <=( A266  and  (not A265) );
 a82444a <=( a82443a  and  a82440a );
 a82447a <=( A269  and  A267 );
 a82450a <=( (not A299)  and  (not A298) );
 a82451a <=( a82450a  and  a82447a );
 a82452a <=( a82451a  and  a82444a );
 a82456a <=( (not A167)  and  A168 );
 a82457a <=( A169  and  a82456a );
 a82460a <=( (not A199)  and  A166 );
 a82463a <=( (not A201)  and  A200 );
 a82464a <=( a82463a  and  a82460a );
 a82465a <=( a82464a  and  a82457a );
 a82468a <=( (not A203)  and  (not A202) );
 a82471a <=( (not A266)  and  A265 );
 a82472a <=( a82471a  and  a82468a );
 a82475a <=( A268  and  A267 );
 a82478a <=( A301  and  (not A300) );
 a82479a <=( a82478a  and  a82475a );
 a82480a <=( a82479a  and  a82472a );
 a82484a <=( (not A167)  and  A168 );
 a82485a <=( A169  and  a82484a );
 a82488a <=( (not A199)  and  A166 );
 a82491a <=( (not A201)  and  A200 );
 a82492a <=( a82491a  and  a82488a );
 a82493a <=( a82492a  and  a82485a );
 a82496a <=( (not A203)  and  (not A202) );
 a82499a <=( (not A266)  and  A265 );
 a82500a <=( a82499a  and  a82496a );
 a82503a <=( A268  and  A267 );
 a82506a <=( A302  and  (not A300) );
 a82507a <=( a82506a  and  a82503a );
 a82508a <=( a82507a  and  a82500a );
 a82512a <=( (not A167)  and  A168 );
 a82513a <=( A169  and  a82512a );
 a82516a <=( (not A199)  and  A166 );
 a82519a <=( (not A201)  and  A200 );
 a82520a <=( a82519a  and  a82516a );
 a82521a <=( a82520a  and  a82513a );
 a82524a <=( (not A203)  and  (not A202) );
 a82527a <=( (not A266)  and  A265 );
 a82528a <=( a82527a  and  a82524a );
 a82531a <=( A268  and  A267 );
 a82534a <=( A299  and  A298 );
 a82535a <=( a82534a  and  a82531a );
 a82536a <=( a82535a  and  a82528a );
 a82540a <=( (not A167)  and  A168 );
 a82541a <=( A169  and  a82540a );
 a82544a <=( (not A199)  and  A166 );
 a82547a <=( (not A201)  and  A200 );
 a82548a <=( a82547a  and  a82544a );
 a82549a <=( a82548a  and  a82541a );
 a82552a <=( (not A203)  and  (not A202) );
 a82555a <=( (not A266)  and  A265 );
 a82556a <=( a82555a  and  a82552a );
 a82559a <=( A268  and  A267 );
 a82562a <=( (not A299)  and  (not A298) );
 a82563a <=( a82562a  and  a82559a );
 a82564a <=( a82563a  and  a82556a );
 a82568a <=( (not A167)  and  A168 );
 a82569a <=( A169  and  a82568a );
 a82572a <=( (not A199)  and  A166 );
 a82575a <=( (not A201)  and  A200 );
 a82576a <=( a82575a  and  a82572a );
 a82577a <=( a82576a  and  a82569a );
 a82580a <=( (not A203)  and  (not A202) );
 a82583a <=( (not A266)  and  A265 );
 a82584a <=( a82583a  and  a82580a );
 a82587a <=( A269  and  A267 );
 a82590a <=( A301  and  (not A300) );
 a82591a <=( a82590a  and  a82587a );
 a82592a <=( a82591a  and  a82584a );
 a82596a <=( (not A167)  and  A168 );
 a82597a <=( A169  and  a82596a );
 a82600a <=( (not A199)  and  A166 );
 a82603a <=( (not A201)  and  A200 );
 a82604a <=( a82603a  and  a82600a );
 a82605a <=( a82604a  and  a82597a );
 a82608a <=( (not A203)  and  (not A202) );
 a82611a <=( (not A266)  and  A265 );
 a82612a <=( a82611a  and  a82608a );
 a82615a <=( A269  and  A267 );
 a82618a <=( A302  and  (not A300) );
 a82619a <=( a82618a  and  a82615a );
 a82620a <=( a82619a  and  a82612a );
 a82624a <=( (not A167)  and  A168 );
 a82625a <=( A169  and  a82624a );
 a82628a <=( (not A199)  and  A166 );
 a82631a <=( (not A201)  and  A200 );
 a82632a <=( a82631a  and  a82628a );
 a82633a <=( a82632a  and  a82625a );
 a82636a <=( (not A203)  and  (not A202) );
 a82639a <=( (not A266)  and  A265 );
 a82640a <=( a82639a  and  a82636a );
 a82643a <=( A269  and  A267 );
 a82646a <=( A299  and  A298 );
 a82647a <=( a82646a  and  a82643a );
 a82648a <=( a82647a  and  a82640a );
 a82652a <=( (not A167)  and  A168 );
 a82653a <=( A169  and  a82652a );
 a82656a <=( (not A199)  and  A166 );
 a82659a <=( (not A201)  and  A200 );
 a82660a <=( a82659a  and  a82656a );
 a82661a <=( a82660a  and  a82653a );
 a82664a <=( (not A203)  and  (not A202) );
 a82667a <=( (not A266)  and  A265 );
 a82668a <=( a82667a  and  a82664a );
 a82671a <=( A269  and  A267 );
 a82674a <=( (not A299)  and  (not A298) );
 a82675a <=( a82674a  and  a82671a );
 a82676a <=( a82675a  and  a82668a );
 a82680a <=( (not A167)  and  A168 );
 a82681a <=( A169  and  a82680a );
 a82684a <=( A199  and  A166 );
 a82687a <=( A201  and  (not A200) );
 a82688a <=( a82687a  and  a82684a );
 a82689a <=( a82688a  and  a82681a );
 a82692a <=( (not A265)  and  A202 );
 a82695a <=( A267  and  A266 );
 a82696a <=( a82695a  and  a82692a );
 a82699a <=( A300  and  A268 );
 a82702a <=( (not A302)  and  (not A301) );
 a82703a <=( a82702a  and  a82699a );
 a82704a <=( a82703a  and  a82696a );
 a82708a <=( (not A167)  and  A168 );
 a82709a <=( A169  and  a82708a );
 a82712a <=( A199  and  A166 );
 a82715a <=( A201  and  (not A200) );
 a82716a <=( a82715a  and  a82712a );
 a82717a <=( a82716a  and  a82709a );
 a82720a <=( (not A265)  and  A202 );
 a82723a <=( A267  and  A266 );
 a82724a <=( a82723a  and  a82720a );
 a82727a <=( A300  and  A269 );
 a82730a <=( (not A302)  and  (not A301) );
 a82731a <=( a82730a  and  a82727a );
 a82732a <=( a82731a  and  a82724a );
 a82736a <=( (not A167)  and  A168 );
 a82737a <=( A169  and  a82736a );
 a82740a <=( A199  and  A166 );
 a82743a <=( A201  and  (not A200) );
 a82744a <=( a82743a  and  a82740a );
 a82745a <=( a82744a  and  a82737a );
 a82748a <=( (not A265)  and  A202 );
 a82751a <=( (not A267)  and  A266 );
 a82752a <=( a82751a  and  a82748a );
 a82755a <=( (not A269)  and  (not A268) );
 a82758a <=( A301  and  (not A300) );
 a82759a <=( a82758a  and  a82755a );
 a82760a <=( a82759a  and  a82752a );
 a82764a <=( (not A167)  and  A168 );
 a82765a <=( A169  and  a82764a );
 a82768a <=( A199  and  A166 );
 a82771a <=( A201  and  (not A200) );
 a82772a <=( a82771a  and  a82768a );
 a82773a <=( a82772a  and  a82765a );
 a82776a <=( (not A265)  and  A202 );
 a82779a <=( (not A267)  and  A266 );
 a82780a <=( a82779a  and  a82776a );
 a82783a <=( (not A269)  and  (not A268) );
 a82786a <=( A302  and  (not A300) );
 a82787a <=( a82786a  and  a82783a );
 a82788a <=( a82787a  and  a82780a );
 a82792a <=( (not A167)  and  A168 );
 a82793a <=( A169  and  a82792a );
 a82796a <=( A199  and  A166 );
 a82799a <=( A201  and  (not A200) );
 a82800a <=( a82799a  and  a82796a );
 a82801a <=( a82800a  and  a82793a );
 a82804a <=( (not A265)  and  A202 );
 a82807a <=( (not A267)  and  A266 );
 a82808a <=( a82807a  and  a82804a );
 a82811a <=( (not A269)  and  (not A268) );
 a82814a <=( A299  and  A298 );
 a82815a <=( a82814a  and  a82811a );
 a82816a <=( a82815a  and  a82808a );
 a82820a <=( (not A167)  and  A168 );
 a82821a <=( A169  and  a82820a );
 a82824a <=( A199  and  A166 );
 a82827a <=( A201  and  (not A200) );
 a82828a <=( a82827a  and  a82824a );
 a82829a <=( a82828a  and  a82821a );
 a82832a <=( (not A265)  and  A202 );
 a82835a <=( (not A267)  and  A266 );
 a82836a <=( a82835a  and  a82832a );
 a82839a <=( (not A269)  and  (not A268) );
 a82842a <=( (not A299)  and  (not A298) );
 a82843a <=( a82842a  and  a82839a );
 a82844a <=( a82843a  and  a82836a );
 a82848a <=( (not A167)  and  A168 );
 a82849a <=( A169  and  a82848a );
 a82852a <=( A199  and  A166 );
 a82855a <=( A201  and  (not A200) );
 a82856a <=( a82855a  and  a82852a );
 a82857a <=( a82856a  and  a82849a );
 a82860a <=( A265  and  A202 );
 a82863a <=( A267  and  (not A266) );
 a82864a <=( a82863a  and  a82860a );
 a82867a <=( A300  and  A268 );
 a82870a <=( (not A302)  and  (not A301) );
 a82871a <=( a82870a  and  a82867a );
 a82872a <=( a82871a  and  a82864a );
 a82876a <=( (not A167)  and  A168 );
 a82877a <=( A169  and  a82876a );
 a82880a <=( A199  and  A166 );
 a82883a <=( A201  and  (not A200) );
 a82884a <=( a82883a  and  a82880a );
 a82885a <=( a82884a  and  a82877a );
 a82888a <=( A265  and  A202 );
 a82891a <=( A267  and  (not A266) );
 a82892a <=( a82891a  and  a82888a );
 a82895a <=( A300  and  A269 );
 a82898a <=( (not A302)  and  (not A301) );
 a82899a <=( a82898a  and  a82895a );
 a82900a <=( a82899a  and  a82892a );
 a82904a <=( (not A167)  and  A168 );
 a82905a <=( A169  and  a82904a );
 a82908a <=( A199  and  A166 );
 a82911a <=( A201  and  (not A200) );
 a82912a <=( a82911a  and  a82908a );
 a82913a <=( a82912a  and  a82905a );
 a82916a <=( A265  and  A202 );
 a82919a <=( (not A267)  and  (not A266) );
 a82920a <=( a82919a  and  a82916a );
 a82923a <=( (not A269)  and  (not A268) );
 a82926a <=( A301  and  (not A300) );
 a82927a <=( a82926a  and  a82923a );
 a82928a <=( a82927a  and  a82920a );
 a82932a <=( (not A167)  and  A168 );
 a82933a <=( A169  and  a82932a );
 a82936a <=( A199  and  A166 );
 a82939a <=( A201  and  (not A200) );
 a82940a <=( a82939a  and  a82936a );
 a82941a <=( a82940a  and  a82933a );
 a82944a <=( A265  and  A202 );
 a82947a <=( (not A267)  and  (not A266) );
 a82948a <=( a82947a  and  a82944a );
 a82951a <=( (not A269)  and  (not A268) );
 a82954a <=( A302  and  (not A300) );
 a82955a <=( a82954a  and  a82951a );
 a82956a <=( a82955a  and  a82948a );
 a82960a <=( (not A167)  and  A168 );
 a82961a <=( A169  and  a82960a );
 a82964a <=( A199  and  A166 );
 a82967a <=( A201  and  (not A200) );
 a82968a <=( a82967a  and  a82964a );
 a82969a <=( a82968a  and  a82961a );
 a82972a <=( A265  and  A202 );
 a82975a <=( (not A267)  and  (not A266) );
 a82976a <=( a82975a  and  a82972a );
 a82979a <=( (not A269)  and  (not A268) );
 a82982a <=( A299  and  A298 );
 a82983a <=( a82982a  and  a82979a );
 a82984a <=( a82983a  and  a82976a );
 a82988a <=( (not A167)  and  A168 );
 a82989a <=( A169  and  a82988a );
 a82992a <=( A199  and  A166 );
 a82995a <=( A201  and  (not A200) );
 a82996a <=( a82995a  and  a82992a );
 a82997a <=( a82996a  and  a82989a );
 a83000a <=( A265  and  A202 );
 a83003a <=( (not A267)  and  (not A266) );
 a83004a <=( a83003a  and  a83000a );
 a83007a <=( (not A269)  and  (not A268) );
 a83010a <=( (not A299)  and  (not A298) );
 a83011a <=( a83010a  and  a83007a );
 a83012a <=( a83011a  and  a83004a );
 a83016a <=( (not A167)  and  A168 );
 a83017a <=( A169  and  a83016a );
 a83020a <=( A199  and  A166 );
 a83023a <=( A201  and  (not A200) );
 a83024a <=( a83023a  and  a83020a );
 a83025a <=( a83024a  and  a83017a );
 a83028a <=( (not A265)  and  A203 );
 a83031a <=( A267  and  A266 );
 a83032a <=( a83031a  and  a83028a );
 a83035a <=( A300  and  A268 );
 a83038a <=( (not A302)  and  (not A301) );
 a83039a <=( a83038a  and  a83035a );
 a83040a <=( a83039a  and  a83032a );
 a83044a <=( (not A167)  and  A168 );
 a83045a <=( A169  and  a83044a );
 a83048a <=( A199  and  A166 );
 a83051a <=( A201  and  (not A200) );
 a83052a <=( a83051a  and  a83048a );
 a83053a <=( a83052a  and  a83045a );
 a83056a <=( (not A265)  and  A203 );
 a83059a <=( A267  and  A266 );
 a83060a <=( a83059a  and  a83056a );
 a83063a <=( A300  and  A269 );
 a83066a <=( (not A302)  and  (not A301) );
 a83067a <=( a83066a  and  a83063a );
 a83068a <=( a83067a  and  a83060a );
 a83072a <=( (not A167)  and  A168 );
 a83073a <=( A169  and  a83072a );
 a83076a <=( A199  and  A166 );
 a83079a <=( A201  and  (not A200) );
 a83080a <=( a83079a  and  a83076a );
 a83081a <=( a83080a  and  a83073a );
 a83084a <=( (not A265)  and  A203 );
 a83087a <=( (not A267)  and  A266 );
 a83088a <=( a83087a  and  a83084a );
 a83091a <=( (not A269)  and  (not A268) );
 a83094a <=( A301  and  (not A300) );
 a83095a <=( a83094a  and  a83091a );
 a83096a <=( a83095a  and  a83088a );
 a83100a <=( (not A167)  and  A168 );
 a83101a <=( A169  and  a83100a );
 a83104a <=( A199  and  A166 );
 a83107a <=( A201  and  (not A200) );
 a83108a <=( a83107a  and  a83104a );
 a83109a <=( a83108a  and  a83101a );
 a83112a <=( (not A265)  and  A203 );
 a83115a <=( (not A267)  and  A266 );
 a83116a <=( a83115a  and  a83112a );
 a83119a <=( (not A269)  and  (not A268) );
 a83122a <=( A302  and  (not A300) );
 a83123a <=( a83122a  and  a83119a );
 a83124a <=( a83123a  and  a83116a );
 a83128a <=( (not A167)  and  A168 );
 a83129a <=( A169  and  a83128a );
 a83132a <=( A199  and  A166 );
 a83135a <=( A201  and  (not A200) );
 a83136a <=( a83135a  and  a83132a );
 a83137a <=( a83136a  and  a83129a );
 a83140a <=( (not A265)  and  A203 );
 a83143a <=( (not A267)  and  A266 );
 a83144a <=( a83143a  and  a83140a );
 a83147a <=( (not A269)  and  (not A268) );
 a83150a <=( A299  and  A298 );
 a83151a <=( a83150a  and  a83147a );
 a83152a <=( a83151a  and  a83144a );
 a83156a <=( (not A167)  and  A168 );
 a83157a <=( A169  and  a83156a );
 a83160a <=( A199  and  A166 );
 a83163a <=( A201  and  (not A200) );
 a83164a <=( a83163a  and  a83160a );
 a83165a <=( a83164a  and  a83157a );
 a83168a <=( (not A265)  and  A203 );
 a83171a <=( (not A267)  and  A266 );
 a83172a <=( a83171a  and  a83168a );
 a83175a <=( (not A269)  and  (not A268) );
 a83178a <=( (not A299)  and  (not A298) );
 a83179a <=( a83178a  and  a83175a );
 a83180a <=( a83179a  and  a83172a );
 a83184a <=( (not A167)  and  A168 );
 a83185a <=( A169  and  a83184a );
 a83188a <=( A199  and  A166 );
 a83191a <=( A201  and  (not A200) );
 a83192a <=( a83191a  and  a83188a );
 a83193a <=( a83192a  and  a83185a );
 a83196a <=( A265  and  A203 );
 a83199a <=( A267  and  (not A266) );
 a83200a <=( a83199a  and  a83196a );
 a83203a <=( A300  and  A268 );
 a83206a <=( (not A302)  and  (not A301) );
 a83207a <=( a83206a  and  a83203a );
 a83208a <=( a83207a  and  a83200a );
 a83212a <=( (not A167)  and  A168 );
 a83213a <=( A169  and  a83212a );
 a83216a <=( A199  and  A166 );
 a83219a <=( A201  and  (not A200) );
 a83220a <=( a83219a  and  a83216a );
 a83221a <=( a83220a  and  a83213a );
 a83224a <=( A265  and  A203 );
 a83227a <=( A267  and  (not A266) );
 a83228a <=( a83227a  and  a83224a );
 a83231a <=( A300  and  A269 );
 a83234a <=( (not A302)  and  (not A301) );
 a83235a <=( a83234a  and  a83231a );
 a83236a <=( a83235a  and  a83228a );
 a83240a <=( (not A167)  and  A168 );
 a83241a <=( A169  and  a83240a );
 a83244a <=( A199  and  A166 );
 a83247a <=( A201  and  (not A200) );
 a83248a <=( a83247a  and  a83244a );
 a83249a <=( a83248a  and  a83241a );
 a83252a <=( A265  and  A203 );
 a83255a <=( (not A267)  and  (not A266) );
 a83256a <=( a83255a  and  a83252a );
 a83259a <=( (not A269)  and  (not A268) );
 a83262a <=( A301  and  (not A300) );
 a83263a <=( a83262a  and  a83259a );
 a83264a <=( a83263a  and  a83256a );
 a83268a <=( (not A167)  and  A168 );
 a83269a <=( A169  and  a83268a );
 a83272a <=( A199  and  A166 );
 a83275a <=( A201  and  (not A200) );
 a83276a <=( a83275a  and  a83272a );
 a83277a <=( a83276a  and  a83269a );
 a83280a <=( A265  and  A203 );
 a83283a <=( (not A267)  and  (not A266) );
 a83284a <=( a83283a  and  a83280a );
 a83287a <=( (not A269)  and  (not A268) );
 a83290a <=( A302  and  (not A300) );
 a83291a <=( a83290a  and  a83287a );
 a83292a <=( a83291a  and  a83284a );
 a83296a <=( (not A167)  and  A168 );
 a83297a <=( A169  and  a83296a );
 a83300a <=( A199  and  A166 );
 a83303a <=( A201  and  (not A200) );
 a83304a <=( a83303a  and  a83300a );
 a83305a <=( a83304a  and  a83297a );
 a83308a <=( A265  and  A203 );
 a83311a <=( (not A267)  and  (not A266) );
 a83312a <=( a83311a  and  a83308a );
 a83315a <=( (not A269)  and  (not A268) );
 a83318a <=( A299  and  A298 );
 a83319a <=( a83318a  and  a83315a );
 a83320a <=( a83319a  and  a83312a );
 a83324a <=( (not A167)  and  A168 );
 a83325a <=( A169  and  a83324a );
 a83328a <=( A199  and  A166 );
 a83331a <=( A201  and  (not A200) );
 a83332a <=( a83331a  and  a83328a );
 a83333a <=( a83332a  and  a83325a );
 a83336a <=( A265  and  A203 );
 a83339a <=( (not A267)  and  (not A266) );
 a83340a <=( a83339a  and  a83336a );
 a83343a <=( (not A269)  and  (not A268) );
 a83346a <=( (not A299)  and  (not A298) );
 a83347a <=( a83346a  and  a83343a );
 a83348a <=( a83347a  and  a83340a );
 a83352a <=( (not A167)  and  A168 );
 a83353a <=( A169  and  a83352a );
 a83356a <=( A199  and  A166 );
 a83359a <=( (not A201)  and  (not A200) );
 a83360a <=( a83359a  and  a83356a );
 a83361a <=( a83360a  and  a83353a );
 a83364a <=( (not A203)  and  (not A202) );
 a83367a <=( A266  and  (not A265) );
 a83368a <=( a83367a  and  a83364a );
 a83371a <=( A268  and  A267 );
 a83374a <=( A301  and  (not A300) );
 a83375a <=( a83374a  and  a83371a );
 a83376a <=( a83375a  and  a83368a );
 a83380a <=( (not A167)  and  A168 );
 a83381a <=( A169  and  a83380a );
 a83384a <=( A199  and  A166 );
 a83387a <=( (not A201)  and  (not A200) );
 a83388a <=( a83387a  and  a83384a );
 a83389a <=( a83388a  and  a83381a );
 a83392a <=( (not A203)  and  (not A202) );
 a83395a <=( A266  and  (not A265) );
 a83396a <=( a83395a  and  a83392a );
 a83399a <=( A268  and  A267 );
 a83402a <=( A302  and  (not A300) );
 a83403a <=( a83402a  and  a83399a );
 a83404a <=( a83403a  and  a83396a );
 a83408a <=( (not A167)  and  A168 );
 a83409a <=( A169  and  a83408a );
 a83412a <=( A199  and  A166 );
 a83415a <=( (not A201)  and  (not A200) );
 a83416a <=( a83415a  and  a83412a );
 a83417a <=( a83416a  and  a83409a );
 a83420a <=( (not A203)  and  (not A202) );
 a83423a <=( A266  and  (not A265) );
 a83424a <=( a83423a  and  a83420a );
 a83427a <=( A268  and  A267 );
 a83430a <=( A299  and  A298 );
 a83431a <=( a83430a  and  a83427a );
 a83432a <=( a83431a  and  a83424a );
 a83436a <=( (not A167)  and  A168 );
 a83437a <=( A169  and  a83436a );
 a83440a <=( A199  and  A166 );
 a83443a <=( (not A201)  and  (not A200) );
 a83444a <=( a83443a  and  a83440a );
 a83445a <=( a83444a  and  a83437a );
 a83448a <=( (not A203)  and  (not A202) );
 a83451a <=( A266  and  (not A265) );
 a83452a <=( a83451a  and  a83448a );
 a83455a <=( A268  and  A267 );
 a83458a <=( (not A299)  and  (not A298) );
 a83459a <=( a83458a  and  a83455a );
 a83460a <=( a83459a  and  a83452a );
 a83464a <=( (not A167)  and  A168 );
 a83465a <=( A169  and  a83464a );
 a83468a <=( A199  and  A166 );
 a83471a <=( (not A201)  and  (not A200) );
 a83472a <=( a83471a  and  a83468a );
 a83473a <=( a83472a  and  a83465a );
 a83476a <=( (not A203)  and  (not A202) );
 a83479a <=( A266  and  (not A265) );
 a83480a <=( a83479a  and  a83476a );
 a83483a <=( A269  and  A267 );
 a83486a <=( A301  and  (not A300) );
 a83487a <=( a83486a  and  a83483a );
 a83488a <=( a83487a  and  a83480a );
 a83492a <=( (not A167)  and  A168 );
 a83493a <=( A169  and  a83492a );
 a83496a <=( A199  and  A166 );
 a83499a <=( (not A201)  and  (not A200) );
 a83500a <=( a83499a  and  a83496a );
 a83501a <=( a83500a  and  a83493a );
 a83504a <=( (not A203)  and  (not A202) );
 a83507a <=( A266  and  (not A265) );
 a83508a <=( a83507a  and  a83504a );
 a83511a <=( A269  and  A267 );
 a83514a <=( A302  and  (not A300) );
 a83515a <=( a83514a  and  a83511a );
 a83516a <=( a83515a  and  a83508a );
 a83520a <=( (not A167)  and  A168 );
 a83521a <=( A169  and  a83520a );
 a83524a <=( A199  and  A166 );
 a83527a <=( (not A201)  and  (not A200) );
 a83528a <=( a83527a  and  a83524a );
 a83529a <=( a83528a  and  a83521a );
 a83532a <=( (not A203)  and  (not A202) );
 a83535a <=( A266  and  (not A265) );
 a83536a <=( a83535a  and  a83532a );
 a83539a <=( A269  and  A267 );
 a83542a <=( A299  and  A298 );
 a83543a <=( a83542a  and  a83539a );
 a83544a <=( a83543a  and  a83536a );
 a83548a <=( (not A167)  and  A168 );
 a83549a <=( A169  and  a83548a );
 a83552a <=( A199  and  A166 );
 a83555a <=( (not A201)  and  (not A200) );
 a83556a <=( a83555a  and  a83552a );
 a83557a <=( a83556a  and  a83549a );
 a83560a <=( (not A203)  and  (not A202) );
 a83563a <=( A266  and  (not A265) );
 a83564a <=( a83563a  and  a83560a );
 a83567a <=( A269  and  A267 );
 a83570a <=( (not A299)  and  (not A298) );
 a83571a <=( a83570a  and  a83567a );
 a83572a <=( a83571a  and  a83564a );
 a83576a <=( (not A167)  and  A168 );
 a83577a <=( A169  and  a83576a );
 a83580a <=( A199  and  A166 );
 a83583a <=( (not A201)  and  (not A200) );
 a83584a <=( a83583a  and  a83580a );
 a83585a <=( a83584a  and  a83577a );
 a83588a <=( (not A203)  and  (not A202) );
 a83591a <=( (not A266)  and  A265 );
 a83592a <=( a83591a  and  a83588a );
 a83595a <=( A268  and  A267 );
 a83598a <=( A301  and  (not A300) );
 a83599a <=( a83598a  and  a83595a );
 a83600a <=( a83599a  and  a83592a );
 a83604a <=( (not A167)  and  A168 );
 a83605a <=( A169  and  a83604a );
 a83608a <=( A199  and  A166 );
 a83611a <=( (not A201)  and  (not A200) );
 a83612a <=( a83611a  and  a83608a );
 a83613a <=( a83612a  and  a83605a );
 a83616a <=( (not A203)  and  (not A202) );
 a83619a <=( (not A266)  and  A265 );
 a83620a <=( a83619a  and  a83616a );
 a83623a <=( A268  and  A267 );
 a83626a <=( A302  and  (not A300) );
 a83627a <=( a83626a  and  a83623a );
 a83628a <=( a83627a  and  a83620a );
 a83632a <=( (not A167)  and  A168 );
 a83633a <=( A169  and  a83632a );
 a83636a <=( A199  and  A166 );
 a83639a <=( (not A201)  and  (not A200) );
 a83640a <=( a83639a  and  a83636a );
 a83641a <=( a83640a  and  a83633a );
 a83644a <=( (not A203)  and  (not A202) );
 a83647a <=( (not A266)  and  A265 );
 a83648a <=( a83647a  and  a83644a );
 a83651a <=( A268  and  A267 );
 a83654a <=( A299  and  A298 );
 a83655a <=( a83654a  and  a83651a );
 a83656a <=( a83655a  and  a83648a );
 a83660a <=( (not A167)  and  A168 );
 a83661a <=( A169  and  a83660a );
 a83664a <=( A199  and  A166 );
 a83667a <=( (not A201)  and  (not A200) );
 a83668a <=( a83667a  and  a83664a );
 a83669a <=( a83668a  and  a83661a );
 a83672a <=( (not A203)  and  (not A202) );
 a83675a <=( (not A266)  and  A265 );
 a83676a <=( a83675a  and  a83672a );
 a83679a <=( A268  and  A267 );
 a83682a <=( (not A299)  and  (not A298) );
 a83683a <=( a83682a  and  a83679a );
 a83684a <=( a83683a  and  a83676a );
 a83688a <=( (not A167)  and  A168 );
 a83689a <=( A169  and  a83688a );
 a83692a <=( A199  and  A166 );
 a83695a <=( (not A201)  and  (not A200) );
 a83696a <=( a83695a  and  a83692a );
 a83697a <=( a83696a  and  a83689a );
 a83700a <=( (not A203)  and  (not A202) );
 a83703a <=( (not A266)  and  A265 );
 a83704a <=( a83703a  and  a83700a );
 a83707a <=( A269  and  A267 );
 a83710a <=( A301  and  (not A300) );
 a83711a <=( a83710a  and  a83707a );
 a83712a <=( a83711a  and  a83704a );
 a83716a <=( (not A167)  and  A168 );
 a83717a <=( A169  and  a83716a );
 a83720a <=( A199  and  A166 );
 a83723a <=( (not A201)  and  (not A200) );
 a83724a <=( a83723a  and  a83720a );
 a83725a <=( a83724a  and  a83717a );
 a83728a <=( (not A203)  and  (not A202) );
 a83731a <=( (not A266)  and  A265 );
 a83732a <=( a83731a  and  a83728a );
 a83735a <=( A269  and  A267 );
 a83738a <=( A302  and  (not A300) );
 a83739a <=( a83738a  and  a83735a );
 a83740a <=( a83739a  and  a83732a );
 a83744a <=( (not A167)  and  A168 );
 a83745a <=( A169  and  a83744a );
 a83748a <=( A199  and  A166 );
 a83751a <=( (not A201)  and  (not A200) );
 a83752a <=( a83751a  and  a83748a );
 a83753a <=( a83752a  and  a83745a );
 a83756a <=( (not A203)  and  (not A202) );
 a83759a <=( (not A266)  and  A265 );
 a83760a <=( a83759a  and  a83756a );
 a83763a <=( A269  and  A267 );
 a83766a <=( A299  and  A298 );
 a83767a <=( a83766a  and  a83763a );
 a83768a <=( a83767a  and  a83760a );
 a83772a <=( (not A167)  and  A168 );
 a83773a <=( A169  and  a83772a );
 a83776a <=( A199  and  A166 );
 a83779a <=( (not A201)  and  (not A200) );
 a83780a <=( a83779a  and  a83776a );
 a83781a <=( a83780a  and  a83773a );
 a83784a <=( (not A203)  and  (not A202) );
 a83787a <=( (not A266)  and  A265 );
 a83788a <=( a83787a  and  a83784a );
 a83791a <=( A269  and  A267 );
 a83794a <=( (not A299)  and  (not A298) );
 a83795a <=( a83794a  and  a83791a );
 a83796a <=( a83795a  and  a83788a );
 a83800a <=( (not A199)  and  (not A168) );
 a83801a <=( A169  and  a83800a );
 a83804a <=( (not A201)  and  A200 );
 a83807a <=( (not A203)  and  (not A202) );
 a83808a <=( a83807a  and  a83804a );
 a83809a <=( a83808a  and  a83801a );
 a83812a <=( (not A268)  and  A267 );
 a83815a <=( A298  and  (not A269) );
 a83816a <=( a83815a  and  a83812a );
 a83819a <=( (not A300)  and  (not A299) );
 a83822a <=( (not A302)  and  (not A301) );
 a83823a <=( a83822a  and  a83819a );
 a83824a <=( a83823a  and  a83816a );
 a83828a <=( (not A199)  and  (not A168) );
 a83829a <=( A169  and  a83828a );
 a83832a <=( (not A201)  and  A200 );
 a83835a <=( (not A203)  and  (not A202) );
 a83836a <=( a83835a  and  a83832a );
 a83837a <=( a83836a  and  a83829a );
 a83840a <=( (not A268)  and  A267 );
 a83843a <=( (not A298)  and  (not A269) );
 a83844a <=( a83843a  and  a83840a );
 a83847a <=( (not A300)  and  A299 );
 a83850a <=( (not A302)  and  (not A301) );
 a83851a <=( a83850a  and  a83847a );
 a83852a <=( a83851a  and  a83844a );
 a83856a <=( A199  and  (not A168) );
 a83857a <=( A169  and  a83856a );
 a83860a <=( (not A201)  and  (not A200) );
 a83863a <=( (not A203)  and  (not A202) );
 a83864a <=( a83863a  and  a83860a );
 a83865a <=( a83864a  and  a83857a );
 a83868a <=( (not A268)  and  A267 );
 a83871a <=( A298  and  (not A269) );
 a83872a <=( a83871a  and  a83868a );
 a83875a <=( (not A300)  and  (not A299) );
 a83878a <=( (not A302)  and  (not A301) );
 a83879a <=( a83878a  and  a83875a );
 a83880a <=( a83879a  and  a83872a );
 a83884a <=( A199  and  (not A168) );
 a83885a <=( A169  and  a83884a );
 a83888a <=( (not A201)  and  (not A200) );
 a83891a <=( (not A203)  and  (not A202) );
 a83892a <=( a83891a  and  a83888a );
 a83893a <=( a83892a  and  a83885a );
 a83896a <=( (not A268)  and  A267 );
 a83899a <=( (not A298)  and  (not A269) );
 a83900a <=( a83899a  and  a83896a );
 a83903a <=( (not A300)  and  A299 );
 a83906a <=( (not A302)  and  (not A301) );
 a83907a <=( a83906a  and  a83903a );
 a83908a <=( a83907a  and  a83900a );
 a83912a <=( A168  and  (not A169) );
 a83913a <=( A170  and  a83912a );
 a83916a <=( A200  and  (not A199) );
 a83919a <=( A202  and  A201 );
 a83920a <=( a83919a  and  a83916a );
 a83921a <=( a83920a  and  a83913a );
 a83924a <=( (not A268)  and  A267 );
 a83927a <=( A298  and  (not A269) );
 a83928a <=( a83927a  and  a83924a );
 a83931a <=( (not A300)  and  (not A299) );
 a83934a <=( (not A302)  and  (not A301) );
 a83935a <=( a83934a  and  a83931a );
 a83936a <=( a83935a  and  a83928a );
 a83940a <=( A168  and  (not A169) );
 a83941a <=( A170  and  a83940a );
 a83944a <=( A200  and  (not A199) );
 a83947a <=( A202  and  A201 );
 a83948a <=( a83947a  and  a83944a );
 a83949a <=( a83948a  and  a83941a );
 a83952a <=( (not A268)  and  A267 );
 a83955a <=( (not A298)  and  (not A269) );
 a83956a <=( a83955a  and  a83952a );
 a83959a <=( (not A300)  and  A299 );
 a83962a <=( (not A302)  and  (not A301) );
 a83963a <=( a83962a  and  a83959a );
 a83964a <=( a83963a  and  a83956a );
 a83968a <=( A168  and  (not A169) );
 a83969a <=( A170  and  a83968a );
 a83972a <=( A200  and  (not A199) );
 a83975a <=( A203  and  A201 );
 a83976a <=( a83975a  and  a83972a );
 a83977a <=( a83976a  and  a83969a );
 a83980a <=( (not A268)  and  A267 );
 a83983a <=( A298  and  (not A269) );
 a83984a <=( a83983a  and  a83980a );
 a83987a <=( (not A300)  and  (not A299) );
 a83990a <=( (not A302)  and  (not A301) );
 a83991a <=( a83990a  and  a83987a );
 a83992a <=( a83991a  and  a83984a );
 a83996a <=( A168  and  (not A169) );
 a83997a <=( A170  and  a83996a );
 a84000a <=( A200  and  (not A199) );
 a84003a <=( A203  and  A201 );
 a84004a <=( a84003a  and  a84000a );
 a84005a <=( a84004a  and  a83997a );
 a84008a <=( (not A268)  and  A267 );
 a84011a <=( (not A298)  and  (not A269) );
 a84012a <=( a84011a  and  a84008a );
 a84015a <=( (not A300)  and  A299 );
 a84018a <=( (not A302)  and  (not A301) );
 a84019a <=( a84018a  and  a84015a );
 a84020a <=( a84019a  and  a84012a );
 a84024a <=( A168  and  (not A169) );
 a84025a <=( A170  and  a84024a );
 a84028a <=( A200  and  (not A199) );
 a84031a <=( (not A202)  and  (not A201) );
 a84032a <=( a84031a  and  a84028a );
 a84033a <=( a84032a  and  a84025a );
 a84036a <=( A267  and  (not A203) );
 a84039a <=( (not A269)  and  (not A268) );
 a84040a <=( a84039a  and  a84036a );
 a84043a <=( (not A299)  and  A298 );
 a84046a <=( A301  and  A300 );
 a84047a <=( a84046a  and  a84043a );
 a84048a <=( a84047a  and  a84040a );
 a84052a <=( A168  and  (not A169) );
 a84053a <=( A170  and  a84052a );
 a84056a <=( A200  and  (not A199) );
 a84059a <=( (not A202)  and  (not A201) );
 a84060a <=( a84059a  and  a84056a );
 a84061a <=( a84060a  and  a84053a );
 a84064a <=( A267  and  (not A203) );
 a84067a <=( (not A269)  and  (not A268) );
 a84068a <=( a84067a  and  a84064a );
 a84071a <=( (not A299)  and  A298 );
 a84074a <=( A302  and  A300 );
 a84075a <=( a84074a  and  a84071a );
 a84076a <=( a84075a  and  a84068a );
 a84080a <=( A168  and  (not A169) );
 a84081a <=( A170  and  a84080a );
 a84084a <=( A200  and  (not A199) );
 a84087a <=( (not A202)  and  (not A201) );
 a84088a <=( a84087a  and  a84084a );
 a84089a <=( a84088a  and  a84081a );
 a84092a <=( A267  and  (not A203) );
 a84095a <=( (not A269)  and  (not A268) );
 a84096a <=( a84095a  and  a84092a );
 a84099a <=( A299  and  (not A298) );
 a84102a <=( A301  and  A300 );
 a84103a <=( a84102a  and  a84099a );
 a84104a <=( a84103a  and  a84096a );
 a84108a <=( A168  and  (not A169) );
 a84109a <=( A170  and  a84108a );
 a84112a <=( A200  and  (not A199) );
 a84115a <=( (not A202)  and  (not A201) );
 a84116a <=( a84115a  and  a84112a );
 a84117a <=( a84116a  and  a84109a );
 a84120a <=( A267  and  (not A203) );
 a84123a <=( (not A269)  and  (not A268) );
 a84124a <=( a84123a  and  a84120a );
 a84127a <=( A299  and  (not A298) );
 a84130a <=( A302  and  A300 );
 a84131a <=( a84130a  and  a84127a );
 a84132a <=( a84131a  and  a84124a );
 a84136a <=( A168  and  (not A169) );
 a84137a <=( A170  and  a84136a );
 a84140a <=( A200  and  (not A199) );
 a84143a <=( (not A202)  and  (not A201) );
 a84144a <=( a84143a  and  a84140a );
 a84145a <=( a84144a  and  a84137a );
 a84148a <=( (not A267)  and  (not A203) );
 a84151a <=( A298  and  A268 );
 a84152a <=( a84151a  and  a84148a );
 a84155a <=( (not A300)  and  (not A299) );
 a84158a <=( (not A302)  and  (not A301) );
 a84159a <=( a84158a  and  a84155a );
 a84160a <=( a84159a  and  a84152a );
 a84164a <=( A168  and  (not A169) );
 a84165a <=( A170  and  a84164a );
 a84168a <=( A200  and  (not A199) );
 a84171a <=( (not A202)  and  (not A201) );
 a84172a <=( a84171a  and  a84168a );
 a84173a <=( a84172a  and  a84165a );
 a84176a <=( (not A267)  and  (not A203) );
 a84179a <=( (not A298)  and  A268 );
 a84180a <=( a84179a  and  a84176a );
 a84183a <=( (not A300)  and  A299 );
 a84186a <=( (not A302)  and  (not A301) );
 a84187a <=( a84186a  and  a84183a );
 a84188a <=( a84187a  and  a84180a );
 a84192a <=( A168  and  (not A169) );
 a84193a <=( A170  and  a84192a );
 a84196a <=( A200  and  (not A199) );
 a84199a <=( (not A202)  and  (not A201) );
 a84200a <=( a84199a  and  a84196a );
 a84201a <=( a84200a  and  a84193a );
 a84204a <=( (not A267)  and  (not A203) );
 a84207a <=( A298  and  A269 );
 a84208a <=( a84207a  and  a84204a );
 a84211a <=( (not A300)  and  (not A299) );
 a84214a <=( (not A302)  and  (not A301) );
 a84215a <=( a84214a  and  a84211a );
 a84216a <=( a84215a  and  a84208a );
 a84220a <=( A168  and  (not A169) );
 a84221a <=( A170  and  a84220a );
 a84224a <=( A200  and  (not A199) );
 a84227a <=( (not A202)  and  (not A201) );
 a84228a <=( a84227a  and  a84224a );
 a84229a <=( a84228a  and  a84221a );
 a84232a <=( (not A267)  and  (not A203) );
 a84235a <=( (not A298)  and  A269 );
 a84236a <=( a84235a  and  a84232a );
 a84239a <=( (not A300)  and  A299 );
 a84242a <=( (not A302)  and  (not A301) );
 a84243a <=( a84242a  and  a84239a );
 a84244a <=( a84243a  and  a84236a );
 a84248a <=( A168  and  (not A169) );
 a84249a <=( A170  and  a84248a );
 a84252a <=( A200  and  (not A199) );
 a84255a <=( (not A202)  and  (not A201) );
 a84256a <=( a84255a  and  a84252a );
 a84257a <=( a84256a  and  a84249a );
 a84260a <=( A265  and  (not A203) );
 a84263a <=( A298  and  A266 );
 a84264a <=( a84263a  and  a84260a );
 a84267a <=( (not A300)  and  (not A299) );
 a84270a <=( (not A302)  and  (not A301) );
 a84271a <=( a84270a  and  a84267a );
 a84272a <=( a84271a  and  a84264a );
 a84276a <=( A168  and  (not A169) );
 a84277a <=( A170  and  a84276a );
 a84280a <=( A200  and  (not A199) );
 a84283a <=( (not A202)  and  (not A201) );
 a84284a <=( a84283a  and  a84280a );
 a84285a <=( a84284a  and  a84277a );
 a84288a <=( A265  and  (not A203) );
 a84291a <=( (not A298)  and  A266 );
 a84292a <=( a84291a  and  a84288a );
 a84295a <=( (not A300)  and  A299 );
 a84298a <=( (not A302)  and  (not A301) );
 a84299a <=( a84298a  and  a84295a );
 a84300a <=( a84299a  and  a84292a );
 a84304a <=( A168  and  (not A169) );
 a84305a <=( A170  and  a84304a );
 a84308a <=( A200  and  (not A199) );
 a84311a <=( (not A202)  and  (not A201) );
 a84312a <=( a84311a  and  a84308a );
 a84313a <=( a84312a  and  a84305a );
 a84316a <=( (not A265)  and  (not A203) );
 a84319a <=( A298  and  (not A266) );
 a84320a <=( a84319a  and  a84316a );
 a84323a <=( (not A300)  and  (not A299) );
 a84326a <=( (not A302)  and  (not A301) );
 a84327a <=( a84326a  and  a84323a );
 a84328a <=( a84327a  and  a84320a );
 a84332a <=( A168  and  (not A169) );
 a84333a <=( A170  and  a84332a );
 a84336a <=( A200  and  (not A199) );
 a84339a <=( (not A202)  and  (not A201) );
 a84340a <=( a84339a  and  a84336a );
 a84341a <=( a84340a  and  a84333a );
 a84344a <=( (not A265)  and  (not A203) );
 a84347a <=( (not A298)  and  (not A266) );
 a84348a <=( a84347a  and  a84344a );
 a84351a <=( (not A300)  and  A299 );
 a84354a <=( (not A302)  and  (not A301) );
 a84355a <=( a84354a  and  a84351a );
 a84356a <=( a84355a  and  a84348a );
 a84360a <=( A168  and  (not A169) );
 a84361a <=( A170  and  a84360a );
 a84364a <=( (not A200)  and  A199 );
 a84367a <=( A202  and  A201 );
 a84368a <=( a84367a  and  a84364a );
 a84369a <=( a84368a  and  a84361a );
 a84372a <=( (not A268)  and  A267 );
 a84375a <=( A298  and  (not A269) );
 a84376a <=( a84375a  and  a84372a );
 a84379a <=( (not A300)  and  (not A299) );
 a84382a <=( (not A302)  and  (not A301) );
 a84383a <=( a84382a  and  a84379a );
 a84384a <=( a84383a  and  a84376a );
 a84388a <=( A168  and  (not A169) );
 a84389a <=( A170  and  a84388a );
 a84392a <=( (not A200)  and  A199 );
 a84395a <=( A202  and  A201 );
 a84396a <=( a84395a  and  a84392a );
 a84397a <=( a84396a  and  a84389a );
 a84400a <=( (not A268)  and  A267 );
 a84403a <=( (not A298)  and  (not A269) );
 a84404a <=( a84403a  and  a84400a );
 a84407a <=( (not A300)  and  A299 );
 a84410a <=( (not A302)  and  (not A301) );
 a84411a <=( a84410a  and  a84407a );
 a84412a <=( a84411a  and  a84404a );
 a84416a <=( A168  and  (not A169) );
 a84417a <=( A170  and  a84416a );
 a84420a <=( (not A200)  and  A199 );
 a84423a <=( A203  and  A201 );
 a84424a <=( a84423a  and  a84420a );
 a84425a <=( a84424a  and  a84417a );
 a84428a <=( (not A268)  and  A267 );
 a84431a <=( A298  and  (not A269) );
 a84432a <=( a84431a  and  a84428a );
 a84435a <=( (not A300)  and  (not A299) );
 a84438a <=( (not A302)  and  (not A301) );
 a84439a <=( a84438a  and  a84435a );
 a84440a <=( a84439a  and  a84432a );
 a84444a <=( A168  and  (not A169) );
 a84445a <=( A170  and  a84444a );
 a84448a <=( (not A200)  and  A199 );
 a84451a <=( A203  and  A201 );
 a84452a <=( a84451a  and  a84448a );
 a84453a <=( a84452a  and  a84445a );
 a84456a <=( (not A268)  and  A267 );
 a84459a <=( (not A298)  and  (not A269) );
 a84460a <=( a84459a  and  a84456a );
 a84463a <=( (not A300)  and  A299 );
 a84466a <=( (not A302)  and  (not A301) );
 a84467a <=( a84466a  and  a84463a );
 a84468a <=( a84467a  and  a84460a );
 a84472a <=( A168  and  (not A169) );
 a84473a <=( A170  and  a84472a );
 a84476a <=( (not A200)  and  A199 );
 a84479a <=( (not A202)  and  (not A201) );
 a84480a <=( a84479a  and  a84476a );
 a84481a <=( a84480a  and  a84473a );
 a84484a <=( A267  and  (not A203) );
 a84487a <=( (not A269)  and  (not A268) );
 a84488a <=( a84487a  and  a84484a );
 a84491a <=( (not A299)  and  A298 );
 a84494a <=( A301  and  A300 );
 a84495a <=( a84494a  and  a84491a );
 a84496a <=( a84495a  and  a84488a );
 a84500a <=( A168  and  (not A169) );
 a84501a <=( A170  and  a84500a );
 a84504a <=( (not A200)  and  A199 );
 a84507a <=( (not A202)  and  (not A201) );
 a84508a <=( a84507a  and  a84504a );
 a84509a <=( a84508a  and  a84501a );
 a84512a <=( A267  and  (not A203) );
 a84515a <=( (not A269)  and  (not A268) );
 a84516a <=( a84515a  and  a84512a );
 a84519a <=( (not A299)  and  A298 );
 a84522a <=( A302  and  A300 );
 a84523a <=( a84522a  and  a84519a );
 a84524a <=( a84523a  and  a84516a );
 a84528a <=( A168  and  (not A169) );
 a84529a <=( A170  and  a84528a );
 a84532a <=( (not A200)  and  A199 );
 a84535a <=( (not A202)  and  (not A201) );
 a84536a <=( a84535a  and  a84532a );
 a84537a <=( a84536a  and  a84529a );
 a84540a <=( A267  and  (not A203) );
 a84543a <=( (not A269)  and  (not A268) );
 a84544a <=( a84543a  and  a84540a );
 a84547a <=( A299  and  (not A298) );
 a84550a <=( A301  and  A300 );
 a84551a <=( a84550a  and  a84547a );
 a84552a <=( a84551a  and  a84544a );
 a84556a <=( A168  and  (not A169) );
 a84557a <=( A170  and  a84556a );
 a84560a <=( (not A200)  and  A199 );
 a84563a <=( (not A202)  and  (not A201) );
 a84564a <=( a84563a  and  a84560a );
 a84565a <=( a84564a  and  a84557a );
 a84568a <=( A267  and  (not A203) );
 a84571a <=( (not A269)  and  (not A268) );
 a84572a <=( a84571a  and  a84568a );
 a84575a <=( A299  and  (not A298) );
 a84578a <=( A302  and  A300 );
 a84579a <=( a84578a  and  a84575a );
 a84580a <=( a84579a  and  a84572a );
 a84584a <=( A168  and  (not A169) );
 a84585a <=( A170  and  a84584a );
 a84588a <=( (not A200)  and  A199 );
 a84591a <=( (not A202)  and  (not A201) );
 a84592a <=( a84591a  and  a84588a );
 a84593a <=( a84592a  and  a84585a );
 a84596a <=( (not A267)  and  (not A203) );
 a84599a <=( A298  and  A268 );
 a84600a <=( a84599a  and  a84596a );
 a84603a <=( (not A300)  and  (not A299) );
 a84606a <=( (not A302)  and  (not A301) );
 a84607a <=( a84606a  and  a84603a );
 a84608a <=( a84607a  and  a84600a );
 a84612a <=( A168  and  (not A169) );
 a84613a <=( A170  and  a84612a );
 a84616a <=( (not A200)  and  A199 );
 a84619a <=( (not A202)  and  (not A201) );
 a84620a <=( a84619a  and  a84616a );
 a84621a <=( a84620a  and  a84613a );
 a84624a <=( (not A267)  and  (not A203) );
 a84627a <=( (not A298)  and  A268 );
 a84628a <=( a84627a  and  a84624a );
 a84631a <=( (not A300)  and  A299 );
 a84634a <=( (not A302)  and  (not A301) );
 a84635a <=( a84634a  and  a84631a );
 a84636a <=( a84635a  and  a84628a );
 a84640a <=( A168  and  (not A169) );
 a84641a <=( A170  and  a84640a );
 a84644a <=( (not A200)  and  A199 );
 a84647a <=( (not A202)  and  (not A201) );
 a84648a <=( a84647a  and  a84644a );
 a84649a <=( a84648a  and  a84641a );
 a84652a <=( (not A267)  and  (not A203) );
 a84655a <=( A298  and  A269 );
 a84656a <=( a84655a  and  a84652a );
 a84659a <=( (not A300)  and  (not A299) );
 a84662a <=( (not A302)  and  (not A301) );
 a84663a <=( a84662a  and  a84659a );
 a84664a <=( a84663a  and  a84656a );
 a84668a <=( A168  and  (not A169) );
 a84669a <=( A170  and  a84668a );
 a84672a <=( (not A200)  and  A199 );
 a84675a <=( (not A202)  and  (not A201) );
 a84676a <=( a84675a  and  a84672a );
 a84677a <=( a84676a  and  a84669a );
 a84680a <=( (not A267)  and  (not A203) );
 a84683a <=( (not A298)  and  A269 );
 a84684a <=( a84683a  and  a84680a );
 a84687a <=( (not A300)  and  A299 );
 a84690a <=( (not A302)  and  (not A301) );
 a84691a <=( a84690a  and  a84687a );
 a84692a <=( a84691a  and  a84684a );
 a84696a <=( A168  and  (not A169) );
 a84697a <=( A170  and  a84696a );
 a84700a <=( (not A200)  and  A199 );
 a84703a <=( (not A202)  and  (not A201) );
 a84704a <=( a84703a  and  a84700a );
 a84705a <=( a84704a  and  a84697a );
 a84708a <=( A265  and  (not A203) );
 a84711a <=( A298  and  A266 );
 a84712a <=( a84711a  and  a84708a );
 a84715a <=( (not A300)  and  (not A299) );
 a84718a <=( (not A302)  and  (not A301) );
 a84719a <=( a84718a  and  a84715a );
 a84720a <=( a84719a  and  a84712a );
 a84724a <=( A168  and  (not A169) );
 a84725a <=( A170  and  a84724a );
 a84728a <=( (not A200)  and  A199 );
 a84731a <=( (not A202)  and  (not A201) );
 a84732a <=( a84731a  and  a84728a );
 a84733a <=( a84732a  and  a84725a );
 a84736a <=( A265  and  (not A203) );
 a84739a <=( (not A298)  and  A266 );
 a84740a <=( a84739a  and  a84736a );
 a84743a <=( (not A300)  and  A299 );
 a84746a <=( (not A302)  and  (not A301) );
 a84747a <=( a84746a  and  a84743a );
 a84748a <=( a84747a  and  a84740a );
 a84752a <=( A168  and  (not A169) );
 a84753a <=( A170  and  a84752a );
 a84756a <=( (not A200)  and  A199 );
 a84759a <=( (not A202)  and  (not A201) );
 a84760a <=( a84759a  and  a84756a );
 a84761a <=( a84760a  and  a84753a );
 a84764a <=( (not A265)  and  (not A203) );
 a84767a <=( A298  and  (not A266) );
 a84768a <=( a84767a  and  a84764a );
 a84771a <=( (not A300)  and  (not A299) );
 a84774a <=( (not A302)  and  (not A301) );
 a84775a <=( a84774a  and  a84771a );
 a84776a <=( a84775a  and  a84768a );
 a84780a <=( A168  and  (not A169) );
 a84781a <=( A170  and  a84780a );
 a84784a <=( (not A200)  and  A199 );
 a84787a <=( (not A202)  and  (not A201) );
 a84788a <=( a84787a  and  a84784a );
 a84789a <=( a84788a  and  a84781a );
 a84792a <=( (not A265)  and  (not A203) );
 a84795a <=( (not A298)  and  (not A266) );
 a84796a <=( a84795a  and  a84792a );
 a84799a <=( (not A300)  and  A299 );
 a84802a <=( (not A302)  and  (not A301) );
 a84803a <=( a84802a  and  a84799a );
 a84804a <=( a84803a  and  a84796a );
 a84808a <=( (not A168)  and  (not A169) );
 a84809a <=( A170  and  a84808a );
 a84812a <=( (not A166)  and  A167 );
 a84815a <=( (not A202)  and  A201 );
 a84816a <=( a84815a  and  a84812a );
 a84817a <=( a84816a  and  a84809a );
 a84820a <=( A267  and  (not A203) );
 a84823a <=( (not A269)  and  (not A268) );
 a84824a <=( a84823a  and  a84820a );
 a84827a <=( (not A299)  and  A298 );
 a84830a <=( A301  and  A300 );
 a84831a <=( a84830a  and  a84827a );
 a84832a <=( a84831a  and  a84824a );
 a84836a <=( (not A168)  and  (not A169) );
 a84837a <=( A170  and  a84836a );
 a84840a <=( (not A166)  and  A167 );
 a84843a <=( (not A202)  and  A201 );
 a84844a <=( a84843a  and  a84840a );
 a84845a <=( a84844a  and  a84837a );
 a84848a <=( A267  and  (not A203) );
 a84851a <=( (not A269)  and  (not A268) );
 a84852a <=( a84851a  and  a84848a );
 a84855a <=( (not A299)  and  A298 );
 a84858a <=( A302  and  A300 );
 a84859a <=( a84858a  and  a84855a );
 a84860a <=( a84859a  and  a84852a );
 a84864a <=( (not A168)  and  (not A169) );
 a84865a <=( A170  and  a84864a );
 a84868a <=( (not A166)  and  A167 );
 a84871a <=( (not A202)  and  A201 );
 a84872a <=( a84871a  and  a84868a );
 a84873a <=( a84872a  and  a84865a );
 a84876a <=( A267  and  (not A203) );
 a84879a <=( (not A269)  and  (not A268) );
 a84880a <=( a84879a  and  a84876a );
 a84883a <=( A299  and  (not A298) );
 a84886a <=( A301  and  A300 );
 a84887a <=( a84886a  and  a84883a );
 a84888a <=( a84887a  and  a84880a );
 a84892a <=( (not A168)  and  (not A169) );
 a84893a <=( A170  and  a84892a );
 a84896a <=( (not A166)  and  A167 );
 a84899a <=( (not A202)  and  A201 );
 a84900a <=( a84899a  and  a84896a );
 a84901a <=( a84900a  and  a84893a );
 a84904a <=( A267  and  (not A203) );
 a84907a <=( (not A269)  and  (not A268) );
 a84908a <=( a84907a  and  a84904a );
 a84911a <=( A299  and  (not A298) );
 a84914a <=( A302  and  A300 );
 a84915a <=( a84914a  and  a84911a );
 a84916a <=( a84915a  and  a84908a );
 a84920a <=( (not A168)  and  (not A169) );
 a84921a <=( A170  and  a84920a );
 a84924a <=( (not A166)  and  A167 );
 a84927a <=( (not A202)  and  A201 );
 a84928a <=( a84927a  and  a84924a );
 a84929a <=( a84928a  and  a84921a );
 a84932a <=( (not A267)  and  (not A203) );
 a84935a <=( A298  and  A268 );
 a84936a <=( a84935a  and  a84932a );
 a84939a <=( (not A300)  and  (not A299) );
 a84942a <=( (not A302)  and  (not A301) );
 a84943a <=( a84942a  and  a84939a );
 a84944a <=( a84943a  and  a84936a );
 a84948a <=( (not A168)  and  (not A169) );
 a84949a <=( A170  and  a84948a );
 a84952a <=( (not A166)  and  A167 );
 a84955a <=( (not A202)  and  A201 );
 a84956a <=( a84955a  and  a84952a );
 a84957a <=( a84956a  and  a84949a );
 a84960a <=( (not A267)  and  (not A203) );
 a84963a <=( (not A298)  and  A268 );
 a84964a <=( a84963a  and  a84960a );
 a84967a <=( (not A300)  and  A299 );
 a84970a <=( (not A302)  and  (not A301) );
 a84971a <=( a84970a  and  a84967a );
 a84972a <=( a84971a  and  a84964a );
 a84976a <=( (not A168)  and  (not A169) );
 a84977a <=( A170  and  a84976a );
 a84980a <=( (not A166)  and  A167 );
 a84983a <=( (not A202)  and  A201 );
 a84984a <=( a84983a  and  a84980a );
 a84985a <=( a84984a  and  a84977a );
 a84988a <=( (not A267)  and  (not A203) );
 a84991a <=( A298  and  A269 );
 a84992a <=( a84991a  and  a84988a );
 a84995a <=( (not A300)  and  (not A299) );
 a84998a <=( (not A302)  and  (not A301) );
 a84999a <=( a84998a  and  a84995a );
 a85000a <=( a84999a  and  a84992a );
 a85004a <=( (not A168)  and  (not A169) );
 a85005a <=( A170  and  a85004a );
 a85008a <=( (not A166)  and  A167 );
 a85011a <=( (not A202)  and  A201 );
 a85012a <=( a85011a  and  a85008a );
 a85013a <=( a85012a  and  a85005a );
 a85016a <=( (not A267)  and  (not A203) );
 a85019a <=( (not A298)  and  A269 );
 a85020a <=( a85019a  and  a85016a );
 a85023a <=( (not A300)  and  A299 );
 a85026a <=( (not A302)  and  (not A301) );
 a85027a <=( a85026a  and  a85023a );
 a85028a <=( a85027a  and  a85020a );
 a85032a <=( (not A168)  and  (not A169) );
 a85033a <=( A170  and  a85032a );
 a85036a <=( (not A166)  and  A167 );
 a85039a <=( (not A202)  and  A201 );
 a85040a <=( a85039a  and  a85036a );
 a85041a <=( a85040a  and  a85033a );
 a85044a <=( A265  and  (not A203) );
 a85047a <=( A298  and  A266 );
 a85048a <=( a85047a  and  a85044a );
 a85051a <=( (not A300)  and  (not A299) );
 a85054a <=( (not A302)  and  (not A301) );
 a85055a <=( a85054a  and  a85051a );
 a85056a <=( a85055a  and  a85048a );
 a85060a <=( (not A168)  and  (not A169) );
 a85061a <=( A170  and  a85060a );
 a85064a <=( (not A166)  and  A167 );
 a85067a <=( (not A202)  and  A201 );
 a85068a <=( a85067a  and  a85064a );
 a85069a <=( a85068a  and  a85061a );
 a85072a <=( A265  and  (not A203) );
 a85075a <=( (not A298)  and  A266 );
 a85076a <=( a85075a  and  a85072a );
 a85079a <=( (not A300)  and  A299 );
 a85082a <=( (not A302)  and  (not A301) );
 a85083a <=( a85082a  and  a85079a );
 a85084a <=( a85083a  and  a85076a );
 a85088a <=( (not A168)  and  (not A169) );
 a85089a <=( A170  and  a85088a );
 a85092a <=( (not A166)  and  A167 );
 a85095a <=( (not A202)  and  A201 );
 a85096a <=( a85095a  and  a85092a );
 a85097a <=( a85096a  and  a85089a );
 a85100a <=( (not A265)  and  (not A203) );
 a85103a <=( A298  and  (not A266) );
 a85104a <=( a85103a  and  a85100a );
 a85107a <=( (not A300)  and  (not A299) );
 a85110a <=( (not A302)  and  (not A301) );
 a85111a <=( a85110a  and  a85107a );
 a85112a <=( a85111a  and  a85104a );
 a85116a <=( (not A168)  and  (not A169) );
 a85117a <=( A170  and  a85116a );
 a85120a <=( (not A166)  and  A167 );
 a85123a <=( (not A202)  and  A201 );
 a85124a <=( a85123a  and  a85120a );
 a85125a <=( a85124a  and  a85117a );
 a85128a <=( (not A265)  and  (not A203) );
 a85131a <=( (not A298)  and  (not A266) );
 a85132a <=( a85131a  and  a85128a );
 a85135a <=( (not A300)  and  A299 );
 a85138a <=( (not A302)  and  (not A301) );
 a85139a <=( a85138a  and  a85135a );
 a85140a <=( a85139a  and  a85132a );
 a85144a <=( (not A168)  and  (not A169) );
 a85145a <=( A170  and  a85144a );
 a85148a <=( (not A166)  and  A167 );
 a85151a <=( A202  and  (not A201) );
 a85152a <=( a85151a  and  a85148a );
 a85153a <=( a85152a  and  a85145a );
 a85156a <=( (not A268)  and  A267 );
 a85159a <=( A298  and  (not A269) );
 a85160a <=( a85159a  and  a85156a );
 a85163a <=( (not A300)  and  (not A299) );
 a85166a <=( (not A302)  and  (not A301) );
 a85167a <=( a85166a  and  a85163a );
 a85168a <=( a85167a  and  a85160a );
 a85172a <=( (not A168)  and  (not A169) );
 a85173a <=( A170  and  a85172a );
 a85176a <=( (not A166)  and  A167 );
 a85179a <=( A202  and  (not A201) );
 a85180a <=( a85179a  and  a85176a );
 a85181a <=( a85180a  and  a85173a );
 a85184a <=( (not A268)  and  A267 );
 a85187a <=( (not A298)  and  (not A269) );
 a85188a <=( a85187a  and  a85184a );
 a85191a <=( (not A300)  and  A299 );
 a85194a <=( (not A302)  and  (not A301) );
 a85195a <=( a85194a  and  a85191a );
 a85196a <=( a85195a  and  a85188a );
 a85200a <=( (not A168)  and  (not A169) );
 a85201a <=( A170  and  a85200a );
 a85204a <=( (not A166)  and  A167 );
 a85207a <=( A203  and  (not A201) );
 a85208a <=( a85207a  and  a85204a );
 a85209a <=( a85208a  and  a85201a );
 a85212a <=( (not A268)  and  A267 );
 a85215a <=( A298  and  (not A269) );
 a85216a <=( a85215a  and  a85212a );
 a85219a <=( (not A300)  and  (not A299) );
 a85222a <=( (not A302)  and  (not A301) );
 a85223a <=( a85222a  and  a85219a );
 a85224a <=( a85223a  and  a85216a );
 a85228a <=( (not A168)  and  (not A169) );
 a85229a <=( A170  and  a85228a );
 a85232a <=( (not A166)  and  A167 );
 a85235a <=( A203  and  (not A201) );
 a85236a <=( a85235a  and  a85232a );
 a85237a <=( a85236a  and  a85229a );
 a85240a <=( (not A268)  and  A267 );
 a85243a <=( (not A298)  and  (not A269) );
 a85244a <=( a85243a  and  a85240a );
 a85247a <=( (not A300)  and  A299 );
 a85250a <=( (not A302)  and  (not A301) );
 a85251a <=( a85250a  and  a85247a );
 a85252a <=( a85251a  and  a85244a );
 a85256a <=( (not A168)  and  (not A169) );
 a85257a <=( A170  and  a85256a );
 a85260a <=( (not A166)  and  A167 );
 a85263a <=( A200  and  A199 );
 a85264a <=( a85263a  and  a85260a );
 a85265a <=( a85264a  and  a85257a );
 a85268a <=( (not A268)  and  A267 );
 a85271a <=( A298  and  (not A269) );
 a85272a <=( a85271a  and  a85268a );
 a85275a <=( (not A300)  and  (not A299) );
 a85278a <=( (not A302)  and  (not A301) );
 a85279a <=( a85278a  and  a85275a );
 a85280a <=( a85279a  and  a85272a );
 a85284a <=( (not A168)  and  (not A169) );
 a85285a <=( A170  and  a85284a );
 a85288a <=( (not A166)  and  A167 );
 a85291a <=( A200  and  A199 );
 a85292a <=( a85291a  and  a85288a );
 a85293a <=( a85292a  and  a85285a );
 a85296a <=( (not A268)  and  A267 );
 a85299a <=( (not A298)  and  (not A269) );
 a85300a <=( a85299a  and  a85296a );
 a85303a <=( (not A300)  and  A299 );
 a85306a <=( (not A302)  and  (not A301) );
 a85307a <=( a85306a  and  a85303a );
 a85308a <=( a85307a  and  a85300a );
 a85312a <=( (not A168)  and  (not A169) );
 a85313a <=( A170  and  a85312a );
 a85316a <=( (not A166)  and  A167 );
 a85319a <=( A200  and  (not A199) );
 a85320a <=( a85319a  and  a85316a );
 a85321a <=( a85320a  and  a85313a );
 a85324a <=( A202  and  A201 );
 a85327a <=( A266  and  (not A265) );
 a85328a <=( a85327a  and  a85324a );
 a85331a <=( A268  and  A267 );
 a85334a <=( A301  and  (not A300) );
 a85335a <=( a85334a  and  a85331a );
 a85336a <=( a85335a  and  a85328a );
 a85340a <=( (not A168)  and  (not A169) );
 a85341a <=( A170  and  a85340a );
 a85344a <=( (not A166)  and  A167 );
 a85347a <=( A200  and  (not A199) );
 a85348a <=( a85347a  and  a85344a );
 a85349a <=( a85348a  and  a85341a );
 a85352a <=( A202  and  A201 );
 a85355a <=( A266  and  (not A265) );
 a85356a <=( a85355a  and  a85352a );
 a85359a <=( A268  and  A267 );
 a85362a <=( A302  and  (not A300) );
 a85363a <=( a85362a  and  a85359a );
 a85364a <=( a85363a  and  a85356a );
 a85368a <=( (not A168)  and  (not A169) );
 a85369a <=( A170  and  a85368a );
 a85372a <=( (not A166)  and  A167 );
 a85375a <=( A200  and  (not A199) );
 a85376a <=( a85375a  and  a85372a );
 a85377a <=( a85376a  and  a85369a );
 a85380a <=( A202  and  A201 );
 a85383a <=( A266  and  (not A265) );
 a85384a <=( a85383a  and  a85380a );
 a85387a <=( A268  and  A267 );
 a85390a <=( A299  and  A298 );
 a85391a <=( a85390a  and  a85387a );
 a85392a <=( a85391a  and  a85384a );
 a85396a <=( (not A168)  and  (not A169) );
 a85397a <=( A170  and  a85396a );
 a85400a <=( (not A166)  and  A167 );
 a85403a <=( A200  and  (not A199) );
 a85404a <=( a85403a  and  a85400a );
 a85405a <=( a85404a  and  a85397a );
 a85408a <=( A202  and  A201 );
 a85411a <=( A266  and  (not A265) );
 a85412a <=( a85411a  and  a85408a );
 a85415a <=( A268  and  A267 );
 a85418a <=( (not A299)  and  (not A298) );
 a85419a <=( a85418a  and  a85415a );
 a85420a <=( a85419a  and  a85412a );
 a85424a <=( (not A168)  and  (not A169) );
 a85425a <=( A170  and  a85424a );
 a85428a <=( (not A166)  and  A167 );
 a85431a <=( A200  and  (not A199) );
 a85432a <=( a85431a  and  a85428a );
 a85433a <=( a85432a  and  a85425a );
 a85436a <=( A202  and  A201 );
 a85439a <=( A266  and  (not A265) );
 a85440a <=( a85439a  and  a85436a );
 a85443a <=( A269  and  A267 );
 a85446a <=( A301  and  (not A300) );
 a85447a <=( a85446a  and  a85443a );
 a85448a <=( a85447a  and  a85440a );
 a85452a <=( (not A168)  and  (not A169) );
 a85453a <=( A170  and  a85452a );
 a85456a <=( (not A166)  and  A167 );
 a85459a <=( A200  and  (not A199) );
 a85460a <=( a85459a  and  a85456a );
 a85461a <=( a85460a  and  a85453a );
 a85464a <=( A202  and  A201 );
 a85467a <=( A266  and  (not A265) );
 a85468a <=( a85467a  and  a85464a );
 a85471a <=( A269  and  A267 );
 a85474a <=( A302  and  (not A300) );
 a85475a <=( a85474a  and  a85471a );
 a85476a <=( a85475a  and  a85468a );
 a85480a <=( (not A168)  and  (not A169) );
 a85481a <=( A170  and  a85480a );
 a85484a <=( (not A166)  and  A167 );
 a85487a <=( A200  and  (not A199) );
 a85488a <=( a85487a  and  a85484a );
 a85489a <=( a85488a  and  a85481a );
 a85492a <=( A202  and  A201 );
 a85495a <=( A266  and  (not A265) );
 a85496a <=( a85495a  and  a85492a );
 a85499a <=( A269  and  A267 );
 a85502a <=( A299  and  A298 );
 a85503a <=( a85502a  and  a85499a );
 a85504a <=( a85503a  and  a85496a );
 a85508a <=( (not A168)  and  (not A169) );
 a85509a <=( A170  and  a85508a );
 a85512a <=( (not A166)  and  A167 );
 a85515a <=( A200  and  (not A199) );
 a85516a <=( a85515a  and  a85512a );
 a85517a <=( a85516a  and  a85509a );
 a85520a <=( A202  and  A201 );
 a85523a <=( A266  and  (not A265) );
 a85524a <=( a85523a  and  a85520a );
 a85527a <=( A269  and  A267 );
 a85530a <=( (not A299)  and  (not A298) );
 a85531a <=( a85530a  and  a85527a );
 a85532a <=( a85531a  and  a85524a );
 a85536a <=( (not A168)  and  (not A169) );
 a85537a <=( A170  and  a85536a );
 a85540a <=( (not A166)  and  A167 );
 a85543a <=( A200  and  (not A199) );
 a85544a <=( a85543a  and  a85540a );
 a85545a <=( a85544a  and  a85537a );
 a85548a <=( A202  and  A201 );
 a85551a <=( (not A266)  and  A265 );
 a85552a <=( a85551a  and  a85548a );
 a85555a <=( A268  and  A267 );
 a85558a <=( A301  and  (not A300) );
 a85559a <=( a85558a  and  a85555a );
 a85560a <=( a85559a  and  a85552a );
 a85564a <=( (not A168)  and  (not A169) );
 a85565a <=( A170  and  a85564a );
 a85568a <=( (not A166)  and  A167 );
 a85571a <=( A200  and  (not A199) );
 a85572a <=( a85571a  and  a85568a );
 a85573a <=( a85572a  and  a85565a );
 a85576a <=( A202  and  A201 );
 a85579a <=( (not A266)  and  A265 );
 a85580a <=( a85579a  and  a85576a );
 a85583a <=( A268  and  A267 );
 a85586a <=( A302  and  (not A300) );
 a85587a <=( a85586a  and  a85583a );
 a85588a <=( a85587a  and  a85580a );
 a85592a <=( (not A168)  and  (not A169) );
 a85593a <=( A170  and  a85592a );
 a85596a <=( (not A166)  and  A167 );
 a85599a <=( A200  and  (not A199) );
 a85600a <=( a85599a  and  a85596a );
 a85601a <=( a85600a  and  a85593a );
 a85604a <=( A202  and  A201 );
 a85607a <=( (not A266)  and  A265 );
 a85608a <=( a85607a  and  a85604a );
 a85611a <=( A268  and  A267 );
 a85614a <=( A299  and  A298 );
 a85615a <=( a85614a  and  a85611a );
 a85616a <=( a85615a  and  a85608a );
 a85620a <=( (not A168)  and  (not A169) );
 a85621a <=( A170  and  a85620a );
 a85624a <=( (not A166)  and  A167 );
 a85627a <=( A200  and  (not A199) );
 a85628a <=( a85627a  and  a85624a );
 a85629a <=( a85628a  and  a85621a );
 a85632a <=( A202  and  A201 );
 a85635a <=( (not A266)  and  A265 );
 a85636a <=( a85635a  and  a85632a );
 a85639a <=( A268  and  A267 );
 a85642a <=( (not A299)  and  (not A298) );
 a85643a <=( a85642a  and  a85639a );
 a85644a <=( a85643a  and  a85636a );
 a85648a <=( (not A168)  and  (not A169) );
 a85649a <=( A170  and  a85648a );
 a85652a <=( (not A166)  and  A167 );
 a85655a <=( A200  and  (not A199) );
 a85656a <=( a85655a  and  a85652a );
 a85657a <=( a85656a  and  a85649a );
 a85660a <=( A202  and  A201 );
 a85663a <=( (not A266)  and  A265 );
 a85664a <=( a85663a  and  a85660a );
 a85667a <=( A269  and  A267 );
 a85670a <=( A301  and  (not A300) );
 a85671a <=( a85670a  and  a85667a );
 a85672a <=( a85671a  and  a85664a );
 a85676a <=( (not A168)  and  (not A169) );
 a85677a <=( A170  and  a85676a );
 a85680a <=( (not A166)  and  A167 );
 a85683a <=( A200  and  (not A199) );
 a85684a <=( a85683a  and  a85680a );
 a85685a <=( a85684a  and  a85677a );
 a85688a <=( A202  and  A201 );
 a85691a <=( (not A266)  and  A265 );
 a85692a <=( a85691a  and  a85688a );
 a85695a <=( A269  and  A267 );
 a85698a <=( A302  and  (not A300) );
 a85699a <=( a85698a  and  a85695a );
 a85700a <=( a85699a  and  a85692a );
 a85704a <=( (not A168)  and  (not A169) );
 a85705a <=( A170  and  a85704a );
 a85708a <=( (not A166)  and  A167 );
 a85711a <=( A200  and  (not A199) );
 a85712a <=( a85711a  and  a85708a );
 a85713a <=( a85712a  and  a85705a );
 a85716a <=( A202  and  A201 );
 a85719a <=( (not A266)  and  A265 );
 a85720a <=( a85719a  and  a85716a );
 a85723a <=( A269  and  A267 );
 a85726a <=( A299  and  A298 );
 a85727a <=( a85726a  and  a85723a );
 a85728a <=( a85727a  and  a85720a );
 a85732a <=( (not A168)  and  (not A169) );
 a85733a <=( A170  and  a85732a );
 a85736a <=( (not A166)  and  A167 );
 a85739a <=( A200  and  (not A199) );
 a85740a <=( a85739a  and  a85736a );
 a85741a <=( a85740a  and  a85733a );
 a85744a <=( A202  and  A201 );
 a85747a <=( (not A266)  and  A265 );
 a85748a <=( a85747a  and  a85744a );
 a85751a <=( A269  and  A267 );
 a85754a <=( (not A299)  and  (not A298) );
 a85755a <=( a85754a  and  a85751a );
 a85756a <=( a85755a  and  a85748a );
 a85760a <=( (not A168)  and  (not A169) );
 a85761a <=( A170  and  a85760a );
 a85764a <=( (not A166)  and  A167 );
 a85767a <=( A200  and  (not A199) );
 a85768a <=( a85767a  and  a85764a );
 a85769a <=( a85768a  and  a85761a );
 a85772a <=( A203  and  A201 );
 a85775a <=( A266  and  (not A265) );
 a85776a <=( a85775a  and  a85772a );
 a85779a <=( A268  and  A267 );
 a85782a <=( A301  and  (not A300) );
 a85783a <=( a85782a  and  a85779a );
 a85784a <=( a85783a  and  a85776a );
 a85788a <=( (not A168)  and  (not A169) );
 a85789a <=( A170  and  a85788a );
 a85792a <=( (not A166)  and  A167 );
 a85795a <=( A200  and  (not A199) );
 a85796a <=( a85795a  and  a85792a );
 a85797a <=( a85796a  and  a85789a );
 a85800a <=( A203  and  A201 );
 a85803a <=( A266  and  (not A265) );
 a85804a <=( a85803a  and  a85800a );
 a85807a <=( A268  and  A267 );
 a85810a <=( A302  and  (not A300) );
 a85811a <=( a85810a  and  a85807a );
 a85812a <=( a85811a  and  a85804a );
 a85816a <=( (not A168)  and  (not A169) );
 a85817a <=( A170  and  a85816a );
 a85820a <=( (not A166)  and  A167 );
 a85823a <=( A200  and  (not A199) );
 a85824a <=( a85823a  and  a85820a );
 a85825a <=( a85824a  and  a85817a );
 a85828a <=( A203  and  A201 );
 a85831a <=( A266  and  (not A265) );
 a85832a <=( a85831a  and  a85828a );
 a85835a <=( A268  and  A267 );
 a85838a <=( A299  and  A298 );
 a85839a <=( a85838a  and  a85835a );
 a85840a <=( a85839a  and  a85832a );
 a85844a <=( (not A168)  and  (not A169) );
 a85845a <=( A170  and  a85844a );
 a85848a <=( (not A166)  and  A167 );
 a85851a <=( A200  and  (not A199) );
 a85852a <=( a85851a  and  a85848a );
 a85853a <=( a85852a  and  a85845a );
 a85856a <=( A203  and  A201 );
 a85859a <=( A266  and  (not A265) );
 a85860a <=( a85859a  and  a85856a );
 a85863a <=( A268  and  A267 );
 a85866a <=( (not A299)  and  (not A298) );
 a85867a <=( a85866a  and  a85863a );
 a85868a <=( a85867a  and  a85860a );
 a85872a <=( (not A168)  and  (not A169) );
 a85873a <=( A170  and  a85872a );
 a85876a <=( (not A166)  and  A167 );
 a85879a <=( A200  and  (not A199) );
 a85880a <=( a85879a  and  a85876a );
 a85881a <=( a85880a  and  a85873a );
 a85884a <=( A203  and  A201 );
 a85887a <=( A266  and  (not A265) );
 a85888a <=( a85887a  and  a85884a );
 a85891a <=( A269  and  A267 );
 a85894a <=( A301  and  (not A300) );
 a85895a <=( a85894a  and  a85891a );
 a85896a <=( a85895a  and  a85888a );
 a85900a <=( (not A168)  and  (not A169) );
 a85901a <=( A170  and  a85900a );
 a85904a <=( (not A166)  and  A167 );
 a85907a <=( A200  and  (not A199) );
 a85908a <=( a85907a  and  a85904a );
 a85909a <=( a85908a  and  a85901a );
 a85912a <=( A203  and  A201 );
 a85915a <=( A266  and  (not A265) );
 a85916a <=( a85915a  and  a85912a );
 a85919a <=( A269  and  A267 );
 a85922a <=( A302  and  (not A300) );
 a85923a <=( a85922a  and  a85919a );
 a85924a <=( a85923a  and  a85916a );
 a85928a <=( (not A168)  and  (not A169) );
 a85929a <=( A170  and  a85928a );
 a85932a <=( (not A166)  and  A167 );
 a85935a <=( A200  and  (not A199) );
 a85936a <=( a85935a  and  a85932a );
 a85937a <=( a85936a  and  a85929a );
 a85940a <=( A203  and  A201 );
 a85943a <=( A266  and  (not A265) );
 a85944a <=( a85943a  and  a85940a );
 a85947a <=( A269  and  A267 );
 a85950a <=( A299  and  A298 );
 a85951a <=( a85950a  and  a85947a );
 a85952a <=( a85951a  and  a85944a );
 a85956a <=( (not A168)  and  (not A169) );
 a85957a <=( A170  and  a85956a );
 a85960a <=( (not A166)  and  A167 );
 a85963a <=( A200  and  (not A199) );
 a85964a <=( a85963a  and  a85960a );
 a85965a <=( a85964a  and  a85957a );
 a85968a <=( A203  and  A201 );
 a85971a <=( A266  and  (not A265) );
 a85972a <=( a85971a  and  a85968a );
 a85975a <=( A269  and  A267 );
 a85978a <=( (not A299)  and  (not A298) );
 a85979a <=( a85978a  and  a85975a );
 a85980a <=( a85979a  and  a85972a );
 a85984a <=( (not A168)  and  (not A169) );
 a85985a <=( A170  and  a85984a );
 a85988a <=( (not A166)  and  A167 );
 a85991a <=( A200  and  (not A199) );
 a85992a <=( a85991a  and  a85988a );
 a85993a <=( a85992a  and  a85985a );
 a85996a <=( A203  and  A201 );
 a85999a <=( (not A266)  and  A265 );
 a86000a <=( a85999a  and  a85996a );
 a86003a <=( A268  and  A267 );
 a86006a <=( A301  and  (not A300) );
 a86007a <=( a86006a  and  a86003a );
 a86008a <=( a86007a  and  a86000a );
 a86012a <=( (not A168)  and  (not A169) );
 a86013a <=( A170  and  a86012a );
 a86016a <=( (not A166)  and  A167 );
 a86019a <=( A200  and  (not A199) );
 a86020a <=( a86019a  and  a86016a );
 a86021a <=( a86020a  and  a86013a );
 a86024a <=( A203  and  A201 );
 a86027a <=( (not A266)  and  A265 );
 a86028a <=( a86027a  and  a86024a );
 a86031a <=( A268  and  A267 );
 a86034a <=( A302  and  (not A300) );
 a86035a <=( a86034a  and  a86031a );
 a86036a <=( a86035a  and  a86028a );
 a86040a <=( (not A168)  and  (not A169) );
 a86041a <=( A170  and  a86040a );
 a86044a <=( (not A166)  and  A167 );
 a86047a <=( A200  and  (not A199) );
 a86048a <=( a86047a  and  a86044a );
 a86049a <=( a86048a  and  a86041a );
 a86052a <=( A203  and  A201 );
 a86055a <=( (not A266)  and  A265 );
 a86056a <=( a86055a  and  a86052a );
 a86059a <=( A268  and  A267 );
 a86062a <=( A299  and  A298 );
 a86063a <=( a86062a  and  a86059a );
 a86064a <=( a86063a  and  a86056a );
 a86068a <=( (not A168)  and  (not A169) );
 a86069a <=( A170  and  a86068a );
 a86072a <=( (not A166)  and  A167 );
 a86075a <=( A200  and  (not A199) );
 a86076a <=( a86075a  and  a86072a );
 a86077a <=( a86076a  and  a86069a );
 a86080a <=( A203  and  A201 );
 a86083a <=( (not A266)  and  A265 );
 a86084a <=( a86083a  and  a86080a );
 a86087a <=( A268  and  A267 );
 a86090a <=( (not A299)  and  (not A298) );
 a86091a <=( a86090a  and  a86087a );
 a86092a <=( a86091a  and  a86084a );
 a86096a <=( (not A168)  and  (not A169) );
 a86097a <=( A170  and  a86096a );
 a86100a <=( (not A166)  and  A167 );
 a86103a <=( A200  and  (not A199) );
 a86104a <=( a86103a  and  a86100a );
 a86105a <=( a86104a  and  a86097a );
 a86108a <=( A203  and  A201 );
 a86111a <=( (not A266)  and  A265 );
 a86112a <=( a86111a  and  a86108a );
 a86115a <=( A269  and  A267 );
 a86118a <=( A301  and  (not A300) );
 a86119a <=( a86118a  and  a86115a );
 a86120a <=( a86119a  and  a86112a );
 a86124a <=( (not A168)  and  (not A169) );
 a86125a <=( A170  and  a86124a );
 a86128a <=( (not A166)  and  A167 );
 a86131a <=( A200  and  (not A199) );
 a86132a <=( a86131a  and  a86128a );
 a86133a <=( a86132a  and  a86125a );
 a86136a <=( A203  and  A201 );
 a86139a <=( (not A266)  and  A265 );
 a86140a <=( a86139a  and  a86136a );
 a86143a <=( A269  and  A267 );
 a86146a <=( A302  and  (not A300) );
 a86147a <=( a86146a  and  a86143a );
 a86148a <=( a86147a  and  a86140a );
 a86152a <=( (not A168)  and  (not A169) );
 a86153a <=( A170  and  a86152a );
 a86156a <=( (not A166)  and  A167 );
 a86159a <=( A200  and  (not A199) );
 a86160a <=( a86159a  and  a86156a );
 a86161a <=( a86160a  and  a86153a );
 a86164a <=( A203  and  A201 );
 a86167a <=( (not A266)  and  A265 );
 a86168a <=( a86167a  and  a86164a );
 a86171a <=( A269  and  A267 );
 a86174a <=( A299  and  A298 );
 a86175a <=( a86174a  and  a86171a );
 a86176a <=( a86175a  and  a86168a );
 a86180a <=( (not A168)  and  (not A169) );
 a86181a <=( A170  and  a86180a );
 a86184a <=( (not A166)  and  A167 );
 a86187a <=( A200  and  (not A199) );
 a86188a <=( a86187a  and  a86184a );
 a86189a <=( a86188a  and  a86181a );
 a86192a <=( A203  and  A201 );
 a86195a <=( (not A266)  and  A265 );
 a86196a <=( a86195a  and  a86192a );
 a86199a <=( A269  and  A267 );
 a86202a <=( (not A299)  and  (not A298) );
 a86203a <=( a86202a  and  a86199a );
 a86204a <=( a86203a  and  a86196a );
 a86208a <=( (not A168)  and  (not A169) );
 a86209a <=( A170  and  a86208a );
 a86212a <=( (not A166)  and  A167 );
 a86215a <=( (not A200)  and  A199 );
 a86216a <=( a86215a  and  a86212a );
 a86217a <=( a86216a  and  a86209a );
 a86220a <=( A202  and  A201 );
 a86223a <=( A266  and  (not A265) );
 a86224a <=( a86223a  and  a86220a );
 a86227a <=( A268  and  A267 );
 a86230a <=( A301  and  (not A300) );
 a86231a <=( a86230a  and  a86227a );
 a86232a <=( a86231a  and  a86224a );
 a86236a <=( (not A168)  and  (not A169) );
 a86237a <=( A170  and  a86236a );
 a86240a <=( (not A166)  and  A167 );
 a86243a <=( (not A200)  and  A199 );
 a86244a <=( a86243a  and  a86240a );
 a86245a <=( a86244a  and  a86237a );
 a86248a <=( A202  and  A201 );
 a86251a <=( A266  and  (not A265) );
 a86252a <=( a86251a  and  a86248a );
 a86255a <=( A268  and  A267 );
 a86258a <=( A302  and  (not A300) );
 a86259a <=( a86258a  and  a86255a );
 a86260a <=( a86259a  and  a86252a );
 a86264a <=( (not A168)  and  (not A169) );
 a86265a <=( A170  and  a86264a );
 a86268a <=( (not A166)  and  A167 );
 a86271a <=( (not A200)  and  A199 );
 a86272a <=( a86271a  and  a86268a );
 a86273a <=( a86272a  and  a86265a );
 a86276a <=( A202  and  A201 );
 a86279a <=( A266  and  (not A265) );
 a86280a <=( a86279a  and  a86276a );
 a86283a <=( A268  and  A267 );
 a86286a <=( A299  and  A298 );
 a86287a <=( a86286a  and  a86283a );
 a86288a <=( a86287a  and  a86280a );
 a86292a <=( (not A168)  and  (not A169) );
 a86293a <=( A170  and  a86292a );
 a86296a <=( (not A166)  and  A167 );
 a86299a <=( (not A200)  and  A199 );
 a86300a <=( a86299a  and  a86296a );
 a86301a <=( a86300a  and  a86293a );
 a86304a <=( A202  and  A201 );
 a86307a <=( A266  and  (not A265) );
 a86308a <=( a86307a  and  a86304a );
 a86311a <=( A268  and  A267 );
 a86314a <=( (not A299)  and  (not A298) );
 a86315a <=( a86314a  and  a86311a );
 a86316a <=( a86315a  and  a86308a );
 a86320a <=( (not A168)  and  (not A169) );
 a86321a <=( A170  and  a86320a );
 a86324a <=( (not A166)  and  A167 );
 a86327a <=( (not A200)  and  A199 );
 a86328a <=( a86327a  and  a86324a );
 a86329a <=( a86328a  and  a86321a );
 a86332a <=( A202  and  A201 );
 a86335a <=( A266  and  (not A265) );
 a86336a <=( a86335a  and  a86332a );
 a86339a <=( A269  and  A267 );
 a86342a <=( A301  and  (not A300) );
 a86343a <=( a86342a  and  a86339a );
 a86344a <=( a86343a  and  a86336a );
 a86348a <=( (not A168)  and  (not A169) );
 a86349a <=( A170  and  a86348a );
 a86352a <=( (not A166)  and  A167 );
 a86355a <=( (not A200)  and  A199 );
 a86356a <=( a86355a  and  a86352a );
 a86357a <=( a86356a  and  a86349a );
 a86360a <=( A202  and  A201 );
 a86363a <=( A266  and  (not A265) );
 a86364a <=( a86363a  and  a86360a );
 a86367a <=( A269  and  A267 );
 a86370a <=( A302  and  (not A300) );
 a86371a <=( a86370a  and  a86367a );
 a86372a <=( a86371a  and  a86364a );
 a86376a <=( (not A168)  and  (not A169) );
 a86377a <=( A170  and  a86376a );
 a86380a <=( (not A166)  and  A167 );
 a86383a <=( (not A200)  and  A199 );
 a86384a <=( a86383a  and  a86380a );
 a86385a <=( a86384a  and  a86377a );
 a86388a <=( A202  and  A201 );
 a86391a <=( A266  and  (not A265) );
 a86392a <=( a86391a  and  a86388a );
 a86395a <=( A269  and  A267 );
 a86398a <=( A299  and  A298 );
 a86399a <=( a86398a  and  a86395a );
 a86400a <=( a86399a  and  a86392a );
 a86404a <=( (not A168)  and  (not A169) );
 a86405a <=( A170  and  a86404a );
 a86408a <=( (not A166)  and  A167 );
 a86411a <=( (not A200)  and  A199 );
 a86412a <=( a86411a  and  a86408a );
 a86413a <=( a86412a  and  a86405a );
 a86416a <=( A202  and  A201 );
 a86419a <=( A266  and  (not A265) );
 a86420a <=( a86419a  and  a86416a );
 a86423a <=( A269  and  A267 );
 a86426a <=( (not A299)  and  (not A298) );
 a86427a <=( a86426a  and  a86423a );
 a86428a <=( a86427a  and  a86420a );
 a86432a <=( (not A168)  and  (not A169) );
 a86433a <=( A170  and  a86432a );
 a86436a <=( (not A166)  and  A167 );
 a86439a <=( (not A200)  and  A199 );
 a86440a <=( a86439a  and  a86436a );
 a86441a <=( a86440a  and  a86433a );
 a86444a <=( A202  and  A201 );
 a86447a <=( (not A266)  and  A265 );
 a86448a <=( a86447a  and  a86444a );
 a86451a <=( A268  and  A267 );
 a86454a <=( A301  and  (not A300) );
 a86455a <=( a86454a  and  a86451a );
 a86456a <=( a86455a  and  a86448a );
 a86460a <=( (not A168)  and  (not A169) );
 a86461a <=( A170  and  a86460a );
 a86464a <=( (not A166)  and  A167 );
 a86467a <=( (not A200)  and  A199 );
 a86468a <=( a86467a  and  a86464a );
 a86469a <=( a86468a  and  a86461a );
 a86472a <=( A202  and  A201 );
 a86475a <=( (not A266)  and  A265 );
 a86476a <=( a86475a  and  a86472a );
 a86479a <=( A268  and  A267 );
 a86482a <=( A302  and  (not A300) );
 a86483a <=( a86482a  and  a86479a );
 a86484a <=( a86483a  and  a86476a );
 a86488a <=( (not A168)  and  (not A169) );
 a86489a <=( A170  and  a86488a );
 a86492a <=( (not A166)  and  A167 );
 a86495a <=( (not A200)  and  A199 );
 a86496a <=( a86495a  and  a86492a );
 a86497a <=( a86496a  and  a86489a );
 a86500a <=( A202  and  A201 );
 a86503a <=( (not A266)  and  A265 );
 a86504a <=( a86503a  and  a86500a );
 a86507a <=( A268  and  A267 );
 a86510a <=( A299  and  A298 );
 a86511a <=( a86510a  and  a86507a );
 a86512a <=( a86511a  and  a86504a );
 a86516a <=( (not A168)  and  (not A169) );
 a86517a <=( A170  and  a86516a );
 a86520a <=( (not A166)  and  A167 );
 a86523a <=( (not A200)  and  A199 );
 a86524a <=( a86523a  and  a86520a );
 a86525a <=( a86524a  and  a86517a );
 a86528a <=( A202  and  A201 );
 a86531a <=( (not A266)  and  A265 );
 a86532a <=( a86531a  and  a86528a );
 a86535a <=( A268  and  A267 );
 a86538a <=( (not A299)  and  (not A298) );
 a86539a <=( a86538a  and  a86535a );
 a86540a <=( a86539a  and  a86532a );
 a86544a <=( (not A168)  and  (not A169) );
 a86545a <=( A170  and  a86544a );
 a86548a <=( (not A166)  and  A167 );
 a86551a <=( (not A200)  and  A199 );
 a86552a <=( a86551a  and  a86548a );
 a86553a <=( a86552a  and  a86545a );
 a86556a <=( A202  and  A201 );
 a86559a <=( (not A266)  and  A265 );
 a86560a <=( a86559a  and  a86556a );
 a86563a <=( A269  and  A267 );
 a86566a <=( A301  and  (not A300) );
 a86567a <=( a86566a  and  a86563a );
 a86568a <=( a86567a  and  a86560a );
 a86572a <=( (not A168)  and  (not A169) );
 a86573a <=( A170  and  a86572a );
 a86576a <=( (not A166)  and  A167 );
 a86579a <=( (not A200)  and  A199 );
 a86580a <=( a86579a  and  a86576a );
 a86581a <=( a86580a  and  a86573a );
 a86584a <=( A202  and  A201 );
 a86587a <=( (not A266)  and  A265 );
 a86588a <=( a86587a  and  a86584a );
 a86591a <=( A269  and  A267 );
 a86594a <=( A302  and  (not A300) );
 a86595a <=( a86594a  and  a86591a );
 a86596a <=( a86595a  and  a86588a );
 a86600a <=( (not A168)  and  (not A169) );
 a86601a <=( A170  and  a86600a );
 a86604a <=( (not A166)  and  A167 );
 a86607a <=( (not A200)  and  A199 );
 a86608a <=( a86607a  and  a86604a );
 a86609a <=( a86608a  and  a86601a );
 a86612a <=( A202  and  A201 );
 a86615a <=( (not A266)  and  A265 );
 a86616a <=( a86615a  and  a86612a );
 a86619a <=( A269  and  A267 );
 a86622a <=( A299  and  A298 );
 a86623a <=( a86622a  and  a86619a );
 a86624a <=( a86623a  and  a86616a );
 a86628a <=( (not A168)  and  (not A169) );
 a86629a <=( A170  and  a86628a );
 a86632a <=( (not A166)  and  A167 );
 a86635a <=( (not A200)  and  A199 );
 a86636a <=( a86635a  and  a86632a );
 a86637a <=( a86636a  and  a86629a );
 a86640a <=( A202  and  A201 );
 a86643a <=( (not A266)  and  A265 );
 a86644a <=( a86643a  and  a86640a );
 a86647a <=( A269  and  A267 );
 a86650a <=( (not A299)  and  (not A298) );
 a86651a <=( a86650a  and  a86647a );
 a86652a <=( a86651a  and  a86644a );
 a86656a <=( (not A168)  and  (not A169) );
 a86657a <=( A170  and  a86656a );
 a86660a <=( (not A166)  and  A167 );
 a86663a <=( (not A200)  and  A199 );
 a86664a <=( a86663a  and  a86660a );
 a86665a <=( a86664a  and  a86657a );
 a86668a <=( A203  and  A201 );
 a86671a <=( A266  and  (not A265) );
 a86672a <=( a86671a  and  a86668a );
 a86675a <=( A268  and  A267 );
 a86678a <=( A301  and  (not A300) );
 a86679a <=( a86678a  and  a86675a );
 a86680a <=( a86679a  and  a86672a );
 a86684a <=( (not A168)  and  (not A169) );
 a86685a <=( A170  and  a86684a );
 a86688a <=( (not A166)  and  A167 );
 a86691a <=( (not A200)  and  A199 );
 a86692a <=( a86691a  and  a86688a );
 a86693a <=( a86692a  and  a86685a );
 a86696a <=( A203  and  A201 );
 a86699a <=( A266  and  (not A265) );
 a86700a <=( a86699a  and  a86696a );
 a86703a <=( A268  and  A267 );
 a86706a <=( A302  and  (not A300) );
 a86707a <=( a86706a  and  a86703a );
 a86708a <=( a86707a  and  a86700a );
 a86712a <=( (not A168)  and  (not A169) );
 a86713a <=( A170  and  a86712a );
 a86716a <=( (not A166)  and  A167 );
 a86719a <=( (not A200)  and  A199 );
 a86720a <=( a86719a  and  a86716a );
 a86721a <=( a86720a  and  a86713a );
 a86724a <=( A203  and  A201 );
 a86727a <=( A266  and  (not A265) );
 a86728a <=( a86727a  and  a86724a );
 a86731a <=( A268  and  A267 );
 a86734a <=( A299  and  A298 );
 a86735a <=( a86734a  and  a86731a );
 a86736a <=( a86735a  and  a86728a );
 a86740a <=( (not A168)  and  (not A169) );
 a86741a <=( A170  and  a86740a );
 a86744a <=( (not A166)  and  A167 );
 a86747a <=( (not A200)  and  A199 );
 a86748a <=( a86747a  and  a86744a );
 a86749a <=( a86748a  and  a86741a );
 a86752a <=( A203  and  A201 );
 a86755a <=( A266  and  (not A265) );
 a86756a <=( a86755a  and  a86752a );
 a86759a <=( A268  and  A267 );
 a86762a <=( (not A299)  and  (not A298) );
 a86763a <=( a86762a  and  a86759a );
 a86764a <=( a86763a  and  a86756a );
 a86768a <=( (not A168)  and  (not A169) );
 a86769a <=( A170  and  a86768a );
 a86772a <=( (not A166)  and  A167 );
 a86775a <=( (not A200)  and  A199 );
 a86776a <=( a86775a  and  a86772a );
 a86777a <=( a86776a  and  a86769a );
 a86780a <=( A203  and  A201 );
 a86783a <=( A266  and  (not A265) );
 a86784a <=( a86783a  and  a86780a );
 a86787a <=( A269  and  A267 );
 a86790a <=( A301  and  (not A300) );
 a86791a <=( a86790a  and  a86787a );
 a86792a <=( a86791a  and  a86784a );
 a86796a <=( (not A168)  and  (not A169) );
 a86797a <=( A170  and  a86796a );
 a86800a <=( (not A166)  and  A167 );
 a86803a <=( (not A200)  and  A199 );
 a86804a <=( a86803a  and  a86800a );
 a86805a <=( a86804a  and  a86797a );
 a86808a <=( A203  and  A201 );
 a86811a <=( A266  and  (not A265) );
 a86812a <=( a86811a  and  a86808a );
 a86815a <=( A269  and  A267 );
 a86818a <=( A302  and  (not A300) );
 a86819a <=( a86818a  and  a86815a );
 a86820a <=( a86819a  and  a86812a );
 a86824a <=( (not A168)  and  (not A169) );
 a86825a <=( A170  and  a86824a );
 a86828a <=( (not A166)  and  A167 );
 a86831a <=( (not A200)  and  A199 );
 a86832a <=( a86831a  and  a86828a );
 a86833a <=( a86832a  and  a86825a );
 a86836a <=( A203  and  A201 );
 a86839a <=( A266  and  (not A265) );
 a86840a <=( a86839a  and  a86836a );
 a86843a <=( A269  and  A267 );
 a86846a <=( A299  and  A298 );
 a86847a <=( a86846a  and  a86843a );
 a86848a <=( a86847a  and  a86840a );
 a86852a <=( (not A168)  and  (not A169) );
 a86853a <=( A170  and  a86852a );
 a86856a <=( (not A166)  and  A167 );
 a86859a <=( (not A200)  and  A199 );
 a86860a <=( a86859a  and  a86856a );
 a86861a <=( a86860a  and  a86853a );
 a86864a <=( A203  and  A201 );
 a86867a <=( A266  and  (not A265) );
 a86868a <=( a86867a  and  a86864a );
 a86871a <=( A269  and  A267 );
 a86874a <=( (not A299)  and  (not A298) );
 a86875a <=( a86874a  and  a86871a );
 a86876a <=( a86875a  and  a86868a );
 a86880a <=( (not A168)  and  (not A169) );
 a86881a <=( A170  and  a86880a );
 a86884a <=( (not A166)  and  A167 );
 a86887a <=( (not A200)  and  A199 );
 a86888a <=( a86887a  and  a86884a );
 a86889a <=( a86888a  and  a86881a );
 a86892a <=( A203  and  A201 );
 a86895a <=( (not A266)  and  A265 );
 a86896a <=( a86895a  and  a86892a );
 a86899a <=( A268  and  A267 );
 a86902a <=( A301  and  (not A300) );
 a86903a <=( a86902a  and  a86899a );
 a86904a <=( a86903a  and  a86896a );
 a86908a <=( (not A168)  and  (not A169) );
 a86909a <=( A170  and  a86908a );
 a86912a <=( (not A166)  and  A167 );
 a86915a <=( (not A200)  and  A199 );
 a86916a <=( a86915a  and  a86912a );
 a86917a <=( a86916a  and  a86909a );
 a86920a <=( A203  and  A201 );
 a86923a <=( (not A266)  and  A265 );
 a86924a <=( a86923a  and  a86920a );
 a86927a <=( A268  and  A267 );
 a86930a <=( A302  and  (not A300) );
 a86931a <=( a86930a  and  a86927a );
 a86932a <=( a86931a  and  a86924a );
 a86936a <=( (not A168)  and  (not A169) );
 a86937a <=( A170  and  a86936a );
 a86940a <=( (not A166)  and  A167 );
 a86943a <=( (not A200)  and  A199 );
 a86944a <=( a86943a  and  a86940a );
 a86945a <=( a86944a  and  a86937a );
 a86948a <=( A203  and  A201 );
 a86951a <=( (not A266)  and  A265 );
 a86952a <=( a86951a  and  a86948a );
 a86955a <=( A268  and  A267 );
 a86958a <=( A299  and  A298 );
 a86959a <=( a86958a  and  a86955a );
 a86960a <=( a86959a  and  a86952a );
 a86964a <=( (not A168)  and  (not A169) );
 a86965a <=( A170  and  a86964a );
 a86968a <=( (not A166)  and  A167 );
 a86971a <=( (not A200)  and  A199 );
 a86972a <=( a86971a  and  a86968a );
 a86973a <=( a86972a  and  a86965a );
 a86976a <=( A203  and  A201 );
 a86979a <=( (not A266)  and  A265 );
 a86980a <=( a86979a  and  a86976a );
 a86983a <=( A268  and  A267 );
 a86986a <=( (not A299)  and  (not A298) );
 a86987a <=( a86986a  and  a86983a );
 a86988a <=( a86987a  and  a86980a );
 a86992a <=( (not A168)  and  (not A169) );
 a86993a <=( A170  and  a86992a );
 a86996a <=( (not A166)  and  A167 );
 a86999a <=( (not A200)  and  A199 );
 a87000a <=( a86999a  and  a86996a );
 a87001a <=( a87000a  and  a86993a );
 a87004a <=( A203  and  A201 );
 a87007a <=( (not A266)  and  A265 );
 a87008a <=( a87007a  and  a87004a );
 a87011a <=( A269  and  A267 );
 a87014a <=( A301  and  (not A300) );
 a87015a <=( a87014a  and  a87011a );
 a87016a <=( a87015a  and  a87008a );
 a87020a <=( (not A168)  and  (not A169) );
 a87021a <=( A170  and  a87020a );
 a87024a <=( (not A166)  and  A167 );
 a87027a <=( (not A200)  and  A199 );
 a87028a <=( a87027a  and  a87024a );
 a87029a <=( a87028a  and  a87021a );
 a87032a <=( A203  and  A201 );
 a87035a <=( (not A266)  and  A265 );
 a87036a <=( a87035a  and  a87032a );
 a87039a <=( A269  and  A267 );
 a87042a <=( A302  and  (not A300) );
 a87043a <=( a87042a  and  a87039a );
 a87044a <=( a87043a  and  a87036a );
 a87048a <=( (not A168)  and  (not A169) );
 a87049a <=( A170  and  a87048a );
 a87052a <=( (not A166)  and  A167 );
 a87055a <=( (not A200)  and  A199 );
 a87056a <=( a87055a  and  a87052a );
 a87057a <=( a87056a  and  a87049a );
 a87060a <=( A203  and  A201 );
 a87063a <=( (not A266)  and  A265 );
 a87064a <=( a87063a  and  a87060a );
 a87067a <=( A269  and  A267 );
 a87070a <=( A299  and  A298 );
 a87071a <=( a87070a  and  a87067a );
 a87072a <=( a87071a  and  a87064a );
 a87076a <=( (not A168)  and  (not A169) );
 a87077a <=( A170  and  a87076a );
 a87080a <=( (not A166)  and  A167 );
 a87083a <=( (not A200)  and  A199 );
 a87084a <=( a87083a  and  a87080a );
 a87085a <=( a87084a  and  a87077a );
 a87088a <=( A203  and  A201 );
 a87091a <=( (not A266)  and  A265 );
 a87092a <=( a87091a  and  a87088a );
 a87095a <=( A269  and  A267 );
 a87098a <=( (not A299)  and  (not A298) );
 a87099a <=( a87098a  and  a87095a );
 a87100a <=( a87099a  and  a87092a );
 a87104a <=( (not A168)  and  (not A169) );
 a87105a <=( A170  and  a87104a );
 a87108a <=( (not A166)  and  A167 );
 a87111a <=( (not A200)  and  (not A199) );
 a87112a <=( a87111a  and  a87108a );
 a87113a <=( a87112a  and  a87105a );
 a87116a <=( (not A268)  and  A267 );
 a87119a <=( A298  and  (not A269) );
 a87120a <=( a87119a  and  a87116a );
 a87123a <=( (not A300)  and  (not A299) );
 a87126a <=( (not A302)  and  (not A301) );
 a87127a <=( a87126a  and  a87123a );
 a87128a <=( a87127a  and  a87120a );
 a87132a <=( (not A168)  and  (not A169) );
 a87133a <=( A170  and  a87132a );
 a87136a <=( (not A166)  and  A167 );
 a87139a <=( (not A200)  and  (not A199) );
 a87140a <=( a87139a  and  a87136a );
 a87141a <=( a87140a  and  a87133a );
 a87144a <=( (not A268)  and  A267 );
 a87147a <=( (not A298)  and  (not A269) );
 a87148a <=( a87147a  and  a87144a );
 a87151a <=( (not A300)  and  A299 );
 a87154a <=( (not A302)  and  (not A301) );
 a87155a <=( a87154a  and  a87151a );
 a87156a <=( a87155a  and  a87148a );
 a87160a <=( (not A168)  and  (not A169) );
 a87161a <=( A170  and  a87160a );
 a87164a <=( A166  and  (not A167) );
 a87167a <=( (not A202)  and  A201 );
 a87168a <=( a87167a  and  a87164a );
 a87169a <=( a87168a  and  a87161a );
 a87172a <=( A267  and  (not A203) );
 a87175a <=( (not A269)  and  (not A268) );
 a87176a <=( a87175a  and  a87172a );
 a87179a <=( (not A299)  and  A298 );
 a87182a <=( A301  and  A300 );
 a87183a <=( a87182a  and  a87179a );
 a87184a <=( a87183a  and  a87176a );
 a87188a <=( (not A168)  and  (not A169) );
 a87189a <=( A170  and  a87188a );
 a87192a <=( A166  and  (not A167) );
 a87195a <=( (not A202)  and  A201 );
 a87196a <=( a87195a  and  a87192a );
 a87197a <=( a87196a  and  a87189a );
 a87200a <=( A267  and  (not A203) );
 a87203a <=( (not A269)  and  (not A268) );
 a87204a <=( a87203a  and  a87200a );
 a87207a <=( (not A299)  and  A298 );
 a87210a <=( A302  and  A300 );
 a87211a <=( a87210a  and  a87207a );
 a87212a <=( a87211a  and  a87204a );
 a87216a <=( (not A168)  and  (not A169) );
 a87217a <=( A170  and  a87216a );
 a87220a <=( A166  and  (not A167) );
 a87223a <=( (not A202)  and  A201 );
 a87224a <=( a87223a  and  a87220a );
 a87225a <=( a87224a  and  a87217a );
 a87228a <=( A267  and  (not A203) );
 a87231a <=( (not A269)  and  (not A268) );
 a87232a <=( a87231a  and  a87228a );
 a87235a <=( A299  and  (not A298) );
 a87238a <=( A301  and  A300 );
 a87239a <=( a87238a  and  a87235a );
 a87240a <=( a87239a  and  a87232a );
 a87244a <=( (not A168)  and  (not A169) );
 a87245a <=( A170  and  a87244a );
 a87248a <=( A166  and  (not A167) );
 a87251a <=( (not A202)  and  A201 );
 a87252a <=( a87251a  and  a87248a );
 a87253a <=( a87252a  and  a87245a );
 a87256a <=( A267  and  (not A203) );
 a87259a <=( (not A269)  and  (not A268) );
 a87260a <=( a87259a  and  a87256a );
 a87263a <=( A299  and  (not A298) );
 a87266a <=( A302  and  A300 );
 a87267a <=( a87266a  and  a87263a );
 a87268a <=( a87267a  and  a87260a );
 a87272a <=( (not A168)  and  (not A169) );
 a87273a <=( A170  and  a87272a );
 a87276a <=( A166  and  (not A167) );
 a87279a <=( (not A202)  and  A201 );
 a87280a <=( a87279a  and  a87276a );
 a87281a <=( a87280a  and  a87273a );
 a87284a <=( (not A267)  and  (not A203) );
 a87287a <=( A298  and  A268 );
 a87288a <=( a87287a  and  a87284a );
 a87291a <=( (not A300)  and  (not A299) );
 a87294a <=( (not A302)  and  (not A301) );
 a87295a <=( a87294a  and  a87291a );
 a87296a <=( a87295a  and  a87288a );
 a87300a <=( (not A168)  and  (not A169) );
 a87301a <=( A170  and  a87300a );
 a87304a <=( A166  and  (not A167) );
 a87307a <=( (not A202)  and  A201 );
 a87308a <=( a87307a  and  a87304a );
 a87309a <=( a87308a  and  a87301a );
 a87312a <=( (not A267)  and  (not A203) );
 a87315a <=( (not A298)  and  A268 );
 a87316a <=( a87315a  and  a87312a );
 a87319a <=( (not A300)  and  A299 );
 a87322a <=( (not A302)  and  (not A301) );
 a87323a <=( a87322a  and  a87319a );
 a87324a <=( a87323a  and  a87316a );
 a87328a <=( (not A168)  and  (not A169) );
 a87329a <=( A170  and  a87328a );
 a87332a <=( A166  and  (not A167) );
 a87335a <=( (not A202)  and  A201 );
 a87336a <=( a87335a  and  a87332a );
 a87337a <=( a87336a  and  a87329a );
 a87340a <=( (not A267)  and  (not A203) );
 a87343a <=( A298  and  A269 );
 a87344a <=( a87343a  and  a87340a );
 a87347a <=( (not A300)  and  (not A299) );
 a87350a <=( (not A302)  and  (not A301) );
 a87351a <=( a87350a  and  a87347a );
 a87352a <=( a87351a  and  a87344a );
 a87356a <=( (not A168)  and  (not A169) );
 a87357a <=( A170  and  a87356a );
 a87360a <=( A166  and  (not A167) );
 a87363a <=( (not A202)  and  A201 );
 a87364a <=( a87363a  and  a87360a );
 a87365a <=( a87364a  and  a87357a );
 a87368a <=( (not A267)  and  (not A203) );
 a87371a <=( (not A298)  and  A269 );
 a87372a <=( a87371a  and  a87368a );
 a87375a <=( (not A300)  and  A299 );
 a87378a <=( (not A302)  and  (not A301) );
 a87379a <=( a87378a  and  a87375a );
 a87380a <=( a87379a  and  a87372a );
 a87384a <=( (not A168)  and  (not A169) );
 a87385a <=( A170  and  a87384a );
 a87388a <=( A166  and  (not A167) );
 a87391a <=( (not A202)  and  A201 );
 a87392a <=( a87391a  and  a87388a );
 a87393a <=( a87392a  and  a87385a );
 a87396a <=( A265  and  (not A203) );
 a87399a <=( A298  and  A266 );
 a87400a <=( a87399a  and  a87396a );
 a87403a <=( (not A300)  and  (not A299) );
 a87406a <=( (not A302)  and  (not A301) );
 a87407a <=( a87406a  and  a87403a );
 a87408a <=( a87407a  and  a87400a );
 a87412a <=( (not A168)  and  (not A169) );
 a87413a <=( A170  and  a87412a );
 a87416a <=( A166  and  (not A167) );
 a87419a <=( (not A202)  and  A201 );
 a87420a <=( a87419a  and  a87416a );
 a87421a <=( a87420a  and  a87413a );
 a87424a <=( A265  and  (not A203) );
 a87427a <=( (not A298)  and  A266 );
 a87428a <=( a87427a  and  a87424a );
 a87431a <=( (not A300)  and  A299 );
 a87434a <=( (not A302)  and  (not A301) );
 a87435a <=( a87434a  and  a87431a );
 a87436a <=( a87435a  and  a87428a );
 a87440a <=( (not A168)  and  (not A169) );
 a87441a <=( A170  and  a87440a );
 a87444a <=( A166  and  (not A167) );
 a87447a <=( (not A202)  and  A201 );
 a87448a <=( a87447a  and  a87444a );
 a87449a <=( a87448a  and  a87441a );
 a87452a <=( (not A265)  and  (not A203) );
 a87455a <=( A298  and  (not A266) );
 a87456a <=( a87455a  and  a87452a );
 a87459a <=( (not A300)  and  (not A299) );
 a87462a <=( (not A302)  and  (not A301) );
 a87463a <=( a87462a  and  a87459a );
 a87464a <=( a87463a  and  a87456a );
 a87468a <=( (not A168)  and  (not A169) );
 a87469a <=( A170  and  a87468a );
 a87472a <=( A166  and  (not A167) );
 a87475a <=( (not A202)  and  A201 );
 a87476a <=( a87475a  and  a87472a );
 a87477a <=( a87476a  and  a87469a );
 a87480a <=( (not A265)  and  (not A203) );
 a87483a <=( (not A298)  and  (not A266) );
 a87484a <=( a87483a  and  a87480a );
 a87487a <=( (not A300)  and  A299 );
 a87490a <=( (not A302)  and  (not A301) );
 a87491a <=( a87490a  and  a87487a );
 a87492a <=( a87491a  and  a87484a );
 a87496a <=( (not A168)  and  (not A169) );
 a87497a <=( A170  and  a87496a );
 a87500a <=( A166  and  (not A167) );
 a87503a <=( A202  and  (not A201) );
 a87504a <=( a87503a  and  a87500a );
 a87505a <=( a87504a  and  a87497a );
 a87508a <=( (not A268)  and  A267 );
 a87511a <=( A298  and  (not A269) );
 a87512a <=( a87511a  and  a87508a );
 a87515a <=( (not A300)  and  (not A299) );
 a87518a <=( (not A302)  and  (not A301) );
 a87519a <=( a87518a  and  a87515a );
 a87520a <=( a87519a  and  a87512a );
 a87524a <=( (not A168)  and  (not A169) );
 a87525a <=( A170  and  a87524a );
 a87528a <=( A166  and  (not A167) );
 a87531a <=( A202  and  (not A201) );
 a87532a <=( a87531a  and  a87528a );
 a87533a <=( a87532a  and  a87525a );
 a87536a <=( (not A268)  and  A267 );
 a87539a <=( (not A298)  and  (not A269) );
 a87540a <=( a87539a  and  a87536a );
 a87543a <=( (not A300)  and  A299 );
 a87546a <=( (not A302)  and  (not A301) );
 a87547a <=( a87546a  and  a87543a );
 a87548a <=( a87547a  and  a87540a );
 a87552a <=( (not A168)  and  (not A169) );
 a87553a <=( A170  and  a87552a );
 a87556a <=( A166  and  (not A167) );
 a87559a <=( A203  and  (not A201) );
 a87560a <=( a87559a  and  a87556a );
 a87561a <=( a87560a  and  a87553a );
 a87564a <=( (not A268)  and  A267 );
 a87567a <=( A298  and  (not A269) );
 a87568a <=( a87567a  and  a87564a );
 a87571a <=( (not A300)  and  (not A299) );
 a87574a <=( (not A302)  and  (not A301) );
 a87575a <=( a87574a  and  a87571a );
 a87576a <=( a87575a  and  a87568a );
 a87580a <=( (not A168)  and  (not A169) );
 a87581a <=( A170  and  a87580a );
 a87584a <=( A166  and  (not A167) );
 a87587a <=( A203  and  (not A201) );
 a87588a <=( a87587a  and  a87584a );
 a87589a <=( a87588a  and  a87581a );
 a87592a <=( (not A268)  and  A267 );
 a87595a <=( (not A298)  and  (not A269) );
 a87596a <=( a87595a  and  a87592a );
 a87599a <=( (not A300)  and  A299 );
 a87602a <=( (not A302)  and  (not A301) );
 a87603a <=( a87602a  and  a87599a );
 a87604a <=( a87603a  and  a87596a );
 a87608a <=( (not A168)  and  (not A169) );
 a87609a <=( A170  and  a87608a );
 a87612a <=( A166  and  (not A167) );
 a87615a <=( A200  and  A199 );
 a87616a <=( a87615a  and  a87612a );
 a87617a <=( a87616a  and  a87609a );
 a87620a <=( (not A268)  and  A267 );
 a87623a <=( A298  and  (not A269) );
 a87624a <=( a87623a  and  a87620a );
 a87627a <=( (not A300)  and  (not A299) );
 a87630a <=( (not A302)  and  (not A301) );
 a87631a <=( a87630a  and  a87627a );
 a87632a <=( a87631a  and  a87624a );
 a87636a <=( (not A168)  and  (not A169) );
 a87637a <=( A170  and  a87636a );
 a87640a <=( A166  and  (not A167) );
 a87643a <=( A200  and  A199 );
 a87644a <=( a87643a  and  a87640a );
 a87645a <=( a87644a  and  a87637a );
 a87648a <=( (not A268)  and  A267 );
 a87651a <=( (not A298)  and  (not A269) );
 a87652a <=( a87651a  and  a87648a );
 a87655a <=( (not A300)  and  A299 );
 a87658a <=( (not A302)  and  (not A301) );
 a87659a <=( a87658a  and  a87655a );
 a87660a <=( a87659a  and  a87652a );
 a87664a <=( (not A168)  and  (not A169) );
 a87665a <=( A170  and  a87664a );
 a87668a <=( A166  and  (not A167) );
 a87671a <=( A200  and  (not A199) );
 a87672a <=( a87671a  and  a87668a );
 a87673a <=( a87672a  and  a87665a );
 a87676a <=( A202  and  A201 );
 a87679a <=( A266  and  (not A265) );
 a87680a <=( a87679a  and  a87676a );
 a87683a <=( A268  and  A267 );
 a87686a <=( A301  and  (not A300) );
 a87687a <=( a87686a  and  a87683a );
 a87688a <=( a87687a  and  a87680a );
 a87692a <=( (not A168)  and  (not A169) );
 a87693a <=( A170  and  a87692a );
 a87696a <=( A166  and  (not A167) );
 a87699a <=( A200  and  (not A199) );
 a87700a <=( a87699a  and  a87696a );
 a87701a <=( a87700a  and  a87693a );
 a87704a <=( A202  and  A201 );
 a87707a <=( A266  and  (not A265) );
 a87708a <=( a87707a  and  a87704a );
 a87711a <=( A268  and  A267 );
 a87714a <=( A302  and  (not A300) );
 a87715a <=( a87714a  and  a87711a );
 a87716a <=( a87715a  and  a87708a );
 a87720a <=( (not A168)  and  (not A169) );
 a87721a <=( A170  and  a87720a );
 a87724a <=( A166  and  (not A167) );
 a87727a <=( A200  and  (not A199) );
 a87728a <=( a87727a  and  a87724a );
 a87729a <=( a87728a  and  a87721a );
 a87732a <=( A202  and  A201 );
 a87735a <=( A266  and  (not A265) );
 a87736a <=( a87735a  and  a87732a );
 a87739a <=( A268  and  A267 );
 a87742a <=( A299  and  A298 );
 a87743a <=( a87742a  and  a87739a );
 a87744a <=( a87743a  and  a87736a );
 a87748a <=( (not A168)  and  (not A169) );
 a87749a <=( A170  and  a87748a );
 a87752a <=( A166  and  (not A167) );
 a87755a <=( A200  and  (not A199) );
 a87756a <=( a87755a  and  a87752a );
 a87757a <=( a87756a  and  a87749a );
 a87760a <=( A202  and  A201 );
 a87763a <=( A266  and  (not A265) );
 a87764a <=( a87763a  and  a87760a );
 a87767a <=( A268  and  A267 );
 a87770a <=( (not A299)  and  (not A298) );
 a87771a <=( a87770a  and  a87767a );
 a87772a <=( a87771a  and  a87764a );
 a87776a <=( (not A168)  and  (not A169) );
 a87777a <=( A170  and  a87776a );
 a87780a <=( A166  and  (not A167) );
 a87783a <=( A200  and  (not A199) );
 a87784a <=( a87783a  and  a87780a );
 a87785a <=( a87784a  and  a87777a );
 a87788a <=( A202  and  A201 );
 a87791a <=( A266  and  (not A265) );
 a87792a <=( a87791a  and  a87788a );
 a87795a <=( A269  and  A267 );
 a87798a <=( A301  and  (not A300) );
 a87799a <=( a87798a  and  a87795a );
 a87800a <=( a87799a  and  a87792a );
 a87804a <=( (not A168)  and  (not A169) );
 a87805a <=( A170  and  a87804a );
 a87808a <=( A166  and  (not A167) );
 a87811a <=( A200  and  (not A199) );
 a87812a <=( a87811a  and  a87808a );
 a87813a <=( a87812a  and  a87805a );
 a87816a <=( A202  and  A201 );
 a87819a <=( A266  and  (not A265) );
 a87820a <=( a87819a  and  a87816a );
 a87823a <=( A269  and  A267 );
 a87826a <=( A302  and  (not A300) );
 a87827a <=( a87826a  and  a87823a );
 a87828a <=( a87827a  and  a87820a );
 a87832a <=( (not A168)  and  (not A169) );
 a87833a <=( A170  and  a87832a );
 a87836a <=( A166  and  (not A167) );
 a87839a <=( A200  and  (not A199) );
 a87840a <=( a87839a  and  a87836a );
 a87841a <=( a87840a  and  a87833a );
 a87844a <=( A202  and  A201 );
 a87847a <=( A266  and  (not A265) );
 a87848a <=( a87847a  and  a87844a );
 a87851a <=( A269  and  A267 );
 a87854a <=( A299  and  A298 );
 a87855a <=( a87854a  and  a87851a );
 a87856a <=( a87855a  and  a87848a );
 a87860a <=( (not A168)  and  (not A169) );
 a87861a <=( A170  and  a87860a );
 a87864a <=( A166  and  (not A167) );
 a87867a <=( A200  and  (not A199) );
 a87868a <=( a87867a  and  a87864a );
 a87869a <=( a87868a  and  a87861a );
 a87872a <=( A202  and  A201 );
 a87875a <=( A266  and  (not A265) );
 a87876a <=( a87875a  and  a87872a );
 a87879a <=( A269  and  A267 );
 a87882a <=( (not A299)  and  (not A298) );
 a87883a <=( a87882a  and  a87879a );
 a87884a <=( a87883a  and  a87876a );
 a87888a <=( (not A168)  and  (not A169) );
 a87889a <=( A170  and  a87888a );
 a87892a <=( A166  and  (not A167) );
 a87895a <=( A200  and  (not A199) );
 a87896a <=( a87895a  and  a87892a );
 a87897a <=( a87896a  and  a87889a );
 a87900a <=( A202  and  A201 );
 a87903a <=( (not A266)  and  A265 );
 a87904a <=( a87903a  and  a87900a );
 a87907a <=( A268  and  A267 );
 a87910a <=( A301  and  (not A300) );
 a87911a <=( a87910a  and  a87907a );
 a87912a <=( a87911a  and  a87904a );
 a87916a <=( (not A168)  and  (not A169) );
 a87917a <=( A170  and  a87916a );
 a87920a <=( A166  and  (not A167) );
 a87923a <=( A200  and  (not A199) );
 a87924a <=( a87923a  and  a87920a );
 a87925a <=( a87924a  and  a87917a );
 a87928a <=( A202  and  A201 );
 a87931a <=( (not A266)  and  A265 );
 a87932a <=( a87931a  and  a87928a );
 a87935a <=( A268  and  A267 );
 a87938a <=( A302  and  (not A300) );
 a87939a <=( a87938a  and  a87935a );
 a87940a <=( a87939a  and  a87932a );
 a87944a <=( (not A168)  and  (not A169) );
 a87945a <=( A170  and  a87944a );
 a87948a <=( A166  and  (not A167) );
 a87951a <=( A200  and  (not A199) );
 a87952a <=( a87951a  and  a87948a );
 a87953a <=( a87952a  and  a87945a );
 a87956a <=( A202  and  A201 );
 a87959a <=( (not A266)  and  A265 );
 a87960a <=( a87959a  and  a87956a );
 a87963a <=( A268  and  A267 );
 a87966a <=( A299  and  A298 );
 a87967a <=( a87966a  and  a87963a );
 a87968a <=( a87967a  and  a87960a );
 a87972a <=( (not A168)  and  (not A169) );
 a87973a <=( A170  and  a87972a );
 a87976a <=( A166  and  (not A167) );
 a87979a <=( A200  and  (not A199) );
 a87980a <=( a87979a  and  a87976a );
 a87981a <=( a87980a  and  a87973a );
 a87984a <=( A202  and  A201 );
 a87987a <=( (not A266)  and  A265 );
 a87988a <=( a87987a  and  a87984a );
 a87991a <=( A268  and  A267 );
 a87994a <=( (not A299)  and  (not A298) );
 a87995a <=( a87994a  and  a87991a );
 a87996a <=( a87995a  and  a87988a );
 a88000a <=( (not A168)  and  (not A169) );
 a88001a <=( A170  and  a88000a );
 a88004a <=( A166  and  (not A167) );
 a88007a <=( A200  and  (not A199) );
 a88008a <=( a88007a  and  a88004a );
 a88009a <=( a88008a  and  a88001a );
 a88012a <=( A202  and  A201 );
 a88015a <=( (not A266)  and  A265 );
 a88016a <=( a88015a  and  a88012a );
 a88019a <=( A269  and  A267 );
 a88022a <=( A301  and  (not A300) );
 a88023a <=( a88022a  and  a88019a );
 a88024a <=( a88023a  and  a88016a );
 a88028a <=( (not A168)  and  (not A169) );
 a88029a <=( A170  and  a88028a );
 a88032a <=( A166  and  (not A167) );
 a88035a <=( A200  and  (not A199) );
 a88036a <=( a88035a  and  a88032a );
 a88037a <=( a88036a  and  a88029a );
 a88040a <=( A202  and  A201 );
 a88043a <=( (not A266)  and  A265 );
 a88044a <=( a88043a  and  a88040a );
 a88047a <=( A269  and  A267 );
 a88050a <=( A302  and  (not A300) );
 a88051a <=( a88050a  and  a88047a );
 a88052a <=( a88051a  and  a88044a );
 a88056a <=( (not A168)  and  (not A169) );
 a88057a <=( A170  and  a88056a );
 a88060a <=( A166  and  (not A167) );
 a88063a <=( A200  and  (not A199) );
 a88064a <=( a88063a  and  a88060a );
 a88065a <=( a88064a  and  a88057a );
 a88068a <=( A202  and  A201 );
 a88071a <=( (not A266)  and  A265 );
 a88072a <=( a88071a  and  a88068a );
 a88075a <=( A269  and  A267 );
 a88078a <=( A299  and  A298 );
 a88079a <=( a88078a  and  a88075a );
 a88080a <=( a88079a  and  a88072a );
 a88084a <=( (not A168)  and  (not A169) );
 a88085a <=( A170  and  a88084a );
 a88088a <=( A166  and  (not A167) );
 a88091a <=( A200  and  (not A199) );
 a88092a <=( a88091a  and  a88088a );
 a88093a <=( a88092a  and  a88085a );
 a88096a <=( A202  and  A201 );
 a88099a <=( (not A266)  and  A265 );
 a88100a <=( a88099a  and  a88096a );
 a88103a <=( A269  and  A267 );
 a88106a <=( (not A299)  and  (not A298) );
 a88107a <=( a88106a  and  a88103a );
 a88108a <=( a88107a  and  a88100a );
 a88112a <=( (not A168)  and  (not A169) );
 a88113a <=( A170  and  a88112a );
 a88116a <=( A166  and  (not A167) );
 a88119a <=( A200  and  (not A199) );
 a88120a <=( a88119a  and  a88116a );
 a88121a <=( a88120a  and  a88113a );
 a88124a <=( A203  and  A201 );
 a88127a <=( A266  and  (not A265) );
 a88128a <=( a88127a  and  a88124a );
 a88131a <=( A268  and  A267 );
 a88134a <=( A301  and  (not A300) );
 a88135a <=( a88134a  and  a88131a );
 a88136a <=( a88135a  and  a88128a );
 a88140a <=( (not A168)  and  (not A169) );
 a88141a <=( A170  and  a88140a );
 a88144a <=( A166  and  (not A167) );
 a88147a <=( A200  and  (not A199) );
 a88148a <=( a88147a  and  a88144a );
 a88149a <=( a88148a  and  a88141a );
 a88152a <=( A203  and  A201 );
 a88155a <=( A266  and  (not A265) );
 a88156a <=( a88155a  and  a88152a );
 a88159a <=( A268  and  A267 );
 a88162a <=( A302  and  (not A300) );
 a88163a <=( a88162a  and  a88159a );
 a88164a <=( a88163a  and  a88156a );
 a88168a <=( (not A168)  and  (not A169) );
 a88169a <=( A170  and  a88168a );
 a88172a <=( A166  and  (not A167) );
 a88175a <=( A200  and  (not A199) );
 a88176a <=( a88175a  and  a88172a );
 a88177a <=( a88176a  and  a88169a );
 a88180a <=( A203  and  A201 );
 a88183a <=( A266  and  (not A265) );
 a88184a <=( a88183a  and  a88180a );
 a88187a <=( A268  and  A267 );
 a88190a <=( A299  and  A298 );
 a88191a <=( a88190a  and  a88187a );
 a88192a <=( a88191a  and  a88184a );
 a88196a <=( (not A168)  and  (not A169) );
 a88197a <=( A170  and  a88196a );
 a88200a <=( A166  and  (not A167) );
 a88203a <=( A200  and  (not A199) );
 a88204a <=( a88203a  and  a88200a );
 a88205a <=( a88204a  and  a88197a );
 a88208a <=( A203  and  A201 );
 a88211a <=( A266  and  (not A265) );
 a88212a <=( a88211a  and  a88208a );
 a88215a <=( A268  and  A267 );
 a88218a <=( (not A299)  and  (not A298) );
 a88219a <=( a88218a  and  a88215a );
 a88220a <=( a88219a  and  a88212a );
 a88224a <=( (not A168)  and  (not A169) );
 a88225a <=( A170  and  a88224a );
 a88228a <=( A166  and  (not A167) );
 a88231a <=( A200  and  (not A199) );
 a88232a <=( a88231a  and  a88228a );
 a88233a <=( a88232a  and  a88225a );
 a88236a <=( A203  and  A201 );
 a88239a <=( A266  and  (not A265) );
 a88240a <=( a88239a  and  a88236a );
 a88243a <=( A269  and  A267 );
 a88246a <=( A301  and  (not A300) );
 a88247a <=( a88246a  and  a88243a );
 a88248a <=( a88247a  and  a88240a );
 a88252a <=( (not A168)  and  (not A169) );
 a88253a <=( A170  and  a88252a );
 a88256a <=( A166  and  (not A167) );
 a88259a <=( A200  and  (not A199) );
 a88260a <=( a88259a  and  a88256a );
 a88261a <=( a88260a  and  a88253a );
 a88264a <=( A203  and  A201 );
 a88267a <=( A266  and  (not A265) );
 a88268a <=( a88267a  and  a88264a );
 a88271a <=( A269  and  A267 );
 a88274a <=( A302  and  (not A300) );
 a88275a <=( a88274a  and  a88271a );
 a88276a <=( a88275a  and  a88268a );
 a88280a <=( (not A168)  and  (not A169) );
 a88281a <=( A170  and  a88280a );
 a88284a <=( A166  and  (not A167) );
 a88287a <=( A200  and  (not A199) );
 a88288a <=( a88287a  and  a88284a );
 a88289a <=( a88288a  and  a88281a );
 a88292a <=( A203  and  A201 );
 a88295a <=( A266  and  (not A265) );
 a88296a <=( a88295a  and  a88292a );
 a88299a <=( A269  and  A267 );
 a88302a <=( A299  and  A298 );
 a88303a <=( a88302a  and  a88299a );
 a88304a <=( a88303a  and  a88296a );
 a88308a <=( (not A168)  and  (not A169) );
 a88309a <=( A170  and  a88308a );
 a88312a <=( A166  and  (not A167) );
 a88315a <=( A200  and  (not A199) );
 a88316a <=( a88315a  and  a88312a );
 a88317a <=( a88316a  and  a88309a );
 a88320a <=( A203  and  A201 );
 a88323a <=( A266  and  (not A265) );
 a88324a <=( a88323a  and  a88320a );
 a88327a <=( A269  and  A267 );
 a88330a <=( (not A299)  and  (not A298) );
 a88331a <=( a88330a  and  a88327a );
 a88332a <=( a88331a  and  a88324a );
 a88336a <=( (not A168)  and  (not A169) );
 a88337a <=( A170  and  a88336a );
 a88340a <=( A166  and  (not A167) );
 a88343a <=( A200  and  (not A199) );
 a88344a <=( a88343a  and  a88340a );
 a88345a <=( a88344a  and  a88337a );
 a88348a <=( A203  and  A201 );
 a88351a <=( (not A266)  and  A265 );
 a88352a <=( a88351a  and  a88348a );
 a88355a <=( A268  and  A267 );
 a88358a <=( A301  and  (not A300) );
 a88359a <=( a88358a  and  a88355a );
 a88360a <=( a88359a  and  a88352a );
 a88364a <=( (not A168)  and  (not A169) );
 a88365a <=( A170  and  a88364a );
 a88368a <=( A166  and  (not A167) );
 a88371a <=( A200  and  (not A199) );
 a88372a <=( a88371a  and  a88368a );
 a88373a <=( a88372a  and  a88365a );
 a88376a <=( A203  and  A201 );
 a88379a <=( (not A266)  and  A265 );
 a88380a <=( a88379a  and  a88376a );
 a88383a <=( A268  and  A267 );
 a88386a <=( A302  and  (not A300) );
 a88387a <=( a88386a  and  a88383a );
 a88388a <=( a88387a  and  a88380a );
 a88392a <=( (not A168)  and  (not A169) );
 a88393a <=( A170  and  a88392a );
 a88396a <=( A166  and  (not A167) );
 a88399a <=( A200  and  (not A199) );
 a88400a <=( a88399a  and  a88396a );
 a88401a <=( a88400a  and  a88393a );
 a88404a <=( A203  and  A201 );
 a88407a <=( (not A266)  and  A265 );
 a88408a <=( a88407a  and  a88404a );
 a88411a <=( A268  and  A267 );
 a88414a <=( A299  and  A298 );
 a88415a <=( a88414a  and  a88411a );
 a88416a <=( a88415a  and  a88408a );
 a88420a <=( (not A168)  and  (not A169) );
 a88421a <=( A170  and  a88420a );
 a88424a <=( A166  and  (not A167) );
 a88427a <=( A200  and  (not A199) );
 a88428a <=( a88427a  and  a88424a );
 a88429a <=( a88428a  and  a88421a );
 a88432a <=( A203  and  A201 );
 a88435a <=( (not A266)  and  A265 );
 a88436a <=( a88435a  and  a88432a );
 a88439a <=( A268  and  A267 );
 a88442a <=( (not A299)  and  (not A298) );
 a88443a <=( a88442a  and  a88439a );
 a88444a <=( a88443a  and  a88436a );
 a88448a <=( (not A168)  and  (not A169) );
 a88449a <=( A170  and  a88448a );
 a88452a <=( A166  and  (not A167) );
 a88455a <=( A200  and  (not A199) );
 a88456a <=( a88455a  and  a88452a );
 a88457a <=( a88456a  and  a88449a );
 a88460a <=( A203  and  A201 );
 a88463a <=( (not A266)  and  A265 );
 a88464a <=( a88463a  and  a88460a );
 a88467a <=( A269  and  A267 );
 a88470a <=( A301  and  (not A300) );
 a88471a <=( a88470a  and  a88467a );
 a88472a <=( a88471a  and  a88464a );
 a88476a <=( (not A168)  and  (not A169) );
 a88477a <=( A170  and  a88476a );
 a88480a <=( A166  and  (not A167) );
 a88483a <=( A200  and  (not A199) );
 a88484a <=( a88483a  and  a88480a );
 a88485a <=( a88484a  and  a88477a );
 a88488a <=( A203  and  A201 );
 a88491a <=( (not A266)  and  A265 );
 a88492a <=( a88491a  and  a88488a );
 a88495a <=( A269  and  A267 );
 a88498a <=( A302  and  (not A300) );
 a88499a <=( a88498a  and  a88495a );
 a88500a <=( a88499a  and  a88492a );
 a88504a <=( (not A168)  and  (not A169) );
 a88505a <=( A170  and  a88504a );
 a88508a <=( A166  and  (not A167) );
 a88511a <=( A200  and  (not A199) );
 a88512a <=( a88511a  and  a88508a );
 a88513a <=( a88512a  and  a88505a );
 a88516a <=( A203  and  A201 );
 a88519a <=( (not A266)  and  A265 );
 a88520a <=( a88519a  and  a88516a );
 a88523a <=( A269  and  A267 );
 a88526a <=( A299  and  A298 );
 a88527a <=( a88526a  and  a88523a );
 a88528a <=( a88527a  and  a88520a );
 a88532a <=( (not A168)  and  (not A169) );
 a88533a <=( A170  and  a88532a );
 a88536a <=( A166  and  (not A167) );
 a88539a <=( A200  and  (not A199) );
 a88540a <=( a88539a  and  a88536a );
 a88541a <=( a88540a  and  a88533a );
 a88544a <=( A203  and  A201 );
 a88547a <=( (not A266)  and  A265 );
 a88548a <=( a88547a  and  a88544a );
 a88551a <=( A269  and  A267 );
 a88554a <=( (not A299)  and  (not A298) );
 a88555a <=( a88554a  and  a88551a );
 a88556a <=( a88555a  and  a88548a );
 a88560a <=( (not A168)  and  (not A169) );
 a88561a <=( A170  and  a88560a );
 a88564a <=( A166  and  (not A167) );
 a88567a <=( (not A200)  and  A199 );
 a88568a <=( a88567a  and  a88564a );
 a88569a <=( a88568a  and  a88561a );
 a88572a <=( A202  and  A201 );
 a88575a <=( A266  and  (not A265) );
 a88576a <=( a88575a  and  a88572a );
 a88579a <=( A268  and  A267 );
 a88582a <=( A301  and  (not A300) );
 a88583a <=( a88582a  and  a88579a );
 a88584a <=( a88583a  and  a88576a );
 a88588a <=( (not A168)  and  (not A169) );
 a88589a <=( A170  and  a88588a );
 a88592a <=( A166  and  (not A167) );
 a88595a <=( (not A200)  and  A199 );
 a88596a <=( a88595a  and  a88592a );
 a88597a <=( a88596a  and  a88589a );
 a88600a <=( A202  and  A201 );
 a88603a <=( A266  and  (not A265) );
 a88604a <=( a88603a  and  a88600a );
 a88607a <=( A268  and  A267 );
 a88610a <=( A302  and  (not A300) );
 a88611a <=( a88610a  and  a88607a );
 a88612a <=( a88611a  and  a88604a );
 a88616a <=( (not A168)  and  (not A169) );
 a88617a <=( A170  and  a88616a );
 a88620a <=( A166  and  (not A167) );
 a88623a <=( (not A200)  and  A199 );
 a88624a <=( a88623a  and  a88620a );
 a88625a <=( a88624a  and  a88617a );
 a88628a <=( A202  and  A201 );
 a88631a <=( A266  and  (not A265) );
 a88632a <=( a88631a  and  a88628a );
 a88635a <=( A268  and  A267 );
 a88638a <=( A299  and  A298 );
 a88639a <=( a88638a  and  a88635a );
 a88640a <=( a88639a  and  a88632a );
 a88644a <=( (not A168)  and  (not A169) );
 a88645a <=( A170  and  a88644a );
 a88648a <=( A166  and  (not A167) );
 a88651a <=( (not A200)  and  A199 );
 a88652a <=( a88651a  and  a88648a );
 a88653a <=( a88652a  and  a88645a );
 a88656a <=( A202  and  A201 );
 a88659a <=( A266  and  (not A265) );
 a88660a <=( a88659a  and  a88656a );
 a88663a <=( A268  and  A267 );
 a88666a <=( (not A299)  and  (not A298) );
 a88667a <=( a88666a  and  a88663a );
 a88668a <=( a88667a  and  a88660a );
 a88672a <=( (not A168)  and  (not A169) );
 a88673a <=( A170  and  a88672a );
 a88676a <=( A166  and  (not A167) );
 a88679a <=( (not A200)  and  A199 );
 a88680a <=( a88679a  and  a88676a );
 a88681a <=( a88680a  and  a88673a );
 a88684a <=( A202  and  A201 );
 a88687a <=( A266  and  (not A265) );
 a88688a <=( a88687a  and  a88684a );
 a88691a <=( A269  and  A267 );
 a88694a <=( A301  and  (not A300) );
 a88695a <=( a88694a  and  a88691a );
 a88696a <=( a88695a  and  a88688a );
 a88700a <=( (not A168)  and  (not A169) );
 a88701a <=( A170  and  a88700a );
 a88704a <=( A166  and  (not A167) );
 a88707a <=( (not A200)  and  A199 );
 a88708a <=( a88707a  and  a88704a );
 a88709a <=( a88708a  and  a88701a );
 a88712a <=( A202  and  A201 );
 a88715a <=( A266  and  (not A265) );
 a88716a <=( a88715a  and  a88712a );
 a88719a <=( A269  and  A267 );
 a88722a <=( A302  and  (not A300) );
 a88723a <=( a88722a  and  a88719a );
 a88724a <=( a88723a  and  a88716a );
 a88728a <=( (not A168)  and  (not A169) );
 a88729a <=( A170  and  a88728a );
 a88732a <=( A166  and  (not A167) );
 a88735a <=( (not A200)  and  A199 );
 a88736a <=( a88735a  and  a88732a );
 a88737a <=( a88736a  and  a88729a );
 a88740a <=( A202  and  A201 );
 a88743a <=( A266  and  (not A265) );
 a88744a <=( a88743a  and  a88740a );
 a88747a <=( A269  and  A267 );
 a88750a <=( A299  and  A298 );
 a88751a <=( a88750a  and  a88747a );
 a88752a <=( a88751a  and  a88744a );
 a88756a <=( (not A168)  and  (not A169) );
 a88757a <=( A170  and  a88756a );
 a88760a <=( A166  and  (not A167) );
 a88763a <=( (not A200)  and  A199 );
 a88764a <=( a88763a  and  a88760a );
 a88765a <=( a88764a  and  a88757a );
 a88768a <=( A202  and  A201 );
 a88771a <=( A266  and  (not A265) );
 a88772a <=( a88771a  and  a88768a );
 a88775a <=( A269  and  A267 );
 a88778a <=( (not A299)  and  (not A298) );
 a88779a <=( a88778a  and  a88775a );
 a88780a <=( a88779a  and  a88772a );
 a88784a <=( (not A168)  and  (not A169) );
 a88785a <=( A170  and  a88784a );
 a88788a <=( A166  and  (not A167) );
 a88791a <=( (not A200)  and  A199 );
 a88792a <=( a88791a  and  a88788a );
 a88793a <=( a88792a  and  a88785a );
 a88796a <=( A202  and  A201 );
 a88799a <=( (not A266)  and  A265 );
 a88800a <=( a88799a  and  a88796a );
 a88803a <=( A268  and  A267 );
 a88806a <=( A301  and  (not A300) );
 a88807a <=( a88806a  and  a88803a );
 a88808a <=( a88807a  and  a88800a );
 a88812a <=( (not A168)  and  (not A169) );
 a88813a <=( A170  and  a88812a );
 a88816a <=( A166  and  (not A167) );
 a88819a <=( (not A200)  and  A199 );
 a88820a <=( a88819a  and  a88816a );
 a88821a <=( a88820a  and  a88813a );
 a88824a <=( A202  and  A201 );
 a88827a <=( (not A266)  and  A265 );
 a88828a <=( a88827a  and  a88824a );
 a88831a <=( A268  and  A267 );
 a88834a <=( A302  and  (not A300) );
 a88835a <=( a88834a  and  a88831a );
 a88836a <=( a88835a  and  a88828a );
 a88840a <=( (not A168)  and  (not A169) );
 a88841a <=( A170  and  a88840a );
 a88844a <=( A166  and  (not A167) );
 a88847a <=( (not A200)  and  A199 );
 a88848a <=( a88847a  and  a88844a );
 a88849a <=( a88848a  and  a88841a );
 a88852a <=( A202  and  A201 );
 a88855a <=( (not A266)  and  A265 );
 a88856a <=( a88855a  and  a88852a );
 a88859a <=( A268  and  A267 );
 a88862a <=( A299  and  A298 );
 a88863a <=( a88862a  and  a88859a );
 a88864a <=( a88863a  and  a88856a );
 a88868a <=( (not A168)  and  (not A169) );
 a88869a <=( A170  and  a88868a );
 a88872a <=( A166  and  (not A167) );
 a88875a <=( (not A200)  and  A199 );
 a88876a <=( a88875a  and  a88872a );
 a88877a <=( a88876a  and  a88869a );
 a88880a <=( A202  and  A201 );
 a88883a <=( (not A266)  and  A265 );
 a88884a <=( a88883a  and  a88880a );
 a88887a <=( A268  and  A267 );
 a88890a <=( (not A299)  and  (not A298) );
 a88891a <=( a88890a  and  a88887a );
 a88892a <=( a88891a  and  a88884a );
 a88896a <=( (not A168)  and  (not A169) );
 a88897a <=( A170  and  a88896a );
 a88900a <=( A166  and  (not A167) );
 a88903a <=( (not A200)  and  A199 );
 a88904a <=( a88903a  and  a88900a );
 a88905a <=( a88904a  and  a88897a );
 a88908a <=( A202  and  A201 );
 a88911a <=( (not A266)  and  A265 );
 a88912a <=( a88911a  and  a88908a );
 a88915a <=( A269  and  A267 );
 a88918a <=( A301  and  (not A300) );
 a88919a <=( a88918a  and  a88915a );
 a88920a <=( a88919a  and  a88912a );
 a88924a <=( (not A168)  and  (not A169) );
 a88925a <=( A170  and  a88924a );
 a88928a <=( A166  and  (not A167) );
 a88931a <=( (not A200)  and  A199 );
 a88932a <=( a88931a  and  a88928a );
 a88933a <=( a88932a  and  a88925a );
 a88936a <=( A202  and  A201 );
 a88939a <=( (not A266)  and  A265 );
 a88940a <=( a88939a  and  a88936a );
 a88943a <=( A269  and  A267 );
 a88946a <=( A302  and  (not A300) );
 a88947a <=( a88946a  and  a88943a );
 a88948a <=( a88947a  and  a88940a );
 a88952a <=( (not A168)  and  (not A169) );
 a88953a <=( A170  and  a88952a );
 a88956a <=( A166  and  (not A167) );
 a88959a <=( (not A200)  and  A199 );
 a88960a <=( a88959a  and  a88956a );
 a88961a <=( a88960a  and  a88953a );
 a88964a <=( A202  and  A201 );
 a88967a <=( (not A266)  and  A265 );
 a88968a <=( a88967a  and  a88964a );
 a88971a <=( A269  and  A267 );
 a88974a <=( A299  and  A298 );
 a88975a <=( a88974a  and  a88971a );
 a88976a <=( a88975a  and  a88968a );
 a88980a <=( (not A168)  and  (not A169) );
 a88981a <=( A170  and  a88980a );
 a88984a <=( A166  and  (not A167) );
 a88987a <=( (not A200)  and  A199 );
 a88988a <=( a88987a  and  a88984a );
 a88989a <=( a88988a  and  a88981a );
 a88992a <=( A202  and  A201 );
 a88995a <=( (not A266)  and  A265 );
 a88996a <=( a88995a  and  a88992a );
 a88999a <=( A269  and  A267 );
 a89002a <=( (not A299)  and  (not A298) );
 a89003a <=( a89002a  and  a88999a );
 a89004a <=( a89003a  and  a88996a );
 a89008a <=( (not A168)  and  (not A169) );
 a89009a <=( A170  and  a89008a );
 a89012a <=( A166  and  (not A167) );
 a89015a <=( (not A200)  and  A199 );
 a89016a <=( a89015a  and  a89012a );
 a89017a <=( a89016a  and  a89009a );
 a89020a <=( A203  and  A201 );
 a89023a <=( A266  and  (not A265) );
 a89024a <=( a89023a  and  a89020a );
 a89027a <=( A268  and  A267 );
 a89030a <=( A301  and  (not A300) );
 a89031a <=( a89030a  and  a89027a );
 a89032a <=( a89031a  and  a89024a );
 a89036a <=( (not A168)  and  (not A169) );
 a89037a <=( A170  and  a89036a );
 a89040a <=( A166  and  (not A167) );
 a89043a <=( (not A200)  and  A199 );
 a89044a <=( a89043a  and  a89040a );
 a89045a <=( a89044a  and  a89037a );
 a89048a <=( A203  and  A201 );
 a89051a <=( A266  and  (not A265) );
 a89052a <=( a89051a  and  a89048a );
 a89055a <=( A268  and  A267 );
 a89058a <=( A302  and  (not A300) );
 a89059a <=( a89058a  and  a89055a );
 a89060a <=( a89059a  and  a89052a );
 a89064a <=( (not A168)  and  (not A169) );
 a89065a <=( A170  and  a89064a );
 a89068a <=( A166  and  (not A167) );
 a89071a <=( (not A200)  and  A199 );
 a89072a <=( a89071a  and  a89068a );
 a89073a <=( a89072a  and  a89065a );
 a89076a <=( A203  and  A201 );
 a89079a <=( A266  and  (not A265) );
 a89080a <=( a89079a  and  a89076a );
 a89083a <=( A268  and  A267 );
 a89086a <=( A299  and  A298 );
 a89087a <=( a89086a  and  a89083a );
 a89088a <=( a89087a  and  a89080a );
 a89092a <=( (not A168)  and  (not A169) );
 a89093a <=( A170  and  a89092a );
 a89096a <=( A166  and  (not A167) );
 a89099a <=( (not A200)  and  A199 );
 a89100a <=( a89099a  and  a89096a );
 a89101a <=( a89100a  and  a89093a );
 a89104a <=( A203  and  A201 );
 a89107a <=( A266  and  (not A265) );
 a89108a <=( a89107a  and  a89104a );
 a89111a <=( A268  and  A267 );
 a89114a <=( (not A299)  and  (not A298) );
 a89115a <=( a89114a  and  a89111a );
 a89116a <=( a89115a  and  a89108a );
 a89120a <=( (not A168)  and  (not A169) );
 a89121a <=( A170  and  a89120a );
 a89124a <=( A166  and  (not A167) );
 a89127a <=( (not A200)  and  A199 );
 a89128a <=( a89127a  and  a89124a );
 a89129a <=( a89128a  and  a89121a );
 a89132a <=( A203  and  A201 );
 a89135a <=( A266  and  (not A265) );
 a89136a <=( a89135a  and  a89132a );
 a89139a <=( A269  and  A267 );
 a89142a <=( A301  and  (not A300) );
 a89143a <=( a89142a  and  a89139a );
 a89144a <=( a89143a  and  a89136a );
 a89148a <=( (not A168)  and  (not A169) );
 a89149a <=( A170  and  a89148a );
 a89152a <=( A166  and  (not A167) );
 a89155a <=( (not A200)  and  A199 );
 a89156a <=( a89155a  and  a89152a );
 a89157a <=( a89156a  and  a89149a );
 a89160a <=( A203  and  A201 );
 a89163a <=( A266  and  (not A265) );
 a89164a <=( a89163a  and  a89160a );
 a89167a <=( A269  and  A267 );
 a89170a <=( A302  and  (not A300) );
 a89171a <=( a89170a  and  a89167a );
 a89172a <=( a89171a  and  a89164a );
 a89176a <=( (not A168)  and  (not A169) );
 a89177a <=( A170  and  a89176a );
 a89180a <=( A166  and  (not A167) );
 a89183a <=( (not A200)  and  A199 );
 a89184a <=( a89183a  and  a89180a );
 a89185a <=( a89184a  and  a89177a );
 a89188a <=( A203  and  A201 );
 a89191a <=( A266  and  (not A265) );
 a89192a <=( a89191a  and  a89188a );
 a89195a <=( A269  and  A267 );
 a89198a <=( A299  and  A298 );
 a89199a <=( a89198a  and  a89195a );
 a89200a <=( a89199a  and  a89192a );
 a89204a <=( (not A168)  and  (not A169) );
 a89205a <=( A170  and  a89204a );
 a89208a <=( A166  and  (not A167) );
 a89211a <=( (not A200)  and  A199 );
 a89212a <=( a89211a  and  a89208a );
 a89213a <=( a89212a  and  a89205a );
 a89216a <=( A203  and  A201 );
 a89219a <=( A266  and  (not A265) );
 a89220a <=( a89219a  and  a89216a );
 a89223a <=( A269  and  A267 );
 a89226a <=( (not A299)  and  (not A298) );
 a89227a <=( a89226a  and  a89223a );
 a89228a <=( a89227a  and  a89220a );
 a89232a <=( (not A168)  and  (not A169) );
 a89233a <=( A170  and  a89232a );
 a89236a <=( A166  and  (not A167) );
 a89239a <=( (not A200)  and  A199 );
 a89240a <=( a89239a  and  a89236a );
 a89241a <=( a89240a  and  a89233a );
 a89244a <=( A203  and  A201 );
 a89247a <=( (not A266)  and  A265 );
 a89248a <=( a89247a  and  a89244a );
 a89251a <=( A268  and  A267 );
 a89254a <=( A301  and  (not A300) );
 a89255a <=( a89254a  and  a89251a );
 a89256a <=( a89255a  and  a89248a );
 a89260a <=( (not A168)  and  (not A169) );
 a89261a <=( A170  and  a89260a );
 a89264a <=( A166  and  (not A167) );
 a89267a <=( (not A200)  and  A199 );
 a89268a <=( a89267a  and  a89264a );
 a89269a <=( a89268a  and  a89261a );
 a89272a <=( A203  and  A201 );
 a89275a <=( (not A266)  and  A265 );
 a89276a <=( a89275a  and  a89272a );
 a89279a <=( A268  and  A267 );
 a89282a <=( A302  and  (not A300) );
 a89283a <=( a89282a  and  a89279a );
 a89284a <=( a89283a  and  a89276a );
 a89288a <=( (not A168)  and  (not A169) );
 a89289a <=( A170  and  a89288a );
 a89292a <=( A166  and  (not A167) );
 a89295a <=( (not A200)  and  A199 );
 a89296a <=( a89295a  and  a89292a );
 a89297a <=( a89296a  and  a89289a );
 a89300a <=( A203  and  A201 );
 a89303a <=( (not A266)  and  A265 );
 a89304a <=( a89303a  and  a89300a );
 a89307a <=( A268  and  A267 );
 a89310a <=( A299  and  A298 );
 a89311a <=( a89310a  and  a89307a );
 a89312a <=( a89311a  and  a89304a );
 a89316a <=( (not A168)  and  (not A169) );
 a89317a <=( A170  and  a89316a );
 a89320a <=( A166  and  (not A167) );
 a89323a <=( (not A200)  and  A199 );
 a89324a <=( a89323a  and  a89320a );
 a89325a <=( a89324a  and  a89317a );
 a89328a <=( A203  and  A201 );
 a89331a <=( (not A266)  and  A265 );
 a89332a <=( a89331a  and  a89328a );
 a89335a <=( A268  and  A267 );
 a89338a <=( (not A299)  and  (not A298) );
 a89339a <=( a89338a  and  a89335a );
 a89340a <=( a89339a  and  a89332a );
 a89344a <=( (not A168)  and  (not A169) );
 a89345a <=( A170  and  a89344a );
 a89348a <=( A166  and  (not A167) );
 a89351a <=( (not A200)  and  A199 );
 a89352a <=( a89351a  and  a89348a );
 a89353a <=( a89352a  and  a89345a );
 a89356a <=( A203  and  A201 );
 a89359a <=( (not A266)  and  A265 );
 a89360a <=( a89359a  and  a89356a );
 a89363a <=( A269  and  A267 );
 a89366a <=( A301  and  (not A300) );
 a89367a <=( a89366a  and  a89363a );
 a89368a <=( a89367a  and  a89360a );
 a89372a <=( (not A168)  and  (not A169) );
 a89373a <=( A170  and  a89372a );
 a89376a <=( A166  and  (not A167) );
 a89379a <=( (not A200)  and  A199 );
 a89380a <=( a89379a  and  a89376a );
 a89381a <=( a89380a  and  a89373a );
 a89384a <=( A203  and  A201 );
 a89387a <=( (not A266)  and  A265 );
 a89388a <=( a89387a  and  a89384a );
 a89391a <=( A269  and  A267 );
 a89394a <=( A302  and  (not A300) );
 a89395a <=( a89394a  and  a89391a );
 a89396a <=( a89395a  and  a89388a );
 a89400a <=( (not A168)  and  (not A169) );
 a89401a <=( A170  and  a89400a );
 a89404a <=( A166  and  (not A167) );
 a89407a <=( (not A200)  and  A199 );
 a89408a <=( a89407a  and  a89404a );
 a89409a <=( a89408a  and  a89401a );
 a89412a <=( A203  and  A201 );
 a89415a <=( (not A266)  and  A265 );
 a89416a <=( a89415a  and  a89412a );
 a89419a <=( A269  and  A267 );
 a89422a <=( A299  and  A298 );
 a89423a <=( a89422a  and  a89419a );
 a89424a <=( a89423a  and  a89416a );
 a89428a <=( (not A168)  and  (not A169) );
 a89429a <=( A170  and  a89428a );
 a89432a <=( A166  and  (not A167) );
 a89435a <=( (not A200)  and  A199 );
 a89436a <=( a89435a  and  a89432a );
 a89437a <=( a89436a  and  a89429a );
 a89440a <=( A203  and  A201 );
 a89443a <=( (not A266)  and  A265 );
 a89444a <=( a89443a  and  a89440a );
 a89447a <=( A269  and  A267 );
 a89450a <=( (not A299)  and  (not A298) );
 a89451a <=( a89450a  and  a89447a );
 a89452a <=( a89451a  and  a89444a );
 a89456a <=( (not A168)  and  (not A169) );
 a89457a <=( A170  and  a89456a );
 a89460a <=( A166  and  (not A167) );
 a89463a <=( (not A200)  and  (not A199) );
 a89464a <=( a89463a  and  a89460a );
 a89465a <=( a89464a  and  a89457a );
 a89468a <=( (not A268)  and  A267 );
 a89471a <=( A298  and  (not A269) );
 a89472a <=( a89471a  and  a89468a );
 a89475a <=( (not A300)  and  (not A299) );
 a89478a <=( (not A302)  and  (not A301) );
 a89479a <=( a89478a  and  a89475a );
 a89480a <=( a89479a  and  a89472a );
 a89484a <=( (not A168)  and  (not A169) );
 a89485a <=( A170  and  a89484a );
 a89488a <=( A166  and  (not A167) );
 a89491a <=( (not A200)  and  (not A199) );
 a89492a <=( a89491a  and  a89488a );
 a89493a <=( a89492a  and  a89485a );
 a89496a <=( (not A268)  and  A267 );
 a89499a <=( (not A298)  and  (not A269) );
 a89500a <=( a89499a  and  a89496a );
 a89503a <=( (not A300)  and  A299 );
 a89506a <=( (not A302)  and  (not A301) );
 a89507a <=( a89506a  and  a89503a );
 a89508a <=( a89507a  and  a89500a );
 a89511a <=( A168  and  (not A170) );
 a89514a <=( (not A166)  and  A167 );
 a89515a <=( a89514a  and  a89511a );
 a89518a <=( A200  and  (not A199) );
 a89521a <=( A202  and  A201 );
 a89522a <=( a89521a  and  a89518a );
 a89523a <=( a89522a  and  a89515a );
 a89526a <=( A266  and  (not A265) );
 a89529a <=( (not A268)  and  (not A267) );
 a89530a <=( a89529a  and  a89526a );
 a89533a <=( A300  and  (not A269) );
 a89536a <=( (not A302)  and  (not A301) );
 a89537a <=( a89536a  and  a89533a );
 a89538a <=( a89537a  and  a89530a );
 a89541a <=( A168  and  (not A170) );
 a89544a <=( (not A166)  and  A167 );
 a89545a <=( a89544a  and  a89541a );
 a89548a <=( A200  and  (not A199) );
 a89551a <=( A202  and  A201 );
 a89552a <=( a89551a  and  a89548a );
 a89553a <=( a89552a  and  a89545a );
 a89556a <=( (not A266)  and  A265 );
 a89559a <=( (not A268)  and  (not A267) );
 a89560a <=( a89559a  and  a89556a );
 a89563a <=( A300  and  (not A269) );
 a89566a <=( (not A302)  and  (not A301) );
 a89567a <=( a89566a  and  a89563a );
 a89568a <=( a89567a  and  a89560a );
 a89571a <=( A168  and  (not A170) );
 a89574a <=( (not A166)  and  A167 );
 a89575a <=( a89574a  and  a89571a );
 a89578a <=( A200  and  (not A199) );
 a89581a <=( A203  and  A201 );
 a89582a <=( a89581a  and  a89578a );
 a89583a <=( a89582a  and  a89575a );
 a89586a <=( A266  and  (not A265) );
 a89589a <=( (not A268)  and  (not A267) );
 a89590a <=( a89589a  and  a89586a );
 a89593a <=( A300  and  (not A269) );
 a89596a <=( (not A302)  and  (not A301) );
 a89597a <=( a89596a  and  a89593a );
 a89598a <=( a89597a  and  a89590a );
 a89601a <=( A168  and  (not A170) );
 a89604a <=( (not A166)  and  A167 );
 a89605a <=( a89604a  and  a89601a );
 a89608a <=( A200  and  (not A199) );
 a89611a <=( A203  and  A201 );
 a89612a <=( a89611a  and  a89608a );
 a89613a <=( a89612a  and  a89605a );
 a89616a <=( (not A266)  and  A265 );
 a89619a <=( (not A268)  and  (not A267) );
 a89620a <=( a89619a  and  a89616a );
 a89623a <=( A300  and  (not A269) );
 a89626a <=( (not A302)  and  (not A301) );
 a89627a <=( a89626a  and  a89623a );
 a89628a <=( a89627a  and  a89620a );
 a89631a <=( A168  and  (not A170) );
 a89634a <=( (not A166)  and  A167 );
 a89635a <=( a89634a  and  a89631a );
 a89638a <=( A200  and  (not A199) );
 a89641a <=( (not A202)  and  (not A201) );
 a89642a <=( a89641a  and  a89638a );
 a89643a <=( a89642a  and  a89635a );
 a89646a <=( (not A265)  and  (not A203) );
 a89649a <=( A267  and  A266 );
 a89650a <=( a89649a  and  a89646a );
 a89653a <=( A300  and  A268 );
 a89656a <=( (not A302)  and  (not A301) );
 a89657a <=( a89656a  and  a89653a );
 a89658a <=( a89657a  and  a89650a );
 a89661a <=( A168  and  (not A170) );
 a89664a <=( (not A166)  and  A167 );
 a89665a <=( a89664a  and  a89661a );
 a89668a <=( A200  and  (not A199) );
 a89671a <=( (not A202)  and  (not A201) );
 a89672a <=( a89671a  and  a89668a );
 a89673a <=( a89672a  and  a89665a );
 a89676a <=( (not A265)  and  (not A203) );
 a89679a <=( A267  and  A266 );
 a89680a <=( a89679a  and  a89676a );
 a89683a <=( A300  and  A269 );
 a89686a <=( (not A302)  and  (not A301) );
 a89687a <=( a89686a  and  a89683a );
 a89688a <=( a89687a  and  a89680a );
 a89691a <=( A168  and  (not A170) );
 a89694a <=( (not A166)  and  A167 );
 a89695a <=( a89694a  and  a89691a );
 a89698a <=( A200  and  (not A199) );
 a89701a <=( (not A202)  and  (not A201) );
 a89702a <=( a89701a  and  a89698a );
 a89703a <=( a89702a  and  a89695a );
 a89706a <=( (not A265)  and  (not A203) );
 a89709a <=( (not A267)  and  A266 );
 a89710a <=( a89709a  and  a89706a );
 a89713a <=( (not A269)  and  (not A268) );
 a89716a <=( A301  and  (not A300) );
 a89717a <=( a89716a  and  a89713a );
 a89718a <=( a89717a  and  a89710a );
 a89721a <=( A168  and  (not A170) );
 a89724a <=( (not A166)  and  A167 );
 a89725a <=( a89724a  and  a89721a );
 a89728a <=( A200  and  (not A199) );
 a89731a <=( (not A202)  and  (not A201) );
 a89732a <=( a89731a  and  a89728a );
 a89733a <=( a89732a  and  a89725a );
 a89736a <=( (not A265)  and  (not A203) );
 a89739a <=( (not A267)  and  A266 );
 a89740a <=( a89739a  and  a89736a );
 a89743a <=( (not A269)  and  (not A268) );
 a89746a <=( A302  and  (not A300) );
 a89747a <=( a89746a  and  a89743a );
 a89748a <=( a89747a  and  a89740a );
 a89751a <=( A168  and  (not A170) );
 a89754a <=( (not A166)  and  A167 );
 a89755a <=( a89754a  and  a89751a );
 a89758a <=( A200  and  (not A199) );
 a89761a <=( (not A202)  and  (not A201) );
 a89762a <=( a89761a  and  a89758a );
 a89763a <=( a89762a  and  a89755a );
 a89766a <=( (not A265)  and  (not A203) );
 a89769a <=( (not A267)  and  A266 );
 a89770a <=( a89769a  and  a89766a );
 a89773a <=( (not A269)  and  (not A268) );
 a89776a <=( A299  and  A298 );
 a89777a <=( a89776a  and  a89773a );
 a89778a <=( a89777a  and  a89770a );
 a89781a <=( A168  and  (not A170) );
 a89784a <=( (not A166)  and  A167 );
 a89785a <=( a89784a  and  a89781a );
 a89788a <=( A200  and  (not A199) );
 a89791a <=( (not A202)  and  (not A201) );
 a89792a <=( a89791a  and  a89788a );
 a89793a <=( a89792a  and  a89785a );
 a89796a <=( (not A265)  and  (not A203) );
 a89799a <=( (not A267)  and  A266 );
 a89800a <=( a89799a  and  a89796a );
 a89803a <=( (not A269)  and  (not A268) );
 a89806a <=( (not A299)  and  (not A298) );
 a89807a <=( a89806a  and  a89803a );
 a89808a <=( a89807a  and  a89800a );
 a89811a <=( A168  and  (not A170) );
 a89814a <=( (not A166)  and  A167 );
 a89815a <=( a89814a  and  a89811a );
 a89818a <=( A200  and  (not A199) );
 a89821a <=( (not A202)  and  (not A201) );
 a89822a <=( a89821a  and  a89818a );
 a89823a <=( a89822a  and  a89815a );
 a89826a <=( A265  and  (not A203) );
 a89829a <=( A267  and  (not A266) );
 a89830a <=( a89829a  and  a89826a );
 a89833a <=( A300  and  A268 );
 a89836a <=( (not A302)  and  (not A301) );
 a89837a <=( a89836a  and  a89833a );
 a89838a <=( a89837a  and  a89830a );
 a89841a <=( A168  and  (not A170) );
 a89844a <=( (not A166)  and  A167 );
 a89845a <=( a89844a  and  a89841a );
 a89848a <=( A200  and  (not A199) );
 a89851a <=( (not A202)  and  (not A201) );
 a89852a <=( a89851a  and  a89848a );
 a89853a <=( a89852a  and  a89845a );
 a89856a <=( A265  and  (not A203) );
 a89859a <=( A267  and  (not A266) );
 a89860a <=( a89859a  and  a89856a );
 a89863a <=( A300  and  A269 );
 a89866a <=( (not A302)  and  (not A301) );
 a89867a <=( a89866a  and  a89863a );
 a89868a <=( a89867a  and  a89860a );
 a89871a <=( A168  and  (not A170) );
 a89874a <=( (not A166)  and  A167 );
 a89875a <=( a89874a  and  a89871a );
 a89878a <=( A200  and  (not A199) );
 a89881a <=( (not A202)  and  (not A201) );
 a89882a <=( a89881a  and  a89878a );
 a89883a <=( a89882a  and  a89875a );
 a89886a <=( A265  and  (not A203) );
 a89889a <=( (not A267)  and  (not A266) );
 a89890a <=( a89889a  and  a89886a );
 a89893a <=( (not A269)  and  (not A268) );
 a89896a <=( A301  and  (not A300) );
 a89897a <=( a89896a  and  a89893a );
 a89898a <=( a89897a  and  a89890a );
 a89901a <=( A168  and  (not A170) );
 a89904a <=( (not A166)  and  A167 );
 a89905a <=( a89904a  and  a89901a );
 a89908a <=( A200  and  (not A199) );
 a89911a <=( (not A202)  and  (not A201) );
 a89912a <=( a89911a  and  a89908a );
 a89913a <=( a89912a  and  a89905a );
 a89916a <=( A265  and  (not A203) );
 a89919a <=( (not A267)  and  (not A266) );
 a89920a <=( a89919a  and  a89916a );
 a89923a <=( (not A269)  and  (not A268) );
 a89926a <=( A302  and  (not A300) );
 a89927a <=( a89926a  and  a89923a );
 a89928a <=( a89927a  and  a89920a );
 a89931a <=( A168  and  (not A170) );
 a89934a <=( (not A166)  and  A167 );
 a89935a <=( a89934a  and  a89931a );
 a89938a <=( A200  and  (not A199) );
 a89941a <=( (not A202)  and  (not A201) );
 a89942a <=( a89941a  and  a89938a );
 a89943a <=( a89942a  and  a89935a );
 a89946a <=( A265  and  (not A203) );
 a89949a <=( (not A267)  and  (not A266) );
 a89950a <=( a89949a  and  a89946a );
 a89953a <=( (not A269)  and  (not A268) );
 a89956a <=( A299  and  A298 );
 a89957a <=( a89956a  and  a89953a );
 a89958a <=( a89957a  and  a89950a );
 a89961a <=( A168  and  (not A170) );
 a89964a <=( (not A166)  and  A167 );
 a89965a <=( a89964a  and  a89961a );
 a89968a <=( A200  and  (not A199) );
 a89971a <=( (not A202)  and  (not A201) );
 a89972a <=( a89971a  and  a89968a );
 a89973a <=( a89972a  and  a89965a );
 a89976a <=( A265  and  (not A203) );
 a89979a <=( (not A267)  and  (not A266) );
 a89980a <=( a89979a  and  a89976a );
 a89983a <=( (not A269)  and  (not A268) );
 a89986a <=( (not A299)  and  (not A298) );
 a89987a <=( a89986a  and  a89983a );
 a89988a <=( a89987a  and  a89980a );
 a89991a <=( A168  and  (not A170) );
 a89994a <=( (not A166)  and  A167 );
 a89995a <=( a89994a  and  a89991a );
 a89998a <=( (not A200)  and  A199 );
 a90001a <=( A202  and  A201 );
 a90002a <=( a90001a  and  a89998a );
 a90003a <=( a90002a  and  a89995a );
 a90006a <=( A266  and  (not A265) );
 a90009a <=( (not A268)  and  (not A267) );
 a90010a <=( a90009a  and  a90006a );
 a90013a <=( A300  and  (not A269) );
 a90016a <=( (not A302)  and  (not A301) );
 a90017a <=( a90016a  and  a90013a );
 a90018a <=( a90017a  and  a90010a );
 a90021a <=( A168  and  (not A170) );
 a90024a <=( (not A166)  and  A167 );
 a90025a <=( a90024a  and  a90021a );
 a90028a <=( (not A200)  and  A199 );
 a90031a <=( A202  and  A201 );
 a90032a <=( a90031a  and  a90028a );
 a90033a <=( a90032a  and  a90025a );
 a90036a <=( (not A266)  and  A265 );
 a90039a <=( (not A268)  and  (not A267) );
 a90040a <=( a90039a  and  a90036a );
 a90043a <=( A300  and  (not A269) );
 a90046a <=( (not A302)  and  (not A301) );
 a90047a <=( a90046a  and  a90043a );
 a90048a <=( a90047a  and  a90040a );
 a90051a <=( A168  and  (not A170) );
 a90054a <=( (not A166)  and  A167 );
 a90055a <=( a90054a  and  a90051a );
 a90058a <=( (not A200)  and  A199 );
 a90061a <=( A203  and  A201 );
 a90062a <=( a90061a  and  a90058a );
 a90063a <=( a90062a  and  a90055a );
 a90066a <=( A266  and  (not A265) );
 a90069a <=( (not A268)  and  (not A267) );
 a90070a <=( a90069a  and  a90066a );
 a90073a <=( A300  and  (not A269) );
 a90076a <=( (not A302)  and  (not A301) );
 a90077a <=( a90076a  and  a90073a );
 a90078a <=( a90077a  and  a90070a );
 a90081a <=( A168  and  (not A170) );
 a90084a <=( (not A166)  and  A167 );
 a90085a <=( a90084a  and  a90081a );
 a90088a <=( (not A200)  and  A199 );
 a90091a <=( A203  and  A201 );
 a90092a <=( a90091a  and  a90088a );
 a90093a <=( a90092a  and  a90085a );
 a90096a <=( (not A266)  and  A265 );
 a90099a <=( (not A268)  and  (not A267) );
 a90100a <=( a90099a  and  a90096a );
 a90103a <=( A300  and  (not A269) );
 a90106a <=( (not A302)  and  (not A301) );
 a90107a <=( a90106a  and  a90103a );
 a90108a <=( a90107a  and  a90100a );
 a90111a <=( A168  and  (not A170) );
 a90114a <=( (not A166)  and  A167 );
 a90115a <=( a90114a  and  a90111a );
 a90118a <=( (not A200)  and  A199 );
 a90121a <=( (not A202)  and  (not A201) );
 a90122a <=( a90121a  and  a90118a );
 a90123a <=( a90122a  and  a90115a );
 a90126a <=( (not A265)  and  (not A203) );
 a90129a <=( A267  and  A266 );
 a90130a <=( a90129a  and  a90126a );
 a90133a <=( A300  and  A268 );
 a90136a <=( (not A302)  and  (not A301) );
 a90137a <=( a90136a  and  a90133a );
 a90138a <=( a90137a  and  a90130a );
 a90141a <=( A168  and  (not A170) );
 a90144a <=( (not A166)  and  A167 );
 a90145a <=( a90144a  and  a90141a );
 a90148a <=( (not A200)  and  A199 );
 a90151a <=( (not A202)  and  (not A201) );
 a90152a <=( a90151a  and  a90148a );
 a90153a <=( a90152a  and  a90145a );
 a90156a <=( (not A265)  and  (not A203) );
 a90159a <=( A267  and  A266 );
 a90160a <=( a90159a  and  a90156a );
 a90163a <=( A300  and  A269 );
 a90166a <=( (not A302)  and  (not A301) );
 a90167a <=( a90166a  and  a90163a );
 a90168a <=( a90167a  and  a90160a );
 a90171a <=( A168  and  (not A170) );
 a90174a <=( (not A166)  and  A167 );
 a90175a <=( a90174a  and  a90171a );
 a90178a <=( (not A200)  and  A199 );
 a90181a <=( (not A202)  and  (not A201) );
 a90182a <=( a90181a  and  a90178a );
 a90183a <=( a90182a  and  a90175a );
 a90186a <=( (not A265)  and  (not A203) );
 a90189a <=( (not A267)  and  A266 );
 a90190a <=( a90189a  and  a90186a );
 a90193a <=( (not A269)  and  (not A268) );
 a90196a <=( A301  and  (not A300) );
 a90197a <=( a90196a  and  a90193a );
 a90198a <=( a90197a  and  a90190a );
 a90201a <=( A168  and  (not A170) );
 a90204a <=( (not A166)  and  A167 );
 a90205a <=( a90204a  and  a90201a );
 a90208a <=( (not A200)  and  A199 );
 a90211a <=( (not A202)  and  (not A201) );
 a90212a <=( a90211a  and  a90208a );
 a90213a <=( a90212a  and  a90205a );
 a90216a <=( (not A265)  and  (not A203) );
 a90219a <=( (not A267)  and  A266 );
 a90220a <=( a90219a  and  a90216a );
 a90223a <=( (not A269)  and  (not A268) );
 a90226a <=( A302  and  (not A300) );
 a90227a <=( a90226a  and  a90223a );
 a90228a <=( a90227a  and  a90220a );
 a90231a <=( A168  and  (not A170) );
 a90234a <=( (not A166)  and  A167 );
 a90235a <=( a90234a  and  a90231a );
 a90238a <=( (not A200)  and  A199 );
 a90241a <=( (not A202)  and  (not A201) );
 a90242a <=( a90241a  and  a90238a );
 a90243a <=( a90242a  and  a90235a );
 a90246a <=( (not A265)  and  (not A203) );
 a90249a <=( (not A267)  and  A266 );
 a90250a <=( a90249a  and  a90246a );
 a90253a <=( (not A269)  and  (not A268) );
 a90256a <=( A299  and  A298 );
 a90257a <=( a90256a  and  a90253a );
 a90258a <=( a90257a  and  a90250a );
 a90261a <=( A168  and  (not A170) );
 a90264a <=( (not A166)  and  A167 );
 a90265a <=( a90264a  and  a90261a );
 a90268a <=( (not A200)  and  A199 );
 a90271a <=( (not A202)  and  (not A201) );
 a90272a <=( a90271a  and  a90268a );
 a90273a <=( a90272a  and  a90265a );
 a90276a <=( (not A265)  and  (not A203) );
 a90279a <=( (not A267)  and  A266 );
 a90280a <=( a90279a  and  a90276a );
 a90283a <=( (not A269)  and  (not A268) );
 a90286a <=( (not A299)  and  (not A298) );
 a90287a <=( a90286a  and  a90283a );
 a90288a <=( a90287a  and  a90280a );
 a90291a <=( A168  and  (not A170) );
 a90294a <=( (not A166)  and  A167 );
 a90295a <=( a90294a  and  a90291a );
 a90298a <=( (not A200)  and  A199 );
 a90301a <=( (not A202)  and  (not A201) );
 a90302a <=( a90301a  and  a90298a );
 a90303a <=( a90302a  and  a90295a );
 a90306a <=( A265  and  (not A203) );
 a90309a <=( A267  and  (not A266) );
 a90310a <=( a90309a  and  a90306a );
 a90313a <=( A300  and  A268 );
 a90316a <=( (not A302)  and  (not A301) );
 a90317a <=( a90316a  and  a90313a );
 a90318a <=( a90317a  and  a90310a );
 a90321a <=( A168  and  (not A170) );
 a90324a <=( (not A166)  and  A167 );
 a90325a <=( a90324a  and  a90321a );
 a90328a <=( (not A200)  and  A199 );
 a90331a <=( (not A202)  and  (not A201) );
 a90332a <=( a90331a  and  a90328a );
 a90333a <=( a90332a  and  a90325a );
 a90336a <=( A265  and  (not A203) );
 a90339a <=( A267  and  (not A266) );
 a90340a <=( a90339a  and  a90336a );
 a90343a <=( A300  and  A269 );
 a90346a <=( (not A302)  and  (not A301) );
 a90347a <=( a90346a  and  a90343a );
 a90348a <=( a90347a  and  a90340a );
 a90351a <=( A168  and  (not A170) );
 a90354a <=( (not A166)  and  A167 );
 a90355a <=( a90354a  and  a90351a );
 a90358a <=( (not A200)  and  A199 );
 a90361a <=( (not A202)  and  (not A201) );
 a90362a <=( a90361a  and  a90358a );
 a90363a <=( a90362a  and  a90355a );
 a90366a <=( A265  and  (not A203) );
 a90369a <=( (not A267)  and  (not A266) );
 a90370a <=( a90369a  and  a90366a );
 a90373a <=( (not A269)  and  (not A268) );
 a90376a <=( A301  and  (not A300) );
 a90377a <=( a90376a  and  a90373a );
 a90378a <=( a90377a  and  a90370a );
 a90381a <=( A168  and  (not A170) );
 a90384a <=( (not A166)  and  A167 );
 a90385a <=( a90384a  and  a90381a );
 a90388a <=( (not A200)  and  A199 );
 a90391a <=( (not A202)  and  (not A201) );
 a90392a <=( a90391a  and  a90388a );
 a90393a <=( a90392a  and  a90385a );
 a90396a <=( A265  and  (not A203) );
 a90399a <=( (not A267)  and  (not A266) );
 a90400a <=( a90399a  and  a90396a );
 a90403a <=( (not A269)  and  (not A268) );
 a90406a <=( A302  and  (not A300) );
 a90407a <=( a90406a  and  a90403a );
 a90408a <=( a90407a  and  a90400a );
 a90411a <=( A168  and  (not A170) );
 a90414a <=( (not A166)  and  A167 );
 a90415a <=( a90414a  and  a90411a );
 a90418a <=( (not A200)  and  A199 );
 a90421a <=( (not A202)  and  (not A201) );
 a90422a <=( a90421a  and  a90418a );
 a90423a <=( a90422a  and  a90415a );
 a90426a <=( A265  and  (not A203) );
 a90429a <=( (not A267)  and  (not A266) );
 a90430a <=( a90429a  and  a90426a );
 a90433a <=( (not A269)  and  (not A268) );
 a90436a <=( A299  and  A298 );
 a90437a <=( a90436a  and  a90433a );
 a90438a <=( a90437a  and  a90430a );
 a90441a <=( A168  and  (not A170) );
 a90444a <=( (not A166)  and  A167 );
 a90445a <=( a90444a  and  a90441a );
 a90448a <=( (not A200)  and  A199 );
 a90451a <=( (not A202)  and  (not A201) );
 a90452a <=( a90451a  and  a90448a );
 a90453a <=( a90452a  and  a90445a );
 a90456a <=( A265  and  (not A203) );
 a90459a <=( (not A267)  and  (not A266) );
 a90460a <=( a90459a  and  a90456a );
 a90463a <=( (not A269)  and  (not A268) );
 a90466a <=( (not A299)  and  (not A298) );
 a90467a <=( a90466a  and  a90463a );
 a90468a <=( a90467a  and  a90460a );
 a90471a <=( A168  and  (not A170) );
 a90474a <=( A166  and  (not A167) );
 a90475a <=( a90474a  and  a90471a );
 a90478a <=( A200  and  (not A199) );
 a90481a <=( A202  and  A201 );
 a90482a <=( a90481a  and  a90478a );
 a90483a <=( a90482a  and  a90475a );
 a90486a <=( A266  and  (not A265) );
 a90489a <=( (not A268)  and  (not A267) );
 a90490a <=( a90489a  and  a90486a );
 a90493a <=( A300  and  (not A269) );
 a90496a <=( (not A302)  and  (not A301) );
 a90497a <=( a90496a  and  a90493a );
 a90498a <=( a90497a  and  a90490a );
 a90501a <=( A168  and  (not A170) );
 a90504a <=( A166  and  (not A167) );
 a90505a <=( a90504a  and  a90501a );
 a90508a <=( A200  and  (not A199) );
 a90511a <=( A202  and  A201 );
 a90512a <=( a90511a  and  a90508a );
 a90513a <=( a90512a  and  a90505a );
 a90516a <=( (not A266)  and  A265 );
 a90519a <=( (not A268)  and  (not A267) );
 a90520a <=( a90519a  and  a90516a );
 a90523a <=( A300  and  (not A269) );
 a90526a <=( (not A302)  and  (not A301) );
 a90527a <=( a90526a  and  a90523a );
 a90528a <=( a90527a  and  a90520a );
 a90531a <=( A168  and  (not A170) );
 a90534a <=( A166  and  (not A167) );
 a90535a <=( a90534a  and  a90531a );
 a90538a <=( A200  and  (not A199) );
 a90541a <=( A203  and  A201 );
 a90542a <=( a90541a  and  a90538a );
 a90543a <=( a90542a  and  a90535a );
 a90546a <=( A266  and  (not A265) );
 a90549a <=( (not A268)  and  (not A267) );
 a90550a <=( a90549a  and  a90546a );
 a90553a <=( A300  and  (not A269) );
 a90556a <=( (not A302)  and  (not A301) );
 a90557a <=( a90556a  and  a90553a );
 a90558a <=( a90557a  and  a90550a );
 a90561a <=( A168  and  (not A170) );
 a90564a <=( A166  and  (not A167) );
 a90565a <=( a90564a  and  a90561a );
 a90568a <=( A200  and  (not A199) );
 a90571a <=( A203  and  A201 );
 a90572a <=( a90571a  and  a90568a );
 a90573a <=( a90572a  and  a90565a );
 a90576a <=( (not A266)  and  A265 );
 a90579a <=( (not A268)  and  (not A267) );
 a90580a <=( a90579a  and  a90576a );
 a90583a <=( A300  and  (not A269) );
 a90586a <=( (not A302)  and  (not A301) );
 a90587a <=( a90586a  and  a90583a );
 a90588a <=( a90587a  and  a90580a );
 a90591a <=( A168  and  (not A170) );
 a90594a <=( A166  and  (not A167) );
 a90595a <=( a90594a  and  a90591a );
 a90598a <=( A200  and  (not A199) );
 a90601a <=( (not A202)  and  (not A201) );
 a90602a <=( a90601a  and  a90598a );
 a90603a <=( a90602a  and  a90595a );
 a90606a <=( (not A265)  and  (not A203) );
 a90609a <=( A267  and  A266 );
 a90610a <=( a90609a  and  a90606a );
 a90613a <=( A300  and  A268 );
 a90616a <=( (not A302)  and  (not A301) );
 a90617a <=( a90616a  and  a90613a );
 a90618a <=( a90617a  and  a90610a );
 a90621a <=( A168  and  (not A170) );
 a90624a <=( A166  and  (not A167) );
 a90625a <=( a90624a  and  a90621a );
 a90628a <=( A200  and  (not A199) );
 a90631a <=( (not A202)  and  (not A201) );
 a90632a <=( a90631a  and  a90628a );
 a90633a <=( a90632a  and  a90625a );
 a90636a <=( (not A265)  and  (not A203) );
 a90639a <=( A267  and  A266 );
 a90640a <=( a90639a  and  a90636a );
 a90643a <=( A300  and  A269 );
 a90646a <=( (not A302)  and  (not A301) );
 a90647a <=( a90646a  and  a90643a );
 a90648a <=( a90647a  and  a90640a );
 a90651a <=( A168  and  (not A170) );
 a90654a <=( A166  and  (not A167) );
 a90655a <=( a90654a  and  a90651a );
 a90658a <=( A200  and  (not A199) );
 a90661a <=( (not A202)  and  (not A201) );
 a90662a <=( a90661a  and  a90658a );
 a90663a <=( a90662a  and  a90655a );
 a90666a <=( (not A265)  and  (not A203) );
 a90669a <=( (not A267)  and  A266 );
 a90670a <=( a90669a  and  a90666a );
 a90673a <=( (not A269)  and  (not A268) );
 a90676a <=( A301  and  (not A300) );
 a90677a <=( a90676a  and  a90673a );
 a90678a <=( a90677a  and  a90670a );
 a90681a <=( A168  and  (not A170) );
 a90684a <=( A166  and  (not A167) );
 a90685a <=( a90684a  and  a90681a );
 a90688a <=( A200  and  (not A199) );
 a90691a <=( (not A202)  and  (not A201) );
 a90692a <=( a90691a  and  a90688a );
 a90693a <=( a90692a  and  a90685a );
 a90696a <=( (not A265)  and  (not A203) );
 a90699a <=( (not A267)  and  A266 );
 a90700a <=( a90699a  and  a90696a );
 a90703a <=( (not A269)  and  (not A268) );
 a90706a <=( A302  and  (not A300) );
 a90707a <=( a90706a  and  a90703a );
 a90708a <=( a90707a  and  a90700a );
 a90711a <=( A168  and  (not A170) );
 a90714a <=( A166  and  (not A167) );
 a90715a <=( a90714a  and  a90711a );
 a90718a <=( A200  and  (not A199) );
 a90721a <=( (not A202)  and  (not A201) );
 a90722a <=( a90721a  and  a90718a );
 a90723a <=( a90722a  and  a90715a );
 a90726a <=( (not A265)  and  (not A203) );
 a90729a <=( (not A267)  and  A266 );
 a90730a <=( a90729a  and  a90726a );
 a90733a <=( (not A269)  and  (not A268) );
 a90736a <=( A299  and  A298 );
 a90737a <=( a90736a  and  a90733a );
 a90738a <=( a90737a  and  a90730a );
 a90741a <=( A168  and  (not A170) );
 a90744a <=( A166  and  (not A167) );
 a90745a <=( a90744a  and  a90741a );
 a90748a <=( A200  and  (not A199) );
 a90751a <=( (not A202)  and  (not A201) );
 a90752a <=( a90751a  and  a90748a );
 a90753a <=( a90752a  and  a90745a );
 a90756a <=( (not A265)  and  (not A203) );
 a90759a <=( (not A267)  and  A266 );
 a90760a <=( a90759a  and  a90756a );
 a90763a <=( (not A269)  and  (not A268) );
 a90766a <=( (not A299)  and  (not A298) );
 a90767a <=( a90766a  and  a90763a );
 a90768a <=( a90767a  and  a90760a );
 a90771a <=( A168  and  (not A170) );
 a90774a <=( A166  and  (not A167) );
 a90775a <=( a90774a  and  a90771a );
 a90778a <=( A200  and  (not A199) );
 a90781a <=( (not A202)  and  (not A201) );
 a90782a <=( a90781a  and  a90778a );
 a90783a <=( a90782a  and  a90775a );
 a90786a <=( A265  and  (not A203) );
 a90789a <=( A267  and  (not A266) );
 a90790a <=( a90789a  and  a90786a );
 a90793a <=( A300  and  A268 );
 a90796a <=( (not A302)  and  (not A301) );
 a90797a <=( a90796a  and  a90793a );
 a90798a <=( a90797a  and  a90790a );
 a90801a <=( A168  and  (not A170) );
 a90804a <=( A166  and  (not A167) );
 a90805a <=( a90804a  and  a90801a );
 a90808a <=( A200  and  (not A199) );
 a90811a <=( (not A202)  and  (not A201) );
 a90812a <=( a90811a  and  a90808a );
 a90813a <=( a90812a  and  a90805a );
 a90816a <=( A265  and  (not A203) );
 a90819a <=( A267  and  (not A266) );
 a90820a <=( a90819a  and  a90816a );
 a90823a <=( A300  and  A269 );
 a90826a <=( (not A302)  and  (not A301) );
 a90827a <=( a90826a  and  a90823a );
 a90828a <=( a90827a  and  a90820a );
 a90831a <=( A168  and  (not A170) );
 a90834a <=( A166  and  (not A167) );
 a90835a <=( a90834a  and  a90831a );
 a90838a <=( A200  and  (not A199) );
 a90841a <=( (not A202)  and  (not A201) );
 a90842a <=( a90841a  and  a90838a );
 a90843a <=( a90842a  and  a90835a );
 a90846a <=( A265  and  (not A203) );
 a90849a <=( (not A267)  and  (not A266) );
 a90850a <=( a90849a  and  a90846a );
 a90853a <=( (not A269)  and  (not A268) );
 a90856a <=( A301  and  (not A300) );
 a90857a <=( a90856a  and  a90853a );
 a90858a <=( a90857a  and  a90850a );
 a90861a <=( A168  and  (not A170) );
 a90864a <=( A166  and  (not A167) );
 a90865a <=( a90864a  and  a90861a );
 a90868a <=( A200  and  (not A199) );
 a90871a <=( (not A202)  and  (not A201) );
 a90872a <=( a90871a  and  a90868a );
 a90873a <=( a90872a  and  a90865a );
 a90876a <=( A265  and  (not A203) );
 a90879a <=( (not A267)  and  (not A266) );
 a90880a <=( a90879a  and  a90876a );
 a90883a <=( (not A269)  and  (not A268) );
 a90886a <=( A302  and  (not A300) );
 a90887a <=( a90886a  and  a90883a );
 a90888a <=( a90887a  and  a90880a );
 a90891a <=( A168  and  (not A170) );
 a90894a <=( A166  and  (not A167) );
 a90895a <=( a90894a  and  a90891a );
 a90898a <=( A200  and  (not A199) );
 a90901a <=( (not A202)  and  (not A201) );
 a90902a <=( a90901a  and  a90898a );
 a90903a <=( a90902a  and  a90895a );
 a90906a <=( A265  and  (not A203) );
 a90909a <=( (not A267)  and  (not A266) );
 a90910a <=( a90909a  and  a90906a );
 a90913a <=( (not A269)  and  (not A268) );
 a90916a <=( A299  and  A298 );
 a90917a <=( a90916a  and  a90913a );
 a90918a <=( a90917a  and  a90910a );
 a90921a <=( A168  and  (not A170) );
 a90924a <=( A166  and  (not A167) );
 a90925a <=( a90924a  and  a90921a );
 a90928a <=( A200  and  (not A199) );
 a90931a <=( (not A202)  and  (not A201) );
 a90932a <=( a90931a  and  a90928a );
 a90933a <=( a90932a  and  a90925a );
 a90936a <=( A265  and  (not A203) );
 a90939a <=( (not A267)  and  (not A266) );
 a90940a <=( a90939a  and  a90936a );
 a90943a <=( (not A269)  and  (not A268) );
 a90946a <=( (not A299)  and  (not A298) );
 a90947a <=( a90946a  and  a90943a );
 a90948a <=( a90947a  and  a90940a );
 a90951a <=( A168  and  (not A170) );
 a90954a <=( A166  and  (not A167) );
 a90955a <=( a90954a  and  a90951a );
 a90958a <=( (not A200)  and  A199 );
 a90961a <=( A202  and  A201 );
 a90962a <=( a90961a  and  a90958a );
 a90963a <=( a90962a  and  a90955a );
 a90966a <=( A266  and  (not A265) );
 a90969a <=( (not A268)  and  (not A267) );
 a90970a <=( a90969a  and  a90966a );
 a90973a <=( A300  and  (not A269) );
 a90976a <=( (not A302)  and  (not A301) );
 a90977a <=( a90976a  and  a90973a );
 a90978a <=( a90977a  and  a90970a );
 a90981a <=( A168  and  (not A170) );
 a90984a <=( A166  and  (not A167) );
 a90985a <=( a90984a  and  a90981a );
 a90988a <=( (not A200)  and  A199 );
 a90991a <=( A202  and  A201 );
 a90992a <=( a90991a  and  a90988a );
 a90993a <=( a90992a  and  a90985a );
 a90996a <=( (not A266)  and  A265 );
 a90999a <=( (not A268)  and  (not A267) );
 a91000a <=( a90999a  and  a90996a );
 a91003a <=( A300  and  (not A269) );
 a91006a <=( (not A302)  and  (not A301) );
 a91007a <=( a91006a  and  a91003a );
 a91008a <=( a91007a  and  a91000a );
 a91011a <=( A168  and  (not A170) );
 a91014a <=( A166  and  (not A167) );
 a91015a <=( a91014a  and  a91011a );
 a91018a <=( (not A200)  and  A199 );
 a91021a <=( A203  and  A201 );
 a91022a <=( a91021a  and  a91018a );
 a91023a <=( a91022a  and  a91015a );
 a91026a <=( A266  and  (not A265) );
 a91029a <=( (not A268)  and  (not A267) );
 a91030a <=( a91029a  and  a91026a );
 a91033a <=( A300  and  (not A269) );
 a91036a <=( (not A302)  and  (not A301) );
 a91037a <=( a91036a  and  a91033a );
 a91038a <=( a91037a  and  a91030a );
 a91041a <=( A168  and  (not A170) );
 a91044a <=( A166  and  (not A167) );
 a91045a <=( a91044a  and  a91041a );
 a91048a <=( (not A200)  and  A199 );
 a91051a <=( A203  and  A201 );
 a91052a <=( a91051a  and  a91048a );
 a91053a <=( a91052a  and  a91045a );
 a91056a <=( (not A266)  and  A265 );
 a91059a <=( (not A268)  and  (not A267) );
 a91060a <=( a91059a  and  a91056a );
 a91063a <=( A300  and  (not A269) );
 a91066a <=( (not A302)  and  (not A301) );
 a91067a <=( a91066a  and  a91063a );
 a91068a <=( a91067a  and  a91060a );
 a91071a <=( A168  and  (not A170) );
 a91074a <=( A166  and  (not A167) );
 a91075a <=( a91074a  and  a91071a );
 a91078a <=( (not A200)  and  A199 );
 a91081a <=( (not A202)  and  (not A201) );
 a91082a <=( a91081a  and  a91078a );
 a91083a <=( a91082a  and  a91075a );
 a91086a <=( (not A265)  and  (not A203) );
 a91089a <=( A267  and  A266 );
 a91090a <=( a91089a  and  a91086a );
 a91093a <=( A300  and  A268 );
 a91096a <=( (not A302)  and  (not A301) );
 a91097a <=( a91096a  and  a91093a );
 a91098a <=( a91097a  and  a91090a );
 a91101a <=( A168  and  (not A170) );
 a91104a <=( A166  and  (not A167) );
 a91105a <=( a91104a  and  a91101a );
 a91108a <=( (not A200)  and  A199 );
 a91111a <=( (not A202)  and  (not A201) );
 a91112a <=( a91111a  and  a91108a );
 a91113a <=( a91112a  and  a91105a );
 a91116a <=( (not A265)  and  (not A203) );
 a91119a <=( A267  and  A266 );
 a91120a <=( a91119a  and  a91116a );
 a91123a <=( A300  and  A269 );
 a91126a <=( (not A302)  and  (not A301) );
 a91127a <=( a91126a  and  a91123a );
 a91128a <=( a91127a  and  a91120a );
 a91131a <=( A168  and  (not A170) );
 a91134a <=( A166  and  (not A167) );
 a91135a <=( a91134a  and  a91131a );
 a91138a <=( (not A200)  and  A199 );
 a91141a <=( (not A202)  and  (not A201) );
 a91142a <=( a91141a  and  a91138a );
 a91143a <=( a91142a  and  a91135a );
 a91146a <=( (not A265)  and  (not A203) );
 a91149a <=( (not A267)  and  A266 );
 a91150a <=( a91149a  and  a91146a );
 a91153a <=( (not A269)  and  (not A268) );
 a91156a <=( A301  and  (not A300) );
 a91157a <=( a91156a  and  a91153a );
 a91158a <=( a91157a  and  a91150a );
 a91161a <=( A168  and  (not A170) );
 a91164a <=( A166  and  (not A167) );
 a91165a <=( a91164a  and  a91161a );
 a91168a <=( (not A200)  and  A199 );
 a91171a <=( (not A202)  and  (not A201) );
 a91172a <=( a91171a  and  a91168a );
 a91173a <=( a91172a  and  a91165a );
 a91176a <=( (not A265)  and  (not A203) );
 a91179a <=( (not A267)  and  A266 );
 a91180a <=( a91179a  and  a91176a );
 a91183a <=( (not A269)  and  (not A268) );
 a91186a <=( A302  and  (not A300) );
 a91187a <=( a91186a  and  a91183a );
 a91188a <=( a91187a  and  a91180a );
 a91191a <=( A168  and  (not A170) );
 a91194a <=( A166  and  (not A167) );
 a91195a <=( a91194a  and  a91191a );
 a91198a <=( (not A200)  and  A199 );
 a91201a <=( (not A202)  and  (not A201) );
 a91202a <=( a91201a  and  a91198a );
 a91203a <=( a91202a  and  a91195a );
 a91206a <=( (not A265)  and  (not A203) );
 a91209a <=( (not A267)  and  A266 );
 a91210a <=( a91209a  and  a91206a );
 a91213a <=( (not A269)  and  (not A268) );
 a91216a <=( A299  and  A298 );
 a91217a <=( a91216a  and  a91213a );
 a91218a <=( a91217a  and  a91210a );
 a91221a <=( A168  and  (not A170) );
 a91224a <=( A166  and  (not A167) );
 a91225a <=( a91224a  and  a91221a );
 a91228a <=( (not A200)  and  A199 );
 a91231a <=( (not A202)  and  (not A201) );
 a91232a <=( a91231a  and  a91228a );
 a91233a <=( a91232a  and  a91225a );
 a91236a <=( (not A265)  and  (not A203) );
 a91239a <=( (not A267)  and  A266 );
 a91240a <=( a91239a  and  a91236a );
 a91243a <=( (not A269)  and  (not A268) );
 a91246a <=( (not A299)  and  (not A298) );
 a91247a <=( a91246a  and  a91243a );
 a91248a <=( a91247a  and  a91240a );
 a91251a <=( A168  and  (not A170) );
 a91254a <=( A166  and  (not A167) );
 a91255a <=( a91254a  and  a91251a );
 a91258a <=( (not A200)  and  A199 );
 a91261a <=( (not A202)  and  (not A201) );
 a91262a <=( a91261a  and  a91258a );
 a91263a <=( a91262a  and  a91255a );
 a91266a <=( A265  and  (not A203) );
 a91269a <=( A267  and  (not A266) );
 a91270a <=( a91269a  and  a91266a );
 a91273a <=( A300  and  A268 );
 a91276a <=( (not A302)  and  (not A301) );
 a91277a <=( a91276a  and  a91273a );
 a91278a <=( a91277a  and  a91270a );
 a91281a <=( A168  and  (not A170) );
 a91284a <=( A166  and  (not A167) );
 a91285a <=( a91284a  and  a91281a );
 a91288a <=( (not A200)  and  A199 );
 a91291a <=( (not A202)  and  (not A201) );
 a91292a <=( a91291a  and  a91288a );
 a91293a <=( a91292a  and  a91285a );
 a91296a <=( A265  and  (not A203) );
 a91299a <=( A267  and  (not A266) );
 a91300a <=( a91299a  and  a91296a );
 a91303a <=( A300  and  A269 );
 a91306a <=( (not A302)  and  (not A301) );
 a91307a <=( a91306a  and  a91303a );
 a91308a <=( a91307a  and  a91300a );
 a91311a <=( A168  and  (not A170) );
 a91314a <=( A166  and  (not A167) );
 a91315a <=( a91314a  and  a91311a );
 a91318a <=( (not A200)  and  A199 );
 a91321a <=( (not A202)  and  (not A201) );
 a91322a <=( a91321a  and  a91318a );
 a91323a <=( a91322a  and  a91315a );
 a91326a <=( A265  and  (not A203) );
 a91329a <=( (not A267)  and  (not A266) );
 a91330a <=( a91329a  and  a91326a );
 a91333a <=( (not A269)  and  (not A268) );
 a91336a <=( A301  and  (not A300) );
 a91337a <=( a91336a  and  a91333a );
 a91338a <=( a91337a  and  a91330a );
 a91341a <=( A168  and  (not A170) );
 a91344a <=( A166  and  (not A167) );
 a91345a <=( a91344a  and  a91341a );
 a91348a <=( (not A200)  and  A199 );
 a91351a <=( (not A202)  and  (not A201) );
 a91352a <=( a91351a  and  a91348a );
 a91353a <=( a91352a  and  a91345a );
 a91356a <=( A265  and  (not A203) );
 a91359a <=( (not A267)  and  (not A266) );
 a91360a <=( a91359a  and  a91356a );
 a91363a <=( (not A269)  and  (not A268) );
 a91366a <=( A302  and  (not A300) );
 a91367a <=( a91366a  and  a91363a );
 a91368a <=( a91367a  and  a91360a );
 a91371a <=( A168  and  (not A170) );
 a91374a <=( A166  and  (not A167) );
 a91375a <=( a91374a  and  a91371a );
 a91378a <=( (not A200)  and  A199 );
 a91381a <=( (not A202)  and  (not A201) );
 a91382a <=( a91381a  and  a91378a );
 a91383a <=( a91382a  and  a91375a );
 a91386a <=( A265  and  (not A203) );
 a91389a <=( (not A267)  and  (not A266) );
 a91390a <=( a91389a  and  a91386a );
 a91393a <=( (not A269)  and  (not A268) );
 a91396a <=( A299  and  A298 );
 a91397a <=( a91396a  and  a91393a );
 a91398a <=( a91397a  and  a91390a );
 a91401a <=( A168  and  (not A170) );
 a91404a <=( A166  and  (not A167) );
 a91405a <=( a91404a  and  a91401a );
 a91408a <=( (not A200)  and  A199 );
 a91411a <=( (not A202)  and  (not A201) );
 a91412a <=( a91411a  and  a91408a );
 a91413a <=( a91412a  and  a91405a );
 a91416a <=( A265  and  (not A203) );
 a91419a <=( (not A267)  and  (not A266) );
 a91420a <=( a91419a  and  a91416a );
 a91423a <=( (not A269)  and  (not A268) );
 a91426a <=( (not A299)  and  (not A298) );
 a91427a <=( a91426a  and  a91423a );
 a91428a <=( a91427a  and  a91420a );
 a91431a <=( A168  and  A169 );
 a91434a <=( (not A166)  and  A167 );
 a91435a <=( a91434a  and  a91431a );
 a91438a <=( A200  and  (not A199) );
 a91441a <=( A202  and  A201 );
 a91442a <=( a91441a  and  a91438a );
 a91443a <=( a91442a  and  a91435a );
 a91446a <=( A266  and  (not A265) );
 a91449a <=( (not A268)  and  (not A267) );
 a91450a <=( a91449a  and  a91446a );
 a91453a <=( A300  and  (not A269) );
 a91456a <=( (not A302)  and  (not A301) );
 a91457a <=( a91456a  and  a91453a );
 a91458a <=( a91457a  and  a91450a );
 a91461a <=( A168  and  A169 );
 a91464a <=( (not A166)  and  A167 );
 a91465a <=( a91464a  and  a91461a );
 a91468a <=( A200  and  (not A199) );
 a91471a <=( A202  and  A201 );
 a91472a <=( a91471a  and  a91468a );
 a91473a <=( a91472a  and  a91465a );
 a91476a <=( (not A266)  and  A265 );
 a91479a <=( (not A268)  and  (not A267) );
 a91480a <=( a91479a  and  a91476a );
 a91483a <=( A300  and  (not A269) );
 a91486a <=( (not A302)  and  (not A301) );
 a91487a <=( a91486a  and  a91483a );
 a91488a <=( a91487a  and  a91480a );
 a91491a <=( A168  and  A169 );
 a91494a <=( (not A166)  and  A167 );
 a91495a <=( a91494a  and  a91491a );
 a91498a <=( A200  and  (not A199) );
 a91501a <=( A203  and  A201 );
 a91502a <=( a91501a  and  a91498a );
 a91503a <=( a91502a  and  a91495a );
 a91506a <=( A266  and  (not A265) );
 a91509a <=( (not A268)  and  (not A267) );
 a91510a <=( a91509a  and  a91506a );
 a91513a <=( A300  and  (not A269) );
 a91516a <=( (not A302)  and  (not A301) );
 a91517a <=( a91516a  and  a91513a );
 a91518a <=( a91517a  and  a91510a );
 a91521a <=( A168  and  A169 );
 a91524a <=( (not A166)  and  A167 );
 a91525a <=( a91524a  and  a91521a );
 a91528a <=( A200  and  (not A199) );
 a91531a <=( A203  and  A201 );
 a91532a <=( a91531a  and  a91528a );
 a91533a <=( a91532a  and  a91525a );
 a91536a <=( (not A266)  and  A265 );
 a91539a <=( (not A268)  and  (not A267) );
 a91540a <=( a91539a  and  a91536a );
 a91543a <=( A300  and  (not A269) );
 a91546a <=( (not A302)  and  (not A301) );
 a91547a <=( a91546a  and  a91543a );
 a91548a <=( a91547a  and  a91540a );
 a91551a <=( A168  and  A169 );
 a91554a <=( (not A166)  and  A167 );
 a91555a <=( a91554a  and  a91551a );
 a91558a <=( A200  and  (not A199) );
 a91561a <=( (not A202)  and  (not A201) );
 a91562a <=( a91561a  and  a91558a );
 a91563a <=( a91562a  and  a91555a );
 a91566a <=( (not A265)  and  (not A203) );
 a91569a <=( A267  and  A266 );
 a91570a <=( a91569a  and  a91566a );
 a91573a <=( A300  and  A268 );
 a91576a <=( (not A302)  and  (not A301) );
 a91577a <=( a91576a  and  a91573a );
 a91578a <=( a91577a  and  a91570a );
 a91581a <=( A168  and  A169 );
 a91584a <=( (not A166)  and  A167 );
 a91585a <=( a91584a  and  a91581a );
 a91588a <=( A200  and  (not A199) );
 a91591a <=( (not A202)  and  (not A201) );
 a91592a <=( a91591a  and  a91588a );
 a91593a <=( a91592a  and  a91585a );
 a91596a <=( (not A265)  and  (not A203) );
 a91599a <=( A267  and  A266 );
 a91600a <=( a91599a  and  a91596a );
 a91603a <=( A300  and  A269 );
 a91606a <=( (not A302)  and  (not A301) );
 a91607a <=( a91606a  and  a91603a );
 a91608a <=( a91607a  and  a91600a );
 a91611a <=( A168  and  A169 );
 a91614a <=( (not A166)  and  A167 );
 a91615a <=( a91614a  and  a91611a );
 a91618a <=( A200  and  (not A199) );
 a91621a <=( (not A202)  and  (not A201) );
 a91622a <=( a91621a  and  a91618a );
 a91623a <=( a91622a  and  a91615a );
 a91626a <=( (not A265)  and  (not A203) );
 a91629a <=( (not A267)  and  A266 );
 a91630a <=( a91629a  and  a91626a );
 a91633a <=( (not A269)  and  (not A268) );
 a91636a <=( A301  and  (not A300) );
 a91637a <=( a91636a  and  a91633a );
 a91638a <=( a91637a  and  a91630a );
 a91641a <=( A168  and  A169 );
 a91644a <=( (not A166)  and  A167 );
 a91645a <=( a91644a  and  a91641a );
 a91648a <=( A200  and  (not A199) );
 a91651a <=( (not A202)  and  (not A201) );
 a91652a <=( a91651a  and  a91648a );
 a91653a <=( a91652a  and  a91645a );
 a91656a <=( (not A265)  and  (not A203) );
 a91659a <=( (not A267)  and  A266 );
 a91660a <=( a91659a  and  a91656a );
 a91663a <=( (not A269)  and  (not A268) );
 a91666a <=( A302  and  (not A300) );
 a91667a <=( a91666a  and  a91663a );
 a91668a <=( a91667a  and  a91660a );
 a91671a <=( A168  and  A169 );
 a91674a <=( (not A166)  and  A167 );
 a91675a <=( a91674a  and  a91671a );
 a91678a <=( A200  and  (not A199) );
 a91681a <=( (not A202)  and  (not A201) );
 a91682a <=( a91681a  and  a91678a );
 a91683a <=( a91682a  and  a91675a );
 a91686a <=( (not A265)  and  (not A203) );
 a91689a <=( (not A267)  and  A266 );
 a91690a <=( a91689a  and  a91686a );
 a91693a <=( (not A269)  and  (not A268) );
 a91696a <=( A299  and  A298 );
 a91697a <=( a91696a  and  a91693a );
 a91698a <=( a91697a  and  a91690a );
 a91701a <=( A168  and  A169 );
 a91704a <=( (not A166)  and  A167 );
 a91705a <=( a91704a  and  a91701a );
 a91708a <=( A200  and  (not A199) );
 a91711a <=( (not A202)  and  (not A201) );
 a91712a <=( a91711a  and  a91708a );
 a91713a <=( a91712a  and  a91705a );
 a91716a <=( (not A265)  and  (not A203) );
 a91719a <=( (not A267)  and  A266 );
 a91720a <=( a91719a  and  a91716a );
 a91723a <=( (not A269)  and  (not A268) );
 a91726a <=( (not A299)  and  (not A298) );
 a91727a <=( a91726a  and  a91723a );
 a91728a <=( a91727a  and  a91720a );
 a91731a <=( A168  and  A169 );
 a91734a <=( (not A166)  and  A167 );
 a91735a <=( a91734a  and  a91731a );
 a91738a <=( A200  and  (not A199) );
 a91741a <=( (not A202)  and  (not A201) );
 a91742a <=( a91741a  and  a91738a );
 a91743a <=( a91742a  and  a91735a );
 a91746a <=( A265  and  (not A203) );
 a91749a <=( A267  and  (not A266) );
 a91750a <=( a91749a  and  a91746a );
 a91753a <=( A300  and  A268 );
 a91756a <=( (not A302)  and  (not A301) );
 a91757a <=( a91756a  and  a91753a );
 a91758a <=( a91757a  and  a91750a );
 a91761a <=( A168  and  A169 );
 a91764a <=( (not A166)  and  A167 );
 a91765a <=( a91764a  and  a91761a );
 a91768a <=( A200  and  (not A199) );
 a91771a <=( (not A202)  and  (not A201) );
 a91772a <=( a91771a  and  a91768a );
 a91773a <=( a91772a  and  a91765a );
 a91776a <=( A265  and  (not A203) );
 a91779a <=( A267  and  (not A266) );
 a91780a <=( a91779a  and  a91776a );
 a91783a <=( A300  and  A269 );
 a91786a <=( (not A302)  and  (not A301) );
 a91787a <=( a91786a  and  a91783a );
 a91788a <=( a91787a  and  a91780a );
 a91791a <=( A168  and  A169 );
 a91794a <=( (not A166)  and  A167 );
 a91795a <=( a91794a  and  a91791a );
 a91798a <=( A200  and  (not A199) );
 a91801a <=( (not A202)  and  (not A201) );
 a91802a <=( a91801a  and  a91798a );
 a91803a <=( a91802a  and  a91795a );
 a91806a <=( A265  and  (not A203) );
 a91809a <=( (not A267)  and  (not A266) );
 a91810a <=( a91809a  and  a91806a );
 a91813a <=( (not A269)  and  (not A268) );
 a91816a <=( A301  and  (not A300) );
 a91817a <=( a91816a  and  a91813a );
 a91818a <=( a91817a  and  a91810a );
 a91821a <=( A168  and  A169 );
 a91824a <=( (not A166)  and  A167 );
 a91825a <=( a91824a  and  a91821a );
 a91828a <=( A200  and  (not A199) );
 a91831a <=( (not A202)  and  (not A201) );
 a91832a <=( a91831a  and  a91828a );
 a91833a <=( a91832a  and  a91825a );
 a91836a <=( A265  and  (not A203) );
 a91839a <=( (not A267)  and  (not A266) );
 a91840a <=( a91839a  and  a91836a );
 a91843a <=( (not A269)  and  (not A268) );
 a91846a <=( A302  and  (not A300) );
 a91847a <=( a91846a  and  a91843a );
 a91848a <=( a91847a  and  a91840a );
 a91851a <=( A168  and  A169 );
 a91854a <=( (not A166)  and  A167 );
 a91855a <=( a91854a  and  a91851a );
 a91858a <=( A200  and  (not A199) );
 a91861a <=( (not A202)  and  (not A201) );
 a91862a <=( a91861a  and  a91858a );
 a91863a <=( a91862a  and  a91855a );
 a91866a <=( A265  and  (not A203) );
 a91869a <=( (not A267)  and  (not A266) );
 a91870a <=( a91869a  and  a91866a );
 a91873a <=( (not A269)  and  (not A268) );
 a91876a <=( A299  and  A298 );
 a91877a <=( a91876a  and  a91873a );
 a91878a <=( a91877a  and  a91870a );
 a91881a <=( A168  and  A169 );
 a91884a <=( (not A166)  and  A167 );
 a91885a <=( a91884a  and  a91881a );
 a91888a <=( A200  and  (not A199) );
 a91891a <=( (not A202)  and  (not A201) );
 a91892a <=( a91891a  and  a91888a );
 a91893a <=( a91892a  and  a91885a );
 a91896a <=( A265  and  (not A203) );
 a91899a <=( (not A267)  and  (not A266) );
 a91900a <=( a91899a  and  a91896a );
 a91903a <=( (not A269)  and  (not A268) );
 a91906a <=( (not A299)  and  (not A298) );
 a91907a <=( a91906a  and  a91903a );
 a91908a <=( a91907a  and  a91900a );
 a91911a <=( A168  and  A169 );
 a91914a <=( (not A166)  and  A167 );
 a91915a <=( a91914a  and  a91911a );
 a91918a <=( (not A200)  and  A199 );
 a91921a <=( A202  and  A201 );
 a91922a <=( a91921a  and  a91918a );
 a91923a <=( a91922a  and  a91915a );
 a91926a <=( A266  and  (not A265) );
 a91929a <=( (not A268)  and  (not A267) );
 a91930a <=( a91929a  and  a91926a );
 a91933a <=( A300  and  (not A269) );
 a91936a <=( (not A302)  and  (not A301) );
 a91937a <=( a91936a  and  a91933a );
 a91938a <=( a91937a  and  a91930a );
 a91941a <=( A168  and  A169 );
 a91944a <=( (not A166)  and  A167 );
 a91945a <=( a91944a  and  a91941a );
 a91948a <=( (not A200)  and  A199 );
 a91951a <=( A202  and  A201 );
 a91952a <=( a91951a  and  a91948a );
 a91953a <=( a91952a  and  a91945a );
 a91956a <=( (not A266)  and  A265 );
 a91959a <=( (not A268)  and  (not A267) );
 a91960a <=( a91959a  and  a91956a );
 a91963a <=( A300  and  (not A269) );
 a91966a <=( (not A302)  and  (not A301) );
 a91967a <=( a91966a  and  a91963a );
 a91968a <=( a91967a  and  a91960a );
 a91971a <=( A168  and  A169 );
 a91974a <=( (not A166)  and  A167 );
 a91975a <=( a91974a  and  a91971a );
 a91978a <=( (not A200)  and  A199 );
 a91981a <=( A203  and  A201 );
 a91982a <=( a91981a  and  a91978a );
 a91983a <=( a91982a  and  a91975a );
 a91986a <=( A266  and  (not A265) );
 a91989a <=( (not A268)  and  (not A267) );
 a91990a <=( a91989a  and  a91986a );
 a91993a <=( A300  and  (not A269) );
 a91996a <=( (not A302)  and  (not A301) );
 a91997a <=( a91996a  and  a91993a );
 a91998a <=( a91997a  and  a91990a );
 a92001a <=( A168  and  A169 );
 a92004a <=( (not A166)  and  A167 );
 a92005a <=( a92004a  and  a92001a );
 a92008a <=( (not A200)  and  A199 );
 a92011a <=( A203  and  A201 );
 a92012a <=( a92011a  and  a92008a );
 a92013a <=( a92012a  and  a92005a );
 a92016a <=( (not A266)  and  A265 );
 a92019a <=( (not A268)  and  (not A267) );
 a92020a <=( a92019a  and  a92016a );
 a92023a <=( A300  and  (not A269) );
 a92026a <=( (not A302)  and  (not A301) );
 a92027a <=( a92026a  and  a92023a );
 a92028a <=( a92027a  and  a92020a );
 a92031a <=( A168  and  A169 );
 a92034a <=( (not A166)  and  A167 );
 a92035a <=( a92034a  and  a92031a );
 a92038a <=( (not A200)  and  A199 );
 a92041a <=( (not A202)  and  (not A201) );
 a92042a <=( a92041a  and  a92038a );
 a92043a <=( a92042a  and  a92035a );
 a92046a <=( (not A265)  and  (not A203) );
 a92049a <=( A267  and  A266 );
 a92050a <=( a92049a  and  a92046a );
 a92053a <=( A300  and  A268 );
 a92056a <=( (not A302)  and  (not A301) );
 a92057a <=( a92056a  and  a92053a );
 a92058a <=( a92057a  and  a92050a );
 a92061a <=( A168  and  A169 );
 a92064a <=( (not A166)  and  A167 );
 a92065a <=( a92064a  and  a92061a );
 a92068a <=( (not A200)  and  A199 );
 a92071a <=( (not A202)  and  (not A201) );
 a92072a <=( a92071a  and  a92068a );
 a92073a <=( a92072a  and  a92065a );
 a92076a <=( (not A265)  and  (not A203) );
 a92079a <=( A267  and  A266 );
 a92080a <=( a92079a  and  a92076a );
 a92083a <=( A300  and  A269 );
 a92086a <=( (not A302)  and  (not A301) );
 a92087a <=( a92086a  and  a92083a );
 a92088a <=( a92087a  and  a92080a );
 a92091a <=( A168  and  A169 );
 a92094a <=( (not A166)  and  A167 );
 a92095a <=( a92094a  and  a92091a );
 a92098a <=( (not A200)  and  A199 );
 a92101a <=( (not A202)  and  (not A201) );
 a92102a <=( a92101a  and  a92098a );
 a92103a <=( a92102a  and  a92095a );
 a92106a <=( (not A265)  and  (not A203) );
 a92109a <=( (not A267)  and  A266 );
 a92110a <=( a92109a  and  a92106a );
 a92113a <=( (not A269)  and  (not A268) );
 a92116a <=( A301  and  (not A300) );
 a92117a <=( a92116a  and  a92113a );
 a92118a <=( a92117a  and  a92110a );
 a92121a <=( A168  and  A169 );
 a92124a <=( (not A166)  and  A167 );
 a92125a <=( a92124a  and  a92121a );
 a92128a <=( (not A200)  and  A199 );
 a92131a <=( (not A202)  and  (not A201) );
 a92132a <=( a92131a  and  a92128a );
 a92133a <=( a92132a  and  a92125a );
 a92136a <=( (not A265)  and  (not A203) );
 a92139a <=( (not A267)  and  A266 );
 a92140a <=( a92139a  and  a92136a );
 a92143a <=( (not A269)  and  (not A268) );
 a92146a <=( A302  and  (not A300) );
 a92147a <=( a92146a  and  a92143a );
 a92148a <=( a92147a  and  a92140a );
 a92151a <=( A168  and  A169 );
 a92154a <=( (not A166)  and  A167 );
 a92155a <=( a92154a  and  a92151a );
 a92158a <=( (not A200)  and  A199 );
 a92161a <=( (not A202)  and  (not A201) );
 a92162a <=( a92161a  and  a92158a );
 a92163a <=( a92162a  and  a92155a );
 a92166a <=( (not A265)  and  (not A203) );
 a92169a <=( (not A267)  and  A266 );
 a92170a <=( a92169a  and  a92166a );
 a92173a <=( (not A269)  and  (not A268) );
 a92176a <=( A299  and  A298 );
 a92177a <=( a92176a  and  a92173a );
 a92178a <=( a92177a  and  a92170a );
 a92181a <=( A168  and  A169 );
 a92184a <=( (not A166)  and  A167 );
 a92185a <=( a92184a  and  a92181a );
 a92188a <=( (not A200)  and  A199 );
 a92191a <=( (not A202)  and  (not A201) );
 a92192a <=( a92191a  and  a92188a );
 a92193a <=( a92192a  and  a92185a );
 a92196a <=( (not A265)  and  (not A203) );
 a92199a <=( (not A267)  and  A266 );
 a92200a <=( a92199a  and  a92196a );
 a92203a <=( (not A269)  and  (not A268) );
 a92206a <=( (not A299)  and  (not A298) );
 a92207a <=( a92206a  and  a92203a );
 a92208a <=( a92207a  and  a92200a );
 a92211a <=( A168  and  A169 );
 a92214a <=( (not A166)  and  A167 );
 a92215a <=( a92214a  and  a92211a );
 a92218a <=( (not A200)  and  A199 );
 a92221a <=( (not A202)  and  (not A201) );
 a92222a <=( a92221a  and  a92218a );
 a92223a <=( a92222a  and  a92215a );
 a92226a <=( A265  and  (not A203) );
 a92229a <=( A267  and  (not A266) );
 a92230a <=( a92229a  and  a92226a );
 a92233a <=( A300  and  A268 );
 a92236a <=( (not A302)  and  (not A301) );
 a92237a <=( a92236a  and  a92233a );
 a92238a <=( a92237a  and  a92230a );
 a92241a <=( A168  and  A169 );
 a92244a <=( (not A166)  and  A167 );
 a92245a <=( a92244a  and  a92241a );
 a92248a <=( (not A200)  and  A199 );
 a92251a <=( (not A202)  and  (not A201) );
 a92252a <=( a92251a  and  a92248a );
 a92253a <=( a92252a  and  a92245a );
 a92256a <=( A265  and  (not A203) );
 a92259a <=( A267  and  (not A266) );
 a92260a <=( a92259a  and  a92256a );
 a92263a <=( A300  and  A269 );
 a92266a <=( (not A302)  and  (not A301) );
 a92267a <=( a92266a  and  a92263a );
 a92268a <=( a92267a  and  a92260a );
 a92271a <=( A168  and  A169 );
 a92274a <=( (not A166)  and  A167 );
 a92275a <=( a92274a  and  a92271a );
 a92278a <=( (not A200)  and  A199 );
 a92281a <=( (not A202)  and  (not A201) );
 a92282a <=( a92281a  and  a92278a );
 a92283a <=( a92282a  and  a92275a );
 a92286a <=( A265  and  (not A203) );
 a92289a <=( (not A267)  and  (not A266) );
 a92290a <=( a92289a  and  a92286a );
 a92293a <=( (not A269)  and  (not A268) );
 a92296a <=( A301  and  (not A300) );
 a92297a <=( a92296a  and  a92293a );
 a92298a <=( a92297a  and  a92290a );
 a92301a <=( A168  and  A169 );
 a92304a <=( (not A166)  and  A167 );
 a92305a <=( a92304a  and  a92301a );
 a92308a <=( (not A200)  and  A199 );
 a92311a <=( (not A202)  and  (not A201) );
 a92312a <=( a92311a  and  a92308a );
 a92313a <=( a92312a  and  a92305a );
 a92316a <=( A265  and  (not A203) );
 a92319a <=( (not A267)  and  (not A266) );
 a92320a <=( a92319a  and  a92316a );
 a92323a <=( (not A269)  and  (not A268) );
 a92326a <=( A302  and  (not A300) );
 a92327a <=( a92326a  and  a92323a );
 a92328a <=( a92327a  and  a92320a );
 a92331a <=( A168  and  A169 );
 a92334a <=( (not A166)  and  A167 );
 a92335a <=( a92334a  and  a92331a );
 a92338a <=( (not A200)  and  A199 );
 a92341a <=( (not A202)  and  (not A201) );
 a92342a <=( a92341a  and  a92338a );
 a92343a <=( a92342a  and  a92335a );
 a92346a <=( A265  and  (not A203) );
 a92349a <=( (not A267)  and  (not A266) );
 a92350a <=( a92349a  and  a92346a );
 a92353a <=( (not A269)  and  (not A268) );
 a92356a <=( A299  and  A298 );
 a92357a <=( a92356a  and  a92353a );
 a92358a <=( a92357a  and  a92350a );
 a92361a <=( A168  and  A169 );
 a92364a <=( (not A166)  and  A167 );
 a92365a <=( a92364a  and  a92361a );
 a92368a <=( (not A200)  and  A199 );
 a92371a <=( (not A202)  and  (not A201) );
 a92372a <=( a92371a  and  a92368a );
 a92373a <=( a92372a  and  a92365a );
 a92376a <=( A265  and  (not A203) );
 a92379a <=( (not A267)  and  (not A266) );
 a92380a <=( a92379a  and  a92376a );
 a92383a <=( (not A269)  and  (not A268) );
 a92386a <=( (not A299)  and  (not A298) );
 a92387a <=( a92386a  and  a92383a );
 a92388a <=( a92387a  and  a92380a );
 a92391a <=( A168  and  A169 );
 a92394a <=( A166  and  (not A167) );
 a92395a <=( a92394a  and  a92391a );
 a92398a <=( A200  and  (not A199) );
 a92401a <=( A202  and  A201 );
 a92402a <=( a92401a  and  a92398a );
 a92403a <=( a92402a  and  a92395a );
 a92406a <=( A266  and  (not A265) );
 a92409a <=( (not A268)  and  (not A267) );
 a92410a <=( a92409a  and  a92406a );
 a92413a <=( A300  and  (not A269) );
 a92416a <=( (not A302)  and  (not A301) );
 a92417a <=( a92416a  and  a92413a );
 a92418a <=( a92417a  and  a92410a );
 a92421a <=( A168  and  A169 );
 a92424a <=( A166  and  (not A167) );
 a92425a <=( a92424a  and  a92421a );
 a92428a <=( A200  and  (not A199) );
 a92431a <=( A202  and  A201 );
 a92432a <=( a92431a  and  a92428a );
 a92433a <=( a92432a  and  a92425a );
 a92436a <=( (not A266)  and  A265 );
 a92439a <=( (not A268)  and  (not A267) );
 a92440a <=( a92439a  and  a92436a );
 a92443a <=( A300  and  (not A269) );
 a92446a <=( (not A302)  and  (not A301) );
 a92447a <=( a92446a  and  a92443a );
 a92448a <=( a92447a  and  a92440a );
 a92451a <=( A168  and  A169 );
 a92454a <=( A166  and  (not A167) );
 a92455a <=( a92454a  and  a92451a );
 a92458a <=( A200  and  (not A199) );
 a92461a <=( A203  and  A201 );
 a92462a <=( a92461a  and  a92458a );
 a92463a <=( a92462a  and  a92455a );
 a92466a <=( A266  and  (not A265) );
 a92469a <=( (not A268)  and  (not A267) );
 a92470a <=( a92469a  and  a92466a );
 a92473a <=( A300  and  (not A269) );
 a92476a <=( (not A302)  and  (not A301) );
 a92477a <=( a92476a  and  a92473a );
 a92478a <=( a92477a  and  a92470a );
 a92481a <=( A168  and  A169 );
 a92484a <=( A166  and  (not A167) );
 a92485a <=( a92484a  and  a92481a );
 a92488a <=( A200  and  (not A199) );
 a92491a <=( A203  and  A201 );
 a92492a <=( a92491a  and  a92488a );
 a92493a <=( a92492a  and  a92485a );
 a92496a <=( (not A266)  and  A265 );
 a92499a <=( (not A268)  and  (not A267) );
 a92500a <=( a92499a  and  a92496a );
 a92503a <=( A300  and  (not A269) );
 a92506a <=( (not A302)  and  (not A301) );
 a92507a <=( a92506a  and  a92503a );
 a92508a <=( a92507a  and  a92500a );
 a92511a <=( A168  and  A169 );
 a92514a <=( A166  and  (not A167) );
 a92515a <=( a92514a  and  a92511a );
 a92518a <=( A200  and  (not A199) );
 a92521a <=( (not A202)  and  (not A201) );
 a92522a <=( a92521a  and  a92518a );
 a92523a <=( a92522a  and  a92515a );
 a92526a <=( (not A265)  and  (not A203) );
 a92529a <=( A267  and  A266 );
 a92530a <=( a92529a  and  a92526a );
 a92533a <=( A300  and  A268 );
 a92536a <=( (not A302)  and  (not A301) );
 a92537a <=( a92536a  and  a92533a );
 a92538a <=( a92537a  and  a92530a );
 a92541a <=( A168  and  A169 );
 a92544a <=( A166  and  (not A167) );
 a92545a <=( a92544a  and  a92541a );
 a92548a <=( A200  and  (not A199) );
 a92551a <=( (not A202)  and  (not A201) );
 a92552a <=( a92551a  and  a92548a );
 a92553a <=( a92552a  and  a92545a );
 a92556a <=( (not A265)  and  (not A203) );
 a92559a <=( A267  and  A266 );
 a92560a <=( a92559a  and  a92556a );
 a92563a <=( A300  and  A269 );
 a92566a <=( (not A302)  and  (not A301) );
 a92567a <=( a92566a  and  a92563a );
 a92568a <=( a92567a  and  a92560a );
 a92571a <=( A168  and  A169 );
 a92574a <=( A166  and  (not A167) );
 a92575a <=( a92574a  and  a92571a );
 a92578a <=( A200  and  (not A199) );
 a92581a <=( (not A202)  and  (not A201) );
 a92582a <=( a92581a  and  a92578a );
 a92583a <=( a92582a  and  a92575a );
 a92586a <=( (not A265)  and  (not A203) );
 a92589a <=( (not A267)  and  A266 );
 a92590a <=( a92589a  and  a92586a );
 a92593a <=( (not A269)  and  (not A268) );
 a92596a <=( A301  and  (not A300) );
 a92597a <=( a92596a  and  a92593a );
 a92598a <=( a92597a  and  a92590a );
 a92601a <=( A168  and  A169 );
 a92604a <=( A166  and  (not A167) );
 a92605a <=( a92604a  and  a92601a );
 a92608a <=( A200  and  (not A199) );
 a92611a <=( (not A202)  and  (not A201) );
 a92612a <=( a92611a  and  a92608a );
 a92613a <=( a92612a  and  a92605a );
 a92616a <=( (not A265)  and  (not A203) );
 a92619a <=( (not A267)  and  A266 );
 a92620a <=( a92619a  and  a92616a );
 a92623a <=( (not A269)  and  (not A268) );
 a92626a <=( A302  and  (not A300) );
 a92627a <=( a92626a  and  a92623a );
 a92628a <=( a92627a  and  a92620a );
 a92631a <=( A168  and  A169 );
 a92634a <=( A166  and  (not A167) );
 a92635a <=( a92634a  and  a92631a );
 a92638a <=( A200  and  (not A199) );
 a92641a <=( (not A202)  and  (not A201) );
 a92642a <=( a92641a  and  a92638a );
 a92643a <=( a92642a  and  a92635a );
 a92646a <=( (not A265)  and  (not A203) );
 a92649a <=( (not A267)  and  A266 );
 a92650a <=( a92649a  and  a92646a );
 a92653a <=( (not A269)  and  (not A268) );
 a92656a <=( A299  and  A298 );
 a92657a <=( a92656a  and  a92653a );
 a92658a <=( a92657a  and  a92650a );
 a92661a <=( A168  and  A169 );
 a92664a <=( A166  and  (not A167) );
 a92665a <=( a92664a  and  a92661a );
 a92668a <=( A200  and  (not A199) );
 a92671a <=( (not A202)  and  (not A201) );
 a92672a <=( a92671a  and  a92668a );
 a92673a <=( a92672a  and  a92665a );
 a92676a <=( (not A265)  and  (not A203) );
 a92679a <=( (not A267)  and  A266 );
 a92680a <=( a92679a  and  a92676a );
 a92683a <=( (not A269)  and  (not A268) );
 a92686a <=( (not A299)  and  (not A298) );
 a92687a <=( a92686a  and  a92683a );
 a92688a <=( a92687a  and  a92680a );
 a92691a <=( A168  and  A169 );
 a92694a <=( A166  and  (not A167) );
 a92695a <=( a92694a  and  a92691a );
 a92698a <=( A200  and  (not A199) );
 a92701a <=( (not A202)  and  (not A201) );
 a92702a <=( a92701a  and  a92698a );
 a92703a <=( a92702a  and  a92695a );
 a92706a <=( A265  and  (not A203) );
 a92709a <=( A267  and  (not A266) );
 a92710a <=( a92709a  and  a92706a );
 a92713a <=( A300  and  A268 );
 a92716a <=( (not A302)  and  (not A301) );
 a92717a <=( a92716a  and  a92713a );
 a92718a <=( a92717a  and  a92710a );
 a92721a <=( A168  and  A169 );
 a92724a <=( A166  and  (not A167) );
 a92725a <=( a92724a  and  a92721a );
 a92728a <=( A200  and  (not A199) );
 a92731a <=( (not A202)  and  (not A201) );
 a92732a <=( a92731a  and  a92728a );
 a92733a <=( a92732a  and  a92725a );
 a92736a <=( A265  and  (not A203) );
 a92739a <=( A267  and  (not A266) );
 a92740a <=( a92739a  and  a92736a );
 a92743a <=( A300  and  A269 );
 a92746a <=( (not A302)  and  (not A301) );
 a92747a <=( a92746a  and  a92743a );
 a92748a <=( a92747a  and  a92740a );
 a92751a <=( A168  and  A169 );
 a92754a <=( A166  and  (not A167) );
 a92755a <=( a92754a  and  a92751a );
 a92758a <=( A200  and  (not A199) );
 a92761a <=( (not A202)  and  (not A201) );
 a92762a <=( a92761a  and  a92758a );
 a92763a <=( a92762a  and  a92755a );
 a92766a <=( A265  and  (not A203) );
 a92769a <=( (not A267)  and  (not A266) );
 a92770a <=( a92769a  and  a92766a );
 a92773a <=( (not A269)  and  (not A268) );
 a92776a <=( A301  and  (not A300) );
 a92777a <=( a92776a  and  a92773a );
 a92778a <=( a92777a  and  a92770a );
 a92781a <=( A168  and  A169 );
 a92784a <=( A166  and  (not A167) );
 a92785a <=( a92784a  and  a92781a );
 a92788a <=( A200  and  (not A199) );
 a92791a <=( (not A202)  and  (not A201) );
 a92792a <=( a92791a  and  a92788a );
 a92793a <=( a92792a  and  a92785a );
 a92796a <=( A265  and  (not A203) );
 a92799a <=( (not A267)  and  (not A266) );
 a92800a <=( a92799a  and  a92796a );
 a92803a <=( (not A269)  and  (not A268) );
 a92806a <=( A302  and  (not A300) );
 a92807a <=( a92806a  and  a92803a );
 a92808a <=( a92807a  and  a92800a );
 a92811a <=( A168  and  A169 );
 a92814a <=( A166  and  (not A167) );
 a92815a <=( a92814a  and  a92811a );
 a92818a <=( A200  and  (not A199) );
 a92821a <=( (not A202)  and  (not A201) );
 a92822a <=( a92821a  and  a92818a );
 a92823a <=( a92822a  and  a92815a );
 a92826a <=( A265  and  (not A203) );
 a92829a <=( (not A267)  and  (not A266) );
 a92830a <=( a92829a  and  a92826a );
 a92833a <=( (not A269)  and  (not A268) );
 a92836a <=( A299  and  A298 );
 a92837a <=( a92836a  and  a92833a );
 a92838a <=( a92837a  and  a92830a );
 a92841a <=( A168  and  A169 );
 a92844a <=( A166  and  (not A167) );
 a92845a <=( a92844a  and  a92841a );
 a92848a <=( A200  and  (not A199) );
 a92851a <=( (not A202)  and  (not A201) );
 a92852a <=( a92851a  and  a92848a );
 a92853a <=( a92852a  and  a92845a );
 a92856a <=( A265  and  (not A203) );
 a92859a <=( (not A267)  and  (not A266) );
 a92860a <=( a92859a  and  a92856a );
 a92863a <=( (not A269)  and  (not A268) );
 a92866a <=( (not A299)  and  (not A298) );
 a92867a <=( a92866a  and  a92863a );
 a92868a <=( a92867a  and  a92860a );
 a92871a <=( A168  and  A169 );
 a92874a <=( A166  and  (not A167) );
 a92875a <=( a92874a  and  a92871a );
 a92878a <=( (not A200)  and  A199 );
 a92881a <=( A202  and  A201 );
 a92882a <=( a92881a  and  a92878a );
 a92883a <=( a92882a  and  a92875a );
 a92886a <=( A266  and  (not A265) );
 a92889a <=( (not A268)  and  (not A267) );
 a92890a <=( a92889a  and  a92886a );
 a92893a <=( A300  and  (not A269) );
 a92896a <=( (not A302)  and  (not A301) );
 a92897a <=( a92896a  and  a92893a );
 a92898a <=( a92897a  and  a92890a );
 a92901a <=( A168  and  A169 );
 a92904a <=( A166  and  (not A167) );
 a92905a <=( a92904a  and  a92901a );
 a92908a <=( (not A200)  and  A199 );
 a92911a <=( A202  and  A201 );
 a92912a <=( a92911a  and  a92908a );
 a92913a <=( a92912a  and  a92905a );
 a92916a <=( (not A266)  and  A265 );
 a92919a <=( (not A268)  and  (not A267) );
 a92920a <=( a92919a  and  a92916a );
 a92923a <=( A300  and  (not A269) );
 a92926a <=( (not A302)  and  (not A301) );
 a92927a <=( a92926a  and  a92923a );
 a92928a <=( a92927a  and  a92920a );
 a92931a <=( A168  and  A169 );
 a92934a <=( A166  and  (not A167) );
 a92935a <=( a92934a  and  a92931a );
 a92938a <=( (not A200)  and  A199 );
 a92941a <=( A203  and  A201 );
 a92942a <=( a92941a  and  a92938a );
 a92943a <=( a92942a  and  a92935a );
 a92946a <=( A266  and  (not A265) );
 a92949a <=( (not A268)  and  (not A267) );
 a92950a <=( a92949a  and  a92946a );
 a92953a <=( A300  and  (not A269) );
 a92956a <=( (not A302)  and  (not A301) );
 a92957a <=( a92956a  and  a92953a );
 a92958a <=( a92957a  and  a92950a );
 a92961a <=( A168  and  A169 );
 a92964a <=( A166  and  (not A167) );
 a92965a <=( a92964a  and  a92961a );
 a92968a <=( (not A200)  and  A199 );
 a92971a <=( A203  and  A201 );
 a92972a <=( a92971a  and  a92968a );
 a92973a <=( a92972a  and  a92965a );
 a92976a <=( (not A266)  and  A265 );
 a92979a <=( (not A268)  and  (not A267) );
 a92980a <=( a92979a  and  a92976a );
 a92983a <=( A300  and  (not A269) );
 a92986a <=( (not A302)  and  (not A301) );
 a92987a <=( a92986a  and  a92983a );
 a92988a <=( a92987a  and  a92980a );
 a92991a <=( A168  and  A169 );
 a92994a <=( A166  and  (not A167) );
 a92995a <=( a92994a  and  a92991a );
 a92998a <=( (not A200)  and  A199 );
 a93001a <=( (not A202)  and  (not A201) );
 a93002a <=( a93001a  and  a92998a );
 a93003a <=( a93002a  and  a92995a );
 a93006a <=( (not A265)  and  (not A203) );
 a93009a <=( A267  and  A266 );
 a93010a <=( a93009a  and  a93006a );
 a93013a <=( A300  and  A268 );
 a93016a <=( (not A302)  and  (not A301) );
 a93017a <=( a93016a  and  a93013a );
 a93018a <=( a93017a  and  a93010a );
 a93021a <=( A168  and  A169 );
 a93024a <=( A166  and  (not A167) );
 a93025a <=( a93024a  and  a93021a );
 a93028a <=( (not A200)  and  A199 );
 a93031a <=( (not A202)  and  (not A201) );
 a93032a <=( a93031a  and  a93028a );
 a93033a <=( a93032a  and  a93025a );
 a93036a <=( (not A265)  and  (not A203) );
 a93039a <=( A267  and  A266 );
 a93040a <=( a93039a  and  a93036a );
 a93043a <=( A300  and  A269 );
 a93046a <=( (not A302)  and  (not A301) );
 a93047a <=( a93046a  and  a93043a );
 a93048a <=( a93047a  and  a93040a );
 a93051a <=( A168  and  A169 );
 a93054a <=( A166  and  (not A167) );
 a93055a <=( a93054a  and  a93051a );
 a93058a <=( (not A200)  and  A199 );
 a93061a <=( (not A202)  and  (not A201) );
 a93062a <=( a93061a  and  a93058a );
 a93063a <=( a93062a  and  a93055a );
 a93066a <=( (not A265)  and  (not A203) );
 a93069a <=( (not A267)  and  A266 );
 a93070a <=( a93069a  and  a93066a );
 a93073a <=( (not A269)  and  (not A268) );
 a93076a <=( A301  and  (not A300) );
 a93077a <=( a93076a  and  a93073a );
 a93078a <=( a93077a  and  a93070a );
 a93081a <=( A168  and  A169 );
 a93084a <=( A166  and  (not A167) );
 a93085a <=( a93084a  and  a93081a );
 a93088a <=( (not A200)  and  A199 );
 a93091a <=( (not A202)  and  (not A201) );
 a93092a <=( a93091a  and  a93088a );
 a93093a <=( a93092a  and  a93085a );
 a93096a <=( (not A265)  and  (not A203) );
 a93099a <=( (not A267)  and  A266 );
 a93100a <=( a93099a  and  a93096a );
 a93103a <=( (not A269)  and  (not A268) );
 a93106a <=( A302  and  (not A300) );
 a93107a <=( a93106a  and  a93103a );
 a93108a <=( a93107a  and  a93100a );
 a93111a <=( A168  and  A169 );
 a93114a <=( A166  and  (not A167) );
 a93115a <=( a93114a  and  a93111a );
 a93118a <=( (not A200)  and  A199 );
 a93121a <=( (not A202)  and  (not A201) );
 a93122a <=( a93121a  and  a93118a );
 a93123a <=( a93122a  and  a93115a );
 a93126a <=( (not A265)  and  (not A203) );
 a93129a <=( (not A267)  and  A266 );
 a93130a <=( a93129a  and  a93126a );
 a93133a <=( (not A269)  and  (not A268) );
 a93136a <=( A299  and  A298 );
 a93137a <=( a93136a  and  a93133a );
 a93138a <=( a93137a  and  a93130a );
 a93141a <=( A168  and  A169 );
 a93144a <=( A166  and  (not A167) );
 a93145a <=( a93144a  and  a93141a );
 a93148a <=( (not A200)  and  A199 );
 a93151a <=( (not A202)  and  (not A201) );
 a93152a <=( a93151a  and  a93148a );
 a93153a <=( a93152a  and  a93145a );
 a93156a <=( (not A265)  and  (not A203) );
 a93159a <=( (not A267)  and  A266 );
 a93160a <=( a93159a  and  a93156a );
 a93163a <=( (not A269)  and  (not A268) );
 a93166a <=( (not A299)  and  (not A298) );
 a93167a <=( a93166a  and  a93163a );
 a93168a <=( a93167a  and  a93160a );
 a93171a <=( A168  and  A169 );
 a93174a <=( A166  and  (not A167) );
 a93175a <=( a93174a  and  a93171a );
 a93178a <=( (not A200)  and  A199 );
 a93181a <=( (not A202)  and  (not A201) );
 a93182a <=( a93181a  and  a93178a );
 a93183a <=( a93182a  and  a93175a );
 a93186a <=( A265  and  (not A203) );
 a93189a <=( A267  and  (not A266) );
 a93190a <=( a93189a  and  a93186a );
 a93193a <=( A300  and  A268 );
 a93196a <=( (not A302)  and  (not A301) );
 a93197a <=( a93196a  and  a93193a );
 a93198a <=( a93197a  and  a93190a );
 a93201a <=( A168  and  A169 );
 a93204a <=( A166  and  (not A167) );
 a93205a <=( a93204a  and  a93201a );
 a93208a <=( (not A200)  and  A199 );
 a93211a <=( (not A202)  and  (not A201) );
 a93212a <=( a93211a  and  a93208a );
 a93213a <=( a93212a  and  a93205a );
 a93216a <=( A265  and  (not A203) );
 a93219a <=( A267  and  (not A266) );
 a93220a <=( a93219a  and  a93216a );
 a93223a <=( A300  and  A269 );
 a93226a <=( (not A302)  and  (not A301) );
 a93227a <=( a93226a  and  a93223a );
 a93228a <=( a93227a  and  a93220a );
 a93231a <=( A168  and  A169 );
 a93234a <=( A166  and  (not A167) );
 a93235a <=( a93234a  and  a93231a );
 a93238a <=( (not A200)  and  A199 );
 a93241a <=( (not A202)  and  (not A201) );
 a93242a <=( a93241a  and  a93238a );
 a93243a <=( a93242a  and  a93235a );
 a93246a <=( A265  and  (not A203) );
 a93249a <=( (not A267)  and  (not A266) );
 a93250a <=( a93249a  and  a93246a );
 a93253a <=( (not A269)  and  (not A268) );
 a93256a <=( A301  and  (not A300) );
 a93257a <=( a93256a  and  a93253a );
 a93258a <=( a93257a  and  a93250a );
 a93261a <=( A168  and  A169 );
 a93264a <=( A166  and  (not A167) );
 a93265a <=( a93264a  and  a93261a );
 a93268a <=( (not A200)  and  A199 );
 a93271a <=( (not A202)  and  (not A201) );
 a93272a <=( a93271a  and  a93268a );
 a93273a <=( a93272a  and  a93265a );
 a93276a <=( A265  and  (not A203) );
 a93279a <=( (not A267)  and  (not A266) );
 a93280a <=( a93279a  and  a93276a );
 a93283a <=( (not A269)  and  (not A268) );
 a93286a <=( A302  and  (not A300) );
 a93287a <=( a93286a  and  a93283a );
 a93288a <=( a93287a  and  a93280a );
 a93291a <=( A168  and  A169 );
 a93294a <=( A166  and  (not A167) );
 a93295a <=( a93294a  and  a93291a );
 a93298a <=( (not A200)  and  A199 );
 a93301a <=( (not A202)  and  (not A201) );
 a93302a <=( a93301a  and  a93298a );
 a93303a <=( a93302a  and  a93295a );
 a93306a <=( A265  and  (not A203) );
 a93309a <=( (not A267)  and  (not A266) );
 a93310a <=( a93309a  and  a93306a );
 a93313a <=( (not A269)  and  (not A268) );
 a93316a <=( A299  and  A298 );
 a93317a <=( a93316a  and  a93313a );
 a93318a <=( a93317a  and  a93310a );
 a93321a <=( A168  and  A169 );
 a93324a <=( A166  and  (not A167) );
 a93325a <=( a93324a  and  a93321a );
 a93328a <=( (not A200)  and  A199 );
 a93331a <=( (not A202)  and  (not A201) );
 a93332a <=( a93331a  and  a93328a );
 a93333a <=( a93332a  and  a93325a );
 a93336a <=( A265  and  (not A203) );
 a93339a <=( (not A267)  and  (not A266) );
 a93340a <=( a93339a  and  a93336a );
 a93343a <=( (not A269)  and  (not A268) );
 a93346a <=( (not A299)  and  (not A298) );
 a93347a <=( a93346a  and  a93343a );
 a93348a <=( a93347a  and  a93340a );
 a93351a <=( (not A169)  and  A170 );
 a93354a <=( (not A199)  and  A168 );
 a93355a <=( a93354a  and  a93351a );
 a93358a <=( (not A201)  and  A200 );
 a93361a <=( (not A203)  and  (not A202) );
 a93362a <=( a93361a  and  a93358a );
 a93363a <=( a93362a  and  a93355a );
 a93366a <=( (not A268)  and  A267 );
 a93369a <=( A298  and  (not A269) );
 a93370a <=( a93369a  and  a93366a );
 a93373a <=( (not A300)  and  (not A299) );
 a93376a <=( (not A302)  and  (not A301) );
 a93377a <=( a93376a  and  a93373a );
 a93378a <=( a93377a  and  a93370a );
 a93381a <=( (not A169)  and  A170 );
 a93384a <=( (not A199)  and  A168 );
 a93385a <=( a93384a  and  a93381a );
 a93388a <=( (not A201)  and  A200 );
 a93391a <=( (not A203)  and  (not A202) );
 a93392a <=( a93391a  and  a93388a );
 a93393a <=( a93392a  and  a93385a );
 a93396a <=( (not A268)  and  A267 );
 a93399a <=( (not A298)  and  (not A269) );
 a93400a <=( a93399a  and  a93396a );
 a93403a <=( (not A300)  and  A299 );
 a93406a <=( (not A302)  and  (not A301) );
 a93407a <=( a93406a  and  a93403a );
 a93408a <=( a93407a  and  a93400a );
 a93411a <=( (not A169)  and  A170 );
 a93414a <=( A199  and  A168 );
 a93415a <=( a93414a  and  a93411a );
 a93418a <=( (not A201)  and  (not A200) );
 a93421a <=( (not A203)  and  (not A202) );
 a93422a <=( a93421a  and  a93418a );
 a93423a <=( a93422a  and  a93415a );
 a93426a <=( (not A268)  and  A267 );
 a93429a <=( A298  and  (not A269) );
 a93430a <=( a93429a  and  a93426a );
 a93433a <=( (not A300)  and  (not A299) );
 a93436a <=( (not A302)  and  (not A301) );
 a93437a <=( a93436a  and  a93433a );
 a93438a <=( a93437a  and  a93430a );
 a93441a <=( (not A169)  and  A170 );
 a93444a <=( A199  and  A168 );
 a93445a <=( a93444a  and  a93441a );
 a93448a <=( (not A201)  and  (not A200) );
 a93451a <=( (not A203)  and  (not A202) );
 a93452a <=( a93451a  and  a93448a );
 a93453a <=( a93452a  and  a93445a );
 a93456a <=( (not A268)  and  A267 );
 a93459a <=( (not A298)  and  (not A269) );
 a93460a <=( a93459a  and  a93456a );
 a93463a <=( (not A300)  and  A299 );
 a93466a <=( (not A302)  and  (not A301) );
 a93467a <=( a93466a  and  a93463a );
 a93468a <=( a93467a  and  a93460a );
 a93471a <=( (not A169)  and  A170 );
 a93474a <=( A167  and  (not A168) );
 a93475a <=( a93474a  and  a93471a );
 a93478a <=( A201  and  (not A166) );
 a93481a <=( (not A203)  and  (not A202) );
 a93482a <=( a93481a  and  a93478a );
 a93483a <=( a93482a  and  a93475a );
 a93486a <=( (not A268)  and  A267 );
 a93489a <=( A298  and  (not A269) );
 a93490a <=( a93489a  and  a93486a );
 a93493a <=( (not A300)  and  (not A299) );
 a93496a <=( (not A302)  and  (not A301) );
 a93497a <=( a93496a  and  a93493a );
 a93498a <=( a93497a  and  a93490a );
 a93501a <=( (not A169)  and  A170 );
 a93504a <=( A167  and  (not A168) );
 a93505a <=( a93504a  and  a93501a );
 a93508a <=( A201  and  (not A166) );
 a93511a <=( (not A203)  and  (not A202) );
 a93512a <=( a93511a  and  a93508a );
 a93513a <=( a93512a  and  a93505a );
 a93516a <=( (not A268)  and  A267 );
 a93519a <=( (not A298)  and  (not A269) );
 a93520a <=( a93519a  and  a93516a );
 a93523a <=( (not A300)  and  A299 );
 a93526a <=( (not A302)  and  (not A301) );
 a93527a <=( a93526a  and  a93523a );
 a93528a <=( a93527a  and  a93520a );
 a93531a <=( (not A169)  and  A170 );
 a93534a <=( A167  and  (not A168) );
 a93535a <=( a93534a  and  a93531a );
 a93538a <=( (not A199)  and  (not A166) );
 a93541a <=( A201  and  A200 );
 a93542a <=( a93541a  and  a93538a );
 a93543a <=( a93542a  and  a93535a );
 a93546a <=( (not A265)  and  A202 );
 a93549a <=( A267  and  A266 );
 a93550a <=( a93549a  and  a93546a );
 a93553a <=( A300  and  A268 );
 a93556a <=( (not A302)  and  (not A301) );
 a93557a <=( a93556a  and  a93553a );
 a93558a <=( a93557a  and  a93550a );
 a93561a <=( (not A169)  and  A170 );
 a93564a <=( A167  and  (not A168) );
 a93565a <=( a93564a  and  a93561a );
 a93568a <=( (not A199)  and  (not A166) );
 a93571a <=( A201  and  A200 );
 a93572a <=( a93571a  and  a93568a );
 a93573a <=( a93572a  and  a93565a );
 a93576a <=( (not A265)  and  A202 );
 a93579a <=( A267  and  A266 );
 a93580a <=( a93579a  and  a93576a );
 a93583a <=( A300  and  A269 );
 a93586a <=( (not A302)  and  (not A301) );
 a93587a <=( a93586a  and  a93583a );
 a93588a <=( a93587a  and  a93580a );
 a93591a <=( (not A169)  and  A170 );
 a93594a <=( A167  and  (not A168) );
 a93595a <=( a93594a  and  a93591a );
 a93598a <=( (not A199)  and  (not A166) );
 a93601a <=( A201  and  A200 );
 a93602a <=( a93601a  and  a93598a );
 a93603a <=( a93602a  and  a93595a );
 a93606a <=( (not A265)  and  A202 );
 a93609a <=( (not A267)  and  A266 );
 a93610a <=( a93609a  and  a93606a );
 a93613a <=( (not A269)  and  (not A268) );
 a93616a <=( A301  and  (not A300) );
 a93617a <=( a93616a  and  a93613a );
 a93618a <=( a93617a  and  a93610a );
 a93621a <=( (not A169)  and  A170 );
 a93624a <=( A167  and  (not A168) );
 a93625a <=( a93624a  and  a93621a );
 a93628a <=( (not A199)  and  (not A166) );
 a93631a <=( A201  and  A200 );
 a93632a <=( a93631a  and  a93628a );
 a93633a <=( a93632a  and  a93625a );
 a93636a <=( (not A265)  and  A202 );
 a93639a <=( (not A267)  and  A266 );
 a93640a <=( a93639a  and  a93636a );
 a93643a <=( (not A269)  and  (not A268) );
 a93646a <=( A302  and  (not A300) );
 a93647a <=( a93646a  and  a93643a );
 a93648a <=( a93647a  and  a93640a );
 a93651a <=( (not A169)  and  A170 );
 a93654a <=( A167  and  (not A168) );
 a93655a <=( a93654a  and  a93651a );
 a93658a <=( (not A199)  and  (not A166) );
 a93661a <=( A201  and  A200 );
 a93662a <=( a93661a  and  a93658a );
 a93663a <=( a93662a  and  a93655a );
 a93666a <=( (not A265)  and  A202 );
 a93669a <=( (not A267)  and  A266 );
 a93670a <=( a93669a  and  a93666a );
 a93673a <=( (not A269)  and  (not A268) );
 a93676a <=( A299  and  A298 );
 a93677a <=( a93676a  and  a93673a );
 a93678a <=( a93677a  and  a93670a );
 a93681a <=( (not A169)  and  A170 );
 a93684a <=( A167  and  (not A168) );
 a93685a <=( a93684a  and  a93681a );
 a93688a <=( (not A199)  and  (not A166) );
 a93691a <=( A201  and  A200 );
 a93692a <=( a93691a  and  a93688a );
 a93693a <=( a93692a  and  a93685a );
 a93696a <=( (not A265)  and  A202 );
 a93699a <=( (not A267)  and  A266 );
 a93700a <=( a93699a  and  a93696a );
 a93703a <=( (not A269)  and  (not A268) );
 a93706a <=( (not A299)  and  (not A298) );
 a93707a <=( a93706a  and  a93703a );
 a93708a <=( a93707a  and  a93700a );
 a93711a <=( (not A169)  and  A170 );
 a93714a <=( A167  and  (not A168) );
 a93715a <=( a93714a  and  a93711a );
 a93718a <=( (not A199)  and  (not A166) );
 a93721a <=( A201  and  A200 );
 a93722a <=( a93721a  and  a93718a );
 a93723a <=( a93722a  and  a93715a );
 a93726a <=( A265  and  A202 );
 a93729a <=( A267  and  (not A266) );
 a93730a <=( a93729a  and  a93726a );
 a93733a <=( A300  and  A268 );
 a93736a <=( (not A302)  and  (not A301) );
 a93737a <=( a93736a  and  a93733a );
 a93738a <=( a93737a  and  a93730a );
 a93741a <=( (not A169)  and  A170 );
 a93744a <=( A167  and  (not A168) );
 a93745a <=( a93744a  and  a93741a );
 a93748a <=( (not A199)  and  (not A166) );
 a93751a <=( A201  and  A200 );
 a93752a <=( a93751a  and  a93748a );
 a93753a <=( a93752a  and  a93745a );
 a93756a <=( A265  and  A202 );
 a93759a <=( A267  and  (not A266) );
 a93760a <=( a93759a  and  a93756a );
 a93763a <=( A300  and  A269 );
 a93766a <=( (not A302)  and  (not A301) );
 a93767a <=( a93766a  and  a93763a );
 a93768a <=( a93767a  and  a93760a );
 a93771a <=( (not A169)  and  A170 );
 a93774a <=( A167  and  (not A168) );
 a93775a <=( a93774a  and  a93771a );
 a93778a <=( (not A199)  and  (not A166) );
 a93781a <=( A201  and  A200 );
 a93782a <=( a93781a  and  a93778a );
 a93783a <=( a93782a  and  a93775a );
 a93786a <=( A265  and  A202 );
 a93789a <=( (not A267)  and  (not A266) );
 a93790a <=( a93789a  and  a93786a );
 a93793a <=( (not A269)  and  (not A268) );
 a93796a <=( A301  and  (not A300) );
 a93797a <=( a93796a  and  a93793a );
 a93798a <=( a93797a  and  a93790a );
 a93801a <=( (not A169)  and  A170 );
 a93804a <=( A167  and  (not A168) );
 a93805a <=( a93804a  and  a93801a );
 a93808a <=( (not A199)  and  (not A166) );
 a93811a <=( A201  and  A200 );
 a93812a <=( a93811a  and  a93808a );
 a93813a <=( a93812a  and  a93805a );
 a93816a <=( A265  and  A202 );
 a93819a <=( (not A267)  and  (not A266) );
 a93820a <=( a93819a  and  a93816a );
 a93823a <=( (not A269)  and  (not A268) );
 a93826a <=( A302  and  (not A300) );
 a93827a <=( a93826a  and  a93823a );
 a93828a <=( a93827a  and  a93820a );
 a93831a <=( (not A169)  and  A170 );
 a93834a <=( A167  and  (not A168) );
 a93835a <=( a93834a  and  a93831a );
 a93838a <=( (not A199)  and  (not A166) );
 a93841a <=( A201  and  A200 );
 a93842a <=( a93841a  and  a93838a );
 a93843a <=( a93842a  and  a93835a );
 a93846a <=( A265  and  A202 );
 a93849a <=( (not A267)  and  (not A266) );
 a93850a <=( a93849a  and  a93846a );
 a93853a <=( (not A269)  and  (not A268) );
 a93856a <=( A299  and  A298 );
 a93857a <=( a93856a  and  a93853a );
 a93858a <=( a93857a  and  a93850a );
 a93861a <=( (not A169)  and  A170 );
 a93864a <=( A167  and  (not A168) );
 a93865a <=( a93864a  and  a93861a );
 a93868a <=( (not A199)  and  (not A166) );
 a93871a <=( A201  and  A200 );
 a93872a <=( a93871a  and  a93868a );
 a93873a <=( a93872a  and  a93865a );
 a93876a <=( A265  and  A202 );
 a93879a <=( (not A267)  and  (not A266) );
 a93880a <=( a93879a  and  a93876a );
 a93883a <=( (not A269)  and  (not A268) );
 a93886a <=( (not A299)  and  (not A298) );
 a93887a <=( a93886a  and  a93883a );
 a93888a <=( a93887a  and  a93880a );
 a93891a <=( (not A169)  and  A170 );
 a93894a <=( A167  and  (not A168) );
 a93895a <=( a93894a  and  a93891a );
 a93898a <=( (not A199)  and  (not A166) );
 a93901a <=( A201  and  A200 );
 a93902a <=( a93901a  and  a93898a );
 a93903a <=( a93902a  and  a93895a );
 a93906a <=( (not A265)  and  A203 );
 a93909a <=( A267  and  A266 );
 a93910a <=( a93909a  and  a93906a );
 a93913a <=( A300  and  A268 );
 a93916a <=( (not A302)  and  (not A301) );
 a93917a <=( a93916a  and  a93913a );
 a93918a <=( a93917a  and  a93910a );
 a93921a <=( (not A169)  and  A170 );
 a93924a <=( A167  and  (not A168) );
 a93925a <=( a93924a  and  a93921a );
 a93928a <=( (not A199)  and  (not A166) );
 a93931a <=( A201  and  A200 );
 a93932a <=( a93931a  and  a93928a );
 a93933a <=( a93932a  and  a93925a );
 a93936a <=( (not A265)  and  A203 );
 a93939a <=( A267  and  A266 );
 a93940a <=( a93939a  and  a93936a );
 a93943a <=( A300  and  A269 );
 a93946a <=( (not A302)  and  (not A301) );
 a93947a <=( a93946a  and  a93943a );
 a93948a <=( a93947a  and  a93940a );
 a93951a <=( (not A169)  and  A170 );
 a93954a <=( A167  and  (not A168) );
 a93955a <=( a93954a  and  a93951a );
 a93958a <=( (not A199)  and  (not A166) );
 a93961a <=( A201  and  A200 );
 a93962a <=( a93961a  and  a93958a );
 a93963a <=( a93962a  and  a93955a );
 a93966a <=( (not A265)  and  A203 );
 a93969a <=( (not A267)  and  A266 );
 a93970a <=( a93969a  and  a93966a );
 a93973a <=( (not A269)  and  (not A268) );
 a93976a <=( A301  and  (not A300) );
 a93977a <=( a93976a  and  a93973a );
 a93978a <=( a93977a  and  a93970a );
 a93981a <=( (not A169)  and  A170 );
 a93984a <=( A167  and  (not A168) );
 a93985a <=( a93984a  and  a93981a );
 a93988a <=( (not A199)  and  (not A166) );
 a93991a <=( A201  and  A200 );
 a93992a <=( a93991a  and  a93988a );
 a93993a <=( a93992a  and  a93985a );
 a93996a <=( (not A265)  and  A203 );
 a93999a <=( (not A267)  and  A266 );
 a94000a <=( a93999a  and  a93996a );
 a94003a <=( (not A269)  and  (not A268) );
 a94006a <=( A302  and  (not A300) );
 a94007a <=( a94006a  and  a94003a );
 a94008a <=( a94007a  and  a94000a );
 a94011a <=( (not A169)  and  A170 );
 a94014a <=( A167  and  (not A168) );
 a94015a <=( a94014a  and  a94011a );
 a94018a <=( (not A199)  and  (not A166) );
 a94021a <=( A201  and  A200 );
 a94022a <=( a94021a  and  a94018a );
 a94023a <=( a94022a  and  a94015a );
 a94026a <=( (not A265)  and  A203 );
 a94029a <=( (not A267)  and  A266 );
 a94030a <=( a94029a  and  a94026a );
 a94033a <=( (not A269)  and  (not A268) );
 a94036a <=( A299  and  A298 );
 a94037a <=( a94036a  and  a94033a );
 a94038a <=( a94037a  and  a94030a );
 a94041a <=( (not A169)  and  A170 );
 a94044a <=( A167  and  (not A168) );
 a94045a <=( a94044a  and  a94041a );
 a94048a <=( (not A199)  and  (not A166) );
 a94051a <=( A201  and  A200 );
 a94052a <=( a94051a  and  a94048a );
 a94053a <=( a94052a  and  a94045a );
 a94056a <=( (not A265)  and  A203 );
 a94059a <=( (not A267)  and  A266 );
 a94060a <=( a94059a  and  a94056a );
 a94063a <=( (not A269)  and  (not A268) );
 a94066a <=( (not A299)  and  (not A298) );
 a94067a <=( a94066a  and  a94063a );
 a94068a <=( a94067a  and  a94060a );
 a94071a <=( (not A169)  and  A170 );
 a94074a <=( A167  and  (not A168) );
 a94075a <=( a94074a  and  a94071a );
 a94078a <=( (not A199)  and  (not A166) );
 a94081a <=( A201  and  A200 );
 a94082a <=( a94081a  and  a94078a );
 a94083a <=( a94082a  and  a94075a );
 a94086a <=( A265  and  A203 );
 a94089a <=( A267  and  (not A266) );
 a94090a <=( a94089a  and  a94086a );
 a94093a <=( A300  and  A268 );
 a94096a <=( (not A302)  and  (not A301) );
 a94097a <=( a94096a  and  a94093a );
 a94098a <=( a94097a  and  a94090a );
 a94101a <=( (not A169)  and  A170 );
 a94104a <=( A167  and  (not A168) );
 a94105a <=( a94104a  and  a94101a );
 a94108a <=( (not A199)  and  (not A166) );
 a94111a <=( A201  and  A200 );
 a94112a <=( a94111a  and  a94108a );
 a94113a <=( a94112a  and  a94105a );
 a94116a <=( A265  and  A203 );
 a94119a <=( A267  and  (not A266) );
 a94120a <=( a94119a  and  a94116a );
 a94123a <=( A300  and  A269 );
 a94126a <=( (not A302)  and  (not A301) );
 a94127a <=( a94126a  and  a94123a );
 a94128a <=( a94127a  and  a94120a );
 a94131a <=( (not A169)  and  A170 );
 a94134a <=( A167  and  (not A168) );
 a94135a <=( a94134a  and  a94131a );
 a94138a <=( (not A199)  and  (not A166) );
 a94141a <=( A201  and  A200 );
 a94142a <=( a94141a  and  a94138a );
 a94143a <=( a94142a  and  a94135a );
 a94146a <=( A265  and  A203 );
 a94149a <=( (not A267)  and  (not A266) );
 a94150a <=( a94149a  and  a94146a );
 a94153a <=( (not A269)  and  (not A268) );
 a94156a <=( A301  and  (not A300) );
 a94157a <=( a94156a  and  a94153a );
 a94158a <=( a94157a  and  a94150a );
 a94161a <=( (not A169)  and  A170 );
 a94164a <=( A167  and  (not A168) );
 a94165a <=( a94164a  and  a94161a );
 a94168a <=( (not A199)  and  (not A166) );
 a94171a <=( A201  and  A200 );
 a94172a <=( a94171a  and  a94168a );
 a94173a <=( a94172a  and  a94165a );
 a94176a <=( A265  and  A203 );
 a94179a <=( (not A267)  and  (not A266) );
 a94180a <=( a94179a  and  a94176a );
 a94183a <=( (not A269)  and  (not A268) );
 a94186a <=( A302  and  (not A300) );
 a94187a <=( a94186a  and  a94183a );
 a94188a <=( a94187a  and  a94180a );
 a94191a <=( (not A169)  and  A170 );
 a94194a <=( A167  and  (not A168) );
 a94195a <=( a94194a  and  a94191a );
 a94198a <=( (not A199)  and  (not A166) );
 a94201a <=( A201  and  A200 );
 a94202a <=( a94201a  and  a94198a );
 a94203a <=( a94202a  and  a94195a );
 a94206a <=( A265  and  A203 );
 a94209a <=( (not A267)  and  (not A266) );
 a94210a <=( a94209a  and  a94206a );
 a94213a <=( (not A269)  and  (not A268) );
 a94216a <=( A299  and  A298 );
 a94217a <=( a94216a  and  a94213a );
 a94218a <=( a94217a  and  a94210a );
 a94221a <=( (not A169)  and  A170 );
 a94224a <=( A167  and  (not A168) );
 a94225a <=( a94224a  and  a94221a );
 a94228a <=( (not A199)  and  (not A166) );
 a94231a <=( A201  and  A200 );
 a94232a <=( a94231a  and  a94228a );
 a94233a <=( a94232a  and  a94225a );
 a94236a <=( A265  and  A203 );
 a94239a <=( (not A267)  and  (not A266) );
 a94240a <=( a94239a  and  a94236a );
 a94243a <=( (not A269)  and  (not A268) );
 a94246a <=( (not A299)  and  (not A298) );
 a94247a <=( a94246a  and  a94243a );
 a94248a <=( a94247a  and  a94240a );
 a94251a <=( (not A169)  and  A170 );
 a94254a <=( A167  and  (not A168) );
 a94255a <=( a94254a  and  a94251a );
 a94258a <=( (not A199)  and  (not A166) );
 a94261a <=( (not A201)  and  A200 );
 a94262a <=( a94261a  and  a94258a );
 a94263a <=( a94262a  and  a94255a );
 a94266a <=( (not A203)  and  (not A202) );
 a94269a <=( A266  and  (not A265) );
 a94270a <=( a94269a  and  a94266a );
 a94273a <=( A268  and  A267 );
 a94276a <=( A301  and  (not A300) );
 a94277a <=( a94276a  and  a94273a );
 a94278a <=( a94277a  and  a94270a );
 a94281a <=( (not A169)  and  A170 );
 a94284a <=( A167  and  (not A168) );
 a94285a <=( a94284a  and  a94281a );
 a94288a <=( (not A199)  and  (not A166) );
 a94291a <=( (not A201)  and  A200 );
 a94292a <=( a94291a  and  a94288a );
 a94293a <=( a94292a  and  a94285a );
 a94296a <=( (not A203)  and  (not A202) );
 a94299a <=( A266  and  (not A265) );
 a94300a <=( a94299a  and  a94296a );
 a94303a <=( A268  and  A267 );
 a94306a <=( A302  and  (not A300) );
 a94307a <=( a94306a  and  a94303a );
 a94308a <=( a94307a  and  a94300a );
 a94311a <=( (not A169)  and  A170 );
 a94314a <=( A167  and  (not A168) );
 a94315a <=( a94314a  and  a94311a );
 a94318a <=( (not A199)  and  (not A166) );
 a94321a <=( (not A201)  and  A200 );
 a94322a <=( a94321a  and  a94318a );
 a94323a <=( a94322a  and  a94315a );
 a94326a <=( (not A203)  and  (not A202) );
 a94329a <=( A266  and  (not A265) );
 a94330a <=( a94329a  and  a94326a );
 a94333a <=( A268  and  A267 );
 a94336a <=( A299  and  A298 );
 a94337a <=( a94336a  and  a94333a );
 a94338a <=( a94337a  and  a94330a );
 a94341a <=( (not A169)  and  A170 );
 a94344a <=( A167  and  (not A168) );
 a94345a <=( a94344a  and  a94341a );
 a94348a <=( (not A199)  and  (not A166) );
 a94351a <=( (not A201)  and  A200 );
 a94352a <=( a94351a  and  a94348a );
 a94353a <=( a94352a  and  a94345a );
 a94356a <=( (not A203)  and  (not A202) );
 a94359a <=( A266  and  (not A265) );
 a94360a <=( a94359a  and  a94356a );
 a94363a <=( A268  and  A267 );
 a94366a <=( (not A299)  and  (not A298) );
 a94367a <=( a94366a  and  a94363a );
 a94368a <=( a94367a  and  a94360a );
 a94371a <=( (not A169)  and  A170 );
 a94374a <=( A167  and  (not A168) );
 a94375a <=( a94374a  and  a94371a );
 a94378a <=( (not A199)  and  (not A166) );
 a94381a <=( (not A201)  and  A200 );
 a94382a <=( a94381a  and  a94378a );
 a94383a <=( a94382a  and  a94375a );
 a94386a <=( (not A203)  and  (not A202) );
 a94389a <=( A266  and  (not A265) );
 a94390a <=( a94389a  and  a94386a );
 a94393a <=( A269  and  A267 );
 a94396a <=( A301  and  (not A300) );
 a94397a <=( a94396a  and  a94393a );
 a94398a <=( a94397a  and  a94390a );
 a94401a <=( (not A169)  and  A170 );
 a94404a <=( A167  and  (not A168) );
 a94405a <=( a94404a  and  a94401a );
 a94408a <=( (not A199)  and  (not A166) );
 a94411a <=( (not A201)  and  A200 );
 a94412a <=( a94411a  and  a94408a );
 a94413a <=( a94412a  and  a94405a );
 a94416a <=( (not A203)  and  (not A202) );
 a94419a <=( A266  and  (not A265) );
 a94420a <=( a94419a  and  a94416a );
 a94423a <=( A269  and  A267 );
 a94426a <=( A302  and  (not A300) );
 a94427a <=( a94426a  and  a94423a );
 a94428a <=( a94427a  and  a94420a );
 a94431a <=( (not A169)  and  A170 );
 a94434a <=( A167  and  (not A168) );
 a94435a <=( a94434a  and  a94431a );
 a94438a <=( (not A199)  and  (not A166) );
 a94441a <=( (not A201)  and  A200 );
 a94442a <=( a94441a  and  a94438a );
 a94443a <=( a94442a  and  a94435a );
 a94446a <=( (not A203)  and  (not A202) );
 a94449a <=( A266  and  (not A265) );
 a94450a <=( a94449a  and  a94446a );
 a94453a <=( A269  and  A267 );
 a94456a <=( A299  and  A298 );
 a94457a <=( a94456a  and  a94453a );
 a94458a <=( a94457a  and  a94450a );
 a94461a <=( (not A169)  and  A170 );
 a94464a <=( A167  and  (not A168) );
 a94465a <=( a94464a  and  a94461a );
 a94468a <=( (not A199)  and  (not A166) );
 a94471a <=( (not A201)  and  A200 );
 a94472a <=( a94471a  and  a94468a );
 a94473a <=( a94472a  and  a94465a );
 a94476a <=( (not A203)  and  (not A202) );
 a94479a <=( A266  and  (not A265) );
 a94480a <=( a94479a  and  a94476a );
 a94483a <=( A269  and  A267 );
 a94486a <=( (not A299)  and  (not A298) );
 a94487a <=( a94486a  and  a94483a );
 a94488a <=( a94487a  and  a94480a );
 a94491a <=( (not A169)  and  A170 );
 a94494a <=( A167  and  (not A168) );
 a94495a <=( a94494a  and  a94491a );
 a94498a <=( (not A199)  and  (not A166) );
 a94501a <=( (not A201)  and  A200 );
 a94502a <=( a94501a  and  a94498a );
 a94503a <=( a94502a  and  a94495a );
 a94506a <=( (not A203)  and  (not A202) );
 a94509a <=( (not A266)  and  A265 );
 a94510a <=( a94509a  and  a94506a );
 a94513a <=( A268  and  A267 );
 a94516a <=( A301  and  (not A300) );
 a94517a <=( a94516a  and  a94513a );
 a94518a <=( a94517a  and  a94510a );
 a94521a <=( (not A169)  and  A170 );
 a94524a <=( A167  and  (not A168) );
 a94525a <=( a94524a  and  a94521a );
 a94528a <=( (not A199)  and  (not A166) );
 a94531a <=( (not A201)  and  A200 );
 a94532a <=( a94531a  and  a94528a );
 a94533a <=( a94532a  and  a94525a );
 a94536a <=( (not A203)  and  (not A202) );
 a94539a <=( (not A266)  and  A265 );
 a94540a <=( a94539a  and  a94536a );
 a94543a <=( A268  and  A267 );
 a94546a <=( A302  and  (not A300) );
 a94547a <=( a94546a  and  a94543a );
 a94548a <=( a94547a  and  a94540a );
 a94551a <=( (not A169)  and  A170 );
 a94554a <=( A167  and  (not A168) );
 a94555a <=( a94554a  and  a94551a );
 a94558a <=( (not A199)  and  (not A166) );
 a94561a <=( (not A201)  and  A200 );
 a94562a <=( a94561a  and  a94558a );
 a94563a <=( a94562a  and  a94555a );
 a94566a <=( (not A203)  and  (not A202) );
 a94569a <=( (not A266)  and  A265 );
 a94570a <=( a94569a  and  a94566a );
 a94573a <=( A268  and  A267 );
 a94576a <=( A299  and  A298 );
 a94577a <=( a94576a  and  a94573a );
 a94578a <=( a94577a  and  a94570a );
 a94581a <=( (not A169)  and  A170 );
 a94584a <=( A167  and  (not A168) );
 a94585a <=( a94584a  and  a94581a );
 a94588a <=( (not A199)  and  (not A166) );
 a94591a <=( (not A201)  and  A200 );
 a94592a <=( a94591a  and  a94588a );
 a94593a <=( a94592a  and  a94585a );
 a94596a <=( (not A203)  and  (not A202) );
 a94599a <=( (not A266)  and  A265 );
 a94600a <=( a94599a  and  a94596a );
 a94603a <=( A268  and  A267 );
 a94606a <=( (not A299)  and  (not A298) );
 a94607a <=( a94606a  and  a94603a );
 a94608a <=( a94607a  and  a94600a );
 a94611a <=( (not A169)  and  A170 );
 a94614a <=( A167  and  (not A168) );
 a94615a <=( a94614a  and  a94611a );
 a94618a <=( (not A199)  and  (not A166) );
 a94621a <=( (not A201)  and  A200 );
 a94622a <=( a94621a  and  a94618a );
 a94623a <=( a94622a  and  a94615a );
 a94626a <=( (not A203)  and  (not A202) );
 a94629a <=( (not A266)  and  A265 );
 a94630a <=( a94629a  and  a94626a );
 a94633a <=( A269  and  A267 );
 a94636a <=( A301  and  (not A300) );
 a94637a <=( a94636a  and  a94633a );
 a94638a <=( a94637a  and  a94630a );
 a94641a <=( (not A169)  and  A170 );
 a94644a <=( A167  and  (not A168) );
 a94645a <=( a94644a  and  a94641a );
 a94648a <=( (not A199)  and  (not A166) );
 a94651a <=( (not A201)  and  A200 );
 a94652a <=( a94651a  and  a94648a );
 a94653a <=( a94652a  and  a94645a );
 a94656a <=( (not A203)  and  (not A202) );
 a94659a <=( (not A266)  and  A265 );
 a94660a <=( a94659a  and  a94656a );
 a94663a <=( A269  and  A267 );
 a94666a <=( A302  and  (not A300) );
 a94667a <=( a94666a  and  a94663a );
 a94668a <=( a94667a  and  a94660a );
 a94671a <=( (not A169)  and  A170 );
 a94674a <=( A167  and  (not A168) );
 a94675a <=( a94674a  and  a94671a );
 a94678a <=( (not A199)  and  (not A166) );
 a94681a <=( (not A201)  and  A200 );
 a94682a <=( a94681a  and  a94678a );
 a94683a <=( a94682a  and  a94675a );
 a94686a <=( (not A203)  and  (not A202) );
 a94689a <=( (not A266)  and  A265 );
 a94690a <=( a94689a  and  a94686a );
 a94693a <=( A269  and  A267 );
 a94696a <=( A299  and  A298 );
 a94697a <=( a94696a  and  a94693a );
 a94698a <=( a94697a  and  a94690a );
 a94701a <=( (not A169)  and  A170 );
 a94704a <=( A167  and  (not A168) );
 a94705a <=( a94704a  and  a94701a );
 a94708a <=( (not A199)  and  (not A166) );
 a94711a <=( (not A201)  and  A200 );
 a94712a <=( a94711a  and  a94708a );
 a94713a <=( a94712a  and  a94705a );
 a94716a <=( (not A203)  and  (not A202) );
 a94719a <=( (not A266)  and  A265 );
 a94720a <=( a94719a  and  a94716a );
 a94723a <=( A269  and  A267 );
 a94726a <=( (not A299)  and  (not A298) );
 a94727a <=( a94726a  and  a94723a );
 a94728a <=( a94727a  and  a94720a );
 a94731a <=( (not A169)  and  A170 );
 a94734a <=( A167  and  (not A168) );
 a94735a <=( a94734a  and  a94731a );
 a94738a <=( A199  and  (not A166) );
 a94741a <=( A201  and  (not A200) );
 a94742a <=( a94741a  and  a94738a );
 a94743a <=( a94742a  and  a94735a );
 a94746a <=( (not A265)  and  A202 );
 a94749a <=( A267  and  A266 );
 a94750a <=( a94749a  and  a94746a );
 a94753a <=( A300  and  A268 );
 a94756a <=( (not A302)  and  (not A301) );
 a94757a <=( a94756a  and  a94753a );
 a94758a <=( a94757a  and  a94750a );
 a94761a <=( (not A169)  and  A170 );
 a94764a <=( A167  and  (not A168) );
 a94765a <=( a94764a  and  a94761a );
 a94768a <=( A199  and  (not A166) );
 a94771a <=( A201  and  (not A200) );
 a94772a <=( a94771a  and  a94768a );
 a94773a <=( a94772a  and  a94765a );
 a94776a <=( (not A265)  and  A202 );
 a94779a <=( A267  and  A266 );
 a94780a <=( a94779a  and  a94776a );
 a94783a <=( A300  and  A269 );
 a94786a <=( (not A302)  and  (not A301) );
 a94787a <=( a94786a  and  a94783a );
 a94788a <=( a94787a  and  a94780a );
 a94791a <=( (not A169)  and  A170 );
 a94794a <=( A167  and  (not A168) );
 a94795a <=( a94794a  and  a94791a );
 a94798a <=( A199  and  (not A166) );
 a94801a <=( A201  and  (not A200) );
 a94802a <=( a94801a  and  a94798a );
 a94803a <=( a94802a  and  a94795a );
 a94806a <=( (not A265)  and  A202 );
 a94809a <=( (not A267)  and  A266 );
 a94810a <=( a94809a  and  a94806a );
 a94813a <=( (not A269)  and  (not A268) );
 a94816a <=( A301  and  (not A300) );
 a94817a <=( a94816a  and  a94813a );
 a94818a <=( a94817a  and  a94810a );
 a94821a <=( (not A169)  and  A170 );
 a94824a <=( A167  and  (not A168) );
 a94825a <=( a94824a  and  a94821a );
 a94828a <=( A199  and  (not A166) );
 a94831a <=( A201  and  (not A200) );
 a94832a <=( a94831a  and  a94828a );
 a94833a <=( a94832a  and  a94825a );
 a94836a <=( (not A265)  and  A202 );
 a94839a <=( (not A267)  and  A266 );
 a94840a <=( a94839a  and  a94836a );
 a94843a <=( (not A269)  and  (not A268) );
 a94846a <=( A302  and  (not A300) );
 a94847a <=( a94846a  and  a94843a );
 a94848a <=( a94847a  and  a94840a );
 a94851a <=( (not A169)  and  A170 );
 a94854a <=( A167  and  (not A168) );
 a94855a <=( a94854a  and  a94851a );
 a94858a <=( A199  and  (not A166) );
 a94861a <=( A201  and  (not A200) );
 a94862a <=( a94861a  and  a94858a );
 a94863a <=( a94862a  and  a94855a );
 a94866a <=( (not A265)  and  A202 );
 a94869a <=( (not A267)  and  A266 );
 a94870a <=( a94869a  and  a94866a );
 a94873a <=( (not A269)  and  (not A268) );
 a94876a <=( A299  and  A298 );
 a94877a <=( a94876a  and  a94873a );
 a94878a <=( a94877a  and  a94870a );
 a94881a <=( (not A169)  and  A170 );
 a94884a <=( A167  and  (not A168) );
 a94885a <=( a94884a  and  a94881a );
 a94888a <=( A199  and  (not A166) );
 a94891a <=( A201  and  (not A200) );
 a94892a <=( a94891a  and  a94888a );
 a94893a <=( a94892a  and  a94885a );
 a94896a <=( (not A265)  and  A202 );
 a94899a <=( (not A267)  and  A266 );
 a94900a <=( a94899a  and  a94896a );
 a94903a <=( (not A269)  and  (not A268) );
 a94906a <=( (not A299)  and  (not A298) );
 a94907a <=( a94906a  and  a94903a );
 a94908a <=( a94907a  and  a94900a );
 a94911a <=( (not A169)  and  A170 );
 a94914a <=( A167  and  (not A168) );
 a94915a <=( a94914a  and  a94911a );
 a94918a <=( A199  and  (not A166) );
 a94921a <=( A201  and  (not A200) );
 a94922a <=( a94921a  and  a94918a );
 a94923a <=( a94922a  and  a94915a );
 a94926a <=( A265  and  A202 );
 a94929a <=( A267  and  (not A266) );
 a94930a <=( a94929a  and  a94926a );
 a94933a <=( A300  and  A268 );
 a94936a <=( (not A302)  and  (not A301) );
 a94937a <=( a94936a  and  a94933a );
 a94938a <=( a94937a  and  a94930a );
 a94941a <=( (not A169)  and  A170 );
 a94944a <=( A167  and  (not A168) );
 a94945a <=( a94944a  and  a94941a );
 a94948a <=( A199  and  (not A166) );
 a94951a <=( A201  and  (not A200) );
 a94952a <=( a94951a  and  a94948a );
 a94953a <=( a94952a  and  a94945a );
 a94956a <=( A265  and  A202 );
 a94959a <=( A267  and  (not A266) );
 a94960a <=( a94959a  and  a94956a );
 a94963a <=( A300  and  A269 );
 a94966a <=( (not A302)  and  (not A301) );
 a94967a <=( a94966a  and  a94963a );
 a94968a <=( a94967a  and  a94960a );
 a94971a <=( (not A169)  and  A170 );
 a94974a <=( A167  and  (not A168) );
 a94975a <=( a94974a  and  a94971a );
 a94978a <=( A199  and  (not A166) );
 a94981a <=( A201  and  (not A200) );
 a94982a <=( a94981a  and  a94978a );
 a94983a <=( a94982a  and  a94975a );
 a94986a <=( A265  and  A202 );
 a94989a <=( (not A267)  and  (not A266) );
 a94990a <=( a94989a  and  a94986a );
 a94993a <=( (not A269)  and  (not A268) );
 a94996a <=( A301  and  (not A300) );
 a94997a <=( a94996a  and  a94993a );
 a94998a <=( a94997a  and  a94990a );
 a95001a <=( (not A169)  and  A170 );
 a95004a <=( A167  and  (not A168) );
 a95005a <=( a95004a  and  a95001a );
 a95008a <=( A199  and  (not A166) );
 a95011a <=( A201  and  (not A200) );
 a95012a <=( a95011a  and  a95008a );
 a95013a <=( a95012a  and  a95005a );
 a95016a <=( A265  and  A202 );
 a95019a <=( (not A267)  and  (not A266) );
 a95020a <=( a95019a  and  a95016a );
 a95023a <=( (not A269)  and  (not A268) );
 a95026a <=( A302  and  (not A300) );
 a95027a <=( a95026a  and  a95023a );
 a95028a <=( a95027a  and  a95020a );
 a95031a <=( (not A169)  and  A170 );
 a95034a <=( A167  and  (not A168) );
 a95035a <=( a95034a  and  a95031a );
 a95038a <=( A199  and  (not A166) );
 a95041a <=( A201  and  (not A200) );
 a95042a <=( a95041a  and  a95038a );
 a95043a <=( a95042a  and  a95035a );
 a95046a <=( A265  and  A202 );
 a95049a <=( (not A267)  and  (not A266) );
 a95050a <=( a95049a  and  a95046a );
 a95053a <=( (not A269)  and  (not A268) );
 a95056a <=( A299  and  A298 );
 a95057a <=( a95056a  and  a95053a );
 a95058a <=( a95057a  and  a95050a );
 a95061a <=( (not A169)  and  A170 );
 a95064a <=( A167  and  (not A168) );
 a95065a <=( a95064a  and  a95061a );
 a95068a <=( A199  and  (not A166) );
 a95071a <=( A201  and  (not A200) );
 a95072a <=( a95071a  and  a95068a );
 a95073a <=( a95072a  and  a95065a );
 a95076a <=( A265  and  A202 );
 a95079a <=( (not A267)  and  (not A266) );
 a95080a <=( a95079a  and  a95076a );
 a95083a <=( (not A269)  and  (not A268) );
 a95086a <=( (not A299)  and  (not A298) );
 a95087a <=( a95086a  and  a95083a );
 a95088a <=( a95087a  and  a95080a );
 a95091a <=( (not A169)  and  A170 );
 a95094a <=( A167  and  (not A168) );
 a95095a <=( a95094a  and  a95091a );
 a95098a <=( A199  and  (not A166) );
 a95101a <=( A201  and  (not A200) );
 a95102a <=( a95101a  and  a95098a );
 a95103a <=( a95102a  and  a95095a );
 a95106a <=( (not A265)  and  A203 );
 a95109a <=( A267  and  A266 );
 a95110a <=( a95109a  and  a95106a );
 a95113a <=( A300  and  A268 );
 a95116a <=( (not A302)  and  (not A301) );
 a95117a <=( a95116a  and  a95113a );
 a95118a <=( a95117a  and  a95110a );
 a95121a <=( (not A169)  and  A170 );
 a95124a <=( A167  and  (not A168) );
 a95125a <=( a95124a  and  a95121a );
 a95128a <=( A199  and  (not A166) );
 a95131a <=( A201  and  (not A200) );
 a95132a <=( a95131a  and  a95128a );
 a95133a <=( a95132a  and  a95125a );
 a95136a <=( (not A265)  and  A203 );
 a95139a <=( A267  and  A266 );
 a95140a <=( a95139a  and  a95136a );
 a95143a <=( A300  and  A269 );
 a95146a <=( (not A302)  and  (not A301) );
 a95147a <=( a95146a  and  a95143a );
 a95148a <=( a95147a  and  a95140a );
 a95151a <=( (not A169)  and  A170 );
 a95154a <=( A167  and  (not A168) );
 a95155a <=( a95154a  and  a95151a );
 a95158a <=( A199  and  (not A166) );
 a95161a <=( A201  and  (not A200) );
 a95162a <=( a95161a  and  a95158a );
 a95163a <=( a95162a  and  a95155a );
 a95166a <=( (not A265)  and  A203 );
 a95169a <=( (not A267)  and  A266 );
 a95170a <=( a95169a  and  a95166a );
 a95173a <=( (not A269)  and  (not A268) );
 a95176a <=( A301  and  (not A300) );
 a95177a <=( a95176a  and  a95173a );
 a95178a <=( a95177a  and  a95170a );
 a95181a <=( (not A169)  and  A170 );
 a95184a <=( A167  and  (not A168) );
 a95185a <=( a95184a  and  a95181a );
 a95188a <=( A199  and  (not A166) );
 a95191a <=( A201  and  (not A200) );
 a95192a <=( a95191a  and  a95188a );
 a95193a <=( a95192a  and  a95185a );
 a95196a <=( (not A265)  and  A203 );
 a95199a <=( (not A267)  and  A266 );
 a95200a <=( a95199a  and  a95196a );
 a95203a <=( (not A269)  and  (not A268) );
 a95206a <=( A302  and  (not A300) );
 a95207a <=( a95206a  and  a95203a );
 a95208a <=( a95207a  and  a95200a );
 a95211a <=( (not A169)  and  A170 );
 a95214a <=( A167  and  (not A168) );
 a95215a <=( a95214a  and  a95211a );
 a95218a <=( A199  and  (not A166) );
 a95221a <=( A201  and  (not A200) );
 a95222a <=( a95221a  and  a95218a );
 a95223a <=( a95222a  and  a95215a );
 a95226a <=( (not A265)  and  A203 );
 a95229a <=( (not A267)  and  A266 );
 a95230a <=( a95229a  and  a95226a );
 a95233a <=( (not A269)  and  (not A268) );
 a95236a <=( A299  and  A298 );
 a95237a <=( a95236a  and  a95233a );
 a95238a <=( a95237a  and  a95230a );
 a95241a <=( (not A169)  and  A170 );
 a95244a <=( A167  and  (not A168) );
 a95245a <=( a95244a  and  a95241a );
 a95248a <=( A199  and  (not A166) );
 a95251a <=( A201  and  (not A200) );
 a95252a <=( a95251a  and  a95248a );
 a95253a <=( a95252a  and  a95245a );
 a95256a <=( (not A265)  and  A203 );
 a95259a <=( (not A267)  and  A266 );
 a95260a <=( a95259a  and  a95256a );
 a95263a <=( (not A269)  and  (not A268) );
 a95266a <=( (not A299)  and  (not A298) );
 a95267a <=( a95266a  and  a95263a );
 a95268a <=( a95267a  and  a95260a );
 a95271a <=( (not A169)  and  A170 );
 a95274a <=( A167  and  (not A168) );
 a95275a <=( a95274a  and  a95271a );
 a95278a <=( A199  and  (not A166) );
 a95281a <=( A201  and  (not A200) );
 a95282a <=( a95281a  and  a95278a );
 a95283a <=( a95282a  and  a95275a );
 a95286a <=( A265  and  A203 );
 a95289a <=( A267  and  (not A266) );
 a95290a <=( a95289a  and  a95286a );
 a95293a <=( A300  and  A268 );
 a95296a <=( (not A302)  and  (not A301) );
 a95297a <=( a95296a  and  a95293a );
 a95298a <=( a95297a  and  a95290a );
 a95301a <=( (not A169)  and  A170 );
 a95304a <=( A167  and  (not A168) );
 a95305a <=( a95304a  and  a95301a );
 a95308a <=( A199  and  (not A166) );
 a95311a <=( A201  and  (not A200) );
 a95312a <=( a95311a  and  a95308a );
 a95313a <=( a95312a  and  a95305a );
 a95316a <=( A265  and  A203 );
 a95319a <=( A267  and  (not A266) );
 a95320a <=( a95319a  and  a95316a );
 a95323a <=( A300  and  A269 );
 a95326a <=( (not A302)  and  (not A301) );
 a95327a <=( a95326a  and  a95323a );
 a95328a <=( a95327a  and  a95320a );
 a95331a <=( (not A169)  and  A170 );
 a95334a <=( A167  and  (not A168) );
 a95335a <=( a95334a  and  a95331a );
 a95338a <=( A199  and  (not A166) );
 a95341a <=( A201  and  (not A200) );
 a95342a <=( a95341a  and  a95338a );
 a95343a <=( a95342a  and  a95335a );
 a95346a <=( A265  and  A203 );
 a95349a <=( (not A267)  and  (not A266) );
 a95350a <=( a95349a  and  a95346a );
 a95353a <=( (not A269)  and  (not A268) );
 a95356a <=( A301  and  (not A300) );
 a95357a <=( a95356a  and  a95353a );
 a95358a <=( a95357a  and  a95350a );
 a95361a <=( (not A169)  and  A170 );
 a95364a <=( A167  and  (not A168) );
 a95365a <=( a95364a  and  a95361a );
 a95368a <=( A199  and  (not A166) );
 a95371a <=( A201  and  (not A200) );
 a95372a <=( a95371a  and  a95368a );
 a95373a <=( a95372a  and  a95365a );
 a95376a <=( A265  and  A203 );
 a95379a <=( (not A267)  and  (not A266) );
 a95380a <=( a95379a  and  a95376a );
 a95383a <=( (not A269)  and  (not A268) );
 a95386a <=( A302  and  (not A300) );
 a95387a <=( a95386a  and  a95383a );
 a95388a <=( a95387a  and  a95380a );
 a95391a <=( (not A169)  and  A170 );
 a95394a <=( A167  and  (not A168) );
 a95395a <=( a95394a  and  a95391a );
 a95398a <=( A199  and  (not A166) );
 a95401a <=( A201  and  (not A200) );
 a95402a <=( a95401a  and  a95398a );
 a95403a <=( a95402a  and  a95395a );
 a95406a <=( A265  and  A203 );
 a95409a <=( (not A267)  and  (not A266) );
 a95410a <=( a95409a  and  a95406a );
 a95413a <=( (not A269)  and  (not A268) );
 a95416a <=( A299  and  A298 );
 a95417a <=( a95416a  and  a95413a );
 a95418a <=( a95417a  and  a95410a );
 a95421a <=( (not A169)  and  A170 );
 a95424a <=( A167  and  (not A168) );
 a95425a <=( a95424a  and  a95421a );
 a95428a <=( A199  and  (not A166) );
 a95431a <=( A201  and  (not A200) );
 a95432a <=( a95431a  and  a95428a );
 a95433a <=( a95432a  and  a95425a );
 a95436a <=( A265  and  A203 );
 a95439a <=( (not A267)  and  (not A266) );
 a95440a <=( a95439a  and  a95436a );
 a95443a <=( (not A269)  and  (not A268) );
 a95446a <=( (not A299)  and  (not A298) );
 a95447a <=( a95446a  and  a95443a );
 a95448a <=( a95447a  and  a95440a );
 a95451a <=( (not A169)  and  A170 );
 a95454a <=( A167  and  (not A168) );
 a95455a <=( a95454a  and  a95451a );
 a95458a <=( A199  and  (not A166) );
 a95461a <=( (not A201)  and  (not A200) );
 a95462a <=( a95461a  and  a95458a );
 a95463a <=( a95462a  and  a95455a );
 a95466a <=( (not A203)  and  (not A202) );
 a95469a <=( A266  and  (not A265) );
 a95470a <=( a95469a  and  a95466a );
 a95473a <=( A268  and  A267 );
 a95476a <=( A301  and  (not A300) );
 a95477a <=( a95476a  and  a95473a );
 a95478a <=( a95477a  and  a95470a );
 a95481a <=( (not A169)  and  A170 );
 a95484a <=( A167  and  (not A168) );
 a95485a <=( a95484a  and  a95481a );
 a95488a <=( A199  and  (not A166) );
 a95491a <=( (not A201)  and  (not A200) );
 a95492a <=( a95491a  and  a95488a );
 a95493a <=( a95492a  and  a95485a );
 a95496a <=( (not A203)  and  (not A202) );
 a95499a <=( A266  and  (not A265) );
 a95500a <=( a95499a  and  a95496a );
 a95503a <=( A268  and  A267 );
 a95506a <=( A302  and  (not A300) );
 a95507a <=( a95506a  and  a95503a );
 a95508a <=( a95507a  and  a95500a );
 a95511a <=( (not A169)  and  A170 );
 a95514a <=( A167  and  (not A168) );
 a95515a <=( a95514a  and  a95511a );
 a95518a <=( A199  and  (not A166) );
 a95521a <=( (not A201)  and  (not A200) );
 a95522a <=( a95521a  and  a95518a );
 a95523a <=( a95522a  and  a95515a );
 a95526a <=( (not A203)  and  (not A202) );
 a95529a <=( A266  and  (not A265) );
 a95530a <=( a95529a  and  a95526a );
 a95533a <=( A268  and  A267 );
 a95536a <=( A299  and  A298 );
 a95537a <=( a95536a  and  a95533a );
 a95538a <=( a95537a  and  a95530a );
 a95541a <=( (not A169)  and  A170 );
 a95544a <=( A167  and  (not A168) );
 a95545a <=( a95544a  and  a95541a );
 a95548a <=( A199  and  (not A166) );
 a95551a <=( (not A201)  and  (not A200) );
 a95552a <=( a95551a  and  a95548a );
 a95553a <=( a95552a  and  a95545a );
 a95556a <=( (not A203)  and  (not A202) );
 a95559a <=( A266  and  (not A265) );
 a95560a <=( a95559a  and  a95556a );
 a95563a <=( A268  and  A267 );
 a95566a <=( (not A299)  and  (not A298) );
 a95567a <=( a95566a  and  a95563a );
 a95568a <=( a95567a  and  a95560a );
 a95571a <=( (not A169)  and  A170 );
 a95574a <=( A167  and  (not A168) );
 a95575a <=( a95574a  and  a95571a );
 a95578a <=( A199  and  (not A166) );
 a95581a <=( (not A201)  and  (not A200) );
 a95582a <=( a95581a  and  a95578a );
 a95583a <=( a95582a  and  a95575a );
 a95586a <=( (not A203)  and  (not A202) );
 a95589a <=( A266  and  (not A265) );
 a95590a <=( a95589a  and  a95586a );
 a95593a <=( A269  and  A267 );
 a95596a <=( A301  and  (not A300) );
 a95597a <=( a95596a  and  a95593a );
 a95598a <=( a95597a  and  a95590a );
 a95601a <=( (not A169)  and  A170 );
 a95604a <=( A167  and  (not A168) );
 a95605a <=( a95604a  and  a95601a );
 a95608a <=( A199  and  (not A166) );
 a95611a <=( (not A201)  and  (not A200) );
 a95612a <=( a95611a  and  a95608a );
 a95613a <=( a95612a  and  a95605a );
 a95616a <=( (not A203)  and  (not A202) );
 a95619a <=( A266  and  (not A265) );
 a95620a <=( a95619a  and  a95616a );
 a95623a <=( A269  and  A267 );
 a95626a <=( A302  and  (not A300) );
 a95627a <=( a95626a  and  a95623a );
 a95628a <=( a95627a  and  a95620a );
 a95631a <=( (not A169)  and  A170 );
 a95634a <=( A167  and  (not A168) );
 a95635a <=( a95634a  and  a95631a );
 a95638a <=( A199  and  (not A166) );
 a95641a <=( (not A201)  and  (not A200) );
 a95642a <=( a95641a  and  a95638a );
 a95643a <=( a95642a  and  a95635a );
 a95646a <=( (not A203)  and  (not A202) );
 a95649a <=( A266  and  (not A265) );
 a95650a <=( a95649a  and  a95646a );
 a95653a <=( A269  and  A267 );
 a95656a <=( A299  and  A298 );
 a95657a <=( a95656a  and  a95653a );
 a95658a <=( a95657a  and  a95650a );
 a95661a <=( (not A169)  and  A170 );
 a95664a <=( A167  and  (not A168) );
 a95665a <=( a95664a  and  a95661a );
 a95668a <=( A199  and  (not A166) );
 a95671a <=( (not A201)  and  (not A200) );
 a95672a <=( a95671a  and  a95668a );
 a95673a <=( a95672a  and  a95665a );
 a95676a <=( (not A203)  and  (not A202) );
 a95679a <=( A266  and  (not A265) );
 a95680a <=( a95679a  and  a95676a );
 a95683a <=( A269  and  A267 );
 a95686a <=( (not A299)  and  (not A298) );
 a95687a <=( a95686a  and  a95683a );
 a95688a <=( a95687a  and  a95680a );
 a95691a <=( (not A169)  and  A170 );
 a95694a <=( A167  and  (not A168) );
 a95695a <=( a95694a  and  a95691a );
 a95698a <=( A199  and  (not A166) );
 a95701a <=( (not A201)  and  (not A200) );
 a95702a <=( a95701a  and  a95698a );
 a95703a <=( a95702a  and  a95695a );
 a95706a <=( (not A203)  and  (not A202) );
 a95709a <=( (not A266)  and  A265 );
 a95710a <=( a95709a  and  a95706a );
 a95713a <=( A268  and  A267 );
 a95716a <=( A301  and  (not A300) );
 a95717a <=( a95716a  and  a95713a );
 a95718a <=( a95717a  and  a95710a );
 a95721a <=( (not A169)  and  A170 );
 a95724a <=( A167  and  (not A168) );
 a95725a <=( a95724a  and  a95721a );
 a95728a <=( A199  and  (not A166) );
 a95731a <=( (not A201)  and  (not A200) );
 a95732a <=( a95731a  and  a95728a );
 a95733a <=( a95732a  and  a95725a );
 a95736a <=( (not A203)  and  (not A202) );
 a95739a <=( (not A266)  and  A265 );
 a95740a <=( a95739a  and  a95736a );
 a95743a <=( A268  and  A267 );
 a95746a <=( A302  and  (not A300) );
 a95747a <=( a95746a  and  a95743a );
 a95748a <=( a95747a  and  a95740a );
 a95751a <=( (not A169)  and  A170 );
 a95754a <=( A167  and  (not A168) );
 a95755a <=( a95754a  and  a95751a );
 a95758a <=( A199  and  (not A166) );
 a95761a <=( (not A201)  and  (not A200) );
 a95762a <=( a95761a  and  a95758a );
 a95763a <=( a95762a  and  a95755a );
 a95766a <=( (not A203)  and  (not A202) );
 a95769a <=( (not A266)  and  A265 );
 a95770a <=( a95769a  and  a95766a );
 a95773a <=( A268  and  A267 );
 a95776a <=( A299  and  A298 );
 a95777a <=( a95776a  and  a95773a );
 a95778a <=( a95777a  and  a95770a );
 a95781a <=( (not A169)  and  A170 );
 a95784a <=( A167  and  (not A168) );
 a95785a <=( a95784a  and  a95781a );
 a95788a <=( A199  and  (not A166) );
 a95791a <=( (not A201)  and  (not A200) );
 a95792a <=( a95791a  and  a95788a );
 a95793a <=( a95792a  and  a95785a );
 a95796a <=( (not A203)  and  (not A202) );
 a95799a <=( (not A266)  and  A265 );
 a95800a <=( a95799a  and  a95796a );
 a95803a <=( A268  and  A267 );
 a95806a <=( (not A299)  and  (not A298) );
 a95807a <=( a95806a  and  a95803a );
 a95808a <=( a95807a  and  a95800a );
 a95811a <=( (not A169)  and  A170 );
 a95814a <=( A167  and  (not A168) );
 a95815a <=( a95814a  and  a95811a );
 a95818a <=( A199  and  (not A166) );
 a95821a <=( (not A201)  and  (not A200) );
 a95822a <=( a95821a  and  a95818a );
 a95823a <=( a95822a  and  a95815a );
 a95826a <=( (not A203)  and  (not A202) );
 a95829a <=( (not A266)  and  A265 );
 a95830a <=( a95829a  and  a95826a );
 a95833a <=( A269  and  A267 );
 a95836a <=( A301  and  (not A300) );
 a95837a <=( a95836a  and  a95833a );
 a95838a <=( a95837a  and  a95830a );
 a95841a <=( (not A169)  and  A170 );
 a95844a <=( A167  and  (not A168) );
 a95845a <=( a95844a  and  a95841a );
 a95848a <=( A199  and  (not A166) );
 a95851a <=( (not A201)  and  (not A200) );
 a95852a <=( a95851a  and  a95848a );
 a95853a <=( a95852a  and  a95845a );
 a95856a <=( (not A203)  and  (not A202) );
 a95859a <=( (not A266)  and  A265 );
 a95860a <=( a95859a  and  a95856a );
 a95863a <=( A269  and  A267 );
 a95866a <=( A302  and  (not A300) );
 a95867a <=( a95866a  and  a95863a );
 a95868a <=( a95867a  and  a95860a );
 a95871a <=( (not A169)  and  A170 );
 a95874a <=( A167  and  (not A168) );
 a95875a <=( a95874a  and  a95871a );
 a95878a <=( A199  and  (not A166) );
 a95881a <=( (not A201)  and  (not A200) );
 a95882a <=( a95881a  and  a95878a );
 a95883a <=( a95882a  and  a95875a );
 a95886a <=( (not A203)  and  (not A202) );
 a95889a <=( (not A266)  and  A265 );
 a95890a <=( a95889a  and  a95886a );
 a95893a <=( A269  and  A267 );
 a95896a <=( A299  and  A298 );
 a95897a <=( a95896a  and  a95893a );
 a95898a <=( a95897a  and  a95890a );
 a95901a <=( (not A169)  and  A170 );
 a95904a <=( A167  and  (not A168) );
 a95905a <=( a95904a  and  a95901a );
 a95908a <=( A199  and  (not A166) );
 a95911a <=( (not A201)  and  (not A200) );
 a95912a <=( a95911a  and  a95908a );
 a95913a <=( a95912a  and  a95905a );
 a95916a <=( (not A203)  and  (not A202) );
 a95919a <=( (not A266)  and  A265 );
 a95920a <=( a95919a  and  a95916a );
 a95923a <=( A269  and  A267 );
 a95926a <=( (not A299)  and  (not A298) );
 a95927a <=( a95926a  and  a95923a );
 a95928a <=( a95927a  and  a95920a );
 a95931a <=( (not A169)  and  A170 );
 a95934a <=( (not A167)  and  (not A168) );
 a95935a <=( a95934a  and  a95931a );
 a95938a <=( A201  and  A166 );
 a95941a <=( (not A203)  and  (not A202) );
 a95942a <=( a95941a  and  a95938a );
 a95943a <=( a95942a  and  a95935a );
 a95946a <=( (not A268)  and  A267 );
 a95949a <=( A298  and  (not A269) );
 a95950a <=( a95949a  and  a95946a );
 a95953a <=( (not A300)  and  (not A299) );
 a95956a <=( (not A302)  and  (not A301) );
 a95957a <=( a95956a  and  a95953a );
 a95958a <=( a95957a  and  a95950a );
 a95961a <=( (not A169)  and  A170 );
 a95964a <=( (not A167)  and  (not A168) );
 a95965a <=( a95964a  and  a95961a );
 a95968a <=( A201  and  A166 );
 a95971a <=( (not A203)  and  (not A202) );
 a95972a <=( a95971a  and  a95968a );
 a95973a <=( a95972a  and  a95965a );
 a95976a <=( (not A268)  and  A267 );
 a95979a <=( (not A298)  and  (not A269) );
 a95980a <=( a95979a  and  a95976a );
 a95983a <=( (not A300)  and  A299 );
 a95986a <=( (not A302)  and  (not A301) );
 a95987a <=( a95986a  and  a95983a );
 a95988a <=( a95987a  and  a95980a );
 a95991a <=( (not A169)  and  A170 );
 a95994a <=( (not A167)  and  (not A168) );
 a95995a <=( a95994a  and  a95991a );
 a95998a <=( (not A199)  and  A166 );
 a96001a <=( A201  and  A200 );
 a96002a <=( a96001a  and  a95998a );
 a96003a <=( a96002a  and  a95995a );
 a96006a <=( (not A265)  and  A202 );
 a96009a <=( A267  and  A266 );
 a96010a <=( a96009a  and  a96006a );
 a96013a <=( A300  and  A268 );
 a96016a <=( (not A302)  and  (not A301) );
 a96017a <=( a96016a  and  a96013a );
 a96018a <=( a96017a  and  a96010a );
 a96021a <=( (not A169)  and  A170 );
 a96024a <=( (not A167)  and  (not A168) );
 a96025a <=( a96024a  and  a96021a );
 a96028a <=( (not A199)  and  A166 );
 a96031a <=( A201  and  A200 );
 a96032a <=( a96031a  and  a96028a );
 a96033a <=( a96032a  and  a96025a );
 a96036a <=( (not A265)  and  A202 );
 a96039a <=( A267  and  A266 );
 a96040a <=( a96039a  and  a96036a );
 a96043a <=( A300  and  A269 );
 a96046a <=( (not A302)  and  (not A301) );
 a96047a <=( a96046a  and  a96043a );
 a96048a <=( a96047a  and  a96040a );
 a96051a <=( (not A169)  and  A170 );
 a96054a <=( (not A167)  and  (not A168) );
 a96055a <=( a96054a  and  a96051a );
 a96058a <=( (not A199)  and  A166 );
 a96061a <=( A201  and  A200 );
 a96062a <=( a96061a  and  a96058a );
 a96063a <=( a96062a  and  a96055a );
 a96066a <=( (not A265)  and  A202 );
 a96069a <=( (not A267)  and  A266 );
 a96070a <=( a96069a  and  a96066a );
 a96073a <=( (not A269)  and  (not A268) );
 a96076a <=( A301  and  (not A300) );
 a96077a <=( a96076a  and  a96073a );
 a96078a <=( a96077a  and  a96070a );
 a96081a <=( (not A169)  and  A170 );
 a96084a <=( (not A167)  and  (not A168) );
 a96085a <=( a96084a  and  a96081a );
 a96088a <=( (not A199)  and  A166 );
 a96091a <=( A201  and  A200 );
 a96092a <=( a96091a  and  a96088a );
 a96093a <=( a96092a  and  a96085a );
 a96096a <=( (not A265)  and  A202 );
 a96099a <=( (not A267)  and  A266 );
 a96100a <=( a96099a  and  a96096a );
 a96103a <=( (not A269)  and  (not A268) );
 a96106a <=( A302  and  (not A300) );
 a96107a <=( a96106a  and  a96103a );
 a96108a <=( a96107a  and  a96100a );
 a96111a <=( (not A169)  and  A170 );
 a96114a <=( (not A167)  and  (not A168) );
 a96115a <=( a96114a  and  a96111a );
 a96118a <=( (not A199)  and  A166 );
 a96121a <=( A201  and  A200 );
 a96122a <=( a96121a  and  a96118a );
 a96123a <=( a96122a  and  a96115a );
 a96126a <=( (not A265)  and  A202 );
 a96129a <=( (not A267)  and  A266 );
 a96130a <=( a96129a  and  a96126a );
 a96133a <=( (not A269)  and  (not A268) );
 a96136a <=( A299  and  A298 );
 a96137a <=( a96136a  and  a96133a );
 a96138a <=( a96137a  and  a96130a );
 a96141a <=( (not A169)  and  A170 );
 a96144a <=( (not A167)  and  (not A168) );
 a96145a <=( a96144a  and  a96141a );
 a96148a <=( (not A199)  and  A166 );
 a96151a <=( A201  and  A200 );
 a96152a <=( a96151a  and  a96148a );
 a96153a <=( a96152a  and  a96145a );
 a96156a <=( (not A265)  and  A202 );
 a96159a <=( (not A267)  and  A266 );
 a96160a <=( a96159a  and  a96156a );
 a96163a <=( (not A269)  and  (not A268) );
 a96166a <=( (not A299)  and  (not A298) );
 a96167a <=( a96166a  and  a96163a );
 a96168a <=( a96167a  and  a96160a );
 a96171a <=( (not A169)  and  A170 );
 a96174a <=( (not A167)  and  (not A168) );
 a96175a <=( a96174a  and  a96171a );
 a96178a <=( (not A199)  and  A166 );
 a96181a <=( A201  and  A200 );
 a96182a <=( a96181a  and  a96178a );
 a96183a <=( a96182a  and  a96175a );
 a96186a <=( A265  and  A202 );
 a96189a <=( A267  and  (not A266) );
 a96190a <=( a96189a  and  a96186a );
 a96193a <=( A300  and  A268 );
 a96196a <=( (not A302)  and  (not A301) );
 a96197a <=( a96196a  and  a96193a );
 a96198a <=( a96197a  and  a96190a );
 a96201a <=( (not A169)  and  A170 );
 a96204a <=( (not A167)  and  (not A168) );
 a96205a <=( a96204a  and  a96201a );
 a96208a <=( (not A199)  and  A166 );
 a96211a <=( A201  and  A200 );
 a96212a <=( a96211a  and  a96208a );
 a96213a <=( a96212a  and  a96205a );
 a96216a <=( A265  and  A202 );
 a96219a <=( A267  and  (not A266) );
 a96220a <=( a96219a  and  a96216a );
 a96223a <=( A300  and  A269 );
 a96226a <=( (not A302)  and  (not A301) );
 a96227a <=( a96226a  and  a96223a );
 a96228a <=( a96227a  and  a96220a );
 a96231a <=( (not A169)  and  A170 );
 a96234a <=( (not A167)  and  (not A168) );
 a96235a <=( a96234a  and  a96231a );
 a96238a <=( (not A199)  and  A166 );
 a96241a <=( A201  and  A200 );
 a96242a <=( a96241a  and  a96238a );
 a96243a <=( a96242a  and  a96235a );
 a96246a <=( A265  and  A202 );
 a96249a <=( (not A267)  and  (not A266) );
 a96250a <=( a96249a  and  a96246a );
 a96253a <=( (not A269)  and  (not A268) );
 a96256a <=( A301  and  (not A300) );
 a96257a <=( a96256a  and  a96253a );
 a96258a <=( a96257a  and  a96250a );
 a96261a <=( (not A169)  and  A170 );
 a96264a <=( (not A167)  and  (not A168) );
 a96265a <=( a96264a  and  a96261a );
 a96268a <=( (not A199)  and  A166 );
 a96271a <=( A201  and  A200 );
 a96272a <=( a96271a  and  a96268a );
 a96273a <=( a96272a  and  a96265a );
 a96276a <=( A265  and  A202 );
 a96279a <=( (not A267)  and  (not A266) );
 a96280a <=( a96279a  and  a96276a );
 a96283a <=( (not A269)  and  (not A268) );
 a96286a <=( A302  and  (not A300) );
 a96287a <=( a96286a  and  a96283a );
 a96288a <=( a96287a  and  a96280a );
 a96291a <=( (not A169)  and  A170 );
 a96294a <=( (not A167)  and  (not A168) );
 a96295a <=( a96294a  and  a96291a );
 a96298a <=( (not A199)  and  A166 );
 a96301a <=( A201  and  A200 );
 a96302a <=( a96301a  and  a96298a );
 a96303a <=( a96302a  and  a96295a );
 a96306a <=( A265  and  A202 );
 a96309a <=( (not A267)  and  (not A266) );
 a96310a <=( a96309a  and  a96306a );
 a96313a <=( (not A269)  and  (not A268) );
 a96316a <=( A299  and  A298 );
 a96317a <=( a96316a  and  a96313a );
 a96318a <=( a96317a  and  a96310a );
 a96321a <=( (not A169)  and  A170 );
 a96324a <=( (not A167)  and  (not A168) );
 a96325a <=( a96324a  and  a96321a );
 a96328a <=( (not A199)  and  A166 );
 a96331a <=( A201  and  A200 );
 a96332a <=( a96331a  and  a96328a );
 a96333a <=( a96332a  and  a96325a );
 a96336a <=( A265  and  A202 );
 a96339a <=( (not A267)  and  (not A266) );
 a96340a <=( a96339a  and  a96336a );
 a96343a <=( (not A269)  and  (not A268) );
 a96346a <=( (not A299)  and  (not A298) );
 a96347a <=( a96346a  and  a96343a );
 a96348a <=( a96347a  and  a96340a );
 a96351a <=( (not A169)  and  A170 );
 a96354a <=( (not A167)  and  (not A168) );
 a96355a <=( a96354a  and  a96351a );
 a96358a <=( (not A199)  and  A166 );
 a96361a <=( A201  and  A200 );
 a96362a <=( a96361a  and  a96358a );
 a96363a <=( a96362a  and  a96355a );
 a96366a <=( (not A265)  and  A203 );
 a96369a <=( A267  and  A266 );
 a96370a <=( a96369a  and  a96366a );
 a96373a <=( A300  and  A268 );
 a96376a <=( (not A302)  and  (not A301) );
 a96377a <=( a96376a  and  a96373a );
 a96378a <=( a96377a  and  a96370a );
 a96381a <=( (not A169)  and  A170 );
 a96384a <=( (not A167)  and  (not A168) );
 a96385a <=( a96384a  and  a96381a );
 a96388a <=( (not A199)  and  A166 );
 a96391a <=( A201  and  A200 );
 a96392a <=( a96391a  and  a96388a );
 a96393a <=( a96392a  and  a96385a );
 a96396a <=( (not A265)  and  A203 );
 a96399a <=( A267  and  A266 );
 a96400a <=( a96399a  and  a96396a );
 a96403a <=( A300  and  A269 );
 a96406a <=( (not A302)  and  (not A301) );
 a96407a <=( a96406a  and  a96403a );
 a96408a <=( a96407a  and  a96400a );
 a96411a <=( (not A169)  and  A170 );
 a96414a <=( (not A167)  and  (not A168) );
 a96415a <=( a96414a  and  a96411a );
 a96418a <=( (not A199)  and  A166 );
 a96421a <=( A201  and  A200 );
 a96422a <=( a96421a  and  a96418a );
 a96423a <=( a96422a  and  a96415a );
 a96426a <=( (not A265)  and  A203 );
 a96429a <=( (not A267)  and  A266 );
 a96430a <=( a96429a  and  a96426a );
 a96433a <=( (not A269)  and  (not A268) );
 a96436a <=( A301  and  (not A300) );
 a96437a <=( a96436a  and  a96433a );
 a96438a <=( a96437a  and  a96430a );
 a96441a <=( (not A169)  and  A170 );
 a96444a <=( (not A167)  and  (not A168) );
 a96445a <=( a96444a  and  a96441a );
 a96448a <=( (not A199)  and  A166 );
 a96451a <=( A201  and  A200 );
 a96452a <=( a96451a  and  a96448a );
 a96453a <=( a96452a  and  a96445a );
 a96456a <=( (not A265)  and  A203 );
 a96459a <=( (not A267)  and  A266 );
 a96460a <=( a96459a  and  a96456a );
 a96463a <=( (not A269)  and  (not A268) );
 a96466a <=( A302  and  (not A300) );
 a96467a <=( a96466a  and  a96463a );
 a96468a <=( a96467a  and  a96460a );
 a96471a <=( (not A169)  and  A170 );
 a96474a <=( (not A167)  and  (not A168) );
 a96475a <=( a96474a  and  a96471a );
 a96478a <=( (not A199)  and  A166 );
 a96481a <=( A201  and  A200 );
 a96482a <=( a96481a  and  a96478a );
 a96483a <=( a96482a  and  a96475a );
 a96486a <=( (not A265)  and  A203 );
 a96489a <=( (not A267)  and  A266 );
 a96490a <=( a96489a  and  a96486a );
 a96493a <=( (not A269)  and  (not A268) );
 a96496a <=( A299  and  A298 );
 a96497a <=( a96496a  and  a96493a );
 a96498a <=( a96497a  and  a96490a );
 a96501a <=( (not A169)  and  A170 );
 a96504a <=( (not A167)  and  (not A168) );
 a96505a <=( a96504a  and  a96501a );
 a96508a <=( (not A199)  and  A166 );
 a96511a <=( A201  and  A200 );
 a96512a <=( a96511a  and  a96508a );
 a96513a <=( a96512a  and  a96505a );
 a96516a <=( (not A265)  and  A203 );
 a96519a <=( (not A267)  and  A266 );
 a96520a <=( a96519a  and  a96516a );
 a96523a <=( (not A269)  and  (not A268) );
 a96526a <=( (not A299)  and  (not A298) );
 a96527a <=( a96526a  and  a96523a );
 a96528a <=( a96527a  and  a96520a );
 a96531a <=( (not A169)  and  A170 );
 a96534a <=( (not A167)  and  (not A168) );
 a96535a <=( a96534a  and  a96531a );
 a96538a <=( (not A199)  and  A166 );
 a96541a <=( A201  and  A200 );
 a96542a <=( a96541a  and  a96538a );
 a96543a <=( a96542a  and  a96535a );
 a96546a <=( A265  and  A203 );
 a96549a <=( A267  and  (not A266) );
 a96550a <=( a96549a  and  a96546a );
 a96553a <=( A300  and  A268 );
 a96556a <=( (not A302)  and  (not A301) );
 a96557a <=( a96556a  and  a96553a );
 a96558a <=( a96557a  and  a96550a );
 a96561a <=( (not A169)  and  A170 );
 a96564a <=( (not A167)  and  (not A168) );
 a96565a <=( a96564a  and  a96561a );
 a96568a <=( (not A199)  and  A166 );
 a96571a <=( A201  and  A200 );
 a96572a <=( a96571a  and  a96568a );
 a96573a <=( a96572a  and  a96565a );
 a96576a <=( A265  and  A203 );
 a96579a <=( A267  and  (not A266) );
 a96580a <=( a96579a  and  a96576a );
 a96583a <=( A300  and  A269 );
 a96586a <=( (not A302)  and  (not A301) );
 a96587a <=( a96586a  and  a96583a );
 a96588a <=( a96587a  and  a96580a );
 a96591a <=( (not A169)  and  A170 );
 a96594a <=( (not A167)  and  (not A168) );
 a96595a <=( a96594a  and  a96591a );
 a96598a <=( (not A199)  and  A166 );
 a96601a <=( A201  and  A200 );
 a96602a <=( a96601a  and  a96598a );
 a96603a <=( a96602a  and  a96595a );
 a96606a <=( A265  and  A203 );
 a96609a <=( (not A267)  and  (not A266) );
 a96610a <=( a96609a  and  a96606a );
 a96613a <=( (not A269)  and  (not A268) );
 a96616a <=( A301  and  (not A300) );
 a96617a <=( a96616a  and  a96613a );
 a96618a <=( a96617a  and  a96610a );
 a96621a <=( (not A169)  and  A170 );
 a96624a <=( (not A167)  and  (not A168) );
 a96625a <=( a96624a  and  a96621a );
 a96628a <=( (not A199)  and  A166 );
 a96631a <=( A201  and  A200 );
 a96632a <=( a96631a  and  a96628a );
 a96633a <=( a96632a  and  a96625a );
 a96636a <=( A265  and  A203 );
 a96639a <=( (not A267)  and  (not A266) );
 a96640a <=( a96639a  and  a96636a );
 a96643a <=( (not A269)  and  (not A268) );
 a96646a <=( A302  and  (not A300) );
 a96647a <=( a96646a  and  a96643a );
 a96648a <=( a96647a  and  a96640a );
 a96651a <=( (not A169)  and  A170 );
 a96654a <=( (not A167)  and  (not A168) );
 a96655a <=( a96654a  and  a96651a );
 a96658a <=( (not A199)  and  A166 );
 a96661a <=( A201  and  A200 );
 a96662a <=( a96661a  and  a96658a );
 a96663a <=( a96662a  and  a96655a );
 a96666a <=( A265  and  A203 );
 a96669a <=( (not A267)  and  (not A266) );
 a96670a <=( a96669a  and  a96666a );
 a96673a <=( (not A269)  and  (not A268) );
 a96676a <=( A299  and  A298 );
 a96677a <=( a96676a  and  a96673a );
 a96678a <=( a96677a  and  a96670a );
 a96681a <=( (not A169)  and  A170 );
 a96684a <=( (not A167)  and  (not A168) );
 a96685a <=( a96684a  and  a96681a );
 a96688a <=( (not A199)  and  A166 );
 a96691a <=( A201  and  A200 );
 a96692a <=( a96691a  and  a96688a );
 a96693a <=( a96692a  and  a96685a );
 a96696a <=( A265  and  A203 );
 a96699a <=( (not A267)  and  (not A266) );
 a96700a <=( a96699a  and  a96696a );
 a96703a <=( (not A269)  and  (not A268) );
 a96706a <=( (not A299)  and  (not A298) );
 a96707a <=( a96706a  and  a96703a );
 a96708a <=( a96707a  and  a96700a );
 a96711a <=( (not A169)  and  A170 );
 a96714a <=( (not A167)  and  (not A168) );
 a96715a <=( a96714a  and  a96711a );
 a96718a <=( (not A199)  and  A166 );
 a96721a <=( (not A201)  and  A200 );
 a96722a <=( a96721a  and  a96718a );
 a96723a <=( a96722a  and  a96715a );
 a96726a <=( (not A203)  and  (not A202) );
 a96729a <=( A266  and  (not A265) );
 a96730a <=( a96729a  and  a96726a );
 a96733a <=( A268  and  A267 );
 a96736a <=( A301  and  (not A300) );
 a96737a <=( a96736a  and  a96733a );
 a96738a <=( a96737a  and  a96730a );
 a96741a <=( (not A169)  and  A170 );
 a96744a <=( (not A167)  and  (not A168) );
 a96745a <=( a96744a  and  a96741a );
 a96748a <=( (not A199)  and  A166 );
 a96751a <=( (not A201)  and  A200 );
 a96752a <=( a96751a  and  a96748a );
 a96753a <=( a96752a  and  a96745a );
 a96756a <=( (not A203)  and  (not A202) );
 a96759a <=( A266  and  (not A265) );
 a96760a <=( a96759a  and  a96756a );
 a96763a <=( A268  and  A267 );
 a96766a <=( A302  and  (not A300) );
 a96767a <=( a96766a  and  a96763a );
 a96768a <=( a96767a  and  a96760a );
 a96771a <=( (not A169)  and  A170 );
 a96774a <=( (not A167)  and  (not A168) );
 a96775a <=( a96774a  and  a96771a );
 a96778a <=( (not A199)  and  A166 );
 a96781a <=( (not A201)  and  A200 );
 a96782a <=( a96781a  and  a96778a );
 a96783a <=( a96782a  and  a96775a );
 a96786a <=( (not A203)  and  (not A202) );
 a96789a <=( A266  and  (not A265) );
 a96790a <=( a96789a  and  a96786a );
 a96793a <=( A268  and  A267 );
 a96796a <=( A299  and  A298 );
 a96797a <=( a96796a  and  a96793a );
 a96798a <=( a96797a  and  a96790a );
 a96801a <=( (not A169)  and  A170 );
 a96804a <=( (not A167)  and  (not A168) );
 a96805a <=( a96804a  and  a96801a );
 a96808a <=( (not A199)  and  A166 );
 a96811a <=( (not A201)  and  A200 );
 a96812a <=( a96811a  and  a96808a );
 a96813a <=( a96812a  and  a96805a );
 a96816a <=( (not A203)  and  (not A202) );
 a96819a <=( A266  and  (not A265) );
 a96820a <=( a96819a  and  a96816a );
 a96823a <=( A268  and  A267 );
 a96826a <=( (not A299)  and  (not A298) );
 a96827a <=( a96826a  and  a96823a );
 a96828a <=( a96827a  and  a96820a );
 a96831a <=( (not A169)  and  A170 );
 a96834a <=( (not A167)  and  (not A168) );
 a96835a <=( a96834a  and  a96831a );
 a96838a <=( (not A199)  and  A166 );
 a96841a <=( (not A201)  and  A200 );
 a96842a <=( a96841a  and  a96838a );
 a96843a <=( a96842a  and  a96835a );
 a96846a <=( (not A203)  and  (not A202) );
 a96849a <=( A266  and  (not A265) );
 a96850a <=( a96849a  and  a96846a );
 a96853a <=( A269  and  A267 );
 a96856a <=( A301  and  (not A300) );
 a96857a <=( a96856a  and  a96853a );
 a96858a <=( a96857a  and  a96850a );
 a96861a <=( (not A169)  and  A170 );
 a96864a <=( (not A167)  and  (not A168) );
 a96865a <=( a96864a  and  a96861a );
 a96868a <=( (not A199)  and  A166 );
 a96871a <=( (not A201)  and  A200 );
 a96872a <=( a96871a  and  a96868a );
 a96873a <=( a96872a  and  a96865a );
 a96876a <=( (not A203)  and  (not A202) );
 a96879a <=( A266  and  (not A265) );
 a96880a <=( a96879a  and  a96876a );
 a96883a <=( A269  and  A267 );
 a96886a <=( A302  and  (not A300) );
 a96887a <=( a96886a  and  a96883a );
 a96888a <=( a96887a  and  a96880a );
 a96891a <=( (not A169)  and  A170 );
 a96894a <=( (not A167)  and  (not A168) );
 a96895a <=( a96894a  and  a96891a );
 a96898a <=( (not A199)  and  A166 );
 a96901a <=( (not A201)  and  A200 );
 a96902a <=( a96901a  and  a96898a );
 a96903a <=( a96902a  and  a96895a );
 a96906a <=( (not A203)  and  (not A202) );
 a96909a <=( A266  and  (not A265) );
 a96910a <=( a96909a  and  a96906a );
 a96913a <=( A269  and  A267 );
 a96916a <=( A299  and  A298 );
 a96917a <=( a96916a  and  a96913a );
 a96918a <=( a96917a  and  a96910a );
 a96921a <=( (not A169)  and  A170 );
 a96924a <=( (not A167)  and  (not A168) );
 a96925a <=( a96924a  and  a96921a );
 a96928a <=( (not A199)  and  A166 );
 a96931a <=( (not A201)  and  A200 );
 a96932a <=( a96931a  and  a96928a );
 a96933a <=( a96932a  and  a96925a );
 a96936a <=( (not A203)  and  (not A202) );
 a96939a <=( A266  and  (not A265) );
 a96940a <=( a96939a  and  a96936a );
 a96943a <=( A269  and  A267 );
 a96946a <=( (not A299)  and  (not A298) );
 a96947a <=( a96946a  and  a96943a );
 a96948a <=( a96947a  and  a96940a );
 a96951a <=( (not A169)  and  A170 );
 a96954a <=( (not A167)  and  (not A168) );
 a96955a <=( a96954a  and  a96951a );
 a96958a <=( (not A199)  and  A166 );
 a96961a <=( (not A201)  and  A200 );
 a96962a <=( a96961a  and  a96958a );
 a96963a <=( a96962a  and  a96955a );
 a96966a <=( (not A203)  and  (not A202) );
 a96969a <=( (not A266)  and  A265 );
 a96970a <=( a96969a  and  a96966a );
 a96973a <=( A268  and  A267 );
 a96976a <=( A301  and  (not A300) );
 a96977a <=( a96976a  and  a96973a );
 a96978a <=( a96977a  and  a96970a );
 a96981a <=( (not A169)  and  A170 );
 a96984a <=( (not A167)  and  (not A168) );
 a96985a <=( a96984a  and  a96981a );
 a96988a <=( (not A199)  and  A166 );
 a96991a <=( (not A201)  and  A200 );
 a96992a <=( a96991a  and  a96988a );
 a96993a <=( a96992a  and  a96985a );
 a96996a <=( (not A203)  and  (not A202) );
 a96999a <=( (not A266)  and  A265 );
 a97000a <=( a96999a  and  a96996a );
 a97003a <=( A268  and  A267 );
 a97006a <=( A302  and  (not A300) );
 a97007a <=( a97006a  and  a97003a );
 a97008a <=( a97007a  and  a97000a );
 a97011a <=( (not A169)  and  A170 );
 a97014a <=( (not A167)  and  (not A168) );
 a97015a <=( a97014a  and  a97011a );
 a97018a <=( (not A199)  and  A166 );
 a97021a <=( (not A201)  and  A200 );
 a97022a <=( a97021a  and  a97018a );
 a97023a <=( a97022a  and  a97015a );
 a97026a <=( (not A203)  and  (not A202) );
 a97029a <=( (not A266)  and  A265 );
 a97030a <=( a97029a  and  a97026a );
 a97033a <=( A268  and  A267 );
 a97036a <=( A299  and  A298 );
 a97037a <=( a97036a  and  a97033a );
 a97038a <=( a97037a  and  a97030a );
 a97041a <=( (not A169)  and  A170 );
 a97044a <=( (not A167)  and  (not A168) );
 a97045a <=( a97044a  and  a97041a );
 a97048a <=( (not A199)  and  A166 );
 a97051a <=( (not A201)  and  A200 );
 a97052a <=( a97051a  and  a97048a );
 a97053a <=( a97052a  and  a97045a );
 a97056a <=( (not A203)  and  (not A202) );
 a97059a <=( (not A266)  and  A265 );
 a97060a <=( a97059a  and  a97056a );
 a97063a <=( A268  and  A267 );
 a97066a <=( (not A299)  and  (not A298) );
 a97067a <=( a97066a  and  a97063a );
 a97068a <=( a97067a  and  a97060a );
 a97071a <=( (not A169)  and  A170 );
 a97074a <=( (not A167)  and  (not A168) );
 a97075a <=( a97074a  and  a97071a );
 a97078a <=( (not A199)  and  A166 );
 a97081a <=( (not A201)  and  A200 );
 a97082a <=( a97081a  and  a97078a );
 a97083a <=( a97082a  and  a97075a );
 a97086a <=( (not A203)  and  (not A202) );
 a97089a <=( (not A266)  and  A265 );
 a97090a <=( a97089a  and  a97086a );
 a97093a <=( A269  and  A267 );
 a97096a <=( A301  and  (not A300) );
 a97097a <=( a97096a  and  a97093a );
 a97098a <=( a97097a  and  a97090a );
 a97101a <=( (not A169)  and  A170 );
 a97104a <=( (not A167)  and  (not A168) );
 a97105a <=( a97104a  and  a97101a );
 a97108a <=( (not A199)  and  A166 );
 a97111a <=( (not A201)  and  A200 );
 a97112a <=( a97111a  and  a97108a );
 a97113a <=( a97112a  and  a97105a );
 a97116a <=( (not A203)  and  (not A202) );
 a97119a <=( (not A266)  and  A265 );
 a97120a <=( a97119a  and  a97116a );
 a97123a <=( A269  and  A267 );
 a97126a <=( A302  and  (not A300) );
 a97127a <=( a97126a  and  a97123a );
 a97128a <=( a97127a  and  a97120a );
 a97131a <=( (not A169)  and  A170 );
 a97134a <=( (not A167)  and  (not A168) );
 a97135a <=( a97134a  and  a97131a );
 a97138a <=( (not A199)  and  A166 );
 a97141a <=( (not A201)  and  A200 );
 a97142a <=( a97141a  and  a97138a );
 a97143a <=( a97142a  and  a97135a );
 a97146a <=( (not A203)  and  (not A202) );
 a97149a <=( (not A266)  and  A265 );
 a97150a <=( a97149a  and  a97146a );
 a97153a <=( A269  and  A267 );
 a97156a <=( A299  and  A298 );
 a97157a <=( a97156a  and  a97153a );
 a97158a <=( a97157a  and  a97150a );
 a97161a <=( (not A169)  and  A170 );
 a97164a <=( (not A167)  and  (not A168) );
 a97165a <=( a97164a  and  a97161a );
 a97168a <=( (not A199)  and  A166 );
 a97171a <=( (not A201)  and  A200 );
 a97172a <=( a97171a  and  a97168a );
 a97173a <=( a97172a  and  a97165a );
 a97176a <=( (not A203)  and  (not A202) );
 a97179a <=( (not A266)  and  A265 );
 a97180a <=( a97179a  and  a97176a );
 a97183a <=( A269  and  A267 );
 a97186a <=( (not A299)  and  (not A298) );
 a97187a <=( a97186a  and  a97183a );
 a97188a <=( a97187a  and  a97180a );
 a97191a <=( (not A169)  and  A170 );
 a97194a <=( (not A167)  and  (not A168) );
 a97195a <=( a97194a  and  a97191a );
 a97198a <=( A199  and  A166 );
 a97201a <=( A201  and  (not A200) );
 a97202a <=( a97201a  and  a97198a );
 a97203a <=( a97202a  and  a97195a );
 a97206a <=( (not A265)  and  A202 );
 a97209a <=( A267  and  A266 );
 a97210a <=( a97209a  and  a97206a );
 a97213a <=( A300  and  A268 );
 a97216a <=( (not A302)  and  (not A301) );
 a97217a <=( a97216a  and  a97213a );
 a97218a <=( a97217a  and  a97210a );
 a97221a <=( (not A169)  and  A170 );
 a97224a <=( (not A167)  and  (not A168) );
 a97225a <=( a97224a  and  a97221a );
 a97228a <=( A199  and  A166 );
 a97231a <=( A201  and  (not A200) );
 a97232a <=( a97231a  and  a97228a );
 a97233a <=( a97232a  and  a97225a );
 a97236a <=( (not A265)  and  A202 );
 a97239a <=( A267  and  A266 );
 a97240a <=( a97239a  and  a97236a );
 a97243a <=( A300  and  A269 );
 a97246a <=( (not A302)  and  (not A301) );
 a97247a <=( a97246a  and  a97243a );
 a97248a <=( a97247a  and  a97240a );
 a97251a <=( (not A169)  and  A170 );
 a97254a <=( (not A167)  and  (not A168) );
 a97255a <=( a97254a  and  a97251a );
 a97258a <=( A199  and  A166 );
 a97261a <=( A201  and  (not A200) );
 a97262a <=( a97261a  and  a97258a );
 a97263a <=( a97262a  and  a97255a );
 a97266a <=( (not A265)  and  A202 );
 a97269a <=( (not A267)  and  A266 );
 a97270a <=( a97269a  and  a97266a );
 a97273a <=( (not A269)  and  (not A268) );
 a97276a <=( A301  and  (not A300) );
 a97277a <=( a97276a  and  a97273a );
 a97278a <=( a97277a  and  a97270a );
 a97281a <=( (not A169)  and  A170 );
 a97284a <=( (not A167)  and  (not A168) );
 a97285a <=( a97284a  and  a97281a );
 a97288a <=( A199  and  A166 );
 a97291a <=( A201  and  (not A200) );
 a97292a <=( a97291a  and  a97288a );
 a97293a <=( a97292a  and  a97285a );
 a97296a <=( (not A265)  and  A202 );
 a97299a <=( (not A267)  and  A266 );
 a97300a <=( a97299a  and  a97296a );
 a97303a <=( (not A269)  and  (not A268) );
 a97306a <=( A302  and  (not A300) );
 a97307a <=( a97306a  and  a97303a );
 a97308a <=( a97307a  and  a97300a );
 a97311a <=( (not A169)  and  A170 );
 a97314a <=( (not A167)  and  (not A168) );
 a97315a <=( a97314a  and  a97311a );
 a97318a <=( A199  and  A166 );
 a97321a <=( A201  and  (not A200) );
 a97322a <=( a97321a  and  a97318a );
 a97323a <=( a97322a  and  a97315a );
 a97326a <=( (not A265)  and  A202 );
 a97329a <=( (not A267)  and  A266 );
 a97330a <=( a97329a  and  a97326a );
 a97333a <=( (not A269)  and  (not A268) );
 a97336a <=( A299  and  A298 );
 a97337a <=( a97336a  and  a97333a );
 a97338a <=( a97337a  and  a97330a );
 a97341a <=( (not A169)  and  A170 );
 a97344a <=( (not A167)  and  (not A168) );
 a97345a <=( a97344a  and  a97341a );
 a97348a <=( A199  and  A166 );
 a97351a <=( A201  and  (not A200) );
 a97352a <=( a97351a  and  a97348a );
 a97353a <=( a97352a  and  a97345a );
 a97356a <=( (not A265)  and  A202 );
 a97359a <=( (not A267)  and  A266 );
 a97360a <=( a97359a  and  a97356a );
 a97363a <=( (not A269)  and  (not A268) );
 a97366a <=( (not A299)  and  (not A298) );
 a97367a <=( a97366a  and  a97363a );
 a97368a <=( a97367a  and  a97360a );
 a97371a <=( (not A169)  and  A170 );
 a97374a <=( (not A167)  and  (not A168) );
 a97375a <=( a97374a  and  a97371a );
 a97378a <=( A199  and  A166 );
 a97381a <=( A201  and  (not A200) );
 a97382a <=( a97381a  and  a97378a );
 a97383a <=( a97382a  and  a97375a );
 a97386a <=( A265  and  A202 );
 a97389a <=( A267  and  (not A266) );
 a97390a <=( a97389a  and  a97386a );
 a97393a <=( A300  and  A268 );
 a97396a <=( (not A302)  and  (not A301) );
 a97397a <=( a97396a  and  a97393a );
 a97398a <=( a97397a  and  a97390a );
 a97401a <=( (not A169)  and  A170 );
 a97404a <=( (not A167)  and  (not A168) );
 a97405a <=( a97404a  and  a97401a );
 a97408a <=( A199  and  A166 );
 a97411a <=( A201  and  (not A200) );
 a97412a <=( a97411a  and  a97408a );
 a97413a <=( a97412a  and  a97405a );
 a97416a <=( A265  and  A202 );
 a97419a <=( A267  and  (not A266) );
 a97420a <=( a97419a  and  a97416a );
 a97423a <=( A300  and  A269 );
 a97426a <=( (not A302)  and  (not A301) );
 a97427a <=( a97426a  and  a97423a );
 a97428a <=( a97427a  and  a97420a );
 a97431a <=( (not A169)  and  A170 );
 a97434a <=( (not A167)  and  (not A168) );
 a97435a <=( a97434a  and  a97431a );
 a97438a <=( A199  and  A166 );
 a97441a <=( A201  and  (not A200) );
 a97442a <=( a97441a  and  a97438a );
 a97443a <=( a97442a  and  a97435a );
 a97446a <=( A265  and  A202 );
 a97449a <=( (not A267)  and  (not A266) );
 a97450a <=( a97449a  and  a97446a );
 a97453a <=( (not A269)  and  (not A268) );
 a97456a <=( A301  and  (not A300) );
 a97457a <=( a97456a  and  a97453a );
 a97458a <=( a97457a  and  a97450a );
 a97461a <=( (not A169)  and  A170 );
 a97464a <=( (not A167)  and  (not A168) );
 a97465a <=( a97464a  and  a97461a );
 a97468a <=( A199  and  A166 );
 a97471a <=( A201  and  (not A200) );
 a97472a <=( a97471a  and  a97468a );
 a97473a <=( a97472a  and  a97465a );
 a97476a <=( A265  and  A202 );
 a97479a <=( (not A267)  and  (not A266) );
 a97480a <=( a97479a  and  a97476a );
 a97483a <=( (not A269)  and  (not A268) );
 a97486a <=( A302  and  (not A300) );
 a97487a <=( a97486a  and  a97483a );
 a97488a <=( a97487a  and  a97480a );
 a97491a <=( (not A169)  and  A170 );
 a97494a <=( (not A167)  and  (not A168) );
 a97495a <=( a97494a  and  a97491a );
 a97498a <=( A199  and  A166 );
 a97501a <=( A201  and  (not A200) );
 a97502a <=( a97501a  and  a97498a );
 a97503a <=( a97502a  and  a97495a );
 a97506a <=( A265  and  A202 );
 a97509a <=( (not A267)  and  (not A266) );
 a97510a <=( a97509a  and  a97506a );
 a97513a <=( (not A269)  and  (not A268) );
 a97516a <=( A299  and  A298 );
 a97517a <=( a97516a  and  a97513a );
 a97518a <=( a97517a  and  a97510a );
 a97521a <=( (not A169)  and  A170 );
 a97524a <=( (not A167)  and  (not A168) );
 a97525a <=( a97524a  and  a97521a );
 a97528a <=( A199  and  A166 );
 a97531a <=( A201  and  (not A200) );
 a97532a <=( a97531a  and  a97528a );
 a97533a <=( a97532a  and  a97525a );
 a97536a <=( A265  and  A202 );
 a97539a <=( (not A267)  and  (not A266) );
 a97540a <=( a97539a  and  a97536a );
 a97543a <=( (not A269)  and  (not A268) );
 a97546a <=( (not A299)  and  (not A298) );
 a97547a <=( a97546a  and  a97543a );
 a97548a <=( a97547a  and  a97540a );
 a97551a <=( (not A169)  and  A170 );
 a97554a <=( (not A167)  and  (not A168) );
 a97555a <=( a97554a  and  a97551a );
 a97558a <=( A199  and  A166 );
 a97561a <=( A201  and  (not A200) );
 a97562a <=( a97561a  and  a97558a );
 a97563a <=( a97562a  and  a97555a );
 a97566a <=( (not A265)  and  A203 );
 a97569a <=( A267  and  A266 );
 a97570a <=( a97569a  and  a97566a );
 a97573a <=( A300  and  A268 );
 a97576a <=( (not A302)  and  (not A301) );
 a97577a <=( a97576a  and  a97573a );
 a97578a <=( a97577a  and  a97570a );
 a97581a <=( (not A169)  and  A170 );
 a97584a <=( (not A167)  and  (not A168) );
 a97585a <=( a97584a  and  a97581a );
 a97588a <=( A199  and  A166 );
 a97591a <=( A201  and  (not A200) );
 a97592a <=( a97591a  and  a97588a );
 a97593a <=( a97592a  and  a97585a );
 a97596a <=( (not A265)  and  A203 );
 a97599a <=( A267  and  A266 );
 a97600a <=( a97599a  and  a97596a );
 a97603a <=( A300  and  A269 );
 a97606a <=( (not A302)  and  (not A301) );
 a97607a <=( a97606a  and  a97603a );
 a97608a <=( a97607a  and  a97600a );
 a97611a <=( (not A169)  and  A170 );
 a97614a <=( (not A167)  and  (not A168) );
 a97615a <=( a97614a  and  a97611a );
 a97618a <=( A199  and  A166 );
 a97621a <=( A201  and  (not A200) );
 a97622a <=( a97621a  and  a97618a );
 a97623a <=( a97622a  and  a97615a );
 a97626a <=( (not A265)  and  A203 );
 a97629a <=( (not A267)  and  A266 );
 a97630a <=( a97629a  and  a97626a );
 a97633a <=( (not A269)  and  (not A268) );
 a97636a <=( A301  and  (not A300) );
 a97637a <=( a97636a  and  a97633a );
 a97638a <=( a97637a  and  a97630a );
 a97641a <=( (not A169)  and  A170 );
 a97644a <=( (not A167)  and  (not A168) );
 a97645a <=( a97644a  and  a97641a );
 a97648a <=( A199  and  A166 );
 a97651a <=( A201  and  (not A200) );
 a97652a <=( a97651a  and  a97648a );
 a97653a <=( a97652a  and  a97645a );
 a97656a <=( (not A265)  and  A203 );
 a97659a <=( (not A267)  and  A266 );
 a97660a <=( a97659a  and  a97656a );
 a97663a <=( (not A269)  and  (not A268) );
 a97666a <=( A302  and  (not A300) );
 a97667a <=( a97666a  and  a97663a );
 a97668a <=( a97667a  and  a97660a );
 a97671a <=( (not A169)  and  A170 );
 a97674a <=( (not A167)  and  (not A168) );
 a97675a <=( a97674a  and  a97671a );
 a97678a <=( A199  and  A166 );
 a97681a <=( A201  and  (not A200) );
 a97682a <=( a97681a  and  a97678a );
 a97683a <=( a97682a  and  a97675a );
 a97686a <=( (not A265)  and  A203 );
 a97689a <=( (not A267)  and  A266 );
 a97690a <=( a97689a  and  a97686a );
 a97693a <=( (not A269)  and  (not A268) );
 a97696a <=( A299  and  A298 );
 a97697a <=( a97696a  and  a97693a );
 a97698a <=( a97697a  and  a97690a );
 a97701a <=( (not A169)  and  A170 );
 a97704a <=( (not A167)  and  (not A168) );
 a97705a <=( a97704a  and  a97701a );
 a97708a <=( A199  and  A166 );
 a97711a <=( A201  and  (not A200) );
 a97712a <=( a97711a  and  a97708a );
 a97713a <=( a97712a  and  a97705a );
 a97716a <=( (not A265)  and  A203 );
 a97719a <=( (not A267)  and  A266 );
 a97720a <=( a97719a  and  a97716a );
 a97723a <=( (not A269)  and  (not A268) );
 a97726a <=( (not A299)  and  (not A298) );
 a97727a <=( a97726a  and  a97723a );
 a97728a <=( a97727a  and  a97720a );
 a97731a <=( (not A169)  and  A170 );
 a97734a <=( (not A167)  and  (not A168) );
 a97735a <=( a97734a  and  a97731a );
 a97738a <=( A199  and  A166 );
 a97741a <=( A201  and  (not A200) );
 a97742a <=( a97741a  and  a97738a );
 a97743a <=( a97742a  and  a97735a );
 a97746a <=( A265  and  A203 );
 a97749a <=( A267  and  (not A266) );
 a97750a <=( a97749a  and  a97746a );
 a97753a <=( A300  and  A268 );
 a97756a <=( (not A302)  and  (not A301) );
 a97757a <=( a97756a  and  a97753a );
 a97758a <=( a97757a  and  a97750a );
 a97761a <=( (not A169)  and  A170 );
 a97764a <=( (not A167)  and  (not A168) );
 a97765a <=( a97764a  and  a97761a );
 a97768a <=( A199  and  A166 );
 a97771a <=( A201  and  (not A200) );
 a97772a <=( a97771a  and  a97768a );
 a97773a <=( a97772a  and  a97765a );
 a97776a <=( A265  and  A203 );
 a97779a <=( A267  and  (not A266) );
 a97780a <=( a97779a  and  a97776a );
 a97783a <=( A300  and  A269 );
 a97786a <=( (not A302)  and  (not A301) );
 a97787a <=( a97786a  and  a97783a );
 a97788a <=( a97787a  and  a97780a );
 a97791a <=( (not A169)  and  A170 );
 a97794a <=( (not A167)  and  (not A168) );
 a97795a <=( a97794a  and  a97791a );
 a97798a <=( A199  and  A166 );
 a97801a <=( A201  and  (not A200) );
 a97802a <=( a97801a  and  a97798a );
 a97803a <=( a97802a  and  a97795a );
 a97806a <=( A265  and  A203 );
 a97809a <=( (not A267)  and  (not A266) );
 a97810a <=( a97809a  and  a97806a );
 a97813a <=( (not A269)  and  (not A268) );
 a97816a <=( A301  and  (not A300) );
 a97817a <=( a97816a  and  a97813a );
 a97818a <=( a97817a  and  a97810a );
 a97821a <=( (not A169)  and  A170 );
 a97824a <=( (not A167)  and  (not A168) );
 a97825a <=( a97824a  and  a97821a );
 a97828a <=( A199  and  A166 );
 a97831a <=( A201  and  (not A200) );
 a97832a <=( a97831a  and  a97828a );
 a97833a <=( a97832a  and  a97825a );
 a97836a <=( A265  and  A203 );
 a97839a <=( (not A267)  and  (not A266) );
 a97840a <=( a97839a  and  a97836a );
 a97843a <=( (not A269)  and  (not A268) );
 a97846a <=( A302  and  (not A300) );
 a97847a <=( a97846a  and  a97843a );
 a97848a <=( a97847a  and  a97840a );
 a97851a <=( (not A169)  and  A170 );
 a97854a <=( (not A167)  and  (not A168) );
 a97855a <=( a97854a  and  a97851a );
 a97858a <=( A199  and  A166 );
 a97861a <=( A201  and  (not A200) );
 a97862a <=( a97861a  and  a97858a );
 a97863a <=( a97862a  and  a97855a );
 a97866a <=( A265  and  A203 );
 a97869a <=( (not A267)  and  (not A266) );
 a97870a <=( a97869a  and  a97866a );
 a97873a <=( (not A269)  and  (not A268) );
 a97876a <=( A299  and  A298 );
 a97877a <=( a97876a  and  a97873a );
 a97878a <=( a97877a  and  a97870a );
 a97881a <=( (not A169)  and  A170 );
 a97884a <=( (not A167)  and  (not A168) );
 a97885a <=( a97884a  and  a97881a );
 a97888a <=( A199  and  A166 );
 a97891a <=( A201  and  (not A200) );
 a97892a <=( a97891a  and  a97888a );
 a97893a <=( a97892a  and  a97885a );
 a97896a <=( A265  and  A203 );
 a97899a <=( (not A267)  and  (not A266) );
 a97900a <=( a97899a  and  a97896a );
 a97903a <=( (not A269)  and  (not A268) );
 a97906a <=( (not A299)  and  (not A298) );
 a97907a <=( a97906a  and  a97903a );
 a97908a <=( a97907a  and  a97900a );
 a97911a <=( (not A169)  and  A170 );
 a97914a <=( (not A167)  and  (not A168) );
 a97915a <=( a97914a  and  a97911a );
 a97918a <=( A199  and  A166 );
 a97921a <=( (not A201)  and  (not A200) );
 a97922a <=( a97921a  and  a97918a );
 a97923a <=( a97922a  and  a97915a );
 a97926a <=( (not A203)  and  (not A202) );
 a97929a <=( A266  and  (not A265) );
 a97930a <=( a97929a  and  a97926a );
 a97933a <=( A268  and  A267 );
 a97936a <=( A301  and  (not A300) );
 a97937a <=( a97936a  and  a97933a );
 a97938a <=( a97937a  and  a97930a );
 a97941a <=( (not A169)  and  A170 );
 a97944a <=( (not A167)  and  (not A168) );
 a97945a <=( a97944a  and  a97941a );
 a97948a <=( A199  and  A166 );
 a97951a <=( (not A201)  and  (not A200) );
 a97952a <=( a97951a  and  a97948a );
 a97953a <=( a97952a  and  a97945a );
 a97956a <=( (not A203)  and  (not A202) );
 a97959a <=( A266  and  (not A265) );
 a97960a <=( a97959a  and  a97956a );
 a97963a <=( A268  and  A267 );
 a97966a <=( A302  and  (not A300) );
 a97967a <=( a97966a  and  a97963a );
 a97968a <=( a97967a  and  a97960a );
 a97971a <=( (not A169)  and  A170 );
 a97974a <=( (not A167)  and  (not A168) );
 a97975a <=( a97974a  and  a97971a );
 a97978a <=( A199  and  A166 );
 a97981a <=( (not A201)  and  (not A200) );
 a97982a <=( a97981a  and  a97978a );
 a97983a <=( a97982a  and  a97975a );
 a97986a <=( (not A203)  and  (not A202) );
 a97989a <=( A266  and  (not A265) );
 a97990a <=( a97989a  and  a97986a );
 a97993a <=( A268  and  A267 );
 a97996a <=( A299  and  A298 );
 a97997a <=( a97996a  and  a97993a );
 a97998a <=( a97997a  and  a97990a );
 a98001a <=( (not A169)  and  A170 );
 a98004a <=( (not A167)  and  (not A168) );
 a98005a <=( a98004a  and  a98001a );
 a98008a <=( A199  and  A166 );
 a98011a <=( (not A201)  and  (not A200) );
 a98012a <=( a98011a  and  a98008a );
 a98013a <=( a98012a  and  a98005a );
 a98016a <=( (not A203)  and  (not A202) );
 a98019a <=( A266  and  (not A265) );
 a98020a <=( a98019a  and  a98016a );
 a98023a <=( A268  and  A267 );
 a98026a <=( (not A299)  and  (not A298) );
 a98027a <=( a98026a  and  a98023a );
 a98028a <=( a98027a  and  a98020a );
 a98031a <=( (not A169)  and  A170 );
 a98034a <=( (not A167)  and  (not A168) );
 a98035a <=( a98034a  and  a98031a );
 a98038a <=( A199  and  A166 );
 a98041a <=( (not A201)  and  (not A200) );
 a98042a <=( a98041a  and  a98038a );
 a98043a <=( a98042a  and  a98035a );
 a98046a <=( (not A203)  and  (not A202) );
 a98049a <=( A266  and  (not A265) );
 a98050a <=( a98049a  and  a98046a );
 a98053a <=( A269  and  A267 );
 a98056a <=( A301  and  (not A300) );
 a98057a <=( a98056a  and  a98053a );
 a98058a <=( a98057a  and  a98050a );
 a98061a <=( (not A169)  and  A170 );
 a98064a <=( (not A167)  and  (not A168) );
 a98065a <=( a98064a  and  a98061a );
 a98068a <=( A199  and  A166 );
 a98071a <=( (not A201)  and  (not A200) );
 a98072a <=( a98071a  and  a98068a );
 a98073a <=( a98072a  and  a98065a );
 a98076a <=( (not A203)  and  (not A202) );
 a98079a <=( A266  and  (not A265) );
 a98080a <=( a98079a  and  a98076a );
 a98083a <=( A269  and  A267 );
 a98086a <=( A302  and  (not A300) );
 a98087a <=( a98086a  and  a98083a );
 a98088a <=( a98087a  and  a98080a );
 a98091a <=( (not A169)  and  A170 );
 a98094a <=( (not A167)  and  (not A168) );
 a98095a <=( a98094a  and  a98091a );
 a98098a <=( A199  and  A166 );
 a98101a <=( (not A201)  and  (not A200) );
 a98102a <=( a98101a  and  a98098a );
 a98103a <=( a98102a  and  a98095a );
 a98106a <=( (not A203)  and  (not A202) );
 a98109a <=( A266  and  (not A265) );
 a98110a <=( a98109a  and  a98106a );
 a98113a <=( A269  and  A267 );
 a98116a <=( A299  and  A298 );
 a98117a <=( a98116a  and  a98113a );
 a98118a <=( a98117a  and  a98110a );
 a98121a <=( (not A169)  and  A170 );
 a98124a <=( (not A167)  and  (not A168) );
 a98125a <=( a98124a  and  a98121a );
 a98128a <=( A199  and  A166 );
 a98131a <=( (not A201)  and  (not A200) );
 a98132a <=( a98131a  and  a98128a );
 a98133a <=( a98132a  and  a98125a );
 a98136a <=( (not A203)  and  (not A202) );
 a98139a <=( A266  and  (not A265) );
 a98140a <=( a98139a  and  a98136a );
 a98143a <=( A269  and  A267 );
 a98146a <=( (not A299)  and  (not A298) );
 a98147a <=( a98146a  and  a98143a );
 a98148a <=( a98147a  and  a98140a );
 a98151a <=( (not A169)  and  A170 );
 a98154a <=( (not A167)  and  (not A168) );
 a98155a <=( a98154a  and  a98151a );
 a98158a <=( A199  and  A166 );
 a98161a <=( (not A201)  and  (not A200) );
 a98162a <=( a98161a  and  a98158a );
 a98163a <=( a98162a  and  a98155a );
 a98166a <=( (not A203)  and  (not A202) );
 a98169a <=( (not A266)  and  A265 );
 a98170a <=( a98169a  and  a98166a );
 a98173a <=( A268  and  A267 );
 a98176a <=( A301  and  (not A300) );
 a98177a <=( a98176a  and  a98173a );
 a98178a <=( a98177a  and  a98170a );
 a98181a <=( (not A169)  and  A170 );
 a98184a <=( (not A167)  and  (not A168) );
 a98185a <=( a98184a  and  a98181a );
 a98188a <=( A199  and  A166 );
 a98191a <=( (not A201)  and  (not A200) );
 a98192a <=( a98191a  and  a98188a );
 a98193a <=( a98192a  and  a98185a );
 a98196a <=( (not A203)  and  (not A202) );
 a98199a <=( (not A266)  and  A265 );
 a98200a <=( a98199a  and  a98196a );
 a98203a <=( A268  and  A267 );
 a98206a <=( A302  and  (not A300) );
 a98207a <=( a98206a  and  a98203a );
 a98208a <=( a98207a  and  a98200a );
 a98211a <=( (not A169)  and  A170 );
 a98214a <=( (not A167)  and  (not A168) );
 a98215a <=( a98214a  and  a98211a );
 a98218a <=( A199  and  A166 );
 a98221a <=( (not A201)  and  (not A200) );
 a98222a <=( a98221a  and  a98218a );
 a98223a <=( a98222a  and  a98215a );
 a98226a <=( (not A203)  and  (not A202) );
 a98229a <=( (not A266)  and  A265 );
 a98230a <=( a98229a  and  a98226a );
 a98233a <=( A268  and  A267 );
 a98236a <=( A299  and  A298 );
 a98237a <=( a98236a  and  a98233a );
 a98238a <=( a98237a  and  a98230a );
 a98241a <=( (not A169)  and  A170 );
 a98244a <=( (not A167)  and  (not A168) );
 a98245a <=( a98244a  and  a98241a );
 a98248a <=( A199  and  A166 );
 a98251a <=( (not A201)  and  (not A200) );
 a98252a <=( a98251a  and  a98248a );
 a98253a <=( a98252a  and  a98245a );
 a98256a <=( (not A203)  and  (not A202) );
 a98259a <=( (not A266)  and  A265 );
 a98260a <=( a98259a  and  a98256a );
 a98263a <=( A268  and  A267 );
 a98266a <=( (not A299)  and  (not A298) );
 a98267a <=( a98266a  and  a98263a );
 a98268a <=( a98267a  and  a98260a );
 a98271a <=( (not A169)  and  A170 );
 a98274a <=( (not A167)  and  (not A168) );
 a98275a <=( a98274a  and  a98271a );
 a98278a <=( A199  and  A166 );
 a98281a <=( (not A201)  and  (not A200) );
 a98282a <=( a98281a  and  a98278a );
 a98283a <=( a98282a  and  a98275a );
 a98286a <=( (not A203)  and  (not A202) );
 a98289a <=( (not A266)  and  A265 );
 a98290a <=( a98289a  and  a98286a );
 a98293a <=( A269  and  A267 );
 a98296a <=( A301  and  (not A300) );
 a98297a <=( a98296a  and  a98293a );
 a98298a <=( a98297a  and  a98290a );
 a98301a <=( (not A169)  and  A170 );
 a98304a <=( (not A167)  and  (not A168) );
 a98305a <=( a98304a  and  a98301a );
 a98308a <=( A199  and  A166 );
 a98311a <=( (not A201)  and  (not A200) );
 a98312a <=( a98311a  and  a98308a );
 a98313a <=( a98312a  and  a98305a );
 a98316a <=( (not A203)  and  (not A202) );
 a98319a <=( (not A266)  and  A265 );
 a98320a <=( a98319a  and  a98316a );
 a98323a <=( A269  and  A267 );
 a98326a <=( A302  and  (not A300) );
 a98327a <=( a98326a  and  a98323a );
 a98328a <=( a98327a  and  a98320a );
 a98331a <=( (not A169)  and  A170 );
 a98334a <=( (not A167)  and  (not A168) );
 a98335a <=( a98334a  and  a98331a );
 a98338a <=( A199  and  A166 );
 a98341a <=( (not A201)  and  (not A200) );
 a98342a <=( a98341a  and  a98338a );
 a98343a <=( a98342a  and  a98335a );
 a98346a <=( (not A203)  and  (not A202) );
 a98349a <=( (not A266)  and  A265 );
 a98350a <=( a98349a  and  a98346a );
 a98353a <=( A269  and  A267 );
 a98356a <=( A299  and  A298 );
 a98357a <=( a98356a  and  a98353a );
 a98358a <=( a98357a  and  a98350a );
 a98361a <=( (not A169)  and  A170 );
 a98364a <=( (not A167)  and  (not A168) );
 a98365a <=( a98364a  and  a98361a );
 a98368a <=( A199  and  A166 );
 a98371a <=( (not A201)  and  (not A200) );
 a98372a <=( a98371a  and  a98368a );
 a98373a <=( a98372a  and  a98365a );
 a98376a <=( (not A203)  and  (not A202) );
 a98379a <=( (not A266)  and  A265 );
 a98380a <=( a98379a  and  a98376a );
 a98383a <=( A269  and  A267 );
 a98386a <=( (not A299)  and  (not A298) );
 a98387a <=( a98386a  and  a98383a );
 a98388a <=( a98387a  and  a98380a );
 a98391a <=( A168  and  (not A170) );
 a98394a <=( (not A166)  and  A167 );
 a98395a <=( a98394a  and  a98391a );
 a98398a <=( A200  and  (not A199) );
 a98401a <=( (not A202)  and  (not A201) );
 a98402a <=( a98401a  and  a98398a );
 a98403a <=( a98402a  and  a98395a );
 a98406a <=( (not A265)  and  (not A203) );
 a98409a <=( (not A267)  and  A266 );
 a98410a <=( a98409a  and  a98406a );
 a98413a <=( (not A269)  and  (not A268) );
 a98417a <=( (not A302)  and  (not A301) );
 a98418a <=( A300  and  a98417a );
 a98419a <=( a98418a  and  a98413a );
 a98420a <=( a98419a  and  a98410a );
 a98423a <=( A168  and  (not A170) );
 a98426a <=( (not A166)  and  A167 );
 a98427a <=( a98426a  and  a98423a );
 a98430a <=( A200  and  (not A199) );
 a98433a <=( (not A202)  and  (not A201) );
 a98434a <=( a98433a  and  a98430a );
 a98435a <=( a98434a  and  a98427a );
 a98438a <=( A265  and  (not A203) );
 a98441a <=( (not A267)  and  (not A266) );
 a98442a <=( a98441a  and  a98438a );
 a98445a <=( (not A269)  and  (not A268) );
 a98449a <=( (not A302)  and  (not A301) );
 a98450a <=( A300  and  a98449a );
 a98451a <=( a98450a  and  a98445a );
 a98452a <=( a98451a  and  a98442a );
 a98455a <=( A168  and  (not A170) );
 a98458a <=( (not A166)  and  A167 );
 a98459a <=( a98458a  and  a98455a );
 a98462a <=( (not A200)  and  A199 );
 a98465a <=( (not A202)  and  (not A201) );
 a98466a <=( a98465a  and  a98462a );
 a98467a <=( a98466a  and  a98459a );
 a98470a <=( (not A265)  and  (not A203) );
 a98473a <=( (not A267)  and  A266 );
 a98474a <=( a98473a  and  a98470a );
 a98477a <=( (not A269)  and  (not A268) );
 a98481a <=( (not A302)  and  (not A301) );
 a98482a <=( A300  and  a98481a );
 a98483a <=( a98482a  and  a98477a );
 a98484a <=( a98483a  and  a98474a );
 a98487a <=( A168  and  (not A170) );
 a98490a <=( (not A166)  and  A167 );
 a98491a <=( a98490a  and  a98487a );
 a98494a <=( (not A200)  and  A199 );
 a98497a <=( (not A202)  and  (not A201) );
 a98498a <=( a98497a  and  a98494a );
 a98499a <=( a98498a  and  a98491a );
 a98502a <=( A265  and  (not A203) );
 a98505a <=( (not A267)  and  (not A266) );
 a98506a <=( a98505a  and  a98502a );
 a98509a <=( (not A269)  and  (not A268) );
 a98513a <=( (not A302)  and  (not A301) );
 a98514a <=( A300  and  a98513a );
 a98515a <=( a98514a  and  a98509a );
 a98516a <=( a98515a  and  a98506a );
 a98519a <=( A168  and  (not A170) );
 a98522a <=( A166  and  (not A167) );
 a98523a <=( a98522a  and  a98519a );
 a98526a <=( A200  and  (not A199) );
 a98529a <=( (not A202)  and  (not A201) );
 a98530a <=( a98529a  and  a98526a );
 a98531a <=( a98530a  and  a98523a );
 a98534a <=( (not A265)  and  (not A203) );
 a98537a <=( (not A267)  and  A266 );
 a98538a <=( a98537a  and  a98534a );
 a98541a <=( (not A269)  and  (not A268) );
 a98545a <=( (not A302)  and  (not A301) );
 a98546a <=( A300  and  a98545a );
 a98547a <=( a98546a  and  a98541a );
 a98548a <=( a98547a  and  a98538a );
 a98551a <=( A168  and  (not A170) );
 a98554a <=( A166  and  (not A167) );
 a98555a <=( a98554a  and  a98551a );
 a98558a <=( A200  and  (not A199) );
 a98561a <=( (not A202)  and  (not A201) );
 a98562a <=( a98561a  and  a98558a );
 a98563a <=( a98562a  and  a98555a );
 a98566a <=( A265  and  (not A203) );
 a98569a <=( (not A267)  and  (not A266) );
 a98570a <=( a98569a  and  a98566a );
 a98573a <=( (not A269)  and  (not A268) );
 a98577a <=( (not A302)  and  (not A301) );
 a98578a <=( A300  and  a98577a );
 a98579a <=( a98578a  and  a98573a );
 a98580a <=( a98579a  and  a98570a );
 a98583a <=( A168  and  (not A170) );
 a98586a <=( A166  and  (not A167) );
 a98587a <=( a98586a  and  a98583a );
 a98590a <=( (not A200)  and  A199 );
 a98593a <=( (not A202)  and  (not A201) );
 a98594a <=( a98593a  and  a98590a );
 a98595a <=( a98594a  and  a98587a );
 a98598a <=( (not A265)  and  (not A203) );
 a98601a <=( (not A267)  and  A266 );
 a98602a <=( a98601a  and  a98598a );
 a98605a <=( (not A269)  and  (not A268) );
 a98609a <=( (not A302)  and  (not A301) );
 a98610a <=( A300  and  a98609a );
 a98611a <=( a98610a  and  a98605a );
 a98612a <=( a98611a  and  a98602a );
 a98615a <=( A168  and  (not A170) );
 a98618a <=( A166  and  (not A167) );
 a98619a <=( a98618a  and  a98615a );
 a98622a <=( (not A200)  and  A199 );
 a98625a <=( (not A202)  and  (not A201) );
 a98626a <=( a98625a  and  a98622a );
 a98627a <=( a98626a  and  a98619a );
 a98630a <=( A265  and  (not A203) );
 a98633a <=( (not A267)  and  (not A266) );
 a98634a <=( a98633a  and  a98630a );
 a98637a <=( (not A269)  and  (not A268) );
 a98641a <=( (not A302)  and  (not A301) );
 a98642a <=( A300  and  a98641a );
 a98643a <=( a98642a  and  a98637a );
 a98644a <=( a98643a  and  a98634a );
 a98647a <=( A168  and  A169 );
 a98650a <=( (not A166)  and  A167 );
 a98651a <=( a98650a  and  a98647a );
 a98654a <=( A200  and  (not A199) );
 a98657a <=( (not A202)  and  (not A201) );
 a98658a <=( a98657a  and  a98654a );
 a98659a <=( a98658a  and  a98651a );
 a98662a <=( (not A265)  and  (not A203) );
 a98665a <=( (not A267)  and  A266 );
 a98666a <=( a98665a  and  a98662a );
 a98669a <=( (not A269)  and  (not A268) );
 a98673a <=( (not A302)  and  (not A301) );
 a98674a <=( A300  and  a98673a );
 a98675a <=( a98674a  and  a98669a );
 a98676a <=( a98675a  and  a98666a );
 a98679a <=( A168  and  A169 );
 a98682a <=( (not A166)  and  A167 );
 a98683a <=( a98682a  and  a98679a );
 a98686a <=( A200  and  (not A199) );
 a98689a <=( (not A202)  and  (not A201) );
 a98690a <=( a98689a  and  a98686a );
 a98691a <=( a98690a  and  a98683a );
 a98694a <=( A265  and  (not A203) );
 a98697a <=( (not A267)  and  (not A266) );
 a98698a <=( a98697a  and  a98694a );
 a98701a <=( (not A269)  and  (not A268) );
 a98705a <=( (not A302)  and  (not A301) );
 a98706a <=( A300  and  a98705a );
 a98707a <=( a98706a  and  a98701a );
 a98708a <=( a98707a  and  a98698a );
 a98711a <=( A168  and  A169 );
 a98714a <=( (not A166)  and  A167 );
 a98715a <=( a98714a  and  a98711a );
 a98718a <=( (not A200)  and  A199 );
 a98721a <=( (not A202)  and  (not A201) );
 a98722a <=( a98721a  and  a98718a );
 a98723a <=( a98722a  and  a98715a );
 a98726a <=( (not A265)  and  (not A203) );
 a98729a <=( (not A267)  and  A266 );
 a98730a <=( a98729a  and  a98726a );
 a98733a <=( (not A269)  and  (not A268) );
 a98737a <=( (not A302)  and  (not A301) );
 a98738a <=( A300  and  a98737a );
 a98739a <=( a98738a  and  a98733a );
 a98740a <=( a98739a  and  a98730a );
 a98743a <=( A168  and  A169 );
 a98746a <=( (not A166)  and  A167 );
 a98747a <=( a98746a  and  a98743a );
 a98750a <=( (not A200)  and  A199 );
 a98753a <=( (not A202)  and  (not A201) );
 a98754a <=( a98753a  and  a98750a );
 a98755a <=( a98754a  and  a98747a );
 a98758a <=( A265  and  (not A203) );
 a98761a <=( (not A267)  and  (not A266) );
 a98762a <=( a98761a  and  a98758a );
 a98765a <=( (not A269)  and  (not A268) );
 a98769a <=( (not A302)  and  (not A301) );
 a98770a <=( A300  and  a98769a );
 a98771a <=( a98770a  and  a98765a );
 a98772a <=( a98771a  and  a98762a );
 a98775a <=( A168  and  A169 );
 a98778a <=( A166  and  (not A167) );
 a98779a <=( a98778a  and  a98775a );
 a98782a <=( A200  and  (not A199) );
 a98785a <=( (not A202)  and  (not A201) );
 a98786a <=( a98785a  and  a98782a );
 a98787a <=( a98786a  and  a98779a );
 a98790a <=( (not A265)  and  (not A203) );
 a98793a <=( (not A267)  and  A266 );
 a98794a <=( a98793a  and  a98790a );
 a98797a <=( (not A269)  and  (not A268) );
 a98801a <=( (not A302)  and  (not A301) );
 a98802a <=( A300  and  a98801a );
 a98803a <=( a98802a  and  a98797a );
 a98804a <=( a98803a  and  a98794a );
 a98807a <=( A168  and  A169 );
 a98810a <=( A166  and  (not A167) );
 a98811a <=( a98810a  and  a98807a );
 a98814a <=( A200  and  (not A199) );
 a98817a <=( (not A202)  and  (not A201) );
 a98818a <=( a98817a  and  a98814a );
 a98819a <=( a98818a  and  a98811a );
 a98822a <=( A265  and  (not A203) );
 a98825a <=( (not A267)  and  (not A266) );
 a98826a <=( a98825a  and  a98822a );
 a98829a <=( (not A269)  and  (not A268) );
 a98833a <=( (not A302)  and  (not A301) );
 a98834a <=( A300  and  a98833a );
 a98835a <=( a98834a  and  a98829a );
 a98836a <=( a98835a  and  a98826a );
 a98839a <=( A168  and  A169 );
 a98842a <=( A166  and  (not A167) );
 a98843a <=( a98842a  and  a98839a );
 a98846a <=( (not A200)  and  A199 );
 a98849a <=( (not A202)  and  (not A201) );
 a98850a <=( a98849a  and  a98846a );
 a98851a <=( a98850a  and  a98843a );
 a98854a <=( (not A265)  and  (not A203) );
 a98857a <=( (not A267)  and  A266 );
 a98858a <=( a98857a  and  a98854a );
 a98861a <=( (not A269)  and  (not A268) );
 a98865a <=( (not A302)  and  (not A301) );
 a98866a <=( A300  and  a98865a );
 a98867a <=( a98866a  and  a98861a );
 a98868a <=( a98867a  and  a98858a );
 a98871a <=( A168  and  A169 );
 a98874a <=( A166  and  (not A167) );
 a98875a <=( a98874a  and  a98871a );
 a98878a <=( (not A200)  and  A199 );
 a98881a <=( (not A202)  and  (not A201) );
 a98882a <=( a98881a  and  a98878a );
 a98883a <=( a98882a  and  a98875a );
 a98886a <=( A265  and  (not A203) );
 a98889a <=( (not A267)  and  (not A266) );
 a98890a <=( a98889a  and  a98886a );
 a98893a <=( (not A269)  and  (not A268) );
 a98897a <=( (not A302)  and  (not A301) );
 a98898a <=( A300  and  a98897a );
 a98899a <=( a98898a  and  a98893a );
 a98900a <=( a98899a  and  a98890a );
 a98903a <=( (not A169)  and  A170 );
 a98906a <=( A167  and  (not A168) );
 a98907a <=( a98906a  and  a98903a );
 a98910a <=( (not A199)  and  (not A166) );
 a98913a <=( A201  and  A200 );
 a98914a <=( a98913a  and  a98910a );
 a98915a <=( a98914a  and  a98907a );
 a98918a <=( (not A265)  and  A202 );
 a98921a <=( (not A267)  and  A266 );
 a98922a <=( a98921a  and  a98918a );
 a98925a <=( (not A269)  and  (not A268) );
 a98929a <=( (not A302)  and  (not A301) );
 a98930a <=( A300  and  a98929a );
 a98931a <=( a98930a  and  a98925a );
 a98932a <=( a98931a  and  a98922a );
 a98935a <=( (not A169)  and  A170 );
 a98938a <=( A167  and  (not A168) );
 a98939a <=( a98938a  and  a98935a );
 a98942a <=( (not A199)  and  (not A166) );
 a98945a <=( A201  and  A200 );
 a98946a <=( a98945a  and  a98942a );
 a98947a <=( a98946a  and  a98939a );
 a98950a <=( A265  and  A202 );
 a98953a <=( (not A267)  and  (not A266) );
 a98954a <=( a98953a  and  a98950a );
 a98957a <=( (not A269)  and  (not A268) );
 a98961a <=( (not A302)  and  (not A301) );
 a98962a <=( A300  and  a98961a );
 a98963a <=( a98962a  and  a98957a );
 a98964a <=( a98963a  and  a98954a );
 a98967a <=( (not A169)  and  A170 );
 a98970a <=( A167  and  (not A168) );
 a98971a <=( a98970a  and  a98967a );
 a98974a <=( (not A199)  and  (not A166) );
 a98977a <=( A201  and  A200 );
 a98978a <=( a98977a  and  a98974a );
 a98979a <=( a98978a  and  a98971a );
 a98982a <=( (not A265)  and  A203 );
 a98985a <=( (not A267)  and  A266 );
 a98986a <=( a98985a  and  a98982a );
 a98989a <=( (not A269)  and  (not A268) );
 a98993a <=( (not A302)  and  (not A301) );
 a98994a <=( A300  and  a98993a );
 a98995a <=( a98994a  and  a98989a );
 a98996a <=( a98995a  and  a98986a );
 a98999a <=( (not A169)  and  A170 );
 a99002a <=( A167  and  (not A168) );
 a99003a <=( a99002a  and  a98999a );
 a99006a <=( (not A199)  and  (not A166) );
 a99009a <=( A201  and  A200 );
 a99010a <=( a99009a  and  a99006a );
 a99011a <=( a99010a  and  a99003a );
 a99014a <=( A265  and  A203 );
 a99017a <=( (not A267)  and  (not A266) );
 a99018a <=( a99017a  and  a99014a );
 a99021a <=( (not A269)  and  (not A268) );
 a99025a <=( (not A302)  and  (not A301) );
 a99026a <=( A300  and  a99025a );
 a99027a <=( a99026a  and  a99021a );
 a99028a <=( a99027a  and  a99018a );
 a99031a <=( (not A169)  and  A170 );
 a99034a <=( A167  and  (not A168) );
 a99035a <=( a99034a  and  a99031a );
 a99038a <=( (not A199)  and  (not A166) );
 a99041a <=( (not A201)  and  A200 );
 a99042a <=( a99041a  and  a99038a );
 a99043a <=( a99042a  and  a99035a );
 a99046a <=( (not A203)  and  (not A202) );
 a99049a <=( A266  and  (not A265) );
 a99050a <=( a99049a  and  a99046a );
 a99053a <=( A268  and  A267 );
 a99057a <=( (not A302)  and  (not A301) );
 a99058a <=( A300  and  a99057a );
 a99059a <=( a99058a  and  a99053a );
 a99060a <=( a99059a  and  a99050a );
 a99063a <=( (not A169)  and  A170 );
 a99066a <=( A167  and  (not A168) );
 a99067a <=( a99066a  and  a99063a );
 a99070a <=( (not A199)  and  (not A166) );
 a99073a <=( (not A201)  and  A200 );
 a99074a <=( a99073a  and  a99070a );
 a99075a <=( a99074a  and  a99067a );
 a99078a <=( (not A203)  and  (not A202) );
 a99081a <=( A266  and  (not A265) );
 a99082a <=( a99081a  and  a99078a );
 a99085a <=( A269  and  A267 );
 a99089a <=( (not A302)  and  (not A301) );
 a99090a <=( A300  and  a99089a );
 a99091a <=( a99090a  and  a99085a );
 a99092a <=( a99091a  and  a99082a );
 a99095a <=( (not A169)  and  A170 );
 a99098a <=( A167  and  (not A168) );
 a99099a <=( a99098a  and  a99095a );
 a99102a <=( (not A199)  and  (not A166) );
 a99105a <=( (not A201)  and  A200 );
 a99106a <=( a99105a  and  a99102a );
 a99107a <=( a99106a  and  a99099a );
 a99110a <=( (not A203)  and  (not A202) );
 a99113a <=( A266  and  (not A265) );
 a99114a <=( a99113a  and  a99110a );
 a99117a <=( (not A268)  and  (not A267) );
 a99121a <=( A301  and  (not A300) );
 a99122a <=( (not A269)  and  a99121a );
 a99123a <=( a99122a  and  a99117a );
 a99124a <=( a99123a  and  a99114a );
 a99127a <=( (not A169)  and  A170 );
 a99130a <=( A167  and  (not A168) );
 a99131a <=( a99130a  and  a99127a );
 a99134a <=( (not A199)  and  (not A166) );
 a99137a <=( (not A201)  and  A200 );
 a99138a <=( a99137a  and  a99134a );
 a99139a <=( a99138a  and  a99131a );
 a99142a <=( (not A203)  and  (not A202) );
 a99145a <=( A266  and  (not A265) );
 a99146a <=( a99145a  and  a99142a );
 a99149a <=( (not A268)  and  (not A267) );
 a99153a <=( A302  and  (not A300) );
 a99154a <=( (not A269)  and  a99153a );
 a99155a <=( a99154a  and  a99149a );
 a99156a <=( a99155a  and  a99146a );
 a99159a <=( (not A169)  and  A170 );
 a99162a <=( A167  and  (not A168) );
 a99163a <=( a99162a  and  a99159a );
 a99166a <=( (not A199)  and  (not A166) );
 a99169a <=( (not A201)  and  A200 );
 a99170a <=( a99169a  and  a99166a );
 a99171a <=( a99170a  and  a99163a );
 a99174a <=( (not A203)  and  (not A202) );
 a99177a <=( A266  and  (not A265) );
 a99178a <=( a99177a  and  a99174a );
 a99181a <=( (not A268)  and  (not A267) );
 a99185a <=( A299  and  A298 );
 a99186a <=( (not A269)  and  a99185a );
 a99187a <=( a99186a  and  a99181a );
 a99188a <=( a99187a  and  a99178a );
 a99191a <=( (not A169)  and  A170 );
 a99194a <=( A167  and  (not A168) );
 a99195a <=( a99194a  and  a99191a );
 a99198a <=( (not A199)  and  (not A166) );
 a99201a <=( (not A201)  and  A200 );
 a99202a <=( a99201a  and  a99198a );
 a99203a <=( a99202a  and  a99195a );
 a99206a <=( (not A203)  and  (not A202) );
 a99209a <=( A266  and  (not A265) );
 a99210a <=( a99209a  and  a99206a );
 a99213a <=( (not A268)  and  (not A267) );
 a99217a <=( (not A299)  and  (not A298) );
 a99218a <=( (not A269)  and  a99217a );
 a99219a <=( a99218a  and  a99213a );
 a99220a <=( a99219a  and  a99210a );
 a99223a <=( (not A169)  and  A170 );
 a99226a <=( A167  and  (not A168) );
 a99227a <=( a99226a  and  a99223a );
 a99230a <=( (not A199)  and  (not A166) );
 a99233a <=( (not A201)  and  A200 );
 a99234a <=( a99233a  and  a99230a );
 a99235a <=( a99234a  and  a99227a );
 a99238a <=( (not A203)  and  (not A202) );
 a99241a <=( (not A266)  and  A265 );
 a99242a <=( a99241a  and  a99238a );
 a99245a <=( A268  and  A267 );
 a99249a <=( (not A302)  and  (not A301) );
 a99250a <=( A300  and  a99249a );
 a99251a <=( a99250a  and  a99245a );
 a99252a <=( a99251a  and  a99242a );
 a99255a <=( (not A169)  and  A170 );
 a99258a <=( A167  and  (not A168) );
 a99259a <=( a99258a  and  a99255a );
 a99262a <=( (not A199)  and  (not A166) );
 a99265a <=( (not A201)  and  A200 );
 a99266a <=( a99265a  and  a99262a );
 a99267a <=( a99266a  and  a99259a );
 a99270a <=( (not A203)  and  (not A202) );
 a99273a <=( (not A266)  and  A265 );
 a99274a <=( a99273a  and  a99270a );
 a99277a <=( A269  and  A267 );
 a99281a <=( (not A302)  and  (not A301) );
 a99282a <=( A300  and  a99281a );
 a99283a <=( a99282a  and  a99277a );
 a99284a <=( a99283a  and  a99274a );
 a99287a <=( (not A169)  and  A170 );
 a99290a <=( A167  and  (not A168) );
 a99291a <=( a99290a  and  a99287a );
 a99294a <=( (not A199)  and  (not A166) );
 a99297a <=( (not A201)  and  A200 );
 a99298a <=( a99297a  and  a99294a );
 a99299a <=( a99298a  and  a99291a );
 a99302a <=( (not A203)  and  (not A202) );
 a99305a <=( (not A266)  and  A265 );
 a99306a <=( a99305a  and  a99302a );
 a99309a <=( (not A268)  and  (not A267) );
 a99313a <=( A301  and  (not A300) );
 a99314a <=( (not A269)  and  a99313a );
 a99315a <=( a99314a  and  a99309a );
 a99316a <=( a99315a  and  a99306a );
 a99319a <=( (not A169)  and  A170 );
 a99322a <=( A167  and  (not A168) );
 a99323a <=( a99322a  and  a99319a );
 a99326a <=( (not A199)  and  (not A166) );
 a99329a <=( (not A201)  and  A200 );
 a99330a <=( a99329a  and  a99326a );
 a99331a <=( a99330a  and  a99323a );
 a99334a <=( (not A203)  and  (not A202) );
 a99337a <=( (not A266)  and  A265 );
 a99338a <=( a99337a  and  a99334a );
 a99341a <=( (not A268)  and  (not A267) );
 a99345a <=( A302  and  (not A300) );
 a99346a <=( (not A269)  and  a99345a );
 a99347a <=( a99346a  and  a99341a );
 a99348a <=( a99347a  and  a99338a );
 a99351a <=( (not A169)  and  A170 );
 a99354a <=( A167  and  (not A168) );
 a99355a <=( a99354a  and  a99351a );
 a99358a <=( (not A199)  and  (not A166) );
 a99361a <=( (not A201)  and  A200 );
 a99362a <=( a99361a  and  a99358a );
 a99363a <=( a99362a  and  a99355a );
 a99366a <=( (not A203)  and  (not A202) );
 a99369a <=( (not A266)  and  A265 );
 a99370a <=( a99369a  and  a99366a );
 a99373a <=( (not A268)  and  (not A267) );
 a99377a <=( A299  and  A298 );
 a99378a <=( (not A269)  and  a99377a );
 a99379a <=( a99378a  and  a99373a );
 a99380a <=( a99379a  and  a99370a );
 a99383a <=( (not A169)  and  A170 );
 a99386a <=( A167  and  (not A168) );
 a99387a <=( a99386a  and  a99383a );
 a99390a <=( (not A199)  and  (not A166) );
 a99393a <=( (not A201)  and  A200 );
 a99394a <=( a99393a  and  a99390a );
 a99395a <=( a99394a  and  a99387a );
 a99398a <=( (not A203)  and  (not A202) );
 a99401a <=( (not A266)  and  A265 );
 a99402a <=( a99401a  and  a99398a );
 a99405a <=( (not A268)  and  (not A267) );
 a99409a <=( (not A299)  and  (not A298) );
 a99410a <=( (not A269)  and  a99409a );
 a99411a <=( a99410a  and  a99405a );
 a99412a <=( a99411a  and  a99402a );
 a99415a <=( (not A169)  and  A170 );
 a99418a <=( A167  and  (not A168) );
 a99419a <=( a99418a  and  a99415a );
 a99422a <=( A199  and  (not A166) );
 a99425a <=( A201  and  (not A200) );
 a99426a <=( a99425a  and  a99422a );
 a99427a <=( a99426a  and  a99419a );
 a99430a <=( (not A265)  and  A202 );
 a99433a <=( (not A267)  and  A266 );
 a99434a <=( a99433a  and  a99430a );
 a99437a <=( (not A269)  and  (not A268) );
 a99441a <=( (not A302)  and  (not A301) );
 a99442a <=( A300  and  a99441a );
 a99443a <=( a99442a  and  a99437a );
 a99444a <=( a99443a  and  a99434a );
 a99447a <=( (not A169)  and  A170 );
 a99450a <=( A167  and  (not A168) );
 a99451a <=( a99450a  and  a99447a );
 a99454a <=( A199  and  (not A166) );
 a99457a <=( A201  and  (not A200) );
 a99458a <=( a99457a  and  a99454a );
 a99459a <=( a99458a  and  a99451a );
 a99462a <=( A265  and  A202 );
 a99465a <=( (not A267)  and  (not A266) );
 a99466a <=( a99465a  and  a99462a );
 a99469a <=( (not A269)  and  (not A268) );
 a99473a <=( (not A302)  and  (not A301) );
 a99474a <=( A300  and  a99473a );
 a99475a <=( a99474a  and  a99469a );
 a99476a <=( a99475a  and  a99466a );
 a99479a <=( (not A169)  and  A170 );
 a99482a <=( A167  and  (not A168) );
 a99483a <=( a99482a  and  a99479a );
 a99486a <=( A199  and  (not A166) );
 a99489a <=( A201  and  (not A200) );
 a99490a <=( a99489a  and  a99486a );
 a99491a <=( a99490a  and  a99483a );
 a99494a <=( (not A265)  and  A203 );
 a99497a <=( (not A267)  and  A266 );
 a99498a <=( a99497a  and  a99494a );
 a99501a <=( (not A269)  and  (not A268) );
 a99505a <=( (not A302)  and  (not A301) );
 a99506a <=( A300  and  a99505a );
 a99507a <=( a99506a  and  a99501a );
 a99508a <=( a99507a  and  a99498a );
 a99511a <=( (not A169)  and  A170 );
 a99514a <=( A167  and  (not A168) );
 a99515a <=( a99514a  and  a99511a );
 a99518a <=( A199  and  (not A166) );
 a99521a <=( A201  and  (not A200) );
 a99522a <=( a99521a  and  a99518a );
 a99523a <=( a99522a  and  a99515a );
 a99526a <=( A265  and  A203 );
 a99529a <=( (not A267)  and  (not A266) );
 a99530a <=( a99529a  and  a99526a );
 a99533a <=( (not A269)  and  (not A268) );
 a99537a <=( (not A302)  and  (not A301) );
 a99538a <=( A300  and  a99537a );
 a99539a <=( a99538a  and  a99533a );
 a99540a <=( a99539a  and  a99530a );
 a99543a <=( (not A169)  and  A170 );
 a99546a <=( A167  and  (not A168) );
 a99547a <=( a99546a  and  a99543a );
 a99550a <=( A199  and  (not A166) );
 a99553a <=( (not A201)  and  (not A200) );
 a99554a <=( a99553a  and  a99550a );
 a99555a <=( a99554a  and  a99547a );
 a99558a <=( (not A203)  and  (not A202) );
 a99561a <=( A266  and  (not A265) );
 a99562a <=( a99561a  and  a99558a );
 a99565a <=( A268  and  A267 );
 a99569a <=( (not A302)  and  (not A301) );
 a99570a <=( A300  and  a99569a );
 a99571a <=( a99570a  and  a99565a );
 a99572a <=( a99571a  and  a99562a );
 a99575a <=( (not A169)  and  A170 );
 a99578a <=( A167  and  (not A168) );
 a99579a <=( a99578a  and  a99575a );
 a99582a <=( A199  and  (not A166) );
 a99585a <=( (not A201)  and  (not A200) );
 a99586a <=( a99585a  and  a99582a );
 a99587a <=( a99586a  and  a99579a );
 a99590a <=( (not A203)  and  (not A202) );
 a99593a <=( A266  and  (not A265) );
 a99594a <=( a99593a  and  a99590a );
 a99597a <=( A269  and  A267 );
 a99601a <=( (not A302)  and  (not A301) );
 a99602a <=( A300  and  a99601a );
 a99603a <=( a99602a  and  a99597a );
 a99604a <=( a99603a  and  a99594a );
 a99607a <=( (not A169)  and  A170 );
 a99610a <=( A167  and  (not A168) );
 a99611a <=( a99610a  and  a99607a );
 a99614a <=( A199  and  (not A166) );
 a99617a <=( (not A201)  and  (not A200) );
 a99618a <=( a99617a  and  a99614a );
 a99619a <=( a99618a  and  a99611a );
 a99622a <=( (not A203)  and  (not A202) );
 a99625a <=( A266  and  (not A265) );
 a99626a <=( a99625a  and  a99622a );
 a99629a <=( (not A268)  and  (not A267) );
 a99633a <=( A301  and  (not A300) );
 a99634a <=( (not A269)  and  a99633a );
 a99635a <=( a99634a  and  a99629a );
 a99636a <=( a99635a  and  a99626a );
 a99639a <=( (not A169)  and  A170 );
 a99642a <=( A167  and  (not A168) );
 a99643a <=( a99642a  and  a99639a );
 a99646a <=( A199  and  (not A166) );
 a99649a <=( (not A201)  and  (not A200) );
 a99650a <=( a99649a  and  a99646a );
 a99651a <=( a99650a  and  a99643a );
 a99654a <=( (not A203)  and  (not A202) );
 a99657a <=( A266  and  (not A265) );
 a99658a <=( a99657a  and  a99654a );
 a99661a <=( (not A268)  and  (not A267) );
 a99665a <=( A302  and  (not A300) );
 a99666a <=( (not A269)  and  a99665a );
 a99667a <=( a99666a  and  a99661a );
 a99668a <=( a99667a  and  a99658a );
 a99671a <=( (not A169)  and  A170 );
 a99674a <=( A167  and  (not A168) );
 a99675a <=( a99674a  and  a99671a );
 a99678a <=( A199  and  (not A166) );
 a99681a <=( (not A201)  and  (not A200) );
 a99682a <=( a99681a  and  a99678a );
 a99683a <=( a99682a  and  a99675a );
 a99686a <=( (not A203)  and  (not A202) );
 a99689a <=( A266  and  (not A265) );
 a99690a <=( a99689a  and  a99686a );
 a99693a <=( (not A268)  and  (not A267) );
 a99697a <=( A299  and  A298 );
 a99698a <=( (not A269)  and  a99697a );
 a99699a <=( a99698a  and  a99693a );
 a99700a <=( a99699a  and  a99690a );
 a99703a <=( (not A169)  and  A170 );
 a99706a <=( A167  and  (not A168) );
 a99707a <=( a99706a  and  a99703a );
 a99710a <=( A199  and  (not A166) );
 a99713a <=( (not A201)  and  (not A200) );
 a99714a <=( a99713a  and  a99710a );
 a99715a <=( a99714a  and  a99707a );
 a99718a <=( (not A203)  and  (not A202) );
 a99721a <=( A266  and  (not A265) );
 a99722a <=( a99721a  and  a99718a );
 a99725a <=( (not A268)  and  (not A267) );
 a99729a <=( (not A299)  and  (not A298) );
 a99730a <=( (not A269)  and  a99729a );
 a99731a <=( a99730a  and  a99725a );
 a99732a <=( a99731a  and  a99722a );
 a99735a <=( (not A169)  and  A170 );
 a99738a <=( A167  and  (not A168) );
 a99739a <=( a99738a  and  a99735a );
 a99742a <=( A199  and  (not A166) );
 a99745a <=( (not A201)  and  (not A200) );
 a99746a <=( a99745a  and  a99742a );
 a99747a <=( a99746a  and  a99739a );
 a99750a <=( (not A203)  and  (not A202) );
 a99753a <=( (not A266)  and  A265 );
 a99754a <=( a99753a  and  a99750a );
 a99757a <=( A268  and  A267 );
 a99761a <=( (not A302)  and  (not A301) );
 a99762a <=( A300  and  a99761a );
 a99763a <=( a99762a  and  a99757a );
 a99764a <=( a99763a  and  a99754a );
 a99767a <=( (not A169)  and  A170 );
 a99770a <=( A167  and  (not A168) );
 a99771a <=( a99770a  and  a99767a );
 a99774a <=( A199  and  (not A166) );
 a99777a <=( (not A201)  and  (not A200) );
 a99778a <=( a99777a  and  a99774a );
 a99779a <=( a99778a  and  a99771a );
 a99782a <=( (not A203)  and  (not A202) );
 a99785a <=( (not A266)  and  A265 );
 a99786a <=( a99785a  and  a99782a );
 a99789a <=( A269  and  A267 );
 a99793a <=( (not A302)  and  (not A301) );
 a99794a <=( A300  and  a99793a );
 a99795a <=( a99794a  and  a99789a );
 a99796a <=( a99795a  and  a99786a );
 a99799a <=( (not A169)  and  A170 );
 a99802a <=( A167  and  (not A168) );
 a99803a <=( a99802a  and  a99799a );
 a99806a <=( A199  and  (not A166) );
 a99809a <=( (not A201)  and  (not A200) );
 a99810a <=( a99809a  and  a99806a );
 a99811a <=( a99810a  and  a99803a );
 a99814a <=( (not A203)  and  (not A202) );
 a99817a <=( (not A266)  and  A265 );
 a99818a <=( a99817a  and  a99814a );
 a99821a <=( (not A268)  and  (not A267) );
 a99825a <=( A301  and  (not A300) );
 a99826a <=( (not A269)  and  a99825a );
 a99827a <=( a99826a  and  a99821a );
 a99828a <=( a99827a  and  a99818a );
 a99831a <=( (not A169)  and  A170 );
 a99834a <=( A167  and  (not A168) );
 a99835a <=( a99834a  and  a99831a );
 a99838a <=( A199  and  (not A166) );
 a99841a <=( (not A201)  and  (not A200) );
 a99842a <=( a99841a  and  a99838a );
 a99843a <=( a99842a  and  a99835a );
 a99846a <=( (not A203)  and  (not A202) );
 a99849a <=( (not A266)  and  A265 );
 a99850a <=( a99849a  and  a99846a );
 a99853a <=( (not A268)  and  (not A267) );
 a99857a <=( A302  and  (not A300) );
 a99858a <=( (not A269)  and  a99857a );
 a99859a <=( a99858a  and  a99853a );
 a99860a <=( a99859a  and  a99850a );
 a99863a <=( (not A169)  and  A170 );
 a99866a <=( A167  and  (not A168) );
 a99867a <=( a99866a  and  a99863a );
 a99870a <=( A199  and  (not A166) );
 a99873a <=( (not A201)  and  (not A200) );
 a99874a <=( a99873a  and  a99870a );
 a99875a <=( a99874a  and  a99867a );
 a99878a <=( (not A203)  and  (not A202) );
 a99881a <=( (not A266)  and  A265 );
 a99882a <=( a99881a  and  a99878a );
 a99885a <=( (not A268)  and  (not A267) );
 a99889a <=( A299  and  A298 );
 a99890a <=( (not A269)  and  a99889a );
 a99891a <=( a99890a  and  a99885a );
 a99892a <=( a99891a  and  a99882a );
 a99895a <=( (not A169)  and  A170 );
 a99898a <=( A167  and  (not A168) );
 a99899a <=( a99898a  and  a99895a );
 a99902a <=( A199  and  (not A166) );
 a99905a <=( (not A201)  and  (not A200) );
 a99906a <=( a99905a  and  a99902a );
 a99907a <=( a99906a  and  a99899a );
 a99910a <=( (not A203)  and  (not A202) );
 a99913a <=( (not A266)  and  A265 );
 a99914a <=( a99913a  and  a99910a );
 a99917a <=( (not A268)  and  (not A267) );
 a99921a <=( (not A299)  and  (not A298) );
 a99922a <=( (not A269)  and  a99921a );
 a99923a <=( a99922a  and  a99917a );
 a99924a <=( a99923a  and  a99914a );
 a99927a <=( (not A169)  and  A170 );
 a99930a <=( (not A167)  and  (not A168) );
 a99931a <=( a99930a  and  a99927a );
 a99934a <=( (not A199)  and  A166 );
 a99937a <=( A201  and  A200 );
 a99938a <=( a99937a  and  a99934a );
 a99939a <=( a99938a  and  a99931a );
 a99942a <=( (not A265)  and  A202 );
 a99945a <=( (not A267)  and  A266 );
 a99946a <=( a99945a  and  a99942a );
 a99949a <=( (not A269)  and  (not A268) );
 a99953a <=( (not A302)  and  (not A301) );
 a99954a <=( A300  and  a99953a );
 a99955a <=( a99954a  and  a99949a );
 a99956a <=( a99955a  and  a99946a );
 a99959a <=( (not A169)  and  A170 );
 a99962a <=( (not A167)  and  (not A168) );
 a99963a <=( a99962a  and  a99959a );
 a99966a <=( (not A199)  and  A166 );
 a99969a <=( A201  and  A200 );
 a99970a <=( a99969a  and  a99966a );
 a99971a <=( a99970a  and  a99963a );
 a99974a <=( A265  and  A202 );
 a99977a <=( (not A267)  and  (not A266) );
 a99978a <=( a99977a  and  a99974a );
 a99981a <=( (not A269)  and  (not A268) );
 a99985a <=( (not A302)  and  (not A301) );
 a99986a <=( A300  and  a99985a );
 a99987a <=( a99986a  and  a99981a );
 a99988a <=( a99987a  and  a99978a );
 a99991a <=( (not A169)  and  A170 );
 a99994a <=( (not A167)  and  (not A168) );
 a99995a <=( a99994a  and  a99991a );
 a99998a <=( (not A199)  and  A166 );
 a100001a <=( A201  and  A200 );
 a100002a <=( a100001a  and  a99998a );
 a100003a <=( a100002a  and  a99995a );
 a100006a <=( (not A265)  and  A203 );
 a100009a <=( (not A267)  and  A266 );
 a100010a <=( a100009a  and  a100006a );
 a100013a <=( (not A269)  and  (not A268) );
 a100017a <=( (not A302)  and  (not A301) );
 a100018a <=( A300  and  a100017a );
 a100019a <=( a100018a  and  a100013a );
 a100020a <=( a100019a  and  a100010a );
 a100023a <=( (not A169)  and  A170 );
 a100026a <=( (not A167)  and  (not A168) );
 a100027a <=( a100026a  and  a100023a );
 a100030a <=( (not A199)  and  A166 );
 a100033a <=( A201  and  A200 );
 a100034a <=( a100033a  and  a100030a );
 a100035a <=( a100034a  and  a100027a );
 a100038a <=( A265  and  A203 );
 a100041a <=( (not A267)  and  (not A266) );
 a100042a <=( a100041a  and  a100038a );
 a100045a <=( (not A269)  and  (not A268) );
 a100049a <=( (not A302)  and  (not A301) );
 a100050a <=( A300  and  a100049a );
 a100051a <=( a100050a  and  a100045a );
 a100052a <=( a100051a  and  a100042a );
 a100055a <=( (not A169)  and  A170 );
 a100058a <=( (not A167)  and  (not A168) );
 a100059a <=( a100058a  and  a100055a );
 a100062a <=( (not A199)  and  A166 );
 a100065a <=( (not A201)  and  A200 );
 a100066a <=( a100065a  and  a100062a );
 a100067a <=( a100066a  and  a100059a );
 a100070a <=( (not A203)  and  (not A202) );
 a100073a <=( A266  and  (not A265) );
 a100074a <=( a100073a  and  a100070a );
 a100077a <=( A268  and  A267 );
 a100081a <=( (not A302)  and  (not A301) );
 a100082a <=( A300  and  a100081a );
 a100083a <=( a100082a  and  a100077a );
 a100084a <=( a100083a  and  a100074a );
 a100087a <=( (not A169)  and  A170 );
 a100090a <=( (not A167)  and  (not A168) );
 a100091a <=( a100090a  and  a100087a );
 a100094a <=( (not A199)  and  A166 );
 a100097a <=( (not A201)  and  A200 );
 a100098a <=( a100097a  and  a100094a );
 a100099a <=( a100098a  and  a100091a );
 a100102a <=( (not A203)  and  (not A202) );
 a100105a <=( A266  and  (not A265) );
 a100106a <=( a100105a  and  a100102a );
 a100109a <=( A269  and  A267 );
 a100113a <=( (not A302)  and  (not A301) );
 a100114a <=( A300  and  a100113a );
 a100115a <=( a100114a  and  a100109a );
 a100116a <=( a100115a  and  a100106a );
 a100119a <=( (not A169)  and  A170 );
 a100122a <=( (not A167)  and  (not A168) );
 a100123a <=( a100122a  and  a100119a );
 a100126a <=( (not A199)  and  A166 );
 a100129a <=( (not A201)  and  A200 );
 a100130a <=( a100129a  and  a100126a );
 a100131a <=( a100130a  and  a100123a );
 a100134a <=( (not A203)  and  (not A202) );
 a100137a <=( A266  and  (not A265) );
 a100138a <=( a100137a  and  a100134a );
 a100141a <=( (not A268)  and  (not A267) );
 a100145a <=( A301  and  (not A300) );
 a100146a <=( (not A269)  and  a100145a );
 a100147a <=( a100146a  and  a100141a );
 a100148a <=( a100147a  and  a100138a );
 a100151a <=( (not A169)  and  A170 );
 a100154a <=( (not A167)  and  (not A168) );
 a100155a <=( a100154a  and  a100151a );
 a100158a <=( (not A199)  and  A166 );
 a100161a <=( (not A201)  and  A200 );
 a100162a <=( a100161a  and  a100158a );
 a100163a <=( a100162a  and  a100155a );
 a100166a <=( (not A203)  and  (not A202) );
 a100169a <=( A266  and  (not A265) );
 a100170a <=( a100169a  and  a100166a );
 a100173a <=( (not A268)  and  (not A267) );
 a100177a <=( A302  and  (not A300) );
 a100178a <=( (not A269)  and  a100177a );
 a100179a <=( a100178a  and  a100173a );
 a100180a <=( a100179a  and  a100170a );
 a100183a <=( (not A169)  and  A170 );
 a100186a <=( (not A167)  and  (not A168) );
 a100187a <=( a100186a  and  a100183a );
 a100190a <=( (not A199)  and  A166 );
 a100193a <=( (not A201)  and  A200 );
 a100194a <=( a100193a  and  a100190a );
 a100195a <=( a100194a  and  a100187a );
 a100198a <=( (not A203)  and  (not A202) );
 a100201a <=( A266  and  (not A265) );
 a100202a <=( a100201a  and  a100198a );
 a100205a <=( (not A268)  and  (not A267) );
 a100209a <=( A299  and  A298 );
 a100210a <=( (not A269)  and  a100209a );
 a100211a <=( a100210a  and  a100205a );
 a100212a <=( a100211a  and  a100202a );
 a100215a <=( (not A169)  and  A170 );
 a100218a <=( (not A167)  and  (not A168) );
 a100219a <=( a100218a  and  a100215a );
 a100222a <=( (not A199)  and  A166 );
 a100225a <=( (not A201)  and  A200 );
 a100226a <=( a100225a  and  a100222a );
 a100227a <=( a100226a  and  a100219a );
 a100230a <=( (not A203)  and  (not A202) );
 a100233a <=( A266  and  (not A265) );
 a100234a <=( a100233a  and  a100230a );
 a100237a <=( (not A268)  and  (not A267) );
 a100241a <=( (not A299)  and  (not A298) );
 a100242a <=( (not A269)  and  a100241a );
 a100243a <=( a100242a  and  a100237a );
 a100244a <=( a100243a  and  a100234a );
 a100247a <=( (not A169)  and  A170 );
 a100250a <=( (not A167)  and  (not A168) );
 a100251a <=( a100250a  and  a100247a );
 a100254a <=( (not A199)  and  A166 );
 a100257a <=( (not A201)  and  A200 );
 a100258a <=( a100257a  and  a100254a );
 a100259a <=( a100258a  and  a100251a );
 a100262a <=( (not A203)  and  (not A202) );
 a100265a <=( (not A266)  and  A265 );
 a100266a <=( a100265a  and  a100262a );
 a100269a <=( A268  and  A267 );
 a100273a <=( (not A302)  and  (not A301) );
 a100274a <=( A300  and  a100273a );
 a100275a <=( a100274a  and  a100269a );
 a100276a <=( a100275a  and  a100266a );
 a100279a <=( (not A169)  and  A170 );
 a100282a <=( (not A167)  and  (not A168) );
 a100283a <=( a100282a  and  a100279a );
 a100286a <=( (not A199)  and  A166 );
 a100289a <=( (not A201)  and  A200 );
 a100290a <=( a100289a  and  a100286a );
 a100291a <=( a100290a  and  a100283a );
 a100294a <=( (not A203)  and  (not A202) );
 a100297a <=( (not A266)  and  A265 );
 a100298a <=( a100297a  and  a100294a );
 a100301a <=( A269  and  A267 );
 a100305a <=( (not A302)  and  (not A301) );
 a100306a <=( A300  and  a100305a );
 a100307a <=( a100306a  and  a100301a );
 a100308a <=( a100307a  and  a100298a );
 a100311a <=( (not A169)  and  A170 );
 a100314a <=( (not A167)  and  (not A168) );
 a100315a <=( a100314a  and  a100311a );
 a100318a <=( (not A199)  and  A166 );
 a100321a <=( (not A201)  and  A200 );
 a100322a <=( a100321a  and  a100318a );
 a100323a <=( a100322a  and  a100315a );
 a100326a <=( (not A203)  and  (not A202) );
 a100329a <=( (not A266)  and  A265 );
 a100330a <=( a100329a  and  a100326a );
 a100333a <=( (not A268)  and  (not A267) );
 a100337a <=( A301  and  (not A300) );
 a100338a <=( (not A269)  and  a100337a );
 a100339a <=( a100338a  and  a100333a );
 a100340a <=( a100339a  and  a100330a );
 a100343a <=( (not A169)  and  A170 );
 a100346a <=( (not A167)  and  (not A168) );
 a100347a <=( a100346a  and  a100343a );
 a100350a <=( (not A199)  and  A166 );
 a100353a <=( (not A201)  and  A200 );
 a100354a <=( a100353a  and  a100350a );
 a100355a <=( a100354a  and  a100347a );
 a100358a <=( (not A203)  and  (not A202) );
 a100361a <=( (not A266)  and  A265 );
 a100362a <=( a100361a  and  a100358a );
 a100365a <=( (not A268)  and  (not A267) );
 a100369a <=( A302  and  (not A300) );
 a100370a <=( (not A269)  and  a100369a );
 a100371a <=( a100370a  and  a100365a );
 a100372a <=( a100371a  and  a100362a );
 a100375a <=( (not A169)  and  A170 );
 a100378a <=( (not A167)  and  (not A168) );
 a100379a <=( a100378a  and  a100375a );
 a100382a <=( (not A199)  and  A166 );
 a100385a <=( (not A201)  and  A200 );
 a100386a <=( a100385a  and  a100382a );
 a100387a <=( a100386a  and  a100379a );
 a100390a <=( (not A203)  and  (not A202) );
 a100393a <=( (not A266)  and  A265 );
 a100394a <=( a100393a  and  a100390a );
 a100397a <=( (not A268)  and  (not A267) );
 a100401a <=( A299  and  A298 );
 a100402a <=( (not A269)  and  a100401a );
 a100403a <=( a100402a  and  a100397a );
 a100404a <=( a100403a  and  a100394a );
 a100407a <=( (not A169)  and  A170 );
 a100410a <=( (not A167)  and  (not A168) );
 a100411a <=( a100410a  and  a100407a );
 a100414a <=( (not A199)  and  A166 );
 a100417a <=( (not A201)  and  A200 );
 a100418a <=( a100417a  and  a100414a );
 a100419a <=( a100418a  and  a100411a );
 a100422a <=( (not A203)  and  (not A202) );
 a100425a <=( (not A266)  and  A265 );
 a100426a <=( a100425a  and  a100422a );
 a100429a <=( (not A268)  and  (not A267) );
 a100433a <=( (not A299)  and  (not A298) );
 a100434a <=( (not A269)  and  a100433a );
 a100435a <=( a100434a  and  a100429a );
 a100436a <=( a100435a  and  a100426a );
 a100439a <=( (not A169)  and  A170 );
 a100442a <=( (not A167)  and  (not A168) );
 a100443a <=( a100442a  and  a100439a );
 a100446a <=( A199  and  A166 );
 a100449a <=( A201  and  (not A200) );
 a100450a <=( a100449a  and  a100446a );
 a100451a <=( a100450a  and  a100443a );
 a100454a <=( (not A265)  and  A202 );
 a100457a <=( (not A267)  and  A266 );
 a100458a <=( a100457a  and  a100454a );
 a100461a <=( (not A269)  and  (not A268) );
 a100465a <=( (not A302)  and  (not A301) );
 a100466a <=( A300  and  a100465a );
 a100467a <=( a100466a  and  a100461a );
 a100468a <=( a100467a  and  a100458a );
 a100471a <=( (not A169)  and  A170 );
 a100474a <=( (not A167)  and  (not A168) );
 a100475a <=( a100474a  and  a100471a );
 a100478a <=( A199  and  A166 );
 a100481a <=( A201  and  (not A200) );
 a100482a <=( a100481a  and  a100478a );
 a100483a <=( a100482a  and  a100475a );
 a100486a <=( A265  and  A202 );
 a100489a <=( (not A267)  and  (not A266) );
 a100490a <=( a100489a  and  a100486a );
 a100493a <=( (not A269)  and  (not A268) );
 a100497a <=( (not A302)  and  (not A301) );
 a100498a <=( A300  and  a100497a );
 a100499a <=( a100498a  and  a100493a );
 a100500a <=( a100499a  and  a100490a );
 a100503a <=( (not A169)  and  A170 );
 a100506a <=( (not A167)  and  (not A168) );
 a100507a <=( a100506a  and  a100503a );
 a100510a <=( A199  and  A166 );
 a100513a <=( A201  and  (not A200) );
 a100514a <=( a100513a  and  a100510a );
 a100515a <=( a100514a  and  a100507a );
 a100518a <=( (not A265)  and  A203 );
 a100521a <=( (not A267)  and  A266 );
 a100522a <=( a100521a  and  a100518a );
 a100525a <=( (not A269)  and  (not A268) );
 a100529a <=( (not A302)  and  (not A301) );
 a100530a <=( A300  and  a100529a );
 a100531a <=( a100530a  and  a100525a );
 a100532a <=( a100531a  and  a100522a );
 a100535a <=( (not A169)  and  A170 );
 a100538a <=( (not A167)  and  (not A168) );
 a100539a <=( a100538a  and  a100535a );
 a100542a <=( A199  and  A166 );
 a100545a <=( A201  and  (not A200) );
 a100546a <=( a100545a  and  a100542a );
 a100547a <=( a100546a  and  a100539a );
 a100550a <=( A265  and  A203 );
 a100553a <=( (not A267)  and  (not A266) );
 a100554a <=( a100553a  and  a100550a );
 a100557a <=( (not A269)  and  (not A268) );
 a100561a <=( (not A302)  and  (not A301) );
 a100562a <=( A300  and  a100561a );
 a100563a <=( a100562a  and  a100557a );
 a100564a <=( a100563a  and  a100554a );
 a100567a <=( (not A169)  and  A170 );
 a100570a <=( (not A167)  and  (not A168) );
 a100571a <=( a100570a  and  a100567a );
 a100574a <=( A199  and  A166 );
 a100577a <=( (not A201)  and  (not A200) );
 a100578a <=( a100577a  and  a100574a );
 a100579a <=( a100578a  and  a100571a );
 a100582a <=( (not A203)  and  (not A202) );
 a100585a <=( A266  and  (not A265) );
 a100586a <=( a100585a  and  a100582a );
 a100589a <=( A268  and  A267 );
 a100593a <=( (not A302)  and  (not A301) );
 a100594a <=( A300  and  a100593a );
 a100595a <=( a100594a  and  a100589a );
 a100596a <=( a100595a  and  a100586a );
 a100599a <=( (not A169)  and  A170 );
 a100602a <=( (not A167)  and  (not A168) );
 a100603a <=( a100602a  and  a100599a );
 a100606a <=( A199  and  A166 );
 a100609a <=( (not A201)  and  (not A200) );
 a100610a <=( a100609a  and  a100606a );
 a100611a <=( a100610a  and  a100603a );
 a100614a <=( (not A203)  and  (not A202) );
 a100617a <=( A266  and  (not A265) );
 a100618a <=( a100617a  and  a100614a );
 a100621a <=( A269  and  A267 );
 a100625a <=( (not A302)  and  (not A301) );
 a100626a <=( A300  and  a100625a );
 a100627a <=( a100626a  and  a100621a );
 a100628a <=( a100627a  and  a100618a );
 a100631a <=( (not A169)  and  A170 );
 a100634a <=( (not A167)  and  (not A168) );
 a100635a <=( a100634a  and  a100631a );
 a100638a <=( A199  and  A166 );
 a100641a <=( (not A201)  and  (not A200) );
 a100642a <=( a100641a  and  a100638a );
 a100643a <=( a100642a  and  a100635a );
 a100646a <=( (not A203)  and  (not A202) );
 a100649a <=( A266  and  (not A265) );
 a100650a <=( a100649a  and  a100646a );
 a100653a <=( (not A268)  and  (not A267) );
 a100657a <=( A301  and  (not A300) );
 a100658a <=( (not A269)  and  a100657a );
 a100659a <=( a100658a  and  a100653a );
 a100660a <=( a100659a  and  a100650a );
 a100663a <=( (not A169)  and  A170 );
 a100666a <=( (not A167)  and  (not A168) );
 a100667a <=( a100666a  and  a100663a );
 a100670a <=( A199  and  A166 );
 a100673a <=( (not A201)  and  (not A200) );
 a100674a <=( a100673a  and  a100670a );
 a100675a <=( a100674a  and  a100667a );
 a100678a <=( (not A203)  and  (not A202) );
 a100681a <=( A266  and  (not A265) );
 a100682a <=( a100681a  and  a100678a );
 a100685a <=( (not A268)  and  (not A267) );
 a100689a <=( A302  and  (not A300) );
 a100690a <=( (not A269)  and  a100689a );
 a100691a <=( a100690a  and  a100685a );
 a100692a <=( a100691a  and  a100682a );
 a100695a <=( (not A169)  and  A170 );
 a100698a <=( (not A167)  and  (not A168) );
 a100699a <=( a100698a  and  a100695a );
 a100702a <=( A199  and  A166 );
 a100705a <=( (not A201)  and  (not A200) );
 a100706a <=( a100705a  and  a100702a );
 a100707a <=( a100706a  and  a100699a );
 a100710a <=( (not A203)  and  (not A202) );
 a100713a <=( A266  and  (not A265) );
 a100714a <=( a100713a  and  a100710a );
 a100717a <=( (not A268)  and  (not A267) );
 a100721a <=( A299  and  A298 );
 a100722a <=( (not A269)  and  a100721a );
 a100723a <=( a100722a  and  a100717a );
 a100724a <=( a100723a  and  a100714a );
 a100727a <=( (not A169)  and  A170 );
 a100730a <=( (not A167)  and  (not A168) );
 a100731a <=( a100730a  and  a100727a );
 a100734a <=( A199  and  A166 );
 a100737a <=( (not A201)  and  (not A200) );
 a100738a <=( a100737a  and  a100734a );
 a100739a <=( a100738a  and  a100731a );
 a100742a <=( (not A203)  and  (not A202) );
 a100745a <=( A266  and  (not A265) );
 a100746a <=( a100745a  and  a100742a );
 a100749a <=( (not A268)  and  (not A267) );
 a100753a <=( (not A299)  and  (not A298) );
 a100754a <=( (not A269)  and  a100753a );
 a100755a <=( a100754a  and  a100749a );
 a100756a <=( a100755a  and  a100746a );
 a100759a <=( (not A169)  and  A170 );
 a100762a <=( (not A167)  and  (not A168) );
 a100763a <=( a100762a  and  a100759a );
 a100766a <=( A199  and  A166 );
 a100769a <=( (not A201)  and  (not A200) );
 a100770a <=( a100769a  and  a100766a );
 a100771a <=( a100770a  and  a100763a );
 a100774a <=( (not A203)  and  (not A202) );
 a100777a <=( (not A266)  and  A265 );
 a100778a <=( a100777a  and  a100774a );
 a100781a <=( A268  and  A267 );
 a100785a <=( (not A302)  and  (not A301) );
 a100786a <=( A300  and  a100785a );
 a100787a <=( a100786a  and  a100781a );
 a100788a <=( a100787a  and  a100778a );
 a100791a <=( (not A169)  and  A170 );
 a100794a <=( (not A167)  and  (not A168) );
 a100795a <=( a100794a  and  a100791a );
 a100798a <=( A199  and  A166 );
 a100801a <=( (not A201)  and  (not A200) );
 a100802a <=( a100801a  and  a100798a );
 a100803a <=( a100802a  and  a100795a );
 a100806a <=( (not A203)  and  (not A202) );
 a100809a <=( (not A266)  and  A265 );
 a100810a <=( a100809a  and  a100806a );
 a100813a <=( A269  and  A267 );
 a100817a <=( (not A302)  and  (not A301) );
 a100818a <=( A300  and  a100817a );
 a100819a <=( a100818a  and  a100813a );
 a100820a <=( a100819a  and  a100810a );
 a100823a <=( (not A169)  and  A170 );
 a100826a <=( (not A167)  and  (not A168) );
 a100827a <=( a100826a  and  a100823a );
 a100830a <=( A199  and  A166 );
 a100833a <=( (not A201)  and  (not A200) );
 a100834a <=( a100833a  and  a100830a );
 a100835a <=( a100834a  and  a100827a );
 a100838a <=( (not A203)  and  (not A202) );
 a100841a <=( (not A266)  and  A265 );
 a100842a <=( a100841a  and  a100838a );
 a100845a <=( (not A268)  and  (not A267) );
 a100849a <=( A301  and  (not A300) );
 a100850a <=( (not A269)  and  a100849a );
 a100851a <=( a100850a  and  a100845a );
 a100852a <=( a100851a  and  a100842a );
 a100855a <=( (not A169)  and  A170 );
 a100858a <=( (not A167)  and  (not A168) );
 a100859a <=( a100858a  and  a100855a );
 a100862a <=( A199  and  A166 );
 a100865a <=( (not A201)  and  (not A200) );
 a100866a <=( a100865a  and  a100862a );
 a100867a <=( a100866a  and  a100859a );
 a100870a <=( (not A203)  and  (not A202) );
 a100873a <=( (not A266)  and  A265 );
 a100874a <=( a100873a  and  a100870a );
 a100877a <=( (not A268)  and  (not A267) );
 a100881a <=( A302  and  (not A300) );
 a100882a <=( (not A269)  and  a100881a );
 a100883a <=( a100882a  and  a100877a );
 a100884a <=( a100883a  and  a100874a );
 a100887a <=( (not A169)  and  A170 );
 a100890a <=( (not A167)  and  (not A168) );
 a100891a <=( a100890a  and  a100887a );
 a100894a <=( A199  and  A166 );
 a100897a <=( (not A201)  and  (not A200) );
 a100898a <=( a100897a  and  a100894a );
 a100899a <=( a100898a  and  a100891a );
 a100902a <=( (not A203)  and  (not A202) );
 a100905a <=( (not A266)  and  A265 );
 a100906a <=( a100905a  and  a100902a );
 a100909a <=( (not A268)  and  (not A267) );
 a100913a <=( A299  and  A298 );
 a100914a <=( (not A269)  and  a100913a );
 a100915a <=( a100914a  and  a100909a );
 a100916a <=( a100915a  and  a100906a );
 a100919a <=( (not A169)  and  A170 );
 a100922a <=( (not A167)  and  (not A168) );
 a100923a <=( a100922a  and  a100919a );
 a100926a <=( A199  and  A166 );
 a100929a <=( (not A201)  and  (not A200) );
 a100930a <=( a100929a  and  a100926a );
 a100931a <=( a100930a  and  a100923a );
 a100934a <=( (not A203)  and  (not A202) );
 a100937a <=( (not A266)  and  A265 );
 a100938a <=( a100937a  and  a100934a );
 a100941a <=( (not A268)  and  (not A267) );
 a100945a <=( (not A299)  and  (not A298) );
 a100946a <=( (not A269)  and  a100945a );
 a100947a <=( a100946a  and  a100941a );
 a100948a <=( a100947a  and  a100938a );
 a100951a <=( (not A169)  and  A170 );
 a100954a <=( A167  and  (not A168) );
 a100955a <=( a100954a  and  a100951a );
 a100958a <=( (not A199)  and  (not A166) );
 a100962a <=( (not A202)  and  (not A201) );
 a100963a <=( A200  and  a100962a );
 a100964a <=( a100963a  and  a100958a );
 a100965a <=( a100964a  and  a100955a );
 a100968a <=( (not A265)  and  (not A203) );
 a100971a <=( (not A267)  and  A266 );
 a100972a <=( a100971a  and  a100968a );
 a100975a <=( (not A269)  and  (not A268) );
 a100979a <=( (not A302)  and  (not A301) );
 a100980a <=( A300  and  a100979a );
 a100981a <=( a100980a  and  a100975a );
 a100982a <=( a100981a  and  a100972a );
 a100985a <=( (not A169)  and  A170 );
 a100988a <=( A167  and  (not A168) );
 a100989a <=( a100988a  and  a100985a );
 a100992a <=( (not A199)  and  (not A166) );
 a100996a <=( (not A202)  and  (not A201) );
 a100997a <=( A200  and  a100996a );
 a100998a <=( a100997a  and  a100992a );
 a100999a <=( a100998a  and  a100989a );
 a101002a <=( A265  and  (not A203) );
 a101005a <=( (not A267)  and  (not A266) );
 a101006a <=( a101005a  and  a101002a );
 a101009a <=( (not A269)  and  (not A268) );
 a101013a <=( (not A302)  and  (not A301) );
 a101014a <=( A300  and  a101013a );
 a101015a <=( a101014a  and  a101009a );
 a101016a <=( a101015a  and  a101006a );
 a101019a <=( (not A169)  and  A170 );
 a101022a <=( A167  and  (not A168) );
 a101023a <=( a101022a  and  a101019a );
 a101026a <=( A199  and  (not A166) );
 a101030a <=( (not A202)  and  (not A201) );
 a101031a <=( (not A200)  and  a101030a );
 a101032a <=( a101031a  and  a101026a );
 a101033a <=( a101032a  and  a101023a );
 a101036a <=( (not A265)  and  (not A203) );
 a101039a <=( (not A267)  and  A266 );
 a101040a <=( a101039a  and  a101036a );
 a101043a <=( (not A269)  and  (not A268) );
 a101047a <=( (not A302)  and  (not A301) );
 a101048a <=( A300  and  a101047a );
 a101049a <=( a101048a  and  a101043a );
 a101050a <=( a101049a  and  a101040a );
 a101053a <=( (not A169)  and  A170 );
 a101056a <=( A167  and  (not A168) );
 a101057a <=( a101056a  and  a101053a );
 a101060a <=( A199  and  (not A166) );
 a101064a <=( (not A202)  and  (not A201) );
 a101065a <=( (not A200)  and  a101064a );
 a101066a <=( a101065a  and  a101060a );
 a101067a <=( a101066a  and  a101057a );
 a101070a <=( A265  and  (not A203) );
 a101073a <=( (not A267)  and  (not A266) );
 a101074a <=( a101073a  and  a101070a );
 a101077a <=( (not A269)  and  (not A268) );
 a101081a <=( (not A302)  and  (not A301) );
 a101082a <=( A300  and  a101081a );
 a101083a <=( a101082a  and  a101077a );
 a101084a <=( a101083a  and  a101074a );
 a101087a <=( (not A169)  and  A170 );
 a101090a <=( (not A167)  and  (not A168) );
 a101091a <=( a101090a  and  a101087a );
 a101094a <=( (not A199)  and  A166 );
 a101098a <=( (not A202)  and  (not A201) );
 a101099a <=( A200  and  a101098a );
 a101100a <=( a101099a  and  a101094a );
 a101101a <=( a101100a  and  a101091a );
 a101104a <=( (not A265)  and  (not A203) );
 a101107a <=( (not A267)  and  A266 );
 a101108a <=( a101107a  and  a101104a );
 a101111a <=( (not A269)  and  (not A268) );
 a101115a <=( (not A302)  and  (not A301) );
 a101116a <=( A300  and  a101115a );
 a101117a <=( a101116a  and  a101111a );
 a101118a <=( a101117a  and  a101108a );
 a101121a <=( (not A169)  and  A170 );
 a101124a <=( (not A167)  and  (not A168) );
 a101125a <=( a101124a  and  a101121a );
 a101128a <=( (not A199)  and  A166 );
 a101132a <=( (not A202)  and  (not A201) );
 a101133a <=( A200  and  a101132a );
 a101134a <=( a101133a  and  a101128a );
 a101135a <=( a101134a  and  a101125a );
 a101138a <=( A265  and  (not A203) );
 a101141a <=( (not A267)  and  (not A266) );
 a101142a <=( a101141a  and  a101138a );
 a101145a <=( (not A269)  and  (not A268) );
 a101149a <=( (not A302)  and  (not A301) );
 a101150a <=( A300  and  a101149a );
 a101151a <=( a101150a  and  a101145a );
 a101152a <=( a101151a  and  a101142a );
 a101155a <=( (not A169)  and  A170 );
 a101158a <=( (not A167)  and  (not A168) );
 a101159a <=( a101158a  and  a101155a );
 a101162a <=( A199  and  A166 );
 a101166a <=( (not A202)  and  (not A201) );
 a101167a <=( (not A200)  and  a101166a );
 a101168a <=( a101167a  and  a101162a );
 a101169a <=( a101168a  and  a101159a );
 a101172a <=( (not A265)  and  (not A203) );
 a101175a <=( (not A267)  and  A266 );
 a101176a <=( a101175a  and  a101172a );
 a101179a <=( (not A269)  and  (not A268) );
 a101183a <=( (not A302)  and  (not A301) );
 a101184a <=( A300  and  a101183a );
 a101185a <=( a101184a  and  a101179a );
 a101186a <=( a101185a  and  a101176a );
 a101189a <=( (not A169)  and  A170 );
 a101192a <=( (not A167)  and  (not A168) );
 a101193a <=( a101192a  and  a101189a );
 a101196a <=( A199  and  A166 );
 a101200a <=( (not A202)  and  (not A201) );
 a101201a <=( (not A200)  and  a101200a );
 a101202a <=( a101201a  and  a101196a );
 a101203a <=( a101202a  and  a101193a );
 a101206a <=( A265  and  (not A203) );
 a101209a <=( (not A267)  and  (not A266) );
 a101210a <=( a101209a  and  a101206a );
 a101213a <=( (not A269)  and  (not A268) );
 a101217a <=( (not A302)  and  (not A301) );
 a101218a <=( A300  and  a101217a );
 a101219a <=( a101218a  and  a101213a );
 a101220a <=( a101219a  and  a101210a );


end x25_4x_behav;
