Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_2x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A141: buffer std_logic
);
end x25_2x;

architecture x25_2x_behav of x25_2x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2193a,a2196a,a2197a,a2200a,a2203a,a2204a,a2205a,a2208a,a2211a,a2212a,a2215a,a2219a,a2220a,a2221a,a2222a,a2223a,a2226a,a2229a,a2230a,a2233a,a2236a,a2237a,a2238a,a2241a,a2244a,a2245a,a2248a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2260a,a2263a,a2264a,a2267a,a2270a,a2271a,a2272a,a2275a,a2278a,a2279a,a2282a,a2286a,a2287a,a2288a,a2289a,a2290a,a2293a,a2296a,a2297a,a2300a,a2303a,a2304a,a2305a,a2308a,a2311a,a2312a,a2315a,a2319a,a2320a,a2321a,a2322a,a2323a,a2324a,a2325a,a2328a,a2331a,a2332a,a2335a,a2338a,a2339a,a2340a,a2343a,a2346a,a2347a,a2350a,a2354a,a2355a,a2356a,a2357a,a2358a,a2361a,a2364a,a2365a,a2368a,a2371a,a2372a,a2373a,a2376a,a2379a,a2380a,a2383a,a2387a,a2388a,a2389a,a2390a,a2391a,a2392a,a2395a,a2398a,a2399a,a2402a,a2405a,a2406a,a2407a,a2410a,a2413a,a2414a,a2417a,a2421a,a2422a,a2423a,a2424a,a2425a,a2428a,a2431a,a2432a,a2435a,a2438a,a2439a,a2440a,a2443a,a2446a,a2447a,a2450a,a2454a,a2455a,a2456a,a2457a,a2458a,a2459a,a2460a,a2461a,a2464a,a2467a,a2468a,a2471a,a2474a,a2475a,a2476a,a2479a,a2482a,a2483a,a2486a,a2490a,a2491a,a2492a,a2493a,a2494a,a2497a,a2500a,a2501a,a2504a,a2507a,a2508a,a2509a,a2512a,a2515a,a2516a,a2519a,a2523a,a2524a,a2525a,a2526a,a2527a,a2528a,a2531a,a2534a,a2535a,a2538a,a2541a,a2542a,a2543a,a2546a,a2549a,a2550a,a2553a,a2557a,a2558a,a2559a,a2560a,a2561a,a2564a,a2567a,a2568a,a2571a,a2574a,a2575a,a2576a,a2579a,a2582a,a2583a,a2586a,a2590a,a2591a,a2592a,a2593a,a2594a,a2595a,a2596a,a2599a,a2602a,a2603a,a2606a,a2609a,a2610a,a2611a,a2614a,a2617a,a2618a,a2621a,a2625a,a2626a,a2627a,a2628a,a2629a,a2632a,a2635a,a2636a,a2639a,a2642a,a2643a,a2644a,a2647a,a2650a,a2651a,a2654a,a2658a,a2659a,a2660a,a2661a,a2662a,a2663a,a2666a,a2669a,a2670a,a2673a,a2676a,a2677a,a2678a,a2681a,a2684a,a2685a,a2688a,a2692a,a2693a,a2694a,a2695a,a2696a,a2699a,a2702a,a2703a,a2706a,a2710a,a2711a,a2712a,a2713a,a2716a,a2719a,a2720a,a2723a,a2727a,a2728a,a2729a,a2730a,a2731a,a2732a,a2733a,a2734a,a2735a,a2738a,a2741a,a2742a,a2745a,a2748a,a2749a,a2750a,a2753a,a2756a,a2757a,a2760a,a2764a,a2765a,a2766a,a2767a,a2768a,a2771a,a2774a,a2775a,a2778a,a2781a,a2782a,a2783a,a2786a,a2789a,a2790a,a2793a,a2797a,a2798a,a2799a,a2800a,a2801a,a2802a,a2805a,a2808a,a2809a,a2812a,a2815a,a2816a,a2817a,a2820a,a2823a,a2824a,a2827a,a2831a,a2832a,a2833a,a2834a,a2835a,a2838a,a2841a,a2842a,a2845a,a2848a,a2849a,a2850a,a2853a,a2856a,a2857a,a2860a,a2864a,a2865a,a2866a,a2867a,a2868a,a2869a,a2870a,a2873a,a2876a,a2877a,a2880a,a2883a,a2884a,a2885a,a2888a,a2891a,a2892a,a2895a,a2899a,a2900a,a2901a,a2902a,a2903a,a2906a,a2909a,a2910a,a2913a,a2916a,a2917a,a2918a,a2921a,a2924a,a2925a,a2928a,a2932a,a2933a,a2934a,a2935a,a2936a,a2937a,a2940a,a2943a,a2944a,a2947a,a2950a,a2951a,a2952a,a2955a,a2958a,a2959a,a2962a,a2966a,a2967a,a2968a,a2969a,a2970a,a2973a,a2976a,a2977a,a2980a,a2984a,a2985a,a2986a,a2987a,a2990a,a2993a,a2994a,a2997a,a3001a,a3002a,a3003a,a3004a,a3005a,a3006a,a3007a,a3008a,a3011a,a3014a,a3015a,a3018a,a3021a,a3022a,a3023a,a3026a,a3029a,a3030a,a3033a,a3037a,a3038a,a3039a,a3040a,a3041a,a3044a,a3047a,a3048a,a3051a,a3054a,a3055a,a3056a,a3059a,a3062a,a3063a,a3066a,a3070a,a3071a,a3072a,a3073a,a3074a,a3075a,a3078a,a3081a,a3082a,a3085a,a3088a,a3089a,a3090a,a3093a,a3096a,a3097a,a3100a,a3104a,a3105a,a3106a,a3107a,a3108a,a3111a,a3114a,a3115a,a3118a,a3121a,a3122a,a3123a,a3126a,a3129a,a3130a,a3133a,a3137a,a3138a,a3139a,a3140a,a3141a,a3142a,a3143a,a3146a,a3149a,a3150a,a3153a,a3156a,a3157a,a3158a,a3161a,a3164a,a3165a,a3168a,a3172a,a3173a,a3174a,a3175a,a3176a,a3179a,a3182a,a3183a,a3186a,a3189a,a3190a,a3191a,a3194a,a3197a,a3198a,a3201a,a3205a,a3206a,a3207a,a3208a,a3209a,a3210a,a3213a,a3216a,a3217a,a3220a,a3223a,a3224a,a3225a,a3228a,a3231a,a3232a,a3235a,a3239a,a3240a,a3241a,a3242a,a3243a,a3246a,a3249a,a3250a,a3253a,a3257a,a3258a,a3259a,a3260a,a3263a,a3266a,a3267a,a3270a,a3274a,a3275a,a3276a,a3277a,a3278a,a3279a,a3280a,a3281a,a3282a,a3283a,a3286a,a3289a,a3290a,a3293a,a3296a,a3297a,a3298a,a3301a,a3304a,a3305a,a3308a,a3312a,a3313a,a3314a,a3315a,a3316a,a3319a,a3322a,a3323a,a3326a,a3329a,a3330a,a3331a,a3334a,a3337a,a3338a,a3341a,a3345a,a3346a,a3347a,a3348a,a3349a,a3350a,a3353a,a3356a,a3357a,a3360a,a3363a,a3364a,a3365a,a3368a,a3371a,a3372a,a3375a,a3379a,a3380a,a3381a,a3382a,a3383a,a3386a,a3389a,a3390a,a3393a,a3396a,a3397a,a3398a,a3401a,a3404a,a3405a,a3408a,a3412a,a3413a,a3414a,a3415a,a3416a,a3417a,a3418a,a3421a,a3424a,a3425a,a3428a,a3431a,a3432a,a3433a,a3436a,a3439a,a3440a,a3443a,a3447a,a3448a,a3449a,a3450a,a3451a,a3454a,a3457a,a3458a,a3461a,a3464a,a3465a,a3466a,a3469a,a3472a,a3473a,a3476a,a3480a,a3481a,a3482a,a3483a,a3484a,a3485a,a3488a,a3491a,a3492a,a3495a,a3498a,a3499a,a3500a,a3503a,a3506a,a3507a,a3510a,a3514a,a3515a,a3516a,a3517a,a3518a,a3521a,a3524a,a3525a,a3528a,a3532a,a3533a,a3534a,a3535a,a3538a,a3541a,a3542a,a3545a,a3549a,a3550a,a3551a,a3552a,a3553a,a3554a,a3555a,a3556a,a3559a,a3562a,a3563a,a3566a,a3569a,a3570a,a3571a,a3574a,a3577a,a3578a,a3581a,a3585a,a3586a,a3587a,a3588a,a3589a,a3592a,a3595a,a3596a,a3599a,a3602a,a3603a,a3604a,a3607a,a3610a,a3611a,a3614a,a3618a,a3619a,a3620a,a3621a,a3622a,a3623a,a3626a,a3629a,a3630a,a3633a,a3636a,a3637a,a3638a,a3641a,a3644a,a3645a,a3648a,a3652a,a3653a,a3654a,a3655a,a3656a,a3659a,a3662a,a3663a,a3666a,a3669a,a3670a,a3671a,a3674a,a3677a,a3678a,a3681a,a3685a,a3686a,a3687a,a3688a,a3689a,a3690a,a3691a,a3694a,a3697a,a3698a,a3701a,a3704a,a3705a,a3706a,a3709a,a3712a,a3713a,a3716a,a3720a,a3721a,a3722a,a3723a,a3724a,a3727a,a3730a,a3731a,a3734a,a3737a,a3738a,a3739a,a3742a,a3745a,a3746a,a3749a,a3753a,a3754a,a3755a,a3756a,a3757a,a3758a,a3761a,a3764a,a3765a,a3768a,a3771a,a3772a,a3773a,a3776a,a3779a,a3780a,a3783a,a3787a,a3788a,a3789a,a3790a,a3791a,a3794a,a3797a,a3798a,a3801a,a3805a,a3806a,a3807a,a3808a,a3811a,a3814a,a3815a,a3818a,a3822a,a3823a,a3824a,a3825a,a3826a,a3827a,a3828a,a3829a,a3830a,a3833a,a3836a,a3837a,a3840a,a3843a,a3844a,a3845a,a3848a,a3851a,a3852a,a3855a,a3859a,a3860a,a3861a,a3862a,a3863a,a3866a,a3869a,a3870a,a3873a,a3876a,a3877a,a3878a,a3881a,a3884a,a3885a,a3888a,a3892a,a3893a,a3894a,a3895a,a3896a,a3897a,a3900a,a3903a,a3904a,a3907a,a3910a,a3911a,a3912a,a3915a,a3918a,a3919a,a3922a,a3926a,a3927a,a3928a,a3929a,a3930a,a3933a,a3936a,a3937a,a3940a,a3943a,a3944a,a3945a,a3948a,a3951a,a3952a,a3955a,a3959a,a3960a,a3961a,a3962a,a3963a,a3964a,a3965a,a3968a,a3971a,a3972a,a3975a,a3978a,a3979a,a3980a,a3983a,a3986a,a3987a,a3990a,a3994a,a3995a,a3996a,a3997a,a3998a,a4001a,a4004a,a4005a,a4008a,a4011a,a4012a,a4013a,a4016a,a4019a,a4020a,a4023a,a4027a,a4028a,a4029a,a4030a,a4031a,a4032a,a4035a,a4038a,a4039a,a4042a,a4045a,a4046a,a4047a,a4050a,a4053a,a4054a,a4057a,a4061a,a4062a,a4063a,a4064a,a4065a,a4068a,a4071a,a4072a,a4075a,a4079a,a4080a,a4081a,a4082a,a4085a,a4088a,a4089a,a4092a,a4096a,a4097a,a4098a,a4099a,a4100a,a4101a,a4102a,a4103a,a4106a,a4109a,a4110a,a4113a,a4116a,a4117a,a4118a,a4121a,a4124a,a4125a,a4128a,a4132a,a4133a,a4134a,a4135a,a4136a,a4139a,a4142a,a4143a,a4146a,a4149a,a4150a,a4151a,a4154a,a4157a,a4158a,a4161a,a4165a,a4166a,a4167a,a4168a,a4169a,a4170a,a4173a,a4176a,a4177a,a4180a,a4183a,a4184a,a4185a,a4188a,a4191a,a4192a,a4195a,a4199a,a4200a,a4201a,a4202a,a4203a,a4206a,a4209a,a4210a,a4213a,a4216a,a4217a,a4218a,a4221a,a4224a,a4225a,a4228a,a4232a,a4233a,a4234a,a4235a,a4236a,a4237a,a4238a,a4241a,a4244a,a4245a,a4248a,a4251a,a4252a,a4253a,a4256a,a4259a,a4260a,a4263a,a4267a,a4268a,a4269a,a4270a,a4271a,a4274a,a4277a,a4278a,a4281a,a4284a,a4285a,a4286a,a4289a,a4292a,a4293a,a4296a,a4300a,a4301a,a4302a,a4303a,a4304a,a4305a,a4308a,a4311a,a4312a,a4315a,a4318a,a4319a,a4320a,a4323a,a4326a,a4327a,a4330a,a4334a,a4335a,a4336a,a4337a,a4338a,a4341a,a4344a,a4345a,a4348a,a4352a,a4353a,a4354a,a4355a,a4358a,a4361a,a4362a,a4365a,a4369a,a4370a,a4371a,a4372a,a4373a,a4374a,a4375a,a4376a,a4377a,a4378a,a4379a,a4382a,a4385a,a4386a,a4389a,a4392a,a4393a,a4394a,a4397a,a4400a,a4401a,a4404a,a4408a,a4409a,a4410a,a4411a,a4412a,a4415a,a4418a,a4419a,a4422a,a4425a,a4426a,a4427a,a4430a,a4433a,a4434a,a4437a,a4441a,a4442a,a4443a,a4444a,a4445a,a4446a,a4449a,a4452a,a4453a,a4456a,a4459a,a4460a,a4461a,a4464a,a4467a,a4468a,a4471a,a4475a,a4476a,a4477a,a4478a,a4479a,a4482a,a4485a,a4486a,a4489a,a4492a,a4493a,a4494a,a4497a,a4500a,a4501a,a4504a,a4508a,a4509a,a4510a,a4511a,a4512a,a4513a,a4514a,a4517a,a4520a,a4521a,a4524a,a4527a,a4528a,a4529a,a4532a,a4535a,a4536a,a4539a,a4543a,a4544a,a4545a,a4546a,a4547a,a4550a,a4553a,a4554a,a4557a,a4560a,a4561a,a4562a,a4565a,a4568a,a4569a,a4572a,a4576a,a4577a,a4578a,a4579a,a4580a,a4581a,a4584a,a4587a,a4588a,a4591a,a4594a,a4595a,a4596a,a4599a,a4602a,a4603a,a4606a,a4610a,a4611a,a4612a,a4613a,a4614a,a4617a,a4620a,a4621a,a4624a,a4627a,a4628a,a4629a,a4632a,a4635a,a4636a,a4639a,a4643a,a4644a,a4645a,a4646a,a4647a,a4648a,a4649a,a4650a,a4653a,a4656a,a4657a,a4660a,a4663a,a4664a,a4665a,a4668a,a4671a,a4672a,a4675a,a4679a,a4680a,a4681a,a4682a,a4683a,a4686a,a4689a,a4690a,a4693a,a4696a,a4697a,a4698a,a4701a,a4704a,a4705a,a4708a,a4712a,a4713a,a4714a,a4715a,a4716a,a4717a,a4720a,a4723a,a4724a,a4727a,a4730a,a4731a,a4732a,a4735a,a4738a,a4739a,a4742a,a4746a,a4747a,a4748a,a4749a,a4750a,a4753a,a4756a,a4757a,a4760a,a4763a,a4764a,a4765a,a4768a,a4771a,a4772a,a4775a,a4779a,a4780a,a4781a,a4782a,a4783a,a4784a,a4785a,a4788a,a4791a,a4792a,a4795a,a4798a,a4799a,a4800a,a4803a,a4806a,a4807a,a4810a,a4814a,a4815a,a4816a,a4817a,a4818a,a4821a,a4824a,a4825a,a4828a,a4831a,a4832a,a4833a,a4836a,a4839a,a4840a,a4843a,a4847a,a4848a,a4849a,a4850a,a4851a,a4852a,a4855a,a4858a,a4859a,a4862a,a4865a,a4866a,a4867a,a4870a,a4873a,a4874a,a4877a,a4881a,a4882a,a4883a,a4884a,a4885a,a4888a,a4891a,a4892a,a4895a,a4899a,a4900a,a4901a,a4902a,a4905a,a4908a,a4909a,a4912a,a4916a,a4917a,a4918a,a4919a,a4920a,a4921a,a4922a,a4923a,a4924a,a4927a,a4930a,a4931a,a4934a,a4937a,a4938a,a4939a,a4942a,a4945a,a4946a,a4949a,a4953a,a4954a,a4955a,a4956a,a4957a,a4960a,a4963a,a4964a,a4967a,a4970a,a4971a,a4972a,a4975a,a4978a,a4979a,a4982a,a4986a,a4987a,a4988a,a4989a,a4990a,a4991a,a4994a,a4997a,a4998a,a5001a,a5004a,a5005a,a5006a,a5009a,a5012a,a5013a,a5016a,a5020a,a5021a,a5022a,a5023a,a5024a,a5027a,a5030a,a5031a,a5034a,a5037a,a5038a,a5039a,a5042a,a5045a,a5046a,a5049a,a5053a,a5054a,a5055a,a5056a,a5057a,a5058a,a5059a,a5062a,a5065a,a5066a,a5069a,a5072a,a5073a,a5074a,a5077a,a5080a,a5081a,a5084a,a5088a,a5089a,a5090a,a5091a,a5092a,a5095a,a5098a,a5099a,a5102a,a5105a,a5106a,a5107a,a5110a,a5113a,a5114a,a5117a,a5121a,a5122a,a5123a,a5124a,a5125a,a5126a,a5129a,a5132a,a5133a,a5136a,a5139a,a5140a,a5141a,a5144a,a5147a,a5148a,a5151a,a5155a,a5156a,a5157a,a5158a,a5159a,a5162a,a5165a,a5166a,a5169a,a5173a,a5174a,a5175a,a5176a,a5179a,a5182a,a5183a,a5186a,a5190a,a5191a,a5192a,a5193a,a5194a,a5195a,a5196a,a5197a,a5200a,a5203a,a5204a,a5207a,a5210a,a5211a,a5212a,a5215a,a5218a,a5219a,a5222a,a5226a,a5227a,a5228a,a5229a,a5230a,a5233a,a5236a,a5237a,a5240a,a5243a,a5244a,a5245a,a5248a,a5251a,a5252a,a5255a,a5259a,a5260a,a5261a,a5262a,a5263a,a5264a,a5267a,a5270a,a5271a,a5274a,a5277a,a5278a,a5279a,a5282a,a5285a,a5286a,a5289a,a5293a,a5294a,a5295a,a5296a,a5297a,a5300a,a5303a,a5304a,a5307a,a5310a,a5311a,a5312a,a5315a,a5318a,a5319a,a5322a,a5326a,a5327a,a5328a,a5329a,a5330a,a5331a,a5332a,a5335a,a5338a,a5339a,a5342a,a5345a,a5346a,a5347a,a5350a,a5353a,a5354a,a5357a,a5361a,a5362a,a5363a,a5364a,a5365a,a5368a,a5371a,a5372a,a5375a,a5378a,a5379a,a5380a,a5383a,a5386a,a5387a,a5390a,a5394a,a5395a,a5396a,a5397a,a5398a,a5399a,a5402a,a5405a,a5406a,a5409a,a5412a,a5413a,a5414a,a5417a,a5420a,a5421a,a5424a,a5428a,a5429a,a5430a,a5431a,a5432a,a5435a,a5438a,a5439a,a5442a,a5446a,a5447a,a5448a,a5449a,a5452a,a5455a,a5456a,a5459a,a5463a,a5464a,a5465a,a5466a,a5467a,a5468a,a5469a,a5470a,a5471a,a5472a,a5475a,a5478a,a5479a,a5482a,a5485a,a5486a,a5487a,a5490a,a5493a,a5494a,a5497a,a5501a,a5502a,a5503a,a5504a,a5505a,a5508a,a5511a,a5512a,a5515a,a5518a,a5519a,a5520a,a5523a,a5526a,a5527a,a5530a,a5534a,a5535a,a5536a,a5537a,a5538a,a5539a,a5542a,a5545a,a5546a,a5549a,a5552a,a5553a,a5554a,a5557a,a5560a,a5561a,a5564a,a5568a,a5569a,a5570a,a5571a,a5572a,a5575a,a5578a,a5579a,a5582a,a5585a,a5586a,a5587a,a5590a,a5593a,a5594a,a5597a,a5601a,a5602a,a5603a,a5604a,a5605a,a5606a,a5607a,a5610a,a5613a,a5614a,a5617a,a5620a,a5621a,a5622a,a5625a,a5628a,a5629a,a5632a,a5636a,a5637a,a5638a,a5639a,a5640a,a5643a,a5646a,a5647a,a5650a,a5653a,a5654a,a5655a,a5658a,a5661a,a5662a,a5665a,a5669a,a5670a,a5671a,a5672a,a5673a,a5674a,a5677a,a5680a,a5681a,a5684a,a5687a,a5688a,a5689a,a5692a,a5695a,a5696a,a5699a,a5703a,a5704a,a5705a,a5706a,a5707a,a5710a,a5713a,a5714a,a5717a,a5721a,a5722a,a5723a,a5724a,a5727a,a5730a,a5731a,a5734a,a5738a,a5739a,a5740a,a5741a,a5742a,a5743a,a5744a,a5745a,a5748a,a5751a,a5752a,a5755a,a5758a,a5759a,a5760a,a5763a,a5766a,a5767a,a5770a,a5774a,a5775a,a5776a,a5777a,a5778a,a5781a,a5784a,a5785a,a5788a,a5791a,a5792a,a5793a,a5796a,a5799a,a5800a,a5803a,a5807a,a5808a,a5809a,a5810a,a5811a,a5812a,a5815a,a5818a,a5819a,a5822a,a5825a,a5826a,a5827a,a5830a,a5833a,a5834a,a5837a,a5841a,a5842a,a5843a,a5844a,a5845a,a5848a,a5851a,a5852a,a5855a,a5858a,a5859a,a5860a,a5863a,a5866a,a5867a,a5870a,a5874a,a5875a,a5876a,a5877a,a5878a,a5879a,a5880a,a5883a,a5886a,a5887a,a5890a,a5893a,a5894a,a5895a,a5898a,a5901a,a5902a,a5905a,a5909a,a5910a,a5911a,a5912a,a5913a,a5916a,a5919a,a5920a,a5923a,a5926a,a5927a,a5928a,a5931a,a5934a,a5935a,a5938a,a5942a,a5943a,a5944a,a5945a,a5946a,a5947a,a5950a,a5953a,a5954a,a5957a,a5960a,a5961a,a5962a,a5965a,a5968a,a5969a,a5972a,a5976a,a5977a,a5978a,a5979a,a5980a,a5983a,a5986a,a5987a,a5990a,a5994a,a5995a,a5996a,a5997a,a6000a,a6003a,a6004a,a6007a,a6011a,a6012a,a6013a,a6014a,a6015a,a6016a,a6017a,a6018a,a6019a,a6022a,a6025a,a6026a,a6029a,a6032a,a6033a,a6034a,a6037a,a6040a,a6041a,a6044a,a6048a,a6049a,a6050a,a6051a,a6052a,a6055a,a6058a,a6059a,a6062a,a6065a,a6066a,a6067a,a6070a,a6073a,a6074a,a6077a,a6081a,a6082a,a6083a,a6084a,a6085a,a6086a,a6089a,a6092a,a6093a,a6096a,a6099a,a6100a,a6101a,a6104a,a6107a,a6108a,a6111a,a6115a,a6116a,a6117a,a6118a,a6119a,a6122a,a6125a,a6126a,a6129a,a6132a,a6133a,a6134a,a6137a,a6140a,a6141a,a6144a,a6148a,a6149a,a6150a,a6151a,a6152a,a6153a,a6154a,a6157a,a6160a,a6161a,a6164a,a6167a,a6168a,a6169a,a6172a,a6175a,a6176a,a6179a,a6183a,a6184a,a6185a,a6186a,a6187a,a6190a,a6193a,a6194a,a6197a,a6200a,a6201a,a6202a,a6205a,a6208a,a6209a,a6212a,a6216a,a6217a,a6218a,a6219a,a6220a,a6221a,a6224a,a6227a,a6228a,a6231a,a6234a,a6235a,a6236a,a6239a,a6242a,a6243a,a6246a,a6250a,a6251a,a6252a,a6253a,a6254a,a6257a,a6260a,a6261a,a6264a,a6268a,a6269a,a6270a,a6271a,a6274a,a6277a,a6278a,a6281a,a6285a,a6286a,a6287a,a6288a,a6289a,a6290a,a6291a,a6292a,a6295a,a6298a,a6299a,a6302a,a6305a,a6306a,a6307a,a6310a,a6313a,a6314a,a6317a,a6321a,a6322a,a6323a,a6324a,a6325a,a6328a,a6331a,a6332a,a6335a,a6338a,a6339a,a6340a,a6343a,a6346a,a6347a,a6350a,a6354a,a6355a,a6356a,a6357a,a6358a,a6359a,a6362a,a6365a,a6366a,a6369a,a6372a,a6373a,a6374a,a6377a,a6380a,a6381a,a6384a,a6388a,a6389a,a6390a,a6391a,a6392a,a6395a,a6398a,a6399a,a6402a,a6405a,a6406a,a6407a,a6410a,a6413a,a6414a,a6417a,a6421a,a6422a,a6423a,a6424a,a6425a,a6426a,a6427a,a6430a,a6433a,a6434a,a6437a,a6440a,a6441a,a6442a,a6445a,a6448a,a6449a,a6452a,a6456a,a6457a,a6458a,a6459a,a6460a,a6463a,a6466a,a6467a,a6470a,a6473a,a6474a,a6475a,a6478a,a6481a,a6482a,a6485a,a6489a,a6490a,a6491a,a6492a,a6493a,a6494a,a6497a,a6500a,a6501a,a6504a,a6507a,a6508a,a6509a,a6512a,a6515a,a6516a,a6519a,a6523a,a6524a,a6525a,a6526a,a6527a,a6530a,a6533a,a6534a,a6537a,a6541a,a6542a,a6543a,a6544a,a6547a,a6550a,a6551a,a6554a,a6558a,a6559a,a6560a,a6561a,a6562a,a6563a,a6564a,a6565a,a6566a,a6567a,a6568a,a6572a,a6573a,a6577a,a6578a,a6582a,a6583a,a6587a,a6588a,a6592a,a6593a,a6597a,a6598a,a6602a,a6603a,a6607a,a6608a,a6612a,a6613a,a6617a,a6618a,a6622a,a6623a,a6627a,a6628a,a6632a,a6633a,a6637a,a6638a,a6642a,a6643a,a6647a,a6648a,a6652a,a6653a,a6657a,a6658a,a6662a,a6663a,a6667a,a6668a,a6672a,a6673a,a6677a,a6678a,a6682a,a6683a,a6687a,a6688a,a6692a,a6693a,a6697a,a6698a,a6702a,a6703a,a6707a,a6708a,a6712a,a6713a,a6717a,a6718a,a6722a,a6723a,a6727a,a6728a,a6732a,a6733a,a6736a,a6739a,a6740a,a6744a,a6745a,a6748a,a6751a,a6752a,a6756a,a6757a,a6760a,a6763a,a6764a,a6768a,a6769a,a6772a,a6775a,a6776a,a6780a,a6781a,a6784a,a6787a,a6788a,a6792a,a6793a,a6796a,a6799a,a6800a,a6804a,a6805a,a6808a,a6811a,a6812a,a6816a,a6817a,a6820a,a6823a,a6824a,a6828a,a6829a,a6832a,a6835a,a6836a,a6840a,a6841a,a6844a,a6847a,a6848a,a6852a,a6853a,a6856a,a6859a,a6860a,a6864a,a6865a,a6868a,a6871a,a6872a,a6875a,a6878a,a6879a,a6882a,a6885a,a6886a,a6889a,a6892a,a6893a,a6896a,a6899a,a6900a,a6904a,a6905a,a6908a,a6911a,a6912a,a6913a,a6917a,a6918a,a6921a,a6924a,a6925a,a6926a,a6930a,a6931a,a6934a,a6937a,a6938a,a6939a,a6943a,a6944a,a6947a,a6950a,a6951a,a6952a,a6956a,a6957a,a6960a,a6963a,a6964a,a6965a,a6969a,a6970a,a6973a,a6976a,a6977a,a6978a,a6982a,a6983a,a6986a,a6989a,a6990a,a6991a,a6995a,a6996a,a6999a,a7002a,a7003a,a7004a,a7008a,a7009a,a7012a,a7015a,a7016a,a7017a,a7021a,a7022a,a7025a,a7028a,a7029a,a7030a,a7034a,a7035a,a7038a,a7041a,a7042a,a7043a,a7047a,a7048a,a7051a,a7054a,a7055a,a7056a,a7060a,a7061a,a7064a,a7067a,a7068a,a7069a,a7073a,a7074a,a7077a,a7080a,a7081a,a7082a,a7086a,a7087a,a7090a,a7093a,a7094a,a7095a,a7099a,a7100a,a7103a,a7106a,a7107a,a7108a,a7112a,a7113a,a7116a,a7119a,a7120a,a7121a,a7125a,a7126a,a7129a,a7132a,a7133a,a7134a,a7138a,a7139a,a7142a,a7145a,a7146a,a7147a,a7151a,a7152a,a7155a,a7158a,a7159a,a7160a,a7164a,a7165a,a7168a,a7171a,a7172a,a7173a,a7177a,a7178a,a7181a,a7184a,a7185a,a7186a,a7190a,a7191a,a7194a,a7197a,a7198a,a7199a,a7203a,a7204a,a7207a,a7210a,a7211a,a7212a,a7216a,a7217a,a7220a,a7223a,a7224a,a7225a,a7229a,a7230a,a7233a,a7236a,a7237a,a7238a,a7242a,a7243a,a7246a,a7249a,a7250a,a7251a,a7255a,a7256a,a7259a,a7262a,a7263a,a7264a,a7268a,a7269a,a7272a,a7275a,a7276a,a7277a,a7281a,a7282a,a7285a,a7288a,a7289a,a7290a,a7294a,a7295a,a7298a,a7301a,a7302a,a7303a,a7307a,a7308a,a7311a,a7314a,a7315a,a7316a,a7320a,a7321a,a7324a,a7327a,a7328a,a7329a,a7333a,a7334a,a7337a,a7340a,a7341a,a7342a,a7346a,a7347a,a7350a,a7353a,a7354a,a7355a,a7359a,a7360a,a7363a,a7366a,a7367a,a7368a,a7372a,a7373a,a7376a,a7379a,a7380a,a7381a,a7385a,a7386a,a7389a,a7392a,a7393a,a7394a,a7398a,a7399a,a7402a,a7405a,a7406a,a7407a,a7411a,a7412a,a7415a,a7418a,a7419a,a7420a,a7424a,a7425a,a7428a,a7431a,a7432a,a7433a,a7437a,a7438a,a7441a,a7444a,a7445a,a7446a,a7450a,a7451a,a7454a,a7457a,a7458a,a7459a,a7463a,a7464a,a7467a,a7470a,a7471a,a7472a,a7476a,a7477a,a7480a,a7483a,a7484a,a7485a,a7489a,a7490a,a7493a,a7496a,a7497a,a7498a,a7502a,a7503a,a7506a,a7509a,a7510a,a7511a,a7515a,a7516a,a7519a,a7522a,a7523a,a7524a,a7528a,a7529a,a7532a,a7535a,a7536a,a7537a,a7541a,a7542a,a7545a,a7548a,a7549a,a7550a,a7554a,a7555a,a7558a,a7561a,a7562a,a7563a,a7567a,a7568a,a7571a,a7574a,a7575a,a7576a,a7580a,a7581a,a7584a,a7587a,a7588a,a7589a,a7593a,a7594a,a7597a,a7600a,a7601a,a7602a,a7606a,a7607a,a7610a,a7613a,a7614a,a7615a,a7619a,a7620a,a7623a,a7626a,a7627a,a7628a,a7632a,a7633a,a7636a,a7639a,a7640a,a7641a,a7645a,a7646a,a7649a,a7652a,a7653a,a7654a,a7658a,a7659a,a7662a,a7665a,a7666a,a7667a,a7671a,a7672a,a7675a,a7678a,a7679a,a7680a,a7684a,a7685a,a7688a,a7691a,a7692a,a7693a,a7697a,a7698a,a7701a,a7704a,a7705a,a7706a,a7710a,a7711a,a7714a,a7717a,a7718a,a7719a,a7723a,a7724a,a7727a,a7730a,a7731a,a7732a,a7736a,a7737a,a7740a,a7743a,a7744a,a7745a,a7749a,a7750a,a7753a,a7756a,a7757a,a7758a,a7762a,a7763a,a7766a,a7769a,a7770a,a7771a,a7775a,a7776a,a7779a,a7782a,a7783a,a7784a,a7788a,a7789a,a7792a,a7795a,a7796a,a7797a,a7801a,a7802a,a7805a,a7808a,a7809a,a7810a,a7814a,a7815a,a7818a,a7821a,a7822a,a7823a,a7827a,a7828a,a7831a,a7834a,a7835a,a7836a,a7840a,a7841a,a7844a,a7847a,a7848a,a7849a,a7853a,a7854a,a7857a,a7860a,a7861a,a7862a,a7866a,a7867a,a7870a,a7873a,a7874a,a7875a,a7879a,a7880a,a7883a,a7886a,a7887a,a7888a,a7892a,a7893a,a7896a,a7899a,a7900a,a7901a,a7905a,a7906a,a7909a,a7912a,a7913a,a7914a,a7918a,a7919a,a7922a,a7925a,a7926a,a7927a,a7931a,a7932a,a7935a,a7938a,a7939a,a7940a,a7944a,a7945a,a7948a,a7951a,a7952a,a7953a,a7957a,a7958a,a7961a,a7964a,a7965a,a7966a,a7970a,a7971a,a7974a,a7977a,a7978a,a7979a,a7983a,a7984a,a7987a,a7990a,a7991a,a7992a,a7996a,a7997a,a8000a,a8003a,a8004a,a8005a,a8009a,a8010a,a8013a,a8016a,a8017a,a8018a,a8022a,a8023a,a8026a,a8029a,a8030a,a8031a,a8035a,a8036a,a8039a,a8042a,a8043a,a8044a,a8048a,a8049a,a8052a,a8055a,a8056a,a8057a,a8061a,a8062a,a8065a,a8068a,a8069a,a8070a,a8074a,a8075a,a8078a,a8081a,a8082a,a8083a,a8087a,a8088a,a8091a,a8094a,a8095a,a8096a,a8100a,a8101a,a8104a,a8107a,a8108a,a8109a,a8113a,a8114a,a8117a,a8120a,a8121a,a8122a,a8126a,a8127a,a8130a,a8133a,a8134a,a8135a,a8139a,a8140a,a8143a,a8146a,a8147a,a8148a,a8152a,a8153a,a8156a,a8159a,a8160a,a8161a,a8165a,a8166a,a8169a,a8172a,a8173a,a8174a,a8178a,a8179a,a8182a,a8185a,a8186a,a8187a,a8191a,a8192a,a8195a,a8198a,a8199a,a8200a,a8204a,a8205a,a8208a,a8211a,a8212a,a8213a,a8217a,a8218a,a8221a,a8224a,a8225a,a8226a,a8230a,a8231a,a8234a,a8237a,a8238a,a8239a,a8243a,a8244a,a8247a,a8250a,a8251a,a8252a,a8256a,a8257a,a8260a,a8263a,a8264a,a8265a,a8269a,a8270a,a8273a,a8276a,a8277a,a8278a,a8282a,a8283a,a8286a,a8289a,a8290a,a8291a,a8295a,a8296a,a8299a,a8302a,a8303a,a8304a,a8308a,a8309a,a8312a,a8315a,a8316a,a8317a,a8321a,a8322a,a8325a,a8328a,a8329a,a8330a,a8334a,a8335a,a8338a,a8341a,a8342a,a8343a,a8347a,a8348a,a8351a,a8354a,a8355a,a8356a,a8360a,a8361a,a8364a,a8367a,a8368a,a8369a,a8373a,a8374a,a8377a,a8380a,a8381a,a8382a,a8386a,a8387a,a8390a,a8393a,a8394a,a8395a,a8399a,a8400a,a8403a,a8406a,a8407a,a8408a,a8412a,a8413a,a8416a,a8419a,a8420a,a8421a,a8425a,a8426a,a8429a,a8432a,a8433a,a8434a,a8438a,a8439a,a8442a,a8445a,a8446a,a8447a,a8451a,a8452a,a8455a,a8458a,a8459a,a8460a,a8464a,a8465a,a8468a,a8471a,a8472a,a8473a,a8477a,a8478a,a8481a,a8484a,a8485a,a8486a,a8490a,a8491a,a8494a,a8497a,a8498a,a8499a,a8503a,a8504a,a8507a,a8510a,a8511a,a8512a,a8516a,a8517a,a8520a,a8523a,a8524a,a8525a,a8529a,a8530a,a8533a,a8536a,a8537a,a8538a,a8542a,a8543a,a8546a,a8549a,a8550a,a8551a,a8555a,a8556a,a8559a,a8562a,a8563a,a8564a,a8568a,a8569a,a8572a,a8575a,a8576a,a8577a,a8581a,a8582a,a8585a,a8588a,a8589a,a8590a,a8594a,a8595a,a8598a,a8601a,a8602a,a8603a,a8607a,a8608a,a8611a,a8614a,a8615a,a8616a,a8620a,a8621a,a8624a,a8627a,a8628a,a8629a,a8633a,a8634a,a8637a,a8640a,a8641a,a8642a,a8646a,a8647a,a8650a,a8653a,a8654a,a8655a,a8659a,a8660a,a8663a,a8666a,a8667a,a8668a,a8672a,a8673a,a8676a,a8679a,a8680a,a8681a,a8685a,a8686a,a8689a,a8692a,a8693a,a8694a,a8698a,a8699a,a8702a,a8705a,a8706a,a8707a,a8711a,a8712a,a8715a,a8718a,a8719a,a8720a,a8724a,a8725a,a8728a,a8731a,a8732a,a8733a,a8737a,a8738a,a8741a,a8744a,a8745a,a8746a,a8750a,a8751a,a8754a,a8757a,a8758a,a8759a,a8763a,a8764a,a8767a,a8770a,a8771a,a8772a,a8776a,a8777a,a8780a,a8783a,a8784a,a8785a,a8789a,a8790a,a8793a,a8796a,a8797a,a8798a,a8802a,a8803a,a8806a,a8809a,a8810a,a8811a,a8815a,a8816a,a8819a,a8822a,a8823a,a8824a,a8828a,a8829a,a8832a,a8835a,a8836a,a8837a,a8841a,a8842a,a8845a,a8848a,a8849a,a8850a,a8854a,a8855a,a8858a,a8861a,a8862a,a8863a,a8867a,a8868a,a8871a,a8874a,a8875a,a8876a,a8880a,a8881a,a8884a,a8887a,a8888a,a8889a,a8893a,a8894a,a8897a,a8900a,a8901a,a8902a,a8906a,a8907a,a8910a,a8913a,a8914a,a8915a,a8919a,a8920a,a8923a,a8926a,a8927a,a8928a,a8932a,a8933a,a8936a,a8939a,a8940a,a8941a,a8945a,a8946a,a8949a,a8952a,a8953a,a8954a,a8958a,a8959a,a8962a,a8965a,a8966a,a8967a,a8971a,a8972a,a8975a,a8978a,a8979a,a8980a,a8984a,a8985a,a8988a,a8991a,a8992a,a8993a,a8997a,a8998a,a9001a,a9004a,a9005a,a9006a,a9010a,a9011a,a9014a,a9017a,a9018a,a9019a,a9023a,a9024a,a9027a,a9030a,a9031a,a9032a,a9036a,a9037a,a9040a,a9043a,a9044a,a9045a,a9049a,a9050a,a9053a,a9056a,a9057a,a9058a,a9062a,a9063a,a9066a,a9069a,a9070a,a9071a,a9075a,a9076a,a9079a,a9082a,a9083a,a9084a,a9088a,a9089a,a9092a,a9095a,a9096a,a9097a,a9101a,a9102a,a9105a,a9108a,a9109a,a9110a,a9114a,a9115a,a9118a,a9121a,a9122a,a9123a,a9127a,a9128a,a9131a,a9134a,a9135a,a9136a,a9140a,a9141a,a9144a,a9147a,a9148a,a9149a,a9153a,a9154a,a9157a,a9160a,a9161a,a9162a,a9166a,a9167a,a9170a,a9173a,a9174a,a9175a,a9179a,a9180a,a9183a,a9186a,a9187a,a9188a,a9192a,a9193a,a9196a,a9199a,a9200a,a9201a,a9205a,a9206a,a9209a,a9212a,a9213a,a9214a,a9218a,a9219a,a9222a,a9225a,a9226a,a9227a,a9231a,a9232a,a9235a,a9238a,a9239a,a9240a,a9244a,a9245a,a9248a,a9251a,a9252a,a9253a,a9257a,a9258a,a9261a,a9264a,a9265a,a9266a,a9270a,a9271a,a9274a,a9277a,a9278a,a9279a,a9283a,a9284a,a9287a,a9290a,a9291a,a9292a,a9296a,a9297a,a9300a,a9303a,a9304a,a9305a,a9309a,a9310a,a9313a,a9316a,a9317a,a9318a,a9322a,a9323a,a9326a,a9329a,a9330a,a9331a,a9335a,a9336a,a9339a,a9342a,a9343a,a9344a,a9348a,a9349a,a9352a,a9355a,a9356a,a9357a,a9361a,a9362a,a9365a,a9368a,a9369a,a9370a,a9374a,a9375a,a9378a,a9381a,a9382a,a9383a,a9387a,a9388a,a9391a,a9394a,a9395a,a9396a,a9400a,a9401a,a9404a,a9407a,a9408a,a9409a,a9413a,a9414a,a9417a,a9420a,a9421a,a9422a,a9426a,a9427a,a9430a,a9433a,a9434a,a9435a,a9439a,a9440a,a9443a,a9446a,a9447a,a9448a,a9452a,a9453a,a9456a,a9459a,a9460a,a9461a,a9465a,a9466a,a9469a,a9472a,a9473a,a9474a,a9478a,a9479a,a9482a,a9485a,a9486a,a9487a,a9491a,a9492a,a9495a,a9498a,a9499a,a9500a,a9504a,a9505a,a9508a,a9511a,a9512a,a9513a,a9517a,a9518a,a9521a,a9524a,a9525a,a9526a,a9530a,a9531a,a9534a,a9537a,a9538a,a9539a,a9543a,a9544a,a9547a,a9550a,a9551a,a9552a,a9556a,a9557a,a9560a,a9563a,a9564a,a9565a,a9569a,a9570a,a9573a,a9576a,a9577a,a9578a,a9582a,a9583a,a9586a,a9589a,a9590a,a9591a,a9595a,a9596a,a9599a,a9602a,a9603a,a9604a,a9608a,a9609a,a9612a,a9615a,a9616a,a9617a,a9621a,a9622a,a9625a,a9628a,a9629a,a9630a,a9634a,a9635a,a9638a,a9641a,a9642a,a9643a,a9647a,a9648a,a9651a,a9654a,a9655a,a9656a,a9660a,a9661a,a9664a,a9667a,a9668a,a9669a,a9673a,a9674a,a9677a,a9680a,a9681a,a9682a,a9686a,a9687a,a9690a,a9693a,a9694a,a9695a,a9699a,a9700a,a9703a,a9706a,a9707a,a9708a,a9712a,a9713a,a9716a,a9719a,a9720a,a9721a,a9725a,a9726a,a9729a,a9732a,a9733a,a9734a,a9738a,a9739a,a9742a,a9745a,a9746a,a9747a,a9751a,a9752a,a9755a,a9758a,a9759a,a9760a,a9764a,a9765a,a9768a,a9771a,a9772a,a9773a,a9777a,a9778a,a9781a,a9784a,a9785a,a9786a,a9790a,a9791a,a9794a,a9797a,a9798a,a9799a,a9803a,a9804a,a9807a,a9810a,a9811a,a9812a,a9816a,a9817a,a9820a,a9823a,a9824a,a9825a,a9829a,a9830a,a9833a,a9836a,a9837a,a9838a,a9842a,a9843a,a9846a,a9849a,a9850a,a9851a,a9855a,a9856a,a9859a,a9862a,a9863a,a9864a,a9868a,a9869a,a9872a,a9875a,a9876a,a9877a,a9881a,a9882a,a9885a,a9888a,a9889a,a9890a,a9894a,a9895a,a9898a,a9901a,a9902a,a9903a,a9907a,a9908a,a9911a,a9914a,a9915a,a9916a,a9920a,a9921a,a9924a,a9927a,a9928a,a9929a,a9933a,a9934a,a9937a,a9940a,a9941a,a9942a,a9946a,a9947a,a9950a,a9953a,a9954a,a9955a,a9959a,a9960a,a9963a,a9966a,a9967a,a9968a,a9972a,a9973a,a9976a,a9979a,a9980a,a9981a,a9985a,a9986a,a9989a,a9992a,a9993a,a9994a,a9998a,a9999a,a10002a,a10005a,a10006a,a10007a,a10011a,a10012a,a10015a,a10018a,a10019a,a10020a,a10024a,a10025a,a10028a,a10031a,a10032a,a10033a,a10037a,a10038a,a10041a,a10044a,a10045a,a10046a,a10050a,a10051a,a10054a,a10057a,a10058a,a10059a,a10063a,a10064a,a10067a,a10070a,a10071a,a10072a,a10076a,a10077a,a10080a,a10083a,a10084a,a10085a,a10089a,a10090a,a10093a,a10096a,a10097a,a10098a,a10102a,a10103a,a10106a,a10109a,a10110a,a10111a,a10115a,a10116a,a10119a,a10122a,a10123a,a10124a,a10128a,a10129a,a10132a,a10135a,a10136a,a10137a,a10141a,a10142a,a10145a,a10148a,a10149a,a10150a,a10154a,a10155a,a10158a,a10161a,a10162a,a10163a,a10167a,a10168a,a10171a,a10174a,a10175a,a10176a,a10180a,a10181a,a10184a,a10187a,a10188a,a10189a,a10193a,a10194a,a10197a,a10200a,a10201a,a10202a,a10206a,a10207a,a10210a,a10213a,a10214a,a10215a,a10219a,a10220a,a10223a,a10226a,a10227a,a10228a,a10232a,a10233a,a10236a,a10239a,a10240a,a10241a,a10245a,a10246a,a10249a,a10252a,a10253a,a10254a,a10258a,a10259a,a10262a,a10265a,a10266a,a10267a,a10271a,a10272a,a10275a,a10278a,a10279a,a10280a,a10284a,a10285a,a10288a,a10291a,a10292a,a10293a,a10297a,a10298a,a10301a,a10304a,a10305a,a10306a,a10310a,a10311a,a10314a,a10317a,a10318a,a10319a,a10323a,a10324a,a10327a,a10330a,a10331a,a10332a,a10336a,a10337a,a10340a,a10343a,a10344a,a10345a,a10349a,a10350a,a10353a,a10356a,a10357a,a10358a,a10362a,a10363a,a10366a,a10369a,a10370a,a10371a,a10375a,a10376a,a10379a,a10382a,a10383a,a10384a,a10388a,a10389a,a10392a,a10395a,a10396a,a10397a,a10401a,a10402a,a10405a,a10408a,a10409a,a10410a,a10414a,a10415a,a10418a,a10421a,a10422a,a10423a,a10427a,a10428a,a10431a,a10434a,a10435a,a10436a,a10440a,a10441a,a10444a,a10447a,a10448a,a10449a,a10453a,a10454a,a10457a,a10460a,a10461a,a10462a,a10466a,a10467a,a10470a,a10473a,a10474a,a10475a,a10479a,a10480a,a10483a,a10486a,a10487a,a10488a,a10492a,a10493a,a10496a,a10499a,a10500a,a10501a,a10505a,a10506a,a10509a,a10512a,a10513a,a10514a,a10518a,a10519a,a10522a,a10525a,a10526a,a10527a,a10531a,a10532a,a10535a,a10538a,a10539a,a10540a,a10544a,a10545a,a10548a,a10551a,a10552a,a10553a,a10557a,a10558a,a10561a,a10564a,a10565a,a10566a,a10570a,a10571a,a10574a,a10577a,a10578a,a10579a,a10583a,a10584a,a10587a,a10590a,a10591a,a10592a,a10596a,a10597a,a10600a,a10603a,a10604a,a10605a,a10609a,a10610a,a10613a,a10616a,a10617a,a10618a,a10622a,a10623a,a10626a,a10629a,a10630a,a10631a,a10635a,a10636a,a10639a,a10642a,a10643a,a10644a,a10648a,a10649a,a10652a,a10655a,a10656a,a10657a,a10661a,a10662a,a10665a,a10668a,a10669a,a10670a,a10674a,a10675a,a10678a,a10681a,a10682a,a10683a,a10687a,a10688a,a10691a,a10694a,a10695a,a10696a,a10700a,a10701a,a10704a,a10707a,a10708a,a10709a,a10713a,a10714a,a10717a,a10720a,a10721a,a10722a,a10726a,a10727a,a10730a,a10733a,a10734a,a10735a,a10739a,a10740a,a10743a,a10746a,a10747a,a10748a,a10752a,a10753a,a10756a,a10759a,a10760a,a10761a,a10765a,a10766a,a10769a,a10772a,a10773a,a10774a,a10778a,a10779a,a10782a,a10785a,a10786a,a10787a,a10791a,a10792a,a10795a,a10798a,a10799a,a10800a,a10804a,a10805a,a10808a,a10811a,a10812a,a10813a,a10817a,a10818a,a10821a,a10824a,a10825a,a10826a,a10830a,a10831a,a10834a,a10837a,a10838a,a10839a,a10843a,a10844a,a10847a,a10850a,a10851a,a10852a,a10856a,a10857a,a10860a,a10863a,a10864a,a10865a,a10869a,a10870a,a10873a,a10876a,a10877a,a10878a,a10882a,a10883a,a10886a,a10889a,a10890a,a10891a,a10895a,a10896a,a10899a,a10902a,a10903a,a10904a,a10908a,a10909a,a10912a,a10915a,a10916a,a10917a,a10921a,a10922a,a10925a,a10928a,a10929a,a10930a,a10934a,a10935a,a10938a,a10941a,a10942a,a10943a,a10947a,a10948a,a10951a,a10954a,a10955a,a10956a,a10960a,a10961a,a10964a,a10967a,a10968a,a10969a,a10973a,a10974a,a10977a,a10980a,a10981a,a10982a,a10986a,a10987a,a10990a,a10993a,a10994a,a10995a,a10999a,a11000a,a11003a,a11006a,a11007a,a11008a,a11012a,a11013a,a11016a,a11019a,a11020a,a11021a,a11025a,a11026a,a11029a,a11032a,a11033a,a11034a,a11038a,a11039a,a11042a,a11045a,a11046a,a11047a,a11051a,a11052a,a11055a,a11058a,a11059a,a11060a,a11064a,a11065a,a11068a,a11071a,a11072a,a11073a,a11077a,a11078a,a11081a,a11084a,a11085a,a11086a,a11090a,a11091a,a11094a,a11097a,a11098a,a11099a,a11103a,a11104a,a11107a,a11110a,a11111a,a11112a,a11116a,a11117a,a11120a,a11123a,a11124a,a11125a,a11129a,a11130a,a11133a,a11136a,a11137a,a11138a,a11142a,a11143a,a11146a,a11149a,a11150a,a11151a,a11155a,a11156a,a11159a,a11162a,a11163a,a11164a,a11168a,a11169a,a11172a,a11175a,a11176a,a11177a,a11181a,a11182a,a11185a,a11188a,a11189a,a11190a,a11194a,a11195a,a11198a,a11201a,a11202a,a11203a,a11207a,a11208a,a11211a,a11214a,a11215a,a11216a,a11220a,a11221a,a11224a,a11227a,a11228a,a11229a,a11233a,a11234a,a11237a,a11240a,a11241a,a11242a,a11246a,a11247a,a11250a,a11253a,a11254a,a11255a,a11259a,a11260a,a11263a,a11266a,a11267a,a11268a,a11272a,a11273a,a11276a,a11279a,a11280a,a11281a,a11285a,a11286a,a11289a,a11292a,a11293a,a11294a,a11298a,a11299a,a11302a,a11305a,a11306a,a11307a,a11311a,a11312a,a11315a,a11318a,a11319a,a11320a,a11324a,a11325a,a11328a,a11331a,a11332a,a11333a,a11337a,a11338a,a11341a,a11344a,a11345a,a11346a,a11350a,a11351a,a11354a,a11357a,a11358a,a11359a,a11363a,a11364a,a11367a,a11370a,a11371a,a11372a,a11376a,a11377a,a11380a,a11383a,a11384a,a11385a,a11389a,a11390a,a11393a,a11396a,a11397a,a11398a,a11402a,a11403a,a11406a,a11409a,a11410a,a11411a,a11415a,a11416a,a11419a,a11422a,a11423a,a11424a,a11428a,a11429a,a11432a,a11435a,a11436a,a11437a,a11441a,a11442a,a11445a,a11448a,a11449a,a11450a,a11454a,a11455a,a11458a,a11461a,a11462a,a11463a,a11467a,a11468a,a11471a,a11474a,a11475a,a11476a,a11480a,a11481a,a11484a,a11487a,a11488a,a11489a,a11493a,a11494a,a11497a,a11500a,a11501a,a11502a,a11506a,a11507a,a11510a,a11513a,a11514a,a11515a,a11519a,a11520a,a11523a,a11526a,a11527a,a11528a,a11532a,a11533a,a11536a,a11539a,a11540a,a11541a,a11545a,a11546a,a11549a,a11552a,a11553a,a11554a,a11558a,a11559a,a11562a,a11565a,a11566a,a11567a,a11571a,a11572a,a11575a,a11578a,a11579a,a11580a,a11584a,a11585a,a11588a,a11591a,a11592a,a11593a,a11597a,a11598a,a11601a,a11604a,a11605a,a11606a,a11610a,a11611a,a11614a,a11617a,a11618a,a11619a,a11623a,a11624a,a11627a,a11630a,a11631a,a11632a,a11636a,a11637a,a11640a,a11643a,a11644a,a11645a,a11649a,a11650a,a11653a,a11656a,a11657a,a11658a,a11662a,a11663a,a11666a,a11669a,a11670a,a11671a,a11675a,a11676a,a11679a,a11682a,a11683a,a11684a,a11688a,a11689a,a11692a,a11695a,a11696a,a11697a,a11701a,a11702a,a11705a,a11708a,a11709a,a11710a,a11714a,a11715a,a11718a,a11721a,a11722a,a11723a,a11727a,a11728a,a11731a,a11734a,a11735a,a11736a,a11740a,a11741a,a11744a,a11747a,a11748a,a11749a,a11753a,a11754a,a11757a,a11760a,a11761a,a11762a,a11766a,a11767a,a11770a,a11773a,a11774a,a11775a,a11779a,a11780a,a11783a,a11786a,a11787a,a11788a,a11792a,a11793a,a11796a,a11799a,a11800a,a11801a,a11805a,a11806a,a11809a,a11812a,a11813a,a11814a,a11818a,a11819a,a11822a,a11825a,a11826a,a11827a,a11831a,a11832a,a11835a,a11838a,a11839a,a11840a,a11844a,a11845a,a11848a,a11851a,a11852a,a11853a,a11857a,a11858a,a11861a,a11864a,a11865a,a11866a,a11870a,a11871a,a11874a,a11877a,a11878a,a11879a,a11883a,a11884a,a11887a,a11890a,a11891a,a11892a,a11896a,a11897a,a11900a,a11903a,a11904a,a11905a,a11909a,a11910a,a11913a,a11916a,a11917a,a11918a,a11922a,a11923a,a11926a,a11929a,a11930a,a11931a,a11935a,a11936a,a11939a,a11942a,a11943a,a11944a,a11948a,a11949a,a11952a,a11955a,a11956a,a11957a,a11961a,a11962a,a11965a,a11968a,a11969a,a11970a,a11974a,a11975a,a11978a,a11981a,a11982a,a11983a,a11987a,a11988a,a11991a,a11994a,a11995a,a11996a,a12000a,a12001a,a12004a,a12007a,a12008a,a12009a,a12013a,a12014a,a12017a,a12020a,a12021a,a12022a,a12026a,a12027a,a12030a,a12033a,a12034a,a12035a,a12039a,a12040a,a12043a,a12046a,a12047a,a12048a,a12052a,a12053a,a12056a,a12059a,a12060a,a12061a,a12065a,a12066a,a12069a,a12072a,a12073a,a12074a,a12078a,a12079a,a12082a,a12085a,a12086a,a12087a,a12091a,a12092a,a12095a,a12098a,a12099a,a12100a,a12104a,a12105a,a12108a,a12111a,a12112a,a12113a,a12117a,a12118a,a12121a,a12124a,a12125a,a12126a,a12130a,a12131a,a12134a,a12137a,a12138a,a12139a,a12143a,a12144a,a12147a,a12150a,a12151a,a12152a,a12156a,a12157a,a12160a,a12163a,a12164a,a12165a,a12169a,a12170a,a12173a,a12176a,a12177a,a12178a,a12182a,a12183a,a12186a,a12189a,a12190a,a12191a,a12195a,a12196a,a12199a,a12202a,a12203a,a12204a,a12208a,a12209a,a12212a,a12215a,a12216a,a12217a,a12221a,a12222a,a12225a,a12228a,a12229a,a12230a,a12234a,a12235a,a12238a,a12241a,a12242a,a12243a,a12247a,a12248a,a12251a,a12254a,a12255a,a12256a,a12260a,a12261a,a12264a,a12267a,a12268a,a12269a,a12273a,a12274a,a12277a,a12280a,a12281a,a12282a,a12286a,a12287a,a12290a,a12293a,a12294a,a12295a,a12299a,a12300a,a12303a,a12306a,a12307a,a12308a,a12312a,a12313a,a12316a,a12319a,a12320a,a12321a,a12325a,a12326a,a12329a,a12332a,a12333a,a12334a,a12338a,a12339a,a12342a,a12345a,a12346a,a12347a,a12351a,a12352a,a12355a,a12358a,a12359a,a12360a,a12364a,a12365a,a12368a,a12371a,a12372a,a12373a,a12377a,a12378a,a12381a,a12384a,a12385a,a12386a,a12390a,a12391a,a12394a,a12397a,a12398a,a12399a,a12403a,a12404a,a12407a,a12410a,a12411a,a12412a,a12416a,a12417a,a12420a,a12423a,a12424a,a12425a,a12429a,a12430a,a12433a,a12436a,a12437a,a12438a,a12442a,a12443a,a12446a,a12449a,a12450a,a12451a,a12455a,a12456a,a12459a,a12462a,a12463a,a12464a,a12468a,a12469a,a12472a,a12475a,a12476a,a12477a,a12481a,a12482a,a12485a,a12488a,a12489a,a12490a,a12494a,a12495a,a12498a,a12501a,a12502a,a12503a,a12507a,a12508a,a12511a,a12514a,a12515a,a12516a,a12520a,a12521a,a12524a,a12527a,a12528a,a12529a,a12533a,a12534a,a12537a,a12540a,a12541a,a12542a,a12546a,a12547a,a12550a,a12553a,a12554a,a12555a,a12559a,a12560a,a12563a,a12566a,a12567a,a12568a,a12572a,a12573a,a12576a,a12579a,a12580a,a12581a,a12585a,a12586a,a12589a,a12592a,a12593a,a12594a,a12598a,a12599a,a12602a,a12605a,a12606a,a12607a,a12611a,a12612a,a12615a,a12618a,a12619a,a12620a,a12624a,a12625a,a12628a,a12631a,a12632a,a12633a,a12637a,a12638a,a12641a,a12644a,a12645a,a12646a,a12650a,a12651a,a12654a,a12657a,a12658a,a12659a,a12663a,a12664a,a12667a,a12670a,a12671a,a12672a,a12676a,a12677a,a12680a,a12683a,a12684a,a12685a,a12689a,a12690a,a12693a,a12696a,a12697a,a12698a,a12702a,a12703a,a12706a,a12709a,a12710a,a12711a,a12715a,a12716a,a12719a,a12722a,a12723a,a12724a,a12728a,a12729a,a12732a,a12735a,a12736a,a12737a,a12741a,a12742a,a12745a,a12748a,a12749a,a12750a,a12754a,a12755a,a12758a,a12761a,a12762a,a12763a,a12767a,a12768a,a12771a,a12774a,a12775a,a12776a,a12780a,a12781a,a12784a,a12787a,a12788a,a12789a,a12793a,a12794a,a12797a,a12800a,a12801a,a12802a,a12806a,a12807a,a12810a,a12813a,a12814a,a12815a,a12819a,a12820a,a12823a,a12826a,a12827a,a12828a,a12832a,a12833a,a12836a,a12839a,a12840a,a12841a,a12845a,a12846a,a12849a,a12852a,a12853a,a12854a,a12858a,a12859a,a12862a,a12865a,a12866a,a12867a,a12871a,a12872a,a12875a,a12878a,a12879a,a12880a,a12884a,a12885a,a12888a,a12891a,a12892a,a12893a,a12897a,a12898a,a12901a,a12904a,a12905a,a12906a,a12910a,a12911a,a12914a,a12917a,a12918a,a12919a,a12923a,a12924a,a12927a,a12930a,a12931a,a12932a,a12936a,a12937a,a12940a,a12943a,a12944a,a12945a,a12949a,a12950a,a12953a,a12956a,a12957a,a12958a,a12962a,a12963a,a12966a,a12969a,a12970a,a12971a,a12975a,a12976a,a12979a,a12982a,a12983a,a12984a,a12988a,a12989a,a12992a,a12995a,a12996a,a12997a,a13001a,a13002a,a13005a,a13008a,a13009a,a13010a,a13014a,a13015a,a13018a,a13021a,a13022a,a13023a,a13027a,a13028a,a13031a,a13034a,a13035a,a13036a,a13040a,a13041a,a13044a,a13047a,a13048a,a13049a,a13053a,a13054a,a13057a,a13060a,a13061a,a13062a,a13066a,a13067a,a13070a,a13073a,a13074a,a13075a,a13079a,a13080a,a13083a,a13086a,a13087a,a13088a,a13092a,a13093a,a13096a,a13099a,a13100a,a13101a,a13105a,a13106a,a13109a,a13112a,a13113a,a13114a,a13118a,a13119a,a13122a,a13125a,a13126a,a13127a,a13131a,a13132a,a13135a,a13138a,a13139a,a13140a,a13144a,a13145a,a13148a,a13151a,a13152a,a13153a,a13157a,a13158a,a13161a,a13164a,a13165a,a13166a,a13170a,a13171a,a13174a,a13177a,a13178a,a13179a,a13183a,a13184a,a13187a,a13190a,a13191a,a13192a,a13196a,a13197a,a13200a,a13203a,a13204a,a13205a,a13209a,a13210a,a13213a,a13216a,a13217a,a13218a,a13222a,a13223a,a13226a,a13229a,a13230a,a13231a,a13235a,a13236a,a13239a,a13242a,a13243a,a13244a,a13248a,a13249a,a13252a,a13255a,a13256a,a13257a,a13261a,a13262a,a13265a,a13268a,a13269a,a13270a,a13274a,a13275a,a13278a,a13281a,a13282a,a13283a,a13287a,a13288a,a13291a,a13294a,a13295a,a13296a,a13300a,a13301a,a13304a,a13307a,a13308a,a13309a,a13313a,a13314a,a13317a,a13320a,a13321a,a13322a,a13326a,a13327a,a13330a,a13333a,a13334a,a13335a,a13339a,a13340a,a13343a,a13346a,a13347a,a13348a,a13352a,a13353a,a13356a,a13359a,a13360a,a13361a,a13365a,a13366a,a13369a,a13372a,a13373a,a13374a,a13378a,a13379a,a13382a,a13385a,a13386a,a13387a,a13391a,a13392a,a13395a,a13398a,a13399a,a13400a,a13404a,a13405a,a13408a,a13411a,a13412a,a13413a,a13417a,a13418a,a13421a,a13424a,a13425a,a13426a,a13430a,a13431a,a13434a,a13437a,a13438a,a13439a,a13443a,a13444a,a13447a,a13450a,a13451a,a13452a,a13456a,a13457a,a13460a,a13463a,a13464a,a13465a,a13469a,a13470a,a13473a,a13476a,a13477a,a13478a,a13482a,a13483a,a13486a,a13489a,a13490a,a13491a,a13495a,a13496a,a13499a,a13502a,a13503a,a13504a,a13508a,a13509a,a13512a,a13515a,a13516a,a13517a,a13521a,a13522a,a13525a,a13528a,a13529a,a13530a,a13534a,a13535a,a13538a,a13541a,a13542a,a13543a,a13547a,a13548a,a13551a,a13554a,a13555a,a13556a,a13560a,a13561a,a13564a,a13567a,a13568a,a13569a,a13573a,a13574a,a13577a,a13580a,a13581a,a13582a,a13586a,a13587a,a13590a,a13593a,a13594a,a13595a,a13599a,a13600a,a13603a,a13606a,a13607a,a13608a,a13612a,a13613a,a13616a,a13619a,a13620a,a13621a,a13625a,a13626a,a13629a,a13632a,a13633a,a13634a,a13638a,a13639a,a13642a,a13645a,a13646a,a13647a,a13651a,a13652a,a13655a,a13658a,a13659a,a13660a,a13664a,a13665a,a13668a,a13671a,a13672a,a13673a,a13677a,a13678a,a13681a,a13684a,a13685a,a13686a,a13690a,a13691a,a13694a,a13697a,a13698a,a13699a,a13703a,a13704a,a13707a,a13710a,a13711a,a13712a,a13716a,a13717a,a13720a,a13723a,a13724a,a13725a,a13729a,a13730a,a13733a,a13736a,a13737a,a13738a,a13742a,a13743a,a13746a,a13749a,a13750a,a13751a,a13755a,a13756a,a13759a,a13762a,a13763a,a13764a,a13768a,a13769a,a13772a,a13775a,a13776a,a13777a,a13781a,a13782a,a13785a,a13788a,a13789a,a13790a,a13794a,a13795a,a13798a,a13801a,a13802a,a13803a,a13807a,a13808a,a13811a,a13814a,a13815a,a13816a,a13820a,a13821a,a13824a,a13827a,a13828a,a13829a,a13833a,a13834a,a13837a,a13840a,a13841a,a13842a,a13846a,a13847a,a13850a,a13853a,a13854a,a13855a,a13859a,a13860a,a13863a,a13866a,a13867a,a13868a,a13872a,a13873a,a13876a,a13879a,a13880a,a13881a,a13885a,a13886a,a13889a,a13892a,a13893a,a13894a,a13898a,a13899a,a13902a,a13905a,a13906a,a13907a,a13911a,a13912a,a13915a,a13918a,a13919a,a13920a,a13924a,a13925a,a13928a,a13931a,a13932a,a13933a,a13937a,a13938a,a13941a,a13944a,a13945a,a13946a,a13950a,a13951a,a13954a,a13957a,a13958a,a13959a,a13963a,a13964a,a13967a,a13970a,a13971a,a13972a,a13976a,a13977a,a13980a,a13983a,a13984a,a13985a,a13989a,a13990a,a13993a,a13996a,a13997a,a13998a,a14002a,a14003a,a14006a,a14009a,a14010a,a14011a,a14015a,a14016a,a14019a,a14022a,a14023a,a14024a,a14028a,a14029a,a14032a,a14035a,a14036a,a14037a,a14041a,a14042a,a14045a,a14048a,a14049a,a14050a,a14054a,a14055a,a14058a,a14061a,a14062a,a14063a,a14067a,a14068a,a14071a,a14074a,a14075a,a14076a,a14080a,a14081a,a14084a,a14087a,a14088a,a14089a,a14093a,a14094a,a14097a,a14100a,a14101a,a14102a,a14106a,a14107a,a14110a,a14113a,a14114a,a14115a,a14119a,a14120a,a14123a,a14126a,a14127a,a14128a,a14132a,a14133a,a14136a,a14139a,a14140a,a14141a,a14145a,a14146a,a14149a,a14152a,a14153a,a14154a,a14158a,a14159a,a14162a,a14165a,a14166a,a14167a,a14171a,a14172a,a14175a,a14178a,a14179a,a14180a,a14184a,a14185a,a14188a,a14191a,a14192a,a14193a,a14197a,a14198a,a14201a,a14204a,a14205a,a14206a,a14210a,a14211a,a14214a,a14217a,a14218a,a14219a,a14223a,a14224a,a14227a,a14230a,a14231a,a14232a,a14236a,a14237a,a14240a,a14243a,a14244a,a14245a,a14249a,a14250a,a14253a,a14256a,a14257a,a14258a,a14262a,a14263a,a14266a,a14269a,a14270a,a14271a,a14275a,a14276a,a14279a,a14282a,a14283a,a14284a,a14288a,a14289a,a14292a,a14295a,a14296a,a14297a,a14301a,a14302a,a14305a,a14308a,a14309a,a14310a,a14314a,a14315a,a14318a,a14321a,a14322a,a14323a,a14327a,a14328a,a14331a,a14334a,a14335a,a14336a,a14340a,a14341a,a14344a,a14347a,a14348a,a14349a,a14353a,a14354a,a14357a,a14360a,a14361a,a14362a,a14366a,a14367a,a14370a,a14373a,a14374a,a14375a,a14379a,a14380a,a14383a,a14386a,a14387a,a14388a,a14392a,a14393a,a14396a,a14399a,a14400a,a14401a,a14405a,a14406a,a14409a,a14412a,a14413a,a14414a,a14418a,a14419a,a14422a,a14425a,a14426a,a14427a,a14431a,a14432a,a14435a,a14438a,a14439a,a14440a,a14444a,a14445a,a14448a,a14451a,a14452a,a14453a,a14457a,a14458a,a14461a,a14464a,a14465a,a14466a,a14470a,a14471a,a14474a,a14477a,a14478a,a14479a,a14483a,a14484a,a14487a,a14490a,a14491a,a14492a,a14496a,a14497a,a14500a,a14503a,a14504a,a14505a,a14509a,a14510a,a14513a,a14516a,a14517a,a14518a,a14522a,a14523a,a14526a,a14529a,a14530a,a14531a,a14535a,a14536a,a14539a,a14542a,a14543a,a14544a,a14548a,a14549a,a14552a,a14555a,a14556a,a14557a,a14561a,a14562a,a14565a,a14568a,a14569a,a14570a,a14574a,a14575a,a14578a,a14581a,a14582a,a14583a,a14587a,a14588a,a14591a,a14594a,a14595a,a14596a,a14600a,a14601a,a14604a,a14607a,a14608a,a14609a,a14613a,a14614a,a14617a,a14620a,a14621a,a14622a,a14626a,a14627a,a14630a,a14633a,a14634a,a14635a,a14639a,a14640a,a14643a,a14646a,a14647a,a14648a,a14652a,a14653a,a14656a,a14659a,a14660a,a14661a,a14665a,a14666a,a14669a,a14672a,a14673a,a14674a,a14678a,a14679a,a14682a,a14685a,a14686a,a14687a,a14691a,a14692a,a14695a,a14698a,a14699a,a14700a,a14704a,a14705a,a14708a,a14711a,a14712a,a14713a,a14717a,a14718a,a14721a,a14724a,a14725a,a14726a,a14730a,a14731a,a14734a,a14737a,a14738a,a14739a,a14743a,a14744a,a14747a,a14750a,a14751a,a14752a,a14756a,a14757a,a14760a,a14763a,a14764a,a14765a,a14769a,a14770a,a14773a,a14776a,a14777a,a14778a,a14782a,a14783a,a14786a,a14789a,a14790a,a14791a,a14795a,a14796a,a14799a,a14802a,a14803a,a14804a,a14808a,a14809a,a14812a,a14815a,a14816a,a14817a,a14821a,a14822a,a14825a,a14828a,a14829a,a14830a,a14834a,a14835a,a14838a,a14841a,a14842a,a14843a,a14847a,a14848a,a14851a,a14854a,a14855a,a14856a,a14860a,a14861a,a14864a,a14867a,a14868a,a14869a,a14873a,a14874a,a14877a,a14880a,a14881a,a14882a,a14886a,a14887a,a14890a,a14893a,a14894a,a14895a,a14899a,a14900a,a14903a,a14906a,a14907a,a14908a,a14912a,a14913a,a14916a,a14919a,a14920a,a14921a,a14925a,a14926a,a14929a,a14932a,a14933a,a14934a,a14938a,a14939a,a14942a,a14945a,a14946a,a14947a,a14951a,a14952a,a14955a,a14958a,a14959a,a14960a,a14964a,a14965a,a14968a,a14971a,a14972a,a14973a,a14977a,a14978a,a14981a,a14984a,a14985a,a14986a,a14990a,a14991a,a14994a,a14997a,a14998a,a14999a,a15003a,a15004a,a15007a,a15010a,a15011a,a15012a,a15016a,a15017a,a15020a,a15023a,a15024a,a15025a,a15029a,a15030a,a15033a,a15036a,a15037a,a15038a,a15042a,a15043a,a15046a,a15049a,a15050a,a15051a,a15055a,a15056a,a15059a,a15062a,a15063a,a15064a,a15068a,a15069a,a15072a,a15075a,a15076a,a15077a,a15081a,a15082a,a15085a,a15088a,a15089a,a15090a,a15094a,a15095a,a15098a,a15101a,a15102a,a15103a,a15107a,a15108a,a15111a,a15114a,a15115a,a15116a,a15120a,a15121a,a15124a,a15127a,a15128a,a15129a,a15133a,a15134a,a15137a,a15140a,a15141a,a15142a,a15146a,a15147a,a15150a,a15153a,a15154a,a15155a,a15159a,a15160a,a15163a,a15166a,a15167a,a15168a,a15172a,a15173a,a15176a,a15179a,a15180a,a15181a,a15185a,a15186a,a15189a,a15192a,a15193a,a15194a,a15198a,a15199a,a15202a,a15205a,a15206a,a15207a,a15211a,a15212a,a15215a,a15218a,a15219a,a15220a,a15224a,a15225a,a15228a,a15231a,a15232a,a15233a,a15237a,a15238a,a15241a,a15244a,a15245a,a15246a,a15250a,a15251a,a15254a,a15257a,a15258a,a15259a,a15263a,a15264a,a15267a,a15270a,a15271a,a15272a,a15276a,a15277a,a15280a,a15283a,a15284a,a15285a,a15289a,a15290a,a15293a,a15296a,a15297a,a15298a,a15302a,a15303a,a15306a,a15309a,a15310a,a15311a,a15315a,a15316a,a15319a,a15322a,a15323a,a15324a,a15328a,a15329a,a15332a,a15335a,a15336a,a15337a,a15341a,a15342a,a15345a,a15348a,a15349a,a15350a,a15354a,a15355a,a15358a,a15361a,a15362a,a15363a,a15367a,a15368a,a15371a,a15374a,a15375a,a15376a,a15380a,a15381a,a15384a,a15387a,a15388a,a15389a,a15393a,a15394a,a15397a,a15400a,a15401a,a15402a,a15406a,a15407a,a15410a,a15413a,a15414a,a15415a,a15419a,a15420a,a15423a,a15426a,a15427a,a15428a,a15432a,a15433a,a15436a,a15439a,a15440a,a15441a,a15445a,a15446a,a15449a,a15452a,a15453a,a15454a,a15458a,a15459a,a15462a,a15465a,a15466a,a15467a,a15471a,a15472a,a15475a,a15478a,a15479a,a15480a,a15484a,a15485a,a15488a,a15491a,a15492a,a15493a,a15497a,a15498a,a15501a,a15504a,a15505a,a15506a,a15510a,a15511a,a15514a,a15517a,a15518a,a15519a,a15523a,a15524a,a15527a,a15530a,a15531a,a15532a,a15536a,a15537a,a15540a,a15543a,a15544a,a15545a,a15549a,a15550a,a15553a,a15556a,a15557a,a15558a,a15562a,a15563a,a15566a,a15569a,a15570a,a15571a,a15575a,a15576a,a15579a,a15582a,a15583a,a15584a,a15588a,a15589a,a15592a,a15595a,a15596a,a15597a,a15601a,a15602a,a15605a,a15608a,a15609a,a15610a,a15614a,a15615a,a15618a,a15621a,a15622a,a15623a,a15627a,a15628a,a15631a,a15634a,a15635a,a15636a,a15640a,a15641a,a15644a,a15647a,a15648a,a15649a,a15653a,a15654a,a15657a,a15660a,a15661a,a15662a,a15666a,a15667a,a15670a,a15673a,a15674a,a15675a,a15679a,a15680a,a15683a,a15686a,a15687a,a15688a,a15692a,a15693a,a15696a,a15699a,a15700a,a15701a,a15705a,a15706a,a15709a,a15712a,a15713a,a15714a,a15718a,a15719a,a15722a,a15725a,a15726a,a15727a,a15731a,a15732a,a15735a,a15738a,a15739a,a15740a,a15744a,a15745a,a15748a,a15751a,a15752a,a15753a,a15757a,a15758a,a15761a,a15764a,a15765a,a15766a,a15770a,a15771a,a15774a,a15777a,a15778a,a15779a,a15783a,a15784a,a15787a,a15790a,a15791a,a15792a,a15796a,a15797a,a15800a,a15803a,a15804a,a15805a,a15809a,a15810a,a15813a,a15816a,a15817a,a15818a,a15822a,a15823a,a15826a,a15829a,a15830a,a15831a,a15835a,a15836a,a15839a,a15842a,a15843a,a15844a,a15848a,a15849a,a15852a,a15855a,a15856a,a15857a,a15861a,a15862a,a15865a,a15868a,a15869a,a15870a,a15874a,a15875a,a15878a,a15881a,a15882a,a15883a,a15887a,a15888a,a15891a,a15894a,a15895a,a15896a,a15900a,a15901a,a15904a,a15907a,a15908a,a15909a,a15913a,a15914a,a15917a,a15920a,a15921a,a15922a,a15926a,a15927a,a15930a,a15933a,a15934a,a15935a,a15939a,a15940a,a15943a,a15946a,a15947a,a15948a,a15952a,a15953a,a15956a,a15959a,a15960a,a15961a,a15965a,a15966a,a15969a,a15972a,a15973a,a15974a,a15978a,a15979a,a15982a,a15985a,a15986a,a15987a,a15991a,a15992a,a15995a,a15998a,a15999a,a16000a,a16004a,a16005a,a16008a,a16011a,a16012a,a16013a,a16017a,a16018a,a16021a,a16024a,a16025a,a16026a,a16030a,a16031a,a16034a,a16037a,a16038a,a16039a,a16043a,a16044a,a16047a,a16050a,a16051a,a16052a,a16056a,a16057a,a16060a,a16063a,a16064a,a16065a,a16069a,a16070a,a16073a,a16076a,a16077a,a16078a,a16082a,a16083a,a16086a,a16089a,a16090a,a16091a,a16095a,a16096a,a16099a,a16102a,a16103a,a16104a,a16108a,a16109a,a16112a,a16115a,a16116a,a16117a,a16121a,a16122a,a16125a,a16128a,a16129a,a16130a,a16134a,a16135a,a16138a,a16141a,a16142a,a16143a,a16147a,a16148a,a16151a,a16154a,a16155a,a16156a,a16160a,a16161a,a16164a,a16167a,a16168a,a16169a,a16173a,a16174a,a16177a,a16180a,a16181a,a16182a,a16186a,a16187a,a16190a,a16193a,a16194a,a16195a,a16199a,a16200a,a16203a,a16206a,a16207a,a16208a,a16212a,a16213a,a16216a,a16219a,a16220a,a16221a,a16225a,a16226a,a16229a,a16232a,a16233a,a16234a,a16238a,a16239a,a16242a,a16245a,a16246a,a16247a,a16251a,a16252a,a16255a,a16258a,a16259a,a16260a,a16264a,a16265a,a16268a,a16271a,a16272a,a16273a,a16277a,a16278a,a16281a,a16284a,a16285a,a16286a,a16290a,a16291a,a16294a,a16297a,a16298a,a16299a,a16303a,a16304a,a16307a,a16310a,a16311a,a16312a,a16316a,a16317a,a16320a,a16323a,a16324a,a16325a,a16329a,a16330a,a16333a,a16336a,a16337a,a16338a,a16342a,a16343a,a16346a,a16349a,a16350a,a16351a,a16355a,a16356a,a16359a,a16362a,a16363a,a16364a,a16368a,a16369a,a16372a,a16375a,a16376a,a16377a,a16381a,a16382a,a16385a,a16388a,a16389a,a16390a,a16394a,a16395a,a16398a,a16401a,a16402a,a16403a,a16407a,a16408a,a16411a,a16414a,a16415a,a16416a,a16420a,a16421a,a16424a,a16427a,a16428a,a16429a,a16433a,a16434a,a16437a,a16440a,a16441a,a16442a,a16446a,a16447a,a16450a,a16453a,a16454a,a16455a,a16459a,a16460a,a16463a,a16466a,a16467a,a16468a,a16472a,a16473a,a16476a,a16479a,a16480a,a16481a,a16485a,a16486a,a16489a,a16492a,a16493a,a16494a,a16498a,a16499a,a16502a,a16505a,a16506a,a16507a,a16511a,a16512a,a16515a,a16518a,a16519a,a16520a,a16524a,a16525a,a16528a,a16531a,a16532a,a16533a,a16537a,a16538a,a16541a,a16544a,a16545a,a16546a,a16550a,a16551a,a16554a,a16557a,a16558a,a16559a,a16563a,a16564a,a16567a,a16570a,a16571a,a16572a,a16576a,a16577a,a16580a,a16583a,a16584a,a16585a,a16589a,a16590a,a16593a,a16596a,a16597a,a16598a,a16602a,a16603a,a16606a,a16609a,a16610a,a16611a,a16615a,a16616a,a16619a,a16622a,a16623a,a16624a,a16628a,a16629a,a16632a,a16635a,a16636a,a16637a,a16641a,a16642a,a16645a,a16648a,a16649a,a16650a,a16654a,a16655a,a16658a,a16661a,a16662a,a16663a,a16667a,a16668a,a16671a,a16674a,a16675a,a16676a,a16680a,a16681a,a16684a,a16687a,a16688a,a16689a,a16693a,a16694a,a16697a,a16700a,a16701a,a16702a,a16706a,a16707a,a16710a,a16713a,a16714a,a16715a,a16719a,a16720a,a16723a,a16726a,a16727a,a16728a,a16732a,a16733a,a16736a,a16739a,a16740a,a16741a,a16745a,a16746a,a16749a,a16752a,a16753a,a16754a,a16758a,a16759a,a16762a,a16765a,a16766a,a16767a,a16771a,a16772a,a16775a,a16778a,a16779a,a16780a,a16784a,a16785a,a16788a,a16791a,a16792a,a16793a,a16797a,a16798a,a16801a,a16804a,a16805a,a16806a,a16810a,a16811a,a16814a,a16817a,a16818a,a16819a,a16823a,a16824a,a16827a,a16830a,a16831a,a16832a,a16836a,a16837a,a16840a,a16843a,a16844a,a16845a,a16849a,a16850a,a16853a,a16856a,a16857a,a16858a,a16862a,a16863a,a16866a,a16869a,a16870a,a16871a,a16875a,a16876a,a16879a,a16882a,a16883a,a16884a,a16888a,a16889a,a16892a,a16895a,a16896a,a16897a,a16901a,a16902a,a16905a,a16908a,a16909a,a16910a,a16914a,a16915a,a16918a,a16921a,a16922a,a16923a,a16927a,a16928a,a16931a,a16934a,a16935a,a16936a,a16940a,a16941a,a16944a,a16947a,a16948a,a16949a,a16953a,a16954a,a16957a,a16960a,a16961a,a16962a,a16966a,a16967a,a16970a,a16973a,a16974a,a16975a,a16979a,a16980a,a16983a,a16986a,a16987a,a16988a,a16992a,a16993a,a16996a,a16999a,a17000a,a17001a,a17005a,a17006a,a17009a,a17012a,a17013a,a17014a,a17018a,a17019a,a17022a,a17025a,a17026a,a17027a,a17031a,a17032a,a17035a,a17038a,a17039a,a17040a,a17044a,a17045a,a17048a,a17051a,a17052a,a17053a,a17057a,a17058a,a17061a,a17064a,a17065a,a17066a,a17070a,a17071a,a17074a,a17077a,a17078a,a17079a,a17083a,a17084a,a17087a,a17090a,a17091a,a17092a,a17096a,a17097a,a17100a,a17103a,a17104a,a17105a,a17109a,a17110a,a17113a,a17116a,a17117a,a17118a,a17122a,a17123a,a17126a,a17129a,a17130a,a17131a,a17135a,a17136a,a17139a,a17142a,a17143a,a17144a,a17148a,a17149a,a17152a,a17155a,a17156a,a17157a,a17161a,a17162a,a17165a,a17168a,a17169a,a17170a,a17174a,a17175a,a17178a,a17181a,a17182a,a17183a,a17187a,a17188a,a17191a,a17194a,a17195a,a17196a,a17200a,a17201a,a17204a,a17207a,a17208a,a17209a,a17213a,a17214a,a17217a,a17220a,a17221a,a17222a,a17226a,a17227a,a17230a,a17233a,a17234a,a17235a,a17239a,a17240a,a17243a,a17246a,a17247a,a17248a,a17252a,a17253a,a17256a,a17259a,a17260a,a17261a,a17265a,a17266a,a17269a,a17272a,a17273a,a17274a,a17278a,a17279a,a17282a,a17285a,a17286a,a17287a,a17291a,a17292a,a17295a,a17298a,a17299a,a17300a,a17304a,a17305a,a17308a,a17311a,a17312a,a17313a,a17317a,a17318a,a17321a,a17324a,a17325a,a17326a,a17330a,a17331a,a17334a,a17337a,a17338a,a17339a,a17343a,a17344a,a17347a,a17350a,a17351a,a17352a,a17356a,a17357a,a17360a,a17363a,a17364a,a17365a,a17369a,a17370a,a17373a,a17376a,a17377a,a17378a,a17382a,a17383a,a17386a,a17389a,a17390a,a17391a,a17395a,a17396a,a17399a,a17402a,a17403a,a17404a,a17408a,a17409a,a17412a,a17415a,a17416a,a17417a,a17421a,a17422a,a17425a,a17428a,a17429a,a17430a,a17434a,a17435a,a17438a,a17441a,a17442a,a17443a,a17447a,a17448a,a17451a,a17454a,a17455a,a17456a,a17460a,a17461a,a17464a,a17467a,a17468a,a17469a,a17473a,a17474a,a17477a,a17480a,a17481a,a17482a,a17486a,a17487a,a17490a,a17493a,a17494a,a17495a,a17499a,a17500a,a17503a,a17506a,a17507a,a17508a,a17512a,a17513a,a17516a,a17519a,a17520a,a17521a,a17525a,a17526a,a17529a,a17532a,a17533a,a17534a,a17538a,a17539a,a17542a,a17545a,a17546a,a17547a,a17551a,a17552a,a17555a,a17558a,a17559a,a17560a,a17564a,a17565a,a17568a,a17571a,a17572a,a17573a,a17577a,a17578a,a17581a,a17584a,a17585a,a17586a,a17590a,a17591a,a17594a,a17597a,a17598a,a17599a,a17603a,a17604a,a17607a,a17610a,a17611a,a17612a,a17616a,a17617a,a17620a,a17623a,a17624a,a17625a,a17629a,a17630a,a17633a,a17636a,a17637a,a17638a,a17642a,a17643a,a17646a,a17649a,a17650a,a17651a,a17655a,a17656a,a17659a,a17662a,a17663a,a17664a,a17668a,a17669a,a17672a,a17675a,a17676a,a17677a,a17681a,a17682a,a17685a,a17688a,a17689a,a17690a,a17694a,a17695a,a17698a,a17701a,a17702a,a17703a,a17707a,a17708a,a17711a,a17714a,a17715a,a17716a,a17720a,a17721a,a17724a,a17727a,a17728a,a17729a,a17733a,a17734a,a17737a,a17740a,a17741a,a17742a,a17746a,a17747a,a17750a,a17753a,a17754a,a17755a,a17759a,a17760a,a17763a,a17766a,a17767a,a17768a,a17772a,a17773a,a17776a,a17779a,a17780a,a17781a,a17785a,a17786a,a17789a,a17792a,a17793a,a17794a,a17798a,a17799a,a17802a,a17805a,a17806a,a17807a,a17811a,a17812a,a17815a,a17818a,a17819a,a17820a,a17824a,a17825a,a17828a,a17831a,a17832a,a17833a,a17837a,a17838a,a17841a,a17844a,a17845a,a17846a,a17850a,a17851a,a17854a,a17857a,a17858a,a17859a,a17863a,a17864a,a17867a,a17870a,a17871a,a17872a,a17876a,a17877a,a17880a,a17883a,a17884a,a17885a,a17889a,a17890a,a17893a,a17896a,a17897a,a17898a,a17902a,a17903a,a17906a,a17909a,a17910a,a17911a,a17915a,a17916a,a17919a,a17922a,a17923a,a17924a,a17928a,a17929a,a17932a,a17935a,a17936a,a17937a,a17941a,a17942a,a17945a,a17948a,a17949a,a17950a,a17954a,a17955a,a17958a,a17961a,a17962a,a17963a,a17967a,a17968a,a17971a,a17974a,a17975a,a17976a,a17980a,a17981a,a17984a,a17987a,a17988a,a17989a,a17993a,a17994a,a17997a,a18000a,a18001a,a18002a,a18006a,a18007a,a18010a,a18013a,a18014a,a18015a,a18019a,a18020a,a18023a,a18026a,a18027a,a18028a,a18032a,a18033a,a18036a,a18039a,a18040a,a18041a,a18045a,a18046a,a18049a,a18052a,a18053a,a18054a,a18058a,a18059a,a18062a,a18065a,a18066a,a18067a,a18071a,a18072a,a18075a,a18078a,a18079a,a18080a,a18084a,a18085a,a18088a,a18091a,a18092a,a18093a,a18097a,a18098a,a18101a,a18104a,a18105a,a18106a,a18110a,a18111a,a18114a,a18117a,a18118a,a18119a,a18123a,a18124a,a18127a,a18130a,a18131a,a18132a,a18136a,a18137a,a18140a,a18143a,a18144a,a18145a,a18149a,a18150a,a18153a,a18156a,a18157a,a18158a,a18162a,a18163a,a18166a,a18169a,a18170a,a18171a,a18175a,a18176a,a18179a,a18182a,a18183a,a18184a,a18188a,a18189a,a18192a,a18195a,a18196a,a18197a,a18201a,a18202a,a18205a,a18208a,a18209a,a18210a,a18214a,a18215a,a18218a,a18221a,a18222a,a18223a,a18227a,a18228a,a18231a,a18234a,a18235a,a18236a,a18240a,a18241a,a18244a,a18247a,a18248a,a18249a,a18253a,a18254a,a18257a,a18260a,a18261a,a18262a,a18266a,a18267a,a18270a,a18273a,a18274a,a18275a,a18279a,a18280a,a18283a,a18286a,a18287a,a18288a,a18292a,a18293a,a18296a,a18299a,a18300a,a18301a,a18305a,a18306a,a18309a,a18312a,a18313a,a18314a,a18318a,a18319a,a18322a,a18325a,a18326a,a18327a,a18331a,a18332a,a18335a,a18338a,a18339a,a18340a,a18344a,a18345a,a18348a,a18351a,a18352a,a18353a,a18357a,a18358a,a18361a,a18364a,a18365a,a18366a,a18370a,a18371a,a18374a,a18377a,a18378a,a18379a,a18383a,a18384a,a18387a,a18390a,a18391a,a18392a,a18396a,a18397a,a18400a,a18403a,a18404a,a18405a,a18409a,a18410a,a18413a,a18416a,a18417a,a18418a,a18422a,a18423a,a18426a,a18429a,a18430a,a18431a,a18435a,a18436a,a18439a,a18442a,a18443a,a18444a,a18448a,a18449a,a18452a,a18455a,a18456a,a18457a,a18461a,a18462a,a18465a,a18468a,a18469a,a18470a,a18474a,a18475a,a18478a,a18481a,a18482a,a18483a,a18487a,a18488a,a18491a,a18494a,a18495a,a18496a,a18500a,a18501a,a18504a,a18507a,a18508a,a18509a,a18513a,a18514a,a18517a,a18520a,a18521a,a18522a,a18526a,a18527a,a18530a,a18533a,a18534a,a18535a,a18539a,a18540a,a18543a,a18546a,a18547a,a18548a,a18552a,a18553a,a18556a,a18559a,a18560a,a18561a,a18565a,a18566a,a18569a,a18572a,a18573a,a18574a,a18578a,a18579a,a18582a,a18585a,a18586a,a18587a,a18591a,a18592a,a18595a,a18598a,a18599a,a18600a,a18604a,a18605a,a18608a,a18611a,a18612a,a18613a,a18617a,a18618a,a18621a,a18624a,a18625a,a18626a,a18630a,a18631a,a18634a,a18637a,a18638a,a18639a,a18643a,a18644a,a18647a,a18650a,a18651a,a18652a,a18656a,a18657a,a18660a,a18663a,a18664a,a18665a,a18669a,a18670a,a18673a,a18676a,a18677a,a18678a,a18682a,a18683a,a18686a,a18689a,a18690a,a18691a,a18695a,a18696a,a18699a,a18702a,a18703a,a18704a,a18708a,a18709a,a18712a,a18715a,a18716a,a18717a,a18721a,a18722a,a18725a,a18728a,a18729a,a18730a,a18734a,a18735a,a18738a,a18741a,a18742a,a18743a,a18747a,a18748a,a18751a,a18754a,a18755a,a18756a,a18760a,a18761a,a18764a,a18767a,a18768a,a18769a,a18773a,a18774a,a18777a,a18780a,a18781a,a18782a,a18786a,a18787a,a18790a,a18793a,a18794a,a18795a,a18799a,a18800a,a18803a,a18806a,a18807a,a18808a,a18812a,a18813a,a18816a,a18819a,a18820a,a18821a,a18825a,a18826a,a18829a,a18832a,a18833a,a18834a,a18838a,a18839a,a18842a,a18845a,a18846a,a18847a,a18851a,a18852a,a18855a,a18858a,a18859a,a18860a,a18864a,a18865a,a18868a,a18871a,a18872a,a18873a,a18877a,a18878a,a18881a,a18884a,a18885a,a18886a,a18890a,a18891a,a18894a,a18897a,a18898a,a18899a,a18903a,a18904a,a18907a,a18910a,a18911a,a18912a,a18916a,a18917a,a18920a,a18923a,a18924a,a18925a,a18929a,a18930a,a18933a,a18936a,a18937a,a18938a,a18942a,a18943a,a18946a,a18949a,a18950a,a18951a,a18955a,a18956a,a18959a,a18962a,a18963a,a18964a,a18968a,a18969a,a18972a,a18975a,a18976a,a18977a,a18981a,a18982a,a18985a,a18988a,a18989a,a18990a,a18994a,a18995a,a18998a,a19001a,a19002a,a19003a,a19007a,a19008a,a19011a,a19014a,a19015a,a19016a,a19020a,a19021a,a19024a,a19027a,a19028a,a19029a,a19033a,a19034a,a19037a,a19040a,a19041a,a19042a,a19046a,a19047a,a19050a,a19053a,a19054a,a19055a,a19059a,a19060a,a19063a,a19066a,a19067a,a19068a,a19072a,a19073a,a19076a,a19079a,a19080a,a19081a,a19085a,a19086a,a19089a,a19092a,a19093a,a19094a,a19098a,a19099a,a19102a,a19105a,a19106a,a19107a,a19111a,a19112a,a19115a,a19118a,a19119a,a19120a,a19124a,a19125a,a19128a,a19131a,a19132a,a19133a,a19137a,a19138a,a19141a,a19144a,a19145a,a19146a,a19150a,a19151a,a19154a,a19157a,a19158a,a19159a,a19163a,a19164a,a19167a,a19170a,a19171a,a19172a,a19176a,a19177a,a19180a,a19183a,a19184a,a19185a,a19189a,a19190a,a19193a,a19196a,a19197a,a19198a,a19202a,a19203a,a19206a,a19209a,a19210a,a19211a,a19215a,a19216a,a19219a,a19222a,a19223a,a19224a,a19228a,a19229a,a19232a,a19235a,a19236a,a19237a,a19241a,a19242a,a19245a,a19248a,a19249a,a19250a,a19254a,a19255a,a19258a,a19261a,a19262a,a19263a,a19267a,a19268a,a19271a,a19274a,a19275a,a19276a,a19280a,a19281a,a19284a,a19287a,a19288a,a19289a,a19293a,a19294a,a19297a,a19300a,a19301a,a19302a,a19306a,a19307a,a19310a,a19313a,a19314a,a19315a,a19319a,a19320a,a19323a,a19326a,a19327a,a19328a,a19332a,a19333a,a19336a,a19339a,a19340a,a19341a,a19345a,a19346a,a19349a,a19352a,a19353a,a19354a,a19358a,a19359a,a19362a,a19365a,a19366a,a19367a,a19371a,a19372a,a19375a,a19378a,a19379a,a19380a,a19384a,a19385a,a19388a,a19391a,a19392a,a19393a,a19397a,a19398a,a19401a,a19404a,a19405a,a19406a,a19410a,a19411a,a19414a,a19417a,a19418a,a19419a,a19423a,a19424a,a19427a,a19430a,a19431a,a19432a,a19436a,a19437a,a19440a,a19443a,a19444a,a19445a,a19449a,a19450a,a19453a,a19456a,a19457a,a19458a,a19462a,a19463a,a19466a,a19469a,a19470a,a19471a,a19475a,a19476a,a19479a,a19482a,a19483a,a19484a,a19488a,a19489a,a19492a,a19495a,a19496a,a19497a,a19501a,a19502a,a19505a,a19508a,a19509a,a19510a,a19514a,a19515a,a19518a,a19521a,a19522a,a19523a,a19527a,a19528a,a19531a,a19534a,a19535a,a19536a,a19540a,a19541a,a19544a,a19547a,a19548a,a19549a,a19553a,a19554a,a19557a,a19560a,a19561a,a19562a,a19566a,a19567a,a19570a,a19573a,a19574a,a19575a,a19579a,a19580a,a19583a,a19586a,a19587a,a19588a,a19592a,a19593a,a19596a,a19599a,a19600a,a19601a,a19605a,a19606a,a19609a,a19612a,a19613a,a19614a,a19618a,a19619a,a19622a,a19625a,a19626a,a19627a,a19631a,a19632a,a19635a,a19638a,a19639a,a19640a,a19644a,a19645a,a19648a,a19651a,a19652a,a19653a,a19657a,a19658a,a19661a,a19664a,a19665a,a19666a,a19670a,a19671a,a19674a,a19677a,a19678a,a19679a,a19683a,a19684a,a19687a,a19690a,a19691a,a19692a,a19696a,a19697a,a19700a,a19703a,a19704a,a19705a,a19709a,a19710a,a19713a,a19716a,a19717a,a19718a,a19722a,a19723a,a19726a,a19729a,a19730a,a19731a,a19735a,a19736a,a19739a,a19742a,a19743a,a19744a,a19748a,a19749a,a19752a,a19755a,a19756a,a19757a,a19761a,a19762a,a19765a,a19768a,a19769a,a19770a,a19774a,a19775a,a19778a,a19781a,a19782a,a19783a,a19787a,a19788a,a19791a,a19794a,a19795a,a19796a,a19800a,a19801a,a19804a,a19807a,a19808a,a19809a,a19813a,a19814a,a19817a,a19820a,a19821a,a19822a,a19826a,a19827a,a19830a,a19833a,a19834a,a19835a,a19839a,a19840a,a19843a,a19846a,a19847a,a19848a,a19852a,a19853a,a19856a,a19859a,a19860a,a19861a,a19865a,a19866a,a19869a,a19872a,a19873a,a19874a,a19878a,a19879a,a19882a,a19885a,a19886a,a19887a,a19891a,a19892a,a19895a,a19898a,a19899a,a19900a,a19904a,a19905a,a19908a,a19911a,a19912a,a19913a,a19917a,a19918a,a19921a,a19924a,a19925a,a19926a,a19930a,a19931a,a19934a,a19937a,a19938a,a19939a,a19943a,a19944a,a19947a,a19950a,a19951a,a19952a,a19956a,a19957a,a19960a,a19963a,a19964a,a19965a,a19969a,a19970a,a19973a,a19976a,a19977a,a19978a,a19982a,a19983a,a19986a,a19989a,a19990a,a19991a,a19995a,a19996a,a19999a,a20002a,a20003a,a20004a,a20008a,a20009a,a20012a,a20015a,a20016a,a20017a,a20021a,a20022a,a20025a,a20028a,a20029a,a20030a,a20034a,a20035a,a20038a,a20041a,a20042a,a20043a,a20047a,a20048a,a20051a,a20054a,a20055a,a20056a,a20060a,a20061a,a20064a,a20067a,a20068a,a20069a,a20073a,a20074a,a20077a,a20080a,a20081a,a20082a,a20086a,a20087a,a20090a,a20093a,a20094a,a20095a,a20099a,a20100a,a20103a,a20106a,a20107a,a20108a,a20112a,a20113a,a20116a,a20119a,a20120a,a20121a,a20125a,a20126a,a20129a,a20132a,a20133a,a20134a,a20138a,a20139a,a20142a,a20145a,a20146a,a20147a,a20151a,a20152a,a20155a,a20158a,a20159a,a20160a,a20164a,a20165a,a20168a,a20171a,a20172a,a20173a,a20177a,a20178a,a20181a,a20184a,a20185a,a20186a,a20190a,a20191a,a20194a,a20197a,a20198a,a20199a,a20203a,a20204a,a20207a,a20210a,a20211a,a20212a,a20216a,a20217a,a20220a,a20223a,a20224a,a20225a,a20228a,a20231a,a20232a,a20235a,a20238a,a20239a,a20240a,a20244a,a20245a,a20248a,a20251a,a20252a,a20253a,a20256a,a20259a,a20260a,a20263a,a20266a,a20267a,a20268a,a20272a,a20273a,a20276a,a20279a,a20280a,a20281a,a20284a,a20287a,a20288a,a20291a,a20294a,a20295a,a20296a,a20300a,a20301a,a20304a,a20307a,a20308a,a20309a,a20312a,a20315a,a20316a,a20319a,a20322a,a20323a,a20324a,a20328a,a20329a,a20332a,a20335a,a20336a,a20337a,a20340a,a20343a,a20344a,a20347a,a20350a,a20351a,a20352a,a20356a,a20357a,a20360a,a20363a,a20364a,a20365a,a20368a,a20371a,a20372a,a20375a,a20378a,a20379a,a20380a,a20384a,a20385a,a20388a,a20391a,a20392a,a20393a,a20396a,a20399a,a20400a,a20403a,a20406a,a20407a,a20408a,a20412a,a20413a,a20416a,a20419a,a20420a,a20421a,a20424a,a20427a,a20428a,a20431a,a20434a,a20435a,a20436a,a20440a,a20441a,a20444a,a20447a,a20448a,a20449a,a20452a,a20455a,a20456a,a20459a,a20462a,a20463a,a20464a,a20468a,a20469a,a20472a,a20475a,a20476a,a20477a,a20480a,a20483a,a20484a,a20487a,a20490a,a20491a,a20492a,a20496a,a20497a,a20500a,a20503a,a20504a,a20505a,a20508a,a20511a,a20512a,a20515a,a20518a,a20519a,a20520a,a20524a,a20525a,a20528a,a20531a,a20532a,a20533a,a20536a,a20539a,a20540a,a20543a,a20546a,a20547a,a20548a,a20552a,a20553a,a20556a,a20559a,a20560a,a20561a,a20564a,a20567a,a20568a,a20571a,a20574a,a20575a,a20576a,a20580a,a20581a,a20584a,a20587a,a20588a,a20589a,a20592a,a20595a,a20596a,a20599a,a20602a,a20603a,a20604a,a20608a,a20609a,a20612a,a20615a,a20616a,a20617a,a20620a,a20623a,a20624a,a20627a,a20630a,a20631a,a20632a,a20636a,a20637a,a20640a,a20643a,a20644a,a20645a,a20648a,a20651a,a20652a,a20655a,a20658a,a20659a,a20660a,a20664a,a20665a,a20668a,a20671a,a20672a,a20673a,a20676a,a20679a,a20680a,a20683a,a20686a,a20687a,a20688a,a20692a,a20693a,a20696a,a20699a,a20700a,a20701a,a20704a,a20707a,a20708a,a20711a,a20714a,a20715a,a20716a,a20720a,a20721a,a20724a,a20727a,a20728a,a20729a,a20732a,a20735a,a20736a,a20739a,a20742a,a20743a,a20744a,a20748a,a20749a,a20752a,a20755a,a20756a,a20757a,a20760a,a20763a,a20764a,a20767a,a20770a,a20771a,a20772a,a20776a,a20777a,a20780a,a20783a,a20784a,a20785a,a20788a,a20791a,a20792a,a20795a,a20798a,a20799a,a20800a,a20804a,a20805a,a20808a,a20811a,a20812a,a20813a,a20816a,a20819a,a20820a,a20823a,a20826a,a20827a,a20828a,a20832a,a20833a,a20836a,a20839a,a20840a,a20841a,a20844a,a20847a,a20848a,a20851a,a20854a,a20855a,a20856a,a20860a,a20861a,a20864a,a20867a,a20868a,a20869a,a20872a,a20875a,a20876a,a20879a,a20882a,a20883a,a20884a,a20888a,a20889a,a20892a,a20895a,a20896a,a20897a,a20900a,a20903a,a20904a,a20907a,a20910a,a20911a,a20912a,a20916a,a20917a,a20920a,a20923a,a20924a,a20925a,a20928a,a20931a,a20932a,a20935a,a20938a,a20939a,a20940a,a20944a,a20945a,a20948a,a20951a,a20952a,a20953a,a20956a,a20959a,a20960a,a20963a,a20966a,a20967a,a20968a,a20972a,a20973a,a20976a,a20979a,a20980a,a20981a,a20984a,a20987a,a20988a,a20991a,a20994a,a20995a,a20996a,a21000a,a21001a,a21004a,a21007a,a21008a,a21009a,a21012a,a21015a,a21016a,a21019a,a21022a,a21023a,a21024a,a21028a,a21029a,a21032a,a21035a,a21036a,a21037a,a21040a,a21043a,a21044a,a21047a,a21050a,a21051a,a21052a,a21056a,a21057a,a21060a,a21063a,a21064a,a21065a,a21068a,a21071a,a21072a,a21075a,a21078a,a21079a,a21080a,a21084a,a21085a,a21088a,a21091a,a21092a,a21093a,a21096a,a21099a,a21100a,a21103a,a21106a,a21107a,a21108a,a21112a,a21113a,a21116a,a21119a,a21120a,a21121a,a21124a,a21127a,a21128a,a21131a,a21134a,a21135a,a21136a,a21140a,a21141a,a21144a,a21147a,a21148a,a21149a,a21152a,a21155a,a21156a,a21159a,a21162a,a21163a,a21164a,a21168a,a21169a,a21172a,a21175a,a21176a,a21177a,a21180a,a21183a,a21184a,a21187a,a21190a,a21191a,a21192a,a21196a,a21197a,a21200a,a21203a,a21204a,a21205a,a21208a,a21211a,a21212a,a21215a,a21218a,a21219a,a21220a,a21224a,a21225a,a21228a,a21231a,a21232a,a21233a,a21236a,a21239a,a21240a,a21243a,a21246a,a21247a,a21248a,a21252a,a21253a,a21256a,a21259a,a21260a,a21261a,a21264a,a21267a,a21268a,a21271a,a21274a,a21275a,a21276a,a21280a,a21281a,a21284a,a21287a,a21288a,a21289a,a21292a,a21295a,a21296a,a21299a,a21302a,a21303a,a21304a,a21308a,a21309a,a21312a,a21315a,a21316a,a21317a,a21320a,a21323a,a21324a,a21327a,a21330a,a21331a,a21332a,a21336a,a21337a,a21340a,a21343a,a21344a,a21345a,a21348a,a21351a,a21352a,a21355a,a21358a,a21359a,a21360a,a21364a,a21365a,a21368a,a21371a,a21372a,a21373a,a21376a,a21379a,a21380a,a21383a,a21386a,a21387a,a21388a,a21392a,a21393a,a21396a,a21399a,a21400a,a21401a,a21404a,a21407a,a21408a,a21411a,a21414a,a21415a,a21416a,a21420a,a21421a,a21424a,a21427a,a21428a,a21429a,a21432a,a21435a,a21436a,a21439a,a21442a,a21443a,a21444a,a21448a,a21449a,a21452a,a21455a,a21456a,a21457a,a21460a,a21463a,a21464a,a21467a,a21470a,a21471a,a21472a,a21476a,a21477a,a21480a,a21483a,a21484a,a21485a,a21488a,a21491a,a21492a,a21495a,a21498a,a21499a,a21500a,a21504a,a21505a,a21508a,a21511a,a21512a,a21513a,a21516a,a21519a,a21520a,a21523a,a21526a,a21527a,a21528a,a21532a,a21533a,a21536a,a21539a,a21540a,a21541a,a21544a,a21547a,a21548a,a21551a,a21554a,a21555a,a21556a,a21560a,a21561a,a21564a,a21567a,a21568a,a21569a,a21572a,a21575a,a21576a,a21579a,a21582a,a21583a,a21584a,a21588a,a21589a,a21592a,a21595a,a21596a,a21597a,a21600a,a21603a,a21604a,a21607a,a21610a,a21611a,a21612a,a21616a,a21617a,a21620a,a21623a,a21624a,a21625a,a21628a,a21631a,a21632a,a21635a,a21638a,a21639a,a21640a,a21644a,a21645a,a21648a,a21651a,a21652a,a21653a,a21656a,a21659a,a21660a,a21663a,a21666a,a21667a,a21668a,a21672a,a21673a,a21676a,a21679a,a21680a,a21681a,a21684a,a21687a,a21688a,a21691a,a21694a,a21695a,a21696a,a21700a,a21701a,a21704a,a21707a,a21708a,a21709a,a21712a,a21715a,a21716a,a21719a,a21722a,a21723a,a21724a,a21728a,a21729a,a21732a,a21735a,a21736a,a21737a,a21740a,a21743a,a21744a,a21747a,a21750a,a21751a,a21752a,a21756a,a21757a,a21760a,a21763a,a21764a,a21765a,a21768a,a21771a,a21772a,a21775a,a21778a,a21779a,a21780a,a21784a,a21785a,a21788a,a21791a,a21792a,a21793a,a21796a,a21799a,a21800a,a21803a,a21806a,a21807a,a21808a,a21812a,a21813a,a21816a,a21819a,a21820a,a21821a,a21824a,a21827a,a21828a,a21831a,a21834a,a21835a,a21836a,a21840a,a21841a,a21844a,a21847a,a21848a,a21849a,a21852a,a21855a,a21856a,a21859a,a21862a,a21863a,a21864a,a21868a,a21869a,a21872a,a21875a,a21876a,a21877a,a21880a,a21883a,a21884a,a21887a,a21890a,a21891a,a21892a,a21896a,a21897a,a21900a,a21903a,a21904a,a21905a,a21908a,a21911a,a21912a,a21915a,a21918a,a21919a,a21920a,a21924a,a21925a,a21928a,a21931a,a21932a,a21933a,a21936a,a21939a,a21940a,a21943a,a21946a,a21947a,a21948a,a21952a,a21953a,a21956a,a21959a,a21960a,a21961a,a21964a,a21967a,a21968a,a21971a,a21974a,a21975a,a21976a,a21980a,a21981a,a21984a,a21987a,a21988a,a21989a,a21992a,a21995a,a21996a,a21999a,a22002a,a22003a,a22004a,a22008a,a22009a,a22012a,a22015a,a22016a,a22017a,a22020a,a22023a,a22024a,a22027a,a22030a,a22031a,a22032a,a22036a,a22037a,a22040a,a22043a,a22044a,a22045a,a22048a,a22051a,a22052a,a22055a,a22058a,a22059a,a22060a,a22064a,a22065a,a22068a,a22071a,a22072a,a22073a,a22076a,a22079a,a22080a,a22083a,a22086a,a22087a,a22088a,a22092a,a22093a,a22096a,a22099a,a22100a,a22101a,a22104a,a22107a,a22108a,a22111a,a22114a,a22115a,a22116a,a22120a,a22121a,a22124a,a22127a,a22128a,a22129a,a22132a,a22135a,a22136a,a22139a,a22142a,a22143a,a22144a,a22148a,a22149a,a22152a,a22155a,a22156a,a22157a,a22160a,a22163a,a22164a,a22167a,a22170a,a22171a,a22172a,a22176a,a22177a,a22180a,a22183a,a22184a,a22185a,a22188a,a22191a,a22192a,a22195a,a22198a,a22199a,a22200a,a22204a,a22205a,a22208a,a22211a,a22212a,a22213a,a22216a,a22219a,a22220a,a22223a,a22226a,a22227a,a22228a,a22232a,a22233a,a22236a,a22239a,a22240a,a22241a,a22244a,a22247a,a22248a,a22251a,a22254a,a22255a,a22256a,a22260a,a22261a,a22264a,a22267a,a22268a,a22269a,a22272a,a22275a,a22276a,a22279a,a22282a,a22283a,a22284a,a22288a,a22289a,a22292a,a22295a,a22296a,a22297a,a22300a,a22303a,a22304a,a22307a,a22310a,a22311a,a22312a,a22316a,a22317a,a22320a,a22323a,a22324a,a22325a,a22328a,a22331a,a22332a,a22335a,a22338a,a22339a,a22340a,a22344a,a22345a,a22348a,a22351a,a22352a,a22353a,a22356a,a22359a,a22360a,a22363a,a22366a,a22367a,a22368a,a22372a,a22373a,a22376a,a22379a,a22380a,a22381a,a22384a,a22387a,a22388a,a22391a,a22394a,a22395a,a22396a,a22400a,a22401a,a22404a,a22407a,a22408a,a22409a,a22412a,a22415a,a22416a,a22419a,a22422a,a22423a,a22424a,a22428a,a22429a,a22432a,a22435a,a22436a,a22437a,a22440a,a22443a,a22444a,a22447a,a22450a,a22451a,a22452a,a22456a,a22457a,a22460a,a22463a,a22464a,a22465a,a22468a,a22471a,a22472a,a22475a,a22478a,a22479a,a22480a,a22484a,a22485a,a22488a,a22491a,a22492a,a22493a,a22496a,a22499a,a22500a,a22503a,a22506a,a22507a,a22508a,a22512a,a22513a,a22516a,a22519a,a22520a,a22521a,a22524a,a22527a,a22528a,a22531a,a22534a,a22535a,a22536a,a22540a,a22541a,a22544a,a22547a,a22548a,a22549a,a22552a,a22555a,a22556a,a22559a,a22562a,a22563a,a22564a,a22568a,a22569a,a22572a,a22575a,a22576a,a22577a,a22580a,a22583a,a22584a,a22587a,a22590a,a22591a,a22592a,a22596a,a22597a,a22600a,a22603a,a22604a,a22605a,a22608a,a22611a,a22612a,a22615a,a22618a,a22619a,a22620a,a22624a,a22625a,a22628a,a22631a,a22632a,a22633a,a22636a,a22639a,a22640a,a22643a,a22646a,a22647a,a22648a,a22652a,a22653a,a22656a,a22659a,a22660a,a22661a,a22664a,a22667a,a22668a,a22671a,a22674a,a22675a,a22676a,a22680a,a22681a,a22684a,a22687a,a22688a,a22689a,a22692a,a22695a,a22696a,a22699a,a22702a,a22703a,a22704a,a22708a,a22709a,a22712a,a22715a,a22716a,a22717a,a22720a,a22723a,a22724a,a22727a,a22730a,a22731a,a22732a,a22736a,a22737a,a22740a,a22743a,a22744a,a22745a,a22748a,a22751a,a22752a,a22755a,a22758a,a22759a,a22760a,a22764a,a22765a,a22768a,a22771a,a22772a,a22773a,a22776a,a22779a,a22780a,a22783a,a22786a,a22787a,a22788a,a22792a,a22793a,a22796a,a22799a,a22800a,a22801a,a22804a,a22807a,a22808a,a22811a,a22814a,a22815a,a22816a,a22820a,a22821a,a22824a,a22827a,a22828a,a22829a,a22832a,a22835a,a22836a,a22839a,a22842a,a22843a,a22844a,a22848a,a22849a,a22852a,a22855a,a22856a,a22857a,a22860a,a22863a,a22864a,a22867a,a22870a,a22871a,a22872a,a22876a,a22877a,a22880a,a22883a,a22884a,a22885a,a22888a,a22891a,a22892a,a22895a,a22898a,a22899a,a22900a,a22904a,a22905a,a22908a,a22911a,a22912a,a22913a,a22916a,a22919a,a22920a,a22923a,a22926a,a22927a,a22928a,a22932a,a22933a,a22936a,a22939a,a22940a,a22941a,a22944a,a22947a,a22948a,a22951a,a22954a,a22955a,a22956a,a22960a,a22961a,a22964a,a22967a,a22968a,a22969a,a22972a,a22975a,a22976a,a22979a,a22982a,a22983a,a22984a,a22988a,a22989a,a22992a,a22995a,a22996a,a22997a,a23000a,a23003a,a23004a,a23007a,a23010a,a23011a,a23012a,a23016a,a23017a,a23020a,a23023a,a23024a,a23025a,a23028a,a23031a,a23032a,a23035a,a23038a,a23039a,a23040a,a23044a,a23045a,a23048a,a23051a,a23052a,a23053a,a23056a,a23059a,a23060a,a23063a,a23066a,a23067a,a23068a,a23072a,a23073a,a23076a,a23079a,a23080a,a23081a,a23084a,a23087a,a23088a,a23091a,a23094a,a23095a,a23096a,a23100a,a23101a,a23104a,a23107a,a23108a,a23109a,a23112a,a23115a,a23116a,a23119a,a23122a,a23123a,a23124a,a23128a,a23129a,a23132a,a23135a,a23136a,a23137a,a23140a,a23143a,a23144a,a23147a,a23150a,a23151a,a23152a,a23156a,a23157a,a23160a,a23163a,a23164a,a23165a,a23168a,a23171a,a23172a,a23175a,a23178a,a23179a,a23180a,a23184a,a23185a,a23188a,a23191a,a23192a,a23193a,a23196a,a23199a,a23200a,a23203a,a23206a,a23207a,a23208a,a23212a,a23213a,a23216a,a23219a,a23220a,a23221a,a23224a,a23227a,a23228a,a23231a,a23234a,a23235a,a23236a,a23240a,a23241a,a23244a,a23247a,a23248a,a23249a,a23252a,a23255a,a23256a,a23259a,a23262a,a23263a,a23264a,a23268a,a23269a,a23272a,a23275a,a23276a,a23277a,a23280a,a23283a,a23284a,a23287a,a23290a,a23291a,a23292a,a23296a,a23297a,a23300a,a23303a,a23304a,a23305a,a23308a,a23311a,a23312a,a23315a,a23318a,a23319a,a23320a,a23324a,a23325a,a23328a,a23331a,a23332a,a23333a,a23336a,a23339a,a23340a,a23343a,a23346a,a23347a,a23348a,a23352a,a23353a,a23356a,a23359a,a23360a,a23361a,a23364a,a23367a,a23368a,a23371a,a23374a,a23375a,a23376a,a23380a,a23381a,a23384a,a23387a,a23388a,a23389a,a23392a,a23395a,a23396a,a23399a,a23402a,a23403a,a23404a,a23408a,a23409a,a23412a,a23415a,a23416a,a23417a,a23420a,a23423a,a23424a,a23427a,a23430a,a23431a,a23432a,a23436a,a23437a,a23440a,a23443a,a23444a,a23445a,a23448a,a23451a,a23452a,a23455a,a23458a,a23459a,a23460a,a23464a,a23465a,a23468a,a23471a,a23472a,a23473a,a23476a,a23479a,a23480a,a23483a,a23486a,a23487a,a23488a,a23492a,a23493a,a23496a,a23499a,a23500a,a23501a,a23504a,a23507a,a23508a,a23511a,a23514a,a23515a,a23516a,a23520a,a23521a,a23524a,a23527a,a23528a,a23529a,a23532a,a23535a,a23536a,a23539a,a23542a,a23543a,a23544a,a23548a,a23549a,a23552a,a23555a,a23556a,a23557a,a23560a,a23563a,a23564a,a23567a,a23570a,a23571a,a23572a,a23576a,a23577a,a23580a,a23583a,a23584a,a23585a,a23588a,a23591a,a23592a,a23595a,a23598a,a23599a,a23600a,a23604a,a23605a,a23608a,a23611a,a23612a,a23613a,a23616a,a23619a,a23620a,a23623a,a23626a,a23627a,a23628a,a23632a,a23633a,a23636a,a23639a,a23640a,a23641a,a23644a,a23647a,a23648a,a23651a,a23654a,a23655a,a23656a,a23660a,a23661a,a23664a,a23667a,a23668a,a23669a,a23672a,a23675a,a23676a,a23679a,a23682a,a23683a,a23684a,a23688a,a23689a,a23692a,a23695a,a23696a,a23697a,a23700a,a23703a,a23704a,a23707a,a23710a,a23711a,a23712a,a23716a,a23717a,a23720a,a23723a,a23724a,a23725a,a23728a,a23731a,a23732a,a23735a,a23738a,a23739a,a23740a,a23744a,a23745a,a23748a,a23751a,a23752a,a23753a,a23756a,a23759a,a23760a,a23763a,a23766a,a23767a,a23768a,a23772a,a23773a,a23776a,a23779a,a23780a,a23781a,a23784a,a23787a,a23788a,a23791a,a23794a,a23795a,a23796a,a23800a,a23801a,a23804a,a23807a,a23808a,a23809a,a23812a,a23815a,a23816a,a23819a,a23822a,a23823a,a23824a,a23828a,a23829a,a23832a,a23835a,a23836a,a23837a,a23840a,a23843a,a23844a,a23847a,a23850a,a23851a,a23852a,a23856a,a23857a,a23860a,a23863a,a23864a,a23865a,a23868a,a23871a,a23872a,a23875a,a23878a,a23879a,a23880a,a23884a,a23885a,a23888a,a23891a,a23892a,a23893a,a23896a,a23899a,a23900a,a23903a,a23906a,a23907a,a23908a,a23912a,a23913a,a23916a,a23919a,a23920a,a23921a,a23924a,a23927a,a23928a,a23931a,a23934a,a23935a,a23936a,a23940a,a23941a,a23944a,a23947a,a23948a,a23949a,a23952a,a23955a,a23956a,a23959a,a23962a,a23963a,a23964a,a23968a,a23969a,a23972a,a23975a,a23976a,a23977a,a23980a,a23983a,a23984a,a23987a,a23990a,a23991a,a23992a,a23996a,a23997a,a24000a,a24003a,a24004a,a24005a,a24008a,a24011a,a24012a,a24015a,a24018a,a24019a,a24020a,a24024a,a24025a,a24028a,a24031a,a24032a,a24033a,a24036a,a24039a,a24040a,a24043a,a24046a,a24047a,a24048a,a24052a,a24053a,a24056a,a24059a,a24060a,a24061a,a24064a,a24067a,a24068a,a24071a,a24074a,a24075a,a24076a,a24080a,a24081a,a24084a,a24087a,a24088a,a24089a,a24092a,a24095a,a24096a,a24099a,a24102a,a24103a,a24104a,a24108a,a24109a,a24112a,a24115a,a24116a,a24117a,a24120a,a24123a,a24124a,a24127a,a24130a,a24131a,a24132a,a24136a,a24137a,a24140a,a24143a,a24144a,a24145a,a24148a,a24151a,a24152a,a24155a,a24158a,a24159a,a24160a,a24164a,a24165a,a24168a,a24171a,a24172a,a24173a,a24176a,a24179a,a24180a,a24183a,a24186a,a24187a,a24188a,a24192a,a24193a,a24196a,a24199a,a24200a,a24201a,a24204a,a24207a,a24208a,a24211a,a24214a,a24215a,a24216a,a24220a,a24221a,a24224a,a24227a,a24228a,a24229a,a24232a,a24235a,a24236a,a24239a,a24242a,a24243a,a24244a,a24248a,a24249a,a24252a,a24255a,a24256a,a24257a,a24260a,a24263a,a24264a,a24267a,a24270a,a24271a,a24272a,a24276a,a24277a,a24280a,a24283a,a24284a,a24285a,a24288a,a24291a,a24292a,a24295a,a24298a,a24299a,a24300a,a24304a,a24305a,a24308a,a24311a,a24312a,a24313a,a24316a,a24319a,a24320a,a24323a,a24326a,a24327a,a24328a,a24332a,a24333a,a24336a,a24339a,a24340a,a24341a,a24344a,a24347a,a24348a,a24351a,a24354a,a24355a,a24356a,a24360a,a24361a,a24364a,a24367a,a24368a,a24369a,a24372a,a24375a,a24376a,a24379a,a24382a,a24383a,a24384a,a24388a,a24389a,a24392a,a24395a,a24396a,a24397a,a24400a,a24403a,a24404a,a24407a,a24410a,a24411a,a24412a,a24416a,a24417a,a24420a,a24423a,a24424a,a24425a,a24428a,a24431a,a24432a,a24435a,a24438a,a24439a,a24440a,a24444a,a24445a,a24448a,a24451a,a24452a,a24453a,a24456a,a24459a,a24460a,a24463a,a24466a,a24467a,a24468a,a24472a,a24473a,a24476a,a24479a,a24480a,a24481a,a24484a,a24487a,a24488a,a24491a,a24494a,a24495a,a24496a,a24500a,a24501a,a24504a,a24507a,a24508a,a24509a,a24512a,a24515a,a24516a,a24519a,a24522a,a24523a,a24524a,a24528a,a24529a,a24532a,a24535a,a24536a,a24537a,a24540a,a24543a,a24544a,a24547a,a24550a,a24551a,a24552a,a24556a,a24557a,a24560a,a24563a,a24564a,a24565a,a24568a,a24571a,a24572a,a24575a,a24578a,a24579a,a24580a,a24584a,a24585a,a24588a,a24591a,a24592a,a24593a,a24596a,a24599a,a24600a,a24603a,a24606a,a24607a,a24608a,a24612a,a24613a,a24616a,a24619a,a24620a,a24621a,a24624a,a24627a,a24628a,a24631a,a24634a,a24635a,a24636a,a24640a,a24641a,a24644a,a24647a,a24648a,a24649a,a24652a,a24655a,a24656a,a24659a,a24662a,a24663a,a24664a,a24668a,a24669a,a24672a,a24675a,a24676a,a24677a,a24680a,a24683a,a24684a,a24687a,a24690a,a24691a,a24692a,a24696a,a24697a,a24700a,a24703a,a24704a,a24705a,a24708a,a24711a,a24712a,a24715a,a24718a,a24719a,a24720a,a24724a,a24725a,a24728a,a24731a,a24732a,a24733a,a24736a,a24739a,a24740a,a24743a,a24746a,a24747a,a24748a,a24752a,a24753a,a24756a,a24759a,a24760a,a24761a,a24764a,a24767a,a24768a,a24771a,a24774a,a24775a,a24776a,a24780a,a24781a,a24784a,a24787a,a24788a,a24789a,a24792a,a24795a,a24796a,a24799a,a24802a,a24803a,a24804a,a24808a,a24809a,a24812a,a24815a,a24816a,a24817a,a24820a,a24823a,a24824a,a24827a,a24830a,a24831a,a24832a,a24836a,a24837a,a24840a,a24843a,a24844a,a24845a,a24848a,a24851a,a24852a,a24855a,a24858a,a24859a,a24860a,a24864a,a24865a,a24868a,a24871a,a24872a,a24873a,a24876a,a24879a,a24880a,a24883a,a24886a,a24887a,a24888a,a24892a,a24893a,a24896a,a24899a,a24900a,a24901a,a24904a,a24907a,a24908a,a24911a,a24914a,a24915a,a24916a,a24920a,a24921a,a24924a,a24927a,a24928a,a24929a,a24932a,a24935a,a24936a,a24939a,a24942a,a24943a,a24944a,a24948a,a24949a,a24952a,a24955a,a24956a,a24957a,a24960a,a24963a,a24964a,a24967a,a24970a,a24971a,a24972a,a24976a,a24977a,a24980a,a24983a,a24984a,a24985a,a24988a,a24991a,a24992a,a24995a,a24998a,a24999a,a25000a,a25004a,a25005a,a25008a,a25011a,a25012a,a25013a,a25016a,a25019a,a25020a,a25023a,a25026a,a25027a,a25028a,a25032a,a25033a,a25036a,a25039a,a25040a,a25041a,a25044a,a25047a,a25048a,a25051a,a25054a,a25055a,a25056a,a25060a,a25061a,a25064a,a25067a,a25068a,a25069a,a25072a,a25075a,a25076a,a25079a,a25082a,a25083a,a25084a,a25088a,a25089a,a25092a,a25095a,a25096a,a25097a,a25100a,a25103a,a25104a,a25107a,a25110a,a25111a,a25112a,a25116a,a25117a,a25120a,a25123a,a25124a,a25125a,a25128a,a25131a,a25132a,a25135a,a25138a,a25139a,a25140a,a25144a,a25145a,a25148a,a25151a,a25152a,a25153a,a25156a,a25159a,a25160a,a25163a,a25166a,a25167a,a25168a,a25172a,a25173a,a25176a,a25179a,a25180a,a25181a,a25184a,a25187a,a25188a,a25191a,a25194a,a25195a,a25196a,a25200a,a25201a,a25204a,a25207a,a25208a,a25209a,a25212a,a25215a,a25216a,a25219a,a25222a,a25223a,a25224a,a25228a,a25229a,a25232a,a25235a,a25236a,a25237a,a25240a,a25243a,a25244a,a25247a,a25250a,a25251a,a25252a,a25256a,a25257a,a25260a,a25263a,a25264a,a25265a,a25268a,a25271a,a25272a,a25275a,a25278a,a25279a,a25280a,a25284a,a25285a,a25288a,a25291a,a25292a,a25293a,a25296a,a25299a,a25300a,a25303a,a25306a,a25307a,a25308a,a25312a,a25313a,a25316a,a25319a,a25320a,a25321a,a25324a,a25327a,a25328a,a25331a,a25334a,a25335a,a25336a,a25340a,a25341a,a25344a,a25347a,a25348a,a25349a,a25352a,a25355a,a25356a,a25359a,a25362a,a25363a,a25364a,a25368a,a25369a,a25372a,a25375a,a25376a,a25377a,a25380a,a25383a,a25384a,a25387a,a25390a,a25391a,a25392a,a25396a,a25397a,a25400a,a25403a,a25404a,a25405a,a25408a,a25411a,a25412a,a25415a,a25418a,a25419a,a25420a,a25424a,a25425a,a25428a,a25431a,a25432a,a25433a,a25436a,a25439a,a25440a,a25443a,a25446a,a25447a,a25448a,a25452a,a25453a,a25456a,a25459a,a25460a,a25461a,a25464a,a25467a,a25468a,a25471a,a25474a,a25475a,a25476a,a25480a,a25481a,a25484a,a25487a,a25488a,a25489a,a25492a,a25495a,a25496a,a25499a,a25502a,a25503a,a25504a,a25508a,a25509a,a25512a,a25515a,a25516a,a25517a,a25520a,a25523a,a25524a,a25527a,a25530a,a25531a,a25532a,a25536a,a25537a,a25540a,a25543a,a25544a,a25545a,a25548a,a25551a,a25552a,a25555a,a25558a,a25559a,a25560a,a25564a,a25565a,a25568a,a25571a,a25572a,a25573a,a25576a,a25579a,a25580a,a25583a,a25586a,a25587a,a25588a,a25592a,a25593a,a25596a,a25599a,a25600a,a25601a,a25604a,a25607a,a25608a,a25611a,a25614a,a25615a,a25616a,a25620a,a25621a,a25624a,a25627a,a25628a,a25629a,a25632a,a25635a,a25636a,a25639a,a25642a,a25643a,a25644a,a25648a,a25649a,a25652a,a25655a,a25656a,a25657a,a25660a,a25663a,a25664a,a25667a,a25670a,a25671a,a25672a,a25676a,a25677a,a25680a,a25683a,a25684a,a25685a,a25688a,a25691a,a25692a,a25695a,a25698a,a25699a,a25700a,a25704a,a25705a,a25708a,a25711a,a25712a,a25713a,a25716a,a25719a,a25720a,a25723a,a25726a,a25727a,a25728a,a25732a,a25733a,a25736a,a25739a,a25740a,a25741a,a25744a,a25747a,a25748a,a25751a,a25754a,a25755a,a25756a,a25760a,a25761a,a25764a,a25767a,a25768a,a25769a,a25772a,a25775a,a25776a,a25779a,a25782a,a25783a,a25784a,a25788a,a25789a,a25792a,a25795a,a25796a,a25797a,a25800a,a25803a,a25804a,a25807a,a25810a,a25811a,a25812a,a25816a,a25817a,a25820a,a25823a,a25824a,a25825a,a25828a,a25831a,a25832a,a25835a,a25838a,a25839a,a25840a,a25844a,a25845a,a25848a,a25851a,a25852a,a25853a,a25856a,a25859a,a25860a,a25863a,a25866a,a25867a,a25868a,a25872a,a25873a,a25876a,a25879a,a25880a,a25881a,a25884a,a25887a,a25888a,a25891a,a25894a,a25895a,a25896a,a25900a,a25901a,a25904a,a25907a,a25908a,a25909a,a25912a,a25915a,a25916a,a25919a,a25922a,a25923a,a25924a,a25928a,a25929a,a25932a,a25935a,a25936a,a25937a,a25940a,a25943a,a25944a,a25947a,a25950a,a25951a,a25952a,a25956a,a25957a,a25960a,a25963a,a25964a,a25965a,a25968a,a25971a,a25972a,a25975a,a25978a,a25979a,a25980a,a25984a,a25985a,a25988a,a25991a,a25992a,a25993a,a25996a,a25999a,a26000a,a26003a,a26006a,a26007a,a26008a,a26012a,a26013a,a26016a,a26019a,a26020a,a26021a,a26024a,a26027a,a26028a,a26031a,a26034a,a26035a,a26036a,a26040a,a26041a,a26044a,a26047a,a26048a,a26049a,a26052a,a26055a,a26056a,a26059a,a26062a,a26063a,a26064a,a26068a,a26069a,a26072a,a26075a,a26076a,a26077a,a26080a,a26083a,a26084a,a26087a,a26090a,a26091a,a26092a,a26096a,a26097a,a26100a,a26103a,a26104a,a26105a,a26108a,a26111a,a26112a,a26115a,a26118a,a26119a,a26120a,a26124a,a26125a,a26128a,a26131a,a26132a,a26133a,a26136a,a26139a,a26140a,a26143a,a26146a,a26147a,a26148a,a26152a,a26153a,a26156a,a26159a,a26160a,a26161a,a26164a,a26167a,a26168a,a26171a,a26174a,a26175a,a26176a,a26180a,a26181a,a26184a,a26187a,a26188a,a26189a,a26192a,a26195a,a26196a,a26199a,a26202a,a26203a,a26204a,a26208a,a26209a,a26212a,a26215a,a26216a,a26217a,a26220a,a26223a,a26224a,a26227a,a26230a,a26231a,a26232a,a26236a,a26237a,a26240a,a26243a,a26244a,a26245a,a26248a,a26251a,a26252a,a26255a,a26258a,a26259a,a26260a,a26264a,a26265a,a26268a,a26271a,a26272a,a26273a,a26276a,a26279a,a26280a,a26283a,a26286a,a26287a,a26288a,a26292a,a26293a,a26296a,a26299a,a26300a,a26301a,a26304a,a26307a,a26308a,a26311a,a26314a,a26315a,a26316a,a26320a,a26321a,a26324a,a26327a,a26328a,a26329a,a26332a,a26335a,a26336a,a26339a,a26342a,a26343a,a26344a,a26348a,a26349a,a26352a,a26355a,a26356a,a26357a,a26360a,a26363a,a26364a,a26367a,a26370a,a26371a,a26372a,a26376a,a26377a,a26380a,a26383a,a26384a,a26385a,a26388a,a26391a,a26392a,a26395a,a26398a,a26399a,a26400a,a26404a,a26405a,a26408a,a26411a,a26412a,a26413a,a26416a,a26419a,a26420a,a26423a,a26426a,a26427a,a26428a,a26432a,a26433a,a26436a,a26439a,a26440a,a26441a,a26444a,a26447a,a26448a,a26451a,a26454a,a26455a,a26456a,a26460a,a26461a,a26464a,a26467a,a26468a,a26469a,a26472a,a26475a,a26476a,a26479a,a26482a,a26483a,a26484a,a26488a,a26489a,a26492a,a26495a,a26496a,a26497a,a26500a,a26503a,a26504a,a26507a,a26510a,a26511a,a26512a,a26516a,a26517a,a26520a,a26523a,a26524a,a26525a,a26528a,a26531a,a26532a,a26535a,a26538a,a26539a,a26540a,a26544a,a26545a,a26548a,a26551a,a26552a,a26553a,a26556a,a26559a,a26560a,a26563a,a26566a,a26567a,a26568a,a26572a,a26573a,a26576a,a26579a,a26580a,a26581a,a26584a,a26587a,a26588a,a26591a,a26594a,a26595a,a26596a,a26600a,a26601a,a26604a,a26607a,a26608a,a26609a,a26612a,a26615a,a26616a,a26619a,a26622a,a26623a,a26624a,a26628a,a26629a,a26632a,a26635a,a26636a,a26637a,a26640a,a26643a,a26644a,a26647a,a26650a,a26651a,a26652a,a26656a,a26657a,a26660a,a26663a,a26664a,a26665a,a26668a,a26671a,a26672a,a26675a,a26678a,a26679a,a26680a,a26684a,a26685a,a26688a,a26691a,a26692a,a26693a,a26696a,a26699a,a26700a,a26703a,a26706a,a26707a,a26708a,a26712a,a26713a,a26716a,a26719a,a26720a,a26721a,a26724a,a26727a,a26728a,a26731a,a26734a,a26735a,a26736a,a26740a,a26741a,a26744a,a26747a,a26748a,a26749a,a26752a,a26755a,a26756a,a26759a,a26762a,a26763a,a26764a,a26768a,a26769a,a26772a,a26775a,a26776a,a26777a,a26780a,a26783a,a26784a,a26787a,a26790a,a26791a,a26792a,a26796a,a26797a,a26800a,a26803a,a26804a,a26805a,a26808a,a26811a,a26812a,a26815a,a26818a,a26819a,a26820a,a26824a,a26825a,a26828a,a26831a,a26832a,a26833a,a26836a,a26839a,a26840a,a26843a,a26846a,a26847a,a26848a,a26852a,a26853a,a26856a,a26859a,a26860a,a26861a,a26864a,a26867a,a26868a,a26871a,a26874a,a26875a,a26876a,a26880a,a26881a,a26884a,a26887a,a26888a,a26889a,a26892a,a26895a,a26896a,a26899a,a26902a,a26903a,a26904a,a26908a,a26909a,a26912a,a26915a,a26916a,a26917a,a26920a,a26923a,a26924a,a26927a,a26930a,a26931a,a26932a,a26936a,a26937a,a26940a,a26943a,a26944a,a26945a,a26948a,a26951a,a26952a,a26955a,a26958a,a26959a,a26960a,a26964a,a26965a,a26968a,a26971a,a26972a,a26973a,a26976a,a26979a,a26980a,a26983a,a26986a,a26987a,a26988a,a26992a,a26993a,a26996a,a26999a,a27000a,a27001a,a27004a,a27007a,a27008a,a27011a,a27014a,a27015a,a27016a,a27020a,a27021a,a27024a,a27027a,a27028a,a27029a,a27032a,a27035a,a27036a,a27039a,a27042a,a27043a,a27044a,a27048a,a27049a,a27052a,a27055a,a27056a,a27057a,a27060a,a27063a,a27064a,a27067a,a27070a,a27071a,a27072a,a27076a,a27077a,a27080a,a27083a,a27084a,a27085a,a27088a,a27091a,a27092a,a27095a,a27098a,a27099a,a27100a,a27104a,a27105a,a27108a,a27111a,a27112a,a27113a,a27116a,a27119a,a27120a,a27123a,a27126a,a27127a,a27128a,a27132a,a27133a,a27136a,a27139a,a27140a,a27141a,a27144a,a27147a,a27148a,a27151a,a27154a,a27155a,a27156a,a27160a,a27161a,a27164a,a27167a,a27168a,a27169a,a27172a,a27175a,a27176a,a27179a,a27182a,a27183a,a27184a,a27188a,a27189a,a27192a,a27195a,a27196a,a27197a,a27200a,a27203a,a27204a,a27207a,a27210a,a27211a,a27212a,a27216a,a27217a,a27220a,a27223a,a27224a,a27225a,a27228a,a27231a,a27232a,a27235a,a27238a,a27239a,a27240a,a27244a,a27245a,a27248a,a27251a,a27252a,a27253a,a27256a,a27259a,a27260a,a27263a,a27266a,a27267a,a27268a,a27272a,a27273a,a27276a,a27279a,a27280a,a27281a,a27284a,a27287a,a27288a,a27291a,a27294a,a27295a,a27296a,a27300a,a27301a,a27304a,a27307a,a27308a,a27309a,a27312a,a27315a,a27316a,a27319a,a27322a,a27323a,a27324a,a27328a,a27329a,a27332a,a27335a,a27336a,a27337a,a27340a,a27343a,a27344a,a27347a,a27350a,a27351a,a27352a,a27356a,a27357a,a27360a,a27363a,a27364a,a27365a,a27368a,a27371a,a27372a,a27375a,a27378a,a27379a,a27380a,a27384a,a27385a,a27388a,a27391a,a27392a,a27393a,a27396a,a27399a,a27400a,a27403a,a27406a,a27407a,a27408a,a27412a,a27413a,a27416a,a27419a,a27420a,a27421a,a27424a,a27427a,a27428a,a27431a,a27434a,a27435a,a27436a,a27440a,a27441a,a27444a,a27447a,a27448a,a27449a,a27452a,a27455a,a27456a,a27459a,a27462a,a27463a,a27464a,a27468a,a27469a,a27472a,a27475a,a27476a,a27477a,a27480a,a27483a,a27484a,a27487a,a27490a,a27491a,a27492a,a27496a,a27497a,a27500a,a27503a,a27504a,a27505a,a27508a,a27511a,a27512a,a27515a,a27518a,a27519a,a27520a,a27524a,a27525a,a27528a,a27531a,a27532a,a27533a,a27536a,a27539a,a27540a,a27543a,a27546a,a27547a,a27548a,a27552a,a27553a,a27556a,a27559a,a27560a,a27561a,a27564a,a27567a,a27568a,a27571a,a27574a,a27575a,a27576a,a27580a,a27581a,a27584a,a27587a,a27588a,a27589a,a27592a,a27595a,a27596a,a27599a,a27602a,a27603a,a27604a,a27608a,a27609a,a27612a,a27615a,a27616a,a27617a,a27620a,a27623a,a27624a,a27627a,a27630a,a27631a,a27632a,a27636a,a27637a,a27640a,a27643a,a27644a,a27645a,a27648a,a27651a,a27652a,a27655a,a27658a,a27659a,a27660a,a27664a,a27665a,a27668a,a27671a,a27672a,a27673a,a27676a,a27679a,a27680a,a27683a,a27686a,a27687a,a27688a,a27692a,a27693a,a27696a,a27699a,a27700a,a27701a,a27704a,a27707a,a27708a,a27711a,a27714a,a27715a,a27716a,a27720a,a27721a,a27724a,a27727a,a27728a,a27729a,a27732a,a27735a,a27736a,a27739a,a27742a,a27743a,a27744a,a27748a,a27749a,a27752a,a27755a,a27756a,a27757a,a27760a,a27763a,a27764a,a27767a,a27770a,a27771a,a27772a,a27776a,a27777a,a27780a,a27783a,a27784a,a27785a,a27788a,a27791a,a27792a,a27795a,a27798a,a27799a,a27800a,a27804a,a27805a,a27808a,a27811a,a27812a,a27813a,a27816a,a27819a,a27820a,a27823a,a27826a,a27827a,a27828a,a27832a,a27833a,a27836a,a27839a,a27840a,a27841a,a27844a,a27847a,a27848a,a27851a,a27854a,a27855a,a27856a,a27860a,a27861a,a27864a,a27867a,a27868a,a27869a,a27872a,a27875a,a27876a,a27879a,a27882a,a27883a,a27884a,a27888a,a27889a,a27892a,a27895a,a27896a,a27897a,a27900a,a27903a,a27904a,a27907a,a27910a,a27911a,a27912a,a27916a,a27917a,a27920a,a27923a,a27924a,a27925a,a27928a,a27931a,a27932a,a27935a,a27938a,a27939a,a27940a,a27944a,a27945a,a27948a,a27951a,a27952a,a27953a,a27956a,a27959a,a27960a,a27963a,a27966a,a27967a,a27968a,a27972a,a27973a,a27976a,a27979a,a27980a,a27981a,a27984a,a27987a,a27988a,a27991a,a27994a,a27995a,a27996a,a28000a,a28001a,a28004a,a28007a,a28008a,a28009a,a28012a,a28015a,a28016a,a28019a,a28022a,a28023a,a28024a,a28028a,a28029a,a28032a,a28035a,a28036a,a28037a,a28040a,a28043a,a28044a,a28047a,a28050a,a28051a,a28052a,a28056a,a28057a,a28060a,a28063a,a28064a,a28065a,a28068a,a28071a,a28072a,a28075a,a28078a,a28079a,a28080a,a28084a,a28085a,a28088a,a28091a,a28092a,a28093a,a28096a,a28099a,a28100a,a28103a,a28106a,a28107a,a28108a,a28112a,a28113a,a28116a,a28119a,a28120a,a28121a,a28124a,a28127a,a28128a,a28131a,a28134a,a28135a,a28136a,a28140a,a28141a,a28144a,a28147a,a28148a,a28149a,a28152a,a28155a,a28156a,a28159a,a28162a,a28163a,a28164a,a28168a,a28169a,a28172a,a28175a,a28176a,a28177a,a28180a,a28183a,a28184a,a28187a,a28190a,a28191a,a28192a,a28196a,a28197a,a28200a,a28203a,a28204a,a28205a,a28208a,a28211a,a28212a,a28215a,a28218a,a28219a,a28220a,a28224a,a28225a,a28228a,a28231a,a28232a,a28233a,a28236a,a28239a,a28240a,a28243a,a28246a,a28247a,a28248a,a28252a,a28253a,a28256a,a28259a,a28260a,a28261a,a28264a,a28267a,a28268a,a28271a,a28274a,a28275a,a28276a,a28280a,a28281a,a28284a,a28287a,a28288a,a28289a,a28292a,a28295a,a28296a,a28299a,a28302a,a28303a,a28304a,a28308a,a28309a,a28312a,a28315a,a28316a,a28317a,a28320a,a28323a,a28324a,a28327a,a28330a,a28331a,a28332a,a28336a,a28337a,a28340a,a28343a,a28344a,a28345a,a28348a,a28351a,a28352a,a28355a,a28358a,a28359a,a28360a,a28364a,a28365a,a28368a,a28371a,a28372a,a28373a,a28376a,a28379a,a28380a,a28383a,a28386a,a28387a,a28388a,a28392a,a28393a,a28396a,a28399a,a28400a,a28401a,a28404a,a28407a,a28408a,a28411a,a28414a,a28415a,a28416a,a28420a,a28421a,a28424a,a28427a,a28428a,a28429a,a28432a,a28435a,a28436a,a28439a,a28442a,a28443a,a28444a,a28448a,a28449a,a28452a,a28455a,a28456a,a28457a,a28460a,a28463a,a28464a,a28467a,a28470a,a28471a,a28472a,a28476a,a28477a,a28480a,a28483a,a28484a,a28485a,a28488a,a28491a,a28492a,a28495a,a28498a,a28499a,a28500a,a28504a,a28505a,a28508a,a28511a,a28512a,a28513a,a28516a,a28519a,a28520a,a28523a,a28526a,a28527a,a28528a,a28532a,a28533a,a28536a,a28539a,a28540a,a28541a,a28544a,a28547a,a28548a,a28551a,a28554a,a28555a,a28556a,a28560a,a28561a,a28564a,a28567a,a28568a,a28569a,a28572a,a28575a,a28576a,a28579a,a28582a,a28583a,a28584a,a28588a,a28589a,a28592a,a28595a,a28596a,a28597a,a28600a,a28603a,a28604a,a28607a,a28610a,a28611a,a28612a,a28616a,a28617a,a28620a,a28623a,a28624a,a28625a,a28628a,a28631a,a28632a,a28635a,a28638a,a28639a,a28640a,a28644a,a28645a,a28648a,a28651a,a28652a,a28653a,a28656a,a28659a,a28660a,a28663a,a28666a,a28667a,a28668a,a28672a,a28673a,a28676a,a28679a,a28680a,a28681a,a28684a,a28687a,a28688a,a28691a,a28694a,a28695a,a28696a,a28700a,a28701a,a28704a,a28707a,a28708a,a28709a,a28712a,a28715a,a28716a,a28719a,a28722a,a28723a,a28724a,a28728a,a28729a,a28732a,a28735a,a28736a,a28737a,a28740a,a28743a,a28744a,a28747a,a28750a,a28751a,a28752a,a28756a,a28757a,a28760a,a28763a,a28764a,a28765a,a28768a,a28771a,a28772a,a28775a,a28778a,a28779a,a28780a,a28784a,a28785a,a28788a,a28791a,a28792a,a28793a,a28796a,a28799a,a28800a,a28803a,a28806a,a28807a,a28808a,a28812a,a28813a,a28816a,a28819a,a28820a,a28821a,a28824a,a28827a,a28828a,a28831a,a28834a,a28835a,a28836a,a28840a,a28841a,a28844a,a28847a,a28848a,a28849a,a28852a,a28855a,a28856a,a28859a,a28862a,a28863a,a28864a,a28868a,a28869a,a28872a,a28875a,a28876a,a28877a,a28880a,a28883a,a28884a,a28887a,a28890a,a28891a,a28892a,a28896a,a28897a,a28900a,a28903a,a28904a,a28905a,a28908a,a28911a,a28912a,a28915a,a28918a,a28919a,a28920a,a28924a,a28925a,a28928a,a28931a,a28932a,a28933a,a28936a,a28939a,a28940a,a28943a,a28946a,a28947a,a28948a,a28952a,a28953a,a28956a,a28959a,a28960a,a28961a,a28964a,a28967a,a28968a,a28971a,a28974a,a28975a,a28976a,a28980a,a28981a,a28984a,a28987a,a28988a,a28989a,a28992a,a28995a,a28996a,a28999a,a29002a,a29003a,a29004a,a29008a,a29009a,a29012a,a29015a,a29016a,a29017a,a29020a,a29023a,a29024a,a29027a,a29030a,a29031a,a29032a,a29036a,a29037a,a29040a,a29043a,a29044a,a29045a,a29048a,a29051a,a29052a,a29055a,a29058a,a29059a,a29060a,a29064a,a29065a,a29068a,a29071a,a29072a,a29073a,a29076a,a29079a,a29080a,a29083a,a29086a,a29087a,a29088a,a29092a,a29093a,a29096a,a29099a,a29100a,a29101a,a29104a,a29107a,a29108a,a29111a,a29114a,a29115a,a29116a,a29120a,a29121a,a29124a,a29127a,a29128a,a29129a,a29132a,a29135a,a29136a,a29139a,a29142a,a29143a,a29144a,a29148a,a29149a,a29152a,a29155a,a29156a,a29157a,a29160a,a29163a,a29164a,a29167a,a29170a,a29171a,a29172a,a29176a,a29177a,a29180a,a29183a,a29184a,a29185a,a29188a,a29191a,a29192a,a29195a,a29198a,a29199a,a29200a,a29204a,a29205a,a29208a,a29211a,a29212a,a29213a,a29216a,a29219a,a29220a,a29223a,a29226a,a29227a,a29228a,a29232a,a29233a,a29236a,a29239a,a29240a,a29241a,a29244a,a29247a,a29248a,a29251a,a29254a,a29255a,a29256a,a29260a,a29261a,a29264a,a29267a,a29268a,a29269a,a29272a,a29275a,a29276a,a29279a,a29282a,a29283a,a29284a,a29288a,a29289a,a29292a,a29295a,a29296a,a29297a,a29300a,a29303a,a29304a,a29307a,a29310a,a29311a,a29312a,a29316a,a29317a,a29320a,a29323a,a29324a,a29325a,a29328a,a29331a,a29332a,a29335a,a29338a,a29339a,a29340a,a29344a,a29345a,a29348a,a29351a,a29352a,a29353a,a29356a,a29359a,a29360a,a29363a,a29366a,a29367a,a29368a,a29372a,a29373a,a29376a,a29379a,a29380a,a29381a,a29384a,a29387a,a29388a,a29391a,a29394a,a29395a,a29396a,a29400a,a29401a,a29404a,a29407a,a29408a,a29409a,a29412a,a29415a,a29416a,a29419a,a29422a,a29423a,a29424a,a29428a,a29429a,a29432a,a29435a,a29436a,a29437a,a29440a,a29443a,a29444a,a29447a,a29450a,a29451a,a29452a,a29456a,a29457a,a29460a,a29463a,a29464a,a29465a,a29468a,a29471a,a29472a,a29475a,a29478a,a29479a,a29480a,a29484a,a29485a,a29488a,a29491a,a29492a,a29493a,a29496a,a29499a,a29500a,a29503a,a29506a,a29507a,a29508a,a29512a,a29513a,a29516a,a29519a,a29520a,a29521a,a29524a,a29527a,a29528a,a29531a,a29534a,a29535a,a29536a,a29540a,a29541a,a29544a,a29547a,a29548a,a29549a,a29552a,a29555a,a29556a,a29559a,a29562a,a29563a,a29564a,a29568a,a29569a,a29572a,a29575a,a29576a,a29577a,a29580a,a29583a,a29584a,a29587a,a29590a,a29591a,a29592a,a29596a,a29597a,a29600a,a29603a,a29604a,a29605a,a29608a,a29611a,a29612a,a29615a,a29618a,a29619a,a29620a,a29624a,a29625a,a29628a,a29631a,a29632a,a29633a,a29636a,a29639a,a29640a,a29643a,a29646a,a29647a,a29648a,a29652a,a29653a,a29656a,a29659a,a29660a,a29661a,a29664a,a29667a,a29668a,a29671a,a29674a,a29675a,a29676a,a29680a,a29681a,a29684a,a29687a,a29688a,a29689a,a29692a,a29695a,a29696a,a29699a,a29702a,a29703a,a29704a,a29708a,a29709a,a29712a,a29715a,a29716a,a29717a,a29720a,a29723a,a29724a,a29727a,a29730a,a29731a,a29732a,a29736a,a29737a,a29740a,a29743a,a29744a,a29745a,a29748a,a29751a,a29752a,a29755a,a29758a,a29759a,a29760a,a29764a,a29765a,a29768a,a29771a,a29772a,a29773a,a29776a,a29779a,a29780a,a29783a,a29786a,a29787a,a29788a,a29792a,a29793a,a29796a,a29799a,a29800a,a29801a,a29804a,a29807a,a29808a,a29811a,a29814a,a29815a,a29816a,a29820a,a29821a,a29824a,a29827a,a29828a,a29829a,a29832a,a29835a,a29836a,a29839a,a29842a,a29843a,a29844a,a29848a,a29849a,a29852a,a29855a,a29856a,a29857a,a29860a,a29863a,a29864a,a29867a,a29870a,a29871a,a29872a,a29876a,a29877a,a29880a,a29883a,a29884a,a29885a,a29888a,a29891a,a29892a,a29895a,a29898a,a29899a,a29900a,a29904a,a29905a,a29908a,a29911a,a29912a,a29913a,a29916a,a29919a,a29920a,a29923a,a29926a,a29927a,a29928a,a29932a,a29933a,a29936a,a29939a,a29940a,a29941a,a29944a,a29947a,a29948a,a29951a,a29954a,a29955a,a29956a,a29960a,a29961a,a29964a,a29967a,a29968a,a29969a,a29972a,a29975a,a29976a,a29979a,a29982a,a29983a,a29984a,a29988a,a29989a,a29992a,a29995a,a29996a,a29997a,a30000a,a30003a,a30004a,a30007a,a30010a,a30011a,a30012a,a30016a,a30017a,a30020a,a30023a,a30024a,a30025a,a30028a,a30031a,a30032a,a30035a,a30038a,a30039a,a30040a,a30044a,a30045a,a30048a,a30051a,a30052a,a30053a,a30056a,a30059a,a30060a,a30063a,a30066a,a30067a,a30068a,a30072a,a30073a,a30076a,a30079a,a30080a,a30081a,a30084a,a30087a,a30088a,a30091a,a30094a,a30095a,a30096a,a30100a,a30101a,a30104a,a30107a,a30108a,a30109a,a30112a,a30115a,a30116a,a30119a,a30122a,a30123a,a30124a,a30128a,a30129a,a30132a,a30135a,a30136a,a30137a,a30140a,a30143a,a30144a,a30147a,a30150a,a30151a,a30152a,a30156a,a30157a,a30160a,a30163a,a30164a,a30165a,a30168a,a30171a,a30172a,a30175a,a30178a,a30179a,a30180a,a30184a,a30185a,a30188a,a30191a,a30192a,a30193a,a30196a,a30199a,a30200a,a30203a,a30206a,a30207a,a30208a,a30212a,a30213a,a30216a,a30219a,a30220a,a30221a,a30224a,a30227a,a30228a,a30231a,a30234a,a30235a,a30236a,a30240a,a30241a,a30244a,a30247a,a30248a,a30249a,a30252a,a30255a,a30256a,a30259a,a30262a,a30263a,a30264a,a30268a,a30269a,a30272a,a30275a,a30276a,a30277a,a30280a,a30283a,a30284a,a30287a,a30290a,a30291a,a30292a,a30296a,a30297a,a30300a,a30303a,a30304a,a30305a,a30308a,a30311a,a30312a,a30315a,a30318a,a30319a,a30320a,a30324a,a30325a,a30328a,a30331a,a30332a,a30333a,a30336a,a30339a,a30340a,a30343a,a30346a,a30347a,a30348a,a30352a,a30353a,a30356a,a30359a,a30360a,a30361a,a30364a,a30367a,a30368a,a30371a,a30374a,a30375a,a30376a,a30380a,a30381a,a30384a,a30387a,a30388a,a30389a,a30392a,a30395a,a30396a,a30399a,a30402a,a30403a,a30404a,a30408a,a30409a,a30412a,a30415a,a30416a,a30417a,a30420a,a30423a,a30424a,a30427a,a30430a,a30431a,a30432a,a30436a,a30437a,a30440a,a30443a,a30444a,a30445a,a30448a,a30451a,a30452a,a30455a,a30458a,a30459a,a30460a,a30464a,a30465a,a30468a,a30471a,a30472a,a30473a,a30476a,a30479a,a30480a,a30483a,a30486a,a30487a,a30488a,a30492a,a30493a,a30496a,a30499a,a30500a,a30501a,a30504a,a30507a,a30508a,a30511a,a30514a,a30515a,a30516a,a30520a,a30521a,a30524a,a30527a,a30528a,a30529a,a30532a,a30535a,a30536a,a30539a,a30542a,a30543a,a30544a,a30548a,a30549a,a30552a,a30555a,a30556a,a30557a,a30560a,a30563a,a30564a,a30567a,a30570a,a30571a,a30572a,a30576a,a30577a,a30580a,a30583a,a30584a,a30585a,a30588a,a30591a,a30592a,a30595a,a30598a,a30599a,a30600a,a30604a,a30605a,a30608a,a30611a,a30612a,a30613a,a30616a,a30619a,a30620a,a30623a,a30626a,a30627a,a30628a,a30632a,a30633a,a30636a,a30639a,a30640a,a30641a,a30644a,a30647a,a30648a,a30651a,a30654a,a30655a,a30656a,a30660a,a30661a,a30664a,a30667a,a30668a,a30669a,a30672a,a30675a,a30676a,a30679a,a30682a,a30683a,a30684a,a30688a,a30689a,a30692a,a30695a,a30696a,a30697a,a30700a,a30703a,a30704a,a30707a,a30710a,a30711a,a30712a,a30716a,a30717a,a30720a,a30723a,a30724a,a30725a,a30728a,a30731a,a30732a,a30735a,a30738a,a30739a,a30740a,a30744a,a30745a,a30748a,a30751a,a30752a,a30753a,a30756a,a30759a,a30760a,a30763a,a30766a,a30767a,a30768a,a30772a,a30773a,a30776a,a30779a,a30780a,a30781a,a30784a,a30787a,a30788a,a30791a,a30794a,a30795a,a30796a,a30800a,a30801a,a30804a,a30807a,a30808a,a30809a,a30812a,a30815a,a30816a,a30819a,a30822a,a30823a,a30824a,a30828a,a30829a,a30832a,a30835a,a30836a,a30837a,a30840a,a30843a,a30844a,a30847a,a30850a,a30851a,a30852a,a30856a,a30857a,a30860a,a30863a,a30864a,a30865a,a30868a,a30871a,a30872a,a30875a,a30878a,a30879a,a30880a,a30884a,a30885a,a30888a,a30891a,a30892a,a30893a,a30896a,a30899a,a30900a,a30903a,a30906a,a30907a,a30908a,a30912a,a30913a,a30916a,a30919a,a30920a,a30921a,a30924a,a30927a,a30928a,a30931a,a30934a,a30935a,a30936a,a30940a,a30941a,a30944a,a30947a,a30948a,a30949a,a30952a,a30955a,a30956a,a30959a,a30962a,a30963a,a30964a,a30968a,a30969a,a30972a,a30975a,a30976a,a30977a,a30980a,a30983a,a30984a,a30987a,a30990a,a30991a,a30992a,a30996a,a30997a,a31000a,a31003a,a31004a,a31005a,a31008a,a31011a,a31012a,a31015a,a31018a,a31019a,a31020a,a31024a,a31025a,a31028a,a31031a,a31032a,a31033a,a31036a,a31039a,a31040a,a31043a,a31046a,a31047a,a31048a,a31052a,a31053a,a31056a,a31059a,a31060a,a31061a,a31064a,a31067a,a31068a,a31071a,a31074a,a31075a,a31076a,a31080a,a31081a,a31084a,a31087a,a31088a,a31089a,a31092a,a31095a,a31096a,a31099a,a31102a,a31103a,a31104a,a31108a,a31109a,a31112a,a31115a,a31116a,a31117a,a31120a,a31123a,a31124a,a31127a,a31130a,a31131a,a31132a,a31136a,a31137a,a31140a,a31143a,a31144a,a31145a,a31148a,a31151a,a31152a,a31155a,a31158a,a31159a,a31160a,a31164a,a31165a,a31168a,a31171a,a31172a,a31173a,a31176a,a31179a,a31180a,a31183a,a31186a,a31187a,a31188a,a31192a,a31193a,a31196a,a31199a,a31200a,a31201a,a31204a,a31207a,a31208a,a31211a,a31214a,a31215a,a31216a,a31220a,a31221a,a31224a,a31227a,a31228a,a31229a,a31232a,a31235a,a31236a,a31239a,a31242a,a31243a,a31244a,a31248a,a31249a,a31252a,a31255a,a31256a,a31257a,a31260a,a31263a,a31264a,a31267a,a31270a,a31271a,a31272a,a31276a,a31277a,a31280a,a31283a,a31284a,a31285a,a31288a,a31291a,a31292a,a31295a,a31298a,a31299a,a31300a,a31304a,a31305a,a31308a,a31311a,a31312a,a31313a,a31316a,a31319a,a31320a,a31323a,a31326a,a31327a,a31328a,a31332a,a31333a,a31336a,a31339a,a31340a,a31341a,a31344a,a31347a,a31348a,a31351a,a31354a,a31355a,a31356a,a31360a,a31361a,a31364a,a31367a,a31368a,a31369a,a31372a,a31375a,a31376a,a31379a,a31382a,a31383a,a31384a,a31388a,a31389a,a31392a,a31395a,a31396a,a31397a,a31400a,a31403a,a31404a,a31407a,a31410a,a31411a,a31412a,a31416a,a31417a,a31420a,a31423a,a31424a,a31425a,a31428a,a31431a,a31432a,a31435a,a31438a,a31439a,a31440a,a31444a,a31445a,a31448a,a31451a,a31452a,a31453a,a31456a,a31459a,a31460a,a31463a,a31466a,a31467a,a31468a,a31472a,a31473a,a31476a,a31479a,a31480a,a31481a,a31484a,a31487a,a31488a,a31491a,a31494a,a31495a,a31496a,a31500a,a31501a,a31504a,a31507a,a31508a,a31509a,a31512a,a31515a,a31516a,a31519a,a31522a,a31523a,a31524a,a31528a,a31529a,a31532a,a31535a,a31536a,a31537a,a31540a,a31543a,a31544a,a31547a,a31550a,a31551a,a31552a,a31556a,a31557a,a31560a,a31563a,a31564a,a31565a,a31568a,a31571a,a31572a,a31575a,a31578a,a31579a,a31580a,a31584a,a31585a,a31588a,a31591a,a31592a,a31593a,a31596a,a31599a,a31600a,a31603a,a31606a,a31607a,a31608a,a31612a,a31613a,a31616a,a31619a,a31620a,a31621a,a31624a,a31627a,a31628a,a31631a,a31634a,a31635a,a31636a,a31640a,a31641a,a31644a,a31647a,a31648a,a31649a,a31652a,a31655a,a31656a,a31659a,a31662a,a31663a,a31664a,a31668a,a31669a,a31672a,a31675a,a31676a,a31677a,a31680a,a31683a,a31684a,a31687a,a31690a,a31691a,a31692a,a31696a,a31697a,a31700a,a31703a,a31704a,a31705a,a31708a,a31711a,a31712a,a31715a,a31718a,a31719a,a31720a,a31724a,a31725a,a31728a,a31731a,a31732a,a31733a,a31736a,a31739a,a31740a,a31743a,a31746a,a31747a,a31748a,a31752a,a31753a,a31756a,a31759a,a31760a,a31761a,a31764a,a31767a,a31768a,a31771a,a31774a,a31775a,a31776a,a31780a,a31781a,a31784a,a31787a,a31788a,a31789a,a31792a,a31795a,a31796a,a31799a,a31802a,a31803a,a31804a,a31808a,a31809a,a31812a,a31815a,a31816a,a31817a,a31820a,a31823a,a31824a,a31827a,a31830a,a31831a,a31832a,a31836a,a31837a,a31840a,a31843a,a31844a,a31845a,a31848a,a31851a,a31852a,a31855a,a31858a,a31859a,a31860a,a31864a,a31865a,a31868a,a31871a,a31872a,a31873a,a31876a,a31879a,a31880a,a31883a,a31886a,a31887a,a31888a,a31892a,a31893a,a31896a,a31899a,a31900a,a31901a,a31904a,a31907a,a31908a,a31911a,a31914a,a31915a,a31916a,a31920a,a31921a,a31924a,a31927a,a31928a,a31929a,a31932a,a31935a,a31936a,a31939a,a31942a,a31943a,a31944a,a31948a,a31949a,a31952a,a31955a,a31956a,a31957a,a31960a,a31963a,a31964a,a31967a,a31970a,a31971a,a31972a,a31976a,a31977a,a31980a,a31983a,a31984a,a31985a,a31988a,a31991a,a31992a,a31995a,a31998a,a31999a,a32000a,a32004a,a32005a,a32008a,a32011a,a32012a,a32013a,a32016a,a32019a,a32020a,a32023a,a32026a,a32027a,a32028a,a32032a,a32033a,a32036a,a32039a,a32040a,a32041a,a32044a,a32047a,a32048a,a32051a,a32054a,a32055a,a32056a,a32060a,a32061a,a32064a,a32067a,a32068a,a32069a,a32072a,a32075a,a32076a,a32079a,a32082a,a32083a,a32084a,a32088a,a32089a,a32092a,a32095a,a32096a,a32097a,a32100a,a32103a,a32104a,a32107a,a32110a,a32111a,a32112a,a32116a,a32117a,a32120a,a32123a,a32124a,a32125a,a32128a,a32131a,a32132a,a32135a,a32138a,a32139a,a32140a,a32144a,a32145a,a32148a,a32151a,a32152a,a32153a,a32156a,a32159a,a32160a,a32163a,a32166a,a32167a,a32168a,a32172a,a32173a,a32176a,a32179a,a32180a,a32181a,a32184a,a32187a,a32188a,a32191a,a32194a,a32195a,a32196a,a32200a,a32201a,a32204a,a32207a,a32208a,a32209a,a32212a,a32215a,a32216a,a32219a,a32222a,a32223a,a32224a,a32228a,a32229a,a32232a,a32235a,a32236a,a32237a,a32240a,a32243a,a32244a,a32247a,a32250a,a32251a,a32252a,a32256a,a32257a,a32260a,a32263a,a32264a,a32265a,a32268a,a32271a,a32272a,a32275a,a32278a,a32279a,a32280a,a32284a,a32285a,a32288a,a32291a,a32292a,a32293a,a32296a,a32299a,a32300a,a32303a,a32306a,a32307a,a32308a,a32312a,a32313a,a32316a,a32319a,a32320a,a32321a,a32324a,a32327a,a32328a,a32331a,a32334a,a32335a,a32336a,a32340a,a32341a,a32344a,a32347a,a32348a,a32349a,a32352a,a32355a,a32356a,a32359a,a32362a,a32363a,a32364a,a32368a,a32369a,a32372a,a32375a,a32376a,a32377a,a32380a,a32383a,a32384a,a32387a,a32390a,a32391a,a32392a,a32396a,a32397a,a32400a,a32403a,a32404a,a32405a,a32408a,a32411a,a32412a,a32415a,a32418a,a32419a,a32420a,a32424a,a32425a,a32428a,a32431a,a32432a,a32433a,a32436a,a32439a,a32440a,a32443a,a32446a,a32447a,a32448a,a32452a,a32453a,a32456a,a32459a,a32460a,a32461a,a32464a,a32467a,a32468a,a32471a,a32474a,a32475a,a32476a,a32480a,a32481a,a32484a,a32487a,a32488a,a32489a,a32492a,a32495a,a32496a,a32499a,a32502a,a32503a,a32504a,a32508a,a32509a,a32512a,a32515a,a32516a,a32517a,a32520a,a32523a,a32524a,a32527a,a32530a,a32531a,a32532a,a32536a,a32537a,a32540a,a32543a,a32544a,a32545a,a32548a,a32551a,a32552a,a32555a,a32558a,a32559a,a32560a,a32564a,a32565a,a32568a,a32571a,a32572a,a32573a,a32576a,a32579a,a32580a,a32583a,a32586a,a32587a,a32588a,a32592a,a32593a,a32596a,a32599a,a32600a,a32601a,a32604a,a32607a,a32608a,a32611a,a32614a,a32615a,a32616a,a32620a,a32621a,a32624a,a32627a,a32628a,a32629a,a32632a,a32635a,a32636a,a32639a,a32642a,a32643a,a32644a,a32648a,a32649a,a32652a,a32655a,a32656a,a32657a,a32660a,a32663a,a32664a,a32667a,a32670a,a32671a,a32672a,a32676a,a32677a,a32680a,a32683a,a32684a,a32685a,a32688a,a32691a,a32692a,a32695a,a32698a,a32699a,a32700a,a32704a,a32705a,a32708a,a32711a,a32712a,a32713a,a32716a,a32719a,a32720a,a32723a,a32726a,a32727a,a32728a,a32732a,a32733a,a32736a,a32739a,a32740a,a32741a,a32744a,a32747a,a32748a,a32751a,a32754a,a32755a,a32756a,a32760a,a32761a,a32764a,a32767a,a32768a,a32769a,a32772a,a32775a,a32776a,a32779a,a32782a,a32783a,a32784a,a32788a,a32789a,a32792a,a32795a,a32796a,a32797a,a32800a,a32803a,a32804a,a32807a,a32810a,a32811a,a32812a,a32816a,a32817a,a32820a,a32823a,a32824a,a32825a,a32828a,a32831a,a32832a,a32835a,a32838a,a32839a,a32840a,a32844a,a32845a,a32848a,a32851a,a32852a,a32853a,a32856a,a32859a,a32860a,a32863a,a32866a,a32867a,a32868a,a32872a,a32873a,a32876a,a32879a,a32880a,a32881a,a32884a,a32887a,a32888a,a32891a,a32894a,a32895a,a32896a,a32900a,a32901a,a32904a,a32907a,a32908a,a32909a,a32912a,a32915a,a32916a,a32919a,a32922a,a32923a,a32924a,a32928a,a32929a,a32932a,a32935a,a32936a,a32937a,a32940a,a32943a,a32944a,a32947a,a32950a,a32951a,a32952a,a32956a,a32957a,a32960a,a32963a,a32964a,a32965a,a32968a,a32971a,a32972a,a32975a,a32978a,a32979a,a32980a,a32984a,a32985a,a32988a,a32991a,a32992a,a32993a,a32996a,a32999a,a33000a,a33003a,a33006a,a33007a,a33008a,a33012a,a33013a,a33016a,a33019a,a33020a,a33021a,a33024a,a33027a,a33028a,a33031a,a33034a,a33035a,a33036a,a33040a,a33041a,a33044a,a33047a,a33048a,a33049a,a33052a,a33055a,a33056a,a33059a,a33062a,a33063a,a33064a,a33068a,a33069a,a33072a,a33075a,a33076a,a33077a,a33080a,a33083a,a33084a,a33087a,a33090a,a33091a,a33092a,a33096a,a33097a,a33100a,a33103a,a33104a,a33105a,a33108a,a33111a,a33112a,a33115a,a33118a,a33119a,a33120a,a33124a,a33125a,a33128a,a33131a,a33132a,a33133a,a33136a,a33139a,a33140a,a33143a,a33146a,a33147a,a33148a,a33152a,a33153a,a33156a,a33159a,a33160a,a33161a,a33164a,a33167a,a33168a,a33171a,a33174a,a33175a,a33176a,a33180a,a33181a,a33184a,a33187a,a33188a,a33189a,a33192a,a33195a,a33196a,a33199a,a33202a,a33203a,a33204a,a33208a,a33209a,a33212a,a33215a,a33216a,a33217a,a33220a,a33223a,a33224a,a33227a,a33230a,a33231a,a33232a,a33236a,a33237a,a33240a,a33243a,a33244a,a33245a,a33248a,a33251a,a33252a,a33255a,a33258a,a33259a,a33260a,a33264a,a33265a,a33268a,a33271a,a33272a,a33273a,a33276a,a33279a,a33280a,a33283a,a33286a,a33287a,a33288a,a33292a,a33293a,a33296a,a33299a,a33300a,a33301a,a33304a,a33307a,a33308a,a33311a,a33314a,a33315a,a33316a,a33320a,a33321a,a33324a,a33327a,a33328a,a33329a,a33332a,a33335a,a33336a,a33339a,a33342a,a33343a,a33344a,a33348a,a33349a,a33352a,a33355a,a33356a,a33357a,a33360a,a33363a,a33364a,a33367a,a33370a,a33371a,a33372a,a33376a,a33377a,a33380a,a33383a,a33384a,a33385a,a33388a,a33391a,a33392a,a33395a,a33398a,a33399a,a33400a,a33404a,a33405a,a33408a,a33411a,a33412a,a33413a,a33416a,a33419a,a33420a,a33423a,a33426a,a33427a,a33428a,a33432a,a33433a,a33436a,a33439a,a33440a,a33441a,a33444a,a33447a,a33448a,a33451a,a33454a,a33455a,a33456a,a33460a,a33461a,a33464a,a33467a,a33468a,a33469a,a33472a,a33475a,a33476a,a33479a,a33482a,a33483a,a33484a,a33488a,a33489a,a33492a,a33495a,a33496a,a33497a,a33500a,a33503a,a33504a,a33507a,a33510a,a33511a,a33512a,a33516a,a33517a,a33520a,a33523a,a33524a,a33525a,a33528a,a33531a,a33532a,a33535a,a33538a,a33539a,a33540a,a33544a,a33545a,a33548a,a33551a,a33552a,a33553a,a33556a,a33559a,a33560a,a33563a,a33566a,a33567a,a33568a,a33572a,a33573a,a33576a,a33579a,a33580a,a33581a,a33584a,a33587a,a33588a,a33591a,a33594a,a33595a,a33596a,a33600a,a33601a,a33604a,a33607a,a33608a,a33609a,a33612a,a33615a,a33616a,a33619a,a33622a,a33623a,a33624a,a33628a,a33629a,a33632a,a33635a,a33636a,a33637a,a33640a,a33643a,a33644a,a33647a,a33650a,a33651a,a33652a,a33656a,a33657a,a33660a,a33663a,a33664a,a33665a,a33668a,a33671a,a33672a,a33675a,a33678a,a33679a,a33680a,a33684a,a33685a,a33688a,a33691a,a33692a,a33693a,a33696a,a33699a,a33700a,a33703a,a33706a,a33707a,a33708a,a33712a,a33713a,a33716a,a33719a,a33720a,a33721a,a33724a,a33727a,a33728a,a33731a,a33734a,a33735a,a33736a,a33740a,a33741a,a33744a,a33747a,a33748a,a33749a,a33752a,a33755a,a33756a,a33759a,a33762a,a33763a,a33764a,a33768a,a33769a,a33772a,a33775a,a33776a,a33777a,a33780a,a33783a,a33784a,a33787a,a33790a,a33791a,a33792a,a33796a,a33797a,a33800a,a33803a,a33804a,a33805a,a33808a,a33811a,a33812a,a33815a,a33818a,a33819a,a33820a,a33824a,a33825a,a33828a,a33831a,a33832a,a33833a,a33836a,a33839a,a33840a,a33843a,a33846a,a33847a,a33848a,a33852a,a33853a,a33856a,a33859a,a33860a,a33861a,a33864a,a33867a,a33868a,a33871a,a33874a,a33875a,a33876a,a33880a,a33881a,a33884a,a33887a,a33888a,a33889a,a33892a,a33895a,a33896a,a33899a,a33902a,a33903a,a33904a,a33908a,a33909a,a33912a,a33915a,a33916a,a33917a,a33920a,a33923a,a33924a,a33927a,a33930a,a33931a,a33932a,a33936a,a33937a,a33940a,a33943a,a33944a,a33945a,a33948a,a33951a,a33952a,a33955a,a33958a,a33959a,a33960a,a33964a,a33965a,a33968a,a33971a,a33972a,a33973a,a33976a,a33979a,a33980a,a33983a,a33986a,a33987a,a33988a,a33992a,a33993a,a33996a,a33999a,a34000a,a34001a,a34004a,a34007a,a34008a,a34011a,a34014a,a34015a,a34016a,a34020a,a34021a,a34024a,a34027a,a34028a,a34029a,a34032a,a34035a,a34036a,a34039a,a34042a,a34043a,a34044a,a34048a,a34049a,a34052a,a34055a,a34056a,a34057a,a34060a,a34063a,a34064a,a34067a,a34070a,a34071a,a34072a,a34076a,a34077a,a34080a,a34083a,a34084a,a34085a,a34088a,a34091a,a34092a,a34095a,a34098a,a34099a,a34100a,a34104a,a34105a,a34108a,a34111a,a34112a,a34113a,a34116a,a34119a,a34120a,a34123a,a34126a,a34127a,a34128a,a34132a,a34133a,a34136a,a34139a,a34140a,a34141a,a34144a,a34147a,a34148a,a34151a,a34154a,a34155a,a34156a,a34160a,a34161a,a34164a,a34167a,a34168a,a34169a,a34172a,a34175a,a34176a,a34179a,a34182a,a34183a,a34184a,a34188a,a34189a,a34192a,a34195a,a34196a,a34197a,a34200a,a34203a,a34204a,a34207a,a34210a,a34211a,a34212a,a34216a,a34217a,a34220a,a34223a,a34224a,a34225a,a34228a,a34231a,a34232a,a34235a,a34238a,a34239a,a34240a,a34244a,a34245a,a34248a,a34251a,a34252a,a34253a,a34256a,a34259a,a34260a,a34263a,a34266a,a34267a,a34268a,a34272a,a34273a,a34276a,a34279a,a34280a,a34281a,a34284a,a34287a,a34288a,a34291a,a34294a,a34295a,a34296a,a34300a,a34301a,a34304a,a34307a,a34308a,a34309a,a34312a,a34315a,a34316a,a34319a,a34322a,a34323a,a34324a,a34328a,a34329a,a34332a,a34335a,a34336a,a34337a,a34340a,a34343a,a34344a,a34347a,a34350a,a34351a,a34352a,a34356a,a34357a,a34360a,a34363a,a34364a,a34365a,a34368a,a34371a,a34372a,a34375a,a34378a,a34379a,a34380a,a34384a,a34385a,a34388a,a34391a,a34392a,a34393a,a34396a,a34399a,a34400a,a34403a,a34406a,a34407a,a34408a,a34412a,a34413a,a34416a,a34419a,a34420a,a34421a,a34424a,a34427a,a34428a,a34431a,a34434a,a34435a,a34436a,a34440a,a34441a,a34444a,a34447a,a34448a,a34449a,a34452a,a34455a,a34456a,a34459a,a34462a,a34463a,a34464a,a34468a,a34469a,a34472a,a34475a,a34476a,a34477a,a34480a,a34483a,a34484a,a34487a,a34490a,a34491a,a34492a,a34496a,a34497a,a34500a,a34503a,a34504a,a34505a,a34508a,a34511a,a34512a,a34515a,a34518a,a34519a,a34520a,a34524a,a34525a,a34528a,a34531a,a34532a,a34533a,a34536a,a34539a,a34540a,a34543a,a34546a,a34547a,a34548a,a34552a,a34553a,a34556a,a34559a,a34560a,a34561a,a34564a,a34567a,a34568a,a34571a,a34574a,a34575a,a34576a,a34580a,a34581a,a34584a,a34587a,a34588a,a34589a,a34592a,a34595a,a34596a,a34599a,a34602a,a34603a,a34604a,a34608a,a34609a,a34612a,a34615a,a34616a,a34617a,a34620a,a34623a,a34624a,a34627a,a34630a,a34631a,a34632a,a34636a,a34637a,a34640a,a34643a,a34644a,a34645a,a34648a,a34651a,a34652a,a34655a,a34658a,a34659a,a34660a,a34664a,a34665a,a34668a,a34671a,a34672a,a34673a,a34676a,a34679a,a34680a,a34683a,a34686a,a34687a,a34688a,a34692a,a34693a,a34696a,a34699a,a34700a,a34701a,a34704a,a34707a,a34708a,a34711a,a34714a,a34715a,a34716a,a34720a,a34721a,a34724a,a34727a,a34728a,a34729a,a34732a,a34735a,a34736a,a34739a,a34742a,a34743a,a34744a,a34748a,a34749a,a34752a,a34755a,a34756a,a34757a,a34760a,a34763a,a34764a,a34767a,a34770a,a34771a,a34772a,a34776a,a34777a,a34780a,a34783a,a34784a,a34785a,a34788a,a34791a,a34792a,a34795a,a34798a,a34799a,a34800a,a34804a,a34805a,a34808a,a34811a,a34812a,a34813a,a34816a,a34819a,a34820a,a34823a,a34826a,a34827a,a34828a,a34832a,a34833a,a34836a,a34839a,a34840a,a34841a,a34844a,a34847a,a34848a,a34851a,a34854a,a34855a,a34856a,a34860a,a34861a,a34864a,a34867a,a34868a,a34869a,a34872a,a34875a,a34876a,a34879a,a34882a,a34883a,a34884a,a34888a,a34889a,a34892a,a34895a,a34896a,a34897a,a34900a,a34903a,a34904a,a34907a,a34910a,a34911a,a34912a,a34916a,a34917a,a34920a,a34923a,a34924a,a34925a,a34928a,a34931a,a34932a,a34935a,a34938a,a34939a,a34940a,a34944a,a34945a,a34948a,a34951a,a34952a,a34953a,a34956a,a34959a,a34960a,a34963a,a34966a,a34967a,a34968a,a34972a,a34973a,a34976a,a34979a,a34980a,a34981a,a34984a,a34987a,a34988a,a34991a,a34994a,a34995a,a34996a,a35000a,a35001a,a35004a,a35007a,a35008a,a35009a,a35012a,a35015a,a35016a,a35019a,a35022a,a35023a,a35024a,a35028a,a35029a,a35032a,a35035a,a35036a,a35037a,a35040a,a35043a,a35044a,a35047a,a35050a,a35051a,a35052a,a35056a,a35057a,a35060a,a35063a,a35064a,a35065a,a35068a,a35071a,a35072a,a35075a,a35078a,a35079a,a35080a,a35084a,a35085a,a35088a,a35091a,a35092a,a35093a,a35096a,a35099a,a35100a,a35103a,a35106a,a35107a,a35108a,a35112a,a35113a,a35116a,a35119a,a35120a,a35121a,a35124a,a35127a,a35128a,a35131a,a35134a,a35135a,a35136a,a35140a,a35141a,a35144a,a35147a,a35148a,a35149a,a35152a,a35155a,a35156a,a35159a,a35162a,a35163a,a35164a,a35168a,a35169a,a35172a,a35175a,a35176a,a35177a,a35180a,a35183a,a35184a,a35187a,a35190a,a35191a,a35192a,a35196a,a35197a,a35200a,a35203a,a35204a,a35205a,a35208a,a35211a,a35212a,a35215a,a35218a,a35219a,a35220a,a35224a,a35225a,a35228a,a35231a,a35232a,a35233a,a35236a,a35239a,a35240a,a35243a,a35246a,a35247a,a35248a,a35252a,a35253a,a35256a,a35259a,a35260a,a35261a,a35264a,a35267a,a35268a,a35271a,a35274a,a35275a,a35276a,a35280a,a35281a,a35284a,a35287a,a35288a,a35289a,a35292a,a35295a,a35296a,a35299a,a35302a,a35303a,a35304a,a35308a,a35309a,a35312a,a35315a,a35316a,a35317a,a35320a,a35323a,a35324a,a35327a,a35330a,a35331a,a35332a,a35336a,a35337a,a35340a,a35343a,a35344a,a35345a,a35348a,a35351a,a35352a,a35355a,a35358a,a35359a,a35360a,a35364a,a35365a,a35368a,a35371a,a35372a,a35373a,a35376a,a35379a,a35380a,a35383a,a35386a,a35387a,a35388a,a35392a,a35393a,a35396a,a35399a,a35400a,a35401a,a35404a,a35407a,a35408a,a35411a,a35414a,a35415a,a35416a,a35420a,a35421a,a35424a,a35427a,a35428a,a35429a,a35432a,a35435a,a35436a,a35439a,a35442a,a35443a,a35444a,a35448a,a35449a,a35452a,a35455a,a35456a,a35457a,a35460a,a35463a,a35464a,a35467a,a35470a,a35471a,a35472a,a35476a,a35477a,a35480a,a35483a,a35484a,a35485a,a35488a,a35491a,a35492a,a35495a,a35498a,a35499a,a35500a,a35504a,a35505a,a35508a,a35511a,a35512a,a35513a,a35516a,a35519a,a35520a,a35523a,a35526a,a35527a,a35528a,a35532a,a35533a,a35536a,a35539a,a35540a,a35541a,a35544a,a35547a,a35548a,a35551a,a35554a,a35555a,a35556a,a35560a,a35561a,a35564a,a35567a,a35568a,a35569a,a35572a,a35575a,a35576a,a35579a,a35582a,a35583a,a35584a,a35588a,a35589a,a35592a,a35595a,a35596a,a35597a,a35600a,a35603a,a35604a,a35607a,a35610a,a35611a,a35612a,a35616a,a35617a,a35620a,a35623a,a35624a,a35625a,a35628a,a35631a,a35632a,a35635a,a35638a,a35639a,a35640a,a35644a,a35645a,a35648a,a35651a,a35652a,a35653a,a35656a,a35659a,a35660a,a35663a,a35666a,a35667a,a35668a,a35672a,a35673a,a35676a,a35679a,a35680a,a35681a,a35684a,a35687a,a35688a,a35691a,a35694a,a35695a,a35696a,a35700a,a35701a,a35704a,a35707a,a35708a,a35709a,a35712a,a35715a,a35716a,a35719a,a35722a,a35723a,a35724a,a35728a,a35729a,a35732a,a35735a,a35736a,a35737a,a35740a,a35743a,a35744a,a35747a,a35750a,a35751a,a35752a,a35756a,a35757a,a35760a,a35763a,a35764a,a35765a,a35768a,a35771a,a35772a,a35775a,a35778a,a35779a,a35780a,a35784a,a35785a,a35788a,a35791a,a35792a,a35793a,a35796a,a35799a,a35800a,a35803a,a35806a,a35807a,a35808a,a35812a,a35813a,a35816a,a35819a,a35820a,a35821a,a35824a,a35827a,a35828a,a35831a,a35834a,a35835a,a35836a,a35840a,a35841a,a35844a,a35847a,a35848a,a35849a,a35852a,a35855a,a35856a,a35859a,a35862a,a35863a,a35864a,a35868a,a35869a,a35872a,a35875a,a35876a,a35877a,a35880a,a35883a,a35884a,a35887a,a35890a,a35891a,a35892a,a35896a,a35897a,a35900a,a35903a,a35904a,a35905a,a35908a,a35911a,a35912a,a35915a,a35918a,a35919a,a35920a,a35924a,a35925a,a35928a,a35931a,a35932a,a35933a,a35936a,a35939a,a35940a,a35943a,a35946a,a35947a,a35948a,a35952a,a35953a,a35956a,a35959a,a35960a,a35961a,a35964a,a35967a,a35968a,a35971a,a35974a,a35975a,a35976a,a35980a,a35981a,a35984a,a35987a,a35988a,a35989a,a35992a,a35995a,a35996a,a35999a,a36002a,a36003a,a36004a,a36008a,a36009a,a36012a,a36015a,a36016a,a36017a,a36020a,a36023a,a36024a,a36027a,a36030a,a36031a,a36032a,a36036a,a36037a,a36040a,a36043a,a36044a,a36045a,a36048a,a36051a,a36052a,a36055a,a36058a,a36059a,a36060a,a36064a,a36065a,a36068a,a36071a,a36072a,a36073a,a36076a,a36079a,a36080a,a36083a,a36086a,a36087a,a36088a,a36092a,a36093a,a36096a,a36099a,a36100a,a36101a,a36104a,a36107a,a36108a,a36111a,a36114a,a36115a,a36116a,a36120a,a36121a,a36124a,a36127a,a36128a,a36129a,a36132a,a36135a,a36136a,a36139a,a36142a,a36143a,a36144a,a36148a,a36149a,a36152a,a36155a,a36156a,a36157a,a36160a,a36163a,a36164a,a36167a,a36170a,a36171a,a36172a,a36176a,a36177a,a36180a,a36183a,a36184a,a36185a,a36188a,a36191a,a36192a,a36195a,a36198a,a36199a,a36200a,a36204a,a36205a,a36208a,a36211a,a36212a,a36213a,a36216a,a36219a,a36220a,a36223a,a36226a,a36227a,a36228a,a36232a,a36233a,a36236a,a36239a,a36240a,a36241a,a36244a,a36247a,a36248a,a36251a,a36254a,a36255a,a36256a,a36260a,a36261a,a36264a,a36267a,a36268a,a36269a,a36272a,a36275a,a36276a,a36279a,a36282a,a36283a,a36284a,a36288a,a36289a,a36292a,a36295a,a36296a,a36297a,a36300a,a36303a,a36304a,a36307a,a36310a,a36311a,a36312a,a36316a,a36317a,a36320a,a36323a,a36324a,a36325a,a36328a,a36331a,a36332a,a36335a,a36338a,a36339a,a36340a,a36344a,a36345a,a36348a,a36351a,a36352a,a36353a,a36356a,a36359a,a36360a,a36363a,a36366a,a36367a,a36368a,a36372a,a36373a,a36376a,a36379a,a36380a,a36381a,a36384a,a36387a,a36388a,a36391a,a36394a,a36395a,a36396a,a36400a,a36401a,a36404a,a36407a,a36408a,a36409a,a36412a,a36415a,a36416a,a36419a,a36422a,a36423a,a36424a,a36428a,a36429a,a36432a,a36435a,a36436a,a36437a,a36440a,a36443a,a36444a,a36447a,a36450a,a36451a,a36452a,a36456a,a36457a,a36460a,a36463a,a36464a,a36465a,a36468a,a36471a,a36472a,a36475a,a36478a,a36479a,a36480a,a36484a,a36485a,a36488a,a36491a,a36492a,a36493a,a36496a,a36499a,a36500a,a36503a,a36506a,a36507a,a36508a,a36512a,a36513a,a36516a,a36519a,a36520a,a36521a,a36524a,a36527a,a36528a,a36531a,a36534a,a36535a,a36536a,a36540a,a36541a,a36544a,a36547a,a36548a,a36549a,a36552a,a36555a,a36556a,a36559a,a36562a,a36563a,a36564a,a36568a,a36569a,a36572a,a36575a,a36576a,a36577a,a36580a,a36583a,a36584a,a36587a,a36590a,a36591a,a36592a,a36596a,a36597a,a36600a,a36603a,a36604a,a36605a,a36608a,a36611a,a36612a,a36615a,a36618a,a36619a,a36620a,a36624a,a36625a,a36628a,a36631a,a36632a,a36633a,a36636a,a36639a,a36640a,a36643a,a36646a,a36647a,a36648a,a36652a,a36653a,a36656a,a36659a,a36660a,a36661a,a36664a,a36667a,a36668a,a36671a,a36674a,a36675a,a36676a,a36680a,a36681a,a36684a,a36687a,a36688a,a36689a,a36692a,a36695a,a36696a,a36699a,a36702a,a36703a,a36704a,a36708a,a36709a,a36712a,a36715a,a36716a,a36717a,a36720a,a36723a,a36724a,a36727a,a36730a,a36731a,a36732a,a36736a,a36737a,a36740a,a36743a,a36744a,a36745a,a36748a,a36751a,a36752a,a36755a,a36758a,a36759a,a36760a,a36764a,a36765a,a36768a,a36771a,a36772a,a36773a,a36776a,a36779a,a36780a,a36783a,a36786a,a36787a,a36788a,a36792a,a36793a,a36796a,a36799a,a36800a,a36801a,a36804a,a36807a,a36808a,a36811a,a36814a,a36815a,a36816a,a36820a,a36821a,a36824a,a36827a,a36828a,a36829a,a36832a,a36835a,a36836a,a36839a,a36842a,a36843a,a36844a,a36848a,a36849a,a36852a,a36855a,a36856a,a36857a,a36860a,a36863a,a36864a,a36867a,a36870a,a36871a,a36872a,a36876a,a36877a,a36880a,a36883a,a36884a,a36885a,a36888a,a36891a,a36892a,a36895a,a36898a,a36899a,a36900a,a36904a,a36905a,a36908a,a36911a,a36912a,a36913a,a36916a,a36919a,a36920a,a36923a,a36926a,a36927a,a36928a,a36932a,a36933a,a36936a,a36939a,a36940a,a36941a,a36944a,a36947a,a36948a,a36951a,a36954a,a36955a,a36956a,a36960a,a36961a,a36964a,a36967a,a36968a,a36969a,a36972a,a36975a,a36976a,a36979a,a36982a,a36983a,a36984a,a36988a,a36989a,a36992a,a36995a,a36996a,a36997a,a37000a,a37003a,a37004a,a37007a,a37010a,a37011a,a37012a,a37016a,a37017a,a37020a,a37023a,a37024a,a37025a,a37028a,a37031a,a37032a,a37035a,a37038a,a37039a,a37040a,a37044a,a37045a,a37048a,a37051a,a37052a,a37053a,a37056a,a37059a,a37060a,a37063a,a37066a,a37067a,a37068a,a37072a,a37073a,a37076a,a37079a,a37080a,a37081a,a37084a,a37087a,a37088a,a37091a,a37094a,a37095a,a37096a,a37100a,a37101a,a37104a,a37107a,a37108a,a37109a,a37112a,a37115a,a37116a,a37119a,a37122a,a37123a,a37124a,a37128a,a37129a,a37132a,a37135a,a37136a,a37137a,a37140a,a37143a,a37144a,a37147a,a37150a,a37151a,a37152a,a37156a,a37157a,a37160a,a37163a,a37164a,a37165a,a37168a,a37171a,a37172a,a37175a,a37178a,a37179a,a37180a,a37184a,a37185a,a37188a,a37191a,a37192a,a37193a,a37196a,a37199a,a37200a,a37203a,a37206a,a37207a,a37208a,a37212a,a37213a,a37216a,a37219a,a37220a,a37221a,a37224a,a37227a,a37228a,a37231a,a37234a,a37235a,a37236a,a37240a,a37241a,a37244a,a37247a,a37248a,a37249a,a37252a,a37255a,a37256a,a37259a,a37262a,a37263a,a37264a,a37268a,a37269a,a37272a,a37275a,a37276a,a37277a,a37280a,a37283a,a37284a,a37287a,a37290a,a37291a,a37292a,a37296a,a37297a,a37300a,a37303a,a37304a,a37305a,a37308a,a37311a,a37312a,a37315a,a37318a,a37319a,a37320a,a37324a,a37325a,a37328a,a37331a,a37332a,a37333a,a37336a,a37339a,a37340a,a37343a,a37346a,a37347a,a37348a,a37352a,a37353a,a37356a,a37359a,a37360a,a37361a,a37364a,a37367a,a37368a,a37371a,a37374a,a37375a,a37376a,a37380a,a37381a,a37384a,a37387a,a37388a,a37389a,a37392a,a37395a,a37396a,a37399a,a37402a,a37403a,a37404a,a37408a,a37409a,a37412a,a37415a,a37416a,a37417a,a37420a,a37423a,a37424a,a37427a,a37430a,a37431a,a37432a,a37436a,a37437a,a37440a,a37443a,a37444a,a37445a,a37448a,a37451a,a37452a,a37455a,a37458a,a37459a,a37460a,a37464a,a37465a,a37468a,a37471a,a37472a,a37473a,a37476a,a37479a,a37480a,a37483a,a37486a,a37487a,a37488a,a37492a,a37493a,a37496a,a37499a,a37500a,a37501a,a37504a,a37507a,a37508a,a37511a,a37514a,a37515a,a37516a,a37520a,a37521a,a37524a,a37527a,a37528a,a37529a,a37532a,a37535a,a37536a,a37539a,a37542a,a37543a,a37544a,a37548a,a37549a,a37552a,a37555a,a37556a,a37557a,a37560a,a37563a,a37564a,a37567a,a37570a,a37571a,a37572a,a37576a,a37577a,a37580a,a37583a,a37584a,a37585a,a37588a,a37591a,a37592a,a37595a,a37598a,a37599a,a37600a,a37604a,a37605a,a37608a,a37611a,a37612a,a37613a,a37616a,a37619a,a37620a,a37623a,a37626a,a37627a,a37628a,a37632a,a37633a,a37636a,a37639a,a37640a,a37641a,a37644a,a37647a,a37648a,a37651a,a37654a,a37655a,a37656a,a37660a,a37661a,a37664a,a37667a,a37668a,a37669a,a37672a,a37675a,a37676a,a37679a,a37682a,a37683a,a37684a,a37688a,a37689a,a37692a,a37695a,a37696a,a37697a,a37700a,a37703a,a37704a,a37707a,a37710a,a37711a,a37712a,a37716a,a37717a,a37720a,a37723a,a37724a,a37725a,a37728a,a37731a,a37732a,a37735a,a37738a,a37739a,a37740a,a37744a,a37745a,a37748a,a37751a,a37752a,a37753a,a37756a,a37759a,a37760a,a37763a,a37766a,a37767a,a37768a,a37772a,a37773a,a37776a,a37779a,a37780a,a37781a,a37784a,a37787a,a37788a,a37791a,a37794a,a37795a,a37796a,a37800a,a37801a,a37804a,a37807a,a37808a,a37809a,a37812a,a37815a,a37816a,a37819a,a37822a,a37823a,a37824a,a37828a,a37829a,a37832a,a37835a,a37836a,a37837a,a37840a,a37843a,a37844a,a37847a,a37850a,a37851a,a37852a,a37856a,a37857a,a37860a,a37863a,a37864a,a37865a,a37868a,a37871a,a37872a,a37875a,a37878a,a37879a,a37880a,a37884a,a37885a,a37888a,a37891a,a37892a,a37893a,a37896a,a37899a,a37900a,a37903a,a37906a,a37907a,a37908a,a37912a,a37913a,a37916a,a37919a,a37920a,a37921a,a37924a,a37927a,a37928a,a37931a,a37934a,a37935a,a37936a,a37940a,a37941a,a37944a,a37947a,a37948a,a37949a,a37952a,a37955a,a37956a,a37959a,a37962a,a37963a,a37964a,a37968a,a37969a,a37972a,a37975a,a37976a,a37977a,a37980a,a37983a,a37984a,a37987a,a37990a,a37991a,a37992a,a37996a,a37997a,a38000a,a38003a,a38004a,a38005a,a38008a,a38011a,a38012a,a38015a,a38018a,a38019a,a38020a,a38024a,a38025a,a38028a,a38031a,a38032a,a38033a,a38036a,a38039a,a38040a,a38043a,a38046a,a38047a,a38048a,a38052a,a38053a,a38056a,a38059a,a38060a,a38061a,a38064a,a38067a,a38068a,a38071a,a38074a,a38075a,a38076a,a38080a,a38081a,a38084a,a38087a,a38088a,a38089a,a38092a,a38095a,a38096a,a38099a,a38102a,a38103a,a38104a,a38108a,a38109a,a38112a,a38115a,a38116a,a38117a,a38120a,a38123a,a38124a,a38127a,a38130a,a38131a,a38132a,a38136a,a38137a,a38140a,a38143a,a38144a,a38145a,a38148a,a38151a,a38152a,a38155a,a38158a,a38159a,a38160a,a38164a,a38165a,a38168a,a38171a,a38172a,a38173a,a38176a,a38179a,a38180a,a38183a,a38186a,a38187a,a38188a,a38192a,a38193a,a38196a,a38199a,a38200a,a38201a,a38204a,a38207a,a38208a,a38211a,a38214a,a38215a,a38216a,a38220a,a38221a,a38224a,a38227a,a38228a,a38229a,a38232a,a38235a,a38236a,a38239a,a38242a,a38243a,a38244a,a38248a,a38249a,a38252a,a38255a,a38256a,a38257a,a38260a,a38263a,a38264a,a38267a,a38270a,a38271a,a38272a,a38276a,a38277a,a38280a,a38283a,a38284a,a38285a,a38288a,a38291a,a38292a,a38295a,a38298a,a38299a,a38300a,a38304a,a38305a,a38308a,a38311a,a38312a,a38313a,a38316a,a38319a,a38320a,a38323a,a38326a,a38327a,a38328a,a38332a,a38333a,a38336a,a38339a,a38340a,a38341a,a38344a,a38347a,a38348a,a38351a,a38354a,a38355a,a38356a,a38360a,a38361a,a38364a,a38367a,a38368a,a38369a,a38372a,a38375a,a38376a,a38379a,a38382a,a38383a,a38384a,a38388a,a38389a,a38392a,a38395a,a38396a,a38397a,a38400a,a38403a,a38404a,a38407a,a38410a,a38411a,a38412a,a38416a,a38417a,a38420a,a38423a,a38424a,a38425a,a38428a,a38431a,a38432a,a38435a,a38438a,a38439a,a38440a,a38444a,a38445a,a38448a,a38451a,a38452a,a38453a,a38456a,a38459a,a38460a,a38463a,a38466a,a38467a,a38468a,a38472a,a38473a,a38476a,a38479a,a38480a,a38481a,a38484a,a38487a,a38488a,a38491a,a38494a,a38495a,a38496a,a38500a,a38501a,a38504a,a38507a,a38508a,a38509a,a38512a,a38515a,a38516a,a38519a,a38522a,a38523a,a38524a,a38528a,a38529a,a38532a,a38535a,a38536a,a38537a,a38540a,a38543a,a38544a,a38547a,a38550a,a38551a,a38552a,a38556a,a38557a,a38560a,a38563a,a38564a,a38565a,a38568a,a38571a,a38572a,a38575a,a38578a,a38579a,a38580a,a38584a,a38585a,a38588a,a38591a,a38592a,a38593a,a38596a,a38599a,a38600a,a38603a,a38606a,a38607a,a38608a,a38612a,a38613a,a38616a,a38619a,a38620a,a38621a,a38624a,a38627a,a38628a,a38631a,a38634a,a38635a,a38636a,a38640a,a38641a,a38644a,a38647a,a38648a,a38649a,a38652a,a38655a,a38656a,a38659a,a38662a,a38663a,a38664a,a38668a,a38669a,a38672a,a38675a,a38676a,a38677a,a38680a,a38683a,a38684a,a38687a,a38690a,a38691a,a38692a,a38696a,a38697a,a38700a,a38703a,a38704a,a38705a,a38708a,a38711a,a38712a,a38715a,a38718a,a38719a,a38720a,a38724a,a38725a,a38728a,a38731a,a38732a,a38733a,a38736a,a38739a,a38740a,a38743a,a38746a,a38747a,a38748a,a38752a,a38753a,a38756a,a38759a,a38760a,a38761a,a38764a,a38767a,a38768a,a38771a,a38774a,a38775a,a38776a,a38780a,a38781a,a38784a,a38787a,a38788a,a38789a,a38792a,a38795a,a38796a,a38799a,a38802a,a38803a,a38804a,a38808a,a38809a,a38812a,a38815a,a38816a,a38817a,a38820a,a38823a,a38824a,a38827a,a38830a,a38831a,a38832a,a38836a,a38837a,a38840a,a38843a,a38844a,a38845a,a38848a,a38851a,a38852a,a38855a,a38858a,a38859a,a38860a,a38864a,a38865a,a38868a,a38871a,a38872a,a38873a,a38876a,a38879a,a38880a,a38883a,a38886a,a38887a,a38888a,a38892a,a38893a,a38896a,a38899a,a38900a,a38901a,a38904a,a38907a,a38908a,a38911a,a38914a,a38915a,a38916a,a38920a,a38921a,a38924a,a38927a,a38928a,a38929a,a38932a,a38935a,a38936a,a38939a,a38942a,a38943a,a38944a,a38948a,a38949a,a38952a,a38955a,a38956a,a38957a,a38960a,a38963a,a38964a,a38967a,a38970a,a38971a,a38972a,a38976a,a38977a,a38980a,a38983a,a38984a,a38985a,a38988a,a38991a,a38992a,a38995a,a38998a,a38999a,a39000a,a39004a,a39005a,a39008a,a39011a,a39012a,a39013a,a39016a,a39019a,a39020a,a39023a,a39026a,a39027a,a39028a,a39032a,a39033a,a39036a,a39039a,a39040a,a39041a,a39044a,a39047a,a39048a,a39051a,a39054a,a39055a,a39056a,a39060a,a39061a,a39064a,a39067a,a39068a,a39069a,a39072a,a39075a,a39076a,a39079a,a39082a,a39083a,a39084a,a39088a,a39089a,a39092a,a39095a,a39096a,a39097a,a39100a,a39103a,a39104a,a39107a,a39110a,a39111a,a39112a,a39116a,a39117a,a39120a,a39123a,a39124a,a39125a,a39128a,a39131a,a39132a,a39135a,a39138a,a39139a,a39140a,a39144a,a39145a,a39148a,a39151a,a39152a,a39153a,a39156a,a39159a,a39160a,a39163a,a39166a,a39167a,a39168a,a39172a,a39173a,a39176a,a39179a,a39180a,a39181a,a39184a,a39187a,a39188a,a39191a,a39194a,a39195a,a39196a,a39200a,a39201a,a39204a,a39207a,a39208a,a39209a,a39212a,a39215a,a39216a,a39219a,a39222a,a39223a,a39224a,a39228a,a39229a,a39232a,a39235a,a39236a,a39237a,a39240a,a39243a,a39244a,a39247a,a39250a,a39251a,a39252a,a39256a,a39257a,a39260a,a39263a,a39264a,a39265a,a39268a,a39271a,a39272a,a39275a,a39278a,a39279a,a39280a,a39284a,a39285a,a39288a,a39291a,a39292a,a39293a,a39296a,a39299a,a39300a,a39303a,a39306a,a39307a,a39308a,a39312a,a39313a,a39316a,a39319a,a39320a,a39321a,a39324a,a39327a,a39328a,a39331a,a39334a,a39335a,a39336a,a39340a,a39341a,a39344a,a39347a,a39348a,a39349a,a39352a,a39355a,a39356a,a39359a,a39362a,a39363a,a39364a,a39368a,a39369a,a39372a,a39375a,a39376a,a39377a,a39380a,a39383a,a39384a,a39387a,a39390a,a39391a,a39392a,a39396a,a39397a,a39400a,a39403a,a39404a,a39405a,a39408a,a39411a,a39412a,a39415a,a39418a,a39419a,a39420a,a39424a,a39425a,a39428a,a39431a,a39432a,a39433a,a39436a,a39439a,a39440a,a39443a,a39446a,a39447a,a39448a,a39452a,a39453a,a39456a,a39459a,a39460a,a39461a,a39464a,a39467a,a39468a,a39471a,a39474a,a39475a,a39476a,a39480a,a39481a,a39484a,a39487a,a39488a,a39489a,a39492a,a39495a,a39496a,a39499a,a39502a,a39503a,a39504a,a39508a,a39509a,a39512a,a39515a,a39516a,a39517a,a39520a,a39523a,a39524a,a39527a,a39530a,a39531a,a39532a,a39536a,a39537a,a39540a,a39543a,a39544a,a39545a,a39548a,a39551a,a39552a,a39555a,a39558a,a39559a,a39560a,a39564a,a39565a,a39568a,a39571a,a39572a,a39573a,a39576a,a39579a,a39580a,a39583a,a39586a,a39587a,a39588a,a39592a,a39593a,a39596a,a39599a,a39600a,a39601a,a39604a,a39607a,a39608a,a39611a,a39614a,a39615a,a39616a,a39620a,a39621a,a39624a,a39627a,a39628a,a39629a,a39632a,a39635a,a39636a,a39639a,a39642a,a39643a,a39644a,a39648a,a39649a,a39652a,a39655a,a39656a,a39657a,a39660a,a39663a,a39664a,a39667a,a39670a,a39671a,a39672a,a39676a,a39677a,a39680a,a39683a,a39684a,a39685a,a39688a,a39691a,a39692a,a39695a,a39698a,a39699a,a39700a,a39704a,a39705a,a39708a,a39711a,a39712a,a39713a,a39716a,a39719a,a39720a,a39723a,a39726a,a39727a,a39728a,a39732a,a39733a,a39736a,a39739a,a39740a,a39741a,a39744a,a39747a,a39748a,a39751a,a39754a,a39755a,a39756a,a39760a,a39761a,a39764a,a39767a,a39768a,a39769a,a39772a,a39775a,a39776a,a39779a,a39782a,a39783a,a39784a,a39788a,a39789a,a39792a,a39795a,a39796a,a39797a,a39800a,a39803a,a39804a,a39807a,a39810a,a39811a,a39812a,a39816a,a39817a,a39820a,a39823a,a39824a,a39825a,a39828a,a39831a,a39832a,a39835a,a39838a,a39839a,a39840a,a39844a,a39845a,a39848a,a39851a,a39852a,a39853a,a39856a,a39859a,a39860a,a39863a,a39866a,a39867a,a39868a,a39872a,a39873a,a39876a,a39879a,a39880a,a39881a,a39884a,a39887a,a39888a,a39891a,a39894a,a39895a,a39896a,a39900a,a39901a,a39904a,a39907a,a39908a,a39909a,a39912a,a39915a,a39916a,a39919a,a39922a,a39923a,a39924a,a39928a,a39929a,a39932a,a39935a,a39936a,a39937a,a39940a,a39943a,a39944a,a39947a,a39950a,a39951a,a39952a,a39956a,a39957a,a39960a,a39963a,a39964a,a39965a,a39968a,a39971a,a39972a,a39975a,a39978a,a39979a,a39980a,a39984a,a39985a,a39988a,a39991a,a39992a,a39993a,a39996a,a39999a,a40000a,a40003a,a40006a,a40007a,a40008a,a40012a,a40013a,a40016a,a40019a,a40020a,a40021a,a40024a,a40027a,a40028a,a40031a,a40034a,a40035a,a40036a,a40040a,a40041a,a40044a,a40047a,a40048a,a40049a,a40052a,a40055a,a40056a,a40059a,a40062a,a40063a,a40064a,a40068a,a40069a,a40072a,a40075a,a40076a,a40077a,a40080a,a40083a,a40084a,a40087a,a40090a,a40091a,a40092a,a40096a,a40097a,a40100a,a40103a,a40104a,a40105a,a40108a,a40111a,a40112a,a40115a,a40118a,a40119a,a40120a,a40124a,a40125a,a40128a,a40131a,a40132a,a40133a,a40136a,a40139a,a40140a,a40143a,a40146a,a40147a,a40148a,a40152a,a40153a,a40156a,a40159a,a40160a,a40161a,a40164a,a40167a,a40168a,a40171a,a40174a,a40175a,a40176a,a40180a,a40181a,a40184a,a40187a,a40188a,a40189a,a40192a,a40195a,a40196a,a40199a,a40202a,a40203a,a40204a,a40208a,a40209a,a40212a,a40215a,a40216a,a40217a,a40220a,a40223a,a40224a,a40227a,a40230a,a40231a,a40232a,a40236a,a40237a,a40240a,a40243a,a40244a,a40245a,a40248a,a40251a,a40252a,a40255a,a40258a,a40259a,a40260a,a40264a,a40265a,a40268a,a40271a,a40272a,a40273a,a40276a,a40279a,a40280a,a40283a,a40286a,a40287a,a40288a,a40292a,a40293a,a40296a,a40299a,a40300a,a40301a,a40304a,a40307a,a40308a,a40311a,a40314a,a40315a,a40316a,a40320a,a40321a,a40324a,a40327a,a40328a,a40329a,a40332a,a40335a,a40336a,a40339a,a40342a,a40343a,a40344a,a40348a,a40349a,a40352a,a40355a,a40356a,a40357a,a40360a,a40363a,a40364a,a40367a,a40370a,a40371a,a40372a,a40376a,a40377a,a40380a,a40383a,a40384a,a40385a,a40388a,a40391a,a40392a,a40395a,a40398a,a40399a,a40400a,a40404a,a40405a,a40408a,a40411a,a40412a,a40413a,a40416a,a40419a,a40420a,a40423a,a40426a,a40427a,a40428a,a40432a,a40433a,a40436a,a40439a,a40440a,a40441a,a40444a,a40447a,a40448a,a40451a,a40454a,a40455a,a40456a,a40460a,a40461a,a40464a,a40467a,a40468a,a40469a,a40472a,a40475a,a40476a,a40479a,a40482a,a40483a,a40484a,a40488a,a40489a,a40492a,a40495a,a40496a,a40497a,a40500a,a40503a,a40504a,a40507a,a40510a,a40511a,a40512a,a40516a,a40517a,a40520a,a40523a,a40524a,a40525a,a40528a,a40531a,a40532a,a40535a,a40538a,a40539a,a40540a,a40544a,a40545a,a40548a,a40551a,a40552a,a40553a,a40556a,a40559a,a40560a,a40563a,a40566a,a40567a,a40568a,a40572a,a40573a,a40576a,a40579a,a40580a,a40581a,a40584a,a40587a,a40588a,a40591a,a40594a,a40595a,a40596a,a40600a,a40601a,a40604a,a40607a,a40608a,a40609a,a40612a,a40615a,a40616a,a40619a,a40622a,a40623a,a40624a,a40628a,a40629a,a40632a,a40635a,a40636a,a40637a,a40640a,a40643a,a40644a,a40647a,a40650a,a40651a,a40652a,a40656a,a40657a,a40660a,a40663a,a40664a,a40665a,a40668a,a40671a,a40672a,a40675a,a40678a,a40679a,a40680a,a40684a,a40685a,a40688a,a40691a,a40692a,a40693a,a40696a,a40699a,a40700a,a40703a,a40706a,a40707a,a40708a,a40712a,a40713a,a40716a,a40719a,a40720a,a40721a,a40724a,a40727a,a40728a,a40731a,a40734a,a40735a,a40736a,a40740a,a40741a,a40744a,a40747a,a40748a,a40749a,a40752a,a40755a,a40756a,a40759a,a40762a,a40763a,a40764a,a40768a,a40769a,a40772a,a40775a,a40776a,a40777a,a40780a,a40783a,a40784a,a40787a,a40790a,a40791a,a40792a,a40796a,a40797a,a40800a,a40803a,a40804a,a40805a,a40808a,a40811a,a40812a,a40815a,a40818a,a40819a,a40820a,a40824a,a40825a,a40828a,a40831a,a40832a,a40833a,a40836a,a40839a,a40840a,a40843a,a40846a,a40847a,a40848a,a40852a,a40853a,a40856a,a40859a,a40860a,a40861a,a40864a,a40867a,a40868a,a40871a,a40874a,a40875a,a40876a,a40880a,a40881a,a40884a,a40887a,a40888a,a40889a,a40892a,a40895a,a40896a,a40899a,a40902a,a40903a,a40904a,a40908a,a40909a,a40912a,a40915a,a40916a,a40917a,a40920a,a40923a,a40924a,a40927a,a40930a,a40931a,a40932a,a40936a,a40937a,a40940a,a40943a,a40944a,a40945a,a40948a,a40951a,a40952a,a40955a,a40958a,a40959a,a40960a,a40964a,a40965a,a40968a,a40971a,a40972a,a40973a,a40976a,a40979a,a40980a,a40983a,a40986a,a40987a,a40988a,a40992a,a40993a,a40996a,a40999a,a41000a,a41001a,a41004a,a41007a,a41008a,a41011a,a41014a,a41015a,a41016a,a41020a,a41021a,a41024a,a41027a,a41028a,a41029a,a41032a,a41035a,a41036a,a41039a,a41042a,a41043a,a41044a,a41048a,a41049a,a41052a,a41055a,a41056a,a41057a,a41060a,a41063a,a41064a,a41067a,a41070a,a41071a,a41072a,a41076a,a41077a,a41080a,a41083a,a41084a,a41085a,a41088a,a41091a,a41092a,a41095a,a41098a,a41099a,a41100a,a41104a,a41105a,a41108a,a41111a,a41112a,a41113a,a41116a,a41119a,a41120a,a41123a,a41126a,a41127a,a41128a,a41132a,a41133a,a41136a,a41139a,a41140a,a41141a,a41144a,a41147a,a41148a,a41151a,a41154a,a41155a,a41156a,a41160a,a41161a,a41164a,a41167a,a41168a,a41169a,a41172a,a41175a,a41176a,a41179a,a41182a,a41183a,a41184a,a41188a,a41189a,a41192a,a41195a,a41196a,a41197a,a41200a,a41203a,a41204a,a41207a,a41210a,a41211a,a41212a,a41216a,a41217a,a41220a,a41223a,a41224a,a41225a,a41228a,a41231a,a41232a,a41235a,a41238a,a41239a,a41240a,a41244a,a41245a,a41248a,a41251a,a41252a,a41253a,a41256a,a41259a,a41260a,a41263a,a41266a,a41267a,a41268a,a41272a,a41273a,a41276a,a41279a,a41280a,a41281a,a41284a,a41287a,a41288a,a41291a,a41294a,a41295a,a41296a,a41300a,a41301a,a41304a,a41307a,a41308a,a41309a,a41312a,a41315a,a41316a,a41319a,a41322a,a41323a,a41324a,a41328a,a41329a,a41332a,a41335a,a41336a,a41337a,a41340a,a41343a,a41344a,a41347a,a41350a,a41351a,a41352a,a41356a,a41357a,a41360a,a41363a,a41364a,a41365a,a41368a,a41371a,a41372a,a41375a,a41378a,a41379a,a41380a,a41384a,a41385a,a41388a,a41391a,a41392a,a41393a,a41396a,a41399a,a41400a,a41403a,a41406a,a41407a,a41408a,a41412a,a41413a,a41416a,a41419a,a41420a,a41421a,a41424a,a41427a,a41428a,a41431a,a41434a,a41435a,a41436a,a41440a,a41441a,a41444a,a41447a,a41448a,a41449a,a41452a,a41455a,a41456a,a41459a,a41462a,a41463a,a41464a,a41468a,a41469a,a41472a,a41475a,a41476a,a41477a,a41480a,a41483a,a41484a,a41487a,a41490a,a41491a,a41492a,a41496a,a41497a,a41500a,a41503a,a41504a,a41505a,a41508a,a41511a,a41512a,a41515a,a41518a,a41519a,a41520a,a41524a,a41525a,a41528a,a41531a,a41532a,a41533a,a41536a,a41539a,a41540a,a41543a,a41546a,a41547a,a41548a,a41552a,a41553a,a41556a,a41559a,a41560a,a41561a,a41564a,a41567a,a41568a,a41571a,a41574a,a41575a,a41576a,a41580a,a41581a,a41584a,a41587a,a41588a,a41589a,a41592a,a41595a,a41596a,a41599a,a41602a,a41603a,a41604a,a41608a,a41609a,a41612a,a41615a,a41616a,a41617a,a41620a,a41623a,a41624a,a41627a,a41630a,a41631a,a41632a,a41636a,a41637a,a41640a,a41643a,a41644a,a41645a,a41648a,a41651a,a41652a,a41655a,a41658a,a41659a,a41660a,a41664a,a41665a,a41668a,a41671a,a41672a,a41673a,a41676a,a41679a,a41680a,a41683a,a41686a,a41687a,a41688a,a41692a,a41693a,a41696a,a41699a,a41700a,a41701a,a41704a,a41707a,a41708a,a41711a,a41714a,a41715a,a41716a,a41720a,a41721a,a41724a,a41727a,a41728a,a41729a,a41732a,a41735a,a41736a,a41739a,a41742a,a41743a,a41744a,a41748a,a41749a,a41752a,a41755a,a41756a,a41757a,a41760a,a41763a,a41764a,a41767a,a41770a,a41771a,a41772a,a41776a,a41777a,a41780a,a41783a,a41784a,a41785a,a41788a,a41791a,a41792a,a41795a,a41798a,a41799a,a41800a,a41804a,a41805a,a41808a,a41811a,a41812a,a41813a,a41816a,a41819a,a41820a,a41823a,a41826a,a41827a,a41828a,a41832a,a41833a,a41836a,a41839a,a41840a,a41841a,a41844a,a41847a,a41848a,a41851a,a41854a,a41855a,a41856a,a41860a,a41861a,a41864a,a41867a,a41868a,a41869a,a41872a,a41875a,a41876a,a41879a,a41882a,a41883a,a41884a,a41888a,a41889a,a41892a,a41895a,a41896a,a41897a,a41900a,a41903a,a41904a,a41907a,a41910a,a41911a,a41912a,a41916a,a41917a,a41920a,a41923a,a41924a,a41925a,a41928a,a41931a,a41932a,a41935a,a41938a,a41939a,a41940a,a41944a,a41945a,a41948a,a41951a,a41952a,a41953a,a41956a,a41959a,a41960a,a41963a,a41966a,a41967a,a41968a,a41972a,a41973a,a41976a,a41979a,a41980a,a41981a,a41984a,a41987a,a41988a,a41991a,a41994a,a41995a,a41996a,a42000a,a42001a,a42004a,a42007a,a42008a,a42009a,a42012a,a42015a,a42016a,a42019a,a42022a,a42023a,a42024a,a42028a,a42029a,a42032a,a42035a,a42036a,a42037a,a42040a,a42043a,a42044a,a42047a,a42050a,a42051a,a42052a,a42056a,a42057a,a42060a,a42063a,a42064a,a42065a,a42068a,a42071a,a42072a,a42075a,a42078a,a42079a,a42080a,a42084a,a42085a,a42088a,a42091a,a42092a,a42093a,a42096a,a42099a,a42100a,a42103a,a42106a,a42107a,a42108a,a42112a,a42113a,a42116a,a42119a,a42120a,a42121a,a42124a,a42127a,a42128a,a42131a,a42134a,a42135a,a42136a,a42140a,a42141a,a42144a,a42147a,a42148a,a42149a,a42152a,a42155a,a42156a,a42159a,a42162a,a42163a,a42164a,a42168a,a42169a,a42172a,a42175a,a42176a,a42177a,a42180a,a42183a,a42184a,a42187a,a42190a,a42191a,a42192a,a42196a,a42197a,a42200a,a42203a,a42204a,a42205a,a42208a,a42211a,a42212a,a42215a,a42218a,a42219a,a42220a,a42224a,a42225a,a42228a,a42231a,a42232a,a42233a,a42236a,a42239a,a42240a,a42243a,a42246a,a42247a,a42248a,a42252a,a42253a,a42256a,a42259a,a42260a,a42261a,a42264a,a42267a,a42268a,a42271a,a42274a,a42275a,a42276a,a42280a,a42281a,a42284a,a42287a,a42288a,a42289a,a42292a,a42295a,a42296a,a42299a,a42302a,a42303a,a42304a,a42308a,a42309a,a42312a,a42315a,a42316a,a42317a,a42320a,a42323a,a42324a,a42327a,a42330a,a42331a,a42332a,a42336a,a42337a,a42340a,a42343a,a42344a,a42345a,a42348a,a42351a,a42352a,a42355a,a42358a,a42359a,a42360a,a42364a,a42365a,a42368a,a42371a,a42372a,a42373a,a42376a,a42379a,a42380a,a42383a,a42386a,a42387a,a42388a,a42392a,a42393a,a42396a,a42399a,a42400a,a42401a,a42404a,a42407a,a42408a,a42411a,a42414a,a42415a,a42416a,a42420a,a42421a,a42424a,a42427a,a42428a,a42429a,a42432a,a42435a,a42436a,a42439a,a42442a,a42443a,a42444a,a42448a,a42449a,a42452a,a42455a,a42456a,a42457a,a42460a,a42463a,a42464a,a42467a,a42470a,a42471a,a42472a,a42476a,a42477a,a42480a,a42483a,a42484a,a42485a,a42488a,a42491a,a42492a,a42495a,a42498a,a42499a,a42500a,a42504a,a42505a,a42508a,a42511a,a42512a,a42513a,a42516a,a42519a,a42520a,a42523a,a42526a,a42527a,a42528a,a42532a,a42533a,a42536a,a42539a,a42540a,a42541a,a42544a,a42547a,a42548a,a42551a,a42554a,a42555a,a42556a,a42560a,a42561a,a42564a,a42567a,a42568a,a42569a,a42572a,a42575a,a42576a,a42579a,a42582a,a42583a,a42584a,a42588a,a42589a,a42592a,a42595a,a42596a,a42597a,a42600a,a42603a,a42604a,a42607a,a42610a,a42611a,a42612a,a42616a,a42617a,a42620a,a42623a,a42624a,a42625a,a42628a,a42631a,a42632a,a42635a,a42638a,a42639a,a42640a,a42644a,a42645a,a42648a,a42651a,a42652a,a42653a,a42656a,a42659a,a42660a,a42663a,a42666a,a42667a,a42668a,a42672a,a42673a,a42676a,a42679a,a42680a,a42681a,a42684a,a42687a,a42688a,a42691a,a42694a,a42695a,a42696a,a42700a,a42701a,a42704a,a42707a,a42708a,a42709a,a42712a,a42715a,a42716a,a42719a,a42722a,a42723a,a42724a,a42728a,a42729a,a42732a,a42735a,a42736a,a42737a,a42740a,a42743a,a42744a,a42747a,a42750a,a42751a,a42752a,a42756a,a42757a,a42760a,a42763a,a42764a,a42765a,a42768a,a42771a,a42772a,a42775a,a42778a,a42779a,a42780a,a42784a,a42785a,a42788a,a42791a,a42792a,a42793a,a42796a,a42799a,a42800a,a42803a,a42806a,a42807a,a42808a,a42812a,a42813a,a42816a,a42819a,a42820a,a42821a,a42824a,a42827a,a42828a,a42831a,a42834a,a42835a,a42836a,a42840a,a42841a,a42844a,a42847a,a42848a,a42849a,a42852a,a42855a,a42856a,a42859a,a42862a,a42863a,a42864a,a42868a,a42869a,a42872a,a42875a,a42876a,a42877a,a42880a,a42883a,a42884a,a42887a,a42890a,a42891a,a42892a,a42896a,a42897a,a42900a,a42903a,a42904a,a42905a,a42908a,a42911a,a42912a,a42915a,a42918a,a42919a,a42920a,a42924a,a42925a,a42928a,a42931a,a42932a,a42933a,a42936a,a42939a,a42940a,a42943a,a42946a,a42947a,a42948a,a42952a,a42953a,a42956a,a42959a,a42960a,a42961a,a42964a,a42967a,a42968a,a42971a,a42974a,a42975a,a42976a,a42980a,a42981a,a42984a,a42987a,a42988a,a42989a,a42992a,a42995a,a42996a,a42999a,a43002a,a43003a,a43004a,a43008a,a43009a,a43012a,a43015a,a43016a,a43017a,a43020a,a43023a,a43024a,a43027a,a43030a,a43031a,a43032a,a43036a,a43037a,a43040a,a43043a,a43044a,a43045a,a43048a,a43051a,a43052a,a43055a,a43058a,a43059a,a43060a,a43064a,a43065a,a43068a,a43071a,a43072a,a43073a,a43076a,a43079a,a43080a,a43083a,a43086a,a43087a,a43088a,a43092a,a43093a,a43096a,a43099a,a43100a,a43101a,a43104a,a43107a,a43108a,a43111a,a43114a,a43115a,a43116a,a43120a,a43121a,a43124a,a43127a,a43128a,a43129a,a43132a,a43135a,a43136a,a43139a,a43142a,a43143a,a43144a,a43148a,a43149a,a43152a,a43155a,a43156a,a43157a,a43160a,a43163a,a43164a,a43167a,a43170a,a43171a,a43172a,a43176a,a43177a,a43180a,a43183a,a43184a,a43185a,a43188a,a43191a,a43192a,a43195a,a43198a,a43199a,a43200a,a43204a,a43205a,a43208a,a43211a,a43212a,a43213a,a43216a,a43219a,a43220a,a43223a,a43226a,a43227a,a43228a,a43232a,a43233a,a43236a,a43239a,a43240a,a43241a,a43244a,a43247a,a43248a,a43251a,a43254a,a43255a,a43256a,a43260a,a43261a,a43264a,a43267a,a43268a,a43269a,a43272a,a43275a,a43276a,a43279a,a43282a,a43283a,a43284a,a43288a,a43289a,a43292a,a43295a,a43296a,a43297a,a43300a,a43303a,a43304a,a43307a,a43310a,a43311a,a43312a,a43316a,a43317a,a43320a,a43323a,a43324a,a43325a,a43328a,a43331a,a43332a,a43335a,a43338a,a43339a,a43340a,a43344a,a43345a,a43348a,a43351a,a43352a,a43353a,a43356a,a43359a,a43360a,a43363a,a43366a,a43367a,a43368a,a43372a,a43373a,a43376a,a43379a,a43380a,a43381a,a43384a,a43387a,a43388a,a43391a,a43394a,a43395a,a43396a,a43400a,a43401a,a43404a,a43407a,a43408a,a43409a,a43412a,a43415a,a43416a,a43419a,a43422a,a43423a,a43424a,a43428a,a43429a,a43432a,a43435a,a43436a,a43437a,a43440a,a43443a,a43444a,a43447a,a43450a,a43451a,a43452a,a43456a,a43457a,a43460a,a43463a,a43464a,a43465a,a43468a,a43471a,a43472a,a43475a,a43478a,a43479a,a43480a,a43484a,a43485a,a43488a,a43491a,a43492a,a43493a,a43496a,a43499a,a43500a,a43503a,a43506a,a43507a,a43508a,a43512a,a43513a,a43516a,a43519a,a43520a,a43521a,a43524a,a43527a,a43528a,a43531a,a43534a,a43535a,a43536a,a43540a,a43541a,a43544a,a43547a,a43548a,a43549a,a43552a,a43555a,a43556a,a43559a,a43562a,a43563a,a43564a,a43568a,a43569a,a43572a,a43575a,a43576a,a43577a,a43580a,a43583a,a43584a,a43587a,a43590a,a43591a,a43592a,a43596a,a43597a,a43600a,a43603a,a43604a,a43605a,a43608a,a43611a,a43612a,a43615a,a43618a,a43619a,a43620a,a43624a,a43625a,a43628a,a43631a,a43632a,a43633a,a43636a,a43639a,a43640a,a43643a,a43646a,a43647a,a43648a,a43652a,a43653a,a43656a,a43659a,a43660a,a43661a,a43664a,a43667a,a43668a,a43671a,a43674a,a43675a,a43676a,a43680a,a43681a,a43684a,a43687a,a43688a,a43689a,a43692a,a43695a,a43696a,a43699a,a43702a,a43703a,a43704a,a43708a,a43709a,a43712a,a43715a,a43716a,a43717a,a43720a,a43723a,a43724a,a43727a,a43730a,a43731a,a43732a,a43736a,a43737a,a43740a,a43743a,a43744a,a43745a,a43748a,a43751a,a43752a,a43755a,a43758a,a43759a,a43760a,a43764a,a43765a,a43768a,a43771a,a43772a,a43773a,a43776a,a43779a,a43780a,a43783a,a43786a,a43787a,a43788a,a43792a,a43793a,a43796a,a43799a,a43800a,a43801a,a43804a,a43807a,a43808a,a43811a,a43814a,a43815a,a43816a,a43820a,a43821a,a43824a,a43827a,a43828a,a43829a,a43832a,a43835a,a43836a,a43839a,a43842a,a43843a,a43844a,a43848a,a43849a,a43852a,a43855a,a43856a,a43857a,a43860a,a43863a,a43864a,a43867a,a43870a,a43871a,a43872a,a43876a,a43877a,a43880a,a43883a,a43884a,a43885a,a43888a,a43891a,a43892a,a43895a,a43898a,a43899a,a43900a,a43904a,a43905a,a43908a,a43911a,a43912a,a43913a,a43916a,a43919a,a43920a,a43923a,a43926a,a43927a,a43928a,a43932a,a43933a,a43936a,a43939a,a43940a,a43941a,a43944a,a43947a,a43948a,a43951a,a43954a,a43955a,a43956a,a43960a,a43961a,a43964a,a43967a,a43968a,a43969a,a43972a,a43975a,a43976a,a43979a,a43982a,a43983a,a43984a,a43988a,a43989a,a43992a,a43995a,a43996a,a43997a,a44000a,a44003a,a44004a,a44007a,a44010a,a44011a,a44012a,a44016a,a44017a,a44020a,a44023a,a44024a,a44025a,a44028a,a44031a,a44032a,a44035a,a44038a,a44039a,a44040a,a44044a,a44045a,a44048a,a44051a,a44052a,a44053a,a44056a,a44059a,a44060a,a44063a,a44066a,a44067a,a44068a,a44072a,a44073a,a44076a,a44079a,a44080a,a44081a,a44084a,a44087a,a44088a,a44091a,a44094a,a44095a,a44096a,a44100a,a44101a,a44104a,a44107a,a44108a,a44109a,a44112a,a44115a,a44116a,a44119a,a44122a,a44123a,a44124a,a44128a,a44129a,a44132a,a44135a,a44136a,a44137a,a44140a,a44143a,a44144a,a44147a,a44150a,a44151a,a44152a,a44156a,a44157a,a44160a,a44163a,a44164a,a44165a,a44168a,a44171a,a44172a,a44175a,a44178a,a44179a,a44180a,a44184a,a44185a,a44188a,a44191a,a44192a,a44193a,a44196a,a44199a,a44200a,a44203a,a44206a,a44207a,a44208a,a44212a,a44213a,a44216a,a44219a,a44220a,a44221a,a44224a,a44227a,a44228a,a44231a,a44234a,a44235a,a44236a,a44240a,a44241a,a44244a,a44247a,a44248a,a44249a,a44252a,a44255a,a44256a,a44259a,a44262a,a44263a,a44264a,a44268a,a44269a,a44272a,a44275a,a44276a,a44277a,a44280a,a44283a,a44284a,a44287a,a44290a,a44291a,a44292a,a44296a,a44297a,a44300a,a44303a,a44304a,a44305a,a44308a,a44311a,a44312a,a44315a,a44318a,a44319a,a44320a,a44324a,a44325a,a44328a,a44331a,a44332a,a44333a,a44336a,a44339a,a44340a,a44343a,a44346a,a44347a,a44348a,a44352a,a44353a,a44356a,a44359a,a44360a,a44361a,a44364a,a44367a,a44368a,a44371a,a44374a,a44375a,a44376a,a44380a,a44381a,a44384a,a44387a,a44388a,a44389a,a44392a,a44395a,a44396a,a44399a,a44402a,a44403a,a44404a,a44408a,a44409a,a44412a,a44415a,a44416a,a44417a,a44420a,a44423a,a44424a,a44427a,a44430a,a44431a,a44432a,a44436a,a44437a,a44440a,a44443a,a44444a,a44445a,a44448a,a44451a,a44452a,a44455a,a44458a,a44459a,a44460a,a44464a,a44465a,a44468a,a44471a,a44472a,a44473a,a44476a,a44479a,a44480a,a44483a,a44486a,a44487a,a44488a,a44492a,a44493a,a44496a,a44499a,a44500a,a44501a,a44504a,a44507a,a44508a,a44511a,a44514a,a44515a,a44516a,a44520a,a44521a,a44524a,a44527a,a44528a,a44529a,a44532a,a44535a,a44536a,a44539a,a44542a,a44543a,a44544a,a44548a,a44549a,a44552a,a44555a,a44556a,a44557a,a44560a,a44563a,a44564a,a44567a,a44570a,a44571a,a44572a,a44576a,a44577a,a44580a,a44583a,a44584a,a44585a,a44588a,a44591a,a44592a,a44595a,a44598a,a44599a,a44600a,a44604a,a44605a,a44608a,a44611a,a44612a,a44613a,a44616a,a44619a,a44620a,a44623a,a44626a,a44627a,a44628a,a44632a,a44633a,a44636a,a44639a,a44640a,a44641a,a44644a,a44647a,a44648a,a44651a,a44654a,a44655a,a44656a,a44660a,a44661a,a44664a,a44667a,a44668a,a44669a,a44672a,a44675a,a44676a,a44679a,a44682a,a44683a,a44684a,a44688a,a44689a,a44692a,a44695a,a44696a,a44697a,a44700a,a44703a,a44704a,a44707a,a44710a,a44711a,a44712a,a44716a,a44717a,a44720a,a44723a,a44724a,a44725a,a44728a,a44731a,a44732a,a44735a,a44738a,a44739a,a44740a,a44744a,a44745a,a44748a,a44751a,a44752a,a44753a,a44756a,a44759a,a44760a,a44763a,a44766a,a44767a,a44768a,a44772a,a44773a,a44776a,a44779a,a44780a,a44781a,a44784a,a44787a,a44788a,a44791a,a44794a,a44795a,a44796a,a44800a,a44801a,a44804a,a44807a,a44808a,a44809a,a44812a,a44815a,a44816a,a44819a,a44822a,a44823a,a44824a,a44828a,a44829a,a44832a,a44835a,a44836a,a44837a,a44840a,a44843a,a44844a,a44847a,a44850a,a44851a,a44852a,a44856a,a44857a,a44860a,a44863a,a44864a,a44865a,a44868a,a44871a,a44872a,a44875a,a44878a,a44879a,a44880a,a44884a,a44885a,a44888a,a44891a,a44892a,a44893a,a44896a,a44899a,a44900a,a44903a,a44906a,a44907a,a44908a,a44912a,a44913a,a44916a,a44919a,a44920a,a44921a,a44924a,a44927a,a44928a,a44931a,a44934a,a44935a,a44936a,a44940a,a44941a,a44944a,a44947a,a44948a,a44949a,a44952a,a44955a,a44956a,a44959a,a44962a,a44963a,a44964a,a44968a,a44969a,a44972a,a44975a,a44976a,a44977a,a44980a,a44983a,a44984a,a44987a,a44990a,a44991a,a44992a,a44996a,a44997a,a45000a,a45003a,a45004a,a45005a,a45008a,a45011a,a45012a,a45015a,a45018a,a45019a,a45020a,a45024a,a45025a,a45028a,a45031a,a45032a,a45033a,a45036a,a45039a,a45040a,a45043a,a45046a,a45047a,a45048a,a45052a,a45053a,a45056a,a45059a,a45060a,a45061a,a45064a,a45067a,a45068a,a45071a,a45074a,a45075a,a45076a,a45080a,a45081a,a45084a,a45087a,a45088a,a45089a,a45092a,a45095a,a45096a,a45099a,a45102a,a45103a,a45104a,a45108a,a45109a,a45112a,a45115a,a45116a,a45117a,a45120a,a45123a,a45124a,a45127a,a45130a,a45131a,a45132a,a45136a,a45137a,a45140a,a45143a,a45144a,a45145a,a45148a,a45151a,a45152a,a45155a,a45158a,a45159a,a45160a,a45164a,a45165a,a45168a,a45171a,a45172a,a45173a,a45176a,a45179a,a45180a,a45183a,a45186a,a45187a,a45188a,a45192a,a45193a,a45196a,a45199a,a45200a,a45201a,a45204a,a45207a,a45208a,a45211a,a45214a,a45215a,a45216a,a45220a,a45221a,a45224a,a45227a,a45228a,a45229a,a45232a,a45235a,a45236a,a45239a,a45242a,a45243a,a45244a,a45248a,a45249a,a45252a,a45255a,a45256a,a45257a,a45260a,a45263a,a45264a,a45267a,a45270a,a45271a,a45272a,a45276a,a45277a,a45280a,a45283a,a45284a,a45285a,a45288a,a45291a,a45292a,a45295a,a45298a,a45299a,a45300a,a45303a,a45306a,a45307a,a45310a,a45313a,a45314a,a45315a,a45318a,a45321a,a45322a,a45325a,a45328a,a45329a,a45330a,a45333a,a45336a,a45337a,a45340a,a45343a,a45344a,a45345a,a45348a,a45351a,a45352a,a45355a,a45358a,a45359a,a45360a,a45363a,a45366a,a45367a,a45370a,a45373a,a45374a,a45375a,a45378a,a45381a,a45382a,a45385a,a45388a,a45389a,a45390a,a45393a,a45396a,a45397a,a45400a,a45403a,a45404a,a45405a,a45408a,a45411a,a45412a,a45415a,a45418a,a45419a,a45420a,a45423a,a45426a,a45427a,a45430a,a45433a,a45434a,a45435a,a45438a,a45441a,a45442a,a45445a,a45448a,a45449a,a45450a,a45453a,a45456a,a45457a,a45460a,a45463a,a45464a,a45465a,a45468a,a45471a,a45472a,a45475a,a45478a,a45479a,a45480a,a45483a,a45486a,a45487a,a45490a,a45493a,a45494a,a45495a,a45498a,a45501a,a45502a,a45505a,a45508a,a45509a,a45510a,a45513a,a45516a,a45517a,a45520a,a45523a,a45524a,a45525a,a45528a,a45531a,a45532a,a45535a,a45538a,a45539a,a45540a,a45543a,a45546a,a45547a,a45550a,a45553a,a45554a,a45555a,a45558a,a45561a,a45562a,a45565a,a45568a,a45569a,a45570a,a45573a,a45576a,a45577a,a45580a,a45583a,a45584a,a45585a,a45588a,a45591a,a45592a,a45595a,a45598a,a45599a,a45600a,a45603a,a45606a,a45607a,a45610a,a45613a,a45614a,a45615a,a45618a,a45621a,a45622a,a45625a,a45628a,a45629a,a45630a,a45633a,a45636a,a45637a,a45640a,a45643a,a45644a,a45645a,a45648a,a45651a,a45652a,a45655a,a45658a,a45659a,a45660a,a45663a,a45666a,a45667a,a45670a,a45673a,a45674a,a45675a,a45678a,a45681a,a45682a,a45685a,a45688a,a45689a,a45690a,a45693a,a45696a,a45697a,a45700a,a45703a,a45704a,a45705a,a45708a,a45711a,a45712a,a45715a,a45718a,a45719a,a45720a,a45723a,a45726a,a45727a,a45730a,a45733a,a45734a,a45735a,a45738a,a45741a,a45742a,a45745a,a45748a,a45749a,a45750a,a45753a,a45756a,a45757a,a45760a,a45763a,a45764a,a45765a,a45768a,a45771a,a45772a,a45775a,a45778a,a45779a,a45780a,a45783a,a45786a,a45787a,a45790a,a45793a,a45794a,a45795a,a45798a,a45801a,a45802a,a45805a,a45808a,a45809a,a45810a,a45813a,a45816a,a45817a,a45820a,a45823a,a45824a,a45825a,a45828a,a45831a,a45832a,a45835a,a45838a,a45839a,a45840a,a45843a,a45846a,a45847a,a45850a,a45853a,a45854a,a45855a,a45858a,a45861a,a45862a,a45865a,a45868a,a45869a,a45870a,a45873a,a45876a,a45877a,a45880a,a45883a,a45884a,a45885a,a45888a,a45891a,a45892a,a45895a,a45898a,a45899a,a45900a,a45903a,a45906a,a45907a,a45910a,a45913a,a45914a,a45915a,a45918a,a45921a,a45922a,a45925a,a45928a,a45929a,a45930a,a45933a,a45936a,a45937a,a45940a,a45943a,a45944a,a45945a,a45948a,a45951a,a45952a,a45955a,a45958a,a45959a,a45960a,a45963a,a45966a,a45967a,a45970a,a45973a,a45974a,a45975a,a45978a,a45981a,a45982a,a45985a,a45988a,a45989a,a45990a,a45993a,a45996a,a45997a,a46000a,a46003a,a46004a,a46005a,a46008a,a46011a,a46012a,a46015a,a46018a,a46019a,a46020a,a46023a,a46026a,a46027a,a46030a,a46033a,a46034a,a46035a,a46038a,a46041a,a46042a,a46045a,a46048a,a46049a,a46050a,a46053a,a46056a,a46057a,a46060a,a46063a,a46064a,a46065a,a46068a,a46071a,a46072a,a46075a,a46078a,a46079a,a46080a,a46083a,a46086a,a46087a,a46090a,a46093a,a46094a,a46095a,a46098a,a46101a,a46102a,a46105a,a46108a,a46109a,a46110a,a46113a,a46116a,a46117a,a46120a,a46123a,a46124a,a46125a,a46128a,a46131a,a46132a,a46135a,a46138a,a46139a,a46140a,a46143a,a46146a,a46147a,a46150a,a46153a,a46154a,a46155a,a46158a,a46161a,a46162a,a46165a,a46168a,a46169a,a46170a,a46173a,a46176a,a46177a,a46180a,a46183a,a46184a,a46185a,a46188a,a46191a,a46192a,a46195a,a46198a,a46199a,a46200a,a46203a,a46206a,a46207a,a46210a,a46213a,a46214a,a46215a,a46218a,a46221a,a46222a,a46225a,a46228a,a46229a,a46230a,a46233a,a46236a,a46237a,a46240a,a46243a,a46244a,a46245a,a46248a,a46251a,a46252a,a46255a,a46258a,a46259a,a46260a,a46263a,a46266a,a46267a,a46270a,a46273a,a46274a,a46275a,a46278a,a46281a,a46282a,a46285a,a46288a,a46289a,a46290a,a46293a,a46296a,a46297a,a46300a,a46303a,a46304a,a46305a,a46308a,a46311a,a46312a,a46315a,a46318a,a46319a,a46320a,a46323a,a46326a,a46327a,a46330a,a46333a,a46334a,a46335a,a46338a,a46341a,a46342a,a46345a,a46348a,a46349a,a46350a,a46353a,a46356a,a46357a,a46360a,a46363a,a46364a,a46365a,a46368a,a46371a,a46372a,a46375a,a46378a,a46379a,a46380a,a46383a,a46386a,a46387a,a46390a,a46393a,a46394a,a46395a,a46398a,a46401a,a46402a,a46405a,a46408a,a46409a,a46410a,a46413a,a46416a,a46417a,a46420a,a46423a,a46424a,a46425a,a46428a,a46431a,a46432a,a46435a,a46438a,a46439a,a46440a,a46443a,a46446a,a46447a,a46450a,a46453a,a46454a,a46455a,a46458a,a46461a,a46462a,a46465a,a46468a,a46469a,a46470a,a46473a,a46476a,a46477a,a46480a,a46483a,a46484a,a46485a,a46488a,a46491a,a46492a,a46495a,a46498a,a46499a,a46500a,a46503a,a46506a,a46507a,a46510a,a46513a,a46514a,a46515a,a46518a,a46521a,a46522a,a46525a,a46528a,a46529a,a46530a,a46533a,a46536a,a46537a,a46540a,a46543a,a46544a,a46545a,a46548a,a46551a,a46552a,a46555a,a46558a,a46559a,a46560a,a46563a,a46566a,a46567a,a46570a,a46573a,a46574a,a46575a,a46578a,a46581a,a46582a,a46585a,a46588a,a46589a,a46590a,a46593a,a46596a,a46597a,a46600a,a46603a,a46604a,a46605a,a46608a,a46611a,a46612a,a46615a,a46618a,a46619a,a46620a,a46623a,a46626a,a46627a,a46630a,a46633a,a46634a,a46635a,a46638a,a46641a,a46642a,a46645a,a46648a,a46649a,a46650a,a46653a,a46656a,a46657a,a46660a,a46663a,a46664a,a46665a,a46668a,a46671a,a46672a,a46675a,a46678a,a46679a,a46680a,a46683a,a46686a,a46687a,a46690a,a46693a,a46694a,a46695a,a46698a,a46701a,a46702a,a46705a,a46708a,a46709a,a46710a,a46713a,a46716a,a46717a,a46720a,a46723a,a46724a,a46725a,a46728a,a46731a,a46732a,a46735a,a46738a,a46739a,a46740a,a46743a,a46746a,a46747a,a46750a,a46753a,a46754a,a46755a,a46758a,a46761a,a46762a,a46765a,a46768a,a46769a,a46770a,a46773a,a46776a,a46777a,a46780a,a46783a,a46784a,a46785a,a46788a,a46791a,a46792a,a46795a,a46798a,a46799a,a46800a,a46803a,a46806a,a46807a,a46810a,a46813a,a46814a,a46815a,a46818a,a46821a,a46822a,a46825a,a46828a,a46829a,a46830a,a46833a,a46836a,a46837a,a46840a,a46843a,a46844a,a46845a,a46848a,a46851a,a46852a,a46855a,a46858a,a46859a,a46860a,a46863a,a46866a,a46867a,a46870a,a46873a,a46874a,a46875a,a46878a,a46881a,a46882a,a46885a,a46888a,a46889a,a46890a,a46893a,a46896a,a46897a,a46900a,a46903a,a46904a,a46905a,a46908a,a46911a,a46912a,a46915a,a46918a,a46919a,a46920a,a46923a,a46926a,a46927a,a46930a,a46933a,a46934a,a46935a,a46938a,a46941a,a46942a,a46945a,a46948a,a46949a,a46950a,a46953a,a46956a,a46957a,a46960a,a46963a,a46964a,a46965a,a46968a,a46971a,a46972a,a46975a,a46978a,a46979a,a46980a,a46983a,a46986a,a46987a,a46990a,a46993a,a46994a,a46995a,a46998a,a47001a,a47002a,a47005a,a47008a,a47009a,a47010a,a47013a,a47016a,a47017a,a47020a,a47023a,a47024a,a47025a,a47028a,a47031a,a47032a,a47035a,a47038a,a47039a,a47040a,a47043a,a47046a,a47047a,a47050a,a47053a,a47054a,a47055a,a47058a,a47061a,a47062a,a47065a,a47068a,a47069a,a47070a,a47073a,a47076a,a47077a,a47080a,a47083a,a47084a,a47085a,a47088a,a47091a,a47092a,a47095a,a47098a,a47099a,a47100a,a47103a,a47106a,a47107a,a47110a,a47113a,a47114a,a47115a,a47118a,a47121a,a47122a,a47125a,a47128a,a47129a,a47130a,a47133a,a47136a,a47137a,a47140a,a47143a,a47144a,a47145a,a47148a,a47151a,a47152a,a47155a,a47158a,a47159a,a47160a,a47163a,a47166a,a47167a,a47170a,a47173a,a47174a,a47175a,a47178a,a47181a,a47182a,a47185a,a47188a,a47189a,a47190a,a47193a,a47196a,a47197a,a47200a,a47203a,a47204a,a47205a,a47208a,a47211a,a47212a,a47215a,a47218a,a47219a,a47220a,a47223a,a47226a,a47227a,a47230a,a47233a,a47234a,a47235a,a47238a,a47241a,a47242a,a47245a,a47248a,a47249a,a47250a,a47253a,a47256a,a47257a,a47260a,a47263a,a47264a,a47265a,a47268a,a47271a,a47272a,a47275a,a47278a,a47279a,a47280a,a47283a,a47286a,a47287a,a47290a,a47293a,a47294a,a47295a,a47298a,a47301a,a47302a,a47305a,a47308a,a47309a,a47310a,a47313a,a47316a,a47317a,a47320a,a47323a,a47324a,a47325a,a47328a,a47331a,a47332a,a47335a,a47338a,a47339a,a47340a,a47343a,a47346a,a47347a,a47350a,a47353a,a47354a,a47355a,a47358a,a47361a,a47362a,a47365a,a47368a,a47369a,a47370a,a47373a,a47376a,a47377a,a47380a,a47383a,a47384a,a47385a,a47388a,a47391a,a47392a,a47395a,a47398a,a47399a,a47400a,a47403a,a47406a,a47407a,a47410a,a47413a,a47414a,a47415a,a47418a,a47421a,a47422a,a47425a,a47428a,a47429a,a47430a,a47433a,a47436a,a47437a,a47440a,a47443a,a47444a,a47445a,a47448a,a47451a,a47452a,a47455a,a47458a,a47459a,a47460a,a47463a,a47466a,a47467a,a47470a,a47473a,a47474a,a47475a,a47478a,a47481a,a47482a,a47485a,a47488a,a47489a,a47490a,a47493a,a47496a,a47497a,a47500a,a47503a,a47504a,a47505a,a47508a,a47511a,a47512a,a47515a,a47518a,a47519a,a47520a,a47523a,a47526a,a47527a,a47530a,a47533a,a47534a,a47535a,a47538a,a47541a,a47542a,a47545a,a47548a,a47549a,a47550a,a47553a,a47556a,a47557a,a47560a,a47563a,a47564a,a47565a,a47568a,a47571a,a47572a,a47575a,a47578a,a47579a,a47580a,a47583a,a47586a,a47587a,a47590a,a47593a,a47594a,a47595a,a47598a,a47601a,a47602a,a47605a,a47608a,a47609a,a47610a,a47613a,a47616a,a47617a,a47620a,a47623a,a47624a,a47625a,a47628a,a47631a,a47632a,a47635a,a47638a,a47639a,a47640a,a47643a,a47646a,a47647a,a47650a,a47653a,a47654a,a47655a,a47658a,a47661a,a47662a,a47665a,a47668a,a47669a,a47670a,a47673a,a47676a,a47677a,a47680a,a47683a,a47684a,a47685a,a47688a,a47691a,a47692a,a47695a,a47698a,a47699a,a47700a,a47703a,a47706a,a47707a,a47710a,a47713a,a47714a,a47715a,a47718a,a47721a,a47722a,a47725a,a47728a,a47729a,a47730a,a47733a,a47736a,a47737a,a47740a,a47743a,a47744a,a47745a,a47748a,a47751a,a47752a,a47755a,a47758a,a47759a,a47760a,a47763a,a47766a,a47767a,a47770a,a47773a,a47774a,a47775a,a47778a,a47781a,a47782a,a47785a,a47788a,a47789a,a47790a,a47793a,a47796a,a47797a,a47800a,a47803a,a47804a,a47805a,a47808a,a47811a,a47812a,a47815a,a47818a,a47819a,a47820a,a47823a,a47826a,a47827a,a47830a,a47833a,a47834a,a47835a,a47838a,a47841a,a47842a,a47845a,a47848a,a47849a,a47850a,a47853a,a47856a,a47857a,a47860a,a47863a,a47864a,a47865a,a47868a,a47871a,a47872a,a47875a,a47878a,a47879a,a47880a,a47883a,a47886a,a47887a,a47890a,a47893a,a47894a,a47895a,a47898a,a47901a,a47902a,a47905a,a47908a,a47909a,a47910a,a47913a,a47916a,a47917a,a47920a,a47923a,a47924a,a47925a,a47928a,a47931a,a47932a,a47935a,a47938a,a47939a,a47940a,a47943a,a47946a,a47947a,a47950a,a47953a,a47954a,a47955a,a47958a,a47961a,a47962a,a47965a,a47968a,a47969a,a47970a,a47973a,a47976a,a47977a,a47980a,a47983a,a47984a,a47985a,a47988a,a47991a,a47992a,a47995a,a47998a,a47999a,a48000a,a48003a,a48006a,a48007a,a48010a,a48013a,a48014a,a48015a,a48018a,a48021a,a48022a,a48025a,a48028a,a48029a,a48030a,a48033a,a48036a,a48037a,a48040a,a48043a,a48044a,a48045a,a48048a,a48051a,a48052a,a48055a,a48058a,a48059a,a48060a,a48063a,a48066a,a48067a,a48070a,a48073a,a48074a,a48075a,a48078a,a48081a,a48082a,a48085a,a48088a,a48089a,a48090a,a48093a,a48096a,a48097a,a48100a,a48103a,a48104a,a48105a,a48108a,a48111a,a48112a,a48115a,a48118a,a48119a,a48120a,a48123a,a48126a,a48127a,a48130a,a48133a,a48134a,a48135a,a48138a,a48141a,a48142a,a48145a,a48148a,a48149a,a48150a,a48153a,a48156a,a48157a,a48160a,a48163a,a48164a,a48165a,a48168a,a48171a,a48172a,a48175a,a48178a,a48179a,a48180a,a48183a,a48186a,a48187a,a48190a,a48193a,a48194a,a48195a,a48198a,a48201a,a48202a,a48205a,a48208a,a48209a,a48210a,a48213a,a48216a,a48217a,a48220a,a48223a,a48224a,a48225a,a48228a,a48231a,a48232a,a48235a,a48238a,a48239a,a48240a,a48243a,a48246a,a48247a,a48250a,a48253a,a48254a,a48255a,a48258a,a48261a,a48262a,a48265a,a48268a,a48269a,a48270a,a48273a,a48276a,a48277a,a48280a,a48283a,a48284a,a48285a,a48288a,a48291a,a48292a,a48295a,a48298a,a48299a,a48300a,a48303a,a48306a,a48307a,a48310a,a48313a,a48314a,a48315a,a48318a,a48321a,a48322a,a48325a,a48328a,a48329a,a48330a,a48333a,a48336a,a48337a,a48340a,a48343a,a48344a,a48345a,a48348a,a48351a,a48352a,a48355a,a48358a,a48359a,a48360a,a48363a,a48366a,a48367a,a48370a,a48373a,a48374a,a48375a,a48378a,a48381a,a48382a,a48385a,a48388a,a48389a,a48390a,a48393a,a48396a,a48397a,a48400a,a48403a,a48404a,a48405a,a48408a,a48411a,a48412a,a48415a,a48418a,a48419a,a48420a,a48423a,a48426a,a48427a,a48430a,a48433a,a48434a,a48435a,a48438a,a48441a,a48442a,a48445a,a48448a,a48449a,a48450a,a48453a,a48456a,a48457a,a48460a,a48463a,a48464a,a48465a,a48468a,a48471a,a48472a,a48475a,a48478a,a48479a,a48480a,a48483a,a48486a,a48487a,a48490a,a48493a,a48494a,a48495a,a48498a,a48501a,a48502a,a48505a,a48508a,a48509a,a48510a,a48513a,a48516a,a48517a,a48520a,a48523a,a48524a,a48525a,a48528a,a48531a,a48532a,a48535a,a48538a,a48539a,a48540a,a48543a,a48546a,a48547a,a48550a,a48553a,a48554a,a48555a,a48558a,a48561a,a48562a,a48565a,a48568a,a48569a,a48570a,a48573a,a48576a,a48577a,a48580a,a48583a,a48584a,a48585a,a48588a,a48591a,a48592a,a48595a,a48598a,a48599a,a48600a,a48603a,a48606a,a48607a,a48610a,a48613a,a48614a,a48615a,a48618a,a48621a,a48622a,a48625a,a48628a,a48629a,a48630a,a48633a,a48636a,a48637a,a48640a,a48643a,a48644a,a48645a,a48648a,a48651a,a48652a,a48655a,a48658a,a48659a,a48660a,a48663a,a48666a,a48667a,a48670a,a48673a,a48674a,a48675a,a48678a,a48681a,a48682a,a48685a,a48688a,a48689a,a48690a,a48693a,a48696a,a48697a,a48700a,a48703a,a48704a,a48705a,a48708a,a48711a,a48712a,a48715a,a48718a,a48719a,a48720a,a48723a,a48726a,a48727a,a48730a,a48733a,a48734a,a48735a,a48738a,a48741a,a48742a,a48745a,a48748a,a48749a,a48750a,a48753a,a48756a,a48757a,a48760a,a48763a,a48764a,a48765a,a48768a,a48771a,a48772a,a48775a,a48778a,a48779a,a48780a,a48783a,a48786a,a48787a,a48790a,a48793a,a48794a,a48795a,a48798a,a48801a,a48802a,a48805a,a48808a,a48809a,a48810a,a48813a,a48816a,a48817a,a48820a,a48823a,a48824a,a48825a,a48828a,a48831a,a48832a,a48835a,a48838a,a48839a,a48840a,a48843a,a48846a,a48847a,a48850a,a48853a,a48854a,a48855a,a48858a,a48861a,a48862a,a48865a,a48868a,a48869a,a48870a,a48873a,a48876a,a48877a,a48880a,a48883a,a48884a,a48885a,a48888a,a48891a,a48892a,a48895a,a48898a,a48899a,a48900a,a48903a,a48906a,a48907a,a48910a,a48913a,a48914a,a48915a,a48918a,a48921a,a48922a,a48925a,a48928a,a48929a,a48930a,a48933a,a48936a,a48937a,a48940a,a48943a,a48944a,a48945a,a48948a,a48951a,a48952a,a48955a,a48958a,a48959a,a48960a,a48963a,a48966a,a48967a,a48970a,a48973a,a48974a,a48975a,a48978a,a48981a,a48982a,a48985a,a48988a,a48989a,a48990a,a48993a,a48996a,a48997a,a49000a,a49003a,a49004a,a49005a,a49008a,a49011a,a49012a,a49015a,a49018a,a49019a,a49020a,a49023a,a49026a,a49027a,a49030a,a49033a,a49034a,a49035a,a49038a,a49041a,a49042a,a49045a,a49048a,a49049a,a49050a,a49053a,a49056a,a49057a,a49060a,a49063a,a49064a,a49065a,a49068a,a49071a,a49072a,a49075a,a49078a,a49079a,a49080a,a49083a,a49086a,a49087a,a49090a,a49093a,a49094a,a49095a,a49098a,a49101a,a49102a,a49105a,a49108a,a49109a,a49110a,a49113a,a49116a,a49117a,a49120a,a49123a,a49124a,a49125a,a49128a,a49131a,a49132a,a49135a,a49138a,a49139a,a49140a,a49143a,a49146a,a49147a,a49150a,a49153a,a49154a,a49155a,a49158a,a49161a,a49162a,a49165a,a49168a,a49169a,a49170a,a49173a,a49176a,a49177a,a49180a,a49183a,a49184a,a49185a,a49188a,a49191a,a49192a,a49195a,a49198a,a49199a,a49200a,a49203a,a49206a,a49207a,a49210a,a49213a,a49214a,a49215a,a49218a,a49221a,a49222a,a49225a,a49228a,a49229a,a49230a,a49233a,a49236a,a49237a,a49240a,a49243a,a49244a,a49245a,a49248a,a49251a,a49252a,a49255a,a49258a,a49259a,a49260a,a49263a,a49266a,a49267a,a49270a,a49273a,a49274a,a49275a,a49278a,a49281a,a49282a,a49285a,a49288a,a49289a,a49290a,a49293a,a49296a,a49297a,a49300a,a49303a,a49304a,a49305a,a49308a,a49311a,a49312a,a49315a,a49318a,a49319a,a49320a,a49323a,a49326a,a49327a,a49330a,a49333a,a49334a,a49335a,a49338a,a49341a,a49342a,a49345a,a49348a,a49349a,a49350a,a49353a,a49356a,a49357a,a49360a,a49363a,a49364a,a49365a,a49368a,a49371a,a49372a,a49375a,a49378a,a49379a,a49380a,a49383a,a49386a,a49387a,a49390a,a49393a,a49394a,a49395a,a49398a,a49401a,a49402a,a49405a,a49408a,a49409a,a49410a,a49413a,a49416a,a49417a,a49420a,a49423a,a49424a,a49425a,a49428a,a49431a,a49432a,a49435a,a49438a,a49439a,a49440a,a49443a,a49446a,a49447a,a49450a,a49453a,a49454a,a49455a,a49458a,a49461a,a49462a,a49465a,a49468a,a49469a,a49470a,a49473a,a49476a,a49477a,a49480a,a49483a,a49484a,a49485a,a49488a,a49491a,a49492a,a49495a,a49498a,a49499a,a49500a,a49503a,a49506a,a49507a,a49510a,a49513a,a49514a,a49515a,a49518a,a49521a,a49522a,a49525a,a49528a,a49529a,a49530a,a49533a,a49536a,a49537a,a49540a,a49543a,a49544a,a49545a,a49548a,a49551a,a49552a,a49555a,a49558a,a49559a,a49560a,a49563a,a49566a,a49567a,a49570a,a49573a,a49574a,a49575a,a49578a,a49581a,a49582a,a49585a,a49588a,a49589a,a49590a,a49593a,a49596a,a49597a,a49600a,a49603a,a49604a,a49605a,a49608a,a49611a,a49612a,a49615a,a49618a,a49619a,a49620a,a49623a,a49626a,a49627a,a49630a,a49633a,a49634a,a49635a,a49638a,a49641a,a49642a,a49645a,a49648a,a49649a,a49650a,a49653a,a49656a,a49657a,a49660a,a49663a,a49664a,a49665a,a49668a,a49671a,a49672a,a49675a,a49678a,a49679a,a49680a,a49683a,a49686a,a49687a,a49690a,a49693a,a49694a,a49695a,a49698a,a49701a,a49702a,a49705a,a49708a,a49709a,a49710a,a49713a,a49716a,a49717a,a49720a,a49723a,a49724a,a49725a,a49728a,a49731a,a49732a,a49735a,a49738a,a49739a,a49740a,a49743a,a49746a,a49747a,a49750a,a49753a,a49754a,a49755a,a49758a,a49761a,a49762a,a49765a,a49768a,a49769a,a49770a,a49773a,a49776a,a49777a,a49780a,a49783a,a49784a,a49785a,a49788a,a49791a,a49792a,a49795a,a49798a,a49799a,a49800a,a49803a,a49806a,a49807a,a49810a,a49813a,a49814a,a49815a,a49818a,a49821a,a49822a,a49825a,a49828a,a49829a,a49830a,a49833a,a49836a,a49837a,a49840a,a49843a,a49844a,a49845a,a49848a,a49851a,a49852a,a49855a,a49858a,a49859a,a49860a,a49863a,a49866a,a49867a,a49870a,a49873a,a49874a,a49875a,a49878a,a49881a,a49882a,a49885a,a49888a,a49889a,a49890a,a49893a,a49896a,a49897a,a49900a,a49903a,a49904a,a49905a,a49908a,a49911a,a49912a,a49915a,a49918a,a49919a,a49920a,a49923a,a49926a,a49927a,a49930a,a49933a,a49934a,a49935a,a49938a,a49941a,a49942a,a49945a,a49948a,a49949a,a49950a,a49953a,a49956a,a49957a,a49960a,a49963a,a49964a,a49965a,a49968a,a49971a,a49972a,a49975a,a49978a,a49979a,a49980a,a49983a,a49986a,a49987a,a49990a,a49993a,a49994a,a49995a,a49998a,a50001a,a50002a,a50005a,a50008a,a50009a,a50010a,a50013a,a50016a,a50017a,a50020a,a50023a,a50024a,a50025a,a50028a,a50031a,a50032a,a50035a,a50038a,a50039a,a50040a,a50043a,a50046a,a50047a,a50050a,a50053a,a50054a,a50055a,a50058a,a50061a,a50062a,a50065a,a50068a,a50069a,a50070a,a50073a,a50076a,a50077a,a50080a,a50083a,a50084a,a50085a,a50088a,a50091a,a50092a,a50095a,a50098a,a50099a,a50100a,a50103a,a50106a,a50107a,a50110a,a50113a,a50114a,a50115a,a50118a,a50121a,a50122a,a50125a,a50128a,a50129a,a50130a,a50133a,a50136a,a50137a,a50140a,a50143a,a50144a,a50145a,a50148a,a50151a,a50152a,a50155a,a50158a,a50159a,a50160a,a50163a,a50166a,a50167a,a50170a,a50173a,a50174a,a50175a,a50178a,a50181a,a50182a,a50185a,a50188a,a50189a,a50190a,a50193a,a50196a,a50197a,a50200a,a50203a,a50204a,a50205a,a50208a,a50211a,a50212a,a50215a,a50218a,a50219a,a50220a,a50223a,a50226a,a50227a,a50230a,a50233a,a50234a,a50235a,a50238a,a50241a,a50242a,a50245a,a50248a,a50249a,a50250a,a50253a,a50256a,a50257a,a50260a,a50263a,a50264a,a50265a,a50268a,a50271a,a50272a,a50275a,a50278a,a50279a,a50280a,a50283a,a50286a,a50287a,a50290a,a50293a,a50294a,a50295a,a50298a,a50301a,a50302a,a50305a,a50308a,a50309a,a50310a,a50313a,a50316a,a50317a,a50320a,a50323a,a50324a,a50325a,a50328a,a50331a,a50332a,a50335a,a50338a,a50339a,a50340a,a50343a,a50346a,a50347a,a50350a,a50353a,a50354a,a50355a,a50358a,a50361a,a50362a,a50365a,a50368a,a50369a,a50370a,a50373a,a50376a,a50377a,a50380a,a50383a,a50384a,a50385a,a50388a,a50391a,a50392a,a50395a,a50398a,a50399a,a50400a,a50403a,a50406a,a50407a,a50410a,a50413a,a50414a,a50415a,a50418a,a50421a,a50422a,a50425a,a50428a,a50429a,a50430a,a50433a,a50436a,a50437a,a50440a,a50443a,a50444a,a50445a,a50448a,a50451a,a50452a,a50455a,a50458a,a50459a,a50460a,a50463a,a50466a,a50467a,a50470a,a50473a,a50474a,a50475a,a50478a,a50481a,a50482a,a50485a,a50488a,a50489a,a50490a,a50493a,a50496a,a50497a,a50500a,a50503a,a50504a,a50505a,a50508a,a50511a,a50512a,a50515a,a50518a,a50519a,a50520a,a50523a,a50526a,a50527a,a50530a,a50533a,a50534a,a50535a,a50538a,a50541a,a50542a,a50545a,a50548a,a50549a,a50550a,a50553a,a50556a,a50557a,a50560a,a50563a,a50564a,a50565a,a50568a,a50571a,a50572a,a50575a,a50578a,a50579a,a50580a,a50583a,a50586a,a50587a,a50590a,a50593a,a50594a,a50595a,a50598a,a50601a,a50602a,a50605a,a50608a,a50609a,a50610a,a50613a,a50616a,a50617a,a50620a,a50623a,a50624a,a50625a,a50628a,a50631a,a50632a,a50635a,a50638a,a50639a,a50640a,a50643a,a50646a,a50647a,a50650a,a50653a,a50654a,a50655a,a50658a,a50661a,a50662a,a50665a,a50668a,a50669a,a50670a,a50673a,a50676a,a50677a,a50680a,a50683a,a50684a,a50685a,a50688a,a50691a,a50692a,a50695a,a50698a,a50699a,a50700a,a50703a,a50706a,a50707a,a50710a,a50713a,a50714a,a50715a,a50718a,a50721a,a50722a,a50725a,a50728a,a50729a,a50730a,a50733a,a50736a,a50737a,a50740a,a50743a,a50744a,a50745a,a50748a,a50751a,a50752a,a50755a,a50758a,a50759a,a50760a,a50763a,a50766a,a50767a,a50770a,a50773a,a50774a,a50775a,a50778a,a50781a,a50782a,a50785a,a50788a,a50789a,a50790a,a50793a,a50796a,a50797a,a50800a,a50803a,a50804a,a50805a,a50808a,a50811a,a50812a,a50815a,a50818a,a50819a,a50820a,a50823a,a50826a,a50827a,a50830a,a50833a,a50834a,a50835a,a50838a,a50841a,a50842a,a50845a,a50848a,a50849a,a50850a,a50853a,a50856a,a50857a,a50860a,a50863a,a50864a,a50865a,a50868a,a50871a,a50872a,a50875a,a50878a,a50879a,a50880a,a50883a,a50886a,a50887a,a50890a,a50893a,a50894a,a50895a,a50898a,a50901a,a50902a,a50905a,a50908a,a50909a,a50910a,a50913a,a50916a,a50917a,a50920a,a50923a,a50924a,a50925a,a50928a,a50931a,a50932a,a50935a,a50938a,a50939a,a50940a,a50943a,a50946a,a50947a,a50950a,a50953a,a50954a,a50955a,a50958a,a50961a,a50962a,a50965a,a50968a,a50969a,a50970a,a50973a,a50976a,a50977a,a50980a,a50983a,a50984a,a50985a,a50988a,a50991a,a50992a,a50995a,a50998a,a50999a,a51000a,a51003a,a51006a,a51007a,a51010a,a51013a,a51014a,a51015a,a51018a,a51021a,a51022a,a51025a,a51028a,a51029a,a51030a,a51033a,a51036a,a51037a,a51040a,a51043a,a51044a,a51045a,a51048a,a51051a,a51052a,a51055a,a51058a,a51059a,a51060a,a51063a,a51066a,a51067a,a51070a,a51073a,a51074a,a51075a,a51078a,a51081a,a51082a,a51085a,a51088a,a51089a,a51090a,a51093a,a51096a,a51097a,a51100a,a51103a,a51104a,a51105a,a51108a,a51111a,a51112a,a51115a,a51118a,a51119a,a51120a,a51123a,a51126a,a51127a,a51130a,a51133a,a51134a,a51135a,a51138a,a51141a,a51142a,a51145a,a51148a,a51149a,a51150a,a51153a,a51156a,a51157a,a51160a,a51163a,a51164a,a51165a,a51168a,a51171a,a51172a,a51175a,a51178a,a51179a,a51180a,a51183a,a51186a,a51187a,a51190a,a51193a,a51194a,a51195a,a51198a,a51201a,a51202a,a51205a,a51208a,a51209a,a51210a,a51213a,a51216a,a51217a,a51220a,a51223a,a51224a,a51225a,a51228a,a51231a,a51232a,a51235a,a51238a,a51239a,a51240a,a51243a,a51246a,a51247a,a51250a,a51253a,a51254a,a51255a,a51258a,a51261a,a51262a,a51265a,a51268a,a51269a,a51270a,a51273a,a51276a,a51277a,a51280a,a51283a,a51284a,a51285a,a51288a,a51291a,a51292a,a51295a,a51298a,a51299a,a51300a,a51303a,a51306a,a51307a,a51310a,a51313a,a51314a,a51315a,a51318a,a51321a,a51322a,a51325a,a51328a,a51329a,a51330a,a51333a,a51336a,a51337a,a51340a,a51343a,a51344a,a51345a,a51348a,a51351a,a51352a,a51355a,a51358a,a51359a,a51360a,a51363a,a51366a,a51367a,a51370a,a51373a,a51374a,a51375a,a51378a,a51381a,a51382a,a51385a,a51388a,a51389a,a51390a,a51393a,a51396a,a51397a,a51400a,a51403a,a51404a,a51405a,a51408a,a51411a,a51412a,a51415a,a51418a,a51419a,a51420a,a51423a,a51426a,a51427a,a51430a,a51433a,a51434a,a51435a,a51438a,a51441a,a51442a,a51445a,a51448a,a51449a,a51450a,a51453a,a51456a,a51457a,a51460a,a51463a,a51464a,a51465a,a51468a,a51471a,a51472a,a51475a,a51478a,a51479a,a51480a,a51483a,a51486a,a51487a,a51490a,a51493a,a51494a,a51495a,a51498a,a51501a,a51502a,a51505a,a51508a,a51509a,a51510a,a51513a,a51516a,a51517a,a51520a,a51523a,a51524a,a51525a,a51528a,a51531a,a51532a,a51535a,a51538a,a51539a,a51540a,a51543a,a51546a,a51547a,a51550a,a51553a,a51554a,a51555a,a51558a,a51561a,a51562a,a51565a,a51568a,a51569a,a51570a,a51573a,a51576a,a51577a,a51580a,a51583a,a51584a,a51585a,a51588a,a51591a,a51592a,a51595a,a51598a,a51599a,a51600a,a51603a,a51606a,a51607a,a51610a,a51613a,a51614a,a51615a,a51618a,a51621a,a51622a,a51625a,a51628a,a51629a,a51630a,a51633a,a51636a,a51637a,a51640a,a51643a,a51644a,a51645a,a51648a,a51651a,a51652a,a51655a,a51658a,a51659a,a51660a,a51663a,a51666a,a51667a,a51670a,a51673a,a51674a,a51675a,a51678a,a51681a,a51682a,a51685a,a51688a,a51689a,a51690a,a51693a,a51696a,a51697a,a51700a,a51703a,a51704a,a51705a,a51708a,a51711a,a51712a,a51715a,a51718a,a51719a,a51720a,a51723a,a51726a,a51727a,a51730a,a51733a,a51734a,a51735a,a51738a,a51741a,a51742a,a51745a,a51748a,a51749a,a51750a,a51753a,a51756a,a51757a,a51760a,a51763a,a51764a,a51765a,a51768a,a51771a,a51772a,a51775a,a51778a,a51779a,a51780a,a51783a,a51786a,a51787a,a51790a,a51793a,a51794a,a51795a,a51798a,a51801a,a51802a,a51805a,a51808a,a51809a,a51810a,a51813a,a51816a,a51817a,a51820a,a51823a,a51824a,a51825a,a51828a,a51831a,a51832a,a51835a,a51838a,a51839a,a51840a,a51843a,a51846a,a51847a,a51850a,a51853a,a51854a,a51855a,a51858a,a51861a,a51862a,a51865a,a51868a,a51869a,a51870a,a51873a,a51876a,a51877a,a51880a,a51883a,a51884a,a51885a,a51888a,a51891a,a51892a,a51895a,a51898a,a51899a,a51900a,a51903a,a51906a,a51907a,a51910a,a51913a,a51914a,a51915a,a51918a,a51921a,a51922a,a51925a,a51928a,a51929a,a51930a,a51933a,a51936a,a51937a,a51940a,a51943a,a51944a,a51945a,a51948a,a51951a,a51952a,a51955a,a51958a,a51959a,a51960a,a51963a,a51966a,a51967a,a51970a,a51973a,a51974a,a51975a,a51978a,a51981a,a51982a,a51985a,a51988a,a51989a,a51990a,a51993a,a51996a,a51997a,a52000a,a52003a,a52004a,a52005a,a52008a,a52011a,a52012a,a52015a,a52018a,a52019a,a52020a,a52023a,a52026a,a52027a,a52030a,a52033a,a52034a,a52035a,a52038a,a52041a,a52042a,a52045a,a52048a,a52049a,a52050a,a52053a,a52056a,a52057a,a52060a,a52063a,a52064a,a52065a,a52068a,a52071a,a52072a,a52075a,a52078a,a52079a,a52080a,a52083a,a52086a,a52087a,a52090a,a52093a,a52094a,a52095a,a52098a,a52101a,a52102a,a52105a,a52108a,a52109a,a52110a,a52113a,a52116a,a52117a,a52120a,a52123a,a52124a,a52125a,a52128a,a52131a,a52132a,a52135a,a52138a,a52139a,a52140a,a52143a,a52146a,a52147a,a52150a,a52153a,a52154a,a52155a,a52158a,a52161a,a52162a,a52165a,a52168a,a52169a,a52170a,a52173a,a52176a,a52177a,a52180a,a52183a,a52184a,a52185a,a52188a,a52191a,a52192a,a52195a,a52198a,a52199a,a52200a,a52203a,a52206a,a52207a,a52210a,a52213a,a52214a,a52215a,a52218a,a52221a,a52222a,a52225a,a52228a,a52229a,a52230a,a52233a,a52236a,a52237a,a52240a,a52243a,a52244a,a52245a,a52248a,a52251a,a52252a,a52255a,a52258a,a52259a,a52260a,a52263a,a52266a,a52267a,a52270a,a52273a,a52274a,a52275a,a52278a,a52281a,a52282a,a52285a,a52288a,a52289a,a52290a,a52293a,a52296a,a52297a,a52300a,a52303a,a52304a,a52305a,a52308a,a52311a,a52312a,a52315a,a52318a,a52319a,a52320a,a52323a,a52326a,a52327a,a52330a,a52333a,a52334a,a52335a,a52338a,a52341a,a52342a,a52345a,a52348a,a52349a,a52350a,a52353a,a52356a,a52357a,a52360a,a52363a,a52364a,a52365a,a52368a,a52371a,a52372a,a52375a,a52378a,a52379a,a52380a,a52383a,a52386a,a52387a,a52390a,a52393a,a52394a,a52395a,a52398a,a52401a,a52402a,a52405a,a52408a,a52409a,a52410a,a52413a,a52416a,a52417a,a52420a,a52423a,a52424a,a52425a,a52428a,a52431a,a52432a,a52435a,a52438a,a52439a,a52440a,a52443a,a52446a,a52447a,a52450a,a52453a,a52454a,a52455a,a52458a,a52461a,a52462a,a52465a,a52468a,a52469a,a52470a,a52473a,a52476a,a52477a,a52480a,a52483a,a52484a,a52485a,a52488a,a52491a,a52492a,a52495a,a52498a,a52499a,a52500a,a52503a,a52506a,a52507a,a52510a,a52513a,a52514a,a52515a,a52518a,a52521a,a52522a,a52525a,a52528a,a52529a,a52530a,a52533a,a52536a,a52537a,a52540a,a52543a,a52544a,a52545a,a52548a,a52551a,a52552a,a52555a,a52558a,a52559a,a52560a,a52563a,a52566a,a52567a,a52570a,a52573a,a52574a,a52575a,a52578a,a52581a,a52582a,a52585a,a52588a,a52589a,a52590a,a52593a,a52596a,a52597a,a52600a,a52603a,a52604a,a52605a,a52608a,a52611a,a52612a,a52615a,a52618a,a52619a,a52620a,a52623a,a52626a,a52627a,a52630a,a52633a,a52634a,a52635a,a52638a,a52641a,a52642a,a52645a,a52648a,a52649a,a52650a,a52653a,a52656a,a52657a,a52660a,a52663a,a52664a,a52665a,a52668a,a52671a,a52672a,a52675a,a52678a,a52679a,a52680a,a52683a,a52686a,a52687a,a52690a,a52693a,a52694a,a52695a,a52698a,a52701a,a52702a,a52705a,a52708a,a52709a,a52710a,a52713a,a52716a,a52717a,a52720a,a52723a,a52724a,a52725a,a52728a,a52731a,a52732a,a52735a,a52738a,a52739a,a52740a,a52743a,a52746a,a52747a,a52750a,a52753a,a52754a,a52755a,a52758a,a52761a,a52762a,a52765a,a52768a,a52769a,a52770a,a52773a,a52776a,a52777a,a52780a,a52783a,a52784a,a52785a,a52788a,a52791a,a52792a,a52795a,a52798a,a52799a,a52800a,a52803a,a52806a,a52807a,a52810a,a52813a,a52814a,a52815a,a52818a,a52821a,a52822a,a52825a,a52828a,a52829a,a52830a,a52833a,a52836a,a52837a,a52840a,a52843a,a52844a,a52845a,a52848a,a52851a,a52852a,a52855a,a52858a,a52859a,a52860a,a52863a,a52866a,a52867a,a52870a,a52873a,a52874a,a52875a,a52878a,a52881a,a52882a,a52885a,a52888a,a52889a,a52890a,a52893a,a52896a,a52897a,a52900a,a52903a,a52904a,a52905a,a52908a,a52911a,a52912a,a52915a,a52918a,a52919a,a52920a,a52923a,a52926a,a52927a,a52930a,a52933a,a52934a,a52935a,a52938a,a52941a,a52942a,a52945a,a52948a,a52949a,a52950a,a52953a,a52956a,a52957a,a52960a,a52963a,a52964a,a52965a,a52968a,a52971a,a52972a,a52975a,a52978a,a52979a,a52980a,a52983a,a52986a,a52987a,a52990a,a52993a,a52994a,a52995a,a52998a,a53001a,a53002a,a53005a,a53008a,a53009a,a53010a,a53013a,a53016a,a53017a,a53020a,a53023a,a53024a,a53025a,a53028a,a53031a,a53032a,a53035a,a53038a,a53039a,a53040a,a53043a,a53046a,a53047a,a53050a,a53053a,a53054a,a53055a,a53058a,a53061a,a53062a,a53065a,a53068a,a53069a,a53070a,a53073a,a53076a,a53077a,a53080a,a53083a,a53084a,a53085a,a53088a,a53091a,a53092a,a53095a,a53098a,a53099a,a53100a,a53103a,a53106a,a53107a,a53110a,a53113a,a53114a,a53115a,a53118a,a53121a,a53122a,a53125a,a53128a,a53129a,a53130a,a53133a,a53136a,a53137a,a53140a,a53143a,a53144a,a53145a,a53148a,a53151a,a53152a,a53155a,a53158a,a53159a,a53160a,a53163a,a53166a,a53167a,a53170a,a53173a,a53174a,a53175a,a53178a,a53181a,a53182a,a53185a,a53188a,a53189a,a53190a,a53193a,a53196a,a53197a,a53200a,a53203a,a53204a,a53205a,a53208a,a53211a,a53212a,a53215a,a53218a,a53219a,a53220a,a53223a,a53226a,a53227a,a53230a,a53233a,a53234a,a53235a,a53238a,a53241a,a53242a,a53245a,a53248a,a53249a,a53250a,a53253a,a53256a,a53257a,a53260a,a53263a,a53264a,a53265a,a53268a,a53271a,a53272a,a53275a,a53278a,a53279a,a53280a,a53283a,a53286a,a53287a,a53290a,a53293a,a53294a,a53295a,a53298a,a53301a,a53302a,a53305a,a53308a,a53309a,a53310a,a53313a,a53316a,a53317a,a53320a,a53323a,a53324a,a53325a,a53328a,a53331a,a53332a,a53335a,a53338a,a53339a,a53340a,a53343a,a53346a,a53347a,a53350a,a53353a,a53354a,a53355a,a53358a,a53361a,a53362a,a53365a,a53368a,a53369a,a53370a,a53373a,a53376a,a53377a,a53380a,a53383a,a53384a,a53385a,a53388a,a53391a,a53392a,a53395a,a53398a,a53399a,a53400a,a53403a,a53406a,a53407a,a53410a,a53413a,a53414a,a53415a,a53418a,a53421a,a53422a,a53425a,a53428a,a53429a,a53430a,a53433a,a53436a,a53437a,a53440a,a53443a,a53444a,a53445a,a53448a,a53451a,a53452a,a53455a,a53458a,a53459a,a53460a,a53463a,a53466a,a53467a,a53470a,a53473a,a53474a,a53475a,a53478a,a53481a,a53482a,a53485a,a53488a,a53489a,a53490a,a53493a,a53496a,a53497a,a53500a,a53503a,a53504a,a53505a,a53508a,a53511a,a53512a,a53515a,a53518a,a53519a,a53520a,a53523a,a53526a,a53527a,a53530a,a53533a,a53534a,a53535a,a53538a,a53541a,a53542a,a53545a,a53548a,a53549a,a53550a,a53553a,a53556a,a53557a,a53560a,a53563a,a53564a,a53565a,a53568a,a53571a,a53572a,a53575a,a53578a,a53579a,a53580a,a53583a,a53586a,a53587a,a53590a,a53593a,a53594a,a53595a,a53598a,a53601a,a53602a,a53605a,a53608a,a53609a,a53610a,a53613a,a53616a,a53617a,a53620a,a53623a,a53624a,a53625a,a53628a,a53631a,a53632a,a53635a,a53638a,a53639a,a53640a,a53643a,a53646a,a53647a,a53650a,a53653a,a53654a,a53655a,a53658a,a53661a,a53662a,a53665a,a53668a,a53669a,a53670a,a53673a,a53676a,a53677a,a53680a,a53683a,a53684a,a53685a,a53688a,a53691a,a53692a,a53695a,a53698a,a53699a,a53700a,a53703a,a53706a,a53707a,a53710a,a53713a,a53714a,a53715a,a53718a,a53721a,a53722a,a53725a,a53728a,a53729a,a53730a,a53733a,a53736a,a53737a,a53740a,a53743a,a53744a,a53745a,a53748a,a53751a,a53752a,a53755a,a53758a,a53759a,a53760a,a53763a,a53766a,a53767a,a53770a,a53773a,a53774a,a53775a,a53778a,a53781a,a53782a,a53785a,a53788a,a53789a,a53790a,a53793a,a53796a,a53797a,a53800a,a53803a,a53804a,a53805a,a53808a,a53811a,a53812a,a53815a,a53818a,a53819a,a53820a,a53823a,a53826a,a53827a,a53830a,a53833a,a53834a,a53835a,a53838a,a53841a,a53842a,a53845a,a53848a,a53849a,a53850a,a53853a,a53856a,a53857a,a53860a,a53863a,a53864a,a53865a,a53868a,a53871a,a53872a,a53875a,a53878a,a53879a,a53880a,a53883a,a53886a,a53887a,a53890a,a53893a,a53894a,a53895a,a53898a,a53901a,a53902a,a53905a,a53908a,a53909a,a53910a,a53913a,a53916a,a53917a,a53920a,a53923a,a53924a,a53925a,a53928a,a53931a,a53932a,a53935a,a53938a,a53939a,a53940a,a53943a,a53946a,a53947a,a53950a,a53953a,a53954a,a53955a,a53958a,a53961a,a53962a,a53965a,a53968a,a53969a,a53970a,a53973a,a53976a,a53977a,a53980a,a53983a,a53984a,a53985a,a53988a,a53991a,a53992a,a53995a,a53998a,a53999a,a54000a,a54003a,a54006a,a54007a,a54010a,a54013a,a54014a,a54015a,a54018a,a54021a,a54022a,a54025a,a54028a,a54029a,a54030a,a54033a,a54036a,a54037a,a54040a,a54043a,a54044a,a54045a,a54048a,a54051a,a54052a,a54055a,a54058a,a54059a,a54060a,a54063a,a54066a,a54067a,a54070a,a54073a,a54074a,a54075a,a54078a,a54081a,a54082a,a54085a,a54088a,a54089a,a54090a,a54093a,a54096a,a54097a,a54100a,a54103a,a54104a,a54105a,a54108a,a54111a,a54112a,a54115a,a54118a,a54119a,a54120a,a54123a,a54126a,a54127a,a54130a,a54133a,a54134a,a54135a,a54138a,a54141a,a54142a,a54145a,a54148a,a54149a,a54150a,a54153a,a54156a,a54157a,a54160a,a54163a,a54164a,a54165a,a54168a,a54171a,a54172a,a54175a,a54178a,a54179a,a54180a,a54183a,a54186a,a54187a,a54190a,a54193a,a54194a,a54195a,a54198a,a54201a,a54202a,a54205a,a54208a,a54209a,a54210a,a54213a,a54216a,a54217a,a54220a,a54223a,a54224a,a54225a,a54228a,a54231a,a54232a,a54235a,a54238a,a54239a,a54240a,a54243a,a54246a,a54247a,a54250a,a54253a,a54254a,a54255a,a54258a,a54261a,a54262a,a54265a,a54268a,a54269a,a54270a,a54273a,a54276a,a54277a,a54280a,a54283a,a54284a,a54285a,a54288a,a54291a,a54292a,a54295a,a54298a,a54299a,a54300a,a54303a,a54306a,a54307a,a54310a,a54313a,a54314a,a54315a,a54318a,a54321a,a54322a,a54325a,a54328a,a54329a,a54330a,a54333a,a54336a,a54337a,a54340a,a54343a,a54344a,a54345a,a54348a,a54351a,a54352a,a54355a,a54358a,a54359a,a54360a,a54363a,a54366a,a54367a,a54370a,a54373a,a54374a,a54375a,a54378a,a54381a,a54382a,a54385a,a54388a,a54389a,a54390a,a54393a,a54396a,a54397a,a54400a,a54403a,a54404a,a54405a,a54408a,a54411a,a54412a,a54415a,a54418a,a54419a,a54420a,a54423a,a54426a,a54427a,a54430a,a54433a,a54434a,a54435a,a54438a,a54441a,a54442a,a54445a,a54448a,a54449a,a54450a,a54453a,a54456a,a54457a,a54460a,a54463a,a54464a,a54465a,a54468a,a54471a,a54472a,a54475a,a54478a,a54479a,a54480a,a54483a,a54486a,a54487a,a54490a,a54493a,a54494a,a54495a,a54498a,a54501a,a54502a,a54505a,a54508a,a54509a,a54510a,a54513a,a54516a,a54517a,a54520a,a54523a,a54524a,a54525a,a54528a,a54531a,a54532a,a54535a,a54538a,a54539a,a54540a,a54543a,a54546a,a54547a,a54550a,a54553a,a54554a,a54555a,a54558a,a54561a,a54562a,a54565a,a54568a,a54569a,a54570a,a54573a,a54576a,a54577a,a54580a,a54583a,a54584a,a54585a,a54588a,a54591a,a54592a,a54595a,a54598a,a54599a,a54600a,a54603a,a54606a,a54607a,a54610a,a54613a,a54614a,a54615a,a54618a,a54621a,a54622a,a54625a,a54628a,a54629a,a54630a,a54633a,a54636a,a54637a,a54640a,a54643a,a54644a,a54645a,a54648a,a54651a,a54652a,a54655a,a54658a,a54659a,a54660a,a54663a,a54666a,a54667a,a54670a,a54673a,a54674a,a54675a,a54678a,a54681a,a54682a,a54685a,a54688a,a54689a,a54690a,a54693a,a54696a,a54697a,a54700a,a54703a,a54704a,a54705a,a54708a,a54711a,a54712a,a54715a,a54718a,a54719a,a54720a,a54723a,a54726a,a54727a,a54730a,a54733a,a54734a,a54735a,a54738a,a54741a,a54742a,a54745a,a54748a,a54749a,a54750a,a54753a,a54756a,a54757a,a54760a,a54763a,a54764a,a54765a,a54768a,a54771a,a54772a,a54775a,a54778a,a54779a,a54780a,a54783a,a54786a,a54787a,a54790a,a54793a,a54794a,a54795a,a54798a,a54801a,a54802a,a54805a,a54808a,a54809a,a54810a,a54813a,a54816a,a54817a,a54820a,a54823a,a54824a,a54825a,a54828a,a54831a,a54832a,a54835a,a54838a,a54839a,a54840a,a54843a,a54846a,a54847a,a54850a,a54853a,a54854a,a54855a,a54858a,a54861a,a54862a,a54865a,a54868a,a54869a,a54870a,a54873a,a54876a,a54877a,a54880a,a54883a,a54884a,a54885a,a54888a,a54891a,a54892a,a54895a,a54898a,a54899a,a54900a,a54903a,a54906a,a54907a,a54910a,a54913a,a54914a,a54915a,a54918a,a54921a,a54922a,a54925a,a54928a,a54929a,a54930a,a54933a,a54936a,a54937a,a54940a,a54943a,a54944a,a54945a,a54948a,a54951a,a54952a,a54955a,a54958a,a54959a,a54960a,a54963a,a54966a,a54967a,a54970a,a54973a,a54974a,a54975a,a54978a,a54981a,a54982a,a54985a,a54988a,a54989a,a54990a,a54993a,a54996a,a54997a,a55000a,a55003a,a55004a,a55005a,a55008a,a55011a,a55012a,a55015a,a55018a,a55019a,a55020a,a55023a,a55026a,a55027a,a55030a,a55033a,a55034a,a55035a,a55038a,a55041a,a55042a,a55045a,a55048a,a55049a,a55050a,a55053a,a55056a,a55057a,a55060a,a55063a,a55064a,a55065a,a55068a,a55071a,a55072a,a55075a,a55078a,a55079a,a55080a,a55083a,a55086a,a55087a,a55090a,a55093a,a55094a,a55095a,a55098a,a55101a,a55102a,a55105a,a55108a,a55109a,a55110a,a55113a,a55116a,a55117a,a55120a,a55123a,a55124a,a55125a,a55128a,a55131a,a55132a,a55135a,a55138a,a55139a,a55140a,a55143a,a55146a,a55147a,a55150a,a55153a,a55154a,a55155a,a55158a,a55161a,a55162a,a55165a,a55168a,a55169a,a55170a,a55173a,a55176a,a55177a,a55180a,a55183a,a55184a,a55185a,a55188a,a55191a,a55192a,a55195a,a55198a,a55199a,a55200a,a55203a,a55206a,a55207a,a55210a,a55213a,a55214a,a55215a,a55218a,a55221a,a55222a,a55225a,a55228a,a55229a,a55230a,a55233a,a55236a,a55237a,a55240a,a55243a,a55244a,a55245a,a55248a,a55251a,a55252a,a55255a,a55258a,a55259a,a55260a,a55263a,a55266a,a55267a,a55270a,a55273a,a55274a,a55275a,a55278a,a55281a,a55282a,a55285a,a55288a,a55289a,a55290a,a55293a,a55296a,a55297a,a55300a,a55303a,a55304a,a55305a,a55308a,a55311a,a55312a,a55315a,a55318a,a55319a,a55320a,a55323a,a55326a,a55327a,a55330a,a55333a,a55334a,a55335a,a55338a,a55341a,a55342a,a55345a,a55348a,a55349a,a55350a,a55353a,a55356a,a55357a,a55360a,a55363a,a55364a,a55365a,a55368a,a55371a,a55372a,a55375a,a55378a,a55379a,a55380a,a55383a,a55386a,a55387a,a55390a,a55393a,a55394a,a55395a,a55398a,a55401a,a55402a,a55405a,a55408a,a55409a,a55410a,a55413a,a55416a,a55417a,a55420a,a55423a,a55424a,a55425a,a55428a,a55431a,a55432a,a55435a,a55438a,a55439a,a55440a,a55443a,a55446a,a55447a,a55450a,a55453a,a55454a,a55455a,a55458a,a55461a,a55462a,a55465a,a55468a,a55469a,a55470a,a55473a,a55476a,a55477a,a55480a,a55483a,a55484a,a55485a,a55488a,a55491a,a55492a,a55495a,a55498a,a55499a,a55500a,a55503a,a55506a,a55507a,a55510a,a55513a,a55514a,a55515a,a55518a,a55521a,a55522a,a55525a,a55528a,a55529a,a55530a,a55533a,a55536a,a55537a,a55540a,a55543a,a55544a,a55545a,a55548a,a55551a,a55552a,a55555a,a55558a,a55559a,a55560a,a55563a,a55566a,a55567a,a55570a,a55573a,a55574a,a55575a,a55578a,a55581a,a55582a,a55585a,a55588a,a55589a,a55590a,a55593a,a55596a,a55597a,a55600a,a55603a,a55604a,a55605a,a55608a,a55611a,a55612a,a55615a,a55618a,a55619a,a55620a,a55623a,a55626a,a55627a,a55630a,a55633a,a55634a,a55635a,a55638a,a55641a,a55642a,a55645a,a55648a,a55649a,a55650a,a55653a,a55656a,a55657a,a55660a,a55663a,a55664a,a55665a,a55668a,a55671a,a55672a,a55675a,a55678a,a55679a,a55680a,a55683a,a55686a,a55687a,a55690a,a55693a,a55694a,a55695a,a55698a,a55701a,a55702a,a55705a,a55708a,a55709a,a55710a,a55713a,a55716a,a55717a,a55720a,a55723a,a55724a,a55725a,a55728a,a55731a,a55732a,a55735a,a55738a,a55739a,a55740a,a55743a,a55746a,a55747a,a55750a,a55753a,a55754a,a55755a,a55758a,a55761a,a55762a,a55765a,a55768a,a55769a,a55770a,a55773a,a55776a,a55777a,a55780a,a55783a,a55784a,a55785a,a55788a,a55791a,a55792a,a55795a,a55798a,a55799a,a55800a,a55803a,a55806a,a55807a,a55810a,a55813a,a55814a,a55815a,a55818a,a55821a,a55822a,a55825a,a55828a,a55829a,a55830a,a55833a,a55836a,a55837a,a55840a,a55843a,a55844a,a55845a,a55848a,a55851a,a55852a,a55855a,a55858a,a55859a,a55860a,a55863a,a55866a,a55867a,a55870a,a55873a,a55874a,a55875a,a55878a,a55881a,a55882a,a55885a,a55888a,a55889a,a55890a,a55893a,a55896a,a55897a,a55900a,a55903a,a55904a,a55905a,a55908a,a55911a,a55912a,a55915a,a55918a,a55919a,a55920a,a55923a,a55926a,a55927a,a55930a,a55933a,a55934a,a55935a,a55938a,a55941a,a55942a,a55945a,a55948a,a55949a,a55950a,a55953a,a55956a,a55957a,a55960a,a55963a,a55964a,a55965a,a55968a,a55971a,a55972a,a55975a,a55978a,a55979a,a55980a,a55983a,a55986a,a55987a,a55990a,a55993a,a55994a,a55995a,a55998a,a56001a,a56002a,a56005a,a56008a,a56009a,a56010a,a56013a,a56016a,a56017a,a56020a,a56023a,a56024a,a56025a,a56028a,a56031a,a56032a,a56035a,a56038a,a56039a,a56040a,a56043a,a56046a,a56047a,a56050a,a56053a,a56054a,a56055a,a56058a,a56061a,a56062a,a56065a,a56068a,a56069a,a56070a,a56073a,a56076a,a56077a,a56080a,a56083a,a56084a,a56085a,a56088a,a56091a,a56092a,a56095a,a56098a,a56099a,a56100a,a56103a,a56106a,a56107a,a56110a,a56113a,a56114a,a56115a,a56118a,a56121a,a56122a,a56125a,a56128a,a56129a,a56130a,a56133a,a56136a,a56137a,a56140a,a56143a,a56144a,a56145a,a56148a,a56151a,a56152a,a56155a,a56158a,a56159a,a56160a,a56163a,a56166a,a56167a,a56170a,a56173a,a56174a,a56175a,a56178a,a56181a,a56182a,a56185a,a56188a,a56189a,a56190a,a56193a,a56196a,a56197a,a56200a,a56203a,a56204a,a56205a,a56208a,a56211a,a56212a,a56215a,a56218a,a56219a,a56220a,a56223a,a56226a,a56227a,a56230a,a56233a,a56234a,a56235a,a56238a,a56241a,a56242a,a56245a,a56248a,a56249a,a56250a,a56253a,a56256a,a56257a,a56260a,a56263a,a56264a,a56265a,a56268a,a56271a,a56272a,a56275a,a56278a,a56279a,a56280a,a56283a,a56286a,a56287a,a56290a,a56293a,a56294a,a56295a,a56298a,a56301a,a56302a,a56305a,a56308a,a56309a,a56310a,a56313a,a56316a,a56317a,a56320a,a56323a,a56324a,a56325a,a56328a,a56331a,a56332a,a56335a,a56338a,a56339a,a56340a,a56343a,a56346a,a56347a,a56350a,a56353a,a56354a,a56355a,a56358a,a56361a,a56362a,a56365a,a56368a,a56369a,a56370a,a56373a,a56376a,a56377a,a56380a,a56383a,a56384a,a56385a,a56388a,a56391a,a56392a,a56395a,a56398a,a56399a,a56400a,a56403a,a56406a,a56407a,a56410a,a56413a,a56414a,a56415a,a56418a,a56421a,a56422a,a56425a,a56428a,a56429a,a56430a,a56433a,a56436a,a56437a,a56440a,a56443a,a56444a,a56445a,a56448a,a56451a,a56452a,a56455a,a56458a,a56459a,a56460a,a56463a,a56466a,a56467a,a56470a,a56473a,a56474a,a56475a,a56478a,a56481a,a56482a,a56485a,a56488a,a56489a,a56490a,a56493a,a56496a,a56497a,a56500a,a56503a,a56504a,a56505a,a56508a,a56511a,a56512a,a56515a,a56518a,a56519a,a56520a,a56523a,a56526a,a56527a,a56530a,a56533a,a56534a,a56535a,a56538a,a56541a,a56542a,a56545a,a56548a,a56549a,a56550a,a56553a,a56556a,a56557a,a56560a,a56563a,a56564a,a56565a,a56568a,a56571a,a56572a,a56575a,a56578a,a56579a,a56580a,a56583a,a56586a,a56587a,a56590a,a56593a,a56594a,a56595a,a56598a,a56601a,a56602a,a56605a,a56608a,a56609a,a56610a,a56613a,a56616a,a56617a,a56620a,a56623a,a56624a,a56625a,a56628a,a56631a,a56632a,a56635a,a56638a,a56639a,a56640a,a56643a,a56646a,a56647a,a56650a,a56653a,a56654a,a56655a,a56658a,a56661a,a56662a,a56665a,a56668a,a56669a,a56670a,a56673a,a56676a,a56677a,a56680a,a56683a,a56684a,a56685a,a56688a,a56691a,a56692a,a56695a,a56698a,a56699a,a56700a,a56703a,a56706a,a56707a,a56710a,a56713a,a56714a,a56715a,a56718a,a56721a,a56722a,a56725a,a56728a,a56729a,a56730a,a56733a,a56736a,a56737a,a56740a,a56743a,a56744a,a56745a,a56748a,a56751a,a56752a,a56755a,a56758a,a56759a,a56760a,a56763a,a56766a,a56767a,a56770a,a56773a,a56774a,a56775a,a56778a,a56781a,a56782a,a56785a,a56788a,a56789a,a56790a,a56793a,a56796a,a56797a,a56800a,a56803a,a56804a,a56805a,a56808a,a56811a,a56812a,a56815a,a56818a,a56819a,a56820a,a56823a,a56826a,a56827a,a56830a,a56833a,a56834a,a56835a,a56838a,a56841a,a56842a,a56845a,a56848a,a56849a,a56850a,a56853a,a56856a,a56857a,a56860a,a56863a,a56864a,a56865a,a56868a,a56871a,a56872a,a56875a,a56878a,a56879a,a56880a,a56883a,a56886a,a56887a,a56890a,a56893a,a56894a,a56895a,a56898a,a56901a,a56902a,a56905a,a56908a,a56909a,a56910a,a56913a,a56916a,a56917a,a56920a,a56923a,a56924a,a56925a,a56928a,a56931a,a56932a,a56935a,a56938a,a56939a,a56940a,a56943a,a56946a,a56947a,a56950a,a56953a,a56954a,a56955a,a56958a,a56961a,a56962a,a56965a,a56968a,a56969a,a56970a,a56973a,a56976a,a56977a,a56980a,a56983a,a56984a,a56985a,a56988a,a56991a,a56992a,a56995a,a56998a,a56999a,a57000a,a57003a,a57006a,a57007a,a57010a,a57013a,a57014a,a57015a,a57018a,a57021a,a57022a,a57025a,a57028a,a57029a,a57030a,a57033a,a57036a,a57037a,a57040a,a57043a,a57044a,a57045a,a57048a,a57051a,a57052a,a57055a,a57058a,a57059a,a57060a,a57063a,a57066a,a57067a,a57070a,a57073a,a57074a,a57075a,a57078a,a57081a,a57082a,a57085a,a57088a,a57089a,a57090a,a57093a,a57096a,a57097a,a57100a,a57103a,a57104a,a57105a,a57108a,a57111a,a57112a,a57115a,a57118a,a57119a,a57120a,a57123a,a57126a,a57127a,a57130a,a57133a,a57134a,a57135a,a57138a,a57141a,a57142a,a57145a,a57148a,a57149a,a57150a,a57153a,a57156a,a57157a,a57160a,a57163a,a57164a,a57165a,a57168a,a57171a,a57172a,a57175a,a57178a,a57179a,a57180a,a57183a,a57186a,a57187a,a57190a,a57193a,a57194a,a57195a,a57198a,a57201a,a57202a,a57205a,a57208a,a57209a,a57210a,a57213a,a57216a,a57217a,a57220a,a57223a,a57224a,a57225a,a57228a,a57231a,a57232a,a57235a,a57238a,a57239a,a57240a,a57243a,a57246a,a57247a,a57250a,a57253a,a57254a,a57255a,a57258a,a57261a,a57262a,a57265a,a57268a,a57269a,a57270a,a57273a,a57276a,a57277a,a57280a,a57283a,a57284a,a57285a,a57288a,a57291a,a57292a,a57295a,a57298a,a57299a,a57300a,a57303a,a57306a,a57307a,a57310a,a57313a,a57314a,a57315a,a57318a,a57321a,a57322a,a57325a,a57328a,a57329a,a57330a,a57333a,a57336a,a57337a,a57340a,a57343a,a57344a,a57345a,a57348a,a57351a,a57352a,a57355a,a57358a,a57359a,a57360a,a57363a,a57366a,a57367a,a57370a,a57373a,a57374a,a57375a,a57378a,a57381a,a57382a,a57385a,a57388a,a57389a,a57390a,a57393a,a57396a,a57397a,a57400a,a57403a,a57404a,a57405a,a57408a,a57411a,a57412a,a57415a,a57418a,a57419a,a57420a,a57423a,a57426a,a57427a,a57430a,a57433a,a57434a,a57435a,a57438a,a57441a,a57442a,a57445a,a57448a,a57449a,a57450a,a57453a,a57456a,a57457a,a57460a,a57463a,a57464a,a57465a,a57468a,a57471a,a57472a,a57475a,a57478a,a57479a,a57480a,a57483a,a57486a,a57487a,a57490a,a57493a,a57494a,a57495a,a57498a,a57501a,a57502a,a57505a,a57508a,a57509a,a57510a,a57513a,a57516a,a57517a,a57520a,a57523a,a57524a,a57525a,a57528a,a57531a,a57532a,a57535a,a57538a,a57539a,a57540a,a57543a,a57546a,a57547a,a57550a,a57553a,a57554a,a57555a,a57558a,a57561a,a57562a,a57565a,a57568a,a57569a,a57570a,a57573a,a57576a,a57577a,a57580a,a57583a,a57584a,a57585a,a57588a,a57591a,a57592a,a57595a,a57598a,a57599a,a57600a,a57603a,a57606a,a57607a,a57610a,a57613a,a57614a,a57615a,a57618a,a57621a,a57622a,a57625a,a57628a,a57629a,a57630a,a57633a,a57636a,a57637a,a57640a,a57643a,a57644a,a57645a,a57648a,a57651a,a57652a,a57655a,a57658a,a57659a,a57660a,a57663a,a57666a,a57667a,a57670a,a57673a,a57674a,a57675a,a57678a,a57681a,a57682a,a57685a,a57688a,a57689a,a57690a,a57693a,a57696a,a57697a,a57700a,a57703a,a57704a,a57705a,a57708a,a57711a,a57712a,a57715a,a57718a,a57719a,a57720a,a57723a,a57726a,a57727a,a57730a,a57733a,a57734a,a57735a,a57738a,a57741a,a57742a,a57745a,a57748a,a57749a,a57750a,a57753a,a57756a,a57757a,a57760a,a57763a,a57764a,a57765a,a57768a,a57771a,a57772a,a57775a,a57778a,a57779a,a57780a,a57783a,a57786a,a57787a,a57790a,a57793a,a57794a,a57795a,a57798a,a57801a,a57802a,a57805a,a57808a,a57809a,a57810a,a57813a,a57816a,a57817a,a57820a,a57823a,a57824a,a57825a,a57828a,a57831a,a57832a,a57835a,a57838a,a57839a,a57840a,a57843a,a57846a,a57847a,a57850a,a57853a,a57854a,a57855a,a57858a,a57861a,a57862a,a57865a,a57868a,a57869a,a57870a,a57873a,a57876a,a57877a,a57880a,a57883a,a57884a,a57885a,a57888a,a57891a,a57892a,a57895a,a57898a,a57899a,a57900a,a57903a,a57906a,a57907a,a57910a,a57913a,a57914a,a57915a,a57918a,a57921a,a57922a,a57925a,a57928a,a57929a,a57930a,a57933a,a57936a,a57937a,a57940a,a57943a,a57944a,a57945a,a57948a,a57951a,a57952a,a57955a,a57958a,a57959a,a57960a,a57963a,a57966a,a57967a,a57970a,a57973a,a57974a,a57975a,a57978a,a57981a,a57982a,a57985a,a57988a,a57989a,a57990a,a57993a,a57996a,a57997a,a58000a,a58003a,a58004a,a58005a,a58008a,a58011a,a58012a,a58015a,a58018a,a58019a,a58020a,a58023a,a58026a,a58027a,a58030a,a58033a,a58034a,a58035a,a58038a,a58041a,a58042a,a58045a,a58048a,a58049a,a58050a,a58053a,a58056a,a58057a,a58060a,a58063a,a58064a,a58065a,a58068a,a58071a,a58072a,a58075a,a58078a,a58079a,a58080a,a58083a,a58086a,a58087a,a58090a,a58093a,a58094a,a58095a,a58098a,a58101a,a58102a,a58105a,a58108a,a58109a,a58110a,a58113a,a58116a,a58117a,a58120a,a58123a,a58124a,a58125a,a58128a,a58131a,a58132a,a58135a,a58138a,a58139a,a58140a,a58143a,a58146a,a58147a,a58150a,a58153a,a58154a,a58155a,a58158a,a58161a,a58162a,a58165a,a58168a,a58169a,a58170a,a58173a,a58176a,a58177a,a58180a,a58183a,a58184a,a58185a,a58188a,a58191a,a58192a,a58195a,a58198a,a58199a,a58200a,a58203a,a58206a,a58207a,a58210a,a58213a,a58214a,a58215a,a58218a,a58221a,a58222a,a58225a,a58228a,a58229a,a58230a,a58233a,a58236a,a58237a,a58240a,a58243a,a58244a,a58245a,a58248a,a58251a,a58252a,a58255a,a58258a,a58259a,a58260a,a58263a,a58266a,a58267a,a58270a,a58273a,a58274a,a58275a,a58278a,a58281a,a58282a,a58285a,a58288a,a58289a,a58290a,a58293a,a58296a,a58297a,a58300a,a58303a,a58304a,a58305a,a58308a,a58311a,a58312a,a58315a,a58318a,a58319a,a58320a,a58323a,a58326a,a58327a,a58330a,a58333a,a58334a,a58335a,a58338a,a58341a,a58342a,a58345a,a58348a,a58349a,a58350a,a58353a,a58356a,a58357a,a58360a,a58363a,a58364a,a58365a,a58368a,a58371a,a58372a,a58375a,a58378a,a58379a,a58380a,a58383a,a58386a,a58387a,a58390a,a58393a,a58394a,a58395a,a58398a,a58401a,a58402a,a58405a,a58408a,a58409a,a58410a,a58413a,a58416a,a58417a,a58420a,a58423a,a58424a,a58425a,a58428a,a58431a,a58432a,a58435a,a58438a,a58439a,a58440a,a58443a,a58446a,a58447a,a58450a,a58453a,a58454a,a58455a,a58458a,a58461a,a58462a,a58465a,a58468a,a58469a,a58470a,a58473a,a58476a,a58477a,a58480a,a58483a,a58484a,a58485a,a58488a,a58491a,a58492a,a58495a,a58498a,a58499a,a58500a,a58503a,a58506a,a58507a,a58510a,a58513a,a58514a,a58515a,a58518a,a58521a,a58522a,a58525a,a58528a,a58529a,a58530a,a58533a,a58536a,a58537a,a58540a,a58543a,a58544a,a58545a,a58548a,a58551a,a58552a,a58555a,a58558a,a58559a,a58560a,a58563a,a58566a,a58567a,a58570a,a58573a,a58574a,a58575a,a58578a,a58581a,a58582a,a58585a,a58588a,a58589a,a58590a,a58593a,a58596a,a58597a,a58600a,a58603a,a58604a,a58605a,a58608a,a58611a,a58612a,a58615a,a58618a,a58619a,a58620a,a58623a,a58626a,a58627a,a58630a,a58633a,a58634a,a58635a,a58638a,a58641a,a58642a,a58645a,a58648a,a58649a,a58650a,a58653a,a58656a,a58657a,a58660a,a58663a,a58664a,a58665a,a58668a,a58671a,a58672a,a58675a,a58678a,a58679a,a58680a,a58683a,a58686a,a58687a,a58690a,a58693a,a58694a,a58695a,a58698a,a58701a,a58702a,a58705a,a58708a,a58709a,a58710a,a58713a,a58716a,a58717a,a58720a,a58723a,a58724a,a58725a,a58728a,a58731a,a58732a,a58735a,a58738a,a58739a,a58740a,a58743a,a58746a,a58747a,a58750a,a58753a,a58754a,a58755a,a58758a,a58761a,a58762a,a58765a,a58768a,a58769a,a58770a,a58773a,a58776a,a58777a,a58780a,a58783a,a58784a,a58785a,a58788a,a58791a,a58792a,a58795a,a58798a,a58799a,a58800a,a58803a,a58806a,a58807a,a58810a,a58813a,a58814a,a58815a,a58818a,a58821a,a58822a,a58825a,a58828a,a58829a,a58830a,a58833a,a58836a,a58837a,a58840a,a58843a,a58844a,a58845a,a58848a,a58851a,a58852a,a58855a,a58858a,a58859a,a58860a,a58863a,a58866a,a58867a,a58870a,a58873a,a58874a,a58875a,a58878a,a58881a,a58882a,a58885a,a58888a,a58889a,a58890a,a58893a,a58896a,a58897a,a58900a,a58903a,a58904a,a58905a,a58908a,a58911a,a58912a,a58915a,a58918a,a58919a,a58920a,a58923a,a58926a,a58927a,a58930a,a58933a,a58934a,a58935a,a58938a,a58941a,a58942a,a58945a,a58948a,a58949a,a58950a,a58953a,a58956a,a58957a,a58960a,a58963a,a58964a,a58965a,a58968a,a58971a,a58972a,a58975a,a58978a,a58979a,a58980a,a58983a,a58986a,a58987a,a58990a,a58993a,a58994a,a58995a,a58998a,a59001a,a59002a,a59005a,a59008a,a59009a,a59010a,a59013a,a59016a,a59017a,a59020a,a59023a,a59024a,a59025a,a59028a,a59031a,a59032a,a59035a,a59038a,a59039a,a59040a,a59043a,a59046a,a59047a,a59050a,a59053a,a59054a,a59055a,a59058a,a59061a,a59062a,a59065a,a59068a,a59069a,a59070a,a59073a,a59076a,a59077a,a59080a,a59083a,a59084a,a59085a,a59088a,a59091a,a59092a,a59095a,a59098a,a59099a,a59100a,a59103a,a59106a,a59107a,a59110a,a59113a,a59114a,a59115a,a59118a,a59121a,a59122a,a59125a,a59128a,a59129a,a59130a,a59133a,a59136a,a59137a,a59140a,a59143a,a59144a,a59145a,a59148a,a59151a,a59152a,a59155a,a59158a,a59159a,a59160a,a59163a,a59166a,a59167a,a59170a,a59173a,a59174a,a59175a,a59178a,a59181a,a59182a,a59185a,a59188a,a59189a,a59190a,a59193a,a59196a,a59197a,a59200a,a59203a,a59204a,a59205a,a59208a,a59211a,a59212a,a59215a,a59218a,a59219a,a59220a,a59223a,a59226a,a59227a,a59230a,a59233a,a59234a,a59235a,a59238a,a59241a,a59242a,a59245a,a59248a,a59249a,a59250a,a59253a,a59256a,a59257a,a59260a,a59263a,a59264a,a59265a,a59268a,a59271a,a59272a,a59275a,a59278a,a59279a,a59280a,a59283a,a59286a,a59287a,a59290a,a59293a,a59294a,a59295a,a59298a,a59301a,a59302a,a59305a,a59308a,a59309a,a59310a,a59313a,a59316a,a59317a,a59320a,a59323a,a59324a,a59325a,a59328a,a59331a,a59332a,a59335a,a59338a,a59339a,a59340a,a59343a,a59346a,a59347a,a59350a,a59353a,a59354a,a59355a,a59358a,a59361a,a59362a,a59365a,a59368a,a59369a,a59370a,a59373a,a59376a,a59377a,a59380a,a59383a,a59384a,a59385a,a59388a,a59391a,a59392a,a59395a,a59398a,a59399a,a59400a,a59403a,a59406a,a59407a,a59410a,a59413a,a59414a,a59415a,a59418a,a59421a,a59422a,a59425a,a59428a,a59429a,a59430a,a59433a,a59436a,a59437a,a59440a,a59443a,a59444a,a59445a,a59448a,a59451a,a59452a,a59455a,a59458a,a59459a,a59460a,a59463a,a59466a,a59467a,a59470a,a59473a,a59474a,a59475a,a59478a,a59481a,a59482a,a59485a,a59488a,a59489a,a59490a,a59493a,a59496a,a59497a,a59500a,a59503a,a59504a,a59505a,a59508a,a59511a,a59512a,a59515a,a59518a,a59519a,a59520a,a59523a,a59526a,a59527a,a59530a,a59533a,a59534a,a59535a,a59538a,a59541a,a59542a,a59545a,a59548a,a59549a,a59550a,a59553a,a59556a,a59557a,a59560a,a59563a,a59564a,a59565a,a59568a,a59571a,a59572a,a59575a,a59578a,a59579a,a59580a,a59583a,a59586a,a59587a,a59590a,a59593a,a59594a,a59595a,a59598a,a59601a,a59602a,a59605a,a59608a,a59609a,a59610a,a59613a,a59616a,a59617a,a59620a,a59623a,a59624a,a59625a,a59628a,a59631a,a59632a,a59635a,a59638a,a59639a,a59640a,a59643a,a59646a,a59647a,a59650a,a59653a,a59654a,a59655a,a59658a,a59661a,a59662a,a59665a,a59668a,a59669a,a59670a,a59673a,a59676a,a59677a,a59680a,a59683a,a59684a,a59685a,a59688a,a59691a,a59692a,a59695a,a59698a,a59699a,a59700a,a59703a,a59706a,a59707a,a59710a,a59713a,a59714a,a59715a,a59718a,a59721a,a59722a,a59725a,a59728a,a59729a,a59730a,a59733a,a59736a,a59737a,a59740a,a59743a,a59744a,a59745a,a59748a,a59751a,a59752a,a59755a,a59758a,a59759a,a59760a,a59763a,a59766a,a59767a,a59770a,a59773a,a59774a,a59775a,a59778a,a59781a,a59782a,a59785a,a59788a,a59789a,a59790a,a59793a,a59796a,a59797a,a59800a,a59803a,a59804a,a59805a,a59808a,a59811a,a59812a,a59815a,a59818a,a59819a,a59820a,a59823a,a59826a,a59827a,a59830a,a59833a,a59834a,a59835a,a59838a,a59841a,a59842a,a59845a,a59848a,a59849a,a59850a,a59853a,a59856a,a59857a,a59860a,a59863a,a59864a,a59865a,a59868a,a59871a,a59872a,a59875a,a59878a,a59879a,a59880a,a59883a,a59886a,a59887a,a59890a,a59893a,a59894a,a59895a,a59898a,a59901a,a59902a,a59905a,a59908a,a59909a,a59910a,a59913a,a59916a,a59917a,a59920a,a59923a,a59924a,a59925a,a59928a,a59931a,a59932a,a59935a,a59938a,a59939a,a59940a,a59943a,a59946a,a59947a,a59950a,a59953a,a59954a,a59955a,a59958a,a59961a,a59962a,a59965a,a59968a,a59969a,a59970a,a59973a,a59976a,a59977a,a59980a,a59983a,a59984a,a59985a,a59988a,a59991a,a59992a,a59995a,a59998a,a59999a,a60000a,a60003a,a60006a,a60007a,a60010a,a60013a,a60014a,a60015a,a60018a,a60021a,a60022a,a60025a,a60028a,a60029a,a60030a,a60033a,a60036a,a60037a,a60040a,a60043a,a60044a,a60045a,a60048a,a60051a,a60052a,a60055a,a60058a,a60059a,a60060a,a60063a,a60066a,a60067a,a60070a,a60073a,a60074a,a60075a,a60078a,a60081a,a60082a,a60085a,a60088a,a60089a,a60090a,a60093a,a60096a,a60097a,a60100a,a60103a,a60104a,a60105a,a60108a,a60111a,a60112a,a60115a,a60118a,a60119a,a60120a,a60123a,a60126a,a60127a,a60130a,a60133a,a60134a,a60135a,a60138a,a60141a,a60142a,a60145a,a60148a,a60149a,a60150a,a60153a,a60156a,a60157a,a60160a,a60163a,a60164a,a60165a,a60168a,a60171a,a60172a,a60175a,a60178a,a60179a,a60180a,a60183a,a60186a,a60187a,a60190a,a60193a,a60194a,a60195a,a60198a,a60201a,a60202a,a60205a,a60208a,a60209a,a60210a,a60213a,a60216a,a60217a,a60220a,a60223a,a60224a,a60225a,a60228a,a60231a,a60232a,a60235a,a60238a,a60239a,a60240a,a60243a,a60246a,a60247a,a60250a,a60253a,a60254a,a60255a,a60258a,a60261a,a60262a,a60265a,a60268a,a60269a,a60270a,a60273a,a60276a,a60277a,a60280a,a60283a,a60284a,a60285a,a60288a,a60291a,a60292a,a60295a,a60298a,a60299a,a60300a,a60303a,a60306a,a60307a,a60310a,a60313a,a60314a,a60315a,a60318a,a60321a,a60322a,a60325a,a60328a,a60329a,a60330a,a60333a,a60336a,a60337a,a60340a,a60343a,a60344a,a60345a,a60348a,a60351a,a60352a,a60355a,a60358a,a60359a,a60360a,a60363a,a60366a,a60367a,a60370a,a60373a,a60374a,a60375a,a60378a,a60381a,a60382a,a60385a,a60388a,a60389a,a60390a,a60393a,a60396a,a60397a,a60400a,a60403a,a60404a,a60405a,a60408a,a60411a,a60412a,a60415a,a60418a,a60419a,a60420a,a60423a,a60426a,a60427a,a60430a,a60433a,a60434a,a60435a,a60438a,a60441a,a60442a,a60445a,a60448a,a60449a,a60450a,a60453a,a60456a,a60457a,a60460a,a60463a,a60464a,a60465a,a60468a,a60471a,a60472a,a60475a,a60478a,a60479a,a60480a,a60483a,a60486a,a60487a,a60490a,a60493a,a60494a,a60495a,a60498a,a60501a,a60502a,a60505a,a60508a,a60509a,a60510a,a60513a,a60516a,a60517a,a60520a,a60523a,a60524a,a60525a,a60528a,a60531a,a60532a,a60535a,a60538a,a60539a,a60540a,a60543a,a60546a,a60547a,a60550a,a60553a,a60554a,a60555a,a60558a,a60561a,a60562a,a60565a,a60568a,a60569a,a60570a,a60573a,a60576a,a60577a,a60580a,a60583a,a60584a,a60585a,a60588a,a60591a,a60592a,a60595a,a60598a,a60599a,a60600a,a60603a,a60606a,a60607a,a60610a,a60613a,a60614a,a60615a,a60618a,a60621a,a60622a,a60625a,a60628a,a60629a,a60630a,a60633a,a60636a,a60637a,a60640a,a60643a,a60644a,a60645a,a60648a,a60651a,a60652a,a60655a,a60658a,a60659a,a60660a,a60663a,a60666a,a60667a,a60670a,a60673a,a60674a,a60675a,a60678a,a60681a,a60682a,a60685a,a60688a,a60689a,a60690a,a60693a,a60696a,a60697a,a60700a,a60703a,a60704a,a60705a,a60708a,a60711a,a60712a,a60715a,a60718a,a60719a,a60720a,a60723a,a60726a,a60727a,a60730a,a60733a,a60734a,a60735a,a60738a,a60741a,a60742a,a60745a,a60748a,a60749a,a60750a,a60753a,a60756a,a60757a,a60760a,a60763a,a60764a,a60765a,a60768a,a60771a,a60772a,a60775a,a60778a,a60779a,a60780a,a60783a,a60786a,a60787a,a60790a,a60793a,a60794a,a60795a,a60798a,a60801a,a60802a,a60805a,a60808a,a60809a,a60810a,a60813a,a60816a,a60817a,a60820a,a60823a,a60824a,a60825a,a60828a,a60831a,a60832a,a60835a,a60838a,a60839a,a60840a,a60843a,a60846a,a60847a,a60850a,a60853a,a60854a,a60855a,a60858a,a60861a,a60862a,a60865a,a60868a,a60869a,a60870a,a60873a,a60876a,a60877a,a60880a,a60883a,a60884a,a60885a,a60888a,a60891a,a60892a,a60895a,a60898a,a60899a,a60900a,a60903a,a60906a,a60907a,a60910a,a60913a,a60914a,a60915a,a60918a,a60921a,a60922a,a60925a,a60928a,a60929a,a60930a,a60933a,a60936a,a60937a,a60940a,a60943a,a60944a,a60945a,a60948a,a60951a,a60952a,a60955a,a60958a,a60959a,a60960a,a60963a,a60966a,a60967a,a60970a,a60973a,a60974a,a60975a,a60978a,a60981a,a60982a,a60985a,a60988a,a60989a,a60990a,a60993a,a60996a,a60997a,a61000a,a61003a,a61004a,a61005a,a61008a,a61011a,a61012a,a61015a,a61018a,a61019a,a61020a,a61023a,a61026a,a61027a,a61030a,a61033a,a61034a,a61035a,a61038a,a61041a,a61042a,a61045a,a61048a,a61049a,a61050a,a61053a,a61056a,a61057a,a61060a,a61063a,a61064a,a61065a,a61068a,a61071a,a61072a,a61075a,a61078a,a61079a,a61080a,a61083a,a61086a,a61087a,a61090a,a61093a,a61094a,a61095a,a61098a,a61101a,a61102a,a61105a,a61108a,a61109a,a61110a,a61113a,a61116a,a61117a,a61120a,a61123a,a61124a,a61125a,a61128a,a61131a,a61132a,a61135a,a61138a,a61139a,a61140a,a61143a,a61146a,a61147a,a61150a,a61153a,a61154a,a61155a,a61158a,a61161a,a61162a,a61165a,a61168a,a61169a,a61170a,a61173a,a61176a,a61177a,a61180a,a61183a,a61184a,a61185a,a61188a,a61191a,a61192a,a61195a,a61198a,a61199a,a61200a,a61203a,a61206a,a61207a,a61210a,a61213a,a61214a,a61215a,a61218a,a61221a,a61222a,a61225a,a61228a,a61229a,a61230a,a61233a,a61236a,a61237a,a61240a,a61243a,a61244a,a61245a,a61248a,a61251a,a61252a,a61255a,a61258a,a61259a,a61260a,a61263a,a61266a,a61267a,a61270a,a61273a,a61274a,a61275a,a61278a,a61281a,a61282a,a61285a,a61288a,a61289a,a61290a,a61293a,a61296a,a61297a,a61300a,a61303a,a61304a,a61305a,a61308a,a61311a,a61312a,a61315a,a61318a,a61319a,a61320a,a61323a,a61326a,a61327a,a61330a,a61333a,a61334a,a61335a,a61338a,a61341a,a61342a,a61345a,a61348a,a61349a,a61350a,a61353a,a61356a,a61357a,a61360a,a61363a,a61364a,a61365a,a61368a,a61371a,a61372a,a61375a,a61378a,a61379a,a61380a,a61383a,a61386a,a61387a,a61390a,a61393a,a61394a,a61395a,a61398a,a61401a,a61402a,a61405a,a61408a,a61409a,a61410a,a61413a,a61416a,a61417a,a61420a,a61423a,a61424a,a61425a,a61428a,a61431a,a61432a,a61435a,a61438a,a61439a,a61440a,a61443a,a61446a,a61447a,a61450a,a61453a,a61454a,a61455a,a61458a,a61461a,a61462a,a61465a,a61468a,a61469a,a61470a,a61473a,a61476a,a61477a,a61480a,a61483a,a61484a,a61485a,a61488a,a61491a,a61492a,a61495a,a61498a,a61499a,a61500a,a61503a,a61506a,a61507a,a61510a,a61513a,a61514a,a61515a,a61518a,a61521a,a61522a,a61525a,a61528a,a61529a,a61530a,a61533a,a61536a,a61537a,a61540a,a61543a,a61544a,a61545a,a61548a,a61551a,a61552a,a61555a,a61558a,a61559a,a61560a,a61563a,a61566a,a61567a,a61570a,a61573a,a61574a,a61575a,a61578a,a61581a,a61582a,a61585a,a61588a,a61589a,a61590a,a61593a,a61596a,a61597a,a61600a,a61603a,a61604a,a61605a,a61608a,a61611a,a61612a,a61615a,a61618a,a61619a,a61620a,a61623a,a61626a,a61627a,a61630a,a61633a,a61634a,a61635a,a61638a,a61641a,a61642a,a61645a,a61648a,a61649a,a61650a,a61653a,a61656a,a61657a,a61660a,a61663a,a61664a,a61665a,a61668a,a61671a,a61672a,a61675a,a61678a,a61679a,a61680a,a61683a,a61686a,a61687a,a61690a,a61693a,a61694a,a61695a,a61698a,a61701a,a61702a,a61705a,a61708a,a61709a,a61710a,a61713a,a61716a,a61717a,a61720a,a61723a,a61724a,a61725a,a61728a,a61731a,a61732a,a61735a,a61738a,a61739a,a61740a,a61743a,a61746a,a61747a,a61750a,a61753a,a61754a,a61755a,a61758a,a61761a,a61762a,a61765a,a61768a,a61769a,a61770a,a61773a,a61776a,a61777a,a61780a,a61783a,a61784a,a61785a,a61788a,a61791a,a61792a,a61795a,a61798a,a61799a,a61800a,a61803a,a61806a,a61807a,a61810a,a61813a,a61814a,a61815a,a61818a,a61821a,a61822a,a61825a,a61828a,a61829a,a61830a,a61833a,a61836a,a61837a,a61840a,a61843a,a61844a,a61845a,a61848a,a61851a,a61852a,a61855a,a61858a,a61859a,a61860a,a61863a,a61866a,a61867a,a61870a,a61873a,a61874a,a61875a,a61878a,a61881a,a61882a,a61885a,a61888a,a61889a,a61890a,a61893a,a61896a,a61897a,a61900a,a61903a,a61904a,a61905a,a61908a,a61911a,a61912a,a61915a,a61918a,a61919a,a61920a,a61923a,a61926a,a61927a,a61930a,a61933a,a61934a,a61935a,a61938a,a61941a,a61942a,a61945a,a61948a,a61949a,a61950a,a61953a,a61956a,a61957a,a61960a,a61963a,a61964a,a61965a,a61968a,a61971a,a61972a,a61975a,a61978a,a61979a,a61980a,a61983a,a61986a,a61987a,a61990a,a61993a,a61994a,a61995a,a61998a,a62001a,a62002a,a62005a,a62008a,a62009a,a62010a,a62013a,a62016a,a62017a,a62020a,a62023a,a62024a,a62025a,a62028a,a62031a,a62032a,a62035a,a62038a,a62039a,a62040a,a62043a,a62046a,a62047a,a62050a,a62053a,a62054a,a62055a,a62058a,a62061a,a62062a,a62065a,a62068a,a62069a,a62070a,a62073a,a62076a,a62077a,a62080a,a62083a,a62084a,a62085a,a62088a,a62091a,a62092a,a62095a,a62098a,a62099a,a62100a,a62103a,a62106a,a62107a,a62110a,a62113a,a62114a,a62115a,a62118a,a62121a,a62122a,a62125a,a62128a,a62129a,a62130a,a62133a,a62136a,a62137a,a62140a,a62143a,a62144a,a62145a,a62148a,a62151a,a62152a,a62155a,a62158a,a62159a,a62160a,a62163a,a62166a,a62167a,a62170a,a62173a,a62174a,a62175a,a62178a,a62181a,a62182a,a62185a,a62188a,a62189a,a62190a,a62193a,a62196a,a62197a,a62200a,a62203a,a62204a,a62205a,a62208a,a62211a,a62212a,a62215a,a62218a,a62219a,a62220a,a62223a,a62226a,a62227a,a62230a,a62233a,a62234a,a62235a,a62238a,a62241a,a62242a,a62245a,a62248a,a62249a,a62250a,a62253a,a62256a,a62257a,a62260a,a62263a,a62264a,a62265a,a62268a,a62271a,a62272a,a62275a,a62278a,a62279a,a62280a,a62283a,a62286a,a62287a,a62290a,a62293a,a62294a,a62295a,a62298a,a62301a,a62302a,a62305a,a62308a,a62309a,a62310a,a62313a,a62316a,a62317a,a62320a,a62323a,a62324a,a62325a,a62328a,a62331a,a62332a,a62335a,a62338a,a62339a,a62340a,a62343a,a62346a,a62347a,a62350a,a62353a,a62354a,a62355a,a62358a,a62361a,a62362a,a62365a,a62368a,a62369a,a62370a,a62373a,a62376a,a62377a,a62380a,a62383a,a62384a,a62385a,a62388a,a62391a,a62392a,a62395a,a62398a,a62399a,a62400a,a62403a,a62406a,a62407a,a62410a,a62413a,a62414a,a62415a,a62418a,a62421a,a62422a,a62425a,a62428a,a62429a,a62430a,a62433a,a62436a,a62437a,a62440a,a62443a,a62444a,a62445a,a62448a,a62451a,a62452a,a62455a,a62458a,a62459a,a62460a,a62463a,a62466a,a62467a,a62470a,a62473a,a62474a,a62475a,a62478a,a62481a,a62482a,a62485a,a62488a,a62489a,a62490a,a62493a,a62496a,a62497a,a62500a,a62503a,a62504a,a62505a,a62508a,a62511a,a62512a,a62515a,a62518a,a62519a,a62520a,a62523a,a62526a,a62527a,a62530a,a62533a,a62534a,a62535a,a62538a,a62541a,a62542a,a62545a,a62548a,a62549a,a62550a,a62553a,a62556a,a62557a,a62560a,a62563a,a62564a,a62565a,a62568a,a62571a,a62572a,a62575a,a62578a,a62579a,a62580a,a62583a,a62586a,a62587a,a62590a,a62593a,a62594a,a62595a,a62598a,a62601a,a62602a,a62605a,a62609a,a62610a,a62611a,a62612a,a62615a,a62618a,a62619a,a62622a,a62625a,a62626a,a62627a,a62630a,a62633a,a62634a,a62637a,a62641a,a62642a,a62643a,a62644a,a62647a,a62650a,a62651a,a62654a,a62657a,a62658a,a62659a,a62662a,a62665a,a62666a,a62669a,a62673a,a62674a,a62675a,a62676a,a62679a,a62682a,a62683a,a62686a,a62689a,a62690a,a62691a,a62694a,a62697a,a62698a,a62701a,a62705a,a62706a,a62707a,a62708a,a62711a,a62714a,a62715a,a62718a,a62721a,a62722a,a62723a,a62726a,a62729a,a62730a,a62733a,a62737a,a62738a,a62739a,a62740a,a62743a,a62746a,a62747a,a62750a,a62753a,a62754a,a62755a,a62758a,a62761a,a62762a,a62765a,a62769a,a62770a,a62771a,a62772a,a62775a,a62778a,a62779a,a62782a,a62785a,a62786a,a62787a,a62790a,a62793a,a62794a,a62797a,a62801a,a62802a,a62803a,a62804a,a62807a,a62810a,a62811a,a62814a,a62817a,a62818a,a62819a,a62822a,a62825a,a62826a,a62829a,a62833a,a62834a,a62835a,a62836a,a62839a,a62842a,a62843a,a62846a,a62849a,a62850a,a62851a,a62854a,a62857a,a62858a,a62861a,a62865a,a62866a,a62867a,a62868a,a62871a,a62874a,a62875a,a62878a,a62881a,a62882a,a62883a,a62886a,a62889a,a62890a,a62893a,a62897a,a62898a,a62899a,a62900a,a62903a,a62906a,a62907a,a62910a,a62913a,a62914a,a62915a,a62918a,a62921a,a62922a,a62925a,a62929a,a62930a,a62931a,a62932a,a62935a,a62938a,a62939a,a62942a,a62945a,a62946a,a62947a,a62950a,a62953a,a62954a,a62957a,a62961a,a62962a,a62963a,a62964a,a62967a,a62970a,a62971a,a62974a,a62977a,a62978a,a62979a,a62982a,a62985a,a62986a,a62989a,a62993a,a62994a,a62995a,a62996a,a62999a,a63002a,a63003a,a63006a,a63009a,a63010a,a63011a,a63014a,a63017a,a63018a,a63021a,a63025a,a63026a,a63027a,a63028a,a63031a,a63034a,a63035a,a63038a,a63041a,a63042a,a63043a,a63046a,a63049a,a63050a,a63053a,a63057a,a63058a,a63059a,a63060a,a63063a,a63066a,a63067a,a63070a,a63073a,a63074a,a63075a,a63078a,a63081a,a63082a,a63085a,a63089a,a63090a,a63091a,a63092a,a63095a,a63098a,a63099a,a63102a,a63105a,a63106a,a63107a,a63110a,a63113a,a63114a,a63117a,a63121a,a63122a,a63123a,a63124a,a63127a,a63130a,a63131a,a63134a,a63137a,a63138a,a63139a,a63142a,a63145a,a63146a,a63149a,a63153a,a63154a,a63155a,a63156a,a63159a,a63162a,a63163a,a63166a,a63169a,a63170a,a63171a,a63174a,a63177a,a63178a,a63181a,a63185a,a63186a,a63187a,a63188a,a63191a,a63194a,a63195a,a63198a,a63201a,a63202a,a63203a,a63206a,a63209a,a63210a,a63213a,a63217a,a63218a,a63219a,a63220a,a63223a,a63226a,a63227a,a63230a,a63233a,a63234a,a63235a,a63238a,a63241a,a63242a,a63245a,a63249a,a63250a,a63251a,a63252a,a63255a,a63258a,a63259a,a63262a,a63265a,a63266a,a63267a,a63270a,a63273a,a63274a,a63277a,a63281a,a63282a,a63283a,a63284a,a63287a,a63290a,a63291a,a63294a,a63297a,a63298a,a63299a,a63302a,a63305a,a63306a,a63309a,a63313a,a63314a,a63315a,a63316a,a63319a,a63322a,a63323a,a63326a,a63329a,a63330a,a63331a,a63334a,a63337a,a63338a,a63341a,a63345a,a63346a,a63347a,a63348a,a63351a,a63354a,a63355a,a63358a,a63361a,a63362a,a63363a,a63366a,a63369a,a63370a,a63373a,a63377a,a63378a,a63379a,a63380a,a63383a,a63386a,a63387a,a63390a,a63393a,a63394a,a63395a,a63398a,a63401a,a63402a,a63405a,a63409a,a63410a,a63411a,a63412a,a63415a,a63418a,a63419a,a63422a,a63425a,a63426a,a63427a,a63430a,a63433a,a63434a,a63437a,a63441a,a63442a,a63443a,a63444a,a63447a,a63450a,a63451a,a63454a,a63457a,a63458a,a63459a,a63462a,a63465a,a63466a,a63469a,a63473a,a63474a,a63475a,a63476a,a63479a,a63482a,a63483a,a63486a,a63489a,a63490a,a63491a,a63494a,a63497a,a63498a,a63501a,a63505a,a63506a,a63507a,a63508a,a63511a,a63514a,a63515a,a63518a,a63521a,a63522a,a63523a,a63526a,a63529a,a63530a,a63533a,a63537a,a63538a,a63539a,a63540a,a63543a,a63546a,a63547a,a63550a,a63553a,a63554a,a63555a,a63558a,a63561a,a63562a,a63565a,a63569a,a63570a,a63571a,a63572a,a63575a,a63578a,a63579a,a63582a,a63585a,a63586a,a63587a,a63590a,a63593a,a63594a,a63597a,a63601a,a63602a,a63603a,a63604a,a63607a,a63610a,a63611a,a63614a,a63617a,a63618a,a63619a,a63622a,a63625a,a63626a,a63629a,a63633a,a63634a,a63635a,a63636a,a63639a,a63642a,a63643a,a63646a,a63649a,a63650a,a63651a,a63654a,a63657a,a63658a,a63661a,a63665a,a63666a,a63667a,a63668a,a63671a,a63674a,a63675a,a63678a,a63681a,a63682a,a63683a,a63686a,a63689a,a63690a,a63693a,a63697a,a63698a,a63699a,a63700a,a63703a,a63706a,a63707a,a63710a,a63713a,a63714a,a63715a,a63718a,a63721a,a63722a,a63725a,a63729a,a63730a,a63731a,a63732a,a63735a,a63738a,a63739a,a63742a,a63745a,a63746a,a63747a,a63750a,a63753a,a63754a,a63757a,a63761a,a63762a,a63763a,a63764a,a63767a,a63770a,a63771a,a63774a,a63777a,a63778a,a63779a,a63782a,a63785a,a63786a,a63789a,a63793a,a63794a,a63795a,a63796a,a63799a,a63802a,a63803a,a63806a,a63809a,a63810a,a63811a,a63814a,a63817a,a63818a,a63821a,a63825a,a63826a,a63827a,a63828a,a63831a,a63834a,a63835a,a63838a,a63841a,a63842a,a63843a,a63846a,a63849a,a63850a,a63853a,a63857a,a63858a,a63859a,a63860a,a63863a,a63866a,a63867a,a63870a,a63873a,a63874a,a63875a,a63878a,a63881a,a63882a,a63885a,a63889a,a63890a,a63891a,a63892a,a63895a,a63898a,a63899a,a63902a,a63905a,a63906a,a63907a,a63910a,a63913a,a63914a,a63917a,a63921a,a63922a,a63923a,a63924a,a63927a,a63930a,a63931a,a63934a,a63937a,a63938a,a63939a,a63942a,a63945a,a63946a,a63949a,a63953a,a63954a,a63955a,a63956a,a63959a,a63962a,a63963a,a63966a,a63969a,a63970a,a63971a,a63974a,a63977a,a63978a,a63981a,a63985a,a63986a,a63987a,a63988a,a63991a,a63994a,a63995a,a63998a,a64001a,a64002a,a64003a,a64006a,a64009a,a64010a,a64013a,a64017a,a64018a,a64019a,a64020a,a64023a,a64026a,a64027a,a64030a,a64033a,a64034a,a64035a,a64038a,a64041a,a64042a,a64045a,a64049a,a64050a,a64051a,a64052a,a64055a,a64058a,a64059a,a64062a,a64065a,a64066a,a64067a,a64070a,a64073a,a64074a,a64077a,a64081a,a64082a,a64083a,a64084a,a64087a,a64090a,a64091a,a64094a,a64097a,a64098a,a64099a,a64102a,a64105a,a64106a,a64109a,a64113a,a64114a,a64115a,a64116a,a64119a,a64122a,a64123a,a64126a,a64129a,a64130a,a64131a,a64134a,a64137a,a64138a,a64141a,a64145a,a64146a,a64147a,a64148a,a64151a,a64154a,a64155a,a64158a,a64161a,a64162a,a64163a,a64166a,a64169a,a64170a,a64173a,a64177a,a64178a,a64179a,a64180a,a64183a,a64186a,a64187a,a64190a,a64193a,a64194a,a64195a,a64198a,a64201a,a64202a,a64205a,a64209a,a64210a,a64211a,a64212a,a64215a,a64218a,a64219a,a64222a,a64225a,a64226a,a64227a,a64230a,a64233a,a64234a,a64237a,a64241a,a64242a,a64243a,a64244a,a64247a,a64250a,a64251a,a64254a,a64257a,a64258a,a64259a,a64262a,a64265a,a64266a,a64269a,a64273a,a64274a,a64275a,a64276a,a64279a,a64282a,a64283a,a64286a,a64289a,a64290a,a64291a,a64294a,a64297a,a64298a,a64301a,a64305a,a64306a,a64307a,a64308a,a64311a,a64314a,a64315a,a64318a,a64321a,a64322a,a64323a,a64326a,a64329a,a64330a,a64333a,a64337a,a64338a,a64339a,a64340a,a64343a,a64346a,a64347a,a64350a,a64353a,a64354a,a64355a,a64358a,a64361a,a64362a,a64365a,a64369a,a64370a,a64371a,a64372a,a64375a,a64378a,a64379a,a64382a,a64385a,a64386a,a64387a,a64390a,a64393a,a64394a,a64397a,a64401a,a64402a,a64403a,a64404a,a64407a,a64410a,a64411a,a64414a,a64417a,a64418a,a64419a,a64422a,a64425a,a64426a,a64429a,a64433a,a64434a,a64435a,a64436a,a64439a,a64442a,a64443a,a64446a,a64449a,a64450a,a64451a,a64454a,a64457a,a64458a,a64461a,a64465a,a64466a,a64467a,a64468a,a64471a,a64474a,a64475a,a64478a,a64481a,a64482a,a64483a,a64486a,a64489a,a64490a,a64493a,a64497a,a64498a,a64499a,a64500a,a64503a,a64506a,a64507a,a64510a,a64513a,a64514a,a64515a,a64518a,a64521a,a64522a,a64525a,a64529a,a64530a,a64531a,a64532a,a64535a,a64538a,a64539a,a64542a,a64545a,a64546a,a64547a,a64550a,a64553a,a64554a,a64557a,a64561a,a64562a,a64563a,a64564a,a64567a,a64570a,a64571a,a64574a,a64577a,a64578a,a64579a,a64582a,a64585a,a64586a,a64589a,a64593a,a64594a,a64595a,a64596a,a64599a,a64602a,a64603a,a64606a,a64609a,a64610a,a64611a,a64614a,a64617a,a64618a,a64621a,a64625a,a64626a,a64627a,a64628a,a64631a,a64634a,a64635a,a64638a,a64641a,a64642a,a64643a,a64646a,a64649a,a64650a,a64653a,a64657a,a64658a,a64659a,a64660a,a64663a,a64666a,a64667a,a64670a,a64673a,a64674a,a64675a,a64678a,a64681a,a64682a,a64685a,a64689a,a64690a,a64691a,a64692a,a64695a,a64698a,a64699a,a64702a,a64705a,a64706a,a64707a,a64710a,a64713a,a64714a,a64717a,a64721a,a64722a,a64723a,a64724a,a64727a,a64730a,a64731a,a64734a,a64737a,a64738a,a64739a,a64742a,a64745a,a64746a,a64749a,a64753a,a64754a,a64755a,a64756a,a64759a,a64762a,a64763a,a64766a,a64769a,a64770a,a64771a,a64774a,a64777a,a64778a,a64781a,a64785a,a64786a,a64787a,a64788a,a64791a,a64794a,a64795a,a64798a,a64801a,a64802a,a64803a,a64806a,a64809a,a64810a,a64813a,a64817a,a64818a,a64819a,a64820a,a64823a,a64826a,a64827a,a64830a,a64833a,a64834a,a64835a,a64838a,a64841a,a64842a,a64845a,a64849a,a64850a,a64851a,a64852a,a64855a,a64858a,a64859a,a64862a,a64865a,a64866a,a64867a,a64870a,a64873a,a64874a,a64877a,a64881a,a64882a,a64883a,a64884a,a64887a,a64890a,a64891a,a64894a,a64897a,a64898a,a64899a,a64902a,a64905a,a64906a,a64909a,a64913a,a64914a,a64915a,a64916a,a64919a,a64922a,a64923a,a64926a,a64929a,a64930a,a64931a,a64934a,a64937a,a64938a,a64941a,a64945a,a64946a,a64947a,a64948a,a64951a,a64954a,a64955a,a64958a,a64961a,a64962a,a64963a,a64966a,a64969a,a64970a,a64973a,a64977a,a64978a,a64979a,a64980a,a64983a,a64986a,a64987a,a64990a,a64993a,a64994a,a64995a,a64998a,a65001a,a65002a,a65005a,a65009a,a65010a,a65011a,a65012a,a65015a,a65018a,a65019a,a65022a,a65025a,a65026a,a65027a,a65030a,a65033a,a65034a,a65037a,a65041a,a65042a,a65043a,a65044a,a65047a,a65050a,a65051a,a65054a,a65057a,a65058a,a65059a,a65062a,a65065a,a65066a,a65069a,a65073a,a65074a,a65075a,a65076a,a65079a,a65082a,a65083a,a65086a,a65089a,a65090a,a65091a,a65094a,a65097a,a65098a,a65101a,a65105a,a65106a,a65107a,a65108a,a65111a,a65114a,a65115a,a65118a,a65121a,a65122a,a65123a,a65126a,a65129a,a65130a,a65133a,a65137a,a65138a,a65139a,a65140a,a65143a,a65146a,a65147a,a65150a,a65153a,a65154a,a65155a,a65158a,a65161a,a65162a,a65165a,a65169a,a65170a,a65171a,a65172a,a65175a,a65178a,a65179a,a65182a,a65185a,a65186a,a65187a,a65190a,a65193a,a65194a,a65197a,a65201a,a65202a,a65203a,a65204a,a65207a,a65210a,a65211a,a65214a,a65217a,a65218a,a65219a,a65222a,a65225a,a65226a,a65229a,a65233a,a65234a,a65235a,a65236a,a65239a,a65242a,a65243a,a65246a,a65249a,a65250a,a65251a,a65254a,a65257a,a65258a,a65261a,a65265a,a65266a,a65267a,a65268a,a65271a,a65274a,a65275a,a65278a,a65281a,a65282a,a65283a,a65286a,a65289a,a65290a,a65293a,a65297a,a65298a,a65299a,a65300a,a65303a,a65306a,a65307a,a65310a,a65313a,a65314a,a65315a,a65318a,a65321a,a65322a,a65325a,a65329a,a65330a,a65331a,a65332a,a65335a,a65338a,a65339a,a65342a,a65345a,a65346a,a65347a,a65350a,a65353a,a65354a,a65357a,a65361a,a65362a,a65363a,a65364a,a65367a,a65370a,a65371a,a65374a,a65377a,a65378a,a65379a,a65382a,a65385a,a65386a,a65389a,a65393a,a65394a,a65395a,a65396a,a65399a,a65402a,a65403a,a65406a,a65409a,a65410a,a65411a,a65414a,a65417a,a65418a,a65421a,a65425a,a65426a,a65427a,a65428a,a65431a,a65434a,a65435a,a65438a,a65441a,a65442a,a65443a,a65446a,a65449a,a65450a,a65453a,a65457a,a65458a,a65459a,a65460a,a65463a,a65466a,a65467a,a65470a,a65473a,a65474a,a65475a,a65478a,a65481a,a65482a,a65485a,a65489a,a65490a,a65491a,a65492a,a65495a,a65498a,a65499a,a65502a,a65505a,a65506a,a65507a,a65510a,a65513a,a65514a,a65517a,a65521a,a65522a,a65523a,a65524a,a65527a,a65530a,a65531a,a65534a,a65537a,a65538a,a65539a,a65542a,a65545a,a65546a,a65549a,a65553a,a65554a,a65555a,a65556a,a65559a,a65562a,a65563a,a65566a,a65569a,a65570a,a65571a,a65574a,a65577a,a65578a,a65581a,a65585a,a65586a,a65587a,a65588a,a65591a,a65594a,a65595a,a65598a,a65601a,a65602a,a65603a,a65606a,a65609a,a65610a,a65613a,a65617a,a65618a,a65619a,a65620a,a65623a,a65626a,a65627a,a65630a,a65633a,a65634a,a65635a,a65638a,a65641a,a65642a,a65645a,a65649a,a65650a,a65651a,a65652a,a65655a,a65658a,a65659a,a65662a,a65665a,a65666a,a65667a,a65670a,a65673a,a65674a,a65677a,a65681a,a65682a,a65683a,a65684a,a65687a,a65690a,a65691a,a65694a,a65697a,a65698a,a65699a,a65702a,a65705a,a65706a,a65709a,a65713a,a65714a,a65715a,a65716a,a65719a,a65722a,a65723a,a65726a,a65729a,a65730a,a65731a,a65734a,a65737a,a65738a,a65741a,a65745a,a65746a,a65747a,a65748a,a65751a,a65754a,a65755a,a65758a,a65761a,a65762a,a65763a,a65766a,a65769a,a65770a,a65773a,a65777a,a65778a,a65779a,a65780a,a65783a,a65786a,a65787a,a65790a,a65793a,a65794a,a65795a,a65798a,a65801a,a65802a,a65805a,a65809a,a65810a,a65811a,a65812a,a65815a,a65818a,a65819a,a65822a,a65825a,a65826a,a65827a,a65830a,a65833a,a65834a,a65837a,a65841a,a65842a,a65843a,a65844a,a65847a,a65850a,a65851a,a65854a,a65857a,a65858a,a65859a,a65862a,a65865a,a65866a,a65869a,a65873a,a65874a,a65875a,a65876a,a65879a,a65882a,a65883a,a65886a,a65889a,a65890a,a65891a,a65894a,a65897a,a65898a,a65901a,a65905a,a65906a,a65907a,a65908a,a65911a,a65914a,a65915a,a65918a,a65921a,a65922a,a65923a,a65926a,a65929a,a65930a,a65933a,a65937a,a65938a,a65939a,a65940a,a65943a,a65946a,a65947a,a65950a,a65953a,a65954a,a65955a,a65958a,a65961a,a65962a,a65965a,a65969a,a65970a,a65971a,a65972a,a65975a,a65978a,a65979a,a65982a,a65985a,a65986a,a65987a,a65990a,a65993a,a65994a,a65997a,a66001a,a66002a,a66003a,a66004a,a66007a,a66010a,a66011a,a66014a,a66017a,a66018a,a66019a,a66022a,a66025a,a66026a,a66029a,a66033a,a66034a,a66035a,a66036a,a66039a,a66042a,a66043a,a66046a,a66049a,a66050a,a66051a,a66054a,a66057a,a66058a,a66061a,a66065a,a66066a,a66067a,a66068a,a66071a,a66074a,a66075a,a66078a,a66081a,a66082a,a66083a,a66086a,a66089a,a66090a,a66093a,a66097a,a66098a,a66099a,a66100a,a66103a,a66106a,a66107a,a66110a,a66113a,a66114a,a66115a,a66118a,a66121a,a66122a,a66125a,a66129a,a66130a,a66131a,a66132a,a66135a,a66138a,a66139a,a66142a,a66145a,a66146a,a66147a,a66150a,a66153a,a66154a,a66157a,a66161a,a66162a,a66163a,a66164a,a66167a,a66170a,a66171a,a66174a,a66177a,a66178a,a66179a,a66182a,a66185a,a66186a,a66189a,a66193a,a66194a,a66195a,a66196a,a66199a,a66202a,a66203a,a66206a,a66209a,a66210a,a66211a,a66214a,a66217a,a66218a,a66221a,a66225a,a66226a,a66227a,a66228a,a66231a,a66234a,a66235a,a66238a,a66241a,a66242a,a66243a,a66246a,a66249a,a66250a,a66253a,a66257a,a66258a,a66259a,a66260a,a66263a,a66266a,a66267a,a66270a,a66273a,a66274a,a66275a,a66278a,a66281a,a66282a,a66285a,a66289a,a66290a,a66291a,a66292a,a66295a,a66298a,a66299a,a66302a,a66305a,a66306a,a66307a,a66310a,a66313a,a66314a,a66317a,a66321a,a66322a,a66323a,a66324a,a66327a,a66330a,a66331a,a66334a,a66337a,a66338a,a66339a,a66342a,a66345a,a66346a,a66349a,a66353a,a66354a,a66355a,a66356a,a66359a,a66362a,a66363a,a66366a,a66369a,a66370a,a66371a,a66374a,a66377a,a66378a,a66381a,a66385a,a66386a,a66387a,a66388a,a66391a,a66394a,a66395a,a66398a,a66401a,a66402a,a66403a,a66406a,a66409a,a66410a,a66413a,a66417a,a66418a,a66419a,a66420a,a66423a,a66426a,a66427a,a66430a,a66433a,a66434a,a66435a,a66438a,a66441a,a66442a,a66445a,a66449a,a66450a,a66451a,a66452a,a66455a,a66458a,a66459a,a66462a,a66465a,a66466a,a66467a,a66470a,a66473a,a66474a,a66477a,a66481a,a66482a,a66483a,a66484a,a66487a,a66490a,a66491a,a66494a,a66497a,a66498a,a66499a,a66502a,a66505a,a66506a,a66509a,a66513a,a66514a,a66515a,a66516a,a66519a,a66522a,a66523a,a66526a,a66529a,a66530a,a66531a,a66534a,a66537a,a66538a,a66541a,a66545a,a66546a,a66547a,a66548a,a66551a,a66554a,a66555a,a66558a,a66561a,a66562a,a66563a,a66566a,a66569a,a66570a,a66573a,a66577a,a66578a,a66579a,a66580a,a66583a,a66586a,a66587a,a66590a,a66593a,a66594a,a66595a,a66598a,a66601a,a66602a,a66605a,a66609a,a66610a,a66611a,a66612a,a66615a,a66618a,a66619a,a66622a,a66625a,a66626a,a66627a,a66630a,a66633a,a66634a,a66637a,a66641a,a66642a,a66643a,a66644a,a66647a,a66650a,a66651a,a66654a,a66657a,a66658a,a66659a,a66662a,a66665a,a66666a,a66669a,a66673a,a66674a,a66675a,a66676a,a66679a,a66682a,a66683a,a66686a,a66689a,a66690a,a66691a,a66694a,a66697a,a66698a,a66701a,a66705a,a66706a,a66707a,a66708a,a66711a,a66714a,a66715a,a66718a,a66721a,a66722a,a66723a,a66726a,a66729a,a66730a,a66733a,a66737a,a66738a,a66739a,a66740a,a66743a,a66746a,a66747a,a66750a,a66753a,a66754a,a66755a,a66758a,a66761a,a66762a,a66765a,a66769a,a66770a,a66771a,a66772a,a66775a,a66778a,a66779a,a66782a,a66785a,a66786a,a66787a,a66790a,a66793a,a66794a,a66797a,a66801a,a66802a,a66803a,a66804a,a66807a,a66810a,a66811a,a66814a,a66817a,a66818a,a66819a,a66822a,a66825a,a66826a,a66829a,a66833a,a66834a,a66835a,a66836a,a66839a,a66842a,a66843a,a66846a,a66849a,a66850a,a66851a,a66854a,a66857a,a66858a,a66861a,a66865a,a66866a,a66867a,a66868a,a66871a,a66874a,a66875a,a66878a,a66881a,a66882a,a66883a,a66886a,a66889a,a66890a,a66893a,a66897a,a66898a,a66899a,a66900a,a66903a,a66906a,a66907a,a66910a,a66913a,a66914a,a66915a,a66918a,a66921a,a66922a,a66925a,a66929a,a66930a,a66931a,a66932a,a66935a,a66938a,a66939a,a66942a,a66945a,a66946a,a66947a,a66950a,a66953a,a66954a,a66957a,a66961a,a66962a,a66963a,a66964a,a66967a,a66970a,a66971a,a66974a,a66977a,a66978a,a66979a,a66982a,a66985a,a66986a,a66989a,a66993a,a66994a,a66995a,a66996a,a66999a,a67002a,a67003a,a67006a,a67009a,a67010a,a67011a,a67014a,a67017a,a67018a,a67021a,a67025a,a67026a,a67027a,a67028a,a67031a,a67034a,a67035a,a67038a,a67041a,a67042a,a67043a,a67046a,a67049a,a67050a,a67053a,a67057a,a67058a,a67059a,a67060a,a67063a,a67066a,a67067a,a67070a,a67073a,a67074a,a67075a,a67078a,a67081a,a67082a,a67085a,a67089a,a67090a,a67091a,a67092a,a67095a,a67098a,a67099a,a67102a,a67105a,a67106a,a67107a,a67110a,a67113a,a67114a,a67117a,a67121a,a67122a,a67123a,a67124a,a67127a,a67130a,a67131a,a67134a,a67137a,a67138a,a67139a,a67142a,a67145a,a67146a,a67149a,a67153a,a67154a,a67155a,a67156a,a67159a,a67162a,a67163a,a67166a,a67169a,a67170a,a67171a,a67174a,a67177a,a67178a,a67181a,a67185a,a67186a,a67187a,a67188a,a67191a,a67194a,a67195a,a67198a,a67201a,a67202a,a67203a,a67206a,a67209a,a67210a,a67213a,a67217a,a67218a,a67219a,a67220a,a67223a,a67226a,a67227a,a67230a,a67233a,a67234a,a67235a,a67238a,a67241a,a67242a,a67245a,a67249a,a67250a,a67251a,a67252a,a67255a,a67258a,a67259a,a67262a,a67265a,a67266a,a67267a,a67270a,a67273a,a67274a,a67277a,a67281a,a67282a,a67283a,a67284a,a67287a,a67290a,a67291a,a67294a,a67297a,a67298a,a67299a,a67302a,a67305a,a67306a,a67309a,a67313a,a67314a,a67315a,a67316a,a67319a,a67322a,a67323a,a67326a,a67329a,a67330a,a67331a,a67334a,a67337a,a67338a,a67341a,a67345a,a67346a,a67347a,a67348a,a67351a,a67354a,a67355a,a67358a,a67361a,a67362a,a67363a,a67366a,a67369a,a67370a,a67373a,a67377a,a67378a,a67379a,a67380a,a67383a,a67386a,a67387a,a67390a,a67393a,a67394a,a67395a,a67398a,a67401a,a67402a,a67405a,a67409a,a67410a,a67411a,a67412a,a67415a,a67418a,a67419a,a67422a,a67425a,a67426a,a67427a,a67430a,a67433a,a67434a,a67437a,a67441a,a67442a,a67443a,a67444a,a67447a,a67450a,a67451a,a67454a,a67457a,a67458a,a67459a,a67462a,a67465a,a67466a,a67469a,a67473a,a67474a,a67475a,a67476a,a67479a,a67482a,a67483a,a67486a,a67489a,a67490a,a67491a,a67494a,a67497a,a67498a,a67501a,a67505a,a67506a,a67507a,a67508a,a67511a,a67514a,a67515a,a67518a,a67521a,a67522a,a67523a,a67526a,a67529a,a67530a,a67533a,a67537a,a67538a,a67539a,a67540a,a67543a,a67546a,a67547a,a67550a,a67553a,a67554a,a67555a,a67558a,a67561a,a67562a,a67565a,a67569a,a67570a,a67571a,a67572a,a67575a,a67578a,a67579a,a67582a,a67585a,a67586a,a67587a,a67590a,a67593a,a67594a,a67597a,a67601a,a67602a,a67603a,a67604a,a67607a,a67610a,a67611a,a67614a,a67617a,a67618a,a67619a,a67622a,a67625a,a67626a,a67629a,a67633a,a67634a,a67635a,a67636a,a67639a,a67642a,a67643a,a67646a,a67649a,a67650a,a67651a,a67654a,a67657a,a67658a,a67661a,a67665a,a67666a,a67667a,a67668a,a67671a,a67674a,a67675a,a67678a,a67681a,a67682a,a67683a,a67686a,a67689a,a67690a,a67693a,a67697a,a67698a,a67699a,a67700a,a67703a,a67706a,a67707a,a67710a,a67714a,a67715a,a67716a,a67717a,a67720a,a67723a,a67724a,a67727a,a67731a,a67732a,a67733a,a67734a,a67737a,a67740a,a67741a,a67744a,a67748a,a67749a,a67750a,a67751a,a67754a,a67757a,a67758a,a67761a,a67765a,a67766a,a67767a,a67768a,a67771a,a67774a,a67775a,a67778a,a67782a,a67783a,a67784a,a67785a,a67788a,a67791a,a67792a,a67795a,a67799a,a67800a,a67801a,a67802a,a67805a,a67808a,a67809a,a67812a,a67816a,a67817a,a67818a,a67819a,a67822a,a67825a,a67826a,a67829a,a67833a,a67834a,a67835a,a67836a,a67839a,a67842a,a67843a,a67846a,a67850a,a67851a,a67852a,a67853a,a67856a,a67859a,a67860a,a67863a,a67867a,a67868a,a67869a,a67870a,a67873a,a67876a,a67877a,a67880a,a67884a,a67885a,a67886a,a67887a,a67890a,a67893a,a67894a,a67897a,a67901a,a67902a,a67903a,a67904a,a67907a,a67910a,a67911a,a67914a,a67918a,a67919a,a67920a,a67921a,a67924a,a67927a,a67928a,a67931a,a67935a,a67936a,a67937a,a67938a,a67941a,a67944a,a67945a,a67948a,a67952a,a67953a,a67954a,a67955a,a67958a,a67961a,a67962a,a67965a,a67969a,a67970a,a67971a,a67972a,a67975a,a67978a,a67979a,a67982a,a67986a,a67987a,a67988a,a67989a,a67992a,a67995a,a67996a,a67999a,a68003a,a68004a,a68005a,a68006a,a68009a,a68012a,a68013a,a68016a,a68020a,a68021a,a68022a,a68023a,a68026a,a68029a,a68030a,a68033a,a68037a,a68038a,a68039a,a68040a,a68043a,a68046a,a68047a,a68050a,a68054a,a68055a,a68056a,a68057a,a68060a,a68063a,a68064a,a68067a,a68071a,a68072a,a68073a,a68074a,a68077a,a68080a,a68081a,a68084a,a68088a,a68089a,a68090a,a68091a,a68094a,a68097a,a68098a,a68101a,a68105a,a68106a,a68107a,a68108a,a68111a,a68114a,a68115a,a68118a,a68122a,a68123a,a68124a,a68125a,a68128a,a68131a,a68132a,a68135a,a68139a,a68140a,a68141a,a68142a,a68145a,a68148a,a68149a,a68152a,a68156a,a68157a,a68158a,a68159a,a68162a,a68165a,a68166a,a68169a,a68173a,a68174a,a68175a,a68176a,a68179a,a68182a,a68183a,a68186a,a68190a,a68191a,a68192a,a68193a,a68196a,a68199a,a68200a,a68203a,a68207a,a68208a,a68209a,a68210a,a68213a,a68216a,a68217a,a68220a,a68224a,a68225a,a68226a,a68227a,a68230a,a68233a,a68234a,a68237a,a68241a,a68242a,a68243a,a68244a: std_logic;
begin

A141 <=( a6568a ) or ( a4379a );
 a1a <=( a68244a  and  a68227a );
 a2a <=( a68210a  and  a68193a );
 a3a <=( a68176a  and  a68159a );
 a4a <=( a68142a  and  a68125a );
 a5a <=( a68108a  and  a68091a );
 a6a <=( a68074a  and  a68057a );
 a7a <=( a68040a  and  a68023a );
 a8a <=( a68006a  and  a67989a );
 a9a <=( a67972a  and  a67955a );
 a10a <=( a67938a  and  a67921a );
 a11a <=( a67904a  and  a67887a );
 a12a <=( a67870a  and  a67853a );
 a13a <=( a67836a  and  a67819a );
 a14a <=( a67802a  and  a67785a );
 a15a <=( a67768a  and  a67751a );
 a16a <=( a67734a  and  a67717a );
 a17a <=( a67700a  and  a67683a );
 a18a <=( a67668a  and  a67651a );
 a19a <=( a67636a  and  a67619a );
 a20a <=( a67604a  and  a67587a );
 a21a <=( a67572a  and  a67555a );
 a22a <=( a67540a  and  a67523a );
 a23a <=( a67508a  and  a67491a );
 a24a <=( a67476a  and  a67459a );
 a25a <=( a67444a  and  a67427a );
 a26a <=( a67412a  and  a67395a );
 a27a <=( a67380a  and  a67363a );
 a28a <=( a67348a  and  a67331a );
 a29a <=( a67316a  and  a67299a );
 a30a <=( a67284a  and  a67267a );
 a31a <=( a67252a  and  a67235a );
 a32a <=( a67220a  and  a67203a );
 a33a <=( a67188a  and  a67171a );
 a34a <=( a67156a  and  a67139a );
 a35a <=( a67124a  and  a67107a );
 a36a <=( a67092a  and  a67075a );
 a37a <=( a67060a  and  a67043a );
 a38a <=( a67028a  and  a67011a );
 a39a <=( a66996a  and  a66979a );
 a40a <=( a66964a  and  a66947a );
 a41a <=( a66932a  and  a66915a );
 a42a <=( a66900a  and  a66883a );
 a43a <=( a66868a  and  a66851a );
 a44a <=( a66836a  and  a66819a );
 a45a <=( a66804a  and  a66787a );
 a46a <=( a66772a  and  a66755a );
 a47a <=( a66740a  and  a66723a );
 a48a <=( a66708a  and  a66691a );
 a49a <=( a66676a  and  a66659a );
 a50a <=( a66644a  and  a66627a );
 a51a <=( a66612a  and  a66595a );
 a52a <=( a66580a  and  a66563a );
 a53a <=( a66548a  and  a66531a );
 a54a <=( a66516a  and  a66499a );
 a55a <=( a66484a  and  a66467a );
 a56a <=( a66452a  and  a66435a );
 a57a <=( a66420a  and  a66403a );
 a58a <=( a66388a  and  a66371a );
 a59a <=( a66356a  and  a66339a );
 a60a <=( a66324a  and  a66307a );
 a61a <=( a66292a  and  a66275a );
 a62a <=( a66260a  and  a66243a );
 a63a <=( a66228a  and  a66211a );
 a64a <=( a66196a  and  a66179a );
 a65a <=( a66164a  and  a66147a );
 a66a <=( a66132a  and  a66115a );
 a67a <=( a66100a  and  a66083a );
 a68a <=( a66068a  and  a66051a );
 a69a <=( a66036a  and  a66019a );
 a70a <=( a66004a  and  a65987a );
 a71a <=( a65972a  and  a65955a );
 a72a <=( a65940a  and  a65923a );
 a73a <=( a65908a  and  a65891a );
 a74a <=( a65876a  and  a65859a );
 a75a <=( a65844a  and  a65827a );
 a76a <=( a65812a  and  a65795a );
 a77a <=( a65780a  and  a65763a );
 a78a <=( a65748a  and  a65731a );
 a79a <=( a65716a  and  a65699a );
 a80a <=( a65684a  and  a65667a );
 a81a <=( a65652a  and  a65635a );
 a82a <=( a65620a  and  a65603a );
 a83a <=( a65588a  and  a65571a );
 a84a <=( a65556a  and  a65539a );
 a85a <=( a65524a  and  a65507a );
 a86a <=( a65492a  and  a65475a );
 a87a <=( a65460a  and  a65443a );
 a88a <=( a65428a  and  a65411a );
 a89a <=( a65396a  and  a65379a );
 a90a <=( a65364a  and  a65347a );
 a91a <=( a65332a  and  a65315a );
 a92a <=( a65300a  and  a65283a );
 a93a <=( a65268a  and  a65251a );
 a94a <=( a65236a  and  a65219a );
 a95a <=( a65204a  and  a65187a );
 a96a <=( a65172a  and  a65155a );
 a97a <=( a65140a  and  a65123a );
 a98a <=( a65108a  and  a65091a );
 a99a <=( a65076a  and  a65059a );
 a100a <=( a65044a  and  a65027a );
 a101a <=( a65012a  and  a64995a );
 a102a <=( a64980a  and  a64963a );
 a103a <=( a64948a  and  a64931a );
 a104a <=( a64916a  and  a64899a );
 a105a <=( a64884a  and  a64867a );
 a106a <=( a64852a  and  a64835a );
 a107a <=( a64820a  and  a64803a );
 a108a <=( a64788a  and  a64771a );
 a109a <=( a64756a  and  a64739a );
 a110a <=( a64724a  and  a64707a );
 a111a <=( a64692a  and  a64675a );
 a112a <=( a64660a  and  a64643a );
 a113a <=( a64628a  and  a64611a );
 a114a <=( a64596a  and  a64579a );
 a115a <=( a64564a  and  a64547a );
 a116a <=( a64532a  and  a64515a );
 a117a <=( a64500a  and  a64483a );
 a118a <=( a64468a  and  a64451a );
 a119a <=( a64436a  and  a64419a );
 a120a <=( a64404a  and  a64387a );
 a121a <=( a64372a  and  a64355a );
 a122a <=( a64340a  and  a64323a );
 a123a <=( a64308a  and  a64291a );
 a124a <=( a64276a  and  a64259a );
 a125a <=( a64244a  and  a64227a );
 a126a <=( a64212a  and  a64195a );
 a127a <=( a64180a  and  a64163a );
 a128a <=( a64148a  and  a64131a );
 a129a <=( a64116a  and  a64099a );
 a130a <=( a64084a  and  a64067a );
 a131a <=( a64052a  and  a64035a );
 a132a <=( a64020a  and  a64003a );
 a133a <=( a63988a  and  a63971a );
 a134a <=( a63956a  and  a63939a );
 a135a <=( a63924a  and  a63907a );
 a136a <=( a63892a  and  a63875a );
 a137a <=( a63860a  and  a63843a );
 a138a <=( a63828a  and  a63811a );
 a139a <=( a63796a  and  a63779a );
 a140a <=( a63764a  and  a63747a );
 a141a <=( a63732a  and  a63715a );
 a142a <=( a63700a  and  a63683a );
 a143a <=( a63668a  and  a63651a );
 a144a <=( a63636a  and  a63619a );
 a145a <=( a63604a  and  a63587a );
 a146a <=( a63572a  and  a63555a );
 a147a <=( a63540a  and  a63523a );
 a148a <=( a63508a  and  a63491a );
 a149a <=( a63476a  and  a63459a );
 a150a <=( a63444a  and  a63427a );
 a151a <=( a63412a  and  a63395a );
 a152a <=( a63380a  and  a63363a );
 a153a <=( a63348a  and  a63331a );
 a154a <=( a63316a  and  a63299a );
 a155a <=( a63284a  and  a63267a );
 a156a <=( a63252a  and  a63235a );
 a157a <=( a63220a  and  a63203a );
 a158a <=( a63188a  and  a63171a );
 a159a <=( a63156a  and  a63139a );
 a160a <=( a63124a  and  a63107a );
 a161a <=( a63092a  and  a63075a );
 a162a <=( a63060a  and  a63043a );
 a163a <=( a63028a  and  a63011a );
 a164a <=( a62996a  and  a62979a );
 a165a <=( a62964a  and  a62947a );
 a166a <=( a62932a  and  a62915a );
 a167a <=( a62900a  and  a62883a );
 a168a <=( a62868a  and  a62851a );
 a169a <=( a62836a  and  a62819a );
 a170a <=( a62804a  and  a62787a );
 a171a <=( a62772a  and  a62755a );
 a172a <=( a62740a  and  a62723a );
 a173a <=( a62708a  and  a62691a );
 a174a <=( a62676a  and  a62659a );
 a175a <=( a62644a  and  a62627a );
 a176a <=( a62612a  and  a62595a );
 a177a <=( a62580a  and  a62565a );
 a178a <=( a62550a  and  a62535a );
 a179a <=( a62520a  and  a62505a );
 a180a <=( a62490a  and  a62475a );
 a181a <=( a62460a  and  a62445a );
 a182a <=( a62430a  and  a62415a );
 a183a <=( a62400a  and  a62385a );
 a184a <=( a62370a  and  a62355a );
 a185a <=( a62340a  and  a62325a );
 a186a <=( a62310a  and  a62295a );
 a187a <=( a62280a  and  a62265a );
 a188a <=( a62250a  and  a62235a );
 a189a <=( a62220a  and  a62205a );
 a190a <=( a62190a  and  a62175a );
 a191a <=( a62160a  and  a62145a );
 a192a <=( a62130a  and  a62115a );
 a193a <=( a62100a  and  a62085a );
 a194a <=( a62070a  and  a62055a );
 a195a <=( a62040a  and  a62025a );
 a196a <=( a62010a  and  a61995a );
 a197a <=( a61980a  and  a61965a );
 a198a <=( a61950a  and  a61935a );
 a199a <=( a61920a  and  a61905a );
 a200a <=( a61890a  and  a61875a );
 a201a <=( a61860a  and  a61845a );
 a202a <=( a61830a  and  a61815a );
 a203a <=( a61800a  and  a61785a );
 a204a <=( a61770a  and  a61755a );
 a205a <=( a61740a  and  a61725a );
 a206a <=( a61710a  and  a61695a );
 a207a <=( a61680a  and  a61665a );
 a208a <=( a61650a  and  a61635a );
 a209a <=( a61620a  and  a61605a );
 a210a <=( a61590a  and  a61575a );
 a211a <=( a61560a  and  a61545a );
 a212a <=( a61530a  and  a61515a );
 a213a <=( a61500a  and  a61485a );
 a214a <=( a61470a  and  a61455a );
 a215a <=( a61440a  and  a61425a );
 a216a <=( a61410a  and  a61395a );
 a217a <=( a61380a  and  a61365a );
 a218a <=( a61350a  and  a61335a );
 a219a <=( a61320a  and  a61305a );
 a220a <=( a61290a  and  a61275a );
 a221a <=( a61260a  and  a61245a );
 a222a <=( a61230a  and  a61215a );
 a223a <=( a61200a  and  a61185a );
 a224a <=( a61170a  and  a61155a );
 a225a <=( a61140a  and  a61125a );
 a226a <=( a61110a  and  a61095a );
 a227a <=( a61080a  and  a61065a );
 a228a <=( a61050a  and  a61035a );
 a229a <=( a61020a  and  a61005a );
 a230a <=( a60990a  and  a60975a );
 a231a <=( a60960a  and  a60945a );
 a232a <=( a60930a  and  a60915a );
 a233a <=( a60900a  and  a60885a );
 a234a <=( a60870a  and  a60855a );
 a235a <=( a60840a  and  a60825a );
 a236a <=( a60810a  and  a60795a );
 a237a <=( a60780a  and  a60765a );
 a238a <=( a60750a  and  a60735a );
 a239a <=( a60720a  and  a60705a );
 a240a <=( a60690a  and  a60675a );
 a241a <=( a60660a  and  a60645a );
 a242a <=( a60630a  and  a60615a );
 a243a <=( a60600a  and  a60585a );
 a244a <=( a60570a  and  a60555a );
 a245a <=( a60540a  and  a60525a );
 a246a <=( a60510a  and  a60495a );
 a247a <=( a60480a  and  a60465a );
 a248a <=( a60450a  and  a60435a );
 a249a <=( a60420a  and  a60405a );
 a250a <=( a60390a  and  a60375a );
 a251a <=( a60360a  and  a60345a );
 a252a <=( a60330a  and  a60315a );
 a253a <=( a60300a  and  a60285a );
 a254a <=( a60270a  and  a60255a );
 a255a <=( a60240a  and  a60225a );
 a256a <=( a60210a  and  a60195a );
 a257a <=( a60180a  and  a60165a );
 a258a <=( a60150a  and  a60135a );
 a259a <=( a60120a  and  a60105a );
 a260a <=( a60090a  and  a60075a );
 a261a <=( a60060a  and  a60045a );
 a262a <=( a60030a  and  a60015a );
 a263a <=( a60000a  and  a59985a );
 a264a <=( a59970a  and  a59955a );
 a265a <=( a59940a  and  a59925a );
 a266a <=( a59910a  and  a59895a );
 a267a <=( a59880a  and  a59865a );
 a268a <=( a59850a  and  a59835a );
 a269a <=( a59820a  and  a59805a );
 a270a <=( a59790a  and  a59775a );
 a271a <=( a59760a  and  a59745a );
 a272a <=( a59730a  and  a59715a );
 a273a <=( a59700a  and  a59685a );
 a274a <=( a59670a  and  a59655a );
 a275a <=( a59640a  and  a59625a );
 a276a <=( a59610a  and  a59595a );
 a277a <=( a59580a  and  a59565a );
 a278a <=( a59550a  and  a59535a );
 a279a <=( a59520a  and  a59505a );
 a280a <=( a59490a  and  a59475a );
 a281a <=( a59460a  and  a59445a );
 a282a <=( a59430a  and  a59415a );
 a283a <=( a59400a  and  a59385a );
 a284a <=( a59370a  and  a59355a );
 a285a <=( a59340a  and  a59325a );
 a286a <=( a59310a  and  a59295a );
 a287a <=( a59280a  and  a59265a );
 a288a <=( a59250a  and  a59235a );
 a289a <=( a59220a  and  a59205a );
 a290a <=( a59190a  and  a59175a );
 a291a <=( a59160a  and  a59145a );
 a292a <=( a59130a  and  a59115a );
 a293a <=( a59100a  and  a59085a );
 a294a <=( a59070a  and  a59055a );
 a295a <=( a59040a  and  a59025a );
 a296a <=( a59010a  and  a58995a );
 a297a <=( a58980a  and  a58965a );
 a298a <=( a58950a  and  a58935a );
 a299a <=( a58920a  and  a58905a );
 a300a <=( a58890a  and  a58875a );
 a301a <=( a58860a  and  a58845a );
 a302a <=( a58830a  and  a58815a );
 a303a <=( a58800a  and  a58785a );
 a304a <=( a58770a  and  a58755a );
 a305a <=( a58740a  and  a58725a );
 a306a <=( a58710a  and  a58695a );
 a307a <=( a58680a  and  a58665a );
 a308a <=( a58650a  and  a58635a );
 a309a <=( a58620a  and  a58605a );
 a310a <=( a58590a  and  a58575a );
 a311a <=( a58560a  and  a58545a );
 a312a <=( a58530a  and  a58515a );
 a313a <=( a58500a  and  a58485a );
 a314a <=( a58470a  and  a58455a );
 a315a <=( a58440a  and  a58425a );
 a316a <=( a58410a  and  a58395a );
 a317a <=( a58380a  and  a58365a );
 a318a <=( a58350a  and  a58335a );
 a319a <=( a58320a  and  a58305a );
 a320a <=( a58290a  and  a58275a );
 a321a <=( a58260a  and  a58245a );
 a322a <=( a58230a  and  a58215a );
 a323a <=( a58200a  and  a58185a );
 a324a <=( a58170a  and  a58155a );
 a325a <=( a58140a  and  a58125a );
 a326a <=( a58110a  and  a58095a );
 a327a <=( a58080a  and  a58065a );
 a328a <=( a58050a  and  a58035a );
 a329a <=( a58020a  and  a58005a );
 a330a <=( a57990a  and  a57975a );
 a331a <=( a57960a  and  a57945a );
 a332a <=( a57930a  and  a57915a );
 a333a <=( a57900a  and  a57885a );
 a334a <=( a57870a  and  a57855a );
 a335a <=( a57840a  and  a57825a );
 a336a <=( a57810a  and  a57795a );
 a337a <=( a57780a  and  a57765a );
 a338a <=( a57750a  and  a57735a );
 a339a <=( a57720a  and  a57705a );
 a340a <=( a57690a  and  a57675a );
 a341a <=( a57660a  and  a57645a );
 a342a <=( a57630a  and  a57615a );
 a343a <=( a57600a  and  a57585a );
 a344a <=( a57570a  and  a57555a );
 a345a <=( a57540a  and  a57525a );
 a346a <=( a57510a  and  a57495a );
 a347a <=( a57480a  and  a57465a );
 a348a <=( a57450a  and  a57435a );
 a349a <=( a57420a  and  a57405a );
 a350a <=( a57390a  and  a57375a );
 a351a <=( a57360a  and  a57345a );
 a352a <=( a57330a  and  a57315a );
 a353a <=( a57300a  and  a57285a );
 a354a <=( a57270a  and  a57255a );
 a355a <=( a57240a  and  a57225a );
 a356a <=( a57210a  and  a57195a );
 a357a <=( a57180a  and  a57165a );
 a358a <=( a57150a  and  a57135a );
 a359a <=( a57120a  and  a57105a );
 a360a <=( a57090a  and  a57075a );
 a361a <=( a57060a  and  a57045a );
 a362a <=( a57030a  and  a57015a );
 a363a <=( a57000a  and  a56985a );
 a364a <=( a56970a  and  a56955a );
 a365a <=( a56940a  and  a56925a );
 a366a <=( a56910a  and  a56895a );
 a367a <=( a56880a  and  a56865a );
 a368a <=( a56850a  and  a56835a );
 a369a <=( a56820a  and  a56805a );
 a370a <=( a56790a  and  a56775a );
 a371a <=( a56760a  and  a56745a );
 a372a <=( a56730a  and  a56715a );
 a373a <=( a56700a  and  a56685a );
 a374a <=( a56670a  and  a56655a );
 a375a <=( a56640a  and  a56625a );
 a376a <=( a56610a  and  a56595a );
 a377a <=( a56580a  and  a56565a );
 a378a <=( a56550a  and  a56535a );
 a379a <=( a56520a  and  a56505a );
 a380a <=( a56490a  and  a56475a );
 a381a <=( a56460a  and  a56445a );
 a382a <=( a56430a  and  a56415a );
 a383a <=( a56400a  and  a56385a );
 a384a <=( a56370a  and  a56355a );
 a385a <=( a56340a  and  a56325a );
 a386a <=( a56310a  and  a56295a );
 a387a <=( a56280a  and  a56265a );
 a388a <=( a56250a  and  a56235a );
 a389a <=( a56220a  and  a56205a );
 a390a <=( a56190a  and  a56175a );
 a391a <=( a56160a  and  a56145a );
 a392a <=( a56130a  and  a56115a );
 a393a <=( a56100a  and  a56085a );
 a394a <=( a56070a  and  a56055a );
 a395a <=( a56040a  and  a56025a );
 a396a <=( a56010a  and  a55995a );
 a397a <=( a55980a  and  a55965a );
 a398a <=( a55950a  and  a55935a );
 a399a <=( a55920a  and  a55905a );
 a400a <=( a55890a  and  a55875a );
 a401a <=( a55860a  and  a55845a );
 a402a <=( a55830a  and  a55815a );
 a403a <=( a55800a  and  a55785a );
 a404a <=( a55770a  and  a55755a );
 a405a <=( a55740a  and  a55725a );
 a406a <=( a55710a  and  a55695a );
 a407a <=( a55680a  and  a55665a );
 a408a <=( a55650a  and  a55635a );
 a409a <=( a55620a  and  a55605a );
 a410a <=( a55590a  and  a55575a );
 a411a <=( a55560a  and  a55545a );
 a412a <=( a55530a  and  a55515a );
 a413a <=( a55500a  and  a55485a );
 a414a <=( a55470a  and  a55455a );
 a415a <=( a55440a  and  a55425a );
 a416a <=( a55410a  and  a55395a );
 a417a <=( a55380a  and  a55365a );
 a418a <=( a55350a  and  a55335a );
 a419a <=( a55320a  and  a55305a );
 a420a <=( a55290a  and  a55275a );
 a421a <=( a55260a  and  a55245a );
 a422a <=( a55230a  and  a55215a );
 a423a <=( a55200a  and  a55185a );
 a424a <=( a55170a  and  a55155a );
 a425a <=( a55140a  and  a55125a );
 a426a <=( a55110a  and  a55095a );
 a427a <=( a55080a  and  a55065a );
 a428a <=( a55050a  and  a55035a );
 a429a <=( a55020a  and  a55005a );
 a430a <=( a54990a  and  a54975a );
 a431a <=( a54960a  and  a54945a );
 a432a <=( a54930a  and  a54915a );
 a433a <=( a54900a  and  a54885a );
 a434a <=( a54870a  and  a54855a );
 a435a <=( a54840a  and  a54825a );
 a436a <=( a54810a  and  a54795a );
 a437a <=( a54780a  and  a54765a );
 a438a <=( a54750a  and  a54735a );
 a439a <=( a54720a  and  a54705a );
 a440a <=( a54690a  and  a54675a );
 a441a <=( a54660a  and  a54645a );
 a442a <=( a54630a  and  a54615a );
 a443a <=( a54600a  and  a54585a );
 a444a <=( a54570a  and  a54555a );
 a445a <=( a54540a  and  a54525a );
 a446a <=( a54510a  and  a54495a );
 a447a <=( a54480a  and  a54465a );
 a448a <=( a54450a  and  a54435a );
 a449a <=( a54420a  and  a54405a );
 a450a <=( a54390a  and  a54375a );
 a451a <=( a54360a  and  a54345a );
 a452a <=( a54330a  and  a54315a );
 a453a <=( a54300a  and  a54285a );
 a454a <=( a54270a  and  a54255a );
 a455a <=( a54240a  and  a54225a );
 a456a <=( a54210a  and  a54195a );
 a457a <=( a54180a  and  a54165a );
 a458a <=( a54150a  and  a54135a );
 a459a <=( a54120a  and  a54105a );
 a460a <=( a54090a  and  a54075a );
 a461a <=( a54060a  and  a54045a );
 a462a <=( a54030a  and  a54015a );
 a463a <=( a54000a  and  a53985a );
 a464a <=( a53970a  and  a53955a );
 a465a <=( a53940a  and  a53925a );
 a466a <=( a53910a  and  a53895a );
 a467a <=( a53880a  and  a53865a );
 a468a <=( a53850a  and  a53835a );
 a469a <=( a53820a  and  a53805a );
 a470a <=( a53790a  and  a53775a );
 a471a <=( a53760a  and  a53745a );
 a472a <=( a53730a  and  a53715a );
 a473a <=( a53700a  and  a53685a );
 a474a <=( a53670a  and  a53655a );
 a475a <=( a53640a  and  a53625a );
 a476a <=( a53610a  and  a53595a );
 a477a <=( a53580a  and  a53565a );
 a478a <=( a53550a  and  a53535a );
 a479a <=( a53520a  and  a53505a );
 a480a <=( a53490a  and  a53475a );
 a481a <=( a53460a  and  a53445a );
 a482a <=( a53430a  and  a53415a );
 a483a <=( a53400a  and  a53385a );
 a484a <=( a53370a  and  a53355a );
 a485a <=( a53340a  and  a53325a );
 a486a <=( a53310a  and  a53295a );
 a487a <=( a53280a  and  a53265a );
 a488a <=( a53250a  and  a53235a );
 a489a <=( a53220a  and  a53205a );
 a490a <=( a53190a  and  a53175a );
 a491a <=( a53160a  and  a53145a );
 a492a <=( a53130a  and  a53115a );
 a493a <=( a53100a  and  a53085a );
 a494a <=( a53070a  and  a53055a );
 a495a <=( a53040a  and  a53025a );
 a496a <=( a53010a  and  a52995a );
 a497a <=( a52980a  and  a52965a );
 a498a <=( a52950a  and  a52935a );
 a499a <=( a52920a  and  a52905a );
 a500a <=( a52890a  and  a52875a );
 a501a <=( a52860a  and  a52845a );
 a502a <=( a52830a  and  a52815a );
 a503a <=( a52800a  and  a52785a );
 a504a <=( a52770a  and  a52755a );
 a505a <=( a52740a  and  a52725a );
 a506a <=( a52710a  and  a52695a );
 a507a <=( a52680a  and  a52665a );
 a508a <=( a52650a  and  a52635a );
 a509a <=( a52620a  and  a52605a );
 a510a <=( a52590a  and  a52575a );
 a511a <=( a52560a  and  a52545a );
 a512a <=( a52530a  and  a52515a );
 a513a <=( a52500a  and  a52485a );
 a514a <=( a52470a  and  a52455a );
 a515a <=( a52440a  and  a52425a );
 a516a <=( a52410a  and  a52395a );
 a517a <=( a52380a  and  a52365a );
 a518a <=( a52350a  and  a52335a );
 a519a <=( a52320a  and  a52305a );
 a520a <=( a52290a  and  a52275a );
 a521a <=( a52260a  and  a52245a );
 a522a <=( a52230a  and  a52215a );
 a523a <=( a52200a  and  a52185a );
 a524a <=( a52170a  and  a52155a );
 a525a <=( a52140a  and  a52125a );
 a526a <=( a52110a  and  a52095a );
 a527a <=( a52080a  and  a52065a );
 a528a <=( a52050a  and  a52035a );
 a529a <=( a52020a  and  a52005a );
 a530a <=( a51990a  and  a51975a );
 a531a <=( a51960a  and  a51945a );
 a532a <=( a51930a  and  a51915a );
 a533a <=( a51900a  and  a51885a );
 a534a <=( a51870a  and  a51855a );
 a535a <=( a51840a  and  a51825a );
 a536a <=( a51810a  and  a51795a );
 a537a <=( a51780a  and  a51765a );
 a538a <=( a51750a  and  a51735a );
 a539a <=( a51720a  and  a51705a );
 a540a <=( a51690a  and  a51675a );
 a541a <=( a51660a  and  a51645a );
 a542a <=( a51630a  and  a51615a );
 a543a <=( a51600a  and  a51585a );
 a544a <=( a51570a  and  a51555a );
 a545a <=( a51540a  and  a51525a );
 a546a <=( a51510a  and  a51495a );
 a547a <=( a51480a  and  a51465a );
 a548a <=( a51450a  and  a51435a );
 a549a <=( a51420a  and  a51405a );
 a550a <=( a51390a  and  a51375a );
 a551a <=( a51360a  and  a51345a );
 a552a <=( a51330a  and  a51315a );
 a553a <=( a51300a  and  a51285a );
 a554a <=( a51270a  and  a51255a );
 a555a <=( a51240a  and  a51225a );
 a556a <=( a51210a  and  a51195a );
 a557a <=( a51180a  and  a51165a );
 a558a <=( a51150a  and  a51135a );
 a559a <=( a51120a  and  a51105a );
 a560a <=( a51090a  and  a51075a );
 a561a <=( a51060a  and  a51045a );
 a562a <=( a51030a  and  a51015a );
 a563a <=( a51000a  and  a50985a );
 a564a <=( a50970a  and  a50955a );
 a565a <=( a50940a  and  a50925a );
 a566a <=( a50910a  and  a50895a );
 a567a <=( a50880a  and  a50865a );
 a568a <=( a50850a  and  a50835a );
 a569a <=( a50820a  and  a50805a );
 a570a <=( a50790a  and  a50775a );
 a571a <=( a50760a  and  a50745a );
 a572a <=( a50730a  and  a50715a );
 a573a <=( a50700a  and  a50685a );
 a574a <=( a50670a  and  a50655a );
 a575a <=( a50640a  and  a50625a );
 a576a <=( a50610a  and  a50595a );
 a577a <=( a50580a  and  a50565a );
 a578a <=( a50550a  and  a50535a );
 a579a <=( a50520a  and  a50505a );
 a580a <=( a50490a  and  a50475a );
 a581a <=( a50460a  and  a50445a );
 a582a <=( a50430a  and  a50415a );
 a583a <=( a50400a  and  a50385a );
 a584a <=( a50370a  and  a50355a );
 a585a <=( a50340a  and  a50325a );
 a586a <=( a50310a  and  a50295a );
 a587a <=( a50280a  and  a50265a );
 a588a <=( a50250a  and  a50235a );
 a589a <=( a50220a  and  a50205a );
 a590a <=( a50190a  and  a50175a );
 a591a <=( a50160a  and  a50145a );
 a592a <=( a50130a  and  a50115a );
 a593a <=( a50100a  and  a50085a );
 a594a <=( a50070a  and  a50055a );
 a595a <=( a50040a  and  a50025a );
 a596a <=( a50010a  and  a49995a );
 a597a <=( a49980a  and  a49965a );
 a598a <=( a49950a  and  a49935a );
 a599a <=( a49920a  and  a49905a );
 a600a <=( a49890a  and  a49875a );
 a601a <=( a49860a  and  a49845a );
 a602a <=( a49830a  and  a49815a );
 a603a <=( a49800a  and  a49785a );
 a604a <=( a49770a  and  a49755a );
 a605a <=( a49740a  and  a49725a );
 a606a <=( a49710a  and  a49695a );
 a607a <=( a49680a  and  a49665a );
 a608a <=( a49650a  and  a49635a );
 a609a <=( a49620a  and  a49605a );
 a610a <=( a49590a  and  a49575a );
 a611a <=( a49560a  and  a49545a );
 a612a <=( a49530a  and  a49515a );
 a613a <=( a49500a  and  a49485a );
 a614a <=( a49470a  and  a49455a );
 a615a <=( a49440a  and  a49425a );
 a616a <=( a49410a  and  a49395a );
 a617a <=( a49380a  and  a49365a );
 a618a <=( a49350a  and  a49335a );
 a619a <=( a49320a  and  a49305a );
 a620a <=( a49290a  and  a49275a );
 a621a <=( a49260a  and  a49245a );
 a622a <=( a49230a  and  a49215a );
 a623a <=( a49200a  and  a49185a );
 a624a <=( a49170a  and  a49155a );
 a625a <=( a49140a  and  a49125a );
 a626a <=( a49110a  and  a49095a );
 a627a <=( a49080a  and  a49065a );
 a628a <=( a49050a  and  a49035a );
 a629a <=( a49020a  and  a49005a );
 a630a <=( a48990a  and  a48975a );
 a631a <=( a48960a  and  a48945a );
 a632a <=( a48930a  and  a48915a );
 a633a <=( a48900a  and  a48885a );
 a634a <=( a48870a  and  a48855a );
 a635a <=( a48840a  and  a48825a );
 a636a <=( a48810a  and  a48795a );
 a637a <=( a48780a  and  a48765a );
 a638a <=( a48750a  and  a48735a );
 a639a <=( a48720a  and  a48705a );
 a640a <=( a48690a  and  a48675a );
 a641a <=( a48660a  and  a48645a );
 a642a <=( a48630a  and  a48615a );
 a643a <=( a48600a  and  a48585a );
 a644a <=( a48570a  and  a48555a );
 a645a <=( a48540a  and  a48525a );
 a646a <=( a48510a  and  a48495a );
 a647a <=( a48480a  and  a48465a );
 a648a <=( a48450a  and  a48435a );
 a649a <=( a48420a  and  a48405a );
 a650a <=( a48390a  and  a48375a );
 a651a <=( a48360a  and  a48345a );
 a652a <=( a48330a  and  a48315a );
 a653a <=( a48300a  and  a48285a );
 a654a <=( a48270a  and  a48255a );
 a655a <=( a48240a  and  a48225a );
 a656a <=( a48210a  and  a48195a );
 a657a <=( a48180a  and  a48165a );
 a658a <=( a48150a  and  a48135a );
 a659a <=( a48120a  and  a48105a );
 a660a <=( a48090a  and  a48075a );
 a661a <=( a48060a  and  a48045a );
 a662a <=( a48030a  and  a48015a );
 a663a <=( a48000a  and  a47985a );
 a664a <=( a47970a  and  a47955a );
 a665a <=( a47940a  and  a47925a );
 a666a <=( a47910a  and  a47895a );
 a667a <=( a47880a  and  a47865a );
 a668a <=( a47850a  and  a47835a );
 a669a <=( a47820a  and  a47805a );
 a670a <=( a47790a  and  a47775a );
 a671a <=( a47760a  and  a47745a );
 a672a <=( a47730a  and  a47715a );
 a673a <=( a47700a  and  a47685a );
 a674a <=( a47670a  and  a47655a );
 a675a <=( a47640a  and  a47625a );
 a676a <=( a47610a  and  a47595a );
 a677a <=( a47580a  and  a47565a );
 a678a <=( a47550a  and  a47535a );
 a679a <=( a47520a  and  a47505a );
 a680a <=( a47490a  and  a47475a );
 a681a <=( a47460a  and  a47445a );
 a682a <=( a47430a  and  a47415a );
 a683a <=( a47400a  and  a47385a );
 a684a <=( a47370a  and  a47355a );
 a685a <=( a47340a  and  a47325a );
 a686a <=( a47310a  and  a47295a );
 a687a <=( a47280a  and  a47265a );
 a688a <=( a47250a  and  a47235a );
 a689a <=( a47220a  and  a47205a );
 a690a <=( a47190a  and  a47175a );
 a691a <=( a47160a  and  a47145a );
 a692a <=( a47130a  and  a47115a );
 a693a <=( a47100a  and  a47085a );
 a694a <=( a47070a  and  a47055a );
 a695a <=( a47040a  and  a47025a );
 a696a <=( a47010a  and  a46995a );
 a697a <=( a46980a  and  a46965a );
 a698a <=( a46950a  and  a46935a );
 a699a <=( a46920a  and  a46905a );
 a700a <=( a46890a  and  a46875a );
 a701a <=( a46860a  and  a46845a );
 a702a <=( a46830a  and  a46815a );
 a703a <=( a46800a  and  a46785a );
 a704a <=( a46770a  and  a46755a );
 a705a <=( a46740a  and  a46725a );
 a706a <=( a46710a  and  a46695a );
 a707a <=( a46680a  and  a46665a );
 a708a <=( a46650a  and  a46635a );
 a709a <=( a46620a  and  a46605a );
 a710a <=( a46590a  and  a46575a );
 a711a <=( a46560a  and  a46545a );
 a712a <=( a46530a  and  a46515a );
 a713a <=( a46500a  and  a46485a );
 a714a <=( a46470a  and  a46455a );
 a715a <=( a46440a  and  a46425a );
 a716a <=( a46410a  and  a46395a );
 a717a <=( a46380a  and  a46365a );
 a718a <=( a46350a  and  a46335a );
 a719a <=( a46320a  and  a46305a );
 a720a <=( a46290a  and  a46275a );
 a721a <=( a46260a  and  a46245a );
 a722a <=( a46230a  and  a46215a );
 a723a <=( a46200a  and  a46185a );
 a724a <=( a46170a  and  a46155a );
 a725a <=( a46140a  and  a46125a );
 a726a <=( a46110a  and  a46095a );
 a727a <=( a46080a  and  a46065a );
 a728a <=( a46050a  and  a46035a );
 a729a <=( a46020a  and  a46005a );
 a730a <=( a45990a  and  a45975a );
 a731a <=( a45960a  and  a45945a );
 a732a <=( a45930a  and  a45915a );
 a733a <=( a45900a  and  a45885a );
 a734a <=( a45870a  and  a45855a );
 a735a <=( a45840a  and  a45825a );
 a736a <=( a45810a  and  a45795a );
 a737a <=( a45780a  and  a45765a );
 a738a <=( a45750a  and  a45735a );
 a739a <=( a45720a  and  a45705a );
 a740a <=( a45690a  and  a45675a );
 a741a <=( a45660a  and  a45645a );
 a742a <=( a45630a  and  a45615a );
 a743a <=( a45600a  and  a45585a );
 a744a <=( a45570a  and  a45555a );
 a745a <=( a45540a  and  a45525a );
 a746a <=( a45510a  and  a45495a );
 a747a <=( a45480a  and  a45465a );
 a748a <=( a45450a  and  a45435a );
 a749a <=( a45420a  and  a45405a );
 a750a <=( a45390a  and  a45375a );
 a751a <=( a45360a  and  a45345a );
 a752a <=( a45330a  and  a45315a );
 a753a <=( a45300a  and  a45285a );
 a754a <=( a45272a  and  a45257a );
 a755a <=( a45244a  and  a45229a );
 a756a <=( a45216a  and  a45201a );
 a757a <=( a45188a  and  a45173a );
 a758a <=( a45160a  and  a45145a );
 a759a <=( a45132a  and  a45117a );
 a760a <=( a45104a  and  a45089a );
 a761a <=( a45076a  and  a45061a );
 a762a <=( a45048a  and  a45033a );
 a763a <=( a45020a  and  a45005a );
 a764a <=( a44992a  and  a44977a );
 a765a <=( a44964a  and  a44949a );
 a766a <=( a44936a  and  a44921a );
 a767a <=( a44908a  and  a44893a );
 a768a <=( a44880a  and  a44865a );
 a769a <=( a44852a  and  a44837a );
 a770a <=( a44824a  and  a44809a );
 a771a <=( a44796a  and  a44781a );
 a772a <=( a44768a  and  a44753a );
 a773a <=( a44740a  and  a44725a );
 a774a <=( a44712a  and  a44697a );
 a775a <=( a44684a  and  a44669a );
 a776a <=( a44656a  and  a44641a );
 a777a <=( a44628a  and  a44613a );
 a778a <=( a44600a  and  a44585a );
 a779a <=( a44572a  and  a44557a );
 a780a <=( a44544a  and  a44529a );
 a781a <=( a44516a  and  a44501a );
 a782a <=( a44488a  and  a44473a );
 a783a <=( a44460a  and  a44445a );
 a784a <=( a44432a  and  a44417a );
 a785a <=( a44404a  and  a44389a );
 a786a <=( a44376a  and  a44361a );
 a787a <=( a44348a  and  a44333a );
 a788a <=( a44320a  and  a44305a );
 a789a <=( a44292a  and  a44277a );
 a790a <=( a44264a  and  a44249a );
 a791a <=( a44236a  and  a44221a );
 a792a <=( a44208a  and  a44193a );
 a793a <=( a44180a  and  a44165a );
 a794a <=( a44152a  and  a44137a );
 a795a <=( a44124a  and  a44109a );
 a796a <=( a44096a  and  a44081a );
 a797a <=( a44068a  and  a44053a );
 a798a <=( a44040a  and  a44025a );
 a799a <=( a44012a  and  a43997a );
 a800a <=( a43984a  and  a43969a );
 a801a <=( a43956a  and  a43941a );
 a802a <=( a43928a  and  a43913a );
 a803a <=( a43900a  and  a43885a );
 a804a <=( a43872a  and  a43857a );
 a805a <=( a43844a  and  a43829a );
 a806a <=( a43816a  and  a43801a );
 a807a <=( a43788a  and  a43773a );
 a808a <=( a43760a  and  a43745a );
 a809a <=( a43732a  and  a43717a );
 a810a <=( a43704a  and  a43689a );
 a811a <=( a43676a  and  a43661a );
 a812a <=( a43648a  and  a43633a );
 a813a <=( a43620a  and  a43605a );
 a814a <=( a43592a  and  a43577a );
 a815a <=( a43564a  and  a43549a );
 a816a <=( a43536a  and  a43521a );
 a817a <=( a43508a  and  a43493a );
 a818a <=( a43480a  and  a43465a );
 a819a <=( a43452a  and  a43437a );
 a820a <=( a43424a  and  a43409a );
 a821a <=( a43396a  and  a43381a );
 a822a <=( a43368a  and  a43353a );
 a823a <=( a43340a  and  a43325a );
 a824a <=( a43312a  and  a43297a );
 a825a <=( a43284a  and  a43269a );
 a826a <=( a43256a  and  a43241a );
 a827a <=( a43228a  and  a43213a );
 a828a <=( a43200a  and  a43185a );
 a829a <=( a43172a  and  a43157a );
 a830a <=( a43144a  and  a43129a );
 a831a <=( a43116a  and  a43101a );
 a832a <=( a43088a  and  a43073a );
 a833a <=( a43060a  and  a43045a );
 a834a <=( a43032a  and  a43017a );
 a835a <=( a43004a  and  a42989a );
 a836a <=( a42976a  and  a42961a );
 a837a <=( a42948a  and  a42933a );
 a838a <=( a42920a  and  a42905a );
 a839a <=( a42892a  and  a42877a );
 a840a <=( a42864a  and  a42849a );
 a841a <=( a42836a  and  a42821a );
 a842a <=( a42808a  and  a42793a );
 a843a <=( a42780a  and  a42765a );
 a844a <=( a42752a  and  a42737a );
 a845a <=( a42724a  and  a42709a );
 a846a <=( a42696a  and  a42681a );
 a847a <=( a42668a  and  a42653a );
 a848a <=( a42640a  and  a42625a );
 a849a <=( a42612a  and  a42597a );
 a850a <=( a42584a  and  a42569a );
 a851a <=( a42556a  and  a42541a );
 a852a <=( a42528a  and  a42513a );
 a853a <=( a42500a  and  a42485a );
 a854a <=( a42472a  and  a42457a );
 a855a <=( a42444a  and  a42429a );
 a856a <=( a42416a  and  a42401a );
 a857a <=( a42388a  and  a42373a );
 a858a <=( a42360a  and  a42345a );
 a859a <=( a42332a  and  a42317a );
 a860a <=( a42304a  and  a42289a );
 a861a <=( a42276a  and  a42261a );
 a862a <=( a42248a  and  a42233a );
 a863a <=( a42220a  and  a42205a );
 a864a <=( a42192a  and  a42177a );
 a865a <=( a42164a  and  a42149a );
 a866a <=( a42136a  and  a42121a );
 a867a <=( a42108a  and  a42093a );
 a868a <=( a42080a  and  a42065a );
 a869a <=( a42052a  and  a42037a );
 a870a <=( a42024a  and  a42009a );
 a871a <=( a41996a  and  a41981a );
 a872a <=( a41968a  and  a41953a );
 a873a <=( a41940a  and  a41925a );
 a874a <=( a41912a  and  a41897a );
 a875a <=( a41884a  and  a41869a );
 a876a <=( a41856a  and  a41841a );
 a877a <=( a41828a  and  a41813a );
 a878a <=( a41800a  and  a41785a );
 a879a <=( a41772a  and  a41757a );
 a880a <=( a41744a  and  a41729a );
 a881a <=( a41716a  and  a41701a );
 a882a <=( a41688a  and  a41673a );
 a883a <=( a41660a  and  a41645a );
 a884a <=( a41632a  and  a41617a );
 a885a <=( a41604a  and  a41589a );
 a886a <=( a41576a  and  a41561a );
 a887a <=( a41548a  and  a41533a );
 a888a <=( a41520a  and  a41505a );
 a889a <=( a41492a  and  a41477a );
 a890a <=( a41464a  and  a41449a );
 a891a <=( a41436a  and  a41421a );
 a892a <=( a41408a  and  a41393a );
 a893a <=( a41380a  and  a41365a );
 a894a <=( a41352a  and  a41337a );
 a895a <=( a41324a  and  a41309a );
 a896a <=( a41296a  and  a41281a );
 a897a <=( a41268a  and  a41253a );
 a898a <=( a41240a  and  a41225a );
 a899a <=( a41212a  and  a41197a );
 a900a <=( a41184a  and  a41169a );
 a901a <=( a41156a  and  a41141a );
 a902a <=( a41128a  and  a41113a );
 a903a <=( a41100a  and  a41085a );
 a904a <=( a41072a  and  a41057a );
 a905a <=( a41044a  and  a41029a );
 a906a <=( a41016a  and  a41001a );
 a907a <=( a40988a  and  a40973a );
 a908a <=( a40960a  and  a40945a );
 a909a <=( a40932a  and  a40917a );
 a910a <=( a40904a  and  a40889a );
 a911a <=( a40876a  and  a40861a );
 a912a <=( a40848a  and  a40833a );
 a913a <=( a40820a  and  a40805a );
 a914a <=( a40792a  and  a40777a );
 a915a <=( a40764a  and  a40749a );
 a916a <=( a40736a  and  a40721a );
 a917a <=( a40708a  and  a40693a );
 a918a <=( a40680a  and  a40665a );
 a919a <=( a40652a  and  a40637a );
 a920a <=( a40624a  and  a40609a );
 a921a <=( a40596a  and  a40581a );
 a922a <=( a40568a  and  a40553a );
 a923a <=( a40540a  and  a40525a );
 a924a <=( a40512a  and  a40497a );
 a925a <=( a40484a  and  a40469a );
 a926a <=( a40456a  and  a40441a );
 a927a <=( a40428a  and  a40413a );
 a928a <=( a40400a  and  a40385a );
 a929a <=( a40372a  and  a40357a );
 a930a <=( a40344a  and  a40329a );
 a931a <=( a40316a  and  a40301a );
 a932a <=( a40288a  and  a40273a );
 a933a <=( a40260a  and  a40245a );
 a934a <=( a40232a  and  a40217a );
 a935a <=( a40204a  and  a40189a );
 a936a <=( a40176a  and  a40161a );
 a937a <=( a40148a  and  a40133a );
 a938a <=( a40120a  and  a40105a );
 a939a <=( a40092a  and  a40077a );
 a940a <=( a40064a  and  a40049a );
 a941a <=( a40036a  and  a40021a );
 a942a <=( a40008a  and  a39993a );
 a943a <=( a39980a  and  a39965a );
 a944a <=( a39952a  and  a39937a );
 a945a <=( a39924a  and  a39909a );
 a946a <=( a39896a  and  a39881a );
 a947a <=( a39868a  and  a39853a );
 a948a <=( a39840a  and  a39825a );
 a949a <=( a39812a  and  a39797a );
 a950a <=( a39784a  and  a39769a );
 a951a <=( a39756a  and  a39741a );
 a952a <=( a39728a  and  a39713a );
 a953a <=( a39700a  and  a39685a );
 a954a <=( a39672a  and  a39657a );
 a955a <=( a39644a  and  a39629a );
 a956a <=( a39616a  and  a39601a );
 a957a <=( a39588a  and  a39573a );
 a958a <=( a39560a  and  a39545a );
 a959a <=( a39532a  and  a39517a );
 a960a <=( a39504a  and  a39489a );
 a961a <=( a39476a  and  a39461a );
 a962a <=( a39448a  and  a39433a );
 a963a <=( a39420a  and  a39405a );
 a964a <=( a39392a  and  a39377a );
 a965a <=( a39364a  and  a39349a );
 a966a <=( a39336a  and  a39321a );
 a967a <=( a39308a  and  a39293a );
 a968a <=( a39280a  and  a39265a );
 a969a <=( a39252a  and  a39237a );
 a970a <=( a39224a  and  a39209a );
 a971a <=( a39196a  and  a39181a );
 a972a <=( a39168a  and  a39153a );
 a973a <=( a39140a  and  a39125a );
 a974a <=( a39112a  and  a39097a );
 a975a <=( a39084a  and  a39069a );
 a976a <=( a39056a  and  a39041a );
 a977a <=( a39028a  and  a39013a );
 a978a <=( a39000a  and  a38985a );
 a979a <=( a38972a  and  a38957a );
 a980a <=( a38944a  and  a38929a );
 a981a <=( a38916a  and  a38901a );
 a982a <=( a38888a  and  a38873a );
 a983a <=( a38860a  and  a38845a );
 a984a <=( a38832a  and  a38817a );
 a985a <=( a38804a  and  a38789a );
 a986a <=( a38776a  and  a38761a );
 a987a <=( a38748a  and  a38733a );
 a988a <=( a38720a  and  a38705a );
 a989a <=( a38692a  and  a38677a );
 a990a <=( a38664a  and  a38649a );
 a991a <=( a38636a  and  a38621a );
 a992a <=( a38608a  and  a38593a );
 a993a <=( a38580a  and  a38565a );
 a994a <=( a38552a  and  a38537a );
 a995a <=( a38524a  and  a38509a );
 a996a <=( a38496a  and  a38481a );
 a997a <=( a38468a  and  a38453a );
 a998a <=( a38440a  and  a38425a );
 a999a <=( a38412a  and  a38397a );
 a1000a <=( a38384a  and  a38369a );
 a1001a <=( a38356a  and  a38341a );
 a1002a <=( a38328a  and  a38313a );
 a1003a <=( a38300a  and  a38285a );
 a1004a <=( a38272a  and  a38257a );
 a1005a <=( a38244a  and  a38229a );
 a1006a <=( a38216a  and  a38201a );
 a1007a <=( a38188a  and  a38173a );
 a1008a <=( a38160a  and  a38145a );
 a1009a <=( a38132a  and  a38117a );
 a1010a <=( a38104a  and  a38089a );
 a1011a <=( a38076a  and  a38061a );
 a1012a <=( a38048a  and  a38033a );
 a1013a <=( a38020a  and  a38005a );
 a1014a <=( a37992a  and  a37977a );
 a1015a <=( a37964a  and  a37949a );
 a1016a <=( a37936a  and  a37921a );
 a1017a <=( a37908a  and  a37893a );
 a1018a <=( a37880a  and  a37865a );
 a1019a <=( a37852a  and  a37837a );
 a1020a <=( a37824a  and  a37809a );
 a1021a <=( a37796a  and  a37781a );
 a1022a <=( a37768a  and  a37753a );
 a1023a <=( a37740a  and  a37725a );
 a1024a <=( a37712a  and  a37697a );
 a1025a <=( a37684a  and  a37669a );
 a1026a <=( a37656a  and  a37641a );
 a1027a <=( a37628a  and  a37613a );
 a1028a <=( a37600a  and  a37585a );
 a1029a <=( a37572a  and  a37557a );
 a1030a <=( a37544a  and  a37529a );
 a1031a <=( a37516a  and  a37501a );
 a1032a <=( a37488a  and  a37473a );
 a1033a <=( a37460a  and  a37445a );
 a1034a <=( a37432a  and  a37417a );
 a1035a <=( a37404a  and  a37389a );
 a1036a <=( a37376a  and  a37361a );
 a1037a <=( a37348a  and  a37333a );
 a1038a <=( a37320a  and  a37305a );
 a1039a <=( a37292a  and  a37277a );
 a1040a <=( a37264a  and  a37249a );
 a1041a <=( a37236a  and  a37221a );
 a1042a <=( a37208a  and  a37193a );
 a1043a <=( a37180a  and  a37165a );
 a1044a <=( a37152a  and  a37137a );
 a1045a <=( a37124a  and  a37109a );
 a1046a <=( a37096a  and  a37081a );
 a1047a <=( a37068a  and  a37053a );
 a1048a <=( a37040a  and  a37025a );
 a1049a <=( a37012a  and  a36997a );
 a1050a <=( a36984a  and  a36969a );
 a1051a <=( a36956a  and  a36941a );
 a1052a <=( a36928a  and  a36913a );
 a1053a <=( a36900a  and  a36885a );
 a1054a <=( a36872a  and  a36857a );
 a1055a <=( a36844a  and  a36829a );
 a1056a <=( a36816a  and  a36801a );
 a1057a <=( a36788a  and  a36773a );
 a1058a <=( a36760a  and  a36745a );
 a1059a <=( a36732a  and  a36717a );
 a1060a <=( a36704a  and  a36689a );
 a1061a <=( a36676a  and  a36661a );
 a1062a <=( a36648a  and  a36633a );
 a1063a <=( a36620a  and  a36605a );
 a1064a <=( a36592a  and  a36577a );
 a1065a <=( a36564a  and  a36549a );
 a1066a <=( a36536a  and  a36521a );
 a1067a <=( a36508a  and  a36493a );
 a1068a <=( a36480a  and  a36465a );
 a1069a <=( a36452a  and  a36437a );
 a1070a <=( a36424a  and  a36409a );
 a1071a <=( a36396a  and  a36381a );
 a1072a <=( a36368a  and  a36353a );
 a1073a <=( a36340a  and  a36325a );
 a1074a <=( a36312a  and  a36297a );
 a1075a <=( a36284a  and  a36269a );
 a1076a <=( a36256a  and  a36241a );
 a1077a <=( a36228a  and  a36213a );
 a1078a <=( a36200a  and  a36185a );
 a1079a <=( a36172a  and  a36157a );
 a1080a <=( a36144a  and  a36129a );
 a1081a <=( a36116a  and  a36101a );
 a1082a <=( a36088a  and  a36073a );
 a1083a <=( a36060a  and  a36045a );
 a1084a <=( a36032a  and  a36017a );
 a1085a <=( a36004a  and  a35989a );
 a1086a <=( a35976a  and  a35961a );
 a1087a <=( a35948a  and  a35933a );
 a1088a <=( a35920a  and  a35905a );
 a1089a <=( a35892a  and  a35877a );
 a1090a <=( a35864a  and  a35849a );
 a1091a <=( a35836a  and  a35821a );
 a1092a <=( a35808a  and  a35793a );
 a1093a <=( a35780a  and  a35765a );
 a1094a <=( a35752a  and  a35737a );
 a1095a <=( a35724a  and  a35709a );
 a1096a <=( a35696a  and  a35681a );
 a1097a <=( a35668a  and  a35653a );
 a1098a <=( a35640a  and  a35625a );
 a1099a <=( a35612a  and  a35597a );
 a1100a <=( a35584a  and  a35569a );
 a1101a <=( a35556a  and  a35541a );
 a1102a <=( a35528a  and  a35513a );
 a1103a <=( a35500a  and  a35485a );
 a1104a <=( a35472a  and  a35457a );
 a1105a <=( a35444a  and  a35429a );
 a1106a <=( a35416a  and  a35401a );
 a1107a <=( a35388a  and  a35373a );
 a1108a <=( a35360a  and  a35345a );
 a1109a <=( a35332a  and  a35317a );
 a1110a <=( a35304a  and  a35289a );
 a1111a <=( a35276a  and  a35261a );
 a1112a <=( a35248a  and  a35233a );
 a1113a <=( a35220a  and  a35205a );
 a1114a <=( a35192a  and  a35177a );
 a1115a <=( a35164a  and  a35149a );
 a1116a <=( a35136a  and  a35121a );
 a1117a <=( a35108a  and  a35093a );
 a1118a <=( a35080a  and  a35065a );
 a1119a <=( a35052a  and  a35037a );
 a1120a <=( a35024a  and  a35009a );
 a1121a <=( a34996a  and  a34981a );
 a1122a <=( a34968a  and  a34953a );
 a1123a <=( a34940a  and  a34925a );
 a1124a <=( a34912a  and  a34897a );
 a1125a <=( a34884a  and  a34869a );
 a1126a <=( a34856a  and  a34841a );
 a1127a <=( a34828a  and  a34813a );
 a1128a <=( a34800a  and  a34785a );
 a1129a <=( a34772a  and  a34757a );
 a1130a <=( a34744a  and  a34729a );
 a1131a <=( a34716a  and  a34701a );
 a1132a <=( a34688a  and  a34673a );
 a1133a <=( a34660a  and  a34645a );
 a1134a <=( a34632a  and  a34617a );
 a1135a <=( a34604a  and  a34589a );
 a1136a <=( a34576a  and  a34561a );
 a1137a <=( a34548a  and  a34533a );
 a1138a <=( a34520a  and  a34505a );
 a1139a <=( a34492a  and  a34477a );
 a1140a <=( a34464a  and  a34449a );
 a1141a <=( a34436a  and  a34421a );
 a1142a <=( a34408a  and  a34393a );
 a1143a <=( a34380a  and  a34365a );
 a1144a <=( a34352a  and  a34337a );
 a1145a <=( a34324a  and  a34309a );
 a1146a <=( a34296a  and  a34281a );
 a1147a <=( a34268a  and  a34253a );
 a1148a <=( a34240a  and  a34225a );
 a1149a <=( a34212a  and  a34197a );
 a1150a <=( a34184a  and  a34169a );
 a1151a <=( a34156a  and  a34141a );
 a1152a <=( a34128a  and  a34113a );
 a1153a <=( a34100a  and  a34085a );
 a1154a <=( a34072a  and  a34057a );
 a1155a <=( a34044a  and  a34029a );
 a1156a <=( a34016a  and  a34001a );
 a1157a <=( a33988a  and  a33973a );
 a1158a <=( a33960a  and  a33945a );
 a1159a <=( a33932a  and  a33917a );
 a1160a <=( a33904a  and  a33889a );
 a1161a <=( a33876a  and  a33861a );
 a1162a <=( a33848a  and  a33833a );
 a1163a <=( a33820a  and  a33805a );
 a1164a <=( a33792a  and  a33777a );
 a1165a <=( a33764a  and  a33749a );
 a1166a <=( a33736a  and  a33721a );
 a1167a <=( a33708a  and  a33693a );
 a1168a <=( a33680a  and  a33665a );
 a1169a <=( a33652a  and  a33637a );
 a1170a <=( a33624a  and  a33609a );
 a1171a <=( a33596a  and  a33581a );
 a1172a <=( a33568a  and  a33553a );
 a1173a <=( a33540a  and  a33525a );
 a1174a <=( a33512a  and  a33497a );
 a1175a <=( a33484a  and  a33469a );
 a1176a <=( a33456a  and  a33441a );
 a1177a <=( a33428a  and  a33413a );
 a1178a <=( a33400a  and  a33385a );
 a1179a <=( a33372a  and  a33357a );
 a1180a <=( a33344a  and  a33329a );
 a1181a <=( a33316a  and  a33301a );
 a1182a <=( a33288a  and  a33273a );
 a1183a <=( a33260a  and  a33245a );
 a1184a <=( a33232a  and  a33217a );
 a1185a <=( a33204a  and  a33189a );
 a1186a <=( a33176a  and  a33161a );
 a1187a <=( a33148a  and  a33133a );
 a1188a <=( a33120a  and  a33105a );
 a1189a <=( a33092a  and  a33077a );
 a1190a <=( a33064a  and  a33049a );
 a1191a <=( a33036a  and  a33021a );
 a1192a <=( a33008a  and  a32993a );
 a1193a <=( a32980a  and  a32965a );
 a1194a <=( a32952a  and  a32937a );
 a1195a <=( a32924a  and  a32909a );
 a1196a <=( a32896a  and  a32881a );
 a1197a <=( a32868a  and  a32853a );
 a1198a <=( a32840a  and  a32825a );
 a1199a <=( a32812a  and  a32797a );
 a1200a <=( a32784a  and  a32769a );
 a1201a <=( a32756a  and  a32741a );
 a1202a <=( a32728a  and  a32713a );
 a1203a <=( a32700a  and  a32685a );
 a1204a <=( a32672a  and  a32657a );
 a1205a <=( a32644a  and  a32629a );
 a1206a <=( a32616a  and  a32601a );
 a1207a <=( a32588a  and  a32573a );
 a1208a <=( a32560a  and  a32545a );
 a1209a <=( a32532a  and  a32517a );
 a1210a <=( a32504a  and  a32489a );
 a1211a <=( a32476a  and  a32461a );
 a1212a <=( a32448a  and  a32433a );
 a1213a <=( a32420a  and  a32405a );
 a1214a <=( a32392a  and  a32377a );
 a1215a <=( a32364a  and  a32349a );
 a1216a <=( a32336a  and  a32321a );
 a1217a <=( a32308a  and  a32293a );
 a1218a <=( a32280a  and  a32265a );
 a1219a <=( a32252a  and  a32237a );
 a1220a <=( a32224a  and  a32209a );
 a1221a <=( a32196a  and  a32181a );
 a1222a <=( a32168a  and  a32153a );
 a1223a <=( a32140a  and  a32125a );
 a1224a <=( a32112a  and  a32097a );
 a1225a <=( a32084a  and  a32069a );
 a1226a <=( a32056a  and  a32041a );
 a1227a <=( a32028a  and  a32013a );
 a1228a <=( a32000a  and  a31985a );
 a1229a <=( a31972a  and  a31957a );
 a1230a <=( a31944a  and  a31929a );
 a1231a <=( a31916a  and  a31901a );
 a1232a <=( a31888a  and  a31873a );
 a1233a <=( a31860a  and  a31845a );
 a1234a <=( a31832a  and  a31817a );
 a1235a <=( a31804a  and  a31789a );
 a1236a <=( a31776a  and  a31761a );
 a1237a <=( a31748a  and  a31733a );
 a1238a <=( a31720a  and  a31705a );
 a1239a <=( a31692a  and  a31677a );
 a1240a <=( a31664a  and  a31649a );
 a1241a <=( a31636a  and  a31621a );
 a1242a <=( a31608a  and  a31593a );
 a1243a <=( a31580a  and  a31565a );
 a1244a <=( a31552a  and  a31537a );
 a1245a <=( a31524a  and  a31509a );
 a1246a <=( a31496a  and  a31481a );
 a1247a <=( a31468a  and  a31453a );
 a1248a <=( a31440a  and  a31425a );
 a1249a <=( a31412a  and  a31397a );
 a1250a <=( a31384a  and  a31369a );
 a1251a <=( a31356a  and  a31341a );
 a1252a <=( a31328a  and  a31313a );
 a1253a <=( a31300a  and  a31285a );
 a1254a <=( a31272a  and  a31257a );
 a1255a <=( a31244a  and  a31229a );
 a1256a <=( a31216a  and  a31201a );
 a1257a <=( a31188a  and  a31173a );
 a1258a <=( a31160a  and  a31145a );
 a1259a <=( a31132a  and  a31117a );
 a1260a <=( a31104a  and  a31089a );
 a1261a <=( a31076a  and  a31061a );
 a1262a <=( a31048a  and  a31033a );
 a1263a <=( a31020a  and  a31005a );
 a1264a <=( a30992a  and  a30977a );
 a1265a <=( a30964a  and  a30949a );
 a1266a <=( a30936a  and  a30921a );
 a1267a <=( a30908a  and  a30893a );
 a1268a <=( a30880a  and  a30865a );
 a1269a <=( a30852a  and  a30837a );
 a1270a <=( a30824a  and  a30809a );
 a1271a <=( a30796a  and  a30781a );
 a1272a <=( a30768a  and  a30753a );
 a1273a <=( a30740a  and  a30725a );
 a1274a <=( a30712a  and  a30697a );
 a1275a <=( a30684a  and  a30669a );
 a1276a <=( a30656a  and  a30641a );
 a1277a <=( a30628a  and  a30613a );
 a1278a <=( a30600a  and  a30585a );
 a1279a <=( a30572a  and  a30557a );
 a1280a <=( a30544a  and  a30529a );
 a1281a <=( a30516a  and  a30501a );
 a1282a <=( a30488a  and  a30473a );
 a1283a <=( a30460a  and  a30445a );
 a1284a <=( a30432a  and  a30417a );
 a1285a <=( a30404a  and  a30389a );
 a1286a <=( a30376a  and  a30361a );
 a1287a <=( a30348a  and  a30333a );
 a1288a <=( a30320a  and  a30305a );
 a1289a <=( a30292a  and  a30277a );
 a1290a <=( a30264a  and  a30249a );
 a1291a <=( a30236a  and  a30221a );
 a1292a <=( a30208a  and  a30193a );
 a1293a <=( a30180a  and  a30165a );
 a1294a <=( a30152a  and  a30137a );
 a1295a <=( a30124a  and  a30109a );
 a1296a <=( a30096a  and  a30081a );
 a1297a <=( a30068a  and  a30053a );
 a1298a <=( a30040a  and  a30025a );
 a1299a <=( a30012a  and  a29997a );
 a1300a <=( a29984a  and  a29969a );
 a1301a <=( a29956a  and  a29941a );
 a1302a <=( a29928a  and  a29913a );
 a1303a <=( a29900a  and  a29885a );
 a1304a <=( a29872a  and  a29857a );
 a1305a <=( a29844a  and  a29829a );
 a1306a <=( a29816a  and  a29801a );
 a1307a <=( a29788a  and  a29773a );
 a1308a <=( a29760a  and  a29745a );
 a1309a <=( a29732a  and  a29717a );
 a1310a <=( a29704a  and  a29689a );
 a1311a <=( a29676a  and  a29661a );
 a1312a <=( a29648a  and  a29633a );
 a1313a <=( a29620a  and  a29605a );
 a1314a <=( a29592a  and  a29577a );
 a1315a <=( a29564a  and  a29549a );
 a1316a <=( a29536a  and  a29521a );
 a1317a <=( a29508a  and  a29493a );
 a1318a <=( a29480a  and  a29465a );
 a1319a <=( a29452a  and  a29437a );
 a1320a <=( a29424a  and  a29409a );
 a1321a <=( a29396a  and  a29381a );
 a1322a <=( a29368a  and  a29353a );
 a1323a <=( a29340a  and  a29325a );
 a1324a <=( a29312a  and  a29297a );
 a1325a <=( a29284a  and  a29269a );
 a1326a <=( a29256a  and  a29241a );
 a1327a <=( a29228a  and  a29213a );
 a1328a <=( a29200a  and  a29185a );
 a1329a <=( a29172a  and  a29157a );
 a1330a <=( a29144a  and  a29129a );
 a1331a <=( a29116a  and  a29101a );
 a1332a <=( a29088a  and  a29073a );
 a1333a <=( a29060a  and  a29045a );
 a1334a <=( a29032a  and  a29017a );
 a1335a <=( a29004a  and  a28989a );
 a1336a <=( a28976a  and  a28961a );
 a1337a <=( a28948a  and  a28933a );
 a1338a <=( a28920a  and  a28905a );
 a1339a <=( a28892a  and  a28877a );
 a1340a <=( a28864a  and  a28849a );
 a1341a <=( a28836a  and  a28821a );
 a1342a <=( a28808a  and  a28793a );
 a1343a <=( a28780a  and  a28765a );
 a1344a <=( a28752a  and  a28737a );
 a1345a <=( a28724a  and  a28709a );
 a1346a <=( a28696a  and  a28681a );
 a1347a <=( a28668a  and  a28653a );
 a1348a <=( a28640a  and  a28625a );
 a1349a <=( a28612a  and  a28597a );
 a1350a <=( a28584a  and  a28569a );
 a1351a <=( a28556a  and  a28541a );
 a1352a <=( a28528a  and  a28513a );
 a1353a <=( a28500a  and  a28485a );
 a1354a <=( a28472a  and  a28457a );
 a1355a <=( a28444a  and  a28429a );
 a1356a <=( a28416a  and  a28401a );
 a1357a <=( a28388a  and  a28373a );
 a1358a <=( a28360a  and  a28345a );
 a1359a <=( a28332a  and  a28317a );
 a1360a <=( a28304a  and  a28289a );
 a1361a <=( a28276a  and  a28261a );
 a1362a <=( a28248a  and  a28233a );
 a1363a <=( a28220a  and  a28205a );
 a1364a <=( a28192a  and  a28177a );
 a1365a <=( a28164a  and  a28149a );
 a1366a <=( a28136a  and  a28121a );
 a1367a <=( a28108a  and  a28093a );
 a1368a <=( a28080a  and  a28065a );
 a1369a <=( a28052a  and  a28037a );
 a1370a <=( a28024a  and  a28009a );
 a1371a <=( a27996a  and  a27981a );
 a1372a <=( a27968a  and  a27953a );
 a1373a <=( a27940a  and  a27925a );
 a1374a <=( a27912a  and  a27897a );
 a1375a <=( a27884a  and  a27869a );
 a1376a <=( a27856a  and  a27841a );
 a1377a <=( a27828a  and  a27813a );
 a1378a <=( a27800a  and  a27785a );
 a1379a <=( a27772a  and  a27757a );
 a1380a <=( a27744a  and  a27729a );
 a1381a <=( a27716a  and  a27701a );
 a1382a <=( a27688a  and  a27673a );
 a1383a <=( a27660a  and  a27645a );
 a1384a <=( a27632a  and  a27617a );
 a1385a <=( a27604a  and  a27589a );
 a1386a <=( a27576a  and  a27561a );
 a1387a <=( a27548a  and  a27533a );
 a1388a <=( a27520a  and  a27505a );
 a1389a <=( a27492a  and  a27477a );
 a1390a <=( a27464a  and  a27449a );
 a1391a <=( a27436a  and  a27421a );
 a1392a <=( a27408a  and  a27393a );
 a1393a <=( a27380a  and  a27365a );
 a1394a <=( a27352a  and  a27337a );
 a1395a <=( a27324a  and  a27309a );
 a1396a <=( a27296a  and  a27281a );
 a1397a <=( a27268a  and  a27253a );
 a1398a <=( a27240a  and  a27225a );
 a1399a <=( a27212a  and  a27197a );
 a1400a <=( a27184a  and  a27169a );
 a1401a <=( a27156a  and  a27141a );
 a1402a <=( a27128a  and  a27113a );
 a1403a <=( a27100a  and  a27085a );
 a1404a <=( a27072a  and  a27057a );
 a1405a <=( a27044a  and  a27029a );
 a1406a <=( a27016a  and  a27001a );
 a1407a <=( a26988a  and  a26973a );
 a1408a <=( a26960a  and  a26945a );
 a1409a <=( a26932a  and  a26917a );
 a1410a <=( a26904a  and  a26889a );
 a1411a <=( a26876a  and  a26861a );
 a1412a <=( a26848a  and  a26833a );
 a1413a <=( a26820a  and  a26805a );
 a1414a <=( a26792a  and  a26777a );
 a1415a <=( a26764a  and  a26749a );
 a1416a <=( a26736a  and  a26721a );
 a1417a <=( a26708a  and  a26693a );
 a1418a <=( a26680a  and  a26665a );
 a1419a <=( a26652a  and  a26637a );
 a1420a <=( a26624a  and  a26609a );
 a1421a <=( a26596a  and  a26581a );
 a1422a <=( a26568a  and  a26553a );
 a1423a <=( a26540a  and  a26525a );
 a1424a <=( a26512a  and  a26497a );
 a1425a <=( a26484a  and  a26469a );
 a1426a <=( a26456a  and  a26441a );
 a1427a <=( a26428a  and  a26413a );
 a1428a <=( a26400a  and  a26385a );
 a1429a <=( a26372a  and  a26357a );
 a1430a <=( a26344a  and  a26329a );
 a1431a <=( a26316a  and  a26301a );
 a1432a <=( a26288a  and  a26273a );
 a1433a <=( a26260a  and  a26245a );
 a1434a <=( a26232a  and  a26217a );
 a1435a <=( a26204a  and  a26189a );
 a1436a <=( a26176a  and  a26161a );
 a1437a <=( a26148a  and  a26133a );
 a1438a <=( a26120a  and  a26105a );
 a1439a <=( a26092a  and  a26077a );
 a1440a <=( a26064a  and  a26049a );
 a1441a <=( a26036a  and  a26021a );
 a1442a <=( a26008a  and  a25993a );
 a1443a <=( a25980a  and  a25965a );
 a1444a <=( a25952a  and  a25937a );
 a1445a <=( a25924a  and  a25909a );
 a1446a <=( a25896a  and  a25881a );
 a1447a <=( a25868a  and  a25853a );
 a1448a <=( a25840a  and  a25825a );
 a1449a <=( a25812a  and  a25797a );
 a1450a <=( a25784a  and  a25769a );
 a1451a <=( a25756a  and  a25741a );
 a1452a <=( a25728a  and  a25713a );
 a1453a <=( a25700a  and  a25685a );
 a1454a <=( a25672a  and  a25657a );
 a1455a <=( a25644a  and  a25629a );
 a1456a <=( a25616a  and  a25601a );
 a1457a <=( a25588a  and  a25573a );
 a1458a <=( a25560a  and  a25545a );
 a1459a <=( a25532a  and  a25517a );
 a1460a <=( a25504a  and  a25489a );
 a1461a <=( a25476a  and  a25461a );
 a1462a <=( a25448a  and  a25433a );
 a1463a <=( a25420a  and  a25405a );
 a1464a <=( a25392a  and  a25377a );
 a1465a <=( a25364a  and  a25349a );
 a1466a <=( a25336a  and  a25321a );
 a1467a <=( a25308a  and  a25293a );
 a1468a <=( a25280a  and  a25265a );
 a1469a <=( a25252a  and  a25237a );
 a1470a <=( a25224a  and  a25209a );
 a1471a <=( a25196a  and  a25181a );
 a1472a <=( a25168a  and  a25153a );
 a1473a <=( a25140a  and  a25125a );
 a1474a <=( a25112a  and  a25097a );
 a1475a <=( a25084a  and  a25069a );
 a1476a <=( a25056a  and  a25041a );
 a1477a <=( a25028a  and  a25013a );
 a1478a <=( a25000a  and  a24985a );
 a1479a <=( a24972a  and  a24957a );
 a1480a <=( a24944a  and  a24929a );
 a1481a <=( a24916a  and  a24901a );
 a1482a <=( a24888a  and  a24873a );
 a1483a <=( a24860a  and  a24845a );
 a1484a <=( a24832a  and  a24817a );
 a1485a <=( a24804a  and  a24789a );
 a1486a <=( a24776a  and  a24761a );
 a1487a <=( a24748a  and  a24733a );
 a1488a <=( a24720a  and  a24705a );
 a1489a <=( a24692a  and  a24677a );
 a1490a <=( a24664a  and  a24649a );
 a1491a <=( a24636a  and  a24621a );
 a1492a <=( a24608a  and  a24593a );
 a1493a <=( a24580a  and  a24565a );
 a1494a <=( a24552a  and  a24537a );
 a1495a <=( a24524a  and  a24509a );
 a1496a <=( a24496a  and  a24481a );
 a1497a <=( a24468a  and  a24453a );
 a1498a <=( a24440a  and  a24425a );
 a1499a <=( a24412a  and  a24397a );
 a1500a <=( a24384a  and  a24369a );
 a1501a <=( a24356a  and  a24341a );
 a1502a <=( a24328a  and  a24313a );
 a1503a <=( a24300a  and  a24285a );
 a1504a <=( a24272a  and  a24257a );
 a1505a <=( a24244a  and  a24229a );
 a1506a <=( a24216a  and  a24201a );
 a1507a <=( a24188a  and  a24173a );
 a1508a <=( a24160a  and  a24145a );
 a1509a <=( a24132a  and  a24117a );
 a1510a <=( a24104a  and  a24089a );
 a1511a <=( a24076a  and  a24061a );
 a1512a <=( a24048a  and  a24033a );
 a1513a <=( a24020a  and  a24005a );
 a1514a <=( a23992a  and  a23977a );
 a1515a <=( a23964a  and  a23949a );
 a1516a <=( a23936a  and  a23921a );
 a1517a <=( a23908a  and  a23893a );
 a1518a <=( a23880a  and  a23865a );
 a1519a <=( a23852a  and  a23837a );
 a1520a <=( a23824a  and  a23809a );
 a1521a <=( a23796a  and  a23781a );
 a1522a <=( a23768a  and  a23753a );
 a1523a <=( a23740a  and  a23725a );
 a1524a <=( a23712a  and  a23697a );
 a1525a <=( a23684a  and  a23669a );
 a1526a <=( a23656a  and  a23641a );
 a1527a <=( a23628a  and  a23613a );
 a1528a <=( a23600a  and  a23585a );
 a1529a <=( a23572a  and  a23557a );
 a1530a <=( a23544a  and  a23529a );
 a1531a <=( a23516a  and  a23501a );
 a1532a <=( a23488a  and  a23473a );
 a1533a <=( a23460a  and  a23445a );
 a1534a <=( a23432a  and  a23417a );
 a1535a <=( a23404a  and  a23389a );
 a1536a <=( a23376a  and  a23361a );
 a1537a <=( a23348a  and  a23333a );
 a1538a <=( a23320a  and  a23305a );
 a1539a <=( a23292a  and  a23277a );
 a1540a <=( a23264a  and  a23249a );
 a1541a <=( a23236a  and  a23221a );
 a1542a <=( a23208a  and  a23193a );
 a1543a <=( a23180a  and  a23165a );
 a1544a <=( a23152a  and  a23137a );
 a1545a <=( a23124a  and  a23109a );
 a1546a <=( a23096a  and  a23081a );
 a1547a <=( a23068a  and  a23053a );
 a1548a <=( a23040a  and  a23025a );
 a1549a <=( a23012a  and  a22997a );
 a1550a <=( a22984a  and  a22969a );
 a1551a <=( a22956a  and  a22941a );
 a1552a <=( a22928a  and  a22913a );
 a1553a <=( a22900a  and  a22885a );
 a1554a <=( a22872a  and  a22857a );
 a1555a <=( a22844a  and  a22829a );
 a1556a <=( a22816a  and  a22801a );
 a1557a <=( a22788a  and  a22773a );
 a1558a <=( a22760a  and  a22745a );
 a1559a <=( a22732a  and  a22717a );
 a1560a <=( a22704a  and  a22689a );
 a1561a <=( a22676a  and  a22661a );
 a1562a <=( a22648a  and  a22633a );
 a1563a <=( a22620a  and  a22605a );
 a1564a <=( a22592a  and  a22577a );
 a1565a <=( a22564a  and  a22549a );
 a1566a <=( a22536a  and  a22521a );
 a1567a <=( a22508a  and  a22493a );
 a1568a <=( a22480a  and  a22465a );
 a1569a <=( a22452a  and  a22437a );
 a1570a <=( a22424a  and  a22409a );
 a1571a <=( a22396a  and  a22381a );
 a1572a <=( a22368a  and  a22353a );
 a1573a <=( a22340a  and  a22325a );
 a1574a <=( a22312a  and  a22297a );
 a1575a <=( a22284a  and  a22269a );
 a1576a <=( a22256a  and  a22241a );
 a1577a <=( a22228a  and  a22213a );
 a1578a <=( a22200a  and  a22185a );
 a1579a <=( a22172a  and  a22157a );
 a1580a <=( a22144a  and  a22129a );
 a1581a <=( a22116a  and  a22101a );
 a1582a <=( a22088a  and  a22073a );
 a1583a <=( a22060a  and  a22045a );
 a1584a <=( a22032a  and  a22017a );
 a1585a <=( a22004a  and  a21989a );
 a1586a <=( a21976a  and  a21961a );
 a1587a <=( a21948a  and  a21933a );
 a1588a <=( a21920a  and  a21905a );
 a1589a <=( a21892a  and  a21877a );
 a1590a <=( a21864a  and  a21849a );
 a1591a <=( a21836a  and  a21821a );
 a1592a <=( a21808a  and  a21793a );
 a1593a <=( a21780a  and  a21765a );
 a1594a <=( a21752a  and  a21737a );
 a1595a <=( a21724a  and  a21709a );
 a1596a <=( a21696a  and  a21681a );
 a1597a <=( a21668a  and  a21653a );
 a1598a <=( a21640a  and  a21625a );
 a1599a <=( a21612a  and  a21597a );
 a1600a <=( a21584a  and  a21569a );
 a1601a <=( a21556a  and  a21541a );
 a1602a <=( a21528a  and  a21513a );
 a1603a <=( a21500a  and  a21485a );
 a1604a <=( a21472a  and  a21457a );
 a1605a <=( a21444a  and  a21429a );
 a1606a <=( a21416a  and  a21401a );
 a1607a <=( a21388a  and  a21373a );
 a1608a <=( a21360a  and  a21345a );
 a1609a <=( a21332a  and  a21317a );
 a1610a <=( a21304a  and  a21289a );
 a1611a <=( a21276a  and  a21261a );
 a1612a <=( a21248a  and  a21233a );
 a1613a <=( a21220a  and  a21205a );
 a1614a <=( a21192a  and  a21177a );
 a1615a <=( a21164a  and  a21149a );
 a1616a <=( a21136a  and  a21121a );
 a1617a <=( a21108a  and  a21093a );
 a1618a <=( a21080a  and  a21065a );
 a1619a <=( a21052a  and  a21037a );
 a1620a <=( a21024a  and  a21009a );
 a1621a <=( a20996a  and  a20981a );
 a1622a <=( a20968a  and  a20953a );
 a1623a <=( a20940a  and  a20925a );
 a1624a <=( a20912a  and  a20897a );
 a1625a <=( a20884a  and  a20869a );
 a1626a <=( a20856a  and  a20841a );
 a1627a <=( a20828a  and  a20813a );
 a1628a <=( a20800a  and  a20785a );
 a1629a <=( a20772a  and  a20757a );
 a1630a <=( a20744a  and  a20729a );
 a1631a <=( a20716a  and  a20701a );
 a1632a <=( a20688a  and  a20673a );
 a1633a <=( a20660a  and  a20645a );
 a1634a <=( a20632a  and  a20617a );
 a1635a <=( a20604a  and  a20589a );
 a1636a <=( a20576a  and  a20561a );
 a1637a <=( a20548a  and  a20533a );
 a1638a <=( a20520a  and  a20505a );
 a1639a <=( a20492a  and  a20477a );
 a1640a <=( a20464a  and  a20449a );
 a1641a <=( a20436a  and  a20421a );
 a1642a <=( a20408a  and  a20393a );
 a1643a <=( a20380a  and  a20365a );
 a1644a <=( a20352a  and  a20337a );
 a1645a <=( a20324a  and  a20309a );
 a1646a <=( a20296a  and  a20281a );
 a1647a <=( a20268a  and  a20253a );
 a1648a <=( a20240a  and  a20225a );
 a1649a <=( a20212a  and  a20199a );
 a1650a <=( a20186a  and  a20173a );
 a1651a <=( a20160a  and  a20147a );
 a1652a <=( a20134a  and  a20121a );
 a1653a <=( a20108a  and  a20095a );
 a1654a <=( a20082a  and  a20069a );
 a1655a <=( a20056a  and  a20043a );
 a1656a <=( a20030a  and  a20017a );
 a1657a <=( a20004a  and  a19991a );
 a1658a <=( a19978a  and  a19965a );
 a1659a <=( a19952a  and  a19939a );
 a1660a <=( a19926a  and  a19913a );
 a1661a <=( a19900a  and  a19887a );
 a1662a <=( a19874a  and  a19861a );
 a1663a <=( a19848a  and  a19835a );
 a1664a <=( a19822a  and  a19809a );
 a1665a <=( a19796a  and  a19783a );
 a1666a <=( a19770a  and  a19757a );
 a1667a <=( a19744a  and  a19731a );
 a1668a <=( a19718a  and  a19705a );
 a1669a <=( a19692a  and  a19679a );
 a1670a <=( a19666a  and  a19653a );
 a1671a <=( a19640a  and  a19627a );
 a1672a <=( a19614a  and  a19601a );
 a1673a <=( a19588a  and  a19575a );
 a1674a <=( a19562a  and  a19549a );
 a1675a <=( a19536a  and  a19523a );
 a1676a <=( a19510a  and  a19497a );
 a1677a <=( a19484a  and  a19471a );
 a1678a <=( a19458a  and  a19445a );
 a1679a <=( a19432a  and  a19419a );
 a1680a <=( a19406a  and  a19393a );
 a1681a <=( a19380a  and  a19367a );
 a1682a <=( a19354a  and  a19341a );
 a1683a <=( a19328a  and  a19315a );
 a1684a <=( a19302a  and  a19289a );
 a1685a <=( a19276a  and  a19263a );
 a1686a <=( a19250a  and  a19237a );
 a1687a <=( a19224a  and  a19211a );
 a1688a <=( a19198a  and  a19185a );
 a1689a <=( a19172a  and  a19159a );
 a1690a <=( a19146a  and  a19133a );
 a1691a <=( a19120a  and  a19107a );
 a1692a <=( a19094a  and  a19081a );
 a1693a <=( a19068a  and  a19055a );
 a1694a <=( a19042a  and  a19029a );
 a1695a <=( a19016a  and  a19003a );
 a1696a <=( a18990a  and  a18977a );
 a1697a <=( a18964a  and  a18951a );
 a1698a <=( a18938a  and  a18925a );
 a1699a <=( a18912a  and  a18899a );
 a1700a <=( a18886a  and  a18873a );
 a1701a <=( a18860a  and  a18847a );
 a1702a <=( a18834a  and  a18821a );
 a1703a <=( a18808a  and  a18795a );
 a1704a <=( a18782a  and  a18769a );
 a1705a <=( a18756a  and  a18743a );
 a1706a <=( a18730a  and  a18717a );
 a1707a <=( a18704a  and  a18691a );
 a1708a <=( a18678a  and  a18665a );
 a1709a <=( a18652a  and  a18639a );
 a1710a <=( a18626a  and  a18613a );
 a1711a <=( a18600a  and  a18587a );
 a1712a <=( a18574a  and  a18561a );
 a1713a <=( a18548a  and  a18535a );
 a1714a <=( a18522a  and  a18509a );
 a1715a <=( a18496a  and  a18483a );
 a1716a <=( a18470a  and  a18457a );
 a1717a <=( a18444a  and  a18431a );
 a1718a <=( a18418a  and  a18405a );
 a1719a <=( a18392a  and  a18379a );
 a1720a <=( a18366a  and  a18353a );
 a1721a <=( a18340a  and  a18327a );
 a1722a <=( a18314a  and  a18301a );
 a1723a <=( a18288a  and  a18275a );
 a1724a <=( a18262a  and  a18249a );
 a1725a <=( a18236a  and  a18223a );
 a1726a <=( a18210a  and  a18197a );
 a1727a <=( a18184a  and  a18171a );
 a1728a <=( a18158a  and  a18145a );
 a1729a <=( a18132a  and  a18119a );
 a1730a <=( a18106a  and  a18093a );
 a1731a <=( a18080a  and  a18067a );
 a1732a <=( a18054a  and  a18041a );
 a1733a <=( a18028a  and  a18015a );
 a1734a <=( a18002a  and  a17989a );
 a1735a <=( a17976a  and  a17963a );
 a1736a <=( a17950a  and  a17937a );
 a1737a <=( a17924a  and  a17911a );
 a1738a <=( a17898a  and  a17885a );
 a1739a <=( a17872a  and  a17859a );
 a1740a <=( a17846a  and  a17833a );
 a1741a <=( a17820a  and  a17807a );
 a1742a <=( a17794a  and  a17781a );
 a1743a <=( a17768a  and  a17755a );
 a1744a <=( a17742a  and  a17729a );
 a1745a <=( a17716a  and  a17703a );
 a1746a <=( a17690a  and  a17677a );
 a1747a <=( a17664a  and  a17651a );
 a1748a <=( a17638a  and  a17625a );
 a1749a <=( a17612a  and  a17599a );
 a1750a <=( a17586a  and  a17573a );
 a1751a <=( a17560a  and  a17547a );
 a1752a <=( a17534a  and  a17521a );
 a1753a <=( a17508a  and  a17495a );
 a1754a <=( a17482a  and  a17469a );
 a1755a <=( a17456a  and  a17443a );
 a1756a <=( a17430a  and  a17417a );
 a1757a <=( a17404a  and  a17391a );
 a1758a <=( a17378a  and  a17365a );
 a1759a <=( a17352a  and  a17339a );
 a1760a <=( a17326a  and  a17313a );
 a1761a <=( a17300a  and  a17287a );
 a1762a <=( a17274a  and  a17261a );
 a1763a <=( a17248a  and  a17235a );
 a1764a <=( a17222a  and  a17209a );
 a1765a <=( a17196a  and  a17183a );
 a1766a <=( a17170a  and  a17157a );
 a1767a <=( a17144a  and  a17131a );
 a1768a <=( a17118a  and  a17105a );
 a1769a <=( a17092a  and  a17079a );
 a1770a <=( a17066a  and  a17053a );
 a1771a <=( a17040a  and  a17027a );
 a1772a <=( a17014a  and  a17001a );
 a1773a <=( a16988a  and  a16975a );
 a1774a <=( a16962a  and  a16949a );
 a1775a <=( a16936a  and  a16923a );
 a1776a <=( a16910a  and  a16897a );
 a1777a <=( a16884a  and  a16871a );
 a1778a <=( a16858a  and  a16845a );
 a1779a <=( a16832a  and  a16819a );
 a1780a <=( a16806a  and  a16793a );
 a1781a <=( a16780a  and  a16767a );
 a1782a <=( a16754a  and  a16741a );
 a1783a <=( a16728a  and  a16715a );
 a1784a <=( a16702a  and  a16689a );
 a1785a <=( a16676a  and  a16663a );
 a1786a <=( a16650a  and  a16637a );
 a1787a <=( a16624a  and  a16611a );
 a1788a <=( a16598a  and  a16585a );
 a1789a <=( a16572a  and  a16559a );
 a1790a <=( a16546a  and  a16533a );
 a1791a <=( a16520a  and  a16507a );
 a1792a <=( a16494a  and  a16481a );
 a1793a <=( a16468a  and  a16455a );
 a1794a <=( a16442a  and  a16429a );
 a1795a <=( a16416a  and  a16403a );
 a1796a <=( a16390a  and  a16377a );
 a1797a <=( a16364a  and  a16351a );
 a1798a <=( a16338a  and  a16325a );
 a1799a <=( a16312a  and  a16299a );
 a1800a <=( a16286a  and  a16273a );
 a1801a <=( a16260a  and  a16247a );
 a1802a <=( a16234a  and  a16221a );
 a1803a <=( a16208a  and  a16195a );
 a1804a <=( a16182a  and  a16169a );
 a1805a <=( a16156a  and  a16143a );
 a1806a <=( a16130a  and  a16117a );
 a1807a <=( a16104a  and  a16091a );
 a1808a <=( a16078a  and  a16065a );
 a1809a <=( a16052a  and  a16039a );
 a1810a <=( a16026a  and  a16013a );
 a1811a <=( a16000a  and  a15987a );
 a1812a <=( a15974a  and  a15961a );
 a1813a <=( a15948a  and  a15935a );
 a1814a <=( a15922a  and  a15909a );
 a1815a <=( a15896a  and  a15883a );
 a1816a <=( a15870a  and  a15857a );
 a1817a <=( a15844a  and  a15831a );
 a1818a <=( a15818a  and  a15805a );
 a1819a <=( a15792a  and  a15779a );
 a1820a <=( a15766a  and  a15753a );
 a1821a <=( a15740a  and  a15727a );
 a1822a <=( a15714a  and  a15701a );
 a1823a <=( a15688a  and  a15675a );
 a1824a <=( a15662a  and  a15649a );
 a1825a <=( a15636a  and  a15623a );
 a1826a <=( a15610a  and  a15597a );
 a1827a <=( a15584a  and  a15571a );
 a1828a <=( a15558a  and  a15545a );
 a1829a <=( a15532a  and  a15519a );
 a1830a <=( a15506a  and  a15493a );
 a1831a <=( a15480a  and  a15467a );
 a1832a <=( a15454a  and  a15441a );
 a1833a <=( a15428a  and  a15415a );
 a1834a <=( a15402a  and  a15389a );
 a1835a <=( a15376a  and  a15363a );
 a1836a <=( a15350a  and  a15337a );
 a1837a <=( a15324a  and  a15311a );
 a1838a <=( a15298a  and  a15285a );
 a1839a <=( a15272a  and  a15259a );
 a1840a <=( a15246a  and  a15233a );
 a1841a <=( a15220a  and  a15207a );
 a1842a <=( a15194a  and  a15181a );
 a1843a <=( a15168a  and  a15155a );
 a1844a <=( a15142a  and  a15129a );
 a1845a <=( a15116a  and  a15103a );
 a1846a <=( a15090a  and  a15077a );
 a1847a <=( a15064a  and  a15051a );
 a1848a <=( a15038a  and  a15025a );
 a1849a <=( a15012a  and  a14999a );
 a1850a <=( a14986a  and  a14973a );
 a1851a <=( a14960a  and  a14947a );
 a1852a <=( a14934a  and  a14921a );
 a1853a <=( a14908a  and  a14895a );
 a1854a <=( a14882a  and  a14869a );
 a1855a <=( a14856a  and  a14843a );
 a1856a <=( a14830a  and  a14817a );
 a1857a <=( a14804a  and  a14791a );
 a1858a <=( a14778a  and  a14765a );
 a1859a <=( a14752a  and  a14739a );
 a1860a <=( a14726a  and  a14713a );
 a1861a <=( a14700a  and  a14687a );
 a1862a <=( a14674a  and  a14661a );
 a1863a <=( a14648a  and  a14635a );
 a1864a <=( a14622a  and  a14609a );
 a1865a <=( a14596a  and  a14583a );
 a1866a <=( a14570a  and  a14557a );
 a1867a <=( a14544a  and  a14531a );
 a1868a <=( a14518a  and  a14505a );
 a1869a <=( a14492a  and  a14479a );
 a1870a <=( a14466a  and  a14453a );
 a1871a <=( a14440a  and  a14427a );
 a1872a <=( a14414a  and  a14401a );
 a1873a <=( a14388a  and  a14375a );
 a1874a <=( a14362a  and  a14349a );
 a1875a <=( a14336a  and  a14323a );
 a1876a <=( a14310a  and  a14297a );
 a1877a <=( a14284a  and  a14271a );
 a1878a <=( a14258a  and  a14245a );
 a1879a <=( a14232a  and  a14219a );
 a1880a <=( a14206a  and  a14193a );
 a1881a <=( a14180a  and  a14167a );
 a1882a <=( a14154a  and  a14141a );
 a1883a <=( a14128a  and  a14115a );
 a1884a <=( a14102a  and  a14089a );
 a1885a <=( a14076a  and  a14063a );
 a1886a <=( a14050a  and  a14037a );
 a1887a <=( a14024a  and  a14011a );
 a1888a <=( a13998a  and  a13985a );
 a1889a <=( a13972a  and  a13959a );
 a1890a <=( a13946a  and  a13933a );
 a1891a <=( a13920a  and  a13907a );
 a1892a <=( a13894a  and  a13881a );
 a1893a <=( a13868a  and  a13855a );
 a1894a <=( a13842a  and  a13829a );
 a1895a <=( a13816a  and  a13803a );
 a1896a <=( a13790a  and  a13777a );
 a1897a <=( a13764a  and  a13751a );
 a1898a <=( a13738a  and  a13725a );
 a1899a <=( a13712a  and  a13699a );
 a1900a <=( a13686a  and  a13673a );
 a1901a <=( a13660a  and  a13647a );
 a1902a <=( a13634a  and  a13621a );
 a1903a <=( a13608a  and  a13595a );
 a1904a <=( a13582a  and  a13569a );
 a1905a <=( a13556a  and  a13543a );
 a1906a <=( a13530a  and  a13517a );
 a1907a <=( a13504a  and  a13491a );
 a1908a <=( a13478a  and  a13465a );
 a1909a <=( a13452a  and  a13439a );
 a1910a <=( a13426a  and  a13413a );
 a1911a <=( a13400a  and  a13387a );
 a1912a <=( a13374a  and  a13361a );
 a1913a <=( a13348a  and  a13335a );
 a1914a <=( a13322a  and  a13309a );
 a1915a <=( a13296a  and  a13283a );
 a1916a <=( a13270a  and  a13257a );
 a1917a <=( a13244a  and  a13231a );
 a1918a <=( a13218a  and  a13205a );
 a1919a <=( a13192a  and  a13179a );
 a1920a <=( a13166a  and  a13153a );
 a1921a <=( a13140a  and  a13127a );
 a1922a <=( a13114a  and  a13101a );
 a1923a <=( a13088a  and  a13075a );
 a1924a <=( a13062a  and  a13049a );
 a1925a <=( a13036a  and  a13023a );
 a1926a <=( a13010a  and  a12997a );
 a1927a <=( a12984a  and  a12971a );
 a1928a <=( a12958a  and  a12945a );
 a1929a <=( a12932a  and  a12919a );
 a1930a <=( a12906a  and  a12893a );
 a1931a <=( a12880a  and  a12867a );
 a1932a <=( a12854a  and  a12841a );
 a1933a <=( a12828a  and  a12815a );
 a1934a <=( a12802a  and  a12789a );
 a1935a <=( a12776a  and  a12763a );
 a1936a <=( a12750a  and  a12737a );
 a1937a <=( a12724a  and  a12711a );
 a1938a <=( a12698a  and  a12685a );
 a1939a <=( a12672a  and  a12659a );
 a1940a <=( a12646a  and  a12633a );
 a1941a <=( a12620a  and  a12607a );
 a1942a <=( a12594a  and  a12581a );
 a1943a <=( a12568a  and  a12555a );
 a1944a <=( a12542a  and  a12529a );
 a1945a <=( a12516a  and  a12503a );
 a1946a <=( a12490a  and  a12477a );
 a1947a <=( a12464a  and  a12451a );
 a1948a <=( a12438a  and  a12425a );
 a1949a <=( a12412a  and  a12399a );
 a1950a <=( a12386a  and  a12373a );
 a1951a <=( a12360a  and  a12347a );
 a1952a <=( a12334a  and  a12321a );
 a1953a <=( a12308a  and  a12295a );
 a1954a <=( a12282a  and  a12269a );
 a1955a <=( a12256a  and  a12243a );
 a1956a <=( a12230a  and  a12217a );
 a1957a <=( a12204a  and  a12191a );
 a1958a <=( a12178a  and  a12165a );
 a1959a <=( a12152a  and  a12139a );
 a1960a <=( a12126a  and  a12113a );
 a1961a <=( a12100a  and  a12087a );
 a1962a <=( a12074a  and  a12061a );
 a1963a <=( a12048a  and  a12035a );
 a1964a <=( a12022a  and  a12009a );
 a1965a <=( a11996a  and  a11983a );
 a1966a <=( a11970a  and  a11957a );
 a1967a <=( a11944a  and  a11931a );
 a1968a <=( a11918a  and  a11905a );
 a1969a <=( a11892a  and  a11879a );
 a1970a <=( a11866a  and  a11853a );
 a1971a <=( a11840a  and  a11827a );
 a1972a <=( a11814a  and  a11801a );
 a1973a <=( a11788a  and  a11775a );
 a1974a <=( a11762a  and  a11749a );
 a1975a <=( a11736a  and  a11723a );
 a1976a <=( a11710a  and  a11697a );
 a1977a <=( a11684a  and  a11671a );
 a1978a <=( a11658a  and  a11645a );
 a1979a <=( a11632a  and  a11619a );
 a1980a <=( a11606a  and  a11593a );
 a1981a <=( a11580a  and  a11567a );
 a1982a <=( a11554a  and  a11541a );
 a1983a <=( a11528a  and  a11515a );
 a1984a <=( a11502a  and  a11489a );
 a1985a <=( a11476a  and  a11463a );
 a1986a <=( a11450a  and  a11437a );
 a1987a <=( a11424a  and  a11411a );
 a1988a <=( a11398a  and  a11385a );
 a1989a <=( a11372a  and  a11359a );
 a1990a <=( a11346a  and  a11333a );
 a1991a <=( a11320a  and  a11307a );
 a1992a <=( a11294a  and  a11281a );
 a1993a <=( a11268a  and  a11255a );
 a1994a <=( a11242a  and  a11229a );
 a1995a <=( a11216a  and  a11203a );
 a1996a <=( a11190a  and  a11177a );
 a1997a <=( a11164a  and  a11151a );
 a1998a <=( a11138a  and  a11125a );
 a1999a <=( a11112a  and  a11099a );
 a2000a <=( a11086a  and  a11073a );
 a2001a <=( a11060a  and  a11047a );
 a2002a <=( a11034a  and  a11021a );
 a2003a <=( a11008a  and  a10995a );
 a2004a <=( a10982a  and  a10969a );
 a2005a <=( a10956a  and  a10943a );
 a2006a <=( a10930a  and  a10917a );
 a2007a <=( a10904a  and  a10891a );
 a2008a <=( a10878a  and  a10865a );
 a2009a <=( a10852a  and  a10839a );
 a2010a <=( a10826a  and  a10813a );
 a2011a <=( a10800a  and  a10787a );
 a2012a <=( a10774a  and  a10761a );
 a2013a <=( a10748a  and  a10735a );
 a2014a <=( a10722a  and  a10709a );
 a2015a <=( a10696a  and  a10683a );
 a2016a <=( a10670a  and  a10657a );
 a2017a <=( a10644a  and  a10631a );
 a2018a <=( a10618a  and  a10605a );
 a2019a <=( a10592a  and  a10579a );
 a2020a <=( a10566a  and  a10553a );
 a2021a <=( a10540a  and  a10527a );
 a2022a <=( a10514a  and  a10501a );
 a2023a <=( a10488a  and  a10475a );
 a2024a <=( a10462a  and  a10449a );
 a2025a <=( a10436a  and  a10423a );
 a2026a <=( a10410a  and  a10397a );
 a2027a <=( a10384a  and  a10371a );
 a2028a <=( a10358a  and  a10345a );
 a2029a <=( a10332a  and  a10319a );
 a2030a <=( a10306a  and  a10293a );
 a2031a <=( a10280a  and  a10267a );
 a2032a <=( a10254a  and  a10241a );
 a2033a <=( a10228a  and  a10215a );
 a2034a <=( a10202a  and  a10189a );
 a2035a <=( a10176a  and  a10163a );
 a2036a <=( a10150a  and  a10137a );
 a2037a <=( a10124a  and  a10111a );
 a2038a <=( a10098a  and  a10085a );
 a2039a <=( a10072a  and  a10059a );
 a2040a <=( a10046a  and  a10033a );
 a2041a <=( a10020a  and  a10007a );
 a2042a <=( a9994a  and  a9981a );
 a2043a <=( a9968a  and  a9955a );
 a2044a <=( a9942a  and  a9929a );
 a2045a <=( a9916a  and  a9903a );
 a2046a <=( a9890a  and  a9877a );
 a2047a <=( a9864a  and  a9851a );
 a2048a <=( a9838a  and  a9825a );
 a2049a <=( a9812a  and  a9799a );
 a2050a <=( a9786a  and  a9773a );
 a2051a <=( a9760a  and  a9747a );
 a2052a <=( a9734a  and  a9721a );
 a2053a <=( a9708a  and  a9695a );
 a2054a <=( a9682a  and  a9669a );
 a2055a <=( a9656a  and  a9643a );
 a2056a <=( a9630a  and  a9617a );
 a2057a <=( a9604a  and  a9591a );
 a2058a <=( a9578a  and  a9565a );
 a2059a <=( a9552a  and  a9539a );
 a2060a <=( a9526a  and  a9513a );
 a2061a <=( a9500a  and  a9487a );
 a2062a <=( a9474a  and  a9461a );
 a2063a <=( a9448a  and  a9435a );
 a2064a <=( a9422a  and  a9409a );
 a2065a <=( a9396a  and  a9383a );
 a2066a <=( a9370a  and  a9357a );
 a2067a <=( a9344a  and  a9331a );
 a2068a <=( a9318a  and  a9305a );
 a2069a <=( a9292a  and  a9279a );
 a2070a <=( a9266a  and  a9253a );
 a2071a <=( a9240a  and  a9227a );
 a2072a <=( a9214a  and  a9201a );
 a2073a <=( a9188a  and  a9175a );
 a2074a <=( a9162a  and  a9149a );
 a2075a <=( a9136a  and  a9123a );
 a2076a <=( a9110a  and  a9097a );
 a2077a <=( a9084a  and  a9071a );
 a2078a <=( a9058a  and  a9045a );
 a2079a <=( a9032a  and  a9019a );
 a2080a <=( a9006a  and  a8993a );
 a2081a <=( a8980a  and  a8967a );
 a2082a <=( a8954a  and  a8941a );
 a2083a <=( a8928a  and  a8915a );
 a2084a <=( a8902a  and  a8889a );
 a2085a <=( a8876a  and  a8863a );
 a2086a <=( a8850a  and  a8837a );
 a2087a <=( a8824a  and  a8811a );
 a2088a <=( a8798a  and  a8785a );
 a2089a <=( a8772a  and  a8759a );
 a2090a <=( a8746a  and  a8733a );
 a2091a <=( a8720a  and  a8707a );
 a2092a <=( a8694a  and  a8681a );
 a2093a <=( a8668a  and  a8655a );
 a2094a <=( a8642a  and  a8629a );
 a2095a <=( a8616a  and  a8603a );
 a2096a <=( a8590a  and  a8577a );
 a2097a <=( a8564a  and  a8551a );
 a2098a <=( a8538a  and  a8525a );
 a2099a <=( a8512a  and  a8499a );
 a2100a <=( a8486a  and  a8473a );
 a2101a <=( a8460a  and  a8447a );
 a2102a <=( a8434a  and  a8421a );
 a2103a <=( a8408a  and  a8395a );
 a2104a <=( a8382a  and  a8369a );
 a2105a <=( a8356a  and  a8343a );
 a2106a <=( a8330a  and  a8317a );
 a2107a <=( a8304a  and  a8291a );
 a2108a <=( a8278a  and  a8265a );
 a2109a <=( a8252a  and  a8239a );
 a2110a <=( a8226a  and  a8213a );
 a2111a <=( a8200a  and  a8187a );
 a2112a <=( a8174a  and  a8161a );
 a2113a <=( a8148a  and  a8135a );
 a2114a <=( a8122a  and  a8109a );
 a2115a <=( a8096a  and  a8083a );
 a2116a <=( a8070a  and  a8057a );
 a2117a <=( a8044a  and  a8031a );
 a2118a <=( a8018a  and  a8005a );
 a2119a <=( a7992a  and  a7979a );
 a2120a <=( a7966a  and  a7953a );
 a2121a <=( a7940a  and  a7927a );
 a2122a <=( a7914a  and  a7901a );
 a2123a <=( a7888a  and  a7875a );
 a2124a <=( a7862a  and  a7849a );
 a2125a <=( a7836a  and  a7823a );
 a2126a <=( a7810a  and  a7797a );
 a2127a <=( a7784a  and  a7771a );
 a2128a <=( a7758a  and  a7745a );
 a2129a <=( a7732a  and  a7719a );
 a2130a <=( a7706a  and  a7693a );
 a2131a <=( a7680a  and  a7667a );
 a2132a <=( a7654a  and  a7641a );
 a2133a <=( a7628a  and  a7615a );
 a2134a <=( a7602a  and  a7589a );
 a2135a <=( a7576a  and  a7563a );
 a2136a <=( a7550a  and  a7537a );
 a2137a <=( a7524a  and  a7511a );
 a2138a <=( a7498a  and  a7485a );
 a2139a <=( a7472a  and  a7459a );
 a2140a <=( a7446a  and  a7433a );
 a2141a <=( a7420a  and  a7407a );
 a2142a <=( a7394a  and  a7381a );
 a2143a <=( a7368a  and  a7355a );
 a2144a <=( a7342a  and  a7329a );
 a2145a <=( a7316a  and  a7303a );
 a2146a <=( a7290a  and  a7277a );
 a2147a <=( a7264a  and  a7251a );
 a2148a <=( a7238a  and  a7225a );
 a2149a <=( a7212a  and  a7199a );
 a2150a <=( a7186a  and  a7173a );
 a2151a <=( a7160a  and  a7147a );
 a2152a <=( a7134a  and  a7121a );
 a2153a <=( a7108a  and  a7095a );
 a2154a <=( a7082a  and  a7069a );
 a2155a <=( a7056a  and  a7043a );
 a2156a <=( a7030a  and  a7017a );
 a2157a <=( a7004a  and  a6991a );
 a2158a <=( a6978a  and  a6965a );
 a2159a <=( a6952a  and  a6939a );
 a2160a <=( a6926a  and  a6913a );
 a2161a <=( a6900a  and  a6893a );
 a2162a <=( a6886a  and  a6879a );
 a2163a <=( a6872a  and  a6865a );
 a2164a <=( a6860a  and  a6853a );
 a2165a <=( a6848a  and  a6841a );
 a2166a <=( a6836a  and  a6829a );
 a2167a <=( a6824a  and  a6817a );
 a2168a <=( a6812a  and  a6805a );
 a2169a <=( a6800a  and  a6793a );
 a2170a <=( a6788a  and  a6781a );
 a2171a <=( a6776a  and  a6769a );
 a2172a <=( a6764a  and  a6757a );
 a2173a <=( a6752a  and  a6745a );
 a2174a <=( a6740a  and  a6733a );
 a2175a <=( a6728a  and  a6723a );
 a2176a <=( a6718a  and  a6713a );
 a2177a <=( a6708a  and  a6703a );
 a2178a <=( a6698a  and  a6693a );
 a2179a <=( a6688a  and  a6683a );
 a2180a <=( a6678a  and  a6673a );
 a2181a <=( a6668a  and  a6663a );
 a2182a <=( a6658a  and  a6653a );
 a2183a <=( a6648a  and  a6643a );
 a2184a <=( a6638a  and  a6633a );
 a2185a <=( a6628a  and  a6623a );
 a2186a <=( a6618a  and  a6613a );
 a2187a <=( a6608a  and  a6603a );
 a2188a <=( a6598a  and  a6593a );
 a2189a <=( a6588a  and  a6583a );
 a2190a <=( a6578a  and  a6573a );
 a2193a <=( a2189a ) or ( a2190a );
 a2196a <=( a2187a ) or ( a2188a );
 a2197a <=( a2196a ) or ( a2193a );
 a2200a <=( a2185a ) or ( a2186a );
 a2203a <=( a2183a ) or ( a2184a );
 a2204a <=( a2203a ) or ( a2200a );
 a2205a <=( a2204a ) or ( a2197a );
 a2208a <=( a2181a ) or ( a2182a );
 a2211a <=( a2179a ) or ( a2180a );
 a2212a <=( a2211a ) or ( a2208a );
 a2215a <=( a2177a ) or ( a2178a );
 a2219a <=( a2174a ) or ( a2175a );
 a2220a <=( a2176a ) or ( a2219a );
 a2221a <=( a2220a ) or ( a2215a );
 a2222a <=( a2221a ) or ( a2212a );
 a2223a <=( a2222a ) or ( a2205a );
 a2226a <=( a2172a ) or ( a2173a );
 a2229a <=( a2170a ) or ( a2171a );
 a2230a <=( a2229a ) or ( a2226a );
 a2233a <=( a2168a ) or ( a2169a );
 a2236a <=( a2166a ) or ( a2167a );
 a2237a <=( a2236a ) or ( a2233a );
 a2238a <=( a2237a ) or ( a2230a );
 a2241a <=( a2164a ) or ( a2165a );
 a2244a <=( a2162a ) or ( a2163a );
 a2245a <=( a2244a ) or ( a2241a );
 a2248a <=( a2160a ) or ( a2161a );
 a2252a <=( a2157a ) or ( a2158a );
 a2253a <=( a2159a ) or ( a2252a );
 a2254a <=( a2253a ) or ( a2248a );
 a2255a <=( a2254a ) or ( a2245a );
 a2256a <=( a2255a ) or ( a2238a );
 a2257a <=( a2256a ) or ( a2223a );
 a2260a <=( a2155a ) or ( a2156a );
 a2263a <=( a2153a ) or ( a2154a );
 a2264a <=( a2263a ) or ( a2260a );
 a2267a <=( a2151a ) or ( a2152a );
 a2270a <=( a2149a ) or ( a2150a );
 a2271a <=( a2270a ) or ( a2267a );
 a2272a <=( a2271a ) or ( a2264a );
 a2275a <=( a2147a ) or ( a2148a );
 a2278a <=( a2145a ) or ( a2146a );
 a2279a <=( a2278a ) or ( a2275a );
 a2282a <=( a2143a ) or ( a2144a );
 a2286a <=( a2140a ) or ( a2141a );
 a2287a <=( a2142a ) or ( a2286a );
 a2288a <=( a2287a ) or ( a2282a );
 a2289a <=( a2288a ) or ( a2279a );
 a2290a <=( a2289a ) or ( a2272a );
 a2293a <=( a2138a ) or ( a2139a );
 a2296a <=( a2136a ) or ( a2137a );
 a2297a <=( a2296a ) or ( a2293a );
 a2300a <=( a2134a ) or ( a2135a );
 a2303a <=( a2132a ) or ( a2133a );
 a2304a <=( a2303a ) or ( a2300a );
 a2305a <=( a2304a ) or ( a2297a );
 a2308a <=( a2130a ) or ( a2131a );
 a2311a <=( a2128a ) or ( a2129a );
 a2312a <=( a2311a ) or ( a2308a );
 a2315a <=( a2126a ) or ( a2127a );
 a2319a <=( a2123a ) or ( a2124a );
 a2320a <=( a2125a ) or ( a2319a );
 a2321a <=( a2320a ) or ( a2315a );
 a2322a <=( a2321a ) or ( a2312a );
 a2323a <=( a2322a ) or ( a2305a );
 a2324a <=( a2323a ) or ( a2290a );
 a2325a <=( a2324a ) or ( a2257a );
 a2328a <=( a2121a ) or ( a2122a );
 a2331a <=( a2119a ) or ( a2120a );
 a2332a <=( a2331a ) or ( a2328a );
 a2335a <=( a2117a ) or ( a2118a );
 a2338a <=( a2115a ) or ( a2116a );
 a2339a <=( a2338a ) or ( a2335a );
 a2340a <=( a2339a ) or ( a2332a );
 a2343a <=( a2113a ) or ( a2114a );
 a2346a <=( a2111a ) or ( a2112a );
 a2347a <=( a2346a ) or ( a2343a );
 a2350a <=( a2109a ) or ( a2110a );
 a2354a <=( a2106a ) or ( a2107a );
 a2355a <=( a2108a ) or ( a2354a );
 a2356a <=( a2355a ) or ( a2350a );
 a2357a <=( a2356a ) or ( a2347a );
 a2358a <=( a2357a ) or ( a2340a );
 a2361a <=( a2104a ) or ( a2105a );
 a2364a <=( a2102a ) or ( a2103a );
 a2365a <=( a2364a ) or ( a2361a );
 a2368a <=( a2100a ) or ( a2101a );
 a2371a <=( a2098a ) or ( a2099a );
 a2372a <=( a2371a ) or ( a2368a );
 a2373a <=( a2372a ) or ( a2365a );
 a2376a <=( a2096a ) or ( a2097a );
 a2379a <=( a2094a ) or ( a2095a );
 a2380a <=( a2379a ) or ( a2376a );
 a2383a <=( a2092a ) or ( a2093a );
 a2387a <=( a2089a ) or ( a2090a );
 a2388a <=( a2091a ) or ( a2387a );
 a2389a <=( a2388a ) or ( a2383a );
 a2390a <=( a2389a ) or ( a2380a );
 a2391a <=( a2390a ) or ( a2373a );
 a2392a <=( a2391a ) or ( a2358a );
 a2395a <=( a2087a ) or ( a2088a );
 a2398a <=( a2085a ) or ( a2086a );
 a2399a <=( a2398a ) or ( a2395a );
 a2402a <=( a2083a ) or ( a2084a );
 a2405a <=( a2081a ) or ( a2082a );
 a2406a <=( a2405a ) or ( a2402a );
 a2407a <=( a2406a ) or ( a2399a );
 a2410a <=( a2079a ) or ( a2080a );
 a2413a <=( a2077a ) or ( a2078a );
 a2414a <=( a2413a ) or ( a2410a );
 a2417a <=( a2075a ) or ( a2076a );
 a2421a <=( a2072a ) or ( a2073a );
 a2422a <=( a2074a ) or ( a2421a );
 a2423a <=( a2422a ) or ( a2417a );
 a2424a <=( a2423a ) or ( a2414a );
 a2425a <=( a2424a ) or ( a2407a );
 a2428a <=( a2070a ) or ( a2071a );
 a2431a <=( a2068a ) or ( a2069a );
 a2432a <=( a2431a ) or ( a2428a );
 a2435a <=( a2066a ) or ( a2067a );
 a2438a <=( a2064a ) or ( a2065a );
 a2439a <=( a2438a ) or ( a2435a );
 a2440a <=( a2439a ) or ( a2432a );
 a2443a <=( a2062a ) or ( a2063a );
 a2446a <=( a2060a ) or ( a2061a );
 a2447a <=( a2446a ) or ( a2443a );
 a2450a <=( a2058a ) or ( a2059a );
 a2454a <=( a2055a ) or ( a2056a );
 a2455a <=( a2057a ) or ( a2454a );
 a2456a <=( a2455a ) or ( a2450a );
 a2457a <=( a2456a ) or ( a2447a );
 a2458a <=( a2457a ) or ( a2440a );
 a2459a <=( a2458a ) or ( a2425a );
 a2460a <=( a2459a ) or ( a2392a );
 a2461a <=( a2460a ) or ( a2325a );
 a2464a <=( a2053a ) or ( a2054a );
 a2467a <=( a2051a ) or ( a2052a );
 a2468a <=( a2467a ) or ( a2464a );
 a2471a <=( a2049a ) or ( a2050a );
 a2474a <=( a2047a ) or ( a2048a );
 a2475a <=( a2474a ) or ( a2471a );
 a2476a <=( a2475a ) or ( a2468a );
 a2479a <=( a2045a ) or ( a2046a );
 a2482a <=( a2043a ) or ( a2044a );
 a2483a <=( a2482a ) or ( a2479a );
 a2486a <=( a2041a ) or ( a2042a );
 a2490a <=( a2038a ) or ( a2039a );
 a2491a <=( a2040a ) or ( a2490a );
 a2492a <=( a2491a ) or ( a2486a );
 a2493a <=( a2492a ) or ( a2483a );
 a2494a <=( a2493a ) or ( a2476a );
 a2497a <=( a2036a ) or ( a2037a );
 a2500a <=( a2034a ) or ( a2035a );
 a2501a <=( a2500a ) or ( a2497a );
 a2504a <=( a2032a ) or ( a2033a );
 a2507a <=( a2030a ) or ( a2031a );
 a2508a <=( a2507a ) or ( a2504a );
 a2509a <=( a2508a ) or ( a2501a );
 a2512a <=( a2028a ) or ( a2029a );
 a2515a <=( a2026a ) or ( a2027a );
 a2516a <=( a2515a ) or ( a2512a );
 a2519a <=( a2024a ) or ( a2025a );
 a2523a <=( a2021a ) or ( a2022a );
 a2524a <=( a2023a ) or ( a2523a );
 a2525a <=( a2524a ) or ( a2519a );
 a2526a <=( a2525a ) or ( a2516a );
 a2527a <=( a2526a ) or ( a2509a );
 a2528a <=( a2527a ) or ( a2494a );
 a2531a <=( a2019a ) or ( a2020a );
 a2534a <=( a2017a ) or ( a2018a );
 a2535a <=( a2534a ) or ( a2531a );
 a2538a <=( a2015a ) or ( a2016a );
 a2541a <=( a2013a ) or ( a2014a );
 a2542a <=( a2541a ) or ( a2538a );
 a2543a <=( a2542a ) or ( a2535a );
 a2546a <=( a2011a ) or ( a2012a );
 a2549a <=( a2009a ) or ( a2010a );
 a2550a <=( a2549a ) or ( a2546a );
 a2553a <=( a2007a ) or ( a2008a );
 a2557a <=( a2004a ) or ( a2005a );
 a2558a <=( a2006a ) or ( a2557a );
 a2559a <=( a2558a ) or ( a2553a );
 a2560a <=( a2559a ) or ( a2550a );
 a2561a <=( a2560a ) or ( a2543a );
 a2564a <=( a2002a ) or ( a2003a );
 a2567a <=( a2000a ) or ( a2001a );
 a2568a <=( a2567a ) or ( a2564a );
 a2571a <=( a1998a ) or ( a1999a );
 a2574a <=( a1996a ) or ( a1997a );
 a2575a <=( a2574a ) or ( a2571a );
 a2576a <=( a2575a ) or ( a2568a );
 a2579a <=( a1994a ) or ( a1995a );
 a2582a <=( a1992a ) or ( a1993a );
 a2583a <=( a2582a ) or ( a2579a );
 a2586a <=( a1990a ) or ( a1991a );
 a2590a <=( a1987a ) or ( a1988a );
 a2591a <=( a1989a ) or ( a2590a );
 a2592a <=( a2591a ) or ( a2586a );
 a2593a <=( a2592a ) or ( a2583a );
 a2594a <=( a2593a ) or ( a2576a );
 a2595a <=( a2594a ) or ( a2561a );
 a2596a <=( a2595a ) or ( a2528a );
 a2599a <=( a1985a ) or ( a1986a );
 a2602a <=( a1983a ) or ( a1984a );
 a2603a <=( a2602a ) or ( a2599a );
 a2606a <=( a1981a ) or ( a1982a );
 a2609a <=( a1979a ) or ( a1980a );
 a2610a <=( a2609a ) or ( a2606a );
 a2611a <=( a2610a ) or ( a2603a );
 a2614a <=( a1977a ) or ( a1978a );
 a2617a <=( a1975a ) or ( a1976a );
 a2618a <=( a2617a ) or ( a2614a );
 a2621a <=( a1973a ) or ( a1974a );
 a2625a <=( a1970a ) or ( a1971a );
 a2626a <=( a1972a ) or ( a2625a );
 a2627a <=( a2626a ) or ( a2621a );
 a2628a <=( a2627a ) or ( a2618a );
 a2629a <=( a2628a ) or ( a2611a );
 a2632a <=( a1968a ) or ( a1969a );
 a2635a <=( a1966a ) or ( a1967a );
 a2636a <=( a2635a ) or ( a2632a );
 a2639a <=( a1964a ) or ( a1965a );
 a2642a <=( a1962a ) or ( a1963a );
 a2643a <=( a2642a ) or ( a2639a );
 a2644a <=( a2643a ) or ( a2636a );
 a2647a <=( a1960a ) or ( a1961a );
 a2650a <=( a1958a ) or ( a1959a );
 a2651a <=( a2650a ) or ( a2647a );
 a2654a <=( a1956a ) or ( a1957a );
 a2658a <=( a1953a ) or ( a1954a );
 a2659a <=( a1955a ) or ( a2658a );
 a2660a <=( a2659a ) or ( a2654a );
 a2661a <=( a2660a ) or ( a2651a );
 a2662a <=( a2661a ) or ( a2644a );
 a2663a <=( a2662a ) or ( a2629a );
 a2666a <=( a1951a ) or ( a1952a );
 a2669a <=( a1949a ) or ( a1950a );
 a2670a <=( a2669a ) or ( a2666a );
 a2673a <=( a1947a ) or ( a1948a );
 a2676a <=( a1945a ) or ( a1946a );
 a2677a <=( a2676a ) or ( a2673a );
 a2678a <=( a2677a ) or ( a2670a );
 a2681a <=( a1943a ) or ( a1944a );
 a2684a <=( a1941a ) or ( a1942a );
 a2685a <=( a2684a ) or ( a2681a );
 a2688a <=( a1939a ) or ( a1940a );
 a2692a <=( a1936a ) or ( a1937a );
 a2693a <=( a1938a ) or ( a2692a );
 a2694a <=( a2693a ) or ( a2688a );
 a2695a <=( a2694a ) or ( a2685a );
 a2696a <=( a2695a ) or ( a2678a );
 a2699a <=( a1934a ) or ( a1935a );
 a2702a <=( a1932a ) or ( a1933a );
 a2703a <=( a2702a ) or ( a2699a );
 a2706a <=( a1930a ) or ( a1931a );
 a2710a <=( a1927a ) or ( a1928a );
 a2711a <=( a1929a ) or ( a2710a );
 a2712a <=( a2711a ) or ( a2706a );
 a2713a <=( a2712a ) or ( a2703a );
 a2716a <=( a1925a ) or ( a1926a );
 a2719a <=( a1923a ) or ( a1924a );
 a2720a <=( a2719a ) or ( a2716a );
 a2723a <=( a1921a ) or ( a1922a );
 a2727a <=( a1918a ) or ( a1919a );
 a2728a <=( a1920a ) or ( a2727a );
 a2729a <=( a2728a ) or ( a2723a );
 a2730a <=( a2729a ) or ( a2720a );
 a2731a <=( a2730a ) or ( a2713a );
 a2732a <=( a2731a ) or ( a2696a );
 a2733a <=( a2732a ) or ( a2663a );
 a2734a <=( a2733a ) or ( a2596a );
 a2735a <=( a2734a ) or ( a2461a );
 a2738a <=( a1916a ) or ( a1917a );
 a2741a <=( a1914a ) or ( a1915a );
 a2742a <=( a2741a ) or ( a2738a );
 a2745a <=( a1912a ) or ( a1913a );
 a2748a <=( a1910a ) or ( a1911a );
 a2749a <=( a2748a ) or ( a2745a );
 a2750a <=( a2749a ) or ( a2742a );
 a2753a <=( a1908a ) or ( a1909a );
 a2756a <=( a1906a ) or ( a1907a );
 a2757a <=( a2756a ) or ( a2753a );
 a2760a <=( a1904a ) or ( a1905a );
 a2764a <=( a1901a ) or ( a1902a );
 a2765a <=( a1903a ) or ( a2764a );
 a2766a <=( a2765a ) or ( a2760a );
 a2767a <=( a2766a ) or ( a2757a );
 a2768a <=( a2767a ) or ( a2750a );
 a2771a <=( a1899a ) or ( a1900a );
 a2774a <=( a1897a ) or ( a1898a );
 a2775a <=( a2774a ) or ( a2771a );
 a2778a <=( a1895a ) or ( a1896a );
 a2781a <=( a1893a ) or ( a1894a );
 a2782a <=( a2781a ) or ( a2778a );
 a2783a <=( a2782a ) or ( a2775a );
 a2786a <=( a1891a ) or ( a1892a );
 a2789a <=( a1889a ) or ( a1890a );
 a2790a <=( a2789a ) or ( a2786a );
 a2793a <=( a1887a ) or ( a1888a );
 a2797a <=( a1884a ) or ( a1885a );
 a2798a <=( a1886a ) or ( a2797a );
 a2799a <=( a2798a ) or ( a2793a );
 a2800a <=( a2799a ) or ( a2790a );
 a2801a <=( a2800a ) or ( a2783a );
 a2802a <=( a2801a ) or ( a2768a );
 a2805a <=( a1882a ) or ( a1883a );
 a2808a <=( a1880a ) or ( a1881a );
 a2809a <=( a2808a ) or ( a2805a );
 a2812a <=( a1878a ) or ( a1879a );
 a2815a <=( a1876a ) or ( a1877a );
 a2816a <=( a2815a ) or ( a2812a );
 a2817a <=( a2816a ) or ( a2809a );
 a2820a <=( a1874a ) or ( a1875a );
 a2823a <=( a1872a ) or ( a1873a );
 a2824a <=( a2823a ) or ( a2820a );
 a2827a <=( a1870a ) or ( a1871a );
 a2831a <=( a1867a ) or ( a1868a );
 a2832a <=( a1869a ) or ( a2831a );
 a2833a <=( a2832a ) or ( a2827a );
 a2834a <=( a2833a ) or ( a2824a );
 a2835a <=( a2834a ) or ( a2817a );
 a2838a <=( a1865a ) or ( a1866a );
 a2841a <=( a1863a ) or ( a1864a );
 a2842a <=( a2841a ) or ( a2838a );
 a2845a <=( a1861a ) or ( a1862a );
 a2848a <=( a1859a ) or ( a1860a );
 a2849a <=( a2848a ) or ( a2845a );
 a2850a <=( a2849a ) or ( a2842a );
 a2853a <=( a1857a ) or ( a1858a );
 a2856a <=( a1855a ) or ( a1856a );
 a2857a <=( a2856a ) or ( a2853a );
 a2860a <=( a1853a ) or ( a1854a );
 a2864a <=( a1850a ) or ( a1851a );
 a2865a <=( a1852a ) or ( a2864a );
 a2866a <=( a2865a ) or ( a2860a );
 a2867a <=( a2866a ) or ( a2857a );
 a2868a <=( a2867a ) or ( a2850a );
 a2869a <=( a2868a ) or ( a2835a );
 a2870a <=( a2869a ) or ( a2802a );
 a2873a <=( a1848a ) or ( a1849a );
 a2876a <=( a1846a ) or ( a1847a );
 a2877a <=( a2876a ) or ( a2873a );
 a2880a <=( a1844a ) or ( a1845a );
 a2883a <=( a1842a ) or ( a1843a );
 a2884a <=( a2883a ) or ( a2880a );
 a2885a <=( a2884a ) or ( a2877a );
 a2888a <=( a1840a ) or ( a1841a );
 a2891a <=( a1838a ) or ( a1839a );
 a2892a <=( a2891a ) or ( a2888a );
 a2895a <=( a1836a ) or ( a1837a );
 a2899a <=( a1833a ) or ( a1834a );
 a2900a <=( a1835a ) or ( a2899a );
 a2901a <=( a2900a ) or ( a2895a );
 a2902a <=( a2901a ) or ( a2892a );
 a2903a <=( a2902a ) or ( a2885a );
 a2906a <=( a1831a ) or ( a1832a );
 a2909a <=( a1829a ) or ( a1830a );
 a2910a <=( a2909a ) or ( a2906a );
 a2913a <=( a1827a ) or ( a1828a );
 a2916a <=( a1825a ) or ( a1826a );
 a2917a <=( a2916a ) or ( a2913a );
 a2918a <=( a2917a ) or ( a2910a );
 a2921a <=( a1823a ) or ( a1824a );
 a2924a <=( a1821a ) or ( a1822a );
 a2925a <=( a2924a ) or ( a2921a );
 a2928a <=( a1819a ) or ( a1820a );
 a2932a <=( a1816a ) or ( a1817a );
 a2933a <=( a1818a ) or ( a2932a );
 a2934a <=( a2933a ) or ( a2928a );
 a2935a <=( a2934a ) or ( a2925a );
 a2936a <=( a2935a ) or ( a2918a );
 a2937a <=( a2936a ) or ( a2903a );
 a2940a <=( a1814a ) or ( a1815a );
 a2943a <=( a1812a ) or ( a1813a );
 a2944a <=( a2943a ) or ( a2940a );
 a2947a <=( a1810a ) or ( a1811a );
 a2950a <=( a1808a ) or ( a1809a );
 a2951a <=( a2950a ) or ( a2947a );
 a2952a <=( a2951a ) or ( a2944a );
 a2955a <=( a1806a ) or ( a1807a );
 a2958a <=( a1804a ) or ( a1805a );
 a2959a <=( a2958a ) or ( a2955a );
 a2962a <=( a1802a ) or ( a1803a );
 a2966a <=( a1799a ) or ( a1800a );
 a2967a <=( a1801a ) or ( a2966a );
 a2968a <=( a2967a ) or ( a2962a );
 a2969a <=( a2968a ) or ( a2959a );
 a2970a <=( a2969a ) or ( a2952a );
 a2973a <=( a1797a ) or ( a1798a );
 a2976a <=( a1795a ) or ( a1796a );
 a2977a <=( a2976a ) or ( a2973a );
 a2980a <=( a1793a ) or ( a1794a );
 a2984a <=( a1790a ) or ( a1791a );
 a2985a <=( a1792a ) or ( a2984a );
 a2986a <=( a2985a ) or ( a2980a );
 a2987a <=( a2986a ) or ( a2977a );
 a2990a <=( a1788a ) or ( a1789a );
 a2993a <=( a1786a ) or ( a1787a );
 a2994a <=( a2993a ) or ( a2990a );
 a2997a <=( a1784a ) or ( a1785a );
 a3001a <=( a1781a ) or ( a1782a );
 a3002a <=( a1783a ) or ( a3001a );
 a3003a <=( a3002a ) or ( a2997a );
 a3004a <=( a3003a ) or ( a2994a );
 a3005a <=( a3004a ) or ( a2987a );
 a3006a <=( a3005a ) or ( a2970a );
 a3007a <=( a3006a ) or ( a2937a );
 a3008a <=( a3007a ) or ( a2870a );
 a3011a <=( a1779a ) or ( a1780a );
 a3014a <=( a1777a ) or ( a1778a );
 a3015a <=( a3014a ) or ( a3011a );
 a3018a <=( a1775a ) or ( a1776a );
 a3021a <=( a1773a ) or ( a1774a );
 a3022a <=( a3021a ) or ( a3018a );
 a3023a <=( a3022a ) or ( a3015a );
 a3026a <=( a1771a ) or ( a1772a );
 a3029a <=( a1769a ) or ( a1770a );
 a3030a <=( a3029a ) or ( a3026a );
 a3033a <=( a1767a ) or ( a1768a );
 a3037a <=( a1764a ) or ( a1765a );
 a3038a <=( a1766a ) or ( a3037a );
 a3039a <=( a3038a ) or ( a3033a );
 a3040a <=( a3039a ) or ( a3030a );
 a3041a <=( a3040a ) or ( a3023a );
 a3044a <=( a1762a ) or ( a1763a );
 a3047a <=( a1760a ) or ( a1761a );
 a3048a <=( a3047a ) or ( a3044a );
 a3051a <=( a1758a ) or ( a1759a );
 a3054a <=( a1756a ) or ( a1757a );
 a3055a <=( a3054a ) or ( a3051a );
 a3056a <=( a3055a ) or ( a3048a );
 a3059a <=( a1754a ) or ( a1755a );
 a3062a <=( a1752a ) or ( a1753a );
 a3063a <=( a3062a ) or ( a3059a );
 a3066a <=( a1750a ) or ( a1751a );
 a3070a <=( a1747a ) or ( a1748a );
 a3071a <=( a1749a ) or ( a3070a );
 a3072a <=( a3071a ) or ( a3066a );
 a3073a <=( a3072a ) or ( a3063a );
 a3074a <=( a3073a ) or ( a3056a );
 a3075a <=( a3074a ) or ( a3041a );
 a3078a <=( a1745a ) or ( a1746a );
 a3081a <=( a1743a ) or ( a1744a );
 a3082a <=( a3081a ) or ( a3078a );
 a3085a <=( a1741a ) or ( a1742a );
 a3088a <=( a1739a ) or ( a1740a );
 a3089a <=( a3088a ) or ( a3085a );
 a3090a <=( a3089a ) or ( a3082a );
 a3093a <=( a1737a ) or ( a1738a );
 a3096a <=( a1735a ) or ( a1736a );
 a3097a <=( a3096a ) or ( a3093a );
 a3100a <=( a1733a ) or ( a1734a );
 a3104a <=( a1730a ) or ( a1731a );
 a3105a <=( a1732a ) or ( a3104a );
 a3106a <=( a3105a ) or ( a3100a );
 a3107a <=( a3106a ) or ( a3097a );
 a3108a <=( a3107a ) or ( a3090a );
 a3111a <=( a1728a ) or ( a1729a );
 a3114a <=( a1726a ) or ( a1727a );
 a3115a <=( a3114a ) or ( a3111a );
 a3118a <=( a1724a ) or ( a1725a );
 a3121a <=( a1722a ) or ( a1723a );
 a3122a <=( a3121a ) or ( a3118a );
 a3123a <=( a3122a ) or ( a3115a );
 a3126a <=( a1720a ) or ( a1721a );
 a3129a <=( a1718a ) or ( a1719a );
 a3130a <=( a3129a ) or ( a3126a );
 a3133a <=( a1716a ) or ( a1717a );
 a3137a <=( a1713a ) or ( a1714a );
 a3138a <=( a1715a ) or ( a3137a );
 a3139a <=( a3138a ) or ( a3133a );
 a3140a <=( a3139a ) or ( a3130a );
 a3141a <=( a3140a ) or ( a3123a );
 a3142a <=( a3141a ) or ( a3108a );
 a3143a <=( a3142a ) or ( a3075a );
 a3146a <=( a1711a ) or ( a1712a );
 a3149a <=( a1709a ) or ( a1710a );
 a3150a <=( a3149a ) or ( a3146a );
 a3153a <=( a1707a ) or ( a1708a );
 a3156a <=( a1705a ) or ( a1706a );
 a3157a <=( a3156a ) or ( a3153a );
 a3158a <=( a3157a ) or ( a3150a );
 a3161a <=( a1703a ) or ( a1704a );
 a3164a <=( a1701a ) or ( a1702a );
 a3165a <=( a3164a ) or ( a3161a );
 a3168a <=( a1699a ) or ( a1700a );
 a3172a <=( a1696a ) or ( a1697a );
 a3173a <=( a1698a ) or ( a3172a );
 a3174a <=( a3173a ) or ( a3168a );
 a3175a <=( a3174a ) or ( a3165a );
 a3176a <=( a3175a ) or ( a3158a );
 a3179a <=( a1694a ) or ( a1695a );
 a3182a <=( a1692a ) or ( a1693a );
 a3183a <=( a3182a ) or ( a3179a );
 a3186a <=( a1690a ) or ( a1691a );
 a3189a <=( a1688a ) or ( a1689a );
 a3190a <=( a3189a ) or ( a3186a );
 a3191a <=( a3190a ) or ( a3183a );
 a3194a <=( a1686a ) or ( a1687a );
 a3197a <=( a1684a ) or ( a1685a );
 a3198a <=( a3197a ) or ( a3194a );
 a3201a <=( a1682a ) or ( a1683a );
 a3205a <=( a1679a ) or ( a1680a );
 a3206a <=( a1681a ) or ( a3205a );
 a3207a <=( a3206a ) or ( a3201a );
 a3208a <=( a3207a ) or ( a3198a );
 a3209a <=( a3208a ) or ( a3191a );
 a3210a <=( a3209a ) or ( a3176a );
 a3213a <=( a1677a ) or ( a1678a );
 a3216a <=( a1675a ) or ( a1676a );
 a3217a <=( a3216a ) or ( a3213a );
 a3220a <=( a1673a ) or ( a1674a );
 a3223a <=( a1671a ) or ( a1672a );
 a3224a <=( a3223a ) or ( a3220a );
 a3225a <=( a3224a ) or ( a3217a );
 a3228a <=( a1669a ) or ( a1670a );
 a3231a <=( a1667a ) or ( a1668a );
 a3232a <=( a3231a ) or ( a3228a );
 a3235a <=( a1665a ) or ( a1666a );
 a3239a <=( a1662a ) or ( a1663a );
 a3240a <=( a1664a ) or ( a3239a );
 a3241a <=( a3240a ) or ( a3235a );
 a3242a <=( a3241a ) or ( a3232a );
 a3243a <=( a3242a ) or ( a3225a );
 a3246a <=( a1660a ) or ( a1661a );
 a3249a <=( a1658a ) or ( a1659a );
 a3250a <=( a3249a ) or ( a3246a );
 a3253a <=( a1656a ) or ( a1657a );
 a3257a <=( a1653a ) or ( a1654a );
 a3258a <=( a1655a ) or ( a3257a );
 a3259a <=( a3258a ) or ( a3253a );
 a3260a <=( a3259a ) or ( a3250a );
 a3263a <=( a1651a ) or ( a1652a );
 a3266a <=( a1649a ) or ( a1650a );
 a3267a <=( a3266a ) or ( a3263a );
 a3270a <=( a1647a ) or ( a1648a );
 a3274a <=( a1644a ) or ( a1645a );
 a3275a <=( a1646a ) or ( a3274a );
 a3276a <=( a3275a ) or ( a3270a );
 a3277a <=( a3276a ) or ( a3267a );
 a3278a <=( a3277a ) or ( a3260a );
 a3279a <=( a3278a ) or ( a3243a );
 a3280a <=( a3279a ) or ( a3210a );
 a3281a <=( a3280a ) or ( a3143a );
 a3282a <=( a3281a ) or ( a3008a );
 a3283a <=( a3282a ) or ( a2735a );
 a3286a <=( a1642a ) or ( a1643a );
 a3289a <=( a1640a ) or ( a1641a );
 a3290a <=( a3289a ) or ( a3286a );
 a3293a <=( a1638a ) or ( a1639a );
 a3296a <=( a1636a ) or ( a1637a );
 a3297a <=( a3296a ) or ( a3293a );
 a3298a <=( a3297a ) or ( a3290a );
 a3301a <=( a1634a ) or ( a1635a );
 a3304a <=( a1632a ) or ( a1633a );
 a3305a <=( a3304a ) or ( a3301a );
 a3308a <=( a1630a ) or ( a1631a );
 a3312a <=( a1627a ) or ( a1628a );
 a3313a <=( a1629a ) or ( a3312a );
 a3314a <=( a3313a ) or ( a3308a );
 a3315a <=( a3314a ) or ( a3305a );
 a3316a <=( a3315a ) or ( a3298a );
 a3319a <=( a1625a ) or ( a1626a );
 a3322a <=( a1623a ) or ( a1624a );
 a3323a <=( a3322a ) or ( a3319a );
 a3326a <=( a1621a ) or ( a1622a );
 a3329a <=( a1619a ) or ( a1620a );
 a3330a <=( a3329a ) or ( a3326a );
 a3331a <=( a3330a ) or ( a3323a );
 a3334a <=( a1617a ) or ( a1618a );
 a3337a <=( a1615a ) or ( a1616a );
 a3338a <=( a3337a ) or ( a3334a );
 a3341a <=( a1613a ) or ( a1614a );
 a3345a <=( a1610a ) or ( a1611a );
 a3346a <=( a1612a ) or ( a3345a );
 a3347a <=( a3346a ) or ( a3341a );
 a3348a <=( a3347a ) or ( a3338a );
 a3349a <=( a3348a ) or ( a3331a );
 a3350a <=( a3349a ) or ( a3316a );
 a3353a <=( a1608a ) or ( a1609a );
 a3356a <=( a1606a ) or ( a1607a );
 a3357a <=( a3356a ) or ( a3353a );
 a3360a <=( a1604a ) or ( a1605a );
 a3363a <=( a1602a ) or ( a1603a );
 a3364a <=( a3363a ) or ( a3360a );
 a3365a <=( a3364a ) or ( a3357a );
 a3368a <=( a1600a ) or ( a1601a );
 a3371a <=( a1598a ) or ( a1599a );
 a3372a <=( a3371a ) or ( a3368a );
 a3375a <=( a1596a ) or ( a1597a );
 a3379a <=( a1593a ) or ( a1594a );
 a3380a <=( a1595a ) or ( a3379a );
 a3381a <=( a3380a ) or ( a3375a );
 a3382a <=( a3381a ) or ( a3372a );
 a3383a <=( a3382a ) or ( a3365a );
 a3386a <=( a1591a ) or ( a1592a );
 a3389a <=( a1589a ) or ( a1590a );
 a3390a <=( a3389a ) or ( a3386a );
 a3393a <=( a1587a ) or ( a1588a );
 a3396a <=( a1585a ) or ( a1586a );
 a3397a <=( a3396a ) or ( a3393a );
 a3398a <=( a3397a ) or ( a3390a );
 a3401a <=( a1583a ) or ( a1584a );
 a3404a <=( a1581a ) or ( a1582a );
 a3405a <=( a3404a ) or ( a3401a );
 a3408a <=( a1579a ) or ( a1580a );
 a3412a <=( a1576a ) or ( a1577a );
 a3413a <=( a1578a ) or ( a3412a );
 a3414a <=( a3413a ) or ( a3408a );
 a3415a <=( a3414a ) or ( a3405a );
 a3416a <=( a3415a ) or ( a3398a );
 a3417a <=( a3416a ) or ( a3383a );
 a3418a <=( a3417a ) or ( a3350a );
 a3421a <=( a1574a ) or ( a1575a );
 a3424a <=( a1572a ) or ( a1573a );
 a3425a <=( a3424a ) or ( a3421a );
 a3428a <=( a1570a ) or ( a1571a );
 a3431a <=( a1568a ) or ( a1569a );
 a3432a <=( a3431a ) or ( a3428a );
 a3433a <=( a3432a ) or ( a3425a );
 a3436a <=( a1566a ) or ( a1567a );
 a3439a <=( a1564a ) or ( a1565a );
 a3440a <=( a3439a ) or ( a3436a );
 a3443a <=( a1562a ) or ( a1563a );
 a3447a <=( a1559a ) or ( a1560a );
 a3448a <=( a1561a ) or ( a3447a );
 a3449a <=( a3448a ) or ( a3443a );
 a3450a <=( a3449a ) or ( a3440a );
 a3451a <=( a3450a ) or ( a3433a );
 a3454a <=( a1557a ) or ( a1558a );
 a3457a <=( a1555a ) or ( a1556a );
 a3458a <=( a3457a ) or ( a3454a );
 a3461a <=( a1553a ) or ( a1554a );
 a3464a <=( a1551a ) or ( a1552a );
 a3465a <=( a3464a ) or ( a3461a );
 a3466a <=( a3465a ) or ( a3458a );
 a3469a <=( a1549a ) or ( a1550a );
 a3472a <=( a1547a ) or ( a1548a );
 a3473a <=( a3472a ) or ( a3469a );
 a3476a <=( a1545a ) or ( a1546a );
 a3480a <=( a1542a ) or ( a1543a );
 a3481a <=( a1544a ) or ( a3480a );
 a3482a <=( a3481a ) or ( a3476a );
 a3483a <=( a3482a ) or ( a3473a );
 a3484a <=( a3483a ) or ( a3466a );
 a3485a <=( a3484a ) or ( a3451a );
 a3488a <=( a1540a ) or ( a1541a );
 a3491a <=( a1538a ) or ( a1539a );
 a3492a <=( a3491a ) or ( a3488a );
 a3495a <=( a1536a ) or ( a1537a );
 a3498a <=( a1534a ) or ( a1535a );
 a3499a <=( a3498a ) or ( a3495a );
 a3500a <=( a3499a ) or ( a3492a );
 a3503a <=( a1532a ) or ( a1533a );
 a3506a <=( a1530a ) or ( a1531a );
 a3507a <=( a3506a ) or ( a3503a );
 a3510a <=( a1528a ) or ( a1529a );
 a3514a <=( a1525a ) or ( a1526a );
 a3515a <=( a1527a ) or ( a3514a );
 a3516a <=( a3515a ) or ( a3510a );
 a3517a <=( a3516a ) or ( a3507a );
 a3518a <=( a3517a ) or ( a3500a );
 a3521a <=( a1523a ) or ( a1524a );
 a3524a <=( a1521a ) or ( a1522a );
 a3525a <=( a3524a ) or ( a3521a );
 a3528a <=( a1519a ) or ( a1520a );
 a3532a <=( a1516a ) or ( a1517a );
 a3533a <=( a1518a ) or ( a3532a );
 a3534a <=( a3533a ) or ( a3528a );
 a3535a <=( a3534a ) or ( a3525a );
 a3538a <=( a1514a ) or ( a1515a );
 a3541a <=( a1512a ) or ( a1513a );
 a3542a <=( a3541a ) or ( a3538a );
 a3545a <=( a1510a ) or ( a1511a );
 a3549a <=( a1507a ) or ( a1508a );
 a3550a <=( a1509a ) or ( a3549a );
 a3551a <=( a3550a ) or ( a3545a );
 a3552a <=( a3551a ) or ( a3542a );
 a3553a <=( a3552a ) or ( a3535a );
 a3554a <=( a3553a ) or ( a3518a );
 a3555a <=( a3554a ) or ( a3485a );
 a3556a <=( a3555a ) or ( a3418a );
 a3559a <=( a1505a ) or ( a1506a );
 a3562a <=( a1503a ) or ( a1504a );
 a3563a <=( a3562a ) or ( a3559a );
 a3566a <=( a1501a ) or ( a1502a );
 a3569a <=( a1499a ) or ( a1500a );
 a3570a <=( a3569a ) or ( a3566a );
 a3571a <=( a3570a ) or ( a3563a );
 a3574a <=( a1497a ) or ( a1498a );
 a3577a <=( a1495a ) or ( a1496a );
 a3578a <=( a3577a ) or ( a3574a );
 a3581a <=( a1493a ) or ( a1494a );
 a3585a <=( a1490a ) or ( a1491a );
 a3586a <=( a1492a ) or ( a3585a );
 a3587a <=( a3586a ) or ( a3581a );
 a3588a <=( a3587a ) or ( a3578a );
 a3589a <=( a3588a ) or ( a3571a );
 a3592a <=( a1488a ) or ( a1489a );
 a3595a <=( a1486a ) or ( a1487a );
 a3596a <=( a3595a ) or ( a3592a );
 a3599a <=( a1484a ) or ( a1485a );
 a3602a <=( a1482a ) or ( a1483a );
 a3603a <=( a3602a ) or ( a3599a );
 a3604a <=( a3603a ) or ( a3596a );
 a3607a <=( a1480a ) or ( a1481a );
 a3610a <=( a1478a ) or ( a1479a );
 a3611a <=( a3610a ) or ( a3607a );
 a3614a <=( a1476a ) or ( a1477a );
 a3618a <=( a1473a ) or ( a1474a );
 a3619a <=( a1475a ) or ( a3618a );
 a3620a <=( a3619a ) or ( a3614a );
 a3621a <=( a3620a ) or ( a3611a );
 a3622a <=( a3621a ) or ( a3604a );
 a3623a <=( a3622a ) or ( a3589a );
 a3626a <=( a1471a ) or ( a1472a );
 a3629a <=( a1469a ) or ( a1470a );
 a3630a <=( a3629a ) or ( a3626a );
 a3633a <=( a1467a ) or ( a1468a );
 a3636a <=( a1465a ) or ( a1466a );
 a3637a <=( a3636a ) or ( a3633a );
 a3638a <=( a3637a ) or ( a3630a );
 a3641a <=( a1463a ) or ( a1464a );
 a3644a <=( a1461a ) or ( a1462a );
 a3645a <=( a3644a ) or ( a3641a );
 a3648a <=( a1459a ) or ( a1460a );
 a3652a <=( a1456a ) or ( a1457a );
 a3653a <=( a1458a ) or ( a3652a );
 a3654a <=( a3653a ) or ( a3648a );
 a3655a <=( a3654a ) or ( a3645a );
 a3656a <=( a3655a ) or ( a3638a );
 a3659a <=( a1454a ) or ( a1455a );
 a3662a <=( a1452a ) or ( a1453a );
 a3663a <=( a3662a ) or ( a3659a );
 a3666a <=( a1450a ) or ( a1451a );
 a3669a <=( a1448a ) or ( a1449a );
 a3670a <=( a3669a ) or ( a3666a );
 a3671a <=( a3670a ) or ( a3663a );
 a3674a <=( a1446a ) or ( a1447a );
 a3677a <=( a1444a ) or ( a1445a );
 a3678a <=( a3677a ) or ( a3674a );
 a3681a <=( a1442a ) or ( a1443a );
 a3685a <=( a1439a ) or ( a1440a );
 a3686a <=( a1441a ) or ( a3685a );
 a3687a <=( a3686a ) or ( a3681a );
 a3688a <=( a3687a ) or ( a3678a );
 a3689a <=( a3688a ) or ( a3671a );
 a3690a <=( a3689a ) or ( a3656a );
 a3691a <=( a3690a ) or ( a3623a );
 a3694a <=( a1437a ) or ( a1438a );
 a3697a <=( a1435a ) or ( a1436a );
 a3698a <=( a3697a ) or ( a3694a );
 a3701a <=( a1433a ) or ( a1434a );
 a3704a <=( a1431a ) or ( a1432a );
 a3705a <=( a3704a ) or ( a3701a );
 a3706a <=( a3705a ) or ( a3698a );
 a3709a <=( a1429a ) or ( a1430a );
 a3712a <=( a1427a ) or ( a1428a );
 a3713a <=( a3712a ) or ( a3709a );
 a3716a <=( a1425a ) or ( a1426a );
 a3720a <=( a1422a ) or ( a1423a );
 a3721a <=( a1424a ) or ( a3720a );
 a3722a <=( a3721a ) or ( a3716a );
 a3723a <=( a3722a ) or ( a3713a );
 a3724a <=( a3723a ) or ( a3706a );
 a3727a <=( a1420a ) or ( a1421a );
 a3730a <=( a1418a ) or ( a1419a );
 a3731a <=( a3730a ) or ( a3727a );
 a3734a <=( a1416a ) or ( a1417a );
 a3737a <=( a1414a ) or ( a1415a );
 a3738a <=( a3737a ) or ( a3734a );
 a3739a <=( a3738a ) or ( a3731a );
 a3742a <=( a1412a ) or ( a1413a );
 a3745a <=( a1410a ) or ( a1411a );
 a3746a <=( a3745a ) or ( a3742a );
 a3749a <=( a1408a ) or ( a1409a );
 a3753a <=( a1405a ) or ( a1406a );
 a3754a <=( a1407a ) or ( a3753a );
 a3755a <=( a3754a ) or ( a3749a );
 a3756a <=( a3755a ) or ( a3746a );
 a3757a <=( a3756a ) or ( a3739a );
 a3758a <=( a3757a ) or ( a3724a );
 a3761a <=( a1403a ) or ( a1404a );
 a3764a <=( a1401a ) or ( a1402a );
 a3765a <=( a3764a ) or ( a3761a );
 a3768a <=( a1399a ) or ( a1400a );
 a3771a <=( a1397a ) or ( a1398a );
 a3772a <=( a3771a ) or ( a3768a );
 a3773a <=( a3772a ) or ( a3765a );
 a3776a <=( a1395a ) or ( a1396a );
 a3779a <=( a1393a ) or ( a1394a );
 a3780a <=( a3779a ) or ( a3776a );
 a3783a <=( a1391a ) or ( a1392a );
 a3787a <=( a1388a ) or ( a1389a );
 a3788a <=( a1390a ) or ( a3787a );
 a3789a <=( a3788a ) or ( a3783a );
 a3790a <=( a3789a ) or ( a3780a );
 a3791a <=( a3790a ) or ( a3773a );
 a3794a <=( a1386a ) or ( a1387a );
 a3797a <=( a1384a ) or ( a1385a );
 a3798a <=( a3797a ) or ( a3794a );
 a3801a <=( a1382a ) or ( a1383a );
 a3805a <=( a1379a ) or ( a1380a );
 a3806a <=( a1381a ) or ( a3805a );
 a3807a <=( a3806a ) or ( a3801a );
 a3808a <=( a3807a ) or ( a3798a );
 a3811a <=( a1377a ) or ( a1378a );
 a3814a <=( a1375a ) or ( a1376a );
 a3815a <=( a3814a ) or ( a3811a );
 a3818a <=( a1373a ) or ( a1374a );
 a3822a <=( a1370a ) or ( a1371a );
 a3823a <=( a1372a ) or ( a3822a );
 a3824a <=( a3823a ) or ( a3818a );
 a3825a <=( a3824a ) or ( a3815a );
 a3826a <=( a3825a ) or ( a3808a );
 a3827a <=( a3826a ) or ( a3791a );
 a3828a <=( a3827a ) or ( a3758a );
 a3829a <=( a3828a ) or ( a3691a );
 a3830a <=( a3829a ) or ( a3556a );
 a3833a <=( a1368a ) or ( a1369a );
 a3836a <=( a1366a ) or ( a1367a );
 a3837a <=( a3836a ) or ( a3833a );
 a3840a <=( a1364a ) or ( a1365a );
 a3843a <=( a1362a ) or ( a1363a );
 a3844a <=( a3843a ) or ( a3840a );
 a3845a <=( a3844a ) or ( a3837a );
 a3848a <=( a1360a ) or ( a1361a );
 a3851a <=( a1358a ) or ( a1359a );
 a3852a <=( a3851a ) or ( a3848a );
 a3855a <=( a1356a ) or ( a1357a );
 a3859a <=( a1353a ) or ( a1354a );
 a3860a <=( a1355a ) or ( a3859a );
 a3861a <=( a3860a ) or ( a3855a );
 a3862a <=( a3861a ) or ( a3852a );
 a3863a <=( a3862a ) or ( a3845a );
 a3866a <=( a1351a ) or ( a1352a );
 a3869a <=( a1349a ) or ( a1350a );
 a3870a <=( a3869a ) or ( a3866a );
 a3873a <=( a1347a ) or ( a1348a );
 a3876a <=( a1345a ) or ( a1346a );
 a3877a <=( a3876a ) or ( a3873a );
 a3878a <=( a3877a ) or ( a3870a );
 a3881a <=( a1343a ) or ( a1344a );
 a3884a <=( a1341a ) or ( a1342a );
 a3885a <=( a3884a ) or ( a3881a );
 a3888a <=( a1339a ) or ( a1340a );
 a3892a <=( a1336a ) or ( a1337a );
 a3893a <=( a1338a ) or ( a3892a );
 a3894a <=( a3893a ) or ( a3888a );
 a3895a <=( a3894a ) or ( a3885a );
 a3896a <=( a3895a ) or ( a3878a );
 a3897a <=( a3896a ) or ( a3863a );
 a3900a <=( a1334a ) or ( a1335a );
 a3903a <=( a1332a ) or ( a1333a );
 a3904a <=( a3903a ) or ( a3900a );
 a3907a <=( a1330a ) or ( a1331a );
 a3910a <=( a1328a ) or ( a1329a );
 a3911a <=( a3910a ) or ( a3907a );
 a3912a <=( a3911a ) or ( a3904a );
 a3915a <=( a1326a ) or ( a1327a );
 a3918a <=( a1324a ) or ( a1325a );
 a3919a <=( a3918a ) or ( a3915a );
 a3922a <=( a1322a ) or ( a1323a );
 a3926a <=( a1319a ) or ( a1320a );
 a3927a <=( a1321a ) or ( a3926a );
 a3928a <=( a3927a ) or ( a3922a );
 a3929a <=( a3928a ) or ( a3919a );
 a3930a <=( a3929a ) or ( a3912a );
 a3933a <=( a1317a ) or ( a1318a );
 a3936a <=( a1315a ) or ( a1316a );
 a3937a <=( a3936a ) or ( a3933a );
 a3940a <=( a1313a ) or ( a1314a );
 a3943a <=( a1311a ) or ( a1312a );
 a3944a <=( a3943a ) or ( a3940a );
 a3945a <=( a3944a ) or ( a3937a );
 a3948a <=( a1309a ) or ( a1310a );
 a3951a <=( a1307a ) or ( a1308a );
 a3952a <=( a3951a ) or ( a3948a );
 a3955a <=( a1305a ) or ( a1306a );
 a3959a <=( a1302a ) or ( a1303a );
 a3960a <=( a1304a ) or ( a3959a );
 a3961a <=( a3960a ) or ( a3955a );
 a3962a <=( a3961a ) or ( a3952a );
 a3963a <=( a3962a ) or ( a3945a );
 a3964a <=( a3963a ) or ( a3930a );
 a3965a <=( a3964a ) or ( a3897a );
 a3968a <=( a1300a ) or ( a1301a );
 a3971a <=( a1298a ) or ( a1299a );
 a3972a <=( a3971a ) or ( a3968a );
 a3975a <=( a1296a ) or ( a1297a );
 a3978a <=( a1294a ) or ( a1295a );
 a3979a <=( a3978a ) or ( a3975a );
 a3980a <=( a3979a ) or ( a3972a );
 a3983a <=( a1292a ) or ( a1293a );
 a3986a <=( a1290a ) or ( a1291a );
 a3987a <=( a3986a ) or ( a3983a );
 a3990a <=( a1288a ) or ( a1289a );
 a3994a <=( a1285a ) or ( a1286a );
 a3995a <=( a1287a ) or ( a3994a );
 a3996a <=( a3995a ) or ( a3990a );
 a3997a <=( a3996a ) or ( a3987a );
 a3998a <=( a3997a ) or ( a3980a );
 a4001a <=( a1283a ) or ( a1284a );
 a4004a <=( a1281a ) or ( a1282a );
 a4005a <=( a4004a ) or ( a4001a );
 a4008a <=( a1279a ) or ( a1280a );
 a4011a <=( a1277a ) or ( a1278a );
 a4012a <=( a4011a ) or ( a4008a );
 a4013a <=( a4012a ) or ( a4005a );
 a4016a <=( a1275a ) or ( a1276a );
 a4019a <=( a1273a ) or ( a1274a );
 a4020a <=( a4019a ) or ( a4016a );
 a4023a <=( a1271a ) or ( a1272a );
 a4027a <=( a1268a ) or ( a1269a );
 a4028a <=( a1270a ) or ( a4027a );
 a4029a <=( a4028a ) or ( a4023a );
 a4030a <=( a4029a ) or ( a4020a );
 a4031a <=( a4030a ) or ( a4013a );
 a4032a <=( a4031a ) or ( a3998a );
 a4035a <=( a1266a ) or ( a1267a );
 a4038a <=( a1264a ) or ( a1265a );
 a4039a <=( a4038a ) or ( a4035a );
 a4042a <=( a1262a ) or ( a1263a );
 a4045a <=( a1260a ) or ( a1261a );
 a4046a <=( a4045a ) or ( a4042a );
 a4047a <=( a4046a ) or ( a4039a );
 a4050a <=( a1258a ) or ( a1259a );
 a4053a <=( a1256a ) or ( a1257a );
 a4054a <=( a4053a ) or ( a4050a );
 a4057a <=( a1254a ) or ( a1255a );
 a4061a <=( a1251a ) or ( a1252a );
 a4062a <=( a1253a ) or ( a4061a );
 a4063a <=( a4062a ) or ( a4057a );
 a4064a <=( a4063a ) or ( a4054a );
 a4065a <=( a4064a ) or ( a4047a );
 a4068a <=( a1249a ) or ( a1250a );
 a4071a <=( a1247a ) or ( a1248a );
 a4072a <=( a4071a ) or ( a4068a );
 a4075a <=( a1245a ) or ( a1246a );
 a4079a <=( a1242a ) or ( a1243a );
 a4080a <=( a1244a ) or ( a4079a );
 a4081a <=( a4080a ) or ( a4075a );
 a4082a <=( a4081a ) or ( a4072a );
 a4085a <=( a1240a ) or ( a1241a );
 a4088a <=( a1238a ) or ( a1239a );
 a4089a <=( a4088a ) or ( a4085a );
 a4092a <=( a1236a ) or ( a1237a );
 a4096a <=( a1233a ) or ( a1234a );
 a4097a <=( a1235a ) or ( a4096a );
 a4098a <=( a4097a ) or ( a4092a );
 a4099a <=( a4098a ) or ( a4089a );
 a4100a <=( a4099a ) or ( a4082a );
 a4101a <=( a4100a ) or ( a4065a );
 a4102a <=( a4101a ) or ( a4032a );
 a4103a <=( a4102a ) or ( a3965a );
 a4106a <=( a1231a ) or ( a1232a );
 a4109a <=( a1229a ) or ( a1230a );
 a4110a <=( a4109a ) or ( a4106a );
 a4113a <=( a1227a ) or ( a1228a );
 a4116a <=( a1225a ) or ( a1226a );
 a4117a <=( a4116a ) or ( a4113a );
 a4118a <=( a4117a ) or ( a4110a );
 a4121a <=( a1223a ) or ( a1224a );
 a4124a <=( a1221a ) or ( a1222a );
 a4125a <=( a4124a ) or ( a4121a );
 a4128a <=( a1219a ) or ( a1220a );
 a4132a <=( a1216a ) or ( a1217a );
 a4133a <=( a1218a ) or ( a4132a );
 a4134a <=( a4133a ) or ( a4128a );
 a4135a <=( a4134a ) or ( a4125a );
 a4136a <=( a4135a ) or ( a4118a );
 a4139a <=( a1214a ) or ( a1215a );
 a4142a <=( a1212a ) or ( a1213a );
 a4143a <=( a4142a ) or ( a4139a );
 a4146a <=( a1210a ) or ( a1211a );
 a4149a <=( a1208a ) or ( a1209a );
 a4150a <=( a4149a ) or ( a4146a );
 a4151a <=( a4150a ) or ( a4143a );
 a4154a <=( a1206a ) or ( a1207a );
 a4157a <=( a1204a ) or ( a1205a );
 a4158a <=( a4157a ) or ( a4154a );
 a4161a <=( a1202a ) or ( a1203a );
 a4165a <=( a1199a ) or ( a1200a );
 a4166a <=( a1201a ) or ( a4165a );
 a4167a <=( a4166a ) or ( a4161a );
 a4168a <=( a4167a ) or ( a4158a );
 a4169a <=( a4168a ) or ( a4151a );
 a4170a <=( a4169a ) or ( a4136a );
 a4173a <=( a1197a ) or ( a1198a );
 a4176a <=( a1195a ) or ( a1196a );
 a4177a <=( a4176a ) or ( a4173a );
 a4180a <=( a1193a ) or ( a1194a );
 a4183a <=( a1191a ) or ( a1192a );
 a4184a <=( a4183a ) or ( a4180a );
 a4185a <=( a4184a ) or ( a4177a );
 a4188a <=( a1189a ) or ( a1190a );
 a4191a <=( a1187a ) or ( a1188a );
 a4192a <=( a4191a ) or ( a4188a );
 a4195a <=( a1185a ) or ( a1186a );
 a4199a <=( a1182a ) or ( a1183a );
 a4200a <=( a1184a ) or ( a4199a );
 a4201a <=( a4200a ) or ( a4195a );
 a4202a <=( a4201a ) or ( a4192a );
 a4203a <=( a4202a ) or ( a4185a );
 a4206a <=( a1180a ) or ( a1181a );
 a4209a <=( a1178a ) or ( a1179a );
 a4210a <=( a4209a ) or ( a4206a );
 a4213a <=( a1176a ) or ( a1177a );
 a4216a <=( a1174a ) or ( a1175a );
 a4217a <=( a4216a ) or ( a4213a );
 a4218a <=( a4217a ) or ( a4210a );
 a4221a <=( a1172a ) or ( a1173a );
 a4224a <=( a1170a ) or ( a1171a );
 a4225a <=( a4224a ) or ( a4221a );
 a4228a <=( a1168a ) or ( a1169a );
 a4232a <=( a1165a ) or ( a1166a );
 a4233a <=( a1167a ) or ( a4232a );
 a4234a <=( a4233a ) or ( a4228a );
 a4235a <=( a4234a ) or ( a4225a );
 a4236a <=( a4235a ) or ( a4218a );
 a4237a <=( a4236a ) or ( a4203a );
 a4238a <=( a4237a ) or ( a4170a );
 a4241a <=( a1163a ) or ( a1164a );
 a4244a <=( a1161a ) or ( a1162a );
 a4245a <=( a4244a ) or ( a4241a );
 a4248a <=( a1159a ) or ( a1160a );
 a4251a <=( a1157a ) or ( a1158a );
 a4252a <=( a4251a ) or ( a4248a );
 a4253a <=( a4252a ) or ( a4245a );
 a4256a <=( a1155a ) or ( a1156a );
 a4259a <=( a1153a ) or ( a1154a );
 a4260a <=( a4259a ) or ( a4256a );
 a4263a <=( a1151a ) or ( a1152a );
 a4267a <=( a1148a ) or ( a1149a );
 a4268a <=( a1150a ) or ( a4267a );
 a4269a <=( a4268a ) or ( a4263a );
 a4270a <=( a4269a ) or ( a4260a );
 a4271a <=( a4270a ) or ( a4253a );
 a4274a <=( a1146a ) or ( a1147a );
 a4277a <=( a1144a ) or ( a1145a );
 a4278a <=( a4277a ) or ( a4274a );
 a4281a <=( a1142a ) or ( a1143a );
 a4284a <=( a1140a ) or ( a1141a );
 a4285a <=( a4284a ) or ( a4281a );
 a4286a <=( a4285a ) or ( a4278a );
 a4289a <=( a1138a ) or ( a1139a );
 a4292a <=( a1136a ) or ( a1137a );
 a4293a <=( a4292a ) or ( a4289a );
 a4296a <=( a1134a ) or ( a1135a );
 a4300a <=( a1131a ) or ( a1132a );
 a4301a <=( a1133a ) or ( a4300a );
 a4302a <=( a4301a ) or ( a4296a );
 a4303a <=( a4302a ) or ( a4293a );
 a4304a <=( a4303a ) or ( a4286a );
 a4305a <=( a4304a ) or ( a4271a );
 a4308a <=( a1129a ) or ( a1130a );
 a4311a <=( a1127a ) or ( a1128a );
 a4312a <=( a4311a ) or ( a4308a );
 a4315a <=( a1125a ) or ( a1126a );
 a4318a <=( a1123a ) or ( a1124a );
 a4319a <=( a4318a ) or ( a4315a );
 a4320a <=( a4319a ) or ( a4312a );
 a4323a <=( a1121a ) or ( a1122a );
 a4326a <=( a1119a ) or ( a1120a );
 a4327a <=( a4326a ) or ( a4323a );
 a4330a <=( a1117a ) or ( a1118a );
 a4334a <=( a1114a ) or ( a1115a );
 a4335a <=( a1116a ) or ( a4334a );
 a4336a <=( a4335a ) or ( a4330a );
 a4337a <=( a4336a ) or ( a4327a );
 a4338a <=( a4337a ) or ( a4320a );
 a4341a <=( a1112a ) or ( a1113a );
 a4344a <=( a1110a ) or ( a1111a );
 a4345a <=( a4344a ) or ( a4341a );
 a4348a <=( a1108a ) or ( a1109a );
 a4352a <=( a1105a ) or ( a1106a );
 a4353a <=( a1107a ) or ( a4352a );
 a4354a <=( a4353a ) or ( a4348a );
 a4355a <=( a4354a ) or ( a4345a );
 a4358a <=( a1103a ) or ( a1104a );
 a4361a <=( a1101a ) or ( a1102a );
 a4362a <=( a4361a ) or ( a4358a );
 a4365a <=( a1099a ) or ( a1100a );
 a4369a <=( a1096a ) or ( a1097a );
 a4370a <=( a1098a ) or ( a4369a );
 a4371a <=( a4370a ) or ( a4365a );
 a4372a <=( a4371a ) or ( a4362a );
 a4373a <=( a4372a ) or ( a4355a );
 a4374a <=( a4373a ) or ( a4338a );
 a4375a <=( a4374a ) or ( a4305a );
 a4376a <=( a4375a ) or ( a4238a );
 a4377a <=( a4376a ) or ( a4103a );
 a4378a <=( a4377a ) or ( a3830a );
 a4379a <=( a4378a ) or ( a3283a );
 a4382a <=( a1094a ) or ( a1095a );
 a4385a <=( a1092a ) or ( a1093a );
 a4386a <=( a4385a ) or ( a4382a );
 a4389a <=( a1090a ) or ( a1091a );
 a4392a <=( a1088a ) or ( a1089a );
 a4393a <=( a4392a ) or ( a4389a );
 a4394a <=( a4393a ) or ( a4386a );
 a4397a <=( a1086a ) or ( a1087a );
 a4400a <=( a1084a ) or ( a1085a );
 a4401a <=( a4400a ) or ( a4397a );
 a4404a <=( a1082a ) or ( a1083a );
 a4408a <=( a1079a ) or ( a1080a );
 a4409a <=( a1081a ) or ( a4408a );
 a4410a <=( a4409a ) or ( a4404a );
 a4411a <=( a4410a ) or ( a4401a );
 a4412a <=( a4411a ) or ( a4394a );
 a4415a <=( a1077a ) or ( a1078a );
 a4418a <=( a1075a ) or ( a1076a );
 a4419a <=( a4418a ) or ( a4415a );
 a4422a <=( a1073a ) or ( a1074a );
 a4425a <=( a1071a ) or ( a1072a );
 a4426a <=( a4425a ) or ( a4422a );
 a4427a <=( a4426a ) or ( a4419a );
 a4430a <=( a1069a ) or ( a1070a );
 a4433a <=( a1067a ) or ( a1068a );
 a4434a <=( a4433a ) or ( a4430a );
 a4437a <=( a1065a ) or ( a1066a );
 a4441a <=( a1062a ) or ( a1063a );
 a4442a <=( a1064a ) or ( a4441a );
 a4443a <=( a4442a ) or ( a4437a );
 a4444a <=( a4443a ) or ( a4434a );
 a4445a <=( a4444a ) or ( a4427a );
 a4446a <=( a4445a ) or ( a4412a );
 a4449a <=( a1060a ) or ( a1061a );
 a4452a <=( a1058a ) or ( a1059a );
 a4453a <=( a4452a ) or ( a4449a );
 a4456a <=( a1056a ) or ( a1057a );
 a4459a <=( a1054a ) or ( a1055a );
 a4460a <=( a4459a ) or ( a4456a );
 a4461a <=( a4460a ) or ( a4453a );
 a4464a <=( a1052a ) or ( a1053a );
 a4467a <=( a1050a ) or ( a1051a );
 a4468a <=( a4467a ) or ( a4464a );
 a4471a <=( a1048a ) or ( a1049a );
 a4475a <=( a1045a ) or ( a1046a );
 a4476a <=( a1047a ) or ( a4475a );
 a4477a <=( a4476a ) or ( a4471a );
 a4478a <=( a4477a ) or ( a4468a );
 a4479a <=( a4478a ) or ( a4461a );
 a4482a <=( a1043a ) or ( a1044a );
 a4485a <=( a1041a ) or ( a1042a );
 a4486a <=( a4485a ) or ( a4482a );
 a4489a <=( a1039a ) or ( a1040a );
 a4492a <=( a1037a ) or ( a1038a );
 a4493a <=( a4492a ) or ( a4489a );
 a4494a <=( a4493a ) or ( a4486a );
 a4497a <=( a1035a ) or ( a1036a );
 a4500a <=( a1033a ) or ( a1034a );
 a4501a <=( a4500a ) or ( a4497a );
 a4504a <=( a1031a ) or ( a1032a );
 a4508a <=( a1028a ) or ( a1029a );
 a4509a <=( a1030a ) or ( a4508a );
 a4510a <=( a4509a ) or ( a4504a );
 a4511a <=( a4510a ) or ( a4501a );
 a4512a <=( a4511a ) or ( a4494a );
 a4513a <=( a4512a ) or ( a4479a );
 a4514a <=( a4513a ) or ( a4446a );
 a4517a <=( a1026a ) or ( a1027a );
 a4520a <=( a1024a ) or ( a1025a );
 a4521a <=( a4520a ) or ( a4517a );
 a4524a <=( a1022a ) or ( a1023a );
 a4527a <=( a1020a ) or ( a1021a );
 a4528a <=( a4527a ) or ( a4524a );
 a4529a <=( a4528a ) or ( a4521a );
 a4532a <=( a1018a ) or ( a1019a );
 a4535a <=( a1016a ) or ( a1017a );
 a4536a <=( a4535a ) or ( a4532a );
 a4539a <=( a1014a ) or ( a1015a );
 a4543a <=( a1011a ) or ( a1012a );
 a4544a <=( a1013a ) or ( a4543a );
 a4545a <=( a4544a ) or ( a4539a );
 a4546a <=( a4545a ) or ( a4536a );
 a4547a <=( a4546a ) or ( a4529a );
 a4550a <=( a1009a ) or ( a1010a );
 a4553a <=( a1007a ) or ( a1008a );
 a4554a <=( a4553a ) or ( a4550a );
 a4557a <=( a1005a ) or ( a1006a );
 a4560a <=( a1003a ) or ( a1004a );
 a4561a <=( a4560a ) or ( a4557a );
 a4562a <=( a4561a ) or ( a4554a );
 a4565a <=( a1001a ) or ( a1002a );
 a4568a <=( a999a ) or ( a1000a );
 a4569a <=( a4568a ) or ( a4565a );
 a4572a <=( a997a ) or ( a998a );
 a4576a <=( a994a ) or ( a995a );
 a4577a <=( a996a ) or ( a4576a );
 a4578a <=( a4577a ) or ( a4572a );
 a4579a <=( a4578a ) or ( a4569a );
 a4580a <=( a4579a ) or ( a4562a );
 a4581a <=( a4580a ) or ( a4547a );
 a4584a <=( a992a ) or ( a993a );
 a4587a <=( a990a ) or ( a991a );
 a4588a <=( a4587a ) or ( a4584a );
 a4591a <=( a988a ) or ( a989a );
 a4594a <=( a986a ) or ( a987a );
 a4595a <=( a4594a ) or ( a4591a );
 a4596a <=( a4595a ) or ( a4588a );
 a4599a <=( a984a ) or ( a985a );
 a4602a <=( a982a ) or ( a983a );
 a4603a <=( a4602a ) or ( a4599a );
 a4606a <=( a980a ) or ( a981a );
 a4610a <=( a977a ) or ( a978a );
 a4611a <=( a979a ) or ( a4610a );
 a4612a <=( a4611a ) or ( a4606a );
 a4613a <=( a4612a ) or ( a4603a );
 a4614a <=( a4613a ) or ( a4596a );
 a4617a <=( a975a ) or ( a976a );
 a4620a <=( a973a ) or ( a974a );
 a4621a <=( a4620a ) or ( a4617a );
 a4624a <=( a971a ) or ( a972a );
 a4627a <=( a969a ) or ( a970a );
 a4628a <=( a4627a ) or ( a4624a );
 a4629a <=( a4628a ) or ( a4621a );
 a4632a <=( a967a ) or ( a968a );
 a4635a <=( a965a ) or ( a966a );
 a4636a <=( a4635a ) or ( a4632a );
 a4639a <=( a963a ) or ( a964a );
 a4643a <=( a960a ) or ( a961a );
 a4644a <=( a962a ) or ( a4643a );
 a4645a <=( a4644a ) or ( a4639a );
 a4646a <=( a4645a ) or ( a4636a );
 a4647a <=( a4646a ) or ( a4629a );
 a4648a <=( a4647a ) or ( a4614a );
 a4649a <=( a4648a ) or ( a4581a );
 a4650a <=( a4649a ) or ( a4514a );
 a4653a <=( a958a ) or ( a959a );
 a4656a <=( a956a ) or ( a957a );
 a4657a <=( a4656a ) or ( a4653a );
 a4660a <=( a954a ) or ( a955a );
 a4663a <=( a952a ) or ( a953a );
 a4664a <=( a4663a ) or ( a4660a );
 a4665a <=( a4664a ) or ( a4657a );
 a4668a <=( a950a ) or ( a951a );
 a4671a <=( a948a ) or ( a949a );
 a4672a <=( a4671a ) or ( a4668a );
 a4675a <=( a946a ) or ( a947a );
 a4679a <=( a943a ) or ( a944a );
 a4680a <=( a945a ) or ( a4679a );
 a4681a <=( a4680a ) or ( a4675a );
 a4682a <=( a4681a ) or ( a4672a );
 a4683a <=( a4682a ) or ( a4665a );
 a4686a <=( a941a ) or ( a942a );
 a4689a <=( a939a ) or ( a940a );
 a4690a <=( a4689a ) or ( a4686a );
 a4693a <=( a937a ) or ( a938a );
 a4696a <=( a935a ) or ( a936a );
 a4697a <=( a4696a ) or ( a4693a );
 a4698a <=( a4697a ) or ( a4690a );
 a4701a <=( a933a ) or ( a934a );
 a4704a <=( a931a ) or ( a932a );
 a4705a <=( a4704a ) or ( a4701a );
 a4708a <=( a929a ) or ( a930a );
 a4712a <=( a926a ) or ( a927a );
 a4713a <=( a928a ) or ( a4712a );
 a4714a <=( a4713a ) or ( a4708a );
 a4715a <=( a4714a ) or ( a4705a );
 a4716a <=( a4715a ) or ( a4698a );
 a4717a <=( a4716a ) or ( a4683a );
 a4720a <=( a924a ) or ( a925a );
 a4723a <=( a922a ) or ( a923a );
 a4724a <=( a4723a ) or ( a4720a );
 a4727a <=( a920a ) or ( a921a );
 a4730a <=( a918a ) or ( a919a );
 a4731a <=( a4730a ) or ( a4727a );
 a4732a <=( a4731a ) or ( a4724a );
 a4735a <=( a916a ) or ( a917a );
 a4738a <=( a914a ) or ( a915a );
 a4739a <=( a4738a ) or ( a4735a );
 a4742a <=( a912a ) or ( a913a );
 a4746a <=( a909a ) or ( a910a );
 a4747a <=( a911a ) or ( a4746a );
 a4748a <=( a4747a ) or ( a4742a );
 a4749a <=( a4748a ) or ( a4739a );
 a4750a <=( a4749a ) or ( a4732a );
 a4753a <=( a907a ) or ( a908a );
 a4756a <=( a905a ) or ( a906a );
 a4757a <=( a4756a ) or ( a4753a );
 a4760a <=( a903a ) or ( a904a );
 a4763a <=( a901a ) or ( a902a );
 a4764a <=( a4763a ) or ( a4760a );
 a4765a <=( a4764a ) or ( a4757a );
 a4768a <=( a899a ) or ( a900a );
 a4771a <=( a897a ) or ( a898a );
 a4772a <=( a4771a ) or ( a4768a );
 a4775a <=( a895a ) or ( a896a );
 a4779a <=( a892a ) or ( a893a );
 a4780a <=( a894a ) or ( a4779a );
 a4781a <=( a4780a ) or ( a4775a );
 a4782a <=( a4781a ) or ( a4772a );
 a4783a <=( a4782a ) or ( a4765a );
 a4784a <=( a4783a ) or ( a4750a );
 a4785a <=( a4784a ) or ( a4717a );
 a4788a <=( a890a ) or ( a891a );
 a4791a <=( a888a ) or ( a889a );
 a4792a <=( a4791a ) or ( a4788a );
 a4795a <=( a886a ) or ( a887a );
 a4798a <=( a884a ) or ( a885a );
 a4799a <=( a4798a ) or ( a4795a );
 a4800a <=( a4799a ) or ( a4792a );
 a4803a <=( a882a ) or ( a883a );
 a4806a <=( a880a ) or ( a881a );
 a4807a <=( a4806a ) or ( a4803a );
 a4810a <=( a878a ) or ( a879a );
 a4814a <=( a875a ) or ( a876a );
 a4815a <=( a877a ) or ( a4814a );
 a4816a <=( a4815a ) or ( a4810a );
 a4817a <=( a4816a ) or ( a4807a );
 a4818a <=( a4817a ) or ( a4800a );
 a4821a <=( a873a ) or ( a874a );
 a4824a <=( a871a ) or ( a872a );
 a4825a <=( a4824a ) or ( a4821a );
 a4828a <=( a869a ) or ( a870a );
 a4831a <=( a867a ) or ( a868a );
 a4832a <=( a4831a ) or ( a4828a );
 a4833a <=( a4832a ) or ( a4825a );
 a4836a <=( a865a ) or ( a866a );
 a4839a <=( a863a ) or ( a864a );
 a4840a <=( a4839a ) or ( a4836a );
 a4843a <=( a861a ) or ( a862a );
 a4847a <=( a858a ) or ( a859a );
 a4848a <=( a860a ) or ( a4847a );
 a4849a <=( a4848a ) or ( a4843a );
 a4850a <=( a4849a ) or ( a4840a );
 a4851a <=( a4850a ) or ( a4833a );
 a4852a <=( a4851a ) or ( a4818a );
 a4855a <=( a856a ) or ( a857a );
 a4858a <=( a854a ) or ( a855a );
 a4859a <=( a4858a ) or ( a4855a );
 a4862a <=( a852a ) or ( a853a );
 a4865a <=( a850a ) or ( a851a );
 a4866a <=( a4865a ) or ( a4862a );
 a4867a <=( a4866a ) or ( a4859a );
 a4870a <=( a848a ) or ( a849a );
 a4873a <=( a846a ) or ( a847a );
 a4874a <=( a4873a ) or ( a4870a );
 a4877a <=( a844a ) or ( a845a );
 a4881a <=( a841a ) or ( a842a );
 a4882a <=( a843a ) or ( a4881a );
 a4883a <=( a4882a ) or ( a4877a );
 a4884a <=( a4883a ) or ( a4874a );
 a4885a <=( a4884a ) or ( a4867a );
 a4888a <=( a839a ) or ( a840a );
 a4891a <=( a837a ) or ( a838a );
 a4892a <=( a4891a ) or ( a4888a );
 a4895a <=( a835a ) or ( a836a );
 a4899a <=( a832a ) or ( a833a );
 a4900a <=( a834a ) or ( a4899a );
 a4901a <=( a4900a ) or ( a4895a );
 a4902a <=( a4901a ) or ( a4892a );
 a4905a <=( a830a ) or ( a831a );
 a4908a <=( a828a ) or ( a829a );
 a4909a <=( a4908a ) or ( a4905a );
 a4912a <=( a826a ) or ( a827a );
 a4916a <=( a823a ) or ( a824a );
 a4917a <=( a825a ) or ( a4916a );
 a4918a <=( a4917a ) or ( a4912a );
 a4919a <=( a4918a ) or ( a4909a );
 a4920a <=( a4919a ) or ( a4902a );
 a4921a <=( a4920a ) or ( a4885a );
 a4922a <=( a4921a ) or ( a4852a );
 a4923a <=( a4922a ) or ( a4785a );
 a4924a <=( a4923a ) or ( a4650a );
 a4927a <=( a821a ) or ( a822a );
 a4930a <=( a819a ) or ( a820a );
 a4931a <=( a4930a ) or ( a4927a );
 a4934a <=( a817a ) or ( a818a );
 a4937a <=( a815a ) or ( a816a );
 a4938a <=( a4937a ) or ( a4934a );
 a4939a <=( a4938a ) or ( a4931a );
 a4942a <=( a813a ) or ( a814a );
 a4945a <=( a811a ) or ( a812a );
 a4946a <=( a4945a ) or ( a4942a );
 a4949a <=( a809a ) or ( a810a );
 a4953a <=( a806a ) or ( a807a );
 a4954a <=( a808a ) or ( a4953a );
 a4955a <=( a4954a ) or ( a4949a );
 a4956a <=( a4955a ) or ( a4946a );
 a4957a <=( a4956a ) or ( a4939a );
 a4960a <=( a804a ) or ( a805a );
 a4963a <=( a802a ) or ( a803a );
 a4964a <=( a4963a ) or ( a4960a );
 a4967a <=( a800a ) or ( a801a );
 a4970a <=( a798a ) or ( a799a );
 a4971a <=( a4970a ) or ( a4967a );
 a4972a <=( a4971a ) or ( a4964a );
 a4975a <=( a796a ) or ( a797a );
 a4978a <=( a794a ) or ( a795a );
 a4979a <=( a4978a ) or ( a4975a );
 a4982a <=( a792a ) or ( a793a );
 a4986a <=( a789a ) or ( a790a );
 a4987a <=( a791a ) or ( a4986a );
 a4988a <=( a4987a ) or ( a4982a );
 a4989a <=( a4988a ) or ( a4979a );
 a4990a <=( a4989a ) or ( a4972a );
 a4991a <=( a4990a ) or ( a4957a );
 a4994a <=( a787a ) or ( a788a );
 a4997a <=( a785a ) or ( a786a );
 a4998a <=( a4997a ) or ( a4994a );
 a5001a <=( a783a ) or ( a784a );
 a5004a <=( a781a ) or ( a782a );
 a5005a <=( a5004a ) or ( a5001a );
 a5006a <=( a5005a ) or ( a4998a );
 a5009a <=( a779a ) or ( a780a );
 a5012a <=( a777a ) or ( a778a );
 a5013a <=( a5012a ) or ( a5009a );
 a5016a <=( a775a ) or ( a776a );
 a5020a <=( a772a ) or ( a773a );
 a5021a <=( a774a ) or ( a5020a );
 a5022a <=( a5021a ) or ( a5016a );
 a5023a <=( a5022a ) or ( a5013a );
 a5024a <=( a5023a ) or ( a5006a );
 a5027a <=( a770a ) or ( a771a );
 a5030a <=( a768a ) or ( a769a );
 a5031a <=( a5030a ) or ( a5027a );
 a5034a <=( a766a ) or ( a767a );
 a5037a <=( a764a ) or ( a765a );
 a5038a <=( a5037a ) or ( a5034a );
 a5039a <=( a5038a ) or ( a5031a );
 a5042a <=( a762a ) or ( a763a );
 a5045a <=( a760a ) or ( a761a );
 a5046a <=( a5045a ) or ( a5042a );
 a5049a <=( a758a ) or ( a759a );
 a5053a <=( a755a ) or ( a756a );
 a5054a <=( a757a ) or ( a5053a );
 a5055a <=( a5054a ) or ( a5049a );
 a5056a <=( a5055a ) or ( a5046a );
 a5057a <=( a5056a ) or ( a5039a );
 a5058a <=( a5057a ) or ( a5024a );
 a5059a <=( a5058a ) or ( a4991a );
 a5062a <=( a753a ) or ( a754a );
 a5065a <=( a751a ) or ( a752a );
 a5066a <=( a5065a ) or ( a5062a );
 a5069a <=( a749a ) or ( a750a );
 a5072a <=( a747a ) or ( a748a );
 a5073a <=( a5072a ) or ( a5069a );
 a5074a <=( a5073a ) or ( a5066a );
 a5077a <=( a745a ) or ( a746a );
 a5080a <=( a743a ) or ( a744a );
 a5081a <=( a5080a ) or ( a5077a );
 a5084a <=( a741a ) or ( a742a );
 a5088a <=( a738a ) or ( a739a );
 a5089a <=( a740a ) or ( a5088a );
 a5090a <=( a5089a ) or ( a5084a );
 a5091a <=( a5090a ) or ( a5081a );
 a5092a <=( a5091a ) or ( a5074a );
 a5095a <=( a736a ) or ( a737a );
 a5098a <=( a734a ) or ( a735a );
 a5099a <=( a5098a ) or ( a5095a );
 a5102a <=( a732a ) or ( a733a );
 a5105a <=( a730a ) or ( a731a );
 a5106a <=( a5105a ) or ( a5102a );
 a5107a <=( a5106a ) or ( a5099a );
 a5110a <=( a728a ) or ( a729a );
 a5113a <=( a726a ) or ( a727a );
 a5114a <=( a5113a ) or ( a5110a );
 a5117a <=( a724a ) or ( a725a );
 a5121a <=( a721a ) or ( a722a );
 a5122a <=( a723a ) or ( a5121a );
 a5123a <=( a5122a ) or ( a5117a );
 a5124a <=( a5123a ) or ( a5114a );
 a5125a <=( a5124a ) or ( a5107a );
 a5126a <=( a5125a ) or ( a5092a );
 a5129a <=( a719a ) or ( a720a );
 a5132a <=( a717a ) or ( a718a );
 a5133a <=( a5132a ) or ( a5129a );
 a5136a <=( a715a ) or ( a716a );
 a5139a <=( a713a ) or ( a714a );
 a5140a <=( a5139a ) or ( a5136a );
 a5141a <=( a5140a ) or ( a5133a );
 a5144a <=( a711a ) or ( a712a );
 a5147a <=( a709a ) or ( a710a );
 a5148a <=( a5147a ) or ( a5144a );
 a5151a <=( a707a ) or ( a708a );
 a5155a <=( a704a ) or ( a705a );
 a5156a <=( a706a ) or ( a5155a );
 a5157a <=( a5156a ) or ( a5151a );
 a5158a <=( a5157a ) or ( a5148a );
 a5159a <=( a5158a ) or ( a5141a );
 a5162a <=( a702a ) or ( a703a );
 a5165a <=( a700a ) or ( a701a );
 a5166a <=( a5165a ) or ( a5162a );
 a5169a <=( a698a ) or ( a699a );
 a5173a <=( a695a ) or ( a696a );
 a5174a <=( a697a ) or ( a5173a );
 a5175a <=( a5174a ) or ( a5169a );
 a5176a <=( a5175a ) or ( a5166a );
 a5179a <=( a693a ) or ( a694a );
 a5182a <=( a691a ) or ( a692a );
 a5183a <=( a5182a ) or ( a5179a );
 a5186a <=( a689a ) or ( a690a );
 a5190a <=( a686a ) or ( a687a );
 a5191a <=( a688a ) or ( a5190a );
 a5192a <=( a5191a ) or ( a5186a );
 a5193a <=( a5192a ) or ( a5183a );
 a5194a <=( a5193a ) or ( a5176a );
 a5195a <=( a5194a ) or ( a5159a );
 a5196a <=( a5195a ) or ( a5126a );
 a5197a <=( a5196a ) or ( a5059a );
 a5200a <=( a684a ) or ( a685a );
 a5203a <=( a682a ) or ( a683a );
 a5204a <=( a5203a ) or ( a5200a );
 a5207a <=( a680a ) or ( a681a );
 a5210a <=( a678a ) or ( a679a );
 a5211a <=( a5210a ) or ( a5207a );
 a5212a <=( a5211a ) or ( a5204a );
 a5215a <=( a676a ) or ( a677a );
 a5218a <=( a674a ) or ( a675a );
 a5219a <=( a5218a ) or ( a5215a );
 a5222a <=( a672a ) or ( a673a );
 a5226a <=( a669a ) or ( a670a );
 a5227a <=( a671a ) or ( a5226a );
 a5228a <=( a5227a ) or ( a5222a );
 a5229a <=( a5228a ) or ( a5219a );
 a5230a <=( a5229a ) or ( a5212a );
 a5233a <=( a667a ) or ( a668a );
 a5236a <=( a665a ) or ( a666a );
 a5237a <=( a5236a ) or ( a5233a );
 a5240a <=( a663a ) or ( a664a );
 a5243a <=( a661a ) or ( a662a );
 a5244a <=( a5243a ) or ( a5240a );
 a5245a <=( a5244a ) or ( a5237a );
 a5248a <=( a659a ) or ( a660a );
 a5251a <=( a657a ) or ( a658a );
 a5252a <=( a5251a ) or ( a5248a );
 a5255a <=( a655a ) or ( a656a );
 a5259a <=( a652a ) or ( a653a );
 a5260a <=( a654a ) or ( a5259a );
 a5261a <=( a5260a ) or ( a5255a );
 a5262a <=( a5261a ) or ( a5252a );
 a5263a <=( a5262a ) or ( a5245a );
 a5264a <=( a5263a ) or ( a5230a );
 a5267a <=( a650a ) or ( a651a );
 a5270a <=( a648a ) or ( a649a );
 a5271a <=( a5270a ) or ( a5267a );
 a5274a <=( a646a ) or ( a647a );
 a5277a <=( a644a ) or ( a645a );
 a5278a <=( a5277a ) or ( a5274a );
 a5279a <=( a5278a ) or ( a5271a );
 a5282a <=( a642a ) or ( a643a );
 a5285a <=( a640a ) or ( a641a );
 a5286a <=( a5285a ) or ( a5282a );
 a5289a <=( a638a ) or ( a639a );
 a5293a <=( a635a ) or ( a636a );
 a5294a <=( a637a ) or ( a5293a );
 a5295a <=( a5294a ) or ( a5289a );
 a5296a <=( a5295a ) or ( a5286a );
 a5297a <=( a5296a ) or ( a5279a );
 a5300a <=( a633a ) or ( a634a );
 a5303a <=( a631a ) or ( a632a );
 a5304a <=( a5303a ) or ( a5300a );
 a5307a <=( a629a ) or ( a630a );
 a5310a <=( a627a ) or ( a628a );
 a5311a <=( a5310a ) or ( a5307a );
 a5312a <=( a5311a ) or ( a5304a );
 a5315a <=( a625a ) or ( a626a );
 a5318a <=( a623a ) or ( a624a );
 a5319a <=( a5318a ) or ( a5315a );
 a5322a <=( a621a ) or ( a622a );
 a5326a <=( a618a ) or ( a619a );
 a5327a <=( a620a ) or ( a5326a );
 a5328a <=( a5327a ) or ( a5322a );
 a5329a <=( a5328a ) or ( a5319a );
 a5330a <=( a5329a ) or ( a5312a );
 a5331a <=( a5330a ) or ( a5297a );
 a5332a <=( a5331a ) or ( a5264a );
 a5335a <=( a616a ) or ( a617a );
 a5338a <=( a614a ) or ( a615a );
 a5339a <=( a5338a ) or ( a5335a );
 a5342a <=( a612a ) or ( a613a );
 a5345a <=( a610a ) or ( a611a );
 a5346a <=( a5345a ) or ( a5342a );
 a5347a <=( a5346a ) or ( a5339a );
 a5350a <=( a608a ) or ( a609a );
 a5353a <=( a606a ) or ( a607a );
 a5354a <=( a5353a ) or ( a5350a );
 a5357a <=( a604a ) or ( a605a );
 a5361a <=( a601a ) or ( a602a );
 a5362a <=( a603a ) or ( a5361a );
 a5363a <=( a5362a ) or ( a5357a );
 a5364a <=( a5363a ) or ( a5354a );
 a5365a <=( a5364a ) or ( a5347a );
 a5368a <=( a599a ) or ( a600a );
 a5371a <=( a597a ) or ( a598a );
 a5372a <=( a5371a ) or ( a5368a );
 a5375a <=( a595a ) or ( a596a );
 a5378a <=( a593a ) or ( a594a );
 a5379a <=( a5378a ) or ( a5375a );
 a5380a <=( a5379a ) or ( a5372a );
 a5383a <=( a591a ) or ( a592a );
 a5386a <=( a589a ) or ( a590a );
 a5387a <=( a5386a ) or ( a5383a );
 a5390a <=( a587a ) or ( a588a );
 a5394a <=( a584a ) or ( a585a );
 a5395a <=( a586a ) or ( a5394a );
 a5396a <=( a5395a ) or ( a5390a );
 a5397a <=( a5396a ) or ( a5387a );
 a5398a <=( a5397a ) or ( a5380a );
 a5399a <=( a5398a ) or ( a5365a );
 a5402a <=( a582a ) or ( a583a );
 a5405a <=( a580a ) or ( a581a );
 a5406a <=( a5405a ) or ( a5402a );
 a5409a <=( a578a ) or ( a579a );
 a5412a <=( a576a ) or ( a577a );
 a5413a <=( a5412a ) or ( a5409a );
 a5414a <=( a5413a ) or ( a5406a );
 a5417a <=( a574a ) or ( a575a );
 a5420a <=( a572a ) or ( a573a );
 a5421a <=( a5420a ) or ( a5417a );
 a5424a <=( a570a ) or ( a571a );
 a5428a <=( a567a ) or ( a568a );
 a5429a <=( a569a ) or ( a5428a );
 a5430a <=( a5429a ) or ( a5424a );
 a5431a <=( a5430a ) or ( a5421a );
 a5432a <=( a5431a ) or ( a5414a );
 a5435a <=( a565a ) or ( a566a );
 a5438a <=( a563a ) or ( a564a );
 a5439a <=( a5438a ) or ( a5435a );
 a5442a <=( a561a ) or ( a562a );
 a5446a <=( a558a ) or ( a559a );
 a5447a <=( a560a ) or ( a5446a );
 a5448a <=( a5447a ) or ( a5442a );
 a5449a <=( a5448a ) or ( a5439a );
 a5452a <=( a556a ) or ( a557a );
 a5455a <=( a554a ) or ( a555a );
 a5456a <=( a5455a ) or ( a5452a );
 a5459a <=( a552a ) or ( a553a );
 a5463a <=( a549a ) or ( a550a );
 a5464a <=( a551a ) or ( a5463a );
 a5465a <=( a5464a ) or ( a5459a );
 a5466a <=( a5465a ) or ( a5456a );
 a5467a <=( a5466a ) or ( a5449a );
 a5468a <=( a5467a ) or ( a5432a );
 a5469a <=( a5468a ) or ( a5399a );
 a5470a <=( a5469a ) or ( a5332a );
 a5471a <=( a5470a ) or ( a5197a );
 a5472a <=( a5471a ) or ( a4924a );
 a5475a <=( a547a ) or ( a548a );
 a5478a <=( a545a ) or ( a546a );
 a5479a <=( a5478a ) or ( a5475a );
 a5482a <=( a543a ) or ( a544a );
 a5485a <=( a541a ) or ( a542a );
 a5486a <=( a5485a ) or ( a5482a );
 a5487a <=( a5486a ) or ( a5479a );
 a5490a <=( a539a ) or ( a540a );
 a5493a <=( a537a ) or ( a538a );
 a5494a <=( a5493a ) or ( a5490a );
 a5497a <=( a535a ) or ( a536a );
 a5501a <=( a532a ) or ( a533a );
 a5502a <=( a534a ) or ( a5501a );
 a5503a <=( a5502a ) or ( a5497a );
 a5504a <=( a5503a ) or ( a5494a );
 a5505a <=( a5504a ) or ( a5487a );
 a5508a <=( a530a ) or ( a531a );
 a5511a <=( a528a ) or ( a529a );
 a5512a <=( a5511a ) or ( a5508a );
 a5515a <=( a526a ) or ( a527a );
 a5518a <=( a524a ) or ( a525a );
 a5519a <=( a5518a ) or ( a5515a );
 a5520a <=( a5519a ) or ( a5512a );
 a5523a <=( a522a ) or ( a523a );
 a5526a <=( a520a ) or ( a521a );
 a5527a <=( a5526a ) or ( a5523a );
 a5530a <=( a518a ) or ( a519a );
 a5534a <=( a515a ) or ( a516a );
 a5535a <=( a517a ) or ( a5534a );
 a5536a <=( a5535a ) or ( a5530a );
 a5537a <=( a5536a ) or ( a5527a );
 a5538a <=( a5537a ) or ( a5520a );
 a5539a <=( a5538a ) or ( a5505a );
 a5542a <=( a513a ) or ( a514a );
 a5545a <=( a511a ) or ( a512a );
 a5546a <=( a5545a ) or ( a5542a );
 a5549a <=( a509a ) or ( a510a );
 a5552a <=( a507a ) or ( a508a );
 a5553a <=( a5552a ) or ( a5549a );
 a5554a <=( a5553a ) or ( a5546a );
 a5557a <=( a505a ) or ( a506a );
 a5560a <=( a503a ) or ( a504a );
 a5561a <=( a5560a ) or ( a5557a );
 a5564a <=( a501a ) or ( a502a );
 a5568a <=( a498a ) or ( a499a );
 a5569a <=( a500a ) or ( a5568a );
 a5570a <=( a5569a ) or ( a5564a );
 a5571a <=( a5570a ) or ( a5561a );
 a5572a <=( a5571a ) or ( a5554a );
 a5575a <=( a496a ) or ( a497a );
 a5578a <=( a494a ) or ( a495a );
 a5579a <=( a5578a ) or ( a5575a );
 a5582a <=( a492a ) or ( a493a );
 a5585a <=( a490a ) or ( a491a );
 a5586a <=( a5585a ) or ( a5582a );
 a5587a <=( a5586a ) or ( a5579a );
 a5590a <=( a488a ) or ( a489a );
 a5593a <=( a486a ) or ( a487a );
 a5594a <=( a5593a ) or ( a5590a );
 a5597a <=( a484a ) or ( a485a );
 a5601a <=( a481a ) or ( a482a );
 a5602a <=( a483a ) or ( a5601a );
 a5603a <=( a5602a ) or ( a5597a );
 a5604a <=( a5603a ) or ( a5594a );
 a5605a <=( a5604a ) or ( a5587a );
 a5606a <=( a5605a ) or ( a5572a );
 a5607a <=( a5606a ) or ( a5539a );
 a5610a <=( a479a ) or ( a480a );
 a5613a <=( a477a ) or ( a478a );
 a5614a <=( a5613a ) or ( a5610a );
 a5617a <=( a475a ) or ( a476a );
 a5620a <=( a473a ) or ( a474a );
 a5621a <=( a5620a ) or ( a5617a );
 a5622a <=( a5621a ) or ( a5614a );
 a5625a <=( a471a ) or ( a472a );
 a5628a <=( a469a ) or ( a470a );
 a5629a <=( a5628a ) or ( a5625a );
 a5632a <=( a467a ) or ( a468a );
 a5636a <=( a464a ) or ( a465a );
 a5637a <=( a466a ) or ( a5636a );
 a5638a <=( a5637a ) or ( a5632a );
 a5639a <=( a5638a ) or ( a5629a );
 a5640a <=( a5639a ) or ( a5622a );
 a5643a <=( a462a ) or ( a463a );
 a5646a <=( a460a ) or ( a461a );
 a5647a <=( a5646a ) or ( a5643a );
 a5650a <=( a458a ) or ( a459a );
 a5653a <=( a456a ) or ( a457a );
 a5654a <=( a5653a ) or ( a5650a );
 a5655a <=( a5654a ) or ( a5647a );
 a5658a <=( a454a ) or ( a455a );
 a5661a <=( a452a ) or ( a453a );
 a5662a <=( a5661a ) or ( a5658a );
 a5665a <=( a450a ) or ( a451a );
 a5669a <=( a447a ) or ( a448a );
 a5670a <=( a449a ) or ( a5669a );
 a5671a <=( a5670a ) or ( a5665a );
 a5672a <=( a5671a ) or ( a5662a );
 a5673a <=( a5672a ) or ( a5655a );
 a5674a <=( a5673a ) or ( a5640a );
 a5677a <=( a445a ) or ( a446a );
 a5680a <=( a443a ) or ( a444a );
 a5681a <=( a5680a ) or ( a5677a );
 a5684a <=( a441a ) or ( a442a );
 a5687a <=( a439a ) or ( a440a );
 a5688a <=( a5687a ) or ( a5684a );
 a5689a <=( a5688a ) or ( a5681a );
 a5692a <=( a437a ) or ( a438a );
 a5695a <=( a435a ) or ( a436a );
 a5696a <=( a5695a ) or ( a5692a );
 a5699a <=( a433a ) or ( a434a );
 a5703a <=( a430a ) or ( a431a );
 a5704a <=( a432a ) or ( a5703a );
 a5705a <=( a5704a ) or ( a5699a );
 a5706a <=( a5705a ) or ( a5696a );
 a5707a <=( a5706a ) or ( a5689a );
 a5710a <=( a428a ) or ( a429a );
 a5713a <=( a426a ) or ( a427a );
 a5714a <=( a5713a ) or ( a5710a );
 a5717a <=( a424a ) or ( a425a );
 a5721a <=( a421a ) or ( a422a );
 a5722a <=( a423a ) or ( a5721a );
 a5723a <=( a5722a ) or ( a5717a );
 a5724a <=( a5723a ) or ( a5714a );
 a5727a <=( a419a ) or ( a420a );
 a5730a <=( a417a ) or ( a418a );
 a5731a <=( a5730a ) or ( a5727a );
 a5734a <=( a415a ) or ( a416a );
 a5738a <=( a412a ) or ( a413a );
 a5739a <=( a414a ) or ( a5738a );
 a5740a <=( a5739a ) or ( a5734a );
 a5741a <=( a5740a ) or ( a5731a );
 a5742a <=( a5741a ) or ( a5724a );
 a5743a <=( a5742a ) or ( a5707a );
 a5744a <=( a5743a ) or ( a5674a );
 a5745a <=( a5744a ) or ( a5607a );
 a5748a <=( a410a ) or ( a411a );
 a5751a <=( a408a ) or ( a409a );
 a5752a <=( a5751a ) or ( a5748a );
 a5755a <=( a406a ) or ( a407a );
 a5758a <=( a404a ) or ( a405a );
 a5759a <=( a5758a ) or ( a5755a );
 a5760a <=( a5759a ) or ( a5752a );
 a5763a <=( a402a ) or ( a403a );
 a5766a <=( a400a ) or ( a401a );
 a5767a <=( a5766a ) or ( a5763a );
 a5770a <=( a398a ) or ( a399a );
 a5774a <=( a395a ) or ( a396a );
 a5775a <=( a397a ) or ( a5774a );
 a5776a <=( a5775a ) or ( a5770a );
 a5777a <=( a5776a ) or ( a5767a );
 a5778a <=( a5777a ) or ( a5760a );
 a5781a <=( a393a ) or ( a394a );
 a5784a <=( a391a ) or ( a392a );
 a5785a <=( a5784a ) or ( a5781a );
 a5788a <=( a389a ) or ( a390a );
 a5791a <=( a387a ) or ( a388a );
 a5792a <=( a5791a ) or ( a5788a );
 a5793a <=( a5792a ) or ( a5785a );
 a5796a <=( a385a ) or ( a386a );
 a5799a <=( a383a ) or ( a384a );
 a5800a <=( a5799a ) or ( a5796a );
 a5803a <=( a381a ) or ( a382a );
 a5807a <=( a378a ) or ( a379a );
 a5808a <=( a380a ) or ( a5807a );
 a5809a <=( a5808a ) or ( a5803a );
 a5810a <=( a5809a ) or ( a5800a );
 a5811a <=( a5810a ) or ( a5793a );
 a5812a <=( a5811a ) or ( a5778a );
 a5815a <=( a376a ) or ( a377a );
 a5818a <=( a374a ) or ( a375a );
 a5819a <=( a5818a ) or ( a5815a );
 a5822a <=( a372a ) or ( a373a );
 a5825a <=( a370a ) or ( a371a );
 a5826a <=( a5825a ) or ( a5822a );
 a5827a <=( a5826a ) or ( a5819a );
 a5830a <=( a368a ) or ( a369a );
 a5833a <=( a366a ) or ( a367a );
 a5834a <=( a5833a ) or ( a5830a );
 a5837a <=( a364a ) or ( a365a );
 a5841a <=( a361a ) or ( a362a );
 a5842a <=( a363a ) or ( a5841a );
 a5843a <=( a5842a ) or ( a5837a );
 a5844a <=( a5843a ) or ( a5834a );
 a5845a <=( a5844a ) or ( a5827a );
 a5848a <=( a359a ) or ( a360a );
 a5851a <=( a357a ) or ( a358a );
 a5852a <=( a5851a ) or ( a5848a );
 a5855a <=( a355a ) or ( a356a );
 a5858a <=( a353a ) or ( a354a );
 a5859a <=( a5858a ) or ( a5855a );
 a5860a <=( a5859a ) or ( a5852a );
 a5863a <=( a351a ) or ( a352a );
 a5866a <=( a349a ) or ( a350a );
 a5867a <=( a5866a ) or ( a5863a );
 a5870a <=( a347a ) or ( a348a );
 a5874a <=( a344a ) or ( a345a );
 a5875a <=( a346a ) or ( a5874a );
 a5876a <=( a5875a ) or ( a5870a );
 a5877a <=( a5876a ) or ( a5867a );
 a5878a <=( a5877a ) or ( a5860a );
 a5879a <=( a5878a ) or ( a5845a );
 a5880a <=( a5879a ) or ( a5812a );
 a5883a <=( a342a ) or ( a343a );
 a5886a <=( a340a ) or ( a341a );
 a5887a <=( a5886a ) or ( a5883a );
 a5890a <=( a338a ) or ( a339a );
 a5893a <=( a336a ) or ( a337a );
 a5894a <=( a5893a ) or ( a5890a );
 a5895a <=( a5894a ) or ( a5887a );
 a5898a <=( a334a ) or ( a335a );
 a5901a <=( a332a ) or ( a333a );
 a5902a <=( a5901a ) or ( a5898a );
 a5905a <=( a330a ) or ( a331a );
 a5909a <=( a327a ) or ( a328a );
 a5910a <=( a329a ) or ( a5909a );
 a5911a <=( a5910a ) or ( a5905a );
 a5912a <=( a5911a ) or ( a5902a );
 a5913a <=( a5912a ) or ( a5895a );
 a5916a <=( a325a ) or ( a326a );
 a5919a <=( a323a ) or ( a324a );
 a5920a <=( a5919a ) or ( a5916a );
 a5923a <=( a321a ) or ( a322a );
 a5926a <=( a319a ) or ( a320a );
 a5927a <=( a5926a ) or ( a5923a );
 a5928a <=( a5927a ) or ( a5920a );
 a5931a <=( a317a ) or ( a318a );
 a5934a <=( a315a ) or ( a316a );
 a5935a <=( a5934a ) or ( a5931a );
 a5938a <=( a313a ) or ( a314a );
 a5942a <=( a310a ) or ( a311a );
 a5943a <=( a312a ) or ( a5942a );
 a5944a <=( a5943a ) or ( a5938a );
 a5945a <=( a5944a ) or ( a5935a );
 a5946a <=( a5945a ) or ( a5928a );
 a5947a <=( a5946a ) or ( a5913a );
 a5950a <=( a308a ) or ( a309a );
 a5953a <=( a306a ) or ( a307a );
 a5954a <=( a5953a ) or ( a5950a );
 a5957a <=( a304a ) or ( a305a );
 a5960a <=( a302a ) or ( a303a );
 a5961a <=( a5960a ) or ( a5957a );
 a5962a <=( a5961a ) or ( a5954a );
 a5965a <=( a300a ) or ( a301a );
 a5968a <=( a298a ) or ( a299a );
 a5969a <=( a5968a ) or ( a5965a );
 a5972a <=( a296a ) or ( a297a );
 a5976a <=( a293a ) or ( a294a );
 a5977a <=( a295a ) or ( a5976a );
 a5978a <=( a5977a ) or ( a5972a );
 a5979a <=( a5978a ) or ( a5969a );
 a5980a <=( a5979a ) or ( a5962a );
 a5983a <=( a291a ) or ( a292a );
 a5986a <=( a289a ) or ( a290a );
 a5987a <=( a5986a ) or ( a5983a );
 a5990a <=( a287a ) or ( a288a );
 a5994a <=( a284a ) or ( a285a );
 a5995a <=( a286a ) or ( a5994a );
 a5996a <=( a5995a ) or ( a5990a );
 a5997a <=( a5996a ) or ( a5987a );
 a6000a <=( a282a ) or ( a283a );
 a6003a <=( a280a ) or ( a281a );
 a6004a <=( a6003a ) or ( a6000a );
 a6007a <=( a278a ) or ( a279a );
 a6011a <=( a275a ) or ( a276a );
 a6012a <=( a277a ) or ( a6011a );
 a6013a <=( a6012a ) or ( a6007a );
 a6014a <=( a6013a ) or ( a6004a );
 a6015a <=( a6014a ) or ( a5997a );
 a6016a <=( a6015a ) or ( a5980a );
 a6017a <=( a6016a ) or ( a5947a );
 a6018a <=( a6017a ) or ( a5880a );
 a6019a <=( a6018a ) or ( a5745a );
 a6022a <=( a273a ) or ( a274a );
 a6025a <=( a271a ) or ( a272a );
 a6026a <=( a6025a ) or ( a6022a );
 a6029a <=( a269a ) or ( a270a );
 a6032a <=( a267a ) or ( a268a );
 a6033a <=( a6032a ) or ( a6029a );
 a6034a <=( a6033a ) or ( a6026a );
 a6037a <=( a265a ) or ( a266a );
 a6040a <=( a263a ) or ( a264a );
 a6041a <=( a6040a ) or ( a6037a );
 a6044a <=( a261a ) or ( a262a );
 a6048a <=( a258a ) or ( a259a );
 a6049a <=( a260a ) or ( a6048a );
 a6050a <=( a6049a ) or ( a6044a );
 a6051a <=( a6050a ) or ( a6041a );
 a6052a <=( a6051a ) or ( a6034a );
 a6055a <=( a256a ) or ( a257a );
 a6058a <=( a254a ) or ( a255a );
 a6059a <=( a6058a ) or ( a6055a );
 a6062a <=( a252a ) or ( a253a );
 a6065a <=( a250a ) or ( a251a );
 a6066a <=( a6065a ) or ( a6062a );
 a6067a <=( a6066a ) or ( a6059a );
 a6070a <=( a248a ) or ( a249a );
 a6073a <=( a246a ) or ( a247a );
 a6074a <=( a6073a ) or ( a6070a );
 a6077a <=( a244a ) or ( a245a );
 a6081a <=( a241a ) or ( a242a );
 a6082a <=( a243a ) or ( a6081a );
 a6083a <=( a6082a ) or ( a6077a );
 a6084a <=( a6083a ) or ( a6074a );
 a6085a <=( a6084a ) or ( a6067a );
 a6086a <=( a6085a ) or ( a6052a );
 a6089a <=( a239a ) or ( a240a );
 a6092a <=( a237a ) or ( a238a );
 a6093a <=( a6092a ) or ( a6089a );
 a6096a <=( a235a ) or ( a236a );
 a6099a <=( a233a ) or ( a234a );
 a6100a <=( a6099a ) or ( a6096a );
 a6101a <=( a6100a ) or ( a6093a );
 a6104a <=( a231a ) or ( a232a );
 a6107a <=( a229a ) or ( a230a );
 a6108a <=( a6107a ) or ( a6104a );
 a6111a <=( a227a ) or ( a228a );
 a6115a <=( a224a ) or ( a225a );
 a6116a <=( a226a ) or ( a6115a );
 a6117a <=( a6116a ) or ( a6111a );
 a6118a <=( a6117a ) or ( a6108a );
 a6119a <=( a6118a ) or ( a6101a );
 a6122a <=( a222a ) or ( a223a );
 a6125a <=( a220a ) or ( a221a );
 a6126a <=( a6125a ) or ( a6122a );
 a6129a <=( a218a ) or ( a219a );
 a6132a <=( a216a ) or ( a217a );
 a6133a <=( a6132a ) or ( a6129a );
 a6134a <=( a6133a ) or ( a6126a );
 a6137a <=( a214a ) or ( a215a );
 a6140a <=( a212a ) or ( a213a );
 a6141a <=( a6140a ) or ( a6137a );
 a6144a <=( a210a ) or ( a211a );
 a6148a <=( a207a ) or ( a208a );
 a6149a <=( a209a ) or ( a6148a );
 a6150a <=( a6149a ) or ( a6144a );
 a6151a <=( a6150a ) or ( a6141a );
 a6152a <=( a6151a ) or ( a6134a );
 a6153a <=( a6152a ) or ( a6119a );
 a6154a <=( a6153a ) or ( a6086a );
 a6157a <=( a205a ) or ( a206a );
 a6160a <=( a203a ) or ( a204a );
 a6161a <=( a6160a ) or ( a6157a );
 a6164a <=( a201a ) or ( a202a );
 a6167a <=( a199a ) or ( a200a );
 a6168a <=( a6167a ) or ( a6164a );
 a6169a <=( a6168a ) or ( a6161a );
 a6172a <=( a197a ) or ( a198a );
 a6175a <=( a195a ) or ( a196a );
 a6176a <=( a6175a ) or ( a6172a );
 a6179a <=( a193a ) or ( a194a );
 a6183a <=( a190a ) or ( a191a );
 a6184a <=( a192a ) or ( a6183a );
 a6185a <=( a6184a ) or ( a6179a );
 a6186a <=( a6185a ) or ( a6176a );
 a6187a <=( a6186a ) or ( a6169a );
 a6190a <=( a188a ) or ( a189a );
 a6193a <=( a186a ) or ( a187a );
 a6194a <=( a6193a ) or ( a6190a );
 a6197a <=( a184a ) or ( a185a );
 a6200a <=( a182a ) or ( a183a );
 a6201a <=( a6200a ) or ( a6197a );
 a6202a <=( a6201a ) or ( a6194a );
 a6205a <=( a180a ) or ( a181a );
 a6208a <=( a178a ) or ( a179a );
 a6209a <=( a6208a ) or ( a6205a );
 a6212a <=( a176a ) or ( a177a );
 a6216a <=( a173a ) or ( a174a );
 a6217a <=( a175a ) or ( a6216a );
 a6218a <=( a6217a ) or ( a6212a );
 a6219a <=( a6218a ) or ( a6209a );
 a6220a <=( a6219a ) or ( a6202a );
 a6221a <=( a6220a ) or ( a6187a );
 a6224a <=( a171a ) or ( a172a );
 a6227a <=( a169a ) or ( a170a );
 a6228a <=( a6227a ) or ( a6224a );
 a6231a <=( a167a ) or ( a168a );
 a6234a <=( a165a ) or ( a166a );
 a6235a <=( a6234a ) or ( a6231a );
 a6236a <=( a6235a ) or ( a6228a );
 a6239a <=( a163a ) or ( a164a );
 a6242a <=( a161a ) or ( a162a );
 a6243a <=( a6242a ) or ( a6239a );
 a6246a <=( a159a ) or ( a160a );
 a6250a <=( a156a ) or ( a157a );
 a6251a <=( a158a ) or ( a6250a );
 a6252a <=( a6251a ) or ( a6246a );
 a6253a <=( a6252a ) or ( a6243a );
 a6254a <=( a6253a ) or ( a6236a );
 a6257a <=( a154a ) or ( a155a );
 a6260a <=( a152a ) or ( a153a );
 a6261a <=( a6260a ) or ( a6257a );
 a6264a <=( a150a ) or ( a151a );
 a6268a <=( a147a ) or ( a148a );
 a6269a <=( a149a ) or ( a6268a );
 a6270a <=( a6269a ) or ( a6264a );
 a6271a <=( a6270a ) or ( a6261a );
 a6274a <=( a145a ) or ( a146a );
 a6277a <=( a143a ) or ( a144a );
 a6278a <=( a6277a ) or ( a6274a );
 a6281a <=( a141a ) or ( a142a );
 a6285a <=( a138a ) or ( a139a );
 a6286a <=( a140a ) or ( a6285a );
 a6287a <=( a6286a ) or ( a6281a );
 a6288a <=( a6287a ) or ( a6278a );
 a6289a <=( a6288a ) or ( a6271a );
 a6290a <=( a6289a ) or ( a6254a );
 a6291a <=( a6290a ) or ( a6221a );
 a6292a <=( a6291a ) or ( a6154a );
 a6295a <=( a136a ) or ( a137a );
 a6298a <=( a134a ) or ( a135a );
 a6299a <=( a6298a ) or ( a6295a );
 a6302a <=( a132a ) or ( a133a );
 a6305a <=( a130a ) or ( a131a );
 a6306a <=( a6305a ) or ( a6302a );
 a6307a <=( a6306a ) or ( a6299a );
 a6310a <=( a128a ) or ( a129a );
 a6313a <=( a126a ) or ( a127a );
 a6314a <=( a6313a ) or ( a6310a );
 a6317a <=( a124a ) or ( a125a );
 a6321a <=( a121a ) or ( a122a );
 a6322a <=( a123a ) or ( a6321a );
 a6323a <=( a6322a ) or ( a6317a );
 a6324a <=( a6323a ) or ( a6314a );
 a6325a <=( a6324a ) or ( a6307a );
 a6328a <=( a119a ) or ( a120a );
 a6331a <=( a117a ) or ( a118a );
 a6332a <=( a6331a ) or ( a6328a );
 a6335a <=( a115a ) or ( a116a );
 a6338a <=( a113a ) or ( a114a );
 a6339a <=( a6338a ) or ( a6335a );
 a6340a <=( a6339a ) or ( a6332a );
 a6343a <=( a111a ) or ( a112a );
 a6346a <=( a109a ) or ( a110a );
 a6347a <=( a6346a ) or ( a6343a );
 a6350a <=( a107a ) or ( a108a );
 a6354a <=( a104a ) or ( a105a );
 a6355a <=( a106a ) or ( a6354a );
 a6356a <=( a6355a ) or ( a6350a );
 a6357a <=( a6356a ) or ( a6347a );
 a6358a <=( a6357a ) or ( a6340a );
 a6359a <=( a6358a ) or ( a6325a );
 a6362a <=( a102a ) or ( a103a );
 a6365a <=( a100a ) or ( a101a );
 a6366a <=( a6365a ) or ( a6362a );
 a6369a <=( a98a ) or ( a99a );
 a6372a <=( a96a ) or ( a97a );
 a6373a <=( a6372a ) or ( a6369a );
 a6374a <=( a6373a ) or ( a6366a );
 a6377a <=( a94a ) or ( a95a );
 a6380a <=( a92a ) or ( a93a );
 a6381a <=( a6380a ) or ( a6377a );
 a6384a <=( a90a ) or ( a91a );
 a6388a <=( a87a ) or ( a88a );
 a6389a <=( a89a ) or ( a6388a );
 a6390a <=( a6389a ) or ( a6384a );
 a6391a <=( a6390a ) or ( a6381a );
 a6392a <=( a6391a ) or ( a6374a );
 a6395a <=( a85a ) or ( a86a );
 a6398a <=( a83a ) or ( a84a );
 a6399a <=( a6398a ) or ( a6395a );
 a6402a <=( a81a ) or ( a82a );
 a6405a <=( a79a ) or ( a80a );
 a6406a <=( a6405a ) or ( a6402a );
 a6407a <=( a6406a ) or ( a6399a );
 a6410a <=( a77a ) or ( a78a );
 a6413a <=( a75a ) or ( a76a );
 a6414a <=( a6413a ) or ( a6410a );
 a6417a <=( a73a ) or ( a74a );
 a6421a <=( a70a ) or ( a71a );
 a6422a <=( a72a ) or ( a6421a );
 a6423a <=( a6422a ) or ( a6417a );
 a6424a <=( a6423a ) or ( a6414a );
 a6425a <=( a6424a ) or ( a6407a );
 a6426a <=( a6425a ) or ( a6392a );
 a6427a <=( a6426a ) or ( a6359a );
 a6430a <=( a68a ) or ( a69a );
 a6433a <=( a66a ) or ( a67a );
 a6434a <=( a6433a ) or ( a6430a );
 a6437a <=( a64a ) or ( a65a );
 a6440a <=( a62a ) or ( a63a );
 a6441a <=( a6440a ) or ( a6437a );
 a6442a <=( a6441a ) or ( a6434a );
 a6445a <=( a60a ) or ( a61a );
 a6448a <=( a58a ) or ( a59a );
 a6449a <=( a6448a ) or ( a6445a );
 a6452a <=( a56a ) or ( a57a );
 a6456a <=( a53a ) or ( a54a );
 a6457a <=( a55a ) or ( a6456a );
 a6458a <=( a6457a ) or ( a6452a );
 a6459a <=( a6458a ) or ( a6449a );
 a6460a <=( a6459a ) or ( a6442a );
 a6463a <=( a51a ) or ( a52a );
 a6466a <=( a49a ) or ( a50a );
 a6467a <=( a6466a ) or ( a6463a );
 a6470a <=( a47a ) or ( a48a );
 a6473a <=( a45a ) or ( a46a );
 a6474a <=( a6473a ) or ( a6470a );
 a6475a <=( a6474a ) or ( a6467a );
 a6478a <=( a43a ) or ( a44a );
 a6481a <=( a41a ) or ( a42a );
 a6482a <=( a6481a ) or ( a6478a );
 a6485a <=( a39a ) or ( a40a );
 a6489a <=( a36a ) or ( a37a );
 a6490a <=( a38a ) or ( a6489a );
 a6491a <=( a6490a ) or ( a6485a );
 a6492a <=( a6491a ) or ( a6482a );
 a6493a <=( a6492a ) or ( a6475a );
 a6494a <=( a6493a ) or ( a6460a );
 a6497a <=( a34a ) or ( a35a );
 a6500a <=( a32a ) or ( a33a );
 a6501a <=( a6500a ) or ( a6497a );
 a6504a <=( a30a ) or ( a31a );
 a6507a <=( a28a ) or ( a29a );
 a6508a <=( a6507a ) or ( a6504a );
 a6509a <=( a6508a ) or ( a6501a );
 a6512a <=( a26a ) or ( a27a );
 a6515a <=( a24a ) or ( a25a );
 a6516a <=( a6515a ) or ( a6512a );
 a6519a <=( a22a ) or ( a23a );
 a6523a <=( a19a ) or ( a20a );
 a6524a <=( a21a ) or ( a6523a );
 a6525a <=( a6524a ) or ( a6519a );
 a6526a <=( a6525a ) or ( a6516a );
 a6527a <=( a6526a ) or ( a6509a );
 a6530a <=( a17a ) or ( a18a );
 a6533a <=( a15a ) or ( a16a );
 a6534a <=( a6533a ) or ( a6530a );
 a6537a <=( a13a ) or ( a14a );
 a6541a <=( a10a ) or ( a11a );
 a6542a <=( a12a ) or ( a6541a );
 a6543a <=( a6542a ) or ( a6537a );
 a6544a <=( a6543a ) or ( a6534a );
 a6547a <=( a8a ) or ( a9a );
 a6550a <=( a6a ) or ( a7a );
 a6551a <=( a6550a ) or ( a6547a );
 a6554a <=( a4a ) or ( a5a );
 a6558a <=( a1a ) or ( a2a );
 a6559a <=( a3a ) or ( a6558a );
 a6560a <=( a6559a ) or ( a6554a );
 a6561a <=( a6560a ) or ( a6551a );
 a6562a <=( a6561a ) or ( a6544a );
 a6563a <=( a6562a ) or ( a6527a );
 a6564a <=( a6563a ) or ( a6494a );
 a6565a <=( a6564a ) or ( a6427a );
 a6566a <=( a6565a ) or ( a6292a );
 a6567a <=( a6566a ) or ( a6019a );
 a6568a <=( a6567a ) or ( a5472a );
 a6572a <=( (not A199)  and  A166 );
 a6573a <=( A167  and  a6572a );
 a6577a <=( A202  and  A201 );
 a6578a <=( A200  and  a6577a );
 a6582a <=( (not A199)  and  A166 );
 a6583a <=( A167  and  a6582a );
 a6587a <=( A203  and  A201 );
 a6588a <=( A200  and  a6587a );
 a6592a <=( A199  and  A166 );
 a6593a <=( A167  and  a6592a );
 a6597a <=( A202  and  A201 );
 a6598a <=( (not A200)  and  a6597a );
 a6602a <=( A199  and  A166 );
 a6603a <=( A167  and  a6602a );
 a6607a <=( A203  and  A201 );
 a6608a <=( (not A200)  and  a6607a );
 a6612a <=( (not A199)  and  (not A166) );
 a6613a <=( (not A167)  and  a6612a );
 a6617a <=( A202  and  A201 );
 a6618a <=( A200  and  a6617a );
 a6622a <=( (not A199)  and  (not A166) );
 a6623a <=( (not A167)  and  a6622a );
 a6627a <=( A203  and  A201 );
 a6628a <=( A200  and  a6627a );
 a6632a <=( A199  and  (not A166) );
 a6633a <=( (not A167)  and  a6632a );
 a6637a <=( A202  and  A201 );
 a6638a <=( (not A200)  and  a6637a );
 a6642a <=( A199  and  (not A166) );
 a6643a <=( (not A167)  and  a6642a );
 a6647a <=( A203  and  A201 );
 a6648a <=( (not A200)  and  a6647a );
 a6652a <=( (not A199)  and  (not A168) );
 a6653a <=( (not A170)  and  a6652a );
 a6657a <=( A202  and  A201 );
 a6658a <=( A200  and  a6657a );
 a6662a <=( (not A199)  and  (not A168) );
 a6663a <=( (not A170)  and  a6662a );
 a6667a <=( A203  and  A201 );
 a6668a <=( A200  and  a6667a );
 a6672a <=( A199  and  (not A168) );
 a6673a <=( (not A170)  and  a6672a );
 a6677a <=( A202  and  A201 );
 a6678a <=( (not A200)  and  a6677a );
 a6682a <=( A199  and  (not A168) );
 a6683a <=( (not A170)  and  a6682a );
 a6687a <=( A203  and  A201 );
 a6688a <=( (not A200)  and  a6687a );
 a6692a <=( (not A199)  and  (not A168) );
 a6693a <=( A169  and  a6692a );
 a6697a <=( A202  and  A201 );
 a6698a <=( A200  and  a6697a );
 a6702a <=( (not A199)  and  (not A168) );
 a6703a <=( A169  and  a6702a );
 a6707a <=( A203  and  A201 );
 a6708a <=( A200  and  a6707a );
 a6712a <=( A199  and  (not A168) );
 a6713a <=( A169  and  a6712a );
 a6717a <=( A202  and  A201 );
 a6718a <=( (not A200)  and  a6717a );
 a6722a <=( A199  and  (not A168) );
 a6723a <=( A169  and  a6722a );
 a6727a <=( A203  and  A201 );
 a6728a <=( (not A200)  and  a6727a );
 a6732a <=( (not A199)  and  A166 );
 a6733a <=( A167  and  a6732a );
 a6736a <=( (not A201)  and  A200 );
 a6739a <=( (not A203)  and  (not A202) );
 a6740a <=( a6739a  and  a6736a );
 a6744a <=( A199  and  A166 );
 a6745a <=( A167  and  a6744a );
 a6748a <=( (not A201)  and  (not A200) );
 a6751a <=( (not A203)  and  (not A202) );
 a6752a <=( a6751a  and  a6748a );
 a6756a <=( (not A199)  and  (not A166) );
 a6757a <=( (not A167)  and  a6756a );
 a6760a <=( (not A201)  and  A200 );
 a6763a <=( (not A203)  and  (not A202) );
 a6764a <=( a6763a  and  a6760a );
 a6768a <=( A199  and  (not A166) );
 a6769a <=( (not A167)  and  a6768a );
 a6772a <=( (not A201)  and  (not A200) );
 a6775a <=( (not A203)  and  (not A202) );
 a6776a <=( a6775a  and  a6772a );
 a6780a <=( (not A199)  and  (not A168) );
 a6781a <=( (not A170)  and  a6780a );
 a6784a <=( (not A201)  and  A200 );
 a6787a <=( (not A203)  and  (not A202) );
 a6788a <=( a6787a  and  a6784a );
 a6792a <=( A199  and  (not A168) );
 a6793a <=( (not A170)  and  a6792a );
 a6796a <=( (not A201)  and  (not A200) );
 a6799a <=( (not A203)  and  (not A202) );
 a6800a <=( a6799a  and  a6796a );
 a6804a <=( (not A199)  and  (not A168) );
 a6805a <=( A169  and  a6804a );
 a6808a <=( (not A201)  and  A200 );
 a6811a <=( (not A203)  and  (not A202) );
 a6812a <=( a6811a  and  a6808a );
 a6816a <=( A199  and  (not A168) );
 a6817a <=( A169  and  a6816a );
 a6820a <=( (not A201)  and  (not A200) );
 a6823a <=( (not A203)  and  (not A202) );
 a6824a <=( a6823a  and  a6820a );
 a6828a <=( A168  and  (not A169) );
 a6829a <=( A170  and  a6828a );
 a6832a <=( A200  and  (not A199) );
 a6835a <=( A202  and  A201 );
 a6836a <=( a6835a  and  a6832a );
 a6840a <=( A168  and  (not A169) );
 a6841a <=( A170  and  a6840a );
 a6844a <=( A200  and  (not A199) );
 a6847a <=( A203  and  A201 );
 a6848a <=( a6847a  and  a6844a );
 a6852a <=( A168  and  (not A169) );
 a6853a <=( A170  and  a6852a );
 a6856a <=( (not A200)  and  A199 );
 a6859a <=( A202  and  A201 );
 a6860a <=( a6859a  and  a6856a );
 a6864a <=( A168  and  (not A169) );
 a6865a <=( A170  and  a6864a );
 a6868a <=( (not A200)  and  A199 );
 a6871a <=( A203  and  A201 );
 a6872a <=( a6871a  and  a6868a );
 a6875a <=( (not A169)  and  A170 );
 a6878a <=( (not A199)  and  A168 );
 a6879a <=( a6878a  and  a6875a );
 a6882a <=( (not A201)  and  A200 );
 a6885a <=( (not A203)  and  (not A202) );
 a6886a <=( a6885a  and  a6882a );
 a6889a <=( (not A169)  and  A170 );
 a6892a <=( A199  and  A168 );
 a6893a <=( a6892a  and  a6889a );
 a6896a <=( (not A201)  and  (not A200) );
 a6899a <=( (not A203)  and  (not A202) );
 a6900a <=( a6899a  and  a6896a );
 a6904a <=( A167  and  A168 );
 a6905a <=( (not A170)  and  a6904a );
 a6908a <=( (not A201)  and  (not A166) );
 a6911a <=( (not A232)  and  A202 );
 a6912a <=( a6911a  and  a6908a );
 a6913a <=( a6912a  and  a6905a );
 a6917a <=( A235  and  A234 );
 a6918a <=( A233  and  a6917a );
 a6921a <=( (not A299)  and  A298 );
 a6924a <=( A301  and  A300 );
 a6925a <=( a6924a  and  a6921a );
 a6926a <=( a6925a  and  a6918a );
 a6930a <=( A167  and  A168 );
 a6931a <=( (not A170)  and  a6930a );
 a6934a <=( (not A201)  and  (not A166) );
 a6937a <=( (not A232)  and  A202 );
 a6938a <=( a6937a  and  a6934a );
 a6939a <=( a6938a  and  a6931a );
 a6943a <=( A235  and  A234 );
 a6944a <=( A233  and  a6943a );
 a6947a <=( (not A299)  and  A298 );
 a6950a <=( A302  and  A300 );
 a6951a <=( a6950a  and  a6947a );
 a6952a <=( a6951a  and  a6944a );
 a6956a <=( A167  and  A168 );
 a6957a <=( (not A170)  and  a6956a );
 a6960a <=( (not A201)  and  (not A166) );
 a6963a <=( (not A232)  and  A202 );
 a6964a <=( a6963a  and  a6960a );
 a6965a <=( a6964a  and  a6957a );
 a6969a <=( A235  and  A234 );
 a6970a <=( A233  and  a6969a );
 a6973a <=( A299  and  (not A298) );
 a6976a <=( A301  and  A300 );
 a6977a <=( a6976a  and  a6973a );
 a6978a <=( a6977a  and  a6970a );
 a6982a <=( A167  and  A168 );
 a6983a <=( (not A170)  and  a6982a );
 a6986a <=( (not A201)  and  (not A166) );
 a6989a <=( (not A232)  and  A202 );
 a6990a <=( a6989a  and  a6986a );
 a6991a <=( a6990a  and  a6983a );
 a6995a <=( A235  and  A234 );
 a6996a <=( A233  and  a6995a );
 a6999a <=( A299  and  (not A298) );
 a7002a <=( A302  and  A300 );
 a7003a <=( a7002a  and  a6999a );
 a7004a <=( a7003a  and  a6996a );
 a7008a <=( A167  and  A168 );
 a7009a <=( (not A170)  and  a7008a );
 a7012a <=( (not A201)  and  (not A166) );
 a7015a <=( (not A232)  and  A202 );
 a7016a <=( a7015a  and  a7012a );
 a7017a <=( a7016a  and  a7009a );
 a7021a <=( A235  and  A234 );
 a7022a <=( A233  and  a7021a );
 a7025a <=( A266  and  (not A265) );
 a7028a <=( A268  and  A267 );
 a7029a <=( a7028a  and  a7025a );
 a7030a <=( a7029a  and  a7022a );
 a7034a <=( A167  and  A168 );
 a7035a <=( (not A170)  and  a7034a );
 a7038a <=( (not A201)  and  (not A166) );
 a7041a <=( (not A232)  and  A202 );
 a7042a <=( a7041a  and  a7038a );
 a7043a <=( a7042a  and  a7035a );
 a7047a <=( A235  and  A234 );
 a7048a <=( A233  and  a7047a );
 a7051a <=( A266  and  (not A265) );
 a7054a <=( A269  and  A267 );
 a7055a <=( a7054a  and  a7051a );
 a7056a <=( a7055a  and  a7048a );
 a7060a <=( A167  and  A168 );
 a7061a <=( (not A170)  and  a7060a );
 a7064a <=( (not A201)  and  (not A166) );
 a7067a <=( (not A232)  and  A202 );
 a7068a <=( a7067a  and  a7064a );
 a7069a <=( a7068a  and  a7061a );
 a7073a <=( A235  and  A234 );
 a7074a <=( A233  and  a7073a );
 a7077a <=( (not A266)  and  A265 );
 a7080a <=( A268  and  A267 );
 a7081a <=( a7080a  and  a7077a );
 a7082a <=( a7081a  and  a7074a );
 a7086a <=( A167  and  A168 );
 a7087a <=( (not A170)  and  a7086a );
 a7090a <=( (not A201)  and  (not A166) );
 a7093a <=( (not A232)  and  A202 );
 a7094a <=( a7093a  and  a7090a );
 a7095a <=( a7094a  and  a7087a );
 a7099a <=( A235  and  A234 );
 a7100a <=( A233  and  a7099a );
 a7103a <=( (not A266)  and  A265 );
 a7106a <=( A269  and  A267 );
 a7107a <=( a7106a  and  a7103a );
 a7108a <=( a7107a  and  a7100a );
 a7112a <=( A167  and  A168 );
 a7113a <=( (not A170)  and  a7112a );
 a7116a <=( (not A201)  and  (not A166) );
 a7119a <=( (not A232)  and  A202 );
 a7120a <=( a7119a  and  a7116a );
 a7121a <=( a7120a  and  a7113a );
 a7125a <=( A236  and  A234 );
 a7126a <=( A233  and  a7125a );
 a7129a <=( (not A299)  and  A298 );
 a7132a <=( A301  and  A300 );
 a7133a <=( a7132a  and  a7129a );
 a7134a <=( a7133a  and  a7126a );
 a7138a <=( A167  and  A168 );
 a7139a <=( (not A170)  and  a7138a );
 a7142a <=( (not A201)  and  (not A166) );
 a7145a <=( (not A232)  and  A202 );
 a7146a <=( a7145a  and  a7142a );
 a7147a <=( a7146a  and  a7139a );
 a7151a <=( A236  and  A234 );
 a7152a <=( A233  and  a7151a );
 a7155a <=( (not A299)  and  A298 );
 a7158a <=( A302  and  A300 );
 a7159a <=( a7158a  and  a7155a );
 a7160a <=( a7159a  and  a7152a );
 a7164a <=( A167  and  A168 );
 a7165a <=( (not A170)  and  a7164a );
 a7168a <=( (not A201)  and  (not A166) );
 a7171a <=( (not A232)  and  A202 );
 a7172a <=( a7171a  and  a7168a );
 a7173a <=( a7172a  and  a7165a );
 a7177a <=( A236  and  A234 );
 a7178a <=( A233  and  a7177a );
 a7181a <=( A299  and  (not A298) );
 a7184a <=( A301  and  A300 );
 a7185a <=( a7184a  and  a7181a );
 a7186a <=( a7185a  and  a7178a );
 a7190a <=( A167  and  A168 );
 a7191a <=( (not A170)  and  a7190a );
 a7194a <=( (not A201)  and  (not A166) );
 a7197a <=( (not A232)  and  A202 );
 a7198a <=( a7197a  and  a7194a );
 a7199a <=( a7198a  and  a7191a );
 a7203a <=( A236  and  A234 );
 a7204a <=( A233  and  a7203a );
 a7207a <=( A299  and  (not A298) );
 a7210a <=( A302  and  A300 );
 a7211a <=( a7210a  and  a7207a );
 a7212a <=( a7211a  and  a7204a );
 a7216a <=( A167  and  A168 );
 a7217a <=( (not A170)  and  a7216a );
 a7220a <=( (not A201)  and  (not A166) );
 a7223a <=( (not A232)  and  A202 );
 a7224a <=( a7223a  and  a7220a );
 a7225a <=( a7224a  and  a7217a );
 a7229a <=( A236  and  A234 );
 a7230a <=( A233  and  a7229a );
 a7233a <=( A266  and  (not A265) );
 a7236a <=( A268  and  A267 );
 a7237a <=( a7236a  and  a7233a );
 a7238a <=( a7237a  and  a7230a );
 a7242a <=( A167  and  A168 );
 a7243a <=( (not A170)  and  a7242a );
 a7246a <=( (not A201)  and  (not A166) );
 a7249a <=( (not A232)  and  A202 );
 a7250a <=( a7249a  and  a7246a );
 a7251a <=( a7250a  and  a7243a );
 a7255a <=( A236  and  A234 );
 a7256a <=( A233  and  a7255a );
 a7259a <=( A266  and  (not A265) );
 a7262a <=( A269  and  A267 );
 a7263a <=( a7262a  and  a7259a );
 a7264a <=( a7263a  and  a7256a );
 a7268a <=( A167  and  A168 );
 a7269a <=( (not A170)  and  a7268a );
 a7272a <=( (not A201)  and  (not A166) );
 a7275a <=( (not A232)  and  A202 );
 a7276a <=( a7275a  and  a7272a );
 a7277a <=( a7276a  and  a7269a );
 a7281a <=( A236  and  A234 );
 a7282a <=( A233  and  a7281a );
 a7285a <=( (not A266)  and  A265 );
 a7288a <=( A268  and  A267 );
 a7289a <=( a7288a  and  a7285a );
 a7290a <=( a7289a  and  a7282a );
 a7294a <=( A167  and  A168 );
 a7295a <=( (not A170)  and  a7294a );
 a7298a <=( (not A201)  and  (not A166) );
 a7301a <=( (not A232)  and  A202 );
 a7302a <=( a7301a  and  a7298a );
 a7303a <=( a7302a  and  a7295a );
 a7307a <=( A236  and  A234 );
 a7308a <=( A233  and  a7307a );
 a7311a <=( (not A266)  and  A265 );
 a7314a <=( A269  and  A267 );
 a7315a <=( a7314a  and  a7311a );
 a7316a <=( a7315a  and  a7308a );
 a7320a <=( A167  and  A168 );
 a7321a <=( (not A170)  and  a7320a );
 a7324a <=( (not A201)  and  (not A166) );
 a7327a <=( A232  and  A202 );
 a7328a <=( a7327a  and  a7324a );
 a7329a <=( a7328a  and  a7321a );
 a7333a <=( A235  and  A234 );
 a7334a <=( (not A233)  and  a7333a );
 a7337a <=( (not A299)  and  A298 );
 a7340a <=( A301  and  A300 );
 a7341a <=( a7340a  and  a7337a );
 a7342a <=( a7341a  and  a7334a );
 a7346a <=( A167  and  A168 );
 a7347a <=( (not A170)  and  a7346a );
 a7350a <=( (not A201)  and  (not A166) );
 a7353a <=( A232  and  A202 );
 a7354a <=( a7353a  and  a7350a );
 a7355a <=( a7354a  and  a7347a );
 a7359a <=( A235  and  A234 );
 a7360a <=( (not A233)  and  a7359a );
 a7363a <=( (not A299)  and  A298 );
 a7366a <=( A302  and  A300 );
 a7367a <=( a7366a  and  a7363a );
 a7368a <=( a7367a  and  a7360a );
 a7372a <=( A167  and  A168 );
 a7373a <=( (not A170)  and  a7372a );
 a7376a <=( (not A201)  and  (not A166) );
 a7379a <=( A232  and  A202 );
 a7380a <=( a7379a  and  a7376a );
 a7381a <=( a7380a  and  a7373a );
 a7385a <=( A235  and  A234 );
 a7386a <=( (not A233)  and  a7385a );
 a7389a <=( A299  and  (not A298) );
 a7392a <=( A301  and  A300 );
 a7393a <=( a7392a  and  a7389a );
 a7394a <=( a7393a  and  a7386a );
 a7398a <=( A167  and  A168 );
 a7399a <=( (not A170)  and  a7398a );
 a7402a <=( (not A201)  and  (not A166) );
 a7405a <=( A232  and  A202 );
 a7406a <=( a7405a  and  a7402a );
 a7407a <=( a7406a  and  a7399a );
 a7411a <=( A235  and  A234 );
 a7412a <=( (not A233)  and  a7411a );
 a7415a <=( A299  and  (not A298) );
 a7418a <=( A302  and  A300 );
 a7419a <=( a7418a  and  a7415a );
 a7420a <=( a7419a  and  a7412a );
 a7424a <=( A167  and  A168 );
 a7425a <=( (not A170)  and  a7424a );
 a7428a <=( (not A201)  and  (not A166) );
 a7431a <=( A232  and  A202 );
 a7432a <=( a7431a  and  a7428a );
 a7433a <=( a7432a  and  a7425a );
 a7437a <=( A235  and  A234 );
 a7438a <=( (not A233)  and  a7437a );
 a7441a <=( A266  and  (not A265) );
 a7444a <=( A268  and  A267 );
 a7445a <=( a7444a  and  a7441a );
 a7446a <=( a7445a  and  a7438a );
 a7450a <=( A167  and  A168 );
 a7451a <=( (not A170)  and  a7450a );
 a7454a <=( (not A201)  and  (not A166) );
 a7457a <=( A232  and  A202 );
 a7458a <=( a7457a  and  a7454a );
 a7459a <=( a7458a  and  a7451a );
 a7463a <=( A235  and  A234 );
 a7464a <=( (not A233)  and  a7463a );
 a7467a <=( A266  and  (not A265) );
 a7470a <=( A269  and  A267 );
 a7471a <=( a7470a  and  a7467a );
 a7472a <=( a7471a  and  a7464a );
 a7476a <=( A167  and  A168 );
 a7477a <=( (not A170)  and  a7476a );
 a7480a <=( (not A201)  and  (not A166) );
 a7483a <=( A232  and  A202 );
 a7484a <=( a7483a  and  a7480a );
 a7485a <=( a7484a  and  a7477a );
 a7489a <=( A235  and  A234 );
 a7490a <=( (not A233)  and  a7489a );
 a7493a <=( (not A266)  and  A265 );
 a7496a <=( A268  and  A267 );
 a7497a <=( a7496a  and  a7493a );
 a7498a <=( a7497a  and  a7490a );
 a7502a <=( A167  and  A168 );
 a7503a <=( (not A170)  and  a7502a );
 a7506a <=( (not A201)  and  (not A166) );
 a7509a <=( A232  and  A202 );
 a7510a <=( a7509a  and  a7506a );
 a7511a <=( a7510a  and  a7503a );
 a7515a <=( A235  and  A234 );
 a7516a <=( (not A233)  and  a7515a );
 a7519a <=( (not A266)  and  A265 );
 a7522a <=( A269  and  A267 );
 a7523a <=( a7522a  and  a7519a );
 a7524a <=( a7523a  and  a7516a );
 a7528a <=( A167  and  A168 );
 a7529a <=( (not A170)  and  a7528a );
 a7532a <=( (not A201)  and  (not A166) );
 a7535a <=( A232  and  A202 );
 a7536a <=( a7535a  and  a7532a );
 a7537a <=( a7536a  and  a7529a );
 a7541a <=( A236  and  A234 );
 a7542a <=( (not A233)  and  a7541a );
 a7545a <=( (not A299)  and  A298 );
 a7548a <=( A301  and  A300 );
 a7549a <=( a7548a  and  a7545a );
 a7550a <=( a7549a  and  a7542a );
 a7554a <=( A167  and  A168 );
 a7555a <=( (not A170)  and  a7554a );
 a7558a <=( (not A201)  and  (not A166) );
 a7561a <=( A232  and  A202 );
 a7562a <=( a7561a  and  a7558a );
 a7563a <=( a7562a  and  a7555a );
 a7567a <=( A236  and  A234 );
 a7568a <=( (not A233)  and  a7567a );
 a7571a <=( (not A299)  and  A298 );
 a7574a <=( A302  and  A300 );
 a7575a <=( a7574a  and  a7571a );
 a7576a <=( a7575a  and  a7568a );
 a7580a <=( A167  and  A168 );
 a7581a <=( (not A170)  and  a7580a );
 a7584a <=( (not A201)  and  (not A166) );
 a7587a <=( A232  and  A202 );
 a7588a <=( a7587a  and  a7584a );
 a7589a <=( a7588a  and  a7581a );
 a7593a <=( A236  and  A234 );
 a7594a <=( (not A233)  and  a7593a );
 a7597a <=( A299  and  (not A298) );
 a7600a <=( A301  and  A300 );
 a7601a <=( a7600a  and  a7597a );
 a7602a <=( a7601a  and  a7594a );
 a7606a <=( A167  and  A168 );
 a7607a <=( (not A170)  and  a7606a );
 a7610a <=( (not A201)  and  (not A166) );
 a7613a <=( A232  and  A202 );
 a7614a <=( a7613a  and  a7610a );
 a7615a <=( a7614a  and  a7607a );
 a7619a <=( A236  and  A234 );
 a7620a <=( (not A233)  and  a7619a );
 a7623a <=( A299  and  (not A298) );
 a7626a <=( A302  and  A300 );
 a7627a <=( a7626a  and  a7623a );
 a7628a <=( a7627a  and  a7620a );
 a7632a <=( A167  and  A168 );
 a7633a <=( (not A170)  and  a7632a );
 a7636a <=( (not A201)  and  (not A166) );
 a7639a <=( A232  and  A202 );
 a7640a <=( a7639a  and  a7636a );
 a7641a <=( a7640a  and  a7633a );
 a7645a <=( A236  and  A234 );
 a7646a <=( (not A233)  and  a7645a );
 a7649a <=( A266  and  (not A265) );
 a7652a <=( A268  and  A267 );
 a7653a <=( a7652a  and  a7649a );
 a7654a <=( a7653a  and  a7646a );
 a7658a <=( A167  and  A168 );
 a7659a <=( (not A170)  and  a7658a );
 a7662a <=( (not A201)  and  (not A166) );
 a7665a <=( A232  and  A202 );
 a7666a <=( a7665a  and  a7662a );
 a7667a <=( a7666a  and  a7659a );
 a7671a <=( A236  and  A234 );
 a7672a <=( (not A233)  and  a7671a );
 a7675a <=( A266  and  (not A265) );
 a7678a <=( A269  and  A267 );
 a7679a <=( a7678a  and  a7675a );
 a7680a <=( a7679a  and  a7672a );
 a7684a <=( A167  and  A168 );
 a7685a <=( (not A170)  and  a7684a );
 a7688a <=( (not A201)  and  (not A166) );
 a7691a <=( A232  and  A202 );
 a7692a <=( a7691a  and  a7688a );
 a7693a <=( a7692a  and  a7685a );
 a7697a <=( A236  and  A234 );
 a7698a <=( (not A233)  and  a7697a );
 a7701a <=( (not A266)  and  A265 );
 a7704a <=( A268  and  A267 );
 a7705a <=( a7704a  and  a7701a );
 a7706a <=( a7705a  and  a7698a );
 a7710a <=( A167  and  A168 );
 a7711a <=( (not A170)  and  a7710a );
 a7714a <=( (not A201)  and  (not A166) );
 a7717a <=( A232  and  A202 );
 a7718a <=( a7717a  and  a7714a );
 a7719a <=( a7718a  and  a7711a );
 a7723a <=( A236  and  A234 );
 a7724a <=( (not A233)  and  a7723a );
 a7727a <=( (not A266)  and  A265 );
 a7730a <=( A269  and  A267 );
 a7731a <=( a7730a  and  a7727a );
 a7732a <=( a7731a  and  a7724a );
 a7736a <=( A167  and  A168 );
 a7737a <=( (not A170)  and  a7736a );
 a7740a <=( (not A201)  and  (not A166) );
 a7743a <=( (not A232)  and  A203 );
 a7744a <=( a7743a  and  a7740a );
 a7745a <=( a7744a  and  a7737a );
 a7749a <=( A235  and  A234 );
 a7750a <=( A233  and  a7749a );
 a7753a <=( (not A299)  and  A298 );
 a7756a <=( A301  and  A300 );
 a7757a <=( a7756a  and  a7753a );
 a7758a <=( a7757a  and  a7750a );
 a7762a <=( A167  and  A168 );
 a7763a <=( (not A170)  and  a7762a );
 a7766a <=( (not A201)  and  (not A166) );
 a7769a <=( (not A232)  and  A203 );
 a7770a <=( a7769a  and  a7766a );
 a7771a <=( a7770a  and  a7763a );
 a7775a <=( A235  and  A234 );
 a7776a <=( A233  and  a7775a );
 a7779a <=( (not A299)  and  A298 );
 a7782a <=( A302  and  A300 );
 a7783a <=( a7782a  and  a7779a );
 a7784a <=( a7783a  and  a7776a );
 a7788a <=( A167  and  A168 );
 a7789a <=( (not A170)  and  a7788a );
 a7792a <=( (not A201)  and  (not A166) );
 a7795a <=( (not A232)  and  A203 );
 a7796a <=( a7795a  and  a7792a );
 a7797a <=( a7796a  and  a7789a );
 a7801a <=( A235  and  A234 );
 a7802a <=( A233  and  a7801a );
 a7805a <=( A299  and  (not A298) );
 a7808a <=( A301  and  A300 );
 a7809a <=( a7808a  and  a7805a );
 a7810a <=( a7809a  and  a7802a );
 a7814a <=( A167  and  A168 );
 a7815a <=( (not A170)  and  a7814a );
 a7818a <=( (not A201)  and  (not A166) );
 a7821a <=( (not A232)  and  A203 );
 a7822a <=( a7821a  and  a7818a );
 a7823a <=( a7822a  and  a7815a );
 a7827a <=( A235  and  A234 );
 a7828a <=( A233  and  a7827a );
 a7831a <=( A299  and  (not A298) );
 a7834a <=( A302  and  A300 );
 a7835a <=( a7834a  and  a7831a );
 a7836a <=( a7835a  and  a7828a );
 a7840a <=( A167  and  A168 );
 a7841a <=( (not A170)  and  a7840a );
 a7844a <=( (not A201)  and  (not A166) );
 a7847a <=( (not A232)  and  A203 );
 a7848a <=( a7847a  and  a7844a );
 a7849a <=( a7848a  and  a7841a );
 a7853a <=( A235  and  A234 );
 a7854a <=( A233  and  a7853a );
 a7857a <=( A266  and  (not A265) );
 a7860a <=( A268  and  A267 );
 a7861a <=( a7860a  and  a7857a );
 a7862a <=( a7861a  and  a7854a );
 a7866a <=( A167  and  A168 );
 a7867a <=( (not A170)  and  a7866a );
 a7870a <=( (not A201)  and  (not A166) );
 a7873a <=( (not A232)  and  A203 );
 a7874a <=( a7873a  and  a7870a );
 a7875a <=( a7874a  and  a7867a );
 a7879a <=( A235  and  A234 );
 a7880a <=( A233  and  a7879a );
 a7883a <=( A266  and  (not A265) );
 a7886a <=( A269  and  A267 );
 a7887a <=( a7886a  and  a7883a );
 a7888a <=( a7887a  and  a7880a );
 a7892a <=( A167  and  A168 );
 a7893a <=( (not A170)  and  a7892a );
 a7896a <=( (not A201)  and  (not A166) );
 a7899a <=( (not A232)  and  A203 );
 a7900a <=( a7899a  and  a7896a );
 a7901a <=( a7900a  and  a7893a );
 a7905a <=( A235  and  A234 );
 a7906a <=( A233  and  a7905a );
 a7909a <=( (not A266)  and  A265 );
 a7912a <=( A268  and  A267 );
 a7913a <=( a7912a  and  a7909a );
 a7914a <=( a7913a  and  a7906a );
 a7918a <=( A167  and  A168 );
 a7919a <=( (not A170)  and  a7918a );
 a7922a <=( (not A201)  and  (not A166) );
 a7925a <=( (not A232)  and  A203 );
 a7926a <=( a7925a  and  a7922a );
 a7927a <=( a7926a  and  a7919a );
 a7931a <=( A235  and  A234 );
 a7932a <=( A233  and  a7931a );
 a7935a <=( (not A266)  and  A265 );
 a7938a <=( A269  and  A267 );
 a7939a <=( a7938a  and  a7935a );
 a7940a <=( a7939a  and  a7932a );
 a7944a <=( A167  and  A168 );
 a7945a <=( (not A170)  and  a7944a );
 a7948a <=( (not A201)  and  (not A166) );
 a7951a <=( (not A232)  and  A203 );
 a7952a <=( a7951a  and  a7948a );
 a7953a <=( a7952a  and  a7945a );
 a7957a <=( A236  and  A234 );
 a7958a <=( A233  and  a7957a );
 a7961a <=( (not A299)  and  A298 );
 a7964a <=( A301  and  A300 );
 a7965a <=( a7964a  and  a7961a );
 a7966a <=( a7965a  and  a7958a );
 a7970a <=( A167  and  A168 );
 a7971a <=( (not A170)  and  a7970a );
 a7974a <=( (not A201)  and  (not A166) );
 a7977a <=( (not A232)  and  A203 );
 a7978a <=( a7977a  and  a7974a );
 a7979a <=( a7978a  and  a7971a );
 a7983a <=( A236  and  A234 );
 a7984a <=( A233  and  a7983a );
 a7987a <=( (not A299)  and  A298 );
 a7990a <=( A302  and  A300 );
 a7991a <=( a7990a  and  a7987a );
 a7992a <=( a7991a  and  a7984a );
 a7996a <=( A167  and  A168 );
 a7997a <=( (not A170)  and  a7996a );
 a8000a <=( (not A201)  and  (not A166) );
 a8003a <=( (not A232)  and  A203 );
 a8004a <=( a8003a  and  a8000a );
 a8005a <=( a8004a  and  a7997a );
 a8009a <=( A236  and  A234 );
 a8010a <=( A233  and  a8009a );
 a8013a <=( A299  and  (not A298) );
 a8016a <=( A301  and  A300 );
 a8017a <=( a8016a  and  a8013a );
 a8018a <=( a8017a  and  a8010a );
 a8022a <=( A167  and  A168 );
 a8023a <=( (not A170)  and  a8022a );
 a8026a <=( (not A201)  and  (not A166) );
 a8029a <=( (not A232)  and  A203 );
 a8030a <=( a8029a  and  a8026a );
 a8031a <=( a8030a  and  a8023a );
 a8035a <=( A236  and  A234 );
 a8036a <=( A233  and  a8035a );
 a8039a <=( A299  and  (not A298) );
 a8042a <=( A302  and  A300 );
 a8043a <=( a8042a  and  a8039a );
 a8044a <=( a8043a  and  a8036a );
 a8048a <=( A167  and  A168 );
 a8049a <=( (not A170)  and  a8048a );
 a8052a <=( (not A201)  and  (not A166) );
 a8055a <=( (not A232)  and  A203 );
 a8056a <=( a8055a  and  a8052a );
 a8057a <=( a8056a  and  a8049a );
 a8061a <=( A236  and  A234 );
 a8062a <=( A233  and  a8061a );
 a8065a <=( A266  and  (not A265) );
 a8068a <=( A268  and  A267 );
 a8069a <=( a8068a  and  a8065a );
 a8070a <=( a8069a  and  a8062a );
 a8074a <=( A167  and  A168 );
 a8075a <=( (not A170)  and  a8074a );
 a8078a <=( (not A201)  and  (not A166) );
 a8081a <=( (not A232)  and  A203 );
 a8082a <=( a8081a  and  a8078a );
 a8083a <=( a8082a  and  a8075a );
 a8087a <=( A236  and  A234 );
 a8088a <=( A233  and  a8087a );
 a8091a <=( A266  and  (not A265) );
 a8094a <=( A269  and  A267 );
 a8095a <=( a8094a  and  a8091a );
 a8096a <=( a8095a  and  a8088a );
 a8100a <=( A167  and  A168 );
 a8101a <=( (not A170)  and  a8100a );
 a8104a <=( (not A201)  and  (not A166) );
 a8107a <=( (not A232)  and  A203 );
 a8108a <=( a8107a  and  a8104a );
 a8109a <=( a8108a  and  a8101a );
 a8113a <=( A236  and  A234 );
 a8114a <=( A233  and  a8113a );
 a8117a <=( (not A266)  and  A265 );
 a8120a <=( A268  and  A267 );
 a8121a <=( a8120a  and  a8117a );
 a8122a <=( a8121a  and  a8114a );
 a8126a <=( A167  and  A168 );
 a8127a <=( (not A170)  and  a8126a );
 a8130a <=( (not A201)  and  (not A166) );
 a8133a <=( (not A232)  and  A203 );
 a8134a <=( a8133a  and  a8130a );
 a8135a <=( a8134a  and  a8127a );
 a8139a <=( A236  and  A234 );
 a8140a <=( A233  and  a8139a );
 a8143a <=( (not A266)  and  A265 );
 a8146a <=( A269  and  A267 );
 a8147a <=( a8146a  and  a8143a );
 a8148a <=( a8147a  and  a8140a );
 a8152a <=( A167  and  A168 );
 a8153a <=( (not A170)  and  a8152a );
 a8156a <=( (not A201)  and  (not A166) );
 a8159a <=( A232  and  A203 );
 a8160a <=( a8159a  and  a8156a );
 a8161a <=( a8160a  and  a8153a );
 a8165a <=( A235  and  A234 );
 a8166a <=( (not A233)  and  a8165a );
 a8169a <=( (not A299)  and  A298 );
 a8172a <=( A301  and  A300 );
 a8173a <=( a8172a  and  a8169a );
 a8174a <=( a8173a  and  a8166a );
 a8178a <=( A167  and  A168 );
 a8179a <=( (not A170)  and  a8178a );
 a8182a <=( (not A201)  and  (not A166) );
 a8185a <=( A232  and  A203 );
 a8186a <=( a8185a  and  a8182a );
 a8187a <=( a8186a  and  a8179a );
 a8191a <=( A235  and  A234 );
 a8192a <=( (not A233)  and  a8191a );
 a8195a <=( (not A299)  and  A298 );
 a8198a <=( A302  and  A300 );
 a8199a <=( a8198a  and  a8195a );
 a8200a <=( a8199a  and  a8192a );
 a8204a <=( A167  and  A168 );
 a8205a <=( (not A170)  and  a8204a );
 a8208a <=( (not A201)  and  (not A166) );
 a8211a <=( A232  and  A203 );
 a8212a <=( a8211a  and  a8208a );
 a8213a <=( a8212a  and  a8205a );
 a8217a <=( A235  and  A234 );
 a8218a <=( (not A233)  and  a8217a );
 a8221a <=( A299  and  (not A298) );
 a8224a <=( A301  and  A300 );
 a8225a <=( a8224a  and  a8221a );
 a8226a <=( a8225a  and  a8218a );
 a8230a <=( A167  and  A168 );
 a8231a <=( (not A170)  and  a8230a );
 a8234a <=( (not A201)  and  (not A166) );
 a8237a <=( A232  and  A203 );
 a8238a <=( a8237a  and  a8234a );
 a8239a <=( a8238a  and  a8231a );
 a8243a <=( A235  and  A234 );
 a8244a <=( (not A233)  and  a8243a );
 a8247a <=( A299  and  (not A298) );
 a8250a <=( A302  and  A300 );
 a8251a <=( a8250a  and  a8247a );
 a8252a <=( a8251a  and  a8244a );
 a8256a <=( A167  and  A168 );
 a8257a <=( (not A170)  and  a8256a );
 a8260a <=( (not A201)  and  (not A166) );
 a8263a <=( A232  and  A203 );
 a8264a <=( a8263a  and  a8260a );
 a8265a <=( a8264a  and  a8257a );
 a8269a <=( A235  and  A234 );
 a8270a <=( (not A233)  and  a8269a );
 a8273a <=( A266  and  (not A265) );
 a8276a <=( A268  and  A267 );
 a8277a <=( a8276a  and  a8273a );
 a8278a <=( a8277a  and  a8270a );
 a8282a <=( A167  and  A168 );
 a8283a <=( (not A170)  and  a8282a );
 a8286a <=( (not A201)  and  (not A166) );
 a8289a <=( A232  and  A203 );
 a8290a <=( a8289a  and  a8286a );
 a8291a <=( a8290a  and  a8283a );
 a8295a <=( A235  and  A234 );
 a8296a <=( (not A233)  and  a8295a );
 a8299a <=( A266  and  (not A265) );
 a8302a <=( A269  and  A267 );
 a8303a <=( a8302a  and  a8299a );
 a8304a <=( a8303a  and  a8296a );
 a8308a <=( A167  and  A168 );
 a8309a <=( (not A170)  and  a8308a );
 a8312a <=( (not A201)  and  (not A166) );
 a8315a <=( A232  and  A203 );
 a8316a <=( a8315a  and  a8312a );
 a8317a <=( a8316a  and  a8309a );
 a8321a <=( A235  and  A234 );
 a8322a <=( (not A233)  and  a8321a );
 a8325a <=( (not A266)  and  A265 );
 a8328a <=( A268  and  A267 );
 a8329a <=( a8328a  and  a8325a );
 a8330a <=( a8329a  and  a8322a );
 a8334a <=( A167  and  A168 );
 a8335a <=( (not A170)  and  a8334a );
 a8338a <=( (not A201)  and  (not A166) );
 a8341a <=( A232  and  A203 );
 a8342a <=( a8341a  and  a8338a );
 a8343a <=( a8342a  and  a8335a );
 a8347a <=( A235  and  A234 );
 a8348a <=( (not A233)  and  a8347a );
 a8351a <=( (not A266)  and  A265 );
 a8354a <=( A269  and  A267 );
 a8355a <=( a8354a  and  a8351a );
 a8356a <=( a8355a  and  a8348a );
 a8360a <=( A167  and  A168 );
 a8361a <=( (not A170)  and  a8360a );
 a8364a <=( (not A201)  and  (not A166) );
 a8367a <=( A232  and  A203 );
 a8368a <=( a8367a  and  a8364a );
 a8369a <=( a8368a  and  a8361a );
 a8373a <=( A236  and  A234 );
 a8374a <=( (not A233)  and  a8373a );
 a8377a <=( (not A299)  and  A298 );
 a8380a <=( A301  and  A300 );
 a8381a <=( a8380a  and  a8377a );
 a8382a <=( a8381a  and  a8374a );
 a8386a <=( A167  and  A168 );
 a8387a <=( (not A170)  and  a8386a );
 a8390a <=( (not A201)  and  (not A166) );
 a8393a <=( A232  and  A203 );
 a8394a <=( a8393a  and  a8390a );
 a8395a <=( a8394a  and  a8387a );
 a8399a <=( A236  and  A234 );
 a8400a <=( (not A233)  and  a8399a );
 a8403a <=( (not A299)  and  A298 );
 a8406a <=( A302  and  A300 );
 a8407a <=( a8406a  and  a8403a );
 a8408a <=( a8407a  and  a8400a );
 a8412a <=( A167  and  A168 );
 a8413a <=( (not A170)  and  a8412a );
 a8416a <=( (not A201)  and  (not A166) );
 a8419a <=( A232  and  A203 );
 a8420a <=( a8419a  and  a8416a );
 a8421a <=( a8420a  and  a8413a );
 a8425a <=( A236  and  A234 );
 a8426a <=( (not A233)  and  a8425a );
 a8429a <=( A299  and  (not A298) );
 a8432a <=( A301  and  A300 );
 a8433a <=( a8432a  and  a8429a );
 a8434a <=( a8433a  and  a8426a );
 a8438a <=( A167  and  A168 );
 a8439a <=( (not A170)  and  a8438a );
 a8442a <=( (not A201)  and  (not A166) );
 a8445a <=( A232  and  A203 );
 a8446a <=( a8445a  and  a8442a );
 a8447a <=( a8446a  and  a8439a );
 a8451a <=( A236  and  A234 );
 a8452a <=( (not A233)  and  a8451a );
 a8455a <=( A299  and  (not A298) );
 a8458a <=( A302  and  A300 );
 a8459a <=( a8458a  and  a8455a );
 a8460a <=( a8459a  and  a8452a );
 a8464a <=( A167  and  A168 );
 a8465a <=( (not A170)  and  a8464a );
 a8468a <=( (not A201)  and  (not A166) );
 a8471a <=( A232  and  A203 );
 a8472a <=( a8471a  and  a8468a );
 a8473a <=( a8472a  and  a8465a );
 a8477a <=( A236  and  A234 );
 a8478a <=( (not A233)  and  a8477a );
 a8481a <=( A266  and  (not A265) );
 a8484a <=( A268  and  A267 );
 a8485a <=( a8484a  and  a8481a );
 a8486a <=( a8485a  and  a8478a );
 a8490a <=( A167  and  A168 );
 a8491a <=( (not A170)  and  a8490a );
 a8494a <=( (not A201)  and  (not A166) );
 a8497a <=( A232  and  A203 );
 a8498a <=( a8497a  and  a8494a );
 a8499a <=( a8498a  and  a8491a );
 a8503a <=( A236  and  A234 );
 a8504a <=( (not A233)  and  a8503a );
 a8507a <=( A266  and  (not A265) );
 a8510a <=( A269  and  A267 );
 a8511a <=( a8510a  and  a8507a );
 a8512a <=( a8511a  and  a8504a );
 a8516a <=( A167  and  A168 );
 a8517a <=( (not A170)  and  a8516a );
 a8520a <=( (not A201)  and  (not A166) );
 a8523a <=( A232  and  A203 );
 a8524a <=( a8523a  and  a8520a );
 a8525a <=( a8524a  and  a8517a );
 a8529a <=( A236  and  A234 );
 a8530a <=( (not A233)  and  a8529a );
 a8533a <=( (not A266)  and  A265 );
 a8536a <=( A268  and  A267 );
 a8537a <=( a8536a  and  a8533a );
 a8538a <=( a8537a  and  a8530a );
 a8542a <=( A167  and  A168 );
 a8543a <=( (not A170)  and  a8542a );
 a8546a <=( (not A201)  and  (not A166) );
 a8549a <=( A232  and  A203 );
 a8550a <=( a8549a  and  a8546a );
 a8551a <=( a8550a  and  a8543a );
 a8555a <=( A236  and  A234 );
 a8556a <=( (not A233)  and  a8555a );
 a8559a <=( (not A266)  and  A265 );
 a8562a <=( A269  and  A267 );
 a8563a <=( a8562a  and  a8559a );
 a8564a <=( a8563a  and  a8556a );
 a8568a <=( A167  and  A168 );
 a8569a <=( (not A170)  and  a8568a );
 a8572a <=( A199  and  (not A166) );
 a8575a <=( (not A232)  and  A200 );
 a8576a <=( a8575a  and  a8572a );
 a8577a <=( a8576a  and  a8569a );
 a8581a <=( A235  and  A234 );
 a8582a <=( A233  and  a8581a );
 a8585a <=( (not A299)  and  A298 );
 a8588a <=( A301  and  A300 );
 a8589a <=( a8588a  and  a8585a );
 a8590a <=( a8589a  and  a8582a );
 a8594a <=( A167  and  A168 );
 a8595a <=( (not A170)  and  a8594a );
 a8598a <=( A199  and  (not A166) );
 a8601a <=( (not A232)  and  A200 );
 a8602a <=( a8601a  and  a8598a );
 a8603a <=( a8602a  and  a8595a );
 a8607a <=( A235  and  A234 );
 a8608a <=( A233  and  a8607a );
 a8611a <=( (not A299)  and  A298 );
 a8614a <=( A302  and  A300 );
 a8615a <=( a8614a  and  a8611a );
 a8616a <=( a8615a  and  a8608a );
 a8620a <=( A167  and  A168 );
 a8621a <=( (not A170)  and  a8620a );
 a8624a <=( A199  and  (not A166) );
 a8627a <=( (not A232)  and  A200 );
 a8628a <=( a8627a  and  a8624a );
 a8629a <=( a8628a  and  a8621a );
 a8633a <=( A235  and  A234 );
 a8634a <=( A233  and  a8633a );
 a8637a <=( A299  and  (not A298) );
 a8640a <=( A301  and  A300 );
 a8641a <=( a8640a  and  a8637a );
 a8642a <=( a8641a  and  a8634a );
 a8646a <=( A167  and  A168 );
 a8647a <=( (not A170)  and  a8646a );
 a8650a <=( A199  and  (not A166) );
 a8653a <=( (not A232)  and  A200 );
 a8654a <=( a8653a  and  a8650a );
 a8655a <=( a8654a  and  a8647a );
 a8659a <=( A235  and  A234 );
 a8660a <=( A233  and  a8659a );
 a8663a <=( A299  and  (not A298) );
 a8666a <=( A302  and  A300 );
 a8667a <=( a8666a  and  a8663a );
 a8668a <=( a8667a  and  a8660a );
 a8672a <=( A167  and  A168 );
 a8673a <=( (not A170)  and  a8672a );
 a8676a <=( A199  and  (not A166) );
 a8679a <=( (not A232)  and  A200 );
 a8680a <=( a8679a  and  a8676a );
 a8681a <=( a8680a  and  a8673a );
 a8685a <=( A235  and  A234 );
 a8686a <=( A233  and  a8685a );
 a8689a <=( A266  and  (not A265) );
 a8692a <=( A268  and  A267 );
 a8693a <=( a8692a  and  a8689a );
 a8694a <=( a8693a  and  a8686a );
 a8698a <=( A167  and  A168 );
 a8699a <=( (not A170)  and  a8698a );
 a8702a <=( A199  and  (not A166) );
 a8705a <=( (not A232)  and  A200 );
 a8706a <=( a8705a  and  a8702a );
 a8707a <=( a8706a  and  a8699a );
 a8711a <=( A235  and  A234 );
 a8712a <=( A233  and  a8711a );
 a8715a <=( A266  and  (not A265) );
 a8718a <=( A269  and  A267 );
 a8719a <=( a8718a  and  a8715a );
 a8720a <=( a8719a  and  a8712a );
 a8724a <=( A167  and  A168 );
 a8725a <=( (not A170)  and  a8724a );
 a8728a <=( A199  and  (not A166) );
 a8731a <=( (not A232)  and  A200 );
 a8732a <=( a8731a  and  a8728a );
 a8733a <=( a8732a  and  a8725a );
 a8737a <=( A235  and  A234 );
 a8738a <=( A233  and  a8737a );
 a8741a <=( (not A266)  and  A265 );
 a8744a <=( A268  and  A267 );
 a8745a <=( a8744a  and  a8741a );
 a8746a <=( a8745a  and  a8738a );
 a8750a <=( A167  and  A168 );
 a8751a <=( (not A170)  and  a8750a );
 a8754a <=( A199  and  (not A166) );
 a8757a <=( (not A232)  and  A200 );
 a8758a <=( a8757a  and  a8754a );
 a8759a <=( a8758a  and  a8751a );
 a8763a <=( A235  and  A234 );
 a8764a <=( A233  and  a8763a );
 a8767a <=( (not A266)  and  A265 );
 a8770a <=( A269  and  A267 );
 a8771a <=( a8770a  and  a8767a );
 a8772a <=( a8771a  and  a8764a );
 a8776a <=( A167  and  A168 );
 a8777a <=( (not A170)  and  a8776a );
 a8780a <=( A199  and  (not A166) );
 a8783a <=( (not A232)  and  A200 );
 a8784a <=( a8783a  and  a8780a );
 a8785a <=( a8784a  and  a8777a );
 a8789a <=( A236  and  A234 );
 a8790a <=( A233  and  a8789a );
 a8793a <=( (not A299)  and  A298 );
 a8796a <=( A301  and  A300 );
 a8797a <=( a8796a  and  a8793a );
 a8798a <=( a8797a  and  a8790a );
 a8802a <=( A167  and  A168 );
 a8803a <=( (not A170)  and  a8802a );
 a8806a <=( A199  and  (not A166) );
 a8809a <=( (not A232)  and  A200 );
 a8810a <=( a8809a  and  a8806a );
 a8811a <=( a8810a  and  a8803a );
 a8815a <=( A236  and  A234 );
 a8816a <=( A233  and  a8815a );
 a8819a <=( (not A299)  and  A298 );
 a8822a <=( A302  and  A300 );
 a8823a <=( a8822a  and  a8819a );
 a8824a <=( a8823a  and  a8816a );
 a8828a <=( A167  and  A168 );
 a8829a <=( (not A170)  and  a8828a );
 a8832a <=( A199  and  (not A166) );
 a8835a <=( (not A232)  and  A200 );
 a8836a <=( a8835a  and  a8832a );
 a8837a <=( a8836a  and  a8829a );
 a8841a <=( A236  and  A234 );
 a8842a <=( A233  and  a8841a );
 a8845a <=( A299  and  (not A298) );
 a8848a <=( A301  and  A300 );
 a8849a <=( a8848a  and  a8845a );
 a8850a <=( a8849a  and  a8842a );
 a8854a <=( A167  and  A168 );
 a8855a <=( (not A170)  and  a8854a );
 a8858a <=( A199  and  (not A166) );
 a8861a <=( (not A232)  and  A200 );
 a8862a <=( a8861a  and  a8858a );
 a8863a <=( a8862a  and  a8855a );
 a8867a <=( A236  and  A234 );
 a8868a <=( A233  and  a8867a );
 a8871a <=( A299  and  (not A298) );
 a8874a <=( A302  and  A300 );
 a8875a <=( a8874a  and  a8871a );
 a8876a <=( a8875a  and  a8868a );
 a8880a <=( A167  and  A168 );
 a8881a <=( (not A170)  and  a8880a );
 a8884a <=( A199  and  (not A166) );
 a8887a <=( (not A232)  and  A200 );
 a8888a <=( a8887a  and  a8884a );
 a8889a <=( a8888a  and  a8881a );
 a8893a <=( A236  and  A234 );
 a8894a <=( A233  and  a8893a );
 a8897a <=( A266  and  (not A265) );
 a8900a <=( A268  and  A267 );
 a8901a <=( a8900a  and  a8897a );
 a8902a <=( a8901a  and  a8894a );
 a8906a <=( A167  and  A168 );
 a8907a <=( (not A170)  and  a8906a );
 a8910a <=( A199  and  (not A166) );
 a8913a <=( (not A232)  and  A200 );
 a8914a <=( a8913a  and  a8910a );
 a8915a <=( a8914a  and  a8907a );
 a8919a <=( A236  and  A234 );
 a8920a <=( A233  and  a8919a );
 a8923a <=( A266  and  (not A265) );
 a8926a <=( A269  and  A267 );
 a8927a <=( a8926a  and  a8923a );
 a8928a <=( a8927a  and  a8920a );
 a8932a <=( A167  and  A168 );
 a8933a <=( (not A170)  and  a8932a );
 a8936a <=( A199  and  (not A166) );
 a8939a <=( (not A232)  and  A200 );
 a8940a <=( a8939a  and  a8936a );
 a8941a <=( a8940a  and  a8933a );
 a8945a <=( A236  and  A234 );
 a8946a <=( A233  and  a8945a );
 a8949a <=( (not A266)  and  A265 );
 a8952a <=( A268  and  A267 );
 a8953a <=( a8952a  and  a8949a );
 a8954a <=( a8953a  and  a8946a );
 a8958a <=( A167  and  A168 );
 a8959a <=( (not A170)  and  a8958a );
 a8962a <=( A199  and  (not A166) );
 a8965a <=( (not A232)  and  A200 );
 a8966a <=( a8965a  and  a8962a );
 a8967a <=( a8966a  and  a8959a );
 a8971a <=( A236  and  A234 );
 a8972a <=( A233  and  a8971a );
 a8975a <=( (not A266)  and  A265 );
 a8978a <=( A269  and  A267 );
 a8979a <=( a8978a  and  a8975a );
 a8980a <=( a8979a  and  a8972a );
 a8984a <=( A167  and  A168 );
 a8985a <=( (not A170)  and  a8984a );
 a8988a <=( A199  and  (not A166) );
 a8991a <=( A232  and  A200 );
 a8992a <=( a8991a  and  a8988a );
 a8993a <=( a8992a  and  a8985a );
 a8997a <=( A235  and  A234 );
 a8998a <=( (not A233)  and  a8997a );
 a9001a <=( (not A299)  and  A298 );
 a9004a <=( A301  and  A300 );
 a9005a <=( a9004a  and  a9001a );
 a9006a <=( a9005a  and  a8998a );
 a9010a <=( A167  and  A168 );
 a9011a <=( (not A170)  and  a9010a );
 a9014a <=( A199  and  (not A166) );
 a9017a <=( A232  and  A200 );
 a9018a <=( a9017a  and  a9014a );
 a9019a <=( a9018a  and  a9011a );
 a9023a <=( A235  and  A234 );
 a9024a <=( (not A233)  and  a9023a );
 a9027a <=( (not A299)  and  A298 );
 a9030a <=( A302  and  A300 );
 a9031a <=( a9030a  and  a9027a );
 a9032a <=( a9031a  and  a9024a );
 a9036a <=( A167  and  A168 );
 a9037a <=( (not A170)  and  a9036a );
 a9040a <=( A199  and  (not A166) );
 a9043a <=( A232  and  A200 );
 a9044a <=( a9043a  and  a9040a );
 a9045a <=( a9044a  and  a9037a );
 a9049a <=( A235  and  A234 );
 a9050a <=( (not A233)  and  a9049a );
 a9053a <=( A299  and  (not A298) );
 a9056a <=( A301  and  A300 );
 a9057a <=( a9056a  and  a9053a );
 a9058a <=( a9057a  and  a9050a );
 a9062a <=( A167  and  A168 );
 a9063a <=( (not A170)  and  a9062a );
 a9066a <=( A199  and  (not A166) );
 a9069a <=( A232  and  A200 );
 a9070a <=( a9069a  and  a9066a );
 a9071a <=( a9070a  and  a9063a );
 a9075a <=( A235  and  A234 );
 a9076a <=( (not A233)  and  a9075a );
 a9079a <=( A299  and  (not A298) );
 a9082a <=( A302  and  A300 );
 a9083a <=( a9082a  and  a9079a );
 a9084a <=( a9083a  and  a9076a );
 a9088a <=( A167  and  A168 );
 a9089a <=( (not A170)  and  a9088a );
 a9092a <=( A199  and  (not A166) );
 a9095a <=( A232  and  A200 );
 a9096a <=( a9095a  and  a9092a );
 a9097a <=( a9096a  and  a9089a );
 a9101a <=( A235  and  A234 );
 a9102a <=( (not A233)  and  a9101a );
 a9105a <=( A266  and  (not A265) );
 a9108a <=( A268  and  A267 );
 a9109a <=( a9108a  and  a9105a );
 a9110a <=( a9109a  and  a9102a );
 a9114a <=( A167  and  A168 );
 a9115a <=( (not A170)  and  a9114a );
 a9118a <=( A199  and  (not A166) );
 a9121a <=( A232  and  A200 );
 a9122a <=( a9121a  and  a9118a );
 a9123a <=( a9122a  and  a9115a );
 a9127a <=( A235  and  A234 );
 a9128a <=( (not A233)  and  a9127a );
 a9131a <=( A266  and  (not A265) );
 a9134a <=( A269  and  A267 );
 a9135a <=( a9134a  and  a9131a );
 a9136a <=( a9135a  and  a9128a );
 a9140a <=( A167  and  A168 );
 a9141a <=( (not A170)  and  a9140a );
 a9144a <=( A199  and  (not A166) );
 a9147a <=( A232  and  A200 );
 a9148a <=( a9147a  and  a9144a );
 a9149a <=( a9148a  and  a9141a );
 a9153a <=( A235  and  A234 );
 a9154a <=( (not A233)  and  a9153a );
 a9157a <=( (not A266)  and  A265 );
 a9160a <=( A268  and  A267 );
 a9161a <=( a9160a  and  a9157a );
 a9162a <=( a9161a  and  a9154a );
 a9166a <=( A167  and  A168 );
 a9167a <=( (not A170)  and  a9166a );
 a9170a <=( A199  and  (not A166) );
 a9173a <=( A232  and  A200 );
 a9174a <=( a9173a  and  a9170a );
 a9175a <=( a9174a  and  a9167a );
 a9179a <=( A235  and  A234 );
 a9180a <=( (not A233)  and  a9179a );
 a9183a <=( (not A266)  and  A265 );
 a9186a <=( A269  and  A267 );
 a9187a <=( a9186a  and  a9183a );
 a9188a <=( a9187a  and  a9180a );
 a9192a <=( A167  and  A168 );
 a9193a <=( (not A170)  and  a9192a );
 a9196a <=( A199  and  (not A166) );
 a9199a <=( A232  and  A200 );
 a9200a <=( a9199a  and  a9196a );
 a9201a <=( a9200a  and  a9193a );
 a9205a <=( A236  and  A234 );
 a9206a <=( (not A233)  and  a9205a );
 a9209a <=( (not A299)  and  A298 );
 a9212a <=( A301  and  A300 );
 a9213a <=( a9212a  and  a9209a );
 a9214a <=( a9213a  and  a9206a );
 a9218a <=( A167  and  A168 );
 a9219a <=( (not A170)  and  a9218a );
 a9222a <=( A199  and  (not A166) );
 a9225a <=( A232  and  A200 );
 a9226a <=( a9225a  and  a9222a );
 a9227a <=( a9226a  and  a9219a );
 a9231a <=( A236  and  A234 );
 a9232a <=( (not A233)  and  a9231a );
 a9235a <=( (not A299)  and  A298 );
 a9238a <=( A302  and  A300 );
 a9239a <=( a9238a  and  a9235a );
 a9240a <=( a9239a  and  a9232a );
 a9244a <=( A167  and  A168 );
 a9245a <=( (not A170)  and  a9244a );
 a9248a <=( A199  and  (not A166) );
 a9251a <=( A232  and  A200 );
 a9252a <=( a9251a  and  a9248a );
 a9253a <=( a9252a  and  a9245a );
 a9257a <=( A236  and  A234 );
 a9258a <=( (not A233)  and  a9257a );
 a9261a <=( A299  and  (not A298) );
 a9264a <=( A301  and  A300 );
 a9265a <=( a9264a  and  a9261a );
 a9266a <=( a9265a  and  a9258a );
 a9270a <=( A167  and  A168 );
 a9271a <=( (not A170)  and  a9270a );
 a9274a <=( A199  and  (not A166) );
 a9277a <=( A232  and  A200 );
 a9278a <=( a9277a  and  a9274a );
 a9279a <=( a9278a  and  a9271a );
 a9283a <=( A236  and  A234 );
 a9284a <=( (not A233)  and  a9283a );
 a9287a <=( A299  and  (not A298) );
 a9290a <=( A302  and  A300 );
 a9291a <=( a9290a  and  a9287a );
 a9292a <=( a9291a  and  a9284a );
 a9296a <=( A167  and  A168 );
 a9297a <=( (not A170)  and  a9296a );
 a9300a <=( A199  and  (not A166) );
 a9303a <=( A232  and  A200 );
 a9304a <=( a9303a  and  a9300a );
 a9305a <=( a9304a  and  a9297a );
 a9309a <=( A236  and  A234 );
 a9310a <=( (not A233)  and  a9309a );
 a9313a <=( A266  and  (not A265) );
 a9316a <=( A268  and  A267 );
 a9317a <=( a9316a  and  a9313a );
 a9318a <=( a9317a  and  a9310a );
 a9322a <=( A167  and  A168 );
 a9323a <=( (not A170)  and  a9322a );
 a9326a <=( A199  and  (not A166) );
 a9329a <=( A232  and  A200 );
 a9330a <=( a9329a  and  a9326a );
 a9331a <=( a9330a  and  a9323a );
 a9335a <=( A236  and  A234 );
 a9336a <=( (not A233)  and  a9335a );
 a9339a <=( A266  and  (not A265) );
 a9342a <=( A269  and  A267 );
 a9343a <=( a9342a  and  a9339a );
 a9344a <=( a9343a  and  a9336a );
 a9348a <=( A167  and  A168 );
 a9349a <=( (not A170)  and  a9348a );
 a9352a <=( A199  and  (not A166) );
 a9355a <=( A232  and  A200 );
 a9356a <=( a9355a  and  a9352a );
 a9357a <=( a9356a  and  a9349a );
 a9361a <=( A236  and  A234 );
 a9362a <=( (not A233)  and  a9361a );
 a9365a <=( (not A266)  and  A265 );
 a9368a <=( A268  and  A267 );
 a9369a <=( a9368a  and  a9365a );
 a9370a <=( a9369a  and  a9362a );
 a9374a <=( A167  and  A168 );
 a9375a <=( (not A170)  and  a9374a );
 a9378a <=( A199  and  (not A166) );
 a9381a <=( A232  and  A200 );
 a9382a <=( a9381a  and  a9378a );
 a9383a <=( a9382a  and  a9375a );
 a9387a <=( A236  and  A234 );
 a9388a <=( (not A233)  and  a9387a );
 a9391a <=( (not A266)  and  A265 );
 a9394a <=( A269  and  A267 );
 a9395a <=( a9394a  and  a9391a );
 a9396a <=( a9395a  and  a9388a );
 a9400a <=( A167  and  A168 );
 a9401a <=( (not A170)  and  a9400a );
 a9404a <=( (not A199)  and  (not A166) );
 a9407a <=( (not A232)  and  (not A200) );
 a9408a <=( a9407a  and  a9404a );
 a9409a <=( a9408a  and  a9401a );
 a9413a <=( A235  and  A234 );
 a9414a <=( A233  and  a9413a );
 a9417a <=( (not A299)  and  A298 );
 a9420a <=( A301  and  A300 );
 a9421a <=( a9420a  and  a9417a );
 a9422a <=( a9421a  and  a9414a );
 a9426a <=( A167  and  A168 );
 a9427a <=( (not A170)  and  a9426a );
 a9430a <=( (not A199)  and  (not A166) );
 a9433a <=( (not A232)  and  (not A200) );
 a9434a <=( a9433a  and  a9430a );
 a9435a <=( a9434a  and  a9427a );
 a9439a <=( A235  and  A234 );
 a9440a <=( A233  and  a9439a );
 a9443a <=( (not A299)  and  A298 );
 a9446a <=( A302  and  A300 );
 a9447a <=( a9446a  and  a9443a );
 a9448a <=( a9447a  and  a9440a );
 a9452a <=( A167  and  A168 );
 a9453a <=( (not A170)  and  a9452a );
 a9456a <=( (not A199)  and  (not A166) );
 a9459a <=( (not A232)  and  (not A200) );
 a9460a <=( a9459a  and  a9456a );
 a9461a <=( a9460a  and  a9453a );
 a9465a <=( A235  and  A234 );
 a9466a <=( A233  and  a9465a );
 a9469a <=( A299  and  (not A298) );
 a9472a <=( A301  and  A300 );
 a9473a <=( a9472a  and  a9469a );
 a9474a <=( a9473a  and  a9466a );
 a9478a <=( A167  and  A168 );
 a9479a <=( (not A170)  and  a9478a );
 a9482a <=( (not A199)  and  (not A166) );
 a9485a <=( (not A232)  and  (not A200) );
 a9486a <=( a9485a  and  a9482a );
 a9487a <=( a9486a  and  a9479a );
 a9491a <=( A235  and  A234 );
 a9492a <=( A233  and  a9491a );
 a9495a <=( A299  and  (not A298) );
 a9498a <=( A302  and  A300 );
 a9499a <=( a9498a  and  a9495a );
 a9500a <=( a9499a  and  a9492a );
 a9504a <=( A167  and  A168 );
 a9505a <=( (not A170)  and  a9504a );
 a9508a <=( (not A199)  and  (not A166) );
 a9511a <=( (not A232)  and  (not A200) );
 a9512a <=( a9511a  and  a9508a );
 a9513a <=( a9512a  and  a9505a );
 a9517a <=( A235  and  A234 );
 a9518a <=( A233  and  a9517a );
 a9521a <=( A266  and  (not A265) );
 a9524a <=( A268  and  A267 );
 a9525a <=( a9524a  and  a9521a );
 a9526a <=( a9525a  and  a9518a );
 a9530a <=( A167  and  A168 );
 a9531a <=( (not A170)  and  a9530a );
 a9534a <=( (not A199)  and  (not A166) );
 a9537a <=( (not A232)  and  (not A200) );
 a9538a <=( a9537a  and  a9534a );
 a9539a <=( a9538a  and  a9531a );
 a9543a <=( A235  and  A234 );
 a9544a <=( A233  and  a9543a );
 a9547a <=( A266  and  (not A265) );
 a9550a <=( A269  and  A267 );
 a9551a <=( a9550a  and  a9547a );
 a9552a <=( a9551a  and  a9544a );
 a9556a <=( A167  and  A168 );
 a9557a <=( (not A170)  and  a9556a );
 a9560a <=( (not A199)  and  (not A166) );
 a9563a <=( (not A232)  and  (not A200) );
 a9564a <=( a9563a  and  a9560a );
 a9565a <=( a9564a  and  a9557a );
 a9569a <=( A235  and  A234 );
 a9570a <=( A233  and  a9569a );
 a9573a <=( (not A266)  and  A265 );
 a9576a <=( A268  and  A267 );
 a9577a <=( a9576a  and  a9573a );
 a9578a <=( a9577a  and  a9570a );
 a9582a <=( A167  and  A168 );
 a9583a <=( (not A170)  and  a9582a );
 a9586a <=( (not A199)  and  (not A166) );
 a9589a <=( (not A232)  and  (not A200) );
 a9590a <=( a9589a  and  a9586a );
 a9591a <=( a9590a  and  a9583a );
 a9595a <=( A235  and  A234 );
 a9596a <=( A233  and  a9595a );
 a9599a <=( (not A266)  and  A265 );
 a9602a <=( A269  and  A267 );
 a9603a <=( a9602a  and  a9599a );
 a9604a <=( a9603a  and  a9596a );
 a9608a <=( A167  and  A168 );
 a9609a <=( (not A170)  and  a9608a );
 a9612a <=( (not A199)  and  (not A166) );
 a9615a <=( (not A232)  and  (not A200) );
 a9616a <=( a9615a  and  a9612a );
 a9617a <=( a9616a  and  a9609a );
 a9621a <=( A236  and  A234 );
 a9622a <=( A233  and  a9621a );
 a9625a <=( (not A299)  and  A298 );
 a9628a <=( A301  and  A300 );
 a9629a <=( a9628a  and  a9625a );
 a9630a <=( a9629a  and  a9622a );
 a9634a <=( A167  and  A168 );
 a9635a <=( (not A170)  and  a9634a );
 a9638a <=( (not A199)  and  (not A166) );
 a9641a <=( (not A232)  and  (not A200) );
 a9642a <=( a9641a  and  a9638a );
 a9643a <=( a9642a  and  a9635a );
 a9647a <=( A236  and  A234 );
 a9648a <=( A233  and  a9647a );
 a9651a <=( (not A299)  and  A298 );
 a9654a <=( A302  and  A300 );
 a9655a <=( a9654a  and  a9651a );
 a9656a <=( a9655a  and  a9648a );
 a9660a <=( A167  and  A168 );
 a9661a <=( (not A170)  and  a9660a );
 a9664a <=( (not A199)  and  (not A166) );
 a9667a <=( (not A232)  and  (not A200) );
 a9668a <=( a9667a  and  a9664a );
 a9669a <=( a9668a  and  a9661a );
 a9673a <=( A236  and  A234 );
 a9674a <=( A233  and  a9673a );
 a9677a <=( A299  and  (not A298) );
 a9680a <=( A301  and  A300 );
 a9681a <=( a9680a  and  a9677a );
 a9682a <=( a9681a  and  a9674a );
 a9686a <=( A167  and  A168 );
 a9687a <=( (not A170)  and  a9686a );
 a9690a <=( (not A199)  and  (not A166) );
 a9693a <=( (not A232)  and  (not A200) );
 a9694a <=( a9693a  and  a9690a );
 a9695a <=( a9694a  and  a9687a );
 a9699a <=( A236  and  A234 );
 a9700a <=( A233  and  a9699a );
 a9703a <=( A299  and  (not A298) );
 a9706a <=( A302  and  A300 );
 a9707a <=( a9706a  and  a9703a );
 a9708a <=( a9707a  and  a9700a );
 a9712a <=( A167  and  A168 );
 a9713a <=( (not A170)  and  a9712a );
 a9716a <=( (not A199)  and  (not A166) );
 a9719a <=( (not A232)  and  (not A200) );
 a9720a <=( a9719a  and  a9716a );
 a9721a <=( a9720a  and  a9713a );
 a9725a <=( A236  and  A234 );
 a9726a <=( A233  and  a9725a );
 a9729a <=( A266  and  (not A265) );
 a9732a <=( A268  and  A267 );
 a9733a <=( a9732a  and  a9729a );
 a9734a <=( a9733a  and  a9726a );
 a9738a <=( A167  and  A168 );
 a9739a <=( (not A170)  and  a9738a );
 a9742a <=( (not A199)  and  (not A166) );
 a9745a <=( (not A232)  and  (not A200) );
 a9746a <=( a9745a  and  a9742a );
 a9747a <=( a9746a  and  a9739a );
 a9751a <=( A236  and  A234 );
 a9752a <=( A233  and  a9751a );
 a9755a <=( A266  and  (not A265) );
 a9758a <=( A269  and  A267 );
 a9759a <=( a9758a  and  a9755a );
 a9760a <=( a9759a  and  a9752a );
 a9764a <=( A167  and  A168 );
 a9765a <=( (not A170)  and  a9764a );
 a9768a <=( (not A199)  and  (not A166) );
 a9771a <=( (not A232)  and  (not A200) );
 a9772a <=( a9771a  and  a9768a );
 a9773a <=( a9772a  and  a9765a );
 a9777a <=( A236  and  A234 );
 a9778a <=( A233  and  a9777a );
 a9781a <=( (not A266)  and  A265 );
 a9784a <=( A268  and  A267 );
 a9785a <=( a9784a  and  a9781a );
 a9786a <=( a9785a  and  a9778a );
 a9790a <=( A167  and  A168 );
 a9791a <=( (not A170)  and  a9790a );
 a9794a <=( (not A199)  and  (not A166) );
 a9797a <=( (not A232)  and  (not A200) );
 a9798a <=( a9797a  and  a9794a );
 a9799a <=( a9798a  and  a9791a );
 a9803a <=( A236  and  A234 );
 a9804a <=( A233  and  a9803a );
 a9807a <=( (not A266)  and  A265 );
 a9810a <=( A269  and  A267 );
 a9811a <=( a9810a  and  a9807a );
 a9812a <=( a9811a  and  a9804a );
 a9816a <=( A167  and  A168 );
 a9817a <=( (not A170)  and  a9816a );
 a9820a <=( (not A199)  and  (not A166) );
 a9823a <=( A232  and  (not A200) );
 a9824a <=( a9823a  and  a9820a );
 a9825a <=( a9824a  and  a9817a );
 a9829a <=( A235  and  A234 );
 a9830a <=( (not A233)  and  a9829a );
 a9833a <=( (not A299)  and  A298 );
 a9836a <=( A301  and  A300 );
 a9837a <=( a9836a  and  a9833a );
 a9838a <=( a9837a  and  a9830a );
 a9842a <=( A167  and  A168 );
 a9843a <=( (not A170)  and  a9842a );
 a9846a <=( (not A199)  and  (not A166) );
 a9849a <=( A232  and  (not A200) );
 a9850a <=( a9849a  and  a9846a );
 a9851a <=( a9850a  and  a9843a );
 a9855a <=( A235  and  A234 );
 a9856a <=( (not A233)  and  a9855a );
 a9859a <=( (not A299)  and  A298 );
 a9862a <=( A302  and  A300 );
 a9863a <=( a9862a  and  a9859a );
 a9864a <=( a9863a  and  a9856a );
 a9868a <=( A167  and  A168 );
 a9869a <=( (not A170)  and  a9868a );
 a9872a <=( (not A199)  and  (not A166) );
 a9875a <=( A232  and  (not A200) );
 a9876a <=( a9875a  and  a9872a );
 a9877a <=( a9876a  and  a9869a );
 a9881a <=( A235  and  A234 );
 a9882a <=( (not A233)  and  a9881a );
 a9885a <=( A299  and  (not A298) );
 a9888a <=( A301  and  A300 );
 a9889a <=( a9888a  and  a9885a );
 a9890a <=( a9889a  and  a9882a );
 a9894a <=( A167  and  A168 );
 a9895a <=( (not A170)  and  a9894a );
 a9898a <=( (not A199)  and  (not A166) );
 a9901a <=( A232  and  (not A200) );
 a9902a <=( a9901a  and  a9898a );
 a9903a <=( a9902a  and  a9895a );
 a9907a <=( A235  and  A234 );
 a9908a <=( (not A233)  and  a9907a );
 a9911a <=( A299  and  (not A298) );
 a9914a <=( A302  and  A300 );
 a9915a <=( a9914a  and  a9911a );
 a9916a <=( a9915a  and  a9908a );
 a9920a <=( A167  and  A168 );
 a9921a <=( (not A170)  and  a9920a );
 a9924a <=( (not A199)  and  (not A166) );
 a9927a <=( A232  and  (not A200) );
 a9928a <=( a9927a  and  a9924a );
 a9929a <=( a9928a  and  a9921a );
 a9933a <=( A235  and  A234 );
 a9934a <=( (not A233)  and  a9933a );
 a9937a <=( A266  and  (not A265) );
 a9940a <=( A268  and  A267 );
 a9941a <=( a9940a  and  a9937a );
 a9942a <=( a9941a  and  a9934a );
 a9946a <=( A167  and  A168 );
 a9947a <=( (not A170)  and  a9946a );
 a9950a <=( (not A199)  and  (not A166) );
 a9953a <=( A232  and  (not A200) );
 a9954a <=( a9953a  and  a9950a );
 a9955a <=( a9954a  and  a9947a );
 a9959a <=( A235  and  A234 );
 a9960a <=( (not A233)  and  a9959a );
 a9963a <=( A266  and  (not A265) );
 a9966a <=( A269  and  A267 );
 a9967a <=( a9966a  and  a9963a );
 a9968a <=( a9967a  and  a9960a );
 a9972a <=( A167  and  A168 );
 a9973a <=( (not A170)  and  a9972a );
 a9976a <=( (not A199)  and  (not A166) );
 a9979a <=( A232  and  (not A200) );
 a9980a <=( a9979a  and  a9976a );
 a9981a <=( a9980a  and  a9973a );
 a9985a <=( A235  and  A234 );
 a9986a <=( (not A233)  and  a9985a );
 a9989a <=( (not A266)  and  A265 );
 a9992a <=( A268  and  A267 );
 a9993a <=( a9992a  and  a9989a );
 a9994a <=( a9993a  and  a9986a );
 a9998a <=( A167  and  A168 );
 a9999a <=( (not A170)  and  a9998a );
 a10002a <=( (not A199)  and  (not A166) );
 a10005a <=( A232  and  (not A200) );
 a10006a <=( a10005a  and  a10002a );
 a10007a <=( a10006a  and  a9999a );
 a10011a <=( A235  and  A234 );
 a10012a <=( (not A233)  and  a10011a );
 a10015a <=( (not A266)  and  A265 );
 a10018a <=( A269  and  A267 );
 a10019a <=( a10018a  and  a10015a );
 a10020a <=( a10019a  and  a10012a );
 a10024a <=( A167  and  A168 );
 a10025a <=( (not A170)  and  a10024a );
 a10028a <=( (not A199)  and  (not A166) );
 a10031a <=( A232  and  (not A200) );
 a10032a <=( a10031a  and  a10028a );
 a10033a <=( a10032a  and  a10025a );
 a10037a <=( A236  and  A234 );
 a10038a <=( (not A233)  and  a10037a );
 a10041a <=( (not A299)  and  A298 );
 a10044a <=( A301  and  A300 );
 a10045a <=( a10044a  and  a10041a );
 a10046a <=( a10045a  and  a10038a );
 a10050a <=( A167  and  A168 );
 a10051a <=( (not A170)  and  a10050a );
 a10054a <=( (not A199)  and  (not A166) );
 a10057a <=( A232  and  (not A200) );
 a10058a <=( a10057a  and  a10054a );
 a10059a <=( a10058a  and  a10051a );
 a10063a <=( A236  and  A234 );
 a10064a <=( (not A233)  and  a10063a );
 a10067a <=( (not A299)  and  A298 );
 a10070a <=( A302  and  A300 );
 a10071a <=( a10070a  and  a10067a );
 a10072a <=( a10071a  and  a10064a );
 a10076a <=( A167  and  A168 );
 a10077a <=( (not A170)  and  a10076a );
 a10080a <=( (not A199)  and  (not A166) );
 a10083a <=( A232  and  (not A200) );
 a10084a <=( a10083a  and  a10080a );
 a10085a <=( a10084a  and  a10077a );
 a10089a <=( A236  and  A234 );
 a10090a <=( (not A233)  and  a10089a );
 a10093a <=( A299  and  (not A298) );
 a10096a <=( A301  and  A300 );
 a10097a <=( a10096a  and  a10093a );
 a10098a <=( a10097a  and  a10090a );
 a10102a <=( A167  and  A168 );
 a10103a <=( (not A170)  and  a10102a );
 a10106a <=( (not A199)  and  (not A166) );
 a10109a <=( A232  and  (not A200) );
 a10110a <=( a10109a  and  a10106a );
 a10111a <=( a10110a  and  a10103a );
 a10115a <=( A236  and  A234 );
 a10116a <=( (not A233)  and  a10115a );
 a10119a <=( A299  and  (not A298) );
 a10122a <=( A302  and  A300 );
 a10123a <=( a10122a  and  a10119a );
 a10124a <=( a10123a  and  a10116a );
 a10128a <=( A167  and  A168 );
 a10129a <=( (not A170)  and  a10128a );
 a10132a <=( (not A199)  and  (not A166) );
 a10135a <=( A232  and  (not A200) );
 a10136a <=( a10135a  and  a10132a );
 a10137a <=( a10136a  and  a10129a );
 a10141a <=( A236  and  A234 );
 a10142a <=( (not A233)  and  a10141a );
 a10145a <=( A266  and  (not A265) );
 a10148a <=( A268  and  A267 );
 a10149a <=( a10148a  and  a10145a );
 a10150a <=( a10149a  and  a10142a );
 a10154a <=( A167  and  A168 );
 a10155a <=( (not A170)  and  a10154a );
 a10158a <=( (not A199)  and  (not A166) );
 a10161a <=( A232  and  (not A200) );
 a10162a <=( a10161a  and  a10158a );
 a10163a <=( a10162a  and  a10155a );
 a10167a <=( A236  and  A234 );
 a10168a <=( (not A233)  and  a10167a );
 a10171a <=( A266  and  (not A265) );
 a10174a <=( A269  and  A267 );
 a10175a <=( a10174a  and  a10171a );
 a10176a <=( a10175a  and  a10168a );
 a10180a <=( A167  and  A168 );
 a10181a <=( (not A170)  and  a10180a );
 a10184a <=( (not A199)  and  (not A166) );
 a10187a <=( A232  and  (not A200) );
 a10188a <=( a10187a  and  a10184a );
 a10189a <=( a10188a  and  a10181a );
 a10193a <=( A236  and  A234 );
 a10194a <=( (not A233)  and  a10193a );
 a10197a <=( (not A266)  and  A265 );
 a10200a <=( A268  and  A267 );
 a10201a <=( a10200a  and  a10197a );
 a10202a <=( a10201a  and  a10194a );
 a10206a <=( A167  and  A168 );
 a10207a <=( (not A170)  and  a10206a );
 a10210a <=( (not A199)  and  (not A166) );
 a10213a <=( A232  and  (not A200) );
 a10214a <=( a10213a  and  a10210a );
 a10215a <=( a10214a  and  a10207a );
 a10219a <=( A236  and  A234 );
 a10220a <=( (not A233)  and  a10219a );
 a10223a <=( (not A266)  and  A265 );
 a10226a <=( A269  and  A267 );
 a10227a <=( a10226a  and  a10223a );
 a10228a <=( a10227a  and  a10220a );
 a10232a <=( (not A167)  and  A168 );
 a10233a <=( (not A170)  and  a10232a );
 a10236a <=( (not A201)  and  A166 );
 a10239a <=( (not A232)  and  A202 );
 a10240a <=( a10239a  and  a10236a );
 a10241a <=( a10240a  and  a10233a );
 a10245a <=( A235  and  A234 );
 a10246a <=( A233  and  a10245a );
 a10249a <=( (not A299)  and  A298 );
 a10252a <=( A301  and  A300 );
 a10253a <=( a10252a  and  a10249a );
 a10254a <=( a10253a  and  a10246a );
 a10258a <=( (not A167)  and  A168 );
 a10259a <=( (not A170)  and  a10258a );
 a10262a <=( (not A201)  and  A166 );
 a10265a <=( (not A232)  and  A202 );
 a10266a <=( a10265a  and  a10262a );
 a10267a <=( a10266a  and  a10259a );
 a10271a <=( A235  and  A234 );
 a10272a <=( A233  and  a10271a );
 a10275a <=( (not A299)  and  A298 );
 a10278a <=( A302  and  A300 );
 a10279a <=( a10278a  and  a10275a );
 a10280a <=( a10279a  and  a10272a );
 a10284a <=( (not A167)  and  A168 );
 a10285a <=( (not A170)  and  a10284a );
 a10288a <=( (not A201)  and  A166 );
 a10291a <=( (not A232)  and  A202 );
 a10292a <=( a10291a  and  a10288a );
 a10293a <=( a10292a  and  a10285a );
 a10297a <=( A235  and  A234 );
 a10298a <=( A233  and  a10297a );
 a10301a <=( A299  and  (not A298) );
 a10304a <=( A301  and  A300 );
 a10305a <=( a10304a  and  a10301a );
 a10306a <=( a10305a  and  a10298a );
 a10310a <=( (not A167)  and  A168 );
 a10311a <=( (not A170)  and  a10310a );
 a10314a <=( (not A201)  and  A166 );
 a10317a <=( (not A232)  and  A202 );
 a10318a <=( a10317a  and  a10314a );
 a10319a <=( a10318a  and  a10311a );
 a10323a <=( A235  and  A234 );
 a10324a <=( A233  and  a10323a );
 a10327a <=( A299  and  (not A298) );
 a10330a <=( A302  and  A300 );
 a10331a <=( a10330a  and  a10327a );
 a10332a <=( a10331a  and  a10324a );
 a10336a <=( (not A167)  and  A168 );
 a10337a <=( (not A170)  and  a10336a );
 a10340a <=( (not A201)  and  A166 );
 a10343a <=( (not A232)  and  A202 );
 a10344a <=( a10343a  and  a10340a );
 a10345a <=( a10344a  and  a10337a );
 a10349a <=( A235  and  A234 );
 a10350a <=( A233  and  a10349a );
 a10353a <=( A266  and  (not A265) );
 a10356a <=( A268  and  A267 );
 a10357a <=( a10356a  and  a10353a );
 a10358a <=( a10357a  and  a10350a );
 a10362a <=( (not A167)  and  A168 );
 a10363a <=( (not A170)  and  a10362a );
 a10366a <=( (not A201)  and  A166 );
 a10369a <=( (not A232)  and  A202 );
 a10370a <=( a10369a  and  a10366a );
 a10371a <=( a10370a  and  a10363a );
 a10375a <=( A235  and  A234 );
 a10376a <=( A233  and  a10375a );
 a10379a <=( A266  and  (not A265) );
 a10382a <=( A269  and  A267 );
 a10383a <=( a10382a  and  a10379a );
 a10384a <=( a10383a  and  a10376a );
 a10388a <=( (not A167)  and  A168 );
 a10389a <=( (not A170)  and  a10388a );
 a10392a <=( (not A201)  and  A166 );
 a10395a <=( (not A232)  and  A202 );
 a10396a <=( a10395a  and  a10392a );
 a10397a <=( a10396a  and  a10389a );
 a10401a <=( A235  and  A234 );
 a10402a <=( A233  and  a10401a );
 a10405a <=( (not A266)  and  A265 );
 a10408a <=( A268  and  A267 );
 a10409a <=( a10408a  and  a10405a );
 a10410a <=( a10409a  and  a10402a );
 a10414a <=( (not A167)  and  A168 );
 a10415a <=( (not A170)  and  a10414a );
 a10418a <=( (not A201)  and  A166 );
 a10421a <=( (not A232)  and  A202 );
 a10422a <=( a10421a  and  a10418a );
 a10423a <=( a10422a  and  a10415a );
 a10427a <=( A235  and  A234 );
 a10428a <=( A233  and  a10427a );
 a10431a <=( (not A266)  and  A265 );
 a10434a <=( A269  and  A267 );
 a10435a <=( a10434a  and  a10431a );
 a10436a <=( a10435a  and  a10428a );
 a10440a <=( (not A167)  and  A168 );
 a10441a <=( (not A170)  and  a10440a );
 a10444a <=( (not A201)  and  A166 );
 a10447a <=( (not A232)  and  A202 );
 a10448a <=( a10447a  and  a10444a );
 a10449a <=( a10448a  and  a10441a );
 a10453a <=( A236  and  A234 );
 a10454a <=( A233  and  a10453a );
 a10457a <=( (not A299)  and  A298 );
 a10460a <=( A301  and  A300 );
 a10461a <=( a10460a  and  a10457a );
 a10462a <=( a10461a  and  a10454a );
 a10466a <=( (not A167)  and  A168 );
 a10467a <=( (not A170)  and  a10466a );
 a10470a <=( (not A201)  and  A166 );
 a10473a <=( (not A232)  and  A202 );
 a10474a <=( a10473a  and  a10470a );
 a10475a <=( a10474a  and  a10467a );
 a10479a <=( A236  and  A234 );
 a10480a <=( A233  and  a10479a );
 a10483a <=( (not A299)  and  A298 );
 a10486a <=( A302  and  A300 );
 a10487a <=( a10486a  and  a10483a );
 a10488a <=( a10487a  and  a10480a );
 a10492a <=( (not A167)  and  A168 );
 a10493a <=( (not A170)  and  a10492a );
 a10496a <=( (not A201)  and  A166 );
 a10499a <=( (not A232)  and  A202 );
 a10500a <=( a10499a  and  a10496a );
 a10501a <=( a10500a  and  a10493a );
 a10505a <=( A236  and  A234 );
 a10506a <=( A233  and  a10505a );
 a10509a <=( A299  and  (not A298) );
 a10512a <=( A301  and  A300 );
 a10513a <=( a10512a  and  a10509a );
 a10514a <=( a10513a  and  a10506a );
 a10518a <=( (not A167)  and  A168 );
 a10519a <=( (not A170)  and  a10518a );
 a10522a <=( (not A201)  and  A166 );
 a10525a <=( (not A232)  and  A202 );
 a10526a <=( a10525a  and  a10522a );
 a10527a <=( a10526a  and  a10519a );
 a10531a <=( A236  and  A234 );
 a10532a <=( A233  and  a10531a );
 a10535a <=( A299  and  (not A298) );
 a10538a <=( A302  and  A300 );
 a10539a <=( a10538a  and  a10535a );
 a10540a <=( a10539a  and  a10532a );
 a10544a <=( (not A167)  and  A168 );
 a10545a <=( (not A170)  and  a10544a );
 a10548a <=( (not A201)  and  A166 );
 a10551a <=( (not A232)  and  A202 );
 a10552a <=( a10551a  and  a10548a );
 a10553a <=( a10552a  and  a10545a );
 a10557a <=( A236  and  A234 );
 a10558a <=( A233  and  a10557a );
 a10561a <=( A266  and  (not A265) );
 a10564a <=( A268  and  A267 );
 a10565a <=( a10564a  and  a10561a );
 a10566a <=( a10565a  and  a10558a );
 a10570a <=( (not A167)  and  A168 );
 a10571a <=( (not A170)  and  a10570a );
 a10574a <=( (not A201)  and  A166 );
 a10577a <=( (not A232)  and  A202 );
 a10578a <=( a10577a  and  a10574a );
 a10579a <=( a10578a  and  a10571a );
 a10583a <=( A236  and  A234 );
 a10584a <=( A233  and  a10583a );
 a10587a <=( A266  and  (not A265) );
 a10590a <=( A269  and  A267 );
 a10591a <=( a10590a  and  a10587a );
 a10592a <=( a10591a  and  a10584a );
 a10596a <=( (not A167)  and  A168 );
 a10597a <=( (not A170)  and  a10596a );
 a10600a <=( (not A201)  and  A166 );
 a10603a <=( (not A232)  and  A202 );
 a10604a <=( a10603a  and  a10600a );
 a10605a <=( a10604a  and  a10597a );
 a10609a <=( A236  and  A234 );
 a10610a <=( A233  and  a10609a );
 a10613a <=( (not A266)  and  A265 );
 a10616a <=( A268  and  A267 );
 a10617a <=( a10616a  and  a10613a );
 a10618a <=( a10617a  and  a10610a );
 a10622a <=( (not A167)  and  A168 );
 a10623a <=( (not A170)  and  a10622a );
 a10626a <=( (not A201)  and  A166 );
 a10629a <=( (not A232)  and  A202 );
 a10630a <=( a10629a  and  a10626a );
 a10631a <=( a10630a  and  a10623a );
 a10635a <=( A236  and  A234 );
 a10636a <=( A233  and  a10635a );
 a10639a <=( (not A266)  and  A265 );
 a10642a <=( A269  and  A267 );
 a10643a <=( a10642a  and  a10639a );
 a10644a <=( a10643a  and  a10636a );
 a10648a <=( (not A167)  and  A168 );
 a10649a <=( (not A170)  and  a10648a );
 a10652a <=( (not A201)  and  A166 );
 a10655a <=( A232  and  A202 );
 a10656a <=( a10655a  and  a10652a );
 a10657a <=( a10656a  and  a10649a );
 a10661a <=( A235  and  A234 );
 a10662a <=( (not A233)  and  a10661a );
 a10665a <=( (not A299)  and  A298 );
 a10668a <=( A301  and  A300 );
 a10669a <=( a10668a  and  a10665a );
 a10670a <=( a10669a  and  a10662a );
 a10674a <=( (not A167)  and  A168 );
 a10675a <=( (not A170)  and  a10674a );
 a10678a <=( (not A201)  and  A166 );
 a10681a <=( A232  and  A202 );
 a10682a <=( a10681a  and  a10678a );
 a10683a <=( a10682a  and  a10675a );
 a10687a <=( A235  and  A234 );
 a10688a <=( (not A233)  and  a10687a );
 a10691a <=( (not A299)  and  A298 );
 a10694a <=( A302  and  A300 );
 a10695a <=( a10694a  and  a10691a );
 a10696a <=( a10695a  and  a10688a );
 a10700a <=( (not A167)  and  A168 );
 a10701a <=( (not A170)  and  a10700a );
 a10704a <=( (not A201)  and  A166 );
 a10707a <=( A232  and  A202 );
 a10708a <=( a10707a  and  a10704a );
 a10709a <=( a10708a  and  a10701a );
 a10713a <=( A235  and  A234 );
 a10714a <=( (not A233)  and  a10713a );
 a10717a <=( A299  and  (not A298) );
 a10720a <=( A301  and  A300 );
 a10721a <=( a10720a  and  a10717a );
 a10722a <=( a10721a  and  a10714a );
 a10726a <=( (not A167)  and  A168 );
 a10727a <=( (not A170)  and  a10726a );
 a10730a <=( (not A201)  and  A166 );
 a10733a <=( A232  and  A202 );
 a10734a <=( a10733a  and  a10730a );
 a10735a <=( a10734a  and  a10727a );
 a10739a <=( A235  and  A234 );
 a10740a <=( (not A233)  and  a10739a );
 a10743a <=( A299  and  (not A298) );
 a10746a <=( A302  and  A300 );
 a10747a <=( a10746a  and  a10743a );
 a10748a <=( a10747a  and  a10740a );
 a10752a <=( (not A167)  and  A168 );
 a10753a <=( (not A170)  and  a10752a );
 a10756a <=( (not A201)  and  A166 );
 a10759a <=( A232  and  A202 );
 a10760a <=( a10759a  and  a10756a );
 a10761a <=( a10760a  and  a10753a );
 a10765a <=( A235  and  A234 );
 a10766a <=( (not A233)  and  a10765a );
 a10769a <=( A266  and  (not A265) );
 a10772a <=( A268  and  A267 );
 a10773a <=( a10772a  and  a10769a );
 a10774a <=( a10773a  and  a10766a );
 a10778a <=( (not A167)  and  A168 );
 a10779a <=( (not A170)  and  a10778a );
 a10782a <=( (not A201)  and  A166 );
 a10785a <=( A232  and  A202 );
 a10786a <=( a10785a  and  a10782a );
 a10787a <=( a10786a  and  a10779a );
 a10791a <=( A235  and  A234 );
 a10792a <=( (not A233)  and  a10791a );
 a10795a <=( A266  and  (not A265) );
 a10798a <=( A269  and  A267 );
 a10799a <=( a10798a  and  a10795a );
 a10800a <=( a10799a  and  a10792a );
 a10804a <=( (not A167)  and  A168 );
 a10805a <=( (not A170)  and  a10804a );
 a10808a <=( (not A201)  and  A166 );
 a10811a <=( A232  and  A202 );
 a10812a <=( a10811a  and  a10808a );
 a10813a <=( a10812a  and  a10805a );
 a10817a <=( A235  and  A234 );
 a10818a <=( (not A233)  and  a10817a );
 a10821a <=( (not A266)  and  A265 );
 a10824a <=( A268  and  A267 );
 a10825a <=( a10824a  and  a10821a );
 a10826a <=( a10825a  and  a10818a );
 a10830a <=( (not A167)  and  A168 );
 a10831a <=( (not A170)  and  a10830a );
 a10834a <=( (not A201)  and  A166 );
 a10837a <=( A232  and  A202 );
 a10838a <=( a10837a  and  a10834a );
 a10839a <=( a10838a  and  a10831a );
 a10843a <=( A235  and  A234 );
 a10844a <=( (not A233)  and  a10843a );
 a10847a <=( (not A266)  and  A265 );
 a10850a <=( A269  and  A267 );
 a10851a <=( a10850a  and  a10847a );
 a10852a <=( a10851a  and  a10844a );
 a10856a <=( (not A167)  and  A168 );
 a10857a <=( (not A170)  and  a10856a );
 a10860a <=( (not A201)  and  A166 );
 a10863a <=( A232  and  A202 );
 a10864a <=( a10863a  and  a10860a );
 a10865a <=( a10864a  and  a10857a );
 a10869a <=( A236  and  A234 );
 a10870a <=( (not A233)  and  a10869a );
 a10873a <=( (not A299)  and  A298 );
 a10876a <=( A301  and  A300 );
 a10877a <=( a10876a  and  a10873a );
 a10878a <=( a10877a  and  a10870a );
 a10882a <=( (not A167)  and  A168 );
 a10883a <=( (not A170)  and  a10882a );
 a10886a <=( (not A201)  and  A166 );
 a10889a <=( A232  and  A202 );
 a10890a <=( a10889a  and  a10886a );
 a10891a <=( a10890a  and  a10883a );
 a10895a <=( A236  and  A234 );
 a10896a <=( (not A233)  and  a10895a );
 a10899a <=( (not A299)  and  A298 );
 a10902a <=( A302  and  A300 );
 a10903a <=( a10902a  and  a10899a );
 a10904a <=( a10903a  and  a10896a );
 a10908a <=( (not A167)  and  A168 );
 a10909a <=( (not A170)  and  a10908a );
 a10912a <=( (not A201)  and  A166 );
 a10915a <=( A232  and  A202 );
 a10916a <=( a10915a  and  a10912a );
 a10917a <=( a10916a  and  a10909a );
 a10921a <=( A236  and  A234 );
 a10922a <=( (not A233)  and  a10921a );
 a10925a <=( A299  and  (not A298) );
 a10928a <=( A301  and  A300 );
 a10929a <=( a10928a  and  a10925a );
 a10930a <=( a10929a  and  a10922a );
 a10934a <=( (not A167)  and  A168 );
 a10935a <=( (not A170)  and  a10934a );
 a10938a <=( (not A201)  and  A166 );
 a10941a <=( A232  and  A202 );
 a10942a <=( a10941a  and  a10938a );
 a10943a <=( a10942a  and  a10935a );
 a10947a <=( A236  and  A234 );
 a10948a <=( (not A233)  and  a10947a );
 a10951a <=( A299  and  (not A298) );
 a10954a <=( A302  and  A300 );
 a10955a <=( a10954a  and  a10951a );
 a10956a <=( a10955a  and  a10948a );
 a10960a <=( (not A167)  and  A168 );
 a10961a <=( (not A170)  and  a10960a );
 a10964a <=( (not A201)  and  A166 );
 a10967a <=( A232  and  A202 );
 a10968a <=( a10967a  and  a10964a );
 a10969a <=( a10968a  and  a10961a );
 a10973a <=( A236  and  A234 );
 a10974a <=( (not A233)  and  a10973a );
 a10977a <=( A266  and  (not A265) );
 a10980a <=( A268  and  A267 );
 a10981a <=( a10980a  and  a10977a );
 a10982a <=( a10981a  and  a10974a );
 a10986a <=( (not A167)  and  A168 );
 a10987a <=( (not A170)  and  a10986a );
 a10990a <=( (not A201)  and  A166 );
 a10993a <=( A232  and  A202 );
 a10994a <=( a10993a  and  a10990a );
 a10995a <=( a10994a  and  a10987a );
 a10999a <=( A236  and  A234 );
 a11000a <=( (not A233)  and  a10999a );
 a11003a <=( A266  and  (not A265) );
 a11006a <=( A269  and  A267 );
 a11007a <=( a11006a  and  a11003a );
 a11008a <=( a11007a  and  a11000a );
 a11012a <=( (not A167)  and  A168 );
 a11013a <=( (not A170)  and  a11012a );
 a11016a <=( (not A201)  and  A166 );
 a11019a <=( A232  and  A202 );
 a11020a <=( a11019a  and  a11016a );
 a11021a <=( a11020a  and  a11013a );
 a11025a <=( A236  and  A234 );
 a11026a <=( (not A233)  and  a11025a );
 a11029a <=( (not A266)  and  A265 );
 a11032a <=( A268  and  A267 );
 a11033a <=( a11032a  and  a11029a );
 a11034a <=( a11033a  and  a11026a );
 a11038a <=( (not A167)  and  A168 );
 a11039a <=( (not A170)  and  a11038a );
 a11042a <=( (not A201)  and  A166 );
 a11045a <=( A232  and  A202 );
 a11046a <=( a11045a  and  a11042a );
 a11047a <=( a11046a  and  a11039a );
 a11051a <=( A236  and  A234 );
 a11052a <=( (not A233)  and  a11051a );
 a11055a <=( (not A266)  and  A265 );
 a11058a <=( A269  and  A267 );
 a11059a <=( a11058a  and  a11055a );
 a11060a <=( a11059a  and  a11052a );
 a11064a <=( (not A167)  and  A168 );
 a11065a <=( (not A170)  and  a11064a );
 a11068a <=( (not A201)  and  A166 );
 a11071a <=( (not A232)  and  A203 );
 a11072a <=( a11071a  and  a11068a );
 a11073a <=( a11072a  and  a11065a );
 a11077a <=( A235  and  A234 );
 a11078a <=( A233  and  a11077a );
 a11081a <=( (not A299)  and  A298 );
 a11084a <=( A301  and  A300 );
 a11085a <=( a11084a  and  a11081a );
 a11086a <=( a11085a  and  a11078a );
 a11090a <=( (not A167)  and  A168 );
 a11091a <=( (not A170)  and  a11090a );
 a11094a <=( (not A201)  and  A166 );
 a11097a <=( (not A232)  and  A203 );
 a11098a <=( a11097a  and  a11094a );
 a11099a <=( a11098a  and  a11091a );
 a11103a <=( A235  and  A234 );
 a11104a <=( A233  and  a11103a );
 a11107a <=( (not A299)  and  A298 );
 a11110a <=( A302  and  A300 );
 a11111a <=( a11110a  and  a11107a );
 a11112a <=( a11111a  and  a11104a );
 a11116a <=( (not A167)  and  A168 );
 a11117a <=( (not A170)  and  a11116a );
 a11120a <=( (not A201)  and  A166 );
 a11123a <=( (not A232)  and  A203 );
 a11124a <=( a11123a  and  a11120a );
 a11125a <=( a11124a  and  a11117a );
 a11129a <=( A235  and  A234 );
 a11130a <=( A233  and  a11129a );
 a11133a <=( A299  and  (not A298) );
 a11136a <=( A301  and  A300 );
 a11137a <=( a11136a  and  a11133a );
 a11138a <=( a11137a  and  a11130a );
 a11142a <=( (not A167)  and  A168 );
 a11143a <=( (not A170)  and  a11142a );
 a11146a <=( (not A201)  and  A166 );
 a11149a <=( (not A232)  and  A203 );
 a11150a <=( a11149a  and  a11146a );
 a11151a <=( a11150a  and  a11143a );
 a11155a <=( A235  and  A234 );
 a11156a <=( A233  and  a11155a );
 a11159a <=( A299  and  (not A298) );
 a11162a <=( A302  and  A300 );
 a11163a <=( a11162a  and  a11159a );
 a11164a <=( a11163a  and  a11156a );
 a11168a <=( (not A167)  and  A168 );
 a11169a <=( (not A170)  and  a11168a );
 a11172a <=( (not A201)  and  A166 );
 a11175a <=( (not A232)  and  A203 );
 a11176a <=( a11175a  and  a11172a );
 a11177a <=( a11176a  and  a11169a );
 a11181a <=( A235  and  A234 );
 a11182a <=( A233  and  a11181a );
 a11185a <=( A266  and  (not A265) );
 a11188a <=( A268  and  A267 );
 a11189a <=( a11188a  and  a11185a );
 a11190a <=( a11189a  and  a11182a );
 a11194a <=( (not A167)  and  A168 );
 a11195a <=( (not A170)  and  a11194a );
 a11198a <=( (not A201)  and  A166 );
 a11201a <=( (not A232)  and  A203 );
 a11202a <=( a11201a  and  a11198a );
 a11203a <=( a11202a  and  a11195a );
 a11207a <=( A235  and  A234 );
 a11208a <=( A233  and  a11207a );
 a11211a <=( A266  and  (not A265) );
 a11214a <=( A269  and  A267 );
 a11215a <=( a11214a  and  a11211a );
 a11216a <=( a11215a  and  a11208a );
 a11220a <=( (not A167)  and  A168 );
 a11221a <=( (not A170)  and  a11220a );
 a11224a <=( (not A201)  and  A166 );
 a11227a <=( (not A232)  and  A203 );
 a11228a <=( a11227a  and  a11224a );
 a11229a <=( a11228a  and  a11221a );
 a11233a <=( A235  and  A234 );
 a11234a <=( A233  and  a11233a );
 a11237a <=( (not A266)  and  A265 );
 a11240a <=( A268  and  A267 );
 a11241a <=( a11240a  and  a11237a );
 a11242a <=( a11241a  and  a11234a );
 a11246a <=( (not A167)  and  A168 );
 a11247a <=( (not A170)  and  a11246a );
 a11250a <=( (not A201)  and  A166 );
 a11253a <=( (not A232)  and  A203 );
 a11254a <=( a11253a  and  a11250a );
 a11255a <=( a11254a  and  a11247a );
 a11259a <=( A235  and  A234 );
 a11260a <=( A233  and  a11259a );
 a11263a <=( (not A266)  and  A265 );
 a11266a <=( A269  and  A267 );
 a11267a <=( a11266a  and  a11263a );
 a11268a <=( a11267a  and  a11260a );
 a11272a <=( (not A167)  and  A168 );
 a11273a <=( (not A170)  and  a11272a );
 a11276a <=( (not A201)  and  A166 );
 a11279a <=( (not A232)  and  A203 );
 a11280a <=( a11279a  and  a11276a );
 a11281a <=( a11280a  and  a11273a );
 a11285a <=( A236  and  A234 );
 a11286a <=( A233  and  a11285a );
 a11289a <=( (not A299)  and  A298 );
 a11292a <=( A301  and  A300 );
 a11293a <=( a11292a  and  a11289a );
 a11294a <=( a11293a  and  a11286a );
 a11298a <=( (not A167)  and  A168 );
 a11299a <=( (not A170)  and  a11298a );
 a11302a <=( (not A201)  and  A166 );
 a11305a <=( (not A232)  and  A203 );
 a11306a <=( a11305a  and  a11302a );
 a11307a <=( a11306a  and  a11299a );
 a11311a <=( A236  and  A234 );
 a11312a <=( A233  and  a11311a );
 a11315a <=( (not A299)  and  A298 );
 a11318a <=( A302  and  A300 );
 a11319a <=( a11318a  and  a11315a );
 a11320a <=( a11319a  and  a11312a );
 a11324a <=( (not A167)  and  A168 );
 a11325a <=( (not A170)  and  a11324a );
 a11328a <=( (not A201)  and  A166 );
 a11331a <=( (not A232)  and  A203 );
 a11332a <=( a11331a  and  a11328a );
 a11333a <=( a11332a  and  a11325a );
 a11337a <=( A236  and  A234 );
 a11338a <=( A233  and  a11337a );
 a11341a <=( A299  and  (not A298) );
 a11344a <=( A301  and  A300 );
 a11345a <=( a11344a  and  a11341a );
 a11346a <=( a11345a  and  a11338a );
 a11350a <=( (not A167)  and  A168 );
 a11351a <=( (not A170)  and  a11350a );
 a11354a <=( (not A201)  and  A166 );
 a11357a <=( (not A232)  and  A203 );
 a11358a <=( a11357a  and  a11354a );
 a11359a <=( a11358a  and  a11351a );
 a11363a <=( A236  and  A234 );
 a11364a <=( A233  and  a11363a );
 a11367a <=( A299  and  (not A298) );
 a11370a <=( A302  and  A300 );
 a11371a <=( a11370a  and  a11367a );
 a11372a <=( a11371a  and  a11364a );
 a11376a <=( (not A167)  and  A168 );
 a11377a <=( (not A170)  and  a11376a );
 a11380a <=( (not A201)  and  A166 );
 a11383a <=( (not A232)  and  A203 );
 a11384a <=( a11383a  and  a11380a );
 a11385a <=( a11384a  and  a11377a );
 a11389a <=( A236  and  A234 );
 a11390a <=( A233  and  a11389a );
 a11393a <=( A266  and  (not A265) );
 a11396a <=( A268  and  A267 );
 a11397a <=( a11396a  and  a11393a );
 a11398a <=( a11397a  and  a11390a );
 a11402a <=( (not A167)  and  A168 );
 a11403a <=( (not A170)  and  a11402a );
 a11406a <=( (not A201)  and  A166 );
 a11409a <=( (not A232)  and  A203 );
 a11410a <=( a11409a  and  a11406a );
 a11411a <=( a11410a  and  a11403a );
 a11415a <=( A236  and  A234 );
 a11416a <=( A233  and  a11415a );
 a11419a <=( A266  and  (not A265) );
 a11422a <=( A269  and  A267 );
 a11423a <=( a11422a  and  a11419a );
 a11424a <=( a11423a  and  a11416a );
 a11428a <=( (not A167)  and  A168 );
 a11429a <=( (not A170)  and  a11428a );
 a11432a <=( (not A201)  and  A166 );
 a11435a <=( (not A232)  and  A203 );
 a11436a <=( a11435a  and  a11432a );
 a11437a <=( a11436a  and  a11429a );
 a11441a <=( A236  and  A234 );
 a11442a <=( A233  and  a11441a );
 a11445a <=( (not A266)  and  A265 );
 a11448a <=( A268  and  A267 );
 a11449a <=( a11448a  and  a11445a );
 a11450a <=( a11449a  and  a11442a );
 a11454a <=( (not A167)  and  A168 );
 a11455a <=( (not A170)  and  a11454a );
 a11458a <=( (not A201)  and  A166 );
 a11461a <=( (not A232)  and  A203 );
 a11462a <=( a11461a  and  a11458a );
 a11463a <=( a11462a  and  a11455a );
 a11467a <=( A236  and  A234 );
 a11468a <=( A233  and  a11467a );
 a11471a <=( (not A266)  and  A265 );
 a11474a <=( A269  and  A267 );
 a11475a <=( a11474a  and  a11471a );
 a11476a <=( a11475a  and  a11468a );
 a11480a <=( (not A167)  and  A168 );
 a11481a <=( (not A170)  and  a11480a );
 a11484a <=( (not A201)  and  A166 );
 a11487a <=( A232  and  A203 );
 a11488a <=( a11487a  and  a11484a );
 a11489a <=( a11488a  and  a11481a );
 a11493a <=( A235  and  A234 );
 a11494a <=( (not A233)  and  a11493a );
 a11497a <=( (not A299)  and  A298 );
 a11500a <=( A301  and  A300 );
 a11501a <=( a11500a  and  a11497a );
 a11502a <=( a11501a  and  a11494a );
 a11506a <=( (not A167)  and  A168 );
 a11507a <=( (not A170)  and  a11506a );
 a11510a <=( (not A201)  and  A166 );
 a11513a <=( A232  and  A203 );
 a11514a <=( a11513a  and  a11510a );
 a11515a <=( a11514a  and  a11507a );
 a11519a <=( A235  and  A234 );
 a11520a <=( (not A233)  and  a11519a );
 a11523a <=( (not A299)  and  A298 );
 a11526a <=( A302  and  A300 );
 a11527a <=( a11526a  and  a11523a );
 a11528a <=( a11527a  and  a11520a );
 a11532a <=( (not A167)  and  A168 );
 a11533a <=( (not A170)  and  a11532a );
 a11536a <=( (not A201)  and  A166 );
 a11539a <=( A232  and  A203 );
 a11540a <=( a11539a  and  a11536a );
 a11541a <=( a11540a  and  a11533a );
 a11545a <=( A235  and  A234 );
 a11546a <=( (not A233)  and  a11545a );
 a11549a <=( A299  and  (not A298) );
 a11552a <=( A301  and  A300 );
 a11553a <=( a11552a  and  a11549a );
 a11554a <=( a11553a  and  a11546a );
 a11558a <=( (not A167)  and  A168 );
 a11559a <=( (not A170)  and  a11558a );
 a11562a <=( (not A201)  and  A166 );
 a11565a <=( A232  and  A203 );
 a11566a <=( a11565a  and  a11562a );
 a11567a <=( a11566a  and  a11559a );
 a11571a <=( A235  and  A234 );
 a11572a <=( (not A233)  and  a11571a );
 a11575a <=( A299  and  (not A298) );
 a11578a <=( A302  and  A300 );
 a11579a <=( a11578a  and  a11575a );
 a11580a <=( a11579a  and  a11572a );
 a11584a <=( (not A167)  and  A168 );
 a11585a <=( (not A170)  and  a11584a );
 a11588a <=( (not A201)  and  A166 );
 a11591a <=( A232  and  A203 );
 a11592a <=( a11591a  and  a11588a );
 a11593a <=( a11592a  and  a11585a );
 a11597a <=( A235  and  A234 );
 a11598a <=( (not A233)  and  a11597a );
 a11601a <=( A266  and  (not A265) );
 a11604a <=( A268  and  A267 );
 a11605a <=( a11604a  and  a11601a );
 a11606a <=( a11605a  and  a11598a );
 a11610a <=( (not A167)  and  A168 );
 a11611a <=( (not A170)  and  a11610a );
 a11614a <=( (not A201)  and  A166 );
 a11617a <=( A232  and  A203 );
 a11618a <=( a11617a  and  a11614a );
 a11619a <=( a11618a  and  a11611a );
 a11623a <=( A235  and  A234 );
 a11624a <=( (not A233)  and  a11623a );
 a11627a <=( A266  and  (not A265) );
 a11630a <=( A269  and  A267 );
 a11631a <=( a11630a  and  a11627a );
 a11632a <=( a11631a  and  a11624a );
 a11636a <=( (not A167)  and  A168 );
 a11637a <=( (not A170)  and  a11636a );
 a11640a <=( (not A201)  and  A166 );
 a11643a <=( A232  and  A203 );
 a11644a <=( a11643a  and  a11640a );
 a11645a <=( a11644a  and  a11637a );
 a11649a <=( A235  and  A234 );
 a11650a <=( (not A233)  and  a11649a );
 a11653a <=( (not A266)  and  A265 );
 a11656a <=( A268  and  A267 );
 a11657a <=( a11656a  and  a11653a );
 a11658a <=( a11657a  and  a11650a );
 a11662a <=( (not A167)  and  A168 );
 a11663a <=( (not A170)  and  a11662a );
 a11666a <=( (not A201)  and  A166 );
 a11669a <=( A232  and  A203 );
 a11670a <=( a11669a  and  a11666a );
 a11671a <=( a11670a  and  a11663a );
 a11675a <=( A235  and  A234 );
 a11676a <=( (not A233)  and  a11675a );
 a11679a <=( (not A266)  and  A265 );
 a11682a <=( A269  and  A267 );
 a11683a <=( a11682a  and  a11679a );
 a11684a <=( a11683a  and  a11676a );
 a11688a <=( (not A167)  and  A168 );
 a11689a <=( (not A170)  and  a11688a );
 a11692a <=( (not A201)  and  A166 );
 a11695a <=( A232  and  A203 );
 a11696a <=( a11695a  and  a11692a );
 a11697a <=( a11696a  and  a11689a );
 a11701a <=( A236  and  A234 );
 a11702a <=( (not A233)  and  a11701a );
 a11705a <=( (not A299)  and  A298 );
 a11708a <=( A301  and  A300 );
 a11709a <=( a11708a  and  a11705a );
 a11710a <=( a11709a  and  a11702a );
 a11714a <=( (not A167)  and  A168 );
 a11715a <=( (not A170)  and  a11714a );
 a11718a <=( (not A201)  and  A166 );
 a11721a <=( A232  and  A203 );
 a11722a <=( a11721a  and  a11718a );
 a11723a <=( a11722a  and  a11715a );
 a11727a <=( A236  and  A234 );
 a11728a <=( (not A233)  and  a11727a );
 a11731a <=( (not A299)  and  A298 );
 a11734a <=( A302  and  A300 );
 a11735a <=( a11734a  and  a11731a );
 a11736a <=( a11735a  and  a11728a );
 a11740a <=( (not A167)  and  A168 );
 a11741a <=( (not A170)  and  a11740a );
 a11744a <=( (not A201)  and  A166 );
 a11747a <=( A232  and  A203 );
 a11748a <=( a11747a  and  a11744a );
 a11749a <=( a11748a  and  a11741a );
 a11753a <=( A236  and  A234 );
 a11754a <=( (not A233)  and  a11753a );
 a11757a <=( A299  and  (not A298) );
 a11760a <=( A301  and  A300 );
 a11761a <=( a11760a  and  a11757a );
 a11762a <=( a11761a  and  a11754a );
 a11766a <=( (not A167)  and  A168 );
 a11767a <=( (not A170)  and  a11766a );
 a11770a <=( (not A201)  and  A166 );
 a11773a <=( A232  and  A203 );
 a11774a <=( a11773a  and  a11770a );
 a11775a <=( a11774a  and  a11767a );
 a11779a <=( A236  and  A234 );
 a11780a <=( (not A233)  and  a11779a );
 a11783a <=( A299  and  (not A298) );
 a11786a <=( A302  and  A300 );
 a11787a <=( a11786a  and  a11783a );
 a11788a <=( a11787a  and  a11780a );
 a11792a <=( (not A167)  and  A168 );
 a11793a <=( (not A170)  and  a11792a );
 a11796a <=( (not A201)  and  A166 );
 a11799a <=( A232  and  A203 );
 a11800a <=( a11799a  and  a11796a );
 a11801a <=( a11800a  and  a11793a );
 a11805a <=( A236  and  A234 );
 a11806a <=( (not A233)  and  a11805a );
 a11809a <=( A266  and  (not A265) );
 a11812a <=( A268  and  A267 );
 a11813a <=( a11812a  and  a11809a );
 a11814a <=( a11813a  and  a11806a );
 a11818a <=( (not A167)  and  A168 );
 a11819a <=( (not A170)  and  a11818a );
 a11822a <=( (not A201)  and  A166 );
 a11825a <=( A232  and  A203 );
 a11826a <=( a11825a  and  a11822a );
 a11827a <=( a11826a  and  a11819a );
 a11831a <=( A236  and  A234 );
 a11832a <=( (not A233)  and  a11831a );
 a11835a <=( A266  and  (not A265) );
 a11838a <=( A269  and  A267 );
 a11839a <=( a11838a  and  a11835a );
 a11840a <=( a11839a  and  a11832a );
 a11844a <=( (not A167)  and  A168 );
 a11845a <=( (not A170)  and  a11844a );
 a11848a <=( (not A201)  and  A166 );
 a11851a <=( A232  and  A203 );
 a11852a <=( a11851a  and  a11848a );
 a11853a <=( a11852a  and  a11845a );
 a11857a <=( A236  and  A234 );
 a11858a <=( (not A233)  and  a11857a );
 a11861a <=( (not A266)  and  A265 );
 a11864a <=( A268  and  A267 );
 a11865a <=( a11864a  and  a11861a );
 a11866a <=( a11865a  and  a11858a );
 a11870a <=( (not A167)  and  A168 );
 a11871a <=( (not A170)  and  a11870a );
 a11874a <=( (not A201)  and  A166 );
 a11877a <=( A232  and  A203 );
 a11878a <=( a11877a  and  a11874a );
 a11879a <=( a11878a  and  a11871a );
 a11883a <=( A236  and  A234 );
 a11884a <=( (not A233)  and  a11883a );
 a11887a <=( (not A266)  and  A265 );
 a11890a <=( A269  and  A267 );
 a11891a <=( a11890a  and  a11887a );
 a11892a <=( a11891a  and  a11884a );
 a11896a <=( (not A167)  and  A168 );
 a11897a <=( (not A170)  and  a11896a );
 a11900a <=( A199  and  A166 );
 a11903a <=( (not A232)  and  A200 );
 a11904a <=( a11903a  and  a11900a );
 a11905a <=( a11904a  and  a11897a );
 a11909a <=( A235  and  A234 );
 a11910a <=( A233  and  a11909a );
 a11913a <=( (not A299)  and  A298 );
 a11916a <=( A301  and  A300 );
 a11917a <=( a11916a  and  a11913a );
 a11918a <=( a11917a  and  a11910a );
 a11922a <=( (not A167)  and  A168 );
 a11923a <=( (not A170)  and  a11922a );
 a11926a <=( A199  and  A166 );
 a11929a <=( (not A232)  and  A200 );
 a11930a <=( a11929a  and  a11926a );
 a11931a <=( a11930a  and  a11923a );
 a11935a <=( A235  and  A234 );
 a11936a <=( A233  and  a11935a );
 a11939a <=( (not A299)  and  A298 );
 a11942a <=( A302  and  A300 );
 a11943a <=( a11942a  and  a11939a );
 a11944a <=( a11943a  and  a11936a );
 a11948a <=( (not A167)  and  A168 );
 a11949a <=( (not A170)  and  a11948a );
 a11952a <=( A199  and  A166 );
 a11955a <=( (not A232)  and  A200 );
 a11956a <=( a11955a  and  a11952a );
 a11957a <=( a11956a  and  a11949a );
 a11961a <=( A235  and  A234 );
 a11962a <=( A233  and  a11961a );
 a11965a <=( A299  and  (not A298) );
 a11968a <=( A301  and  A300 );
 a11969a <=( a11968a  and  a11965a );
 a11970a <=( a11969a  and  a11962a );
 a11974a <=( (not A167)  and  A168 );
 a11975a <=( (not A170)  and  a11974a );
 a11978a <=( A199  and  A166 );
 a11981a <=( (not A232)  and  A200 );
 a11982a <=( a11981a  and  a11978a );
 a11983a <=( a11982a  and  a11975a );
 a11987a <=( A235  and  A234 );
 a11988a <=( A233  and  a11987a );
 a11991a <=( A299  and  (not A298) );
 a11994a <=( A302  and  A300 );
 a11995a <=( a11994a  and  a11991a );
 a11996a <=( a11995a  and  a11988a );
 a12000a <=( (not A167)  and  A168 );
 a12001a <=( (not A170)  and  a12000a );
 a12004a <=( A199  and  A166 );
 a12007a <=( (not A232)  and  A200 );
 a12008a <=( a12007a  and  a12004a );
 a12009a <=( a12008a  and  a12001a );
 a12013a <=( A235  and  A234 );
 a12014a <=( A233  and  a12013a );
 a12017a <=( A266  and  (not A265) );
 a12020a <=( A268  and  A267 );
 a12021a <=( a12020a  and  a12017a );
 a12022a <=( a12021a  and  a12014a );
 a12026a <=( (not A167)  and  A168 );
 a12027a <=( (not A170)  and  a12026a );
 a12030a <=( A199  and  A166 );
 a12033a <=( (not A232)  and  A200 );
 a12034a <=( a12033a  and  a12030a );
 a12035a <=( a12034a  and  a12027a );
 a12039a <=( A235  and  A234 );
 a12040a <=( A233  and  a12039a );
 a12043a <=( A266  and  (not A265) );
 a12046a <=( A269  and  A267 );
 a12047a <=( a12046a  and  a12043a );
 a12048a <=( a12047a  and  a12040a );
 a12052a <=( (not A167)  and  A168 );
 a12053a <=( (not A170)  and  a12052a );
 a12056a <=( A199  and  A166 );
 a12059a <=( (not A232)  and  A200 );
 a12060a <=( a12059a  and  a12056a );
 a12061a <=( a12060a  and  a12053a );
 a12065a <=( A235  and  A234 );
 a12066a <=( A233  and  a12065a );
 a12069a <=( (not A266)  and  A265 );
 a12072a <=( A268  and  A267 );
 a12073a <=( a12072a  and  a12069a );
 a12074a <=( a12073a  and  a12066a );
 a12078a <=( (not A167)  and  A168 );
 a12079a <=( (not A170)  and  a12078a );
 a12082a <=( A199  and  A166 );
 a12085a <=( (not A232)  and  A200 );
 a12086a <=( a12085a  and  a12082a );
 a12087a <=( a12086a  and  a12079a );
 a12091a <=( A235  and  A234 );
 a12092a <=( A233  and  a12091a );
 a12095a <=( (not A266)  and  A265 );
 a12098a <=( A269  and  A267 );
 a12099a <=( a12098a  and  a12095a );
 a12100a <=( a12099a  and  a12092a );
 a12104a <=( (not A167)  and  A168 );
 a12105a <=( (not A170)  and  a12104a );
 a12108a <=( A199  and  A166 );
 a12111a <=( (not A232)  and  A200 );
 a12112a <=( a12111a  and  a12108a );
 a12113a <=( a12112a  and  a12105a );
 a12117a <=( A236  and  A234 );
 a12118a <=( A233  and  a12117a );
 a12121a <=( (not A299)  and  A298 );
 a12124a <=( A301  and  A300 );
 a12125a <=( a12124a  and  a12121a );
 a12126a <=( a12125a  and  a12118a );
 a12130a <=( (not A167)  and  A168 );
 a12131a <=( (not A170)  and  a12130a );
 a12134a <=( A199  and  A166 );
 a12137a <=( (not A232)  and  A200 );
 a12138a <=( a12137a  and  a12134a );
 a12139a <=( a12138a  and  a12131a );
 a12143a <=( A236  and  A234 );
 a12144a <=( A233  and  a12143a );
 a12147a <=( (not A299)  and  A298 );
 a12150a <=( A302  and  A300 );
 a12151a <=( a12150a  and  a12147a );
 a12152a <=( a12151a  and  a12144a );
 a12156a <=( (not A167)  and  A168 );
 a12157a <=( (not A170)  and  a12156a );
 a12160a <=( A199  and  A166 );
 a12163a <=( (not A232)  and  A200 );
 a12164a <=( a12163a  and  a12160a );
 a12165a <=( a12164a  and  a12157a );
 a12169a <=( A236  and  A234 );
 a12170a <=( A233  and  a12169a );
 a12173a <=( A299  and  (not A298) );
 a12176a <=( A301  and  A300 );
 a12177a <=( a12176a  and  a12173a );
 a12178a <=( a12177a  and  a12170a );
 a12182a <=( (not A167)  and  A168 );
 a12183a <=( (not A170)  and  a12182a );
 a12186a <=( A199  and  A166 );
 a12189a <=( (not A232)  and  A200 );
 a12190a <=( a12189a  and  a12186a );
 a12191a <=( a12190a  and  a12183a );
 a12195a <=( A236  and  A234 );
 a12196a <=( A233  and  a12195a );
 a12199a <=( A299  and  (not A298) );
 a12202a <=( A302  and  A300 );
 a12203a <=( a12202a  and  a12199a );
 a12204a <=( a12203a  and  a12196a );
 a12208a <=( (not A167)  and  A168 );
 a12209a <=( (not A170)  and  a12208a );
 a12212a <=( A199  and  A166 );
 a12215a <=( (not A232)  and  A200 );
 a12216a <=( a12215a  and  a12212a );
 a12217a <=( a12216a  and  a12209a );
 a12221a <=( A236  and  A234 );
 a12222a <=( A233  and  a12221a );
 a12225a <=( A266  and  (not A265) );
 a12228a <=( A268  and  A267 );
 a12229a <=( a12228a  and  a12225a );
 a12230a <=( a12229a  and  a12222a );
 a12234a <=( (not A167)  and  A168 );
 a12235a <=( (not A170)  and  a12234a );
 a12238a <=( A199  and  A166 );
 a12241a <=( (not A232)  and  A200 );
 a12242a <=( a12241a  and  a12238a );
 a12243a <=( a12242a  and  a12235a );
 a12247a <=( A236  and  A234 );
 a12248a <=( A233  and  a12247a );
 a12251a <=( A266  and  (not A265) );
 a12254a <=( A269  and  A267 );
 a12255a <=( a12254a  and  a12251a );
 a12256a <=( a12255a  and  a12248a );
 a12260a <=( (not A167)  and  A168 );
 a12261a <=( (not A170)  and  a12260a );
 a12264a <=( A199  and  A166 );
 a12267a <=( (not A232)  and  A200 );
 a12268a <=( a12267a  and  a12264a );
 a12269a <=( a12268a  and  a12261a );
 a12273a <=( A236  and  A234 );
 a12274a <=( A233  and  a12273a );
 a12277a <=( (not A266)  and  A265 );
 a12280a <=( A268  and  A267 );
 a12281a <=( a12280a  and  a12277a );
 a12282a <=( a12281a  and  a12274a );
 a12286a <=( (not A167)  and  A168 );
 a12287a <=( (not A170)  and  a12286a );
 a12290a <=( A199  and  A166 );
 a12293a <=( (not A232)  and  A200 );
 a12294a <=( a12293a  and  a12290a );
 a12295a <=( a12294a  and  a12287a );
 a12299a <=( A236  and  A234 );
 a12300a <=( A233  and  a12299a );
 a12303a <=( (not A266)  and  A265 );
 a12306a <=( A269  and  A267 );
 a12307a <=( a12306a  and  a12303a );
 a12308a <=( a12307a  and  a12300a );
 a12312a <=( (not A167)  and  A168 );
 a12313a <=( (not A170)  and  a12312a );
 a12316a <=( A199  and  A166 );
 a12319a <=( A232  and  A200 );
 a12320a <=( a12319a  and  a12316a );
 a12321a <=( a12320a  and  a12313a );
 a12325a <=( A235  and  A234 );
 a12326a <=( (not A233)  and  a12325a );
 a12329a <=( (not A299)  and  A298 );
 a12332a <=( A301  and  A300 );
 a12333a <=( a12332a  and  a12329a );
 a12334a <=( a12333a  and  a12326a );
 a12338a <=( (not A167)  and  A168 );
 a12339a <=( (not A170)  and  a12338a );
 a12342a <=( A199  and  A166 );
 a12345a <=( A232  and  A200 );
 a12346a <=( a12345a  and  a12342a );
 a12347a <=( a12346a  and  a12339a );
 a12351a <=( A235  and  A234 );
 a12352a <=( (not A233)  and  a12351a );
 a12355a <=( (not A299)  and  A298 );
 a12358a <=( A302  and  A300 );
 a12359a <=( a12358a  and  a12355a );
 a12360a <=( a12359a  and  a12352a );
 a12364a <=( (not A167)  and  A168 );
 a12365a <=( (not A170)  and  a12364a );
 a12368a <=( A199  and  A166 );
 a12371a <=( A232  and  A200 );
 a12372a <=( a12371a  and  a12368a );
 a12373a <=( a12372a  and  a12365a );
 a12377a <=( A235  and  A234 );
 a12378a <=( (not A233)  and  a12377a );
 a12381a <=( A299  and  (not A298) );
 a12384a <=( A301  and  A300 );
 a12385a <=( a12384a  and  a12381a );
 a12386a <=( a12385a  and  a12378a );
 a12390a <=( (not A167)  and  A168 );
 a12391a <=( (not A170)  and  a12390a );
 a12394a <=( A199  and  A166 );
 a12397a <=( A232  and  A200 );
 a12398a <=( a12397a  and  a12394a );
 a12399a <=( a12398a  and  a12391a );
 a12403a <=( A235  and  A234 );
 a12404a <=( (not A233)  and  a12403a );
 a12407a <=( A299  and  (not A298) );
 a12410a <=( A302  and  A300 );
 a12411a <=( a12410a  and  a12407a );
 a12412a <=( a12411a  and  a12404a );
 a12416a <=( (not A167)  and  A168 );
 a12417a <=( (not A170)  and  a12416a );
 a12420a <=( A199  and  A166 );
 a12423a <=( A232  and  A200 );
 a12424a <=( a12423a  and  a12420a );
 a12425a <=( a12424a  and  a12417a );
 a12429a <=( A235  and  A234 );
 a12430a <=( (not A233)  and  a12429a );
 a12433a <=( A266  and  (not A265) );
 a12436a <=( A268  and  A267 );
 a12437a <=( a12436a  and  a12433a );
 a12438a <=( a12437a  and  a12430a );
 a12442a <=( (not A167)  and  A168 );
 a12443a <=( (not A170)  and  a12442a );
 a12446a <=( A199  and  A166 );
 a12449a <=( A232  and  A200 );
 a12450a <=( a12449a  and  a12446a );
 a12451a <=( a12450a  and  a12443a );
 a12455a <=( A235  and  A234 );
 a12456a <=( (not A233)  and  a12455a );
 a12459a <=( A266  and  (not A265) );
 a12462a <=( A269  and  A267 );
 a12463a <=( a12462a  and  a12459a );
 a12464a <=( a12463a  and  a12456a );
 a12468a <=( (not A167)  and  A168 );
 a12469a <=( (not A170)  and  a12468a );
 a12472a <=( A199  and  A166 );
 a12475a <=( A232  and  A200 );
 a12476a <=( a12475a  and  a12472a );
 a12477a <=( a12476a  and  a12469a );
 a12481a <=( A235  and  A234 );
 a12482a <=( (not A233)  and  a12481a );
 a12485a <=( (not A266)  and  A265 );
 a12488a <=( A268  and  A267 );
 a12489a <=( a12488a  and  a12485a );
 a12490a <=( a12489a  and  a12482a );
 a12494a <=( (not A167)  and  A168 );
 a12495a <=( (not A170)  and  a12494a );
 a12498a <=( A199  and  A166 );
 a12501a <=( A232  and  A200 );
 a12502a <=( a12501a  and  a12498a );
 a12503a <=( a12502a  and  a12495a );
 a12507a <=( A235  and  A234 );
 a12508a <=( (not A233)  and  a12507a );
 a12511a <=( (not A266)  and  A265 );
 a12514a <=( A269  and  A267 );
 a12515a <=( a12514a  and  a12511a );
 a12516a <=( a12515a  and  a12508a );
 a12520a <=( (not A167)  and  A168 );
 a12521a <=( (not A170)  and  a12520a );
 a12524a <=( A199  and  A166 );
 a12527a <=( A232  and  A200 );
 a12528a <=( a12527a  and  a12524a );
 a12529a <=( a12528a  and  a12521a );
 a12533a <=( A236  and  A234 );
 a12534a <=( (not A233)  and  a12533a );
 a12537a <=( (not A299)  and  A298 );
 a12540a <=( A301  and  A300 );
 a12541a <=( a12540a  and  a12537a );
 a12542a <=( a12541a  and  a12534a );
 a12546a <=( (not A167)  and  A168 );
 a12547a <=( (not A170)  and  a12546a );
 a12550a <=( A199  and  A166 );
 a12553a <=( A232  and  A200 );
 a12554a <=( a12553a  and  a12550a );
 a12555a <=( a12554a  and  a12547a );
 a12559a <=( A236  and  A234 );
 a12560a <=( (not A233)  and  a12559a );
 a12563a <=( (not A299)  and  A298 );
 a12566a <=( A302  and  A300 );
 a12567a <=( a12566a  and  a12563a );
 a12568a <=( a12567a  and  a12560a );
 a12572a <=( (not A167)  and  A168 );
 a12573a <=( (not A170)  and  a12572a );
 a12576a <=( A199  and  A166 );
 a12579a <=( A232  and  A200 );
 a12580a <=( a12579a  and  a12576a );
 a12581a <=( a12580a  and  a12573a );
 a12585a <=( A236  and  A234 );
 a12586a <=( (not A233)  and  a12585a );
 a12589a <=( A299  and  (not A298) );
 a12592a <=( A301  and  A300 );
 a12593a <=( a12592a  and  a12589a );
 a12594a <=( a12593a  and  a12586a );
 a12598a <=( (not A167)  and  A168 );
 a12599a <=( (not A170)  and  a12598a );
 a12602a <=( A199  and  A166 );
 a12605a <=( A232  and  A200 );
 a12606a <=( a12605a  and  a12602a );
 a12607a <=( a12606a  and  a12599a );
 a12611a <=( A236  and  A234 );
 a12612a <=( (not A233)  and  a12611a );
 a12615a <=( A299  and  (not A298) );
 a12618a <=( A302  and  A300 );
 a12619a <=( a12618a  and  a12615a );
 a12620a <=( a12619a  and  a12612a );
 a12624a <=( (not A167)  and  A168 );
 a12625a <=( (not A170)  and  a12624a );
 a12628a <=( A199  and  A166 );
 a12631a <=( A232  and  A200 );
 a12632a <=( a12631a  and  a12628a );
 a12633a <=( a12632a  and  a12625a );
 a12637a <=( A236  and  A234 );
 a12638a <=( (not A233)  and  a12637a );
 a12641a <=( A266  and  (not A265) );
 a12644a <=( A268  and  A267 );
 a12645a <=( a12644a  and  a12641a );
 a12646a <=( a12645a  and  a12638a );
 a12650a <=( (not A167)  and  A168 );
 a12651a <=( (not A170)  and  a12650a );
 a12654a <=( A199  and  A166 );
 a12657a <=( A232  and  A200 );
 a12658a <=( a12657a  and  a12654a );
 a12659a <=( a12658a  and  a12651a );
 a12663a <=( A236  and  A234 );
 a12664a <=( (not A233)  and  a12663a );
 a12667a <=( A266  and  (not A265) );
 a12670a <=( A269  and  A267 );
 a12671a <=( a12670a  and  a12667a );
 a12672a <=( a12671a  and  a12664a );
 a12676a <=( (not A167)  and  A168 );
 a12677a <=( (not A170)  and  a12676a );
 a12680a <=( A199  and  A166 );
 a12683a <=( A232  and  A200 );
 a12684a <=( a12683a  and  a12680a );
 a12685a <=( a12684a  and  a12677a );
 a12689a <=( A236  and  A234 );
 a12690a <=( (not A233)  and  a12689a );
 a12693a <=( (not A266)  and  A265 );
 a12696a <=( A268  and  A267 );
 a12697a <=( a12696a  and  a12693a );
 a12698a <=( a12697a  and  a12690a );
 a12702a <=( (not A167)  and  A168 );
 a12703a <=( (not A170)  and  a12702a );
 a12706a <=( A199  and  A166 );
 a12709a <=( A232  and  A200 );
 a12710a <=( a12709a  and  a12706a );
 a12711a <=( a12710a  and  a12703a );
 a12715a <=( A236  and  A234 );
 a12716a <=( (not A233)  and  a12715a );
 a12719a <=( (not A266)  and  A265 );
 a12722a <=( A269  and  A267 );
 a12723a <=( a12722a  and  a12719a );
 a12724a <=( a12723a  and  a12716a );
 a12728a <=( (not A167)  and  A168 );
 a12729a <=( (not A170)  and  a12728a );
 a12732a <=( (not A199)  and  A166 );
 a12735a <=( (not A232)  and  (not A200) );
 a12736a <=( a12735a  and  a12732a );
 a12737a <=( a12736a  and  a12729a );
 a12741a <=( A235  and  A234 );
 a12742a <=( A233  and  a12741a );
 a12745a <=( (not A299)  and  A298 );
 a12748a <=( A301  and  A300 );
 a12749a <=( a12748a  and  a12745a );
 a12750a <=( a12749a  and  a12742a );
 a12754a <=( (not A167)  and  A168 );
 a12755a <=( (not A170)  and  a12754a );
 a12758a <=( (not A199)  and  A166 );
 a12761a <=( (not A232)  and  (not A200) );
 a12762a <=( a12761a  and  a12758a );
 a12763a <=( a12762a  and  a12755a );
 a12767a <=( A235  and  A234 );
 a12768a <=( A233  and  a12767a );
 a12771a <=( (not A299)  and  A298 );
 a12774a <=( A302  and  A300 );
 a12775a <=( a12774a  and  a12771a );
 a12776a <=( a12775a  and  a12768a );
 a12780a <=( (not A167)  and  A168 );
 a12781a <=( (not A170)  and  a12780a );
 a12784a <=( (not A199)  and  A166 );
 a12787a <=( (not A232)  and  (not A200) );
 a12788a <=( a12787a  and  a12784a );
 a12789a <=( a12788a  and  a12781a );
 a12793a <=( A235  and  A234 );
 a12794a <=( A233  and  a12793a );
 a12797a <=( A299  and  (not A298) );
 a12800a <=( A301  and  A300 );
 a12801a <=( a12800a  and  a12797a );
 a12802a <=( a12801a  and  a12794a );
 a12806a <=( (not A167)  and  A168 );
 a12807a <=( (not A170)  and  a12806a );
 a12810a <=( (not A199)  and  A166 );
 a12813a <=( (not A232)  and  (not A200) );
 a12814a <=( a12813a  and  a12810a );
 a12815a <=( a12814a  and  a12807a );
 a12819a <=( A235  and  A234 );
 a12820a <=( A233  and  a12819a );
 a12823a <=( A299  and  (not A298) );
 a12826a <=( A302  and  A300 );
 a12827a <=( a12826a  and  a12823a );
 a12828a <=( a12827a  and  a12820a );
 a12832a <=( (not A167)  and  A168 );
 a12833a <=( (not A170)  and  a12832a );
 a12836a <=( (not A199)  and  A166 );
 a12839a <=( (not A232)  and  (not A200) );
 a12840a <=( a12839a  and  a12836a );
 a12841a <=( a12840a  and  a12833a );
 a12845a <=( A235  and  A234 );
 a12846a <=( A233  and  a12845a );
 a12849a <=( A266  and  (not A265) );
 a12852a <=( A268  and  A267 );
 a12853a <=( a12852a  and  a12849a );
 a12854a <=( a12853a  and  a12846a );
 a12858a <=( (not A167)  and  A168 );
 a12859a <=( (not A170)  and  a12858a );
 a12862a <=( (not A199)  and  A166 );
 a12865a <=( (not A232)  and  (not A200) );
 a12866a <=( a12865a  and  a12862a );
 a12867a <=( a12866a  and  a12859a );
 a12871a <=( A235  and  A234 );
 a12872a <=( A233  and  a12871a );
 a12875a <=( A266  and  (not A265) );
 a12878a <=( A269  and  A267 );
 a12879a <=( a12878a  and  a12875a );
 a12880a <=( a12879a  and  a12872a );
 a12884a <=( (not A167)  and  A168 );
 a12885a <=( (not A170)  and  a12884a );
 a12888a <=( (not A199)  and  A166 );
 a12891a <=( (not A232)  and  (not A200) );
 a12892a <=( a12891a  and  a12888a );
 a12893a <=( a12892a  and  a12885a );
 a12897a <=( A235  and  A234 );
 a12898a <=( A233  and  a12897a );
 a12901a <=( (not A266)  and  A265 );
 a12904a <=( A268  and  A267 );
 a12905a <=( a12904a  and  a12901a );
 a12906a <=( a12905a  and  a12898a );
 a12910a <=( (not A167)  and  A168 );
 a12911a <=( (not A170)  and  a12910a );
 a12914a <=( (not A199)  and  A166 );
 a12917a <=( (not A232)  and  (not A200) );
 a12918a <=( a12917a  and  a12914a );
 a12919a <=( a12918a  and  a12911a );
 a12923a <=( A235  and  A234 );
 a12924a <=( A233  and  a12923a );
 a12927a <=( (not A266)  and  A265 );
 a12930a <=( A269  and  A267 );
 a12931a <=( a12930a  and  a12927a );
 a12932a <=( a12931a  and  a12924a );
 a12936a <=( (not A167)  and  A168 );
 a12937a <=( (not A170)  and  a12936a );
 a12940a <=( (not A199)  and  A166 );
 a12943a <=( (not A232)  and  (not A200) );
 a12944a <=( a12943a  and  a12940a );
 a12945a <=( a12944a  and  a12937a );
 a12949a <=( A236  and  A234 );
 a12950a <=( A233  and  a12949a );
 a12953a <=( (not A299)  and  A298 );
 a12956a <=( A301  and  A300 );
 a12957a <=( a12956a  and  a12953a );
 a12958a <=( a12957a  and  a12950a );
 a12962a <=( (not A167)  and  A168 );
 a12963a <=( (not A170)  and  a12962a );
 a12966a <=( (not A199)  and  A166 );
 a12969a <=( (not A232)  and  (not A200) );
 a12970a <=( a12969a  and  a12966a );
 a12971a <=( a12970a  and  a12963a );
 a12975a <=( A236  and  A234 );
 a12976a <=( A233  and  a12975a );
 a12979a <=( (not A299)  and  A298 );
 a12982a <=( A302  and  A300 );
 a12983a <=( a12982a  and  a12979a );
 a12984a <=( a12983a  and  a12976a );
 a12988a <=( (not A167)  and  A168 );
 a12989a <=( (not A170)  and  a12988a );
 a12992a <=( (not A199)  and  A166 );
 a12995a <=( (not A232)  and  (not A200) );
 a12996a <=( a12995a  and  a12992a );
 a12997a <=( a12996a  and  a12989a );
 a13001a <=( A236  and  A234 );
 a13002a <=( A233  and  a13001a );
 a13005a <=( A299  and  (not A298) );
 a13008a <=( A301  and  A300 );
 a13009a <=( a13008a  and  a13005a );
 a13010a <=( a13009a  and  a13002a );
 a13014a <=( (not A167)  and  A168 );
 a13015a <=( (not A170)  and  a13014a );
 a13018a <=( (not A199)  and  A166 );
 a13021a <=( (not A232)  and  (not A200) );
 a13022a <=( a13021a  and  a13018a );
 a13023a <=( a13022a  and  a13015a );
 a13027a <=( A236  and  A234 );
 a13028a <=( A233  and  a13027a );
 a13031a <=( A299  and  (not A298) );
 a13034a <=( A302  and  A300 );
 a13035a <=( a13034a  and  a13031a );
 a13036a <=( a13035a  and  a13028a );
 a13040a <=( (not A167)  and  A168 );
 a13041a <=( (not A170)  and  a13040a );
 a13044a <=( (not A199)  and  A166 );
 a13047a <=( (not A232)  and  (not A200) );
 a13048a <=( a13047a  and  a13044a );
 a13049a <=( a13048a  and  a13041a );
 a13053a <=( A236  and  A234 );
 a13054a <=( A233  and  a13053a );
 a13057a <=( A266  and  (not A265) );
 a13060a <=( A268  and  A267 );
 a13061a <=( a13060a  and  a13057a );
 a13062a <=( a13061a  and  a13054a );
 a13066a <=( (not A167)  and  A168 );
 a13067a <=( (not A170)  and  a13066a );
 a13070a <=( (not A199)  and  A166 );
 a13073a <=( (not A232)  and  (not A200) );
 a13074a <=( a13073a  and  a13070a );
 a13075a <=( a13074a  and  a13067a );
 a13079a <=( A236  and  A234 );
 a13080a <=( A233  and  a13079a );
 a13083a <=( A266  and  (not A265) );
 a13086a <=( A269  and  A267 );
 a13087a <=( a13086a  and  a13083a );
 a13088a <=( a13087a  and  a13080a );
 a13092a <=( (not A167)  and  A168 );
 a13093a <=( (not A170)  and  a13092a );
 a13096a <=( (not A199)  and  A166 );
 a13099a <=( (not A232)  and  (not A200) );
 a13100a <=( a13099a  and  a13096a );
 a13101a <=( a13100a  and  a13093a );
 a13105a <=( A236  and  A234 );
 a13106a <=( A233  and  a13105a );
 a13109a <=( (not A266)  and  A265 );
 a13112a <=( A268  and  A267 );
 a13113a <=( a13112a  and  a13109a );
 a13114a <=( a13113a  and  a13106a );
 a13118a <=( (not A167)  and  A168 );
 a13119a <=( (not A170)  and  a13118a );
 a13122a <=( (not A199)  and  A166 );
 a13125a <=( (not A232)  and  (not A200) );
 a13126a <=( a13125a  and  a13122a );
 a13127a <=( a13126a  and  a13119a );
 a13131a <=( A236  and  A234 );
 a13132a <=( A233  and  a13131a );
 a13135a <=( (not A266)  and  A265 );
 a13138a <=( A269  and  A267 );
 a13139a <=( a13138a  and  a13135a );
 a13140a <=( a13139a  and  a13132a );
 a13144a <=( (not A167)  and  A168 );
 a13145a <=( (not A170)  and  a13144a );
 a13148a <=( (not A199)  and  A166 );
 a13151a <=( A232  and  (not A200) );
 a13152a <=( a13151a  and  a13148a );
 a13153a <=( a13152a  and  a13145a );
 a13157a <=( A235  and  A234 );
 a13158a <=( (not A233)  and  a13157a );
 a13161a <=( (not A299)  and  A298 );
 a13164a <=( A301  and  A300 );
 a13165a <=( a13164a  and  a13161a );
 a13166a <=( a13165a  and  a13158a );
 a13170a <=( (not A167)  and  A168 );
 a13171a <=( (not A170)  and  a13170a );
 a13174a <=( (not A199)  and  A166 );
 a13177a <=( A232  and  (not A200) );
 a13178a <=( a13177a  and  a13174a );
 a13179a <=( a13178a  and  a13171a );
 a13183a <=( A235  and  A234 );
 a13184a <=( (not A233)  and  a13183a );
 a13187a <=( (not A299)  and  A298 );
 a13190a <=( A302  and  A300 );
 a13191a <=( a13190a  and  a13187a );
 a13192a <=( a13191a  and  a13184a );
 a13196a <=( (not A167)  and  A168 );
 a13197a <=( (not A170)  and  a13196a );
 a13200a <=( (not A199)  and  A166 );
 a13203a <=( A232  and  (not A200) );
 a13204a <=( a13203a  and  a13200a );
 a13205a <=( a13204a  and  a13197a );
 a13209a <=( A235  and  A234 );
 a13210a <=( (not A233)  and  a13209a );
 a13213a <=( A299  and  (not A298) );
 a13216a <=( A301  and  A300 );
 a13217a <=( a13216a  and  a13213a );
 a13218a <=( a13217a  and  a13210a );
 a13222a <=( (not A167)  and  A168 );
 a13223a <=( (not A170)  and  a13222a );
 a13226a <=( (not A199)  and  A166 );
 a13229a <=( A232  and  (not A200) );
 a13230a <=( a13229a  and  a13226a );
 a13231a <=( a13230a  and  a13223a );
 a13235a <=( A235  and  A234 );
 a13236a <=( (not A233)  and  a13235a );
 a13239a <=( A299  and  (not A298) );
 a13242a <=( A302  and  A300 );
 a13243a <=( a13242a  and  a13239a );
 a13244a <=( a13243a  and  a13236a );
 a13248a <=( (not A167)  and  A168 );
 a13249a <=( (not A170)  and  a13248a );
 a13252a <=( (not A199)  and  A166 );
 a13255a <=( A232  and  (not A200) );
 a13256a <=( a13255a  and  a13252a );
 a13257a <=( a13256a  and  a13249a );
 a13261a <=( A235  and  A234 );
 a13262a <=( (not A233)  and  a13261a );
 a13265a <=( A266  and  (not A265) );
 a13268a <=( A268  and  A267 );
 a13269a <=( a13268a  and  a13265a );
 a13270a <=( a13269a  and  a13262a );
 a13274a <=( (not A167)  and  A168 );
 a13275a <=( (not A170)  and  a13274a );
 a13278a <=( (not A199)  and  A166 );
 a13281a <=( A232  and  (not A200) );
 a13282a <=( a13281a  and  a13278a );
 a13283a <=( a13282a  and  a13275a );
 a13287a <=( A235  and  A234 );
 a13288a <=( (not A233)  and  a13287a );
 a13291a <=( A266  and  (not A265) );
 a13294a <=( A269  and  A267 );
 a13295a <=( a13294a  and  a13291a );
 a13296a <=( a13295a  and  a13288a );
 a13300a <=( (not A167)  and  A168 );
 a13301a <=( (not A170)  and  a13300a );
 a13304a <=( (not A199)  and  A166 );
 a13307a <=( A232  and  (not A200) );
 a13308a <=( a13307a  and  a13304a );
 a13309a <=( a13308a  and  a13301a );
 a13313a <=( A235  and  A234 );
 a13314a <=( (not A233)  and  a13313a );
 a13317a <=( (not A266)  and  A265 );
 a13320a <=( A268  and  A267 );
 a13321a <=( a13320a  and  a13317a );
 a13322a <=( a13321a  and  a13314a );
 a13326a <=( (not A167)  and  A168 );
 a13327a <=( (not A170)  and  a13326a );
 a13330a <=( (not A199)  and  A166 );
 a13333a <=( A232  and  (not A200) );
 a13334a <=( a13333a  and  a13330a );
 a13335a <=( a13334a  and  a13327a );
 a13339a <=( A235  and  A234 );
 a13340a <=( (not A233)  and  a13339a );
 a13343a <=( (not A266)  and  A265 );
 a13346a <=( A269  and  A267 );
 a13347a <=( a13346a  and  a13343a );
 a13348a <=( a13347a  and  a13340a );
 a13352a <=( (not A167)  and  A168 );
 a13353a <=( (not A170)  and  a13352a );
 a13356a <=( (not A199)  and  A166 );
 a13359a <=( A232  and  (not A200) );
 a13360a <=( a13359a  and  a13356a );
 a13361a <=( a13360a  and  a13353a );
 a13365a <=( A236  and  A234 );
 a13366a <=( (not A233)  and  a13365a );
 a13369a <=( (not A299)  and  A298 );
 a13372a <=( A301  and  A300 );
 a13373a <=( a13372a  and  a13369a );
 a13374a <=( a13373a  and  a13366a );
 a13378a <=( (not A167)  and  A168 );
 a13379a <=( (not A170)  and  a13378a );
 a13382a <=( (not A199)  and  A166 );
 a13385a <=( A232  and  (not A200) );
 a13386a <=( a13385a  and  a13382a );
 a13387a <=( a13386a  and  a13379a );
 a13391a <=( A236  and  A234 );
 a13392a <=( (not A233)  and  a13391a );
 a13395a <=( (not A299)  and  A298 );
 a13398a <=( A302  and  A300 );
 a13399a <=( a13398a  and  a13395a );
 a13400a <=( a13399a  and  a13392a );
 a13404a <=( (not A167)  and  A168 );
 a13405a <=( (not A170)  and  a13404a );
 a13408a <=( (not A199)  and  A166 );
 a13411a <=( A232  and  (not A200) );
 a13412a <=( a13411a  and  a13408a );
 a13413a <=( a13412a  and  a13405a );
 a13417a <=( A236  and  A234 );
 a13418a <=( (not A233)  and  a13417a );
 a13421a <=( A299  and  (not A298) );
 a13424a <=( A301  and  A300 );
 a13425a <=( a13424a  and  a13421a );
 a13426a <=( a13425a  and  a13418a );
 a13430a <=( (not A167)  and  A168 );
 a13431a <=( (not A170)  and  a13430a );
 a13434a <=( (not A199)  and  A166 );
 a13437a <=( A232  and  (not A200) );
 a13438a <=( a13437a  and  a13434a );
 a13439a <=( a13438a  and  a13431a );
 a13443a <=( A236  and  A234 );
 a13444a <=( (not A233)  and  a13443a );
 a13447a <=( A299  and  (not A298) );
 a13450a <=( A302  and  A300 );
 a13451a <=( a13450a  and  a13447a );
 a13452a <=( a13451a  and  a13444a );
 a13456a <=( (not A167)  and  A168 );
 a13457a <=( (not A170)  and  a13456a );
 a13460a <=( (not A199)  and  A166 );
 a13463a <=( A232  and  (not A200) );
 a13464a <=( a13463a  and  a13460a );
 a13465a <=( a13464a  and  a13457a );
 a13469a <=( A236  and  A234 );
 a13470a <=( (not A233)  and  a13469a );
 a13473a <=( A266  and  (not A265) );
 a13476a <=( A268  and  A267 );
 a13477a <=( a13476a  and  a13473a );
 a13478a <=( a13477a  and  a13470a );
 a13482a <=( (not A167)  and  A168 );
 a13483a <=( (not A170)  and  a13482a );
 a13486a <=( (not A199)  and  A166 );
 a13489a <=( A232  and  (not A200) );
 a13490a <=( a13489a  and  a13486a );
 a13491a <=( a13490a  and  a13483a );
 a13495a <=( A236  and  A234 );
 a13496a <=( (not A233)  and  a13495a );
 a13499a <=( A266  and  (not A265) );
 a13502a <=( A269  and  A267 );
 a13503a <=( a13502a  and  a13499a );
 a13504a <=( a13503a  and  a13496a );
 a13508a <=( (not A167)  and  A168 );
 a13509a <=( (not A170)  and  a13508a );
 a13512a <=( (not A199)  and  A166 );
 a13515a <=( A232  and  (not A200) );
 a13516a <=( a13515a  and  a13512a );
 a13517a <=( a13516a  and  a13509a );
 a13521a <=( A236  and  A234 );
 a13522a <=( (not A233)  and  a13521a );
 a13525a <=( (not A266)  and  A265 );
 a13528a <=( A268  and  A267 );
 a13529a <=( a13528a  and  a13525a );
 a13530a <=( a13529a  and  a13522a );
 a13534a <=( (not A167)  and  A168 );
 a13535a <=( (not A170)  and  a13534a );
 a13538a <=( (not A199)  and  A166 );
 a13541a <=( A232  and  (not A200) );
 a13542a <=( a13541a  and  a13538a );
 a13543a <=( a13542a  and  a13535a );
 a13547a <=( A236  and  A234 );
 a13548a <=( (not A233)  and  a13547a );
 a13551a <=( (not A266)  and  A265 );
 a13554a <=( A269  and  A267 );
 a13555a <=( a13554a  and  a13551a );
 a13556a <=( a13555a  and  a13548a );
 a13560a <=( A167  and  A168 );
 a13561a <=( A169  and  a13560a );
 a13564a <=( (not A201)  and  (not A166) );
 a13567a <=( (not A232)  and  A202 );
 a13568a <=( a13567a  and  a13564a );
 a13569a <=( a13568a  and  a13561a );
 a13573a <=( A235  and  A234 );
 a13574a <=( A233  and  a13573a );
 a13577a <=( (not A299)  and  A298 );
 a13580a <=( A301  and  A300 );
 a13581a <=( a13580a  and  a13577a );
 a13582a <=( a13581a  and  a13574a );
 a13586a <=( A167  and  A168 );
 a13587a <=( A169  and  a13586a );
 a13590a <=( (not A201)  and  (not A166) );
 a13593a <=( (not A232)  and  A202 );
 a13594a <=( a13593a  and  a13590a );
 a13595a <=( a13594a  and  a13587a );
 a13599a <=( A235  and  A234 );
 a13600a <=( A233  and  a13599a );
 a13603a <=( (not A299)  and  A298 );
 a13606a <=( A302  and  A300 );
 a13607a <=( a13606a  and  a13603a );
 a13608a <=( a13607a  and  a13600a );
 a13612a <=( A167  and  A168 );
 a13613a <=( A169  and  a13612a );
 a13616a <=( (not A201)  and  (not A166) );
 a13619a <=( (not A232)  and  A202 );
 a13620a <=( a13619a  and  a13616a );
 a13621a <=( a13620a  and  a13613a );
 a13625a <=( A235  and  A234 );
 a13626a <=( A233  and  a13625a );
 a13629a <=( A299  and  (not A298) );
 a13632a <=( A301  and  A300 );
 a13633a <=( a13632a  and  a13629a );
 a13634a <=( a13633a  and  a13626a );
 a13638a <=( A167  and  A168 );
 a13639a <=( A169  and  a13638a );
 a13642a <=( (not A201)  and  (not A166) );
 a13645a <=( (not A232)  and  A202 );
 a13646a <=( a13645a  and  a13642a );
 a13647a <=( a13646a  and  a13639a );
 a13651a <=( A235  and  A234 );
 a13652a <=( A233  and  a13651a );
 a13655a <=( A299  and  (not A298) );
 a13658a <=( A302  and  A300 );
 a13659a <=( a13658a  and  a13655a );
 a13660a <=( a13659a  and  a13652a );
 a13664a <=( A167  and  A168 );
 a13665a <=( A169  and  a13664a );
 a13668a <=( (not A201)  and  (not A166) );
 a13671a <=( (not A232)  and  A202 );
 a13672a <=( a13671a  and  a13668a );
 a13673a <=( a13672a  and  a13665a );
 a13677a <=( A235  and  A234 );
 a13678a <=( A233  and  a13677a );
 a13681a <=( A266  and  (not A265) );
 a13684a <=( A268  and  A267 );
 a13685a <=( a13684a  and  a13681a );
 a13686a <=( a13685a  and  a13678a );
 a13690a <=( A167  and  A168 );
 a13691a <=( A169  and  a13690a );
 a13694a <=( (not A201)  and  (not A166) );
 a13697a <=( (not A232)  and  A202 );
 a13698a <=( a13697a  and  a13694a );
 a13699a <=( a13698a  and  a13691a );
 a13703a <=( A235  and  A234 );
 a13704a <=( A233  and  a13703a );
 a13707a <=( A266  and  (not A265) );
 a13710a <=( A269  and  A267 );
 a13711a <=( a13710a  and  a13707a );
 a13712a <=( a13711a  and  a13704a );
 a13716a <=( A167  and  A168 );
 a13717a <=( A169  and  a13716a );
 a13720a <=( (not A201)  and  (not A166) );
 a13723a <=( (not A232)  and  A202 );
 a13724a <=( a13723a  and  a13720a );
 a13725a <=( a13724a  and  a13717a );
 a13729a <=( A235  and  A234 );
 a13730a <=( A233  and  a13729a );
 a13733a <=( (not A266)  and  A265 );
 a13736a <=( A268  and  A267 );
 a13737a <=( a13736a  and  a13733a );
 a13738a <=( a13737a  and  a13730a );
 a13742a <=( A167  and  A168 );
 a13743a <=( A169  and  a13742a );
 a13746a <=( (not A201)  and  (not A166) );
 a13749a <=( (not A232)  and  A202 );
 a13750a <=( a13749a  and  a13746a );
 a13751a <=( a13750a  and  a13743a );
 a13755a <=( A235  and  A234 );
 a13756a <=( A233  and  a13755a );
 a13759a <=( (not A266)  and  A265 );
 a13762a <=( A269  and  A267 );
 a13763a <=( a13762a  and  a13759a );
 a13764a <=( a13763a  and  a13756a );
 a13768a <=( A167  and  A168 );
 a13769a <=( A169  and  a13768a );
 a13772a <=( (not A201)  and  (not A166) );
 a13775a <=( (not A232)  and  A202 );
 a13776a <=( a13775a  and  a13772a );
 a13777a <=( a13776a  and  a13769a );
 a13781a <=( A236  and  A234 );
 a13782a <=( A233  and  a13781a );
 a13785a <=( (not A299)  and  A298 );
 a13788a <=( A301  and  A300 );
 a13789a <=( a13788a  and  a13785a );
 a13790a <=( a13789a  and  a13782a );
 a13794a <=( A167  and  A168 );
 a13795a <=( A169  and  a13794a );
 a13798a <=( (not A201)  and  (not A166) );
 a13801a <=( (not A232)  and  A202 );
 a13802a <=( a13801a  and  a13798a );
 a13803a <=( a13802a  and  a13795a );
 a13807a <=( A236  and  A234 );
 a13808a <=( A233  and  a13807a );
 a13811a <=( (not A299)  and  A298 );
 a13814a <=( A302  and  A300 );
 a13815a <=( a13814a  and  a13811a );
 a13816a <=( a13815a  and  a13808a );
 a13820a <=( A167  and  A168 );
 a13821a <=( A169  and  a13820a );
 a13824a <=( (not A201)  and  (not A166) );
 a13827a <=( (not A232)  and  A202 );
 a13828a <=( a13827a  and  a13824a );
 a13829a <=( a13828a  and  a13821a );
 a13833a <=( A236  and  A234 );
 a13834a <=( A233  and  a13833a );
 a13837a <=( A299  and  (not A298) );
 a13840a <=( A301  and  A300 );
 a13841a <=( a13840a  and  a13837a );
 a13842a <=( a13841a  and  a13834a );
 a13846a <=( A167  and  A168 );
 a13847a <=( A169  and  a13846a );
 a13850a <=( (not A201)  and  (not A166) );
 a13853a <=( (not A232)  and  A202 );
 a13854a <=( a13853a  and  a13850a );
 a13855a <=( a13854a  and  a13847a );
 a13859a <=( A236  and  A234 );
 a13860a <=( A233  and  a13859a );
 a13863a <=( A299  and  (not A298) );
 a13866a <=( A302  and  A300 );
 a13867a <=( a13866a  and  a13863a );
 a13868a <=( a13867a  and  a13860a );
 a13872a <=( A167  and  A168 );
 a13873a <=( A169  and  a13872a );
 a13876a <=( (not A201)  and  (not A166) );
 a13879a <=( (not A232)  and  A202 );
 a13880a <=( a13879a  and  a13876a );
 a13881a <=( a13880a  and  a13873a );
 a13885a <=( A236  and  A234 );
 a13886a <=( A233  and  a13885a );
 a13889a <=( A266  and  (not A265) );
 a13892a <=( A268  and  A267 );
 a13893a <=( a13892a  and  a13889a );
 a13894a <=( a13893a  and  a13886a );
 a13898a <=( A167  and  A168 );
 a13899a <=( A169  and  a13898a );
 a13902a <=( (not A201)  and  (not A166) );
 a13905a <=( (not A232)  and  A202 );
 a13906a <=( a13905a  and  a13902a );
 a13907a <=( a13906a  and  a13899a );
 a13911a <=( A236  and  A234 );
 a13912a <=( A233  and  a13911a );
 a13915a <=( A266  and  (not A265) );
 a13918a <=( A269  and  A267 );
 a13919a <=( a13918a  and  a13915a );
 a13920a <=( a13919a  and  a13912a );
 a13924a <=( A167  and  A168 );
 a13925a <=( A169  and  a13924a );
 a13928a <=( (not A201)  and  (not A166) );
 a13931a <=( (not A232)  and  A202 );
 a13932a <=( a13931a  and  a13928a );
 a13933a <=( a13932a  and  a13925a );
 a13937a <=( A236  and  A234 );
 a13938a <=( A233  and  a13937a );
 a13941a <=( (not A266)  and  A265 );
 a13944a <=( A268  and  A267 );
 a13945a <=( a13944a  and  a13941a );
 a13946a <=( a13945a  and  a13938a );
 a13950a <=( A167  and  A168 );
 a13951a <=( A169  and  a13950a );
 a13954a <=( (not A201)  and  (not A166) );
 a13957a <=( (not A232)  and  A202 );
 a13958a <=( a13957a  and  a13954a );
 a13959a <=( a13958a  and  a13951a );
 a13963a <=( A236  and  A234 );
 a13964a <=( A233  and  a13963a );
 a13967a <=( (not A266)  and  A265 );
 a13970a <=( A269  and  A267 );
 a13971a <=( a13970a  and  a13967a );
 a13972a <=( a13971a  and  a13964a );
 a13976a <=( A167  and  A168 );
 a13977a <=( A169  and  a13976a );
 a13980a <=( (not A201)  and  (not A166) );
 a13983a <=( A232  and  A202 );
 a13984a <=( a13983a  and  a13980a );
 a13985a <=( a13984a  and  a13977a );
 a13989a <=( A235  and  A234 );
 a13990a <=( (not A233)  and  a13989a );
 a13993a <=( (not A299)  and  A298 );
 a13996a <=( A301  and  A300 );
 a13997a <=( a13996a  and  a13993a );
 a13998a <=( a13997a  and  a13990a );
 a14002a <=( A167  and  A168 );
 a14003a <=( A169  and  a14002a );
 a14006a <=( (not A201)  and  (not A166) );
 a14009a <=( A232  and  A202 );
 a14010a <=( a14009a  and  a14006a );
 a14011a <=( a14010a  and  a14003a );
 a14015a <=( A235  and  A234 );
 a14016a <=( (not A233)  and  a14015a );
 a14019a <=( (not A299)  and  A298 );
 a14022a <=( A302  and  A300 );
 a14023a <=( a14022a  and  a14019a );
 a14024a <=( a14023a  and  a14016a );
 a14028a <=( A167  and  A168 );
 a14029a <=( A169  and  a14028a );
 a14032a <=( (not A201)  and  (not A166) );
 a14035a <=( A232  and  A202 );
 a14036a <=( a14035a  and  a14032a );
 a14037a <=( a14036a  and  a14029a );
 a14041a <=( A235  and  A234 );
 a14042a <=( (not A233)  and  a14041a );
 a14045a <=( A299  and  (not A298) );
 a14048a <=( A301  and  A300 );
 a14049a <=( a14048a  and  a14045a );
 a14050a <=( a14049a  and  a14042a );
 a14054a <=( A167  and  A168 );
 a14055a <=( A169  and  a14054a );
 a14058a <=( (not A201)  and  (not A166) );
 a14061a <=( A232  and  A202 );
 a14062a <=( a14061a  and  a14058a );
 a14063a <=( a14062a  and  a14055a );
 a14067a <=( A235  and  A234 );
 a14068a <=( (not A233)  and  a14067a );
 a14071a <=( A299  and  (not A298) );
 a14074a <=( A302  and  A300 );
 a14075a <=( a14074a  and  a14071a );
 a14076a <=( a14075a  and  a14068a );
 a14080a <=( A167  and  A168 );
 a14081a <=( A169  and  a14080a );
 a14084a <=( (not A201)  and  (not A166) );
 a14087a <=( A232  and  A202 );
 a14088a <=( a14087a  and  a14084a );
 a14089a <=( a14088a  and  a14081a );
 a14093a <=( A235  and  A234 );
 a14094a <=( (not A233)  and  a14093a );
 a14097a <=( A266  and  (not A265) );
 a14100a <=( A268  and  A267 );
 a14101a <=( a14100a  and  a14097a );
 a14102a <=( a14101a  and  a14094a );
 a14106a <=( A167  and  A168 );
 a14107a <=( A169  and  a14106a );
 a14110a <=( (not A201)  and  (not A166) );
 a14113a <=( A232  and  A202 );
 a14114a <=( a14113a  and  a14110a );
 a14115a <=( a14114a  and  a14107a );
 a14119a <=( A235  and  A234 );
 a14120a <=( (not A233)  and  a14119a );
 a14123a <=( A266  and  (not A265) );
 a14126a <=( A269  and  A267 );
 a14127a <=( a14126a  and  a14123a );
 a14128a <=( a14127a  and  a14120a );
 a14132a <=( A167  and  A168 );
 a14133a <=( A169  and  a14132a );
 a14136a <=( (not A201)  and  (not A166) );
 a14139a <=( A232  and  A202 );
 a14140a <=( a14139a  and  a14136a );
 a14141a <=( a14140a  and  a14133a );
 a14145a <=( A235  and  A234 );
 a14146a <=( (not A233)  and  a14145a );
 a14149a <=( (not A266)  and  A265 );
 a14152a <=( A268  and  A267 );
 a14153a <=( a14152a  and  a14149a );
 a14154a <=( a14153a  and  a14146a );
 a14158a <=( A167  and  A168 );
 a14159a <=( A169  and  a14158a );
 a14162a <=( (not A201)  and  (not A166) );
 a14165a <=( A232  and  A202 );
 a14166a <=( a14165a  and  a14162a );
 a14167a <=( a14166a  and  a14159a );
 a14171a <=( A235  and  A234 );
 a14172a <=( (not A233)  and  a14171a );
 a14175a <=( (not A266)  and  A265 );
 a14178a <=( A269  and  A267 );
 a14179a <=( a14178a  and  a14175a );
 a14180a <=( a14179a  and  a14172a );
 a14184a <=( A167  and  A168 );
 a14185a <=( A169  and  a14184a );
 a14188a <=( (not A201)  and  (not A166) );
 a14191a <=( A232  and  A202 );
 a14192a <=( a14191a  and  a14188a );
 a14193a <=( a14192a  and  a14185a );
 a14197a <=( A236  and  A234 );
 a14198a <=( (not A233)  and  a14197a );
 a14201a <=( (not A299)  and  A298 );
 a14204a <=( A301  and  A300 );
 a14205a <=( a14204a  and  a14201a );
 a14206a <=( a14205a  and  a14198a );
 a14210a <=( A167  and  A168 );
 a14211a <=( A169  and  a14210a );
 a14214a <=( (not A201)  and  (not A166) );
 a14217a <=( A232  and  A202 );
 a14218a <=( a14217a  and  a14214a );
 a14219a <=( a14218a  and  a14211a );
 a14223a <=( A236  and  A234 );
 a14224a <=( (not A233)  and  a14223a );
 a14227a <=( (not A299)  and  A298 );
 a14230a <=( A302  and  A300 );
 a14231a <=( a14230a  and  a14227a );
 a14232a <=( a14231a  and  a14224a );
 a14236a <=( A167  and  A168 );
 a14237a <=( A169  and  a14236a );
 a14240a <=( (not A201)  and  (not A166) );
 a14243a <=( A232  and  A202 );
 a14244a <=( a14243a  and  a14240a );
 a14245a <=( a14244a  and  a14237a );
 a14249a <=( A236  and  A234 );
 a14250a <=( (not A233)  and  a14249a );
 a14253a <=( A299  and  (not A298) );
 a14256a <=( A301  and  A300 );
 a14257a <=( a14256a  and  a14253a );
 a14258a <=( a14257a  and  a14250a );
 a14262a <=( A167  and  A168 );
 a14263a <=( A169  and  a14262a );
 a14266a <=( (not A201)  and  (not A166) );
 a14269a <=( A232  and  A202 );
 a14270a <=( a14269a  and  a14266a );
 a14271a <=( a14270a  and  a14263a );
 a14275a <=( A236  and  A234 );
 a14276a <=( (not A233)  and  a14275a );
 a14279a <=( A299  and  (not A298) );
 a14282a <=( A302  and  A300 );
 a14283a <=( a14282a  and  a14279a );
 a14284a <=( a14283a  and  a14276a );
 a14288a <=( A167  and  A168 );
 a14289a <=( A169  and  a14288a );
 a14292a <=( (not A201)  and  (not A166) );
 a14295a <=( A232  and  A202 );
 a14296a <=( a14295a  and  a14292a );
 a14297a <=( a14296a  and  a14289a );
 a14301a <=( A236  and  A234 );
 a14302a <=( (not A233)  and  a14301a );
 a14305a <=( A266  and  (not A265) );
 a14308a <=( A268  and  A267 );
 a14309a <=( a14308a  and  a14305a );
 a14310a <=( a14309a  and  a14302a );
 a14314a <=( A167  and  A168 );
 a14315a <=( A169  and  a14314a );
 a14318a <=( (not A201)  and  (not A166) );
 a14321a <=( A232  and  A202 );
 a14322a <=( a14321a  and  a14318a );
 a14323a <=( a14322a  and  a14315a );
 a14327a <=( A236  and  A234 );
 a14328a <=( (not A233)  and  a14327a );
 a14331a <=( A266  and  (not A265) );
 a14334a <=( A269  and  A267 );
 a14335a <=( a14334a  and  a14331a );
 a14336a <=( a14335a  and  a14328a );
 a14340a <=( A167  and  A168 );
 a14341a <=( A169  and  a14340a );
 a14344a <=( (not A201)  and  (not A166) );
 a14347a <=( A232  and  A202 );
 a14348a <=( a14347a  and  a14344a );
 a14349a <=( a14348a  and  a14341a );
 a14353a <=( A236  and  A234 );
 a14354a <=( (not A233)  and  a14353a );
 a14357a <=( (not A266)  and  A265 );
 a14360a <=( A268  and  A267 );
 a14361a <=( a14360a  and  a14357a );
 a14362a <=( a14361a  and  a14354a );
 a14366a <=( A167  and  A168 );
 a14367a <=( A169  and  a14366a );
 a14370a <=( (not A201)  and  (not A166) );
 a14373a <=( A232  and  A202 );
 a14374a <=( a14373a  and  a14370a );
 a14375a <=( a14374a  and  a14367a );
 a14379a <=( A236  and  A234 );
 a14380a <=( (not A233)  and  a14379a );
 a14383a <=( (not A266)  and  A265 );
 a14386a <=( A269  and  A267 );
 a14387a <=( a14386a  and  a14383a );
 a14388a <=( a14387a  and  a14380a );
 a14392a <=( A167  and  A168 );
 a14393a <=( A169  and  a14392a );
 a14396a <=( (not A201)  and  (not A166) );
 a14399a <=( (not A232)  and  A203 );
 a14400a <=( a14399a  and  a14396a );
 a14401a <=( a14400a  and  a14393a );
 a14405a <=( A235  and  A234 );
 a14406a <=( A233  and  a14405a );
 a14409a <=( (not A299)  and  A298 );
 a14412a <=( A301  and  A300 );
 a14413a <=( a14412a  and  a14409a );
 a14414a <=( a14413a  and  a14406a );
 a14418a <=( A167  and  A168 );
 a14419a <=( A169  and  a14418a );
 a14422a <=( (not A201)  and  (not A166) );
 a14425a <=( (not A232)  and  A203 );
 a14426a <=( a14425a  and  a14422a );
 a14427a <=( a14426a  and  a14419a );
 a14431a <=( A235  and  A234 );
 a14432a <=( A233  and  a14431a );
 a14435a <=( (not A299)  and  A298 );
 a14438a <=( A302  and  A300 );
 a14439a <=( a14438a  and  a14435a );
 a14440a <=( a14439a  and  a14432a );
 a14444a <=( A167  and  A168 );
 a14445a <=( A169  and  a14444a );
 a14448a <=( (not A201)  and  (not A166) );
 a14451a <=( (not A232)  and  A203 );
 a14452a <=( a14451a  and  a14448a );
 a14453a <=( a14452a  and  a14445a );
 a14457a <=( A235  and  A234 );
 a14458a <=( A233  and  a14457a );
 a14461a <=( A299  and  (not A298) );
 a14464a <=( A301  and  A300 );
 a14465a <=( a14464a  and  a14461a );
 a14466a <=( a14465a  and  a14458a );
 a14470a <=( A167  and  A168 );
 a14471a <=( A169  and  a14470a );
 a14474a <=( (not A201)  and  (not A166) );
 a14477a <=( (not A232)  and  A203 );
 a14478a <=( a14477a  and  a14474a );
 a14479a <=( a14478a  and  a14471a );
 a14483a <=( A235  and  A234 );
 a14484a <=( A233  and  a14483a );
 a14487a <=( A299  and  (not A298) );
 a14490a <=( A302  and  A300 );
 a14491a <=( a14490a  and  a14487a );
 a14492a <=( a14491a  and  a14484a );
 a14496a <=( A167  and  A168 );
 a14497a <=( A169  and  a14496a );
 a14500a <=( (not A201)  and  (not A166) );
 a14503a <=( (not A232)  and  A203 );
 a14504a <=( a14503a  and  a14500a );
 a14505a <=( a14504a  and  a14497a );
 a14509a <=( A235  and  A234 );
 a14510a <=( A233  and  a14509a );
 a14513a <=( A266  and  (not A265) );
 a14516a <=( A268  and  A267 );
 a14517a <=( a14516a  and  a14513a );
 a14518a <=( a14517a  and  a14510a );
 a14522a <=( A167  and  A168 );
 a14523a <=( A169  and  a14522a );
 a14526a <=( (not A201)  and  (not A166) );
 a14529a <=( (not A232)  and  A203 );
 a14530a <=( a14529a  and  a14526a );
 a14531a <=( a14530a  and  a14523a );
 a14535a <=( A235  and  A234 );
 a14536a <=( A233  and  a14535a );
 a14539a <=( A266  and  (not A265) );
 a14542a <=( A269  and  A267 );
 a14543a <=( a14542a  and  a14539a );
 a14544a <=( a14543a  and  a14536a );
 a14548a <=( A167  and  A168 );
 a14549a <=( A169  and  a14548a );
 a14552a <=( (not A201)  and  (not A166) );
 a14555a <=( (not A232)  and  A203 );
 a14556a <=( a14555a  and  a14552a );
 a14557a <=( a14556a  and  a14549a );
 a14561a <=( A235  and  A234 );
 a14562a <=( A233  and  a14561a );
 a14565a <=( (not A266)  and  A265 );
 a14568a <=( A268  and  A267 );
 a14569a <=( a14568a  and  a14565a );
 a14570a <=( a14569a  and  a14562a );
 a14574a <=( A167  and  A168 );
 a14575a <=( A169  and  a14574a );
 a14578a <=( (not A201)  and  (not A166) );
 a14581a <=( (not A232)  and  A203 );
 a14582a <=( a14581a  and  a14578a );
 a14583a <=( a14582a  and  a14575a );
 a14587a <=( A235  and  A234 );
 a14588a <=( A233  and  a14587a );
 a14591a <=( (not A266)  and  A265 );
 a14594a <=( A269  and  A267 );
 a14595a <=( a14594a  and  a14591a );
 a14596a <=( a14595a  and  a14588a );
 a14600a <=( A167  and  A168 );
 a14601a <=( A169  and  a14600a );
 a14604a <=( (not A201)  and  (not A166) );
 a14607a <=( (not A232)  and  A203 );
 a14608a <=( a14607a  and  a14604a );
 a14609a <=( a14608a  and  a14601a );
 a14613a <=( A236  and  A234 );
 a14614a <=( A233  and  a14613a );
 a14617a <=( (not A299)  and  A298 );
 a14620a <=( A301  and  A300 );
 a14621a <=( a14620a  and  a14617a );
 a14622a <=( a14621a  and  a14614a );
 a14626a <=( A167  and  A168 );
 a14627a <=( A169  and  a14626a );
 a14630a <=( (not A201)  and  (not A166) );
 a14633a <=( (not A232)  and  A203 );
 a14634a <=( a14633a  and  a14630a );
 a14635a <=( a14634a  and  a14627a );
 a14639a <=( A236  and  A234 );
 a14640a <=( A233  and  a14639a );
 a14643a <=( (not A299)  and  A298 );
 a14646a <=( A302  and  A300 );
 a14647a <=( a14646a  and  a14643a );
 a14648a <=( a14647a  and  a14640a );
 a14652a <=( A167  and  A168 );
 a14653a <=( A169  and  a14652a );
 a14656a <=( (not A201)  and  (not A166) );
 a14659a <=( (not A232)  and  A203 );
 a14660a <=( a14659a  and  a14656a );
 a14661a <=( a14660a  and  a14653a );
 a14665a <=( A236  and  A234 );
 a14666a <=( A233  and  a14665a );
 a14669a <=( A299  and  (not A298) );
 a14672a <=( A301  and  A300 );
 a14673a <=( a14672a  and  a14669a );
 a14674a <=( a14673a  and  a14666a );
 a14678a <=( A167  and  A168 );
 a14679a <=( A169  and  a14678a );
 a14682a <=( (not A201)  and  (not A166) );
 a14685a <=( (not A232)  and  A203 );
 a14686a <=( a14685a  and  a14682a );
 a14687a <=( a14686a  and  a14679a );
 a14691a <=( A236  and  A234 );
 a14692a <=( A233  and  a14691a );
 a14695a <=( A299  and  (not A298) );
 a14698a <=( A302  and  A300 );
 a14699a <=( a14698a  and  a14695a );
 a14700a <=( a14699a  and  a14692a );
 a14704a <=( A167  and  A168 );
 a14705a <=( A169  and  a14704a );
 a14708a <=( (not A201)  and  (not A166) );
 a14711a <=( (not A232)  and  A203 );
 a14712a <=( a14711a  and  a14708a );
 a14713a <=( a14712a  and  a14705a );
 a14717a <=( A236  and  A234 );
 a14718a <=( A233  and  a14717a );
 a14721a <=( A266  and  (not A265) );
 a14724a <=( A268  and  A267 );
 a14725a <=( a14724a  and  a14721a );
 a14726a <=( a14725a  and  a14718a );
 a14730a <=( A167  and  A168 );
 a14731a <=( A169  and  a14730a );
 a14734a <=( (not A201)  and  (not A166) );
 a14737a <=( (not A232)  and  A203 );
 a14738a <=( a14737a  and  a14734a );
 a14739a <=( a14738a  and  a14731a );
 a14743a <=( A236  and  A234 );
 a14744a <=( A233  and  a14743a );
 a14747a <=( A266  and  (not A265) );
 a14750a <=( A269  and  A267 );
 a14751a <=( a14750a  and  a14747a );
 a14752a <=( a14751a  and  a14744a );
 a14756a <=( A167  and  A168 );
 a14757a <=( A169  and  a14756a );
 a14760a <=( (not A201)  and  (not A166) );
 a14763a <=( (not A232)  and  A203 );
 a14764a <=( a14763a  and  a14760a );
 a14765a <=( a14764a  and  a14757a );
 a14769a <=( A236  and  A234 );
 a14770a <=( A233  and  a14769a );
 a14773a <=( (not A266)  and  A265 );
 a14776a <=( A268  and  A267 );
 a14777a <=( a14776a  and  a14773a );
 a14778a <=( a14777a  and  a14770a );
 a14782a <=( A167  and  A168 );
 a14783a <=( A169  and  a14782a );
 a14786a <=( (not A201)  and  (not A166) );
 a14789a <=( (not A232)  and  A203 );
 a14790a <=( a14789a  and  a14786a );
 a14791a <=( a14790a  and  a14783a );
 a14795a <=( A236  and  A234 );
 a14796a <=( A233  and  a14795a );
 a14799a <=( (not A266)  and  A265 );
 a14802a <=( A269  and  A267 );
 a14803a <=( a14802a  and  a14799a );
 a14804a <=( a14803a  and  a14796a );
 a14808a <=( A167  and  A168 );
 a14809a <=( A169  and  a14808a );
 a14812a <=( (not A201)  and  (not A166) );
 a14815a <=( A232  and  A203 );
 a14816a <=( a14815a  and  a14812a );
 a14817a <=( a14816a  and  a14809a );
 a14821a <=( A235  and  A234 );
 a14822a <=( (not A233)  and  a14821a );
 a14825a <=( (not A299)  and  A298 );
 a14828a <=( A301  and  A300 );
 a14829a <=( a14828a  and  a14825a );
 a14830a <=( a14829a  and  a14822a );
 a14834a <=( A167  and  A168 );
 a14835a <=( A169  and  a14834a );
 a14838a <=( (not A201)  and  (not A166) );
 a14841a <=( A232  and  A203 );
 a14842a <=( a14841a  and  a14838a );
 a14843a <=( a14842a  and  a14835a );
 a14847a <=( A235  and  A234 );
 a14848a <=( (not A233)  and  a14847a );
 a14851a <=( (not A299)  and  A298 );
 a14854a <=( A302  and  A300 );
 a14855a <=( a14854a  and  a14851a );
 a14856a <=( a14855a  and  a14848a );
 a14860a <=( A167  and  A168 );
 a14861a <=( A169  and  a14860a );
 a14864a <=( (not A201)  and  (not A166) );
 a14867a <=( A232  and  A203 );
 a14868a <=( a14867a  and  a14864a );
 a14869a <=( a14868a  and  a14861a );
 a14873a <=( A235  and  A234 );
 a14874a <=( (not A233)  and  a14873a );
 a14877a <=( A299  and  (not A298) );
 a14880a <=( A301  and  A300 );
 a14881a <=( a14880a  and  a14877a );
 a14882a <=( a14881a  and  a14874a );
 a14886a <=( A167  and  A168 );
 a14887a <=( A169  and  a14886a );
 a14890a <=( (not A201)  and  (not A166) );
 a14893a <=( A232  and  A203 );
 a14894a <=( a14893a  and  a14890a );
 a14895a <=( a14894a  and  a14887a );
 a14899a <=( A235  and  A234 );
 a14900a <=( (not A233)  and  a14899a );
 a14903a <=( A299  and  (not A298) );
 a14906a <=( A302  and  A300 );
 a14907a <=( a14906a  and  a14903a );
 a14908a <=( a14907a  and  a14900a );
 a14912a <=( A167  and  A168 );
 a14913a <=( A169  and  a14912a );
 a14916a <=( (not A201)  and  (not A166) );
 a14919a <=( A232  and  A203 );
 a14920a <=( a14919a  and  a14916a );
 a14921a <=( a14920a  and  a14913a );
 a14925a <=( A235  and  A234 );
 a14926a <=( (not A233)  and  a14925a );
 a14929a <=( A266  and  (not A265) );
 a14932a <=( A268  and  A267 );
 a14933a <=( a14932a  and  a14929a );
 a14934a <=( a14933a  and  a14926a );
 a14938a <=( A167  and  A168 );
 a14939a <=( A169  and  a14938a );
 a14942a <=( (not A201)  and  (not A166) );
 a14945a <=( A232  and  A203 );
 a14946a <=( a14945a  and  a14942a );
 a14947a <=( a14946a  and  a14939a );
 a14951a <=( A235  and  A234 );
 a14952a <=( (not A233)  and  a14951a );
 a14955a <=( A266  and  (not A265) );
 a14958a <=( A269  and  A267 );
 a14959a <=( a14958a  and  a14955a );
 a14960a <=( a14959a  and  a14952a );
 a14964a <=( A167  and  A168 );
 a14965a <=( A169  and  a14964a );
 a14968a <=( (not A201)  and  (not A166) );
 a14971a <=( A232  and  A203 );
 a14972a <=( a14971a  and  a14968a );
 a14973a <=( a14972a  and  a14965a );
 a14977a <=( A235  and  A234 );
 a14978a <=( (not A233)  and  a14977a );
 a14981a <=( (not A266)  and  A265 );
 a14984a <=( A268  and  A267 );
 a14985a <=( a14984a  and  a14981a );
 a14986a <=( a14985a  and  a14978a );
 a14990a <=( A167  and  A168 );
 a14991a <=( A169  and  a14990a );
 a14994a <=( (not A201)  and  (not A166) );
 a14997a <=( A232  and  A203 );
 a14998a <=( a14997a  and  a14994a );
 a14999a <=( a14998a  and  a14991a );
 a15003a <=( A235  and  A234 );
 a15004a <=( (not A233)  and  a15003a );
 a15007a <=( (not A266)  and  A265 );
 a15010a <=( A269  and  A267 );
 a15011a <=( a15010a  and  a15007a );
 a15012a <=( a15011a  and  a15004a );
 a15016a <=( A167  and  A168 );
 a15017a <=( A169  and  a15016a );
 a15020a <=( (not A201)  and  (not A166) );
 a15023a <=( A232  and  A203 );
 a15024a <=( a15023a  and  a15020a );
 a15025a <=( a15024a  and  a15017a );
 a15029a <=( A236  and  A234 );
 a15030a <=( (not A233)  and  a15029a );
 a15033a <=( (not A299)  and  A298 );
 a15036a <=( A301  and  A300 );
 a15037a <=( a15036a  and  a15033a );
 a15038a <=( a15037a  and  a15030a );
 a15042a <=( A167  and  A168 );
 a15043a <=( A169  and  a15042a );
 a15046a <=( (not A201)  and  (not A166) );
 a15049a <=( A232  and  A203 );
 a15050a <=( a15049a  and  a15046a );
 a15051a <=( a15050a  and  a15043a );
 a15055a <=( A236  and  A234 );
 a15056a <=( (not A233)  and  a15055a );
 a15059a <=( (not A299)  and  A298 );
 a15062a <=( A302  and  A300 );
 a15063a <=( a15062a  and  a15059a );
 a15064a <=( a15063a  and  a15056a );
 a15068a <=( A167  and  A168 );
 a15069a <=( A169  and  a15068a );
 a15072a <=( (not A201)  and  (not A166) );
 a15075a <=( A232  and  A203 );
 a15076a <=( a15075a  and  a15072a );
 a15077a <=( a15076a  and  a15069a );
 a15081a <=( A236  and  A234 );
 a15082a <=( (not A233)  and  a15081a );
 a15085a <=( A299  and  (not A298) );
 a15088a <=( A301  and  A300 );
 a15089a <=( a15088a  and  a15085a );
 a15090a <=( a15089a  and  a15082a );
 a15094a <=( A167  and  A168 );
 a15095a <=( A169  and  a15094a );
 a15098a <=( (not A201)  and  (not A166) );
 a15101a <=( A232  and  A203 );
 a15102a <=( a15101a  and  a15098a );
 a15103a <=( a15102a  and  a15095a );
 a15107a <=( A236  and  A234 );
 a15108a <=( (not A233)  and  a15107a );
 a15111a <=( A299  and  (not A298) );
 a15114a <=( A302  and  A300 );
 a15115a <=( a15114a  and  a15111a );
 a15116a <=( a15115a  and  a15108a );
 a15120a <=( A167  and  A168 );
 a15121a <=( A169  and  a15120a );
 a15124a <=( (not A201)  and  (not A166) );
 a15127a <=( A232  and  A203 );
 a15128a <=( a15127a  and  a15124a );
 a15129a <=( a15128a  and  a15121a );
 a15133a <=( A236  and  A234 );
 a15134a <=( (not A233)  and  a15133a );
 a15137a <=( A266  and  (not A265) );
 a15140a <=( A268  and  A267 );
 a15141a <=( a15140a  and  a15137a );
 a15142a <=( a15141a  and  a15134a );
 a15146a <=( A167  and  A168 );
 a15147a <=( A169  and  a15146a );
 a15150a <=( (not A201)  and  (not A166) );
 a15153a <=( A232  and  A203 );
 a15154a <=( a15153a  and  a15150a );
 a15155a <=( a15154a  and  a15147a );
 a15159a <=( A236  and  A234 );
 a15160a <=( (not A233)  and  a15159a );
 a15163a <=( A266  and  (not A265) );
 a15166a <=( A269  and  A267 );
 a15167a <=( a15166a  and  a15163a );
 a15168a <=( a15167a  and  a15160a );
 a15172a <=( A167  and  A168 );
 a15173a <=( A169  and  a15172a );
 a15176a <=( (not A201)  and  (not A166) );
 a15179a <=( A232  and  A203 );
 a15180a <=( a15179a  and  a15176a );
 a15181a <=( a15180a  and  a15173a );
 a15185a <=( A236  and  A234 );
 a15186a <=( (not A233)  and  a15185a );
 a15189a <=( (not A266)  and  A265 );
 a15192a <=( A268  and  A267 );
 a15193a <=( a15192a  and  a15189a );
 a15194a <=( a15193a  and  a15186a );
 a15198a <=( A167  and  A168 );
 a15199a <=( A169  and  a15198a );
 a15202a <=( (not A201)  and  (not A166) );
 a15205a <=( A232  and  A203 );
 a15206a <=( a15205a  and  a15202a );
 a15207a <=( a15206a  and  a15199a );
 a15211a <=( A236  and  A234 );
 a15212a <=( (not A233)  and  a15211a );
 a15215a <=( (not A266)  and  A265 );
 a15218a <=( A269  and  A267 );
 a15219a <=( a15218a  and  a15215a );
 a15220a <=( a15219a  and  a15212a );
 a15224a <=( A167  and  A168 );
 a15225a <=( A169  and  a15224a );
 a15228a <=( A199  and  (not A166) );
 a15231a <=( (not A232)  and  A200 );
 a15232a <=( a15231a  and  a15228a );
 a15233a <=( a15232a  and  a15225a );
 a15237a <=( A235  and  A234 );
 a15238a <=( A233  and  a15237a );
 a15241a <=( (not A299)  and  A298 );
 a15244a <=( A301  and  A300 );
 a15245a <=( a15244a  and  a15241a );
 a15246a <=( a15245a  and  a15238a );
 a15250a <=( A167  and  A168 );
 a15251a <=( A169  and  a15250a );
 a15254a <=( A199  and  (not A166) );
 a15257a <=( (not A232)  and  A200 );
 a15258a <=( a15257a  and  a15254a );
 a15259a <=( a15258a  and  a15251a );
 a15263a <=( A235  and  A234 );
 a15264a <=( A233  and  a15263a );
 a15267a <=( (not A299)  and  A298 );
 a15270a <=( A302  and  A300 );
 a15271a <=( a15270a  and  a15267a );
 a15272a <=( a15271a  and  a15264a );
 a15276a <=( A167  and  A168 );
 a15277a <=( A169  and  a15276a );
 a15280a <=( A199  and  (not A166) );
 a15283a <=( (not A232)  and  A200 );
 a15284a <=( a15283a  and  a15280a );
 a15285a <=( a15284a  and  a15277a );
 a15289a <=( A235  and  A234 );
 a15290a <=( A233  and  a15289a );
 a15293a <=( A299  and  (not A298) );
 a15296a <=( A301  and  A300 );
 a15297a <=( a15296a  and  a15293a );
 a15298a <=( a15297a  and  a15290a );
 a15302a <=( A167  and  A168 );
 a15303a <=( A169  and  a15302a );
 a15306a <=( A199  and  (not A166) );
 a15309a <=( (not A232)  and  A200 );
 a15310a <=( a15309a  and  a15306a );
 a15311a <=( a15310a  and  a15303a );
 a15315a <=( A235  and  A234 );
 a15316a <=( A233  and  a15315a );
 a15319a <=( A299  and  (not A298) );
 a15322a <=( A302  and  A300 );
 a15323a <=( a15322a  and  a15319a );
 a15324a <=( a15323a  and  a15316a );
 a15328a <=( A167  and  A168 );
 a15329a <=( A169  and  a15328a );
 a15332a <=( A199  and  (not A166) );
 a15335a <=( (not A232)  and  A200 );
 a15336a <=( a15335a  and  a15332a );
 a15337a <=( a15336a  and  a15329a );
 a15341a <=( A235  and  A234 );
 a15342a <=( A233  and  a15341a );
 a15345a <=( A266  and  (not A265) );
 a15348a <=( A268  and  A267 );
 a15349a <=( a15348a  and  a15345a );
 a15350a <=( a15349a  and  a15342a );
 a15354a <=( A167  and  A168 );
 a15355a <=( A169  and  a15354a );
 a15358a <=( A199  and  (not A166) );
 a15361a <=( (not A232)  and  A200 );
 a15362a <=( a15361a  and  a15358a );
 a15363a <=( a15362a  and  a15355a );
 a15367a <=( A235  and  A234 );
 a15368a <=( A233  and  a15367a );
 a15371a <=( A266  and  (not A265) );
 a15374a <=( A269  and  A267 );
 a15375a <=( a15374a  and  a15371a );
 a15376a <=( a15375a  and  a15368a );
 a15380a <=( A167  and  A168 );
 a15381a <=( A169  and  a15380a );
 a15384a <=( A199  and  (not A166) );
 a15387a <=( (not A232)  and  A200 );
 a15388a <=( a15387a  and  a15384a );
 a15389a <=( a15388a  and  a15381a );
 a15393a <=( A235  and  A234 );
 a15394a <=( A233  and  a15393a );
 a15397a <=( (not A266)  and  A265 );
 a15400a <=( A268  and  A267 );
 a15401a <=( a15400a  and  a15397a );
 a15402a <=( a15401a  and  a15394a );
 a15406a <=( A167  and  A168 );
 a15407a <=( A169  and  a15406a );
 a15410a <=( A199  and  (not A166) );
 a15413a <=( (not A232)  and  A200 );
 a15414a <=( a15413a  and  a15410a );
 a15415a <=( a15414a  and  a15407a );
 a15419a <=( A235  and  A234 );
 a15420a <=( A233  and  a15419a );
 a15423a <=( (not A266)  and  A265 );
 a15426a <=( A269  and  A267 );
 a15427a <=( a15426a  and  a15423a );
 a15428a <=( a15427a  and  a15420a );
 a15432a <=( A167  and  A168 );
 a15433a <=( A169  and  a15432a );
 a15436a <=( A199  and  (not A166) );
 a15439a <=( (not A232)  and  A200 );
 a15440a <=( a15439a  and  a15436a );
 a15441a <=( a15440a  and  a15433a );
 a15445a <=( A236  and  A234 );
 a15446a <=( A233  and  a15445a );
 a15449a <=( (not A299)  and  A298 );
 a15452a <=( A301  and  A300 );
 a15453a <=( a15452a  and  a15449a );
 a15454a <=( a15453a  and  a15446a );
 a15458a <=( A167  and  A168 );
 a15459a <=( A169  and  a15458a );
 a15462a <=( A199  and  (not A166) );
 a15465a <=( (not A232)  and  A200 );
 a15466a <=( a15465a  and  a15462a );
 a15467a <=( a15466a  and  a15459a );
 a15471a <=( A236  and  A234 );
 a15472a <=( A233  and  a15471a );
 a15475a <=( (not A299)  and  A298 );
 a15478a <=( A302  and  A300 );
 a15479a <=( a15478a  and  a15475a );
 a15480a <=( a15479a  and  a15472a );
 a15484a <=( A167  and  A168 );
 a15485a <=( A169  and  a15484a );
 a15488a <=( A199  and  (not A166) );
 a15491a <=( (not A232)  and  A200 );
 a15492a <=( a15491a  and  a15488a );
 a15493a <=( a15492a  and  a15485a );
 a15497a <=( A236  and  A234 );
 a15498a <=( A233  and  a15497a );
 a15501a <=( A299  and  (not A298) );
 a15504a <=( A301  and  A300 );
 a15505a <=( a15504a  and  a15501a );
 a15506a <=( a15505a  and  a15498a );
 a15510a <=( A167  and  A168 );
 a15511a <=( A169  and  a15510a );
 a15514a <=( A199  and  (not A166) );
 a15517a <=( (not A232)  and  A200 );
 a15518a <=( a15517a  and  a15514a );
 a15519a <=( a15518a  and  a15511a );
 a15523a <=( A236  and  A234 );
 a15524a <=( A233  and  a15523a );
 a15527a <=( A299  and  (not A298) );
 a15530a <=( A302  and  A300 );
 a15531a <=( a15530a  and  a15527a );
 a15532a <=( a15531a  and  a15524a );
 a15536a <=( A167  and  A168 );
 a15537a <=( A169  and  a15536a );
 a15540a <=( A199  and  (not A166) );
 a15543a <=( (not A232)  and  A200 );
 a15544a <=( a15543a  and  a15540a );
 a15545a <=( a15544a  and  a15537a );
 a15549a <=( A236  and  A234 );
 a15550a <=( A233  and  a15549a );
 a15553a <=( A266  and  (not A265) );
 a15556a <=( A268  and  A267 );
 a15557a <=( a15556a  and  a15553a );
 a15558a <=( a15557a  and  a15550a );
 a15562a <=( A167  and  A168 );
 a15563a <=( A169  and  a15562a );
 a15566a <=( A199  and  (not A166) );
 a15569a <=( (not A232)  and  A200 );
 a15570a <=( a15569a  and  a15566a );
 a15571a <=( a15570a  and  a15563a );
 a15575a <=( A236  and  A234 );
 a15576a <=( A233  and  a15575a );
 a15579a <=( A266  and  (not A265) );
 a15582a <=( A269  and  A267 );
 a15583a <=( a15582a  and  a15579a );
 a15584a <=( a15583a  and  a15576a );
 a15588a <=( A167  and  A168 );
 a15589a <=( A169  and  a15588a );
 a15592a <=( A199  and  (not A166) );
 a15595a <=( (not A232)  and  A200 );
 a15596a <=( a15595a  and  a15592a );
 a15597a <=( a15596a  and  a15589a );
 a15601a <=( A236  and  A234 );
 a15602a <=( A233  and  a15601a );
 a15605a <=( (not A266)  and  A265 );
 a15608a <=( A268  and  A267 );
 a15609a <=( a15608a  and  a15605a );
 a15610a <=( a15609a  and  a15602a );
 a15614a <=( A167  and  A168 );
 a15615a <=( A169  and  a15614a );
 a15618a <=( A199  and  (not A166) );
 a15621a <=( (not A232)  and  A200 );
 a15622a <=( a15621a  and  a15618a );
 a15623a <=( a15622a  and  a15615a );
 a15627a <=( A236  and  A234 );
 a15628a <=( A233  and  a15627a );
 a15631a <=( (not A266)  and  A265 );
 a15634a <=( A269  and  A267 );
 a15635a <=( a15634a  and  a15631a );
 a15636a <=( a15635a  and  a15628a );
 a15640a <=( A167  and  A168 );
 a15641a <=( A169  and  a15640a );
 a15644a <=( A199  and  (not A166) );
 a15647a <=( A232  and  A200 );
 a15648a <=( a15647a  and  a15644a );
 a15649a <=( a15648a  and  a15641a );
 a15653a <=( A235  and  A234 );
 a15654a <=( (not A233)  and  a15653a );
 a15657a <=( (not A299)  and  A298 );
 a15660a <=( A301  and  A300 );
 a15661a <=( a15660a  and  a15657a );
 a15662a <=( a15661a  and  a15654a );
 a15666a <=( A167  and  A168 );
 a15667a <=( A169  and  a15666a );
 a15670a <=( A199  and  (not A166) );
 a15673a <=( A232  and  A200 );
 a15674a <=( a15673a  and  a15670a );
 a15675a <=( a15674a  and  a15667a );
 a15679a <=( A235  and  A234 );
 a15680a <=( (not A233)  and  a15679a );
 a15683a <=( (not A299)  and  A298 );
 a15686a <=( A302  and  A300 );
 a15687a <=( a15686a  and  a15683a );
 a15688a <=( a15687a  and  a15680a );
 a15692a <=( A167  and  A168 );
 a15693a <=( A169  and  a15692a );
 a15696a <=( A199  and  (not A166) );
 a15699a <=( A232  and  A200 );
 a15700a <=( a15699a  and  a15696a );
 a15701a <=( a15700a  and  a15693a );
 a15705a <=( A235  and  A234 );
 a15706a <=( (not A233)  and  a15705a );
 a15709a <=( A299  and  (not A298) );
 a15712a <=( A301  and  A300 );
 a15713a <=( a15712a  and  a15709a );
 a15714a <=( a15713a  and  a15706a );
 a15718a <=( A167  and  A168 );
 a15719a <=( A169  and  a15718a );
 a15722a <=( A199  and  (not A166) );
 a15725a <=( A232  and  A200 );
 a15726a <=( a15725a  and  a15722a );
 a15727a <=( a15726a  and  a15719a );
 a15731a <=( A235  and  A234 );
 a15732a <=( (not A233)  and  a15731a );
 a15735a <=( A299  and  (not A298) );
 a15738a <=( A302  and  A300 );
 a15739a <=( a15738a  and  a15735a );
 a15740a <=( a15739a  and  a15732a );
 a15744a <=( A167  and  A168 );
 a15745a <=( A169  and  a15744a );
 a15748a <=( A199  and  (not A166) );
 a15751a <=( A232  and  A200 );
 a15752a <=( a15751a  and  a15748a );
 a15753a <=( a15752a  and  a15745a );
 a15757a <=( A235  and  A234 );
 a15758a <=( (not A233)  and  a15757a );
 a15761a <=( A266  and  (not A265) );
 a15764a <=( A268  and  A267 );
 a15765a <=( a15764a  and  a15761a );
 a15766a <=( a15765a  and  a15758a );
 a15770a <=( A167  and  A168 );
 a15771a <=( A169  and  a15770a );
 a15774a <=( A199  and  (not A166) );
 a15777a <=( A232  and  A200 );
 a15778a <=( a15777a  and  a15774a );
 a15779a <=( a15778a  and  a15771a );
 a15783a <=( A235  and  A234 );
 a15784a <=( (not A233)  and  a15783a );
 a15787a <=( A266  and  (not A265) );
 a15790a <=( A269  and  A267 );
 a15791a <=( a15790a  and  a15787a );
 a15792a <=( a15791a  and  a15784a );
 a15796a <=( A167  and  A168 );
 a15797a <=( A169  and  a15796a );
 a15800a <=( A199  and  (not A166) );
 a15803a <=( A232  and  A200 );
 a15804a <=( a15803a  and  a15800a );
 a15805a <=( a15804a  and  a15797a );
 a15809a <=( A235  and  A234 );
 a15810a <=( (not A233)  and  a15809a );
 a15813a <=( (not A266)  and  A265 );
 a15816a <=( A268  and  A267 );
 a15817a <=( a15816a  and  a15813a );
 a15818a <=( a15817a  and  a15810a );
 a15822a <=( A167  and  A168 );
 a15823a <=( A169  and  a15822a );
 a15826a <=( A199  and  (not A166) );
 a15829a <=( A232  and  A200 );
 a15830a <=( a15829a  and  a15826a );
 a15831a <=( a15830a  and  a15823a );
 a15835a <=( A235  and  A234 );
 a15836a <=( (not A233)  and  a15835a );
 a15839a <=( (not A266)  and  A265 );
 a15842a <=( A269  and  A267 );
 a15843a <=( a15842a  and  a15839a );
 a15844a <=( a15843a  and  a15836a );
 a15848a <=( A167  and  A168 );
 a15849a <=( A169  and  a15848a );
 a15852a <=( A199  and  (not A166) );
 a15855a <=( A232  and  A200 );
 a15856a <=( a15855a  and  a15852a );
 a15857a <=( a15856a  and  a15849a );
 a15861a <=( A236  and  A234 );
 a15862a <=( (not A233)  and  a15861a );
 a15865a <=( (not A299)  and  A298 );
 a15868a <=( A301  and  A300 );
 a15869a <=( a15868a  and  a15865a );
 a15870a <=( a15869a  and  a15862a );
 a15874a <=( A167  and  A168 );
 a15875a <=( A169  and  a15874a );
 a15878a <=( A199  and  (not A166) );
 a15881a <=( A232  and  A200 );
 a15882a <=( a15881a  and  a15878a );
 a15883a <=( a15882a  and  a15875a );
 a15887a <=( A236  and  A234 );
 a15888a <=( (not A233)  and  a15887a );
 a15891a <=( (not A299)  and  A298 );
 a15894a <=( A302  and  A300 );
 a15895a <=( a15894a  and  a15891a );
 a15896a <=( a15895a  and  a15888a );
 a15900a <=( A167  and  A168 );
 a15901a <=( A169  and  a15900a );
 a15904a <=( A199  and  (not A166) );
 a15907a <=( A232  and  A200 );
 a15908a <=( a15907a  and  a15904a );
 a15909a <=( a15908a  and  a15901a );
 a15913a <=( A236  and  A234 );
 a15914a <=( (not A233)  and  a15913a );
 a15917a <=( A299  and  (not A298) );
 a15920a <=( A301  and  A300 );
 a15921a <=( a15920a  and  a15917a );
 a15922a <=( a15921a  and  a15914a );
 a15926a <=( A167  and  A168 );
 a15927a <=( A169  and  a15926a );
 a15930a <=( A199  and  (not A166) );
 a15933a <=( A232  and  A200 );
 a15934a <=( a15933a  and  a15930a );
 a15935a <=( a15934a  and  a15927a );
 a15939a <=( A236  and  A234 );
 a15940a <=( (not A233)  and  a15939a );
 a15943a <=( A299  and  (not A298) );
 a15946a <=( A302  and  A300 );
 a15947a <=( a15946a  and  a15943a );
 a15948a <=( a15947a  and  a15940a );
 a15952a <=( A167  and  A168 );
 a15953a <=( A169  and  a15952a );
 a15956a <=( A199  and  (not A166) );
 a15959a <=( A232  and  A200 );
 a15960a <=( a15959a  and  a15956a );
 a15961a <=( a15960a  and  a15953a );
 a15965a <=( A236  and  A234 );
 a15966a <=( (not A233)  and  a15965a );
 a15969a <=( A266  and  (not A265) );
 a15972a <=( A268  and  A267 );
 a15973a <=( a15972a  and  a15969a );
 a15974a <=( a15973a  and  a15966a );
 a15978a <=( A167  and  A168 );
 a15979a <=( A169  and  a15978a );
 a15982a <=( A199  and  (not A166) );
 a15985a <=( A232  and  A200 );
 a15986a <=( a15985a  and  a15982a );
 a15987a <=( a15986a  and  a15979a );
 a15991a <=( A236  and  A234 );
 a15992a <=( (not A233)  and  a15991a );
 a15995a <=( A266  and  (not A265) );
 a15998a <=( A269  and  A267 );
 a15999a <=( a15998a  and  a15995a );
 a16000a <=( a15999a  and  a15992a );
 a16004a <=( A167  and  A168 );
 a16005a <=( A169  and  a16004a );
 a16008a <=( A199  and  (not A166) );
 a16011a <=( A232  and  A200 );
 a16012a <=( a16011a  and  a16008a );
 a16013a <=( a16012a  and  a16005a );
 a16017a <=( A236  and  A234 );
 a16018a <=( (not A233)  and  a16017a );
 a16021a <=( (not A266)  and  A265 );
 a16024a <=( A268  and  A267 );
 a16025a <=( a16024a  and  a16021a );
 a16026a <=( a16025a  and  a16018a );
 a16030a <=( A167  and  A168 );
 a16031a <=( A169  and  a16030a );
 a16034a <=( A199  and  (not A166) );
 a16037a <=( A232  and  A200 );
 a16038a <=( a16037a  and  a16034a );
 a16039a <=( a16038a  and  a16031a );
 a16043a <=( A236  and  A234 );
 a16044a <=( (not A233)  and  a16043a );
 a16047a <=( (not A266)  and  A265 );
 a16050a <=( A269  and  A267 );
 a16051a <=( a16050a  and  a16047a );
 a16052a <=( a16051a  and  a16044a );
 a16056a <=( A167  and  A168 );
 a16057a <=( A169  and  a16056a );
 a16060a <=( (not A199)  and  (not A166) );
 a16063a <=( (not A232)  and  (not A200) );
 a16064a <=( a16063a  and  a16060a );
 a16065a <=( a16064a  and  a16057a );
 a16069a <=( A235  and  A234 );
 a16070a <=( A233  and  a16069a );
 a16073a <=( (not A299)  and  A298 );
 a16076a <=( A301  and  A300 );
 a16077a <=( a16076a  and  a16073a );
 a16078a <=( a16077a  and  a16070a );
 a16082a <=( A167  and  A168 );
 a16083a <=( A169  and  a16082a );
 a16086a <=( (not A199)  and  (not A166) );
 a16089a <=( (not A232)  and  (not A200) );
 a16090a <=( a16089a  and  a16086a );
 a16091a <=( a16090a  and  a16083a );
 a16095a <=( A235  and  A234 );
 a16096a <=( A233  and  a16095a );
 a16099a <=( (not A299)  and  A298 );
 a16102a <=( A302  and  A300 );
 a16103a <=( a16102a  and  a16099a );
 a16104a <=( a16103a  and  a16096a );
 a16108a <=( A167  and  A168 );
 a16109a <=( A169  and  a16108a );
 a16112a <=( (not A199)  and  (not A166) );
 a16115a <=( (not A232)  and  (not A200) );
 a16116a <=( a16115a  and  a16112a );
 a16117a <=( a16116a  and  a16109a );
 a16121a <=( A235  and  A234 );
 a16122a <=( A233  and  a16121a );
 a16125a <=( A299  and  (not A298) );
 a16128a <=( A301  and  A300 );
 a16129a <=( a16128a  and  a16125a );
 a16130a <=( a16129a  and  a16122a );
 a16134a <=( A167  and  A168 );
 a16135a <=( A169  and  a16134a );
 a16138a <=( (not A199)  and  (not A166) );
 a16141a <=( (not A232)  and  (not A200) );
 a16142a <=( a16141a  and  a16138a );
 a16143a <=( a16142a  and  a16135a );
 a16147a <=( A235  and  A234 );
 a16148a <=( A233  and  a16147a );
 a16151a <=( A299  and  (not A298) );
 a16154a <=( A302  and  A300 );
 a16155a <=( a16154a  and  a16151a );
 a16156a <=( a16155a  and  a16148a );
 a16160a <=( A167  and  A168 );
 a16161a <=( A169  and  a16160a );
 a16164a <=( (not A199)  and  (not A166) );
 a16167a <=( (not A232)  and  (not A200) );
 a16168a <=( a16167a  and  a16164a );
 a16169a <=( a16168a  and  a16161a );
 a16173a <=( A235  and  A234 );
 a16174a <=( A233  and  a16173a );
 a16177a <=( A266  and  (not A265) );
 a16180a <=( A268  and  A267 );
 a16181a <=( a16180a  and  a16177a );
 a16182a <=( a16181a  and  a16174a );
 a16186a <=( A167  and  A168 );
 a16187a <=( A169  and  a16186a );
 a16190a <=( (not A199)  and  (not A166) );
 a16193a <=( (not A232)  and  (not A200) );
 a16194a <=( a16193a  and  a16190a );
 a16195a <=( a16194a  and  a16187a );
 a16199a <=( A235  and  A234 );
 a16200a <=( A233  and  a16199a );
 a16203a <=( A266  and  (not A265) );
 a16206a <=( A269  and  A267 );
 a16207a <=( a16206a  and  a16203a );
 a16208a <=( a16207a  and  a16200a );
 a16212a <=( A167  and  A168 );
 a16213a <=( A169  and  a16212a );
 a16216a <=( (not A199)  and  (not A166) );
 a16219a <=( (not A232)  and  (not A200) );
 a16220a <=( a16219a  and  a16216a );
 a16221a <=( a16220a  and  a16213a );
 a16225a <=( A235  and  A234 );
 a16226a <=( A233  and  a16225a );
 a16229a <=( (not A266)  and  A265 );
 a16232a <=( A268  and  A267 );
 a16233a <=( a16232a  and  a16229a );
 a16234a <=( a16233a  and  a16226a );
 a16238a <=( A167  and  A168 );
 a16239a <=( A169  and  a16238a );
 a16242a <=( (not A199)  and  (not A166) );
 a16245a <=( (not A232)  and  (not A200) );
 a16246a <=( a16245a  and  a16242a );
 a16247a <=( a16246a  and  a16239a );
 a16251a <=( A235  and  A234 );
 a16252a <=( A233  and  a16251a );
 a16255a <=( (not A266)  and  A265 );
 a16258a <=( A269  and  A267 );
 a16259a <=( a16258a  and  a16255a );
 a16260a <=( a16259a  and  a16252a );
 a16264a <=( A167  and  A168 );
 a16265a <=( A169  and  a16264a );
 a16268a <=( (not A199)  and  (not A166) );
 a16271a <=( (not A232)  and  (not A200) );
 a16272a <=( a16271a  and  a16268a );
 a16273a <=( a16272a  and  a16265a );
 a16277a <=( A236  and  A234 );
 a16278a <=( A233  and  a16277a );
 a16281a <=( (not A299)  and  A298 );
 a16284a <=( A301  and  A300 );
 a16285a <=( a16284a  and  a16281a );
 a16286a <=( a16285a  and  a16278a );
 a16290a <=( A167  and  A168 );
 a16291a <=( A169  and  a16290a );
 a16294a <=( (not A199)  and  (not A166) );
 a16297a <=( (not A232)  and  (not A200) );
 a16298a <=( a16297a  and  a16294a );
 a16299a <=( a16298a  and  a16291a );
 a16303a <=( A236  and  A234 );
 a16304a <=( A233  and  a16303a );
 a16307a <=( (not A299)  and  A298 );
 a16310a <=( A302  and  A300 );
 a16311a <=( a16310a  and  a16307a );
 a16312a <=( a16311a  and  a16304a );
 a16316a <=( A167  and  A168 );
 a16317a <=( A169  and  a16316a );
 a16320a <=( (not A199)  and  (not A166) );
 a16323a <=( (not A232)  and  (not A200) );
 a16324a <=( a16323a  and  a16320a );
 a16325a <=( a16324a  and  a16317a );
 a16329a <=( A236  and  A234 );
 a16330a <=( A233  and  a16329a );
 a16333a <=( A299  and  (not A298) );
 a16336a <=( A301  and  A300 );
 a16337a <=( a16336a  and  a16333a );
 a16338a <=( a16337a  and  a16330a );
 a16342a <=( A167  and  A168 );
 a16343a <=( A169  and  a16342a );
 a16346a <=( (not A199)  and  (not A166) );
 a16349a <=( (not A232)  and  (not A200) );
 a16350a <=( a16349a  and  a16346a );
 a16351a <=( a16350a  and  a16343a );
 a16355a <=( A236  and  A234 );
 a16356a <=( A233  and  a16355a );
 a16359a <=( A299  and  (not A298) );
 a16362a <=( A302  and  A300 );
 a16363a <=( a16362a  and  a16359a );
 a16364a <=( a16363a  and  a16356a );
 a16368a <=( A167  and  A168 );
 a16369a <=( A169  and  a16368a );
 a16372a <=( (not A199)  and  (not A166) );
 a16375a <=( (not A232)  and  (not A200) );
 a16376a <=( a16375a  and  a16372a );
 a16377a <=( a16376a  and  a16369a );
 a16381a <=( A236  and  A234 );
 a16382a <=( A233  and  a16381a );
 a16385a <=( A266  and  (not A265) );
 a16388a <=( A268  and  A267 );
 a16389a <=( a16388a  and  a16385a );
 a16390a <=( a16389a  and  a16382a );
 a16394a <=( A167  and  A168 );
 a16395a <=( A169  and  a16394a );
 a16398a <=( (not A199)  and  (not A166) );
 a16401a <=( (not A232)  and  (not A200) );
 a16402a <=( a16401a  and  a16398a );
 a16403a <=( a16402a  and  a16395a );
 a16407a <=( A236  and  A234 );
 a16408a <=( A233  and  a16407a );
 a16411a <=( A266  and  (not A265) );
 a16414a <=( A269  and  A267 );
 a16415a <=( a16414a  and  a16411a );
 a16416a <=( a16415a  and  a16408a );
 a16420a <=( A167  and  A168 );
 a16421a <=( A169  and  a16420a );
 a16424a <=( (not A199)  and  (not A166) );
 a16427a <=( (not A232)  and  (not A200) );
 a16428a <=( a16427a  and  a16424a );
 a16429a <=( a16428a  and  a16421a );
 a16433a <=( A236  and  A234 );
 a16434a <=( A233  and  a16433a );
 a16437a <=( (not A266)  and  A265 );
 a16440a <=( A268  and  A267 );
 a16441a <=( a16440a  and  a16437a );
 a16442a <=( a16441a  and  a16434a );
 a16446a <=( A167  and  A168 );
 a16447a <=( A169  and  a16446a );
 a16450a <=( (not A199)  and  (not A166) );
 a16453a <=( (not A232)  and  (not A200) );
 a16454a <=( a16453a  and  a16450a );
 a16455a <=( a16454a  and  a16447a );
 a16459a <=( A236  and  A234 );
 a16460a <=( A233  and  a16459a );
 a16463a <=( (not A266)  and  A265 );
 a16466a <=( A269  and  A267 );
 a16467a <=( a16466a  and  a16463a );
 a16468a <=( a16467a  and  a16460a );
 a16472a <=( A167  and  A168 );
 a16473a <=( A169  and  a16472a );
 a16476a <=( (not A199)  and  (not A166) );
 a16479a <=( A232  and  (not A200) );
 a16480a <=( a16479a  and  a16476a );
 a16481a <=( a16480a  and  a16473a );
 a16485a <=( A235  and  A234 );
 a16486a <=( (not A233)  and  a16485a );
 a16489a <=( (not A299)  and  A298 );
 a16492a <=( A301  and  A300 );
 a16493a <=( a16492a  and  a16489a );
 a16494a <=( a16493a  and  a16486a );
 a16498a <=( A167  and  A168 );
 a16499a <=( A169  and  a16498a );
 a16502a <=( (not A199)  and  (not A166) );
 a16505a <=( A232  and  (not A200) );
 a16506a <=( a16505a  and  a16502a );
 a16507a <=( a16506a  and  a16499a );
 a16511a <=( A235  and  A234 );
 a16512a <=( (not A233)  and  a16511a );
 a16515a <=( (not A299)  and  A298 );
 a16518a <=( A302  and  A300 );
 a16519a <=( a16518a  and  a16515a );
 a16520a <=( a16519a  and  a16512a );
 a16524a <=( A167  and  A168 );
 a16525a <=( A169  and  a16524a );
 a16528a <=( (not A199)  and  (not A166) );
 a16531a <=( A232  and  (not A200) );
 a16532a <=( a16531a  and  a16528a );
 a16533a <=( a16532a  and  a16525a );
 a16537a <=( A235  and  A234 );
 a16538a <=( (not A233)  and  a16537a );
 a16541a <=( A299  and  (not A298) );
 a16544a <=( A301  and  A300 );
 a16545a <=( a16544a  and  a16541a );
 a16546a <=( a16545a  and  a16538a );
 a16550a <=( A167  and  A168 );
 a16551a <=( A169  and  a16550a );
 a16554a <=( (not A199)  and  (not A166) );
 a16557a <=( A232  and  (not A200) );
 a16558a <=( a16557a  and  a16554a );
 a16559a <=( a16558a  and  a16551a );
 a16563a <=( A235  and  A234 );
 a16564a <=( (not A233)  and  a16563a );
 a16567a <=( A299  and  (not A298) );
 a16570a <=( A302  and  A300 );
 a16571a <=( a16570a  and  a16567a );
 a16572a <=( a16571a  and  a16564a );
 a16576a <=( A167  and  A168 );
 a16577a <=( A169  and  a16576a );
 a16580a <=( (not A199)  and  (not A166) );
 a16583a <=( A232  and  (not A200) );
 a16584a <=( a16583a  and  a16580a );
 a16585a <=( a16584a  and  a16577a );
 a16589a <=( A235  and  A234 );
 a16590a <=( (not A233)  and  a16589a );
 a16593a <=( A266  and  (not A265) );
 a16596a <=( A268  and  A267 );
 a16597a <=( a16596a  and  a16593a );
 a16598a <=( a16597a  and  a16590a );
 a16602a <=( A167  and  A168 );
 a16603a <=( A169  and  a16602a );
 a16606a <=( (not A199)  and  (not A166) );
 a16609a <=( A232  and  (not A200) );
 a16610a <=( a16609a  and  a16606a );
 a16611a <=( a16610a  and  a16603a );
 a16615a <=( A235  and  A234 );
 a16616a <=( (not A233)  and  a16615a );
 a16619a <=( A266  and  (not A265) );
 a16622a <=( A269  and  A267 );
 a16623a <=( a16622a  and  a16619a );
 a16624a <=( a16623a  and  a16616a );
 a16628a <=( A167  and  A168 );
 a16629a <=( A169  and  a16628a );
 a16632a <=( (not A199)  and  (not A166) );
 a16635a <=( A232  and  (not A200) );
 a16636a <=( a16635a  and  a16632a );
 a16637a <=( a16636a  and  a16629a );
 a16641a <=( A235  and  A234 );
 a16642a <=( (not A233)  and  a16641a );
 a16645a <=( (not A266)  and  A265 );
 a16648a <=( A268  and  A267 );
 a16649a <=( a16648a  and  a16645a );
 a16650a <=( a16649a  and  a16642a );
 a16654a <=( A167  and  A168 );
 a16655a <=( A169  and  a16654a );
 a16658a <=( (not A199)  and  (not A166) );
 a16661a <=( A232  and  (not A200) );
 a16662a <=( a16661a  and  a16658a );
 a16663a <=( a16662a  and  a16655a );
 a16667a <=( A235  and  A234 );
 a16668a <=( (not A233)  and  a16667a );
 a16671a <=( (not A266)  and  A265 );
 a16674a <=( A269  and  A267 );
 a16675a <=( a16674a  and  a16671a );
 a16676a <=( a16675a  and  a16668a );
 a16680a <=( A167  and  A168 );
 a16681a <=( A169  and  a16680a );
 a16684a <=( (not A199)  and  (not A166) );
 a16687a <=( A232  and  (not A200) );
 a16688a <=( a16687a  and  a16684a );
 a16689a <=( a16688a  and  a16681a );
 a16693a <=( A236  and  A234 );
 a16694a <=( (not A233)  and  a16693a );
 a16697a <=( (not A299)  and  A298 );
 a16700a <=( A301  and  A300 );
 a16701a <=( a16700a  and  a16697a );
 a16702a <=( a16701a  and  a16694a );
 a16706a <=( A167  and  A168 );
 a16707a <=( A169  and  a16706a );
 a16710a <=( (not A199)  and  (not A166) );
 a16713a <=( A232  and  (not A200) );
 a16714a <=( a16713a  and  a16710a );
 a16715a <=( a16714a  and  a16707a );
 a16719a <=( A236  and  A234 );
 a16720a <=( (not A233)  and  a16719a );
 a16723a <=( (not A299)  and  A298 );
 a16726a <=( A302  and  A300 );
 a16727a <=( a16726a  and  a16723a );
 a16728a <=( a16727a  and  a16720a );
 a16732a <=( A167  and  A168 );
 a16733a <=( A169  and  a16732a );
 a16736a <=( (not A199)  and  (not A166) );
 a16739a <=( A232  and  (not A200) );
 a16740a <=( a16739a  and  a16736a );
 a16741a <=( a16740a  and  a16733a );
 a16745a <=( A236  and  A234 );
 a16746a <=( (not A233)  and  a16745a );
 a16749a <=( A299  and  (not A298) );
 a16752a <=( A301  and  A300 );
 a16753a <=( a16752a  and  a16749a );
 a16754a <=( a16753a  and  a16746a );
 a16758a <=( A167  and  A168 );
 a16759a <=( A169  and  a16758a );
 a16762a <=( (not A199)  and  (not A166) );
 a16765a <=( A232  and  (not A200) );
 a16766a <=( a16765a  and  a16762a );
 a16767a <=( a16766a  and  a16759a );
 a16771a <=( A236  and  A234 );
 a16772a <=( (not A233)  and  a16771a );
 a16775a <=( A299  and  (not A298) );
 a16778a <=( A302  and  A300 );
 a16779a <=( a16778a  and  a16775a );
 a16780a <=( a16779a  and  a16772a );
 a16784a <=( A167  and  A168 );
 a16785a <=( A169  and  a16784a );
 a16788a <=( (not A199)  and  (not A166) );
 a16791a <=( A232  and  (not A200) );
 a16792a <=( a16791a  and  a16788a );
 a16793a <=( a16792a  and  a16785a );
 a16797a <=( A236  and  A234 );
 a16798a <=( (not A233)  and  a16797a );
 a16801a <=( A266  and  (not A265) );
 a16804a <=( A268  and  A267 );
 a16805a <=( a16804a  and  a16801a );
 a16806a <=( a16805a  and  a16798a );
 a16810a <=( A167  and  A168 );
 a16811a <=( A169  and  a16810a );
 a16814a <=( (not A199)  and  (not A166) );
 a16817a <=( A232  and  (not A200) );
 a16818a <=( a16817a  and  a16814a );
 a16819a <=( a16818a  and  a16811a );
 a16823a <=( A236  and  A234 );
 a16824a <=( (not A233)  and  a16823a );
 a16827a <=( A266  and  (not A265) );
 a16830a <=( A269  and  A267 );
 a16831a <=( a16830a  and  a16827a );
 a16832a <=( a16831a  and  a16824a );
 a16836a <=( A167  and  A168 );
 a16837a <=( A169  and  a16836a );
 a16840a <=( (not A199)  and  (not A166) );
 a16843a <=( A232  and  (not A200) );
 a16844a <=( a16843a  and  a16840a );
 a16845a <=( a16844a  and  a16837a );
 a16849a <=( A236  and  A234 );
 a16850a <=( (not A233)  and  a16849a );
 a16853a <=( (not A266)  and  A265 );
 a16856a <=( A268  and  A267 );
 a16857a <=( a16856a  and  a16853a );
 a16858a <=( a16857a  and  a16850a );
 a16862a <=( A167  and  A168 );
 a16863a <=( A169  and  a16862a );
 a16866a <=( (not A199)  and  (not A166) );
 a16869a <=( A232  and  (not A200) );
 a16870a <=( a16869a  and  a16866a );
 a16871a <=( a16870a  and  a16863a );
 a16875a <=( A236  and  A234 );
 a16876a <=( (not A233)  and  a16875a );
 a16879a <=( (not A266)  and  A265 );
 a16882a <=( A269  and  A267 );
 a16883a <=( a16882a  and  a16879a );
 a16884a <=( a16883a  and  a16876a );
 a16888a <=( (not A167)  and  A168 );
 a16889a <=( A169  and  a16888a );
 a16892a <=( (not A201)  and  A166 );
 a16895a <=( (not A232)  and  A202 );
 a16896a <=( a16895a  and  a16892a );
 a16897a <=( a16896a  and  a16889a );
 a16901a <=( A235  and  A234 );
 a16902a <=( A233  and  a16901a );
 a16905a <=( (not A299)  and  A298 );
 a16908a <=( A301  and  A300 );
 a16909a <=( a16908a  and  a16905a );
 a16910a <=( a16909a  and  a16902a );
 a16914a <=( (not A167)  and  A168 );
 a16915a <=( A169  and  a16914a );
 a16918a <=( (not A201)  and  A166 );
 a16921a <=( (not A232)  and  A202 );
 a16922a <=( a16921a  and  a16918a );
 a16923a <=( a16922a  and  a16915a );
 a16927a <=( A235  and  A234 );
 a16928a <=( A233  and  a16927a );
 a16931a <=( (not A299)  and  A298 );
 a16934a <=( A302  and  A300 );
 a16935a <=( a16934a  and  a16931a );
 a16936a <=( a16935a  and  a16928a );
 a16940a <=( (not A167)  and  A168 );
 a16941a <=( A169  and  a16940a );
 a16944a <=( (not A201)  and  A166 );
 a16947a <=( (not A232)  and  A202 );
 a16948a <=( a16947a  and  a16944a );
 a16949a <=( a16948a  and  a16941a );
 a16953a <=( A235  and  A234 );
 a16954a <=( A233  and  a16953a );
 a16957a <=( A299  and  (not A298) );
 a16960a <=( A301  and  A300 );
 a16961a <=( a16960a  and  a16957a );
 a16962a <=( a16961a  and  a16954a );
 a16966a <=( (not A167)  and  A168 );
 a16967a <=( A169  and  a16966a );
 a16970a <=( (not A201)  and  A166 );
 a16973a <=( (not A232)  and  A202 );
 a16974a <=( a16973a  and  a16970a );
 a16975a <=( a16974a  and  a16967a );
 a16979a <=( A235  and  A234 );
 a16980a <=( A233  and  a16979a );
 a16983a <=( A299  and  (not A298) );
 a16986a <=( A302  and  A300 );
 a16987a <=( a16986a  and  a16983a );
 a16988a <=( a16987a  and  a16980a );
 a16992a <=( (not A167)  and  A168 );
 a16993a <=( A169  and  a16992a );
 a16996a <=( (not A201)  and  A166 );
 a16999a <=( (not A232)  and  A202 );
 a17000a <=( a16999a  and  a16996a );
 a17001a <=( a17000a  and  a16993a );
 a17005a <=( A235  and  A234 );
 a17006a <=( A233  and  a17005a );
 a17009a <=( A266  and  (not A265) );
 a17012a <=( A268  and  A267 );
 a17013a <=( a17012a  and  a17009a );
 a17014a <=( a17013a  and  a17006a );
 a17018a <=( (not A167)  and  A168 );
 a17019a <=( A169  and  a17018a );
 a17022a <=( (not A201)  and  A166 );
 a17025a <=( (not A232)  and  A202 );
 a17026a <=( a17025a  and  a17022a );
 a17027a <=( a17026a  and  a17019a );
 a17031a <=( A235  and  A234 );
 a17032a <=( A233  and  a17031a );
 a17035a <=( A266  and  (not A265) );
 a17038a <=( A269  and  A267 );
 a17039a <=( a17038a  and  a17035a );
 a17040a <=( a17039a  and  a17032a );
 a17044a <=( (not A167)  and  A168 );
 a17045a <=( A169  and  a17044a );
 a17048a <=( (not A201)  and  A166 );
 a17051a <=( (not A232)  and  A202 );
 a17052a <=( a17051a  and  a17048a );
 a17053a <=( a17052a  and  a17045a );
 a17057a <=( A235  and  A234 );
 a17058a <=( A233  and  a17057a );
 a17061a <=( (not A266)  and  A265 );
 a17064a <=( A268  and  A267 );
 a17065a <=( a17064a  and  a17061a );
 a17066a <=( a17065a  and  a17058a );
 a17070a <=( (not A167)  and  A168 );
 a17071a <=( A169  and  a17070a );
 a17074a <=( (not A201)  and  A166 );
 a17077a <=( (not A232)  and  A202 );
 a17078a <=( a17077a  and  a17074a );
 a17079a <=( a17078a  and  a17071a );
 a17083a <=( A235  and  A234 );
 a17084a <=( A233  and  a17083a );
 a17087a <=( (not A266)  and  A265 );
 a17090a <=( A269  and  A267 );
 a17091a <=( a17090a  and  a17087a );
 a17092a <=( a17091a  and  a17084a );
 a17096a <=( (not A167)  and  A168 );
 a17097a <=( A169  and  a17096a );
 a17100a <=( (not A201)  and  A166 );
 a17103a <=( (not A232)  and  A202 );
 a17104a <=( a17103a  and  a17100a );
 a17105a <=( a17104a  and  a17097a );
 a17109a <=( A236  and  A234 );
 a17110a <=( A233  and  a17109a );
 a17113a <=( (not A299)  and  A298 );
 a17116a <=( A301  and  A300 );
 a17117a <=( a17116a  and  a17113a );
 a17118a <=( a17117a  and  a17110a );
 a17122a <=( (not A167)  and  A168 );
 a17123a <=( A169  and  a17122a );
 a17126a <=( (not A201)  and  A166 );
 a17129a <=( (not A232)  and  A202 );
 a17130a <=( a17129a  and  a17126a );
 a17131a <=( a17130a  and  a17123a );
 a17135a <=( A236  and  A234 );
 a17136a <=( A233  and  a17135a );
 a17139a <=( (not A299)  and  A298 );
 a17142a <=( A302  and  A300 );
 a17143a <=( a17142a  and  a17139a );
 a17144a <=( a17143a  and  a17136a );
 a17148a <=( (not A167)  and  A168 );
 a17149a <=( A169  and  a17148a );
 a17152a <=( (not A201)  and  A166 );
 a17155a <=( (not A232)  and  A202 );
 a17156a <=( a17155a  and  a17152a );
 a17157a <=( a17156a  and  a17149a );
 a17161a <=( A236  and  A234 );
 a17162a <=( A233  and  a17161a );
 a17165a <=( A299  and  (not A298) );
 a17168a <=( A301  and  A300 );
 a17169a <=( a17168a  and  a17165a );
 a17170a <=( a17169a  and  a17162a );
 a17174a <=( (not A167)  and  A168 );
 a17175a <=( A169  and  a17174a );
 a17178a <=( (not A201)  and  A166 );
 a17181a <=( (not A232)  and  A202 );
 a17182a <=( a17181a  and  a17178a );
 a17183a <=( a17182a  and  a17175a );
 a17187a <=( A236  and  A234 );
 a17188a <=( A233  and  a17187a );
 a17191a <=( A299  and  (not A298) );
 a17194a <=( A302  and  A300 );
 a17195a <=( a17194a  and  a17191a );
 a17196a <=( a17195a  and  a17188a );
 a17200a <=( (not A167)  and  A168 );
 a17201a <=( A169  and  a17200a );
 a17204a <=( (not A201)  and  A166 );
 a17207a <=( (not A232)  and  A202 );
 a17208a <=( a17207a  and  a17204a );
 a17209a <=( a17208a  and  a17201a );
 a17213a <=( A236  and  A234 );
 a17214a <=( A233  and  a17213a );
 a17217a <=( A266  and  (not A265) );
 a17220a <=( A268  and  A267 );
 a17221a <=( a17220a  and  a17217a );
 a17222a <=( a17221a  and  a17214a );
 a17226a <=( (not A167)  and  A168 );
 a17227a <=( A169  and  a17226a );
 a17230a <=( (not A201)  and  A166 );
 a17233a <=( (not A232)  and  A202 );
 a17234a <=( a17233a  and  a17230a );
 a17235a <=( a17234a  and  a17227a );
 a17239a <=( A236  and  A234 );
 a17240a <=( A233  and  a17239a );
 a17243a <=( A266  and  (not A265) );
 a17246a <=( A269  and  A267 );
 a17247a <=( a17246a  and  a17243a );
 a17248a <=( a17247a  and  a17240a );
 a17252a <=( (not A167)  and  A168 );
 a17253a <=( A169  and  a17252a );
 a17256a <=( (not A201)  and  A166 );
 a17259a <=( (not A232)  and  A202 );
 a17260a <=( a17259a  and  a17256a );
 a17261a <=( a17260a  and  a17253a );
 a17265a <=( A236  and  A234 );
 a17266a <=( A233  and  a17265a );
 a17269a <=( (not A266)  and  A265 );
 a17272a <=( A268  and  A267 );
 a17273a <=( a17272a  and  a17269a );
 a17274a <=( a17273a  and  a17266a );
 a17278a <=( (not A167)  and  A168 );
 a17279a <=( A169  and  a17278a );
 a17282a <=( (not A201)  and  A166 );
 a17285a <=( (not A232)  and  A202 );
 a17286a <=( a17285a  and  a17282a );
 a17287a <=( a17286a  and  a17279a );
 a17291a <=( A236  and  A234 );
 a17292a <=( A233  and  a17291a );
 a17295a <=( (not A266)  and  A265 );
 a17298a <=( A269  and  A267 );
 a17299a <=( a17298a  and  a17295a );
 a17300a <=( a17299a  and  a17292a );
 a17304a <=( (not A167)  and  A168 );
 a17305a <=( A169  and  a17304a );
 a17308a <=( (not A201)  and  A166 );
 a17311a <=( A232  and  A202 );
 a17312a <=( a17311a  and  a17308a );
 a17313a <=( a17312a  and  a17305a );
 a17317a <=( A235  and  A234 );
 a17318a <=( (not A233)  and  a17317a );
 a17321a <=( (not A299)  and  A298 );
 a17324a <=( A301  and  A300 );
 a17325a <=( a17324a  and  a17321a );
 a17326a <=( a17325a  and  a17318a );
 a17330a <=( (not A167)  and  A168 );
 a17331a <=( A169  and  a17330a );
 a17334a <=( (not A201)  and  A166 );
 a17337a <=( A232  and  A202 );
 a17338a <=( a17337a  and  a17334a );
 a17339a <=( a17338a  and  a17331a );
 a17343a <=( A235  and  A234 );
 a17344a <=( (not A233)  and  a17343a );
 a17347a <=( (not A299)  and  A298 );
 a17350a <=( A302  and  A300 );
 a17351a <=( a17350a  and  a17347a );
 a17352a <=( a17351a  and  a17344a );
 a17356a <=( (not A167)  and  A168 );
 a17357a <=( A169  and  a17356a );
 a17360a <=( (not A201)  and  A166 );
 a17363a <=( A232  and  A202 );
 a17364a <=( a17363a  and  a17360a );
 a17365a <=( a17364a  and  a17357a );
 a17369a <=( A235  and  A234 );
 a17370a <=( (not A233)  and  a17369a );
 a17373a <=( A299  and  (not A298) );
 a17376a <=( A301  and  A300 );
 a17377a <=( a17376a  and  a17373a );
 a17378a <=( a17377a  and  a17370a );
 a17382a <=( (not A167)  and  A168 );
 a17383a <=( A169  and  a17382a );
 a17386a <=( (not A201)  and  A166 );
 a17389a <=( A232  and  A202 );
 a17390a <=( a17389a  and  a17386a );
 a17391a <=( a17390a  and  a17383a );
 a17395a <=( A235  and  A234 );
 a17396a <=( (not A233)  and  a17395a );
 a17399a <=( A299  and  (not A298) );
 a17402a <=( A302  and  A300 );
 a17403a <=( a17402a  and  a17399a );
 a17404a <=( a17403a  and  a17396a );
 a17408a <=( (not A167)  and  A168 );
 a17409a <=( A169  and  a17408a );
 a17412a <=( (not A201)  and  A166 );
 a17415a <=( A232  and  A202 );
 a17416a <=( a17415a  and  a17412a );
 a17417a <=( a17416a  and  a17409a );
 a17421a <=( A235  and  A234 );
 a17422a <=( (not A233)  and  a17421a );
 a17425a <=( A266  and  (not A265) );
 a17428a <=( A268  and  A267 );
 a17429a <=( a17428a  and  a17425a );
 a17430a <=( a17429a  and  a17422a );
 a17434a <=( (not A167)  and  A168 );
 a17435a <=( A169  and  a17434a );
 a17438a <=( (not A201)  and  A166 );
 a17441a <=( A232  and  A202 );
 a17442a <=( a17441a  and  a17438a );
 a17443a <=( a17442a  and  a17435a );
 a17447a <=( A235  and  A234 );
 a17448a <=( (not A233)  and  a17447a );
 a17451a <=( A266  and  (not A265) );
 a17454a <=( A269  and  A267 );
 a17455a <=( a17454a  and  a17451a );
 a17456a <=( a17455a  and  a17448a );
 a17460a <=( (not A167)  and  A168 );
 a17461a <=( A169  and  a17460a );
 a17464a <=( (not A201)  and  A166 );
 a17467a <=( A232  and  A202 );
 a17468a <=( a17467a  and  a17464a );
 a17469a <=( a17468a  and  a17461a );
 a17473a <=( A235  and  A234 );
 a17474a <=( (not A233)  and  a17473a );
 a17477a <=( (not A266)  and  A265 );
 a17480a <=( A268  and  A267 );
 a17481a <=( a17480a  and  a17477a );
 a17482a <=( a17481a  and  a17474a );
 a17486a <=( (not A167)  and  A168 );
 a17487a <=( A169  and  a17486a );
 a17490a <=( (not A201)  and  A166 );
 a17493a <=( A232  and  A202 );
 a17494a <=( a17493a  and  a17490a );
 a17495a <=( a17494a  and  a17487a );
 a17499a <=( A235  and  A234 );
 a17500a <=( (not A233)  and  a17499a );
 a17503a <=( (not A266)  and  A265 );
 a17506a <=( A269  and  A267 );
 a17507a <=( a17506a  and  a17503a );
 a17508a <=( a17507a  and  a17500a );
 a17512a <=( (not A167)  and  A168 );
 a17513a <=( A169  and  a17512a );
 a17516a <=( (not A201)  and  A166 );
 a17519a <=( A232  and  A202 );
 a17520a <=( a17519a  and  a17516a );
 a17521a <=( a17520a  and  a17513a );
 a17525a <=( A236  and  A234 );
 a17526a <=( (not A233)  and  a17525a );
 a17529a <=( (not A299)  and  A298 );
 a17532a <=( A301  and  A300 );
 a17533a <=( a17532a  and  a17529a );
 a17534a <=( a17533a  and  a17526a );
 a17538a <=( (not A167)  and  A168 );
 a17539a <=( A169  and  a17538a );
 a17542a <=( (not A201)  and  A166 );
 a17545a <=( A232  and  A202 );
 a17546a <=( a17545a  and  a17542a );
 a17547a <=( a17546a  and  a17539a );
 a17551a <=( A236  and  A234 );
 a17552a <=( (not A233)  and  a17551a );
 a17555a <=( (not A299)  and  A298 );
 a17558a <=( A302  and  A300 );
 a17559a <=( a17558a  and  a17555a );
 a17560a <=( a17559a  and  a17552a );
 a17564a <=( (not A167)  and  A168 );
 a17565a <=( A169  and  a17564a );
 a17568a <=( (not A201)  and  A166 );
 a17571a <=( A232  and  A202 );
 a17572a <=( a17571a  and  a17568a );
 a17573a <=( a17572a  and  a17565a );
 a17577a <=( A236  and  A234 );
 a17578a <=( (not A233)  and  a17577a );
 a17581a <=( A299  and  (not A298) );
 a17584a <=( A301  and  A300 );
 a17585a <=( a17584a  and  a17581a );
 a17586a <=( a17585a  and  a17578a );
 a17590a <=( (not A167)  and  A168 );
 a17591a <=( A169  and  a17590a );
 a17594a <=( (not A201)  and  A166 );
 a17597a <=( A232  and  A202 );
 a17598a <=( a17597a  and  a17594a );
 a17599a <=( a17598a  and  a17591a );
 a17603a <=( A236  and  A234 );
 a17604a <=( (not A233)  and  a17603a );
 a17607a <=( A299  and  (not A298) );
 a17610a <=( A302  and  A300 );
 a17611a <=( a17610a  and  a17607a );
 a17612a <=( a17611a  and  a17604a );
 a17616a <=( (not A167)  and  A168 );
 a17617a <=( A169  and  a17616a );
 a17620a <=( (not A201)  and  A166 );
 a17623a <=( A232  and  A202 );
 a17624a <=( a17623a  and  a17620a );
 a17625a <=( a17624a  and  a17617a );
 a17629a <=( A236  and  A234 );
 a17630a <=( (not A233)  and  a17629a );
 a17633a <=( A266  and  (not A265) );
 a17636a <=( A268  and  A267 );
 a17637a <=( a17636a  and  a17633a );
 a17638a <=( a17637a  and  a17630a );
 a17642a <=( (not A167)  and  A168 );
 a17643a <=( A169  and  a17642a );
 a17646a <=( (not A201)  and  A166 );
 a17649a <=( A232  and  A202 );
 a17650a <=( a17649a  and  a17646a );
 a17651a <=( a17650a  and  a17643a );
 a17655a <=( A236  and  A234 );
 a17656a <=( (not A233)  and  a17655a );
 a17659a <=( A266  and  (not A265) );
 a17662a <=( A269  and  A267 );
 a17663a <=( a17662a  and  a17659a );
 a17664a <=( a17663a  and  a17656a );
 a17668a <=( (not A167)  and  A168 );
 a17669a <=( A169  and  a17668a );
 a17672a <=( (not A201)  and  A166 );
 a17675a <=( A232  and  A202 );
 a17676a <=( a17675a  and  a17672a );
 a17677a <=( a17676a  and  a17669a );
 a17681a <=( A236  and  A234 );
 a17682a <=( (not A233)  and  a17681a );
 a17685a <=( (not A266)  and  A265 );
 a17688a <=( A268  and  A267 );
 a17689a <=( a17688a  and  a17685a );
 a17690a <=( a17689a  and  a17682a );
 a17694a <=( (not A167)  and  A168 );
 a17695a <=( A169  and  a17694a );
 a17698a <=( (not A201)  and  A166 );
 a17701a <=( A232  and  A202 );
 a17702a <=( a17701a  and  a17698a );
 a17703a <=( a17702a  and  a17695a );
 a17707a <=( A236  and  A234 );
 a17708a <=( (not A233)  and  a17707a );
 a17711a <=( (not A266)  and  A265 );
 a17714a <=( A269  and  A267 );
 a17715a <=( a17714a  and  a17711a );
 a17716a <=( a17715a  and  a17708a );
 a17720a <=( (not A167)  and  A168 );
 a17721a <=( A169  and  a17720a );
 a17724a <=( (not A201)  and  A166 );
 a17727a <=( (not A232)  and  A203 );
 a17728a <=( a17727a  and  a17724a );
 a17729a <=( a17728a  and  a17721a );
 a17733a <=( A235  and  A234 );
 a17734a <=( A233  and  a17733a );
 a17737a <=( (not A299)  and  A298 );
 a17740a <=( A301  and  A300 );
 a17741a <=( a17740a  and  a17737a );
 a17742a <=( a17741a  and  a17734a );
 a17746a <=( (not A167)  and  A168 );
 a17747a <=( A169  and  a17746a );
 a17750a <=( (not A201)  and  A166 );
 a17753a <=( (not A232)  and  A203 );
 a17754a <=( a17753a  and  a17750a );
 a17755a <=( a17754a  and  a17747a );
 a17759a <=( A235  and  A234 );
 a17760a <=( A233  and  a17759a );
 a17763a <=( (not A299)  and  A298 );
 a17766a <=( A302  and  A300 );
 a17767a <=( a17766a  and  a17763a );
 a17768a <=( a17767a  and  a17760a );
 a17772a <=( (not A167)  and  A168 );
 a17773a <=( A169  and  a17772a );
 a17776a <=( (not A201)  and  A166 );
 a17779a <=( (not A232)  and  A203 );
 a17780a <=( a17779a  and  a17776a );
 a17781a <=( a17780a  and  a17773a );
 a17785a <=( A235  and  A234 );
 a17786a <=( A233  and  a17785a );
 a17789a <=( A299  and  (not A298) );
 a17792a <=( A301  and  A300 );
 a17793a <=( a17792a  and  a17789a );
 a17794a <=( a17793a  and  a17786a );
 a17798a <=( (not A167)  and  A168 );
 a17799a <=( A169  and  a17798a );
 a17802a <=( (not A201)  and  A166 );
 a17805a <=( (not A232)  and  A203 );
 a17806a <=( a17805a  and  a17802a );
 a17807a <=( a17806a  and  a17799a );
 a17811a <=( A235  and  A234 );
 a17812a <=( A233  and  a17811a );
 a17815a <=( A299  and  (not A298) );
 a17818a <=( A302  and  A300 );
 a17819a <=( a17818a  and  a17815a );
 a17820a <=( a17819a  and  a17812a );
 a17824a <=( (not A167)  and  A168 );
 a17825a <=( A169  and  a17824a );
 a17828a <=( (not A201)  and  A166 );
 a17831a <=( (not A232)  and  A203 );
 a17832a <=( a17831a  and  a17828a );
 a17833a <=( a17832a  and  a17825a );
 a17837a <=( A235  and  A234 );
 a17838a <=( A233  and  a17837a );
 a17841a <=( A266  and  (not A265) );
 a17844a <=( A268  and  A267 );
 a17845a <=( a17844a  and  a17841a );
 a17846a <=( a17845a  and  a17838a );
 a17850a <=( (not A167)  and  A168 );
 a17851a <=( A169  and  a17850a );
 a17854a <=( (not A201)  and  A166 );
 a17857a <=( (not A232)  and  A203 );
 a17858a <=( a17857a  and  a17854a );
 a17859a <=( a17858a  and  a17851a );
 a17863a <=( A235  and  A234 );
 a17864a <=( A233  and  a17863a );
 a17867a <=( A266  and  (not A265) );
 a17870a <=( A269  and  A267 );
 a17871a <=( a17870a  and  a17867a );
 a17872a <=( a17871a  and  a17864a );
 a17876a <=( (not A167)  and  A168 );
 a17877a <=( A169  and  a17876a );
 a17880a <=( (not A201)  and  A166 );
 a17883a <=( (not A232)  and  A203 );
 a17884a <=( a17883a  and  a17880a );
 a17885a <=( a17884a  and  a17877a );
 a17889a <=( A235  and  A234 );
 a17890a <=( A233  and  a17889a );
 a17893a <=( (not A266)  and  A265 );
 a17896a <=( A268  and  A267 );
 a17897a <=( a17896a  and  a17893a );
 a17898a <=( a17897a  and  a17890a );
 a17902a <=( (not A167)  and  A168 );
 a17903a <=( A169  and  a17902a );
 a17906a <=( (not A201)  and  A166 );
 a17909a <=( (not A232)  and  A203 );
 a17910a <=( a17909a  and  a17906a );
 a17911a <=( a17910a  and  a17903a );
 a17915a <=( A235  and  A234 );
 a17916a <=( A233  and  a17915a );
 a17919a <=( (not A266)  and  A265 );
 a17922a <=( A269  and  A267 );
 a17923a <=( a17922a  and  a17919a );
 a17924a <=( a17923a  and  a17916a );
 a17928a <=( (not A167)  and  A168 );
 a17929a <=( A169  and  a17928a );
 a17932a <=( (not A201)  and  A166 );
 a17935a <=( (not A232)  and  A203 );
 a17936a <=( a17935a  and  a17932a );
 a17937a <=( a17936a  and  a17929a );
 a17941a <=( A236  and  A234 );
 a17942a <=( A233  and  a17941a );
 a17945a <=( (not A299)  and  A298 );
 a17948a <=( A301  and  A300 );
 a17949a <=( a17948a  and  a17945a );
 a17950a <=( a17949a  and  a17942a );
 a17954a <=( (not A167)  and  A168 );
 a17955a <=( A169  and  a17954a );
 a17958a <=( (not A201)  and  A166 );
 a17961a <=( (not A232)  and  A203 );
 a17962a <=( a17961a  and  a17958a );
 a17963a <=( a17962a  and  a17955a );
 a17967a <=( A236  and  A234 );
 a17968a <=( A233  and  a17967a );
 a17971a <=( (not A299)  and  A298 );
 a17974a <=( A302  and  A300 );
 a17975a <=( a17974a  and  a17971a );
 a17976a <=( a17975a  and  a17968a );
 a17980a <=( (not A167)  and  A168 );
 a17981a <=( A169  and  a17980a );
 a17984a <=( (not A201)  and  A166 );
 a17987a <=( (not A232)  and  A203 );
 a17988a <=( a17987a  and  a17984a );
 a17989a <=( a17988a  and  a17981a );
 a17993a <=( A236  and  A234 );
 a17994a <=( A233  and  a17993a );
 a17997a <=( A299  and  (not A298) );
 a18000a <=( A301  and  A300 );
 a18001a <=( a18000a  and  a17997a );
 a18002a <=( a18001a  and  a17994a );
 a18006a <=( (not A167)  and  A168 );
 a18007a <=( A169  and  a18006a );
 a18010a <=( (not A201)  and  A166 );
 a18013a <=( (not A232)  and  A203 );
 a18014a <=( a18013a  and  a18010a );
 a18015a <=( a18014a  and  a18007a );
 a18019a <=( A236  and  A234 );
 a18020a <=( A233  and  a18019a );
 a18023a <=( A299  and  (not A298) );
 a18026a <=( A302  and  A300 );
 a18027a <=( a18026a  and  a18023a );
 a18028a <=( a18027a  and  a18020a );
 a18032a <=( (not A167)  and  A168 );
 a18033a <=( A169  and  a18032a );
 a18036a <=( (not A201)  and  A166 );
 a18039a <=( (not A232)  and  A203 );
 a18040a <=( a18039a  and  a18036a );
 a18041a <=( a18040a  and  a18033a );
 a18045a <=( A236  and  A234 );
 a18046a <=( A233  and  a18045a );
 a18049a <=( A266  and  (not A265) );
 a18052a <=( A268  and  A267 );
 a18053a <=( a18052a  and  a18049a );
 a18054a <=( a18053a  and  a18046a );
 a18058a <=( (not A167)  and  A168 );
 a18059a <=( A169  and  a18058a );
 a18062a <=( (not A201)  and  A166 );
 a18065a <=( (not A232)  and  A203 );
 a18066a <=( a18065a  and  a18062a );
 a18067a <=( a18066a  and  a18059a );
 a18071a <=( A236  and  A234 );
 a18072a <=( A233  and  a18071a );
 a18075a <=( A266  and  (not A265) );
 a18078a <=( A269  and  A267 );
 a18079a <=( a18078a  and  a18075a );
 a18080a <=( a18079a  and  a18072a );
 a18084a <=( (not A167)  and  A168 );
 a18085a <=( A169  and  a18084a );
 a18088a <=( (not A201)  and  A166 );
 a18091a <=( (not A232)  and  A203 );
 a18092a <=( a18091a  and  a18088a );
 a18093a <=( a18092a  and  a18085a );
 a18097a <=( A236  and  A234 );
 a18098a <=( A233  and  a18097a );
 a18101a <=( (not A266)  and  A265 );
 a18104a <=( A268  and  A267 );
 a18105a <=( a18104a  and  a18101a );
 a18106a <=( a18105a  and  a18098a );
 a18110a <=( (not A167)  and  A168 );
 a18111a <=( A169  and  a18110a );
 a18114a <=( (not A201)  and  A166 );
 a18117a <=( (not A232)  and  A203 );
 a18118a <=( a18117a  and  a18114a );
 a18119a <=( a18118a  and  a18111a );
 a18123a <=( A236  and  A234 );
 a18124a <=( A233  and  a18123a );
 a18127a <=( (not A266)  and  A265 );
 a18130a <=( A269  and  A267 );
 a18131a <=( a18130a  and  a18127a );
 a18132a <=( a18131a  and  a18124a );
 a18136a <=( (not A167)  and  A168 );
 a18137a <=( A169  and  a18136a );
 a18140a <=( (not A201)  and  A166 );
 a18143a <=( A232  and  A203 );
 a18144a <=( a18143a  and  a18140a );
 a18145a <=( a18144a  and  a18137a );
 a18149a <=( A235  and  A234 );
 a18150a <=( (not A233)  and  a18149a );
 a18153a <=( (not A299)  and  A298 );
 a18156a <=( A301  and  A300 );
 a18157a <=( a18156a  and  a18153a );
 a18158a <=( a18157a  and  a18150a );
 a18162a <=( (not A167)  and  A168 );
 a18163a <=( A169  and  a18162a );
 a18166a <=( (not A201)  and  A166 );
 a18169a <=( A232  and  A203 );
 a18170a <=( a18169a  and  a18166a );
 a18171a <=( a18170a  and  a18163a );
 a18175a <=( A235  and  A234 );
 a18176a <=( (not A233)  and  a18175a );
 a18179a <=( (not A299)  and  A298 );
 a18182a <=( A302  and  A300 );
 a18183a <=( a18182a  and  a18179a );
 a18184a <=( a18183a  and  a18176a );
 a18188a <=( (not A167)  and  A168 );
 a18189a <=( A169  and  a18188a );
 a18192a <=( (not A201)  and  A166 );
 a18195a <=( A232  and  A203 );
 a18196a <=( a18195a  and  a18192a );
 a18197a <=( a18196a  and  a18189a );
 a18201a <=( A235  and  A234 );
 a18202a <=( (not A233)  and  a18201a );
 a18205a <=( A299  and  (not A298) );
 a18208a <=( A301  and  A300 );
 a18209a <=( a18208a  and  a18205a );
 a18210a <=( a18209a  and  a18202a );
 a18214a <=( (not A167)  and  A168 );
 a18215a <=( A169  and  a18214a );
 a18218a <=( (not A201)  and  A166 );
 a18221a <=( A232  and  A203 );
 a18222a <=( a18221a  and  a18218a );
 a18223a <=( a18222a  and  a18215a );
 a18227a <=( A235  and  A234 );
 a18228a <=( (not A233)  and  a18227a );
 a18231a <=( A299  and  (not A298) );
 a18234a <=( A302  and  A300 );
 a18235a <=( a18234a  and  a18231a );
 a18236a <=( a18235a  and  a18228a );
 a18240a <=( (not A167)  and  A168 );
 a18241a <=( A169  and  a18240a );
 a18244a <=( (not A201)  and  A166 );
 a18247a <=( A232  and  A203 );
 a18248a <=( a18247a  and  a18244a );
 a18249a <=( a18248a  and  a18241a );
 a18253a <=( A235  and  A234 );
 a18254a <=( (not A233)  and  a18253a );
 a18257a <=( A266  and  (not A265) );
 a18260a <=( A268  and  A267 );
 a18261a <=( a18260a  and  a18257a );
 a18262a <=( a18261a  and  a18254a );
 a18266a <=( (not A167)  and  A168 );
 a18267a <=( A169  and  a18266a );
 a18270a <=( (not A201)  and  A166 );
 a18273a <=( A232  and  A203 );
 a18274a <=( a18273a  and  a18270a );
 a18275a <=( a18274a  and  a18267a );
 a18279a <=( A235  and  A234 );
 a18280a <=( (not A233)  and  a18279a );
 a18283a <=( A266  and  (not A265) );
 a18286a <=( A269  and  A267 );
 a18287a <=( a18286a  and  a18283a );
 a18288a <=( a18287a  and  a18280a );
 a18292a <=( (not A167)  and  A168 );
 a18293a <=( A169  and  a18292a );
 a18296a <=( (not A201)  and  A166 );
 a18299a <=( A232  and  A203 );
 a18300a <=( a18299a  and  a18296a );
 a18301a <=( a18300a  and  a18293a );
 a18305a <=( A235  and  A234 );
 a18306a <=( (not A233)  and  a18305a );
 a18309a <=( (not A266)  and  A265 );
 a18312a <=( A268  and  A267 );
 a18313a <=( a18312a  and  a18309a );
 a18314a <=( a18313a  and  a18306a );
 a18318a <=( (not A167)  and  A168 );
 a18319a <=( A169  and  a18318a );
 a18322a <=( (not A201)  and  A166 );
 a18325a <=( A232  and  A203 );
 a18326a <=( a18325a  and  a18322a );
 a18327a <=( a18326a  and  a18319a );
 a18331a <=( A235  and  A234 );
 a18332a <=( (not A233)  and  a18331a );
 a18335a <=( (not A266)  and  A265 );
 a18338a <=( A269  and  A267 );
 a18339a <=( a18338a  and  a18335a );
 a18340a <=( a18339a  and  a18332a );
 a18344a <=( (not A167)  and  A168 );
 a18345a <=( A169  and  a18344a );
 a18348a <=( (not A201)  and  A166 );
 a18351a <=( A232  and  A203 );
 a18352a <=( a18351a  and  a18348a );
 a18353a <=( a18352a  and  a18345a );
 a18357a <=( A236  and  A234 );
 a18358a <=( (not A233)  and  a18357a );
 a18361a <=( (not A299)  and  A298 );
 a18364a <=( A301  and  A300 );
 a18365a <=( a18364a  and  a18361a );
 a18366a <=( a18365a  and  a18358a );
 a18370a <=( (not A167)  and  A168 );
 a18371a <=( A169  and  a18370a );
 a18374a <=( (not A201)  and  A166 );
 a18377a <=( A232  and  A203 );
 a18378a <=( a18377a  and  a18374a );
 a18379a <=( a18378a  and  a18371a );
 a18383a <=( A236  and  A234 );
 a18384a <=( (not A233)  and  a18383a );
 a18387a <=( (not A299)  and  A298 );
 a18390a <=( A302  and  A300 );
 a18391a <=( a18390a  and  a18387a );
 a18392a <=( a18391a  and  a18384a );
 a18396a <=( (not A167)  and  A168 );
 a18397a <=( A169  and  a18396a );
 a18400a <=( (not A201)  and  A166 );
 a18403a <=( A232  and  A203 );
 a18404a <=( a18403a  and  a18400a );
 a18405a <=( a18404a  and  a18397a );
 a18409a <=( A236  and  A234 );
 a18410a <=( (not A233)  and  a18409a );
 a18413a <=( A299  and  (not A298) );
 a18416a <=( A301  and  A300 );
 a18417a <=( a18416a  and  a18413a );
 a18418a <=( a18417a  and  a18410a );
 a18422a <=( (not A167)  and  A168 );
 a18423a <=( A169  and  a18422a );
 a18426a <=( (not A201)  and  A166 );
 a18429a <=( A232  and  A203 );
 a18430a <=( a18429a  and  a18426a );
 a18431a <=( a18430a  and  a18423a );
 a18435a <=( A236  and  A234 );
 a18436a <=( (not A233)  and  a18435a );
 a18439a <=( A299  and  (not A298) );
 a18442a <=( A302  and  A300 );
 a18443a <=( a18442a  and  a18439a );
 a18444a <=( a18443a  and  a18436a );
 a18448a <=( (not A167)  and  A168 );
 a18449a <=( A169  and  a18448a );
 a18452a <=( (not A201)  and  A166 );
 a18455a <=( A232  and  A203 );
 a18456a <=( a18455a  and  a18452a );
 a18457a <=( a18456a  and  a18449a );
 a18461a <=( A236  and  A234 );
 a18462a <=( (not A233)  and  a18461a );
 a18465a <=( A266  and  (not A265) );
 a18468a <=( A268  and  A267 );
 a18469a <=( a18468a  and  a18465a );
 a18470a <=( a18469a  and  a18462a );
 a18474a <=( (not A167)  and  A168 );
 a18475a <=( A169  and  a18474a );
 a18478a <=( (not A201)  and  A166 );
 a18481a <=( A232  and  A203 );
 a18482a <=( a18481a  and  a18478a );
 a18483a <=( a18482a  and  a18475a );
 a18487a <=( A236  and  A234 );
 a18488a <=( (not A233)  and  a18487a );
 a18491a <=( A266  and  (not A265) );
 a18494a <=( A269  and  A267 );
 a18495a <=( a18494a  and  a18491a );
 a18496a <=( a18495a  and  a18488a );
 a18500a <=( (not A167)  and  A168 );
 a18501a <=( A169  and  a18500a );
 a18504a <=( (not A201)  and  A166 );
 a18507a <=( A232  and  A203 );
 a18508a <=( a18507a  and  a18504a );
 a18509a <=( a18508a  and  a18501a );
 a18513a <=( A236  and  A234 );
 a18514a <=( (not A233)  and  a18513a );
 a18517a <=( (not A266)  and  A265 );
 a18520a <=( A268  and  A267 );
 a18521a <=( a18520a  and  a18517a );
 a18522a <=( a18521a  and  a18514a );
 a18526a <=( (not A167)  and  A168 );
 a18527a <=( A169  and  a18526a );
 a18530a <=( (not A201)  and  A166 );
 a18533a <=( A232  and  A203 );
 a18534a <=( a18533a  and  a18530a );
 a18535a <=( a18534a  and  a18527a );
 a18539a <=( A236  and  A234 );
 a18540a <=( (not A233)  and  a18539a );
 a18543a <=( (not A266)  and  A265 );
 a18546a <=( A269  and  A267 );
 a18547a <=( a18546a  and  a18543a );
 a18548a <=( a18547a  and  a18540a );
 a18552a <=( (not A167)  and  A168 );
 a18553a <=( A169  and  a18552a );
 a18556a <=( A199  and  A166 );
 a18559a <=( (not A232)  and  A200 );
 a18560a <=( a18559a  and  a18556a );
 a18561a <=( a18560a  and  a18553a );
 a18565a <=( A235  and  A234 );
 a18566a <=( A233  and  a18565a );
 a18569a <=( (not A299)  and  A298 );
 a18572a <=( A301  and  A300 );
 a18573a <=( a18572a  and  a18569a );
 a18574a <=( a18573a  and  a18566a );
 a18578a <=( (not A167)  and  A168 );
 a18579a <=( A169  and  a18578a );
 a18582a <=( A199  and  A166 );
 a18585a <=( (not A232)  and  A200 );
 a18586a <=( a18585a  and  a18582a );
 a18587a <=( a18586a  and  a18579a );
 a18591a <=( A235  and  A234 );
 a18592a <=( A233  and  a18591a );
 a18595a <=( (not A299)  and  A298 );
 a18598a <=( A302  and  A300 );
 a18599a <=( a18598a  and  a18595a );
 a18600a <=( a18599a  and  a18592a );
 a18604a <=( (not A167)  and  A168 );
 a18605a <=( A169  and  a18604a );
 a18608a <=( A199  and  A166 );
 a18611a <=( (not A232)  and  A200 );
 a18612a <=( a18611a  and  a18608a );
 a18613a <=( a18612a  and  a18605a );
 a18617a <=( A235  and  A234 );
 a18618a <=( A233  and  a18617a );
 a18621a <=( A299  and  (not A298) );
 a18624a <=( A301  and  A300 );
 a18625a <=( a18624a  and  a18621a );
 a18626a <=( a18625a  and  a18618a );
 a18630a <=( (not A167)  and  A168 );
 a18631a <=( A169  and  a18630a );
 a18634a <=( A199  and  A166 );
 a18637a <=( (not A232)  and  A200 );
 a18638a <=( a18637a  and  a18634a );
 a18639a <=( a18638a  and  a18631a );
 a18643a <=( A235  and  A234 );
 a18644a <=( A233  and  a18643a );
 a18647a <=( A299  and  (not A298) );
 a18650a <=( A302  and  A300 );
 a18651a <=( a18650a  and  a18647a );
 a18652a <=( a18651a  and  a18644a );
 a18656a <=( (not A167)  and  A168 );
 a18657a <=( A169  and  a18656a );
 a18660a <=( A199  and  A166 );
 a18663a <=( (not A232)  and  A200 );
 a18664a <=( a18663a  and  a18660a );
 a18665a <=( a18664a  and  a18657a );
 a18669a <=( A235  and  A234 );
 a18670a <=( A233  and  a18669a );
 a18673a <=( A266  and  (not A265) );
 a18676a <=( A268  and  A267 );
 a18677a <=( a18676a  and  a18673a );
 a18678a <=( a18677a  and  a18670a );
 a18682a <=( (not A167)  and  A168 );
 a18683a <=( A169  and  a18682a );
 a18686a <=( A199  and  A166 );
 a18689a <=( (not A232)  and  A200 );
 a18690a <=( a18689a  and  a18686a );
 a18691a <=( a18690a  and  a18683a );
 a18695a <=( A235  and  A234 );
 a18696a <=( A233  and  a18695a );
 a18699a <=( A266  and  (not A265) );
 a18702a <=( A269  and  A267 );
 a18703a <=( a18702a  and  a18699a );
 a18704a <=( a18703a  and  a18696a );
 a18708a <=( (not A167)  and  A168 );
 a18709a <=( A169  and  a18708a );
 a18712a <=( A199  and  A166 );
 a18715a <=( (not A232)  and  A200 );
 a18716a <=( a18715a  and  a18712a );
 a18717a <=( a18716a  and  a18709a );
 a18721a <=( A235  and  A234 );
 a18722a <=( A233  and  a18721a );
 a18725a <=( (not A266)  and  A265 );
 a18728a <=( A268  and  A267 );
 a18729a <=( a18728a  and  a18725a );
 a18730a <=( a18729a  and  a18722a );
 a18734a <=( (not A167)  and  A168 );
 a18735a <=( A169  and  a18734a );
 a18738a <=( A199  and  A166 );
 a18741a <=( (not A232)  and  A200 );
 a18742a <=( a18741a  and  a18738a );
 a18743a <=( a18742a  and  a18735a );
 a18747a <=( A235  and  A234 );
 a18748a <=( A233  and  a18747a );
 a18751a <=( (not A266)  and  A265 );
 a18754a <=( A269  and  A267 );
 a18755a <=( a18754a  and  a18751a );
 a18756a <=( a18755a  and  a18748a );
 a18760a <=( (not A167)  and  A168 );
 a18761a <=( A169  and  a18760a );
 a18764a <=( A199  and  A166 );
 a18767a <=( (not A232)  and  A200 );
 a18768a <=( a18767a  and  a18764a );
 a18769a <=( a18768a  and  a18761a );
 a18773a <=( A236  and  A234 );
 a18774a <=( A233  and  a18773a );
 a18777a <=( (not A299)  and  A298 );
 a18780a <=( A301  and  A300 );
 a18781a <=( a18780a  and  a18777a );
 a18782a <=( a18781a  and  a18774a );
 a18786a <=( (not A167)  and  A168 );
 a18787a <=( A169  and  a18786a );
 a18790a <=( A199  and  A166 );
 a18793a <=( (not A232)  and  A200 );
 a18794a <=( a18793a  and  a18790a );
 a18795a <=( a18794a  and  a18787a );
 a18799a <=( A236  and  A234 );
 a18800a <=( A233  and  a18799a );
 a18803a <=( (not A299)  and  A298 );
 a18806a <=( A302  and  A300 );
 a18807a <=( a18806a  and  a18803a );
 a18808a <=( a18807a  and  a18800a );
 a18812a <=( (not A167)  and  A168 );
 a18813a <=( A169  and  a18812a );
 a18816a <=( A199  and  A166 );
 a18819a <=( (not A232)  and  A200 );
 a18820a <=( a18819a  and  a18816a );
 a18821a <=( a18820a  and  a18813a );
 a18825a <=( A236  and  A234 );
 a18826a <=( A233  and  a18825a );
 a18829a <=( A299  and  (not A298) );
 a18832a <=( A301  and  A300 );
 a18833a <=( a18832a  and  a18829a );
 a18834a <=( a18833a  and  a18826a );
 a18838a <=( (not A167)  and  A168 );
 a18839a <=( A169  and  a18838a );
 a18842a <=( A199  and  A166 );
 a18845a <=( (not A232)  and  A200 );
 a18846a <=( a18845a  and  a18842a );
 a18847a <=( a18846a  and  a18839a );
 a18851a <=( A236  and  A234 );
 a18852a <=( A233  and  a18851a );
 a18855a <=( A299  and  (not A298) );
 a18858a <=( A302  and  A300 );
 a18859a <=( a18858a  and  a18855a );
 a18860a <=( a18859a  and  a18852a );
 a18864a <=( (not A167)  and  A168 );
 a18865a <=( A169  and  a18864a );
 a18868a <=( A199  and  A166 );
 a18871a <=( (not A232)  and  A200 );
 a18872a <=( a18871a  and  a18868a );
 a18873a <=( a18872a  and  a18865a );
 a18877a <=( A236  and  A234 );
 a18878a <=( A233  and  a18877a );
 a18881a <=( A266  and  (not A265) );
 a18884a <=( A268  and  A267 );
 a18885a <=( a18884a  and  a18881a );
 a18886a <=( a18885a  and  a18878a );
 a18890a <=( (not A167)  and  A168 );
 a18891a <=( A169  and  a18890a );
 a18894a <=( A199  and  A166 );
 a18897a <=( (not A232)  and  A200 );
 a18898a <=( a18897a  and  a18894a );
 a18899a <=( a18898a  and  a18891a );
 a18903a <=( A236  and  A234 );
 a18904a <=( A233  and  a18903a );
 a18907a <=( A266  and  (not A265) );
 a18910a <=( A269  and  A267 );
 a18911a <=( a18910a  and  a18907a );
 a18912a <=( a18911a  and  a18904a );
 a18916a <=( (not A167)  and  A168 );
 a18917a <=( A169  and  a18916a );
 a18920a <=( A199  and  A166 );
 a18923a <=( (not A232)  and  A200 );
 a18924a <=( a18923a  and  a18920a );
 a18925a <=( a18924a  and  a18917a );
 a18929a <=( A236  and  A234 );
 a18930a <=( A233  and  a18929a );
 a18933a <=( (not A266)  and  A265 );
 a18936a <=( A268  and  A267 );
 a18937a <=( a18936a  and  a18933a );
 a18938a <=( a18937a  and  a18930a );
 a18942a <=( (not A167)  and  A168 );
 a18943a <=( A169  and  a18942a );
 a18946a <=( A199  and  A166 );
 a18949a <=( (not A232)  and  A200 );
 a18950a <=( a18949a  and  a18946a );
 a18951a <=( a18950a  and  a18943a );
 a18955a <=( A236  and  A234 );
 a18956a <=( A233  and  a18955a );
 a18959a <=( (not A266)  and  A265 );
 a18962a <=( A269  and  A267 );
 a18963a <=( a18962a  and  a18959a );
 a18964a <=( a18963a  and  a18956a );
 a18968a <=( (not A167)  and  A168 );
 a18969a <=( A169  and  a18968a );
 a18972a <=( A199  and  A166 );
 a18975a <=( A232  and  A200 );
 a18976a <=( a18975a  and  a18972a );
 a18977a <=( a18976a  and  a18969a );
 a18981a <=( A235  and  A234 );
 a18982a <=( (not A233)  and  a18981a );
 a18985a <=( (not A299)  and  A298 );
 a18988a <=( A301  and  A300 );
 a18989a <=( a18988a  and  a18985a );
 a18990a <=( a18989a  and  a18982a );
 a18994a <=( (not A167)  and  A168 );
 a18995a <=( A169  and  a18994a );
 a18998a <=( A199  and  A166 );
 a19001a <=( A232  and  A200 );
 a19002a <=( a19001a  and  a18998a );
 a19003a <=( a19002a  and  a18995a );
 a19007a <=( A235  and  A234 );
 a19008a <=( (not A233)  and  a19007a );
 a19011a <=( (not A299)  and  A298 );
 a19014a <=( A302  and  A300 );
 a19015a <=( a19014a  and  a19011a );
 a19016a <=( a19015a  and  a19008a );
 a19020a <=( (not A167)  and  A168 );
 a19021a <=( A169  and  a19020a );
 a19024a <=( A199  and  A166 );
 a19027a <=( A232  and  A200 );
 a19028a <=( a19027a  and  a19024a );
 a19029a <=( a19028a  and  a19021a );
 a19033a <=( A235  and  A234 );
 a19034a <=( (not A233)  and  a19033a );
 a19037a <=( A299  and  (not A298) );
 a19040a <=( A301  and  A300 );
 a19041a <=( a19040a  and  a19037a );
 a19042a <=( a19041a  and  a19034a );
 a19046a <=( (not A167)  and  A168 );
 a19047a <=( A169  and  a19046a );
 a19050a <=( A199  and  A166 );
 a19053a <=( A232  and  A200 );
 a19054a <=( a19053a  and  a19050a );
 a19055a <=( a19054a  and  a19047a );
 a19059a <=( A235  and  A234 );
 a19060a <=( (not A233)  and  a19059a );
 a19063a <=( A299  and  (not A298) );
 a19066a <=( A302  and  A300 );
 a19067a <=( a19066a  and  a19063a );
 a19068a <=( a19067a  and  a19060a );
 a19072a <=( (not A167)  and  A168 );
 a19073a <=( A169  and  a19072a );
 a19076a <=( A199  and  A166 );
 a19079a <=( A232  and  A200 );
 a19080a <=( a19079a  and  a19076a );
 a19081a <=( a19080a  and  a19073a );
 a19085a <=( A235  and  A234 );
 a19086a <=( (not A233)  and  a19085a );
 a19089a <=( A266  and  (not A265) );
 a19092a <=( A268  and  A267 );
 a19093a <=( a19092a  and  a19089a );
 a19094a <=( a19093a  and  a19086a );
 a19098a <=( (not A167)  and  A168 );
 a19099a <=( A169  and  a19098a );
 a19102a <=( A199  and  A166 );
 a19105a <=( A232  and  A200 );
 a19106a <=( a19105a  and  a19102a );
 a19107a <=( a19106a  and  a19099a );
 a19111a <=( A235  and  A234 );
 a19112a <=( (not A233)  and  a19111a );
 a19115a <=( A266  and  (not A265) );
 a19118a <=( A269  and  A267 );
 a19119a <=( a19118a  and  a19115a );
 a19120a <=( a19119a  and  a19112a );
 a19124a <=( (not A167)  and  A168 );
 a19125a <=( A169  and  a19124a );
 a19128a <=( A199  and  A166 );
 a19131a <=( A232  and  A200 );
 a19132a <=( a19131a  and  a19128a );
 a19133a <=( a19132a  and  a19125a );
 a19137a <=( A235  and  A234 );
 a19138a <=( (not A233)  and  a19137a );
 a19141a <=( (not A266)  and  A265 );
 a19144a <=( A268  and  A267 );
 a19145a <=( a19144a  and  a19141a );
 a19146a <=( a19145a  and  a19138a );
 a19150a <=( (not A167)  and  A168 );
 a19151a <=( A169  and  a19150a );
 a19154a <=( A199  and  A166 );
 a19157a <=( A232  and  A200 );
 a19158a <=( a19157a  and  a19154a );
 a19159a <=( a19158a  and  a19151a );
 a19163a <=( A235  and  A234 );
 a19164a <=( (not A233)  and  a19163a );
 a19167a <=( (not A266)  and  A265 );
 a19170a <=( A269  and  A267 );
 a19171a <=( a19170a  and  a19167a );
 a19172a <=( a19171a  and  a19164a );
 a19176a <=( (not A167)  and  A168 );
 a19177a <=( A169  and  a19176a );
 a19180a <=( A199  and  A166 );
 a19183a <=( A232  and  A200 );
 a19184a <=( a19183a  and  a19180a );
 a19185a <=( a19184a  and  a19177a );
 a19189a <=( A236  and  A234 );
 a19190a <=( (not A233)  and  a19189a );
 a19193a <=( (not A299)  and  A298 );
 a19196a <=( A301  and  A300 );
 a19197a <=( a19196a  and  a19193a );
 a19198a <=( a19197a  and  a19190a );
 a19202a <=( (not A167)  and  A168 );
 a19203a <=( A169  and  a19202a );
 a19206a <=( A199  and  A166 );
 a19209a <=( A232  and  A200 );
 a19210a <=( a19209a  and  a19206a );
 a19211a <=( a19210a  and  a19203a );
 a19215a <=( A236  and  A234 );
 a19216a <=( (not A233)  and  a19215a );
 a19219a <=( (not A299)  and  A298 );
 a19222a <=( A302  and  A300 );
 a19223a <=( a19222a  and  a19219a );
 a19224a <=( a19223a  and  a19216a );
 a19228a <=( (not A167)  and  A168 );
 a19229a <=( A169  and  a19228a );
 a19232a <=( A199  and  A166 );
 a19235a <=( A232  and  A200 );
 a19236a <=( a19235a  and  a19232a );
 a19237a <=( a19236a  and  a19229a );
 a19241a <=( A236  and  A234 );
 a19242a <=( (not A233)  and  a19241a );
 a19245a <=( A299  and  (not A298) );
 a19248a <=( A301  and  A300 );
 a19249a <=( a19248a  and  a19245a );
 a19250a <=( a19249a  and  a19242a );
 a19254a <=( (not A167)  and  A168 );
 a19255a <=( A169  and  a19254a );
 a19258a <=( A199  and  A166 );
 a19261a <=( A232  and  A200 );
 a19262a <=( a19261a  and  a19258a );
 a19263a <=( a19262a  and  a19255a );
 a19267a <=( A236  and  A234 );
 a19268a <=( (not A233)  and  a19267a );
 a19271a <=( A299  and  (not A298) );
 a19274a <=( A302  and  A300 );
 a19275a <=( a19274a  and  a19271a );
 a19276a <=( a19275a  and  a19268a );
 a19280a <=( (not A167)  and  A168 );
 a19281a <=( A169  and  a19280a );
 a19284a <=( A199  and  A166 );
 a19287a <=( A232  and  A200 );
 a19288a <=( a19287a  and  a19284a );
 a19289a <=( a19288a  and  a19281a );
 a19293a <=( A236  and  A234 );
 a19294a <=( (not A233)  and  a19293a );
 a19297a <=( A266  and  (not A265) );
 a19300a <=( A268  and  A267 );
 a19301a <=( a19300a  and  a19297a );
 a19302a <=( a19301a  and  a19294a );
 a19306a <=( (not A167)  and  A168 );
 a19307a <=( A169  and  a19306a );
 a19310a <=( A199  and  A166 );
 a19313a <=( A232  and  A200 );
 a19314a <=( a19313a  and  a19310a );
 a19315a <=( a19314a  and  a19307a );
 a19319a <=( A236  and  A234 );
 a19320a <=( (not A233)  and  a19319a );
 a19323a <=( A266  and  (not A265) );
 a19326a <=( A269  and  A267 );
 a19327a <=( a19326a  and  a19323a );
 a19328a <=( a19327a  and  a19320a );
 a19332a <=( (not A167)  and  A168 );
 a19333a <=( A169  and  a19332a );
 a19336a <=( A199  and  A166 );
 a19339a <=( A232  and  A200 );
 a19340a <=( a19339a  and  a19336a );
 a19341a <=( a19340a  and  a19333a );
 a19345a <=( A236  and  A234 );
 a19346a <=( (not A233)  and  a19345a );
 a19349a <=( (not A266)  and  A265 );
 a19352a <=( A268  and  A267 );
 a19353a <=( a19352a  and  a19349a );
 a19354a <=( a19353a  and  a19346a );
 a19358a <=( (not A167)  and  A168 );
 a19359a <=( A169  and  a19358a );
 a19362a <=( A199  and  A166 );
 a19365a <=( A232  and  A200 );
 a19366a <=( a19365a  and  a19362a );
 a19367a <=( a19366a  and  a19359a );
 a19371a <=( A236  and  A234 );
 a19372a <=( (not A233)  and  a19371a );
 a19375a <=( (not A266)  and  A265 );
 a19378a <=( A269  and  A267 );
 a19379a <=( a19378a  and  a19375a );
 a19380a <=( a19379a  and  a19372a );
 a19384a <=( (not A167)  and  A168 );
 a19385a <=( A169  and  a19384a );
 a19388a <=( (not A199)  and  A166 );
 a19391a <=( (not A232)  and  (not A200) );
 a19392a <=( a19391a  and  a19388a );
 a19393a <=( a19392a  and  a19385a );
 a19397a <=( A235  and  A234 );
 a19398a <=( A233  and  a19397a );
 a19401a <=( (not A299)  and  A298 );
 a19404a <=( A301  and  A300 );
 a19405a <=( a19404a  and  a19401a );
 a19406a <=( a19405a  and  a19398a );
 a19410a <=( (not A167)  and  A168 );
 a19411a <=( A169  and  a19410a );
 a19414a <=( (not A199)  and  A166 );
 a19417a <=( (not A232)  and  (not A200) );
 a19418a <=( a19417a  and  a19414a );
 a19419a <=( a19418a  and  a19411a );
 a19423a <=( A235  and  A234 );
 a19424a <=( A233  and  a19423a );
 a19427a <=( (not A299)  and  A298 );
 a19430a <=( A302  and  A300 );
 a19431a <=( a19430a  and  a19427a );
 a19432a <=( a19431a  and  a19424a );
 a19436a <=( (not A167)  and  A168 );
 a19437a <=( A169  and  a19436a );
 a19440a <=( (not A199)  and  A166 );
 a19443a <=( (not A232)  and  (not A200) );
 a19444a <=( a19443a  and  a19440a );
 a19445a <=( a19444a  and  a19437a );
 a19449a <=( A235  and  A234 );
 a19450a <=( A233  and  a19449a );
 a19453a <=( A299  and  (not A298) );
 a19456a <=( A301  and  A300 );
 a19457a <=( a19456a  and  a19453a );
 a19458a <=( a19457a  and  a19450a );
 a19462a <=( (not A167)  and  A168 );
 a19463a <=( A169  and  a19462a );
 a19466a <=( (not A199)  and  A166 );
 a19469a <=( (not A232)  and  (not A200) );
 a19470a <=( a19469a  and  a19466a );
 a19471a <=( a19470a  and  a19463a );
 a19475a <=( A235  and  A234 );
 a19476a <=( A233  and  a19475a );
 a19479a <=( A299  and  (not A298) );
 a19482a <=( A302  and  A300 );
 a19483a <=( a19482a  and  a19479a );
 a19484a <=( a19483a  and  a19476a );
 a19488a <=( (not A167)  and  A168 );
 a19489a <=( A169  and  a19488a );
 a19492a <=( (not A199)  and  A166 );
 a19495a <=( (not A232)  and  (not A200) );
 a19496a <=( a19495a  and  a19492a );
 a19497a <=( a19496a  and  a19489a );
 a19501a <=( A235  and  A234 );
 a19502a <=( A233  and  a19501a );
 a19505a <=( A266  and  (not A265) );
 a19508a <=( A268  and  A267 );
 a19509a <=( a19508a  and  a19505a );
 a19510a <=( a19509a  and  a19502a );
 a19514a <=( (not A167)  and  A168 );
 a19515a <=( A169  and  a19514a );
 a19518a <=( (not A199)  and  A166 );
 a19521a <=( (not A232)  and  (not A200) );
 a19522a <=( a19521a  and  a19518a );
 a19523a <=( a19522a  and  a19515a );
 a19527a <=( A235  and  A234 );
 a19528a <=( A233  and  a19527a );
 a19531a <=( A266  and  (not A265) );
 a19534a <=( A269  and  A267 );
 a19535a <=( a19534a  and  a19531a );
 a19536a <=( a19535a  and  a19528a );
 a19540a <=( (not A167)  and  A168 );
 a19541a <=( A169  and  a19540a );
 a19544a <=( (not A199)  and  A166 );
 a19547a <=( (not A232)  and  (not A200) );
 a19548a <=( a19547a  and  a19544a );
 a19549a <=( a19548a  and  a19541a );
 a19553a <=( A235  and  A234 );
 a19554a <=( A233  and  a19553a );
 a19557a <=( (not A266)  and  A265 );
 a19560a <=( A268  and  A267 );
 a19561a <=( a19560a  and  a19557a );
 a19562a <=( a19561a  and  a19554a );
 a19566a <=( (not A167)  and  A168 );
 a19567a <=( A169  and  a19566a );
 a19570a <=( (not A199)  and  A166 );
 a19573a <=( (not A232)  and  (not A200) );
 a19574a <=( a19573a  and  a19570a );
 a19575a <=( a19574a  and  a19567a );
 a19579a <=( A235  and  A234 );
 a19580a <=( A233  and  a19579a );
 a19583a <=( (not A266)  and  A265 );
 a19586a <=( A269  and  A267 );
 a19587a <=( a19586a  and  a19583a );
 a19588a <=( a19587a  and  a19580a );
 a19592a <=( (not A167)  and  A168 );
 a19593a <=( A169  and  a19592a );
 a19596a <=( (not A199)  and  A166 );
 a19599a <=( (not A232)  and  (not A200) );
 a19600a <=( a19599a  and  a19596a );
 a19601a <=( a19600a  and  a19593a );
 a19605a <=( A236  and  A234 );
 a19606a <=( A233  and  a19605a );
 a19609a <=( (not A299)  and  A298 );
 a19612a <=( A301  and  A300 );
 a19613a <=( a19612a  and  a19609a );
 a19614a <=( a19613a  and  a19606a );
 a19618a <=( (not A167)  and  A168 );
 a19619a <=( A169  and  a19618a );
 a19622a <=( (not A199)  and  A166 );
 a19625a <=( (not A232)  and  (not A200) );
 a19626a <=( a19625a  and  a19622a );
 a19627a <=( a19626a  and  a19619a );
 a19631a <=( A236  and  A234 );
 a19632a <=( A233  and  a19631a );
 a19635a <=( (not A299)  and  A298 );
 a19638a <=( A302  and  A300 );
 a19639a <=( a19638a  and  a19635a );
 a19640a <=( a19639a  and  a19632a );
 a19644a <=( (not A167)  and  A168 );
 a19645a <=( A169  and  a19644a );
 a19648a <=( (not A199)  and  A166 );
 a19651a <=( (not A232)  and  (not A200) );
 a19652a <=( a19651a  and  a19648a );
 a19653a <=( a19652a  and  a19645a );
 a19657a <=( A236  and  A234 );
 a19658a <=( A233  and  a19657a );
 a19661a <=( A299  and  (not A298) );
 a19664a <=( A301  and  A300 );
 a19665a <=( a19664a  and  a19661a );
 a19666a <=( a19665a  and  a19658a );
 a19670a <=( (not A167)  and  A168 );
 a19671a <=( A169  and  a19670a );
 a19674a <=( (not A199)  and  A166 );
 a19677a <=( (not A232)  and  (not A200) );
 a19678a <=( a19677a  and  a19674a );
 a19679a <=( a19678a  and  a19671a );
 a19683a <=( A236  and  A234 );
 a19684a <=( A233  and  a19683a );
 a19687a <=( A299  and  (not A298) );
 a19690a <=( A302  and  A300 );
 a19691a <=( a19690a  and  a19687a );
 a19692a <=( a19691a  and  a19684a );
 a19696a <=( (not A167)  and  A168 );
 a19697a <=( A169  and  a19696a );
 a19700a <=( (not A199)  and  A166 );
 a19703a <=( (not A232)  and  (not A200) );
 a19704a <=( a19703a  and  a19700a );
 a19705a <=( a19704a  and  a19697a );
 a19709a <=( A236  and  A234 );
 a19710a <=( A233  and  a19709a );
 a19713a <=( A266  and  (not A265) );
 a19716a <=( A268  and  A267 );
 a19717a <=( a19716a  and  a19713a );
 a19718a <=( a19717a  and  a19710a );
 a19722a <=( (not A167)  and  A168 );
 a19723a <=( A169  and  a19722a );
 a19726a <=( (not A199)  and  A166 );
 a19729a <=( (not A232)  and  (not A200) );
 a19730a <=( a19729a  and  a19726a );
 a19731a <=( a19730a  and  a19723a );
 a19735a <=( A236  and  A234 );
 a19736a <=( A233  and  a19735a );
 a19739a <=( A266  and  (not A265) );
 a19742a <=( A269  and  A267 );
 a19743a <=( a19742a  and  a19739a );
 a19744a <=( a19743a  and  a19736a );
 a19748a <=( (not A167)  and  A168 );
 a19749a <=( A169  and  a19748a );
 a19752a <=( (not A199)  and  A166 );
 a19755a <=( (not A232)  and  (not A200) );
 a19756a <=( a19755a  and  a19752a );
 a19757a <=( a19756a  and  a19749a );
 a19761a <=( A236  and  A234 );
 a19762a <=( A233  and  a19761a );
 a19765a <=( (not A266)  and  A265 );
 a19768a <=( A268  and  A267 );
 a19769a <=( a19768a  and  a19765a );
 a19770a <=( a19769a  and  a19762a );
 a19774a <=( (not A167)  and  A168 );
 a19775a <=( A169  and  a19774a );
 a19778a <=( (not A199)  and  A166 );
 a19781a <=( (not A232)  and  (not A200) );
 a19782a <=( a19781a  and  a19778a );
 a19783a <=( a19782a  and  a19775a );
 a19787a <=( A236  and  A234 );
 a19788a <=( A233  and  a19787a );
 a19791a <=( (not A266)  and  A265 );
 a19794a <=( A269  and  A267 );
 a19795a <=( a19794a  and  a19791a );
 a19796a <=( a19795a  and  a19788a );
 a19800a <=( (not A167)  and  A168 );
 a19801a <=( A169  and  a19800a );
 a19804a <=( (not A199)  and  A166 );
 a19807a <=( A232  and  (not A200) );
 a19808a <=( a19807a  and  a19804a );
 a19809a <=( a19808a  and  a19801a );
 a19813a <=( A235  and  A234 );
 a19814a <=( (not A233)  and  a19813a );
 a19817a <=( (not A299)  and  A298 );
 a19820a <=( A301  and  A300 );
 a19821a <=( a19820a  and  a19817a );
 a19822a <=( a19821a  and  a19814a );
 a19826a <=( (not A167)  and  A168 );
 a19827a <=( A169  and  a19826a );
 a19830a <=( (not A199)  and  A166 );
 a19833a <=( A232  and  (not A200) );
 a19834a <=( a19833a  and  a19830a );
 a19835a <=( a19834a  and  a19827a );
 a19839a <=( A235  and  A234 );
 a19840a <=( (not A233)  and  a19839a );
 a19843a <=( (not A299)  and  A298 );
 a19846a <=( A302  and  A300 );
 a19847a <=( a19846a  and  a19843a );
 a19848a <=( a19847a  and  a19840a );
 a19852a <=( (not A167)  and  A168 );
 a19853a <=( A169  and  a19852a );
 a19856a <=( (not A199)  and  A166 );
 a19859a <=( A232  and  (not A200) );
 a19860a <=( a19859a  and  a19856a );
 a19861a <=( a19860a  and  a19853a );
 a19865a <=( A235  and  A234 );
 a19866a <=( (not A233)  and  a19865a );
 a19869a <=( A299  and  (not A298) );
 a19872a <=( A301  and  A300 );
 a19873a <=( a19872a  and  a19869a );
 a19874a <=( a19873a  and  a19866a );
 a19878a <=( (not A167)  and  A168 );
 a19879a <=( A169  and  a19878a );
 a19882a <=( (not A199)  and  A166 );
 a19885a <=( A232  and  (not A200) );
 a19886a <=( a19885a  and  a19882a );
 a19887a <=( a19886a  and  a19879a );
 a19891a <=( A235  and  A234 );
 a19892a <=( (not A233)  and  a19891a );
 a19895a <=( A299  and  (not A298) );
 a19898a <=( A302  and  A300 );
 a19899a <=( a19898a  and  a19895a );
 a19900a <=( a19899a  and  a19892a );
 a19904a <=( (not A167)  and  A168 );
 a19905a <=( A169  and  a19904a );
 a19908a <=( (not A199)  and  A166 );
 a19911a <=( A232  and  (not A200) );
 a19912a <=( a19911a  and  a19908a );
 a19913a <=( a19912a  and  a19905a );
 a19917a <=( A235  and  A234 );
 a19918a <=( (not A233)  and  a19917a );
 a19921a <=( A266  and  (not A265) );
 a19924a <=( A268  and  A267 );
 a19925a <=( a19924a  and  a19921a );
 a19926a <=( a19925a  and  a19918a );
 a19930a <=( (not A167)  and  A168 );
 a19931a <=( A169  and  a19930a );
 a19934a <=( (not A199)  and  A166 );
 a19937a <=( A232  and  (not A200) );
 a19938a <=( a19937a  and  a19934a );
 a19939a <=( a19938a  and  a19931a );
 a19943a <=( A235  and  A234 );
 a19944a <=( (not A233)  and  a19943a );
 a19947a <=( A266  and  (not A265) );
 a19950a <=( A269  and  A267 );
 a19951a <=( a19950a  and  a19947a );
 a19952a <=( a19951a  and  a19944a );
 a19956a <=( (not A167)  and  A168 );
 a19957a <=( A169  and  a19956a );
 a19960a <=( (not A199)  and  A166 );
 a19963a <=( A232  and  (not A200) );
 a19964a <=( a19963a  and  a19960a );
 a19965a <=( a19964a  and  a19957a );
 a19969a <=( A235  and  A234 );
 a19970a <=( (not A233)  and  a19969a );
 a19973a <=( (not A266)  and  A265 );
 a19976a <=( A268  and  A267 );
 a19977a <=( a19976a  and  a19973a );
 a19978a <=( a19977a  and  a19970a );
 a19982a <=( (not A167)  and  A168 );
 a19983a <=( A169  and  a19982a );
 a19986a <=( (not A199)  and  A166 );
 a19989a <=( A232  and  (not A200) );
 a19990a <=( a19989a  and  a19986a );
 a19991a <=( a19990a  and  a19983a );
 a19995a <=( A235  and  A234 );
 a19996a <=( (not A233)  and  a19995a );
 a19999a <=( (not A266)  and  A265 );
 a20002a <=( A269  and  A267 );
 a20003a <=( a20002a  and  a19999a );
 a20004a <=( a20003a  and  a19996a );
 a20008a <=( (not A167)  and  A168 );
 a20009a <=( A169  and  a20008a );
 a20012a <=( (not A199)  and  A166 );
 a20015a <=( A232  and  (not A200) );
 a20016a <=( a20015a  and  a20012a );
 a20017a <=( a20016a  and  a20009a );
 a20021a <=( A236  and  A234 );
 a20022a <=( (not A233)  and  a20021a );
 a20025a <=( (not A299)  and  A298 );
 a20028a <=( A301  and  A300 );
 a20029a <=( a20028a  and  a20025a );
 a20030a <=( a20029a  and  a20022a );
 a20034a <=( (not A167)  and  A168 );
 a20035a <=( A169  and  a20034a );
 a20038a <=( (not A199)  and  A166 );
 a20041a <=( A232  and  (not A200) );
 a20042a <=( a20041a  and  a20038a );
 a20043a <=( a20042a  and  a20035a );
 a20047a <=( A236  and  A234 );
 a20048a <=( (not A233)  and  a20047a );
 a20051a <=( (not A299)  and  A298 );
 a20054a <=( A302  and  A300 );
 a20055a <=( a20054a  and  a20051a );
 a20056a <=( a20055a  and  a20048a );
 a20060a <=( (not A167)  and  A168 );
 a20061a <=( A169  and  a20060a );
 a20064a <=( (not A199)  and  A166 );
 a20067a <=( A232  and  (not A200) );
 a20068a <=( a20067a  and  a20064a );
 a20069a <=( a20068a  and  a20061a );
 a20073a <=( A236  and  A234 );
 a20074a <=( (not A233)  and  a20073a );
 a20077a <=( A299  and  (not A298) );
 a20080a <=( A301  and  A300 );
 a20081a <=( a20080a  and  a20077a );
 a20082a <=( a20081a  and  a20074a );
 a20086a <=( (not A167)  and  A168 );
 a20087a <=( A169  and  a20086a );
 a20090a <=( (not A199)  and  A166 );
 a20093a <=( A232  and  (not A200) );
 a20094a <=( a20093a  and  a20090a );
 a20095a <=( a20094a  and  a20087a );
 a20099a <=( A236  and  A234 );
 a20100a <=( (not A233)  and  a20099a );
 a20103a <=( A299  and  (not A298) );
 a20106a <=( A302  and  A300 );
 a20107a <=( a20106a  and  a20103a );
 a20108a <=( a20107a  and  a20100a );
 a20112a <=( (not A167)  and  A168 );
 a20113a <=( A169  and  a20112a );
 a20116a <=( (not A199)  and  A166 );
 a20119a <=( A232  and  (not A200) );
 a20120a <=( a20119a  and  a20116a );
 a20121a <=( a20120a  and  a20113a );
 a20125a <=( A236  and  A234 );
 a20126a <=( (not A233)  and  a20125a );
 a20129a <=( A266  and  (not A265) );
 a20132a <=( A268  and  A267 );
 a20133a <=( a20132a  and  a20129a );
 a20134a <=( a20133a  and  a20126a );
 a20138a <=( (not A167)  and  A168 );
 a20139a <=( A169  and  a20138a );
 a20142a <=( (not A199)  and  A166 );
 a20145a <=( A232  and  (not A200) );
 a20146a <=( a20145a  and  a20142a );
 a20147a <=( a20146a  and  a20139a );
 a20151a <=( A236  and  A234 );
 a20152a <=( (not A233)  and  a20151a );
 a20155a <=( A266  and  (not A265) );
 a20158a <=( A269  and  A267 );
 a20159a <=( a20158a  and  a20155a );
 a20160a <=( a20159a  and  a20152a );
 a20164a <=( (not A167)  and  A168 );
 a20165a <=( A169  and  a20164a );
 a20168a <=( (not A199)  and  A166 );
 a20171a <=( A232  and  (not A200) );
 a20172a <=( a20171a  and  a20168a );
 a20173a <=( a20172a  and  a20165a );
 a20177a <=( A236  and  A234 );
 a20178a <=( (not A233)  and  a20177a );
 a20181a <=( (not A266)  and  A265 );
 a20184a <=( A268  and  A267 );
 a20185a <=( a20184a  and  a20181a );
 a20186a <=( a20185a  and  a20178a );
 a20190a <=( (not A167)  and  A168 );
 a20191a <=( A169  and  a20190a );
 a20194a <=( (not A199)  and  A166 );
 a20197a <=( A232  and  (not A200) );
 a20198a <=( a20197a  and  a20194a );
 a20199a <=( a20198a  and  a20191a );
 a20203a <=( A236  and  A234 );
 a20204a <=( (not A233)  and  a20203a );
 a20207a <=( (not A266)  and  A265 );
 a20210a <=( A269  and  A267 );
 a20211a <=( a20210a  and  a20207a );
 a20212a <=( a20211a  and  a20204a );
 a20216a <=( A167  and  A168 );
 a20217a <=( (not A170)  and  a20216a );
 a20220a <=( A201  and  (not A166) );
 a20223a <=( (not A203)  and  (not A202) );
 a20224a <=( a20223a  and  a20220a );
 a20225a <=( a20224a  and  a20217a );
 a20228a <=( A233  and  (not A232) );
 a20231a <=( A235  and  A234 );
 a20232a <=( a20231a  and  a20228a );
 a20235a <=( (not A299)  and  A298 );
 a20238a <=( A301  and  A300 );
 a20239a <=( a20238a  and  a20235a );
 a20240a <=( a20239a  and  a20232a );
 a20244a <=( A167  and  A168 );
 a20245a <=( (not A170)  and  a20244a );
 a20248a <=( A201  and  (not A166) );
 a20251a <=( (not A203)  and  (not A202) );
 a20252a <=( a20251a  and  a20248a );
 a20253a <=( a20252a  and  a20245a );
 a20256a <=( A233  and  (not A232) );
 a20259a <=( A235  and  A234 );
 a20260a <=( a20259a  and  a20256a );
 a20263a <=( (not A299)  and  A298 );
 a20266a <=( A302  and  A300 );
 a20267a <=( a20266a  and  a20263a );
 a20268a <=( a20267a  and  a20260a );
 a20272a <=( A167  and  A168 );
 a20273a <=( (not A170)  and  a20272a );
 a20276a <=( A201  and  (not A166) );
 a20279a <=( (not A203)  and  (not A202) );
 a20280a <=( a20279a  and  a20276a );
 a20281a <=( a20280a  and  a20273a );
 a20284a <=( A233  and  (not A232) );
 a20287a <=( A235  and  A234 );
 a20288a <=( a20287a  and  a20284a );
 a20291a <=( A299  and  (not A298) );
 a20294a <=( A301  and  A300 );
 a20295a <=( a20294a  and  a20291a );
 a20296a <=( a20295a  and  a20288a );
 a20300a <=( A167  and  A168 );
 a20301a <=( (not A170)  and  a20300a );
 a20304a <=( A201  and  (not A166) );
 a20307a <=( (not A203)  and  (not A202) );
 a20308a <=( a20307a  and  a20304a );
 a20309a <=( a20308a  and  a20301a );
 a20312a <=( A233  and  (not A232) );
 a20315a <=( A235  and  A234 );
 a20316a <=( a20315a  and  a20312a );
 a20319a <=( A299  and  (not A298) );
 a20322a <=( A302  and  A300 );
 a20323a <=( a20322a  and  a20319a );
 a20324a <=( a20323a  and  a20316a );
 a20328a <=( A167  and  A168 );
 a20329a <=( (not A170)  and  a20328a );
 a20332a <=( A201  and  (not A166) );
 a20335a <=( (not A203)  and  (not A202) );
 a20336a <=( a20335a  and  a20332a );
 a20337a <=( a20336a  and  a20329a );
 a20340a <=( A233  and  (not A232) );
 a20343a <=( A235  and  A234 );
 a20344a <=( a20343a  and  a20340a );
 a20347a <=( A266  and  (not A265) );
 a20350a <=( A268  and  A267 );
 a20351a <=( a20350a  and  a20347a );
 a20352a <=( a20351a  and  a20344a );
 a20356a <=( A167  and  A168 );
 a20357a <=( (not A170)  and  a20356a );
 a20360a <=( A201  and  (not A166) );
 a20363a <=( (not A203)  and  (not A202) );
 a20364a <=( a20363a  and  a20360a );
 a20365a <=( a20364a  and  a20357a );
 a20368a <=( A233  and  (not A232) );
 a20371a <=( A235  and  A234 );
 a20372a <=( a20371a  and  a20368a );
 a20375a <=( A266  and  (not A265) );
 a20378a <=( A269  and  A267 );
 a20379a <=( a20378a  and  a20375a );
 a20380a <=( a20379a  and  a20372a );
 a20384a <=( A167  and  A168 );
 a20385a <=( (not A170)  and  a20384a );
 a20388a <=( A201  and  (not A166) );
 a20391a <=( (not A203)  and  (not A202) );
 a20392a <=( a20391a  and  a20388a );
 a20393a <=( a20392a  and  a20385a );
 a20396a <=( A233  and  (not A232) );
 a20399a <=( A235  and  A234 );
 a20400a <=( a20399a  and  a20396a );
 a20403a <=( (not A266)  and  A265 );
 a20406a <=( A268  and  A267 );
 a20407a <=( a20406a  and  a20403a );
 a20408a <=( a20407a  and  a20400a );
 a20412a <=( A167  and  A168 );
 a20413a <=( (not A170)  and  a20412a );
 a20416a <=( A201  and  (not A166) );
 a20419a <=( (not A203)  and  (not A202) );
 a20420a <=( a20419a  and  a20416a );
 a20421a <=( a20420a  and  a20413a );
 a20424a <=( A233  and  (not A232) );
 a20427a <=( A235  and  A234 );
 a20428a <=( a20427a  and  a20424a );
 a20431a <=( (not A266)  and  A265 );
 a20434a <=( A269  and  A267 );
 a20435a <=( a20434a  and  a20431a );
 a20436a <=( a20435a  and  a20428a );
 a20440a <=( A167  and  A168 );
 a20441a <=( (not A170)  and  a20440a );
 a20444a <=( A201  and  (not A166) );
 a20447a <=( (not A203)  and  (not A202) );
 a20448a <=( a20447a  and  a20444a );
 a20449a <=( a20448a  and  a20441a );
 a20452a <=( A233  and  (not A232) );
 a20455a <=( A236  and  A234 );
 a20456a <=( a20455a  and  a20452a );
 a20459a <=( (not A299)  and  A298 );
 a20462a <=( A301  and  A300 );
 a20463a <=( a20462a  and  a20459a );
 a20464a <=( a20463a  and  a20456a );
 a20468a <=( A167  and  A168 );
 a20469a <=( (not A170)  and  a20468a );
 a20472a <=( A201  and  (not A166) );
 a20475a <=( (not A203)  and  (not A202) );
 a20476a <=( a20475a  and  a20472a );
 a20477a <=( a20476a  and  a20469a );
 a20480a <=( A233  and  (not A232) );
 a20483a <=( A236  and  A234 );
 a20484a <=( a20483a  and  a20480a );
 a20487a <=( (not A299)  and  A298 );
 a20490a <=( A302  and  A300 );
 a20491a <=( a20490a  and  a20487a );
 a20492a <=( a20491a  and  a20484a );
 a20496a <=( A167  and  A168 );
 a20497a <=( (not A170)  and  a20496a );
 a20500a <=( A201  and  (not A166) );
 a20503a <=( (not A203)  and  (not A202) );
 a20504a <=( a20503a  and  a20500a );
 a20505a <=( a20504a  and  a20497a );
 a20508a <=( A233  and  (not A232) );
 a20511a <=( A236  and  A234 );
 a20512a <=( a20511a  and  a20508a );
 a20515a <=( A299  and  (not A298) );
 a20518a <=( A301  and  A300 );
 a20519a <=( a20518a  and  a20515a );
 a20520a <=( a20519a  and  a20512a );
 a20524a <=( A167  and  A168 );
 a20525a <=( (not A170)  and  a20524a );
 a20528a <=( A201  and  (not A166) );
 a20531a <=( (not A203)  and  (not A202) );
 a20532a <=( a20531a  and  a20528a );
 a20533a <=( a20532a  and  a20525a );
 a20536a <=( A233  and  (not A232) );
 a20539a <=( A236  and  A234 );
 a20540a <=( a20539a  and  a20536a );
 a20543a <=( A299  and  (not A298) );
 a20546a <=( A302  and  A300 );
 a20547a <=( a20546a  and  a20543a );
 a20548a <=( a20547a  and  a20540a );
 a20552a <=( A167  and  A168 );
 a20553a <=( (not A170)  and  a20552a );
 a20556a <=( A201  and  (not A166) );
 a20559a <=( (not A203)  and  (not A202) );
 a20560a <=( a20559a  and  a20556a );
 a20561a <=( a20560a  and  a20553a );
 a20564a <=( A233  and  (not A232) );
 a20567a <=( A236  and  A234 );
 a20568a <=( a20567a  and  a20564a );
 a20571a <=( A266  and  (not A265) );
 a20574a <=( A268  and  A267 );
 a20575a <=( a20574a  and  a20571a );
 a20576a <=( a20575a  and  a20568a );
 a20580a <=( A167  and  A168 );
 a20581a <=( (not A170)  and  a20580a );
 a20584a <=( A201  and  (not A166) );
 a20587a <=( (not A203)  and  (not A202) );
 a20588a <=( a20587a  and  a20584a );
 a20589a <=( a20588a  and  a20581a );
 a20592a <=( A233  and  (not A232) );
 a20595a <=( A236  and  A234 );
 a20596a <=( a20595a  and  a20592a );
 a20599a <=( A266  and  (not A265) );
 a20602a <=( A269  and  A267 );
 a20603a <=( a20602a  and  a20599a );
 a20604a <=( a20603a  and  a20596a );
 a20608a <=( A167  and  A168 );
 a20609a <=( (not A170)  and  a20608a );
 a20612a <=( A201  and  (not A166) );
 a20615a <=( (not A203)  and  (not A202) );
 a20616a <=( a20615a  and  a20612a );
 a20617a <=( a20616a  and  a20609a );
 a20620a <=( A233  and  (not A232) );
 a20623a <=( A236  and  A234 );
 a20624a <=( a20623a  and  a20620a );
 a20627a <=( (not A266)  and  A265 );
 a20630a <=( A268  and  A267 );
 a20631a <=( a20630a  and  a20627a );
 a20632a <=( a20631a  and  a20624a );
 a20636a <=( A167  and  A168 );
 a20637a <=( (not A170)  and  a20636a );
 a20640a <=( A201  and  (not A166) );
 a20643a <=( (not A203)  and  (not A202) );
 a20644a <=( a20643a  and  a20640a );
 a20645a <=( a20644a  and  a20637a );
 a20648a <=( A233  and  (not A232) );
 a20651a <=( A236  and  A234 );
 a20652a <=( a20651a  and  a20648a );
 a20655a <=( (not A266)  and  A265 );
 a20658a <=( A269  and  A267 );
 a20659a <=( a20658a  and  a20655a );
 a20660a <=( a20659a  and  a20652a );
 a20664a <=( A167  and  A168 );
 a20665a <=( (not A170)  and  a20664a );
 a20668a <=( A201  and  (not A166) );
 a20671a <=( (not A203)  and  (not A202) );
 a20672a <=( a20671a  and  a20668a );
 a20673a <=( a20672a  and  a20665a );
 a20676a <=( (not A233)  and  A232 );
 a20679a <=( A235  and  A234 );
 a20680a <=( a20679a  and  a20676a );
 a20683a <=( (not A299)  and  A298 );
 a20686a <=( A301  and  A300 );
 a20687a <=( a20686a  and  a20683a );
 a20688a <=( a20687a  and  a20680a );
 a20692a <=( A167  and  A168 );
 a20693a <=( (not A170)  and  a20692a );
 a20696a <=( A201  and  (not A166) );
 a20699a <=( (not A203)  and  (not A202) );
 a20700a <=( a20699a  and  a20696a );
 a20701a <=( a20700a  and  a20693a );
 a20704a <=( (not A233)  and  A232 );
 a20707a <=( A235  and  A234 );
 a20708a <=( a20707a  and  a20704a );
 a20711a <=( (not A299)  and  A298 );
 a20714a <=( A302  and  A300 );
 a20715a <=( a20714a  and  a20711a );
 a20716a <=( a20715a  and  a20708a );
 a20720a <=( A167  and  A168 );
 a20721a <=( (not A170)  and  a20720a );
 a20724a <=( A201  and  (not A166) );
 a20727a <=( (not A203)  and  (not A202) );
 a20728a <=( a20727a  and  a20724a );
 a20729a <=( a20728a  and  a20721a );
 a20732a <=( (not A233)  and  A232 );
 a20735a <=( A235  and  A234 );
 a20736a <=( a20735a  and  a20732a );
 a20739a <=( A299  and  (not A298) );
 a20742a <=( A301  and  A300 );
 a20743a <=( a20742a  and  a20739a );
 a20744a <=( a20743a  and  a20736a );
 a20748a <=( A167  and  A168 );
 a20749a <=( (not A170)  and  a20748a );
 a20752a <=( A201  and  (not A166) );
 a20755a <=( (not A203)  and  (not A202) );
 a20756a <=( a20755a  and  a20752a );
 a20757a <=( a20756a  and  a20749a );
 a20760a <=( (not A233)  and  A232 );
 a20763a <=( A235  and  A234 );
 a20764a <=( a20763a  and  a20760a );
 a20767a <=( A299  and  (not A298) );
 a20770a <=( A302  and  A300 );
 a20771a <=( a20770a  and  a20767a );
 a20772a <=( a20771a  and  a20764a );
 a20776a <=( A167  and  A168 );
 a20777a <=( (not A170)  and  a20776a );
 a20780a <=( A201  and  (not A166) );
 a20783a <=( (not A203)  and  (not A202) );
 a20784a <=( a20783a  and  a20780a );
 a20785a <=( a20784a  and  a20777a );
 a20788a <=( (not A233)  and  A232 );
 a20791a <=( A235  and  A234 );
 a20792a <=( a20791a  and  a20788a );
 a20795a <=( A266  and  (not A265) );
 a20798a <=( A268  and  A267 );
 a20799a <=( a20798a  and  a20795a );
 a20800a <=( a20799a  and  a20792a );
 a20804a <=( A167  and  A168 );
 a20805a <=( (not A170)  and  a20804a );
 a20808a <=( A201  and  (not A166) );
 a20811a <=( (not A203)  and  (not A202) );
 a20812a <=( a20811a  and  a20808a );
 a20813a <=( a20812a  and  a20805a );
 a20816a <=( (not A233)  and  A232 );
 a20819a <=( A235  and  A234 );
 a20820a <=( a20819a  and  a20816a );
 a20823a <=( A266  and  (not A265) );
 a20826a <=( A269  and  A267 );
 a20827a <=( a20826a  and  a20823a );
 a20828a <=( a20827a  and  a20820a );
 a20832a <=( A167  and  A168 );
 a20833a <=( (not A170)  and  a20832a );
 a20836a <=( A201  and  (not A166) );
 a20839a <=( (not A203)  and  (not A202) );
 a20840a <=( a20839a  and  a20836a );
 a20841a <=( a20840a  and  a20833a );
 a20844a <=( (not A233)  and  A232 );
 a20847a <=( A235  and  A234 );
 a20848a <=( a20847a  and  a20844a );
 a20851a <=( (not A266)  and  A265 );
 a20854a <=( A268  and  A267 );
 a20855a <=( a20854a  and  a20851a );
 a20856a <=( a20855a  and  a20848a );
 a20860a <=( A167  and  A168 );
 a20861a <=( (not A170)  and  a20860a );
 a20864a <=( A201  and  (not A166) );
 a20867a <=( (not A203)  and  (not A202) );
 a20868a <=( a20867a  and  a20864a );
 a20869a <=( a20868a  and  a20861a );
 a20872a <=( (not A233)  and  A232 );
 a20875a <=( A235  and  A234 );
 a20876a <=( a20875a  and  a20872a );
 a20879a <=( (not A266)  and  A265 );
 a20882a <=( A269  and  A267 );
 a20883a <=( a20882a  and  a20879a );
 a20884a <=( a20883a  and  a20876a );
 a20888a <=( A167  and  A168 );
 a20889a <=( (not A170)  and  a20888a );
 a20892a <=( A201  and  (not A166) );
 a20895a <=( (not A203)  and  (not A202) );
 a20896a <=( a20895a  and  a20892a );
 a20897a <=( a20896a  and  a20889a );
 a20900a <=( (not A233)  and  A232 );
 a20903a <=( A236  and  A234 );
 a20904a <=( a20903a  and  a20900a );
 a20907a <=( (not A299)  and  A298 );
 a20910a <=( A301  and  A300 );
 a20911a <=( a20910a  and  a20907a );
 a20912a <=( a20911a  and  a20904a );
 a20916a <=( A167  and  A168 );
 a20917a <=( (not A170)  and  a20916a );
 a20920a <=( A201  and  (not A166) );
 a20923a <=( (not A203)  and  (not A202) );
 a20924a <=( a20923a  and  a20920a );
 a20925a <=( a20924a  and  a20917a );
 a20928a <=( (not A233)  and  A232 );
 a20931a <=( A236  and  A234 );
 a20932a <=( a20931a  and  a20928a );
 a20935a <=( (not A299)  and  A298 );
 a20938a <=( A302  and  A300 );
 a20939a <=( a20938a  and  a20935a );
 a20940a <=( a20939a  and  a20932a );
 a20944a <=( A167  and  A168 );
 a20945a <=( (not A170)  and  a20944a );
 a20948a <=( A201  and  (not A166) );
 a20951a <=( (not A203)  and  (not A202) );
 a20952a <=( a20951a  and  a20948a );
 a20953a <=( a20952a  and  a20945a );
 a20956a <=( (not A233)  and  A232 );
 a20959a <=( A236  and  A234 );
 a20960a <=( a20959a  and  a20956a );
 a20963a <=( A299  and  (not A298) );
 a20966a <=( A301  and  A300 );
 a20967a <=( a20966a  and  a20963a );
 a20968a <=( a20967a  and  a20960a );
 a20972a <=( A167  and  A168 );
 a20973a <=( (not A170)  and  a20972a );
 a20976a <=( A201  and  (not A166) );
 a20979a <=( (not A203)  and  (not A202) );
 a20980a <=( a20979a  and  a20976a );
 a20981a <=( a20980a  and  a20973a );
 a20984a <=( (not A233)  and  A232 );
 a20987a <=( A236  and  A234 );
 a20988a <=( a20987a  and  a20984a );
 a20991a <=( A299  and  (not A298) );
 a20994a <=( A302  and  A300 );
 a20995a <=( a20994a  and  a20991a );
 a20996a <=( a20995a  and  a20988a );
 a21000a <=( A167  and  A168 );
 a21001a <=( (not A170)  and  a21000a );
 a21004a <=( A201  and  (not A166) );
 a21007a <=( (not A203)  and  (not A202) );
 a21008a <=( a21007a  and  a21004a );
 a21009a <=( a21008a  and  a21001a );
 a21012a <=( (not A233)  and  A232 );
 a21015a <=( A236  and  A234 );
 a21016a <=( a21015a  and  a21012a );
 a21019a <=( A266  and  (not A265) );
 a21022a <=( A268  and  A267 );
 a21023a <=( a21022a  and  a21019a );
 a21024a <=( a21023a  and  a21016a );
 a21028a <=( A167  and  A168 );
 a21029a <=( (not A170)  and  a21028a );
 a21032a <=( A201  and  (not A166) );
 a21035a <=( (not A203)  and  (not A202) );
 a21036a <=( a21035a  and  a21032a );
 a21037a <=( a21036a  and  a21029a );
 a21040a <=( (not A233)  and  A232 );
 a21043a <=( A236  and  A234 );
 a21044a <=( a21043a  and  a21040a );
 a21047a <=( A266  and  (not A265) );
 a21050a <=( A269  and  A267 );
 a21051a <=( a21050a  and  a21047a );
 a21052a <=( a21051a  and  a21044a );
 a21056a <=( A167  and  A168 );
 a21057a <=( (not A170)  and  a21056a );
 a21060a <=( A201  and  (not A166) );
 a21063a <=( (not A203)  and  (not A202) );
 a21064a <=( a21063a  and  a21060a );
 a21065a <=( a21064a  and  a21057a );
 a21068a <=( (not A233)  and  A232 );
 a21071a <=( A236  and  A234 );
 a21072a <=( a21071a  and  a21068a );
 a21075a <=( (not A266)  and  A265 );
 a21078a <=( A268  and  A267 );
 a21079a <=( a21078a  and  a21075a );
 a21080a <=( a21079a  and  a21072a );
 a21084a <=( A167  and  A168 );
 a21085a <=( (not A170)  and  a21084a );
 a21088a <=( A201  and  (not A166) );
 a21091a <=( (not A203)  and  (not A202) );
 a21092a <=( a21091a  and  a21088a );
 a21093a <=( a21092a  and  a21085a );
 a21096a <=( (not A233)  and  A232 );
 a21099a <=( A236  and  A234 );
 a21100a <=( a21099a  and  a21096a );
 a21103a <=( (not A266)  and  A265 );
 a21106a <=( A269  and  A267 );
 a21107a <=( a21106a  and  a21103a );
 a21108a <=( a21107a  and  a21100a );
 a21112a <=( A167  and  A168 );
 a21113a <=( (not A170)  and  a21112a );
 a21116a <=( (not A201)  and  (not A166) );
 a21119a <=( (not A232)  and  A202 );
 a21120a <=( a21119a  and  a21116a );
 a21121a <=( a21120a  and  a21113a );
 a21124a <=( A234  and  A233 );
 a21127a <=( A298  and  A235 );
 a21128a <=( a21127a  and  a21124a );
 a21131a <=( (not A300)  and  (not A299) );
 a21134a <=( (not A302)  and  (not A301) );
 a21135a <=( a21134a  and  a21131a );
 a21136a <=( a21135a  and  a21128a );
 a21140a <=( A167  and  A168 );
 a21141a <=( (not A170)  and  a21140a );
 a21144a <=( (not A201)  and  (not A166) );
 a21147a <=( (not A232)  and  A202 );
 a21148a <=( a21147a  and  a21144a );
 a21149a <=( a21148a  and  a21141a );
 a21152a <=( A234  and  A233 );
 a21155a <=( (not A298)  and  A235 );
 a21156a <=( a21155a  and  a21152a );
 a21159a <=( (not A300)  and  A299 );
 a21162a <=( (not A302)  and  (not A301) );
 a21163a <=( a21162a  and  a21159a );
 a21164a <=( a21163a  and  a21156a );
 a21168a <=( A167  and  A168 );
 a21169a <=( (not A170)  and  a21168a );
 a21172a <=( (not A201)  and  (not A166) );
 a21175a <=( (not A232)  and  A202 );
 a21176a <=( a21175a  and  a21172a );
 a21177a <=( a21176a  and  a21169a );
 a21180a <=( A234  and  A233 );
 a21183a <=( (not A265)  and  A235 );
 a21184a <=( a21183a  and  a21180a );
 a21187a <=( (not A267)  and  A266 );
 a21190a <=( (not A269)  and  (not A268) );
 a21191a <=( a21190a  and  a21187a );
 a21192a <=( a21191a  and  a21184a );
 a21196a <=( A167  and  A168 );
 a21197a <=( (not A170)  and  a21196a );
 a21200a <=( (not A201)  and  (not A166) );
 a21203a <=( (not A232)  and  A202 );
 a21204a <=( a21203a  and  a21200a );
 a21205a <=( a21204a  and  a21197a );
 a21208a <=( A234  and  A233 );
 a21211a <=( A265  and  A235 );
 a21212a <=( a21211a  and  a21208a );
 a21215a <=( (not A267)  and  (not A266) );
 a21218a <=( (not A269)  and  (not A268) );
 a21219a <=( a21218a  and  a21215a );
 a21220a <=( a21219a  and  a21212a );
 a21224a <=( A167  and  A168 );
 a21225a <=( (not A170)  and  a21224a );
 a21228a <=( (not A201)  and  (not A166) );
 a21231a <=( (not A232)  and  A202 );
 a21232a <=( a21231a  and  a21228a );
 a21233a <=( a21232a  and  a21225a );
 a21236a <=( A234  and  A233 );
 a21239a <=( A298  and  A236 );
 a21240a <=( a21239a  and  a21236a );
 a21243a <=( (not A300)  and  (not A299) );
 a21246a <=( (not A302)  and  (not A301) );
 a21247a <=( a21246a  and  a21243a );
 a21248a <=( a21247a  and  a21240a );
 a21252a <=( A167  and  A168 );
 a21253a <=( (not A170)  and  a21252a );
 a21256a <=( (not A201)  and  (not A166) );
 a21259a <=( (not A232)  and  A202 );
 a21260a <=( a21259a  and  a21256a );
 a21261a <=( a21260a  and  a21253a );
 a21264a <=( A234  and  A233 );
 a21267a <=( (not A298)  and  A236 );
 a21268a <=( a21267a  and  a21264a );
 a21271a <=( (not A300)  and  A299 );
 a21274a <=( (not A302)  and  (not A301) );
 a21275a <=( a21274a  and  a21271a );
 a21276a <=( a21275a  and  a21268a );
 a21280a <=( A167  and  A168 );
 a21281a <=( (not A170)  and  a21280a );
 a21284a <=( (not A201)  and  (not A166) );
 a21287a <=( (not A232)  and  A202 );
 a21288a <=( a21287a  and  a21284a );
 a21289a <=( a21288a  and  a21281a );
 a21292a <=( A234  and  A233 );
 a21295a <=( (not A265)  and  A236 );
 a21296a <=( a21295a  and  a21292a );
 a21299a <=( (not A267)  and  A266 );
 a21302a <=( (not A269)  and  (not A268) );
 a21303a <=( a21302a  and  a21299a );
 a21304a <=( a21303a  and  a21296a );
 a21308a <=( A167  and  A168 );
 a21309a <=( (not A170)  and  a21308a );
 a21312a <=( (not A201)  and  (not A166) );
 a21315a <=( (not A232)  and  A202 );
 a21316a <=( a21315a  and  a21312a );
 a21317a <=( a21316a  and  a21309a );
 a21320a <=( A234  and  A233 );
 a21323a <=( A265  and  A236 );
 a21324a <=( a21323a  and  a21320a );
 a21327a <=( (not A267)  and  (not A266) );
 a21330a <=( (not A269)  and  (not A268) );
 a21331a <=( a21330a  and  a21327a );
 a21332a <=( a21331a  and  a21324a );
 a21336a <=( A167  and  A168 );
 a21337a <=( (not A170)  and  a21336a );
 a21340a <=( (not A201)  and  (not A166) );
 a21343a <=( (not A232)  and  A202 );
 a21344a <=( a21343a  and  a21340a );
 a21345a <=( a21344a  and  a21337a );
 a21348a <=( (not A234)  and  A233 );
 a21351a <=( (not A236)  and  (not A235) );
 a21352a <=( a21351a  and  a21348a );
 a21355a <=( (not A299)  and  A298 );
 a21358a <=( A301  and  A300 );
 a21359a <=( a21358a  and  a21355a );
 a21360a <=( a21359a  and  a21352a );
 a21364a <=( A167  and  A168 );
 a21365a <=( (not A170)  and  a21364a );
 a21368a <=( (not A201)  and  (not A166) );
 a21371a <=( (not A232)  and  A202 );
 a21372a <=( a21371a  and  a21368a );
 a21373a <=( a21372a  and  a21365a );
 a21376a <=( (not A234)  and  A233 );
 a21379a <=( (not A236)  and  (not A235) );
 a21380a <=( a21379a  and  a21376a );
 a21383a <=( (not A299)  and  A298 );
 a21386a <=( A302  and  A300 );
 a21387a <=( a21386a  and  a21383a );
 a21388a <=( a21387a  and  a21380a );
 a21392a <=( A167  and  A168 );
 a21393a <=( (not A170)  and  a21392a );
 a21396a <=( (not A201)  and  (not A166) );
 a21399a <=( (not A232)  and  A202 );
 a21400a <=( a21399a  and  a21396a );
 a21401a <=( a21400a  and  a21393a );
 a21404a <=( (not A234)  and  A233 );
 a21407a <=( (not A236)  and  (not A235) );
 a21408a <=( a21407a  and  a21404a );
 a21411a <=( A299  and  (not A298) );
 a21414a <=( A301  and  A300 );
 a21415a <=( a21414a  and  a21411a );
 a21416a <=( a21415a  and  a21408a );
 a21420a <=( A167  and  A168 );
 a21421a <=( (not A170)  and  a21420a );
 a21424a <=( (not A201)  and  (not A166) );
 a21427a <=( (not A232)  and  A202 );
 a21428a <=( a21427a  and  a21424a );
 a21429a <=( a21428a  and  a21421a );
 a21432a <=( (not A234)  and  A233 );
 a21435a <=( (not A236)  and  (not A235) );
 a21436a <=( a21435a  and  a21432a );
 a21439a <=( A299  and  (not A298) );
 a21442a <=( A302  and  A300 );
 a21443a <=( a21442a  and  a21439a );
 a21444a <=( a21443a  and  a21436a );
 a21448a <=( A167  and  A168 );
 a21449a <=( (not A170)  and  a21448a );
 a21452a <=( (not A201)  and  (not A166) );
 a21455a <=( (not A232)  and  A202 );
 a21456a <=( a21455a  and  a21452a );
 a21457a <=( a21456a  and  a21449a );
 a21460a <=( (not A234)  and  A233 );
 a21463a <=( (not A236)  and  (not A235) );
 a21464a <=( a21463a  and  a21460a );
 a21467a <=( A266  and  (not A265) );
 a21470a <=( A268  and  A267 );
 a21471a <=( a21470a  and  a21467a );
 a21472a <=( a21471a  and  a21464a );
 a21476a <=( A167  and  A168 );
 a21477a <=( (not A170)  and  a21476a );
 a21480a <=( (not A201)  and  (not A166) );
 a21483a <=( (not A232)  and  A202 );
 a21484a <=( a21483a  and  a21480a );
 a21485a <=( a21484a  and  a21477a );
 a21488a <=( (not A234)  and  A233 );
 a21491a <=( (not A236)  and  (not A235) );
 a21492a <=( a21491a  and  a21488a );
 a21495a <=( A266  and  (not A265) );
 a21498a <=( A269  and  A267 );
 a21499a <=( a21498a  and  a21495a );
 a21500a <=( a21499a  and  a21492a );
 a21504a <=( A167  and  A168 );
 a21505a <=( (not A170)  and  a21504a );
 a21508a <=( (not A201)  and  (not A166) );
 a21511a <=( (not A232)  and  A202 );
 a21512a <=( a21511a  and  a21508a );
 a21513a <=( a21512a  and  a21505a );
 a21516a <=( (not A234)  and  A233 );
 a21519a <=( (not A236)  and  (not A235) );
 a21520a <=( a21519a  and  a21516a );
 a21523a <=( (not A266)  and  A265 );
 a21526a <=( A268  and  A267 );
 a21527a <=( a21526a  and  a21523a );
 a21528a <=( a21527a  and  a21520a );
 a21532a <=( A167  and  A168 );
 a21533a <=( (not A170)  and  a21532a );
 a21536a <=( (not A201)  and  (not A166) );
 a21539a <=( (not A232)  and  A202 );
 a21540a <=( a21539a  and  a21536a );
 a21541a <=( a21540a  and  a21533a );
 a21544a <=( (not A234)  and  A233 );
 a21547a <=( (not A236)  and  (not A235) );
 a21548a <=( a21547a  and  a21544a );
 a21551a <=( (not A266)  and  A265 );
 a21554a <=( A269  and  A267 );
 a21555a <=( a21554a  and  a21551a );
 a21556a <=( a21555a  and  a21548a );
 a21560a <=( A167  and  A168 );
 a21561a <=( (not A170)  and  a21560a );
 a21564a <=( (not A201)  and  (not A166) );
 a21567a <=( A232  and  A202 );
 a21568a <=( a21567a  and  a21564a );
 a21569a <=( a21568a  and  a21561a );
 a21572a <=( A234  and  (not A233) );
 a21575a <=( A298  and  A235 );
 a21576a <=( a21575a  and  a21572a );
 a21579a <=( (not A300)  and  (not A299) );
 a21582a <=( (not A302)  and  (not A301) );
 a21583a <=( a21582a  and  a21579a );
 a21584a <=( a21583a  and  a21576a );
 a21588a <=( A167  and  A168 );
 a21589a <=( (not A170)  and  a21588a );
 a21592a <=( (not A201)  and  (not A166) );
 a21595a <=( A232  and  A202 );
 a21596a <=( a21595a  and  a21592a );
 a21597a <=( a21596a  and  a21589a );
 a21600a <=( A234  and  (not A233) );
 a21603a <=( (not A298)  and  A235 );
 a21604a <=( a21603a  and  a21600a );
 a21607a <=( (not A300)  and  A299 );
 a21610a <=( (not A302)  and  (not A301) );
 a21611a <=( a21610a  and  a21607a );
 a21612a <=( a21611a  and  a21604a );
 a21616a <=( A167  and  A168 );
 a21617a <=( (not A170)  and  a21616a );
 a21620a <=( (not A201)  and  (not A166) );
 a21623a <=( A232  and  A202 );
 a21624a <=( a21623a  and  a21620a );
 a21625a <=( a21624a  and  a21617a );
 a21628a <=( A234  and  (not A233) );
 a21631a <=( (not A265)  and  A235 );
 a21632a <=( a21631a  and  a21628a );
 a21635a <=( (not A267)  and  A266 );
 a21638a <=( (not A269)  and  (not A268) );
 a21639a <=( a21638a  and  a21635a );
 a21640a <=( a21639a  and  a21632a );
 a21644a <=( A167  and  A168 );
 a21645a <=( (not A170)  and  a21644a );
 a21648a <=( (not A201)  and  (not A166) );
 a21651a <=( A232  and  A202 );
 a21652a <=( a21651a  and  a21648a );
 a21653a <=( a21652a  and  a21645a );
 a21656a <=( A234  and  (not A233) );
 a21659a <=( A265  and  A235 );
 a21660a <=( a21659a  and  a21656a );
 a21663a <=( (not A267)  and  (not A266) );
 a21666a <=( (not A269)  and  (not A268) );
 a21667a <=( a21666a  and  a21663a );
 a21668a <=( a21667a  and  a21660a );
 a21672a <=( A167  and  A168 );
 a21673a <=( (not A170)  and  a21672a );
 a21676a <=( (not A201)  and  (not A166) );
 a21679a <=( A232  and  A202 );
 a21680a <=( a21679a  and  a21676a );
 a21681a <=( a21680a  and  a21673a );
 a21684a <=( A234  and  (not A233) );
 a21687a <=( A298  and  A236 );
 a21688a <=( a21687a  and  a21684a );
 a21691a <=( (not A300)  and  (not A299) );
 a21694a <=( (not A302)  and  (not A301) );
 a21695a <=( a21694a  and  a21691a );
 a21696a <=( a21695a  and  a21688a );
 a21700a <=( A167  and  A168 );
 a21701a <=( (not A170)  and  a21700a );
 a21704a <=( (not A201)  and  (not A166) );
 a21707a <=( A232  and  A202 );
 a21708a <=( a21707a  and  a21704a );
 a21709a <=( a21708a  and  a21701a );
 a21712a <=( A234  and  (not A233) );
 a21715a <=( (not A298)  and  A236 );
 a21716a <=( a21715a  and  a21712a );
 a21719a <=( (not A300)  and  A299 );
 a21722a <=( (not A302)  and  (not A301) );
 a21723a <=( a21722a  and  a21719a );
 a21724a <=( a21723a  and  a21716a );
 a21728a <=( A167  and  A168 );
 a21729a <=( (not A170)  and  a21728a );
 a21732a <=( (not A201)  and  (not A166) );
 a21735a <=( A232  and  A202 );
 a21736a <=( a21735a  and  a21732a );
 a21737a <=( a21736a  and  a21729a );
 a21740a <=( A234  and  (not A233) );
 a21743a <=( (not A265)  and  A236 );
 a21744a <=( a21743a  and  a21740a );
 a21747a <=( (not A267)  and  A266 );
 a21750a <=( (not A269)  and  (not A268) );
 a21751a <=( a21750a  and  a21747a );
 a21752a <=( a21751a  and  a21744a );
 a21756a <=( A167  and  A168 );
 a21757a <=( (not A170)  and  a21756a );
 a21760a <=( (not A201)  and  (not A166) );
 a21763a <=( A232  and  A202 );
 a21764a <=( a21763a  and  a21760a );
 a21765a <=( a21764a  and  a21757a );
 a21768a <=( A234  and  (not A233) );
 a21771a <=( A265  and  A236 );
 a21772a <=( a21771a  and  a21768a );
 a21775a <=( (not A267)  and  (not A266) );
 a21778a <=( (not A269)  and  (not A268) );
 a21779a <=( a21778a  and  a21775a );
 a21780a <=( a21779a  and  a21772a );
 a21784a <=( A167  and  A168 );
 a21785a <=( (not A170)  and  a21784a );
 a21788a <=( (not A201)  and  (not A166) );
 a21791a <=( A232  and  A202 );
 a21792a <=( a21791a  and  a21788a );
 a21793a <=( a21792a  and  a21785a );
 a21796a <=( (not A234)  and  (not A233) );
 a21799a <=( (not A236)  and  (not A235) );
 a21800a <=( a21799a  and  a21796a );
 a21803a <=( (not A299)  and  A298 );
 a21806a <=( A301  and  A300 );
 a21807a <=( a21806a  and  a21803a );
 a21808a <=( a21807a  and  a21800a );
 a21812a <=( A167  and  A168 );
 a21813a <=( (not A170)  and  a21812a );
 a21816a <=( (not A201)  and  (not A166) );
 a21819a <=( A232  and  A202 );
 a21820a <=( a21819a  and  a21816a );
 a21821a <=( a21820a  and  a21813a );
 a21824a <=( (not A234)  and  (not A233) );
 a21827a <=( (not A236)  and  (not A235) );
 a21828a <=( a21827a  and  a21824a );
 a21831a <=( (not A299)  and  A298 );
 a21834a <=( A302  and  A300 );
 a21835a <=( a21834a  and  a21831a );
 a21836a <=( a21835a  and  a21828a );
 a21840a <=( A167  and  A168 );
 a21841a <=( (not A170)  and  a21840a );
 a21844a <=( (not A201)  and  (not A166) );
 a21847a <=( A232  and  A202 );
 a21848a <=( a21847a  and  a21844a );
 a21849a <=( a21848a  and  a21841a );
 a21852a <=( (not A234)  and  (not A233) );
 a21855a <=( (not A236)  and  (not A235) );
 a21856a <=( a21855a  and  a21852a );
 a21859a <=( A299  and  (not A298) );
 a21862a <=( A301  and  A300 );
 a21863a <=( a21862a  and  a21859a );
 a21864a <=( a21863a  and  a21856a );
 a21868a <=( A167  and  A168 );
 a21869a <=( (not A170)  and  a21868a );
 a21872a <=( (not A201)  and  (not A166) );
 a21875a <=( A232  and  A202 );
 a21876a <=( a21875a  and  a21872a );
 a21877a <=( a21876a  and  a21869a );
 a21880a <=( (not A234)  and  (not A233) );
 a21883a <=( (not A236)  and  (not A235) );
 a21884a <=( a21883a  and  a21880a );
 a21887a <=( A299  and  (not A298) );
 a21890a <=( A302  and  A300 );
 a21891a <=( a21890a  and  a21887a );
 a21892a <=( a21891a  and  a21884a );
 a21896a <=( A167  and  A168 );
 a21897a <=( (not A170)  and  a21896a );
 a21900a <=( (not A201)  and  (not A166) );
 a21903a <=( A232  and  A202 );
 a21904a <=( a21903a  and  a21900a );
 a21905a <=( a21904a  and  a21897a );
 a21908a <=( (not A234)  and  (not A233) );
 a21911a <=( (not A236)  and  (not A235) );
 a21912a <=( a21911a  and  a21908a );
 a21915a <=( A266  and  (not A265) );
 a21918a <=( A268  and  A267 );
 a21919a <=( a21918a  and  a21915a );
 a21920a <=( a21919a  and  a21912a );
 a21924a <=( A167  and  A168 );
 a21925a <=( (not A170)  and  a21924a );
 a21928a <=( (not A201)  and  (not A166) );
 a21931a <=( A232  and  A202 );
 a21932a <=( a21931a  and  a21928a );
 a21933a <=( a21932a  and  a21925a );
 a21936a <=( (not A234)  and  (not A233) );
 a21939a <=( (not A236)  and  (not A235) );
 a21940a <=( a21939a  and  a21936a );
 a21943a <=( A266  and  (not A265) );
 a21946a <=( A269  and  A267 );
 a21947a <=( a21946a  and  a21943a );
 a21948a <=( a21947a  and  a21940a );
 a21952a <=( A167  and  A168 );
 a21953a <=( (not A170)  and  a21952a );
 a21956a <=( (not A201)  and  (not A166) );
 a21959a <=( A232  and  A202 );
 a21960a <=( a21959a  and  a21956a );
 a21961a <=( a21960a  and  a21953a );
 a21964a <=( (not A234)  and  (not A233) );
 a21967a <=( (not A236)  and  (not A235) );
 a21968a <=( a21967a  and  a21964a );
 a21971a <=( (not A266)  and  A265 );
 a21974a <=( A268  and  A267 );
 a21975a <=( a21974a  and  a21971a );
 a21976a <=( a21975a  and  a21968a );
 a21980a <=( A167  and  A168 );
 a21981a <=( (not A170)  and  a21980a );
 a21984a <=( (not A201)  and  (not A166) );
 a21987a <=( A232  and  A202 );
 a21988a <=( a21987a  and  a21984a );
 a21989a <=( a21988a  and  a21981a );
 a21992a <=( (not A234)  and  (not A233) );
 a21995a <=( (not A236)  and  (not A235) );
 a21996a <=( a21995a  and  a21992a );
 a21999a <=( (not A266)  and  A265 );
 a22002a <=( A269  and  A267 );
 a22003a <=( a22002a  and  a21999a );
 a22004a <=( a22003a  and  a21996a );
 a22008a <=( A167  and  A168 );
 a22009a <=( (not A170)  and  a22008a );
 a22012a <=( (not A201)  and  (not A166) );
 a22015a <=( (not A232)  and  A203 );
 a22016a <=( a22015a  and  a22012a );
 a22017a <=( a22016a  and  a22009a );
 a22020a <=( A234  and  A233 );
 a22023a <=( A298  and  A235 );
 a22024a <=( a22023a  and  a22020a );
 a22027a <=( (not A300)  and  (not A299) );
 a22030a <=( (not A302)  and  (not A301) );
 a22031a <=( a22030a  and  a22027a );
 a22032a <=( a22031a  and  a22024a );
 a22036a <=( A167  and  A168 );
 a22037a <=( (not A170)  and  a22036a );
 a22040a <=( (not A201)  and  (not A166) );
 a22043a <=( (not A232)  and  A203 );
 a22044a <=( a22043a  and  a22040a );
 a22045a <=( a22044a  and  a22037a );
 a22048a <=( A234  and  A233 );
 a22051a <=( (not A298)  and  A235 );
 a22052a <=( a22051a  and  a22048a );
 a22055a <=( (not A300)  and  A299 );
 a22058a <=( (not A302)  and  (not A301) );
 a22059a <=( a22058a  and  a22055a );
 a22060a <=( a22059a  and  a22052a );
 a22064a <=( A167  and  A168 );
 a22065a <=( (not A170)  and  a22064a );
 a22068a <=( (not A201)  and  (not A166) );
 a22071a <=( (not A232)  and  A203 );
 a22072a <=( a22071a  and  a22068a );
 a22073a <=( a22072a  and  a22065a );
 a22076a <=( A234  and  A233 );
 a22079a <=( (not A265)  and  A235 );
 a22080a <=( a22079a  and  a22076a );
 a22083a <=( (not A267)  and  A266 );
 a22086a <=( (not A269)  and  (not A268) );
 a22087a <=( a22086a  and  a22083a );
 a22088a <=( a22087a  and  a22080a );
 a22092a <=( A167  and  A168 );
 a22093a <=( (not A170)  and  a22092a );
 a22096a <=( (not A201)  and  (not A166) );
 a22099a <=( (not A232)  and  A203 );
 a22100a <=( a22099a  and  a22096a );
 a22101a <=( a22100a  and  a22093a );
 a22104a <=( A234  and  A233 );
 a22107a <=( A265  and  A235 );
 a22108a <=( a22107a  and  a22104a );
 a22111a <=( (not A267)  and  (not A266) );
 a22114a <=( (not A269)  and  (not A268) );
 a22115a <=( a22114a  and  a22111a );
 a22116a <=( a22115a  and  a22108a );
 a22120a <=( A167  and  A168 );
 a22121a <=( (not A170)  and  a22120a );
 a22124a <=( (not A201)  and  (not A166) );
 a22127a <=( (not A232)  and  A203 );
 a22128a <=( a22127a  and  a22124a );
 a22129a <=( a22128a  and  a22121a );
 a22132a <=( A234  and  A233 );
 a22135a <=( A298  and  A236 );
 a22136a <=( a22135a  and  a22132a );
 a22139a <=( (not A300)  and  (not A299) );
 a22142a <=( (not A302)  and  (not A301) );
 a22143a <=( a22142a  and  a22139a );
 a22144a <=( a22143a  and  a22136a );
 a22148a <=( A167  and  A168 );
 a22149a <=( (not A170)  and  a22148a );
 a22152a <=( (not A201)  and  (not A166) );
 a22155a <=( (not A232)  and  A203 );
 a22156a <=( a22155a  and  a22152a );
 a22157a <=( a22156a  and  a22149a );
 a22160a <=( A234  and  A233 );
 a22163a <=( (not A298)  and  A236 );
 a22164a <=( a22163a  and  a22160a );
 a22167a <=( (not A300)  and  A299 );
 a22170a <=( (not A302)  and  (not A301) );
 a22171a <=( a22170a  and  a22167a );
 a22172a <=( a22171a  and  a22164a );
 a22176a <=( A167  and  A168 );
 a22177a <=( (not A170)  and  a22176a );
 a22180a <=( (not A201)  and  (not A166) );
 a22183a <=( (not A232)  and  A203 );
 a22184a <=( a22183a  and  a22180a );
 a22185a <=( a22184a  and  a22177a );
 a22188a <=( A234  and  A233 );
 a22191a <=( (not A265)  and  A236 );
 a22192a <=( a22191a  and  a22188a );
 a22195a <=( (not A267)  and  A266 );
 a22198a <=( (not A269)  and  (not A268) );
 a22199a <=( a22198a  and  a22195a );
 a22200a <=( a22199a  and  a22192a );
 a22204a <=( A167  and  A168 );
 a22205a <=( (not A170)  and  a22204a );
 a22208a <=( (not A201)  and  (not A166) );
 a22211a <=( (not A232)  and  A203 );
 a22212a <=( a22211a  and  a22208a );
 a22213a <=( a22212a  and  a22205a );
 a22216a <=( A234  and  A233 );
 a22219a <=( A265  and  A236 );
 a22220a <=( a22219a  and  a22216a );
 a22223a <=( (not A267)  and  (not A266) );
 a22226a <=( (not A269)  and  (not A268) );
 a22227a <=( a22226a  and  a22223a );
 a22228a <=( a22227a  and  a22220a );
 a22232a <=( A167  and  A168 );
 a22233a <=( (not A170)  and  a22232a );
 a22236a <=( (not A201)  and  (not A166) );
 a22239a <=( (not A232)  and  A203 );
 a22240a <=( a22239a  and  a22236a );
 a22241a <=( a22240a  and  a22233a );
 a22244a <=( (not A234)  and  A233 );
 a22247a <=( (not A236)  and  (not A235) );
 a22248a <=( a22247a  and  a22244a );
 a22251a <=( (not A299)  and  A298 );
 a22254a <=( A301  and  A300 );
 a22255a <=( a22254a  and  a22251a );
 a22256a <=( a22255a  and  a22248a );
 a22260a <=( A167  and  A168 );
 a22261a <=( (not A170)  and  a22260a );
 a22264a <=( (not A201)  and  (not A166) );
 a22267a <=( (not A232)  and  A203 );
 a22268a <=( a22267a  and  a22264a );
 a22269a <=( a22268a  and  a22261a );
 a22272a <=( (not A234)  and  A233 );
 a22275a <=( (not A236)  and  (not A235) );
 a22276a <=( a22275a  and  a22272a );
 a22279a <=( (not A299)  and  A298 );
 a22282a <=( A302  and  A300 );
 a22283a <=( a22282a  and  a22279a );
 a22284a <=( a22283a  and  a22276a );
 a22288a <=( A167  and  A168 );
 a22289a <=( (not A170)  and  a22288a );
 a22292a <=( (not A201)  and  (not A166) );
 a22295a <=( (not A232)  and  A203 );
 a22296a <=( a22295a  and  a22292a );
 a22297a <=( a22296a  and  a22289a );
 a22300a <=( (not A234)  and  A233 );
 a22303a <=( (not A236)  and  (not A235) );
 a22304a <=( a22303a  and  a22300a );
 a22307a <=( A299  and  (not A298) );
 a22310a <=( A301  and  A300 );
 a22311a <=( a22310a  and  a22307a );
 a22312a <=( a22311a  and  a22304a );
 a22316a <=( A167  and  A168 );
 a22317a <=( (not A170)  and  a22316a );
 a22320a <=( (not A201)  and  (not A166) );
 a22323a <=( (not A232)  and  A203 );
 a22324a <=( a22323a  and  a22320a );
 a22325a <=( a22324a  and  a22317a );
 a22328a <=( (not A234)  and  A233 );
 a22331a <=( (not A236)  and  (not A235) );
 a22332a <=( a22331a  and  a22328a );
 a22335a <=( A299  and  (not A298) );
 a22338a <=( A302  and  A300 );
 a22339a <=( a22338a  and  a22335a );
 a22340a <=( a22339a  and  a22332a );
 a22344a <=( A167  and  A168 );
 a22345a <=( (not A170)  and  a22344a );
 a22348a <=( (not A201)  and  (not A166) );
 a22351a <=( (not A232)  and  A203 );
 a22352a <=( a22351a  and  a22348a );
 a22353a <=( a22352a  and  a22345a );
 a22356a <=( (not A234)  and  A233 );
 a22359a <=( (not A236)  and  (not A235) );
 a22360a <=( a22359a  and  a22356a );
 a22363a <=( A266  and  (not A265) );
 a22366a <=( A268  and  A267 );
 a22367a <=( a22366a  and  a22363a );
 a22368a <=( a22367a  and  a22360a );
 a22372a <=( A167  and  A168 );
 a22373a <=( (not A170)  and  a22372a );
 a22376a <=( (not A201)  and  (not A166) );
 a22379a <=( (not A232)  and  A203 );
 a22380a <=( a22379a  and  a22376a );
 a22381a <=( a22380a  and  a22373a );
 a22384a <=( (not A234)  and  A233 );
 a22387a <=( (not A236)  and  (not A235) );
 a22388a <=( a22387a  and  a22384a );
 a22391a <=( A266  and  (not A265) );
 a22394a <=( A269  and  A267 );
 a22395a <=( a22394a  and  a22391a );
 a22396a <=( a22395a  and  a22388a );
 a22400a <=( A167  and  A168 );
 a22401a <=( (not A170)  and  a22400a );
 a22404a <=( (not A201)  and  (not A166) );
 a22407a <=( (not A232)  and  A203 );
 a22408a <=( a22407a  and  a22404a );
 a22409a <=( a22408a  and  a22401a );
 a22412a <=( (not A234)  and  A233 );
 a22415a <=( (not A236)  and  (not A235) );
 a22416a <=( a22415a  and  a22412a );
 a22419a <=( (not A266)  and  A265 );
 a22422a <=( A268  and  A267 );
 a22423a <=( a22422a  and  a22419a );
 a22424a <=( a22423a  and  a22416a );
 a22428a <=( A167  and  A168 );
 a22429a <=( (not A170)  and  a22428a );
 a22432a <=( (not A201)  and  (not A166) );
 a22435a <=( (not A232)  and  A203 );
 a22436a <=( a22435a  and  a22432a );
 a22437a <=( a22436a  and  a22429a );
 a22440a <=( (not A234)  and  A233 );
 a22443a <=( (not A236)  and  (not A235) );
 a22444a <=( a22443a  and  a22440a );
 a22447a <=( (not A266)  and  A265 );
 a22450a <=( A269  and  A267 );
 a22451a <=( a22450a  and  a22447a );
 a22452a <=( a22451a  and  a22444a );
 a22456a <=( A167  and  A168 );
 a22457a <=( (not A170)  and  a22456a );
 a22460a <=( (not A201)  and  (not A166) );
 a22463a <=( A232  and  A203 );
 a22464a <=( a22463a  and  a22460a );
 a22465a <=( a22464a  and  a22457a );
 a22468a <=( A234  and  (not A233) );
 a22471a <=( A298  and  A235 );
 a22472a <=( a22471a  and  a22468a );
 a22475a <=( (not A300)  and  (not A299) );
 a22478a <=( (not A302)  and  (not A301) );
 a22479a <=( a22478a  and  a22475a );
 a22480a <=( a22479a  and  a22472a );
 a22484a <=( A167  and  A168 );
 a22485a <=( (not A170)  and  a22484a );
 a22488a <=( (not A201)  and  (not A166) );
 a22491a <=( A232  and  A203 );
 a22492a <=( a22491a  and  a22488a );
 a22493a <=( a22492a  and  a22485a );
 a22496a <=( A234  and  (not A233) );
 a22499a <=( (not A298)  and  A235 );
 a22500a <=( a22499a  and  a22496a );
 a22503a <=( (not A300)  and  A299 );
 a22506a <=( (not A302)  and  (not A301) );
 a22507a <=( a22506a  and  a22503a );
 a22508a <=( a22507a  and  a22500a );
 a22512a <=( A167  and  A168 );
 a22513a <=( (not A170)  and  a22512a );
 a22516a <=( (not A201)  and  (not A166) );
 a22519a <=( A232  and  A203 );
 a22520a <=( a22519a  and  a22516a );
 a22521a <=( a22520a  and  a22513a );
 a22524a <=( A234  and  (not A233) );
 a22527a <=( (not A265)  and  A235 );
 a22528a <=( a22527a  and  a22524a );
 a22531a <=( (not A267)  and  A266 );
 a22534a <=( (not A269)  and  (not A268) );
 a22535a <=( a22534a  and  a22531a );
 a22536a <=( a22535a  and  a22528a );
 a22540a <=( A167  and  A168 );
 a22541a <=( (not A170)  and  a22540a );
 a22544a <=( (not A201)  and  (not A166) );
 a22547a <=( A232  and  A203 );
 a22548a <=( a22547a  and  a22544a );
 a22549a <=( a22548a  and  a22541a );
 a22552a <=( A234  and  (not A233) );
 a22555a <=( A265  and  A235 );
 a22556a <=( a22555a  and  a22552a );
 a22559a <=( (not A267)  and  (not A266) );
 a22562a <=( (not A269)  and  (not A268) );
 a22563a <=( a22562a  and  a22559a );
 a22564a <=( a22563a  and  a22556a );
 a22568a <=( A167  and  A168 );
 a22569a <=( (not A170)  and  a22568a );
 a22572a <=( (not A201)  and  (not A166) );
 a22575a <=( A232  and  A203 );
 a22576a <=( a22575a  and  a22572a );
 a22577a <=( a22576a  and  a22569a );
 a22580a <=( A234  and  (not A233) );
 a22583a <=( A298  and  A236 );
 a22584a <=( a22583a  and  a22580a );
 a22587a <=( (not A300)  and  (not A299) );
 a22590a <=( (not A302)  and  (not A301) );
 a22591a <=( a22590a  and  a22587a );
 a22592a <=( a22591a  and  a22584a );
 a22596a <=( A167  and  A168 );
 a22597a <=( (not A170)  and  a22596a );
 a22600a <=( (not A201)  and  (not A166) );
 a22603a <=( A232  and  A203 );
 a22604a <=( a22603a  and  a22600a );
 a22605a <=( a22604a  and  a22597a );
 a22608a <=( A234  and  (not A233) );
 a22611a <=( (not A298)  and  A236 );
 a22612a <=( a22611a  and  a22608a );
 a22615a <=( (not A300)  and  A299 );
 a22618a <=( (not A302)  and  (not A301) );
 a22619a <=( a22618a  and  a22615a );
 a22620a <=( a22619a  and  a22612a );
 a22624a <=( A167  and  A168 );
 a22625a <=( (not A170)  and  a22624a );
 a22628a <=( (not A201)  and  (not A166) );
 a22631a <=( A232  and  A203 );
 a22632a <=( a22631a  and  a22628a );
 a22633a <=( a22632a  and  a22625a );
 a22636a <=( A234  and  (not A233) );
 a22639a <=( (not A265)  and  A236 );
 a22640a <=( a22639a  and  a22636a );
 a22643a <=( (not A267)  and  A266 );
 a22646a <=( (not A269)  and  (not A268) );
 a22647a <=( a22646a  and  a22643a );
 a22648a <=( a22647a  and  a22640a );
 a22652a <=( A167  and  A168 );
 a22653a <=( (not A170)  and  a22652a );
 a22656a <=( (not A201)  and  (not A166) );
 a22659a <=( A232  and  A203 );
 a22660a <=( a22659a  and  a22656a );
 a22661a <=( a22660a  and  a22653a );
 a22664a <=( A234  and  (not A233) );
 a22667a <=( A265  and  A236 );
 a22668a <=( a22667a  and  a22664a );
 a22671a <=( (not A267)  and  (not A266) );
 a22674a <=( (not A269)  and  (not A268) );
 a22675a <=( a22674a  and  a22671a );
 a22676a <=( a22675a  and  a22668a );
 a22680a <=( A167  and  A168 );
 a22681a <=( (not A170)  and  a22680a );
 a22684a <=( (not A201)  and  (not A166) );
 a22687a <=( A232  and  A203 );
 a22688a <=( a22687a  and  a22684a );
 a22689a <=( a22688a  and  a22681a );
 a22692a <=( (not A234)  and  (not A233) );
 a22695a <=( (not A236)  and  (not A235) );
 a22696a <=( a22695a  and  a22692a );
 a22699a <=( (not A299)  and  A298 );
 a22702a <=( A301  and  A300 );
 a22703a <=( a22702a  and  a22699a );
 a22704a <=( a22703a  and  a22696a );
 a22708a <=( A167  and  A168 );
 a22709a <=( (not A170)  and  a22708a );
 a22712a <=( (not A201)  and  (not A166) );
 a22715a <=( A232  and  A203 );
 a22716a <=( a22715a  and  a22712a );
 a22717a <=( a22716a  and  a22709a );
 a22720a <=( (not A234)  and  (not A233) );
 a22723a <=( (not A236)  and  (not A235) );
 a22724a <=( a22723a  and  a22720a );
 a22727a <=( (not A299)  and  A298 );
 a22730a <=( A302  and  A300 );
 a22731a <=( a22730a  and  a22727a );
 a22732a <=( a22731a  and  a22724a );
 a22736a <=( A167  and  A168 );
 a22737a <=( (not A170)  and  a22736a );
 a22740a <=( (not A201)  and  (not A166) );
 a22743a <=( A232  and  A203 );
 a22744a <=( a22743a  and  a22740a );
 a22745a <=( a22744a  and  a22737a );
 a22748a <=( (not A234)  and  (not A233) );
 a22751a <=( (not A236)  and  (not A235) );
 a22752a <=( a22751a  and  a22748a );
 a22755a <=( A299  and  (not A298) );
 a22758a <=( A301  and  A300 );
 a22759a <=( a22758a  and  a22755a );
 a22760a <=( a22759a  and  a22752a );
 a22764a <=( A167  and  A168 );
 a22765a <=( (not A170)  and  a22764a );
 a22768a <=( (not A201)  and  (not A166) );
 a22771a <=( A232  and  A203 );
 a22772a <=( a22771a  and  a22768a );
 a22773a <=( a22772a  and  a22765a );
 a22776a <=( (not A234)  and  (not A233) );
 a22779a <=( (not A236)  and  (not A235) );
 a22780a <=( a22779a  and  a22776a );
 a22783a <=( A299  and  (not A298) );
 a22786a <=( A302  and  A300 );
 a22787a <=( a22786a  and  a22783a );
 a22788a <=( a22787a  and  a22780a );
 a22792a <=( A167  and  A168 );
 a22793a <=( (not A170)  and  a22792a );
 a22796a <=( (not A201)  and  (not A166) );
 a22799a <=( A232  and  A203 );
 a22800a <=( a22799a  and  a22796a );
 a22801a <=( a22800a  and  a22793a );
 a22804a <=( (not A234)  and  (not A233) );
 a22807a <=( (not A236)  and  (not A235) );
 a22808a <=( a22807a  and  a22804a );
 a22811a <=( A266  and  (not A265) );
 a22814a <=( A268  and  A267 );
 a22815a <=( a22814a  and  a22811a );
 a22816a <=( a22815a  and  a22808a );
 a22820a <=( A167  and  A168 );
 a22821a <=( (not A170)  and  a22820a );
 a22824a <=( (not A201)  and  (not A166) );
 a22827a <=( A232  and  A203 );
 a22828a <=( a22827a  and  a22824a );
 a22829a <=( a22828a  and  a22821a );
 a22832a <=( (not A234)  and  (not A233) );
 a22835a <=( (not A236)  and  (not A235) );
 a22836a <=( a22835a  and  a22832a );
 a22839a <=( A266  and  (not A265) );
 a22842a <=( A269  and  A267 );
 a22843a <=( a22842a  and  a22839a );
 a22844a <=( a22843a  and  a22836a );
 a22848a <=( A167  and  A168 );
 a22849a <=( (not A170)  and  a22848a );
 a22852a <=( (not A201)  and  (not A166) );
 a22855a <=( A232  and  A203 );
 a22856a <=( a22855a  and  a22852a );
 a22857a <=( a22856a  and  a22849a );
 a22860a <=( (not A234)  and  (not A233) );
 a22863a <=( (not A236)  and  (not A235) );
 a22864a <=( a22863a  and  a22860a );
 a22867a <=( (not A266)  and  A265 );
 a22870a <=( A268  and  A267 );
 a22871a <=( a22870a  and  a22867a );
 a22872a <=( a22871a  and  a22864a );
 a22876a <=( A167  and  A168 );
 a22877a <=( (not A170)  and  a22876a );
 a22880a <=( (not A201)  and  (not A166) );
 a22883a <=( A232  and  A203 );
 a22884a <=( a22883a  and  a22880a );
 a22885a <=( a22884a  and  a22877a );
 a22888a <=( (not A234)  and  (not A233) );
 a22891a <=( (not A236)  and  (not A235) );
 a22892a <=( a22891a  and  a22888a );
 a22895a <=( (not A266)  and  A265 );
 a22898a <=( A269  and  A267 );
 a22899a <=( a22898a  and  a22895a );
 a22900a <=( a22899a  and  a22892a );
 a22904a <=( A167  and  A168 );
 a22905a <=( (not A170)  and  a22904a );
 a22908a <=( A199  and  (not A166) );
 a22911a <=( (not A232)  and  A200 );
 a22912a <=( a22911a  and  a22908a );
 a22913a <=( a22912a  and  a22905a );
 a22916a <=( A234  and  A233 );
 a22919a <=( A298  and  A235 );
 a22920a <=( a22919a  and  a22916a );
 a22923a <=( (not A300)  and  (not A299) );
 a22926a <=( (not A302)  and  (not A301) );
 a22927a <=( a22926a  and  a22923a );
 a22928a <=( a22927a  and  a22920a );
 a22932a <=( A167  and  A168 );
 a22933a <=( (not A170)  and  a22932a );
 a22936a <=( A199  and  (not A166) );
 a22939a <=( (not A232)  and  A200 );
 a22940a <=( a22939a  and  a22936a );
 a22941a <=( a22940a  and  a22933a );
 a22944a <=( A234  and  A233 );
 a22947a <=( (not A298)  and  A235 );
 a22948a <=( a22947a  and  a22944a );
 a22951a <=( (not A300)  and  A299 );
 a22954a <=( (not A302)  and  (not A301) );
 a22955a <=( a22954a  and  a22951a );
 a22956a <=( a22955a  and  a22948a );
 a22960a <=( A167  and  A168 );
 a22961a <=( (not A170)  and  a22960a );
 a22964a <=( A199  and  (not A166) );
 a22967a <=( (not A232)  and  A200 );
 a22968a <=( a22967a  and  a22964a );
 a22969a <=( a22968a  and  a22961a );
 a22972a <=( A234  and  A233 );
 a22975a <=( (not A265)  and  A235 );
 a22976a <=( a22975a  and  a22972a );
 a22979a <=( (not A267)  and  A266 );
 a22982a <=( (not A269)  and  (not A268) );
 a22983a <=( a22982a  and  a22979a );
 a22984a <=( a22983a  and  a22976a );
 a22988a <=( A167  and  A168 );
 a22989a <=( (not A170)  and  a22988a );
 a22992a <=( A199  and  (not A166) );
 a22995a <=( (not A232)  and  A200 );
 a22996a <=( a22995a  and  a22992a );
 a22997a <=( a22996a  and  a22989a );
 a23000a <=( A234  and  A233 );
 a23003a <=( A265  and  A235 );
 a23004a <=( a23003a  and  a23000a );
 a23007a <=( (not A267)  and  (not A266) );
 a23010a <=( (not A269)  and  (not A268) );
 a23011a <=( a23010a  and  a23007a );
 a23012a <=( a23011a  and  a23004a );
 a23016a <=( A167  and  A168 );
 a23017a <=( (not A170)  and  a23016a );
 a23020a <=( A199  and  (not A166) );
 a23023a <=( (not A232)  and  A200 );
 a23024a <=( a23023a  and  a23020a );
 a23025a <=( a23024a  and  a23017a );
 a23028a <=( A234  and  A233 );
 a23031a <=( A298  and  A236 );
 a23032a <=( a23031a  and  a23028a );
 a23035a <=( (not A300)  and  (not A299) );
 a23038a <=( (not A302)  and  (not A301) );
 a23039a <=( a23038a  and  a23035a );
 a23040a <=( a23039a  and  a23032a );
 a23044a <=( A167  and  A168 );
 a23045a <=( (not A170)  and  a23044a );
 a23048a <=( A199  and  (not A166) );
 a23051a <=( (not A232)  and  A200 );
 a23052a <=( a23051a  and  a23048a );
 a23053a <=( a23052a  and  a23045a );
 a23056a <=( A234  and  A233 );
 a23059a <=( (not A298)  and  A236 );
 a23060a <=( a23059a  and  a23056a );
 a23063a <=( (not A300)  and  A299 );
 a23066a <=( (not A302)  and  (not A301) );
 a23067a <=( a23066a  and  a23063a );
 a23068a <=( a23067a  and  a23060a );
 a23072a <=( A167  and  A168 );
 a23073a <=( (not A170)  and  a23072a );
 a23076a <=( A199  and  (not A166) );
 a23079a <=( (not A232)  and  A200 );
 a23080a <=( a23079a  and  a23076a );
 a23081a <=( a23080a  and  a23073a );
 a23084a <=( A234  and  A233 );
 a23087a <=( (not A265)  and  A236 );
 a23088a <=( a23087a  and  a23084a );
 a23091a <=( (not A267)  and  A266 );
 a23094a <=( (not A269)  and  (not A268) );
 a23095a <=( a23094a  and  a23091a );
 a23096a <=( a23095a  and  a23088a );
 a23100a <=( A167  and  A168 );
 a23101a <=( (not A170)  and  a23100a );
 a23104a <=( A199  and  (not A166) );
 a23107a <=( (not A232)  and  A200 );
 a23108a <=( a23107a  and  a23104a );
 a23109a <=( a23108a  and  a23101a );
 a23112a <=( A234  and  A233 );
 a23115a <=( A265  and  A236 );
 a23116a <=( a23115a  and  a23112a );
 a23119a <=( (not A267)  and  (not A266) );
 a23122a <=( (not A269)  and  (not A268) );
 a23123a <=( a23122a  and  a23119a );
 a23124a <=( a23123a  and  a23116a );
 a23128a <=( A167  and  A168 );
 a23129a <=( (not A170)  and  a23128a );
 a23132a <=( A199  and  (not A166) );
 a23135a <=( (not A232)  and  A200 );
 a23136a <=( a23135a  and  a23132a );
 a23137a <=( a23136a  and  a23129a );
 a23140a <=( (not A234)  and  A233 );
 a23143a <=( (not A236)  and  (not A235) );
 a23144a <=( a23143a  and  a23140a );
 a23147a <=( (not A299)  and  A298 );
 a23150a <=( A301  and  A300 );
 a23151a <=( a23150a  and  a23147a );
 a23152a <=( a23151a  and  a23144a );
 a23156a <=( A167  and  A168 );
 a23157a <=( (not A170)  and  a23156a );
 a23160a <=( A199  and  (not A166) );
 a23163a <=( (not A232)  and  A200 );
 a23164a <=( a23163a  and  a23160a );
 a23165a <=( a23164a  and  a23157a );
 a23168a <=( (not A234)  and  A233 );
 a23171a <=( (not A236)  and  (not A235) );
 a23172a <=( a23171a  and  a23168a );
 a23175a <=( (not A299)  and  A298 );
 a23178a <=( A302  and  A300 );
 a23179a <=( a23178a  and  a23175a );
 a23180a <=( a23179a  and  a23172a );
 a23184a <=( A167  and  A168 );
 a23185a <=( (not A170)  and  a23184a );
 a23188a <=( A199  and  (not A166) );
 a23191a <=( (not A232)  and  A200 );
 a23192a <=( a23191a  and  a23188a );
 a23193a <=( a23192a  and  a23185a );
 a23196a <=( (not A234)  and  A233 );
 a23199a <=( (not A236)  and  (not A235) );
 a23200a <=( a23199a  and  a23196a );
 a23203a <=( A299  and  (not A298) );
 a23206a <=( A301  and  A300 );
 a23207a <=( a23206a  and  a23203a );
 a23208a <=( a23207a  and  a23200a );
 a23212a <=( A167  and  A168 );
 a23213a <=( (not A170)  and  a23212a );
 a23216a <=( A199  and  (not A166) );
 a23219a <=( (not A232)  and  A200 );
 a23220a <=( a23219a  and  a23216a );
 a23221a <=( a23220a  and  a23213a );
 a23224a <=( (not A234)  and  A233 );
 a23227a <=( (not A236)  and  (not A235) );
 a23228a <=( a23227a  and  a23224a );
 a23231a <=( A299  and  (not A298) );
 a23234a <=( A302  and  A300 );
 a23235a <=( a23234a  and  a23231a );
 a23236a <=( a23235a  and  a23228a );
 a23240a <=( A167  and  A168 );
 a23241a <=( (not A170)  and  a23240a );
 a23244a <=( A199  and  (not A166) );
 a23247a <=( (not A232)  and  A200 );
 a23248a <=( a23247a  and  a23244a );
 a23249a <=( a23248a  and  a23241a );
 a23252a <=( (not A234)  and  A233 );
 a23255a <=( (not A236)  and  (not A235) );
 a23256a <=( a23255a  and  a23252a );
 a23259a <=( A266  and  (not A265) );
 a23262a <=( A268  and  A267 );
 a23263a <=( a23262a  and  a23259a );
 a23264a <=( a23263a  and  a23256a );
 a23268a <=( A167  and  A168 );
 a23269a <=( (not A170)  and  a23268a );
 a23272a <=( A199  and  (not A166) );
 a23275a <=( (not A232)  and  A200 );
 a23276a <=( a23275a  and  a23272a );
 a23277a <=( a23276a  and  a23269a );
 a23280a <=( (not A234)  and  A233 );
 a23283a <=( (not A236)  and  (not A235) );
 a23284a <=( a23283a  and  a23280a );
 a23287a <=( A266  and  (not A265) );
 a23290a <=( A269  and  A267 );
 a23291a <=( a23290a  and  a23287a );
 a23292a <=( a23291a  and  a23284a );
 a23296a <=( A167  and  A168 );
 a23297a <=( (not A170)  and  a23296a );
 a23300a <=( A199  and  (not A166) );
 a23303a <=( (not A232)  and  A200 );
 a23304a <=( a23303a  and  a23300a );
 a23305a <=( a23304a  and  a23297a );
 a23308a <=( (not A234)  and  A233 );
 a23311a <=( (not A236)  and  (not A235) );
 a23312a <=( a23311a  and  a23308a );
 a23315a <=( (not A266)  and  A265 );
 a23318a <=( A268  and  A267 );
 a23319a <=( a23318a  and  a23315a );
 a23320a <=( a23319a  and  a23312a );
 a23324a <=( A167  and  A168 );
 a23325a <=( (not A170)  and  a23324a );
 a23328a <=( A199  and  (not A166) );
 a23331a <=( (not A232)  and  A200 );
 a23332a <=( a23331a  and  a23328a );
 a23333a <=( a23332a  and  a23325a );
 a23336a <=( (not A234)  and  A233 );
 a23339a <=( (not A236)  and  (not A235) );
 a23340a <=( a23339a  and  a23336a );
 a23343a <=( (not A266)  and  A265 );
 a23346a <=( A269  and  A267 );
 a23347a <=( a23346a  and  a23343a );
 a23348a <=( a23347a  and  a23340a );
 a23352a <=( A167  and  A168 );
 a23353a <=( (not A170)  and  a23352a );
 a23356a <=( A199  and  (not A166) );
 a23359a <=( A232  and  A200 );
 a23360a <=( a23359a  and  a23356a );
 a23361a <=( a23360a  and  a23353a );
 a23364a <=( A234  and  (not A233) );
 a23367a <=( A298  and  A235 );
 a23368a <=( a23367a  and  a23364a );
 a23371a <=( (not A300)  and  (not A299) );
 a23374a <=( (not A302)  and  (not A301) );
 a23375a <=( a23374a  and  a23371a );
 a23376a <=( a23375a  and  a23368a );
 a23380a <=( A167  and  A168 );
 a23381a <=( (not A170)  and  a23380a );
 a23384a <=( A199  and  (not A166) );
 a23387a <=( A232  and  A200 );
 a23388a <=( a23387a  and  a23384a );
 a23389a <=( a23388a  and  a23381a );
 a23392a <=( A234  and  (not A233) );
 a23395a <=( (not A298)  and  A235 );
 a23396a <=( a23395a  and  a23392a );
 a23399a <=( (not A300)  and  A299 );
 a23402a <=( (not A302)  and  (not A301) );
 a23403a <=( a23402a  and  a23399a );
 a23404a <=( a23403a  and  a23396a );
 a23408a <=( A167  and  A168 );
 a23409a <=( (not A170)  and  a23408a );
 a23412a <=( A199  and  (not A166) );
 a23415a <=( A232  and  A200 );
 a23416a <=( a23415a  and  a23412a );
 a23417a <=( a23416a  and  a23409a );
 a23420a <=( A234  and  (not A233) );
 a23423a <=( (not A265)  and  A235 );
 a23424a <=( a23423a  and  a23420a );
 a23427a <=( (not A267)  and  A266 );
 a23430a <=( (not A269)  and  (not A268) );
 a23431a <=( a23430a  and  a23427a );
 a23432a <=( a23431a  and  a23424a );
 a23436a <=( A167  and  A168 );
 a23437a <=( (not A170)  and  a23436a );
 a23440a <=( A199  and  (not A166) );
 a23443a <=( A232  and  A200 );
 a23444a <=( a23443a  and  a23440a );
 a23445a <=( a23444a  and  a23437a );
 a23448a <=( A234  and  (not A233) );
 a23451a <=( A265  and  A235 );
 a23452a <=( a23451a  and  a23448a );
 a23455a <=( (not A267)  and  (not A266) );
 a23458a <=( (not A269)  and  (not A268) );
 a23459a <=( a23458a  and  a23455a );
 a23460a <=( a23459a  and  a23452a );
 a23464a <=( A167  and  A168 );
 a23465a <=( (not A170)  and  a23464a );
 a23468a <=( A199  and  (not A166) );
 a23471a <=( A232  and  A200 );
 a23472a <=( a23471a  and  a23468a );
 a23473a <=( a23472a  and  a23465a );
 a23476a <=( A234  and  (not A233) );
 a23479a <=( A298  and  A236 );
 a23480a <=( a23479a  and  a23476a );
 a23483a <=( (not A300)  and  (not A299) );
 a23486a <=( (not A302)  and  (not A301) );
 a23487a <=( a23486a  and  a23483a );
 a23488a <=( a23487a  and  a23480a );
 a23492a <=( A167  and  A168 );
 a23493a <=( (not A170)  and  a23492a );
 a23496a <=( A199  and  (not A166) );
 a23499a <=( A232  and  A200 );
 a23500a <=( a23499a  and  a23496a );
 a23501a <=( a23500a  and  a23493a );
 a23504a <=( A234  and  (not A233) );
 a23507a <=( (not A298)  and  A236 );
 a23508a <=( a23507a  and  a23504a );
 a23511a <=( (not A300)  and  A299 );
 a23514a <=( (not A302)  and  (not A301) );
 a23515a <=( a23514a  and  a23511a );
 a23516a <=( a23515a  and  a23508a );
 a23520a <=( A167  and  A168 );
 a23521a <=( (not A170)  and  a23520a );
 a23524a <=( A199  and  (not A166) );
 a23527a <=( A232  and  A200 );
 a23528a <=( a23527a  and  a23524a );
 a23529a <=( a23528a  and  a23521a );
 a23532a <=( A234  and  (not A233) );
 a23535a <=( (not A265)  and  A236 );
 a23536a <=( a23535a  and  a23532a );
 a23539a <=( (not A267)  and  A266 );
 a23542a <=( (not A269)  and  (not A268) );
 a23543a <=( a23542a  and  a23539a );
 a23544a <=( a23543a  and  a23536a );
 a23548a <=( A167  and  A168 );
 a23549a <=( (not A170)  and  a23548a );
 a23552a <=( A199  and  (not A166) );
 a23555a <=( A232  and  A200 );
 a23556a <=( a23555a  and  a23552a );
 a23557a <=( a23556a  and  a23549a );
 a23560a <=( A234  and  (not A233) );
 a23563a <=( A265  and  A236 );
 a23564a <=( a23563a  and  a23560a );
 a23567a <=( (not A267)  and  (not A266) );
 a23570a <=( (not A269)  and  (not A268) );
 a23571a <=( a23570a  and  a23567a );
 a23572a <=( a23571a  and  a23564a );
 a23576a <=( A167  and  A168 );
 a23577a <=( (not A170)  and  a23576a );
 a23580a <=( A199  and  (not A166) );
 a23583a <=( A232  and  A200 );
 a23584a <=( a23583a  and  a23580a );
 a23585a <=( a23584a  and  a23577a );
 a23588a <=( (not A234)  and  (not A233) );
 a23591a <=( (not A236)  and  (not A235) );
 a23592a <=( a23591a  and  a23588a );
 a23595a <=( (not A299)  and  A298 );
 a23598a <=( A301  and  A300 );
 a23599a <=( a23598a  and  a23595a );
 a23600a <=( a23599a  and  a23592a );
 a23604a <=( A167  and  A168 );
 a23605a <=( (not A170)  and  a23604a );
 a23608a <=( A199  and  (not A166) );
 a23611a <=( A232  and  A200 );
 a23612a <=( a23611a  and  a23608a );
 a23613a <=( a23612a  and  a23605a );
 a23616a <=( (not A234)  and  (not A233) );
 a23619a <=( (not A236)  and  (not A235) );
 a23620a <=( a23619a  and  a23616a );
 a23623a <=( (not A299)  and  A298 );
 a23626a <=( A302  and  A300 );
 a23627a <=( a23626a  and  a23623a );
 a23628a <=( a23627a  and  a23620a );
 a23632a <=( A167  and  A168 );
 a23633a <=( (not A170)  and  a23632a );
 a23636a <=( A199  and  (not A166) );
 a23639a <=( A232  and  A200 );
 a23640a <=( a23639a  and  a23636a );
 a23641a <=( a23640a  and  a23633a );
 a23644a <=( (not A234)  and  (not A233) );
 a23647a <=( (not A236)  and  (not A235) );
 a23648a <=( a23647a  and  a23644a );
 a23651a <=( A299  and  (not A298) );
 a23654a <=( A301  and  A300 );
 a23655a <=( a23654a  and  a23651a );
 a23656a <=( a23655a  and  a23648a );
 a23660a <=( A167  and  A168 );
 a23661a <=( (not A170)  and  a23660a );
 a23664a <=( A199  and  (not A166) );
 a23667a <=( A232  and  A200 );
 a23668a <=( a23667a  and  a23664a );
 a23669a <=( a23668a  and  a23661a );
 a23672a <=( (not A234)  and  (not A233) );
 a23675a <=( (not A236)  and  (not A235) );
 a23676a <=( a23675a  and  a23672a );
 a23679a <=( A299  and  (not A298) );
 a23682a <=( A302  and  A300 );
 a23683a <=( a23682a  and  a23679a );
 a23684a <=( a23683a  and  a23676a );
 a23688a <=( A167  and  A168 );
 a23689a <=( (not A170)  and  a23688a );
 a23692a <=( A199  and  (not A166) );
 a23695a <=( A232  and  A200 );
 a23696a <=( a23695a  and  a23692a );
 a23697a <=( a23696a  and  a23689a );
 a23700a <=( (not A234)  and  (not A233) );
 a23703a <=( (not A236)  and  (not A235) );
 a23704a <=( a23703a  and  a23700a );
 a23707a <=( A266  and  (not A265) );
 a23710a <=( A268  and  A267 );
 a23711a <=( a23710a  and  a23707a );
 a23712a <=( a23711a  and  a23704a );
 a23716a <=( A167  and  A168 );
 a23717a <=( (not A170)  and  a23716a );
 a23720a <=( A199  and  (not A166) );
 a23723a <=( A232  and  A200 );
 a23724a <=( a23723a  and  a23720a );
 a23725a <=( a23724a  and  a23717a );
 a23728a <=( (not A234)  and  (not A233) );
 a23731a <=( (not A236)  and  (not A235) );
 a23732a <=( a23731a  and  a23728a );
 a23735a <=( A266  and  (not A265) );
 a23738a <=( A269  and  A267 );
 a23739a <=( a23738a  and  a23735a );
 a23740a <=( a23739a  and  a23732a );
 a23744a <=( A167  and  A168 );
 a23745a <=( (not A170)  and  a23744a );
 a23748a <=( A199  and  (not A166) );
 a23751a <=( A232  and  A200 );
 a23752a <=( a23751a  and  a23748a );
 a23753a <=( a23752a  and  a23745a );
 a23756a <=( (not A234)  and  (not A233) );
 a23759a <=( (not A236)  and  (not A235) );
 a23760a <=( a23759a  and  a23756a );
 a23763a <=( (not A266)  and  A265 );
 a23766a <=( A268  and  A267 );
 a23767a <=( a23766a  and  a23763a );
 a23768a <=( a23767a  and  a23760a );
 a23772a <=( A167  and  A168 );
 a23773a <=( (not A170)  and  a23772a );
 a23776a <=( A199  and  (not A166) );
 a23779a <=( A232  and  A200 );
 a23780a <=( a23779a  and  a23776a );
 a23781a <=( a23780a  and  a23773a );
 a23784a <=( (not A234)  and  (not A233) );
 a23787a <=( (not A236)  and  (not A235) );
 a23788a <=( a23787a  and  a23784a );
 a23791a <=( (not A266)  and  A265 );
 a23794a <=( A269  and  A267 );
 a23795a <=( a23794a  and  a23791a );
 a23796a <=( a23795a  and  a23788a );
 a23800a <=( A167  and  A168 );
 a23801a <=( (not A170)  and  a23800a );
 a23804a <=( (not A199)  and  (not A166) );
 a23807a <=( (not A232)  and  (not A200) );
 a23808a <=( a23807a  and  a23804a );
 a23809a <=( a23808a  and  a23801a );
 a23812a <=( A234  and  A233 );
 a23815a <=( A298  and  A235 );
 a23816a <=( a23815a  and  a23812a );
 a23819a <=( (not A300)  and  (not A299) );
 a23822a <=( (not A302)  and  (not A301) );
 a23823a <=( a23822a  and  a23819a );
 a23824a <=( a23823a  and  a23816a );
 a23828a <=( A167  and  A168 );
 a23829a <=( (not A170)  and  a23828a );
 a23832a <=( (not A199)  and  (not A166) );
 a23835a <=( (not A232)  and  (not A200) );
 a23836a <=( a23835a  and  a23832a );
 a23837a <=( a23836a  and  a23829a );
 a23840a <=( A234  and  A233 );
 a23843a <=( (not A298)  and  A235 );
 a23844a <=( a23843a  and  a23840a );
 a23847a <=( (not A300)  and  A299 );
 a23850a <=( (not A302)  and  (not A301) );
 a23851a <=( a23850a  and  a23847a );
 a23852a <=( a23851a  and  a23844a );
 a23856a <=( A167  and  A168 );
 a23857a <=( (not A170)  and  a23856a );
 a23860a <=( (not A199)  and  (not A166) );
 a23863a <=( (not A232)  and  (not A200) );
 a23864a <=( a23863a  and  a23860a );
 a23865a <=( a23864a  and  a23857a );
 a23868a <=( A234  and  A233 );
 a23871a <=( (not A265)  and  A235 );
 a23872a <=( a23871a  and  a23868a );
 a23875a <=( (not A267)  and  A266 );
 a23878a <=( (not A269)  and  (not A268) );
 a23879a <=( a23878a  and  a23875a );
 a23880a <=( a23879a  and  a23872a );
 a23884a <=( A167  and  A168 );
 a23885a <=( (not A170)  and  a23884a );
 a23888a <=( (not A199)  and  (not A166) );
 a23891a <=( (not A232)  and  (not A200) );
 a23892a <=( a23891a  and  a23888a );
 a23893a <=( a23892a  and  a23885a );
 a23896a <=( A234  and  A233 );
 a23899a <=( A265  and  A235 );
 a23900a <=( a23899a  and  a23896a );
 a23903a <=( (not A267)  and  (not A266) );
 a23906a <=( (not A269)  and  (not A268) );
 a23907a <=( a23906a  and  a23903a );
 a23908a <=( a23907a  and  a23900a );
 a23912a <=( A167  and  A168 );
 a23913a <=( (not A170)  and  a23912a );
 a23916a <=( (not A199)  and  (not A166) );
 a23919a <=( (not A232)  and  (not A200) );
 a23920a <=( a23919a  and  a23916a );
 a23921a <=( a23920a  and  a23913a );
 a23924a <=( A234  and  A233 );
 a23927a <=( A298  and  A236 );
 a23928a <=( a23927a  and  a23924a );
 a23931a <=( (not A300)  and  (not A299) );
 a23934a <=( (not A302)  and  (not A301) );
 a23935a <=( a23934a  and  a23931a );
 a23936a <=( a23935a  and  a23928a );
 a23940a <=( A167  and  A168 );
 a23941a <=( (not A170)  and  a23940a );
 a23944a <=( (not A199)  and  (not A166) );
 a23947a <=( (not A232)  and  (not A200) );
 a23948a <=( a23947a  and  a23944a );
 a23949a <=( a23948a  and  a23941a );
 a23952a <=( A234  and  A233 );
 a23955a <=( (not A298)  and  A236 );
 a23956a <=( a23955a  and  a23952a );
 a23959a <=( (not A300)  and  A299 );
 a23962a <=( (not A302)  and  (not A301) );
 a23963a <=( a23962a  and  a23959a );
 a23964a <=( a23963a  and  a23956a );
 a23968a <=( A167  and  A168 );
 a23969a <=( (not A170)  and  a23968a );
 a23972a <=( (not A199)  and  (not A166) );
 a23975a <=( (not A232)  and  (not A200) );
 a23976a <=( a23975a  and  a23972a );
 a23977a <=( a23976a  and  a23969a );
 a23980a <=( A234  and  A233 );
 a23983a <=( (not A265)  and  A236 );
 a23984a <=( a23983a  and  a23980a );
 a23987a <=( (not A267)  and  A266 );
 a23990a <=( (not A269)  and  (not A268) );
 a23991a <=( a23990a  and  a23987a );
 a23992a <=( a23991a  and  a23984a );
 a23996a <=( A167  and  A168 );
 a23997a <=( (not A170)  and  a23996a );
 a24000a <=( (not A199)  and  (not A166) );
 a24003a <=( (not A232)  and  (not A200) );
 a24004a <=( a24003a  and  a24000a );
 a24005a <=( a24004a  and  a23997a );
 a24008a <=( A234  and  A233 );
 a24011a <=( A265  and  A236 );
 a24012a <=( a24011a  and  a24008a );
 a24015a <=( (not A267)  and  (not A266) );
 a24018a <=( (not A269)  and  (not A268) );
 a24019a <=( a24018a  and  a24015a );
 a24020a <=( a24019a  and  a24012a );
 a24024a <=( A167  and  A168 );
 a24025a <=( (not A170)  and  a24024a );
 a24028a <=( (not A199)  and  (not A166) );
 a24031a <=( (not A232)  and  (not A200) );
 a24032a <=( a24031a  and  a24028a );
 a24033a <=( a24032a  and  a24025a );
 a24036a <=( (not A234)  and  A233 );
 a24039a <=( (not A236)  and  (not A235) );
 a24040a <=( a24039a  and  a24036a );
 a24043a <=( (not A299)  and  A298 );
 a24046a <=( A301  and  A300 );
 a24047a <=( a24046a  and  a24043a );
 a24048a <=( a24047a  and  a24040a );
 a24052a <=( A167  and  A168 );
 a24053a <=( (not A170)  and  a24052a );
 a24056a <=( (not A199)  and  (not A166) );
 a24059a <=( (not A232)  and  (not A200) );
 a24060a <=( a24059a  and  a24056a );
 a24061a <=( a24060a  and  a24053a );
 a24064a <=( (not A234)  and  A233 );
 a24067a <=( (not A236)  and  (not A235) );
 a24068a <=( a24067a  and  a24064a );
 a24071a <=( (not A299)  and  A298 );
 a24074a <=( A302  and  A300 );
 a24075a <=( a24074a  and  a24071a );
 a24076a <=( a24075a  and  a24068a );
 a24080a <=( A167  and  A168 );
 a24081a <=( (not A170)  and  a24080a );
 a24084a <=( (not A199)  and  (not A166) );
 a24087a <=( (not A232)  and  (not A200) );
 a24088a <=( a24087a  and  a24084a );
 a24089a <=( a24088a  and  a24081a );
 a24092a <=( (not A234)  and  A233 );
 a24095a <=( (not A236)  and  (not A235) );
 a24096a <=( a24095a  and  a24092a );
 a24099a <=( A299  and  (not A298) );
 a24102a <=( A301  and  A300 );
 a24103a <=( a24102a  and  a24099a );
 a24104a <=( a24103a  and  a24096a );
 a24108a <=( A167  and  A168 );
 a24109a <=( (not A170)  and  a24108a );
 a24112a <=( (not A199)  and  (not A166) );
 a24115a <=( (not A232)  and  (not A200) );
 a24116a <=( a24115a  and  a24112a );
 a24117a <=( a24116a  and  a24109a );
 a24120a <=( (not A234)  and  A233 );
 a24123a <=( (not A236)  and  (not A235) );
 a24124a <=( a24123a  and  a24120a );
 a24127a <=( A299  and  (not A298) );
 a24130a <=( A302  and  A300 );
 a24131a <=( a24130a  and  a24127a );
 a24132a <=( a24131a  and  a24124a );
 a24136a <=( A167  and  A168 );
 a24137a <=( (not A170)  and  a24136a );
 a24140a <=( (not A199)  and  (not A166) );
 a24143a <=( (not A232)  and  (not A200) );
 a24144a <=( a24143a  and  a24140a );
 a24145a <=( a24144a  and  a24137a );
 a24148a <=( (not A234)  and  A233 );
 a24151a <=( (not A236)  and  (not A235) );
 a24152a <=( a24151a  and  a24148a );
 a24155a <=( A266  and  (not A265) );
 a24158a <=( A268  and  A267 );
 a24159a <=( a24158a  and  a24155a );
 a24160a <=( a24159a  and  a24152a );
 a24164a <=( A167  and  A168 );
 a24165a <=( (not A170)  and  a24164a );
 a24168a <=( (not A199)  and  (not A166) );
 a24171a <=( (not A232)  and  (not A200) );
 a24172a <=( a24171a  and  a24168a );
 a24173a <=( a24172a  and  a24165a );
 a24176a <=( (not A234)  and  A233 );
 a24179a <=( (not A236)  and  (not A235) );
 a24180a <=( a24179a  and  a24176a );
 a24183a <=( A266  and  (not A265) );
 a24186a <=( A269  and  A267 );
 a24187a <=( a24186a  and  a24183a );
 a24188a <=( a24187a  and  a24180a );
 a24192a <=( A167  and  A168 );
 a24193a <=( (not A170)  and  a24192a );
 a24196a <=( (not A199)  and  (not A166) );
 a24199a <=( (not A232)  and  (not A200) );
 a24200a <=( a24199a  and  a24196a );
 a24201a <=( a24200a  and  a24193a );
 a24204a <=( (not A234)  and  A233 );
 a24207a <=( (not A236)  and  (not A235) );
 a24208a <=( a24207a  and  a24204a );
 a24211a <=( (not A266)  and  A265 );
 a24214a <=( A268  and  A267 );
 a24215a <=( a24214a  and  a24211a );
 a24216a <=( a24215a  and  a24208a );
 a24220a <=( A167  and  A168 );
 a24221a <=( (not A170)  and  a24220a );
 a24224a <=( (not A199)  and  (not A166) );
 a24227a <=( (not A232)  and  (not A200) );
 a24228a <=( a24227a  and  a24224a );
 a24229a <=( a24228a  and  a24221a );
 a24232a <=( (not A234)  and  A233 );
 a24235a <=( (not A236)  and  (not A235) );
 a24236a <=( a24235a  and  a24232a );
 a24239a <=( (not A266)  and  A265 );
 a24242a <=( A269  and  A267 );
 a24243a <=( a24242a  and  a24239a );
 a24244a <=( a24243a  and  a24236a );
 a24248a <=( A167  and  A168 );
 a24249a <=( (not A170)  and  a24248a );
 a24252a <=( (not A199)  and  (not A166) );
 a24255a <=( A232  and  (not A200) );
 a24256a <=( a24255a  and  a24252a );
 a24257a <=( a24256a  and  a24249a );
 a24260a <=( A234  and  (not A233) );
 a24263a <=( A298  and  A235 );
 a24264a <=( a24263a  and  a24260a );
 a24267a <=( (not A300)  and  (not A299) );
 a24270a <=( (not A302)  and  (not A301) );
 a24271a <=( a24270a  and  a24267a );
 a24272a <=( a24271a  and  a24264a );
 a24276a <=( A167  and  A168 );
 a24277a <=( (not A170)  and  a24276a );
 a24280a <=( (not A199)  and  (not A166) );
 a24283a <=( A232  and  (not A200) );
 a24284a <=( a24283a  and  a24280a );
 a24285a <=( a24284a  and  a24277a );
 a24288a <=( A234  and  (not A233) );
 a24291a <=( (not A298)  and  A235 );
 a24292a <=( a24291a  and  a24288a );
 a24295a <=( (not A300)  and  A299 );
 a24298a <=( (not A302)  and  (not A301) );
 a24299a <=( a24298a  and  a24295a );
 a24300a <=( a24299a  and  a24292a );
 a24304a <=( A167  and  A168 );
 a24305a <=( (not A170)  and  a24304a );
 a24308a <=( (not A199)  and  (not A166) );
 a24311a <=( A232  and  (not A200) );
 a24312a <=( a24311a  and  a24308a );
 a24313a <=( a24312a  and  a24305a );
 a24316a <=( A234  and  (not A233) );
 a24319a <=( (not A265)  and  A235 );
 a24320a <=( a24319a  and  a24316a );
 a24323a <=( (not A267)  and  A266 );
 a24326a <=( (not A269)  and  (not A268) );
 a24327a <=( a24326a  and  a24323a );
 a24328a <=( a24327a  and  a24320a );
 a24332a <=( A167  and  A168 );
 a24333a <=( (not A170)  and  a24332a );
 a24336a <=( (not A199)  and  (not A166) );
 a24339a <=( A232  and  (not A200) );
 a24340a <=( a24339a  and  a24336a );
 a24341a <=( a24340a  and  a24333a );
 a24344a <=( A234  and  (not A233) );
 a24347a <=( A265  and  A235 );
 a24348a <=( a24347a  and  a24344a );
 a24351a <=( (not A267)  and  (not A266) );
 a24354a <=( (not A269)  and  (not A268) );
 a24355a <=( a24354a  and  a24351a );
 a24356a <=( a24355a  and  a24348a );
 a24360a <=( A167  and  A168 );
 a24361a <=( (not A170)  and  a24360a );
 a24364a <=( (not A199)  and  (not A166) );
 a24367a <=( A232  and  (not A200) );
 a24368a <=( a24367a  and  a24364a );
 a24369a <=( a24368a  and  a24361a );
 a24372a <=( A234  and  (not A233) );
 a24375a <=( A298  and  A236 );
 a24376a <=( a24375a  and  a24372a );
 a24379a <=( (not A300)  and  (not A299) );
 a24382a <=( (not A302)  and  (not A301) );
 a24383a <=( a24382a  and  a24379a );
 a24384a <=( a24383a  and  a24376a );
 a24388a <=( A167  and  A168 );
 a24389a <=( (not A170)  and  a24388a );
 a24392a <=( (not A199)  and  (not A166) );
 a24395a <=( A232  and  (not A200) );
 a24396a <=( a24395a  and  a24392a );
 a24397a <=( a24396a  and  a24389a );
 a24400a <=( A234  and  (not A233) );
 a24403a <=( (not A298)  and  A236 );
 a24404a <=( a24403a  and  a24400a );
 a24407a <=( (not A300)  and  A299 );
 a24410a <=( (not A302)  and  (not A301) );
 a24411a <=( a24410a  and  a24407a );
 a24412a <=( a24411a  and  a24404a );
 a24416a <=( A167  and  A168 );
 a24417a <=( (not A170)  and  a24416a );
 a24420a <=( (not A199)  and  (not A166) );
 a24423a <=( A232  and  (not A200) );
 a24424a <=( a24423a  and  a24420a );
 a24425a <=( a24424a  and  a24417a );
 a24428a <=( A234  and  (not A233) );
 a24431a <=( (not A265)  and  A236 );
 a24432a <=( a24431a  and  a24428a );
 a24435a <=( (not A267)  and  A266 );
 a24438a <=( (not A269)  and  (not A268) );
 a24439a <=( a24438a  and  a24435a );
 a24440a <=( a24439a  and  a24432a );
 a24444a <=( A167  and  A168 );
 a24445a <=( (not A170)  and  a24444a );
 a24448a <=( (not A199)  and  (not A166) );
 a24451a <=( A232  and  (not A200) );
 a24452a <=( a24451a  and  a24448a );
 a24453a <=( a24452a  and  a24445a );
 a24456a <=( A234  and  (not A233) );
 a24459a <=( A265  and  A236 );
 a24460a <=( a24459a  and  a24456a );
 a24463a <=( (not A267)  and  (not A266) );
 a24466a <=( (not A269)  and  (not A268) );
 a24467a <=( a24466a  and  a24463a );
 a24468a <=( a24467a  and  a24460a );
 a24472a <=( A167  and  A168 );
 a24473a <=( (not A170)  and  a24472a );
 a24476a <=( (not A199)  and  (not A166) );
 a24479a <=( A232  and  (not A200) );
 a24480a <=( a24479a  and  a24476a );
 a24481a <=( a24480a  and  a24473a );
 a24484a <=( (not A234)  and  (not A233) );
 a24487a <=( (not A236)  and  (not A235) );
 a24488a <=( a24487a  and  a24484a );
 a24491a <=( (not A299)  and  A298 );
 a24494a <=( A301  and  A300 );
 a24495a <=( a24494a  and  a24491a );
 a24496a <=( a24495a  and  a24488a );
 a24500a <=( A167  and  A168 );
 a24501a <=( (not A170)  and  a24500a );
 a24504a <=( (not A199)  and  (not A166) );
 a24507a <=( A232  and  (not A200) );
 a24508a <=( a24507a  and  a24504a );
 a24509a <=( a24508a  and  a24501a );
 a24512a <=( (not A234)  and  (not A233) );
 a24515a <=( (not A236)  and  (not A235) );
 a24516a <=( a24515a  and  a24512a );
 a24519a <=( (not A299)  and  A298 );
 a24522a <=( A302  and  A300 );
 a24523a <=( a24522a  and  a24519a );
 a24524a <=( a24523a  and  a24516a );
 a24528a <=( A167  and  A168 );
 a24529a <=( (not A170)  and  a24528a );
 a24532a <=( (not A199)  and  (not A166) );
 a24535a <=( A232  and  (not A200) );
 a24536a <=( a24535a  and  a24532a );
 a24537a <=( a24536a  and  a24529a );
 a24540a <=( (not A234)  and  (not A233) );
 a24543a <=( (not A236)  and  (not A235) );
 a24544a <=( a24543a  and  a24540a );
 a24547a <=( A299  and  (not A298) );
 a24550a <=( A301  and  A300 );
 a24551a <=( a24550a  and  a24547a );
 a24552a <=( a24551a  and  a24544a );
 a24556a <=( A167  and  A168 );
 a24557a <=( (not A170)  and  a24556a );
 a24560a <=( (not A199)  and  (not A166) );
 a24563a <=( A232  and  (not A200) );
 a24564a <=( a24563a  and  a24560a );
 a24565a <=( a24564a  and  a24557a );
 a24568a <=( (not A234)  and  (not A233) );
 a24571a <=( (not A236)  and  (not A235) );
 a24572a <=( a24571a  and  a24568a );
 a24575a <=( A299  and  (not A298) );
 a24578a <=( A302  and  A300 );
 a24579a <=( a24578a  and  a24575a );
 a24580a <=( a24579a  and  a24572a );
 a24584a <=( A167  and  A168 );
 a24585a <=( (not A170)  and  a24584a );
 a24588a <=( (not A199)  and  (not A166) );
 a24591a <=( A232  and  (not A200) );
 a24592a <=( a24591a  and  a24588a );
 a24593a <=( a24592a  and  a24585a );
 a24596a <=( (not A234)  and  (not A233) );
 a24599a <=( (not A236)  and  (not A235) );
 a24600a <=( a24599a  and  a24596a );
 a24603a <=( A266  and  (not A265) );
 a24606a <=( A268  and  A267 );
 a24607a <=( a24606a  and  a24603a );
 a24608a <=( a24607a  and  a24600a );
 a24612a <=( A167  and  A168 );
 a24613a <=( (not A170)  and  a24612a );
 a24616a <=( (not A199)  and  (not A166) );
 a24619a <=( A232  and  (not A200) );
 a24620a <=( a24619a  and  a24616a );
 a24621a <=( a24620a  and  a24613a );
 a24624a <=( (not A234)  and  (not A233) );
 a24627a <=( (not A236)  and  (not A235) );
 a24628a <=( a24627a  and  a24624a );
 a24631a <=( A266  and  (not A265) );
 a24634a <=( A269  and  A267 );
 a24635a <=( a24634a  and  a24631a );
 a24636a <=( a24635a  and  a24628a );
 a24640a <=( A167  and  A168 );
 a24641a <=( (not A170)  and  a24640a );
 a24644a <=( (not A199)  and  (not A166) );
 a24647a <=( A232  and  (not A200) );
 a24648a <=( a24647a  and  a24644a );
 a24649a <=( a24648a  and  a24641a );
 a24652a <=( (not A234)  and  (not A233) );
 a24655a <=( (not A236)  and  (not A235) );
 a24656a <=( a24655a  and  a24652a );
 a24659a <=( (not A266)  and  A265 );
 a24662a <=( A268  and  A267 );
 a24663a <=( a24662a  and  a24659a );
 a24664a <=( a24663a  and  a24656a );
 a24668a <=( A167  and  A168 );
 a24669a <=( (not A170)  and  a24668a );
 a24672a <=( (not A199)  and  (not A166) );
 a24675a <=( A232  and  (not A200) );
 a24676a <=( a24675a  and  a24672a );
 a24677a <=( a24676a  and  a24669a );
 a24680a <=( (not A234)  and  (not A233) );
 a24683a <=( (not A236)  and  (not A235) );
 a24684a <=( a24683a  and  a24680a );
 a24687a <=( (not A266)  and  A265 );
 a24690a <=( A269  and  A267 );
 a24691a <=( a24690a  and  a24687a );
 a24692a <=( a24691a  and  a24684a );
 a24696a <=( (not A167)  and  A168 );
 a24697a <=( (not A170)  and  a24696a );
 a24700a <=( A201  and  A166 );
 a24703a <=( (not A203)  and  (not A202) );
 a24704a <=( a24703a  and  a24700a );
 a24705a <=( a24704a  and  a24697a );
 a24708a <=( A233  and  (not A232) );
 a24711a <=( A235  and  A234 );
 a24712a <=( a24711a  and  a24708a );
 a24715a <=( (not A299)  and  A298 );
 a24718a <=( A301  and  A300 );
 a24719a <=( a24718a  and  a24715a );
 a24720a <=( a24719a  and  a24712a );
 a24724a <=( (not A167)  and  A168 );
 a24725a <=( (not A170)  and  a24724a );
 a24728a <=( A201  and  A166 );
 a24731a <=( (not A203)  and  (not A202) );
 a24732a <=( a24731a  and  a24728a );
 a24733a <=( a24732a  and  a24725a );
 a24736a <=( A233  and  (not A232) );
 a24739a <=( A235  and  A234 );
 a24740a <=( a24739a  and  a24736a );
 a24743a <=( (not A299)  and  A298 );
 a24746a <=( A302  and  A300 );
 a24747a <=( a24746a  and  a24743a );
 a24748a <=( a24747a  and  a24740a );
 a24752a <=( (not A167)  and  A168 );
 a24753a <=( (not A170)  and  a24752a );
 a24756a <=( A201  and  A166 );
 a24759a <=( (not A203)  and  (not A202) );
 a24760a <=( a24759a  and  a24756a );
 a24761a <=( a24760a  and  a24753a );
 a24764a <=( A233  and  (not A232) );
 a24767a <=( A235  and  A234 );
 a24768a <=( a24767a  and  a24764a );
 a24771a <=( A299  and  (not A298) );
 a24774a <=( A301  and  A300 );
 a24775a <=( a24774a  and  a24771a );
 a24776a <=( a24775a  and  a24768a );
 a24780a <=( (not A167)  and  A168 );
 a24781a <=( (not A170)  and  a24780a );
 a24784a <=( A201  and  A166 );
 a24787a <=( (not A203)  and  (not A202) );
 a24788a <=( a24787a  and  a24784a );
 a24789a <=( a24788a  and  a24781a );
 a24792a <=( A233  and  (not A232) );
 a24795a <=( A235  and  A234 );
 a24796a <=( a24795a  and  a24792a );
 a24799a <=( A299  and  (not A298) );
 a24802a <=( A302  and  A300 );
 a24803a <=( a24802a  and  a24799a );
 a24804a <=( a24803a  and  a24796a );
 a24808a <=( (not A167)  and  A168 );
 a24809a <=( (not A170)  and  a24808a );
 a24812a <=( A201  and  A166 );
 a24815a <=( (not A203)  and  (not A202) );
 a24816a <=( a24815a  and  a24812a );
 a24817a <=( a24816a  and  a24809a );
 a24820a <=( A233  and  (not A232) );
 a24823a <=( A235  and  A234 );
 a24824a <=( a24823a  and  a24820a );
 a24827a <=( A266  and  (not A265) );
 a24830a <=( A268  and  A267 );
 a24831a <=( a24830a  and  a24827a );
 a24832a <=( a24831a  and  a24824a );
 a24836a <=( (not A167)  and  A168 );
 a24837a <=( (not A170)  and  a24836a );
 a24840a <=( A201  and  A166 );
 a24843a <=( (not A203)  and  (not A202) );
 a24844a <=( a24843a  and  a24840a );
 a24845a <=( a24844a  and  a24837a );
 a24848a <=( A233  and  (not A232) );
 a24851a <=( A235  and  A234 );
 a24852a <=( a24851a  and  a24848a );
 a24855a <=( A266  and  (not A265) );
 a24858a <=( A269  and  A267 );
 a24859a <=( a24858a  and  a24855a );
 a24860a <=( a24859a  and  a24852a );
 a24864a <=( (not A167)  and  A168 );
 a24865a <=( (not A170)  and  a24864a );
 a24868a <=( A201  and  A166 );
 a24871a <=( (not A203)  and  (not A202) );
 a24872a <=( a24871a  and  a24868a );
 a24873a <=( a24872a  and  a24865a );
 a24876a <=( A233  and  (not A232) );
 a24879a <=( A235  and  A234 );
 a24880a <=( a24879a  and  a24876a );
 a24883a <=( (not A266)  and  A265 );
 a24886a <=( A268  and  A267 );
 a24887a <=( a24886a  and  a24883a );
 a24888a <=( a24887a  and  a24880a );
 a24892a <=( (not A167)  and  A168 );
 a24893a <=( (not A170)  and  a24892a );
 a24896a <=( A201  and  A166 );
 a24899a <=( (not A203)  and  (not A202) );
 a24900a <=( a24899a  and  a24896a );
 a24901a <=( a24900a  and  a24893a );
 a24904a <=( A233  and  (not A232) );
 a24907a <=( A235  and  A234 );
 a24908a <=( a24907a  and  a24904a );
 a24911a <=( (not A266)  and  A265 );
 a24914a <=( A269  and  A267 );
 a24915a <=( a24914a  and  a24911a );
 a24916a <=( a24915a  and  a24908a );
 a24920a <=( (not A167)  and  A168 );
 a24921a <=( (not A170)  and  a24920a );
 a24924a <=( A201  and  A166 );
 a24927a <=( (not A203)  and  (not A202) );
 a24928a <=( a24927a  and  a24924a );
 a24929a <=( a24928a  and  a24921a );
 a24932a <=( A233  and  (not A232) );
 a24935a <=( A236  and  A234 );
 a24936a <=( a24935a  and  a24932a );
 a24939a <=( (not A299)  and  A298 );
 a24942a <=( A301  and  A300 );
 a24943a <=( a24942a  and  a24939a );
 a24944a <=( a24943a  and  a24936a );
 a24948a <=( (not A167)  and  A168 );
 a24949a <=( (not A170)  and  a24948a );
 a24952a <=( A201  and  A166 );
 a24955a <=( (not A203)  and  (not A202) );
 a24956a <=( a24955a  and  a24952a );
 a24957a <=( a24956a  and  a24949a );
 a24960a <=( A233  and  (not A232) );
 a24963a <=( A236  and  A234 );
 a24964a <=( a24963a  and  a24960a );
 a24967a <=( (not A299)  and  A298 );
 a24970a <=( A302  and  A300 );
 a24971a <=( a24970a  and  a24967a );
 a24972a <=( a24971a  and  a24964a );
 a24976a <=( (not A167)  and  A168 );
 a24977a <=( (not A170)  and  a24976a );
 a24980a <=( A201  and  A166 );
 a24983a <=( (not A203)  and  (not A202) );
 a24984a <=( a24983a  and  a24980a );
 a24985a <=( a24984a  and  a24977a );
 a24988a <=( A233  and  (not A232) );
 a24991a <=( A236  and  A234 );
 a24992a <=( a24991a  and  a24988a );
 a24995a <=( A299  and  (not A298) );
 a24998a <=( A301  and  A300 );
 a24999a <=( a24998a  and  a24995a );
 a25000a <=( a24999a  and  a24992a );
 a25004a <=( (not A167)  and  A168 );
 a25005a <=( (not A170)  and  a25004a );
 a25008a <=( A201  and  A166 );
 a25011a <=( (not A203)  and  (not A202) );
 a25012a <=( a25011a  and  a25008a );
 a25013a <=( a25012a  and  a25005a );
 a25016a <=( A233  and  (not A232) );
 a25019a <=( A236  and  A234 );
 a25020a <=( a25019a  and  a25016a );
 a25023a <=( A299  and  (not A298) );
 a25026a <=( A302  and  A300 );
 a25027a <=( a25026a  and  a25023a );
 a25028a <=( a25027a  and  a25020a );
 a25032a <=( (not A167)  and  A168 );
 a25033a <=( (not A170)  and  a25032a );
 a25036a <=( A201  and  A166 );
 a25039a <=( (not A203)  and  (not A202) );
 a25040a <=( a25039a  and  a25036a );
 a25041a <=( a25040a  and  a25033a );
 a25044a <=( A233  and  (not A232) );
 a25047a <=( A236  and  A234 );
 a25048a <=( a25047a  and  a25044a );
 a25051a <=( A266  and  (not A265) );
 a25054a <=( A268  and  A267 );
 a25055a <=( a25054a  and  a25051a );
 a25056a <=( a25055a  and  a25048a );
 a25060a <=( (not A167)  and  A168 );
 a25061a <=( (not A170)  and  a25060a );
 a25064a <=( A201  and  A166 );
 a25067a <=( (not A203)  and  (not A202) );
 a25068a <=( a25067a  and  a25064a );
 a25069a <=( a25068a  and  a25061a );
 a25072a <=( A233  and  (not A232) );
 a25075a <=( A236  and  A234 );
 a25076a <=( a25075a  and  a25072a );
 a25079a <=( A266  and  (not A265) );
 a25082a <=( A269  and  A267 );
 a25083a <=( a25082a  and  a25079a );
 a25084a <=( a25083a  and  a25076a );
 a25088a <=( (not A167)  and  A168 );
 a25089a <=( (not A170)  and  a25088a );
 a25092a <=( A201  and  A166 );
 a25095a <=( (not A203)  and  (not A202) );
 a25096a <=( a25095a  and  a25092a );
 a25097a <=( a25096a  and  a25089a );
 a25100a <=( A233  and  (not A232) );
 a25103a <=( A236  and  A234 );
 a25104a <=( a25103a  and  a25100a );
 a25107a <=( (not A266)  and  A265 );
 a25110a <=( A268  and  A267 );
 a25111a <=( a25110a  and  a25107a );
 a25112a <=( a25111a  and  a25104a );
 a25116a <=( (not A167)  and  A168 );
 a25117a <=( (not A170)  and  a25116a );
 a25120a <=( A201  and  A166 );
 a25123a <=( (not A203)  and  (not A202) );
 a25124a <=( a25123a  and  a25120a );
 a25125a <=( a25124a  and  a25117a );
 a25128a <=( A233  and  (not A232) );
 a25131a <=( A236  and  A234 );
 a25132a <=( a25131a  and  a25128a );
 a25135a <=( (not A266)  and  A265 );
 a25138a <=( A269  and  A267 );
 a25139a <=( a25138a  and  a25135a );
 a25140a <=( a25139a  and  a25132a );
 a25144a <=( (not A167)  and  A168 );
 a25145a <=( (not A170)  and  a25144a );
 a25148a <=( A201  and  A166 );
 a25151a <=( (not A203)  and  (not A202) );
 a25152a <=( a25151a  and  a25148a );
 a25153a <=( a25152a  and  a25145a );
 a25156a <=( (not A233)  and  A232 );
 a25159a <=( A235  and  A234 );
 a25160a <=( a25159a  and  a25156a );
 a25163a <=( (not A299)  and  A298 );
 a25166a <=( A301  and  A300 );
 a25167a <=( a25166a  and  a25163a );
 a25168a <=( a25167a  and  a25160a );
 a25172a <=( (not A167)  and  A168 );
 a25173a <=( (not A170)  and  a25172a );
 a25176a <=( A201  and  A166 );
 a25179a <=( (not A203)  and  (not A202) );
 a25180a <=( a25179a  and  a25176a );
 a25181a <=( a25180a  and  a25173a );
 a25184a <=( (not A233)  and  A232 );
 a25187a <=( A235  and  A234 );
 a25188a <=( a25187a  and  a25184a );
 a25191a <=( (not A299)  and  A298 );
 a25194a <=( A302  and  A300 );
 a25195a <=( a25194a  and  a25191a );
 a25196a <=( a25195a  and  a25188a );
 a25200a <=( (not A167)  and  A168 );
 a25201a <=( (not A170)  and  a25200a );
 a25204a <=( A201  and  A166 );
 a25207a <=( (not A203)  and  (not A202) );
 a25208a <=( a25207a  and  a25204a );
 a25209a <=( a25208a  and  a25201a );
 a25212a <=( (not A233)  and  A232 );
 a25215a <=( A235  and  A234 );
 a25216a <=( a25215a  and  a25212a );
 a25219a <=( A299  and  (not A298) );
 a25222a <=( A301  and  A300 );
 a25223a <=( a25222a  and  a25219a );
 a25224a <=( a25223a  and  a25216a );
 a25228a <=( (not A167)  and  A168 );
 a25229a <=( (not A170)  and  a25228a );
 a25232a <=( A201  and  A166 );
 a25235a <=( (not A203)  and  (not A202) );
 a25236a <=( a25235a  and  a25232a );
 a25237a <=( a25236a  and  a25229a );
 a25240a <=( (not A233)  and  A232 );
 a25243a <=( A235  and  A234 );
 a25244a <=( a25243a  and  a25240a );
 a25247a <=( A299  and  (not A298) );
 a25250a <=( A302  and  A300 );
 a25251a <=( a25250a  and  a25247a );
 a25252a <=( a25251a  and  a25244a );
 a25256a <=( (not A167)  and  A168 );
 a25257a <=( (not A170)  and  a25256a );
 a25260a <=( A201  and  A166 );
 a25263a <=( (not A203)  and  (not A202) );
 a25264a <=( a25263a  and  a25260a );
 a25265a <=( a25264a  and  a25257a );
 a25268a <=( (not A233)  and  A232 );
 a25271a <=( A235  and  A234 );
 a25272a <=( a25271a  and  a25268a );
 a25275a <=( A266  and  (not A265) );
 a25278a <=( A268  and  A267 );
 a25279a <=( a25278a  and  a25275a );
 a25280a <=( a25279a  and  a25272a );
 a25284a <=( (not A167)  and  A168 );
 a25285a <=( (not A170)  and  a25284a );
 a25288a <=( A201  and  A166 );
 a25291a <=( (not A203)  and  (not A202) );
 a25292a <=( a25291a  and  a25288a );
 a25293a <=( a25292a  and  a25285a );
 a25296a <=( (not A233)  and  A232 );
 a25299a <=( A235  and  A234 );
 a25300a <=( a25299a  and  a25296a );
 a25303a <=( A266  and  (not A265) );
 a25306a <=( A269  and  A267 );
 a25307a <=( a25306a  and  a25303a );
 a25308a <=( a25307a  and  a25300a );
 a25312a <=( (not A167)  and  A168 );
 a25313a <=( (not A170)  and  a25312a );
 a25316a <=( A201  and  A166 );
 a25319a <=( (not A203)  and  (not A202) );
 a25320a <=( a25319a  and  a25316a );
 a25321a <=( a25320a  and  a25313a );
 a25324a <=( (not A233)  and  A232 );
 a25327a <=( A235  and  A234 );
 a25328a <=( a25327a  and  a25324a );
 a25331a <=( (not A266)  and  A265 );
 a25334a <=( A268  and  A267 );
 a25335a <=( a25334a  and  a25331a );
 a25336a <=( a25335a  and  a25328a );
 a25340a <=( (not A167)  and  A168 );
 a25341a <=( (not A170)  and  a25340a );
 a25344a <=( A201  and  A166 );
 a25347a <=( (not A203)  and  (not A202) );
 a25348a <=( a25347a  and  a25344a );
 a25349a <=( a25348a  and  a25341a );
 a25352a <=( (not A233)  and  A232 );
 a25355a <=( A235  and  A234 );
 a25356a <=( a25355a  and  a25352a );
 a25359a <=( (not A266)  and  A265 );
 a25362a <=( A269  and  A267 );
 a25363a <=( a25362a  and  a25359a );
 a25364a <=( a25363a  and  a25356a );
 a25368a <=( (not A167)  and  A168 );
 a25369a <=( (not A170)  and  a25368a );
 a25372a <=( A201  and  A166 );
 a25375a <=( (not A203)  and  (not A202) );
 a25376a <=( a25375a  and  a25372a );
 a25377a <=( a25376a  and  a25369a );
 a25380a <=( (not A233)  and  A232 );
 a25383a <=( A236  and  A234 );
 a25384a <=( a25383a  and  a25380a );
 a25387a <=( (not A299)  and  A298 );
 a25390a <=( A301  and  A300 );
 a25391a <=( a25390a  and  a25387a );
 a25392a <=( a25391a  and  a25384a );
 a25396a <=( (not A167)  and  A168 );
 a25397a <=( (not A170)  and  a25396a );
 a25400a <=( A201  and  A166 );
 a25403a <=( (not A203)  and  (not A202) );
 a25404a <=( a25403a  and  a25400a );
 a25405a <=( a25404a  and  a25397a );
 a25408a <=( (not A233)  and  A232 );
 a25411a <=( A236  and  A234 );
 a25412a <=( a25411a  and  a25408a );
 a25415a <=( (not A299)  and  A298 );
 a25418a <=( A302  and  A300 );
 a25419a <=( a25418a  and  a25415a );
 a25420a <=( a25419a  and  a25412a );
 a25424a <=( (not A167)  and  A168 );
 a25425a <=( (not A170)  and  a25424a );
 a25428a <=( A201  and  A166 );
 a25431a <=( (not A203)  and  (not A202) );
 a25432a <=( a25431a  and  a25428a );
 a25433a <=( a25432a  and  a25425a );
 a25436a <=( (not A233)  and  A232 );
 a25439a <=( A236  and  A234 );
 a25440a <=( a25439a  and  a25436a );
 a25443a <=( A299  and  (not A298) );
 a25446a <=( A301  and  A300 );
 a25447a <=( a25446a  and  a25443a );
 a25448a <=( a25447a  and  a25440a );
 a25452a <=( (not A167)  and  A168 );
 a25453a <=( (not A170)  and  a25452a );
 a25456a <=( A201  and  A166 );
 a25459a <=( (not A203)  and  (not A202) );
 a25460a <=( a25459a  and  a25456a );
 a25461a <=( a25460a  and  a25453a );
 a25464a <=( (not A233)  and  A232 );
 a25467a <=( A236  and  A234 );
 a25468a <=( a25467a  and  a25464a );
 a25471a <=( A299  and  (not A298) );
 a25474a <=( A302  and  A300 );
 a25475a <=( a25474a  and  a25471a );
 a25476a <=( a25475a  and  a25468a );
 a25480a <=( (not A167)  and  A168 );
 a25481a <=( (not A170)  and  a25480a );
 a25484a <=( A201  and  A166 );
 a25487a <=( (not A203)  and  (not A202) );
 a25488a <=( a25487a  and  a25484a );
 a25489a <=( a25488a  and  a25481a );
 a25492a <=( (not A233)  and  A232 );
 a25495a <=( A236  and  A234 );
 a25496a <=( a25495a  and  a25492a );
 a25499a <=( A266  and  (not A265) );
 a25502a <=( A268  and  A267 );
 a25503a <=( a25502a  and  a25499a );
 a25504a <=( a25503a  and  a25496a );
 a25508a <=( (not A167)  and  A168 );
 a25509a <=( (not A170)  and  a25508a );
 a25512a <=( A201  and  A166 );
 a25515a <=( (not A203)  and  (not A202) );
 a25516a <=( a25515a  and  a25512a );
 a25517a <=( a25516a  and  a25509a );
 a25520a <=( (not A233)  and  A232 );
 a25523a <=( A236  and  A234 );
 a25524a <=( a25523a  and  a25520a );
 a25527a <=( A266  and  (not A265) );
 a25530a <=( A269  and  A267 );
 a25531a <=( a25530a  and  a25527a );
 a25532a <=( a25531a  and  a25524a );
 a25536a <=( (not A167)  and  A168 );
 a25537a <=( (not A170)  and  a25536a );
 a25540a <=( A201  and  A166 );
 a25543a <=( (not A203)  and  (not A202) );
 a25544a <=( a25543a  and  a25540a );
 a25545a <=( a25544a  and  a25537a );
 a25548a <=( (not A233)  and  A232 );
 a25551a <=( A236  and  A234 );
 a25552a <=( a25551a  and  a25548a );
 a25555a <=( (not A266)  and  A265 );
 a25558a <=( A268  and  A267 );
 a25559a <=( a25558a  and  a25555a );
 a25560a <=( a25559a  and  a25552a );
 a25564a <=( (not A167)  and  A168 );
 a25565a <=( (not A170)  and  a25564a );
 a25568a <=( A201  and  A166 );
 a25571a <=( (not A203)  and  (not A202) );
 a25572a <=( a25571a  and  a25568a );
 a25573a <=( a25572a  and  a25565a );
 a25576a <=( (not A233)  and  A232 );
 a25579a <=( A236  and  A234 );
 a25580a <=( a25579a  and  a25576a );
 a25583a <=( (not A266)  and  A265 );
 a25586a <=( A269  and  A267 );
 a25587a <=( a25586a  and  a25583a );
 a25588a <=( a25587a  and  a25580a );
 a25592a <=( (not A167)  and  A168 );
 a25593a <=( (not A170)  and  a25592a );
 a25596a <=( (not A201)  and  A166 );
 a25599a <=( (not A232)  and  A202 );
 a25600a <=( a25599a  and  a25596a );
 a25601a <=( a25600a  and  a25593a );
 a25604a <=( A234  and  A233 );
 a25607a <=( A298  and  A235 );
 a25608a <=( a25607a  and  a25604a );
 a25611a <=( (not A300)  and  (not A299) );
 a25614a <=( (not A302)  and  (not A301) );
 a25615a <=( a25614a  and  a25611a );
 a25616a <=( a25615a  and  a25608a );
 a25620a <=( (not A167)  and  A168 );
 a25621a <=( (not A170)  and  a25620a );
 a25624a <=( (not A201)  and  A166 );
 a25627a <=( (not A232)  and  A202 );
 a25628a <=( a25627a  and  a25624a );
 a25629a <=( a25628a  and  a25621a );
 a25632a <=( A234  and  A233 );
 a25635a <=( (not A298)  and  A235 );
 a25636a <=( a25635a  and  a25632a );
 a25639a <=( (not A300)  and  A299 );
 a25642a <=( (not A302)  and  (not A301) );
 a25643a <=( a25642a  and  a25639a );
 a25644a <=( a25643a  and  a25636a );
 a25648a <=( (not A167)  and  A168 );
 a25649a <=( (not A170)  and  a25648a );
 a25652a <=( (not A201)  and  A166 );
 a25655a <=( (not A232)  and  A202 );
 a25656a <=( a25655a  and  a25652a );
 a25657a <=( a25656a  and  a25649a );
 a25660a <=( A234  and  A233 );
 a25663a <=( (not A265)  and  A235 );
 a25664a <=( a25663a  and  a25660a );
 a25667a <=( (not A267)  and  A266 );
 a25670a <=( (not A269)  and  (not A268) );
 a25671a <=( a25670a  and  a25667a );
 a25672a <=( a25671a  and  a25664a );
 a25676a <=( (not A167)  and  A168 );
 a25677a <=( (not A170)  and  a25676a );
 a25680a <=( (not A201)  and  A166 );
 a25683a <=( (not A232)  and  A202 );
 a25684a <=( a25683a  and  a25680a );
 a25685a <=( a25684a  and  a25677a );
 a25688a <=( A234  and  A233 );
 a25691a <=( A265  and  A235 );
 a25692a <=( a25691a  and  a25688a );
 a25695a <=( (not A267)  and  (not A266) );
 a25698a <=( (not A269)  and  (not A268) );
 a25699a <=( a25698a  and  a25695a );
 a25700a <=( a25699a  and  a25692a );
 a25704a <=( (not A167)  and  A168 );
 a25705a <=( (not A170)  and  a25704a );
 a25708a <=( (not A201)  and  A166 );
 a25711a <=( (not A232)  and  A202 );
 a25712a <=( a25711a  and  a25708a );
 a25713a <=( a25712a  and  a25705a );
 a25716a <=( A234  and  A233 );
 a25719a <=( A298  and  A236 );
 a25720a <=( a25719a  and  a25716a );
 a25723a <=( (not A300)  and  (not A299) );
 a25726a <=( (not A302)  and  (not A301) );
 a25727a <=( a25726a  and  a25723a );
 a25728a <=( a25727a  and  a25720a );
 a25732a <=( (not A167)  and  A168 );
 a25733a <=( (not A170)  and  a25732a );
 a25736a <=( (not A201)  and  A166 );
 a25739a <=( (not A232)  and  A202 );
 a25740a <=( a25739a  and  a25736a );
 a25741a <=( a25740a  and  a25733a );
 a25744a <=( A234  and  A233 );
 a25747a <=( (not A298)  and  A236 );
 a25748a <=( a25747a  and  a25744a );
 a25751a <=( (not A300)  and  A299 );
 a25754a <=( (not A302)  and  (not A301) );
 a25755a <=( a25754a  and  a25751a );
 a25756a <=( a25755a  and  a25748a );
 a25760a <=( (not A167)  and  A168 );
 a25761a <=( (not A170)  and  a25760a );
 a25764a <=( (not A201)  and  A166 );
 a25767a <=( (not A232)  and  A202 );
 a25768a <=( a25767a  and  a25764a );
 a25769a <=( a25768a  and  a25761a );
 a25772a <=( A234  and  A233 );
 a25775a <=( (not A265)  and  A236 );
 a25776a <=( a25775a  and  a25772a );
 a25779a <=( (not A267)  and  A266 );
 a25782a <=( (not A269)  and  (not A268) );
 a25783a <=( a25782a  and  a25779a );
 a25784a <=( a25783a  and  a25776a );
 a25788a <=( (not A167)  and  A168 );
 a25789a <=( (not A170)  and  a25788a );
 a25792a <=( (not A201)  and  A166 );
 a25795a <=( (not A232)  and  A202 );
 a25796a <=( a25795a  and  a25792a );
 a25797a <=( a25796a  and  a25789a );
 a25800a <=( A234  and  A233 );
 a25803a <=( A265  and  A236 );
 a25804a <=( a25803a  and  a25800a );
 a25807a <=( (not A267)  and  (not A266) );
 a25810a <=( (not A269)  and  (not A268) );
 a25811a <=( a25810a  and  a25807a );
 a25812a <=( a25811a  and  a25804a );
 a25816a <=( (not A167)  and  A168 );
 a25817a <=( (not A170)  and  a25816a );
 a25820a <=( (not A201)  and  A166 );
 a25823a <=( (not A232)  and  A202 );
 a25824a <=( a25823a  and  a25820a );
 a25825a <=( a25824a  and  a25817a );
 a25828a <=( (not A234)  and  A233 );
 a25831a <=( (not A236)  and  (not A235) );
 a25832a <=( a25831a  and  a25828a );
 a25835a <=( (not A299)  and  A298 );
 a25838a <=( A301  and  A300 );
 a25839a <=( a25838a  and  a25835a );
 a25840a <=( a25839a  and  a25832a );
 a25844a <=( (not A167)  and  A168 );
 a25845a <=( (not A170)  and  a25844a );
 a25848a <=( (not A201)  and  A166 );
 a25851a <=( (not A232)  and  A202 );
 a25852a <=( a25851a  and  a25848a );
 a25853a <=( a25852a  and  a25845a );
 a25856a <=( (not A234)  and  A233 );
 a25859a <=( (not A236)  and  (not A235) );
 a25860a <=( a25859a  and  a25856a );
 a25863a <=( (not A299)  and  A298 );
 a25866a <=( A302  and  A300 );
 a25867a <=( a25866a  and  a25863a );
 a25868a <=( a25867a  and  a25860a );
 a25872a <=( (not A167)  and  A168 );
 a25873a <=( (not A170)  and  a25872a );
 a25876a <=( (not A201)  and  A166 );
 a25879a <=( (not A232)  and  A202 );
 a25880a <=( a25879a  and  a25876a );
 a25881a <=( a25880a  and  a25873a );
 a25884a <=( (not A234)  and  A233 );
 a25887a <=( (not A236)  and  (not A235) );
 a25888a <=( a25887a  and  a25884a );
 a25891a <=( A299  and  (not A298) );
 a25894a <=( A301  and  A300 );
 a25895a <=( a25894a  and  a25891a );
 a25896a <=( a25895a  and  a25888a );
 a25900a <=( (not A167)  and  A168 );
 a25901a <=( (not A170)  and  a25900a );
 a25904a <=( (not A201)  and  A166 );
 a25907a <=( (not A232)  and  A202 );
 a25908a <=( a25907a  and  a25904a );
 a25909a <=( a25908a  and  a25901a );
 a25912a <=( (not A234)  and  A233 );
 a25915a <=( (not A236)  and  (not A235) );
 a25916a <=( a25915a  and  a25912a );
 a25919a <=( A299  and  (not A298) );
 a25922a <=( A302  and  A300 );
 a25923a <=( a25922a  and  a25919a );
 a25924a <=( a25923a  and  a25916a );
 a25928a <=( (not A167)  and  A168 );
 a25929a <=( (not A170)  and  a25928a );
 a25932a <=( (not A201)  and  A166 );
 a25935a <=( (not A232)  and  A202 );
 a25936a <=( a25935a  and  a25932a );
 a25937a <=( a25936a  and  a25929a );
 a25940a <=( (not A234)  and  A233 );
 a25943a <=( (not A236)  and  (not A235) );
 a25944a <=( a25943a  and  a25940a );
 a25947a <=( A266  and  (not A265) );
 a25950a <=( A268  and  A267 );
 a25951a <=( a25950a  and  a25947a );
 a25952a <=( a25951a  and  a25944a );
 a25956a <=( (not A167)  and  A168 );
 a25957a <=( (not A170)  and  a25956a );
 a25960a <=( (not A201)  and  A166 );
 a25963a <=( (not A232)  and  A202 );
 a25964a <=( a25963a  and  a25960a );
 a25965a <=( a25964a  and  a25957a );
 a25968a <=( (not A234)  and  A233 );
 a25971a <=( (not A236)  and  (not A235) );
 a25972a <=( a25971a  and  a25968a );
 a25975a <=( A266  and  (not A265) );
 a25978a <=( A269  and  A267 );
 a25979a <=( a25978a  and  a25975a );
 a25980a <=( a25979a  and  a25972a );
 a25984a <=( (not A167)  and  A168 );
 a25985a <=( (not A170)  and  a25984a );
 a25988a <=( (not A201)  and  A166 );
 a25991a <=( (not A232)  and  A202 );
 a25992a <=( a25991a  and  a25988a );
 a25993a <=( a25992a  and  a25985a );
 a25996a <=( (not A234)  and  A233 );
 a25999a <=( (not A236)  and  (not A235) );
 a26000a <=( a25999a  and  a25996a );
 a26003a <=( (not A266)  and  A265 );
 a26006a <=( A268  and  A267 );
 a26007a <=( a26006a  and  a26003a );
 a26008a <=( a26007a  and  a26000a );
 a26012a <=( (not A167)  and  A168 );
 a26013a <=( (not A170)  and  a26012a );
 a26016a <=( (not A201)  and  A166 );
 a26019a <=( (not A232)  and  A202 );
 a26020a <=( a26019a  and  a26016a );
 a26021a <=( a26020a  and  a26013a );
 a26024a <=( (not A234)  and  A233 );
 a26027a <=( (not A236)  and  (not A235) );
 a26028a <=( a26027a  and  a26024a );
 a26031a <=( (not A266)  and  A265 );
 a26034a <=( A269  and  A267 );
 a26035a <=( a26034a  and  a26031a );
 a26036a <=( a26035a  and  a26028a );
 a26040a <=( (not A167)  and  A168 );
 a26041a <=( (not A170)  and  a26040a );
 a26044a <=( (not A201)  and  A166 );
 a26047a <=( A232  and  A202 );
 a26048a <=( a26047a  and  a26044a );
 a26049a <=( a26048a  and  a26041a );
 a26052a <=( A234  and  (not A233) );
 a26055a <=( A298  and  A235 );
 a26056a <=( a26055a  and  a26052a );
 a26059a <=( (not A300)  and  (not A299) );
 a26062a <=( (not A302)  and  (not A301) );
 a26063a <=( a26062a  and  a26059a );
 a26064a <=( a26063a  and  a26056a );
 a26068a <=( (not A167)  and  A168 );
 a26069a <=( (not A170)  and  a26068a );
 a26072a <=( (not A201)  and  A166 );
 a26075a <=( A232  and  A202 );
 a26076a <=( a26075a  and  a26072a );
 a26077a <=( a26076a  and  a26069a );
 a26080a <=( A234  and  (not A233) );
 a26083a <=( (not A298)  and  A235 );
 a26084a <=( a26083a  and  a26080a );
 a26087a <=( (not A300)  and  A299 );
 a26090a <=( (not A302)  and  (not A301) );
 a26091a <=( a26090a  and  a26087a );
 a26092a <=( a26091a  and  a26084a );
 a26096a <=( (not A167)  and  A168 );
 a26097a <=( (not A170)  and  a26096a );
 a26100a <=( (not A201)  and  A166 );
 a26103a <=( A232  and  A202 );
 a26104a <=( a26103a  and  a26100a );
 a26105a <=( a26104a  and  a26097a );
 a26108a <=( A234  and  (not A233) );
 a26111a <=( (not A265)  and  A235 );
 a26112a <=( a26111a  and  a26108a );
 a26115a <=( (not A267)  and  A266 );
 a26118a <=( (not A269)  and  (not A268) );
 a26119a <=( a26118a  and  a26115a );
 a26120a <=( a26119a  and  a26112a );
 a26124a <=( (not A167)  and  A168 );
 a26125a <=( (not A170)  and  a26124a );
 a26128a <=( (not A201)  and  A166 );
 a26131a <=( A232  and  A202 );
 a26132a <=( a26131a  and  a26128a );
 a26133a <=( a26132a  and  a26125a );
 a26136a <=( A234  and  (not A233) );
 a26139a <=( A265  and  A235 );
 a26140a <=( a26139a  and  a26136a );
 a26143a <=( (not A267)  and  (not A266) );
 a26146a <=( (not A269)  and  (not A268) );
 a26147a <=( a26146a  and  a26143a );
 a26148a <=( a26147a  and  a26140a );
 a26152a <=( (not A167)  and  A168 );
 a26153a <=( (not A170)  and  a26152a );
 a26156a <=( (not A201)  and  A166 );
 a26159a <=( A232  and  A202 );
 a26160a <=( a26159a  and  a26156a );
 a26161a <=( a26160a  and  a26153a );
 a26164a <=( A234  and  (not A233) );
 a26167a <=( A298  and  A236 );
 a26168a <=( a26167a  and  a26164a );
 a26171a <=( (not A300)  and  (not A299) );
 a26174a <=( (not A302)  and  (not A301) );
 a26175a <=( a26174a  and  a26171a );
 a26176a <=( a26175a  and  a26168a );
 a26180a <=( (not A167)  and  A168 );
 a26181a <=( (not A170)  and  a26180a );
 a26184a <=( (not A201)  and  A166 );
 a26187a <=( A232  and  A202 );
 a26188a <=( a26187a  and  a26184a );
 a26189a <=( a26188a  and  a26181a );
 a26192a <=( A234  and  (not A233) );
 a26195a <=( (not A298)  and  A236 );
 a26196a <=( a26195a  and  a26192a );
 a26199a <=( (not A300)  and  A299 );
 a26202a <=( (not A302)  and  (not A301) );
 a26203a <=( a26202a  and  a26199a );
 a26204a <=( a26203a  and  a26196a );
 a26208a <=( (not A167)  and  A168 );
 a26209a <=( (not A170)  and  a26208a );
 a26212a <=( (not A201)  and  A166 );
 a26215a <=( A232  and  A202 );
 a26216a <=( a26215a  and  a26212a );
 a26217a <=( a26216a  and  a26209a );
 a26220a <=( A234  and  (not A233) );
 a26223a <=( (not A265)  and  A236 );
 a26224a <=( a26223a  and  a26220a );
 a26227a <=( (not A267)  and  A266 );
 a26230a <=( (not A269)  and  (not A268) );
 a26231a <=( a26230a  and  a26227a );
 a26232a <=( a26231a  and  a26224a );
 a26236a <=( (not A167)  and  A168 );
 a26237a <=( (not A170)  and  a26236a );
 a26240a <=( (not A201)  and  A166 );
 a26243a <=( A232  and  A202 );
 a26244a <=( a26243a  and  a26240a );
 a26245a <=( a26244a  and  a26237a );
 a26248a <=( A234  and  (not A233) );
 a26251a <=( A265  and  A236 );
 a26252a <=( a26251a  and  a26248a );
 a26255a <=( (not A267)  and  (not A266) );
 a26258a <=( (not A269)  and  (not A268) );
 a26259a <=( a26258a  and  a26255a );
 a26260a <=( a26259a  and  a26252a );
 a26264a <=( (not A167)  and  A168 );
 a26265a <=( (not A170)  and  a26264a );
 a26268a <=( (not A201)  and  A166 );
 a26271a <=( A232  and  A202 );
 a26272a <=( a26271a  and  a26268a );
 a26273a <=( a26272a  and  a26265a );
 a26276a <=( (not A234)  and  (not A233) );
 a26279a <=( (not A236)  and  (not A235) );
 a26280a <=( a26279a  and  a26276a );
 a26283a <=( (not A299)  and  A298 );
 a26286a <=( A301  and  A300 );
 a26287a <=( a26286a  and  a26283a );
 a26288a <=( a26287a  and  a26280a );
 a26292a <=( (not A167)  and  A168 );
 a26293a <=( (not A170)  and  a26292a );
 a26296a <=( (not A201)  and  A166 );
 a26299a <=( A232  and  A202 );
 a26300a <=( a26299a  and  a26296a );
 a26301a <=( a26300a  and  a26293a );
 a26304a <=( (not A234)  and  (not A233) );
 a26307a <=( (not A236)  and  (not A235) );
 a26308a <=( a26307a  and  a26304a );
 a26311a <=( (not A299)  and  A298 );
 a26314a <=( A302  and  A300 );
 a26315a <=( a26314a  and  a26311a );
 a26316a <=( a26315a  and  a26308a );
 a26320a <=( (not A167)  and  A168 );
 a26321a <=( (not A170)  and  a26320a );
 a26324a <=( (not A201)  and  A166 );
 a26327a <=( A232  and  A202 );
 a26328a <=( a26327a  and  a26324a );
 a26329a <=( a26328a  and  a26321a );
 a26332a <=( (not A234)  and  (not A233) );
 a26335a <=( (not A236)  and  (not A235) );
 a26336a <=( a26335a  and  a26332a );
 a26339a <=( A299  and  (not A298) );
 a26342a <=( A301  and  A300 );
 a26343a <=( a26342a  and  a26339a );
 a26344a <=( a26343a  and  a26336a );
 a26348a <=( (not A167)  and  A168 );
 a26349a <=( (not A170)  and  a26348a );
 a26352a <=( (not A201)  and  A166 );
 a26355a <=( A232  and  A202 );
 a26356a <=( a26355a  and  a26352a );
 a26357a <=( a26356a  and  a26349a );
 a26360a <=( (not A234)  and  (not A233) );
 a26363a <=( (not A236)  and  (not A235) );
 a26364a <=( a26363a  and  a26360a );
 a26367a <=( A299  and  (not A298) );
 a26370a <=( A302  and  A300 );
 a26371a <=( a26370a  and  a26367a );
 a26372a <=( a26371a  and  a26364a );
 a26376a <=( (not A167)  and  A168 );
 a26377a <=( (not A170)  and  a26376a );
 a26380a <=( (not A201)  and  A166 );
 a26383a <=( A232  and  A202 );
 a26384a <=( a26383a  and  a26380a );
 a26385a <=( a26384a  and  a26377a );
 a26388a <=( (not A234)  and  (not A233) );
 a26391a <=( (not A236)  and  (not A235) );
 a26392a <=( a26391a  and  a26388a );
 a26395a <=( A266  and  (not A265) );
 a26398a <=( A268  and  A267 );
 a26399a <=( a26398a  and  a26395a );
 a26400a <=( a26399a  and  a26392a );
 a26404a <=( (not A167)  and  A168 );
 a26405a <=( (not A170)  and  a26404a );
 a26408a <=( (not A201)  and  A166 );
 a26411a <=( A232  and  A202 );
 a26412a <=( a26411a  and  a26408a );
 a26413a <=( a26412a  and  a26405a );
 a26416a <=( (not A234)  and  (not A233) );
 a26419a <=( (not A236)  and  (not A235) );
 a26420a <=( a26419a  and  a26416a );
 a26423a <=( A266  and  (not A265) );
 a26426a <=( A269  and  A267 );
 a26427a <=( a26426a  and  a26423a );
 a26428a <=( a26427a  and  a26420a );
 a26432a <=( (not A167)  and  A168 );
 a26433a <=( (not A170)  and  a26432a );
 a26436a <=( (not A201)  and  A166 );
 a26439a <=( A232  and  A202 );
 a26440a <=( a26439a  and  a26436a );
 a26441a <=( a26440a  and  a26433a );
 a26444a <=( (not A234)  and  (not A233) );
 a26447a <=( (not A236)  and  (not A235) );
 a26448a <=( a26447a  and  a26444a );
 a26451a <=( (not A266)  and  A265 );
 a26454a <=( A268  and  A267 );
 a26455a <=( a26454a  and  a26451a );
 a26456a <=( a26455a  and  a26448a );
 a26460a <=( (not A167)  and  A168 );
 a26461a <=( (not A170)  and  a26460a );
 a26464a <=( (not A201)  and  A166 );
 a26467a <=( A232  and  A202 );
 a26468a <=( a26467a  and  a26464a );
 a26469a <=( a26468a  and  a26461a );
 a26472a <=( (not A234)  and  (not A233) );
 a26475a <=( (not A236)  and  (not A235) );
 a26476a <=( a26475a  and  a26472a );
 a26479a <=( (not A266)  and  A265 );
 a26482a <=( A269  and  A267 );
 a26483a <=( a26482a  and  a26479a );
 a26484a <=( a26483a  and  a26476a );
 a26488a <=( (not A167)  and  A168 );
 a26489a <=( (not A170)  and  a26488a );
 a26492a <=( (not A201)  and  A166 );
 a26495a <=( (not A232)  and  A203 );
 a26496a <=( a26495a  and  a26492a );
 a26497a <=( a26496a  and  a26489a );
 a26500a <=( A234  and  A233 );
 a26503a <=( A298  and  A235 );
 a26504a <=( a26503a  and  a26500a );
 a26507a <=( (not A300)  and  (not A299) );
 a26510a <=( (not A302)  and  (not A301) );
 a26511a <=( a26510a  and  a26507a );
 a26512a <=( a26511a  and  a26504a );
 a26516a <=( (not A167)  and  A168 );
 a26517a <=( (not A170)  and  a26516a );
 a26520a <=( (not A201)  and  A166 );
 a26523a <=( (not A232)  and  A203 );
 a26524a <=( a26523a  and  a26520a );
 a26525a <=( a26524a  and  a26517a );
 a26528a <=( A234  and  A233 );
 a26531a <=( (not A298)  and  A235 );
 a26532a <=( a26531a  and  a26528a );
 a26535a <=( (not A300)  and  A299 );
 a26538a <=( (not A302)  and  (not A301) );
 a26539a <=( a26538a  and  a26535a );
 a26540a <=( a26539a  and  a26532a );
 a26544a <=( (not A167)  and  A168 );
 a26545a <=( (not A170)  and  a26544a );
 a26548a <=( (not A201)  and  A166 );
 a26551a <=( (not A232)  and  A203 );
 a26552a <=( a26551a  and  a26548a );
 a26553a <=( a26552a  and  a26545a );
 a26556a <=( A234  and  A233 );
 a26559a <=( (not A265)  and  A235 );
 a26560a <=( a26559a  and  a26556a );
 a26563a <=( (not A267)  and  A266 );
 a26566a <=( (not A269)  and  (not A268) );
 a26567a <=( a26566a  and  a26563a );
 a26568a <=( a26567a  and  a26560a );
 a26572a <=( (not A167)  and  A168 );
 a26573a <=( (not A170)  and  a26572a );
 a26576a <=( (not A201)  and  A166 );
 a26579a <=( (not A232)  and  A203 );
 a26580a <=( a26579a  and  a26576a );
 a26581a <=( a26580a  and  a26573a );
 a26584a <=( A234  and  A233 );
 a26587a <=( A265  and  A235 );
 a26588a <=( a26587a  and  a26584a );
 a26591a <=( (not A267)  and  (not A266) );
 a26594a <=( (not A269)  and  (not A268) );
 a26595a <=( a26594a  and  a26591a );
 a26596a <=( a26595a  and  a26588a );
 a26600a <=( (not A167)  and  A168 );
 a26601a <=( (not A170)  and  a26600a );
 a26604a <=( (not A201)  and  A166 );
 a26607a <=( (not A232)  and  A203 );
 a26608a <=( a26607a  and  a26604a );
 a26609a <=( a26608a  and  a26601a );
 a26612a <=( A234  and  A233 );
 a26615a <=( A298  and  A236 );
 a26616a <=( a26615a  and  a26612a );
 a26619a <=( (not A300)  and  (not A299) );
 a26622a <=( (not A302)  and  (not A301) );
 a26623a <=( a26622a  and  a26619a );
 a26624a <=( a26623a  and  a26616a );
 a26628a <=( (not A167)  and  A168 );
 a26629a <=( (not A170)  and  a26628a );
 a26632a <=( (not A201)  and  A166 );
 a26635a <=( (not A232)  and  A203 );
 a26636a <=( a26635a  and  a26632a );
 a26637a <=( a26636a  and  a26629a );
 a26640a <=( A234  and  A233 );
 a26643a <=( (not A298)  and  A236 );
 a26644a <=( a26643a  and  a26640a );
 a26647a <=( (not A300)  and  A299 );
 a26650a <=( (not A302)  and  (not A301) );
 a26651a <=( a26650a  and  a26647a );
 a26652a <=( a26651a  and  a26644a );
 a26656a <=( (not A167)  and  A168 );
 a26657a <=( (not A170)  and  a26656a );
 a26660a <=( (not A201)  and  A166 );
 a26663a <=( (not A232)  and  A203 );
 a26664a <=( a26663a  and  a26660a );
 a26665a <=( a26664a  and  a26657a );
 a26668a <=( A234  and  A233 );
 a26671a <=( (not A265)  and  A236 );
 a26672a <=( a26671a  and  a26668a );
 a26675a <=( (not A267)  and  A266 );
 a26678a <=( (not A269)  and  (not A268) );
 a26679a <=( a26678a  and  a26675a );
 a26680a <=( a26679a  and  a26672a );
 a26684a <=( (not A167)  and  A168 );
 a26685a <=( (not A170)  and  a26684a );
 a26688a <=( (not A201)  and  A166 );
 a26691a <=( (not A232)  and  A203 );
 a26692a <=( a26691a  and  a26688a );
 a26693a <=( a26692a  and  a26685a );
 a26696a <=( A234  and  A233 );
 a26699a <=( A265  and  A236 );
 a26700a <=( a26699a  and  a26696a );
 a26703a <=( (not A267)  and  (not A266) );
 a26706a <=( (not A269)  and  (not A268) );
 a26707a <=( a26706a  and  a26703a );
 a26708a <=( a26707a  and  a26700a );
 a26712a <=( (not A167)  and  A168 );
 a26713a <=( (not A170)  and  a26712a );
 a26716a <=( (not A201)  and  A166 );
 a26719a <=( (not A232)  and  A203 );
 a26720a <=( a26719a  and  a26716a );
 a26721a <=( a26720a  and  a26713a );
 a26724a <=( (not A234)  and  A233 );
 a26727a <=( (not A236)  and  (not A235) );
 a26728a <=( a26727a  and  a26724a );
 a26731a <=( (not A299)  and  A298 );
 a26734a <=( A301  and  A300 );
 a26735a <=( a26734a  and  a26731a );
 a26736a <=( a26735a  and  a26728a );
 a26740a <=( (not A167)  and  A168 );
 a26741a <=( (not A170)  and  a26740a );
 a26744a <=( (not A201)  and  A166 );
 a26747a <=( (not A232)  and  A203 );
 a26748a <=( a26747a  and  a26744a );
 a26749a <=( a26748a  and  a26741a );
 a26752a <=( (not A234)  and  A233 );
 a26755a <=( (not A236)  and  (not A235) );
 a26756a <=( a26755a  and  a26752a );
 a26759a <=( (not A299)  and  A298 );
 a26762a <=( A302  and  A300 );
 a26763a <=( a26762a  and  a26759a );
 a26764a <=( a26763a  and  a26756a );
 a26768a <=( (not A167)  and  A168 );
 a26769a <=( (not A170)  and  a26768a );
 a26772a <=( (not A201)  and  A166 );
 a26775a <=( (not A232)  and  A203 );
 a26776a <=( a26775a  and  a26772a );
 a26777a <=( a26776a  and  a26769a );
 a26780a <=( (not A234)  and  A233 );
 a26783a <=( (not A236)  and  (not A235) );
 a26784a <=( a26783a  and  a26780a );
 a26787a <=( A299  and  (not A298) );
 a26790a <=( A301  and  A300 );
 a26791a <=( a26790a  and  a26787a );
 a26792a <=( a26791a  and  a26784a );
 a26796a <=( (not A167)  and  A168 );
 a26797a <=( (not A170)  and  a26796a );
 a26800a <=( (not A201)  and  A166 );
 a26803a <=( (not A232)  and  A203 );
 a26804a <=( a26803a  and  a26800a );
 a26805a <=( a26804a  and  a26797a );
 a26808a <=( (not A234)  and  A233 );
 a26811a <=( (not A236)  and  (not A235) );
 a26812a <=( a26811a  and  a26808a );
 a26815a <=( A299  and  (not A298) );
 a26818a <=( A302  and  A300 );
 a26819a <=( a26818a  and  a26815a );
 a26820a <=( a26819a  and  a26812a );
 a26824a <=( (not A167)  and  A168 );
 a26825a <=( (not A170)  and  a26824a );
 a26828a <=( (not A201)  and  A166 );
 a26831a <=( (not A232)  and  A203 );
 a26832a <=( a26831a  and  a26828a );
 a26833a <=( a26832a  and  a26825a );
 a26836a <=( (not A234)  and  A233 );
 a26839a <=( (not A236)  and  (not A235) );
 a26840a <=( a26839a  and  a26836a );
 a26843a <=( A266  and  (not A265) );
 a26846a <=( A268  and  A267 );
 a26847a <=( a26846a  and  a26843a );
 a26848a <=( a26847a  and  a26840a );
 a26852a <=( (not A167)  and  A168 );
 a26853a <=( (not A170)  and  a26852a );
 a26856a <=( (not A201)  and  A166 );
 a26859a <=( (not A232)  and  A203 );
 a26860a <=( a26859a  and  a26856a );
 a26861a <=( a26860a  and  a26853a );
 a26864a <=( (not A234)  and  A233 );
 a26867a <=( (not A236)  and  (not A235) );
 a26868a <=( a26867a  and  a26864a );
 a26871a <=( A266  and  (not A265) );
 a26874a <=( A269  and  A267 );
 a26875a <=( a26874a  and  a26871a );
 a26876a <=( a26875a  and  a26868a );
 a26880a <=( (not A167)  and  A168 );
 a26881a <=( (not A170)  and  a26880a );
 a26884a <=( (not A201)  and  A166 );
 a26887a <=( (not A232)  and  A203 );
 a26888a <=( a26887a  and  a26884a );
 a26889a <=( a26888a  and  a26881a );
 a26892a <=( (not A234)  and  A233 );
 a26895a <=( (not A236)  and  (not A235) );
 a26896a <=( a26895a  and  a26892a );
 a26899a <=( (not A266)  and  A265 );
 a26902a <=( A268  and  A267 );
 a26903a <=( a26902a  and  a26899a );
 a26904a <=( a26903a  and  a26896a );
 a26908a <=( (not A167)  and  A168 );
 a26909a <=( (not A170)  and  a26908a );
 a26912a <=( (not A201)  and  A166 );
 a26915a <=( (not A232)  and  A203 );
 a26916a <=( a26915a  and  a26912a );
 a26917a <=( a26916a  and  a26909a );
 a26920a <=( (not A234)  and  A233 );
 a26923a <=( (not A236)  and  (not A235) );
 a26924a <=( a26923a  and  a26920a );
 a26927a <=( (not A266)  and  A265 );
 a26930a <=( A269  and  A267 );
 a26931a <=( a26930a  and  a26927a );
 a26932a <=( a26931a  and  a26924a );
 a26936a <=( (not A167)  and  A168 );
 a26937a <=( (not A170)  and  a26936a );
 a26940a <=( (not A201)  and  A166 );
 a26943a <=( A232  and  A203 );
 a26944a <=( a26943a  and  a26940a );
 a26945a <=( a26944a  and  a26937a );
 a26948a <=( A234  and  (not A233) );
 a26951a <=( A298  and  A235 );
 a26952a <=( a26951a  and  a26948a );
 a26955a <=( (not A300)  and  (not A299) );
 a26958a <=( (not A302)  and  (not A301) );
 a26959a <=( a26958a  and  a26955a );
 a26960a <=( a26959a  and  a26952a );
 a26964a <=( (not A167)  and  A168 );
 a26965a <=( (not A170)  and  a26964a );
 a26968a <=( (not A201)  and  A166 );
 a26971a <=( A232  and  A203 );
 a26972a <=( a26971a  and  a26968a );
 a26973a <=( a26972a  and  a26965a );
 a26976a <=( A234  and  (not A233) );
 a26979a <=( (not A298)  and  A235 );
 a26980a <=( a26979a  and  a26976a );
 a26983a <=( (not A300)  and  A299 );
 a26986a <=( (not A302)  and  (not A301) );
 a26987a <=( a26986a  and  a26983a );
 a26988a <=( a26987a  and  a26980a );
 a26992a <=( (not A167)  and  A168 );
 a26993a <=( (not A170)  and  a26992a );
 a26996a <=( (not A201)  and  A166 );
 a26999a <=( A232  and  A203 );
 a27000a <=( a26999a  and  a26996a );
 a27001a <=( a27000a  and  a26993a );
 a27004a <=( A234  and  (not A233) );
 a27007a <=( (not A265)  and  A235 );
 a27008a <=( a27007a  and  a27004a );
 a27011a <=( (not A267)  and  A266 );
 a27014a <=( (not A269)  and  (not A268) );
 a27015a <=( a27014a  and  a27011a );
 a27016a <=( a27015a  and  a27008a );
 a27020a <=( (not A167)  and  A168 );
 a27021a <=( (not A170)  and  a27020a );
 a27024a <=( (not A201)  and  A166 );
 a27027a <=( A232  and  A203 );
 a27028a <=( a27027a  and  a27024a );
 a27029a <=( a27028a  and  a27021a );
 a27032a <=( A234  and  (not A233) );
 a27035a <=( A265  and  A235 );
 a27036a <=( a27035a  and  a27032a );
 a27039a <=( (not A267)  and  (not A266) );
 a27042a <=( (not A269)  and  (not A268) );
 a27043a <=( a27042a  and  a27039a );
 a27044a <=( a27043a  and  a27036a );
 a27048a <=( (not A167)  and  A168 );
 a27049a <=( (not A170)  and  a27048a );
 a27052a <=( (not A201)  and  A166 );
 a27055a <=( A232  and  A203 );
 a27056a <=( a27055a  and  a27052a );
 a27057a <=( a27056a  and  a27049a );
 a27060a <=( A234  and  (not A233) );
 a27063a <=( A298  and  A236 );
 a27064a <=( a27063a  and  a27060a );
 a27067a <=( (not A300)  and  (not A299) );
 a27070a <=( (not A302)  and  (not A301) );
 a27071a <=( a27070a  and  a27067a );
 a27072a <=( a27071a  and  a27064a );
 a27076a <=( (not A167)  and  A168 );
 a27077a <=( (not A170)  and  a27076a );
 a27080a <=( (not A201)  and  A166 );
 a27083a <=( A232  and  A203 );
 a27084a <=( a27083a  and  a27080a );
 a27085a <=( a27084a  and  a27077a );
 a27088a <=( A234  and  (not A233) );
 a27091a <=( (not A298)  and  A236 );
 a27092a <=( a27091a  and  a27088a );
 a27095a <=( (not A300)  and  A299 );
 a27098a <=( (not A302)  and  (not A301) );
 a27099a <=( a27098a  and  a27095a );
 a27100a <=( a27099a  and  a27092a );
 a27104a <=( (not A167)  and  A168 );
 a27105a <=( (not A170)  and  a27104a );
 a27108a <=( (not A201)  and  A166 );
 a27111a <=( A232  and  A203 );
 a27112a <=( a27111a  and  a27108a );
 a27113a <=( a27112a  and  a27105a );
 a27116a <=( A234  and  (not A233) );
 a27119a <=( (not A265)  and  A236 );
 a27120a <=( a27119a  and  a27116a );
 a27123a <=( (not A267)  and  A266 );
 a27126a <=( (not A269)  and  (not A268) );
 a27127a <=( a27126a  and  a27123a );
 a27128a <=( a27127a  and  a27120a );
 a27132a <=( (not A167)  and  A168 );
 a27133a <=( (not A170)  and  a27132a );
 a27136a <=( (not A201)  and  A166 );
 a27139a <=( A232  and  A203 );
 a27140a <=( a27139a  and  a27136a );
 a27141a <=( a27140a  and  a27133a );
 a27144a <=( A234  and  (not A233) );
 a27147a <=( A265  and  A236 );
 a27148a <=( a27147a  and  a27144a );
 a27151a <=( (not A267)  and  (not A266) );
 a27154a <=( (not A269)  and  (not A268) );
 a27155a <=( a27154a  and  a27151a );
 a27156a <=( a27155a  and  a27148a );
 a27160a <=( (not A167)  and  A168 );
 a27161a <=( (not A170)  and  a27160a );
 a27164a <=( (not A201)  and  A166 );
 a27167a <=( A232  and  A203 );
 a27168a <=( a27167a  and  a27164a );
 a27169a <=( a27168a  and  a27161a );
 a27172a <=( (not A234)  and  (not A233) );
 a27175a <=( (not A236)  and  (not A235) );
 a27176a <=( a27175a  and  a27172a );
 a27179a <=( (not A299)  and  A298 );
 a27182a <=( A301  and  A300 );
 a27183a <=( a27182a  and  a27179a );
 a27184a <=( a27183a  and  a27176a );
 a27188a <=( (not A167)  and  A168 );
 a27189a <=( (not A170)  and  a27188a );
 a27192a <=( (not A201)  and  A166 );
 a27195a <=( A232  and  A203 );
 a27196a <=( a27195a  and  a27192a );
 a27197a <=( a27196a  and  a27189a );
 a27200a <=( (not A234)  and  (not A233) );
 a27203a <=( (not A236)  and  (not A235) );
 a27204a <=( a27203a  and  a27200a );
 a27207a <=( (not A299)  and  A298 );
 a27210a <=( A302  and  A300 );
 a27211a <=( a27210a  and  a27207a );
 a27212a <=( a27211a  and  a27204a );
 a27216a <=( (not A167)  and  A168 );
 a27217a <=( (not A170)  and  a27216a );
 a27220a <=( (not A201)  and  A166 );
 a27223a <=( A232  and  A203 );
 a27224a <=( a27223a  and  a27220a );
 a27225a <=( a27224a  and  a27217a );
 a27228a <=( (not A234)  and  (not A233) );
 a27231a <=( (not A236)  and  (not A235) );
 a27232a <=( a27231a  and  a27228a );
 a27235a <=( A299  and  (not A298) );
 a27238a <=( A301  and  A300 );
 a27239a <=( a27238a  and  a27235a );
 a27240a <=( a27239a  and  a27232a );
 a27244a <=( (not A167)  and  A168 );
 a27245a <=( (not A170)  and  a27244a );
 a27248a <=( (not A201)  and  A166 );
 a27251a <=( A232  and  A203 );
 a27252a <=( a27251a  and  a27248a );
 a27253a <=( a27252a  and  a27245a );
 a27256a <=( (not A234)  and  (not A233) );
 a27259a <=( (not A236)  and  (not A235) );
 a27260a <=( a27259a  and  a27256a );
 a27263a <=( A299  and  (not A298) );
 a27266a <=( A302  and  A300 );
 a27267a <=( a27266a  and  a27263a );
 a27268a <=( a27267a  and  a27260a );
 a27272a <=( (not A167)  and  A168 );
 a27273a <=( (not A170)  and  a27272a );
 a27276a <=( (not A201)  and  A166 );
 a27279a <=( A232  and  A203 );
 a27280a <=( a27279a  and  a27276a );
 a27281a <=( a27280a  and  a27273a );
 a27284a <=( (not A234)  and  (not A233) );
 a27287a <=( (not A236)  and  (not A235) );
 a27288a <=( a27287a  and  a27284a );
 a27291a <=( A266  and  (not A265) );
 a27294a <=( A268  and  A267 );
 a27295a <=( a27294a  and  a27291a );
 a27296a <=( a27295a  and  a27288a );
 a27300a <=( (not A167)  and  A168 );
 a27301a <=( (not A170)  and  a27300a );
 a27304a <=( (not A201)  and  A166 );
 a27307a <=( A232  and  A203 );
 a27308a <=( a27307a  and  a27304a );
 a27309a <=( a27308a  and  a27301a );
 a27312a <=( (not A234)  and  (not A233) );
 a27315a <=( (not A236)  and  (not A235) );
 a27316a <=( a27315a  and  a27312a );
 a27319a <=( A266  and  (not A265) );
 a27322a <=( A269  and  A267 );
 a27323a <=( a27322a  and  a27319a );
 a27324a <=( a27323a  and  a27316a );
 a27328a <=( (not A167)  and  A168 );
 a27329a <=( (not A170)  and  a27328a );
 a27332a <=( (not A201)  and  A166 );
 a27335a <=( A232  and  A203 );
 a27336a <=( a27335a  and  a27332a );
 a27337a <=( a27336a  and  a27329a );
 a27340a <=( (not A234)  and  (not A233) );
 a27343a <=( (not A236)  and  (not A235) );
 a27344a <=( a27343a  and  a27340a );
 a27347a <=( (not A266)  and  A265 );
 a27350a <=( A268  and  A267 );
 a27351a <=( a27350a  and  a27347a );
 a27352a <=( a27351a  and  a27344a );
 a27356a <=( (not A167)  and  A168 );
 a27357a <=( (not A170)  and  a27356a );
 a27360a <=( (not A201)  and  A166 );
 a27363a <=( A232  and  A203 );
 a27364a <=( a27363a  and  a27360a );
 a27365a <=( a27364a  and  a27357a );
 a27368a <=( (not A234)  and  (not A233) );
 a27371a <=( (not A236)  and  (not A235) );
 a27372a <=( a27371a  and  a27368a );
 a27375a <=( (not A266)  and  A265 );
 a27378a <=( A269  and  A267 );
 a27379a <=( a27378a  and  a27375a );
 a27380a <=( a27379a  and  a27372a );
 a27384a <=( (not A167)  and  A168 );
 a27385a <=( (not A170)  and  a27384a );
 a27388a <=( A199  and  A166 );
 a27391a <=( (not A232)  and  A200 );
 a27392a <=( a27391a  and  a27388a );
 a27393a <=( a27392a  and  a27385a );
 a27396a <=( A234  and  A233 );
 a27399a <=( A298  and  A235 );
 a27400a <=( a27399a  and  a27396a );
 a27403a <=( (not A300)  and  (not A299) );
 a27406a <=( (not A302)  and  (not A301) );
 a27407a <=( a27406a  and  a27403a );
 a27408a <=( a27407a  and  a27400a );
 a27412a <=( (not A167)  and  A168 );
 a27413a <=( (not A170)  and  a27412a );
 a27416a <=( A199  and  A166 );
 a27419a <=( (not A232)  and  A200 );
 a27420a <=( a27419a  and  a27416a );
 a27421a <=( a27420a  and  a27413a );
 a27424a <=( A234  and  A233 );
 a27427a <=( (not A298)  and  A235 );
 a27428a <=( a27427a  and  a27424a );
 a27431a <=( (not A300)  and  A299 );
 a27434a <=( (not A302)  and  (not A301) );
 a27435a <=( a27434a  and  a27431a );
 a27436a <=( a27435a  and  a27428a );
 a27440a <=( (not A167)  and  A168 );
 a27441a <=( (not A170)  and  a27440a );
 a27444a <=( A199  and  A166 );
 a27447a <=( (not A232)  and  A200 );
 a27448a <=( a27447a  and  a27444a );
 a27449a <=( a27448a  and  a27441a );
 a27452a <=( A234  and  A233 );
 a27455a <=( (not A265)  and  A235 );
 a27456a <=( a27455a  and  a27452a );
 a27459a <=( (not A267)  and  A266 );
 a27462a <=( (not A269)  and  (not A268) );
 a27463a <=( a27462a  and  a27459a );
 a27464a <=( a27463a  and  a27456a );
 a27468a <=( (not A167)  and  A168 );
 a27469a <=( (not A170)  and  a27468a );
 a27472a <=( A199  and  A166 );
 a27475a <=( (not A232)  and  A200 );
 a27476a <=( a27475a  and  a27472a );
 a27477a <=( a27476a  and  a27469a );
 a27480a <=( A234  and  A233 );
 a27483a <=( A265  and  A235 );
 a27484a <=( a27483a  and  a27480a );
 a27487a <=( (not A267)  and  (not A266) );
 a27490a <=( (not A269)  and  (not A268) );
 a27491a <=( a27490a  and  a27487a );
 a27492a <=( a27491a  and  a27484a );
 a27496a <=( (not A167)  and  A168 );
 a27497a <=( (not A170)  and  a27496a );
 a27500a <=( A199  and  A166 );
 a27503a <=( (not A232)  and  A200 );
 a27504a <=( a27503a  and  a27500a );
 a27505a <=( a27504a  and  a27497a );
 a27508a <=( A234  and  A233 );
 a27511a <=( A298  and  A236 );
 a27512a <=( a27511a  and  a27508a );
 a27515a <=( (not A300)  and  (not A299) );
 a27518a <=( (not A302)  and  (not A301) );
 a27519a <=( a27518a  and  a27515a );
 a27520a <=( a27519a  and  a27512a );
 a27524a <=( (not A167)  and  A168 );
 a27525a <=( (not A170)  and  a27524a );
 a27528a <=( A199  and  A166 );
 a27531a <=( (not A232)  and  A200 );
 a27532a <=( a27531a  and  a27528a );
 a27533a <=( a27532a  and  a27525a );
 a27536a <=( A234  and  A233 );
 a27539a <=( (not A298)  and  A236 );
 a27540a <=( a27539a  and  a27536a );
 a27543a <=( (not A300)  and  A299 );
 a27546a <=( (not A302)  and  (not A301) );
 a27547a <=( a27546a  and  a27543a );
 a27548a <=( a27547a  and  a27540a );
 a27552a <=( (not A167)  and  A168 );
 a27553a <=( (not A170)  and  a27552a );
 a27556a <=( A199  and  A166 );
 a27559a <=( (not A232)  and  A200 );
 a27560a <=( a27559a  and  a27556a );
 a27561a <=( a27560a  and  a27553a );
 a27564a <=( A234  and  A233 );
 a27567a <=( (not A265)  and  A236 );
 a27568a <=( a27567a  and  a27564a );
 a27571a <=( (not A267)  and  A266 );
 a27574a <=( (not A269)  and  (not A268) );
 a27575a <=( a27574a  and  a27571a );
 a27576a <=( a27575a  and  a27568a );
 a27580a <=( (not A167)  and  A168 );
 a27581a <=( (not A170)  and  a27580a );
 a27584a <=( A199  and  A166 );
 a27587a <=( (not A232)  and  A200 );
 a27588a <=( a27587a  and  a27584a );
 a27589a <=( a27588a  and  a27581a );
 a27592a <=( A234  and  A233 );
 a27595a <=( A265  and  A236 );
 a27596a <=( a27595a  and  a27592a );
 a27599a <=( (not A267)  and  (not A266) );
 a27602a <=( (not A269)  and  (not A268) );
 a27603a <=( a27602a  and  a27599a );
 a27604a <=( a27603a  and  a27596a );
 a27608a <=( (not A167)  and  A168 );
 a27609a <=( (not A170)  and  a27608a );
 a27612a <=( A199  and  A166 );
 a27615a <=( (not A232)  and  A200 );
 a27616a <=( a27615a  and  a27612a );
 a27617a <=( a27616a  and  a27609a );
 a27620a <=( (not A234)  and  A233 );
 a27623a <=( (not A236)  and  (not A235) );
 a27624a <=( a27623a  and  a27620a );
 a27627a <=( (not A299)  and  A298 );
 a27630a <=( A301  and  A300 );
 a27631a <=( a27630a  and  a27627a );
 a27632a <=( a27631a  and  a27624a );
 a27636a <=( (not A167)  and  A168 );
 a27637a <=( (not A170)  and  a27636a );
 a27640a <=( A199  and  A166 );
 a27643a <=( (not A232)  and  A200 );
 a27644a <=( a27643a  and  a27640a );
 a27645a <=( a27644a  and  a27637a );
 a27648a <=( (not A234)  and  A233 );
 a27651a <=( (not A236)  and  (not A235) );
 a27652a <=( a27651a  and  a27648a );
 a27655a <=( (not A299)  and  A298 );
 a27658a <=( A302  and  A300 );
 a27659a <=( a27658a  and  a27655a );
 a27660a <=( a27659a  and  a27652a );
 a27664a <=( (not A167)  and  A168 );
 a27665a <=( (not A170)  and  a27664a );
 a27668a <=( A199  and  A166 );
 a27671a <=( (not A232)  and  A200 );
 a27672a <=( a27671a  and  a27668a );
 a27673a <=( a27672a  and  a27665a );
 a27676a <=( (not A234)  and  A233 );
 a27679a <=( (not A236)  and  (not A235) );
 a27680a <=( a27679a  and  a27676a );
 a27683a <=( A299  and  (not A298) );
 a27686a <=( A301  and  A300 );
 a27687a <=( a27686a  and  a27683a );
 a27688a <=( a27687a  and  a27680a );
 a27692a <=( (not A167)  and  A168 );
 a27693a <=( (not A170)  and  a27692a );
 a27696a <=( A199  and  A166 );
 a27699a <=( (not A232)  and  A200 );
 a27700a <=( a27699a  and  a27696a );
 a27701a <=( a27700a  and  a27693a );
 a27704a <=( (not A234)  and  A233 );
 a27707a <=( (not A236)  and  (not A235) );
 a27708a <=( a27707a  and  a27704a );
 a27711a <=( A299  and  (not A298) );
 a27714a <=( A302  and  A300 );
 a27715a <=( a27714a  and  a27711a );
 a27716a <=( a27715a  and  a27708a );
 a27720a <=( (not A167)  and  A168 );
 a27721a <=( (not A170)  and  a27720a );
 a27724a <=( A199  and  A166 );
 a27727a <=( (not A232)  and  A200 );
 a27728a <=( a27727a  and  a27724a );
 a27729a <=( a27728a  and  a27721a );
 a27732a <=( (not A234)  and  A233 );
 a27735a <=( (not A236)  and  (not A235) );
 a27736a <=( a27735a  and  a27732a );
 a27739a <=( A266  and  (not A265) );
 a27742a <=( A268  and  A267 );
 a27743a <=( a27742a  and  a27739a );
 a27744a <=( a27743a  and  a27736a );
 a27748a <=( (not A167)  and  A168 );
 a27749a <=( (not A170)  and  a27748a );
 a27752a <=( A199  and  A166 );
 a27755a <=( (not A232)  and  A200 );
 a27756a <=( a27755a  and  a27752a );
 a27757a <=( a27756a  and  a27749a );
 a27760a <=( (not A234)  and  A233 );
 a27763a <=( (not A236)  and  (not A235) );
 a27764a <=( a27763a  and  a27760a );
 a27767a <=( A266  and  (not A265) );
 a27770a <=( A269  and  A267 );
 a27771a <=( a27770a  and  a27767a );
 a27772a <=( a27771a  and  a27764a );
 a27776a <=( (not A167)  and  A168 );
 a27777a <=( (not A170)  and  a27776a );
 a27780a <=( A199  and  A166 );
 a27783a <=( (not A232)  and  A200 );
 a27784a <=( a27783a  and  a27780a );
 a27785a <=( a27784a  and  a27777a );
 a27788a <=( (not A234)  and  A233 );
 a27791a <=( (not A236)  and  (not A235) );
 a27792a <=( a27791a  and  a27788a );
 a27795a <=( (not A266)  and  A265 );
 a27798a <=( A268  and  A267 );
 a27799a <=( a27798a  and  a27795a );
 a27800a <=( a27799a  and  a27792a );
 a27804a <=( (not A167)  and  A168 );
 a27805a <=( (not A170)  and  a27804a );
 a27808a <=( A199  and  A166 );
 a27811a <=( (not A232)  and  A200 );
 a27812a <=( a27811a  and  a27808a );
 a27813a <=( a27812a  and  a27805a );
 a27816a <=( (not A234)  and  A233 );
 a27819a <=( (not A236)  and  (not A235) );
 a27820a <=( a27819a  and  a27816a );
 a27823a <=( (not A266)  and  A265 );
 a27826a <=( A269  and  A267 );
 a27827a <=( a27826a  and  a27823a );
 a27828a <=( a27827a  and  a27820a );
 a27832a <=( (not A167)  and  A168 );
 a27833a <=( (not A170)  and  a27832a );
 a27836a <=( A199  and  A166 );
 a27839a <=( A232  and  A200 );
 a27840a <=( a27839a  and  a27836a );
 a27841a <=( a27840a  and  a27833a );
 a27844a <=( A234  and  (not A233) );
 a27847a <=( A298  and  A235 );
 a27848a <=( a27847a  and  a27844a );
 a27851a <=( (not A300)  and  (not A299) );
 a27854a <=( (not A302)  and  (not A301) );
 a27855a <=( a27854a  and  a27851a );
 a27856a <=( a27855a  and  a27848a );
 a27860a <=( (not A167)  and  A168 );
 a27861a <=( (not A170)  and  a27860a );
 a27864a <=( A199  and  A166 );
 a27867a <=( A232  and  A200 );
 a27868a <=( a27867a  and  a27864a );
 a27869a <=( a27868a  and  a27861a );
 a27872a <=( A234  and  (not A233) );
 a27875a <=( (not A298)  and  A235 );
 a27876a <=( a27875a  and  a27872a );
 a27879a <=( (not A300)  and  A299 );
 a27882a <=( (not A302)  and  (not A301) );
 a27883a <=( a27882a  and  a27879a );
 a27884a <=( a27883a  and  a27876a );
 a27888a <=( (not A167)  and  A168 );
 a27889a <=( (not A170)  and  a27888a );
 a27892a <=( A199  and  A166 );
 a27895a <=( A232  and  A200 );
 a27896a <=( a27895a  and  a27892a );
 a27897a <=( a27896a  and  a27889a );
 a27900a <=( A234  and  (not A233) );
 a27903a <=( (not A265)  and  A235 );
 a27904a <=( a27903a  and  a27900a );
 a27907a <=( (not A267)  and  A266 );
 a27910a <=( (not A269)  and  (not A268) );
 a27911a <=( a27910a  and  a27907a );
 a27912a <=( a27911a  and  a27904a );
 a27916a <=( (not A167)  and  A168 );
 a27917a <=( (not A170)  and  a27916a );
 a27920a <=( A199  and  A166 );
 a27923a <=( A232  and  A200 );
 a27924a <=( a27923a  and  a27920a );
 a27925a <=( a27924a  and  a27917a );
 a27928a <=( A234  and  (not A233) );
 a27931a <=( A265  and  A235 );
 a27932a <=( a27931a  and  a27928a );
 a27935a <=( (not A267)  and  (not A266) );
 a27938a <=( (not A269)  and  (not A268) );
 a27939a <=( a27938a  and  a27935a );
 a27940a <=( a27939a  and  a27932a );
 a27944a <=( (not A167)  and  A168 );
 a27945a <=( (not A170)  and  a27944a );
 a27948a <=( A199  and  A166 );
 a27951a <=( A232  and  A200 );
 a27952a <=( a27951a  and  a27948a );
 a27953a <=( a27952a  and  a27945a );
 a27956a <=( A234  and  (not A233) );
 a27959a <=( A298  and  A236 );
 a27960a <=( a27959a  and  a27956a );
 a27963a <=( (not A300)  and  (not A299) );
 a27966a <=( (not A302)  and  (not A301) );
 a27967a <=( a27966a  and  a27963a );
 a27968a <=( a27967a  and  a27960a );
 a27972a <=( (not A167)  and  A168 );
 a27973a <=( (not A170)  and  a27972a );
 a27976a <=( A199  and  A166 );
 a27979a <=( A232  and  A200 );
 a27980a <=( a27979a  and  a27976a );
 a27981a <=( a27980a  and  a27973a );
 a27984a <=( A234  and  (not A233) );
 a27987a <=( (not A298)  and  A236 );
 a27988a <=( a27987a  and  a27984a );
 a27991a <=( (not A300)  and  A299 );
 a27994a <=( (not A302)  and  (not A301) );
 a27995a <=( a27994a  and  a27991a );
 a27996a <=( a27995a  and  a27988a );
 a28000a <=( (not A167)  and  A168 );
 a28001a <=( (not A170)  and  a28000a );
 a28004a <=( A199  and  A166 );
 a28007a <=( A232  and  A200 );
 a28008a <=( a28007a  and  a28004a );
 a28009a <=( a28008a  and  a28001a );
 a28012a <=( A234  and  (not A233) );
 a28015a <=( (not A265)  and  A236 );
 a28016a <=( a28015a  and  a28012a );
 a28019a <=( (not A267)  and  A266 );
 a28022a <=( (not A269)  and  (not A268) );
 a28023a <=( a28022a  and  a28019a );
 a28024a <=( a28023a  and  a28016a );
 a28028a <=( (not A167)  and  A168 );
 a28029a <=( (not A170)  and  a28028a );
 a28032a <=( A199  and  A166 );
 a28035a <=( A232  and  A200 );
 a28036a <=( a28035a  and  a28032a );
 a28037a <=( a28036a  and  a28029a );
 a28040a <=( A234  and  (not A233) );
 a28043a <=( A265  and  A236 );
 a28044a <=( a28043a  and  a28040a );
 a28047a <=( (not A267)  and  (not A266) );
 a28050a <=( (not A269)  and  (not A268) );
 a28051a <=( a28050a  and  a28047a );
 a28052a <=( a28051a  and  a28044a );
 a28056a <=( (not A167)  and  A168 );
 a28057a <=( (not A170)  and  a28056a );
 a28060a <=( A199  and  A166 );
 a28063a <=( A232  and  A200 );
 a28064a <=( a28063a  and  a28060a );
 a28065a <=( a28064a  and  a28057a );
 a28068a <=( (not A234)  and  (not A233) );
 a28071a <=( (not A236)  and  (not A235) );
 a28072a <=( a28071a  and  a28068a );
 a28075a <=( (not A299)  and  A298 );
 a28078a <=( A301  and  A300 );
 a28079a <=( a28078a  and  a28075a );
 a28080a <=( a28079a  and  a28072a );
 a28084a <=( (not A167)  and  A168 );
 a28085a <=( (not A170)  and  a28084a );
 a28088a <=( A199  and  A166 );
 a28091a <=( A232  and  A200 );
 a28092a <=( a28091a  and  a28088a );
 a28093a <=( a28092a  and  a28085a );
 a28096a <=( (not A234)  and  (not A233) );
 a28099a <=( (not A236)  and  (not A235) );
 a28100a <=( a28099a  and  a28096a );
 a28103a <=( (not A299)  and  A298 );
 a28106a <=( A302  and  A300 );
 a28107a <=( a28106a  and  a28103a );
 a28108a <=( a28107a  and  a28100a );
 a28112a <=( (not A167)  and  A168 );
 a28113a <=( (not A170)  and  a28112a );
 a28116a <=( A199  and  A166 );
 a28119a <=( A232  and  A200 );
 a28120a <=( a28119a  and  a28116a );
 a28121a <=( a28120a  and  a28113a );
 a28124a <=( (not A234)  and  (not A233) );
 a28127a <=( (not A236)  and  (not A235) );
 a28128a <=( a28127a  and  a28124a );
 a28131a <=( A299  and  (not A298) );
 a28134a <=( A301  and  A300 );
 a28135a <=( a28134a  and  a28131a );
 a28136a <=( a28135a  and  a28128a );
 a28140a <=( (not A167)  and  A168 );
 a28141a <=( (not A170)  and  a28140a );
 a28144a <=( A199  and  A166 );
 a28147a <=( A232  and  A200 );
 a28148a <=( a28147a  and  a28144a );
 a28149a <=( a28148a  and  a28141a );
 a28152a <=( (not A234)  and  (not A233) );
 a28155a <=( (not A236)  and  (not A235) );
 a28156a <=( a28155a  and  a28152a );
 a28159a <=( A299  and  (not A298) );
 a28162a <=( A302  and  A300 );
 a28163a <=( a28162a  and  a28159a );
 a28164a <=( a28163a  and  a28156a );
 a28168a <=( (not A167)  and  A168 );
 a28169a <=( (not A170)  and  a28168a );
 a28172a <=( A199  and  A166 );
 a28175a <=( A232  and  A200 );
 a28176a <=( a28175a  and  a28172a );
 a28177a <=( a28176a  and  a28169a );
 a28180a <=( (not A234)  and  (not A233) );
 a28183a <=( (not A236)  and  (not A235) );
 a28184a <=( a28183a  and  a28180a );
 a28187a <=( A266  and  (not A265) );
 a28190a <=( A268  and  A267 );
 a28191a <=( a28190a  and  a28187a );
 a28192a <=( a28191a  and  a28184a );
 a28196a <=( (not A167)  and  A168 );
 a28197a <=( (not A170)  and  a28196a );
 a28200a <=( A199  and  A166 );
 a28203a <=( A232  and  A200 );
 a28204a <=( a28203a  and  a28200a );
 a28205a <=( a28204a  and  a28197a );
 a28208a <=( (not A234)  and  (not A233) );
 a28211a <=( (not A236)  and  (not A235) );
 a28212a <=( a28211a  and  a28208a );
 a28215a <=( A266  and  (not A265) );
 a28218a <=( A269  and  A267 );
 a28219a <=( a28218a  and  a28215a );
 a28220a <=( a28219a  and  a28212a );
 a28224a <=( (not A167)  and  A168 );
 a28225a <=( (not A170)  and  a28224a );
 a28228a <=( A199  and  A166 );
 a28231a <=( A232  and  A200 );
 a28232a <=( a28231a  and  a28228a );
 a28233a <=( a28232a  and  a28225a );
 a28236a <=( (not A234)  and  (not A233) );
 a28239a <=( (not A236)  and  (not A235) );
 a28240a <=( a28239a  and  a28236a );
 a28243a <=( (not A266)  and  A265 );
 a28246a <=( A268  and  A267 );
 a28247a <=( a28246a  and  a28243a );
 a28248a <=( a28247a  and  a28240a );
 a28252a <=( (not A167)  and  A168 );
 a28253a <=( (not A170)  and  a28252a );
 a28256a <=( A199  and  A166 );
 a28259a <=( A232  and  A200 );
 a28260a <=( a28259a  and  a28256a );
 a28261a <=( a28260a  and  a28253a );
 a28264a <=( (not A234)  and  (not A233) );
 a28267a <=( (not A236)  and  (not A235) );
 a28268a <=( a28267a  and  a28264a );
 a28271a <=( (not A266)  and  A265 );
 a28274a <=( A269  and  A267 );
 a28275a <=( a28274a  and  a28271a );
 a28276a <=( a28275a  and  a28268a );
 a28280a <=( (not A167)  and  A168 );
 a28281a <=( (not A170)  and  a28280a );
 a28284a <=( (not A199)  and  A166 );
 a28287a <=( (not A232)  and  (not A200) );
 a28288a <=( a28287a  and  a28284a );
 a28289a <=( a28288a  and  a28281a );
 a28292a <=( A234  and  A233 );
 a28295a <=( A298  and  A235 );
 a28296a <=( a28295a  and  a28292a );
 a28299a <=( (not A300)  and  (not A299) );
 a28302a <=( (not A302)  and  (not A301) );
 a28303a <=( a28302a  and  a28299a );
 a28304a <=( a28303a  and  a28296a );
 a28308a <=( (not A167)  and  A168 );
 a28309a <=( (not A170)  and  a28308a );
 a28312a <=( (not A199)  and  A166 );
 a28315a <=( (not A232)  and  (not A200) );
 a28316a <=( a28315a  and  a28312a );
 a28317a <=( a28316a  and  a28309a );
 a28320a <=( A234  and  A233 );
 a28323a <=( (not A298)  and  A235 );
 a28324a <=( a28323a  and  a28320a );
 a28327a <=( (not A300)  and  A299 );
 a28330a <=( (not A302)  and  (not A301) );
 a28331a <=( a28330a  and  a28327a );
 a28332a <=( a28331a  and  a28324a );
 a28336a <=( (not A167)  and  A168 );
 a28337a <=( (not A170)  and  a28336a );
 a28340a <=( (not A199)  and  A166 );
 a28343a <=( (not A232)  and  (not A200) );
 a28344a <=( a28343a  and  a28340a );
 a28345a <=( a28344a  and  a28337a );
 a28348a <=( A234  and  A233 );
 a28351a <=( (not A265)  and  A235 );
 a28352a <=( a28351a  and  a28348a );
 a28355a <=( (not A267)  and  A266 );
 a28358a <=( (not A269)  and  (not A268) );
 a28359a <=( a28358a  and  a28355a );
 a28360a <=( a28359a  and  a28352a );
 a28364a <=( (not A167)  and  A168 );
 a28365a <=( (not A170)  and  a28364a );
 a28368a <=( (not A199)  and  A166 );
 a28371a <=( (not A232)  and  (not A200) );
 a28372a <=( a28371a  and  a28368a );
 a28373a <=( a28372a  and  a28365a );
 a28376a <=( A234  and  A233 );
 a28379a <=( A265  and  A235 );
 a28380a <=( a28379a  and  a28376a );
 a28383a <=( (not A267)  and  (not A266) );
 a28386a <=( (not A269)  and  (not A268) );
 a28387a <=( a28386a  and  a28383a );
 a28388a <=( a28387a  and  a28380a );
 a28392a <=( (not A167)  and  A168 );
 a28393a <=( (not A170)  and  a28392a );
 a28396a <=( (not A199)  and  A166 );
 a28399a <=( (not A232)  and  (not A200) );
 a28400a <=( a28399a  and  a28396a );
 a28401a <=( a28400a  and  a28393a );
 a28404a <=( A234  and  A233 );
 a28407a <=( A298  and  A236 );
 a28408a <=( a28407a  and  a28404a );
 a28411a <=( (not A300)  and  (not A299) );
 a28414a <=( (not A302)  and  (not A301) );
 a28415a <=( a28414a  and  a28411a );
 a28416a <=( a28415a  and  a28408a );
 a28420a <=( (not A167)  and  A168 );
 a28421a <=( (not A170)  and  a28420a );
 a28424a <=( (not A199)  and  A166 );
 a28427a <=( (not A232)  and  (not A200) );
 a28428a <=( a28427a  and  a28424a );
 a28429a <=( a28428a  and  a28421a );
 a28432a <=( A234  and  A233 );
 a28435a <=( (not A298)  and  A236 );
 a28436a <=( a28435a  and  a28432a );
 a28439a <=( (not A300)  and  A299 );
 a28442a <=( (not A302)  and  (not A301) );
 a28443a <=( a28442a  and  a28439a );
 a28444a <=( a28443a  and  a28436a );
 a28448a <=( (not A167)  and  A168 );
 a28449a <=( (not A170)  and  a28448a );
 a28452a <=( (not A199)  and  A166 );
 a28455a <=( (not A232)  and  (not A200) );
 a28456a <=( a28455a  and  a28452a );
 a28457a <=( a28456a  and  a28449a );
 a28460a <=( A234  and  A233 );
 a28463a <=( (not A265)  and  A236 );
 a28464a <=( a28463a  and  a28460a );
 a28467a <=( (not A267)  and  A266 );
 a28470a <=( (not A269)  and  (not A268) );
 a28471a <=( a28470a  and  a28467a );
 a28472a <=( a28471a  and  a28464a );
 a28476a <=( (not A167)  and  A168 );
 a28477a <=( (not A170)  and  a28476a );
 a28480a <=( (not A199)  and  A166 );
 a28483a <=( (not A232)  and  (not A200) );
 a28484a <=( a28483a  and  a28480a );
 a28485a <=( a28484a  and  a28477a );
 a28488a <=( A234  and  A233 );
 a28491a <=( A265  and  A236 );
 a28492a <=( a28491a  and  a28488a );
 a28495a <=( (not A267)  and  (not A266) );
 a28498a <=( (not A269)  and  (not A268) );
 a28499a <=( a28498a  and  a28495a );
 a28500a <=( a28499a  and  a28492a );
 a28504a <=( (not A167)  and  A168 );
 a28505a <=( (not A170)  and  a28504a );
 a28508a <=( (not A199)  and  A166 );
 a28511a <=( (not A232)  and  (not A200) );
 a28512a <=( a28511a  and  a28508a );
 a28513a <=( a28512a  and  a28505a );
 a28516a <=( (not A234)  and  A233 );
 a28519a <=( (not A236)  and  (not A235) );
 a28520a <=( a28519a  and  a28516a );
 a28523a <=( (not A299)  and  A298 );
 a28526a <=( A301  and  A300 );
 a28527a <=( a28526a  and  a28523a );
 a28528a <=( a28527a  and  a28520a );
 a28532a <=( (not A167)  and  A168 );
 a28533a <=( (not A170)  and  a28532a );
 a28536a <=( (not A199)  and  A166 );
 a28539a <=( (not A232)  and  (not A200) );
 a28540a <=( a28539a  and  a28536a );
 a28541a <=( a28540a  and  a28533a );
 a28544a <=( (not A234)  and  A233 );
 a28547a <=( (not A236)  and  (not A235) );
 a28548a <=( a28547a  and  a28544a );
 a28551a <=( (not A299)  and  A298 );
 a28554a <=( A302  and  A300 );
 a28555a <=( a28554a  and  a28551a );
 a28556a <=( a28555a  and  a28548a );
 a28560a <=( (not A167)  and  A168 );
 a28561a <=( (not A170)  and  a28560a );
 a28564a <=( (not A199)  and  A166 );
 a28567a <=( (not A232)  and  (not A200) );
 a28568a <=( a28567a  and  a28564a );
 a28569a <=( a28568a  and  a28561a );
 a28572a <=( (not A234)  and  A233 );
 a28575a <=( (not A236)  and  (not A235) );
 a28576a <=( a28575a  and  a28572a );
 a28579a <=( A299  and  (not A298) );
 a28582a <=( A301  and  A300 );
 a28583a <=( a28582a  and  a28579a );
 a28584a <=( a28583a  and  a28576a );
 a28588a <=( (not A167)  and  A168 );
 a28589a <=( (not A170)  and  a28588a );
 a28592a <=( (not A199)  and  A166 );
 a28595a <=( (not A232)  and  (not A200) );
 a28596a <=( a28595a  and  a28592a );
 a28597a <=( a28596a  and  a28589a );
 a28600a <=( (not A234)  and  A233 );
 a28603a <=( (not A236)  and  (not A235) );
 a28604a <=( a28603a  and  a28600a );
 a28607a <=( A299  and  (not A298) );
 a28610a <=( A302  and  A300 );
 a28611a <=( a28610a  and  a28607a );
 a28612a <=( a28611a  and  a28604a );
 a28616a <=( (not A167)  and  A168 );
 a28617a <=( (not A170)  and  a28616a );
 a28620a <=( (not A199)  and  A166 );
 a28623a <=( (not A232)  and  (not A200) );
 a28624a <=( a28623a  and  a28620a );
 a28625a <=( a28624a  and  a28617a );
 a28628a <=( (not A234)  and  A233 );
 a28631a <=( (not A236)  and  (not A235) );
 a28632a <=( a28631a  and  a28628a );
 a28635a <=( A266  and  (not A265) );
 a28638a <=( A268  and  A267 );
 a28639a <=( a28638a  and  a28635a );
 a28640a <=( a28639a  and  a28632a );
 a28644a <=( (not A167)  and  A168 );
 a28645a <=( (not A170)  and  a28644a );
 a28648a <=( (not A199)  and  A166 );
 a28651a <=( (not A232)  and  (not A200) );
 a28652a <=( a28651a  and  a28648a );
 a28653a <=( a28652a  and  a28645a );
 a28656a <=( (not A234)  and  A233 );
 a28659a <=( (not A236)  and  (not A235) );
 a28660a <=( a28659a  and  a28656a );
 a28663a <=( A266  and  (not A265) );
 a28666a <=( A269  and  A267 );
 a28667a <=( a28666a  and  a28663a );
 a28668a <=( a28667a  and  a28660a );
 a28672a <=( (not A167)  and  A168 );
 a28673a <=( (not A170)  and  a28672a );
 a28676a <=( (not A199)  and  A166 );
 a28679a <=( (not A232)  and  (not A200) );
 a28680a <=( a28679a  and  a28676a );
 a28681a <=( a28680a  and  a28673a );
 a28684a <=( (not A234)  and  A233 );
 a28687a <=( (not A236)  and  (not A235) );
 a28688a <=( a28687a  and  a28684a );
 a28691a <=( (not A266)  and  A265 );
 a28694a <=( A268  and  A267 );
 a28695a <=( a28694a  and  a28691a );
 a28696a <=( a28695a  and  a28688a );
 a28700a <=( (not A167)  and  A168 );
 a28701a <=( (not A170)  and  a28700a );
 a28704a <=( (not A199)  and  A166 );
 a28707a <=( (not A232)  and  (not A200) );
 a28708a <=( a28707a  and  a28704a );
 a28709a <=( a28708a  and  a28701a );
 a28712a <=( (not A234)  and  A233 );
 a28715a <=( (not A236)  and  (not A235) );
 a28716a <=( a28715a  and  a28712a );
 a28719a <=( (not A266)  and  A265 );
 a28722a <=( A269  and  A267 );
 a28723a <=( a28722a  and  a28719a );
 a28724a <=( a28723a  and  a28716a );
 a28728a <=( (not A167)  and  A168 );
 a28729a <=( (not A170)  and  a28728a );
 a28732a <=( (not A199)  and  A166 );
 a28735a <=( A232  and  (not A200) );
 a28736a <=( a28735a  and  a28732a );
 a28737a <=( a28736a  and  a28729a );
 a28740a <=( A234  and  (not A233) );
 a28743a <=( A298  and  A235 );
 a28744a <=( a28743a  and  a28740a );
 a28747a <=( (not A300)  and  (not A299) );
 a28750a <=( (not A302)  and  (not A301) );
 a28751a <=( a28750a  and  a28747a );
 a28752a <=( a28751a  and  a28744a );
 a28756a <=( (not A167)  and  A168 );
 a28757a <=( (not A170)  and  a28756a );
 a28760a <=( (not A199)  and  A166 );
 a28763a <=( A232  and  (not A200) );
 a28764a <=( a28763a  and  a28760a );
 a28765a <=( a28764a  and  a28757a );
 a28768a <=( A234  and  (not A233) );
 a28771a <=( (not A298)  and  A235 );
 a28772a <=( a28771a  and  a28768a );
 a28775a <=( (not A300)  and  A299 );
 a28778a <=( (not A302)  and  (not A301) );
 a28779a <=( a28778a  and  a28775a );
 a28780a <=( a28779a  and  a28772a );
 a28784a <=( (not A167)  and  A168 );
 a28785a <=( (not A170)  and  a28784a );
 a28788a <=( (not A199)  and  A166 );
 a28791a <=( A232  and  (not A200) );
 a28792a <=( a28791a  and  a28788a );
 a28793a <=( a28792a  and  a28785a );
 a28796a <=( A234  and  (not A233) );
 a28799a <=( (not A265)  and  A235 );
 a28800a <=( a28799a  and  a28796a );
 a28803a <=( (not A267)  and  A266 );
 a28806a <=( (not A269)  and  (not A268) );
 a28807a <=( a28806a  and  a28803a );
 a28808a <=( a28807a  and  a28800a );
 a28812a <=( (not A167)  and  A168 );
 a28813a <=( (not A170)  and  a28812a );
 a28816a <=( (not A199)  and  A166 );
 a28819a <=( A232  and  (not A200) );
 a28820a <=( a28819a  and  a28816a );
 a28821a <=( a28820a  and  a28813a );
 a28824a <=( A234  and  (not A233) );
 a28827a <=( A265  and  A235 );
 a28828a <=( a28827a  and  a28824a );
 a28831a <=( (not A267)  and  (not A266) );
 a28834a <=( (not A269)  and  (not A268) );
 a28835a <=( a28834a  and  a28831a );
 a28836a <=( a28835a  and  a28828a );
 a28840a <=( (not A167)  and  A168 );
 a28841a <=( (not A170)  and  a28840a );
 a28844a <=( (not A199)  and  A166 );
 a28847a <=( A232  and  (not A200) );
 a28848a <=( a28847a  and  a28844a );
 a28849a <=( a28848a  and  a28841a );
 a28852a <=( A234  and  (not A233) );
 a28855a <=( A298  and  A236 );
 a28856a <=( a28855a  and  a28852a );
 a28859a <=( (not A300)  and  (not A299) );
 a28862a <=( (not A302)  and  (not A301) );
 a28863a <=( a28862a  and  a28859a );
 a28864a <=( a28863a  and  a28856a );
 a28868a <=( (not A167)  and  A168 );
 a28869a <=( (not A170)  and  a28868a );
 a28872a <=( (not A199)  and  A166 );
 a28875a <=( A232  and  (not A200) );
 a28876a <=( a28875a  and  a28872a );
 a28877a <=( a28876a  and  a28869a );
 a28880a <=( A234  and  (not A233) );
 a28883a <=( (not A298)  and  A236 );
 a28884a <=( a28883a  and  a28880a );
 a28887a <=( (not A300)  and  A299 );
 a28890a <=( (not A302)  and  (not A301) );
 a28891a <=( a28890a  and  a28887a );
 a28892a <=( a28891a  and  a28884a );
 a28896a <=( (not A167)  and  A168 );
 a28897a <=( (not A170)  and  a28896a );
 a28900a <=( (not A199)  and  A166 );
 a28903a <=( A232  and  (not A200) );
 a28904a <=( a28903a  and  a28900a );
 a28905a <=( a28904a  and  a28897a );
 a28908a <=( A234  and  (not A233) );
 a28911a <=( (not A265)  and  A236 );
 a28912a <=( a28911a  and  a28908a );
 a28915a <=( (not A267)  and  A266 );
 a28918a <=( (not A269)  and  (not A268) );
 a28919a <=( a28918a  and  a28915a );
 a28920a <=( a28919a  and  a28912a );
 a28924a <=( (not A167)  and  A168 );
 a28925a <=( (not A170)  and  a28924a );
 a28928a <=( (not A199)  and  A166 );
 a28931a <=( A232  and  (not A200) );
 a28932a <=( a28931a  and  a28928a );
 a28933a <=( a28932a  and  a28925a );
 a28936a <=( A234  and  (not A233) );
 a28939a <=( A265  and  A236 );
 a28940a <=( a28939a  and  a28936a );
 a28943a <=( (not A267)  and  (not A266) );
 a28946a <=( (not A269)  and  (not A268) );
 a28947a <=( a28946a  and  a28943a );
 a28948a <=( a28947a  and  a28940a );
 a28952a <=( (not A167)  and  A168 );
 a28953a <=( (not A170)  and  a28952a );
 a28956a <=( (not A199)  and  A166 );
 a28959a <=( A232  and  (not A200) );
 a28960a <=( a28959a  and  a28956a );
 a28961a <=( a28960a  and  a28953a );
 a28964a <=( (not A234)  and  (not A233) );
 a28967a <=( (not A236)  and  (not A235) );
 a28968a <=( a28967a  and  a28964a );
 a28971a <=( (not A299)  and  A298 );
 a28974a <=( A301  and  A300 );
 a28975a <=( a28974a  and  a28971a );
 a28976a <=( a28975a  and  a28968a );
 a28980a <=( (not A167)  and  A168 );
 a28981a <=( (not A170)  and  a28980a );
 a28984a <=( (not A199)  and  A166 );
 a28987a <=( A232  and  (not A200) );
 a28988a <=( a28987a  and  a28984a );
 a28989a <=( a28988a  and  a28981a );
 a28992a <=( (not A234)  and  (not A233) );
 a28995a <=( (not A236)  and  (not A235) );
 a28996a <=( a28995a  and  a28992a );
 a28999a <=( (not A299)  and  A298 );
 a29002a <=( A302  and  A300 );
 a29003a <=( a29002a  and  a28999a );
 a29004a <=( a29003a  and  a28996a );
 a29008a <=( (not A167)  and  A168 );
 a29009a <=( (not A170)  and  a29008a );
 a29012a <=( (not A199)  and  A166 );
 a29015a <=( A232  and  (not A200) );
 a29016a <=( a29015a  and  a29012a );
 a29017a <=( a29016a  and  a29009a );
 a29020a <=( (not A234)  and  (not A233) );
 a29023a <=( (not A236)  and  (not A235) );
 a29024a <=( a29023a  and  a29020a );
 a29027a <=( A299  and  (not A298) );
 a29030a <=( A301  and  A300 );
 a29031a <=( a29030a  and  a29027a );
 a29032a <=( a29031a  and  a29024a );
 a29036a <=( (not A167)  and  A168 );
 a29037a <=( (not A170)  and  a29036a );
 a29040a <=( (not A199)  and  A166 );
 a29043a <=( A232  and  (not A200) );
 a29044a <=( a29043a  and  a29040a );
 a29045a <=( a29044a  and  a29037a );
 a29048a <=( (not A234)  and  (not A233) );
 a29051a <=( (not A236)  and  (not A235) );
 a29052a <=( a29051a  and  a29048a );
 a29055a <=( A299  and  (not A298) );
 a29058a <=( A302  and  A300 );
 a29059a <=( a29058a  and  a29055a );
 a29060a <=( a29059a  and  a29052a );
 a29064a <=( (not A167)  and  A168 );
 a29065a <=( (not A170)  and  a29064a );
 a29068a <=( (not A199)  and  A166 );
 a29071a <=( A232  and  (not A200) );
 a29072a <=( a29071a  and  a29068a );
 a29073a <=( a29072a  and  a29065a );
 a29076a <=( (not A234)  and  (not A233) );
 a29079a <=( (not A236)  and  (not A235) );
 a29080a <=( a29079a  and  a29076a );
 a29083a <=( A266  and  (not A265) );
 a29086a <=( A268  and  A267 );
 a29087a <=( a29086a  and  a29083a );
 a29088a <=( a29087a  and  a29080a );
 a29092a <=( (not A167)  and  A168 );
 a29093a <=( (not A170)  and  a29092a );
 a29096a <=( (not A199)  and  A166 );
 a29099a <=( A232  and  (not A200) );
 a29100a <=( a29099a  and  a29096a );
 a29101a <=( a29100a  and  a29093a );
 a29104a <=( (not A234)  and  (not A233) );
 a29107a <=( (not A236)  and  (not A235) );
 a29108a <=( a29107a  and  a29104a );
 a29111a <=( A266  and  (not A265) );
 a29114a <=( A269  and  A267 );
 a29115a <=( a29114a  and  a29111a );
 a29116a <=( a29115a  and  a29108a );
 a29120a <=( (not A167)  and  A168 );
 a29121a <=( (not A170)  and  a29120a );
 a29124a <=( (not A199)  and  A166 );
 a29127a <=( A232  and  (not A200) );
 a29128a <=( a29127a  and  a29124a );
 a29129a <=( a29128a  and  a29121a );
 a29132a <=( (not A234)  and  (not A233) );
 a29135a <=( (not A236)  and  (not A235) );
 a29136a <=( a29135a  and  a29132a );
 a29139a <=( (not A266)  and  A265 );
 a29142a <=( A268  and  A267 );
 a29143a <=( a29142a  and  a29139a );
 a29144a <=( a29143a  and  a29136a );
 a29148a <=( (not A167)  and  A168 );
 a29149a <=( (not A170)  and  a29148a );
 a29152a <=( (not A199)  and  A166 );
 a29155a <=( A232  and  (not A200) );
 a29156a <=( a29155a  and  a29152a );
 a29157a <=( a29156a  and  a29149a );
 a29160a <=( (not A234)  and  (not A233) );
 a29163a <=( (not A236)  and  (not A235) );
 a29164a <=( a29163a  and  a29160a );
 a29167a <=( (not A266)  and  A265 );
 a29170a <=( A269  and  A267 );
 a29171a <=( a29170a  and  a29167a );
 a29172a <=( a29171a  and  a29164a );
 a29176a <=( A167  and  A168 );
 a29177a <=( A169  and  a29176a );
 a29180a <=( A201  and  (not A166) );
 a29183a <=( (not A203)  and  (not A202) );
 a29184a <=( a29183a  and  a29180a );
 a29185a <=( a29184a  and  a29177a );
 a29188a <=( A233  and  (not A232) );
 a29191a <=( A235  and  A234 );
 a29192a <=( a29191a  and  a29188a );
 a29195a <=( (not A299)  and  A298 );
 a29198a <=( A301  and  A300 );
 a29199a <=( a29198a  and  a29195a );
 a29200a <=( a29199a  and  a29192a );
 a29204a <=( A167  and  A168 );
 a29205a <=( A169  and  a29204a );
 a29208a <=( A201  and  (not A166) );
 a29211a <=( (not A203)  and  (not A202) );
 a29212a <=( a29211a  and  a29208a );
 a29213a <=( a29212a  and  a29205a );
 a29216a <=( A233  and  (not A232) );
 a29219a <=( A235  and  A234 );
 a29220a <=( a29219a  and  a29216a );
 a29223a <=( (not A299)  and  A298 );
 a29226a <=( A302  and  A300 );
 a29227a <=( a29226a  and  a29223a );
 a29228a <=( a29227a  and  a29220a );
 a29232a <=( A167  and  A168 );
 a29233a <=( A169  and  a29232a );
 a29236a <=( A201  and  (not A166) );
 a29239a <=( (not A203)  and  (not A202) );
 a29240a <=( a29239a  and  a29236a );
 a29241a <=( a29240a  and  a29233a );
 a29244a <=( A233  and  (not A232) );
 a29247a <=( A235  and  A234 );
 a29248a <=( a29247a  and  a29244a );
 a29251a <=( A299  and  (not A298) );
 a29254a <=( A301  and  A300 );
 a29255a <=( a29254a  and  a29251a );
 a29256a <=( a29255a  and  a29248a );
 a29260a <=( A167  and  A168 );
 a29261a <=( A169  and  a29260a );
 a29264a <=( A201  and  (not A166) );
 a29267a <=( (not A203)  and  (not A202) );
 a29268a <=( a29267a  and  a29264a );
 a29269a <=( a29268a  and  a29261a );
 a29272a <=( A233  and  (not A232) );
 a29275a <=( A235  and  A234 );
 a29276a <=( a29275a  and  a29272a );
 a29279a <=( A299  and  (not A298) );
 a29282a <=( A302  and  A300 );
 a29283a <=( a29282a  and  a29279a );
 a29284a <=( a29283a  and  a29276a );
 a29288a <=( A167  and  A168 );
 a29289a <=( A169  and  a29288a );
 a29292a <=( A201  and  (not A166) );
 a29295a <=( (not A203)  and  (not A202) );
 a29296a <=( a29295a  and  a29292a );
 a29297a <=( a29296a  and  a29289a );
 a29300a <=( A233  and  (not A232) );
 a29303a <=( A235  and  A234 );
 a29304a <=( a29303a  and  a29300a );
 a29307a <=( A266  and  (not A265) );
 a29310a <=( A268  and  A267 );
 a29311a <=( a29310a  and  a29307a );
 a29312a <=( a29311a  and  a29304a );
 a29316a <=( A167  and  A168 );
 a29317a <=( A169  and  a29316a );
 a29320a <=( A201  and  (not A166) );
 a29323a <=( (not A203)  and  (not A202) );
 a29324a <=( a29323a  and  a29320a );
 a29325a <=( a29324a  and  a29317a );
 a29328a <=( A233  and  (not A232) );
 a29331a <=( A235  and  A234 );
 a29332a <=( a29331a  and  a29328a );
 a29335a <=( A266  and  (not A265) );
 a29338a <=( A269  and  A267 );
 a29339a <=( a29338a  and  a29335a );
 a29340a <=( a29339a  and  a29332a );
 a29344a <=( A167  and  A168 );
 a29345a <=( A169  and  a29344a );
 a29348a <=( A201  and  (not A166) );
 a29351a <=( (not A203)  and  (not A202) );
 a29352a <=( a29351a  and  a29348a );
 a29353a <=( a29352a  and  a29345a );
 a29356a <=( A233  and  (not A232) );
 a29359a <=( A235  and  A234 );
 a29360a <=( a29359a  and  a29356a );
 a29363a <=( (not A266)  and  A265 );
 a29366a <=( A268  and  A267 );
 a29367a <=( a29366a  and  a29363a );
 a29368a <=( a29367a  and  a29360a );
 a29372a <=( A167  and  A168 );
 a29373a <=( A169  and  a29372a );
 a29376a <=( A201  and  (not A166) );
 a29379a <=( (not A203)  and  (not A202) );
 a29380a <=( a29379a  and  a29376a );
 a29381a <=( a29380a  and  a29373a );
 a29384a <=( A233  and  (not A232) );
 a29387a <=( A235  and  A234 );
 a29388a <=( a29387a  and  a29384a );
 a29391a <=( (not A266)  and  A265 );
 a29394a <=( A269  and  A267 );
 a29395a <=( a29394a  and  a29391a );
 a29396a <=( a29395a  and  a29388a );
 a29400a <=( A167  and  A168 );
 a29401a <=( A169  and  a29400a );
 a29404a <=( A201  and  (not A166) );
 a29407a <=( (not A203)  and  (not A202) );
 a29408a <=( a29407a  and  a29404a );
 a29409a <=( a29408a  and  a29401a );
 a29412a <=( A233  and  (not A232) );
 a29415a <=( A236  and  A234 );
 a29416a <=( a29415a  and  a29412a );
 a29419a <=( (not A299)  and  A298 );
 a29422a <=( A301  and  A300 );
 a29423a <=( a29422a  and  a29419a );
 a29424a <=( a29423a  and  a29416a );
 a29428a <=( A167  and  A168 );
 a29429a <=( A169  and  a29428a );
 a29432a <=( A201  and  (not A166) );
 a29435a <=( (not A203)  and  (not A202) );
 a29436a <=( a29435a  and  a29432a );
 a29437a <=( a29436a  and  a29429a );
 a29440a <=( A233  and  (not A232) );
 a29443a <=( A236  and  A234 );
 a29444a <=( a29443a  and  a29440a );
 a29447a <=( (not A299)  and  A298 );
 a29450a <=( A302  and  A300 );
 a29451a <=( a29450a  and  a29447a );
 a29452a <=( a29451a  and  a29444a );
 a29456a <=( A167  and  A168 );
 a29457a <=( A169  and  a29456a );
 a29460a <=( A201  and  (not A166) );
 a29463a <=( (not A203)  and  (not A202) );
 a29464a <=( a29463a  and  a29460a );
 a29465a <=( a29464a  and  a29457a );
 a29468a <=( A233  and  (not A232) );
 a29471a <=( A236  and  A234 );
 a29472a <=( a29471a  and  a29468a );
 a29475a <=( A299  and  (not A298) );
 a29478a <=( A301  and  A300 );
 a29479a <=( a29478a  and  a29475a );
 a29480a <=( a29479a  and  a29472a );
 a29484a <=( A167  and  A168 );
 a29485a <=( A169  and  a29484a );
 a29488a <=( A201  and  (not A166) );
 a29491a <=( (not A203)  and  (not A202) );
 a29492a <=( a29491a  and  a29488a );
 a29493a <=( a29492a  and  a29485a );
 a29496a <=( A233  and  (not A232) );
 a29499a <=( A236  and  A234 );
 a29500a <=( a29499a  and  a29496a );
 a29503a <=( A299  and  (not A298) );
 a29506a <=( A302  and  A300 );
 a29507a <=( a29506a  and  a29503a );
 a29508a <=( a29507a  and  a29500a );
 a29512a <=( A167  and  A168 );
 a29513a <=( A169  and  a29512a );
 a29516a <=( A201  and  (not A166) );
 a29519a <=( (not A203)  and  (not A202) );
 a29520a <=( a29519a  and  a29516a );
 a29521a <=( a29520a  and  a29513a );
 a29524a <=( A233  and  (not A232) );
 a29527a <=( A236  and  A234 );
 a29528a <=( a29527a  and  a29524a );
 a29531a <=( A266  and  (not A265) );
 a29534a <=( A268  and  A267 );
 a29535a <=( a29534a  and  a29531a );
 a29536a <=( a29535a  and  a29528a );
 a29540a <=( A167  and  A168 );
 a29541a <=( A169  and  a29540a );
 a29544a <=( A201  and  (not A166) );
 a29547a <=( (not A203)  and  (not A202) );
 a29548a <=( a29547a  and  a29544a );
 a29549a <=( a29548a  and  a29541a );
 a29552a <=( A233  and  (not A232) );
 a29555a <=( A236  and  A234 );
 a29556a <=( a29555a  and  a29552a );
 a29559a <=( A266  and  (not A265) );
 a29562a <=( A269  and  A267 );
 a29563a <=( a29562a  and  a29559a );
 a29564a <=( a29563a  and  a29556a );
 a29568a <=( A167  and  A168 );
 a29569a <=( A169  and  a29568a );
 a29572a <=( A201  and  (not A166) );
 a29575a <=( (not A203)  and  (not A202) );
 a29576a <=( a29575a  and  a29572a );
 a29577a <=( a29576a  and  a29569a );
 a29580a <=( A233  and  (not A232) );
 a29583a <=( A236  and  A234 );
 a29584a <=( a29583a  and  a29580a );
 a29587a <=( (not A266)  and  A265 );
 a29590a <=( A268  and  A267 );
 a29591a <=( a29590a  and  a29587a );
 a29592a <=( a29591a  and  a29584a );
 a29596a <=( A167  and  A168 );
 a29597a <=( A169  and  a29596a );
 a29600a <=( A201  and  (not A166) );
 a29603a <=( (not A203)  and  (not A202) );
 a29604a <=( a29603a  and  a29600a );
 a29605a <=( a29604a  and  a29597a );
 a29608a <=( A233  and  (not A232) );
 a29611a <=( A236  and  A234 );
 a29612a <=( a29611a  and  a29608a );
 a29615a <=( (not A266)  and  A265 );
 a29618a <=( A269  and  A267 );
 a29619a <=( a29618a  and  a29615a );
 a29620a <=( a29619a  and  a29612a );
 a29624a <=( A167  and  A168 );
 a29625a <=( A169  and  a29624a );
 a29628a <=( A201  and  (not A166) );
 a29631a <=( (not A203)  and  (not A202) );
 a29632a <=( a29631a  and  a29628a );
 a29633a <=( a29632a  and  a29625a );
 a29636a <=( (not A233)  and  A232 );
 a29639a <=( A235  and  A234 );
 a29640a <=( a29639a  and  a29636a );
 a29643a <=( (not A299)  and  A298 );
 a29646a <=( A301  and  A300 );
 a29647a <=( a29646a  and  a29643a );
 a29648a <=( a29647a  and  a29640a );
 a29652a <=( A167  and  A168 );
 a29653a <=( A169  and  a29652a );
 a29656a <=( A201  and  (not A166) );
 a29659a <=( (not A203)  and  (not A202) );
 a29660a <=( a29659a  and  a29656a );
 a29661a <=( a29660a  and  a29653a );
 a29664a <=( (not A233)  and  A232 );
 a29667a <=( A235  and  A234 );
 a29668a <=( a29667a  and  a29664a );
 a29671a <=( (not A299)  and  A298 );
 a29674a <=( A302  and  A300 );
 a29675a <=( a29674a  and  a29671a );
 a29676a <=( a29675a  and  a29668a );
 a29680a <=( A167  and  A168 );
 a29681a <=( A169  and  a29680a );
 a29684a <=( A201  and  (not A166) );
 a29687a <=( (not A203)  and  (not A202) );
 a29688a <=( a29687a  and  a29684a );
 a29689a <=( a29688a  and  a29681a );
 a29692a <=( (not A233)  and  A232 );
 a29695a <=( A235  and  A234 );
 a29696a <=( a29695a  and  a29692a );
 a29699a <=( A299  and  (not A298) );
 a29702a <=( A301  and  A300 );
 a29703a <=( a29702a  and  a29699a );
 a29704a <=( a29703a  and  a29696a );
 a29708a <=( A167  and  A168 );
 a29709a <=( A169  and  a29708a );
 a29712a <=( A201  and  (not A166) );
 a29715a <=( (not A203)  and  (not A202) );
 a29716a <=( a29715a  and  a29712a );
 a29717a <=( a29716a  and  a29709a );
 a29720a <=( (not A233)  and  A232 );
 a29723a <=( A235  and  A234 );
 a29724a <=( a29723a  and  a29720a );
 a29727a <=( A299  and  (not A298) );
 a29730a <=( A302  and  A300 );
 a29731a <=( a29730a  and  a29727a );
 a29732a <=( a29731a  and  a29724a );
 a29736a <=( A167  and  A168 );
 a29737a <=( A169  and  a29736a );
 a29740a <=( A201  and  (not A166) );
 a29743a <=( (not A203)  and  (not A202) );
 a29744a <=( a29743a  and  a29740a );
 a29745a <=( a29744a  and  a29737a );
 a29748a <=( (not A233)  and  A232 );
 a29751a <=( A235  and  A234 );
 a29752a <=( a29751a  and  a29748a );
 a29755a <=( A266  and  (not A265) );
 a29758a <=( A268  and  A267 );
 a29759a <=( a29758a  and  a29755a );
 a29760a <=( a29759a  and  a29752a );
 a29764a <=( A167  and  A168 );
 a29765a <=( A169  and  a29764a );
 a29768a <=( A201  and  (not A166) );
 a29771a <=( (not A203)  and  (not A202) );
 a29772a <=( a29771a  and  a29768a );
 a29773a <=( a29772a  and  a29765a );
 a29776a <=( (not A233)  and  A232 );
 a29779a <=( A235  and  A234 );
 a29780a <=( a29779a  and  a29776a );
 a29783a <=( A266  and  (not A265) );
 a29786a <=( A269  and  A267 );
 a29787a <=( a29786a  and  a29783a );
 a29788a <=( a29787a  and  a29780a );
 a29792a <=( A167  and  A168 );
 a29793a <=( A169  and  a29792a );
 a29796a <=( A201  and  (not A166) );
 a29799a <=( (not A203)  and  (not A202) );
 a29800a <=( a29799a  and  a29796a );
 a29801a <=( a29800a  and  a29793a );
 a29804a <=( (not A233)  and  A232 );
 a29807a <=( A235  and  A234 );
 a29808a <=( a29807a  and  a29804a );
 a29811a <=( (not A266)  and  A265 );
 a29814a <=( A268  and  A267 );
 a29815a <=( a29814a  and  a29811a );
 a29816a <=( a29815a  and  a29808a );
 a29820a <=( A167  and  A168 );
 a29821a <=( A169  and  a29820a );
 a29824a <=( A201  and  (not A166) );
 a29827a <=( (not A203)  and  (not A202) );
 a29828a <=( a29827a  and  a29824a );
 a29829a <=( a29828a  and  a29821a );
 a29832a <=( (not A233)  and  A232 );
 a29835a <=( A235  and  A234 );
 a29836a <=( a29835a  and  a29832a );
 a29839a <=( (not A266)  and  A265 );
 a29842a <=( A269  and  A267 );
 a29843a <=( a29842a  and  a29839a );
 a29844a <=( a29843a  and  a29836a );
 a29848a <=( A167  and  A168 );
 a29849a <=( A169  and  a29848a );
 a29852a <=( A201  and  (not A166) );
 a29855a <=( (not A203)  and  (not A202) );
 a29856a <=( a29855a  and  a29852a );
 a29857a <=( a29856a  and  a29849a );
 a29860a <=( (not A233)  and  A232 );
 a29863a <=( A236  and  A234 );
 a29864a <=( a29863a  and  a29860a );
 a29867a <=( (not A299)  and  A298 );
 a29870a <=( A301  and  A300 );
 a29871a <=( a29870a  and  a29867a );
 a29872a <=( a29871a  and  a29864a );
 a29876a <=( A167  and  A168 );
 a29877a <=( A169  and  a29876a );
 a29880a <=( A201  and  (not A166) );
 a29883a <=( (not A203)  and  (not A202) );
 a29884a <=( a29883a  and  a29880a );
 a29885a <=( a29884a  and  a29877a );
 a29888a <=( (not A233)  and  A232 );
 a29891a <=( A236  and  A234 );
 a29892a <=( a29891a  and  a29888a );
 a29895a <=( (not A299)  and  A298 );
 a29898a <=( A302  and  A300 );
 a29899a <=( a29898a  and  a29895a );
 a29900a <=( a29899a  and  a29892a );
 a29904a <=( A167  and  A168 );
 a29905a <=( A169  and  a29904a );
 a29908a <=( A201  and  (not A166) );
 a29911a <=( (not A203)  and  (not A202) );
 a29912a <=( a29911a  and  a29908a );
 a29913a <=( a29912a  and  a29905a );
 a29916a <=( (not A233)  and  A232 );
 a29919a <=( A236  and  A234 );
 a29920a <=( a29919a  and  a29916a );
 a29923a <=( A299  and  (not A298) );
 a29926a <=( A301  and  A300 );
 a29927a <=( a29926a  and  a29923a );
 a29928a <=( a29927a  and  a29920a );
 a29932a <=( A167  and  A168 );
 a29933a <=( A169  and  a29932a );
 a29936a <=( A201  and  (not A166) );
 a29939a <=( (not A203)  and  (not A202) );
 a29940a <=( a29939a  and  a29936a );
 a29941a <=( a29940a  and  a29933a );
 a29944a <=( (not A233)  and  A232 );
 a29947a <=( A236  and  A234 );
 a29948a <=( a29947a  and  a29944a );
 a29951a <=( A299  and  (not A298) );
 a29954a <=( A302  and  A300 );
 a29955a <=( a29954a  and  a29951a );
 a29956a <=( a29955a  and  a29948a );
 a29960a <=( A167  and  A168 );
 a29961a <=( A169  and  a29960a );
 a29964a <=( A201  and  (not A166) );
 a29967a <=( (not A203)  and  (not A202) );
 a29968a <=( a29967a  and  a29964a );
 a29969a <=( a29968a  and  a29961a );
 a29972a <=( (not A233)  and  A232 );
 a29975a <=( A236  and  A234 );
 a29976a <=( a29975a  and  a29972a );
 a29979a <=( A266  and  (not A265) );
 a29982a <=( A268  and  A267 );
 a29983a <=( a29982a  and  a29979a );
 a29984a <=( a29983a  and  a29976a );
 a29988a <=( A167  and  A168 );
 a29989a <=( A169  and  a29988a );
 a29992a <=( A201  and  (not A166) );
 a29995a <=( (not A203)  and  (not A202) );
 a29996a <=( a29995a  and  a29992a );
 a29997a <=( a29996a  and  a29989a );
 a30000a <=( (not A233)  and  A232 );
 a30003a <=( A236  and  A234 );
 a30004a <=( a30003a  and  a30000a );
 a30007a <=( A266  and  (not A265) );
 a30010a <=( A269  and  A267 );
 a30011a <=( a30010a  and  a30007a );
 a30012a <=( a30011a  and  a30004a );
 a30016a <=( A167  and  A168 );
 a30017a <=( A169  and  a30016a );
 a30020a <=( A201  and  (not A166) );
 a30023a <=( (not A203)  and  (not A202) );
 a30024a <=( a30023a  and  a30020a );
 a30025a <=( a30024a  and  a30017a );
 a30028a <=( (not A233)  and  A232 );
 a30031a <=( A236  and  A234 );
 a30032a <=( a30031a  and  a30028a );
 a30035a <=( (not A266)  and  A265 );
 a30038a <=( A268  and  A267 );
 a30039a <=( a30038a  and  a30035a );
 a30040a <=( a30039a  and  a30032a );
 a30044a <=( A167  and  A168 );
 a30045a <=( A169  and  a30044a );
 a30048a <=( A201  and  (not A166) );
 a30051a <=( (not A203)  and  (not A202) );
 a30052a <=( a30051a  and  a30048a );
 a30053a <=( a30052a  and  a30045a );
 a30056a <=( (not A233)  and  A232 );
 a30059a <=( A236  and  A234 );
 a30060a <=( a30059a  and  a30056a );
 a30063a <=( (not A266)  and  A265 );
 a30066a <=( A269  and  A267 );
 a30067a <=( a30066a  and  a30063a );
 a30068a <=( a30067a  and  a30060a );
 a30072a <=( A167  and  A168 );
 a30073a <=( A169  and  a30072a );
 a30076a <=( (not A201)  and  (not A166) );
 a30079a <=( (not A232)  and  A202 );
 a30080a <=( a30079a  and  a30076a );
 a30081a <=( a30080a  and  a30073a );
 a30084a <=( A234  and  A233 );
 a30087a <=( A298  and  A235 );
 a30088a <=( a30087a  and  a30084a );
 a30091a <=( (not A300)  and  (not A299) );
 a30094a <=( (not A302)  and  (not A301) );
 a30095a <=( a30094a  and  a30091a );
 a30096a <=( a30095a  and  a30088a );
 a30100a <=( A167  and  A168 );
 a30101a <=( A169  and  a30100a );
 a30104a <=( (not A201)  and  (not A166) );
 a30107a <=( (not A232)  and  A202 );
 a30108a <=( a30107a  and  a30104a );
 a30109a <=( a30108a  and  a30101a );
 a30112a <=( A234  and  A233 );
 a30115a <=( (not A298)  and  A235 );
 a30116a <=( a30115a  and  a30112a );
 a30119a <=( (not A300)  and  A299 );
 a30122a <=( (not A302)  and  (not A301) );
 a30123a <=( a30122a  and  a30119a );
 a30124a <=( a30123a  and  a30116a );
 a30128a <=( A167  and  A168 );
 a30129a <=( A169  and  a30128a );
 a30132a <=( (not A201)  and  (not A166) );
 a30135a <=( (not A232)  and  A202 );
 a30136a <=( a30135a  and  a30132a );
 a30137a <=( a30136a  and  a30129a );
 a30140a <=( A234  and  A233 );
 a30143a <=( (not A265)  and  A235 );
 a30144a <=( a30143a  and  a30140a );
 a30147a <=( (not A267)  and  A266 );
 a30150a <=( (not A269)  and  (not A268) );
 a30151a <=( a30150a  and  a30147a );
 a30152a <=( a30151a  and  a30144a );
 a30156a <=( A167  and  A168 );
 a30157a <=( A169  and  a30156a );
 a30160a <=( (not A201)  and  (not A166) );
 a30163a <=( (not A232)  and  A202 );
 a30164a <=( a30163a  and  a30160a );
 a30165a <=( a30164a  and  a30157a );
 a30168a <=( A234  and  A233 );
 a30171a <=( A265  and  A235 );
 a30172a <=( a30171a  and  a30168a );
 a30175a <=( (not A267)  and  (not A266) );
 a30178a <=( (not A269)  and  (not A268) );
 a30179a <=( a30178a  and  a30175a );
 a30180a <=( a30179a  and  a30172a );
 a30184a <=( A167  and  A168 );
 a30185a <=( A169  and  a30184a );
 a30188a <=( (not A201)  and  (not A166) );
 a30191a <=( (not A232)  and  A202 );
 a30192a <=( a30191a  and  a30188a );
 a30193a <=( a30192a  and  a30185a );
 a30196a <=( A234  and  A233 );
 a30199a <=( A298  and  A236 );
 a30200a <=( a30199a  and  a30196a );
 a30203a <=( (not A300)  and  (not A299) );
 a30206a <=( (not A302)  and  (not A301) );
 a30207a <=( a30206a  and  a30203a );
 a30208a <=( a30207a  and  a30200a );
 a30212a <=( A167  and  A168 );
 a30213a <=( A169  and  a30212a );
 a30216a <=( (not A201)  and  (not A166) );
 a30219a <=( (not A232)  and  A202 );
 a30220a <=( a30219a  and  a30216a );
 a30221a <=( a30220a  and  a30213a );
 a30224a <=( A234  and  A233 );
 a30227a <=( (not A298)  and  A236 );
 a30228a <=( a30227a  and  a30224a );
 a30231a <=( (not A300)  and  A299 );
 a30234a <=( (not A302)  and  (not A301) );
 a30235a <=( a30234a  and  a30231a );
 a30236a <=( a30235a  and  a30228a );
 a30240a <=( A167  and  A168 );
 a30241a <=( A169  and  a30240a );
 a30244a <=( (not A201)  and  (not A166) );
 a30247a <=( (not A232)  and  A202 );
 a30248a <=( a30247a  and  a30244a );
 a30249a <=( a30248a  and  a30241a );
 a30252a <=( A234  and  A233 );
 a30255a <=( (not A265)  and  A236 );
 a30256a <=( a30255a  and  a30252a );
 a30259a <=( (not A267)  and  A266 );
 a30262a <=( (not A269)  and  (not A268) );
 a30263a <=( a30262a  and  a30259a );
 a30264a <=( a30263a  and  a30256a );
 a30268a <=( A167  and  A168 );
 a30269a <=( A169  and  a30268a );
 a30272a <=( (not A201)  and  (not A166) );
 a30275a <=( (not A232)  and  A202 );
 a30276a <=( a30275a  and  a30272a );
 a30277a <=( a30276a  and  a30269a );
 a30280a <=( A234  and  A233 );
 a30283a <=( A265  and  A236 );
 a30284a <=( a30283a  and  a30280a );
 a30287a <=( (not A267)  and  (not A266) );
 a30290a <=( (not A269)  and  (not A268) );
 a30291a <=( a30290a  and  a30287a );
 a30292a <=( a30291a  and  a30284a );
 a30296a <=( A167  and  A168 );
 a30297a <=( A169  and  a30296a );
 a30300a <=( (not A201)  and  (not A166) );
 a30303a <=( (not A232)  and  A202 );
 a30304a <=( a30303a  and  a30300a );
 a30305a <=( a30304a  and  a30297a );
 a30308a <=( (not A234)  and  A233 );
 a30311a <=( (not A236)  and  (not A235) );
 a30312a <=( a30311a  and  a30308a );
 a30315a <=( (not A299)  and  A298 );
 a30318a <=( A301  and  A300 );
 a30319a <=( a30318a  and  a30315a );
 a30320a <=( a30319a  and  a30312a );
 a30324a <=( A167  and  A168 );
 a30325a <=( A169  and  a30324a );
 a30328a <=( (not A201)  and  (not A166) );
 a30331a <=( (not A232)  and  A202 );
 a30332a <=( a30331a  and  a30328a );
 a30333a <=( a30332a  and  a30325a );
 a30336a <=( (not A234)  and  A233 );
 a30339a <=( (not A236)  and  (not A235) );
 a30340a <=( a30339a  and  a30336a );
 a30343a <=( (not A299)  and  A298 );
 a30346a <=( A302  and  A300 );
 a30347a <=( a30346a  and  a30343a );
 a30348a <=( a30347a  and  a30340a );
 a30352a <=( A167  and  A168 );
 a30353a <=( A169  and  a30352a );
 a30356a <=( (not A201)  and  (not A166) );
 a30359a <=( (not A232)  and  A202 );
 a30360a <=( a30359a  and  a30356a );
 a30361a <=( a30360a  and  a30353a );
 a30364a <=( (not A234)  and  A233 );
 a30367a <=( (not A236)  and  (not A235) );
 a30368a <=( a30367a  and  a30364a );
 a30371a <=( A299  and  (not A298) );
 a30374a <=( A301  and  A300 );
 a30375a <=( a30374a  and  a30371a );
 a30376a <=( a30375a  and  a30368a );
 a30380a <=( A167  and  A168 );
 a30381a <=( A169  and  a30380a );
 a30384a <=( (not A201)  and  (not A166) );
 a30387a <=( (not A232)  and  A202 );
 a30388a <=( a30387a  and  a30384a );
 a30389a <=( a30388a  and  a30381a );
 a30392a <=( (not A234)  and  A233 );
 a30395a <=( (not A236)  and  (not A235) );
 a30396a <=( a30395a  and  a30392a );
 a30399a <=( A299  and  (not A298) );
 a30402a <=( A302  and  A300 );
 a30403a <=( a30402a  and  a30399a );
 a30404a <=( a30403a  and  a30396a );
 a30408a <=( A167  and  A168 );
 a30409a <=( A169  and  a30408a );
 a30412a <=( (not A201)  and  (not A166) );
 a30415a <=( (not A232)  and  A202 );
 a30416a <=( a30415a  and  a30412a );
 a30417a <=( a30416a  and  a30409a );
 a30420a <=( (not A234)  and  A233 );
 a30423a <=( (not A236)  and  (not A235) );
 a30424a <=( a30423a  and  a30420a );
 a30427a <=( A266  and  (not A265) );
 a30430a <=( A268  and  A267 );
 a30431a <=( a30430a  and  a30427a );
 a30432a <=( a30431a  and  a30424a );
 a30436a <=( A167  and  A168 );
 a30437a <=( A169  and  a30436a );
 a30440a <=( (not A201)  and  (not A166) );
 a30443a <=( (not A232)  and  A202 );
 a30444a <=( a30443a  and  a30440a );
 a30445a <=( a30444a  and  a30437a );
 a30448a <=( (not A234)  and  A233 );
 a30451a <=( (not A236)  and  (not A235) );
 a30452a <=( a30451a  and  a30448a );
 a30455a <=( A266  and  (not A265) );
 a30458a <=( A269  and  A267 );
 a30459a <=( a30458a  and  a30455a );
 a30460a <=( a30459a  and  a30452a );
 a30464a <=( A167  and  A168 );
 a30465a <=( A169  and  a30464a );
 a30468a <=( (not A201)  and  (not A166) );
 a30471a <=( (not A232)  and  A202 );
 a30472a <=( a30471a  and  a30468a );
 a30473a <=( a30472a  and  a30465a );
 a30476a <=( (not A234)  and  A233 );
 a30479a <=( (not A236)  and  (not A235) );
 a30480a <=( a30479a  and  a30476a );
 a30483a <=( (not A266)  and  A265 );
 a30486a <=( A268  and  A267 );
 a30487a <=( a30486a  and  a30483a );
 a30488a <=( a30487a  and  a30480a );
 a30492a <=( A167  and  A168 );
 a30493a <=( A169  and  a30492a );
 a30496a <=( (not A201)  and  (not A166) );
 a30499a <=( (not A232)  and  A202 );
 a30500a <=( a30499a  and  a30496a );
 a30501a <=( a30500a  and  a30493a );
 a30504a <=( (not A234)  and  A233 );
 a30507a <=( (not A236)  and  (not A235) );
 a30508a <=( a30507a  and  a30504a );
 a30511a <=( (not A266)  and  A265 );
 a30514a <=( A269  and  A267 );
 a30515a <=( a30514a  and  a30511a );
 a30516a <=( a30515a  and  a30508a );
 a30520a <=( A167  and  A168 );
 a30521a <=( A169  and  a30520a );
 a30524a <=( (not A201)  and  (not A166) );
 a30527a <=( A232  and  A202 );
 a30528a <=( a30527a  and  a30524a );
 a30529a <=( a30528a  and  a30521a );
 a30532a <=( A234  and  (not A233) );
 a30535a <=( A298  and  A235 );
 a30536a <=( a30535a  and  a30532a );
 a30539a <=( (not A300)  and  (not A299) );
 a30542a <=( (not A302)  and  (not A301) );
 a30543a <=( a30542a  and  a30539a );
 a30544a <=( a30543a  and  a30536a );
 a30548a <=( A167  and  A168 );
 a30549a <=( A169  and  a30548a );
 a30552a <=( (not A201)  and  (not A166) );
 a30555a <=( A232  and  A202 );
 a30556a <=( a30555a  and  a30552a );
 a30557a <=( a30556a  and  a30549a );
 a30560a <=( A234  and  (not A233) );
 a30563a <=( (not A298)  and  A235 );
 a30564a <=( a30563a  and  a30560a );
 a30567a <=( (not A300)  and  A299 );
 a30570a <=( (not A302)  and  (not A301) );
 a30571a <=( a30570a  and  a30567a );
 a30572a <=( a30571a  and  a30564a );
 a30576a <=( A167  and  A168 );
 a30577a <=( A169  and  a30576a );
 a30580a <=( (not A201)  and  (not A166) );
 a30583a <=( A232  and  A202 );
 a30584a <=( a30583a  and  a30580a );
 a30585a <=( a30584a  and  a30577a );
 a30588a <=( A234  and  (not A233) );
 a30591a <=( (not A265)  and  A235 );
 a30592a <=( a30591a  and  a30588a );
 a30595a <=( (not A267)  and  A266 );
 a30598a <=( (not A269)  and  (not A268) );
 a30599a <=( a30598a  and  a30595a );
 a30600a <=( a30599a  and  a30592a );
 a30604a <=( A167  and  A168 );
 a30605a <=( A169  and  a30604a );
 a30608a <=( (not A201)  and  (not A166) );
 a30611a <=( A232  and  A202 );
 a30612a <=( a30611a  and  a30608a );
 a30613a <=( a30612a  and  a30605a );
 a30616a <=( A234  and  (not A233) );
 a30619a <=( A265  and  A235 );
 a30620a <=( a30619a  and  a30616a );
 a30623a <=( (not A267)  and  (not A266) );
 a30626a <=( (not A269)  and  (not A268) );
 a30627a <=( a30626a  and  a30623a );
 a30628a <=( a30627a  and  a30620a );
 a30632a <=( A167  and  A168 );
 a30633a <=( A169  and  a30632a );
 a30636a <=( (not A201)  and  (not A166) );
 a30639a <=( A232  and  A202 );
 a30640a <=( a30639a  and  a30636a );
 a30641a <=( a30640a  and  a30633a );
 a30644a <=( A234  and  (not A233) );
 a30647a <=( A298  and  A236 );
 a30648a <=( a30647a  and  a30644a );
 a30651a <=( (not A300)  and  (not A299) );
 a30654a <=( (not A302)  and  (not A301) );
 a30655a <=( a30654a  and  a30651a );
 a30656a <=( a30655a  and  a30648a );
 a30660a <=( A167  and  A168 );
 a30661a <=( A169  and  a30660a );
 a30664a <=( (not A201)  and  (not A166) );
 a30667a <=( A232  and  A202 );
 a30668a <=( a30667a  and  a30664a );
 a30669a <=( a30668a  and  a30661a );
 a30672a <=( A234  and  (not A233) );
 a30675a <=( (not A298)  and  A236 );
 a30676a <=( a30675a  and  a30672a );
 a30679a <=( (not A300)  and  A299 );
 a30682a <=( (not A302)  and  (not A301) );
 a30683a <=( a30682a  and  a30679a );
 a30684a <=( a30683a  and  a30676a );
 a30688a <=( A167  and  A168 );
 a30689a <=( A169  and  a30688a );
 a30692a <=( (not A201)  and  (not A166) );
 a30695a <=( A232  and  A202 );
 a30696a <=( a30695a  and  a30692a );
 a30697a <=( a30696a  and  a30689a );
 a30700a <=( A234  and  (not A233) );
 a30703a <=( (not A265)  and  A236 );
 a30704a <=( a30703a  and  a30700a );
 a30707a <=( (not A267)  and  A266 );
 a30710a <=( (not A269)  and  (not A268) );
 a30711a <=( a30710a  and  a30707a );
 a30712a <=( a30711a  and  a30704a );
 a30716a <=( A167  and  A168 );
 a30717a <=( A169  and  a30716a );
 a30720a <=( (not A201)  and  (not A166) );
 a30723a <=( A232  and  A202 );
 a30724a <=( a30723a  and  a30720a );
 a30725a <=( a30724a  and  a30717a );
 a30728a <=( A234  and  (not A233) );
 a30731a <=( A265  and  A236 );
 a30732a <=( a30731a  and  a30728a );
 a30735a <=( (not A267)  and  (not A266) );
 a30738a <=( (not A269)  and  (not A268) );
 a30739a <=( a30738a  and  a30735a );
 a30740a <=( a30739a  and  a30732a );
 a30744a <=( A167  and  A168 );
 a30745a <=( A169  and  a30744a );
 a30748a <=( (not A201)  and  (not A166) );
 a30751a <=( A232  and  A202 );
 a30752a <=( a30751a  and  a30748a );
 a30753a <=( a30752a  and  a30745a );
 a30756a <=( (not A234)  and  (not A233) );
 a30759a <=( (not A236)  and  (not A235) );
 a30760a <=( a30759a  and  a30756a );
 a30763a <=( (not A299)  and  A298 );
 a30766a <=( A301  and  A300 );
 a30767a <=( a30766a  and  a30763a );
 a30768a <=( a30767a  and  a30760a );
 a30772a <=( A167  and  A168 );
 a30773a <=( A169  and  a30772a );
 a30776a <=( (not A201)  and  (not A166) );
 a30779a <=( A232  and  A202 );
 a30780a <=( a30779a  and  a30776a );
 a30781a <=( a30780a  and  a30773a );
 a30784a <=( (not A234)  and  (not A233) );
 a30787a <=( (not A236)  and  (not A235) );
 a30788a <=( a30787a  and  a30784a );
 a30791a <=( (not A299)  and  A298 );
 a30794a <=( A302  and  A300 );
 a30795a <=( a30794a  and  a30791a );
 a30796a <=( a30795a  and  a30788a );
 a30800a <=( A167  and  A168 );
 a30801a <=( A169  and  a30800a );
 a30804a <=( (not A201)  and  (not A166) );
 a30807a <=( A232  and  A202 );
 a30808a <=( a30807a  and  a30804a );
 a30809a <=( a30808a  and  a30801a );
 a30812a <=( (not A234)  and  (not A233) );
 a30815a <=( (not A236)  and  (not A235) );
 a30816a <=( a30815a  and  a30812a );
 a30819a <=( A299  and  (not A298) );
 a30822a <=( A301  and  A300 );
 a30823a <=( a30822a  and  a30819a );
 a30824a <=( a30823a  and  a30816a );
 a30828a <=( A167  and  A168 );
 a30829a <=( A169  and  a30828a );
 a30832a <=( (not A201)  and  (not A166) );
 a30835a <=( A232  and  A202 );
 a30836a <=( a30835a  and  a30832a );
 a30837a <=( a30836a  and  a30829a );
 a30840a <=( (not A234)  and  (not A233) );
 a30843a <=( (not A236)  and  (not A235) );
 a30844a <=( a30843a  and  a30840a );
 a30847a <=( A299  and  (not A298) );
 a30850a <=( A302  and  A300 );
 a30851a <=( a30850a  and  a30847a );
 a30852a <=( a30851a  and  a30844a );
 a30856a <=( A167  and  A168 );
 a30857a <=( A169  and  a30856a );
 a30860a <=( (not A201)  and  (not A166) );
 a30863a <=( A232  and  A202 );
 a30864a <=( a30863a  and  a30860a );
 a30865a <=( a30864a  and  a30857a );
 a30868a <=( (not A234)  and  (not A233) );
 a30871a <=( (not A236)  and  (not A235) );
 a30872a <=( a30871a  and  a30868a );
 a30875a <=( A266  and  (not A265) );
 a30878a <=( A268  and  A267 );
 a30879a <=( a30878a  and  a30875a );
 a30880a <=( a30879a  and  a30872a );
 a30884a <=( A167  and  A168 );
 a30885a <=( A169  and  a30884a );
 a30888a <=( (not A201)  and  (not A166) );
 a30891a <=( A232  and  A202 );
 a30892a <=( a30891a  and  a30888a );
 a30893a <=( a30892a  and  a30885a );
 a30896a <=( (not A234)  and  (not A233) );
 a30899a <=( (not A236)  and  (not A235) );
 a30900a <=( a30899a  and  a30896a );
 a30903a <=( A266  and  (not A265) );
 a30906a <=( A269  and  A267 );
 a30907a <=( a30906a  and  a30903a );
 a30908a <=( a30907a  and  a30900a );
 a30912a <=( A167  and  A168 );
 a30913a <=( A169  and  a30912a );
 a30916a <=( (not A201)  and  (not A166) );
 a30919a <=( A232  and  A202 );
 a30920a <=( a30919a  and  a30916a );
 a30921a <=( a30920a  and  a30913a );
 a30924a <=( (not A234)  and  (not A233) );
 a30927a <=( (not A236)  and  (not A235) );
 a30928a <=( a30927a  and  a30924a );
 a30931a <=( (not A266)  and  A265 );
 a30934a <=( A268  and  A267 );
 a30935a <=( a30934a  and  a30931a );
 a30936a <=( a30935a  and  a30928a );
 a30940a <=( A167  and  A168 );
 a30941a <=( A169  and  a30940a );
 a30944a <=( (not A201)  and  (not A166) );
 a30947a <=( A232  and  A202 );
 a30948a <=( a30947a  and  a30944a );
 a30949a <=( a30948a  and  a30941a );
 a30952a <=( (not A234)  and  (not A233) );
 a30955a <=( (not A236)  and  (not A235) );
 a30956a <=( a30955a  and  a30952a );
 a30959a <=( (not A266)  and  A265 );
 a30962a <=( A269  and  A267 );
 a30963a <=( a30962a  and  a30959a );
 a30964a <=( a30963a  and  a30956a );
 a30968a <=( A167  and  A168 );
 a30969a <=( A169  and  a30968a );
 a30972a <=( (not A201)  and  (not A166) );
 a30975a <=( (not A232)  and  A203 );
 a30976a <=( a30975a  and  a30972a );
 a30977a <=( a30976a  and  a30969a );
 a30980a <=( A234  and  A233 );
 a30983a <=( A298  and  A235 );
 a30984a <=( a30983a  and  a30980a );
 a30987a <=( (not A300)  and  (not A299) );
 a30990a <=( (not A302)  and  (not A301) );
 a30991a <=( a30990a  and  a30987a );
 a30992a <=( a30991a  and  a30984a );
 a30996a <=( A167  and  A168 );
 a30997a <=( A169  and  a30996a );
 a31000a <=( (not A201)  and  (not A166) );
 a31003a <=( (not A232)  and  A203 );
 a31004a <=( a31003a  and  a31000a );
 a31005a <=( a31004a  and  a30997a );
 a31008a <=( A234  and  A233 );
 a31011a <=( (not A298)  and  A235 );
 a31012a <=( a31011a  and  a31008a );
 a31015a <=( (not A300)  and  A299 );
 a31018a <=( (not A302)  and  (not A301) );
 a31019a <=( a31018a  and  a31015a );
 a31020a <=( a31019a  and  a31012a );
 a31024a <=( A167  and  A168 );
 a31025a <=( A169  and  a31024a );
 a31028a <=( (not A201)  and  (not A166) );
 a31031a <=( (not A232)  and  A203 );
 a31032a <=( a31031a  and  a31028a );
 a31033a <=( a31032a  and  a31025a );
 a31036a <=( A234  and  A233 );
 a31039a <=( (not A265)  and  A235 );
 a31040a <=( a31039a  and  a31036a );
 a31043a <=( (not A267)  and  A266 );
 a31046a <=( (not A269)  and  (not A268) );
 a31047a <=( a31046a  and  a31043a );
 a31048a <=( a31047a  and  a31040a );
 a31052a <=( A167  and  A168 );
 a31053a <=( A169  and  a31052a );
 a31056a <=( (not A201)  and  (not A166) );
 a31059a <=( (not A232)  and  A203 );
 a31060a <=( a31059a  and  a31056a );
 a31061a <=( a31060a  and  a31053a );
 a31064a <=( A234  and  A233 );
 a31067a <=( A265  and  A235 );
 a31068a <=( a31067a  and  a31064a );
 a31071a <=( (not A267)  and  (not A266) );
 a31074a <=( (not A269)  and  (not A268) );
 a31075a <=( a31074a  and  a31071a );
 a31076a <=( a31075a  and  a31068a );
 a31080a <=( A167  and  A168 );
 a31081a <=( A169  and  a31080a );
 a31084a <=( (not A201)  and  (not A166) );
 a31087a <=( (not A232)  and  A203 );
 a31088a <=( a31087a  and  a31084a );
 a31089a <=( a31088a  and  a31081a );
 a31092a <=( A234  and  A233 );
 a31095a <=( A298  and  A236 );
 a31096a <=( a31095a  and  a31092a );
 a31099a <=( (not A300)  and  (not A299) );
 a31102a <=( (not A302)  and  (not A301) );
 a31103a <=( a31102a  and  a31099a );
 a31104a <=( a31103a  and  a31096a );
 a31108a <=( A167  and  A168 );
 a31109a <=( A169  and  a31108a );
 a31112a <=( (not A201)  and  (not A166) );
 a31115a <=( (not A232)  and  A203 );
 a31116a <=( a31115a  and  a31112a );
 a31117a <=( a31116a  and  a31109a );
 a31120a <=( A234  and  A233 );
 a31123a <=( (not A298)  and  A236 );
 a31124a <=( a31123a  and  a31120a );
 a31127a <=( (not A300)  and  A299 );
 a31130a <=( (not A302)  and  (not A301) );
 a31131a <=( a31130a  and  a31127a );
 a31132a <=( a31131a  and  a31124a );
 a31136a <=( A167  and  A168 );
 a31137a <=( A169  and  a31136a );
 a31140a <=( (not A201)  and  (not A166) );
 a31143a <=( (not A232)  and  A203 );
 a31144a <=( a31143a  and  a31140a );
 a31145a <=( a31144a  and  a31137a );
 a31148a <=( A234  and  A233 );
 a31151a <=( (not A265)  and  A236 );
 a31152a <=( a31151a  and  a31148a );
 a31155a <=( (not A267)  and  A266 );
 a31158a <=( (not A269)  and  (not A268) );
 a31159a <=( a31158a  and  a31155a );
 a31160a <=( a31159a  and  a31152a );
 a31164a <=( A167  and  A168 );
 a31165a <=( A169  and  a31164a );
 a31168a <=( (not A201)  and  (not A166) );
 a31171a <=( (not A232)  and  A203 );
 a31172a <=( a31171a  and  a31168a );
 a31173a <=( a31172a  and  a31165a );
 a31176a <=( A234  and  A233 );
 a31179a <=( A265  and  A236 );
 a31180a <=( a31179a  and  a31176a );
 a31183a <=( (not A267)  and  (not A266) );
 a31186a <=( (not A269)  and  (not A268) );
 a31187a <=( a31186a  and  a31183a );
 a31188a <=( a31187a  and  a31180a );
 a31192a <=( A167  and  A168 );
 a31193a <=( A169  and  a31192a );
 a31196a <=( (not A201)  and  (not A166) );
 a31199a <=( (not A232)  and  A203 );
 a31200a <=( a31199a  and  a31196a );
 a31201a <=( a31200a  and  a31193a );
 a31204a <=( (not A234)  and  A233 );
 a31207a <=( (not A236)  and  (not A235) );
 a31208a <=( a31207a  and  a31204a );
 a31211a <=( (not A299)  and  A298 );
 a31214a <=( A301  and  A300 );
 a31215a <=( a31214a  and  a31211a );
 a31216a <=( a31215a  and  a31208a );
 a31220a <=( A167  and  A168 );
 a31221a <=( A169  and  a31220a );
 a31224a <=( (not A201)  and  (not A166) );
 a31227a <=( (not A232)  and  A203 );
 a31228a <=( a31227a  and  a31224a );
 a31229a <=( a31228a  and  a31221a );
 a31232a <=( (not A234)  and  A233 );
 a31235a <=( (not A236)  and  (not A235) );
 a31236a <=( a31235a  and  a31232a );
 a31239a <=( (not A299)  and  A298 );
 a31242a <=( A302  and  A300 );
 a31243a <=( a31242a  and  a31239a );
 a31244a <=( a31243a  and  a31236a );
 a31248a <=( A167  and  A168 );
 a31249a <=( A169  and  a31248a );
 a31252a <=( (not A201)  and  (not A166) );
 a31255a <=( (not A232)  and  A203 );
 a31256a <=( a31255a  and  a31252a );
 a31257a <=( a31256a  and  a31249a );
 a31260a <=( (not A234)  and  A233 );
 a31263a <=( (not A236)  and  (not A235) );
 a31264a <=( a31263a  and  a31260a );
 a31267a <=( A299  and  (not A298) );
 a31270a <=( A301  and  A300 );
 a31271a <=( a31270a  and  a31267a );
 a31272a <=( a31271a  and  a31264a );
 a31276a <=( A167  and  A168 );
 a31277a <=( A169  and  a31276a );
 a31280a <=( (not A201)  and  (not A166) );
 a31283a <=( (not A232)  and  A203 );
 a31284a <=( a31283a  and  a31280a );
 a31285a <=( a31284a  and  a31277a );
 a31288a <=( (not A234)  and  A233 );
 a31291a <=( (not A236)  and  (not A235) );
 a31292a <=( a31291a  and  a31288a );
 a31295a <=( A299  and  (not A298) );
 a31298a <=( A302  and  A300 );
 a31299a <=( a31298a  and  a31295a );
 a31300a <=( a31299a  and  a31292a );
 a31304a <=( A167  and  A168 );
 a31305a <=( A169  and  a31304a );
 a31308a <=( (not A201)  and  (not A166) );
 a31311a <=( (not A232)  and  A203 );
 a31312a <=( a31311a  and  a31308a );
 a31313a <=( a31312a  and  a31305a );
 a31316a <=( (not A234)  and  A233 );
 a31319a <=( (not A236)  and  (not A235) );
 a31320a <=( a31319a  and  a31316a );
 a31323a <=( A266  and  (not A265) );
 a31326a <=( A268  and  A267 );
 a31327a <=( a31326a  and  a31323a );
 a31328a <=( a31327a  and  a31320a );
 a31332a <=( A167  and  A168 );
 a31333a <=( A169  and  a31332a );
 a31336a <=( (not A201)  and  (not A166) );
 a31339a <=( (not A232)  and  A203 );
 a31340a <=( a31339a  and  a31336a );
 a31341a <=( a31340a  and  a31333a );
 a31344a <=( (not A234)  and  A233 );
 a31347a <=( (not A236)  and  (not A235) );
 a31348a <=( a31347a  and  a31344a );
 a31351a <=( A266  and  (not A265) );
 a31354a <=( A269  and  A267 );
 a31355a <=( a31354a  and  a31351a );
 a31356a <=( a31355a  and  a31348a );
 a31360a <=( A167  and  A168 );
 a31361a <=( A169  and  a31360a );
 a31364a <=( (not A201)  and  (not A166) );
 a31367a <=( (not A232)  and  A203 );
 a31368a <=( a31367a  and  a31364a );
 a31369a <=( a31368a  and  a31361a );
 a31372a <=( (not A234)  and  A233 );
 a31375a <=( (not A236)  and  (not A235) );
 a31376a <=( a31375a  and  a31372a );
 a31379a <=( (not A266)  and  A265 );
 a31382a <=( A268  and  A267 );
 a31383a <=( a31382a  and  a31379a );
 a31384a <=( a31383a  and  a31376a );
 a31388a <=( A167  and  A168 );
 a31389a <=( A169  and  a31388a );
 a31392a <=( (not A201)  and  (not A166) );
 a31395a <=( (not A232)  and  A203 );
 a31396a <=( a31395a  and  a31392a );
 a31397a <=( a31396a  and  a31389a );
 a31400a <=( (not A234)  and  A233 );
 a31403a <=( (not A236)  and  (not A235) );
 a31404a <=( a31403a  and  a31400a );
 a31407a <=( (not A266)  and  A265 );
 a31410a <=( A269  and  A267 );
 a31411a <=( a31410a  and  a31407a );
 a31412a <=( a31411a  and  a31404a );
 a31416a <=( A167  and  A168 );
 a31417a <=( A169  and  a31416a );
 a31420a <=( (not A201)  and  (not A166) );
 a31423a <=( A232  and  A203 );
 a31424a <=( a31423a  and  a31420a );
 a31425a <=( a31424a  and  a31417a );
 a31428a <=( A234  and  (not A233) );
 a31431a <=( A298  and  A235 );
 a31432a <=( a31431a  and  a31428a );
 a31435a <=( (not A300)  and  (not A299) );
 a31438a <=( (not A302)  and  (not A301) );
 a31439a <=( a31438a  and  a31435a );
 a31440a <=( a31439a  and  a31432a );
 a31444a <=( A167  and  A168 );
 a31445a <=( A169  and  a31444a );
 a31448a <=( (not A201)  and  (not A166) );
 a31451a <=( A232  and  A203 );
 a31452a <=( a31451a  and  a31448a );
 a31453a <=( a31452a  and  a31445a );
 a31456a <=( A234  and  (not A233) );
 a31459a <=( (not A298)  and  A235 );
 a31460a <=( a31459a  and  a31456a );
 a31463a <=( (not A300)  and  A299 );
 a31466a <=( (not A302)  and  (not A301) );
 a31467a <=( a31466a  and  a31463a );
 a31468a <=( a31467a  and  a31460a );
 a31472a <=( A167  and  A168 );
 a31473a <=( A169  and  a31472a );
 a31476a <=( (not A201)  and  (not A166) );
 a31479a <=( A232  and  A203 );
 a31480a <=( a31479a  and  a31476a );
 a31481a <=( a31480a  and  a31473a );
 a31484a <=( A234  and  (not A233) );
 a31487a <=( (not A265)  and  A235 );
 a31488a <=( a31487a  and  a31484a );
 a31491a <=( (not A267)  and  A266 );
 a31494a <=( (not A269)  and  (not A268) );
 a31495a <=( a31494a  and  a31491a );
 a31496a <=( a31495a  and  a31488a );
 a31500a <=( A167  and  A168 );
 a31501a <=( A169  and  a31500a );
 a31504a <=( (not A201)  and  (not A166) );
 a31507a <=( A232  and  A203 );
 a31508a <=( a31507a  and  a31504a );
 a31509a <=( a31508a  and  a31501a );
 a31512a <=( A234  and  (not A233) );
 a31515a <=( A265  and  A235 );
 a31516a <=( a31515a  and  a31512a );
 a31519a <=( (not A267)  and  (not A266) );
 a31522a <=( (not A269)  and  (not A268) );
 a31523a <=( a31522a  and  a31519a );
 a31524a <=( a31523a  and  a31516a );
 a31528a <=( A167  and  A168 );
 a31529a <=( A169  and  a31528a );
 a31532a <=( (not A201)  and  (not A166) );
 a31535a <=( A232  and  A203 );
 a31536a <=( a31535a  and  a31532a );
 a31537a <=( a31536a  and  a31529a );
 a31540a <=( A234  and  (not A233) );
 a31543a <=( A298  and  A236 );
 a31544a <=( a31543a  and  a31540a );
 a31547a <=( (not A300)  and  (not A299) );
 a31550a <=( (not A302)  and  (not A301) );
 a31551a <=( a31550a  and  a31547a );
 a31552a <=( a31551a  and  a31544a );
 a31556a <=( A167  and  A168 );
 a31557a <=( A169  and  a31556a );
 a31560a <=( (not A201)  and  (not A166) );
 a31563a <=( A232  and  A203 );
 a31564a <=( a31563a  and  a31560a );
 a31565a <=( a31564a  and  a31557a );
 a31568a <=( A234  and  (not A233) );
 a31571a <=( (not A298)  and  A236 );
 a31572a <=( a31571a  and  a31568a );
 a31575a <=( (not A300)  and  A299 );
 a31578a <=( (not A302)  and  (not A301) );
 a31579a <=( a31578a  and  a31575a );
 a31580a <=( a31579a  and  a31572a );
 a31584a <=( A167  and  A168 );
 a31585a <=( A169  and  a31584a );
 a31588a <=( (not A201)  and  (not A166) );
 a31591a <=( A232  and  A203 );
 a31592a <=( a31591a  and  a31588a );
 a31593a <=( a31592a  and  a31585a );
 a31596a <=( A234  and  (not A233) );
 a31599a <=( (not A265)  and  A236 );
 a31600a <=( a31599a  and  a31596a );
 a31603a <=( (not A267)  and  A266 );
 a31606a <=( (not A269)  and  (not A268) );
 a31607a <=( a31606a  and  a31603a );
 a31608a <=( a31607a  and  a31600a );
 a31612a <=( A167  and  A168 );
 a31613a <=( A169  and  a31612a );
 a31616a <=( (not A201)  and  (not A166) );
 a31619a <=( A232  and  A203 );
 a31620a <=( a31619a  and  a31616a );
 a31621a <=( a31620a  and  a31613a );
 a31624a <=( A234  and  (not A233) );
 a31627a <=( A265  and  A236 );
 a31628a <=( a31627a  and  a31624a );
 a31631a <=( (not A267)  and  (not A266) );
 a31634a <=( (not A269)  and  (not A268) );
 a31635a <=( a31634a  and  a31631a );
 a31636a <=( a31635a  and  a31628a );
 a31640a <=( A167  and  A168 );
 a31641a <=( A169  and  a31640a );
 a31644a <=( (not A201)  and  (not A166) );
 a31647a <=( A232  and  A203 );
 a31648a <=( a31647a  and  a31644a );
 a31649a <=( a31648a  and  a31641a );
 a31652a <=( (not A234)  and  (not A233) );
 a31655a <=( (not A236)  and  (not A235) );
 a31656a <=( a31655a  and  a31652a );
 a31659a <=( (not A299)  and  A298 );
 a31662a <=( A301  and  A300 );
 a31663a <=( a31662a  and  a31659a );
 a31664a <=( a31663a  and  a31656a );
 a31668a <=( A167  and  A168 );
 a31669a <=( A169  and  a31668a );
 a31672a <=( (not A201)  and  (not A166) );
 a31675a <=( A232  and  A203 );
 a31676a <=( a31675a  and  a31672a );
 a31677a <=( a31676a  and  a31669a );
 a31680a <=( (not A234)  and  (not A233) );
 a31683a <=( (not A236)  and  (not A235) );
 a31684a <=( a31683a  and  a31680a );
 a31687a <=( (not A299)  and  A298 );
 a31690a <=( A302  and  A300 );
 a31691a <=( a31690a  and  a31687a );
 a31692a <=( a31691a  and  a31684a );
 a31696a <=( A167  and  A168 );
 a31697a <=( A169  and  a31696a );
 a31700a <=( (not A201)  and  (not A166) );
 a31703a <=( A232  and  A203 );
 a31704a <=( a31703a  and  a31700a );
 a31705a <=( a31704a  and  a31697a );
 a31708a <=( (not A234)  and  (not A233) );
 a31711a <=( (not A236)  and  (not A235) );
 a31712a <=( a31711a  and  a31708a );
 a31715a <=( A299  and  (not A298) );
 a31718a <=( A301  and  A300 );
 a31719a <=( a31718a  and  a31715a );
 a31720a <=( a31719a  and  a31712a );
 a31724a <=( A167  and  A168 );
 a31725a <=( A169  and  a31724a );
 a31728a <=( (not A201)  and  (not A166) );
 a31731a <=( A232  and  A203 );
 a31732a <=( a31731a  and  a31728a );
 a31733a <=( a31732a  and  a31725a );
 a31736a <=( (not A234)  and  (not A233) );
 a31739a <=( (not A236)  and  (not A235) );
 a31740a <=( a31739a  and  a31736a );
 a31743a <=( A299  and  (not A298) );
 a31746a <=( A302  and  A300 );
 a31747a <=( a31746a  and  a31743a );
 a31748a <=( a31747a  and  a31740a );
 a31752a <=( A167  and  A168 );
 a31753a <=( A169  and  a31752a );
 a31756a <=( (not A201)  and  (not A166) );
 a31759a <=( A232  and  A203 );
 a31760a <=( a31759a  and  a31756a );
 a31761a <=( a31760a  and  a31753a );
 a31764a <=( (not A234)  and  (not A233) );
 a31767a <=( (not A236)  and  (not A235) );
 a31768a <=( a31767a  and  a31764a );
 a31771a <=( A266  and  (not A265) );
 a31774a <=( A268  and  A267 );
 a31775a <=( a31774a  and  a31771a );
 a31776a <=( a31775a  and  a31768a );
 a31780a <=( A167  and  A168 );
 a31781a <=( A169  and  a31780a );
 a31784a <=( (not A201)  and  (not A166) );
 a31787a <=( A232  and  A203 );
 a31788a <=( a31787a  and  a31784a );
 a31789a <=( a31788a  and  a31781a );
 a31792a <=( (not A234)  and  (not A233) );
 a31795a <=( (not A236)  and  (not A235) );
 a31796a <=( a31795a  and  a31792a );
 a31799a <=( A266  and  (not A265) );
 a31802a <=( A269  and  A267 );
 a31803a <=( a31802a  and  a31799a );
 a31804a <=( a31803a  and  a31796a );
 a31808a <=( A167  and  A168 );
 a31809a <=( A169  and  a31808a );
 a31812a <=( (not A201)  and  (not A166) );
 a31815a <=( A232  and  A203 );
 a31816a <=( a31815a  and  a31812a );
 a31817a <=( a31816a  and  a31809a );
 a31820a <=( (not A234)  and  (not A233) );
 a31823a <=( (not A236)  and  (not A235) );
 a31824a <=( a31823a  and  a31820a );
 a31827a <=( (not A266)  and  A265 );
 a31830a <=( A268  and  A267 );
 a31831a <=( a31830a  and  a31827a );
 a31832a <=( a31831a  and  a31824a );
 a31836a <=( A167  and  A168 );
 a31837a <=( A169  and  a31836a );
 a31840a <=( (not A201)  and  (not A166) );
 a31843a <=( A232  and  A203 );
 a31844a <=( a31843a  and  a31840a );
 a31845a <=( a31844a  and  a31837a );
 a31848a <=( (not A234)  and  (not A233) );
 a31851a <=( (not A236)  and  (not A235) );
 a31852a <=( a31851a  and  a31848a );
 a31855a <=( (not A266)  and  A265 );
 a31858a <=( A269  and  A267 );
 a31859a <=( a31858a  and  a31855a );
 a31860a <=( a31859a  and  a31852a );
 a31864a <=( A167  and  A168 );
 a31865a <=( A169  and  a31864a );
 a31868a <=( A199  and  (not A166) );
 a31871a <=( (not A232)  and  A200 );
 a31872a <=( a31871a  and  a31868a );
 a31873a <=( a31872a  and  a31865a );
 a31876a <=( A234  and  A233 );
 a31879a <=( A298  and  A235 );
 a31880a <=( a31879a  and  a31876a );
 a31883a <=( (not A300)  and  (not A299) );
 a31886a <=( (not A302)  and  (not A301) );
 a31887a <=( a31886a  and  a31883a );
 a31888a <=( a31887a  and  a31880a );
 a31892a <=( A167  and  A168 );
 a31893a <=( A169  and  a31892a );
 a31896a <=( A199  and  (not A166) );
 a31899a <=( (not A232)  and  A200 );
 a31900a <=( a31899a  and  a31896a );
 a31901a <=( a31900a  and  a31893a );
 a31904a <=( A234  and  A233 );
 a31907a <=( (not A298)  and  A235 );
 a31908a <=( a31907a  and  a31904a );
 a31911a <=( (not A300)  and  A299 );
 a31914a <=( (not A302)  and  (not A301) );
 a31915a <=( a31914a  and  a31911a );
 a31916a <=( a31915a  and  a31908a );
 a31920a <=( A167  and  A168 );
 a31921a <=( A169  and  a31920a );
 a31924a <=( A199  and  (not A166) );
 a31927a <=( (not A232)  and  A200 );
 a31928a <=( a31927a  and  a31924a );
 a31929a <=( a31928a  and  a31921a );
 a31932a <=( A234  and  A233 );
 a31935a <=( (not A265)  and  A235 );
 a31936a <=( a31935a  and  a31932a );
 a31939a <=( (not A267)  and  A266 );
 a31942a <=( (not A269)  and  (not A268) );
 a31943a <=( a31942a  and  a31939a );
 a31944a <=( a31943a  and  a31936a );
 a31948a <=( A167  and  A168 );
 a31949a <=( A169  and  a31948a );
 a31952a <=( A199  and  (not A166) );
 a31955a <=( (not A232)  and  A200 );
 a31956a <=( a31955a  and  a31952a );
 a31957a <=( a31956a  and  a31949a );
 a31960a <=( A234  and  A233 );
 a31963a <=( A265  and  A235 );
 a31964a <=( a31963a  and  a31960a );
 a31967a <=( (not A267)  and  (not A266) );
 a31970a <=( (not A269)  and  (not A268) );
 a31971a <=( a31970a  and  a31967a );
 a31972a <=( a31971a  and  a31964a );
 a31976a <=( A167  and  A168 );
 a31977a <=( A169  and  a31976a );
 a31980a <=( A199  and  (not A166) );
 a31983a <=( (not A232)  and  A200 );
 a31984a <=( a31983a  and  a31980a );
 a31985a <=( a31984a  and  a31977a );
 a31988a <=( A234  and  A233 );
 a31991a <=( A298  and  A236 );
 a31992a <=( a31991a  and  a31988a );
 a31995a <=( (not A300)  and  (not A299) );
 a31998a <=( (not A302)  and  (not A301) );
 a31999a <=( a31998a  and  a31995a );
 a32000a <=( a31999a  and  a31992a );
 a32004a <=( A167  and  A168 );
 a32005a <=( A169  and  a32004a );
 a32008a <=( A199  and  (not A166) );
 a32011a <=( (not A232)  and  A200 );
 a32012a <=( a32011a  and  a32008a );
 a32013a <=( a32012a  and  a32005a );
 a32016a <=( A234  and  A233 );
 a32019a <=( (not A298)  and  A236 );
 a32020a <=( a32019a  and  a32016a );
 a32023a <=( (not A300)  and  A299 );
 a32026a <=( (not A302)  and  (not A301) );
 a32027a <=( a32026a  and  a32023a );
 a32028a <=( a32027a  and  a32020a );
 a32032a <=( A167  and  A168 );
 a32033a <=( A169  and  a32032a );
 a32036a <=( A199  and  (not A166) );
 a32039a <=( (not A232)  and  A200 );
 a32040a <=( a32039a  and  a32036a );
 a32041a <=( a32040a  and  a32033a );
 a32044a <=( A234  and  A233 );
 a32047a <=( (not A265)  and  A236 );
 a32048a <=( a32047a  and  a32044a );
 a32051a <=( (not A267)  and  A266 );
 a32054a <=( (not A269)  and  (not A268) );
 a32055a <=( a32054a  and  a32051a );
 a32056a <=( a32055a  and  a32048a );
 a32060a <=( A167  and  A168 );
 a32061a <=( A169  and  a32060a );
 a32064a <=( A199  and  (not A166) );
 a32067a <=( (not A232)  and  A200 );
 a32068a <=( a32067a  and  a32064a );
 a32069a <=( a32068a  and  a32061a );
 a32072a <=( A234  and  A233 );
 a32075a <=( A265  and  A236 );
 a32076a <=( a32075a  and  a32072a );
 a32079a <=( (not A267)  and  (not A266) );
 a32082a <=( (not A269)  and  (not A268) );
 a32083a <=( a32082a  and  a32079a );
 a32084a <=( a32083a  and  a32076a );
 a32088a <=( A167  and  A168 );
 a32089a <=( A169  and  a32088a );
 a32092a <=( A199  and  (not A166) );
 a32095a <=( (not A232)  and  A200 );
 a32096a <=( a32095a  and  a32092a );
 a32097a <=( a32096a  and  a32089a );
 a32100a <=( (not A234)  and  A233 );
 a32103a <=( (not A236)  and  (not A235) );
 a32104a <=( a32103a  and  a32100a );
 a32107a <=( (not A299)  and  A298 );
 a32110a <=( A301  and  A300 );
 a32111a <=( a32110a  and  a32107a );
 a32112a <=( a32111a  and  a32104a );
 a32116a <=( A167  and  A168 );
 a32117a <=( A169  and  a32116a );
 a32120a <=( A199  and  (not A166) );
 a32123a <=( (not A232)  and  A200 );
 a32124a <=( a32123a  and  a32120a );
 a32125a <=( a32124a  and  a32117a );
 a32128a <=( (not A234)  and  A233 );
 a32131a <=( (not A236)  and  (not A235) );
 a32132a <=( a32131a  and  a32128a );
 a32135a <=( (not A299)  and  A298 );
 a32138a <=( A302  and  A300 );
 a32139a <=( a32138a  and  a32135a );
 a32140a <=( a32139a  and  a32132a );
 a32144a <=( A167  and  A168 );
 a32145a <=( A169  and  a32144a );
 a32148a <=( A199  and  (not A166) );
 a32151a <=( (not A232)  and  A200 );
 a32152a <=( a32151a  and  a32148a );
 a32153a <=( a32152a  and  a32145a );
 a32156a <=( (not A234)  and  A233 );
 a32159a <=( (not A236)  and  (not A235) );
 a32160a <=( a32159a  and  a32156a );
 a32163a <=( A299  and  (not A298) );
 a32166a <=( A301  and  A300 );
 a32167a <=( a32166a  and  a32163a );
 a32168a <=( a32167a  and  a32160a );
 a32172a <=( A167  and  A168 );
 a32173a <=( A169  and  a32172a );
 a32176a <=( A199  and  (not A166) );
 a32179a <=( (not A232)  and  A200 );
 a32180a <=( a32179a  and  a32176a );
 a32181a <=( a32180a  and  a32173a );
 a32184a <=( (not A234)  and  A233 );
 a32187a <=( (not A236)  and  (not A235) );
 a32188a <=( a32187a  and  a32184a );
 a32191a <=( A299  and  (not A298) );
 a32194a <=( A302  and  A300 );
 a32195a <=( a32194a  and  a32191a );
 a32196a <=( a32195a  and  a32188a );
 a32200a <=( A167  and  A168 );
 a32201a <=( A169  and  a32200a );
 a32204a <=( A199  and  (not A166) );
 a32207a <=( (not A232)  and  A200 );
 a32208a <=( a32207a  and  a32204a );
 a32209a <=( a32208a  and  a32201a );
 a32212a <=( (not A234)  and  A233 );
 a32215a <=( (not A236)  and  (not A235) );
 a32216a <=( a32215a  and  a32212a );
 a32219a <=( A266  and  (not A265) );
 a32222a <=( A268  and  A267 );
 a32223a <=( a32222a  and  a32219a );
 a32224a <=( a32223a  and  a32216a );
 a32228a <=( A167  and  A168 );
 a32229a <=( A169  and  a32228a );
 a32232a <=( A199  and  (not A166) );
 a32235a <=( (not A232)  and  A200 );
 a32236a <=( a32235a  and  a32232a );
 a32237a <=( a32236a  and  a32229a );
 a32240a <=( (not A234)  and  A233 );
 a32243a <=( (not A236)  and  (not A235) );
 a32244a <=( a32243a  and  a32240a );
 a32247a <=( A266  and  (not A265) );
 a32250a <=( A269  and  A267 );
 a32251a <=( a32250a  and  a32247a );
 a32252a <=( a32251a  and  a32244a );
 a32256a <=( A167  and  A168 );
 a32257a <=( A169  and  a32256a );
 a32260a <=( A199  and  (not A166) );
 a32263a <=( (not A232)  and  A200 );
 a32264a <=( a32263a  and  a32260a );
 a32265a <=( a32264a  and  a32257a );
 a32268a <=( (not A234)  and  A233 );
 a32271a <=( (not A236)  and  (not A235) );
 a32272a <=( a32271a  and  a32268a );
 a32275a <=( (not A266)  and  A265 );
 a32278a <=( A268  and  A267 );
 a32279a <=( a32278a  and  a32275a );
 a32280a <=( a32279a  and  a32272a );
 a32284a <=( A167  and  A168 );
 a32285a <=( A169  and  a32284a );
 a32288a <=( A199  and  (not A166) );
 a32291a <=( (not A232)  and  A200 );
 a32292a <=( a32291a  and  a32288a );
 a32293a <=( a32292a  and  a32285a );
 a32296a <=( (not A234)  and  A233 );
 a32299a <=( (not A236)  and  (not A235) );
 a32300a <=( a32299a  and  a32296a );
 a32303a <=( (not A266)  and  A265 );
 a32306a <=( A269  and  A267 );
 a32307a <=( a32306a  and  a32303a );
 a32308a <=( a32307a  and  a32300a );
 a32312a <=( A167  and  A168 );
 a32313a <=( A169  and  a32312a );
 a32316a <=( A199  and  (not A166) );
 a32319a <=( A232  and  A200 );
 a32320a <=( a32319a  and  a32316a );
 a32321a <=( a32320a  and  a32313a );
 a32324a <=( A234  and  (not A233) );
 a32327a <=( A298  and  A235 );
 a32328a <=( a32327a  and  a32324a );
 a32331a <=( (not A300)  and  (not A299) );
 a32334a <=( (not A302)  and  (not A301) );
 a32335a <=( a32334a  and  a32331a );
 a32336a <=( a32335a  and  a32328a );
 a32340a <=( A167  and  A168 );
 a32341a <=( A169  and  a32340a );
 a32344a <=( A199  and  (not A166) );
 a32347a <=( A232  and  A200 );
 a32348a <=( a32347a  and  a32344a );
 a32349a <=( a32348a  and  a32341a );
 a32352a <=( A234  and  (not A233) );
 a32355a <=( (not A298)  and  A235 );
 a32356a <=( a32355a  and  a32352a );
 a32359a <=( (not A300)  and  A299 );
 a32362a <=( (not A302)  and  (not A301) );
 a32363a <=( a32362a  and  a32359a );
 a32364a <=( a32363a  and  a32356a );
 a32368a <=( A167  and  A168 );
 a32369a <=( A169  and  a32368a );
 a32372a <=( A199  and  (not A166) );
 a32375a <=( A232  and  A200 );
 a32376a <=( a32375a  and  a32372a );
 a32377a <=( a32376a  and  a32369a );
 a32380a <=( A234  and  (not A233) );
 a32383a <=( (not A265)  and  A235 );
 a32384a <=( a32383a  and  a32380a );
 a32387a <=( (not A267)  and  A266 );
 a32390a <=( (not A269)  and  (not A268) );
 a32391a <=( a32390a  and  a32387a );
 a32392a <=( a32391a  and  a32384a );
 a32396a <=( A167  and  A168 );
 a32397a <=( A169  and  a32396a );
 a32400a <=( A199  and  (not A166) );
 a32403a <=( A232  and  A200 );
 a32404a <=( a32403a  and  a32400a );
 a32405a <=( a32404a  and  a32397a );
 a32408a <=( A234  and  (not A233) );
 a32411a <=( A265  and  A235 );
 a32412a <=( a32411a  and  a32408a );
 a32415a <=( (not A267)  and  (not A266) );
 a32418a <=( (not A269)  and  (not A268) );
 a32419a <=( a32418a  and  a32415a );
 a32420a <=( a32419a  and  a32412a );
 a32424a <=( A167  and  A168 );
 a32425a <=( A169  and  a32424a );
 a32428a <=( A199  and  (not A166) );
 a32431a <=( A232  and  A200 );
 a32432a <=( a32431a  and  a32428a );
 a32433a <=( a32432a  and  a32425a );
 a32436a <=( A234  and  (not A233) );
 a32439a <=( A298  and  A236 );
 a32440a <=( a32439a  and  a32436a );
 a32443a <=( (not A300)  and  (not A299) );
 a32446a <=( (not A302)  and  (not A301) );
 a32447a <=( a32446a  and  a32443a );
 a32448a <=( a32447a  and  a32440a );
 a32452a <=( A167  and  A168 );
 a32453a <=( A169  and  a32452a );
 a32456a <=( A199  and  (not A166) );
 a32459a <=( A232  and  A200 );
 a32460a <=( a32459a  and  a32456a );
 a32461a <=( a32460a  and  a32453a );
 a32464a <=( A234  and  (not A233) );
 a32467a <=( (not A298)  and  A236 );
 a32468a <=( a32467a  and  a32464a );
 a32471a <=( (not A300)  and  A299 );
 a32474a <=( (not A302)  and  (not A301) );
 a32475a <=( a32474a  and  a32471a );
 a32476a <=( a32475a  and  a32468a );
 a32480a <=( A167  and  A168 );
 a32481a <=( A169  and  a32480a );
 a32484a <=( A199  and  (not A166) );
 a32487a <=( A232  and  A200 );
 a32488a <=( a32487a  and  a32484a );
 a32489a <=( a32488a  and  a32481a );
 a32492a <=( A234  and  (not A233) );
 a32495a <=( (not A265)  and  A236 );
 a32496a <=( a32495a  and  a32492a );
 a32499a <=( (not A267)  and  A266 );
 a32502a <=( (not A269)  and  (not A268) );
 a32503a <=( a32502a  and  a32499a );
 a32504a <=( a32503a  and  a32496a );
 a32508a <=( A167  and  A168 );
 a32509a <=( A169  and  a32508a );
 a32512a <=( A199  and  (not A166) );
 a32515a <=( A232  and  A200 );
 a32516a <=( a32515a  and  a32512a );
 a32517a <=( a32516a  and  a32509a );
 a32520a <=( A234  and  (not A233) );
 a32523a <=( A265  and  A236 );
 a32524a <=( a32523a  and  a32520a );
 a32527a <=( (not A267)  and  (not A266) );
 a32530a <=( (not A269)  and  (not A268) );
 a32531a <=( a32530a  and  a32527a );
 a32532a <=( a32531a  and  a32524a );
 a32536a <=( A167  and  A168 );
 a32537a <=( A169  and  a32536a );
 a32540a <=( A199  and  (not A166) );
 a32543a <=( A232  and  A200 );
 a32544a <=( a32543a  and  a32540a );
 a32545a <=( a32544a  and  a32537a );
 a32548a <=( (not A234)  and  (not A233) );
 a32551a <=( (not A236)  and  (not A235) );
 a32552a <=( a32551a  and  a32548a );
 a32555a <=( (not A299)  and  A298 );
 a32558a <=( A301  and  A300 );
 a32559a <=( a32558a  and  a32555a );
 a32560a <=( a32559a  and  a32552a );
 a32564a <=( A167  and  A168 );
 a32565a <=( A169  and  a32564a );
 a32568a <=( A199  and  (not A166) );
 a32571a <=( A232  and  A200 );
 a32572a <=( a32571a  and  a32568a );
 a32573a <=( a32572a  and  a32565a );
 a32576a <=( (not A234)  and  (not A233) );
 a32579a <=( (not A236)  and  (not A235) );
 a32580a <=( a32579a  and  a32576a );
 a32583a <=( (not A299)  and  A298 );
 a32586a <=( A302  and  A300 );
 a32587a <=( a32586a  and  a32583a );
 a32588a <=( a32587a  and  a32580a );
 a32592a <=( A167  and  A168 );
 a32593a <=( A169  and  a32592a );
 a32596a <=( A199  and  (not A166) );
 a32599a <=( A232  and  A200 );
 a32600a <=( a32599a  and  a32596a );
 a32601a <=( a32600a  and  a32593a );
 a32604a <=( (not A234)  and  (not A233) );
 a32607a <=( (not A236)  and  (not A235) );
 a32608a <=( a32607a  and  a32604a );
 a32611a <=( A299  and  (not A298) );
 a32614a <=( A301  and  A300 );
 a32615a <=( a32614a  and  a32611a );
 a32616a <=( a32615a  and  a32608a );
 a32620a <=( A167  and  A168 );
 a32621a <=( A169  and  a32620a );
 a32624a <=( A199  and  (not A166) );
 a32627a <=( A232  and  A200 );
 a32628a <=( a32627a  and  a32624a );
 a32629a <=( a32628a  and  a32621a );
 a32632a <=( (not A234)  and  (not A233) );
 a32635a <=( (not A236)  and  (not A235) );
 a32636a <=( a32635a  and  a32632a );
 a32639a <=( A299  and  (not A298) );
 a32642a <=( A302  and  A300 );
 a32643a <=( a32642a  and  a32639a );
 a32644a <=( a32643a  and  a32636a );
 a32648a <=( A167  and  A168 );
 a32649a <=( A169  and  a32648a );
 a32652a <=( A199  and  (not A166) );
 a32655a <=( A232  and  A200 );
 a32656a <=( a32655a  and  a32652a );
 a32657a <=( a32656a  and  a32649a );
 a32660a <=( (not A234)  and  (not A233) );
 a32663a <=( (not A236)  and  (not A235) );
 a32664a <=( a32663a  and  a32660a );
 a32667a <=( A266  and  (not A265) );
 a32670a <=( A268  and  A267 );
 a32671a <=( a32670a  and  a32667a );
 a32672a <=( a32671a  and  a32664a );
 a32676a <=( A167  and  A168 );
 a32677a <=( A169  and  a32676a );
 a32680a <=( A199  and  (not A166) );
 a32683a <=( A232  and  A200 );
 a32684a <=( a32683a  and  a32680a );
 a32685a <=( a32684a  and  a32677a );
 a32688a <=( (not A234)  and  (not A233) );
 a32691a <=( (not A236)  and  (not A235) );
 a32692a <=( a32691a  and  a32688a );
 a32695a <=( A266  and  (not A265) );
 a32698a <=( A269  and  A267 );
 a32699a <=( a32698a  and  a32695a );
 a32700a <=( a32699a  and  a32692a );
 a32704a <=( A167  and  A168 );
 a32705a <=( A169  and  a32704a );
 a32708a <=( A199  and  (not A166) );
 a32711a <=( A232  and  A200 );
 a32712a <=( a32711a  and  a32708a );
 a32713a <=( a32712a  and  a32705a );
 a32716a <=( (not A234)  and  (not A233) );
 a32719a <=( (not A236)  and  (not A235) );
 a32720a <=( a32719a  and  a32716a );
 a32723a <=( (not A266)  and  A265 );
 a32726a <=( A268  and  A267 );
 a32727a <=( a32726a  and  a32723a );
 a32728a <=( a32727a  and  a32720a );
 a32732a <=( A167  and  A168 );
 a32733a <=( A169  and  a32732a );
 a32736a <=( A199  and  (not A166) );
 a32739a <=( A232  and  A200 );
 a32740a <=( a32739a  and  a32736a );
 a32741a <=( a32740a  and  a32733a );
 a32744a <=( (not A234)  and  (not A233) );
 a32747a <=( (not A236)  and  (not A235) );
 a32748a <=( a32747a  and  a32744a );
 a32751a <=( (not A266)  and  A265 );
 a32754a <=( A269  and  A267 );
 a32755a <=( a32754a  and  a32751a );
 a32756a <=( a32755a  and  a32748a );
 a32760a <=( A167  and  A168 );
 a32761a <=( A169  and  a32760a );
 a32764a <=( (not A199)  and  (not A166) );
 a32767a <=( (not A232)  and  (not A200) );
 a32768a <=( a32767a  and  a32764a );
 a32769a <=( a32768a  and  a32761a );
 a32772a <=( A234  and  A233 );
 a32775a <=( A298  and  A235 );
 a32776a <=( a32775a  and  a32772a );
 a32779a <=( (not A300)  and  (not A299) );
 a32782a <=( (not A302)  and  (not A301) );
 a32783a <=( a32782a  and  a32779a );
 a32784a <=( a32783a  and  a32776a );
 a32788a <=( A167  and  A168 );
 a32789a <=( A169  and  a32788a );
 a32792a <=( (not A199)  and  (not A166) );
 a32795a <=( (not A232)  and  (not A200) );
 a32796a <=( a32795a  and  a32792a );
 a32797a <=( a32796a  and  a32789a );
 a32800a <=( A234  and  A233 );
 a32803a <=( (not A298)  and  A235 );
 a32804a <=( a32803a  and  a32800a );
 a32807a <=( (not A300)  and  A299 );
 a32810a <=( (not A302)  and  (not A301) );
 a32811a <=( a32810a  and  a32807a );
 a32812a <=( a32811a  and  a32804a );
 a32816a <=( A167  and  A168 );
 a32817a <=( A169  and  a32816a );
 a32820a <=( (not A199)  and  (not A166) );
 a32823a <=( (not A232)  and  (not A200) );
 a32824a <=( a32823a  and  a32820a );
 a32825a <=( a32824a  and  a32817a );
 a32828a <=( A234  and  A233 );
 a32831a <=( (not A265)  and  A235 );
 a32832a <=( a32831a  and  a32828a );
 a32835a <=( (not A267)  and  A266 );
 a32838a <=( (not A269)  and  (not A268) );
 a32839a <=( a32838a  and  a32835a );
 a32840a <=( a32839a  and  a32832a );
 a32844a <=( A167  and  A168 );
 a32845a <=( A169  and  a32844a );
 a32848a <=( (not A199)  and  (not A166) );
 a32851a <=( (not A232)  and  (not A200) );
 a32852a <=( a32851a  and  a32848a );
 a32853a <=( a32852a  and  a32845a );
 a32856a <=( A234  and  A233 );
 a32859a <=( A265  and  A235 );
 a32860a <=( a32859a  and  a32856a );
 a32863a <=( (not A267)  and  (not A266) );
 a32866a <=( (not A269)  and  (not A268) );
 a32867a <=( a32866a  and  a32863a );
 a32868a <=( a32867a  and  a32860a );
 a32872a <=( A167  and  A168 );
 a32873a <=( A169  and  a32872a );
 a32876a <=( (not A199)  and  (not A166) );
 a32879a <=( (not A232)  and  (not A200) );
 a32880a <=( a32879a  and  a32876a );
 a32881a <=( a32880a  and  a32873a );
 a32884a <=( A234  and  A233 );
 a32887a <=( A298  and  A236 );
 a32888a <=( a32887a  and  a32884a );
 a32891a <=( (not A300)  and  (not A299) );
 a32894a <=( (not A302)  and  (not A301) );
 a32895a <=( a32894a  and  a32891a );
 a32896a <=( a32895a  and  a32888a );
 a32900a <=( A167  and  A168 );
 a32901a <=( A169  and  a32900a );
 a32904a <=( (not A199)  and  (not A166) );
 a32907a <=( (not A232)  and  (not A200) );
 a32908a <=( a32907a  and  a32904a );
 a32909a <=( a32908a  and  a32901a );
 a32912a <=( A234  and  A233 );
 a32915a <=( (not A298)  and  A236 );
 a32916a <=( a32915a  and  a32912a );
 a32919a <=( (not A300)  and  A299 );
 a32922a <=( (not A302)  and  (not A301) );
 a32923a <=( a32922a  and  a32919a );
 a32924a <=( a32923a  and  a32916a );
 a32928a <=( A167  and  A168 );
 a32929a <=( A169  and  a32928a );
 a32932a <=( (not A199)  and  (not A166) );
 a32935a <=( (not A232)  and  (not A200) );
 a32936a <=( a32935a  and  a32932a );
 a32937a <=( a32936a  and  a32929a );
 a32940a <=( A234  and  A233 );
 a32943a <=( (not A265)  and  A236 );
 a32944a <=( a32943a  and  a32940a );
 a32947a <=( (not A267)  and  A266 );
 a32950a <=( (not A269)  and  (not A268) );
 a32951a <=( a32950a  and  a32947a );
 a32952a <=( a32951a  and  a32944a );
 a32956a <=( A167  and  A168 );
 a32957a <=( A169  and  a32956a );
 a32960a <=( (not A199)  and  (not A166) );
 a32963a <=( (not A232)  and  (not A200) );
 a32964a <=( a32963a  and  a32960a );
 a32965a <=( a32964a  and  a32957a );
 a32968a <=( A234  and  A233 );
 a32971a <=( A265  and  A236 );
 a32972a <=( a32971a  and  a32968a );
 a32975a <=( (not A267)  and  (not A266) );
 a32978a <=( (not A269)  and  (not A268) );
 a32979a <=( a32978a  and  a32975a );
 a32980a <=( a32979a  and  a32972a );
 a32984a <=( A167  and  A168 );
 a32985a <=( A169  and  a32984a );
 a32988a <=( (not A199)  and  (not A166) );
 a32991a <=( (not A232)  and  (not A200) );
 a32992a <=( a32991a  and  a32988a );
 a32993a <=( a32992a  and  a32985a );
 a32996a <=( (not A234)  and  A233 );
 a32999a <=( (not A236)  and  (not A235) );
 a33000a <=( a32999a  and  a32996a );
 a33003a <=( (not A299)  and  A298 );
 a33006a <=( A301  and  A300 );
 a33007a <=( a33006a  and  a33003a );
 a33008a <=( a33007a  and  a33000a );
 a33012a <=( A167  and  A168 );
 a33013a <=( A169  and  a33012a );
 a33016a <=( (not A199)  and  (not A166) );
 a33019a <=( (not A232)  and  (not A200) );
 a33020a <=( a33019a  and  a33016a );
 a33021a <=( a33020a  and  a33013a );
 a33024a <=( (not A234)  and  A233 );
 a33027a <=( (not A236)  and  (not A235) );
 a33028a <=( a33027a  and  a33024a );
 a33031a <=( (not A299)  and  A298 );
 a33034a <=( A302  and  A300 );
 a33035a <=( a33034a  and  a33031a );
 a33036a <=( a33035a  and  a33028a );
 a33040a <=( A167  and  A168 );
 a33041a <=( A169  and  a33040a );
 a33044a <=( (not A199)  and  (not A166) );
 a33047a <=( (not A232)  and  (not A200) );
 a33048a <=( a33047a  and  a33044a );
 a33049a <=( a33048a  and  a33041a );
 a33052a <=( (not A234)  and  A233 );
 a33055a <=( (not A236)  and  (not A235) );
 a33056a <=( a33055a  and  a33052a );
 a33059a <=( A299  and  (not A298) );
 a33062a <=( A301  and  A300 );
 a33063a <=( a33062a  and  a33059a );
 a33064a <=( a33063a  and  a33056a );
 a33068a <=( A167  and  A168 );
 a33069a <=( A169  and  a33068a );
 a33072a <=( (not A199)  and  (not A166) );
 a33075a <=( (not A232)  and  (not A200) );
 a33076a <=( a33075a  and  a33072a );
 a33077a <=( a33076a  and  a33069a );
 a33080a <=( (not A234)  and  A233 );
 a33083a <=( (not A236)  and  (not A235) );
 a33084a <=( a33083a  and  a33080a );
 a33087a <=( A299  and  (not A298) );
 a33090a <=( A302  and  A300 );
 a33091a <=( a33090a  and  a33087a );
 a33092a <=( a33091a  and  a33084a );
 a33096a <=( A167  and  A168 );
 a33097a <=( A169  and  a33096a );
 a33100a <=( (not A199)  and  (not A166) );
 a33103a <=( (not A232)  and  (not A200) );
 a33104a <=( a33103a  and  a33100a );
 a33105a <=( a33104a  and  a33097a );
 a33108a <=( (not A234)  and  A233 );
 a33111a <=( (not A236)  and  (not A235) );
 a33112a <=( a33111a  and  a33108a );
 a33115a <=( A266  and  (not A265) );
 a33118a <=( A268  and  A267 );
 a33119a <=( a33118a  and  a33115a );
 a33120a <=( a33119a  and  a33112a );
 a33124a <=( A167  and  A168 );
 a33125a <=( A169  and  a33124a );
 a33128a <=( (not A199)  and  (not A166) );
 a33131a <=( (not A232)  and  (not A200) );
 a33132a <=( a33131a  and  a33128a );
 a33133a <=( a33132a  and  a33125a );
 a33136a <=( (not A234)  and  A233 );
 a33139a <=( (not A236)  and  (not A235) );
 a33140a <=( a33139a  and  a33136a );
 a33143a <=( A266  and  (not A265) );
 a33146a <=( A269  and  A267 );
 a33147a <=( a33146a  and  a33143a );
 a33148a <=( a33147a  and  a33140a );
 a33152a <=( A167  and  A168 );
 a33153a <=( A169  and  a33152a );
 a33156a <=( (not A199)  and  (not A166) );
 a33159a <=( (not A232)  and  (not A200) );
 a33160a <=( a33159a  and  a33156a );
 a33161a <=( a33160a  and  a33153a );
 a33164a <=( (not A234)  and  A233 );
 a33167a <=( (not A236)  and  (not A235) );
 a33168a <=( a33167a  and  a33164a );
 a33171a <=( (not A266)  and  A265 );
 a33174a <=( A268  and  A267 );
 a33175a <=( a33174a  and  a33171a );
 a33176a <=( a33175a  and  a33168a );
 a33180a <=( A167  and  A168 );
 a33181a <=( A169  and  a33180a );
 a33184a <=( (not A199)  and  (not A166) );
 a33187a <=( (not A232)  and  (not A200) );
 a33188a <=( a33187a  and  a33184a );
 a33189a <=( a33188a  and  a33181a );
 a33192a <=( (not A234)  and  A233 );
 a33195a <=( (not A236)  and  (not A235) );
 a33196a <=( a33195a  and  a33192a );
 a33199a <=( (not A266)  and  A265 );
 a33202a <=( A269  and  A267 );
 a33203a <=( a33202a  and  a33199a );
 a33204a <=( a33203a  and  a33196a );
 a33208a <=( A167  and  A168 );
 a33209a <=( A169  and  a33208a );
 a33212a <=( (not A199)  and  (not A166) );
 a33215a <=( A232  and  (not A200) );
 a33216a <=( a33215a  and  a33212a );
 a33217a <=( a33216a  and  a33209a );
 a33220a <=( A234  and  (not A233) );
 a33223a <=( A298  and  A235 );
 a33224a <=( a33223a  and  a33220a );
 a33227a <=( (not A300)  and  (not A299) );
 a33230a <=( (not A302)  and  (not A301) );
 a33231a <=( a33230a  and  a33227a );
 a33232a <=( a33231a  and  a33224a );
 a33236a <=( A167  and  A168 );
 a33237a <=( A169  and  a33236a );
 a33240a <=( (not A199)  and  (not A166) );
 a33243a <=( A232  and  (not A200) );
 a33244a <=( a33243a  and  a33240a );
 a33245a <=( a33244a  and  a33237a );
 a33248a <=( A234  and  (not A233) );
 a33251a <=( (not A298)  and  A235 );
 a33252a <=( a33251a  and  a33248a );
 a33255a <=( (not A300)  and  A299 );
 a33258a <=( (not A302)  and  (not A301) );
 a33259a <=( a33258a  and  a33255a );
 a33260a <=( a33259a  and  a33252a );
 a33264a <=( A167  and  A168 );
 a33265a <=( A169  and  a33264a );
 a33268a <=( (not A199)  and  (not A166) );
 a33271a <=( A232  and  (not A200) );
 a33272a <=( a33271a  and  a33268a );
 a33273a <=( a33272a  and  a33265a );
 a33276a <=( A234  and  (not A233) );
 a33279a <=( (not A265)  and  A235 );
 a33280a <=( a33279a  and  a33276a );
 a33283a <=( (not A267)  and  A266 );
 a33286a <=( (not A269)  and  (not A268) );
 a33287a <=( a33286a  and  a33283a );
 a33288a <=( a33287a  and  a33280a );
 a33292a <=( A167  and  A168 );
 a33293a <=( A169  and  a33292a );
 a33296a <=( (not A199)  and  (not A166) );
 a33299a <=( A232  and  (not A200) );
 a33300a <=( a33299a  and  a33296a );
 a33301a <=( a33300a  and  a33293a );
 a33304a <=( A234  and  (not A233) );
 a33307a <=( A265  and  A235 );
 a33308a <=( a33307a  and  a33304a );
 a33311a <=( (not A267)  and  (not A266) );
 a33314a <=( (not A269)  and  (not A268) );
 a33315a <=( a33314a  and  a33311a );
 a33316a <=( a33315a  and  a33308a );
 a33320a <=( A167  and  A168 );
 a33321a <=( A169  and  a33320a );
 a33324a <=( (not A199)  and  (not A166) );
 a33327a <=( A232  and  (not A200) );
 a33328a <=( a33327a  and  a33324a );
 a33329a <=( a33328a  and  a33321a );
 a33332a <=( A234  and  (not A233) );
 a33335a <=( A298  and  A236 );
 a33336a <=( a33335a  and  a33332a );
 a33339a <=( (not A300)  and  (not A299) );
 a33342a <=( (not A302)  and  (not A301) );
 a33343a <=( a33342a  and  a33339a );
 a33344a <=( a33343a  and  a33336a );
 a33348a <=( A167  and  A168 );
 a33349a <=( A169  and  a33348a );
 a33352a <=( (not A199)  and  (not A166) );
 a33355a <=( A232  and  (not A200) );
 a33356a <=( a33355a  and  a33352a );
 a33357a <=( a33356a  and  a33349a );
 a33360a <=( A234  and  (not A233) );
 a33363a <=( (not A298)  and  A236 );
 a33364a <=( a33363a  and  a33360a );
 a33367a <=( (not A300)  and  A299 );
 a33370a <=( (not A302)  and  (not A301) );
 a33371a <=( a33370a  and  a33367a );
 a33372a <=( a33371a  and  a33364a );
 a33376a <=( A167  and  A168 );
 a33377a <=( A169  and  a33376a );
 a33380a <=( (not A199)  and  (not A166) );
 a33383a <=( A232  and  (not A200) );
 a33384a <=( a33383a  and  a33380a );
 a33385a <=( a33384a  and  a33377a );
 a33388a <=( A234  and  (not A233) );
 a33391a <=( (not A265)  and  A236 );
 a33392a <=( a33391a  and  a33388a );
 a33395a <=( (not A267)  and  A266 );
 a33398a <=( (not A269)  and  (not A268) );
 a33399a <=( a33398a  and  a33395a );
 a33400a <=( a33399a  and  a33392a );
 a33404a <=( A167  and  A168 );
 a33405a <=( A169  and  a33404a );
 a33408a <=( (not A199)  and  (not A166) );
 a33411a <=( A232  and  (not A200) );
 a33412a <=( a33411a  and  a33408a );
 a33413a <=( a33412a  and  a33405a );
 a33416a <=( A234  and  (not A233) );
 a33419a <=( A265  and  A236 );
 a33420a <=( a33419a  and  a33416a );
 a33423a <=( (not A267)  and  (not A266) );
 a33426a <=( (not A269)  and  (not A268) );
 a33427a <=( a33426a  and  a33423a );
 a33428a <=( a33427a  and  a33420a );
 a33432a <=( A167  and  A168 );
 a33433a <=( A169  and  a33432a );
 a33436a <=( (not A199)  and  (not A166) );
 a33439a <=( A232  and  (not A200) );
 a33440a <=( a33439a  and  a33436a );
 a33441a <=( a33440a  and  a33433a );
 a33444a <=( (not A234)  and  (not A233) );
 a33447a <=( (not A236)  and  (not A235) );
 a33448a <=( a33447a  and  a33444a );
 a33451a <=( (not A299)  and  A298 );
 a33454a <=( A301  and  A300 );
 a33455a <=( a33454a  and  a33451a );
 a33456a <=( a33455a  and  a33448a );
 a33460a <=( A167  and  A168 );
 a33461a <=( A169  and  a33460a );
 a33464a <=( (not A199)  and  (not A166) );
 a33467a <=( A232  and  (not A200) );
 a33468a <=( a33467a  and  a33464a );
 a33469a <=( a33468a  and  a33461a );
 a33472a <=( (not A234)  and  (not A233) );
 a33475a <=( (not A236)  and  (not A235) );
 a33476a <=( a33475a  and  a33472a );
 a33479a <=( (not A299)  and  A298 );
 a33482a <=( A302  and  A300 );
 a33483a <=( a33482a  and  a33479a );
 a33484a <=( a33483a  and  a33476a );
 a33488a <=( A167  and  A168 );
 a33489a <=( A169  and  a33488a );
 a33492a <=( (not A199)  and  (not A166) );
 a33495a <=( A232  and  (not A200) );
 a33496a <=( a33495a  and  a33492a );
 a33497a <=( a33496a  and  a33489a );
 a33500a <=( (not A234)  and  (not A233) );
 a33503a <=( (not A236)  and  (not A235) );
 a33504a <=( a33503a  and  a33500a );
 a33507a <=( A299  and  (not A298) );
 a33510a <=( A301  and  A300 );
 a33511a <=( a33510a  and  a33507a );
 a33512a <=( a33511a  and  a33504a );
 a33516a <=( A167  and  A168 );
 a33517a <=( A169  and  a33516a );
 a33520a <=( (not A199)  and  (not A166) );
 a33523a <=( A232  and  (not A200) );
 a33524a <=( a33523a  and  a33520a );
 a33525a <=( a33524a  and  a33517a );
 a33528a <=( (not A234)  and  (not A233) );
 a33531a <=( (not A236)  and  (not A235) );
 a33532a <=( a33531a  and  a33528a );
 a33535a <=( A299  and  (not A298) );
 a33538a <=( A302  and  A300 );
 a33539a <=( a33538a  and  a33535a );
 a33540a <=( a33539a  and  a33532a );
 a33544a <=( A167  and  A168 );
 a33545a <=( A169  and  a33544a );
 a33548a <=( (not A199)  and  (not A166) );
 a33551a <=( A232  and  (not A200) );
 a33552a <=( a33551a  and  a33548a );
 a33553a <=( a33552a  and  a33545a );
 a33556a <=( (not A234)  and  (not A233) );
 a33559a <=( (not A236)  and  (not A235) );
 a33560a <=( a33559a  and  a33556a );
 a33563a <=( A266  and  (not A265) );
 a33566a <=( A268  and  A267 );
 a33567a <=( a33566a  and  a33563a );
 a33568a <=( a33567a  and  a33560a );
 a33572a <=( A167  and  A168 );
 a33573a <=( A169  and  a33572a );
 a33576a <=( (not A199)  and  (not A166) );
 a33579a <=( A232  and  (not A200) );
 a33580a <=( a33579a  and  a33576a );
 a33581a <=( a33580a  and  a33573a );
 a33584a <=( (not A234)  and  (not A233) );
 a33587a <=( (not A236)  and  (not A235) );
 a33588a <=( a33587a  and  a33584a );
 a33591a <=( A266  and  (not A265) );
 a33594a <=( A269  and  A267 );
 a33595a <=( a33594a  and  a33591a );
 a33596a <=( a33595a  and  a33588a );
 a33600a <=( A167  and  A168 );
 a33601a <=( A169  and  a33600a );
 a33604a <=( (not A199)  and  (not A166) );
 a33607a <=( A232  and  (not A200) );
 a33608a <=( a33607a  and  a33604a );
 a33609a <=( a33608a  and  a33601a );
 a33612a <=( (not A234)  and  (not A233) );
 a33615a <=( (not A236)  and  (not A235) );
 a33616a <=( a33615a  and  a33612a );
 a33619a <=( (not A266)  and  A265 );
 a33622a <=( A268  and  A267 );
 a33623a <=( a33622a  and  a33619a );
 a33624a <=( a33623a  and  a33616a );
 a33628a <=( A167  and  A168 );
 a33629a <=( A169  and  a33628a );
 a33632a <=( (not A199)  and  (not A166) );
 a33635a <=( A232  and  (not A200) );
 a33636a <=( a33635a  and  a33632a );
 a33637a <=( a33636a  and  a33629a );
 a33640a <=( (not A234)  and  (not A233) );
 a33643a <=( (not A236)  and  (not A235) );
 a33644a <=( a33643a  and  a33640a );
 a33647a <=( (not A266)  and  A265 );
 a33650a <=( A269  and  A267 );
 a33651a <=( a33650a  and  a33647a );
 a33652a <=( a33651a  and  a33644a );
 a33656a <=( (not A167)  and  A168 );
 a33657a <=( A169  and  a33656a );
 a33660a <=( A201  and  A166 );
 a33663a <=( (not A203)  and  (not A202) );
 a33664a <=( a33663a  and  a33660a );
 a33665a <=( a33664a  and  a33657a );
 a33668a <=( A233  and  (not A232) );
 a33671a <=( A235  and  A234 );
 a33672a <=( a33671a  and  a33668a );
 a33675a <=( (not A299)  and  A298 );
 a33678a <=( A301  and  A300 );
 a33679a <=( a33678a  and  a33675a );
 a33680a <=( a33679a  and  a33672a );
 a33684a <=( (not A167)  and  A168 );
 a33685a <=( A169  and  a33684a );
 a33688a <=( A201  and  A166 );
 a33691a <=( (not A203)  and  (not A202) );
 a33692a <=( a33691a  and  a33688a );
 a33693a <=( a33692a  and  a33685a );
 a33696a <=( A233  and  (not A232) );
 a33699a <=( A235  and  A234 );
 a33700a <=( a33699a  and  a33696a );
 a33703a <=( (not A299)  and  A298 );
 a33706a <=( A302  and  A300 );
 a33707a <=( a33706a  and  a33703a );
 a33708a <=( a33707a  and  a33700a );
 a33712a <=( (not A167)  and  A168 );
 a33713a <=( A169  and  a33712a );
 a33716a <=( A201  and  A166 );
 a33719a <=( (not A203)  and  (not A202) );
 a33720a <=( a33719a  and  a33716a );
 a33721a <=( a33720a  and  a33713a );
 a33724a <=( A233  and  (not A232) );
 a33727a <=( A235  and  A234 );
 a33728a <=( a33727a  and  a33724a );
 a33731a <=( A299  and  (not A298) );
 a33734a <=( A301  and  A300 );
 a33735a <=( a33734a  and  a33731a );
 a33736a <=( a33735a  and  a33728a );
 a33740a <=( (not A167)  and  A168 );
 a33741a <=( A169  and  a33740a );
 a33744a <=( A201  and  A166 );
 a33747a <=( (not A203)  and  (not A202) );
 a33748a <=( a33747a  and  a33744a );
 a33749a <=( a33748a  and  a33741a );
 a33752a <=( A233  and  (not A232) );
 a33755a <=( A235  and  A234 );
 a33756a <=( a33755a  and  a33752a );
 a33759a <=( A299  and  (not A298) );
 a33762a <=( A302  and  A300 );
 a33763a <=( a33762a  and  a33759a );
 a33764a <=( a33763a  and  a33756a );
 a33768a <=( (not A167)  and  A168 );
 a33769a <=( A169  and  a33768a );
 a33772a <=( A201  and  A166 );
 a33775a <=( (not A203)  and  (not A202) );
 a33776a <=( a33775a  and  a33772a );
 a33777a <=( a33776a  and  a33769a );
 a33780a <=( A233  and  (not A232) );
 a33783a <=( A235  and  A234 );
 a33784a <=( a33783a  and  a33780a );
 a33787a <=( A266  and  (not A265) );
 a33790a <=( A268  and  A267 );
 a33791a <=( a33790a  and  a33787a );
 a33792a <=( a33791a  and  a33784a );
 a33796a <=( (not A167)  and  A168 );
 a33797a <=( A169  and  a33796a );
 a33800a <=( A201  and  A166 );
 a33803a <=( (not A203)  and  (not A202) );
 a33804a <=( a33803a  and  a33800a );
 a33805a <=( a33804a  and  a33797a );
 a33808a <=( A233  and  (not A232) );
 a33811a <=( A235  and  A234 );
 a33812a <=( a33811a  and  a33808a );
 a33815a <=( A266  and  (not A265) );
 a33818a <=( A269  and  A267 );
 a33819a <=( a33818a  and  a33815a );
 a33820a <=( a33819a  and  a33812a );
 a33824a <=( (not A167)  and  A168 );
 a33825a <=( A169  and  a33824a );
 a33828a <=( A201  and  A166 );
 a33831a <=( (not A203)  and  (not A202) );
 a33832a <=( a33831a  and  a33828a );
 a33833a <=( a33832a  and  a33825a );
 a33836a <=( A233  and  (not A232) );
 a33839a <=( A235  and  A234 );
 a33840a <=( a33839a  and  a33836a );
 a33843a <=( (not A266)  and  A265 );
 a33846a <=( A268  and  A267 );
 a33847a <=( a33846a  and  a33843a );
 a33848a <=( a33847a  and  a33840a );
 a33852a <=( (not A167)  and  A168 );
 a33853a <=( A169  and  a33852a );
 a33856a <=( A201  and  A166 );
 a33859a <=( (not A203)  and  (not A202) );
 a33860a <=( a33859a  and  a33856a );
 a33861a <=( a33860a  and  a33853a );
 a33864a <=( A233  and  (not A232) );
 a33867a <=( A235  and  A234 );
 a33868a <=( a33867a  and  a33864a );
 a33871a <=( (not A266)  and  A265 );
 a33874a <=( A269  and  A267 );
 a33875a <=( a33874a  and  a33871a );
 a33876a <=( a33875a  and  a33868a );
 a33880a <=( (not A167)  and  A168 );
 a33881a <=( A169  and  a33880a );
 a33884a <=( A201  and  A166 );
 a33887a <=( (not A203)  and  (not A202) );
 a33888a <=( a33887a  and  a33884a );
 a33889a <=( a33888a  and  a33881a );
 a33892a <=( A233  and  (not A232) );
 a33895a <=( A236  and  A234 );
 a33896a <=( a33895a  and  a33892a );
 a33899a <=( (not A299)  and  A298 );
 a33902a <=( A301  and  A300 );
 a33903a <=( a33902a  and  a33899a );
 a33904a <=( a33903a  and  a33896a );
 a33908a <=( (not A167)  and  A168 );
 a33909a <=( A169  and  a33908a );
 a33912a <=( A201  and  A166 );
 a33915a <=( (not A203)  and  (not A202) );
 a33916a <=( a33915a  and  a33912a );
 a33917a <=( a33916a  and  a33909a );
 a33920a <=( A233  and  (not A232) );
 a33923a <=( A236  and  A234 );
 a33924a <=( a33923a  and  a33920a );
 a33927a <=( (not A299)  and  A298 );
 a33930a <=( A302  and  A300 );
 a33931a <=( a33930a  and  a33927a );
 a33932a <=( a33931a  and  a33924a );
 a33936a <=( (not A167)  and  A168 );
 a33937a <=( A169  and  a33936a );
 a33940a <=( A201  and  A166 );
 a33943a <=( (not A203)  and  (not A202) );
 a33944a <=( a33943a  and  a33940a );
 a33945a <=( a33944a  and  a33937a );
 a33948a <=( A233  and  (not A232) );
 a33951a <=( A236  and  A234 );
 a33952a <=( a33951a  and  a33948a );
 a33955a <=( A299  and  (not A298) );
 a33958a <=( A301  and  A300 );
 a33959a <=( a33958a  and  a33955a );
 a33960a <=( a33959a  and  a33952a );
 a33964a <=( (not A167)  and  A168 );
 a33965a <=( A169  and  a33964a );
 a33968a <=( A201  and  A166 );
 a33971a <=( (not A203)  and  (not A202) );
 a33972a <=( a33971a  and  a33968a );
 a33973a <=( a33972a  and  a33965a );
 a33976a <=( A233  and  (not A232) );
 a33979a <=( A236  and  A234 );
 a33980a <=( a33979a  and  a33976a );
 a33983a <=( A299  and  (not A298) );
 a33986a <=( A302  and  A300 );
 a33987a <=( a33986a  and  a33983a );
 a33988a <=( a33987a  and  a33980a );
 a33992a <=( (not A167)  and  A168 );
 a33993a <=( A169  and  a33992a );
 a33996a <=( A201  and  A166 );
 a33999a <=( (not A203)  and  (not A202) );
 a34000a <=( a33999a  and  a33996a );
 a34001a <=( a34000a  and  a33993a );
 a34004a <=( A233  and  (not A232) );
 a34007a <=( A236  and  A234 );
 a34008a <=( a34007a  and  a34004a );
 a34011a <=( A266  and  (not A265) );
 a34014a <=( A268  and  A267 );
 a34015a <=( a34014a  and  a34011a );
 a34016a <=( a34015a  and  a34008a );
 a34020a <=( (not A167)  and  A168 );
 a34021a <=( A169  and  a34020a );
 a34024a <=( A201  and  A166 );
 a34027a <=( (not A203)  and  (not A202) );
 a34028a <=( a34027a  and  a34024a );
 a34029a <=( a34028a  and  a34021a );
 a34032a <=( A233  and  (not A232) );
 a34035a <=( A236  and  A234 );
 a34036a <=( a34035a  and  a34032a );
 a34039a <=( A266  and  (not A265) );
 a34042a <=( A269  and  A267 );
 a34043a <=( a34042a  and  a34039a );
 a34044a <=( a34043a  and  a34036a );
 a34048a <=( (not A167)  and  A168 );
 a34049a <=( A169  and  a34048a );
 a34052a <=( A201  and  A166 );
 a34055a <=( (not A203)  and  (not A202) );
 a34056a <=( a34055a  and  a34052a );
 a34057a <=( a34056a  and  a34049a );
 a34060a <=( A233  and  (not A232) );
 a34063a <=( A236  and  A234 );
 a34064a <=( a34063a  and  a34060a );
 a34067a <=( (not A266)  and  A265 );
 a34070a <=( A268  and  A267 );
 a34071a <=( a34070a  and  a34067a );
 a34072a <=( a34071a  and  a34064a );
 a34076a <=( (not A167)  and  A168 );
 a34077a <=( A169  and  a34076a );
 a34080a <=( A201  and  A166 );
 a34083a <=( (not A203)  and  (not A202) );
 a34084a <=( a34083a  and  a34080a );
 a34085a <=( a34084a  and  a34077a );
 a34088a <=( A233  and  (not A232) );
 a34091a <=( A236  and  A234 );
 a34092a <=( a34091a  and  a34088a );
 a34095a <=( (not A266)  and  A265 );
 a34098a <=( A269  and  A267 );
 a34099a <=( a34098a  and  a34095a );
 a34100a <=( a34099a  and  a34092a );
 a34104a <=( (not A167)  and  A168 );
 a34105a <=( A169  and  a34104a );
 a34108a <=( A201  and  A166 );
 a34111a <=( (not A203)  and  (not A202) );
 a34112a <=( a34111a  and  a34108a );
 a34113a <=( a34112a  and  a34105a );
 a34116a <=( (not A233)  and  A232 );
 a34119a <=( A235  and  A234 );
 a34120a <=( a34119a  and  a34116a );
 a34123a <=( (not A299)  and  A298 );
 a34126a <=( A301  and  A300 );
 a34127a <=( a34126a  and  a34123a );
 a34128a <=( a34127a  and  a34120a );
 a34132a <=( (not A167)  and  A168 );
 a34133a <=( A169  and  a34132a );
 a34136a <=( A201  and  A166 );
 a34139a <=( (not A203)  and  (not A202) );
 a34140a <=( a34139a  and  a34136a );
 a34141a <=( a34140a  and  a34133a );
 a34144a <=( (not A233)  and  A232 );
 a34147a <=( A235  and  A234 );
 a34148a <=( a34147a  and  a34144a );
 a34151a <=( (not A299)  and  A298 );
 a34154a <=( A302  and  A300 );
 a34155a <=( a34154a  and  a34151a );
 a34156a <=( a34155a  and  a34148a );
 a34160a <=( (not A167)  and  A168 );
 a34161a <=( A169  and  a34160a );
 a34164a <=( A201  and  A166 );
 a34167a <=( (not A203)  and  (not A202) );
 a34168a <=( a34167a  and  a34164a );
 a34169a <=( a34168a  and  a34161a );
 a34172a <=( (not A233)  and  A232 );
 a34175a <=( A235  and  A234 );
 a34176a <=( a34175a  and  a34172a );
 a34179a <=( A299  and  (not A298) );
 a34182a <=( A301  and  A300 );
 a34183a <=( a34182a  and  a34179a );
 a34184a <=( a34183a  and  a34176a );
 a34188a <=( (not A167)  and  A168 );
 a34189a <=( A169  and  a34188a );
 a34192a <=( A201  and  A166 );
 a34195a <=( (not A203)  and  (not A202) );
 a34196a <=( a34195a  and  a34192a );
 a34197a <=( a34196a  and  a34189a );
 a34200a <=( (not A233)  and  A232 );
 a34203a <=( A235  and  A234 );
 a34204a <=( a34203a  and  a34200a );
 a34207a <=( A299  and  (not A298) );
 a34210a <=( A302  and  A300 );
 a34211a <=( a34210a  and  a34207a );
 a34212a <=( a34211a  and  a34204a );
 a34216a <=( (not A167)  and  A168 );
 a34217a <=( A169  and  a34216a );
 a34220a <=( A201  and  A166 );
 a34223a <=( (not A203)  and  (not A202) );
 a34224a <=( a34223a  and  a34220a );
 a34225a <=( a34224a  and  a34217a );
 a34228a <=( (not A233)  and  A232 );
 a34231a <=( A235  and  A234 );
 a34232a <=( a34231a  and  a34228a );
 a34235a <=( A266  and  (not A265) );
 a34238a <=( A268  and  A267 );
 a34239a <=( a34238a  and  a34235a );
 a34240a <=( a34239a  and  a34232a );
 a34244a <=( (not A167)  and  A168 );
 a34245a <=( A169  and  a34244a );
 a34248a <=( A201  and  A166 );
 a34251a <=( (not A203)  and  (not A202) );
 a34252a <=( a34251a  and  a34248a );
 a34253a <=( a34252a  and  a34245a );
 a34256a <=( (not A233)  and  A232 );
 a34259a <=( A235  and  A234 );
 a34260a <=( a34259a  and  a34256a );
 a34263a <=( A266  and  (not A265) );
 a34266a <=( A269  and  A267 );
 a34267a <=( a34266a  and  a34263a );
 a34268a <=( a34267a  and  a34260a );
 a34272a <=( (not A167)  and  A168 );
 a34273a <=( A169  and  a34272a );
 a34276a <=( A201  and  A166 );
 a34279a <=( (not A203)  and  (not A202) );
 a34280a <=( a34279a  and  a34276a );
 a34281a <=( a34280a  and  a34273a );
 a34284a <=( (not A233)  and  A232 );
 a34287a <=( A235  and  A234 );
 a34288a <=( a34287a  and  a34284a );
 a34291a <=( (not A266)  and  A265 );
 a34294a <=( A268  and  A267 );
 a34295a <=( a34294a  and  a34291a );
 a34296a <=( a34295a  and  a34288a );
 a34300a <=( (not A167)  and  A168 );
 a34301a <=( A169  and  a34300a );
 a34304a <=( A201  and  A166 );
 a34307a <=( (not A203)  and  (not A202) );
 a34308a <=( a34307a  and  a34304a );
 a34309a <=( a34308a  and  a34301a );
 a34312a <=( (not A233)  and  A232 );
 a34315a <=( A235  and  A234 );
 a34316a <=( a34315a  and  a34312a );
 a34319a <=( (not A266)  and  A265 );
 a34322a <=( A269  and  A267 );
 a34323a <=( a34322a  and  a34319a );
 a34324a <=( a34323a  and  a34316a );
 a34328a <=( (not A167)  and  A168 );
 a34329a <=( A169  and  a34328a );
 a34332a <=( A201  and  A166 );
 a34335a <=( (not A203)  and  (not A202) );
 a34336a <=( a34335a  and  a34332a );
 a34337a <=( a34336a  and  a34329a );
 a34340a <=( (not A233)  and  A232 );
 a34343a <=( A236  and  A234 );
 a34344a <=( a34343a  and  a34340a );
 a34347a <=( (not A299)  and  A298 );
 a34350a <=( A301  and  A300 );
 a34351a <=( a34350a  and  a34347a );
 a34352a <=( a34351a  and  a34344a );
 a34356a <=( (not A167)  and  A168 );
 a34357a <=( A169  and  a34356a );
 a34360a <=( A201  and  A166 );
 a34363a <=( (not A203)  and  (not A202) );
 a34364a <=( a34363a  and  a34360a );
 a34365a <=( a34364a  and  a34357a );
 a34368a <=( (not A233)  and  A232 );
 a34371a <=( A236  and  A234 );
 a34372a <=( a34371a  and  a34368a );
 a34375a <=( (not A299)  and  A298 );
 a34378a <=( A302  and  A300 );
 a34379a <=( a34378a  and  a34375a );
 a34380a <=( a34379a  and  a34372a );
 a34384a <=( (not A167)  and  A168 );
 a34385a <=( A169  and  a34384a );
 a34388a <=( A201  and  A166 );
 a34391a <=( (not A203)  and  (not A202) );
 a34392a <=( a34391a  and  a34388a );
 a34393a <=( a34392a  and  a34385a );
 a34396a <=( (not A233)  and  A232 );
 a34399a <=( A236  and  A234 );
 a34400a <=( a34399a  and  a34396a );
 a34403a <=( A299  and  (not A298) );
 a34406a <=( A301  and  A300 );
 a34407a <=( a34406a  and  a34403a );
 a34408a <=( a34407a  and  a34400a );
 a34412a <=( (not A167)  and  A168 );
 a34413a <=( A169  and  a34412a );
 a34416a <=( A201  and  A166 );
 a34419a <=( (not A203)  and  (not A202) );
 a34420a <=( a34419a  and  a34416a );
 a34421a <=( a34420a  and  a34413a );
 a34424a <=( (not A233)  and  A232 );
 a34427a <=( A236  and  A234 );
 a34428a <=( a34427a  and  a34424a );
 a34431a <=( A299  and  (not A298) );
 a34434a <=( A302  and  A300 );
 a34435a <=( a34434a  and  a34431a );
 a34436a <=( a34435a  and  a34428a );
 a34440a <=( (not A167)  and  A168 );
 a34441a <=( A169  and  a34440a );
 a34444a <=( A201  and  A166 );
 a34447a <=( (not A203)  and  (not A202) );
 a34448a <=( a34447a  and  a34444a );
 a34449a <=( a34448a  and  a34441a );
 a34452a <=( (not A233)  and  A232 );
 a34455a <=( A236  and  A234 );
 a34456a <=( a34455a  and  a34452a );
 a34459a <=( A266  and  (not A265) );
 a34462a <=( A268  and  A267 );
 a34463a <=( a34462a  and  a34459a );
 a34464a <=( a34463a  and  a34456a );
 a34468a <=( (not A167)  and  A168 );
 a34469a <=( A169  and  a34468a );
 a34472a <=( A201  and  A166 );
 a34475a <=( (not A203)  and  (not A202) );
 a34476a <=( a34475a  and  a34472a );
 a34477a <=( a34476a  and  a34469a );
 a34480a <=( (not A233)  and  A232 );
 a34483a <=( A236  and  A234 );
 a34484a <=( a34483a  and  a34480a );
 a34487a <=( A266  and  (not A265) );
 a34490a <=( A269  and  A267 );
 a34491a <=( a34490a  and  a34487a );
 a34492a <=( a34491a  and  a34484a );
 a34496a <=( (not A167)  and  A168 );
 a34497a <=( A169  and  a34496a );
 a34500a <=( A201  and  A166 );
 a34503a <=( (not A203)  and  (not A202) );
 a34504a <=( a34503a  and  a34500a );
 a34505a <=( a34504a  and  a34497a );
 a34508a <=( (not A233)  and  A232 );
 a34511a <=( A236  and  A234 );
 a34512a <=( a34511a  and  a34508a );
 a34515a <=( (not A266)  and  A265 );
 a34518a <=( A268  and  A267 );
 a34519a <=( a34518a  and  a34515a );
 a34520a <=( a34519a  and  a34512a );
 a34524a <=( (not A167)  and  A168 );
 a34525a <=( A169  and  a34524a );
 a34528a <=( A201  and  A166 );
 a34531a <=( (not A203)  and  (not A202) );
 a34532a <=( a34531a  and  a34528a );
 a34533a <=( a34532a  and  a34525a );
 a34536a <=( (not A233)  and  A232 );
 a34539a <=( A236  and  A234 );
 a34540a <=( a34539a  and  a34536a );
 a34543a <=( (not A266)  and  A265 );
 a34546a <=( A269  and  A267 );
 a34547a <=( a34546a  and  a34543a );
 a34548a <=( a34547a  and  a34540a );
 a34552a <=( (not A167)  and  A168 );
 a34553a <=( A169  and  a34552a );
 a34556a <=( (not A201)  and  A166 );
 a34559a <=( (not A232)  and  A202 );
 a34560a <=( a34559a  and  a34556a );
 a34561a <=( a34560a  and  a34553a );
 a34564a <=( A234  and  A233 );
 a34567a <=( A298  and  A235 );
 a34568a <=( a34567a  and  a34564a );
 a34571a <=( (not A300)  and  (not A299) );
 a34574a <=( (not A302)  and  (not A301) );
 a34575a <=( a34574a  and  a34571a );
 a34576a <=( a34575a  and  a34568a );
 a34580a <=( (not A167)  and  A168 );
 a34581a <=( A169  and  a34580a );
 a34584a <=( (not A201)  and  A166 );
 a34587a <=( (not A232)  and  A202 );
 a34588a <=( a34587a  and  a34584a );
 a34589a <=( a34588a  and  a34581a );
 a34592a <=( A234  and  A233 );
 a34595a <=( (not A298)  and  A235 );
 a34596a <=( a34595a  and  a34592a );
 a34599a <=( (not A300)  and  A299 );
 a34602a <=( (not A302)  and  (not A301) );
 a34603a <=( a34602a  and  a34599a );
 a34604a <=( a34603a  and  a34596a );
 a34608a <=( (not A167)  and  A168 );
 a34609a <=( A169  and  a34608a );
 a34612a <=( (not A201)  and  A166 );
 a34615a <=( (not A232)  and  A202 );
 a34616a <=( a34615a  and  a34612a );
 a34617a <=( a34616a  and  a34609a );
 a34620a <=( A234  and  A233 );
 a34623a <=( (not A265)  and  A235 );
 a34624a <=( a34623a  and  a34620a );
 a34627a <=( (not A267)  and  A266 );
 a34630a <=( (not A269)  and  (not A268) );
 a34631a <=( a34630a  and  a34627a );
 a34632a <=( a34631a  and  a34624a );
 a34636a <=( (not A167)  and  A168 );
 a34637a <=( A169  and  a34636a );
 a34640a <=( (not A201)  and  A166 );
 a34643a <=( (not A232)  and  A202 );
 a34644a <=( a34643a  and  a34640a );
 a34645a <=( a34644a  and  a34637a );
 a34648a <=( A234  and  A233 );
 a34651a <=( A265  and  A235 );
 a34652a <=( a34651a  and  a34648a );
 a34655a <=( (not A267)  and  (not A266) );
 a34658a <=( (not A269)  and  (not A268) );
 a34659a <=( a34658a  and  a34655a );
 a34660a <=( a34659a  and  a34652a );
 a34664a <=( (not A167)  and  A168 );
 a34665a <=( A169  and  a34664a );
 a34668a <=( (not A201)  and  A166 );
 a34671a <=( (not A232)  and  A202 );
 a34672a <=( a34671a  and  a34668a );
 a34673a <=( a34672a  and  a34665a );
 a34676a <=( A234  and  A233 );
 a34679a <=( A298  and  A236 );
 a34680a <=( a34679a  and  a34676a );
 a34683a <=( (not A300)  and  (not A299) );
 a34686a <=( (not A302)  and  (not A301) );
 a34687a <=( a34686a  and  a34683a );
 a34688a <=( a34687a  and  a34680a );
 a34692a <=( (not A167)  and  A168 );
 a34693a <=( A169  and  a34692a );
 a34696a <=( (not A201)  and  A166 );
 a34699a <=( (not A232)  and  A202 );
 a34700a <=( a34699a  and  a34696a );
 a34701a <=( a34700a  and  a34693a );
 a34704a <=( A234  and  A233 );
 a34707a <=( (not A298)  and  A236 );
 a34708a <=( a34707a  and  a34704a );
 a34711a <=( (not A300)  and  A299 );
 a34714a <=( (not A302)  and  (not A301) );
 a34715a <=( a34714a  and  a34711a );
 a34716a <=( a34715a  and  a34708a );
 a34720a <=( (not A167)  and  A168 );
 a34721a <=( A169  and  a34720a );
 a34724a <=( (not A201)  and  A166 );
 a34727a <=( (not A232)  and  A202 );
 a34728a <=( a34727a  and  a34724a );
 a34729a <=( a34728a  and  a34721a );
 a34732a <=( A234  and  A233 );
 a34735a <=( (not A265)  and  A236 );
 a34736a <=( a34735a  and  a34732a );
 a34739a <=( (not A267)  and  A266 );
 a34742a <=( (not A269)  and  (not A268) );
 a34743a <=( a34742a  and  a34739a );
 a34744a <=( a34743a  and  a34736a );
 a34748a <=( (not A167)  and  A168 );
 a34749a <=( A169  and  a34748a );
 a34752a <=( (not A201)  and  A166 );
 a34755a <=( (not A232)  and  A202 );
 a34756a <=( a34755a  and  a34752a );
 a34757a <=( a34756a  and  a34749a );
 a34760a <=( A234  and  A233 );
 a34763a <=( A265  and  A236 );
 a34764a <=( a34763a  and  a34760a );
 a34767a <=( (not A267)  and  (not A266) );
 a34770a <=( (not A269)  and  (not A268) );
 a34771a <=( a34770a  and  a34767a );
 a34772a <=( a34771a  and  a34764a );
 a34776a <=( (not A167)  and  A168 );
 a34777a <=( A169  and  a34776a );
 a34780a <=( (not A201)  and  A166 );
 a34783a <=( (not A232)  and  A202 );
 a34784a <=( a34783a  and  a34780a );
 a34785a <=( a34784a  and  a34777a );
 a34788a <=( (not A234)  and  A233 );
 a34791a <=( (not A236)  and  (not A235) );
 a34792a <=( a34791a  and  a34788a );
 a34795a <=( (not A299)  and  A298 );
 a34798a <=( A301  and  A300 );
 a34799a <=( a34798a  and  a34795a );
 a34800a <=( a34799a  and  a34792a );
 a34804a <=( (not A167)  and  A168 );
 a34805a <=( A169  and  a34804a );
 a34808a <=( (not A201)  and  A166 );
 a34811a <=( (not A232)  and  A202 );
 a34812a <=( a34811a  and  a34808a );
 a34813a <=( a34812a  and  a34805a );
 a34816a <=( (not A234)  and  A233 );
 a34819a <=( (not A236)  and  (not A235) );
 a34820a <=( a34819a  and  a34816a );
 a34823a <=( (not A299)  and  A298 );
 a34826a <=( A302  and  A300 );
 a34827a <=( a34826a  and  a34823a );
 a34828a <=( a34827a  and  a34820a );
 a34832a <=( (not A167)  and  A168 );
 a34833a <=( A169  and  a34832a );
 a34836a <=( (not A201)  and  A166 );
 a34839a <=( (not A232)  and  A202 );
 a34840a <=( a34839a  and  a34836a );
 a34841a <=( a34840a  and  a34833a );
 a34844a <=( (not A234)  and  A233 );
 a34847a <=( (not A236)  and  (not A235) );
 a34848a <=( a34847a  and  a34844a );
 a34851a <=( A299  and  (not A298) );
 a34854a <=( A301  and  A300 );
 a34855a <=( a34854a  and  a34851a );
 a34856a <=( a34855a  and  a34848a );
 a34860a <=( (not A167)  and  A168 );
 a34861a <=( A169  and  a34860a );
 a34864a <=( (not A201)  and  A166 );
 a34867a <=( (not A232)  and  A202 );
 a34868a <=( a34867a  and  a34864a );
 a34869a <=( a34868a  and  a34861a );
 a34872a <=( (not A234)  and  A233 );
 a34875a <=( (not A236)  and  (not A235) );
 a34876a <=( a34875a  and  a34872a );
 a34879a <=( A299  and  (not A298) );
 a34882a <=( A302  and  A300 );
 a34883a <=( a34882a  and  a34879a );
 a34884a <=( a34883a  and  a34876a );
 a34888a <=( (not A167)  and  A168 );
 a34889a <=( A169  and  a34888a );
 a34892a <=( (not A201)  and  A166 );
 a34895a <=( (not A232)  and  A202 );
 a34896a <=( a34895a  and  a34892a );
 a34897a <=( a34896a  and  a34889a );
 a34900a <=( (not A234)  and  A233 );
 a34903a <=( (not A236)  and  (not A235) );
 a34904a <=( a34903a  and  a34900a );
 a34907a <=( A266  and  (not A265) );
 a34910a <=( A268  and  A267 );
 a34911a <=( a34910a  and  a34907a );
 a34912a <=( a34911a  and  a34904a );
 a34916a <=( (not A167)  and  A168 );
 a34917a <=( A169  and  a34916a );
 a34920a <=( (not A201)  and  A166 );
 a34923a <=( (not A232)  and  A202 );
 a34924a <=( a34923a  and  a34920a );
 a34925a <=( a34924a  and  a34917a );
 a34928a <=( (not A234)  and  A233 );
 a34931a <=( (not A236)  and  (not A235) );
 a34932a <=( a34931a  and  a34928a );
 a34935a <=( A266  and  (not A265) );
 a34938a <=( A269  and  A267 );
 a34939a <=( a34938a  and  a34935a );
 a34940a <=( a34939a  and  a34932a );
 a34944a <=( (not A167)  and  A168 );
 a34945a <=( A169  and  a34944a );
 a34948a <=( (not A201)  and  A166 );
 a34951a <=( (not A232)  and  A202 );
 a34952a <=( a34951a  and  a34948a );
 a34953a <=( a34952a  and  a34945a );
 a34956a <=( (not A234)  and  A233 );
 a34959a <=( (not A236)  and  (not A235) );
 a34960a <=( a34959a  and  a34956a );
 a34963a <=( (not A266)  and  A265 );
 a34966a <=( A268  and  A267 );
 a34967a <=( a34966a  and  a34963a );
 a34968a <=( a34967a  and  a34960a );
 a34972a <=( (not A167)  and  A168 );
 a34973a <=( A169  and  a34972a );
 a34976a <=( (not A201)  and  A166 );
 a34979a <=( (not A232)  and  A202 );
 a34980a <=( a34979a  and  a34976a );
 a34981a <=( a34980a  and  a34973a );
 a34984a <=( (not A234)  and  A233 );
 a34987a <=( (not A236)  and  (not A235) );
 a34988a <=( a34987a  and  a34984a );
 a34991a <=( (not A266)  and  A265 );
 a34994a <=( A269  and  A267 );
 a34995a <=( a34994a  and  a34991a );
 a34996a <=( a34995a  and  a34988a );
 a35000a <=( (not A167)  and  A168 );
 a35001a <=( A169  and  a35000a );
 a35004a <=( (not A201)  and  A166 );
 a35007a <=( A232  and  A202 );
 a35008a <=( a35007a  and  a35004a );
 a35009a <=( a35008a  and  a35001a );
 a35012a <=( A234  and  (not A233) );
 a35015a <=( A298  and  A235 );
 a35016a <=( a35015a  and  a35012a );
 a35019a <=( (not A300)  and  (not A299) );
 a35022a <=( (not A302)  and  (not A301) );
 a35023a <=( a35022a  and  a35019a );
 a35024a <=( a35023a  and  a35016a );
 a35028a <=( (not A167)  and  A168 );
 a35029a <=( A169  and  a35028a );
 a35032a <=( (not A201)  and  A166 );
 a35035a <=( A232  and  A202 );
 a35036a <=( a35035a  and  a35032a );
 a35037a <=( a35036a  and  a35029a );
 a35040a <=( A234  and  (not A233) );
 a35043a <=( (not A298)  and  A235 );
 a35044a <=( a35043a  and  a35040a );
 a35047a <=( (not A300)  and  A299 );
 a35050a <=( (not A302)  and  (not A301) );
 a35051a <=( a35050a  and  a35047a );
 a35052a <=( a35051a  and  a35044a );
 a35056a <=( (not A167)  and  A168 );
 a35057a <=( A169  and  a35056a );
 a35060a <=( (not A201)  and  A166 );
 a35063a <=( A232  and  A202 );
 a35064a <=( a35063a  and  a35060a );
 a35065a <=( a35064a  and  a35057a );
 a35068a <=( A234  and  (not A233) );
 a35071a <=( (not A265)  and  A235 );
 a35072a <=( a35071a  and  a35068a );
 a35075a <=( (not A267)  and  A266 );
 a35078a <=( (not A269)  and  (not A268) );
 a35079a <=( a35078a  and  a35075a );
 a35080a <=( a35079a  and  a35072a );
 a35084a <=( (not A167)  and  A168 );
 a35085a <=( A169  and  a35084a );
 a35088a <=( (not A201)  and  A166 );
 a35091a <=( A232  and  A202 );
 a35092a <=( a35091a  and  a35088a );
 a35093a <=( a35092a  and  a35085a );
 a35096a <=( A234  and  (not A233) );
 a35099a <=( A265  and  A235 );
 a35100a <=( a35099a  and  a35096a );
 a35103a <=( (not A267)  and  (not A266) );
 a35106a <=( (not A269)  and  (not A268) );
 a35107a <=( a35106a  and  a35103a );
 a35108a <=( a35107a  and  a35100a );
 a35112a <=( (not A167)  and  A168 );
 a35113a <=( A169  and  a35112a );
 a35116a <=( (not A201)  and  A166 );
 a35119a <=( A232  and  A202 );
 a35120a <=( a35119a  and  a35116a );
 a35121a <=( a35120a  and  a35113a );
 a35124a <=( A234  and  (not A233) );
 a35127a <=( A298  and  A236 );
 a35128a <=( a35127a  and  a35124a );
 a35131a <=( (not A300)  and  (not A299) );
 a35134a <=( (not A302)  and  (not A301) );
 a35135a <=( a35134a  and  a35131a );
 a35136a <=( a35135a  and  a35128a );
 a35140a <=( (not A167)  and  A168 );
 a35141a <=( A169  and  a35140a );
 a35144a <=( (not A201)  and  A166 );
 a35147a <=( A232  and  A202 );
 a35148a <=( a35147a  and  a35144a );
 a35149a <=( a35148a  and  a35141a );
 a35152a <=( A234  and  (not A233) );
 a35155a <=( (not A298)  and  A236 );
 a35156a <=( a35155a  and  a35152a );
 a35159a <=( (not A300)  and  A299 );
 a35162a <=( (not A302)  and  (not A301) );
 a35163a <=( a35162a  and  a35159a );
 a35164a <=( a35163a  and  a35156a );
 a35168a <=( (not A167)  and  A168 );
 a35169a <=( A169  and  a35168a );
 a35172a <=( (not A201)  and  A166 );
 a35175a <=( A232  and  A202 );
 a35176a <=( a35175a  and  a35172a );
 a35177a <=( a35176a  and  a35169a );
 a35180a <=( A234  and  (not A233) );
 a35183a <=( (not A265)  and  A236 );
 a35184a <=( a35183a  and  a35180a );
 a35187a <=( (not A267)  and  A266 );
 a35190a <=( (not A269)  and  (not A268) );
 a35191a <=( a35190a  and  a35187a );
 a35192a <=( a35191a  and  a35184a );
 a35196a <=( (not A167)  and  A168 );
 a35197a <=( A169  and  a35196a );
 a35200a <=( (not A201)  and  A166 );
 a35203a <=( A232  and  A202 );
 a35204a <=( a35203a  and  a35200a );
 a35205a <=( a35204a  and  a35197a );
 a35208a <=( A234  and  (not A233) );
 a35211a <=( A265  and  A236 );
 a35212a <=( a35211a  and  a35208a );
 a35215a <=( (not A267)  and  (not A266) );
 a35218a <=( (not A269)  and  (not A268) );
 a35219a <=( a35218a  and  a35215a );
 a35220a <=( a35219a  and  a35212a );
 a35224a <=( (not A167)  and  A168 );
 a35225a <=( A169  and  a35224a );
 a35228a <=( (not A201)  and  A166 );
 a35231a <=( A232  and  A202 );
 a35232a <=( a35231a  and  a35228a );
 a35233a <=( a35232a  and  a35225a );
 a35236a <=( (not A234)  and  (not A233) );
 a35239a <=( (not A236)  and  (not A235) );
 a35240a <=( a35239a  and  a35236a );
 a35243a <=( (not A299)  and  A298 );
 a35246a <=( A301  and  A300 );
 a35247a <=( a35246a  and  a35243a );
 a35248a <=( a35247a  and  a35240a );
 a35252a <=( (not A167)  and  A168 );
 a35253a <=( A169  and  a35252a );
 a35256a <=( (not A201)  and  A166 );
 a35259a <=( A232  and  A202 );
 a35260a <=( a35259a  and  a35256a );
 a35261a <=( a35260a  and  a35253a );
 a35264a <=( (not A234)  and  (not A233) );
 a35267a <=( (not A236)  and  (not A235) );
 a35268a <=( a35267a  and  a35264a );
 a35271a <=( (not A299)  and  A298 );
 a35274a <=( A302  and  A300 );
 a35275a <=( a35274a  and  a35271a );
 a35276a <=( a35275a  and  a35268a );
 a35280a <=( (not A167)  and  A168 );
 a35281a <=( A169  and  a35280a );
 a35284a <=( (not A201)  and  A166 );
 a35287a <=( A232  and  A202 );
 a35288a <=( a35287a  and  a35284a );
 a35289a <=( a35288a  and  a35281a );
 a35292a <=( (not A234)  and  (not A233) );
 a35295a <=( (not A236)  and  (not A235) );
 a35296a <=( a35295a  and  a35292a );
 a35299a <=( A299  and  (not A298) );
 a35302a <=( A301  and  A300 );
 a35303a <=( a35302a  and  a35299a );
 a35304a <=( a35303a  and  a35296a );
 a35308a <=( (not A167)  and  A168 );
 a35309a <=( A169  and  a35308a );
 a35312a <=( (not A201)  and  A166 );
 a35315a <=( A232  and  A202 );
 a35316a <=( a35315a  and  a35312a );
 a35317a <=( a35316a  and  a35309a );
 a35320a <=( (not A234)  and  (not A233) );
 a35323a <=( (not A236)  and  (not A235) );
 a35324a <=( a35323a  and  a35320a );
 a35327a <=( A299  and  (not A298) );
 a35330a <=( A302  and  A300 );
 a35331a <=( a35330a  and  a35327a );
 a35332a <=( a35331a  and  a35324a );
 a35336a <=( (not A167)  and  A168 );
 a35337a <=( A169  and  a35336a );
 a35340a <=( (not A201)  and  A166 );
 a35343a <=( A232  and  A202 );
 a35344a <=( a35343a  and  a35340a );
 a35345a <=( a35344a  and  a35337a );
 a35348a <=( (not A234)  and  (not A233) );
 a35351a <=( (not A236)  and  (not A235) );
 a35352a <=( a35351a  and  a35348a );
 a35355a <=( A266  and  (not A265) );
 a35358a <=( A268  and  A267 );
 a35359a <=( a35358a  and  a35355a );
 a35360a <=( a35359a  and  a35352a );
 a35364a <=( (not A167)  and  A168 );
 a35365a <=( A169  and  a35364a );
 a35368a <=( (not A201)  and  A166 );
 a35371a <=( A232  and  A202 );
 a35372a <=( a35371a  and  a35368a );
 a35373a <=( a35372a  and  a35365a );
 a35376a <=( (not A234)  and  (not A233) );
 a35379a <=( (not A236)  and  (not A235) );
 a35380a <=( a35379a  and  a35376a );
 a35383a <=( A266  and  (not A265) );
 a35386a <=( A269  and  A267 );
 a35387a <=( a35386a  and  a35383a );
 a35388a <=( a35387a  and  a35380a );
 a35392a <=( (not A167)  and  A168 );
 a35393a <=( A169  and  a35392a );
 a35396a <=( (not A201)  and  A166 );
 a35399a <=( A232  and  A202 );
 a35400a <=( a35399a  and  a35396a );
 a35401a <=( a35400a  and  a35393a );
 a35404a <=( (not A234)  and  (not A233) );
 a35407a <=( (not A236)  and  (not A235) );
 a35408a <=( a35407a  and  a35404a );
 a35411a <=( (not A266)  and  A265 );
 a35414a <=( A268  and  A267 );
 a35415a <=( a35414a  and  a35411a );
 a35416a <=( a35415a  and  a35408a );
 a35420a <=( (not A167)  and  A168 );
 a35421a <=( A169  and  a35420a );
 a35424a <=( (not A201)  and  A166 );
 a35427a <=( A232  and  A202 );
 a35428a <=( a35427a  and  a35424a );
 a35429a <=( a35428a  and  a35421a );
 a35432a <=( (not A234)  and  (not A233) );
 a35435a <=( (not A236)  and  (not A235) );
 a35436a <=( a35435a  and  a35432a );
 a35439a <=( (not A266)  and  A265 );
 a35442a <=( A269  and  A267 );
 a35443a <=( a35442a  and  a35439a );
 a35444a <=( a35443a  and  a35436a );
 a35448a <=( (not A167)  and  A168 );
 a35449a <=( A169  and  a35448a );
 a35452a <=( (not A201)  and  A166 );
 a35455a <=( (not A232)  and  A203 );
 a35456a <=( a35455a  and  a35452a );
 a35457a <=( a35456a  and  a35449a );
 a35460a <=( A234  and  A233 );
 a35463a <=( A298  and  A235 );
 a35464a <=( a35463a  and  a35460a );
 a35467a <=( (not A300)  and  (not A299) );
 a35470a <=( (not A302)  and  (not A301) );
 a35471a <=( a35470a  and  a35467a );
 a35472a <=( a35471a  and  a35464a );
 a35476a <=( (not A167)  and  A168 );
 a35477a <=( A169  and  a35476a );
 a35480a <=( (not A201)  and  A166 );
 a35483a <=( (not A232)  and  A203 );
 a35484a <=( a35483a  and  a35480a );
 a35485a <=( a35484a  and  a35477a );
 a35488a <=( A234  and  A233 );
 a35491a <=( (not A298)  and  A235 );
 a35492a <=( a35491a  and  a35488a );
 a35495a <=( (not A300)  and  A299 );
 a35498a <=( (not A302)  and  (not A301) );
 a35499a <=( a35498a  and  a35495a );
 a35500a <=( a35499a  and  a35492a );
 a35504a <=( (not A167)  and  A168 );
 a35505a <=( A169  and  a35504a );
 a35508a <=( (not A201)  and  A166 );
 a35511a <=( (not A232)  and  A203 );
 a35512a <=( a35511a  and  a35508a );
 a35513a <=( a35512a  and  a35505a );
 a35516a <=( A234  and  A233 );
 a35519a <=( (not A265)  and  A235 );
 a35520a <=( a35519a  and  a35516a );
 a35523a <=( (not A267)  and  A266 );
 a35526a <=( (not A269)  and  (not A268) );
 a35527a <=( a35526a  and  a35523a );
 a35528a <=( a35527a  and  a35520a );
 a35532a <=( (not A167)  and  A168 );
 a35533a <=( A169  and  a35532a );
 a35536a <=( (not A201)  and  A166 );
 a35539a <=( (not A232)  and  A203 );
 a35540a <=( a35539a  and  a35536a );
 a35541a <=( a35540a  and  a35533a );
 a35544a <=( A234  and  A233 );
 a35547a <=( A265  and  A235 );
 a35548a <=( a35547a  and  a35544a );
 a35551a <=( (not A267)  and  (not A266) );
 a35554a <=( (not A269)  and  (not A268) );
 a35555a <=( a35554a  and  a35551a );
 a35556a <=( a35555a  and  a35548a );
 a35560a <=( (not A167)  and  A168 );
 a35561a <=( A169  and  a35560a );
 a35564a <=( (not A201)  and  A166 );
 a35567a <=( (not A232)  and  A203 );
 a35568a <=( a35567a  and  a35564a );
 a35569a <=( a35568a  and  a35561a );
 a35572a <=( A234  and  A233 );
 a35575a <=( A298  and  A236 );
 a35576a <=( a35575a  and  a35572a );
 a35579a <=( (not A300)  and  (not A299) );
 a35582a <=( (not A302)  and  (not A301) );
 a35583a <=( a35582a  and  a35579a );
 a35584a <=( a35583a  and  a35576a );
 a35588a <=( (not A167)  and  A168 );
 a35589a <=( A169  and  a35588a );
 a35592a <=( (not A201)  and  A166 );
 a35595a <=( (not A232)  and  A203 );
 a35596a <=( a35595a  and  a35592a );
 a35597a <=( a35596a  and  a35589a );
 a35600a <=( A234  and  A233 );
 a35603a <=( (not A298)  and  A236 );
 a35604a <=( a35603a  and  a35600a );
 a35607a <=( (not A300)  and  A299 );
 a35610a <=( (not A302)  and  (not A301) );
 a35611a <=( a35610a  and  a35607a );
 a35612a <=( a35611a  and  a35604a );
 a35616a <=( (not A167)  and  A168 );
 a35617a <=( A169  and  a35616a );
 a35620a <=( (not A201)  and  A166 );
 a35623a <=( (not A232)  and  A203 );
 a35624a <=( a35623a  and  a35620a );
 a35625a <=( a35624a  and  a35617a );
 a35628a <=( A234  and  A233 );
 a35631a <=( (not A265)  and  A236 );
 a35632a <=( a35631a  and  a35628a );
 a35635a <=( (not A267)  and  A266 );
 a35638a <=( (not A269)  and  (not A268) );
 a35639a <=( a35638a  and  a35635a );
 a35640a <=( a35639a  and  a35632a );
 a35644a <=( (not A167)  and  A168 );
 a35645a <=( A169  and  a35644a );
 a35648a <=( (not A201)  and  A166 );
 a35651a <=( (not A232)  and  A203 );
 a35652a <=( a35651a  and  a35648a );
 a35653a <=( a35652a  and  a35645a );
 a35656a <=( A234  and  A233 );
 a35659a <=( A265  and  A236 );
 a35660a <=( a35659a  and  a35656a );
 a35663a <=( (not A267)  and  (not A266) );
 a35666a <=( (not A269)  and  (not A268) );
 a35667a <=( a35666a  and  a35663a );
 a35668a <=( a35667a  and  a35660a );
 a35672a <=( (not A167)  and  A168 );
 a35673a <=( A169  and  a35672a );
 a35676a <=( (not A201)  and  A166 );
 a35679a <=( (not A232)  and  A203 );
 a35680a <=( a35679a  and  a35676a );
 a35681a <=( a35680a  and  a35673a );
 a35684a <=( (not A234)  and  A233 );
 a35687a <=( (not A236)  and  (not A235) );
 a35688a <=( a35687a  and  a35684a );
 a35691a <=( (not A299)  and  A298 );
 a35694a <=( A301  and  A300 );
 a35695a <=( a35694a  and  a35691a );
 a35696a <=( a35695a  and  a35688a );
 a35700a <=( (not A167)  and  A168 );
 a35701a <=( A169  and  a35700a );
 a35704a <=( (not A201)  and  A166 );
 a35707a <=( (not A232)  and  A203 );
 a35708a <=( a35707a  and  a35704a );
 a35709a <=( a35708a  and  a35701a );
 a35712a <=( (not A234)  and  A233 );
 a35715a <=( (not A236)  and  (not A235) );
 a35716a <=( a35715a  and  a35712a );
 a35719a <=( (not A299)  and  A298 );
 a35722a <=( A302  and  A300 );
 a35723a <=( a35722a  and  a35719a );
 a35724a <=( a35723a  and  a35716a );
 a35728a <=( (not A167)  and  A168 );
 a35729a <=( A169  and  a35728a );
 a35732a <=( (not A201)  and  A166 );
 a35735a <=( (not A232)  and  A203 );
 a35736a <=( a35735a  and  a35732a );
 a35737a <=( a35736a  and  a35729a );
 a35740a <=( (not A234)  and  A233 );
 a35743a <=( (not A236)  and  (not A235) );
 a35744a <=( a35743a  and  a35740a );
 a35747a <=( A299  and  (not A298) );
 a35750a <=( A301  and  A300 );
 a35751a <=( a35750a  and  a35747a );
 a35752a <=( a35751a  and  a35744a );
 a35756a <=( (not A167)  and  A168 );
 a35757a <=( A169  and  a35756a );
 a35760a <=( (not A201)  and  A166 );
 a35763a <=( (not A232)  and  A203 );
 a35764a <=( a35763a  and  a35760a );
 a35765a <=( a35764a  and  a35757a );
 a35768a <=( (not A234)  and  A233 );
 a35771a <=( (not A236)  and  (not A235) );
 a35772a <=( a35771a  and  a35768a );
 a35775a <=( A299  and  (not A298) );
 a35778a <=( A302  and  A300 );
 a35779a <=( a35778a  and  a35775a );
 a35780a <=( a35779a  and  a35772a );
 a35784a <=( (not A167)  and  A168 );
 a35785a <=( A169  and  a35784a );
 a35788a <=( (not A201)  and  A166 );
 a35791a <=( (not A232)  and  A203 );
 a35792a <=( a35791a  and  a35788a );
 a35793a <=( a35792a  and  a35785a );
 a35796a <=( (not A234)  and  A233 );
 a35799a <=( (not A236)  and  (not A235) );
 a35800a <=( a35799a  and  a35796a );
 a35803a <=( A266  and  (not A265) );
 a35806a <=( A268  and  A267 );
 a35807a <=( a35806a  and  a35803a );
 a35808a <=( a35807a  and  a35800a );
 a35812a <=( (not A167)  and  A168 );
 a35813a <=( A169  and  a35812a );
 a35816a <=( (not A201)  and  A166 );
 a35819a <=( (not A232)  and  A203 );
 a35820a <=( a35819a  and  a35816a );
 a35821a <=( a35820a  and  a35813a );
 a35824a <=( (not A234)  and  A233 );
 a35827a <=( (not A236)  and  (not A235) );
 a35828a <=( a35827a  and  a35824a );
 a35831a <=( A266  and  (not A265) );
 a35834a <=( A269  and  A267 );
 a35835a <=( a35834a  and  a35831a );
 a35836a <=( a35835a  and  a35828a );
 a35840a <=( (not A167)  and  A168 );
 a35841a <=( A169  and  a35840a );
 a35844a <=( (not A201)  and  A166 );
 a35847a <=( (not A232)  and  A203 );
 a35848a <=( a35847a  and  a35844a );
 a35849a <=( a35848a  and  a35841a );
 a35852a <=( (not A234)  and  A233 );
 a35855a <=( (not A236)  and  (not A235) );
 a35856a <=( a35855a  and  a35852a );
 a35859a <=( (not A266)  and  A265 );
 a35862a <=( A268  and  A267 );
 a35863a <=( a35862a  and  a35859a );
 a35864a <=( a35863a  and  a35856a );
 a35868a <=( (not A167)  and  A168 );
 a35869a <=( A169  and  a35868a );
 a35872a <=( (not A201)  and  A166 );
 a35875a <=( (not A232)  and  A203 );
 a35876a <=( a35875a  and  a35872a );
 a35877a <=( a35876a  and  a35869a );
 a35880a <=( (not A234)  and  A233 );
 a35883a <=( (not A236)  and  (not A235) );
 a35884a <=( a35883a  and  a35880a );
 a35887a <=( (not A266)  and  A265 );
 a35890a <=( A269  and  A267 );
 a35891a <=( a35890a  and  a35887a );
 a35892a <=( a35891a  and  a35884a );
 a35896a <=( (not A167)  and  A168 );
 a35897a <=( A169  and  a35896a );
 a35900a <=( (not A201)  and  A166 );
 a35903a <=( A232  and  A203 );
 a35904a <=( a35903a  and  a35900a );
 a35905a <=( a35904a  and  a35897a );
 a35908a <=( A234  and  (not A233) );
 a35911a <=( A298  and  A235 );
 a35912a <=( a35911a  and  a35908a );
 a35915a <=( (not A300)  and  (not A299) );
 a35918a <=( (not A302)  and  (not A301) );
 a35919a <=( a35918a  and  a35915a );
 a35920a <=( a35919a  and  a35912a );
 a35924a <=( (not A167)  and  A168 );
 a35925a <=( A169  and  a35924a );
 a35928a <=( (not A201)  and  A166 );
 a35931a <=( A232  and  A203 );
 a35932a <=( a35931a  and  a35928a );
 a35933a <=( a35932a  and  a35925a );
 a35936a <=( A234  and  (not A233) );
 a35939a <=( (not A298)  and  A235 );
 a35940a <=( a35939a  and  a35936a );
 a35943a <=( (not A300)  and  A299 );
 a35946a <=( (not A302)  and  (not A301) );
 a35947a <=( a35946a  and  a35943a );
 a35948a <=( a35947a  and  a35940a );
 a35952a <=( (not A167)  and  A168 );
 a35953a <=( A169  and  a35952a );
 a35956a <=( (not A201)  and  A166 );
 a35959a <=( A232  and  A203 );
 a35960a <=( a35959a  and  a35956a );
 a35961a <=( a35960a  and  a35953a );
 a35964a <=( A234  and  (not A233) );
 a35967a <=( (not A265)  and  A235 );
 a35968a <=( a35967a  and  a35964a );
 a35971a <=( (not A267)  and  A266 );
 a35974a <=( (not A269)  and  (not A268) );
 a35975a <=( a35974a  and  a35971a );
 a35976a <=( a35975a  and  a35968a );
 a35980a <=( (not A167)  and  A168 );
 a35981a <=( A169  and  a35980a );
 a35984a <=( (not A201)  and  A166 );
 a35987a <=( A232  and  A203 );
 a35988a <=( a35987a  and  a35984a );
 a35989a <=( a35988a  and  a35981a );
 a35992a <=( A234  and  (not A233) );
 a35995a <=( A265  and  A235 );
 a35996a <=( a35995a  and  a35992a );
 a35999a <=( (not A267)  and  (not A266) );
 a36002a <=( (not A269)  and  (not A268) );
 a36003a <=( a36002a  and  a35999a );
 a36004a <=( a36003a  and  a35996a );
 a36008a <=( (not A167)  and  A168 );
 a36009a <=( A169  and  a36008a );
 a36012a <=( (not A201)  and  A166 );
 a36015a <=( A232  and  A203 );
 a36016a <=( a36015a  and  a36012a );
 a36017a <=( a36016a  and  a36009a );
 a36020a <=( A234  and  (not A233) );
 a36023a <=( A298  and  A236 );
 a36024a <=( a36023a  and  a36020a );
 a36027a <=( (not A300)  and  (not A299) );
 a36030a <=( (not A302)  and  (not A301) );
 a36031a <=( a36030a  and  a36027a );
 a36032a <=( a36031a  and  a36024a );
 a36036a <=( (not A167)  and  A168 );
 a36037a <=( A169  and  a36036a );
 a36040a <=( (not A201)  and  A166 );
 a36043a <=( A232  and  A203 );
 a36044a <=( a36043a  and  a36040a );
 a36045a <=( a36044a  and  a36037a );
 a36048a <=( A234  and  (not A233) );
 a36051a <=( (not A298)  and  A236 );
 a36052a <=( a36051a  and  a36048a );
 a36055a <=( (not A300)  and  A299 );
 a36058a <=( (not A302)  and  (not A301) );
 a36059a <=( a36058a  and  a36055a );
 a36060a <=( a36059a  and  a36052a );
 a36064a <=( (not A167)  and  A168 );
 a36065a <=( A169  and  a36064a );
 a36068a <=( (not A201)  and  A166 );
 a36071a <=( A232  and  A203 );
 a36072a <=( a36071a  and  a36068a );
 a36073a <=( a36072a  and  a36065a );
 a36076a <=( A234  and  (not A233) );
 a36079a <=( (not A265)  and  A236 );
 a36080a <=( a36079a  and  a36076a );
 a36083a <=( (not A267)  and  A266 );
 a36086a <=( (not A269)  and  (not A268) );
 a36087a <=( a36086a  and  a36083a );
 a36088a <=( a36087a  and  a36080a );
 a36092a <=( (not A167)  and  A168 );
 a36093a <=( A169  and  a36092a );
 a36096a <=( (not A201)  and  A166 );
 a36099a <=( A232  and  A203 );
 a36100a <=( a36099a  and  a36096a );
 a36101a <=( a36100a  and  a36093a );
 a36104a <=( A234  and  (not A233) );
 a36107a <=( A265  and  A236 );
 a36108a <=( a36107a  and  a36104a );
 a36111a <=( (not A267)  and  (not A266) );
 a36114a <=( (not A269)  and  (not A268) );
 a36115a <=( a36114a  and  a36111a );
 a36116a <=( a36115a  and  a36108a );
 a36120a <=( (not A167)  and  A168 );
 a36121a <=( A169  and  a36120a );
 a36124a <=( (not A201)  and  A166 );
 a36127a <=( A232  and  A203 );
 a36128a <=( a36127a  and  a36124a );
 a36129a <=( a36128a  and  a36121a );
 a36132a <=( (not A234)  and  (not A233) );
 a36135a <=( (not A236)  and  (not A235) );
 a36136a <=( a36135a  and  a36132a );
 a36139a <=( (not A299)  and  A298 );
 a36142a <=( A301  and  A300 );
 a36143a <=( a36142a  and  a36139a );
 a36144a <=( a36143a  and  a36136a );
 a36148a <=( (not A167)  and  A168 );
 a36149a <=( A169  and  a36148a );
 a36152a <=( (not A201)  and  A166 );
 a36155a <=( A232  and  A203 );
 a36156a <=( a36155a  and  a36152a );
 a36157a <=( a36156a  and  a36149a );
 a36160a <=( (not A234)  and  (not A233) );
 a36163a <=( (not A236)  and  (not A235) );
 a36164a <=( a36163a  and  a36160a );
 a36167a <=( (not A299)  and  A298 );
 a36170a <=( A302  and  A300 );
 a36171a <=( a36170a  and  a36167a );
 a36172a <=( a36171a  and  a36164a );
 a36176a <=( (not A167)  and  A168 );
 a36177a <=( A169  and  a36176a );
 a36180a <=( (not A201)  and  A166 );
 a36183a <=( A232  and  A203 );
 a36184a <=( a36183a  and  a36180a );
 a36185a <=( a36184a  and  a36177a );
 a36188a <=( (not A234)  and  (not A233) );
 a36191a <=( (not A236)  and  (not A235) );
 a36192a <=( a36191a  and  a36188a );
 a36195a <=( A299  and  (not A298) );
 a36198a <=( A301  and  A300 );
 a36199a <=( a36198a  and  a36195a );
 a36200a <=( a36199a  and  a36192a );
 a36204a <=( (not A167)  and  A168 );
 a36205a <=( A169  and  a36204a );
 a36208a <=( (not A201)  and  A166 );
 a36211a <=( A232  and  A203 );
 a36212a <=( a36211a  and  a36208a );
 a36213a <=( a36212a  and  a36205a );
 a36216a <=( (not A234)  and  (not A233) );
 a36219a <=( (not A236)  and  (not A235) );
 a36220a <=( a36219a  and  a36216a );
 a36223a <=( A299  and  (not A298) );
 a36226a <=( A302  and  A300 );
 a36227a <=( a36226a  and  a36223a );
 a36228a <=( a36227a  and  a36220a );
 a36232a <=( (not A167)  and  A168 );
 a36233a <=( A169  and  a36232a );
 a36236a <=( (not A201)  and  A166 );
 a36239a <=( A232  and  A203 );
 a36240a <=( a36239a  and  a36236a );
 a36241a <=( a36240a  and  a36233a );
 a36244a <=( (not A234)  and  (not A233) );
 a36247a <=( (not A236)  and  (not A235) );
 a36248a <=( a36247a  and  a36244a );
 a36251a <=( A266  and  (not A265) );
 a36254a <=( A268  and  A267 );
 a36255a <=( a36254a  and  a36251a );
 a36256a <=( a36255a  and  a36248a );
 a36260a <=( (not A167)  and  A168 );
 a36261a <=( A169  and  a36260a );
 a36264a <=( (not A201)  and  A166 );
 a36267a <=( A232  and  A203 );
 a36268a <=( a36267a  and  a36264a );
 a36269a <=( a36268a  and  a36261a );
 a36272a <=( (not A234)  and  (not A233) );
 a36275a <=( (not A236)  and  (not A235) );
 a36276a <=( a36275a  and  a36272a );
 a36279a <=( A266  and  (not A265) );
 a36282a <=( A269  and  A267 );
 a36283a <=( a36282a  and  a36279a );
 a36284a <=( a36283a  and  a36276a );
 a36288a <=( (not A167)  and  A168 );
 a36289a <=( A169  and  a36288a );
 a36292a <=( (not A201)  and  A166 );
 a36295a <=( A232  and  A203 );
 a36296a <=( a36295a  and  a36292a );
 a36297a <=( a36296a  and  a36289a );
 a36300a <=( (not A234)  and  (not A233) );
 a36303a <=( (not A236)  and  (not A235) );
 a36304a <=( a36303a  and  a36300a );
 a36307a <=( (not A266)  and  A265 );
 a36310a <=( A268  and  A267 );
 a36311a <=( a36310a  and  a36307a );
 a36312a <=( a36311a  and  a36304a );
 a36316a <=( (not A167)  and  A168 );
 a36317a <=( A169  and  a36316a );
 a36320a <=( (not A201)  and  A166 );
 a36323a <=( A232  and  A203 );
 a36324a <=( a36323a  and  a36320a );
 a36325a <=( a36324a  and  a36317a );
 a36328a <=( (not A234)  and  (not A233) );
 a36331a <=( (not A236)  and  (not A235) );
 a36332a <=( a36331a  and  a36328a );
 a36335a <=( (not A266)  and  A265 );
 a36338a <=( A269  and  A267 );
 a36339a <=( a36338a  and  a36335a );
 a36340a <=( a36339a  and  a36332a );
 a36344a <=( (not A167)  and  A168 );
 a36345a <=( A169  and  a36344a );
 a36348a <=( A199  and  A166 );
 a36351a <=( (not A232)  and  A200 );
 a36352a <=( a36351a  and  a36348a );
 a36353a <=( a36352a  and  a36345a );
 a36356a <=( A234  and  A233 );
 a36359a <=( A298  and  A235 );
 a36360a <=( a36359a  and  a36356a );
 a36363a <=( (not A300)  and  (not A299) );
 a36366a <=( (not A302)  and  (not A301) );
 a36367a <=( a36366a  and  a36363a );
 a36368a <=( a36367a  and  a36360a );
 a36372a <=( (not A167)  and  A168 );
 a36373a <=( A169  and  a36372a );
 a36376a <=( A199  and  A166 );
 a36379a <=( (not A232)  and  A200 );
 a36380a <=( a36379a  and  a36376a );
 a36381a <=( a36380a  and  a36373a );
 a36384a <=( A234  and  A233 );
 a36387a <=( (not A298)  and  A235 );
 a36388a <=( a36387a  and  a36384a );
 a36391a <=( (not A300)  and  A299 );
 a36394a <=( (not A302)  and  (not A301) );
 a36395a <=( a36394a  and  a36391a );
 a36396a <=( a36395a  and  a36388a );
 a36400a <=( (not A167)  and  A168 );
 a36401a <=( A169  and  a36400a );
 a36404a <=( A199  and  A166 );
 a36407a <=( (not A232)  and  A200 );
 a36408a <=( a36407a  and  a36404a );
 a36409a <=( a36408a  and  a36401a );
 a36412a <=( A234  and  A233 );
 a36415a <=( (not A265)  and  A235 );
 a36416a <=( a36415a  and  a36412a );
 a36419a <=( (not A267)  and  A266 );
 a36422a <=( (not A269)  and  (not A268) );
 a36423a <=( a36422a  and  a36419a );
 a36424a <=( a36423a  and  a36416a );
 a36428a <=( (not A167)  and  A168 );
 a36429a <=( A169  and  a36428a );
 a36432a <=( A199  and  A166 );
 a36435a <=( (not A232)  and  A200 );
 a36436a <=( a36435a  and  a36432a );
 a36437a <=( a36436a  and  a36429a );
 a36440a <=( A234  and  A233 );
 a36443a <=( A265  and  A235 );
 a36444a <=( a36443a  and  a36440a );
 a36447a <=( (not A267)  and  (not A266) );
 a36450a <=( (not A269)  and  (not A268) );
 a36451a <=( a36450a  and  a36447a );
 a36452a <=( a36451a  and  a36444a );
 a36456a <=( (not A167)  and  A168 );
 a36457a <=( A169  and  a36456a );
 a36460a <=( A199  and  A166 );
 a36463a <=( (not A232)  and  A200 );
 a36464a <=( a36463a  and  a36460a );
 a36465a <=( a36464a  and  a36457a );
 a36468a <=( A234  and  A233 );
 a36471a <=( A298  and  A236 );
 a36472a <=( a36471a  and  a36468a );
 a36475a <=( (not A300)  and  (not A299) );
 a36478a <=( (not A302)  and  (not A301) );
 a36479a <=( a36478a  and  a36475a );
 a36480a <=( a36479a  and  a36472a );
 a36484a <=( (not A167)  and  A168 );
 a36485a <=( A169  and  a36484a );
 a36488a <=( A199  and  A166 );
 a36491a <=( (not A232)  and  A200 );
 a36492a <=( a36491a  and  a36488a );
 a36493a <=( a36492a  and  a36485a );
 a36496a <=( A234  and  A233 );
 a36499a <=( (not A298)  and  A236 );
 a36500a <=( a36499a  and  a36496a );
 a36503a <=( (not A300)  and  A299 );
 a36506a <=( (not A302)  and  (not A301) );
 a36507a <=( a36506a  and  a36503a );
 a36508a <=( a36507a  and  a36500a );
 a36512a <=( (not A167)  and  A168 );
 a36513a <=( A169  and  a36512a );
 a36516a <=( A199  and  A166 );
 a36519a <=( (not A232)  and  A200 );
 a36520a <=( a36519a  and  a36516a );
 a36521a <=( a36520a  and  a36513a );
 a36524a <=( A234  and  A233 );
 a36527a <=( (not A265)  and  A236 );
 a36528a <=( a36527a  and  a36524a );
 a36531a <=( (not A267)  and  A266 );
 a36534a <=( (not A269)  and  (not A268) );
 a36535a <=( a36534a  and  a36531a );
 a36536a <=( a36535a  and  a36528a );
 a36540a <=( (not A167)  and  A168 );
 a36541a <=( A169  and  a36540a );
 a36544a <=( A199  and  A166 );
 a36547a <=( (not A232)  and  A200 );
 a36548a <=( a36547a  and  a36544a );
 a36549a <=( a36548a  and  a36541a );
 a36552a <=( A234  and  A233 );
 a36555a <=( A265  and  A236 );
 a36556a <=( a36555a  and  a36552a );
 a36559a <=( (not A267)  and  (not A266) );
 a36562a <=( (not A269)  and  (not A268) );
 a36563a <=( a36562a  and  a36559a );
 a36564a <=( a36563a  and  a36556a );
 a36568a <=( (not A167)  and  A168 );
 a36569a <=( A169  and  a36568a );
 a36572a <=( A199  and  A166 );
 a36575a <=( (not A232)  and  A200 );
 a36576a <=( a36575a  and  a36572a );
 a36577a <=( a36576a  and  a36569a );
 a36580a <=( (not A234)  and  A233 );
 a36583a <=( (not A236)  and  (not A235) );
 a36584a <=( a36583a  and  a36580a );
 a36587a <=( (not A299)  and  A298 );
 a36590a <=( A301  and  A300 );
 a36591a <=( a36590a  and  a36587a );
 a36592a <=( a36591a  and  a36584a );
 a36596a <=( (not A167)  and  A168 );
 a36597a <=( A169  and  a36596a );
 a36600a <=( A199  and  A166 );
 a36603a <=( (not A232)  and  A200 );
 a36604a <=( a36603a  and  a36600a );
 a36605a <=( a36604a  and  a36597a );
 a36608a <=( (not A234)  and  A233 );
 a36611a <=( (not A236)  and  (not A235) );
 a36612a <=( a36611a  and  a36608a );
 a36615a <=( (not A299)  and  A298 );
 a36618a <=( A302  and  A300 );
 a36619a <=( a36618a  and  a36615a );
 a36620a <=( a36619a  and  a36612a );
 a36624a <=( (not A167)  and  A168 );
 a36625a <=( A169  and  a36624a );
 a36628a <=( A199  and  A166 );
 a36631a <=( (not A232)  and  A200 );
 a36632a <=( a36631a  and  a36628a );
 a36633a <=( a36632a  and  a36625a );
 a36636a <=( (not A234)  and  A233 );
 a36639a <=( (not A236)  and  (not A235) );
 a36640a <=( a36639a  and  a36636a );
 a36643a <=( A299  and  (not A298) );
 a36646a <=( A301  and  A300 );
 a36647a <=( a36646a  and  a36643a );
 a36648a <=( a36647a  and  a36640a );
 a36652a <=( (not A167)  and  A168 );
 a36653a <=( A169  and  a36652a );
 a36656a <=( A199  and  A166 );
 a36659a <=( (not A232)  and  A200 );
 a36660a <=( a36659a  and  a36656a );
 a36661a <=( a36660a  and  a36653a );
 a36664a <=( (not A234)  and  A233 );
 a36667a <=( (not A236)  and  (not A235) );
 a36668a <=( a36667a  and  a36664a );
 a36671a <=( A299  and  (not A298) );
 a36674a <=( A302  and  A300 );
 a36675a <=( a36674a  and  a36671a );
 a36676a <=( a36675a  and  a36668a );
 a36680a <=( (not A167)  and  A168 );
 a36681a <=( A169  and  a36680a );
 a36684a <=( A199  and  A166 );
 a36687a <=( (not A232)  and  A200 );
 a36688a <=( a36687a  and  a36684a );
 a36689a <=( a36688a  and  a36681a );
 a36692a <=( (not A234)  and  A233 );
 a36695a <=( (not A236)  and  (not A235) );
 a36696a <=( a36695a  and  a36692a );
 a36699a <=( A266  and  (not A265) );
 a36702a <=( A268  and  A267 );
 a36703a <=( a36702a  and  a36699a );
 a36704a <=( a36703a  and  a36696a );
 a36708a <=( (not A167)  and  A168 );
 a36709a <=( A169  and  a36708a );
 a36712a <=( A199  and  A166 );
 a36715a <=( (not A232)  and  A200 );
 a36716a <=( a36715a  and  a36712a );
 a36717a <=( a36716a  and  a36709a );
 a36720a <=( (not A234)  and  A233 );
 a36723a <=( (not A236)  and  (not A235) );
 a36724a <=( a36723a  and  a36720a );
 a36727a <=( A266  and  (not A265) );
 a36730a <=( A269  and  A267 );
 a36731a <=( a36730a  and  a36727a );
 a36732a <=( a36731a  and  a36724a );
 a36736a <=( (not A167)  and  A168 );
 a36737a <=( A169  and  a36736a );
 a36740a <=( A199  and  A166 );
 a36743a <=( (not A232)  and  A200 );
 a36744a <=( a36743a  and  a36740a );
 a36745a <=( a36744a  and  a36737a );
 a36748a <=( (not A234)  and  A233 );
 a36751a <=( (not A236)  and  (not A235) );
 a36752a <=( a36751a  and  a36748a );
 a36755a <=( (not A266)  and  A265 );
 a36758a <=( A268  and  A267 );
 a36759a <=( a36758a  and  a36755a );
 a36760a <=( a36759a  and  a36752a );
 a36764a <=( (not A167)  and  A168 );
 a36765a <=( A169  and  a36764a );
 a36768a <=( A199  and  A166 );
 a36771a <=( (not A232)  and  A200 );
 a36772a <=( a36771a  and  a36768a );
 a36773a <=( a36772a  and  a36765a );
 a36776a <=( (not A234)  and  A233 );
 a36779a <=( (not A236)  and  (not A235) );
 a36780a <=( a36779a  and  a36776a );
 a36783a <=( (not A266)  and  A265 );
 a36786a <=( A269  and  A267 );
 a36787a <=( a36786a  and  a36783a );
 a36788a <=( a36787a  and  a36780a );
 a36792a <=( (not A167)  and  A168 );
 a36793a <=( A169  and  a36792a );
 a36796a <=( A199  and  A166 );
 a36799a <=( A232  and  A200 );
 a36800a <=( a36799a  and  a36796a );
 a36801a <=( a36800a  and  a36793a );
 a36804a <=( A234  and  (not A233) );
 a36807a <=( A298  and  A235 );
 a36808a <=( a36807a  and  a36804a );
 a36811a <=( (not A300)  and  (not A299) );
 a36814a <=( (not A302)  and  (not A301) );
 a36815a <=( a36814a  and  a36811a );
 a36816a <=( a36815a  and  a36808a );
 a36820a <=( (not A167)  and  A168 );
 a36821a <=( A169  and  a36820a );
 a36824a <=( A199  and  A166 );
 a36827a <=( A232  and  A200 );
 a36828a <=( a36827a  and  a36824a );
 a36829a <=( a36828a  and  a36821a );
 a36832a <=( A234  and  (not A233) );
 a36835a <=( (not A298)  and  A235 );
 a36836a <=( a36835a  and  a36832a );
 a36839a <=( (not A300)  and  A299 );
 a36842a <=( (not A302)  and  (not A301) );
 a36843a <=( a36842a  and  a36839a );
 a36844a <=( a36843a  and  a36836a );
 a36848a <=( (not A167)  and  A168 );
 a36849a <=( A169  and  a36848a );
 a36852a <=( A199  and  A166 );
 a36855a <=( A232  and  A200 );
 a36856a <=( a36855a  and  a36852a );
 a36857a <=( a36856a  and  a36849a );
 a36860a <=( A234  and  (not A233) );
 a36863a <=( (not A265)  and  A235 );
 a36864a <=( a36863a  and  a36860a );
 a36867a <=( (not A267)  and  A266 );
 a36870a <=( (not A269)  and  (not A268) );
 a36871a <=( a36870a  and  a36867a );
 a36872a <=( a36871a  and  a36864a );
 a36876a <=( (not A167)  and  A168 );
 a36877a <=( A169  and  a36876a );
 a36880a <=( A199  and  A166 );
 a36883a <=( A232  and  A200 );
 a36884a <=( a36883a  and  a36880a );
 a36885a <=( a36884a  and  a36877a );
 a36888a <=( A234  and  (not A233) );
 a36891a <=( A265  and  A235 );
 a36892a <=( a36891a  and  a36888a );
 a36895a <=( (not A267)  and  (not A266) );
 a36898a <=( (not A269)  and  (not A268) );
 a36899a <=( a36898a  and  a36895a );
 a36900a <=( a36899a  and  a36892a );
 a36904a <=( (not A167)  and  A168 );
 a36905a <=( A169  and  a36904a );
 a36908a <=( A199  and  A166 );
 a36911a <=( A232  and  A200 );
 a36912a <=( a36911a  and  a36908a );
 a36913a <=( a36912a  and  a36905a );
 a36916a <=( A234  and  (not A233) );
 a36919a <=( A298  and  A236 );
 a36920a <=( a36919a  and  a36916a );
 a36923a <=( (not A300)  and  (not A299) );
 a36926a <=( (not A302)  and  (not A301) );
 a36927a <=( a36926a  and  a36923a );
 a36928a <=( a36927a  and  a36920a );
 a36932a <=( (not A167)  and  A168 );
 a36933a <=( A169  and  a36932a );
 a36936a <=( A199  and  A166 );
 a36939a <=( A232  and  A200 );
 a36940a <=( a36939a  and  a36936a );
 a36941a <=( a36940a  and  a36933a );
 a36944a <=( A234  and  (not A233) );
 a36947a <=( (not A298)  and  A236 );
 a36948a <=( a36947a  and  a36944a );
 a36951a <=( (not A300)  and  A299 );
 a36954a <=( (not A302)  and  (not A301) );
 a36955a <=( a36954a  and  a36951a );
 a36956a <=( a36955a  and  a36948a );
 a36960a <=( (not A167)  and  A168 );
 a36961a <=( A169  and  a36960a );
 a36964a <=( A199  and  A166 );
 a36967a <=( A232  and  A200 );
 a36968a <=( a36967a  and  a36964a );
 a36969a <=( a36968a  and  a36961a );
 a36972a <=( A234  and  (not A233) );
 a36975a <=( (not A265)  and  A236 );
 a36976a <=( a36975a  and  a36972a );
 a36979a <=( (not A267)  and  A266 );
 a36982a <=( (not A269)  and  (not A268) );
 a36983a <=( a36982a  and  a36979a );
 a36984a <=( a36983a  and  a36976a );
 a36988a <=( (not A167)  and  A168 );
 a36989a <=( A169  and  a36988a );
 a36992a <=( A199  and  A166 );
 a36995a <=( A232  and  A200 );
 a36996a <=( a36995a  and  a36992a );
 a36997a <=( a36996a  and  a36989a );
 a37000a <=( A234  and  (not A233) );
 a37003a <=( A265  and  A236 );
 a37004a <=( a37003a  and  a37000a );
 a37007a <=( (not A267)  and  (not A266) );
 a37010a <=( (not A269)  and  (not A268) );
 a37011a <=( a37010a  and  a37007a );
 a37012a <=( a37011a  and  a37004a );
 a37016a <=( (not A167)  and  A168 );
 a37017a <=( A169  and  a37016a );
 a37020a <=( A199  and  A166 );
 a37023a <=( A232  and  A200 );
 a37024a <=( a37023a  and  a37020a );
 a37025a <=( a37024a  and  a37017a );
 a37028a <=( (not A234)  and  (not A233) );
 a37031a <=( (not A236)  and  (not A235) );
 a37032a <=( a37031a  and  a37028a );
 a37035a <=( (not A299)  and  A298 );
 a37038a <=( A301  and  A300 );
 a37039a <=( a37038a  and  a37035a );
 a37040a <=( a37039a  and  a37032a );
 a37044a <=( (not A167)  and  A168 );
 a37045a <=( A169  and  a37044a );
 a37048a <=( A199  and  A166 );
 a37051a <=( A232  and  A200 );
 a37052a <=( a37051a  and  a37048a );
 a37053a <=( a37052a  and  a37045a );
 a37056a <=( (not A234)  and  (not A233) );
 a37059a <=( (not A236)  and  (not A235) );
 a37060a <=( a37059a  and  a37056a );
 a37063a <=( (not A299)  and  A298 );
 a37066a <=( A302  and  A300 );
 a37067a <=( a37066a  and  a37063a );
 a37068a <=( a37067a  and  a37060a );
 a37072a <=( (not A167)  and  A168 );
 a37073a <=( A169  and  a37072a );
 a37076a <=( A199  and  A166 );
 a37079a <=( A232  and  A200 );
 a37080a <=( a37079a  and  a37076a );
 a37081a <=( a37080a  and  a37073a );
 a37084a <=( (not A234)  and  (not A233) );
 a37087a <=( (not A236)  and  (not A235) );
 a37088a <=( a37087a  and  a37084a );
 a37091a <=( A299  and  (not A298) );
 a37094a <=( A301  and  A300 );
 a37095a <=( a37094a  and  a37091a );
 a37096a <=( a37095a  and  a37088a );
 a37100a <=( (not A167)  and  A168 );
 a37101a <=( A169  and  a37100a );
 a37104a <=( A199  and  A166 );
 a37107a <=( A232  and  A200 );
 a37108a <=( a37107a  and  a37104a );
 a37109a <=( a37108a  and  a37101a );
 a37112a <=( (not A234)  and  (not A233) );
 a37115a <=( (not A236)  and  (not A235) );
 a37116a <=( a37115a  and  a37112a );
 a37119a <=( A299  and  (not A298) );
 a37122a <=( A302  and  A300 );
 a37123a <=( a37122a  and  a37119a );
 a37124a <=( a37123a  and  a37116a );
 a37128a <=( (not A167)  and  A168 );
 a37129a <=( A169  and  a37128a );
 a37132a <=( A199  and  A166 );
 a37135a <=( A232  and  A200 );
 a37136a <=( a37135a  and  a37132a );
 a37137a <=( a37136a  and  a37129a );
 a37140a <=( (not A234)  and  (not A233) );
 a37143a <=( (not A236)  and  (not A235) );
 a37144a <=( a37143a  and  a37140a );
 a37147a <=( A266  and  (not A265) );
 a37150a <=( A268  and  A267 );
 a37151a <=( a37150a  and  a37147a );
 a37152a <=( a37151a  and  a37144a );
 a37156a <=( (not A167)  and  A168 );
 a37157a <=( A169  and  a37156a );
 a37160a <=( A199  and  A166 );
 a37163a <=( A232  and  A200 );
 a37164a <=( a37163a  and  a37160a );
 a37165a <=( a37164a  and  a37157a );
 a37168a <=( (not A234)  and  (not A233) );
 a37171a <=( (not A236)  and  (not A235) );
 a37172a <=( a37171a  and  a37168a );
 a37175a <=( A266  and  (not A265) );
 a37178a <=( A269  and  A267 );
 a37179a <=( a37178a  and  a37175a );
 a37180a <=( a37179a  and  a37172a );
 a37184a <=( (not A167)  and  A168 );
 a37185a <=( A169  and  a37184a );
 a37188a <=( A199  and  A166 );
 a37191a <=( A232  and  A200 );
 a37192a <=( a37191a  and  a37188a );
 a37193a <=( a37192a  and  a37185a );
 a37196a <=( (not A234)  and  (not A233) );
 a37199a <=( (not A236)  and  (not A235) );
 a37200a <=( a37199a  and  a37196a );
 a37203a <=( (not A266)  and  A265 );
 a37206a <=( A268  and  A267 );
 a37207a <=( a37206a  and  a37203a );
 a37208a <=( a37207a  and  a37200a );
 a37212a <=( (not A167)  and  A168 );
 a37213a <=( A169  and  a37212a );
 a37216a <=( A199  and  A166 );
 a37219a <=( A232  and  A200 );
 a37220a <=( a37219a  and  a37216a );
 a37221a <=( a37220a  and  a37213a );
 a37224a <=( (not A234)  and  (not A233) );
 a37227a <=( (not A236)  and  (not A235) );
 a37228a <=( a37227a  and  a37224a );
 a37231a <=( (not A266)  and  A265 );
 a37234a <=( A269  and  A267 );
 a37235a <=( a37234a  and  a37231a );
 a37236a <=( a37235a  and  a37228a );
 a37240a <=( (not A167)  and  A168 );
 a37241a <=( A169  and  a37240a );
 a37244a <=( (not A199)  and  A166 );
 a37247a <=( (not A232)  and  (not A200) );
 a37248a <=( a37247a  and  a37244a );
 a37249a <=( a37248a  and  a37241a );
 a37252a <=( A234  and  A233 );
 a37255a <=( A298  and  A235 );
 a37256a <=( a37255a  and  a37252a );
 a37259a <=( (not A300)  and  (not A299) );
 a37262a <=( (not A302)  and  (not A301) );
 a37263a <=( a37262a  and  a37259a );
 a37264a <=( a37263a  and  a37256a );
 a37268a <=( (not A167)  and  A168 );
 a37269a <=( A169  and  a37268a );
 a37272a <=( (not A199)  and  A166 );
 a37275a <=( (not A232)  and  (not A200) );
 a37276a <=( a37275a  and  a37272a );
 a37277a <=( a37276a  and  a37269a );
 a37280a <=( A234  and  A233 );
 a37283a <=( (not A298)  and  A235 );
 a37284a <=( a37283a  and  a37280a );
 a37287a <=( (not A300)  and  A299 );
 a37290a <=( (not A302)  and  (not A301) );
 a37291a <=( a37290a  and  a37287a );
 a37292a <=( a37291a  and  a37284a );
 a37296a <=( (not A167)  and  A168 );
 a37297a <=( A169  and  a37296a );
 a37300a <=( (not A199)  and  A166 );
 a37303a <=( (not A232)  and  (not A200) );
 a37304a <=( a37303a  and  a37300a );
 a37305a <=( a37304a  and  a37297a );
 a37308a <=( A234  and  A233 );
 a37311a <=( (not A265)  and  A235 );
 a37312a <=( a37311a  and  a37308a );
 a37315a <=( (not A267)  and  A266 );
 a37318a <=( (not A269)  and  (not A268) );
 a37319a <=( a37318a  and  a37315a );
 a37320a <=( a37319a  and  a37312a );
 a37324a <=( (not A167)  and  A168 );
 a37325a <=( A169  and  a37324a );
 a37328a <=( (not A199)  and  A166 );
 a37331a <=( (not A232)  and  (not A200) );
 a37332a <=( a37331a  and  a37328a );
 a37333a <=( a37332a  and  a37325a );
 a37336a <=( A234  and  A233 );
 a37339a <=( A265  and  A235 );
 a37340a <=( a37339a  and  a37336a );
 a37343a <=( (not A267)  and  (not A266) );
 a37346a <=( (not A269)  and  (not A268) );
 a37347a <=( a37346a  and  a37343a );
 a37348a <=( a37347a  and  a37340a );
 a37352a <=( (not A167)  and  A168 );
 a37353a <=( A169  and  a37352a );
 a37356a <=( (not A199)  and  A166 );
 a37359a <=( (not A232)  and  (not A200) );
 a37360a <=( a37359a  and  a37356a );
 a37361a <=( a37360a  and  a37353a );
 a37364a <=( A234  and  A233 );
 a37367a <=( A298  and  A236 );
 a37368a <=( a37367a  and  a37364a );
 a37371a <=( (not A300)  and  (not A299) );
 a37374a <=( (not A302)  and  (not A301) );
 a37375a <=( a37374a  and  a37371a );
 a37376a <=( a37375a  and  a37368a );
 a37380a <=( (not A167)  and  A168 );
 a37381a <=( A169  and  a37380a );
 a37384a <=( (not A199)  and  A166 );
 a37387a <=( (not A232)  and  (not A200) );
 a37388a <=( a37387a  and  a37384a );
 a37389a <=( a37388a  and  a37381a );
 a37392a <=( A234  and  A233 );
 a37395a <=( (not A298)  and  A236 );
 a37396a <=( a37395a  and  a37392a );
 a37399a <=( (not A300)  and  A299 );
 a37402a <=( (not A302)  and  (not A301) );
 a37403a <=( a37402a  and  a37399a );
 a37404a <=( a37403a  and  a37396a );
 a37408a <=( (not A167)  and  A168 );
 a37409a <=( A169  and  a37408a );
 a37412a <=( (not A199)  and  A166 );
 a37415a <=( (not A232)  and  (not A200) );
 a37416a <=( a37415a  and  a37412a );
 a37417a <=( a37416a  and  a37409a );
 a37420a <=( A234  and  A233 );
 a37423a <=( (not A265)  and  A236 );
 a37424a <=( a37423a  and  a37420a );
 a37427a <=( (not A267)  and  A266 );
 a37430a <=( (not A269)  and  (not A268) );
 a37431a <=( a37430a  and  a37427a );
 a37432a <=( a37431a  and  a37424a );
 a37436a <=( (not A167)  and  A168 );
 a37437a <=( A169  and  a37436a );
 a37440a <=( (not A199)  and  A166 );
 a37443a <=( (not A232)  and  (not A200) );
 a37444a <=( a37443a  and  a37440a );
 a37445a <=( a37444a  and  a37437a );
 a37448a <=( A234  and  A233 );
 a37451a <=( A265  and  A236 );
 a37452a <=( a37451a  and  a37448a );
 a37455a <=( (not A267)  and  (not A266) );
 a37458a <=( (not A269)  and  (not A268) );
 a37459a <=( a37458a  and  a37455a );
 a37460a <=( a37459a  and  a37452a );
 a37464a <=( (not A167)  and  A168 );
 a37465a <=( A169  and  a37464a );
 a37468a <=( (not A199)  and  A166 );
 a37471a <=( (not A232)  and  (not A200) );
 a37472a <=( a37471a  and  a37468a );
 a37473a <=( a37472a  and  a37465a );
 a37476a <=( (not A234)  and  A233 );
 a37479a <=( (not A236)  and  (not A235) );
 a37480a <=( a37479a  and  a37476a );
 a37483a <=( (not A299)  and  A298 );
 a37486a <=( A301  and  A300 );
 a37487a <=( a37486a  and  a37483a );
 a37488a <=( a37487a  and  a37480a );
 a37492a <=( (not A167)  and  A168 );
 a37493a <=( A169  and  a37492a );
 a37496a <=( (not A199)  and  A166 );
 a37499a <=( (not A232)  and  (not A200) );
 a37500a <=( a37499a  and  a37496a );
 a37501a <=( a37500a  and  a37493a );
 a37504a <=( (not A234)  and  A233 );
 a37507a <=( (not A236)  and  (not A235) );
 a37508a <=( a37507a  and  a37504a );
 a37511a <=( (not A299)  and  A298 );
 a37514a <=( A302  and  A300 );
 a37515a <=( a37514a  and  a37511a );
 a37516a <=( a37515a  and  a37508a );
 a37520a <=( (not A167)  and  A168 );
 a37521a <=( A169  and  a37520a );
 a37524a <=( (not A199)  and  A166 );
 a37527a <=( (not A232)  and  (not A200) );
 a37528a <=( a37527a  and  a37524a );
 a37529a <=( a37528a  and  a37521a );
 a37532a <=( (not A234)  and  A233 );
 a37535a <=( (not A236)  and  (not A235) );
 a37536a <=( a37535a  and  a37532a );
 a37539a <=( A299  and  (not A298) );
 a37542a <=( A301  and  A300 );
 a37543a <=( a37542a  and  a37539a );
 a37544a <=( a37543a  and  a37536a );
 a37548a <=( (not A167)  and  A168 );
 a37549a <=( A169  and  a37548a );
 a37552a <=( (not A199)  and  A166 );
 a37555a <=( (not A232)  and  (not A200) );
 a37556a <=( a37555a  and  a37552a );
 a37557a <=( a37556a  and  a37549a );
 a37560a <=( (not A234)  and  A233 );
 a37563a <=( (not A236)  and  (not A235) );
 a37564a <=( a37563a  and  a37560a );
 a37567a <=( A299  and  (not A298) );
 a37570a <=( A302  and  A300 );
 a37571a <=( a37570a  and  a37567a );
 a37572a <=( a37571a  and  a37564a );
 a37576a <=( (not A167)  and  A168 );
 a37577a <=( A169  and  a37576a );
 a37580a <=( (not A199)  and  A166 );
 a37583a <=( (not A232)  and  (not A200) );
 a37584a <=( a37583a  and  a37580a );
 a37585a <=( a37584a  and  a37577a );
 a37588a <=( (not A234)  and  A233 );
 a37591a <=( (not A236)  and  (not A235) );
 a37592a <=( a37591a  and  a37588a );
 a37595a <=( A266  and  (not A265) );
 a37598a <=( A268  and  A267 );
 a37599a <=( a37598a  and  a37595a );
 a37600a <=( a37599a  and  a37592a );
 a37604a <=( (not A167)  and  A168 );
 a37605a <=( A169  and  a37604a );
 a37608a <=( (not A199)  and  A166 );
 a37611a <=( (not A232)  and  (not A200) );
 a37612a <=( a37611a  and  a37608a );
 a37613a <=( a37612a  and  a37605a );
 a37616a <=( (not A234)  and  A233 );
 a37619a <=( (not A236)  and  (not A235) );
 a37620a <=( a37619a  and  a37616a );
 a37623a <=( A266  and  (not A265) );
 a37626a <=( A269  and  A267 );
 a37627a <=( a37626a  and  a37623a );
 a37628a <=( a37627a  and  a37620a );
 a37632a <=( (not A167)  and  A168 );
 a37633a <=( A169  and  a37632a );
 a37636a <=( (not A199)  and  A166 );
 a37639a <=( (not A232)  and  (not A200) );
 a37640a <=( a37639a  and  a37636a );
 a37641a <=( a37640a  and  a37633a );
 a37644a <=( (not A234)  and  A233 );
 a37647a <=( (not A236)  and  (not A235) );
 a37648a <=( a37647a  and  a37644a );
 a37651a <=( (not A266)  and  A265 );
 a37654a <=( A268  and  A267 );
 a37655a <=( a37654a  and  a37651a );
 a37656a <=( a37655a  and  a37648a );
 a37660a <=( (not A167)  and  A168 );
 a37661a <=( A169  and  a37660a );
 a37664a <=( (not A199)  and  A166 );
 a37667a <=( (not A232)  and  (not A200) );
 a37668a <=( a37667a  and  a37664a );
 a37669a <=( a37668a  and  a37661a );
 a37672a <=( (not A234)  and  A233 );
 a37675a <=( (not A236)  and  (not A235) );
 a37676a <=( a37675a  and  a37672a );
 a37679a <=( (not A266)  and  A265 );
 a37682a <=( A269  and  A267 );
 a37683a <=( a37682a  and  a37679a );
 a37684a <=( a37683a  and  a37676a );
 a37688a <=( (not A167)  and  A168 );
 a37689a <=( A169  and  a37688a );
 a37692a <=( (not A199)  and  A166 );
 a37695a <=( A232  and  (not A200) );
 a37696a <=( a37695a  and  a37692a );
 a37697a <=( a37696a  and  a37689a );
 a37700a <=( A234  and  (not A233) );
 a37703a <=( A298  and  A235 );
 a37704a <=( a37703a  and  a37700a );
 a37707a <=( (not A300)  and  (not A299) );
 a37710a <=( (not A302)  and  (not A301) );
 a37711a <=( a37710a  and  a37707a );
 a37712a <=( a37711a  and  a37704a );
 a37716a <=( (not A167)  and  A168 );
 a37717a <=( A169  and  a37716a );
 a37720a <=( (not A199)  and  A166 );
 a37723a <=( A232  and  (not A200) );
 a37724a <=( a37723a  and  a37720a );
 a37725a <=( a37724a  and  a37717a );
 a37728a <=( A234  and  (not A233) );
 a37731a <=( (not A298)  and  A235 );
 a37732a <=( a37731a  and  a37728a );
 a37735a <=( (not A300)  and  A299 );
 a37738a <=( (not A302)  and  (not A301) );
 a37739a <=( a37738a  and  a37735a );
 a37740a <=( a37739a  and  a37732a );
 a37744a <=( (not A167)  and  A168 );
 a37745a <=( A169  and  a37744a );
 a37748a <=( (not A199)  and  A166 );
 a37751a <=( A232  and  (not A200) );
 a37752a <=( a37751a  and  a37748a );
 a37753a <=( a37752a  and  a37745a );
 a37756a <=( A234  and  (not A233) );
 a37759a <=( (not A265)  and  A235 );
 a37760a <=( a37759a  and  a37756a );
 a37763a <=( (not A267)  and  A266 );
 a37766a <=( (not A269)  and  (not A268) );
 a37767a <=( a37766a  and  a37763a );
 a37768a <=( a37767a  and  a37760a );
 a37772a <=( (not A167)  and  A168 );
 a37773a <=( A169  and  a37772a );
 a37776a <=( (not A199)  and  A166 );
 a37779a <=( A232  and  (not A200) );
 a37780a <=( a37779a  and  a37776a );
 a37781a <=( a37780a  and  a37773a );
 a37784a <=( A234  and  (not A233) );
 a37787a <=( A265  and  A235 );
 a37788a <=( a37787a  and  a37784a );
 a37791a <=( (not A267)  and  (not A266) );
 a37794a <=( (not A269)  and  (not A268) );
 a37795a <=( a37794a  and  a37791a );
 a37796a <=( a37795a  and  a37788a );
 a37800a <=( (not A167)  and  A168 );
 a37801a <=( A169  and  a37800a );
 a37804a <=( (not A199)  and  A166 );
 a37807a <=( A232  and  (not A200) );
 a37808a <=( a37807a  and  a37804a );
 a37809a <=( a37808a  and  a37801a );
 a37812a <=( A234  and  (not A233) );
 a37815a <=( A298  and  A236 );
 a37816a <=( a37815a  and  a37812a );
 a37819a <=( (not A300)  and  (not A299) );
 a37822a <=( (not A302)  and  (not A301) );
 a37823a <=( a37822a  and  a37819a );
 a37824a <=( a37823a  and  a37816a );
 a37828a <=( (not A167)  and  A168 );
 a37829a <=( A169  and  a37828a );
 a37832a <=( (not A199)  and  A166 );
 a37835a <=( A232  and  (not A200) );
 a37836a <=( a37835a  and  a37832a );
 a37837a <=( a37836a  and  a37829a );
 a37840a <=( A234  and  (not A233) );
 a37843a <=( (not A298)  and  A236 );
 a37844a <=( a37843a  and  a37840a );
 a37847a <=( (not A300)  and  A299 );
 a37850a <=( (not A302)  and  (not A301) );
 a37851a <=( a37850a  and  a37847a );
 a37852a <=( a37851a  and  a37844a );
 a37856a <=( (not A167)  and  A168 );
 a37857a <=( A169  and  a37856a );
 a37860a <=( (not A199)  and  A166 );
 a37863a <=( A232  and  (not A200) );
 a37864a <=( a37863a  and  a37860a );
 a37865a <=( a37864a  and  a37857a );
 a37868a <=( A234  and  (not A233) );
 a37871a <=( (not A265)  and  A236 );
 a37872a <=( a37871a  and  a37868a );
 a37875a <=( (not A267)  and  A266 );
 a37878a <=( (not A269)  and  (not A268) );
 a37879a <=( a37878a  and  a37875a );
 a37880a <=( a37879a  and  a37872a );
 a37884a <=( (not A167)  and  A168 );
 a37885a <=( A169  and  a37884a );
 a37888a <=( (not A199)  and  A166 );
 a37891a <=( A232  and  (not A200) );
 a37892a <=( a37891a  and  a37888a );
 a37893a <=( a37892a  and  a37885a );
 a37896a <=( A234  and  (not A233) );
 a37899a <=( A265  and  A236 );
 a37900a <=( a37899a  and  a37896a );
 a37903a <=( (not A267)  and  (not A266) );
 a37906a <=( (not A269)  and  (not A268) );
 a37907a <=( a37906a  and  a37903a );
 a37908a <=( a37907a  and  a37900a );
 a37912a <=( (not A167)  and  A168 );
 a37913a <=( A169  and  a37912a );
 a37916a <=( (not A199)  and  A166 );
 a37919a <=( A232  and  (not A200) );
 a37920a <=( a37919a  and  a37916a );
 a37921a <=( a37920a  and  a37913a );
 a37924a <=( (not A234)  and  (not A233) );
 a37927a <=( (not A236)  and  (not A235) );
 a37928a <=( a37927a  and  a37924a );
 a37931a <=( (not A299)  and  A298 );
 a37934a <=( A301  and  A300 );
 a37935a <=( a37934a  and  a37931a );
 a37936a <=( a37935a  and  a37928a );
 a37940a <=( (not A167)  and  A168 );
 a37941a <=( A169  and  a37940a );
 a37944a <=( (not A199)  and  A166 );
 a37947a <=( A232  and  (not A200) );
 a37948a <=( a37947a  and  a37944a );
 a37949a <=( a37948a  and  a37941a );
 a37952a <=( (not A234)  and  (not A233) );
 a37955a <=( (not A236)  and  (not A235) );
 a37956a <=( a37955a  and  a37952a );
 a37959a <=( (not A299)  and  A298 );
 a37962a <=( A302  and  A300 );
 a37963a <=( a37962a  and  a37959a );
 a37964a <=( a37963a  and  a37956a );
 a37968a <=( (not A167)  and  A168 );
 a37969a <=( A169  and  a37968a );
 a37972a <=( (not A199)  and  A166 );
 a37975a <=( A232  and  (not A200) );
 a37976a <=( a37975a  and  a37972a );
 a37977a <=( a37976a  and  a37969a );
 a37980a <=( (not A234)  and  (not A233) );
 a37983a <=( (not A236)  and  (not A235) );
 a37984a <=( a37983a  and  a37980a );
 a37987a <=( A299  and  (not A298) );
 a37990a <=( A301  and  A300 );
 a37991a <=( a37990a  and  a37987a );
 a37992a <=( a37991a  and  a37984a );
 a37996a <=( (not A167)  and  A168 );
 a37997a <=( A169  and  a37996a );
 a38000a <=( (not A199)  and  A166 );
 a38003a <=( A232  and  (not A200) );
 a38004a <=( a38003a  and  a38000a );
 a38005a <=( a38004a  and  a37997a );
 a38008a <=( (not A234)  and  (not A233) );
 a38011a <=( (not A236)  and  (not A235) );
 a38012a <=( a38011a  and  a38008a );
 a38015a <=( A299  and  (not A298) );
 a38018a <=( A302  and  A300 );
 a38019a <=( a38018a  and  a38015a );
 a38020a <=( a38019a  and  a38012a );
 a38024a <=( (not A167)  and  A168 );
 a38025a <=( A169  and  a38024a );
 a38028a <=( (not A199)  and  A166 );
 a38031a <=( A232  and  (not A200) );
 a38032a <=( a38031a  and  a38028a );
 a38033a <=( a38032a  and  a38025a );
 a38036a <=( (not A234)  and  (not A233) );
 a38039a <=( (not A236)  and  (not A235) );
 a38040a <=( a38039a  and  a38036a );
 a38043a <=( A266  and  (not A265) );
 a38046a <=( A268  and  A267 );
 a38047a <=( a38046a  and  a38043a );
 a38048a <=( a38047a  and  a38040a );
 a38052a <=( (not A167)  and  A168 );
 a38053a <=( A169  and  a38052a );
 a38056a <=( (not A199)  and  A166 );
 a38059a <=( A232  and  (not A200) );
 a38060a <=( a38059a  and  a38056a );
 a38061a <=( a38060a  and  a38053a );
 a38064a <=( (not A234)  and  (not A233) );
 a38067a <=( (not A236)  and  (not A235) );
 a38068a <=( a38067a  and  a38064a );
 a38071a <=( A266  and  (not A265) );
 a38074a <=( A269  and  A267 );
 a38075a <=( a38074a  and  a38071a );
 a38076a <=( a38075a  and  a38068a );
 a38080a <=( (not A167)  and  A168 );
 a38081a <=( A169  and  a38080a );
 a38084a <=( (not A199)  and  A166 );
 a38087a <=( A232  and  (not A200) );
 a38088a <=( a38087a  and  a38084a );
 a38089a <=( a38088a  and  a38081a );
 a38092a <=( (not A234)  and  (not A233) );
 a38095a <=( (not A236)  and  (not A235) );
 a38096a <=( a38095a  and  a38092a );
 a38099a <=( (not A266)  and  A265 );
 a38102a <=( A268  and  A267 );
 a38103a <=( a38102a  and  a38099a );
 a38104a <=( a38103a  and  a38096a );
 a38108a <=( (not A167)  and  A168 );
 a38109a <=( A169  and  a38108a );
 a38112a <=( (not A199)  and  A166 );
 a38115a <=( A232  and  (not A200) );
 a38116a <=( a38115a  and  a38112a );
 a38117a <=( a38116a  and  a38109a );
 a38120a <=( (not A234)  and  (not A233) );
 a38123a <=( (not A236)  and  (not A235) );
 a38124a <=( a38123a  and  a38120a );
 a38127a <=( (not A266)  and  A265 );
 a38130a <=( A269  and  A267 );
 a38131a <=( a38130a  and  a38127a );
 a38132a <=( a38131a  and  a38124a );
 a38136a <=( (not A168)  and  (not A169) );
 a38137a <=( A170  and  a38136a );
 a38140a <=( (not A166)  and  A167 );
 a38143a <=( A202  and  (not A201) );
 a38144a <=( a38143a  and  a38140a );
 a38145a <=( a38144a  and  a38137a );
 a38148a <=( A233  and  (not A232) );
 a38151a <=( A235  and  A234 );
 a38152a <=( a38151a  and  a38148a );
 a38155a <=( (not A299)  and  A298 );
 a38158a <=( A301  and  A300 );
 a38159a <=( a38158a  and  a38155a );
 a38160a <=( a38159a  and  a38152a );
 a38164a <=( (not A168)  and  (not A169) );
 a38165a <=( A170  and  a38164a );
 a38168a <=( (not A166)  and  A167 );
 a38171a <=( A202  and  (not A201) );
 a38172a <=( a38171a  and  a38168a );
 a38173a <=( a38172a  and  a38165a );
 a38176a <=( A233  and  (not A232) );
 a38179a <=( A235  and  A234 );
 a38180a <=( a38179a  and  a38176a );
 a38183a <=( (not A299)  and  A298 );
 a38186a <=( A302  and  A300 );
 a38187a <=( a38186a  and  a38183a );
 a38188a <=( a38187a  and  a38180a );
 a38192a <=( (not A168)  and  (not A169) );
 a38193a <=( A170  and  a38192a );
 a38196a <=( (not A166)  and  A167 );
 a38199a <=( A202  and  (not A201) );
 a38200a <=( a38199a  and  a38196a );
 a38201a <=( a38200a  and  a38193a );
 a38204a <=( A233  and  (not A232) );
 a38207a <=( A235  and  A234 );
 a38208a <=( a38207a  and  a38204a );
 a38211a <=( A299  and  (not A298) );
 a38214a <=( A301  and  A300 );
 a38215a <=( a38214a  and  a38211a );
 a38216a <=( a38215a  and  a38208a );
 a38220a <=( (not A168)  and  (not A169) );
 a38221a <=( A170  and  a38220a );
 a38224a <=( (not A166)  and  A167 );
 a38227a <=( A202  and  (not A201) );
 a38228a <=( a38227a  and  a38224a );
 a38229a <=( a38228a  and  a38221a );
 a38232a <=( A233  and  (not A232) );
 a38235a <=( A235  and  A234 );
 a38236a <=( a38235a  and  a38232a );
 a38239a <=( A299  and  (not A298) );
 a38242a <=( A302  and  A300 );
 a38243a <=( a38242a  and  a38239a );
 a38244a <=( a38243a  and  a38236a );
 a38248a <=( (not A168)  and  (not A169) );
 a38249a <=( A170  and  a38248a );
 a38252a <=( (not A166)  and  A167 );
 a38255a <=( A202  and  (not A201) );
 a38256a <=( a38255a  and  a38252a );
 a38257a <=( a38256a  and  a38249a );
 a38260a <=( A233  and  (not A232) );
 a38263a <=( A235  and  A234 );
 a38264a <=( a38263a  and  a38260a );
 a38267a <=( A266  and  (not A265) );
 a38270a <=( A268  and  A267 );
 a38271a <=( a38270a  and  a38267a );
 a38272a <=( a38271a  and  a38264a );
 a38276a <=( (not A168)  and  (not A169) );
 a38277a <=( A170  and  a38276a );
 a38280a <=( (not A166)  and  A167 );
 a38283a <=( A202  and  (not A201) );
 a38284a <=( a38283a  and  a38280a );
 a38285a <=( a38284a  and  a38277a );
 a38288a <=( A233  and  (not A232) );
 a38291a <=( A235  and  A234 );
 a38292a <=( a38291a  and  a38288a );
 a38295a <=( A266  and  (not A265) );
 a38298a <=( A269  and  A267 );
 a38299a <=( a38298a  and  a38295a );
 a38300a <=( a38299a  and  a38292a );
 a38304a <=( (not A168)  and  (not A169) );
 a38305a <=( A170  and  a38304a );
 a38308a <=( (not A166)  and  A167 );
 a38311a <=( A202  and  (not A201) );
 a38312a <=( a38311a  and  a38308a );
 a38313a <=( a38312a  and  a38305a );
 a38316a <=( A233  and  (not A232) );
 a38319a <=( A235  and  A234 );
 a38320a <=( a38319a  and  a38316a );
 a38323a <=( (not A266)  and  A265 );
 a38326a <=( A268  and  A267 );
 a38327a <=( a38326a  and  a38323a );
 a38328a <=( a38327a  and  a38320a );
 a38332a <=( (not A168)  and  (not A169) );
 a38333a <=( A170  and  a38332a );
 a38336a <=( (not A166)  and  A167 );
 a38339a <=( A202  and  (not A201) );
 a38340a <=( a38339a  and  a38336a );
 a38341a <=( a38340a  and  a38333a );
 a38344a <=( A233  and  (not A232) );
 a38347a <=( A235  and  A234 );
 a38348a <=( a38347a  and  a38344a );
 a38351a <=( (not A266)  and  A265 );
 a38354a <=( A269  and  A267 );
 a38355a <=( a38354a  and  a38351a );
 a38356a <=( a38355a  and  a38348a );
 a38360a <=( (not A168)  and  (not A169) );
 a38361a <=( A170  and  a38360a );
 a38364a <=( (not A166)  and  A167 );
 a38367a <=( A202  and  (not A201) );
 a38368a <=( a38367a  and  a38364a );
 a38369a <=( a38368a  and  a38361a );
 a38372a <=( A233  and  (not A232) );
 a38375a <=( A236  and  A234 );
 a38376a <=( a38375a  and  a38372a );
 a38379a <=( (not A299)  and  A298 );
 a38382a <=( A301  and  A300 );
 a38383a <=( a38382a  and  a38379a );
 a38384a <=( a38383a  and  a38376a );
 a38388a <=( (not A168)  and  (not A169) );
 a38389a <=( A170  and  a38388a );
 a38392a <=( (not A166)  and  A167 );
 a38395a <=( A202  and  (not A201) );
 a38396a <=( a38395a  and  a38392a );
 a38397a <=( a38396a  and  a38389a );
 a38400a <=( A233  and  (not A232) );
 a38403a <=( A236  and  A234 );
 a38404a <=( a38403a  and  a38400a );
 a38407a <=( (not A299)  and  A298 );
 a38410a <=( A302  and  A300 );
 a38411a <=( a38410a  and  a38407a );
 a38412a <=( a38411a  and  a38404a );
 a38416a <=( (not A168)  and  (not A169) );
 a38417a <=( A170  and  a38416a );
 a38420a <=( (not A166)  and  A167 );
 a38423a <=( A202  and  (not A201) );
 a38424a <=( a38423a  and  a38420a );
 a38425a <=( a38424a  and  a38417a );
 a38428a <=( A233  and  (not A232) );
 a38431a <=( A236  and  A234 );
 a38432a <=( a38431a  and  a38428a );
 a38435a <=( A299  and  (not A298) );
 a38438a <=( A301  and  A300 );
 a38439a <=( a38438a  and  a38435a );
 a38440a <=( a38439a  and  a38432a );
 a38444a <=( (not A168)  and  (not A169) );
 a38445a <=( A170  and  a38444a );
 a38448a <=( (not A166)  and  A167 );
 a38451a <=( A202  and  (not A201) );
 a38452a <=( a38451a  and  a38448a );
 a38453a <=( a38452a  and  a38445a );
 a38456a <=( A233  and  (not A232) );
 a38459a <=( A236  and  A234 );
 a38460a <=( a38459a  and  a38456a );
 a38463a <=( A299  and  (not A298) );
 a38466a <=( A302  and  A300 );
 a38467a <=( a38466a  and  a38463a );
 a38468a <=( a38467a  and  a38460a );
 a38472a <=( (not A168)  and  (not A169) );
 a38473a <=( A170  and  a38472a );
 a38476a <=( (not A166)  and  A167 );
 a38479a <=( A202  and  (not A201) );
 a38480a <=( a38479a  and  a38476a );
 a38481a <=( a38480a  and  a38473a );
 a38484a <=( A233  and  (not A232) );
 a38487a <=( A236  and  A234 );
 a38488a <=( a38487a  and  a38484a );
 a38491a <=( A266  and  (not A265) );
 a38494a <=( A268  and  A267 );
 a38495a <=( a38494a  and  a38491a );
 a38496a <=( a38495a  and  a38488a );
 a38500a <=( (not A168)  and  (not A169) );
 a38501a <=( A170  and  a38500a );
 a38504a <=( (not A166)  and  A167 );
 a38507a <=( A202  and  (not A201) );
 a38508a <=( a38507a  and  a38504a );
 a38509a <=( a38508a  and  a38501a );
 a38512a <=( A233  and  (not A232) );
 a38515a <=( A236  and  A234 );
 a38516a <=( a38515a  and  a38512a );
 a38519a <=( A266  and  (not A265) );
 a38522a <=( A269  and  A267 );
 a38523a <=( a38522a  and  a38519a );
 a38524a <=( a38523a  and  a38516a );
 a38528a <=( (not A168)  and  (not A169) );
 a38529a <=( A170  and  a38528a );
 a38532a <=( (not A166)  and  A167 );
 a38535a <=( A202  and  (not A201) );
 a38536a <=( a38535a  and  a38532a );
 a38537a <=( a38536a  and  a38529a );
 a38540a <=( A233  and  (not A232) );
 a38543a <=( A236  and  A234 );
 a38544a <=( a38543a  and  a38540a );
 a38547a <=( (not A266)  and  A265 );
 a38550a <=( A268  and  A267 );
 a38551a <=( a38550a  and  a38547a );
 a38552a <=( a38551a  and  a38544a );
 a38556a <=( (not A168)  and  (not A169) );
 a38557a <=( A170  and  a38556a );
 a38560a <=( (not A166)  and  A167 );
 a38563a <=( A202  and  (not A201) );
 a38564a <=( a38563a  and  a38560a );
 a38565a <=( a38564a  and  a38557a );
 a38568a <=( A233  and  (not A232) );
 a38571a <=( A236  and  A234 );
 a38572a <=( a38571a  and  a38568a );
 a38575a <=( (not A266)  and  A265 );
 a38578a <=( A269  and  A267 );
 a38579a <=( a38578a  and  a38575a );
 a38580a <=( a38579a  and  a38572a );
 a38584a <=( (not A168)  and  (not A169) );
 a38585a <=( A170  and  a38584a );
 a38588a <=( (not A166)  and  A167 );
 a38591a <=( A202  and  (not A201) );
 a38592a <=( a38591a  and  a38588a );
 a38593a <=( a38592a  and  a38585a );
 a38596a <=( (not A233)  and  A232 );
 a38599a <=( A235  and  A234 );
 a38600a <=( a38599a  and  a38596a );
 a38603a <=( (not A299)  and  A298 );
 a38606a <=( A301  and  A300 );
 a38607a <=( a38606a  and  a38603a );
 a38608a <=( a38607a  and  a38600a );
 a38612a <=( (not A168)  and  (not A169) );
 a38613a <=( A170  and  a38612a );
 a38616a <=( (not A166)  and  A167 );
 a38619a <=( A202  and  (not A201) );
 a38620a <=( a38619a  and  a38616a );
 a38621a <=( a38620a  and  a38613a );
 a38624a <=( (not A233)  and  A232 );
 a38627a <=( A235  and  A234 );
 a38628a <=( a38627a  and  a38624a );
 a38631a <=( (not A299)  and  A298 );
 a38634a <=( A302  and  A300 );
 a38635a <=( a38634a  and  a38631a );
 a38636a <=( a38635a  and  a38628a );
 a38640a <=( (not A168)  and  (not A169) );
 a38641a <=( A170  and  a38640a );
 a38644a <=( (not A166)  and  A167 );
 a38647a <=( A202  and  (not A201) );
 a38648a <=( a38647a  and  a38644a );
 a38649a <=( a38648a  and  a38641a );
 a38652a <=( (not A233)  and  A232 );
 a38655a <=( A235  and  A234 );
 a38656a <=( a38655a  and  a38652a );
 a38659a <=( A299  and  (not A298) );
 a38662a <=( A301  and  A300 );
 a38663a <=( a38662a  and  a38659a );
 a38664a <=( a38663a  and  a38656a );
 a38668a <=( (not A168)  and  (not A169) );
 a38669a <=( A170  and  a38668a );
 a38672a <=( (not A166)  and  A167 );
 a38675a <=( A202  and  (not A201) );
 a38676a <=( a38675a  and  a38672a );
 a38677a <=( a38676a  and  a38669a );
 a38680a <=( (not A233)  and  A232 );
 a38683a <=( A235  and  A234 );
 a38684a <=( a38683a  and  a38680a );
 a38687a <=( A299  and  (not A298) );
 a38690a <=( A302  and  A300 );
 a38691a <=( a38690a  and  a38687a );
 a38692a <=( a38691a  and  a38684a );
 a38696a <=( (not A168)  and  (not A169) );
 a38697a <=( A170  and  a38696a );
 a38700a <=( (not A166)  and  A167 );
 a38703a <=( A202  and  (not A201) );
 a38704a <=( a38703a  and  a38700a );
 a38705a <=( a38704a  and  a38697a );
 a38708a <=( (not A233)  and  A232 );
 a38711a <=( A235  and  A234 );
 a38712a <=( a38711a  and  a38708a );
 a38715a <=( A266  and  (not A265) );
 a38718a <=( A268  and  A267 );
 a38719a <=( a38718a  and  a38715a );
 a38720a <=( a38719a  and  a38712a );
 a38724a <=( (not A168)  and  (not A169) );
 a38725a <=( A170  and  a38724a );
 a38728a <=( (not A166)  and  A167 );
 a38731a <=( A202  and  (not A201) );
 a38732a <=( a38731a  and  a38728a );
 a38733a <=( a38732a  and  a38725a );
 a38736a <=( (not A233)  and  A232 );
 a38739a <=( A235  and  A234 );
 a38740a <=( a38739a  and  a38736a );
 a38743a <=( A266  and  (not A265) );
 a38746a <=( A269  and  A267 );
 a38747a <=( a38746a  and  a38743a );
 a38748a <=( a38747a  and  a38740a );
 a38752a <=( (not A168)  and  (not A169) );
 a38753a <=( A170  and  a38752a );
 a38756a <=( (not A166)  and  A167 );
 a38759a <=( A202  and  (not A201) );
 a38760a <=( a38759a  and  a38756a );
 a38761a <=( a38760a  and  a38753a );
 a38764a <=( (not A233)  and  A232 );
 a38767a <=( A235  and  A234 );
 a38768a <=( a38767a  and  a38764a );
 a38771a <=( (not A266)  and  A265 );
 a38774a <=( A268  and  A267 );
 a38775a <=( a38774a  and  a38771a );
 a38776a <=( a38775a  and  a38768a );
 a38780a <=( (not A168)  and  (not A169) );
 a38781a <=( A170  and  a38780a );
 a38784a <=( (not A166)  and  A167 );
 a38787a <=( A202  and  (not A201) );
 a38788a <=( a38787a  and  a38784a );
 a38789a <=( a38788a  and  a38781a );
 a38792a <=( (not A233)  and  A232 );
 a38795a <=( A235  and  A234 );
 a38796a <=( a38795a  and  a38792a );
 a38799a <=( (not A266)  and  A265 );
 a38802a <=( A269  and  A267 );
 a38803a <=( a38802a  and  a38799a );
 a38804a <=( a38803a  and  a38796a );
 a38808a <=( (not A168)  and  (not A169) );
 a38809a <=( A170  and  a38808a );
 a38812a <=( (not A166)  and  A167 );
 a38815a <=( A202  and  (not A201) );
 a38816a <=( a38815a  and  a38812a );
 a38817a <=( a38816a  and  a38809a );
 a38820a <=( (not A233)  and  A232 );
 a38823a <=( A236  and  A234 );
 a38824a <=( a38823a  and  a38820a );
 a38827a <=( (not A299)  and  A298 );
 a38830a <=( A301  and  A300 );
 a38831a <=( a38830a  and  a38827a );
 a38832a <=( a38831a  and  a38824a );
 a38836a <=( (not A168)  and  (not A169) );
 a38837a <=( A170  and  a38836a );
 a38840a <=( (not A166)  and  A167 );
 a38843a <=( A202  and  (not A201) );
 a38844a <=( a38843a  and  a38840a );
 a38845a <=( a38844a  and  a38837a );
 a38848a <=( (not A233)  and  A232 );
 a38851a <=( A236  and  A234 );
 a38852a <=( a38851a  and  a38848a );
 a38855a <=( (not A299)  and  A298 );
 a38858a <=( A302  and  A300 );
 a38859a <=( a38858a  and  a38855a );
 a38860a <=( a38859a  and  a38852a );
 a38864a <=( (not A168)  and  (not A169) );
 a38865a <=( A170  and  a38864a );
 a38868a <=( (not A166)  and  A167 );
 a38871a <=( A202  and  (not A201) );
 a38872a <=( a38871a  and  a38868a );
 a38873a <=( a38872a  and  a38865a );
 a38876a <=( (not A233)  and  A232 );
 a38879a <=( A236  and  A234 );
 a38880a <=( a38879a  and  a38876a );
 a38883a <=( A299  and  (not A298) );
 a38886a <=( A301  and  A300 );
 a38887a <=( a38886a  and  a38883a );
 a38888a <=( a38887a  and  a38880a );
 a38892a <=( (not A168)  and  (not A169) );
 a38893a <=( A170  and  a38892a );
 a38896a <=( (not A166)  and  A167 );
 a38899a <=( A202  and  (not A201) );
 a38900a <=( a38899a  and  a38896a );
 a38901a <=( a38900a  and  a38893a );
 a38904a <=( (not A233)  and  A232 );
 a38907a <=( A236  and  A234 );
 a38908a <=( a38907a  and  a38904a );
 a38911a <=( A299  and  (not A298) );
 a38914a <=( A302  and  A300 );
 a38915a <=( a38914a  and  a38911a );
 a38916a <=( a38915a  and  a38908a );
 a38920a <=( (not A168)  and  (not A169) );
 a38921a <=( A170  and  a38920a );
 a38924a <=( (not A166)  and  A167 );
 a38927a <=( A202  and  (not A201) );
 a38928a <=( a38927a  and  a38924a );
 a38929a <=( a38928a  and  a38921a );
 a38932a <=( (not A233)  and  A232 );
 a38935a <=( A236  and  A234 );
 a38936a <=( a38935a  and  a38932a );
 a38939a <=( A266  and  (not A265) );
 a38942a <=( A268  and  A267 );
 a38943a <=( a38942a  and  a38939a );
 a38944a <=( a38943a  and  a38936a );
 a38948a <=( (not A168)  and  (not A169) );
 a38949a <=( A170  and  a38948a );
 a38952a <=( (not A166)  and  A167 );
 a38955a <=( A202  and  (not A201) );
 a38956a <=( a38955a  and  a38952a );
 a38957a <=( a38956a  and  a38949a );
 a38960a <=( (not A233)  and  A232 );
 a38963a <=( A236  and  A234 );
 a38964a <=( a38963a  and  a38960a );
 a38967a <=( A266  and  (not A265) );
 a38970a <=( A269  and  A267 );
 a38971a <=( a38970a  and  a38967a );
 a38972a <=( a38971a  and  a38964a );
 a38976a <=( (not A168)  and  (not A169) );
 a38977a <=( A170  and  a38976a );
 a38980a <=( (not A166)  and  A167 );
 a38983a <=( A202  and  (not A201) );
 a38984a <=( a38983a  and  a38980a );
 a38985a <=( a38984a  and  a38977a );
 a38988a <=( (not A233)  and  A232 );
 a38991a <=( A236  and  A234 );
 a38992a <=( a38991a  and  a38988a );
 a38995a <=( (not A266)  and  A265 );
 a38998a <=( A268  and  A267 );
 a38999a <=( a38998a  and  a38995a );
 a39000a <=( a38999a  and  a38992a );
 a39004a <=( (not A168)  and  (not A169) );
 a39005a <=( A170  and  a39004a );
 a39008a <=( (not A166)  and  A167 );
 a39011a <=( A202  and  (not A201) );
 a39012a <=( a39011a  and  a39008a );
 a39013a <=( a39012a  and  a39005a );
 a39016a <=( (not A233)  and  A232 );
 a39019a <=( A236  and  A234 );
 a39020a <=( a39019a  and  a39016a );
 a39023a <=( (not A266)  and  A265 );
 a39026a <=( A269  and  A267 );
 a39027a <=( a39026a  and  a39023a );
 a39028a <=( a39027a  and  a39020a );
 a39032a <=( (not A168)  and  (not A169) );
 a39033a <=( A170  and  a39032a );
 a39036a <=( (not A166)  and  A167 );
 a39039a <=( A203  and  (not A201) );
 a39040a <=( a39039a  and  a39036a );
 a39041a <=( a39040a  and  a39033a );
 a39044a <=( A233  and  (not A232) );
 a39047a <=( A235  and  A234 );
 a39048a <=( a39047a  and  a39044a );
 a39051a <=( (not A299)  and  A298 );
 a39054a <=( A301  and  A300 );
 a39055a <=( a39054a  and  a39051a );
 a39056a <=( a39055a  and  a39048a );
 a39060a <=( (not A168)  and  (not A169) );
 a39061a <=( A170  and  a39060a );
 a39064a <=( (not A166)  and  A167 );
 a39067a <=( A203  and  (not A201) );
 a39068a <=( a39067a  and  a39064a );
 a39069a <=( a39068a  and  a39061a );
 a39072a <=( A233  and  (not A232) );
 a39075a <=( A235  and  A234 );
 a39076a <=( a39075a  and  a39072a );
 a39079a <=( (not A299)  and  A298 );
 a39082a <=( A302  and  A300 );
 a39083a <=( a39082a  and  a39079a );
 a39084a <=( a39083a  and  a39076a );
 a39088a <=( (not A168)  and  (not A169) );
 a39089a <=( A170  and  a39088a );
 a39092a <=( (not A166)  and  A167 );
 a39095a <=( A203  and  (not A201) );
 a39096a <=( a39095a  and  a39092a );
 a39097a <=( a39096a  and  a39089a );
 a39100a <=( A233  and  (not A232) );
 a39103a <=( A235  and  A234 );
 a39104a <=( a39103a  and  a39100a );
 a39107a <=( A299  and  (not A298) );
 a39110a <=( A301  and  A300 );
 a39111a <=( a39110a  and  a39107a );
 a39112a <=( a39111a  and  a39104a );
 a39116a <=( (not A168)  and  (not A169) );
 a39117a <=( A170  and  a39116a );
 a39120a <=( (not A166)  and  A167 );
 a39123a <=( A203  and  (not A201) );
 a39124a <=( a39123a  and  a39120a );
 a39125a <=( a39124a  and  a39117a );
 a39128a <=( A233  and  (not A232) );
 a39131a <=( A235  and  A234 );
 a39132a <=( a39131a  and  a39128a );
 a39135a <=( A299  and  (not A298) );
 a39138a <=( A302  and  A300 );
 a39139a <=( a39138a  and  a39135a );
 a39140a <=( a39139a  and  a39132a );
 a39144a <=( (not A168)  and  (not A169) );
 a39145a <=( A170  and  a39144a );
 a39148a <=( (not A166)  and  A167 );
 a39151a <=( A203  and  (not A201) );
 a39152a <=( a39151a  and  a39148a );
 a39153a <=( a39152a  and  a39145a );
 a39156a <=( A233  and  (not A232) );
 a39159a <=( A235  and  A234 );
 a39160a <=( a39159a  and  a39156a );
 a39163a <=( A266  and  (not A265) );
 a39166a <=( A268  and  A267 );
 a39167a <=( a39166a  and  a39163a );
 a39168a <=( a39167a  and  a39160a );
 a39172a <=( (not A168)  and  (not A169) );
 a39173a <=( A170  and  a39172a );
 a39176a <=( (not A166)  and  A167 );
 a39179a <=( A203  and  (not A201) );
 a39180a <=( a39179a  and  a39176a );
 a39181a <=( a39180a  and  a39173a );
 a39184a <=( A233  and  (not A232) );
 a39187a <=( A235  and  A234 );
 a39188a <=( a39187a  and  a39184a );
 a39191a <=( A266  and  (not A265) );
 a39194a <=( A269  and  A267 );
 a39195a <=( a39194a  and  a39191a );
 a39196a <=( a39195a  and  a39188a );
 a39200a <=( (not A168)  and  (not A169) );
 a39201a <=( A170  and  a39200a );
 a39204a <=( (not A166)  and  A167 );
 a39207a <=( A203  and  (not A201) );
 a39208a <=( a39207a  and  a39204a );
 a39209a <=( a39208a  and  a39201a );
 a39212a <=( A233  and  (not A232) );
 a39215a <=( A235  and  A234 );
 a39216a <=( a39215a  and  a39212a );
 a39219a <=( (not A266)  and  A265 );
 a39222a <=( A268  and  A267 );
 a39223a <=( a39222a  and  a39219a );
 a39224a <=( a39223a  and  a39216a );
 a39228a <=( (not A168)  and  (not A169) );
 a39229a <=( A170  and  a39228a );
 a39232a <=( (not A166)  and  A167 );
 a39235a <=( A203  and  (not A201) );
 a39236a <=( a39235a  and  a39232a );
 a39237a <=( a39236a  and  a39229a );
 a39240a <=( A233  and  (not A232) );
 a39243a <=( A235  and  A234 );
 a39244a <=( a39243a  and  a39240a );
 a39247a <=( (not A266)  and  A265 );
 a39250a <=( A269  and  A267 );
 a39251a <=( a39250a  and  a39247a );
 a39252a <=( a39251a  and  a39244a );
 a39256a <=( (not A168)  and  (not A169) );
 a39257a <=( A170  and  a39256a );
 a39260a <=( (not A166)  and  A167 );
 a39263a <=( A203  and  (not A201) );
 a39264a <=( a39263a  and  a39260a );
 a39265a <=( a39264a  and  a39257a );
 a39268a <=( A233  and  (not A232) );
 a39271a <=( A236  and  A234 );
 a39272a <=( a39271a  and  a39268a );
 a39275a <=( (not A299)  and  A298 );
 a39278a <=( A301  and  A300 );
 a39279a <=( a39278a  and  a39275a );
 a39280a <=( a39279a  and  a39272a );
 a39284a <=( (not A168)  and  (not A169) );
 a39285a <=( A170  and  a39284a );
 a39288a <=( (not A166)  and  A167 );
 a39291a <=( A203  and  (not A201) );
 a39292a <=( a39291a  and  a39288a );
 a39293a <=( a39292a  and  a39285a );
 a39296a <=( A233  and  (not A232) );
 a39299a <=( A236  and  A234 );
 a39300a <=( a39299a  and  a39296a );
 a39303a <=( (not A299)  and  A298 );
 a39306a <=( A302  and  A300 );
 a39307a <=( a39306a  and  a39303a );
 a39308a <=( a39307a  and  a39300a );
 a39312a <=( (not A168)  and  (not A169) );
 a39313a <=( A170  and  a39312a );
 a39316a <=( (not A166)  and  A167 );
 a39319a <=( A203  and  (not A201) );
 a39320a <=( a39319a  and  a39316a );
 a39321a <=( a39320a  and  a39313a );
 a39324a <=( A233  and  (not A232) );
 a39327a <=( A236  and  A234 );
 a39328a <=( a39327a  and  a39324a );
 a39331a <=( A299  and  (not A298) );
 a39334a <=( A301  and  A300 );
 a39335a <=( a39334a  and  a39331a );
 a39336a <=( a39335a  and  a39328a );
 a39340a <=( (not A168)  and  (not A169) );
 a39341a <=( A170  and  a39340a );
 a39344a <=( (not A166)  and  A167 );
 a39347a <=( A203  and  (not A201) );
 a39348a <=( a39347a  and  a39344a );
 a39349a <=( a39348a  and  a39341a );
 a39352a <=( A233  and  (not A232) );
 a39355a <=( A236  and  A234 );
 a39356a <=( a39355a  and  a39352a );
 a39359a <=( A299  and  (not A298) );
 a39362a <=( A302  and  A300 );
 a39363a <=( a39362a  and  a39359a );
 a39364a <=( a39363a  and  a39356a );
 a39368a <=( (not A168)  and  (not A169) );
 a39369a <=( A170  and  a39368a );
 a39372a <=( (not A166)  and  A167 );
 a39375a <=( A203  and  (not A201) );
 a39376a <=( a39375a  and  a39372a );
 a39377a <=( a39376a  and  a39369a );
 a39380a <=( A233  and  (not A232) );
 a39383a <=( A236  and  A234 );
 a39384a <=( a39383a  and  a39380a );
 a39387a <=( A266  and  (not A265) );
 a39390a <=( A268  and  A267 );
 a39391a <=( a39390a  and  a39387a );
 a39392a <=( a39391a  and  a39384a );
 a39396a <=( (not A168)  and  (not A169) );
 a39397a <=( A170  and  a39396a );
 a39400a <=( (not A166)  and  A167 );
 a39403a <=( A203  and  (not A201) );
 a39404a <=( a39403a  and  a39400a );
 a39405a <=( a39404a  and  a39397a );
 a39408a <=( A233  and  (not A232) );
 a39411a <=( A236  and  A234 );
 a39412a <=( a39411a  and  a39408a );
 a39415a <=( A266  and  (not A265) );
 a39418a <=( A269  and  A267 );
 a39419a <=( a39418a  and  a39415a );
 a39420a <=( a39419a  and  a39412a );
 a39424a <=( (not A168)  and  (not A169) );
 a39425a <=( A170  and  a39424a );
 a39428a <=( (not A166)  and  A167 );
 a39431a <=( A203  and  (not A201) );
 a39432a <=( a39431a  and  a39428a );
 a39433a <=( a39432a  and  a39425a );
 a39436a <=( A233  and  (not A232) );
 a39439a <=( A236  and  A234 );
 a39440a <=( a39439a  and  a39436a );
 a39443a <=( (not A266)  and  A265 );
 a39446a <=( A268  and  A267 );
 a39447a <=( a39446a  and  a39443a );
 a39448a <=( a39447a  and  a39440a );
 a39452a <=( (not A168)  and  (not A169) );
 a39453a <=( A170  and  a39452a );
 a39456a <=( (not A166)  and  A167 );
 a39459a <=( A203  and  (not A201) );
 a39460a <=( a39459a  and  a39456a );
 a39461a <=( a39460a  and  a39453a );
 a39464a <=( A233  and  (not A232) );
 a39467a <=( A236  and  A234 );
 a39468a <=( a39467a  and  a39464a );
 a39471a <=( (not A266)  and  A265 );
 a39474a <=( A269  and  A267 );
 a39475a <=( a39474a  and  a39471a );
 a39476a <=( a39475a  and  a39468a );
 a39480a <=( (not A168)  and  (not A169) );
 a39481a <=( A170  and  a39480a );
 a39484a <=( (not A166)  and  A167 );
 a39487a <=( A203  and  (not A201) );
 a39488a <=( a39487a  and  a39484a );
 a39489a <=( a39488a  and  a39481a );
 a39492a <=( (not A233)  and  A232 );
 a39495a <=( A235  and  A234 );
 a39496a <=( a39495a  and  a39492a );
 a39499a <=( (not A299)  and  A298 );
 a39502a <=( A301  and  A300 );
 a39503a <=( a39502a  and  a39499a );
 a39504a <=( a39503a  and  a39496a );
 a39508a <=( (not A168)  and  (not A169) );
 a39509a <=( A170  and  a39508a );
 a39512a <=( (not A166)  and  A167 );
 a39515a <=( A203  and  (not A201) );
 a39516a <=( a39515a  and  a39512a );
 a39517a <=( a39516a  and  a39509a );
 a39520a <=( (not A233)  and  A232 );
 a39523a <=( A235  and  A234 );
 a39524a <=( a39523a  and  a39520a );
 a39527a <=( (not A299)  and  A298 );
 a39530a <=( A302  and  A300 );
 a39531a <=( a39530a  and  a39527a );
 a39532a <=( a39531a  and  a39524a );
 a39536a <=( (not A168)  and  (not A169) );
 a39537a <=( A170  and  a39536a );
 a39540a <=( (not A166)  and  A167 );
 a39543a <=( A203  and  (not A201) );
 a39544a <=( a39543a  and  a39540a );
 a39545a <=( a39544a  and  a39537a );
 a39548a <=( (not A233)  and  A232 );
 a39551a <=( A235  and  A234 );
 a39552a <=( a39551a  and  a39548a );
 a39555a <=( A299  and  (not A298) );
 a39558a <=( A301  and  A300 );
 a39559a <=( a39558a  and  a39555a );
 a39560a <=( a39559a  and  a39552a );
 a39564a <=( (not A168)  and  (not A169) );
 a39565a <=( A170  and  a39564a );
 a39568a <=( (not A166)  and  A167 );
 a39571a <=( A203  and  (not A201) );
 a39572a <=( a39571a  and  a39568a );
 a39573a <=( a39572a  and  a39565a );
 a39576a <=( (not A233)  and  A232 );
 a39579a <=( A235  and  A234 );
 a39580a <=( a39579a  and  a39576a );
 a39583a <=( A299  and  (not A298) );
 a39586a <=( A302  and  A300 );
 a39587a <=( a39586a  and  a39583a );
 a39588a <=( a39587a  and  a39580a );
 a39592a <=( (not A168)  and  (not A169) );
 a39593a <=( A170  and  a39592a );
 a39596a <=( (not A166)  and  A167 );
 a39599a <=( A203  and  (not A201) );
 a39600a <=( a39599a  and  a39596a );
 a39601a <=( a39600a  and  a39593a );
 a39604a <=( (not A233)  and  A232 );
 a39607a <=( A235  and  A234 );
 a39608a <=( a39607a  and  a39604a );
 a39611a <=( A266  and  (not A265) );
 a39614a <=( A268  and  A267 );
 a39615a <=( a39614a  and  a39611a );
 a39616a <=( a39615a  and  a39608a );
 a39620a <=( (not A168)  and  (not A169) );
 a39621a <=( A170  and  a39620a );
 a39624a <=( (not A166)  and  A167 );
 a39627a <=( A203  and  (not A201) );
 a39628a <=( a39627a  and  a39624a );
 a39629a <=( a39628a  and  a39621a );
 a39632a <=( (not A233)  and  A232 );
 a39635a <=( A235  and  A234 );
 a39636a <=( a39635a  and  a39632a );
 a39639a <=( A266  and  (not A265) );
 a39642a <=( A269  and  A267 );
 a39643a <=( a39642a  and  a39639a );
 a39644a <=( a39643a  and  a39636a );
 a39648a <=( (not A168)  and  (not A169) );
 a39649a <=( A170  and  a39648a );
 a39652a <=( (not A166)  and  A167 );
 a39655a <=( A203  and  (not A201) );
 a39656a <=( a39655a  and  a39652a );
 a39657a <=( a39656a  and  a39649a );
 a39660a <=( (not A233)  and  A232 );
 a39663a <=( A235  and  A234 );
 a39664a <=( a39663a  and  a39660a );
 a39667a <=( (not A266)  and  A265 );
 a39670a <=( A268  and  A267 );
 a39671a <=( a39670a  and  a39667a );
 a39672a <=( a39671a  and  a39664a );
 a39676a <=( (not A168)  and  (not A169) );
 a39677a <=( A170  and  a39676a );
 a39680a <=( (not A166)  and  A167 );
 a39683a <=( A203  and  (not A201) );
 a39684a <=( a39683a  and  a39680a );
 a39685a <=( a39684a  and  a39677a );
 a39688a <=( (not A233)  and  A232 );
 a39691a <=( A235  and  A234 );
 a39692a <=( a39691a  and  a39688a );
 a39695a <=( (not A266)  and  A265 );
 a39698a <=( A269  and  A267 );
 a39699a <=( a39698a  and  a39695a );
 a39700a <=( a39699a  and  a39692a );
 a39704a <=( (not A168)  and  (not A169) );
 a39705a <=( A170  and  a39704a );
 a39708a <=( (not A166)  and  A167 );
 a39711a <=( A203  and  (not A201) );
 a39712a <=( a39711a  and  a39708a );
 a39713a <=( a39712a  and  a39705a );
 a39716a <=( (not A233)  and  A232 );
 a39719a <=( A236  and  A234 );
 a39720a <=( a39719a  and  a39716a );
 a39723a <=( (not A299)  and  A298 );
 a39726a <=( A301  and  A300 );
 a39727a <=( a39726a  and  a39723a );
 a39728a <=( a39727a  and  a39720a );
 a39732a <=( (not A168)  and  (not A169) );
 a39733a <=( A170  and  a39732a );
 a39736a <=( (not A166)  and  A167 );
 a39739a <=( A203  and  (not A201) );
 a39740a <=( a39739a  and  a39736a );
 a39741a <=( a39740a  and  a39733a );
 a39744a <=( (not A233)  and  A232 );
 a39747a <=( A236  and  A234 );
 a39748a <=( a39747a  and  a39744a );
 a39751a <=( (not A299)  and  A298 );
 a39754a <=( A302  and  A300 );
 a39755a <=( a39754a  and  a39751a );
 a39756a <=( a39755a  and  a39748a );
 a39760a <=( (not A168)  and  (not A169) );
 a39761a <=( A170  and  a39760a );
 a39764a <=( (not A166)  and  A167 );
 a39767a <=( A203  and  (not A201) );
 a39768a <=( a39767a  and  a39764a );
 a39769a <=( a39768a  and  a39761a );
 a39772a <=( (not A233)  and  A232 );
 a39775a <=( A236  and  A234 );
 a39776a <=( a39775a  and  a39772a );
 a39779a <=( A299  and  (not A298) );
 a39782a <=( A301  and  A300 );
 a39783a <=( a39782a  and  a39779a );
 a39784a <=( a39783a  and  a39776a );
 a39788a <=( (not A168)  and  (not A169) );
 a39789a <=( A170  and  a39788a );
 a39792a <=( (not A166)  and  A167 );
 a39795a <=( A203  and  (not A201) );
 a39796a <=( a39795a  and  a39792a );
 a39797a <=( a39796a  and  a39789a );
 a39800a <=( (not A233)  and  A232 );
 a39803a <=( A236  and  A234 );
 a39804a <=( a39803a  and  a39800a );
 a39807a <=( A299  and  (not A298) );
 a39810a <=( A302  and  A300 );
 a39811a <=( a39810a  and  a39807a );
 a39812a <=( a39811a  and  a39804a );
 a39816a <=( (not A168)  and  (not A169) );
 a39817a <=( A170  and  a39816a );
 a39820a <=( (not A166)  and  A167 );
 a39823a <=( A203  and  (not A201) );
 a39824a <=( a39823a  and  a39820a );
 a39825a <=( a39824a  and  a39817a );
 a39828a <=( (not A233)  and  A232 );
 a39831a <=( A236  and  A234 );
 a39832a <=( a39831a  and  a39828a );
 a39835a <=( A266  and  (not A265) );
 a39838a <=( A268  and  A267 );
 a39839a <=( a39838a  and  a39835a );
 a39840a <=( a39839a  and  a39832a );
 a39844a <=( (not A168)  and  (not A169) );
 a39845a <=( A170  and  a39844a );
 a39848a <=( (not A166)  and  A167 );
 a39851a <=( A203  and  (not A201) );
 a39852a <=( a39851a  and  a39848a );
 a39853a <=( a39852a  and  a39845a );
 a39856a <=( (not A233)  and  A232 );
 a39859a <=( A236  and  A234 );
 a39860a <=( a39859a  and  a39856a );
 a39863a <=( A266  and  (not A265) );
 a39866a <=( A269  and  A267 );
 a39867a <=( a39866a  and  a39863a );
 a39868a <=( a39867a  and  a39860a );
 a39872a <=( (not A168)  and  (not A169) );
 a39873a <=( A170  and  a39872a );
 a39876a <=( (not A166)  and  A167 );
 a39879a <=( A203  and  (not A201) );
 a39880a <=( a39879a  and  a39876a );
 a39881a <=( a39880a  and  a39873a );
 a39884a <=( (not A233)  and  A232 );
 a39887a <=( A236  and  A234 );
 a39888a <=( a39887a  and  a39884a );
 a39891a <=( (not A266)  and  A265 );
 a39894a <=( A268  and  A267 );
 a39895a <=( a39894a  and  a39891a );
 a39896a <=( a39895a  and  a39888a );
 a39900a <=( (not A168)  and  (not A169) );
 a39901a <=( A170  and  a39900a );
 a39904a <=( (not A166)  and  A167 );
 a39907a <=( A203  and  (not A201) );
 a39908a <=( a39907a  and  a39904a );
 a39909a <=( a39908a  and  a39901a );
 a39912a <=( (not A233)  and  A232 );
 a39915a <=( A236  and  A234 );
 a39916a <=( a39915a  and  a39912a );
 a39919a <=( (not A266)  and  A265 );
 a39922a <=( A269  and  A267 );
 a39923a <=( a39922a  and  a39919a );
 a39924a <=( a39923a  and  a39916a );
 a39928a <=( (not A168)  and  (not A169) );
 a39929a <=( A170  and  a39928a );
 a39932a <=( (not A166)  and  A167 );
 a39935a <=( A200  and  A199 );
 a39936a <=( a39935a  and  a39932a );
 a39937a <=( a39936a  and  a39929a );
 a39940a <=( A233  and  (not A232) );
 a39943a <=( A235  and  A234 );
 a39944a <=( a39943a  and  a39940a );
 a39947a <=( (not A299)  and  A298 );
 a39950a <=( A301  and  A300 );
 a39951a <=( a39950a  and  a39947a );
 a39952a <=( a39951a  and  a39944a );
 a39956a <=( (not A168)  and  (not A169) );
 a39957a <=( A170  and  a39956a );
 a39960a <=( (not A166)  and  A167 );
 a39963a <=( A200  and  A199 );
 a39964a <=( a39963a  and  a39960a );
 a39965a <=( a39964a  and  a39957a );
 a39968a <=( A233  and  (not A232) );
 a39971a <=( A235  and  A234 );
 a39972a <=( a39971a  and  a39968a );
 a39975a <=( (not A299)  and  A298 );
 a39978a <=( A302  and  A300 );
 a39979a <=( a39978a  and  a39975a );
 a39980a <=( a39979a  and  a39972a );
 a39984a <=( (not A168)  and  (not A169) );
 a39985a <=( A170  and  a39984a );
 a39988a <=( (not A166)  and  A167 );
 a39991a <=( A200  and  A199 );
 a39992a <=( a39991a  and  a39988a );
 a39993a <=( a39992a  and  a39985a );
 a39996a <=( A233  and  (not A232) );
 a39999a <=( A235  and  A234 );
 a40000a <=( a39999a  and  a39996a );
 a40003a <=( A299  and  (not A298) );
 a40006a <=( A301  and  A300 );
 a40007a <=( a40006a  and  a40003a );
 a40008a <=( a40007a  and  a40000a );
 a40012a <=( (not A168)  and  (not A169) );
 a40013a <=( A170  and  a40012a );
 a40016a <=( (not A166)  and  A167 );
 a40019a <=( A200  and  A199 );
 a40020a <=( a40019a  and  a40016a );
 a40021a <=( a40020a  and  a40013a );
 a40024a <=( A233  and  (not A232) );
 a40027a <=( A235  and  A234 );
 a40028a <=( a40027a  and  a40024a );
 a40031a <=( A299  and  (not A298) );
 a40034a <=( A302  and  A300 );
 a40035a <=( a40034a  and  a40031a );
 a40036a <=( a40035a  and  a40028a );
 a40040a <=( (not A168)  and  (not A169) );
 a40041a <=( A170  and  a40040a );
 a40044a <=( (not A166)  and  A167 );
 a40047a <=( A200  and  A199 );
 a40048a <=( a40047a  and  a40044a );
 a40049a <=( a40048a  and  a40041a );
 a40052a <=( A233  and  (not A232) );
 a40055a <=( A235  and  A234 );
 a40056a <=( a40055a  and  a40052a );
 a40059a <=( A266  and  (not A265) );
 a40062a <=( A268  and  A267 );
 a40063a <=( a40062a  and  a40059a );
 a40064a <=( a40063a  and  a40056a );
 a40068a <=( (not A168)  and  (not A169) );
 a40069a <=( A170  and  a40068a );
 a40072a <=( (not A166)  and  A167 );
 a40075a <=( A200  and  A199 );
 a40076a <=( a40075a  and  a40072a );
 a40077a <=( a40076a  and  a40069a );
 a40080a <=( A233  and  (not A232) );
 a40083a <=( A235  and  A234 );
 a40084a <=( a40083a  and  a40080a );
 a40087a <=( A266  and  (not A265) );
 a40090a <=( A269  and  A267 );
 a40091a <=( a40090a  and  a40087a );
 a40092a <=( a40091a  and  a40084a );
 a40096a <=( (not A168)  and  (not A169) );
 a40097a <=( A170  and  a40096a );
 a40100a <=( (not A166)  and  A167 );
 a40103a <=( A200  and  A199 );
 a40104a <=( a40103a  and  a40100a );
 a40105a <=( a40104a  and  a40097a );
 a40108a <=( A233  and  (not A232) );
 a40111a <=( A235  and  A234 );
 a40112a <=( a40111a  and  a40108a );
 a40115a <=( (not A266)  and  A265 );
 a40118a <=( A268  and  A267 );
 a40119a <=( a40118a  and  a40115a );
 a40120a <=( a40119a  and  a40112a );
 a40124a <=( (not A168)  and  (not A169) );
 a40125a <=( A170  and  a40124a );
 a40128a <=( (not A166)  and  A167 );
 a40131a <=( A200  and  A199 );
 a40132a <=( a40131a  and  a40128a );
 a40133a <=( a40132a  and  a40125a );
 a40136a <=( A233  and  (not A232) );
 a40139a <=( A235  and  A234 );
 a40140a <=( a40139a  and  a40136a );
 a40143a <=( (not A266)  and  A265 );
 a40146a <=( A269  and  A267 );
 a40147a <=( a40146a  and  a40143a );
 a40148a <=( a40147a  and  a40140a );
 a40152a <=( (not A168)  and  (not A169) );
 a40153a <=( A170  and  a40152a );
 a40156a <=( (not A166)  and  A167 );
 a40159a <=( A200  and  A199 );
 a40160a <=( a40159a  and  a40156a );
 a40161a <=( a40160a  and  a40153a );
 a40164a <=( A233  and  (not A232) );
 a40167a <=( A236  and  A234 );
 a40168a <=( a40167a  and  a40164a );
 a40171a <=( (not A299)  and  A298 );
 a40174a <=( A301  and  A300 );
 a40175a <=( a40174a  and  a40171a );
 a40176a <=( a40175a  and  a40168a );
 a40180a <=( (not A168)  and  (not A169) );
 a40181a <=( A170  and  a40180a );
 a40184a <=( (not A166)  and  A167 );
 a40187a <=( A200  and  A199 );
 a40188a <=( a40187a  and  a40184a );
 a40189a <=( a40188a  and  a40181a );
 a40192a <=( A233  and  (not A232) );
 a40195a <=( A236  and  A234 );
 a40196a <=( a40195a  and  a40192a );
 a40199a <=( (not A299)  and  A298 );
 a40202a <=( A302  and  A300 );
 a40203a <=( a40202a  and  a40199a );
 a40204a <=( a40203a  and  a40196a );
 a40208a <=( (not A168)  and  (not A169) );
 a40209a <=( A170  and  a40208a );
 a40212a <=( (not A166)  and  A167 );
 a40215a <=( A200  and  A199 );
 a40216a <=( a40215a  and  a40212a );
 a40217a <=( a40216a  and  a40209a );
 a40220a <=( A233  and  (not A232) );
 a40223a <=( A236  and  A234 );
 a40224a <=( a40223a  and  a40220a );
 a40227a <=( A299  and  (not A298) );
 a40230a <=( A301  and  A300 );
 a40231a <=( a40230a  and  a40227a );
 a40232a <=( a40231a  and  a40224a );
 a40236a <=( (not A168)  and  (not A169) );
 a40237a <=( A170  and  a40236a );
 a40240a <=( (not A166)  and  A167 );
 a40243a <=( A200  and  A199 );
 a40244a <=( a40243a  and  a40240a );
 a40245a <=( a40244a  and  a40237a );
 a40248a <=( A233  and  (not A232) );
 a40251a <=( A236  and  A234 );
 a40252a <=( a40251a  and  a40248a );
 a40255a <=( A299  and  (not A298) );
 a40258a <=( A302  and  A300 );
 a40259a <=( a40258a  and  a40255a );
 a40260a <=( a40259a  and  a40252a );
 a40264a <=( (not A168)  and  (not A169) );
 a40265a <=( A170  and  a40264a );
 a40268a <=( (not A166)  and  A167 );
 a40271a <=( A200  and  A199 );
 a40272a <=( a40271a  and  a40268a );
 a40273a <=( a40272a  and  a40265a );
 a40276a <=( A233  and  (not A232) );
 a40279a <=( A236  and  A234 );
 a40280a <=( a40279a  and  a40276a );
 a40283a <=( A266  and  (not A265) );
 a40286a <=( A268  and  A267 );
 a40287a <=( a40286a  and  a40283a );
 a40288a <=( a40287a  and  a40280a );
 a40292a <=( (not A168)  and  (not A169) );
 a40293a <=( A170  and  a40292a );
 a40296a <=( (not A166)  and  A167 );
 a40299a <=( A200  and  A199 );
 a40300a <=( a40299a  and  a40296a );
 a40301a <=( a40300a  and  a40293a );
 a40304a <=( A233  and  (not A232) );
 a40307a <=( A236  and  A234 );
 a40308a <=( a40307a  and  a40304a );
 a40311a <=( A266  and  (not A265) );
 a40314a <=( A269  and  A267 );
 a40315a <=( a40314a  and  a40311a );
 a40316a <=( a40315a  and  a40308a );
 a40320a <=( (not A168)  and  (not A169) );
 a40321a <=( A170  and  a40320a );
 a40324a <=( (not A166)  and  A167 );
 a40327a <=( A200  and  A199 );
 a40328a <=( a40327a  and  a40324a );
 a40329a <=( a40328a  and  a40321a );
 a40332a <=( A233  and  (not A232) );
 a40335a <=( A236  and  A234 );
 a40336a <=( a40335a  and  a40332a );
 a40339a <=( (not A266)  and  A265 );
 a40342a <=( A268  and  A267 );
 a40343a <=( a40342a  and  a40339a );
 a40344a <=( a40343a  and  a40336a );
 a40348a <=( (not A168)  and  (not A169) );
 a40349a <=( A170  and  a40348a );
 a40352a <=( (not A166)  and  A167 );
 a40355a <=( A200  and  A199 );
 a40356a <=( a40355a  and  a40352a );
 a40357a <=( a40356a  and  a40349a );
 a40360a <=( A233  and  (not A232) );
 a40363a <=( A236  and  A234 );
 a40364a <=( a40363a  and  a40360a );
 a40367a <=( (not A266)  and  A265 );
 a40370a <=( A269  and  A267 );
 a40371a <=( a40370a  and  a40367a );
 a40372a <=( a40371a  and  a40364a );
 a40376a <=( (not A168)  and  (not A169) );
 a40377a <=( A170  and  a40376a );
 a40380a <=( (not A166)  and  A167 );
 a40383a <=( A200  and  A199 );
 a40384a <=( a40383a  and  a40380a );
 a40385a <=( a40384a  and  a40377a );
 a40388a <=( (not A233)  and  A232 );
 a40391a <=( A235  and  A234 );
 a40392a <=( a40391a  and  a40388a );
 a40395a <=( (not A299)  and  A298 );
 a40398a <=( A301  and  A300 );
 a40399a <=( a40398a  and  a40395a );
 a40400a <=( a40399a  and  a40392a );
 a40404a <=( (not A168)  and  (not A169) );
 a40405a <=( A170  and  a40404a );
 a40408a <=( (not A166)  and  A167 );
 a40411a <=( A200  and  A199 );
 a40412a <=( a40411a  and  a40408a );
 a40413a <=( a40412a  and  a40405a );
 a40416a <=( (not A233)  and  A232 );
 a40419a <=( A235  and  A234 );
 a40420a <=( a40419a  and  a40416a );
 a40423a <=( (not A299)  and  A298 );
 a40426a <=( A302  and  A300 );
 a40427a <=( a40426a  and  a40423a );
 a40428a <=( a40427a  and  a40420a );
 a40432a <=( (not A168)  and  (not A169) );
 a40433a <=( A170  and  a40432a );
 a40436a <=( (not A166)  and  A167 );
 a40439a <=( A200  and  A199 );
 a40440a <=( a40439a  and  a40436a );
 a40441a <=( a40440a  and  a40433a );
 a40444a <=( (not A233)  and  A232 );
 a40447a <=( A235  and  A234 );
 a40448a <=( a40447a  and  a40444a );
 a40451a <=( A299  and  (not A298) );
 a40454a <=( A301  and  A300 );
 a40455a <=( a40454a  and  a40451a );
 a40456a <=( a40455a  and  a40448a );
 a40460a <=( (not A168)  and  (not A169) );
 a40461a <=( A170  and  a40460a );
 a40464a <=( (not A166)  and  A167 );
 a40467a <=( A200  and  A199 );
 a40468a <=( a40467a  and  a40464a );
 a40469a <=( a40468a  and  a40461a );
 a40472a <=( (not A233)  and  A232 );
 a40475a <=( A235  and  A234 );
 a40476a <=( a40475a  and  a40472a );
 a40479a <=( A299  and  (not A298) );
 a40482a <=( A302  and  A300 );
 a40483a <=( a40482a  and  a40479a );
 a40484a <=( a40483a  and  a40476a );
 a40488a <=( (not A168)  and  (not A169) );
 a40489a <=( A170  and  a40488a );
 a40492a <=( (not A166)  and  A167 );
 a40495a <=( A200  and  A199 );
 a40496a <=( a40495a  and  a40492a );
 a40497a <=( a40496a  and  a40489a );
 a40500a <=( (not A233)  and  A232 );
 a40503a <=( A235  and  A234 );
 a40504a <=( a40503a  and  a40500a );
 a40507a <=( A266  and  (not A265) );
 a40510a <=( A268  and  A267 );
 a40511a <=( a40510a  and  a40507a );
 a40512a <=( a40511a  and  a40504a );
 a40516a <=( (not A168)  and  (not A169) );
 a40517a <=( A170  and  a40516a );
 a40520a <=( (not A166)  and  A167 );
 a40523a <=( A200  and  A199 );
 a40524a <=( a40523a  and  a40520a );
 a40525a <=( a40524a  and  a40517a );
 a40528a <=( (not A233)  and  A232 );
 a40531a <=( A235  and  A234 );
 a40532a <=( a40531a  and  a40528a );
 a40535a <=( A266  and  (not A265) );
 a40538a <=( A269  and  A267 );
 a40539a <=( a40538a  and  a40535a );
 a40540a <=( a40539a  and  a40532a );
 a40544a <=( (not A168)  and  (not A169) );
 a40545a <=( A170  and  a40544a );
 a40548a <=( (not A166)  and  A167 );
 a40551a <=( A200  and  A199 );
 a40552a <=( a40551a  and  a40548a );
 a40553a <=( a40552a  and  a40545a );
 a40556a <=( (not A233)  and  A232 );
 a40559a <=( A235  and  A234 );
 a40560a <=( a40559a  and  a40556a );
 a40563a <=( (not A266)  and  A265 );
 a40566a <=( A268  and  A267 );
 a40567a <=( a40566a  and  a40563a );
 a40568a <=( a40567a  and  a40560a );
 a40572a <=( (not A168)  and  (not A169) );
 a40573a <=( A170  and  a40572a );
 a40576a <=( (not A166)  and  A167 );
 a40579a <=( A200  and  A199 );
 a40580a <=( a40579a  and  a40576a );
 a40581a <=( a40580a  and  a40573a );
 a40584a <=( (not A233)  and  A232 );
 a40587a <=( A235  and  A234 );
 a40588a <=( a40587a  and  a40584a );
 a40591a <=( (not A266)  and  A265 );
 a40594a <=( A269  and  A267 );
 a40595a <=( a40594a  and  a40591a );
 a40596a <=( a40595a  and  a40588a );
 a40600a <=( (not A168)  and  (not A169) );
 a40601a <=( A170  and  a40600a );
 a40604a <=( (not A166)  and  A167 );
 a40607a <=( A200  and  A199 );
 a40608a <=( a40607a  and  a40604a );
 a40609a <=( a40608a  and  a40601a );
 a40612a <=( (not A233)  and  A232 );
 a40615a <=( A236  and  A234 );
 a40616a <=( a40615a  and  a40612a );
 a40619a <=( (not A299)  and  A298 );
 a40622a <=( A301  and  A300 );
 a40623a <=( a40622a  and  a40619a );
 a40624a <=( a40623a  and  a40616a );
 a40628a <=( (not A168)  and  (not A169) );
 a40629a <=( A170  and  a40628a );
 a40632a <=( (not A166)  and  A167 );
 a40635a <=( A200  and  A199 );
 a40636a <=( a40635a  and  a40632a );
 a40637a <=( a40636a  and  a40629a );
 a40640a <=( (not A233)  and  A232 );
 a40643a <=( A236  and  A234 );
 a40644a <=( a40643a  and  a40640a );
 a40647a <=( (not A299)  and  A298 );
 a40650a <=( A302  and  A300 );
 a40651a <=( a40650a  and  a40647a );
 a40652a <=( a40651a  and  a40644a );
 a40656a <=( (not A168)  and  (not A169) );
 a40657a <=( A170  and  a40656a );
 a40660a <=( (not A166)  and  A167 );
 a40663a <=( A200  and  A199 );
 a40664a <=( a40663a  and  a40660a );
 a40665a <=( a40664a  and  a40657a );
 a40668a <=( (not A233)  and  A232 );
 a40671a <=( A236  and  A234 );
 a40672a <=( a40671a  and  a40668a );
 a40675a <=( A299  and  (not A298) );
 a40678a <=( A301  and  A300 );
 a40679a <=( a40678a  and  a40675a );
 a40680a <=( a40679a  and  a40672a );
 a40684a <=( (not A168)  and  (not A169) );
 a40685a <=( A170  and  a40684a );
 a40688a <=( (not A166)  and  A167 );
 a40691a <=( A200  and  A199 );
 a40692a <=( a40691a  and  a40688a );
 a40693a <=( a40692a  and  a40685a );
 a40696a <=( (not A233)  and  A232 );
 a40699a <=( A236  and  A234 );
 a40700a <=( a40699a  and  a40696a );
 a40703a <=( A299  and  (not A298) );
 a40706a <=( A302  and  A300 );
 a40707a <=( a40706a  and  a40703a );
 a40708a <=( a40707a  and  a40700a );
 a40712a <=( (not A168)  and  (not A169) );
 a40713a <=( A170  and  a40712a );
 a40716a <=( (not A166)  and  A167 );
 a40719a <=( A200  and  A199 );
 a40720a <=( a40719a  and  a40716a );
 a40721a <=( a40720a  and  a40713a );
 a40724a <=( (not A233)  and  A232 );
 a40727a <=( A236  and  A234 );
 a40728a <=( a40727a  and  a40724a );
 a40731a <=( A266  and  (not A265) );
 a40734a <=( A268  and  A267 );
 a40735a <=( a40734a  and  a40731a );
 a40736a <=( a40735a  and  a40728a );
 a40740a <=( (not A168)  and  (not A169) );
 a40741a <=( A170  and  a40740a );
 a40744a <=( (not A166)  and  A167 );
 a40747a <=( A200  and  A199 );
 a40748a <=( a40747a  and  a40744a );
 a40749a <=( a40748a  and  a40741a );
 a40752a <=( (not A233)  and  A232 );
 a40755a <=( A236  and  A234 );
 a40756a <=( a40755a  and  a40752a );
 a40759a <=( A266  and  (not A265) );
 a40762a <=( A269  and  A267 );
 a40763a <=( a40762a  and  a40759a );
 a40764a <=( a40763a  and  a40756a );
 a40768a <=( (not A168)  and  (not A169) );
 a40769a <=( A170  and  a40768a );
 a40772a <=( (not A166)  and  A167 );
 a40775a <=( A200  and  A199 );
 a40776a <=( a40775a  and  a40772a );
 a40777a <=( a40776a  and  a40769a );
 a40780a <=( (not A233)  and  A232 );
 a40783a <=( A236  and  A234 );
 a40784a <=( a40783a  and  a40780a );
 a40787a <=( (not A266)  and  A265 );
 a40790a <=( A268  and  A267 );
 a40791a <=( a40790a  and  a40787a );
 a40792a <=( a40791a  and  a40784a );
 a40796a <=( (not A168)  and  (not A169) );
 a40797a <=( A170  and  a40796a );
 a40800a <=( (not A166)  and  A167 );
 a40803a <=( A200  and  A199 );
 a40804a <=( a40803a  and  a40800a );
 a40805a <=( a40804a  and  a40797a );
 a40808a <=( (not A233)  and  A232 );
 a40811a <=( A236  and  A234 );
 a40812a <=( a40811a  and  a40808a );
 a40815a <=( (not A266)  and  A265 );
 a40818a <=( A269  and  A267 );
 a40819a <=( a40818a  and  a40815a );
 a40820a <=( a40819a  and  a40812a );
 a40824a <=( (not A168)  and  (not A169) );
 a40825a <=( A170  and  a40824a );
 a40828a <=( (not A166)  and  A167 );
 a40831a <=( (not A200)  and  (not A199) );
 a40832a <=( a40831a  and  a40828a );
 a40833a <=( a40832a  and  a40825a );
 a40836a <=( A233  and  (not A232) );
 a40839a <=( A235  and  A234 );
 a40840a <=( a40839a  and  a40836a );
 a40843a <=( (not A299)  and  A298 );
 a40846a <=( A301  and  A300 );
 a40847a <=( a40846a  and  a40843a );
 a40848a <=( a40847a  and  a40840a );
 a40852a <=( (not A168)  and  (not A169) );
 a40853a <=( A170  and  a40852a );
 a40856a <=( (not A166)  and  A167 );
 a40859a <=( (not A200)  and  (not A199) );
 a40860a <=( a40859a  and  a40856a );
 a40861a <=( a40860a  and  a40853a );
 a40864a <=( A233  and  (not A232) );
 a40867a <=( A235  and  A234 );
 a40868a <=( a40867a  and  a40864a );
 a40871a <=( (not A299)  and  A298 );
 a40874a <=( A302  and  A300 );
 a40875a <=( a40874a  and  a40871a );
 a40876a <=( a40875a  and  a40868a );
 a40880a <=( (not A168)  and  (not A169) );
 a40881a <=( A170  and  a40880a );
 a40884a <=( (not A166)  and  A167 );
 a40887a <=( (not A200)  and  (not A199) );
 a40888a <=( a40887a  and  a40884a );
 a40889a <=( a40888a  and  a40881a );
 a40892a <=( A233  and  (not A232) );
 a40895a <=( A235  and  A234 );
 a40896a <=( a40895a  and  a40892a );
 a40899a <=( A299  and  (not A298) );
 a40902a <=( A301  and  A300 );
 a40903a <=( a40902a  and  a40899a );
 a40904a <=( a40903a  and  a40896a );
 a40908a <=( (not A168)  and  (not A169) );
 a40909a <=( A170  and  a40908a );
 a40912a <=( (not A166)  and  A167 );
 a40915a <=( (not A200)  and  (not A199) );
 a40916a <=( a40915a  and  a40912a );
 a40917a <=( a40916a  and  a40909a );
 a40920a <=( A233  and  (not A232) );
 a40923a <=( A235  and  A234 );
 a40924a <=( a40923a  and  a40920a );
 a40927a <=( A299  and  (not A298) );
 a40930a <=( A302  and  A300 );
 a40931a <=( a40930a  and  a40927a );
 a40932a <=( a40931a  and  a40924a );
 a40936a <=( (not A168)  and  (not A169) );
 a40937a <=( A170  and  a40936a );
 a40940a <=( (not A166)  and  A167 );
 a40943a <=( (not A200)  and  (not A199) );
 a40944a <=( a40943a  and  a40940a );
 a40945a <=( a40944a  and  a40937a );
 a40948a <=( A233  and  (not A232) );
 a40951a <=( A235  and  A234 );
 a40952a <=( a40951a  and  a40948a );
 a40955a <=( A266  and  (not A265) );
 a40958a <=( A268  and  A267 );
 a40959a <=( a40958a  and  a40955a );
 a40960a <=( a40959a  and  a40952a );
 a40964a <=( (not A168)  and  (not A169) );
 a40965a <=( A170  and  a40964a );
 a40968a <=( (not A166)  and  A167 );
 a40971a <=( (not A200)  and  (not A199) );
 a40972a <=( a40971a  and  a40968a );
 a40973a <=( a40972a  and  a40965a );
 a40976a <=( A233  and  (not A232) );
 a40979a <=( A235  and  A234 );
 a40980a <=( a40979a  and  a40976a );
 a40983a <=( A266  and  (not A265) );
 a40986a <=( A269  and  A267 );
 a40987a <=( a40986a  and  a40983a );
 a40988a <=( a40987a  and  a40980a );
 a40992a <=( (not A168)  and  (not A169) );
 a40993a <=( A170  and  a40992a );
 a40996a <=( (not A166)  and  A167 );
 a40999a <=( (not A200)  and  (not A199) );
 a41000a <=( a40999a  and  a40996a );
 a41001a <=( a41000a  and  a40993a );
 a41004a <=( A233  and  (not A232) );
 a41007a <=( A235  and  A234 );
 a41008a <=( a41007a  and  a41004a );
 a41011a <=( (not A266)  and  A265 );
 a41014a <=( A268  and  A267 );
 a41015a <=( a41014a  and  a41011a );
 a41016a <=( a41015a  and  a41008a );
 a41020a <=( (not A168)  and  (not A169) );
 a41021a <=( A170  and  a41020a );
 a41024a <=( (not A166)  and  A167 );
 a41027a <=( (not A200)  and  (not A199) );
 a41028a <=( a41027a  and  a41024a );
 a41029a <=( a41028a  and  a41021a );
 a41032a <=( A233  and  (not A232) );
 a41035a <=( A235  and  A234 );
 a41036a <=( a41035a  and  a41032a );
 a41039a <=( (not A266)  and  A265 );
 a41042a <=( A269  and  A267 );
 a41043a <=( a41042a  and  a41039a );
 a41044a <=( a41043a  and  a41036a );
 a41048a <=( (not A168)  and  (not A169) );
 a41049a <=( A170  and  a41048a );
 a41052a <=( (not A166)  and  A167 );
 a41055a <=( (not A200)  and  (not A199) );
 a41056a <=( a41055a  and  a41052a );
 a41057a <=( a41056a  and  a41049a );
 a41060a <=( A233  and  (not A232) );
 a41063a <=( A236  and  A234 );
 a41064a <=( a41063a  and  a41060a );
 a41067a <=( (not A299)  and  A298 );
 a41070a <=( A301  and  A300 );
 a41071a <=( a41070a  and  a41067a );
 a41072a <=( a41071a  and  a41064a );
 a41076a <=( (not A168)  and  (not A169) );
 a41077a <=( A170  and  a41076a );
 a41080a <=( (not A166)  and  A167 );
 a41083a <=( (not A200)  and  (not A199) );
 a41084a <=( a41083a  and  a41080a );
 a41085a <=( a41084a  and  a41077a );
 a41088a <=( A233  and  (not A232) );
 a41091a <=( A236  and  A234 );
 a41092a <=( a41091a  and  a41088a );
 a41095a <=( (not A299)  and  A298 );
 a41098a <=( A302  and  A300 );
 a41099a <=( a41098a  and  a41095a );
 a41100a <=( a41099a  and  a41092a );
 a41104a <=( (not A168)  and  (not A169) );
 a41105a <=( A170  and  a41104a );
 a41108a <=( (not A166)  and  A167 );
 a41111a <=( (not A200)  and  (not A199) );
 a41112a <=( a41111a  and  a41108a );
 a41113a <=( a41112a  and  a41105a );
 a41116a <=( A233  and  (not A232) );
 a41119a <=( A236  and  A234 );
 a41120a <=( a41119a  and  a41116a );
 a41123a <=( A299  and  (not A298) );
 a41126a <=( A301  and  A300 );
 a41127a <=( a41126a  and  a41123a );
 a41128a <=( a41127a  and  a41120a );
 a41132a <=( (not A168)  and  (not A169) );
 a41133a <=( A170  and  a41132a );
 a41136a <=( (not A166)  and  A167 );
 a41139a <=( (not A200)  and  (not A199) );
 a41140a <=( a41139a  and  a41136a );
 a41141a <=( a41140a  and  a41133a );
 a41144a <=( A233  and  (not A232) );
 a41147a <=( A236  and  A234 );
 a41148a <=( a41147a  and  a41144a );
 a41151a <=( A299  and  (not A298) );
 a41154a <=( A302  and  A300 );
 a41155a <=( a41154a  and  a41151a );
 a41156a <=( a41155a  and  a41148a );
 a41160a <=( (not A168)  and  (not A169) );
 a41161a <=( A170  and  a41160a );
 a41164a <=( (not A166)  and  A167 );
 a41167a <=( (not A200)  and  (not A199) );
 a41168a <=( a41167a  and  a41164a );
 a41169a <=( a41168a  and  a41161a );
 a41172a <=( A233  and  (not A232) );
 a41175a <=( A236  and  A234 );
 a41176a <=( a41175a  and  a41172a );
 a41179a <=( A266  and  (not A265) );
 a41182a <=( A268  and  A267 );
 a41183a <=( a41182a  and  a41179a );
 a41184a <=( a41183a  and  a41176a );
 a41188a <=( (not A168)  and  (not A169) );
 a41189a <=( A170  and  a41188a );
 a41192a <=( (not A166)  and  A167 );
 a41195a <=( (not A200)  and  (not A199) );
 a41196a <=( a41195a  and  a41192a );
 a41197a <=( a41196a  and  a41189a );
 a41200a <=( A233  and  (not A232) );
 a41203a <=( A236  and  A234 );
 a41204a <=( a41203a  and  a41200a );
 a41207a <=( A266  and  (not A265) );
 a41210a <=( A269  and  A267 );
 a41211a <=( a41210a  and  a41207a );
 a41212a <=( a41211a  and  a41204a );
 a41216a <=( (not A168)  and  (not A169) );
 a41217a <=( A170  and  a41216a );
 a41220a <=( (not A166)  and  A167 );
 a41223a <=( (not A200)  and  (not A199) );
 a41224a <=( a41223a  and  a41220a );
 a41225a <=( a41224a  and  a41217a );
 a41228a <=( A233  and  (not A232) );
 a41231a <=( A236  and  A234 );
 a41232a <=( a41231a  and  a41228a );
 a41235a <=( (not A266)  and  A265 );
 a41238a <=( A268  and  A267 );
 a41239a <=( a41238a  and  a41235a );
 a41240a <=( a41239a  and  a41232a );
 a41244a <=( (not A168)  and  (not A169) );
 a41245a <=( A170  and  a41244a );
 a41248a <=( (not A166)  and  A167 );
 a41251a <=( (not A200)  and  (not A199) );
 a41252a <=( a41251a  and  a41248a );
 a41253a <=( a41252a  and  a41245a );
 a41256a <=( A233  and  (not A232) );
 a41259a <=( A236  and  A234 );
 a41260a <=( a41259a  and  a41256a );
 a41263a <=( (not A266)  and  A265 );
 a41266a <=( A269  and  A267 );
 a41267a <=( a41266a  and  a41263a );
 a41268a <=( a41267a  and  a41260a );
 a41272a <=( (not A168)  and  (not A169) );
 a41273a <=( A170  and  a41272a );
 a41276a <=( (not A166)  and  A167 );
 a41279a <=( (not A200)  and  (not A199) );
 a41280a <=( a41279a  and  a41276a );
 a41281a <=( a41280a  and  a41273a );
 a41284a <=( (not A233)  and  A232 );
 a41287a <=( A235  and  A234 );
 a41288a <=( a41287a  and  a41284a );
 a41291a <=( (not A299)  and  A298 );
 a41294a <=( A301  and  A300 );
 a41295a <=( a41294a  and  a41291a );
 a41296a <=( a41295a  and  a41288a );
 a41300a <=( (not A168)  and  (not A169) );
 a41301a <=( A170  and  a41300a );
 a41304a <=( (not A166)  and  A167 );
 a41307a <=( (not A200)  and  (not A199) );
 a41308a <=( a41307a  and  a41304a );
 a41309a <=( a41308a  and  a41301a );
 a41312a <=( (not A233)  and  A232 );
 a41315a <=( A235  and  A234 );
 a41316a <=( a41315a  and  a41312a );
 a41319a <=( (not A299)  and  A298 );
 a41322a <=( A302  and  A300 );
 a41323a <=( a41322a  and  a41319a );
 a41324a <=( a41323a  and  a41316a );
 a41328a <=( (not A168)  and  (not A169) );
 a41329a <=( A170  and  a41328a );
 a41332a <=( (not A166)  and  A167 );
 a41335a <=( (not A200)  and  (not A199) );
 a41336a <=( a41335a  and  a41332a );
 a41337a <=( a41336a  and  a41329a );
 a41340a <=( (not A233)  and  A232 );
 a41343a <=( A235  and  A234 );
 a41344a <=( a41343a  and  a41340a );
 a41347a <=( A299  and  (not A298) );
 a41350a <=( A301  and  A300 );
 a41351a <=( a41350a  and  a41347a );
 a41352a <=( a41351a  and  a41344a );
 a41356a <=( (not A168)  and  (not A169) );
 a41357a <=( A170  and  a41356a );
 a41360a <=( (not A166)  and  A167 );
 a41363a <=( (not A200)  and  (not A199) );
 a41364a <=( a41363a  and  a41360a );
 a41365a <=( a41364a  and  a41357a );
 a41368a <=( (not A233)  and  A232 );
 a41371a <=( A235  and  A234 );
 a41372a <=( a41371a  and  a41368a );
 a41375a <=( A299  and  (not A298) );
 a41378a <=( A302  and  A300 );
 a41379a <=( a41378a  and  a41375a );
 a41380a <=( a41379a  and  a41372a );
 a41384a <=( (not A168)  and  (not A169) );
 a41385a <=( A170  and  a41384a );
 a41388a <=( (not A166)  and  A167 );
 a41391a <=( (not A200)  and  (not A199) );
 a41392a <=( a41391a  and  a41388a );
 a41393a <=( a41392a  and  a41385a );
 a41396a <=( (not A233)  and  A232 );
 a41399a <=( A235  and  A234 );
 a41400a <=( a41399a  and  a41396a );
 a41403a <=( A266  and  (not A265) );
 a41406a <=( A268  and  A267 );
 a41407a <=( a41406a  and  a41403a );
 a41408a <=( a41407a  and  a41400a );
 a41412a <=( (not A168)  and  (not A169) );
 a41413a <=( A170  and  a41412a );
 a41416a <=( (not A166)  and  A167 );
 a41419a <=( (not A200)  and  (not A199) );
 a41420a <=( a41419a  and  a41416a );
 a41421a <=( a41420a  and  a41413a );
 a41424a <=( (not A233)  and  A232 );
 a41427a <=( A235  and  A234 );
 a41428a <=( a41427a  and  a41424a );
 a41431a <=( A266  and  (not A265) );
 a41434a <=( A269  and  A267 );
 a41435a <=( a41434a  and  a41431a );
 a41436a <=( a41435a  and  a41428a );
 a41440a <=( (not A168)  and  (not A169) );
 a41441a <=( A170  and  a41440a );
 a41444a <=( (not A166)  and  A167 );
 a41447a <=( (not A200)  and  (not A199) );
 a41448a <=( a41447a  and  a41444a );
 a41449a <=( a41448a  and  a41441a );
 a41452a <=( (not A233)  and  A232 );
 a41455a <=( A235  and  A234 );
 a41456a <=( a41455a  and  a41452a );
 a41459a <=( (not A266)  and  A265 );
 a41462a <=( A268  and  A267 );
 a41463a <=( a41462a  and  a41459a );
 a41464a <=( a41463a  and  a41456a );
 a41468a <=( (not A168)  and  (not A169) );
 a41469a <=( A170  and  a41468a );
 a41472a <=( (not A166)  and  A167 );
 a41475a <=( (not A200)  and  (not A199) );
 a41476a <=( a41475a  and  a41472a );
 a41477a <=( a41476a  and  a41469a );
 a41480a <=( (not A233)  and  A232 );
 a41483a <=( A235  and  A234 );
 a41484a <=( a41483a  and  a41480a );
 a41487a <=( (not A266)  and  A265 );
 a41490a <=( A269  and  A267 );
 a41491a <=( a41490a  and  a41487a );
 a41492a <=( a41491a  and  a41484a );
 a41496a <=( (not A168)  and  (not A169) );
 a41497a <=( A170  and  a41496a );
 a41500a <=( (not A166)  and  A167 );
 a41503a <=( (not A200)  and  (not A199) );
 a41504a <=( a41503a  and  a41500a );
 a41505a <=( a41504a  and  a41497a );
 a41508a <=( (not A233)  and  A232 );
 a41511a <=( A236  and  A234 );
 a41512a <=( a41511a  and  a41508a );
 a41515a <=( (not A299)  and  A298 );
 a41518a <=( A301  and  A300 );
 a41519a <=( a41518a  and  a41515a );
 a41520a <=( a41519a  and  a41512a );
 a41524a <=( (not A168)  and  (not A169) );
 a41525a <=( A170  and  a41524a );
 a41528a <=( (not A166)  and  A167 );
 a41531a <=( (not A200)  and  (not A199) );
 a41532a <=( a41531a  and  a41528a );
 a41533a <=( a41532a  and  a41525a );
 a41536a <=( (not A233)  and  A232 );
 a41539a <=( A236  and  A234 );
 a41540a <=( a41539a  and  a41536a );
 a41543a <=( (not A299)  and  A298 );
 a41546a <=( A302  and  A300 );
 a41547a <=( a41546a  and  a41543a );
 a41548a <=( a41547a  and  a41540a );
 a41552a <=( (not A168)  and  (not A169) );
 a41553a <=( A170  and  a41552a );
 a41556a <=( (not A166)  and  A167 );
 a41559a <=( (not A200)  and  (not A199) );
 a41560a <=( a41559a  and  a41556a );
 a41561a <=( a41560a  and  a41553a );
 a41564a <=( (not A233)  and  A232 );
 a41567a <=( A236  and  A234 );
 a41568a <=( a41567a  and  a41564a );
 a41571a <=( A299  and  (not A298) );
 a41574a <=( A301  and  A300 );
 a41575a <=( a41574a  and  a41571a );
 a41576a <=( a41575a  and  a41568a );
 a41580a <=( (not A168)  and  (not A169) );
 a41581a <=( A170  and  a41580a );
 a41584a <=( (not A166)  and  A167 );
 a41587a <=( (not A200)  and  (not A199) );
 a41588a <=( a41587a  and  a41584a );
 a41589a <=( a41588a  and  a41581a );
 a41592a <=( (not A233)  and  A232 );
 a41595a <=( A236  and  A234 );
 a41596a <=( a41595a  and  a41592a );
 a41599a <=( A299  and  (not A298) );
 a41602a <=( A302  and  A300 );
 a41603a <=( a41602a  and  a41599a );
 a41604a <=( a41603a  and  a41596a );
 a41608a <=( (not A168)  and  (not A169) );
 a41609a <=( A170  and  a41608a );
 a41612a <=( (not A166)  and  A167 );
 a41615a <=( (not A200)  and  (not A199) );
 a41616a <=( a41615a  and  a41612a );
 a41617a <=( a41616a  and  a41609a );
 a41620a <=( (not A233)  and  A232 );
 a41623a <=( A236  and  A234 );
 a41624a <=( a41623a  and  a41620a );
 a41627a <=( A266  and  (not A265) );
 a41630a <=( A268  and  A267 );
 a41631a <=( a41630a  and  a41627a );
 a41632a <=( a41631a  and  a41624a );
 a41636a <=( (not A168)  and  (not A169) );
 a41637a <=( A170  and  a41636a );
 a41640a <=( (not A166)  and  A167 );
 a41643a <=( (not A200)  and  (not A199) );
 a41644a <=( a41643a  and  a41640a );
 a41645a <=( a41644a  and  a41637a );
 a41648a <=( (not A233)  and  A232 );
 a41651a <=( A236  and  A234 );
 a41652a <=( a41651a  and  a41648a );
 a41655a <=( A266  and  (not A265) );
 a41658a <=( A269  and  A267 );
 a41659a <=( a41658a  and  a41655a );
 a41660a <=( a41659a  and  a41652a );
 a41664a <=( (not A168)  and  (not A169) );
 a41665a <=( A170  and  a41664a );
 a41668a <=( (not A166)  and  A167 );
 a41671a <=( (not A200)  and  (not A199) );
 a41672a <=( a41671a  and  a41668a );
 a41673a <=( a41672a  and  a41665a );
 a41676a <=( (not A233)  and  A232 );
 a41679a <=( A236  and  A234 );
 a41680a <=( a41679a  and  a41676a );
 a41683a <=( (not A266)  and  A265 );
 a41686a <=( A268  and  A267 );
 a41687a <=( a41686a  and  a41683a );
 a41688a <=( a41687a  and  a41680a );
 a41692a <=( (not A168)  and  (not A169) );
 a41693a <=( A170  and  a41692a );
 a41696a <=( (not A166)  and  A167 );
 a41699a <=( (not A200)  and  (not A199) );
 a41700a <=( a41699a  and  a41696a );
 a41701a <=( a41700a  and  a41693a );
 a41704a <=( (not A233)  and  A232 );
 a41707a <=( A236  and  A234 );
 a41708a <=( a41707a  and  a41704a );
 a41711a <=( (not A266)  and  A265 );
 a41714a <=( A269  and  A267 );
 a41715a <=( a41714a  and  a41711a );
 a41716a <=( a41715a  and  a41708a );
 a41720a <=( (not A168)  and  (not A169) );
 a41721a <=( A170  and  a41720a );
 a41724a <=( A166  and  (not A167) );
 a41727a <=( A202  and  (not A201) );
 a41728a <=( a41727a  and  a41724a );
 a41729a <=( a41728a  and  a41721a );
 a41732a <=( A233  and  (not A232) );
 a41735a <=( A235  and  A234 );
 a41736a <=( a41735a  and  a41732a );
 a41739a <=( (not A299)  and  A298 );
 a41742a <=( A301  and  A300 );
 a41743a <=( a41742a  and  a41739a );
 a41744a <=( a41743a  and  a41736a );
 a41748a <=( (not A168)  and  (not A169) );
 a41749a <=( A170  and  a41748a );
 a41752a <=( A166  and  (not A167) );
 a41755a <=( A202  and  (not A201) );
 a41756a <=( a41755a  and  a41752a );
 a41757a <=( a41756a  and  a41749a );
 a41760a <=( A233  and  (not A232) );
 a41763a <=( A235  and  A234 );
 a41764a <=( a41763a  and  a41760a );
 a41767a <=( (not A299)  and  A298 );
 a41770a <=( A302  and  A300 );
 a41771a <=( a41770a  and  a41767a );
 a41772a <=( a41771a  and  a41764a );
 a41776a <=( (not A168)  and  (not A169) );
 a41777a <=( A170  and  a41776a );
 a41780a <=( A166  and  (not A167) );
 a41783a <=( A202  and  (not A201) );
 a41784a <=( a41783a  and  a41780a );
 a41785a <=( a41784a  and  a41777a );
 a41788a <=( A233  and  (not A232) );
 a41791a <=( A235  and  A234 );
 a41792a <=( a41791a  and  a41788a );
 a41795a <=( A299  and  (not A298) );
 a41798a <=( A301  and  A300 );
 a41799a <=( a41798a  and  a41795a );
 a41800a <=( a41799a  and  a41792a );
 a41804a <=( (not A168)  and  (not A169) );
 a41805a <=( A170  and  a41804a );
 a41808a <=( A166  and  (not A167) );
 a41811a <=( A202  and  (not A201) );
 a41812a <=( a41811a  and  a41808a );
 a41813a <=( a41812a  and  a41805a );
 a41816a <=( A233  and  (not A232) );
 a41819a <=( A235  and  A234 );
 a41820a <=( a41819a  and  a41816a );
 a41823a <=( A299  and  (not A298) );
 a41826a <=( A302  and  A300 );
 a41827a <=( a41826a  and  a41823a );
 a41828a <=( a41827a  and  a41820a );
 a41832a <=( (not A168)  and  (not A169) );
 a41833a <=( A170  and  a41832a );
 a41836a <=( A166  and  (not A167) );
 a41839a <=( A202  and  (not A201) );
 a41840a <=( a41839a  and  a41836a );
 a41841a <=( a41840a  and  a41833a );
 a41844a <=( A233  and  (not A232) );
 a41847a <=( A235  and  A234 );
 a41848a <=( a41847a  and  a41844a );
 a41851a <=( A266  and  (not A265) );
 a41854a <=( A268  and  A267 );
 a41855a <=( a41854a  and  a41851a );
 a41856a <=( a41855a  and  a41848a );
 a41860a <=( (not A168)  and  (not A169) );
 a41861a <=( A170  and  a41860a );
 a41864a <=( A166  and  (not A167) );
 a41867a <=( A202  and  (not A201) );
 a41868a <=( a41867a  and  a41864a );
 a41869a <=( a41868a  and  a41861a );
 a41872a <=( A233  and  (not A232) );
 a41875a <=( A235  and  A234 );
 a41876a <=( a41875a  and  a41872a );
 a41879a <=( A266  and  (not A265) );
 a41882a <=( A269  and  A267 );
 a41883a <=( a41882a  and  a41879a );
 a41884a <=( a41883a  and  a41876a );
 a41888a <=( (not A168)  and  (not A169) );
 a41889a <=( A170  and  a41888a );
 a41892a <=( A166  and  (not A167) );
 a41895a <=( A202  and  (not A201) );
 a41896a <=( a41895a  and  a41892a );
 a41897a <=( a41896a  and  a41889a );
 a41900a <=( A233  and  (not A232) );
 a41903a <=( A235  and  A234 );
 a41904a <=( a41903a  and  a41900a );
 a41907a <=( (not A266)  and  A265 );
 a41910a <=( A268  and  A267 );
 a41911a <=( a41910a  and  a41907a );
 a41912a <=( a41911a  and  a41904a );
 a41916a <=( (not A168)  and  (not A169) );
 a41917a <=( A170  and  a41916a );
 a41920a <=( A166  and  (not A167) );
 a41923a <=( A202  and  (not A201) );
 a41924a <=( a41923a  and  a41920a );
 a41925a <=( a41924a  and  a41917a );
 a41928a <=( A233  and  (not A232) );
 a41931a <=( A235  and  A234 );
 a41932a <=( a41931a  and  a41928a );
 a41935a <=( (not A266)  and  A265 );
 a41938a <=( A269  and  A267 );
 a41939a <=( a41938a  and  a41935a );
 a41940a <=( a41939a  and  a41932a );
 a41944a <=( (not A168)  and  (not A169) );
 a41945a <=( A170  and  a41944a );
 a41948a <=( A166  and  (not A167) );
 a41951a <=( A202  and  (not A201) );
 a41952a <=( a41951a  and  a41948a );
 a41953a <=( a41952a  and  a41945a );
 a41956a <=( A233  and  (not A232) );
 a41959a <=( A236  and  A234 );
 a41960a <=( a41959a  and  a41956a );
 a41963a <=( (not A299)  and  A298 );
 a41966a <=( A301  and  A300 );
 a41967a <=( a41966a  and  a41963a );
 a41968a <=( a41967a  and  a41960a );
 a41972a <=( (not A168)  and  (not A169) );
 a41973a <=( A170  and  a41972a );
 a41976a <=( A166  and  (not A167) );
 a41979a <=( A202  and  (not A201) );
 a41980a <=( a41979a  and  a41976a );
 a41981a <=( a41980a  and  a41973a );
 a41984a <=( A233  and  (not A232) );
 a41987a <=( A236  and  A234 );
 a41988a <=( a41987a  and  a41984a );
 a41991a <=( (not A299)  and  A298 );
 a41994a <=( A302  and  A300 );
 a41995a <=( a41994a  and  a41991a );
 a41996a <=( a41995a  and  a41988a );
 a42000a <=( (not A168)  and  (not A169) );
 a42001a <=( A170  and  a42000a );
 a42004a <=( A166  and  (not A167) );
 a42007a <=( A202  and  (not A201) );
 a42008a <=( a42007a  and  a42004a );
 a42009a <=( a42008a  and  a42001a );
 a42012a <=( A233  and  (not A232) );
 a42015a <=( A236  and  A234 );
 a42016a <=( a42015a  and  a42012a );
 a42019a <=( A299  and  (not A298) );
 a42022a <=( A301  and  A300 );
 a42023a <=( a42022a  and  a42019a );
 a42024a <=( a42023a  and  a42016a );
 a42028a <=( (not A168)  and  (not A169) );
 a42029a <=( A170  and  a42028a );
 a42032a <=( A166  and  (not A167) );
 a42035a <=( A202  and  (not A201) );
 a42036a <=( a42035a  and  a42032a );
 a42037a <=( a42036a  and  a42029a );
 a42040a <=( A233  and  (not A232) );
 a42043a <=( A236  and  A234 );
 a42044a <=( a42043a  and  a42040a );
 a42047a <=( A299  and  (not A298) );
 a42050a <=( A302  and  A300 );
 a42051a <=( a42050a  and  a42047a );
 a42052a <=( a42051a  and  a42044a );
 a42056a <=( (not A168)  and  (not A169) );
 a42057a <=( A170  and  a42056a );
 a42060a <=( A166  and  (not A167) );
 a42063a <=( A202  and  (not A201) );
 a42064a <=( a42063a  and  a42060a );
 a42065a <=( a42064a  and  a42057a );
 a42068a <=( A233  and  (not A232) );
 a42071a <=( A236  and  A234 );
 a42072a <=( a42071a  and  a42068a );
 a42075a <=( A266  and  (not A265) );
 a42078a <=( A268  and  A267 );
 a42079a <=( a42078a  and  a42075a );
 a42080a <=( a42079a  and  a42072a );
 a42084a <=( (not A168)  and  (not A169) );
 a42085a <=( A170  and  a42084a );
 a42088a <=( A166  and  (not A167) );
 a42091a <=( A202  and  (not A201) );
 a42092a <=( a42091a  and  a42088a );
 a42093a <=( a42092a  and  a42085a );
 a42096a <=( A233  and  (not A232) );
 a42099a <=( A236  and  A234 );
 a42100a <=( a42099a  and  a42096a );
 a42103a <=( A266  and  (not A265) );
 a42106a <=( A269  and  A267 );
 a42107a <=( a42106a  and  a42103a );
 a42108a <=( a42107a  and  a42100a );
 a42112a <=( (not A168)  and  (not A169) );
 a42113a <=( A170  and  a42112a );
 a42116a <=( A166  and  (not A167) );
 a42119a <=( A202  and  (not A201) );
 a42120a <=( a42119a  and  a42116a );
 a42121a <=( a42120a  and  a42113a );
 a42124a <=( A233  and  (not A232) );
 a42127a <=( A236  and  A234 );
 a42128a <=( a42127a  and  a42124a );
 a42131a <=( (not A266)  and  A265 );
 a42134a <=( A268  and  A267 );
 a42135a <=( a42134a  and  a42131a );
 a42136a <=( a42135a  and  a42128a );
 a42140a <=( (not A168)  and  (not A169) );
 a42141a <=( A170  and  a42140a );
 a42144a <=( A166  and  (not A167) );
 a42147a <=( A202  and  (not A201) );
 a42148a <=( a42147a  and  a42144a );
 a42149a <=( a42148a  and  a42141a );
 a42152a <=( A233  and  (not A232) );
 a42155a <=( A236  and  A234 );
 a42156a <=( a42155a  and  a42152a );
 a42159a <=( (not A266)  and  A265 );
 a42162a <=( A269  and  A267 );
 a42163a <=( a42162a  and  a42159a );
 a42164a <=( a42163a  and  a42156a );
 a42168a <=( (not A168)  and  (not A169) );
 a42169a <=( A170  and  a42168a );
 a42172a <=( A166  and  (not A167) );
 a42175a <=( A202  and  (not A201) );
 a42176a <=( a42175a  and  a42172a );
 a42177a <=( a42176a  and  a42169a );
 a42180a <=( (not A233)  and  A232 );
 a42183a <=( A235  and  A234 );
 a42184a <=( a42183a  and  a42180a );
 a42187a <=( (not A299)  and  A298 );
 a42190a <=( A301  and  A300 );
 a42191a <=( a42190a  and  a42187a );
 a42192a <=( a42191a  and  a42184a );
 a42196a <=( (not A168)  and  (not A169) );
 a42197a <=( A170  and  a42196a );
 a42200a <=( A166  and  (not A167) );
 a42203a <=( A202  and  (not A201) );
 a42204a <=( a42203a  and  a42200a );
 a42205a <=( a42204a  and  a42197a );
 a42208a <=( (not A233)  and  A232 );
 a42211a <=( A235  and  A234 );
 a42212a <=( a42211a  and  a42208a );
 a42215a <=( (not A299)  and  A298 );
 a42218a <=( A302  and  A300 );
 a42219a <=( a42218a  and  a42215a );
 a42220a <=( a42219a  and  a42212a );
 a42224a <=( (not A168)  and  (not A169) );
 a42225a <=( A170  and  a42224a );
 a42228a <=( A166  and  (not A167) );
 a42231a <=( A202  and  (not A201) );
 a42232a <=( a42231a  and  a42228a );
 a42233a <=( a42232a  and  a42225a );
 a42236a <=( (not A233)  and  A232 );
 a42239a <=( A235  and  A234 );
 a42240a <=( a42239a  and  a42236a );
 a42243a <=( A299  and  (not A298) );
 a42246a <=( A301  and  A300 );
 a42247a <=( a42246a  and  a42243a );
 a42248a <=( a42247a  and  a42240a );
 a42252a <=( (not A168)  and  (not A169) );
 a42253a <=( A170  and  a42252a );
 a42256a <=( A166  and  (not A167) );
 a42259a <=( A202  and  (not A201) );
 a42260a <=( a42259a  and  a42256a );
 a42261a <=( a42260a  and  a42253a );
 a42264a <=( (not A233)  and  A232 );
 a42267a <=( A235  and  A234 );
 a42268a <=( a42267a  and  a42264a );
 a42271a <=( A299  and  (not A298) );
 a42274a <=( A302  and  A300 );
 a42275a <=( a42274a  and  a42271a );
 a42276a <=( a42275a  and  a42268a );
 a42280a <=( (not A168)  and  (not A169) );
 a42281a <=( A170  and  a42280a );
 a42284a <=( A166  and  (not A167) );
 a42287a <=( A202  and  (not A201) );
 a42288a <=( a42287a  and  a42284a );
 a42289a <=( a42288a  and  a42281a );
 a42292a <=( (not A233)  and  A232 );
 a42295a <=( A235  and  A234 );
 a42296a <=( a42295a  and  a42292a );
 a42299a <=( A266  and  (not A265) );
 a42302a <=( A268  and  A267 );
 a42303a <=( a42302a  and  a42299a );
 a42304a <=( a42303a  and  a42296a );
 a42308a <=( (not A168)  and  (not A169) );
 a42309a <=( A170  and  a42308a );
 a42312a <=( A166  and  (not A167) );
 a42315a <=( A202  and  (not A201) );
 a42316a <=( a42315a  and  a42312a );
 a42317a <=( a42316a  and  a42309a );
 a42320a <=( (not A233)  and  A232 );
 a42323a <=( A235  and  A234 );
 a42324a <=( a42323a  and  a42320a );
 a42327a <=( A266  and  (not A265) );
 a42330a <=( A269  and  A267 );
 a42331a <=( a42330a  and  a42327a );
 a42332a <=( a42331a  and  a42324a );
 a42336a <=( (not A168)  and  (not A169) );
 a42337a <=( A170  and  a42336a );
 a42340a <=( A166  and  (not A167) );
 a42343a <=( A202  and  (not A201) );
 a42344a <=( a42343a  and  a42340a );
 a42345a <=( a42344a  and  a42337a );
 a42348a <=( (not A233)  and  A232 );
 a42351a <=( A235  and  A234 );
 a42352a <=( a42351a  and  a42348a );
 a42355a <=( (not A266)  and  A265 );
 a42358a <=( A268  and  A267 );
 a42359a <=( a42358a  and  a42355a );
 a42360a <=( a42359a  and  a42352a );
 a42364a <=( (not A168)  and  (not A169) );
 a42365a <=( A170  and  a42364a );
 a42368a <=( A166  and  (not A167) );
 a42371a <=( A202  and  (not A201) );
 a42372a <=( a42371a  and  a42368a );
 a42373a <=( a42372a  and  a42365a );
 a42376a <=( (not A233)  and  A232 );
 a42379a <=( A235  and  A234 );
 a42380a <=( a42379a  and  a42376a );
 a42383a <=( (not A266)  and  A265 );
 a42386a <=( A269  and  A267 );
 a42387a <=( a42386a  and  a42383a );
 a42388a <=( a42387a  and  a42380a );
 a42392a <=( (not A168)  and  (not A169) );
 a42393a <=( A170  and  a42392a );
 a42396a <=( A166  and  (not A167) );
 a42399a <=( A202  and  (not A201) );
 a42400a <=( a42399a  and  a42396a );
 a42401a <=( a42400a  and  a42393a );
 a42404a <=( (not A233)  and  A232 );
 a42407a <=( A236  and  A234 );
 a42408a <=( a42407a  and  a42404a );
 a42411a <=( (not A299)  and  A298 );
 a42414a <=( A301  and  A300 );
 a42415a <=( a42414a  and  a42411a );
 a42416a <=( a42415a  and  a42408a );
 a42420a <=( (not A168)  and  (not A169) );
 a42421a <=( A170  and  a42420a );
 a42424a <=( A166  and  (not A167) );
 a42427a <=( A202  and  (not A201) );
 a42428a <=( a42427a  and  a42424a );
 a42429a <=( a42428a  and  a42421a );
 a42432a <=( (not A233)  and  A232 );
 a42435a <=( A236  and  A234 );
 a42436a <=( a42435a  and  a42432a );
 a42439a <=( (not A299)  and  A298 );
 a42442a <=( A302  and  A300 );
 a42443a <=( a42442a  and  a42439a );
 a42444a <=( a42443a  and  a42436a );
 a42448a <=( (not A168)  and  (not A169) );
 a42449a <=( A170  and  a42448a );
 a42452a <=( A166  and  (not A167) );
 a42455a <=( A202  and  (not A201) );
 a42456a <=( a42455a  and  a42452a );
 a42457a <=( a42456a  and  a42449a );
 a42460a <=( (not A233)  and  A232 );
 a42463a <=( A236  and  A234 );
 a42464a <=( a42463a  and  a42460a );
 a42467a <=( A299  and  (not A298) );
 a42470a <=( A301  and  A300 );
 a42471a <=( a42470a  and  a42467a );
 a42472a <=( a42471a  and  a42464a );
 a42476a <=( (not A168)  and  (not A169) );
 a42477a <=( A170  and  a42476a );
 a42480a <=( A166  and  (not A167) );
 a42483a <=( A202  and  (not A201) );
 a42484a <=( a42483a  and  a42480a );
 a42485a <=( a42484a  and  a42477a );
 a42488a <=( (not A233)  and  A232 );
 a42491a <=( A236  and  A234 );
 a42492a <=( a42491a  and  a42488a );
 a42495a <=( A299  and  (not A298) );
 a42498a <=( A302  and  A300 );
 a42499a <=( a42498a  and  a42495a );
 a42500a <=( a42499a  and  a42492a );
 a42504a <=( (not A168)  and  (not A169) );
 a42505a <=( A170  and  a42504a );
 a42508a <=( A166  and  (not A167) );
 a42511a <=( A202  and  (not A201) );
 a42512a <=( a42511a  and  a42508a );
 a42513a <=( a42512a  and  a42505a );
 a42516a <=( (not A233)  and  A232 );
 a42519a <=( A236  and  A234 );
 a42520a <=( a42519a  and  a42516a );
 a42523a <=( A266  and  (not A265) );
 a42526a <=( A268  and  A267 );
 a42527a <=( a42526a  and  a42523a );
 a42528a <=( a42527a  and  a42520a );
 a42532a <=( (not A168)  and  (not A169) );
 a42533a <=( A170  and  a42532a );
 a42536a <=( A166  and  (not A167) );
 a42539a <=( A202  and  (not A201) );
 a42540a <=( a42539a  and  a42536a );
 a42541a <=( a42540a  and  a42533a );
 a42544a <=( (not A233)  and  A232 );
 a42547a <=( A236  and  A234 );
 a42548a <=( a42547a  and  a42544a );
 a42551a <=( A266  and  (not A265) );
 a42554a <=( A269  and  A267 );
 a42555a <=( a42554a  and  a42551a );
 a42556a <=( a42555a  and  a42548a );
 a42560a <=( (not A168)  and  (not A169) );
 a42561a <=( A170  and  a42560a );
 a42564a <=( A166  and  (not A167) );
 a42567a <=( A202  and  (not A201) );
 a42568a <=( a42567a  and  a42564a );
 a42569a <=( a42568a  and  a42561a );
 a42572a <=( (not A233)  and  A232 );
 a42575a <=( A236  and  A234 );
 a42576a <=( a42575a  and  a42572a );
 a42579a <=( (not A266)  and  A265 );
 a42582a <=( A268  and  A267 );
 a42583a <=( a42582a  and  a42579a );
 a42584a <=( a42583a  and  a42576a );
 a42588a <=( (not A168)  and  (not A169) );
 a42589a <=( A170  and  a42588a );
 a42592a <=( A166  and  (not A167) );
 a42595a <=( A202  and  (not A201) );
 a42596a <=( a42595a  and  a42592a );
 a42597a <=( a42596a  and  a42589a );
 a42600a <=( (not A233)  and  A232 );
 a42603a <=( A236  and  A234 );
 a42604a <=( a42603a  and  a42600a );
 a42607a <=( (not A266)  and  A265 );
 a42610a <=( A269  and  A267 );
 a42611a <=( a42610a  and  a42607a );
 a42612a <=( a42611a  and  a42604a );
 a42616a <=( (not A168)  and  (not A169) );
 a42617a <=( A170  and  a42616a );
 a42620a <=( A166  and  (not A167) );
 a42623a <=( A203  and  (not A201) );
 a42624a <=( a42623a  and  a42620a );
 a42625a <=( a42624a  and  a42617a );
 a42628a <=( A233  and  (not A232) );
 a42631a <=( A235  and  A234 );
 a42632a <=( a42631a  and  a42628a );
 a42635a <=( (not A299)  and  A298 );
 a42638a <=( A301  and  A300 );
 a42639a <=( a42638a  and  a42635a );
 a42640a <=( a42639a  and  a42632a );
 a42644a <=( (not A168)  and  (not A169) );
 a42645a <=( A170  and  a42644a );
 a42648a <=( A166  and  (not A167) );
 a42651a <=( A203  and  (not A201) );
 a42652a <=( a42651a  and  a42648a );
 a42653a <=( a42652a  and  a42645a );
 a42656a <=( A233  and  (not A232) );
 a42659a <=( A235  and  A234 );
 a42660a <=( a42659a  and  a42656a );
 a42663a <=( (not A299)  and  A298 );
 a42666a <=( A302  and  A300 );
 a42667a <=( a42666a  and  a42663a );
 a42668a <=( a42667a  and  a42660a );
 a42672a <=( (not A168)  and  (not A169) );
 a42673a <=( A170  and  a42672a );
 a42676a <=( A166  and  (not A167) );
 a42679a <=( A203  and  (not A201) );
 a42680a <=( a42679a  and  a42676a );
 a42681a <=( a42680a  and  a42673a );
 a42684a <=( A233  and  (not A232) );
 a42687a <=( A235  and  A234 );
 a42688a <=( a42687a  and  a42684a );
 a42691a <=( A299  and  (not A298) );
 a42694a <=( A301  and  A300 );
 a42695a <=( a42694a  and  a42691a );
 a42696a <=( a42695a  and  a42688a );
 a42700a <=( (not A168)  and  (not A169) );
 a42701a <=( A170  and  a42700a );
 a42704a <=( A166  and  (not A167) );
 a42707a <=( A203  and  (not A201) );
 a42708a <=( a42707a  and  a42704a );
 a42709a <=( a42708a  and  a42701a );
 a42712a <=( A233  and  (not A232) );
 a42715a <=( A235  and  A234 );
 a42716a <=( a42715a  and  a42712a );
 a42719a <=( A299  and  (not A298) );
 a42722a <=( A302  and  A300 );
 a42723a <=( a42722a  and  a42719a );
 a42724a <=( a42723a  and  a42716a );
 a42728a <=( (not A168)  and  (not A169) );
 a42729a <=( A170  and  a42728a );
 a42732a <=( A166  and  (not A167) );
 a42735a <=( A203  and  (not A201) );
 a42736a <=( a42735a  and  a42732a );
 a42737a <=( a42736a  and  a42729a );
 a42740a <=( A233  and  (not A232) );
 a42743a <=( A235  and  A234 );
 a42744a <=( a42743a  and  a42740a );
 a42747a <=( A266  and  (not A265) );
 a42750a <=( A268  and  A267 );
 a42751a <=( a42750a  and  a42747a );
 a42752a <=( a42751a  and  a42744a );
 a42756a <=( (not A168)  and  (not A169) );
 a42757a <=( A170  and  a42756a );
 a42760a <=( A166  and  (not A167) );
 a42763a <=( A203  and  (not A201) );
 a42764a <=( a42763a  and  a42760a );
 a42765a <=( a42764a  and  a42757a );
 a42768a <=( A233  and  (not A232) );
 a42771a <=( A235  and  A234 );
 a42772a <=( a42771a  and  a42768a );
 a42775a <=( A266  and  (not A265) );
 a42778a <=( A269  and  A267 );
 a42779a <=( a42778a  and  a42775a );
 a42780a <=( a42779a  and  a42772a );
 a42784a <=( (not A168)  and  (not A169) );
 a42785a <=( A170  and  a42784a );
 a42788a <=( A166  and  (not A167) );
 a42791a <=( A203  and  (not A201) );
 a42792a <=( a42791a  and  a42788a );
 a42793a <=( a42792a  and  a42785a );
 a42796a <=( A233  and  (not A232) );
 a42799a <=( A235  and  A234 );
 a42800a <=( a42799a  and  a42796a );
 a42803a <=( (not A266)  and  A265 );
 a42806a <=( A268  and  A267 );
 a42807a <=( a42806a  and  a42803a );
 a42808a <=( a42807a  and  a42800a );
 a42812a <=( (not A168)  and  (not A169) );
 a42813a <=( A170  and  a42812a );
 a42816a <=( A166  and  (not A167) );
 a42819a <=( A203  and  (not A201) );
 a42820a <=( a42819a  and  a42816a );
 a42821a <=( a42820a  and  a42813a );
 a42824a <=( A233  and  (not A232) );
 a42827a <=( A235  and  A234 );
 a42828a <=( a42827a  and  a42824a );
 a42831a <=( (not A266)  and  A265 );
 a42834a <=( A269  and  A267 );
 a42835a <=( a42834a  and  a42831a );
 a42836a <=( a42835a  and  a42828a );
 a42840a <=( (not A168)  and  (not A169) );
 a42841a <=( A170  and  a42840a );
 a42844a <=( A166  and  (not A167) );
 a42847a <=( A203  and  (not A201) );
 a42848a <=( a42847a  and  a42844a );
 a42849a <=( a42848a  and  a42841a );
 a42852a <=( A233  and  (not A232) );
 a42855a <=( A236  and  A234 );
 a42856a <=( a42855a  and  a42852a );
 a42859a <=( (not A299)  and  A298 );
 a42862a <=( A301  and  A300 );
 a42863a <=( a42862a  and  a42859a );
 a42864a <=( a42863a  and  a42856a );
 a42868a <=( (not A168)  and  (not A169) );
 a42869a <=( A170  and  a42868a );
 a42872a <=( A166  and  (not A167) );
 a42875a <=( A203  and  (not A201) );
 a42876a <=( a42875a  and  a42872a );
 a42877a <=( a42876a  and  a42869a );
 a42880a <=( A233  and  (not A232) );
 a42883a <=( A236  and  A234 );
 a42884a <=( a42883a  and  a42880a );
 a42887a <=( (not A299)  and  A298 );
 a42890a <=( A302  and  A300 );
 a42891a <=( a42890a  and  a42887a );
 a42892a <=( a42891a  and  a42884a );
 a42896a <=( (not A168)  and  (not A169) );
 a42897a <=( A170  and  a42896a );
 a42900a <=( A166  and  (not A167) );
 a42903a <=( A203  and  (not A201) );
 a42904a <=( a42903a  and  a42900a );
 a42905a <=( a42904a  and  a42897a );
 a42908a <=( A233  and  (not A232) );
 a42911a <=( A236  and  A234 );
 a42912a <=( a42911a  and  a42908a );
 a42915a <=( A299  and  (not A298) );
 a42918a <=( A301  and  A300 );
 a42919a <=( a42918a  and  a42915a );
 a42920a <=( a42919a  and  a42912a );
 a42924a <=( (not A168)  and  (not A169) );
 a42925a <=( A170  and  a42924a );
 a42928a <=( A166  and  (not A167) );
 a42931a <=( A203  and  (not A201) );
 a42932a <=( a42931a  and  a42928a );
 a42933a <=( a42932a  and  a42925a );
 a42936a <=( A233  and  (not A232) );
 a42939a <=( A236  and  A234 );
 a42940a <=( a42939a  and  a42936a );
 a42943a <=( A299  and  (not A298) );
 a42946a <=( A302  and  A300 );
 a42947a <=( a42946a  and  a42943a );
 a42948a <=( a42947a  and  a42940a );
 a42952a <=( (not A168)  and  (not A169) );
 a42953a <=( A170  and  a42952a );
 a42956a <=( A166  and  (not A167) );
 a42959a <=( A203  and  (not A201) );
 a42960a <=( a42959a  and  a42956a );
 a42961a <=( a42960a  and  a42953a );
 a42964a <=( A233  and  (not A232) );
 a42967a <=( A236  and  A234 );
 a42968a <=( a42967a  and  a42964a );
 a42971a <=( A266  and  (not A265) );
 a42974a <=( A268  and  A267 );
 a42975a <=( a42974a  and  a42971a );
 a42976a <=( a42975a  and  a42968a );
 a42980a <=( (not A168)  and  (not A169) );
 a42981a <=( A170  and  a42980a );
 a42984a <=( A166  and  (not A167) );
 a42987a <=( A203  and  (not A201) );
 a42988a <=( a42987a  and  a42984a );
 a42989a <=( a42988a  and  a42981a );
 a42992a <=( A233  and  (not A232) );
 a42995a <=( A236  and  A234 );
 a42996a <=( a42995a  and  a42992a );
 a42999a <=( A266  and  (not A265) );
 a43002a <=( A269  and  A267 );
 a43003a <=( a43002a  and  a42999a );
 a43004a <=( a43003a  and  a42996a );
 a43008a <=( (not A168)  and  (not A169) );
 a43009a <=( A170  and  a43008a );
 a43012a <=( A166  and  (not A167) );
 a43015a <=( A203  and  (not A201) );
 a43016a <=( a43015a  and  a43012a );
 a43017a <=( a43016a  and  a43009a );
 a43020a <=( A233  and  (not A232) );
 a43023a <=( A236  and  A234 );
 a43024a <=( a43023a  and  a43020a );
 a43027a <=( (not A266)  and  A265 );
 a43030a <=( A268  and  A267 );
 a43031a <=( a43030a  and  a43027a );
 a43032a <=( a43031a  and  a43024a );
 a43036a <=( (not A168)  and  (not A169) );
 a43037a <=( A170  and  a43036a );
 a43040a <=( A166  and  (not A167) );
 a43043a <=( A203  and  (not A201) );
 a43044a <=( a43043a  and  a43040a );
 a43045a <=( a43044a  and  a43037a );
 a43048a <=( A233  and  (not A232) );
 a43051a <=( A236  and  A234 );
 a43052a <=( a43051a  and  a43048a );
 a43055a <=( (not A266)  and  A265 );
 a43058a <=( A269  and  A267 );
 a43059a <=( a43058a  and  a43055a );
 a43060a <=( a43059a  and  a43052a );
 a43064a <=( (not A168)  and  (not A169) );
 a43065a <=( A170  and  a43064a );
 a43068a <=( A166  and  (not A167) );
 a43071a <=( A203  and  (not A201) );
 a43072a <=( a43071a  and  a43068a );
 a43073a <=( a43072a  and  a43065a );
 a43076a <=( (not A233)  and  A232 );
 a43079a <=( A235  and  A234 );
 a43080a <=( a43079a  and  a43076a );
 a43083a <=( (not A299)  and  A298 );
 a43086a <=( A301  and  A300 );
 a43087a <=( a43086a  and  a43083a );
 a43088a <=( a43087a  and  a43080a );
 a43092a <=( (not A168)  and  (not A169) );
 a43093a <=( A170  and  a43092a );
 a43096a <=( A166  and  (not A167) );
 a43099a <=( A203  and  (not A201) );
 a43100a <=( a43099a  and  a43096a );
 a43101a <=( a43100a  and  a43093a );
 a43104a <=( (not A233)  and  A232 );
 a43107a <=( A235  and  A234 );
 a43108a <=( a43107a  and  a43104a );
 a43111a <=( (not A299)  and  A298 );
 a43114a <=( A302  and  A300 );
 a43115a <=( a43114a  and  a43111a );
 a43116a <=( a43115a  and  a43108a );
 a43120a <=( (not A168)  and  (not A169) );
 a43121a <=( A170  and  a43120a );
 a43124a <=( A166  and  (not A167) );
 a43127a <=( A203  and  (not A201) );
 a43128a <=( a43127a  and  a43124a );
 a43129a <=( a43128a  and  a43121a );
 a43132a <=( (not A233)  and  A232 );
 a43135a <=( A235  and  A234 );
 a43136a <=( a43135a  and  a43132a );
 a43139a <=( A299  and  (not A298) );
 a43142a <=( A301  and  A300 );
 a43143a <=( a43142a  and  a43139a );
 a43144a <=( a43143a  and  a43136a );
 a43148a <=( (not A168)  and  (not A169) );
 a43149a <=( A170  and  a43148a );
 a43152a <=( A166  and  (not A167) );
 a43155a <=( A203  and  (not A201) );
 a43156a <=( a43155a  and  a43152a );
 a43157a <=( a43156a  and  a43149a );
 a43160a <=( (not A233)  and  A232 );
 a43163a <=( A235  and  A234 );
 a43164a <=( a43163a  and  a43160a );
 a43167a <=( A299  and  (not A298) );
 a43170a <=( A302  and  A300 );
 a43171a <=( a43170a  and  a43167a );
 a43172a <=( a43171a  and  a43164a );
 a43176a <=( (not A168)  and  (not A169) );
 a43177a <=( A170  and  a43176a );
 a43180a <=( A166  and  (not A167) );
 a43183a <=( A203  and  (not A201) );
 a43184a <=( a43183a  and  a43180a );
 a43185a <=( a43184a  and  a43177a );
 a43188a <=( (not A233)  and  A232 );
 a43191a <=( A235  and  A234 );
 a43192a <=( a43191a  and  a43188a );
 a43195a <=( A266  and  (not A265) );
 a43198a <=( A268  and  A267 );
 a43199a <=( a43198a  and  a43195a );
 a43200a <=( a43199a  and  a43192a );
 a43204a <=( (not A168)  and  (not A169) );
 a43205a <=( A170  and  a43204a );
 a43208a <=( A166  and  (not A167) );
 a43211a <=( A203  and  (not A201) );
 a43212a <=( a43211a  and  a43208a );
 a43213a <=( a43212a  and  a43205a );
 a43216a <=( (not A233)  and  A232 );
 a43219a <=( A235  and  A234 );
 a43220a <=( a43219a  and  a43216a );
 a43223a <=( A266  and  (not A265) );
 a43226a <=( A269  and  A267 );
 a43227a <=( a43226a  and  a43223a );
 a43228a <=( a43227a  and  a43220a );
 a43232a <=( (not A168)  and  (not A169) );
 a43233a <=( A170  and  a43232a );
 a43236a <=( A166  and  (not A167) );
 a43239a <=( A203  and  (not A201) );
 a43240a <=( a43239a  and  a43236a );
 a43241a <=( a43240a  and  a43233a );
 a43244a <=( (not A233)  and  A232 );
 a43247a <=( A235  and  A234 );
 a43248a <=( a43247a  and  a43244a );
 a43251a <=( (not A266)  and  A265 );
 a43254a <=( A268  and  A267 );
 a43255a <=( a43254a  and  a43251a );
 a43256a <=( a43255a  and  a43248a );
 a43260a <=( (not A168)  and  (not A169) );
 a43261a <=( A170  and  a43260a );
 a43264a <=( A166  and  (not A167) );
 a43267a <=( A203  and  (not A201) );
 a43268a <=( a43267a  and  a43264a );
 a43269a <=( a43268a  and  a43261a );
 a43272a <=( (not A233)  and  A232 );
 a43275a <=( A235  and  A234 );
 a43276a <=( a43275a  and  a43272a );
 a43279a <=( (not A266)  and  A265 );
 a43282a <=( A269  and  A267 );
 a43283a <=( a43282a  and  a43279a );
 a43284a <=( a43283a  and  a43276a );
 a43288a <=( (not A168)  and  (not A169) );
 a43289a <=( A170  and  a43288a );
 a43292a <=( A166  and  (not A167) );
 a43295a <=( A203  and  (not A201) );
 a43296a <=( a43295a  and  a43292a );
 a43297a <=( a43296a  and  a43289a );
 a43300a <=( (not A233)  and  A232 );
 a43303a <=( A236  and  A234 );
 a43304a <=( a43303a  and  a43300a );
 a43307a <=( (not A299)  and  A298 );
 a43310a <=( A301  and  A300 );
 a43311a <=( a43310a  and  a43307a );
 a43312a <=( a43311a  and  a43304a );
 a43316a <=( (not A168)  and  (not A169) );
 a43317a <=( A170  and  a43316a );
 a43320a <=( A166  and  (not A167) );
 a43323a <=( A203  and  (not A201) );
 a43324a <=( a43323a  and  a43320a );
 a43325a <=( a43324a  and  a43317a );
 a43328a <=( (not A233)  and  A232 );
 a43331a <=( A236  and  A234 );
 a43332a <=( a43331a  and  a43328a );
 a43335a <=( (not A299)  and  A298 );
 a43338a <=( A302  and  A300 );
 a43339a <=( a43338a  and  a43335a );
 a43340a <=( a43339a  and  a43332a );
 a43344a <=( (not A168)  and  (not A169) );
 a43345a <=( A170  and  a43344a );
 a43348a <=( A166  and  (not A167) );
 a43351a <=( A203  and  (not A201) );
 a43352a <=( a43351a  and  a43348a );
 a43353a <=( a43352a  and  a43345a );
 a43356a <=( (not A233)  and  A232 );
 a43359a <=( A236  and  A234 );
 a43360a <=( a43359a  and  a43356a );
 a43363a <=( A299  and  (not A298) );
 a43366a <=( A301  and  A300 );
 a43367a <=( a43366a  and  a43363a );
 a43368a <=( a43367a  and  a43360a );
 a43372a <=( (not A168)  and  (not A169) );
 a43373a <=( A170  and  a43372a );
 a43376a <=( A166  and  (not A167) );
 a43379a <=( A203  and  (not A201) );
 a43380a <=( a43379a  and  a43376a );
 a43381a <=( a43380a  and  a43373a );
 a43384a <=( (not A233)  and  A232 );
 a43387a <=( A236  and  A234 );
 a43388a <=( a43387a  and  a43384a );
 a43391a <=( A299  and  (not A298) );
 a43394a <=( A302  and  A300 );
 a43395a <=( a43394a  and  a43391a );
 a43396a <=( a43395a  and  a43388a );
 a43400a <=( (not A168)  and  (not A169) );
 a43401a <=( A170  and  a43400a );
 a43404a <=( A166  and  (not A167) );
 a43407a <=( A203  and  (not A201) );
 a43408a <=( a43407a  and  a43404a );
 a43409a <=( a43408a  and  a43401a );
 a43412a <=( (not A233)  and  A232 );
 a43415a <=( A236  and  A234 );
 a43416a <=( a43415a  and  a43412a );
 a43419a <=( A266  and  (not A265) );
 a43422a <=( A268  and  A267 );
 a43423a <=( a43422a  and  a43419a );
 a43424a <=( a43423a  and  a43416a );
 a43428a <=( (not A168)  and  (not A169) );
 a43429a <=( A170  and  a43428a );
 a43432a <=( A166  and  (not A167) );
 a43435a <=( A203  and  (not A201) );
 a43436a <=( a43435a  and  a43432a );
 a43437a <=( a43436a  and  a43429a );
 a43440a <=( (not A233)  and  A232 );
 a43443a <=( A236  and  A234 );
 a43444a <=( a43443a  and  a43440a );
 a43447a <=( A266  and  (not A265) );
 a43450a <=( A269  and  A267 );
 a43451a <=( a43450a  and  a43447a );
 a43452a <=( a43451a  and  a43444a );
 a43456a <=( (not A168)  and  (not A169) );
 a43457a <=( A170  and  a43456a );
 a43460a <=( A166  and  (not A167) );
 a43463a <=( A203  and  (not A201) );
 a43464a <=( a43463a  and  a43460a );
 a43465a <=( a43464a  and  a43457a );
 a43468a <=( (not A233)  and  A232 );
 a43471a <=( A236  and  A234 );
 a43472a <=( a43471a  and  a43468a );
 a43475a <=( (not A266)  and  A265 );
 a43478a <=( A268  and  A267 );
 a43479a <=( a43478a  and  a43475a );
 a43480a <=( a43479a  and  a43472a );
 a43484a <=( (not A168)  and  (not A169) );
 a43485a <=( A170  and  a43484a );
 a43488a <=( A166  and  (not A167) );
 a43491a <=( A203  and  (not A201) );
 a43492a <=( a43491a  and  a43488a );
 a43493a <=( a43492a  and  a43485a );
 a43496a <=( (not A233)  and  A232 );
 a43499a <=( A236  and  A234 );
 a43500a <=( a43499a  and  a43496a );
 a43503a <=( (not A266)  and  A265 );
 a43506a <=( A269  and  A267 );
 a43507a <=( a43506a  and  a43503a );
 a43508a <=( a43507a  and  a43500a );
 a43512a <=( (not A168)  and  (not A169) );
 a43513a <=( A170  and  a43512a );
 a43516a <=( A166  and  (not A167) );
 a43519a <=( A200  and  A199 );
 a43520a <=( a43519a  and  a43516a );
 a43521a <=( a43520a  and  a43513a );
 a43524a <=( A233  and  (not A232) );
 a43527a <=( A235  and  A234 );
 a43528a <=( a43527a  and  a43524a );
 a43531a <=( (not A299)  and  A298 );
 a43534a <=( A301  and  A300 );
 a43535a <=( a43534a  and  a43531a );
 a43536a <=( a43535a  and  a43528a );
 a43540a <=( (not A168)  and  (not A169) );
 a43541a <=( A170  and  a43540a );
 a43544a <=( A166  and  (not A167) );
 a43547a <=( A200  and  A199 );
 a43548a <=( a43547a  and  a43544a );
 a43549a <=( a43548a  and  a43541a );
 a43552a <=( A233  and  (not A232) );
 a43555a <=( A235  and  A234 );
 a43556a <=( a43555a  and  a43552a );
 a43559a <=( (not A299)  and  A298 );
 a43562a <=( A302  and  A300 );
 a43563a <=( a43562a  and  a43559a );
 a43564a <=( a43563a  and  a43556a );
 a43568a <=( (not A168)  and  (not A169) );
 a43569a <=( A170  and  a43568a );
 a43572a <=( A166  and  (not A167) );
 a43575a <=( A200  and  A199 );
 a43576a <=( a43575a  and  a43572a );
 a43577a <=( a43576a  and  a43569a );
 a43580a <=( A233  and  (not A232) );
 a43583a <=( A235  and  A234 );
 a43584a <=( a43583a  and  a43580a );
 a43587a <=( A299  and  (not A298) );
 a43590a <=( A301  and  A300 );
 a43591a <=( a43590a  and  a43587a );
 a43592a <=( a43591a  and  a43584a );
 a43596a <=( (not A168)  and  (not A169) );
 a43597a <=( A170  and  a43596a );
 a43600a <=( A166  and  (not A167) );
 a43603a <=( A200  and  A199 );
 a43604a <=( a43603a  and  a43600a );
 a43605a <=( a43604a  and  a43597a );
 a43608a <=( A233  and  (not A232) );
 a43611a <=( A235  and  A234 );
 a43612a <=( a43611a  and  a43608a );
 a43615a <=( A299  and  (not A298) );
 a43618a <=( A302  and  A300 );
 a43619a <=( a43618a  and  a43615a );
 a43620a <=( a43619a  and  a43612a );
 a43624a <=( (not A168)  and  (not A169) );
 a43625a <=( A170  and  a43624a );
 a43628a <=( A166  and  (not A167) );
 a43631a <=( A200  and  A199 );
 a43632a <=( a43631a  and  a43628a );
 a43633a <=( a43632a  and  a43625a );
 a43636a <=( A233  and  (not A232) );
 a43639a <=( A235  and  A234 );
 a43640a <=( a43639a  and  a43636a );
 a43643a <=( A266  and  (not A265) );
 a43646a <=( A268  and  A267 );
 a43647a <=( a43646a  and  a43643a );
 a43648a <=( a43647a  and  a43640a );
 a43652a <=( (not A168)  and  (not A169) );
 a43653a <=( A170  and  a43652a );
 a43656a <=( A166  and  (not A167) );
 a43659a <=( A200  and  A199 );
 a43660a <=( a43659a  and  a43656a );
 a43661a <=( a43660a  and  a43653a );
 a43664a <=( A233  and  (not A232) );
 a43667a <=( A235  and  A234 );
 a43668a <=( a43667a  and  a43664a );
 a43671a <=( A266  and  (not A265) );
 a43674a <=( A269  and  A267 );
 a43675a <=( a43674a  and  a43671a );
 a43676a <=( a43675a  and  a43668a );
 a43680a <=( (not A168)  and  (not A169) );
 a43681a <=( A170  and  a43680a );
 a43684a <=( A166  and  (not A167) );
 a43687a <=( A200  and  A199 );
 a43688a <=( a43687a  and  a43684a );
 a43689a <=( a43688a  and  a43681a );
 a43692a <=( A233  and  (not A232) );
 a43695a <=( A235  and  A234 );
 a43696a <=( a43695a  and  a43692a );
 a43699a <=( (not A266)  and  A265 );
 a43702a <=( A268  and  A267 );
 a43703a <=( a43702a  and  a43699a );
 a43704a <=( a43703a  and  a43696a );
 a43708a <=( (not A168)  and  (not A169) );
 a43709a <=( A170  and  a43708a );
 a43712a <=( A166  and  (not A167) );
 a43715a <=( A200  and  A199 );
 a43716a <=( a43715a  and  a43712a );
 a43717a <=( a43716a  and  a43709a );
 a43720a <=( A233  and  (not A232) );
 a43723a <=( A235  and  A234 );
 a43724a <=( a43723a  and  a43720a );
 a43727a <=( (not A266)  and  A265 );
 a43730a <=( A269  and  A267 );
 a43731a <=( a43730a  and  a43727a );
 a43732a <=( a43731a  and  a43724a );
 a43736a <=( (not A168)  and  (not A169) );
 a43737a <=( A170  and  a43736a );
 a43740a <=( A166  and  (not A167) );
 a43743a <=( A200  and  A199 );
 a43744a <=( a43743a  and  a43740a );
 a43745a <=( a43744a  and  a43737a );
 a43748a <=( A233  and  (not A232) );
 a43751a <=( A236  and  A234 );
 a43752a <=( a43751a  and  a43748a );
 a43755a <=( (not A299)  and  A298 );
 a43758a <=( A301  and  A300 );
 a43759a <=( a43758a  and  a43755a );
 a43760a <=( a43759a  and  a43752a );
 a43764a <=( (not A168)  and  (not A169) );
 a43765a <=( A170  and  a43764a );
 a43768a <=( A166  and  (not A167) );
 a43771a <=( A200  and  A199 );
 a43772a <=( a43771a  and  a43768a );
 a43773a <=( a43772a  and  a43765a );
 a43776a <=( A233  and  (not A232) );
 a43779a <=( A236  and  A234 );
 a43780a <=( a43779a  and  a43776a );
 a43783a <=( (not A299)  and  A298 );
 a43786a <=( A302  and  A300 );
 a43787a <=( a43786a  and  a43783a );
 a43788a <=( a43787a  and  a43780a );
 a43792a <=( (not A168)  and  (not A169) );
 a43793a <=( A170  and  a43792a );
 a43796a <=( A166  and  (not A167) );
 a43799a <=( A200  and  A199 );
 a43800a <=( a43799a  and  a43796a );
 a43801a <=( a43800a  and  a43793a );
 a43804a <=( A233  and  (not A232) );
 a43807a <=( A236  and  A234 );
 a43808a <=( a43807a  and  a43804a );
 a43811a <=( A299  and  (not A298) );
 a43814a <=( A301  and  A300 );
 a43815a <=( a43814a  and  a43811a );
 a43816a <=( a43815a  and  a43808a );
 a43820a <=( (not A168)  and  (not A169) );
 a43821a <=( A170  and  a43820a );
 a43824a <=( A166  and  (not A167) );
 a43827a <=( A200  and  A199 );
 a43828a <=( a43827a  and  a43824a );
 a43829a <=( a43828a  and  a43821a );
 a43832a <=( A233  and  (not A232) );
 a43835a <=( A236  and  A234 );
 a43836a <=( a43835a  and  a43832a );
 a43839a <=( A299  and  (not A298) );
 a43842a <=( A302  and  A300 );
 a43843a <=( a43842a  and  a43839a );
 a43844a <=( a43843a  and  a43836a );
 a43848a <=( (not A168)  and  (not A169) );
 a43849a <=( A170  and  a43848a );
 a43852a <=( A166  and  (not A167) );
 a43855a <=( A200  and  A199 );
 a43856a <=( a43855a  and  a43852a );
 a43857a <=( a43856a  and  a43849a );
 a43860a <=( A233  and  (not A232) );
 a43863a <=( A236  and  A234 );
 a43864a <=( a43863a  and  a43860a );
 a43867a <=( A266  and  (not A265) );
 a43870a <=( A268  and  A267 );
 a43871a <=( a43870a  and  a43867a );
 a43872a <=( a43871a  and  a43864a );
 a43876a <=( (not A168)  and  (not A169) );
 a43877a <=( A170  and  a43876a );
 a43880a <=( A166  and  (not A167) );
 a43883a <=( A200  and  A199 );
 a43884a <=( a43883a  and  a43880a );
 a43885a <=( a43884a  and  a43877a );
 a43888a <=( A233  and  (not A232) );
 a43891a <=( A236  and  A234 );
 a43892a <=( a43891a  and  a43888a );
 a43895a <=( A266  and  (not A265) );
 a43898a <=( A269  and  A267 );
 a43899a <=( a43898a  and  a43895a );
 a43900a <=( a43899a  and  a43892a );
 a43904a <=( (not A168)  and  (not A169) );
 a43905a <=( A170  and  a43904a );
 a43908a <=( A166  and  (not A167) );
 a43911a <=( A200  and  A199 );
 a43912a <=( a43911a  and  a43908a );
 a43913a <=( a43912a  and  a43905a );
 a43916a <=( A233  and  (not A232) );
 a43919a <=( A236  and  A234 );
 a43920a <=( a43919a  and  a43916a );
 a43923a <=( (not A266)  and  A265 );
 a43926a <=( A268  and  A267 );
 a43927a <=( a43926a  and  a43923a );
 a43928a <=( a43927a  and  a43920a );
 a43932a <=( (not A168)  and  (not A169) );
 a43933a <=( A170  and  a43932a );
 a43936a <=( A166  and  (not A167) );
 a43939a <=( A200  and  A199 );
 a43940a <=( a43939a  and  a43936a );
 a43941a <=( a43940a  and  a43933a );
 a43944a <=( A233  and  (not A232) );
 a43947a <=( A236  and  A234 );
 a43948a <=( a43947a  and  a43944a );
 a43951a <=( (not A266)  and  A265 );
 a43954a <=( A269  and  A267 );
 a43955a <=( a43954a  and  a43951a );
 a43956a <=( a43955a  and  a43948a );
 a43960a <=( (not A168)  and  (not A169) );
 a43961a <=( A170  and  a43960a );
 a43964a <=( A166  and  (not A167) );
 a43967a <=( A200  and  A199 );
 a43968a <=( a43967a  and  a43964a );
 a43969a <=( a43968a  and  a43961a );
 a43972a <=( (not A233)  and  A232 );
 a43975a <=( A235  and  A234 );
 a43976a <=( a43975a  and  a43972a );
 a43979a <=( (not A299)  and  A298 );
 a43982a <=( A301  and  A300 );
 a43983a <=( a43982a  and  a43979a );
 a43984a <=( a43983a  and  a43976a );
 a43988a <=( (not A168)  and  (not A169) );
 a43989a <=( A170  and  a43988a );
 a43992a <=( A166  and  (not A167) );
 a43995a <=( A200  and  A199 );
 a43996a <=( a43995a  and  a43992a );
 a43997a <=( a43996a  and  a43989a );
 a44000a <=( (not A233)  and  A232 );
 a44003a <=( A235  and  A234 );
 a44004a <=( a44003a  and  a44000a );
 a44007a <=( (not A299)  and  A298 );
 a44010a <=( A302  and  A300 );
 a44011a <=( a44010a  and  a44007a );
 a44012a <=( a44011a  and  a44004a );
 a44016a <=( (not A168)  and  (not A169) );
 a44017a <=( A170  and  a44016a );
 a44020a <=( A166  and  (not A167) );
 a44023a <=( A200  and  A199 );
 a44024a <=( a44023a  and  a44020a );
 a44025a <=( a44024a  and  a44017a );
 a44028a <=( (not A233)  and  A232 );
 a44031a <=( A235  and  A234 );
 a44032a <=( a44031a  and  a44028a );
 a44035a <=( A299  and  (not A298) );
 a44038a <=( A301  and  A300 );
 a44039a <=( a44038a  and  a44035a );
 a44040a <=( a44039a  and  a44032a );
 a44044a <=( (not A168)  and  (not A169) );
 a44045a <=( A170  and  a44044a );
 a44048a <=( A166  and  (not A167) );
 a44051a <=( A200  and  A199 );
 a44052a <=( a44051a  and  a44048a );
 a44053a <=( a44052a  and  a44045a );
 a44056a <=( (not A233)  and  A232 );
 a44059a <=( A235  and  A234 );
 a44060a <=( a44059a  and  a44056a );
 a44063a <=( A299  and  (not A298) );
 a44066a <=( A302  and  A300 );
 a44067a <=( a44066a  and  a44063a );
 a44068a <=( a44067a  and  a44060a );
 a44072a <=( (not A168)  and  (not A169) );
 a44073a <=( A170  and  a44072a );
 a44076a <=( A166  and  (not A167) );
 a44079a <=( A200  and  A199 );
 a44080a <=( a44079a  and  a44076a );
 a44081a <=( a44080a  and  a44073a );
 a44084a <=( (not A233)  and  A232 );
 a44087a <=( A235  and  A234 );
 a44088a <=( a44087a  and  a44084a );
 a44091a <=( A266  and  (not A265) );
 a44094a <=( A268  and  A267 );
 a44095a <=( a44094a  and  a44091a );
 a44096a <=( a44095a  and  a44088a );
 a44100a <=( (not A168)  and  (not A169) );
 a44101a <=( A170  and  a44100a );
 a44104a <=( A166  and  (not A167) );
 a44107a <=( A200  and  A199 );
 a44108a <=( a44107a  and  a44104a );
 a44109a <=( a44108a  and  a44101a );
 a44112a <=( (not A233)  and  A232 );
 a44115a <=( A235  and  A234 );
 a44116a <=( a44115a  and  a44112a );
 a44119a <=( A266  and  (not A265) );
 a44122a <=( A269  and  A267 );
 a44123a <=( a44122a  and  a44119a );
 a44124a <=( a44123a  and  a44116a );
 a44128a <=( (not A168)  and  (not A169) );
 a44129a <=( A170  and  a44128a );
 a44132a <=( A166  and  (not A167) );
 a44135a <=( A200  and  A199 );
 a44136a <=( a44135a  and  a44132a );
 a44137a <=( a44136a  and  a44129a );
 a44140a <=( (not A233)  and  A232 );
 a44143a <=( A235  and  A234 );
 a44144a <=( a44143a  and  a44140a );
 a44147a <=( (not A266)  and  A265 );
 a44150a <=( A268  and  A267 );
 a44151a <=( a44150a  and  a44147a );
 a44152a <=( a44151a  and  a44144a );
 a44156a <=( (not A168)  and  (not A169) );
 a44157a <=( A170  and  a44156a );
 a44160a <=( A166  and  (not A167) );
 a44163a <=( A200  and  A199 );
 a44164a <=( a44163a  and  a44160a );
 a44165a <=( a44164a  and  a44157a );
 a44168a <=( (not A233)  and  A232 );
 a44171a <=( A235  and  A234 );
 a44172a <=( a44171a  and  a44168a );
 a44175a <=( (not A266)  and  A265 );
 a44178a <=( A269  and  A267 );
 a44179a <=( a44178a  and  a44175a );
 a44180a <=( a44179a  and  a44172a );
 a44184a <=( (not A168)  and  (not A169) );
 a44185a <=( A170  and  a44184a );
 a44188a <=( A166  and  (not A167) );
 a44191a <=( A200  and  A199 );
 a44192a <=( a44191a  and  a44188a );
 a44193a <=( a44192a  and  a44185a );
 a44196a <=( (not A233)  and  A232 );
 a44199a <=( A236  and  A234 );
 a44200a <=( a44199a  and  a44196a );
 a44203a <=( (not A299)  and  A298 );
 a44206a <=( A301  and  A300 );
 a44207a <=( a44206a  and  a44203a );
 a44208a <=( a44207a  and  a44200a );
 a44212a <=( (not A168)  and  (not A169) );
 a44213a <=( A170  and  a44212a );
 a44216a <=( A166  and  (not A167) );
 a44219a <=( A200  and  A199 );
 a44220a <=( a44219a  and  a44216a );
 a44221a <=( a44220a  and  a44213a );
 a44224a <=( (not A233)  and  A232 );
 a44227a <=( A236  and  A234 );
 a44228a <=( a44227a  and  a44224a );
 a44231a <=( (not A299)  and  A298 );
 a44234a <=( A302  and  A300 );
 a44235a <=( a44234a  and  a44231a );
 a44236a <=( a44235a  and  a44228a );
 a44240a <=( (not A168)  and  (not A169) );
 a44241a <=( A170  and  a44240a );
 a44244a <=( A166  and  (not A167) );
 a44247a <=( A200  and  A199 );
 a44248a <=( a44247a  and  a44244a );
 a44249a <=( a44248a  and  a44241a );
 a44252a <=( (not A233)  and  A232 );
 a44255a <=( A236  and  A234 );
 a44256a <=( a44255a  and  a44252a );
 a44259a <=( A299  and  (not A298) );
 a44262a <=( A301  and  A300 );
 a44263a <=( a44262a  and  a44259a );
 a44264a <=( a44263a  and  a44256a );
 a44268a <=( (not A168)  and  (not A169) );
 a44269a <=( A170  and  a44268a );
 a44272a <=( A166  and  (not A167) );
 a44275a <=( A200  and  A199 );
 a44276a <=( a44275a  and  a44272a );
 a44277a <=( a44276a  and  a44269a );
 a44280a <=( (not A233)  and  A232 );
 a44283a <=( A236  and  A234 );
 a44284a <=( a44283a  and  a44280a );
 a44287a <=( A299  and  (not A298) );
 a44290a <=( A302  and  A300 );
 a44291a <=( a44290a  and  a44287a );
 a44292a <=( a44291a  and  a44284a );
 a44296a <=( (not A168)  and  (not A169) );
 a44297a <=( A170  and  a44296a );
 a44300a <=( A166  and  (not A167) );
 a44303a <=( A200  and  A199 );
 a44304a <=( a44303a  and  a44300a );
 a44305a <=( a44304a  and  a44297a );
 a44308a <=( (not A233)  and  A232 );
 a44311a <=( A236  and  A234 );
 a44312a <=( a44311a  and  a44308a );
 a44315a <=( A266  and  (not A265) );
 a44318a <=( A268  and  A267 );
 a44319a <=( a44318a  and  a44315a );
 a44320a <=( a44319a  and  a44312a );
 a44324a <=( (not A168)  and  (not A169) );
 a44325a <=( A170  and  a44324a );
 a44328a <=( A166  and  (not A167) );
 a44331a <=( A200  and  A199 );
 a44332a <=( a44331a  and  a44328a );
 a44333a <=( a44332a  and  a44325a );
 a44336a <=( (not A233)  and  A232 );
 a44339a <=( A236  and  A234 );
 a44340a <=( a44339a  and  a44336a );
 a44343a <=( A266  and  (not A265) );
 a44346a <=( A269  and  A267 );
 a44347a <=( a44346a  and  a44343a );
 a44348a <=( a44347a  and  a44340a );
 a44352a <=( (not A168)  and  (not A169) );
 a44353a <=( A170  and  a44352a );
 a44356a <=( A166  and  (not A167) );
 a44359a <=( A200  and  A199 );
 a44360a <=( a44359a  and  a44356a );
 a44361a <=( a44360a  and  a44353a );
 a44364a <=( (not A233)  and  A232 );
 a44367a <=( A236  and  A234 );
 a44368a <=( a44367a  and  a44364a );
 a44371a <=( (not A266)  and  A265 );
 a44374a <=( A268  and  A267 );
 a44375a <=( a44374a  and  a44371a );
 a44376a <=( a44375a  and  a44368a );
 a44380a <=( (not A168)  and  (not A169) );
 a44381a <=( A170  and  a44380a );
 a44384a <=( A166  and  (not A167) );
 a44387a <=( A200  and  A199 );
 a44388a <=( a44387a  and  a44384a );
 a44389a <=( a44388a  and  a44381a );
 a44392a <=( (not A233)  and  A232 );
 a44395a <=( A236  and  A234 );
 a44396a <=( a44395a  and  a44392a );
 a44399a <=( (not A266)  and  A265 );
 a44402a <=( A269  and  A267 );
 a44403a <=( a44402a  and  a44399a );
 a44404a <=( a44403a  and  a44396a );
 a44408a <=( (not A168)  and  (not A169) );
 a44409a <=( A170  and  a44408a );
 a44412a <=( A166  and  (not A167) );
 a44415a <=( (not A200)  and  (not A199) );
 a44416a <=( a44415a  and  a44412a );
 a44417a <=( a44416a  and  a44409a );
 a44420a <=( A233  and  (not A232) );
 a44423a <=( A235  and  A234 );
 a44424a <=( a44423a  and  a44420a );
 a44427a <=( (not A299)  and  A298 );
 a44430a <=( A301  and  A300 );
 a44431a <=( a44430a  and  a44427a );
 a44432a <=( a44431a  and  a44424a );
 a44436a <=( (not A168)  and  (not A169) );
 a44437a <=( A170  and  a44436a );
 a44440a <=( A166  and  (not A167) );
 a44443a <=( (not A200)  and  (not A199) );
 a44444a <=( a44443a  and  a44440a );
 a44445a <=( a44444a  and  a44437a );
 a44448a <=( A233  and  (not A232) );
 a44451a <=( A235  and  A234 );
 a44452a <=( a44451a  and  a44448a );
 a44455a <=( (not A299)  and  A298 );
 a44458a <=( A302  and  A300 );
 a44459a <=( a44458a  and  a44455a );
 a44460a <=( a44459a  and  a44452a );
 a44464a <=( (not A168)  and  (not A169) );
 a44465a <=( A170  and  a44464a );
 a44468a <=( A166  and  (not A167) );
 a44471a <=( (not A200)  and  (not A199) );
 a44472a <=( a44471a  and  a44468a );
 a44473a <=( a44472a  and  a44465a );
 a44476a <=( A233  and  (not A232) );
 a44479a <=( A235  and  A234 );
 a44480a <=( a44479a  and  a44476a );
 a44483a <=( A299  and  (not A298) );
 a44486a <=( A301  and  A300 );
 a44487a <=( a44486a  and  a44483a );
 a44488a <=( a44487a  and  a44480a );
 a44492a <=( (not A168)  and  (not A169) );
 a44493a <=( A170  and  a44492a );
 a44496a <=( A166  and  (not A167) );
 a44499a <=( (not A200)  and  (not A199) );
 a44500a <=( a44499a  and  a44496a );
 a44501a <=( a44500a  and  a44493a );
 a44504a <=( A233  and  (not A232) );
 a44507a <=( A235  and  A234 );
 a44508a <=( a44507a  and  a44504a );
 a44511a <=( A299  and  (not A298) );
 a44514a <=( A302  and  A300 );
 a44515a <=( a44514a  and  a44511a );
 a44516a <=( a44515a  and  a44508a );
 a44520a <=( (not A168)  and  (not A169) );
 a44521a <=( A170  and  a44520a );
 a44524a <=( A166  and  (not A167) );
 a44527a <=( (not A200)  and  (not A199) );
 a44528a <=( a44527a  and  a44524a );
 a44529a <=( a44528a  and  a44521a );
 a44532a <=( A233  and  (not A232) );
 a44535a <=( A235  and  A234 );
 a44536a <=( a44535a  and  a44532a );
 a44539a <=( A266  and  (not A265) );
 a44542a <=( A268  and  A267 );
 a44543a <=( a44542a  and  a44539a );
 a44544a <=( a44543a  and  a44536a );
 a44548a <=( (not A168)  and  (not A169) );
 a44549a <=( A170  and  a44548a );
 a44552a <=( A166  and  (not A167) );
 a44555a <=( (not A200)  and  (not A199) );
 a44556a <=( a44555a  and  a44552a );
 a44557a <=( a44556a  and  a44549a );
 a44560a <=( A233  and  (not A232) );
 a44563a <=( A235  and  A234 );
 a44564a <=( a44563a  and  a44560a );
 a44567a <=( A266  and  (not A265) );
 a44570a <=( A269  and  A267 );
 a44571a <=( a44570a  and  a44567a );
 a44572a <=( a44571a  and  a44564a );
 a44576a <=( (not A168)  and  (not A169) );
 a44577a <=( A170  and  a44576a );
 a44580a <=( A166  and  (not A167) );
 a44583a <=( (not A200)  and  (not A199) );
 a44584a <=( a44583a  and  a44580a );
 a44585a <=( a44584a  and  a44577a );
 a44588a <=( A233  and  (not A232) );
 a44591a <=( A235  and  A234 );
 a44592a <=( a44591a  and  a44588a );
 a44595a <=( (not A266)  and  A265 );
 a44598a <=( A268  and  A267 );
 a44599a <=( a44598a  and  a44595a );
 a44600a <=( a44599a  and  a44592a );
 a44604a <=( (not A168)  and  (not A169) );
 a44605a <=( A170  and  a44604a );
 a44608a <=( A166  and  (not A167) );
 a44611a <=( (not A200)  and  (not A199) );
 a44612a <=( a44611a  and  a44608a );
 a44613a <=( a44612a  and  a44605a );
 a44616a <=( A233  and  (not A232) );
 a44619a <=( A235  and  A234 );
 a44620a <=( a44619a  and  a44616a );
 a44623a <=( (not A266)  and  A265 );
 a44626a <=( A269  and  A267 );
 a44627a <=( a44626a  and  a44623a );
 a44628a <=( a44627a  and  a44620a );
 a44632a <=( (not A168)  and  (not A169) );
 a44633a <=( A170  and  a44632a );
 a44636a <=( A166  and  (not A167) );
 a44639a <=( (not A200)  and  (not A199) );
 a44640a <=( a44639a  and  a44636a );
 a44641a <=( a44640a  and  a44633a );
 a44644a <=( A233  and  (not A232) );
 a44647a <=( A236  and  A234 );
 a44648a <=( a44647a  and  a44644a );
 a44651a <=( (not A299)  and  A298 );
 a44654a <=( A301  and  A300 );
 a44655a <=( a44654a  and  a44651a );
 a44656a <=( a44655a  and  a44648a );
 a44660a <=( (not A168)  and  (not A169) );
 a44661a <=( A170  and  a44660a );
 a44664a <=( A166  and  (not A167) );
 a44667a <=( (not A200)  and  (not A199) );
 a44668a <=( a44667a  and  a44664a );
 a44669a <=( a44668a  and  a44661a );
 a44672a <=( A233  and  (not A232) );
 a44675a <=( A236  and  A234 );
 a44676a <=( a44675a  and  a44672a );
 a44679a <=( (not A299)  and  A298 );
 a44682a <=( A302  and  A300 );
 a44683a <=( a44682a  and  a44679a );
 a44684a <=( a44683a  and  a44676a );
 a44688a <=( (not A168)  and  (not A169) );
 a44689a <=( A170  and  a44688a );
 a44692a <=( A166  and  (not A167) );
 a44695a <=( (not A200)  and  (not A199) );
 a44696a <=( a44695a  and  a44692a );
 a44697a <=( a44696a  and  a44689a );
 a44700a <=( A233  and  (not A232) );
 a44703a <=( A236  and  A234 );
 a44704a <=( a44703a  and  a44700a );
 a44707a <=( A299  and  (not A298) );
 a44710a <=( A301  and  A300 );
 a44711a <=( a44710a  and  a44707a );
 a44712a <=( a44711a  and  a44704a );
 a44716a <=( (not A168)  and  (not A169) );
 a44717a <=( A170  and  a44716a );
 a44720a <=( A166  and  (not A167) );
 a44723a <=( (not A200)  and  (not A199) );
 a44724a <=( a44723a  and  a44720a );
 a44725a <=( a44724a  and  a44717a );
 a44728a <=( A233  and  (not A232) );
 a44731a <=( A236  and  A234 );
 a44732a <=( a44731a  and  a44728a );
 a44735a <=( A299  and  (not A298) );
 a44738a <=( A302  and  A300 );
 a44739a <=( a44738a  and  a44735a );
 a44740a <=( a44739a  and  a44732a );
 a44744a <=( (not A168)  and  (not A169) );
 a44745a <=( A170  and  a44744a );
 a44748a <=( A166  and  (not A167) );
 a44751a <=( (not A200)  and  (not A199) );
 a44752a <=( a44751a  and  a44748a );
 a44753a <=( a44752a  and  a44745a );
 a44756a <=( A233  and  (not A232) );
 a44759a <=( A236  and  A234 );
 a44760a <=( a44759a  and  a44756a );
 a44763a <=( A266  and  (not A265) );
 a44766a <=( A268  and  A267 );
 a44767a <=( a44766a  and  a44763a );
 a44768a <=( a44767a  and  a44760a );
 a44772a <=( (not A168)  and  (not A169) );
 a44773a <=( A170  and  a44772a );
 a44776a <=( A166  and  (not A167) );
 a44779a <=( (not A200)  and  (not A199) );
 a44780a <=( a44779a  and  a44776a );
 a44781a <=( a44780a  and  a44773a );
 a44784a <=( A233  and  (not A232) );
 a44787a <=( A236  and  A234 );
 a44788a <=( a44787a  and  a44784a );
 a44791a <=( A266  and  (not A265) );
 a44794a <=( A269  and  A267 );
 a44795a <=( a44794a  and  a44791a );
 a44796a <=( a44795a  and  a44788a );
 a44800a <=( (not A168)  and  (not A169) );
 a44801a <=( A170  and  a44800a );
 a44804a <=( A166  and  (not A167) );
 a44807a <=( (not A200)  and  (not A199) );
 a44808a <=( a44807a  and  a44804a );
 a44809a <=( a44808a  and  a44801a );
 a44812a <=( A233  and  (not A232) );
 a44815a <=( A236  and  A234 );
 a44816a <=( a44815a  and  a44812a );
 a44819a <=( (not A266)  and  A265 );
 a44822a <=( A268  and  A267 );
 a44823a <=( a44822a  and  a44819a );
 a44824a <=( a44823a  and  a44816a );
 a44828a <=( (not A168)  and  (not A169) );
 a44829a <=( A170  and  a44828a );
 a44832a <=( A166  and  (not A167) );
 a44835a <=( (not A200)  and  (not A199) );
 a44836a <=( a44835a  and  a44832a );
 a44837a <=( a44836a  and  a44829a );
 a44840a <=( A233  and  (not A232) );
 a44843a <=( A236  and  A234 );
 a44844a <=( a44843a  and  a44840a );
 a44847a <=( (not A266)  and  A265 );
 a44850a <=( A269  and  A267 );
 a44851a <=( a44850a  and  a44847a );
 a44852a <=( a44851a  and  a44844a );
 a44856a <=( (not A168)  and  (not A169) );
 a44857a <=( A170  and  a44856a );
 a44860a <=( A166  and  (not A167) );
 a44863a <=( (not A200)  and  (not A199) );
 a44864a <=( a44863a  and  a44860a );
 a44865a <=( a44864a  and  a44857a );
 a44868a <=( (not A233)  and  A232 );
 a44871a <=( A235  and  A234 );
 a44872a <=( a44871a  and  a44868a );
 a44875a <=( (not A299)  and  A298 );
 a44878a <=( A301  and  A300 );
 a44879a <=( a44878a  and  a44875a );
 a44880a <=( a44879a  and  a44872a );
 a44884a <=( (not A168)  and  (not A169) );
 a44885a <=( A170  and  a44884a );
 a44888a <=( A166  and  (not A167) );
 a44891a <=( (not A200)  and  (not A199) );
 a44892a <=( a44891a  and  a44888a );
 a44893a <=( a44892a  and  a44885a );
 a44896a <=( (not A233)  and  A232 );
 a44899a <=( A235  and  A234 );
 a44900a <=( a44899a  and  a44896a );
 a44903a <=( (not A299)  and  A298 );
 a44906a <=( A302  and  A300 );
 a44907a <=( a44906a  and  a44903a );
 a44908a <=( a44907a  and  a44900a );
 a44912a <=( (not A168)  and  (not A169) );
 a44913a <=( A170  and  a44912a );
 a44916a <=( A166  and  (not A167) );
 a44919a <=( (not A200)  and  (not A199) );
 a44920a <=( a44919a  and  a44916a );
 a44921a <=( a44920a  and  a44913a );
 a44924a <=( (not A233)  and  A232 );
 a44927a <=( A235  and  A234 );
 a44928a <=( a44927a  and  a44924a );
 a44931a <=( A299  and  (not A298) );
 a44934a <=( A301  and  A300 );
 a44935a <=( a44934a  and  a44931a );
 a44936a <=( a44935a  and  a44928a );
 a44940a <=( (not A168)  and  (not A169) );
 a44941a <=( A170  and  a44940a );
 a44944a <=( A166  and  (not A167) );
 a44947a <=( (not A200)  and  (not A199) );
 a44948a <=( a44947a  and  a44944a );
 a44949a <=( a44948a  and  a44941a );
 a44952a <=( (not A233)  and  A232 );
 a44955a <=( A235  and  A234 );
 a44956a <=( a44955a  and  a44952a );
 a44959a <=( A299  and  (not A298) );
 a44962a <=( A302  and  A300 );
 a44963a <=( a44962a  and  a44959a );
 a44964a <=( a44963a  and  a44956a );
 a44968a <=( (not A168)  and  (not A169) );
 a44969a <=( A170  and  a44968a );
 a44972a <=( A166  and  (not A167) );
 a44975a <=( (not A200)  and  (not A199) );
 a44976a <=( a44975a  and  a44972a );
 a44977a <=( a44976a  and  a44969a );
 a44980a <=( (not A233)  and  A232 );
 a44983a <=( A235  and  A234 );
 a44984a <=( a44983a  and  a44980a );
 a44987a <=( A266  and  (not A265) );
 a44990a <=( A268  and  A267 );
 a44991a <=( a44990a  and  a44987a );
 a44992a <=( a44991a  and  a44984a );
 a44996a <=( (not A168)  and  (not A169) );
 a44997a <=( A170  and  a44996a );
 a45000a <=( A166  and  (not A167) );
 a45003a <=( (not A200)  and  (not A199) );
 a45004a <=( a45003a  and  a45000a );
 a45005a <=( a45004a  and  a44997a );
 a45008a <=( (not A233)  and  A232 );
 a45011a <=( A235  and  A234 );
 a45012a <=( a45011a  and  a45008a );
 a45015a <=( A266  and  (not A265) );
 a45018a <=( A269  and  A267 );
 a45019a <=( a45018a  and  a45015a );
 a45020a <=( a45019a  and  a45012a );
 a45024a <=( (not A168)  and  (not A169) );
 a45025a <=( A170  and  a45024a );
 a45028a <=( A166  and  (not A167) );
 a45031a <=( (not A200)  and  (not A199) );
 a45032a <=( a45031a  and  a45028a );
 a45033a <=( a45032a  and  a45025a );
 a45036a <=( (not A233)  and  A232 );
 a45039a <=( A235  and  A234 );
 a45040a <=( a45039a  and  a45036a );
 a45043a <=( (not A266)  and  A265 );
 a45046a <=( A268  and  A267 );
 a45047a <=( a45046a  and  a45043a );
 a45048a <=( a45047a  and  a45040a );
 a45052a <=( (not A168)  and  (not A169) );
 a45053a <=( A170  and  a45052a );
 a45056a <=( A166  and  (not A167) );
 a45059a <=( (not A200)  and  (not A199) );
 a45060a <=( a45059a  and  a45056a );
 a45061a <=( a45060a  and  a45053a );
 a45064a <=( (not A233)  and  A232 );
 a45067a <=( A235  and  A234 );
 a45068a <=( a45067a  and  a45064a );
 a45071a <=( (not A266)  and  A265 );
 a45074a <=( A269  and  A267 );
 a45075a <=( a45074a  and  a45071a );
 a45076a <=( a45075a  and  a45068a );
 a45080a <=( (not A168)  and  (not A169) );
 a45081a <=( A170  and  a45080a );
 a45084a <=( A166  and  (not A167) );
 a45087a <=( (not A200)  and  (not A199) );
 a45088a <=( a45087a  and  a45084a );
 a45089a <=( a45088a  and  a45081a );
 a45092a <=( (not A233)  and  A232 );
 a45095a <=( A236  and  A234 );
 a45096a <=( a45095a  and  a45092a );
 a45099a <=( (not A299)  and  A298 );
 a45102a <=( A301  and  A300 );
 a45103a <=( a45102a  and  a45099a );
 a45104a <=( a45103a  and  a45096a );
 a45108a <=( (not A168)  and  (not A169) );
 a45109a <=( A170  and  a45108a );
 a45112a <=( A166  and  (not A167) );
 a45115a <=( (not A200)  and  (not A199) );
 a45116a <=( a45115a  and  a45112a );
 a45117a <=( a45116a  and  a45109a );
 a45120a <=( (not A233)  and  A232 );
 a45123a <=( A236  and  A234 );
 a45124a <=( a45123a  and  a45120a );
 a45127a <=( (not A299)  and  A298 );
 a45130a <=( A302  and  A300 );
 a45131a <=( a45130a  and  a45127a );
 a45132a <=( a45131a  and  a45124a );
 a45136a <=( (not A168)  and  (not A169) );
 a45137a <=( A170  and  a45136a );
 a45140a <=( A166  and  (not A167) );
 a45143a <=( (not A200)  and  (not A199) );
 a45144a <=( a45143a  and  a45140a );
 a45145a <=( a45144a  and  a45137a );
 a45148a <=( (not A233)  and  A232 );
 a45151a <=( A236  and  A234 );
 a45152a <=( a45151a  and  a45148a );
 a45155a <=( A299  and  (not A298) );
 a45158a <=( A301  and  A300 );
 a45159a <=( a45158a  and  a45155a );
 a45160a <=( a45159a  and  a45152a );
 a45164a <=( (not A168)  and  (not A169) );
 a45165a <=( A170  and  a45164a );
 a45168a <=( A166  and  (not A167) );
 a45171a <=( (not A200)  and  (not A199) );
 a45172a <=( a45171a  and  a45168a );
 a45173a <=( a45172a  and  a45165a );
 a45176a <=( (not A233)  and  A232 );
 a45179a <=( A236  and  A234 );
 a45180a <=( a45179a  and  a45176a );
 a45183a <=( A299  and  (not A298) );
 a45186a <=( A302  and  A300 );
 a45187a <=( a45186a  and  a45183a );
 a45188a <=( a45187a  and  a45180a );
 a45192a <=( (not A168)  and  (not A169) );
 a45193a <=( A170  and  a45192a );
 a45196a <=( A166  and  (not A167) );
 a45199a <=( (not A200)  and  (not A199) );
 a45200a <=( a45199a  and  a45196a );
 a45201a <=( a45200a  and  a45193a );
 a45204a <=( (not A233)  and  A232 );
 a45207a <=( A236  and  A234 );
 a45208a <=( a45207a  and  a45204a );
 a45211a <=( A266  and  (not A265) );
 a45214a <=( A268  and  A267 );
 a45215a <=( a45214a  and  a45211a );
 a45216a <=( a45215a  and  a45208a );
 a45220a <=( (not A168)  and  (not A169) );
 a45221a <=( A170  and  a45220a );
 a45224a <=( A166  and  (not A167) );
 a45227a <=( (not A200)  and  (not A199) );
 a45228a <=( a45227a  and  a45224a );
 a45229a <=( a45228a  and  a45221a );
 a45232a <=( (not A233)  and  A232 );
 a45235a <=( A236  and  A234 );
 a45236a <=( a45235a  and  a45232a );
 a45239a <=( A266  and  (not A265) );
 a45242a <=( A269  and  A267 );
 a45243a <=( a45242a  and  a45239a );
 a45244a <=( a45243a  and  a45236a );
 a45248a <=( (not A168)  and  (not A169) );
 a45249a <=( A170  and  a45248a );
 a45252a <=( A166  and  (not A167) );
 a45255a <=( (not A200)  and  (not A199) );
 a45256a <=( a45255a  and  a45252a );
 a45257a <=( a45256a  and  a45249a );
 a45260a <=( (not A233)  and  A232 );
 a45263a <=( A236  and  A234 );
 a45264a <=( a45263a  and  a45260a );
 a45267a <=( (not A266)  and  A265 );
 a45270a <=( A268  and  A267 );
 a45271a <=( a45270a  and  a45267a );
 a45272a <=( a45271a  and  a45264a );
 a45276a <=( (not A168)  and  (not A169) );
 a45277a <=( A170  and  a45276a );
 a45280a <=( A166  and  (not A167) );
 a45283a <=( (not A200)  and  (not A199) );
 a45284a <=( a45283a  and  a45280a );
 a45285a <=( a45284a  and  a45277a );
 a45288a <=( (not A233)  and  A232 );
 a45291a <=( A236  and  A234 );
 a45292a <=( a45291a  and  a45288a );
 a45295a <=( (not A266)  and  A265 );
 a45298a <=( A269  and  A267 );
 a45299a <=( a45298a  and  a45295a );
 a45300a <=( a45299a  and  a45292a );
 a45303a <=( A168  and  (not A170) );
 a45306a <=( (not A166)  and  A167 );
 a45307a <=( a45306a  and  a45303a );
 a45310a <=( (not A202)  and  A201 );
 a45313a <=( (not A232)  and  (not A203) );
 a45314a <=( a45313a  and  a45310a );
 a45315a <=( a45314a  and  a45307a );
 a45318a <=( A234  and  A233 );
 a45321a <=( A298  and  A235 );
 a45322a <=( a45321a  and  a45318a );
 a45325a <=( (not A300)  and  (not A299) );
 a45328a <=( (not A302)  and  (not A301) );
 a45329a <=( a45328a  and  a45325a );
 a45330a <=( a45329a  and  a45322a );
 a45333a <=( A168  and  (not A170) );
 a45336a <=( (not A166)  and  A167 );
 a45337a <=( a45336a  and  a45333a );
 a45340a <=( (not A202)  and  A201 );
 a45343a <=( (not A232)  and  (not A203) );
 a45344a <=( a45343a  and  a45340a );
 a45345a <=( a45344a  and  a45337a );
 a45348a <=( A234  and  A233 );
 a45351a <=( (not A298)  and  A235 );
 a45352a <=( a45351a  and  a45348a );
 a45355a <=( (not A300)  and  A299 );
 a45358a <=( (not A302)  and  (not A301) );
 a45359a <=( a45358a  and  a45355a );
 a45360a <=( a45359a  and  a45352a );
 a45363a <=( A168  and  (not A170) );
 a45366a <=( (not A166)  and  A167 );
 a45367a <=( a45366a  and  a45363a );
 a45370a <=( (not A202)  and  A201 );
 a45373a <=( (not A232)  and  (not A203) );
 a45374a <=( a45373a  and  a45370a );
 a45375a <=( a45374a  and  a45367a );
 a45378a <=( A234  and  A233 );
 a45381a <=( (not A265)  and  A235 );
 a45382a <=( a45381a  and  a45378a );
 a45385a <=( (not A267)  and  A266 );
 a45388a <=( (not A269)  and  (not A268) );
 a45389a <=( a45388a  and  a45385a );
 a45390a <=( a45389a  and  a45382a );
 a45393a <=( A168  and  (not A170) );
 a45396a <=( (not A166)  and  A167 );
 a45397a <=( a45396a  and  a45393a );
 a45400a <=( (not A202)  and  A201 );
 a45403a <=( (not A232)  and  (not A203) );
 a45404a <=( a45403a  and  a45400a );
 a45405a <=( a45404a  and  a45397a );
 a45408a <=( A234  and  A233 );
 a45411a <=( A265  and  A235 );
 a45412a <=( a45411a  and  a45408a );
 a45415a <=( (not A267)  and  (not A266) );
 a45418a <=( (not A269)  and  (not A268) );
 a45419a <=( a45418a  and  a45415a );
 a45420a <=( a45419a  and  a45412a );
 a45423a <=( A168  and  (not A170) );
 a45426a <=( (not A166)  and  A167 );
 a45427a <=( a45426a  and  a45423a );
 a45430a <=( (not A202)  and  A201 );
 a45433a <=( (not A232)  and  (not A203) );
 a45434a <=( a45433a  and  a45430a );
 a45435a <=( a45434a  and  a45427a );
 a45438a <=( A234  and  A233 );
 a45441a <=( A298  and  A236 );
 a45442a <=( a45441a  and  a45438a );
 a45445a <=( (not A300)  and  (not A299) );
 a45448a <=( (not A302)  and  (not A301) );
 a45449a <=( a45448a  and  a45445a );
 a45450a <=( a45449a  and  a45442a );
 a45453a <=( A168  and  (not A170) );
 a45456a <=( (not A166)  and  A167 );
 a45457a <=( a45456a  and  a45453a );
 a45460a <=( (not A202)  and  A201 );
 a45463a <=( (not A232)  and  (not A203) );
 a45464a <=( a45463a  and  a45460a );
 a45465a <=( a45464a  and  a45457a );
 a45468a <=( A234  and  A233 );
 a45471a <=( (not A298)  and  A236 );
 a45472a <=( a45471a  and  a45468a );
 a45475a <=( (not A300)  and  A299 );
 a45478a <=( (not A302)  and  (not A301) );
 a45479a <=( a45478a  and  a45475a );
 a45480a <=( a45479a  and  a45472a );
 a45483a <=( A168  and  (not A170) );
 a45486a <=( (not A166)  and  A167 );
 a45487a <=( a45486a  and  a45483a );
 a45490a <=( (not A202)  and  A201 );
 a45493a <=( (not A232)  and  (not A203) );
 a45494a <=( a45493a  and  a45490a );
 a45495a <=( a45494a  and  a45487a );
 a45498a <=( A234  and  A233 );
 a45501a <=( (not A265)  and  A236 );
 a45502a <=( a45501a  and  a45498a );
 a45505a <=( (not A267)  and  A266 );
 a45508a <=( (not A269)  and  (not A268) );
 a45509a <=( a45508a  and  a45505a );
 a45510a <=( a45509a  and  a45502a );
 a45513a <=( A168  and  (not A170) );
 a45516a <=( (not A166)  and  A167 );
 a45517a <=( a45516a  and  a45513a );
 a45520a <=( (not A202)  and  A201 );
 a45523a <=( (not A232)  and  (not A203) );
 a45524a <=( a45523a  and  a45520a );
 a45525a <=( a45524a  and  a45517a );
 a45528a <=( A234  and  A233 );
 a45531a <=( A265  and  A236 );
 a45532a <=( a45531a  and  a45528a );
 a45535a <=( (not A267)  and  (not A266) );
 a45538a <=( (not A269)  and  (not A268) );
 a45539a <=( a45538a  and  a45535a );
 a45540a <=( a45539a  and  a45532a );
 a45543a <=( A168  and  (not A170) );
 a45546a <=( (not A166)  and  A167 );
 a45547a <=( a45546a  and  a45543a );
 a45550a <=( (not A202)  and  A201 );
 a45553a <=( (not A232)  and  (not A203) );
 a45554a <=( a45553a  and  a45550a );
 a45555a <=( a45554a  and  a45547a );
 a45558a <=( (not A234)  and  A233 );
 a45561a <=( (not A236)  and  (not A235) );
 a45562a <=( a45561a  and  a45558a );
 a45565a <=( (not A299)  and  A298 );
 a45568a <=( A301  and  A300 );
 a45569a <=( a45568a  and  a45565a );
 a45570a <=( a45569a  and  a45562a );
 a45573a <=( A168  and  (not A170) );
 a45576a <=( (not A166)  and  A167 );
 a45577a <=( a45576a  and  a45573a );
 a45580a <=( (not A202)  and  A201 );
 a45583a <=( (not A232)  and  (not A203) );
 a45584a <=( a45583a  and  a45580a );
 a45585a <=( a45584a  and  a45577a );
 a45588a <=( (not A234)  and  A233 );
 a45591a <=( (not A236)  and  (not A235) );
 a45592a <=( a45591a  and  a45588a );
 a45595a <=( (not A299)  and  A298 );
 a45598a <=( A302  and  A300 );
 a45599a <=( a45598a  and  a45595a );
 a45600a <=( a45599a  and  a45592a );
 a45603a <=( A168  and  (not A170) );
 a45606a <=( (not A166)  and  A167 );
 a45607a <=( a45606a  and  a45603a );
 a45610a <=( (not A202)  and  A201 );
 a45613a <=( (not A232)  and  (not A203) );
 a45614a <=( a45613a  and  a45610a );
 a45615a <=( a45614a  and  a45607a );
 a45618a <=( (not A234)  and  A233 );
 a45621a <=( (not A236)  and  (not A235) );
 a45622a <=( a45621a  and  a45618a );
 a45625a <=( A299  and  (not A298) );
 a45628a <=( A301  and  A300 );
 a45629a <=( a45628a  and  a45625a );
 a45630a <=( a45629a  and  a45622a );
 a45633a <=( A168  and  (not A170) );
 a45636a <=( (not A166)  and  A167 );
 a45637a <=( a45636a  and  a45633a );
 a45640a <=( (not A202)  and  A201 );
 a45643a <=( (not A232)  and  (not A203) );
 a45644a <=( a45643a  and  a45640a );
 a45645a <=( a45644a  and  a45637a );
 a45648a <=( (not A234)  and  A233 );
 a45651a <=( (not A236)  and  (not A235) );
 a45652a <=( a45651a  and  a45648a );
 a45655a <=( A299  and  (not A298) );
 a45658a <=( A302  and  A300 );
 a45659a <=( a45658a  and  a45655a );
 a45660a <=( a45659a  and  a45652a );
 a45663a <=( A168  and  (not A170) );
 a45666a <=( (not A166)  and  A167 );
 a45667a <=( a45666a  and  a45663a );
 a45670a <=( (not A202)  and  A201 );
 a45673a <=( (not A232)  and  (not A203) );
 a45674a <=( a45673a  and  a45670a );
 a45675a <=( a45674a  and  a45667a );
 a45678a <=( (not A234)  and  A233 );
 a45681a <=( (not A236)  and  (not A235) );
 a45682a <=( a45681a  and  a45678a );
 a45685a <=( A266  and  (not A265) );
 a45688a <=( A268  and  A267 );
 a45689a <=( a45688a  and  a45685a );
 a45690a <=( a45689a  and  a45682a );
 a45693a <=( A168  and  (not A170) );
 a45696a <=( (not A166)  and  A167 );
 a45697a <=( a45696a  and  a45693a );
 a45700a <=( (not A202)  and  A201 );
 a45703a <=( (not A232)  and  (not A203) );
 a45704a <=( a45703a  and  a45700a );
 a45705a <=( a45704a  and  a45697a );
 a45708a <=( (not A234)  and  A233 );
 a45711a <=( (not A236)  and  (not A235) );
 a45712a <=( a45711a  and  a45708a );
 a45715a <=( A266  and  (not A265) );
 a45718a <=( A269  and  A267 );
 a45719a <=( a45718a  and  a45715a );
 a45720a <=( a45719a  and  a45712a );
 a45723a <=( A168  and  (not A170) );
 a45726a <=( (not A166)  and  A167 );
 a45727a <=( a45726a  and  a45723a );
 a45730a <=( (not A202)  and  A201 );
 a45733a <=( (not A232)  and  (not A203) );
 a45734a <=( a45733a  and  a45730a );
 a45735a <=( a45734a  and  a45727a );
 a45738a <=( (not A234)  and  A233 );
 a45741a <=( (not A236)  and  (not A235) );
 a45742a <=( a45741a  and  a45738a );
 a45745a <=( (not A266)  and  A265 );
 a45748a <=( A268  and  A267 );
 a45749a <=( a45748a  and  a45745a );
 a45750a <=( a45749a  and  a45742a );
 a45753a <=( A168  and  (not A170) );
 a45756a <=( (not A166)  and  A167 );
 a45757a <=( a45756a  and  a45753a );
 a45760a <=( (not A202)  and  A201 );
 a45763a <=( (not A232)  and  (not A203) );
 a45764a <=( a45763a  and  a45760a );
 a45765a <=( a45764a  and  a45757a );
 a45768a <=( (not A234)  and  A233 );
 a45771a <=( (not A236)  and  (not A235) );
 a45772a <=( a45771a  and  a45768a );
 a45775a <=( (not A266)  and  A265 );
 a45778a <=( A269  and  A267 );
 a45779a <=( a45778a  and  a45775a );
 a45780a <=( a45779a  and  a45772a );
 a45783a <=( A168  and  (not A170) );
 a45786a <=( (not A166)  and  A167 );
 a45787a <=( a45786a  and  a45783a );
 a45790a <=( (not A202)  and  A201 );
 a45793a <=( A232  and  (not A203) );
 a45794a <=( a45793a  and  a45790a );
 a45795a <=( a45794a  and  a45787a );
 a45798a <=( A234  and  (not A233) );
 a45801a <=( A298  and  A235 );
 a45802a <=( a45801a  and  a45798a );
 a45805a <=( (not A300)  and  (not A299) );
 a45808a <=( (not A302)  and  (not A301) );
 a45809a <=( a45808a  and  a45805a );
 a45810a <=( a45809a  and  a45802a );
 a45813a <=( A168  and  (not A170) );
 a45816a <=( (not A166)  and  A167 );
 a45817a <=( a45816a  and  a45813a );
 a45820a <=( (not A202)  and  A201 );
 a45823a <=( A232  and  (not A203) );
 a45824a <=( a45823a  and  a45820a );
 a45825a <=( a45824a  and  a45817a );
 a45828a <=( A234  and  (not A233) );
 a45831a <=( (not A298)  and  A235 );
 a45832a <=( a45831a  and  a45828a );
 a45835a <=( (not A300)  and  A299 );
 a45838a <=( (not A302)  and  (not A301) );
 a45839a <=( a45838a  and  a45835a );
 a45840a <=( a45839a  and  a45832a );
 a45843a <=( A168  and  (not A170) );
 a45846a <=( (not A166)  and  A167 );
 a45847a <=( a45846a  and  a45843a );
 a45850a <=( (not A202)  and  A201 );
 a45853a <=( A232  and  (not A203) );
 a45854a <=( a45853a  and  a45850a );
 a45855a <=( a45854a  and  a45847a );
 a45858a <=( A234  and  (not A233) );
 a45861a <=( (not A265)  and  A235 );
 a45862a <=( a45861a  and  a45858a );
 a45865a <=( (not A267)  and  A266 );
 a45868a <=( (not A269)  and  (not A268) );
 a45869a <=( a45868a  and  a45865a );
 a45870a <=( a45869a  and  a45862a );
 a45873a <=( A168  and  (not A170) );
 a45876a <=( (not A166)  and  A167 );
 a45877a <=( a45876a  and  a45873a );
 a45880a <=( (not A202)  and  A201 );
 a45883a <=( A232  and  (not A203) );
 a45884a <=( a45883a  and  a45880a );
 a45885a <=( a45884a  and  a45877a );
 a45888a <=( A234  and  (not A233) );
 a45891a <=( A265  and  A235 );
 a45892a <=( a45891a  and  a45888a );
 a45895a <=( (not A267)  and  (not A266) );
 a45898a <=( (not A269)  and  (not A268) );
 a45899a <=( a45898a  and  a45895a );
 a45900a <=( a45899a  and  a45892a );
 a45903a <=( A168  and  (not A170) );
 a45906a <=( (not A166)  and  A167 );
 a45907a <=( a45906a  and  a45903a );
 a45910a <=( (not A202)  and  A201 );
 a45913a <=( A232  and  (not A203) );
 a45914a <=( a45913a  and  a45910a );
 a45915a <=( a45914a  and  a45907a );
 a45918a <=( A234  and  (not A233) );
 a45921a <=( A298  and  A236 );
 a45922a <=( a45921a  and  a45918a );
 a45925a <=( (not A300)  and  (not A299) );
 a45928a <=( (not A302)  and  (not A301) );
 a45929a <=( a45928a  and  a45925a );
 a45930a <=( a45929a  and  a45922a );
 a45933a <=( A168  and  (not A170) );
 a45936a <=( (not A166)  and  A167 );
 a45937a <=( a45936a  and  a45933a );
 a45940a <=( (not A202)  and  A201 );
 a45943a <=( A232  and  (not A203) );
 a45944a <=( a45943a  and  a45940a );
 a45945a <=( a45944a  and  a45937a );
 a45948a <=( A234  and  (not A233) );
 a45951a <=( (not A298)  and  A236 );
 a45952a <=( a45951a  and  a45948a );
 a45955a <=( (not A300)  and  A299 );
 a45958a <=( (not A302)  and  (not A301) );
 a45959a <=( a45958a  and  a45955a );
 a45960a <=( a45959a  and  a45952a );
 a45963a <=( A168  and  (not A170) );
 a45966a <=( (not A166)  and  A167 );
 a45967a <=( a45966a  and  a45963a );
 a45970a <=( (not A202)  and  A201 );
 a45973a <=( A232  and  (not A203) );
 a45974a <=( a45973a  and  a45970a );
 a45975a <=( a45974a  and  a45967a );
 a45978a <=( A234  and  (not A233) );
 a45981a <=( (not A265)  and  A236 );
 a45982a <=( a45981a  and  a45978a );
 a45985a <=( (not A267)  and  A266 );
 a45988a <=( (not A269)  and  (not A268) );
 a45989a <=( a45988a  and  a45985a );
 a45990a <=( a45989a  and  a45982a );
 a45993a <=( A168  and  (not A170) );
 a45996a <=( (not A166)  and  A167 );
 a45997a <=( a45996a  and  a45993a );
 a46000a <=( (not A202)  and  A201 );
 a46003a <=( A232  and  (not A203) );
 a46004a <=( a46003a  and  a46000a );
 a46005a <=( a46004a  and  a45997a );
 a46008a <=( A234  and  (not A233) );
 a46011a <=( A265  and  A236 );
 a46012a <=( a46011a  and  a46008a );
 a46015a <=( (not A267)  and  (not A266) );
 a46018a <=( (not A269)  and  (not A268) );
 a46019a <=( a46018a  and  a46015a );
 a46020a <=( a46019a  and  a46012a );
 a46023a <=( A168  and  (not A170) );
 a46026a <=( (not A166)  and  A167 );
 a46027a <=( a46026a  and  a46023a );
 a46030a <=( (not A202)  and  A201 );
 a46033a <=( A232  and  (not A203) );
 a46034a <=( a46033a  and  a46030a );
 a46035a <=( a46034a  and  a46027a );
 a46038a <=( (not A234)  and  (not A233) );
 a46041a <=( (not A236)  and  (not A235) );
 a46042a <=( a46041a  and  a46038a );
 a46045a <=( (not A299)  and  A298 );
 a46048a <=( A301  and  A300 );
 a46049a <=( a46048a  and  a46045a );
 a46050a <=( a46049a  and  a46042a );
 a46053a <=( A168  and  (not A170) );
 a46056a <=( (not A166)  and  A167 );
 a46057a <=( a46056a  and  a46053a );
 a46060a <=( (not A202)  and  A201 );
 a46063a <=( A232  and  (not A203) );
 a46064a <=( a46063a  and  a46060a );
 a46065a <=( a46064a  and  a46057a );
 a46068a <=( (not A234)  and  (not A233) );
 a46071a <=( (not A236)  and  (not A235) );
 a46072a <=( a46071a  and  a46068a );
 a46075a <=( (not A299)  and  A298 );
 a46078a <=( A302  and  A300 );
 a46079a <=( a46078a  and  a46075a );
 a46080a <=( a46079a  and  a46072a );
 a46083a <=( A168  and  (not A170) );
 a46086a <=( (not A166)  and  A167 );
 a46087a <=( a46086a  and  a46083a );
 a46090a <=( (not A202)  and  A201 );
 a46093a <=( A232  and  (not A203) );
 a46094a <=( a46093a  and  a46090a );
 a46095a <=( a46094a  and  a46087a );
 a46098a <=( (not A234)  and  (not A233) );
 a46101a <=( (not A236)  and  (not A235) );
 a46102a <=( a46101a  and  a46098a );
 a46105a <=( A299  and  (not A298) );
 a46108a <=( A301  and  A300 );
 a46109a <=( a46108a  and  a46105a );
 a46110a <=( a46109a  and  a46102a );
 a46113a <=( A168  and  (not A170) );
 a46116a <=( (not A166)  and  A167 );
 a46117a <=( a46116a  and  a46113a );
 a46120a <=( (not A202)  and  A201 );
 a46123a <=( A232  and  (not A203) );
 a46124a <=( a46123a  and  a46120a );
 a46125a <=( a46124a  and  a46117a );
 a46128a <=( (not A234)  and  (not A233) );
 a46131a <=( (not A236)  and  (not A235) );
 a46132a <=( a46131a  and  a46128a );
 a46135a <=( A299  and  (not A298) );
 a46138a <=( A302  and  A300 );
 a46139a <=( a46138a  and  a46135a );
 a46140a <=( a46139a  and  a46132a );
 a46143a <=( A168  and  (not A170) );
 a46146a <=( (not A166)  and  A167 );
 a46147a <=( a46146a  and  a46143a );
 a46150a <=( (not A202)  and  A201 );
 a46153a <=( A232  and  (not A203) );
 a46154a <=( a46153a  and  a46150a );
 a46155a <=( a46154a  and  a46147a );
 a46158a <=( (not A234)  and  (not A233) );
 a46161a <=( (not A236)  and  (not A235) );
 a46162a <=( a46161a  and  a46158a );
 a46165a <=( A266  and  (not A265) );
 a46168a <=( A268  and  A267 );
 a46169a <=( a46168a  and  a46165a );
 a46170a <=( a46169a  and  a46162a );
 a46173a <=( A168  and  (not A170) );
 a46176a <=( (not A166)  and  A167 );
 a46177a <=( a46176a  and  a46173a );
 a46180a <=( (not A202)  and  A201 );
 a46183a <=( A232  and  (not A203) );
 a46184a <=( a46183a  and  a46180a );
 a46185a <=( a46184a  and  a46177a );
 a46188a <=( (not A234)  and  (not A233) );
 a46191a <=( (not A236)  and  (not A235) );
 a46192a <=( a46191a  and  a46188a );
 a46195a <=( A266  and  (not A265) );
 a46198a <=( A269  and  A267 );
 a46199a <=( a46198a  and  a46195a );
 a46200a <=( a46199a  and  a46192a );
 a46203a <=( A168  and  (not A170) );
 a46206a <=( (not A166)  and  A167 );
 a46207a <=( a46206a  and  a46203a );
 a46210a <=( (not A202)  and  A201 );
 a46213a <=( A232  and  (not A203) );
 a46214a <=( a46213a  and  a46210a );
 a46215a <=( a46214a  and  a46207a );
 a46218a <=( (not A234)  and  (not A233) );
 a46221a <=( (not A236)  and  (not A235) );
 a46222a <=( a46221a  and  a46218a );
 a46225a <=( (not A266)  and  A265 );
 a46228a <=( A268  and  A267 );
 a46229a <=( a46228a  and  a46225a );
 a46230a <=( a46229a  and  a46222a );
 a46233a <=( A168  and  (not A170) );
 a46236a <=( (not A166)  and  A167 );
 a46237a <=( a46236a  and  a46233a );
 a46240a <=( (not A202)  and  A201 );
 a46243a <=( A232  and  (not A203) );
 a46244a <=( a46243a  and  a46240a );
 a46245a <=( a46244a  and  a46237a );
 a46248a <=( (not A234)  and  (not A233) );
 a46251a <=( (not A236)  and  (not A235) );
 a46252a <=( a46251a  and  a46248a );
 a46255a <=( (not A266)  and  A265 );
 a46258a <=( A269  and  A267 );
 a46259a <=( a46258a  and  a46255a );
 a46260a <=( a46259a  and  a46252a );
 a46263a <=( A168  and  (not A170) );
 a46266a <=( (not A166)  and  A167 );
 a46267a <=( a46266a  and  a46263a );
 a46270a <=( A202  and  (not A201) );
 a46273a <=( A233  and  (not A232) );
 a46274a <=( a46273a  and  a46270a );
 a46275a <=( a46274a  and  a46267a );
 a46278a <=( (not A235)  and  (not A234) );
 a46281a <=( A298  and  (not A236) );
 a46282a <=( a46281a  and  a46278a );
 a46285a <=( (not A300)  and  (not A299) );
 a46288a <=( (not A302)  and  (not A301) );
 a46289a <=( a46288a  and  a46285a );
 a46290a <=( a46289a  and  a46282a );
 a46293a <=( A168  and  (not A170) );
 a46296a <=( (not A166)  and  A167 );
 a46297a <=( a46296a  and  a46293a );
 a46300a <=( A202  and  (not A201) );
 a46303a <=( A233  and  (not A232) );
 a46304a <=( a46303a  and  a46300a );
 a46305a <=( a46304a  and  a46297a );
 a46308a <=( (not A235)  and  (not A234) );
 a46311a <=( (not A298)  and  (not A236) );
 a46312a <=( a46311a  and  a46308a );
 a46315a <=( (not A300)  and  A299 );
 a46318a <=( (not A302)  and  (not A301) );
 a46319a <=( a46318a  and  a46315a );
 a46320a <=( a46319a  and  a46312a );
 a46323a <=( A168  and  (not A170) );
 a46326a <=( (not A166)  and  A167 );
 a46327a <=( a46326a  and  a46323a );
 a46330a <=( A202  and  (not A201) );
 a46333a <=( A233  and  (not A232) );
 a46334a <=( a46333a  and  a46330a );
 a46335a <=( a46334a  and  a46327a );
 a46338a <=( (not A235)  and  (not A234) );
 a46341a <=( (not A265)  and  (not A236) );
 a46342a <=( a46341a  and  a46338a );
 a46345a <=( (not A267)  and  A266 );
 a46348a <=( (not A269)  and  (not A268) );
 a46349a <=( a46348a  and  a46345a );
 a46350a <=( a46349a  and  a46342a );
 a46353a <=( A168  and  (not A170) );
 a46356a <=( (not A166)  and  A167 );
 a46357a <=( a46356a  and  a46353a );
 a46360a <=( A202  and  (not A201) );
 a46363a <=( A233  and  (not A232) );
 a46364a <=( a46363a  and  a46360a );
 a46365a <=( a46364a  and  a46357a );
 a46368a <=( (not A235)  and  (not A234) );
 a46371a <=( A265  and  (not A236) );
 a46372a <=( a46371a  and  a46368a );
 a46375a <=( (not A267)  and  (not A266) );
 a46378a <=( (not A269)  and  (not A268) );
 a46379a <=( a46378a  and  a46375a );
 a46380a <=( a46379a  and  a46372a );
 a46383a <=( A168  and  (not A170) );
 a46386a <=( (not A166)  and  A167 );
 a46387a <=( a46386a  and  a46383a );
 a46390a <=( A202  and  (not A201) );
 a46393a <=( (not A233)  and  A232 );
 a46394a <=( a46393a  and  a46390a );
 a46395a <=( a46394a  and  a46387a );
 a46398a <=( (not A235)  and  (not A234) );
 a46401a <=( A298  and  (not A236) );
 a46402a <=( a46401a  and  a46398a );
 a46405a <=( (not A300)  and  (not A299) );
 a46408a <=( (not A302)  and  (not A301) );
 a46409a <=( a46408a  and  a46405a );
 a46410a <=( a46409a  and  a46402a );
 a46413a <=( A168  and  (not A170) );
 a46416a <=( (not A166)  and  A167 );
 a46417a <=( a46416a  and  a46413a );
 a46420a <=( A202  and  (not A201) );
 a46423a <=( (not A233)  and  A232 );
 a46424a <=( a46423a  and  a46420a );
 a46425a <=( a46424a  and  a46417a );
 a46428a <=( (not A235)  and  (not A234) );
 a46431a <=( (not A298)  and  (not A236) );
 a46432a <=( a46431a  and  a46428a );
 a46435a <=( (not A300)  and  A299 );
 a46438a <=( (not A302)  and  (not A301) );
 a46439a <=( a46438a  and  a46435a );
 a46440a <=( a46439a  and  a46432a );
 a46443a <=( A168  and  (not A170) );
 a46446a <=( (not A166)  and  A167 );
 a46447a <=( a46446a  and  a46443a );
 a46450a <=( A202  and  (not A201) );
 a46453a <=( (not A233)  and  A232 );
 a46454a <=( a46453a  and  a46450a );
 a46455a <=( a46454a  and  a46447a );
 a46458a <=( (not A235)  and  (not A234) );
 a46461a <=( (not A265)  and  (not A236) );
 a46462a <=( a46461a  and  a46458a );
 a46465a <=( (not A267)  and  A266 );
 a46468a <=( (not A269)  and  (not A268) );
 a46469a <=( a46468a  and  a46465a );
 a46470a <=( a46469a  and  a46462a );
 a46473a <=( A168  and  (not A170) );
 a46476a <=( (not A166)  and  A167 );
 a46477a <=( a46476a  and  a46473a );
 a46480a <=( A202  and  (not A201) );
 a46483a <=( (not A233)  and  A232 );
 a46484a <=( a46483a  and  a46480a );
 a46485a <=( a46484a  and  a46477a );
 a46488a <=( (not A235)  and  (not A234) );
 a46491a <=( A265  and  (not A236) );
 a46492a <=( a46491a  and  a46488a );
 a46495a <=( (not A267)  and  (not A266) );
 a46498a <=( (not A269)  and  (not A268) );
 a46499a <=( a46498a  and  a46495a );
 a46500a <=( a46499a  and  a46492a );
 a46503a <=( A168  and  (not A170) );
 a46506a <=( (not A166)  and  A167 );
 a46507a <=( a46506a  and  a46503a );
 a46510a <=( A203  and  (not A201) );
 a46513a <=( A233  and  (not A232) );
 a46514a <=( a46513a  and  a46510a );
 a46515a <=( a46514a  and  a46507a );
 a46518a <=( (not A235)  and  (not A234) );
 a46521a <=( A298  and  (not A236) );
 a46522a <=( a46521a  and  a46518a );
 a46525a <=( (not A300)  and  (not A299) );
 a46528a <=( (not A302)  and  (not A301) );
 a46529a <=( a46528a  and  a46525a );
 a46530a <=( a46529a  and  a46522a );
 a46533a <=( A168  and  (not A170) );
 a46536a <=( (not A166)  and  A167 );
 a46537a <=( a46536a  and  a46533a );
 a46540a <=( A203  and  (not A201) );
 a46543a <=( A233  and  (not A232) );
 a46544a <=( a46543a  and  a46540a );
 a46545a <=( a46544a  and  a46537a );
 a46548a <=( (not A235)  and  (not A234) );
 a46551a <=( (not A298)  and  (not A236) );
 a46552a <=( a46551a  and  a46548a );
 a46555a <=( (not A300)  and  A299 );
 a46558a <=( (not A302)  and  (not A301) );
 a46559a <=( a46558a  and  a46555a );
 a46560a <=( a46559a  and  a46552a );
 a46563a <=( A168  and  (not A170) );
 a46566a <=( (not A166)  and  A167 );
 a46567a <=( a46566a  and  a46563a );
 a46570a <=( A203  and  (not A201) );
 a46573a <=( A233  and  (not A232) );
 a46574a <=( a46573a  and  a46570a );
 a46575a <=( a46574a  and  a46567a );
 a46578a <=( (not A235)  and  (not A234) );
 a46581a <=( (not A265)  and  (not A236) );
 a46582a <=( a46581a  and  a46578a );
 a46585a <=( (not A267)  and  A266 );
 a46588a <=( (not A269)  and  (not A268) );
 a46589a <=( a46588a  and  a46585a );
 a46590a <=( a46589a  and  a46582a );
 a46593a <=( A168  and  (not A170) );
 a46596a <=( (not A166)  and  A167 );
 a46597a <=( a46596a  and  a46593a );
 a46600a <=( A203  and  (not A201) );
 a46603a <=( A233  and  (not A232) );
 a46604a <=( a46603a  and  a46600a );
 a46605a <=( a46604a  and  a46597a );
 a46608a <=( (not A235)  and  (not A234) );
 a46611a <=( A265  and  (not A236) );
 a46612a <=( a46611a  and  a46608a );
 a46615a <=( (not A267)  and  (not A266) );
 a46618a <=( (not A269)  and  (not A268) );
 a46619a <=( a46618a  and  a46615a );
 a46620a <=( a46619a  and  a46612a );
 a46623a <=( A168  and  (not A170) );
 a46626a <=( (not A166)  and  A167 );
 a46627a <=( a46626a  and  a46623a );
 a46630a <=( A203  and  (not A201) );
 a46633a <=( (not A233)  and  A232 );
 a46634a <=( a46633a  and  a46630a );
 a46635a <=( a46634a  and  a46627a );
 a46638a <=( (not A235)  and  (not A234) );
 a46641a <=( A298  and  (not A236) );
 a46642a <=( a46641a  and  a46638a );
 a46645a <=( (not A300)  and  (not A299) );
 a46648a <=( (not A302)  and  (not A301) );
 a46649a <=( a46648a  and  a46645a );
 a46650a <=( a46649a  and  a46642a );
 a46653a <=( A168  and  (not A170) );
 a46656a <=( (not A166)  and  A167 );
 a46657a <=( a46656a  and  a46653a );
 a46660a <=( A203  and  (not A201) );
 a46663a <=( (not A233)  and  A232 );
 a46664a <=( a46663a  and  a46660a );
 a46665a <=( a46664a  and  a46657a );
 a46668a <=( (not A235)  and  (not A234) );
 a46671a <=( (not A298)  and  (not A236) );
 a46672a <=( a46671a  and  a46668a );
 a46675a <=( (not A300)  and  A299 );
 a46678a <=( (not A302)  and  (not A301) );
 a46679a <=( a46678a  and  a46675a );
 a46680a <=( a46679a  and  a46672a );
 a46683a <=( A168  and  (not A170) );
 a46686a <=( (not A166)  and  A167 );
 a46687a <=( a46686a  and  a46683a );
 a46690a <=( A203  and  (not A201) );
 a46693a <=( (not A233)  and  A232 );
 a46694a <=( a46693a  and  a46690a );
 a46695a <=( a46694a  and  a46687a );
 a46698a <=( (not A235)  and  (not A234) );
 a46701a <=( (not A265)  and  (not A236) );
 a46702a <=( a46701a  and  a46698a );
 a46705a <=( (not A267)  and  A266 );
 a46708a <=( (not A269)  and  (not A268) );
 a46709a <=( a46708a  and  a46705a );
 a46710a <=( a46709a  and  a46702a );
 a46713a <=( A168  and  (not A170) );
 a46716a <=( (not A166)  and  A167 );
 a46717a <=( a46716a  and  a46713a );
 a46720a <=( A203  and  (not A201) );
 a46723a <=( (not A233)  and  A232 );
 a46724a <=( a46723a  and  a46720a );
 a46725a <=( a46724a  and  a46717a );
 a46728a <=( (not A235)  and  (not A234) );
 a46731a <=( A265  and  (not A236) );
 a46732a <=( a46731a  and  a46728a );
 a46735a <=( (not A267)  and  (not A266) );
 a46738a <=( (not A269)  and  (not A268) );
 a46739a <=( a46738a  and  a46735a );
 a46740a <=( a46739a  and  a46732a );
 a46743a <=( A168  and  (not A170) );
 a46746a <=( (not A166)  and  A167 );
 a46747a <=( a46746a  and  a46743a );
 a46750a <=( A200  and  A199 );
 a46753a <=( A233  and  (not A232) );
 a46754a <=( a46753a  and  a46750a );
 a46755a <=( a46754a  and  a46747a );
 a46758a <=( (not A235)  and  (not A234) );
 a46761a <=( A298  and  (not A236) );
 a46762a <=( a46761a  and  a46758a );
 a46765a <=( (not A300)  and  (not A299) );
 a46768a <=( (not A302)  and  (not A301) );
 a46769a <=( a46768a  and  a46765a );
 a46770a <=( a46769a  and  a46762a );
 a46773a <=( A168  and  (not A170) );
 a46776a <=( (not A166)  and  A167 );
 a46777a <=( a46776a  and  a46773a );
 a46780a <=( A200  and  A199 );
 a46783a <=( A233  and  (not A232) );
 a46784a <=( a46783a  and  a46780a );
 a46785a <=( a46784a  and  a46777a );
 a46788a <=( (not A235)  and  (not A234) );
 a46791a <=( (not A298)  and  (not A236) );
 a46792a <=( a46791a  and  a46788a );
 a46795a <=( (not A300)  and  A299 );
 a46798a <=( (not A302)  and  (not A301) );
 a46799a <=( a46798a  and  a46795a );
 a46800a <=( a46799a  and  a46792a );
 a46803a <=( A168  and  (not A170) );
 a46806a <=( (not A166)  and  A167 );
 a46807a <=( a46806a  and  a46803a );
 a46810a <=( A200  and  A199 );
 a46813a <=( A233  and  (not A232) );
 a46814a <=( a46813a  and  a46810a );
 a46815a <=( a46814a  and  a46807a );
 a46818a <=( (not A235)  and  (not A234) );
 a46821a <=( (not A265)  and  (not A236) );
 a46822a <=( a46821a  and  a46818a );
 a46825a <=( (not A267)  and  A266 );
 a46828a <=( (not A269)  and  (not A268) );
 a46829a <=( a46828a  and  a46825a );
 a46830a <=( a46829a  and  a46822a );
 a46833a <=( A168  and  (not A170) );
 a46836a <=( (not A166)  and  A167 );
 a46837a <=( a46836a  and  a46833a );
 a46840a <=( A200  and  A199 );
 a46843a <=( A233  and  (not A232) );
 a46844a <=( a46843a  and  a46840a );
 a46845a <=( a46844a  and  a46837a );
 a46848a <=( (not A235)  and  (not A234) );
 a46851a <=( A265  and  (not A236) );
 a46852a <=( a46851a  and  a46848a );
 a46855a <=( (not A267)  and  (not A266) );
 a46858a <=( (not A269)  and  (not A268) );
 a46859a <=( a46858a  and  a46855a );
 a46860a <=( a46859a  and  a46852a );
 a46863a <=( A168  and  (not A170) );
 a46866a <=( (not A166)  and  A167 );
 a46867a <=( a46866a  and  a46863a );
 a46870a <=( A200  and  A199 );
 a46873a <=( (not A233)  and  A232 );
 a46874a <=( a46873a  and  a46870a );
 a46875a <=( a46874a  and  a46867a );
 a46878a <=( (not A235)  and  (not A234) );
 a46881a <=( A298  and  (not A236) );
 a46882a <=( a46881a  and  a46878a );
 a46885a <=( (not A300)  and  (not A299) );
 a46888a <=( (not A302)  and  (not A301) );
 a46889a <=( a46888a  and  a46885a );
 a46890a <=( a46889a  and  a46882a );
 a46893a <=( A168  and  (not A170) );
 a46896a <=( (not A166)  and  A167 );
 a46897a <=( a46896a  and  a46893a );
 a46900a <=( A200  and  A199 );
 a46903a <=( (not A233)  and  A232 );
 a46904a <=( a46903a  and  a46900a );
 a46905a <=( a46904a  and  a46897a );
 a46908a <=( (not A235)  and  (not A234) );
 a46911a <=( (not A298)  and  (not A236) );
 a46912a <=( a46911a  and  a46908a );
 a46915a <=( (not A300)  and  A299 );
 a46918a <=( (not A302)  and  (not A301) );
 a46919a <=( a46918a  and  a46915a );
 a46920a <=( a46919a  and  a46912a );
 a46923a <=( A168  and  (not A170) );
 a46926a <=( (not A166)  and  A167 );
 a46927a <=( a46926a  and  a46923a );
 a46930a <=( A200  and  A199 );
 a46933a <=( (not A233)  and  A232 );
 a46934a <=( a46933a  and  a46930a );
 a46935a <=( a46934a  and  a46927a );
 a46938a <=( (not A235)  and  (not A234) );
 a46941a <=( (not A265)  and  (not A236) );
 a46942a <=( a46941a  and  a46938a );
 a46945a <=( (not A267)  and  A266 );
 a46948a <=( (not A269)  and  (not A268) );
 a46949a <=( a46948a  and  a46945a );
 a46950a <=( a46949a  and  a46942a );
 a46953a <=( A168  and  (not A170) );
 a46956a <=( (not A166)  and  A167 );
 a46957a <=( a46956a  and  a46953a );
 a46960a <=( A200  and  A199 );
 a46963a <=( (not A233)  and  A232 );
 a46964a <=( a46963a  and  a46960a );
 a46965a <=( a46964a  and  a46957a );
 a46968a <=( (not A235)  and  (not A234) );
 a46971a <=( A265  and  (not A236) );
 a46972a <=( a46971a  and  a46968a );
 a46975a <=( (not A267)  and  (not A266) );
 a46978a <=( (not A269)  and  (not A268) );
 a46979a <=( a46978a  and  a46975a );
 a46980a <=( a46979a  and  a46972a );
 a46983a <=( A168  and  (not A170) );
 a46986a <=( (not A166)  and  A167 );
 a46987a <=( a46986a  and  a46983a );
 a46990a <=( (not A200)  and  (not A199) );
 a46993a <=( A233  and  (not A232) );
 a46994a <=( a46993a  and  a46990a );
 a46995a <=( a46994a  and  a46987a );
 a46998a <=( (not A235)  and  (not A234) );
 a47001a <=( A298  and  (not A236) );
 a47002a <=( a47001a  and  a46998a );
 a47005a <=( (not A300)  and  (not A299) );
 a47008a <=( (not A302)  and  (not A301) );
 a47009a <=( a47008a  and  a47005a );
 a47010a <=( a47009a  and  a47002a );
 a47013a <=( A168  and  (not A170) );
 a47016a <=( (not A166)  and  A167 );
 a47017a <=( a47016a  and  a47013a );
 a47020a <=( (not A200)  and  (not A199) );
 a47023a <=( A233  and  (not A232) );
 a47024a <=( a47023a  and  a47020a );
 a47025a <=( a47024a  and  a47017a );
 a47028a <=( (not A235)  and  (not A234) );
 a47031a <=( (not A298)  and  (not A236) );
 a47032a <=( a47031a  and  a47028a );
 a47035a <=( (not A300)  and  A299 );
 a47038a <=( (not A302)  and  (not A301) );
 a47039a <=( a47038a  and  a47035a );
 a47040a <=( a47039a  and  a47032a );
 a47043a <=( A168  and  (not A170) );
 a47046a <=( (not A166)  and  A167 );
 a47047a <=( a47046a  and  a47043a );
 a47050a <=( (not A200)  and  (not A199) );
 a47053a <=( A233  and  (not A232) );
 a47054a <=( a47053a  and  a47050a );
 a47055a <=( a47054a  and  a47047a );
 a47058a <=( (not A235)  and  (not A234) );
 a47061a <=( (not A265)  and  (not A236) );
 a47062a <=( a47061a  and  a47058a );
 a47065a <=( (not A267)  and  A266 );
 a47068a <=( (not A269)  and  (not A268) );
 a47069a <=( a47068a  and  a47065a );
 a47070a <=( a47069a  and  a47062a );
 a47073a <=( A168  and  (not A170) );
 a47076a <=( (not A166)  and  A167 );
 a47077a <=( a47076a  and  a47073a );
 a47080a <=( (not A200)  and  (not A199) );
 a47083a <=( A233  and  (not A232) );
 a47084a <=( a47083a  and  a47080a );
 a47085a <=( a47084a  and  a47077a );
 a47088a <=( (not A235)  and  (not A234) );
 a47091a <=( A265  and  (not A236) );
 a47092a <=( a47091a  and  a47088a );
 a47095a <=( (not A267)  and  (not A266) );
 a47098a <=( (not A269)  and  (not A268) );
 a47099a <=( a47098a  and  a47095a );
 a47100a <=( a47099a  and  a47092a );
 a47103a <=( A168  and  (not A170) );
 a47106a <=( (not A166)  and  A167 );
 a47107a <=( a47106a  and  a47103a );
 a47110a <=( (not A200)  and  (not A199) );
 a47113a <=( (not A233)  and  A232 );
 a47114a <=( a47113a  and  a47110a );
 a47115a <=( a47114a  and  a47107a );
 a47118a <=( (not A235)  and  (not A234) );
 a47121a <=( A298  and  (not A236) );
 a47122a <=( a47121a  and  a47118a );
 a47125a <=( (not A300)  and  (not A299) );
 a47128a <=( (not A302)  and  (not A301) );
 a47129a <=( a47128a  and  a47125a );
 a47130a <=( a47129a  and  a47122a );
 a47133a <=( A168  and  (not A170) );
 a47136a <=( (not A166)  and  A167 );
 a47137a <=( a47136a  and  a47133a );
 a47140a <=( (not A200)  and  (not A199) );
 a47143a <=( (not A233)  and  A232 );
 a47144a <=( a47143a  and  a47140a );
 a47145a <=( a47144a  and  a47137a );
 a47148a <=( (not A235)  and  (not A234) );
 a47151a <=( (not A298)  and  (not A236) );
 a47152a <=( a47151a  and  a47148a );
 a47155a <=( (not A300)  and  A299 );
 a47158a <=( (not A302)  and  (not A301) );
 a47159a <=( a47158a  and  a47155a );
 a47160a <=( a47159a  and  a47152a );
 a47163a <=( A168  and  (not A170) );
 a47166a <=( (not A166)  and  A167 );
 a47167a <=( a47166a  and  a47163a );
 a47170a <=( (not A200)  and  (not A199) );
 a47173a <=( (not A233)  and  A232 );
 a47174a <=( a47173a  and  a47170a );
 a47175a <=( a47174a  and  a47167a );
 a47178a <=( (not A235)  and  (not A234) );
 a47181a <=( (not A265)  and  (not A236) );
 a47182a <=( a47181a  and  a47178a );
 a47185a <=( (not A267)  and  A266 );
 a47188a <=( (not A269)  and  (not A268) );
 a47189a <=( a47188a  and  a47185a );
 a47190a <=( a47189a  and  a47182a );
 a47193a <=( A168  and  (not A170) );
 a47196a <=( (not A166)  and  A167 );
 a47197a <=( a47196a  and  a47193a );
 a47200a <=( (not A200)  and  (not A199) );
 a47203a <=( (not A233)  and  A232 );
 a47204a <=( a47203a  and  a47200a );
 a47205a <=( a47204a  and  a47197a );
 a47208a <=( (not A235)  and  (not A234) );
 a47211a <=( A265  and  (not A236) );
 a47212a <=( a47211a  and  a47208a );
 a47215a <=( (not A267)  and  (not A266) );
 a47218a <=( (not A269)  and  (not A268) );
 a47219a <=( a47218a  and  a47215a );
 a47220a <=( a47219a  and  a47212a );
 a47223a <=( A168  and  (not A170) );
 a47226a <=( A166  and  (not A167) );
 a47227a <=( a47226a  and  a47223a );
 a47230a <=( (not A202)  and  A201 );
 a47233a <=( (not A232)  and  (not A203) );
 a47234a <=( a47233a  and  a47230a );
 a47235a <=( a47234a  and  a47227a );
 a47238a <=( A234  and  A233 );
 a47241a <=( A298  and  A235 );
 a47242a <=( a47241a  and  a47238a );
 a47245a <=( (not A300)  and  (not A299) );
 a47248a <=( (not A302)  and  (not A301) );
 a47249a <=( a47248a  and  a47245a );
 a47250a <=( a47249a  and  a47242a );
 a47253a <=( A168  and  (not A170) );
 a47256a <=( A166  and  (not A167) );
 a47257a <=( a47256a  and  a47253a );
 a47260a <=( (not A202)  and  A201 );
 a47263a <=( (not A232)  and  (not A203) );
 a47264a <=( a47263a  and  a47260a );
 a47265a <=( a47264a  and  a47257a );
 a47268a <=( A234  and  A233 );
 a47271a <=( (not A298)  and  A235 );
 a47272a <=( a47271a  and  a47268a );
 a47275a <=( (not A300)  and  A299 );
 a47278a <=( (not A302)  and  (not A301) );
 a47279a <=( a47278a  and  a47275a );
 a47280a <=( a47279a  and  a47272a );
 a47283a <=( A168  and  (not A170) );
 a47286a <=( A166  and  (not A167) );
 a47287a <=( a47286a  and  a47283a );
 a47290a <=( (not A202)  and  A201 );
 a47293a <=( (not A232)  and  (not A203) );
 a47294a <=( a47293a  and  a47290a );
 a47295a <=( a47294a  and  a47287a );
 a47298a <=( A234  and  A233 );
 a47301a <=( (not A265)  and  A235 );
 a47302a <=( a47301a  and  a47298a );
 a47305a <=( (not A267)  and  A266 );
 a47308a <=( (not A269)  and  (not A268) );
 a47309a <=( a47308a  and  a47305a );
 a47310a <=( a47309a  and  a47302a );
 a47313a <=( A168  and  (not A170) );
 a47316a <=( A166  and  (not A167) );
 a47317a <=( a47316a  and  a47313a );
 a47320a <=( (not A202)  and  A201 );
 a47323a <=( (not A232)  and  (not A203) );
 a47324a <=( a47323a  and  a47320a );
 a47325a <=( a47324a  and  a47317a );
 a47328a <=( A234  and  A233 );
 a47331a <=( A265  and  A235 );
 a47332a <=( a47331a  and  a47328a );
 a47335a <=( (not A267)  and  (not A266) );
 a47338a <=( (not A269)  and  (not A268) );
 a47339a <=( a47338a  and  a47335a );
 a47340a <=( a47339a  and  a47332a );
 a47343a <=( A168  and  (not A170) );
 a47346a <=( A166  and  (not A167) );
 a47347a <=( a47346a  and  a47343a );
 a47350a <=( (not A202)  and  A201 );
 a47353a <=( (not A232)  and  (not A203) );
 a47354a <=( a47353a  and  a47350a );
 a47355a <=( a47354a  and  a47347a );
 a47358a <=( A234  and  A233 );
 a47361a <=( A298  and  A236 );
 a47362a <=( a47361a  and  a47358a );
 a47365a <=( (not A300)  and  (not A299) );
 a47368a <=( (not A302)  and  (not A301) );
 a47369a <=( a47368a  and  a47365a );
 a47370a <=( a47369a  and  a47362a );
 a47373a <=( A168  and  (not A170) );
 a47376a <=( A166  and  (not A167) );
 a47377a <=( a47376a  and  a47373a );
 a47380a <=( (not A202)  and  A201 );
 a47383a <=( (not A232)  and  (not A203) );
 a47384a <=( a47383a  and  a47380a );
 a47385a <=( a47384a  and  a47377a );
 a47388a <=( A234  and  A233 );
 a47391a <=( (not A298)  and  A236 );
 a47392a <=( a47391a  and  a47388a );
 a47395a <=( (not A300)  and  A299 );
 a47398a <=( (not A302)  and  (not A301) );
 a47399a <=( a47398a  and  a47395a );
 a47400a <=( a47399a  and  a47392a );
 a47403a <=( A168  and  (not A170) );
 a47406a <=( A166  and  (not A167) );
 a47407a <=( a47406a  and  a47403a );
 a47410a <=( (not A202)  and  A201 );
 a47413a <=( (not A232)  and  (not A203) );
 a47414a <=( a47413a  and  a47410a );
 a47415a <=( a47414a  and  a47407a );
 a47418a <=( A234  and  A233 );
 a47421a <=( (not A265)  and  A236 );
 a47422a <=( a47421a  and  a47418a );
 a47425a <=( (not A267)  and  A266 );
 a47428a <=( (not A269)  and  (not A268) );
 a47429a <=( a47428a  and  a47425a );
 a47430a <=( a47429a  and  a47422a );
 a47433a <=( A168  and  (not A170) );
 a47436a <=( A166  and  (not A167) );
 a47437a <=( a47436a  and  a47433a );
 a47440a <=( (not A202)  and  A201 );
 a47443a <=( (not A232)  and  (not A203) );
 a47444a <=( a47443a  and  a47440a );
 a47445a <=( a47444a  and  a47437a );
 a47448a <=( A234  and  A233 );
 a47451a <=( A265  and  A236 );
 a47452a <=( a47451a  and  a47448a );
 a47455a <=( (not A267)  and  (not A266) );
 a47458a <=( (not A269)  and  (not A268) );
 a47459a <=( a47458a  and  a47455a );
 a47460a <=( a47459a  and  a47452a );
 a47463a <=( A168  and  (not A170) );
 a47466a <=( A166  and  (not A167) );
 a47467a <=( a47466a  and  a47463a );
 a47470a <=( (not A202)  and  A201 );
 a47473a <=( (not A232)  and  (not A203) );
 a47474a <=( a47473a  and  a47470a );
 a47475a <=( a47474a  and  a47467a );
 a47478a <=( (not A234)  and  A233 );
 a47481a <=( (not A236)  and  (not A235) );
 a47482a <=( a47481a  and  a47478a );
 a47485a <=( (not A299)  and  A298 );
 a47488a <=( A301  and  A300 );
 a47489a <=( a47488a  and  a47485a );
 a47490a <=( a47489a  and  a47482a );
 a47493a <=( A168  and  (not A170) );
 a47496a <=( A166  and  (not A167) );
 a47497a <=( a47496a  and  a47493a );
 a47500a <=( (not A202)  and  A201 );
 a47503a <=( (not A232)  and  (not A203) );
 a47504a <=( a47503a  and  a47500a );
 a47505a <=( a47504a  and  a47497a );
 a47508a <=( (not A234)  and  A233 );
 a47511a <=( (not A236)  and  (not A235) );
 a47512a <=( a47511a  and  a47508a );
 a47515a <=( (not A299)  and  A298 );
 a47518a <=( A302  and  A300 );
 a47519a <=( a47518a  and  a47515a );
 a47520a <=( a47519a  and  a47512a );
 a47523a <=( A168  and  (not A170) );
 a47526a <=( A166  and  (not A167) );
 a47527a <=( a47526a  and  a47523a );
 a47530a <=( (not A202)  and  A201 );
 a47533a <=( (not A232)  and  (not A203) );
 a47534a <=( a47533a  and  a47530a );
 a47535a <=( a47534a  and  a47527a );
 a47538a <=( (not A234)  and  A233 );
 a47541a <=( (not A236)  and  (not A235) );
 a47542a <=( a47541a  and  a47538a );
 a47545a <=( A299  and  (not A298) );
 a47548a <=( A301  and  A300 );
 a47549a <=( a47548a  and  a47545a );
 a47550a <=( a47549a  and  a47542a );
 a47553a <=( A168  and  (not A170) );
 a47556a <=( A166  and  (not A167) );
 a47557a <=( a47556a  and  a47553a );
 a47560a <=( (not A202)  and  A201 );
 a47563a <=( (not A232)  and  (not A203) );
 a47564a <=( a47563a  and  a47560a );
 a47565a <=( a47564a  and  a47557a );
 a47568a <=( (not A234)  and  A233 );
 a47571a <=( (not A236)  and  (not A235) );
 a47572a <=( a47571a  and  a47568a );
 a47575a <=( A299  and  (not A298) );
 a47578a <=( A302  and  A300 );
 a47579a <=( a47578a  and  a47575a );
 a47580a <=( a47579a  and  a47572a );
 a47583a <=( A168  and  (not A170) );
 a47586a <=( A166  and  (not A167) );
 a47587a <=( a47586a  and  a47583a );
 a47590a <=( (not A202)  and  A201 );
 a47593a <=( (not A232)  and  (not A203) );
 a47594a <=( a47593a  and  a47590a );
 a47595a <=( a47594a  and  a47587a );
 a47598a <=( (not A234)  and  A233 );
 a47601a <=( (not A236)  and  (not A235) );
 a47602a <=( a47601a  and  a47598a );
 a47605a <=( A266  and  (not A265) );
 a47608a <=( A268  and  A267 );
 a47609a <=( a47608a  and  a47605a );
 a47610a <=( a47609a  and  a47602a );
 a47613a <=( A168  and  (not A170) );
 a47616a <=( A166  and  (not A167) );
 a47617a <=( a47616a  and  a47613a );
 a47620a <=( (not A202)  and  A201 );
 a47623a <=( (not A232)  and  (not A203) );
 a47624a <=( a47623a  and  a47620a );
 a47625a <=( a47624a  and  a47617a );
 a47628a <=( (not A234)  and  A233 );
 a47631a <=( (not A236)  and  (not A235) );
 a47632a <=( a47631a  and  a47628a );
 a47635a <=( A266  and  (not A265) );
 a47638a <=( A269  and  A267 );
 a47639a <=( a47638a  and  a47635a );
 a47640a <=( a47639a  and  a47632a );
 a47643a <=( A168  and  (not A170) );
 a47646a <=( A166  and  (not A167) );
 a47647a <=( a47646a  and  a47643a );
 a47650a <=( (not A202)  and  A201 );
 a47653a <=( (not A232)  and  (not A203) );
 a47654a <=( a47653a  and  a47650a );
 a47655a <=( a47654a  and  a47647a );
 a47658a <=( (not A234)  and  A233 );
 a47661a <=( (not A236)  and  (not A235) );
 a47662a <=( a47661a  and  a47658a );
 a47665a <=( (not A266)  and  A265 );
 a47668a <=( A268  and  A267 );
 a47669a <=( a47668a  and  a47665a );
 a47670a <=( a47669a  and  a47662a );
 a47673a <=( A168  and  (not A170) );
 a47676a <=( A166  and  (not A167) );
 a47677a <=( a47676a  and  a47673a );
 a47680a <=( (not A202)  and  A201 );
 a47683a <=( (not A232)  and  (not A203) );
 a47684a <=( a47683a  and  a47680a );
 a47685a <=( a47684a  and  a47677a );
 a47688a <=( (not A234)  and  A233 );
 a47691a <=( (not A236)  and  (not A235) );
 a47692a <=( a47691a  and  a47688a );
 a47695a <=( (not A266)  and  A265 );
 a47698a <=( A269  and  A267 );
 a47699a <=( a47698a  and  a47695a );
 a47700a <=( a47699a  and  a47692a );
 a47703a <=( A168  and  (not A170) );
 a47706a <=( A166  and  (not A167) );
 a47707a <=( a47706a  and  a47703a );
 a47710a <=( (not A202)  and  A201 );
 a47713a <=( A232  and  (not A203) );
 a47714a <=( a47713a  and  a47710a );
 a47715a <=( a47714a  and  a47707a );
 a47718a <=( A234  and  (not A233) );
 a47721a <=( A298  and  A235 );
 a47722a <=( a47721a  and  a47718a );
 a47725a <=( (not A300)  and  (not A299) );
 a47728a <=( (not A302)  and  (not A301) );
 a47729a <=( a47728a  and  a47725a );
 a47730a <=( a47729a  and  a47722a );
 a47733a <=( A168  and  (not A170) );
 a47736a <=( A166  and  (not A167) );
 a47737a <=( a47736a  and  a47733a );
 a47740a <=( (not A202)  and  A201 );
 a47743a <=( A232  and  (not A203) );
 a47744a <=( a47743a  and  a47740a );
 a47745a <=( a47744a  and  a47737a );
 a47748a <=( A234  and  (not A233) );
 a47751a <=( (not A298)  and  A235 );
 a47752a <=( a47751a  and  a47748a );
 a47755a <=( (not A300)  and  A299 );
 a47758a <=( (not A302)  and  (not A301) );
 a47759a <=( a47758a  and  a47755a );
 a47760a <=( a47759a  and  a47752a );
 a47763a <=( A168  and  (not A170) );
 a47766a <=( A166  and  (not A167) );
 a47767a <=( a47766a  and  a47763a );
 a47770a <=( (not A202)  and  A201 );
 a47773a <=( A232  and  (not A203) );
 a47774a <=( a47773a  and  a47770a );
 a47775a <=( a47774a  and  a47767a );
 a47778a <=( A234  and  (not A233) );
 a47781a <=( (not A265)  and  A235 );
 a47782a <=( a47781a  and  a47778a );
 a47785a <=( (not A267)  and  A266 );
 a47788a <=( (not A269)  and  (not A268) );
 a47789a <=( a47788a  and  a47785a );
 a47790a <=( a47789a  and  a47782a );
 a47793a <=( A168  and  (not A170) );
 a47796a <=( A166  and  (not A167) );
 a47797a <=( a47796a  and  a47793a );
 a47800a <=( (not A202)  and  A201 );
 a47803a <=( A232  and  (not A203) );
 a47804a <=( a47803a  and  a47800a );
 a47805a <=( a47804a  and  a47797a );
 a47808a <=( A234  and  (not A233) );
 a47811a <=( A265  and  A235 );
 a47812a <=( a47811a  and  a47808a );
 a47815a <=( (not A267)  and  (not A266) );
 a47818a <=( (not A269)  and  (not A268) );
 a47819a <=( a47818a  and  a47815a );
 a47820a <=( a47819a  and  a47812a );
 a47823a <=( A168  and  (not A170) );
 a47826a <=( A166  and  (not A167) );
 a47827a <=( a47826a  and  a47823a );
 a47830a <=( (not A202)  and  A201 );
 a47833a <=( A232  and  (not A203) );
 a47834a <=( a47833a  and  a47830a );
 a47835a <=( a47834a  and  a47827a );
 a47838a <=( A234  and  (not A233) );
 a47841a <=( A298  and  A236 );
 a47842a <=( a47841a  and  a47838a );
 a47845a <=( (not A300)  and  (not A299) );
 a47848a <=( (not A302)  and  (not A301) );
 a47849a <=( a47848a  and  a47845a );
 a47850a <=( a47849a  and  a47842a );
 a47853a <=( A168  and  (not A170) );
 a47856a <=( A166  and  (not A167) );
 a47857a <=( a47856a  and  a47853a );
 a47860a <=( (not A202)  and  A201 );
 a47863a <=( A232  and  (not A203) );
 a47864a <=( a47863a  and  a47860a );
 a47865a <=( a47864a  and  a47857a );
 a47868a <=( A234  and  (not A233) );
 a47871a <=( (not A298)  and  A236 );
 a47872a <=( a47871a  and  a47868a );
 a47875a <=( (not A300)  and  A299 );
 a47878a <=( (not A302)  and  (not A301) );
 a47879a <=( a47878a  and  a47875a );
 a47880a <=( a47879a  and  a47872a );
 a47883a <=( A168  and  (not A170) );
 a47886a <=( A166  and  (not A167) );
 a47887a <=( a47886a  and  a47883a );
 a47890a <=( (not A202)  and  A201 );
 a47893a <=( A232  and  (not A203) );
 a47894a <=( a47893a  and  a47890a );
 a47895a <=( a47894a  and  a47887a );
 a47898a <=( A234  and  (not A233) );
 a47901a <=( (not A265)  and  A236 );
 a47902a <=( a47901a  and  a47898a );
 a47905a <=( (not A267)  and  A266 );
 a47908a <=( (not A269)  and  (not A268) );
 a47909a <=( a47908a  and  a47905a );
 a47910a <=( a47909a  and  a47902a );
 a47913a <=( A168  and  (not A170) );
 a47916a <=( A166  and  (not A167) );
 a47917a <=( a47916a  and  a47913a );
 a47920a <=( (not A202)  and  A201 );
 a47923a <=( A232  and  (not A203) );
 a47924a <=( a47923a  and  a47920a );
 a47925a <=( a47924a  and  a47917a );
 a47928a <=( A234  and  (not A233) );
 a47931a <=( A265  and  A236 );
 a47932a <=( a47931a  and  a47928a );
 a47935a <=( (not A267)  and  (not A266) );
 a47938a <=( (not A269)  and  (not A268) );
 a47939a <=( a47938a  and  a47935a );
 a47940a <=( a47939a  and  a47932a );
 a47943a <=( A168  and  (not A170) );
 a47946a <=( A166  and  (not A167) );
 a47947a <=( a47946a  and  a47943a );
 a47950a <=( (not A202)  and  A201 );
 a47953a <=( A232  and  (not A203) );
 a47954a <=( a47953a  and  a47950a );
 a47955a <=( a47954a  and  a47947a );
 a47958a <=( (not A234)  and  (not A233) );
 a47961a <=( (not A236)  and  (not A235) );
 a47962a <=( a47961a  and  a47958a );
 a47965a <=( (not A299)  and  A298 );
 a47968a <=( A301  and  A300 );
 a47969a <=( a47968a  and  a47965a );
 a47970a <=( a47969a  and  a47962a );
 a47973a <=( A168  and  (not A170) );
 a47976a <=( A166  and  (not A167) );
 a47977a <=( a47976a  and  a47973a );
 a47980a <=( (not A202)  and  A201 );
 a47983a <=( A232  and  (not A203) );
 a47984a <=( a47983a  and  a47980a );
 a47985a <=( a47984a  and  a47977a );
 a47988a <=( (not A234)  and  (not A233) );
 a47991a <=( (not A236)  and  (not A235) );
 a47992a <=( a47991a  and  a47988a );
 a47995a <=( (not A299)  and  A298 );
 a47998a <=( A302  and  A300 );
 a47999a <=( a47998a  and  a47995a );
 a48000a <=( a47999a  and  a47992a );
 a48003a <=( A168  and  (not A170) );
 a48006a <=( A166  and  (not A167) );
 a48007a <=( a48006a  and  a48003a );
 a48010a <=( (not A202)  and  A201 );
 a48013a <=( A232  and  (not A203) );
 a48014a <=( a48013a  and  a48010a );
 a48015a <=( a48014a  and  a48007a );
 a48018a <=( (not A234)  and  (not A233) );
 a48021a <=( (not A236)  and  (not A235) );
 a48022a <=( a48021a  and  a48018a );
 a48025a <=( A299  and  (not A298) );
 a48028a <=( A301  and  A300 );
 a48029a <=( a48028a  and  a48025a );
 a48030a <=( a48029a  and  a48022a );
 a48033a <=( A168  and  (not A170) );
 a48036a <=( A166  and  (not A167) );
 a48037a <=( a48036a  and  a48033a );
 a48040a <=( (not A202)  and  A201 );
 a48043a <=( A232  and  (not A203) );
 a48044a <=( a48043a  and  a48040a );
 a48045a <=( a48044a  and  a48037a );
 a48048a <=( (not A234)  and  (not A233) );
 a48051a <=( (not A236)  and  (not A235) );
 a48052a <=( a48051a  and  a48048a );
 a48055a <=( A299  and  (not A298) );
 a48058a <=( A302  and  A300 );
 a48059a <=( a48058a  and  a48055a );
 a48060a <=( a48059a  and  a48052a );
 a48063a <=( A168  and  (not A170) );
 a48066a <=( A166  and  (not A167) );
 a48067a <=( a48066a  and  a48063a );
 a48070a <=( (not A202)  and  A201 );
 a48073a <=( A232  and  (not A203) );
 a48074a <=( a48073a  and  a48070a );
 a48075a <=( a48074a  and  a48067a );
 a48078a <=( (not A234)  and  (not A233) );
 a48081a <=( (not A236)  and  (not A235) );
 a48082a <=( a48081a  and  a48078a );
 a48085a <=( A266  and  (not A265) );
 a48088a <=( A268  and  A267 );
 a48089a <=( a48088a  and  a48085a );
 a48090a <=( a48089a  and  a48082a );
 a48093a <=( A168  and  (not A170) );
 a48096a <=( A166  and  (not A167) );
 a48097a <=( a48096a  and  a48093a );
 a48100a <=( (not A202)  and  A201 );
 a48103a <=( A232  and  (not A203) );
 a48104a <=( a48103a  and  a48100a );
 a48105a <=( a48104a  and  a48097a );
 a48108a <=( (not A234)  and  (not A233) );
 a48111a <=( (not A236)  and  (not A235) );
 a48112a <=( a48111a  and  a48108a );
 a48115a <=( A266  and  (not A265) );
 a48118a <=( A269  and  A267 );
 a48119a <=( a48118a  and  a48115a );
 a48120a <=( a48119a  and  a48112a );
 a48123a <=( A168  and  (not A170) );
 a48126a <=( A166  and  (not A167) );
 a48127a <=( a48126a  and  a48123a );
 a48130a <=( (not A202)  and  A201 );
 a48133a <=( A232  and  (not A203) );
 a48134a <=( a48133a  and  a48130a );
 a48135a <=( a48134a  and  a48127a );
 a48138a <=( (not A234)  and  (not A233) );
 a48141a <=( (not A236)  and  (not A235) );
 a48142a <=( a48141a  and  a48138a );
 a48145a <=( (not A266)  and  A265 );
 a48148a <=( A268  and  A267 );
 a48149a <=( a48148a  and  a48145a );
 a48150a <=( a48149a  and  a48142a );
 a48153a <=( A168  and  (not A170) );
 a48156a <=( A166  and  (not A167) );
 a48157a <=( a48156a  and  a48153a );
 a48160a <=( (not A202)  and  A201 );
 a48163a <=( A232  and  (not A203) );
 a48164a <=( a48163a  and  a48160a );
 a48165a <=( a48164a  and  a48157a );
 a48168a <=( (not A234)  and  (not A233) );
 a48171a <=( (not A236)  and  (not A235) );
 a48172a <=( a48171a  and  a48168a );
 a48175a <=( (not A266)  and  A265 );
 a48178a <=( A269  and  A267 );
 a48179a <=( a48178a  and  a48175a );
 a48180a <=( a48179a  and  a48172a );
 a48183a <=( A168  and  (not A170) );
 a48186a <=( A166  and  (not A167) );
 a48187a <=( a48186a  and  a48183a );
 a48190a <=( A202  and  (not A201) );
 a48193a <=( A233  and  (not A232) );
 a48194a <=( a48193a  and  a48190a );
 a48195a <=( a48194a  and  a48187a );
 a48198a <=( (not A235)  and  (not A234) );
 a48201a <=( A298  and  (not A236) );
 a48202a <=( a48201a  and  a48198a );
 a48205a <=( (not A300)  and  (not A299) );
 a48208a <=( (not A302)  and  (not A301) );
 a48209a <=( a48208a  and  a48205a );
 a48210a <=( a48209a  and  a48202a );
 a48213a <=( A168  and  (not A170) );
 a48216a <=( A166  and  (not A167) );
 a48217a <=( a48216a  and  a48213a );
 a48220a <=( A202  and  (not A201) );
 a48223a <=( A233  and  (not A232) );
 a48224a <=( a48223a  and  a48220a );
 a48225a <=( a48224a  and  a48217a );
 a48228a <=( (not A235)  and  (not A234) );
 a48231a <=( (not A298)  and  (not A236) );
 a48232a <=( a48231a  and  a48228a );
 a48235a <=( (not A300)  and  A299 );
 a48238a <=( (not A302)  and  (not A301) );
 a48239a <=( a48238a  and  a48235a );
 a48240a <=( a48239a  and  a48232a );
 a48243a <=( A168  and  (not A170) );
 a48246a <=( A166  and  (not A167) );
 a48247a <=( a48246a  and  a48243a );
 a48250a <=( A202  and  (not A201) );
 a48253a <=( A233  and  (not A232) );
 a48254a <=( a48253a  and  a48250a );
 a48255a <=( a48254a  and  a48247a );
 a48258a <=( (not A235)  and  (not A234) );
 a48261a <=( (not A265)  and  (not A236) );
 a48262a <=( a48261a  and  a48258a );
 a48265a <=( (not A267)  and  A266 );
 a48268a <=( (not A269)  and  (not A268) );
 a48269a <=( a48268a  and  a48265a );
 a48270a <=( a48269a  and  a48262a );
 a48273a <=( A168  and  (not A170) );
 a48276a <=( A166  and  (not A167) );
 a48277a <=( a48276a  and  a48273a );
 a48280a <=( A202  and  (not A201) );
 a48283a <=( A233  and  (not A232) );
 a48284a <=( a48283a  and  a48280a );
 a48285a <=( a48284a  and  a48277a );
 a48288a <=( (not A235)  and  (not A234) );
 a48291a <=( A265  and  (not A236) );
 a48292a <=( a48291a  and  a48288a );
 a48295a <=( (not A267)  and  (not A266) );
 a48298a <=( (not A269)  and  (not A268) );
 a48299a <=( a48298a  and  a48295a );
 a48300a <=( a48299a  and  a48292a );
 a48303a <=( A168  and  (not A170) );
 a48306a <=( A166  and  (not A167) );
 a48307a <=( a48306a  and  a48303a );
 a48310a <=( A202  and  (not A201) );
 a48313a <=( (not A233)  and  A232 );
 a48314a <=( a48313a  and  a48310a );
 a48315a <=( a48314a  and  a48307a );
 a48318a <=( (not A235)  and  (not A234) );
 a48321a <=( A298  and  (not A236) );
 a48322a <=( a48321a  and  a48318a );
 a48325a <=( (not A300)  and  (not A299) );
 a48328a <=( (not A302)  and  (not A301) );
 a48329a <=( a48328a  and  a48325a );
 a48330a <=( a48329a  and  a48322a );
 a48333a <=( A168  and  (not A170) );
 a48336a <=( A166  and  (not A167) );
 a48337a <=( a48336a  and  a48333a );
 a48340a <=( A202  and  (not A201) );
 a48343a <=( (not A233)  and  A232 );
 a48344a <=( a48343a  and  a48340a );
 a48345a <=( a48344a  and  a48337a );
 a48348a <=( (not A235)  and  (not A234) );
 a48351a <=( (not A298)  and  (not A236) );
 a48352a <=( a48351a  and  a48348a );
 a48355a <=( (not A300)  and  A299 );
 a48358a <=( (not A302)  and  (not A301) );
 a48359a <=( a48358a  and  a48355a );
 a48360a <=( a48359a  and  a48352a );
 a48363a <=( A168  and  (not A170) );
 a48366a <=( A166  and  (not A167) );
 a48367a <=( a48366a  and  a48363a );
 a48370a <=( A202  and  (not A201) );
 a48373a <=( (not A233)  and  A232 );
 a48374a <=( a48373a  and  a48370a );
 a48375a <=( a48374a  and  a48367a );
 a48378a <=( (not A235)  and  (not A234) );
 a48381a <=( (not A265)  and  (not A236) );
 a48382a <=( a48381a  and  a48378a );
 a48385a <=( (not A267)  and  A266 );
 a48388a <=( (not A269)  and  (not A268) );
 a48389a <=( a48388a  and  a48385a );
 a48390a <=( a48389a  and  a48382a );
 a48393a <=( A168  and  (not A170) );
 a48396a <=( A166  and  (not A167) );
 a48397a <=( a48396a  and  a48393a );
 a48400a <=( A202  and  (not A201) );
 a48403a <=( (not A233)  and  A232 );
 a48404a <=( a48403a  and  a48400a );
 a48405a <=( a48404a  and  a48397a );
 a48408a <=( (not A235)  and  (not A234) );
 a48411a <=( A265  and  (not A236) );
 a48412a <=( a48411a  and  a48408a );
 a48415a <=( (not A267)  and  (not A266) );
 a48418a <=( (not A269)  and  (not A268) );
 a48419a <=( a48418a  and  a48415a );
 a48420a <=( a48419a  and  a48412a );
 a48423a <=( A168  and  (not A170) );
 a48426a <=( A166  and  (not A167) );
 a48427a <=( a48426a  and  a48423a );
 a48430a <=( A203  and  (not A201) );
 a48433a <=( A233  and  (not A232) );
 a48434a <=( a48433a  and  a48430a );
 a48435a <=( a48434a  and  a48427a );
 a48438a <=( (not A235)  and  (not A234) );
 a48441a <=( A298  and  (not A236) );
 a48442a <=( a48441a  and  a48438a );
 a48445a <=( (not A300)  and  (not A299) );
 a48448a <=( (not A302)  and  (not A301) );
 a48449a <=( a48448a  and  a48445a );
 a48450a <=( a48449a  and  a48442a );
 a48453a <=( A168  and  (not A170) );
 a48456a <=( A166  and  (not A167) );
 a48457a <=( a48456a  and  a48453a );
 a48460a <=( A203  and  (not A201) );
 a48463a <=( A233  and  (not A232) );
 a48464a <=( a48463a  and  a48460a );
 a48465a <=( a48464a  and  a48457a );
 a48468a <=( (not A235)  and  (not A234) );
 a48471a <=( (not A298)  and  (not A236) );
 a48472a <=( a48471a  and  a48468a );
 a48475a <=( (not A300)  and  A299 );
 a48478a <=( (not A302)  and  (not A301) );
 a48479a <=( a48478a  and  a48475a );
 a48480a <=( a48479a  and  a48472a );
 a48483a <=( A168  and  (not A170) );
 a48486a <=( A166  and  (not A167) );
 a48487a <=( a48486a  and  a48483a );
 a48490a <=( A203  and  (not A201) );
 a48493a <=( A233  and  (not A232) );
 a48494a <=( a48493a  and  a48490a );
 a48495a <=( a48494a  and  a48487a );
 a48498a <=( (not A235)  and  (not A234) );
 a48501a <=( (not A265)  and  (not A236) );
 a48502a <=( a48501a  and  a48498a );
 a48505a <=( (not A267)  and  A266 );
 a48508a <=( (not A269)  and  (not A268) );
 a48509a <=( a48508a  and  a48505a );
 a48510a <=( a48509a  and  a48502a );
 a48513a <=( A168  and  (not A170) );
 a48516a <=( A166  and  (not A167) );
 a48517a <=( a48516a  and  a48513a );
 a48520a <=( A203  and  (not A201) );
 a48523a <=( A233  and  (not A232) );
 a48524a <=( a48523a  and  a48520a );
 a48525a <=( a48524a  and  a48517a );
 a48528a <=( (not A235)  and  (not A234) );
 a48531a <=( A265  and  (not A236) );
 a48532a <=( a48531a  and  a48528a );
 a48535a <=( (not A267)  and  (not A266) );
 a48538a <=( (not A269)  and  (not A268) );
 a48539a <=( a48538a  and  a48535a );
 a48540a <=( a48539a  and  a48532a );
 a48543a <=( A168  and  (not A170) );
 a48546a <=( A166  and  (not A167) );
 a48547a <=( a48546a  and  a48543a );
 a48550a <=( A203  and  (not A201) );
 a48553a <=( (not A233)  and  A232 );
 a48554a <=( a48553a  and  a48550a );
 a48555a <=( a48554a  and  a48547a );
 a48558a <=( (not A235)  and  (not A234) );
 a48561a <=( A298  and  (not A236) );
 a48562a <=( a48561a  and  a48558a );
 a48565a <=( (not A300)  and  (not A299) );
 a48568a <=( (not A302)  and  (not A301) );
 a48569a <=( a48568a  and  a48565a );
 a48570a <=( a48569a  and  a48562a );
 a48573a <=( A168  and  (not A170) );
 a48576a <=( A166  and  (not A167) );
 a48577a <=( a48576a  and  a48573a );
 a48580a <=( A203  and  (not A201) );
 a48583a <=( (not A233)  and  A232 );
 a48584a <=( a48583a  and  a48580a );
 a48585a <=( a48584a  and  a48577a );
 a48588a <=( (not A235)  and  (not A234) );
 a48591a <=( (not A298)  and  (not A236) );
 a48592a <=( a48591a  and  a48588a );
 a48595a <=( (not A300)  and  A299 );
 a48598a <=( (not A302)  and  (not A301) );
 a48599a <=( a48598a  and  a48595a );
 a48600a <=( a48599a  and  a48592a );
 a48603a <=( A168  and  (not A170) );
 a48606a <=( A166  and  (not A167) );
 a48607a <=( a48606a  and  a48603a );
 a48610a <=( A203  and  (not A201) );
 a48613a <=( (not A233)  and  A232 );
 a48614a <=( a48613a  and  a48610a );
 a48615a <=( a48614a  and  a48607a );
 a48618a <=( (not A235)  and  (not A234) );
 a48621a <=( (not A265)  and  (not A236) );
 a48622a <=( a48621a  and  a48618a );
 a48625a <=( (not A267)  and  A266 );
 a48628a <=( (not A269)  and  (not A268) );
 a48629a <=( a48628a  and  a48625a );
 a48630a <=( a48629a  and  a48622a );
 a48633a <=( A168  and  (not A170) );
 a48636a <=( A166  and  (not A167) );
 a48637a <=( a48636a  and  a48633a );
 a48640a <=( A203  and  (not A201) );
 a48643a <=( (not A233)  and  A232 );
 a48644a <=( a48643a  and  a48640a );
 a48645a <=( a48644a  and  a48637a );
 a48648a <=( (not A235)  and  (not A234) );
 a48651a <=( A265  and  (not A236) );
 a48652a <=( a48651a  and  a48648a );
 a48655a <=( (not A267)  and  (not A266) );
 a48658a <=( (not A269)  and  (not A268) );
 a48659a <=( a48658a  and  a48655a );
 a48660a <=( a48659a  and  a48652a );
 a48663a <=( A168  and  (not A170) );
 a48666a <=( A166  and  (not A167) );
 a48667a <=( a48666a  and  a48663a );
 a48670a <=( A200  and  A199 );
 a48673a <=( A233  and  (not A232) );
 a48674a <=( a48673a  and  a48670a );
 a48675a <=( a48674a  and  a48667a );
 a48678a <=( (not A235)  and  (not A234) );
 a48681a <=( A298  and  (not A236) );
 a48682a <=( a48681a  and  a48678a );
 a48685a <=( (not A300)  and  (not A299) );
 a48688a <=( (not A302)  and  (not A301) );
 a48689a <=( a48688a  and  a48685a );
 a48690a <=( a48689a  and  a48682a );
 a48693a <=( A168  and  (not A170) );
 a48696a <=( A166  and  (not A167) );
 a48697a <=( a48696a  and  a48693a );
 a48700a <=( A200  and  A199 );
 a48703a <=( A233  and  (not A232) );
 a48704a <=( a48703a  and  a48700a );
 a48705a <=( a48704a  and  a48697a );
 a48708a <=( (not A235)  and  (not A234) );
 a48711a <=( (not A298)  and  (not A236) );
 a48712a <=( a48711a  and  a48708a );
 a48715a <=( (not A300)  and  A299 );
 a48718a <=( (not A302)  and  (not A301) );
 a48719a <=( a48718a  and  a48715a );
 a48720a <=( a48719a  and  a48712a );
 a48723a <=( A168  and  (not A170) );
 a48726a <=( A166  and  (not A167) );
 a48727a <=( a48726a  and  a48723a );
 a48730a <=( A200  and  A199 );
 a48733a <=( A233  and  (not A232) );
 a48734a <=( a48733a  and  a48730a );
 a48735a <=( a48734a  and  a48727a );
 a48738a <=( (not A235)  and  (not A234) );
 a48741a <=( (not A265)  and  (not A236) );
 a48742a <=( a48741a  and  a48738a );
 a48745a <=( (not A267)  and  A266 );
 a48748a <=( (not A269)  and  (not A268) );
 a48749a <=( a48748a  and  a48745a );
 a48750a <=( a48749a  and  a48742a );
 a48753a <=( A168  and  (not A170) );
 a48756a <=( A166  and  (not A167) );
 a48757a <=( a48756a  and  a48753a );
 a48760a <=( A200  and  A199 );
 a48763a <=( A233  and  (not A232) );
 a48764a <=( a48763a  and  a48760a );
 a48765a <=( a48764a  and  a48757a );
 a48768a <=( (not A235)  and  (not A234) );
 a48771a <=( A265  and  (not A236) );
 a48772a <=( a48771a  and  a48768a );
 a48775a <=( (not A267)  and  (not A266) );
 a48778a <=( (not A269)  and  (not A268) );
 a48779a <=( a48778a  and  a48775a );
 a48780a <=( a48779a  and  a48772a );
 a48783a <=( A168  and  (not A170) );
 a48786a <=( A166  and  (not A167) );
 a48787a <=( a48786a  and  a48783a );
 a48790a <=( A200  and  A199 );
 a48793a <=( (not A233)  and  A232 );
 a48794a <=( a48793a  and  a48790a );
 a48795a <=( a48794a  and  a48787a );
 a48798a <=( (not A235)  and  (not A234) );
 a48801a <=( A298  and  (not A236) );
 a48802a <=( a48801a  and  a48798a );
 a48805a <=( (not A300)  and  (not A299) );
 a48808a <=( (not A302)  and  (not A301) );
 a48809a <=( a48808a  and  a48805a );
 a48810a <=( a48809a  and  a48802a );
 a48813a <=( A168  and  (not A170) );
 a48816a <=( A166  and  (not A167) );
 a48817a <=( a48816a  and  a48813a );
 a48820a <=( A200  and  A199 );
 a48823a <=( (not A233)  and  A232 );
 a48824a <=( a48823a  and  a48820a );
 a48825a <=( a48824a  and  a48817a );
 a48828a <=( (not A235)  and  (not A234) );
 a48831a <=( (not A298)  and  (not A236) );
 a48832a <=( a48831a  and  a48828a );
 a48835a <=( (not A300)  and  A299 );
 a48838a <=( (not A302)  and  (not A301) );
 a48839a <=( a48838a  and  a48835a );
 a48840a <=( a48839a  and  a48832a );
 a48843a <=( A168  and  (not A170) );
 a48846a <=( A166  and  (not A167) );
 a48847a <=( a48846a  and  a48843a );
 a48850a <=( A200  and  A199 );
 a48853a <=( (not A233)  and  A232 );
 a48854a <=( a48853a  and  a48850a );
 a48855a <=( a48854a  and  a48847a );
 a48858a <=( (not A235)  and  (not A234) );
 a48861a <=( (not A265)  and  (not A236) );
 a48862a <=( a48861a  and  a48858a );
 a48865a <=( (not A267)  and  A266 );
 a48868a <=( (not A269)  and  (not A268) );
 a48869a <=( a48868a  and  a48865a );
 a48870a <=( a48869a  and  a48862a );
 a48873a <=( A168  and  (not A170) );
 a48876a <=( A166  and  (not A167) );
 a48877a <=( a48876a  and  a48873a );
 a48880a <=( A200  and  A199 );
 a48883a <=( (not A233)  and  A232 );
 a48884a <=( a48883a  and  a48880a );
 a48885a <=( a48884a  and  a48877a );
 a48888a <=( (not A235)  and  (not A234) );
 a48891a <=( A265  and  (not A236) );
 a48892a <=( a48891a  and  a48888a );
 a48895a <=( (not A267)  and  (not A266) );
 a48898a <=( (not A269)  and  (not A268) );
 a48899a <=( a48898a  and  a48895a );
 a48900a <=( a48899a  and  a48892a );
 a48903a <=( A168  and  (not A170) );
 a48906a <=( A166  and  (not A167) );
 a48907a <=( a48906a  and  a48903a );
 a48910a <=( (not A200)  and  (not A199) );
 a48913a <=( A233  and  (not A232) );
 a48914a <=( a48913a  and  a48910a );
 a48915a <=( a48914a  and  a48907a );
 a48918a <=( (not A235)  and  (not A234) );
 a48921a <=( A298  and  (not A236) );
 a48922a <=( a48921a  and  a48918a );
 a48925a <=( (not A300)  and  (not A299) );
 a48928a <=( (not A302)  and  (not A301) );
 a48929a <=( a48928a  and  a48925a );
 a48930a <=( a48929a  and  a48922a );
 a48933a <=( A168  and  (not A170) );
 a48936a <=( A166  and  (not A167) );
 a48937a <=( a48936a  and  a48933a );
 a48940a <=( (not A200)  and  (not A199) );
 a48943a <=( A233  and  (not A232) );
 a48944a <=( a48943a  and  a48940a );
 a48945a <=( a48944a  and  a48937a );
 a48948a <=( (not A235)  and  (not A234) );
 a48951a <=( (not A298)  and  (not A236) );
 a48952a <=( a48951a  and  a48948a );
 a48955a <=( (not A300)  and  A299 );
 a48958a <=( (not A302)  and  (not A301) );
 a48959a <=( a48958a  and  a48955a );
 a48960a <=( a48959a  and  a48952a );
 a48963a <=( A168  and  (not A170) );
 a48966a <=( A166  and  (not A167) );
 a48967a <=( a48966a  and  a48963a );
 a48970a <=( (not A200)  and  (not A199) );
 a48973a <=( A233  and  (not A232) );
 a48974a <=( a48973a  and  a48970a );
 a48975a <=( a48974a  and  a48967a );
 a48978a <=( (not A235)  and  (not A234) );
 a48981a <=( (not A265)  and  (not A236) );
 a48982a <=( a48981a  and  a48978a );
 a48985a <=( (not A267)  and  A266 );
 a48988a <=( (not A269)  and  (not A268) );
 a48989a <=( a48988a  and  a48985a );
 a48990a <=( a48989a  and  a48982a );
 a48993a <=( A168  and  (not A170) );
 a48996a <=( A166  and  (not A167) );
 a48997a <=( a48996a  and  a48993a );
 a49000a <=( (not A200)  and  (not A199) );
 a49003a <=( A233  and  (not A232) );
 a49004a <=( a49003a  and  a49000a );
 a49005a <=( a49004a  and  a48997a );
 a49008a <=( (not A235)  and  (not A234) );
 a49011a <=( A265  and  (not A236) );
 a49012a <=( a49011a  and  a49008a );
 a49015a <=( (not A267)  and  (not A266) );
 a49018a <=( (not A269)  and  (not A268) );
 a49019a <=( a49018a  and  a49015a );
 a49020a <=( a49019a  and  a49012a );
 a49023a <=( A168  and  (not A170) );
 a49026a <=( A166  and  (not A167) );
 a49027a <=( a49026a  and  a49023a );
 a49030a <=( (not A200)  and  (not A199) );
 a49033a <=( (not A233)  and  A232 );
 a49034a <=( a49033a  and  a49030a );
 a49035a <=( a49034a  and  a49027a );
 a49038a <=( (not A235)  and  (not A234) );
 a49041a <=( A298  and  (not A236) );
 a49042a <=( a49041a  and  a49038a );
 a49045a <=( (not A300)  and  (not A299) );
 a49048a <=( (not A302)  and  (not A301) );
 a49049a <=( a49048a  and  a49045a );
 a49050a <=( a49049a  and  a49042a );
 a49053a <=( A168  and  (not A170) );
 a49056a <=( A166  and  (not A167) );
 a49057a <=( a49056a  and  a49053a );
 a49060a <=( (not A200)  and  (not A199) );
 a49063a <=( (not A233)  and  A232 );
 a49064a <=( a49063a  and  a49060a );
 a49065a <=( a49064a  and  a49057a );
 a49068a <=( (not A235)  and  (not A234) );
 a49071a <=( (not A298)  and  (not A236) );
 a49072a <=( a49071a  and  a49068a );
 a49075a <=( (not A300)  and  A299 );
 a49078a <=( (not A302)  and  (not A301) );
 a49079a <=( a49078a  and  a49075a );
 a49080a <=( a49079a  and  a49072a );
 a49083a <=( A168  and  (not A170) );
 a49086a <=( A166  and  (not A167) );
 a49087a <=( a49086a  and  a49083a );
 a49090a <=( (not A200)  and  (not A199) );
 a49093a <=( (not A233)  and  A232 );
 a49094a <=( a49093a  and  a49090a );
 a49095a <=( a49094a  and  a49087a );
 a49098a <=( (not A235)  and  (not A234) );
 a49101a <=( (not A265)  and  (not A236) );
 a49102a <=( a49101a  and  a49098a );
 a49105a <=( (not A267)  and  A266 );
 a49108a <=( (not A269)  and  (not A268) );
 a49109a <=( a49108a  and  a49105a );
 a49110a <=( a49109a  and  a49102a );
 a49113a <=( A168  and  (not A170) );
 a49116a <=( A166  and  (not A167) );
 a49117a <=( a49116a  and  a49113a );
 a49120a <=( (not A200)  and  (not A199) );
 a49123a <=( (not A233)  and  A232 );
 a49124a <=( a49123a  and  a49120a );
 a49125a <=( a49124a  and  a49117a );
 a49128a <=( (not A235)  and  (not A234) );
 a49131a <=( A265  and  (not A236) );
 a49132a <=( a49131a  and  a49128a );
 a49135a <=( (not A267)  and  (not A266) );
 a49138a <=( (not A269)  and  (not A268) );
 a49139a <=( a49138a  and  a49135a );
 a49140a <=( a49139a  and  a49132a );
 a49143a <=( A168  and  A169 );
 a49146a <=( (not A166)  and  A167 );
 a49147a <=( a49146a  and  a49143a );
 a49150a <=( (not A202)  and  A201 );
 a49153a <=( (not A232)  and  (not A203) );
 a49154a <=( a49153a  and  a49150a );
 a49155a <=( a49154a  and  a49147a );
 a49158a <=( A234  and  A233 );
 a49161a <=( A298  and  A235 );
 a49162a <=( a49161a  and  a49158a );
 a49165a <=( (not A300)  and  (not A299) );
 a49168a <=( (not A302)  and  (not A301) );
 a49169a <=( a49168a  and  a49165a );
 a49170a <=( a49169a  and  a49162a );
 a49173a <=( A168  and  A169 );
 a49176a <=( (not A166)  and  A167 );
 a49177a <=( a49176a  and  a49173a );
 a49180a <=( (not A202)  and  A201 );
 a49183a <=( (not A232)  and  (not A203) );
 a49184a <=( a49183a  and  a49180a );
 a49185a <=( a49184a  and  a49177a );
 a49188a <=( A234  and  A233 );
 a49191a <=( (not A298)  and  A235 );
 a49192a <=( a49191a  and  a49188a );
 a49195a <=( (not A300)  and  A299 );
 a49198a <=( (not A302)  and  (not A301) );
 a49199a <=( a49198a  and  a49195a );
 a49200a <=( a49199a  and  a49192a );
 a49203a <=( A168  and  A169 );
 a49206a <=( (not A166)  and  A167 );
 a49207a <=( a49206a  and  a49203a );
 a49210a <=( (not A202)  and  A201 );
 a49213a <=( (not A232)  and  (not A203) );
 a49214a <=( a49213a  and  a49210a );
 a49215a <=( a49214a  and  a49207a );
 a49218a <=( A234  and  A233 );
 a49221a <=( (not A265)  and  A235 );
 a49222a <=( a49221a  and  a49218a );
 a49225a <=( (not A267)  and  A266 );
 a49228a <=( (not A269)  and  (not A268) );
 a49229a <=( a49228a  and  a49225a );
 a49230a <=( a49229a  and  a49222a );
 a49233a <=( A168  and  A169 );
 a49236a <=( (not A166)  and  A167 );
 a49237a <=( a49236a  and  a49233a );
 a49240a <=( (not A202)  and  A201 );
 a49243a <=( (not A232)  and  (not A203) );
 a49244a <=( a49243a  and  a49240a );
 a49245a <=( a49244a  and  a49237a );
 a49248a <=( A234  and  A233 );
 a49251a <=( A265  and  A235 );
 a49252a <=( a49251a  and  a49248a );
 a49255a <=( (not A267)  and  (not A266) );
 a49258a <=( (not A269)  and  (not A268) );
 a49259a <=( a49258a  and  a49255a );
 a49260a <=( a49259a  and  a49252a );
 a49263a <=( A168  and  A169 );
 a49266a <=( (not A166)  and  A167 );
 a49267a <=( a49266a  and  a49263a );
 a49270a <=( (not A202)  and  A201 );
 a49273a <=( (not A232)  and  (not A203) );
 a49274a <=( a49273a  and  a49270a );
 a49275a <=( a49274a  and  a49267a );
 a49278a <=( A234  and  A233 );
 a49281a <=( A298  and  A236 );
 a49282a <=( a49281a  and  a49278a );
 a49285a <=( (not A300)  and  (not A299) );
 a49288a <=( (not A302)  and  (not A301) );
 a49289a <=( a49288a  and  a49285a );
 a49290a <=( a49289a  and  a49282a );
 a49293a <=( A168  and  A169 );
 a49296a <=( (not A166)  and  A167 );
 a49297a <=( a49296a  and  a49293a );
 a49300a <=( (not A202)  and  A201 );
 a49303a <=( (not A232)  and  (not A203) );
 a49304a <=( a49303a  and  a49300a );
 a49305a <=( a49304a  and  a49297a );
 a49308a <=( A234  and  A233 );
 a49311a <=( (not A298)  and  A236 );
 a49312a <=( a49311a  and  a49308a );
 a49315a <=( (not A300)  and  A299 );
 a49318a <=( (not A302)  and  (not A301) );
 a49319a <=( a49318a  and  a49315a );
 a49320a <=( a49319a  and  a49312a );
 a49323a <=( A168  and  A169 );
 a49326a <=( (not A166)  and  A167 );
 a49327a <=( a49326a  and  a49323a );
 a49330a <=( (not A202)  and  A201 );
 a49333a <=( (not A232)  and  (not A203) );
 a49334a <=( a49333a  and  a49330a );
 a49335a <=( a49334a  and  a49327a );
 a49338a <=( A234  and  A233 );
 a49341a <=( (not A265)  and  A236 );
 a49342a <=( a49341a  and  a49338a );
 a49345a <=( (not A267)  and  A266 );
 a49348a <=( (not A269)  and  (not A268) );
 a49349a <=( a49348a  and  a49345a );
 a49350a <=( a49349a  and  a49342a );
 a49353a <=( A168  and  A169 );
 a49356a <=( (not A166)  and  A167 );
 a49357a <=( a49356a  and  a49353a );
 a49360a <=( (not A202)  and  A201 );
 a49363a <=( (not A232)  and  (not A203) );
 a49364a <=( a49363a  and  a49360a );
 a49365a <=( a49364a  and  a49357a );
 a49368a <=( A234  and  A233 );
 a49371a <=( A265  and  A236 );
 a49372a <=( a49371a  and  a49368a );
 a49375a <=( (not A267)  and  (not A266) );
 a49378a <=( (not A269)  and  (not A268) );
 a49379a <=( a49378a  and  a49375a );
 a49380a <=( a49379a  and  a49372a );
 a49383a <=( A168  and  A169 );
 a49386a <=( (not A166)  and  A167 );
 a49387a <=( a49386a  and  a49383a );
 a49390a <=( (not A202)  and  A201 );
 a49393a <=( (not A232)  and  (not A203) );
 a49394a <=( a49393a  and  a49390a );
 a49395a <=( a49394a  and  a49387a );
 a49398a <=( (not A234)  and  A233 );
 a49401a <=( (not A236)  and  (not A235) );
 a49402a <=( a49401a  and  a49398a );
 a49405a <=( (not A299)  and  A298 );
 a49408a <=( A301  and  A300 );
 a49409a <=( a49408a  and  a49405a );
 a49410a <=( a49409a  and  a49402a );
 a49413a <=( A168  and  A169 );
 a49416a <=( (not A166)  and  A167 );
 a49417a <=( a49416a  and  a49413a );
 a49420a <=( (not A202)  and  A201 );
 a49423a <=( (not A232)  and  (not A203) );
 a49424a <=( a49423a  and  a49420a );
 a49425a <=( a49424a  and  a49417a );
 a49428a <=( (not A234)  and  A233 );
 a49431a <=( (not A236)  and  (not A235) );
 a49432a <=( a49431a  and  a49428a );
 a49435a <=( (not A299)  and  A298 );
 a49438a <=( A302  and  A300 );
 a49439a <=( a49438a  and  a49435a );
 a49440a <=( a49439a  and  a49432a );
 a49443a <=( A168  and  A169 );
 a49446a <=( (not A166)  and  A167 );
 a49447a <=( a49446a  and  a49443a );
 a49450a <=( (not A202)  and  A201 );
 a49453a <=( (not A232)  and  (not A203) );
 a49454a <=( a49453a  and  a49450a );
 a49455a <=( a49454a  and  a49447a );
 a49458a <=( (not A234)  and  A233 );
 a49461a <=( (not A236)  and  (not A235) );
 a49462a <=( a49461a  and  a49458a );
 a49465a <=( A299  and  (not A298) );
 a49468a <=( A301  and  A300 );
 a49469a <=( a49468a  and  a49465a );
 a49470a <=( a49469a  and  a49462a );
 a49473a <=( A168  and  A169 );
 a49476a <=( (not A166)  and  A167 );
 a49477a <=( a49476a  and  a49473a );
 a49480a <=( (not A202)  and  A201 );
 a49483a <=( (not A232)  and  (not A203) );
 a49484a <=( a49483a  and  a49480a );
 a49485a <=( a49484a  and  a49477a );
 a49488a <=( (not A234)  and  A233 );
 a49491a <=( (not A236)  and  (not A235) );
 a49492a <=( a49491a  and  a49488a );
 a49495a <=( A299  and  (not A298) );
 a49498a <=( A302  and  A300 );
 a49499a <=( a49498a  and  a49495a );
 a49500a <=( a49499a  and  a49492a );
 a49503a <=( A168  and  A169 );
 a49506a <=( (not A166)  and  A167 );
 a49507a <=( a49506a  and  a49503a );
 a49510a <=( (not A202)  and  A201 );
 a49513a <=( (not A232)  and  (not A203) );
 a49514a <=( a49513a  and  a49510a );
 a49515a <=( a49514a  and  a49507a );
 a49518a <=( (not A234)  and  A233 );
 a49521a <=( (not A236)  and  (not A235) );
 a49522a <=( a49521a  and  a49518a );
 a49525a <=( A266  and  (not A265) );
 a49528a <=( A268  and  A267 );
 a49529a <=( a49528a  and  a49525a );
 a49530a <=( a49529a  and  a49522a );
 a49533a <=( A168  and  A169 );
 a49536a <=( (not A166)  and  A167 );
 a49537a <=( a49536a  and  a49533a );
 a49540a <=( (not A202)  and  A201 );
 a49543a <=( (not A232)  and  (not A203) );
 a49544a <=( a49543a  and  a49540a );
 a49545a <=( a49544a  and  a49537a );
 a49548a <=( (not A234)  and  A233 );
 a49551a <=( (not A236)  and  (not A235) );
 a49552a <=( a49551a  and  a49548a );
 a49555a <=( A266  and  (not A265) );
 a49558a <=( A269  and  A267 );
 a49559a <=( a49558a  and  a49555a );
 a49560a <=( a49559a  and  a49552a );
 a49563a <=( A168  and  A169 );
 a49566a <=( (not A166)  and  A167 );
 a49567a <=( a49566a  and  a49563a );
 a49570a <=( (not A202)  and  A201 );
 a49573a <=( (not A232)  and  (not A203) );
 a49574a <=( a49573a  and  a49570a );
 a49575a <=( a49574a  and  a49567a );
 a49578a <=( (not A234)  and  A233 );
 a49581a <=( (not A236)  and  (not A235) );
 a49582a <=( a49581a  and  a49578a );
 a49585a <=( (not A266)  and  A265 );
 a49588a <=( A268  and  A267 );
 a49589a <=( a49588a  and  a49585a );
 a49590a <=( a49589a  and  a49582a );
 a49593a <=( A168  and  A169 );
 a49596a <=( (not A166)  and  A167 );
 a49597a <=( a49596a  and  a49593a );
 a49600a <=( (not A202)  and  A201 );
 a49603a <=( (not A232)  and  (not A203) );
 a49604a <=( a49603a  and  a49600a );
 a49605a <=( a49604a  and  a49597a );
 a49608a <=( (not A234)  and  A233 );
 a49611a <=( (not A236)  and  (not A235) );
 a49612a <=( a49611a  and  a49608a );
 a49615a <=( (not A266)  and  A265 );
 a49618a <=( A269  and  A267 );
 a49619a <=( a49618a  and  a49615a );
 a49620a <=( a49619a  and  a49612a );
 a49623a <=( A168  and  A169 );
 a49626a <=( (not A166)  and  A167 );
 a49627a <=( a49626a  and  a49623a );
 a49630a <=( (not A202)  and  A201 );
 a49633a <=( A232  and  (not A203) );
 a49634a <=( a49633a  and  a49630a );
 a49635a <=( a49634a  and  a49627a );
 a49638a <=( A234  and  (not A233) );
 a49641a <=( A298  and  A235 );
 a49642a <=( a49641a  and  a49638a );
 a49645a <=( (not A300)  and  (not A299) );
 a49648a <=( (not A302)  and  (not A301) );
 a49649a <=( a49648a  and  a49645a );
 a49650a <=( a49649a  and  a49642a );
 a49653a <=( A168  and  A169 );
 a49656a <=( (not A166)  and  A167 );
 a49657a <=( a49656a  and  a49653a );
 a49660a <=( (not A202)  and  A201 );
 a49663a <=( A232  and  (not A203) );
 a49664a <=( a49663a  and  a49660a );
 a49665a <=( a49664a  and  a49657a );
 a49668a <=( A234  and  (not A233) );
 a49671a <=( (not A298)  and  A235 );
 a49672a <=( a49671a  and  a49668a );
 a49675a <=( (not A300)  and  A299 );
 a49678a <=( (not A302)  and  (not A301) );
 a49679a <=( a49678a  and  a49675a );
 a49680a <=( a49679a  and  a49672a );
 a49683a <=( A168  and  A169 );
 a49686a <=( (not A166)  and  A167 );
 a49687a <=( a49686a  and  a49683a );
 a49690a <=( (not A202)  and  A201 );
 a49693a <=( A232  and  (not A203) );
 a49694a <=( a49693a  and  a49690a );
 a49695a <=( a49694a  and  a49687a );
 a49698a <=( A234  and  (not A233) );
 a49701a <=( (not A265)  and  A235 );
 a49702a <=( a49701a  and  a49698a );
 a49705a <=( (not A267)  and  A266 );
 a49708a <=( (not A269)  and  (not A268) );
 a49709a <=( a49708a  and  a49705a );
 a49710a <=( a49709a  and  a49702a );
 a49713a <=( A168  and  A169 );
 a49716a <=( (not A166)  and  A167 );
 a49717a <=( a49716a  and  a49713a );
 a49720a <=( (not A202)  and  A201 );
 a49723a <=( A232  and  (not A203) );
 a49724a <=( a49723a  and  a49720a );
 a49725a <=( a49724a  and  a49717a );
 a49728a <=( A234  and  (not A233) );
 a49731a <=( A265  and  A235 );
 a49732a <=( a49731a  and  a49728a );
 a49735a <=( (not A267)  and  (not A266) );
 a49738a <=( (not A269)  and  (not A268) );
 a49739a <=( a49738a  and  a49735a );
 a49740a <=( a49739a  and  a49732a );
 a49743a <=( A168  and  A169 );
 a49746a <=( (not A166)  and  A167 );
 a49747a <=( a49746a  and  a49743a );
 a49750a <=( (not A202)  and  A201 );
 a49753a <=( A232  and  (not A203) );
 a49754a <=( a49753a  and  a49750a );
 a49755a <=( a49754a  and  a49747a );
 a49758a <=( A234  and  (not A233) );
 a49761a <=( A298  and  A236 );
 a49762a <=( a49761a  and  a49758a );
 a49765a <=( (not A300)  and  (not A299) );
 a49768a <=( (not A302)  and  (not A301) );
 a49769a <=( a49768a  and  a49765a );
 a49770a <=( a49769a  and  a49762a );
 a49773a <=( A168  and  A169 );
 a49776a <=( (not A166)  and  A167 );
 a49777a <=( a49776a  and  a49773a );
 a49780a <=( (not A202)  and  A201 );
 a49783a <=( A232  and  (not A203) );
 a49784a <=( a49783a  and  a49780a );
 a49785a <=( a49784a  and  a49777a );
 a49788a <=( A234  and  (not A233) );
 a49791a <=( (not A298)  and  A236 );
 a49792a <=( a49791a  and  a49788a );
 a49795a <=( (not A300)  and  A299 );
 a49798a <=( (not A302)  and  (not A301) );
 a49799a <=( a49798a  and  a49795a );
 a49800a <=( a49799a  and  a49792a );
 a49803a <=( A168  and  A169 );
 a49806a <=( (not A166)  and  A167 );
 a49807a <=( a49806a  and  a49803a );
 a49810a <=( (not A202)  and  A201 );
 a49813a <=( A232  and  (not A203) );
 a49814a <=( a49813a  and  a49810a );
 a49815a <=( a49814a  and  a49807a );
 a49818a <=( A234  and  (not A233) );
 a49821a <=( (not A265)  and  A236 );
 a49822a <=( a49821a  and  a49818a );
 a49825a <=( (not A267)  and  A266 );
 a49828a <=( (not A269)  and  (not A268) );
 a49829a <=( a49828a  and  a49825a );
 a49830a <=( a49829a  and  a49822a );
 a49833a <=( A168  and  A169 );
 a49836a <=( (not A166)  and  A167 );
 a49837a <=( a49836a  and  a49833a );
 a49840a <=( (not A202)  and  A201 );
 a49843a <=( A232  and  (not A203) );
 a49844a <=( a49843a  and  a49840a );
 a49845a <=( a49844a  and  a49837a );
 a49848a <=( A234  and  (not A233) );
 a49851a <=( A265  and  A236 );
 a49852a <=( a49851a  and  a49848a );
 a49855a <=( (not A267)  and  (not A266) );
 a49858a <=( (not A269)  and  (not A268) );
 a49859a <=( a49858a  and  a49855a );
 a49860a <=( a49859a  and  a49852a );
 a49863a <=( A168  and  A169 );
 a49866a <=( (not A166)  and  A167 );
 a49867a <=( a49866a  and  a49863a );
 a49870a <=( (not A202)  and  A201 );
 a49873a <=( A232  and  (not A203) );
 a49874a <=( a49873a  and  a49870a );
 a49875a <=( a49874a  and  a49867a );
 a49878a <=( (not A234)  and  (not A233) );
 a49881a <=( (not A236)  and  (not A235) );
 a49882a <=( a49881a  and  a49878a );
 a49885a <=( (not A299)  and  A298 );
 a49888a <=( A301  and  A300 );
 a49889a <=( a49888a  and  a49885a );
 a49890a <=( a49889a  and  a49882a );
 a49893a <=( A168  and  A169 );
 a49896a <=( (not A166)  and  A167 );
 a49897a <=( a49896a  and  a49893a );
 a49900a <=( (not A202)  and  A201 );
 a49903a <=( A232  and  (not A203) );
 a49904a <=( a49903a  and  a49900a );
 a49905a <=( a49904a  and  a49897a );
 a49908a <=( (not A234)  and  (not A233) );
 a49911a <=( (not A236)  and  (not A235) );
 a49912a <=( a49911a  and  a49908a );
 a49915a <=( (not A299)  and  A298 );
 a49918a <=( A302  and  A300 );
 a49919a <=( a49918a  and  a49915a );
 a49920a <=( a49919a  and  a49912a );
 a49923a <=( A168  and  A169 );
 a49926a <=( (not A166)  and  A167 );
 a49927a <=( a49926a  and  a49923a );
 a49930a <=( (not A202)  and  A201 );
 a49933a <=( A232  and  (not A203) );
 a49934a <=( a49933a  and  a49930a );
 a49935a <=( a49934a  and  a49927a );
 a49938a <=( (not A234)  and  (not A233) );
 a49941a <=( (not A236)  and  (not A235) );
 a49942a <=( a49941a  and  a49938a );
 a49945a <=( A299  and  (not A298) );
 a49948a <=( A301  and  A300 );
 a49949a <=( a49948a  and  a49945a );
 a49950a <=( a49949a  and  a49942a );
 a49953a <=( A168  and  A169 );
 a49956a <=( (not A166)  and  A167 );
 a49957a <=( a49956a  and  a49953a );
 a49960a <=( (not A202)  and  A201 );
 a49963a <=( A232  and  (not A203) );
 a49964a <=( a49963a  and  a49960a );
 a49965a <=( a49964a  and  a49957a );
 a49968a <=( (not A234)  and  (not A233) );
 a49971a <=( (not A236)  and  (not A235) );
 a49972a <=( a49971a  and  a49968a );
 a49975a <=( A299  and  (not A298) );
 a49978a <=( A302  and  A300 );
 a49979a <=( a49978a  and  a49975a );
 a49980a <=( a49979a  and  a49972a );
 a49983a <=( A168  and  A169 );
 a49986a <=( (not A166)  and  A167 );
 a49987a <=( a49986a  and  a49983a );
 a49990a <=( (not A202)  and  A201 );
 a49993a <=( A232  and  (not A203) );
 a49994a <=( a49993a  and  a49990a );
 a49995a <=( a49994a  and  a49987a );
 a49998a <=( (not A234)  and  (not A233) );
 a50001a <=( (not A236)  and  (not A235) );
 a50002a <=( a50001a  and  a49998a );
 a50005a <=( A266  and  (not A265) );
 a50008a <=( A268  and  A267 );
 a50009a <=( a50008a  and  a50005a );
 a50010a <=( a50009a  and  a50002a );
 a50013a <=( A168  and  A169 );
 a50016a <=( (not A166)  and  A167 );
 a50017a <=( a50016a  and  a50013a );
 a50020a <=( (not A202)  and  A201 );
 a50023a <=( A232  and  (not A203) );
 a50024a <=( a50023a  and  a50020a );
 a50025a <=( a50024a  and  a50017a );
 a50028a <=( (not A234)  and  (not A233) );
 a50031a <=( (not A236)  and  (not A235) );
 a50032a <=( a50031a  and  a50028a );
 a50035a <=( A266  and  (not A265) );
 a50038a <=( A269  and  A267 );
 a50039a <=( a50038a  and  a50035a );
 a50040a <=( a50039a  and  a50032a );
 a50043a <=( A168  and  A169 );
 a50046a <=( (not A166)  and  A167 );
 a50047a <=( a50046a  and  a50043a );
 a50050a <=( (not A202)  and  A201 );
 a50053a <=( A232  and  (not A203) );
 a50054a <=( a50053a  and  a50050a );
 a50055a <=( a50054a  and  a50047a );
 a50058a <=( (not A234)  and  (not A233) );
 a50061a <=( (not A236)  and  (not A235) );
 a50062a <=( a50061a  and  a50058a );
 a50065a <=( (not A266)  and  A265 );
 a50068a <=( A268  and  A267 );
 a50069a <=( a50068a  and  a50065a );
 a50070a <=( a50069a  and  a50062a );
 a50073a <=( A168  and  A169 );
 a50076a <=( (not A166)  and  A167 );
 a50077a <=( a50076a  and  a50073a );
 a50080a <=( (not A202)  and  A201 );
 a50083a <=( A232  and  (not A203) );
 a50084a <=( a50083a  and  a50080a );
 a50085a <=( a50084a  and  a50077a );
 a50088a <=( (not A234)  and  (not A233) );
 a50091a <=( (not A236)  and  (not A235) );
 a50092a <=( a50091a  and  a50088a );
 a50095a <=( (not A266)  and  A265 );
 a50098a <=( A269  and  A267 );
 a50099a <=( a50098a  and  a50095a );
 a50100a <=( a50099a  and  a50092a );
 a50103a <=( A168  and  A169 );
 a50106a <=( (not A166)  and  A167 );
 a50107a <=( a50106a  and  a50103a );
 a50110a <=( A202  and  (not A201) );
 a50113a <=( A233  and  (not A232) );
 a50114a <=( a50113a  and  a50110a );
 a50115a <=( a50114a  and  a50107a );
 a50118a <=( (not A235)  and  (not A234) );
 a50121a <=( A298  and  (not A236) );
 a50122a <=( a50121a  and  a50118a );
 a50125a <=( (not A300)  and  (not A299) );
 a50128a <=( (not A302)  and  (not A301) );
 a50129a <=( a50128a  and  a50125a );
 a50130a <=( a50129a  and  a50122a );
 a50133a <=( A168  and  A169 );
 a50136a <=( (not A166)  and  A167 );
 a50137a <=( a50136a  and  a50133a );
 a50140a <=( A202  and  (not A201) );
 a50143a <=( A233  and  (not A232) );
 a50144a <=( a50143a  and  a50140a );
 a50145a <=( a50144a  and  a50137a );
 a50148a <=( (not A235)  and  (not A234) );
 a50151a <=( (not A298)  and  (not A236) );
 a50152a <=( a50151a  and  a50148a );
 a50155a <=( (not A300)  and  A299 );
 a50158a <=( (not A302)  and  (not A301) );
 a50159a <=( a50158a  and  a50155a );
 a50160a <=( a50159a  and  a50152a );
 a50163a <=( A168  and  A169 );
 a50166a <=( (not A166)  and  A167 );
 a50167a <=( a50166a  and  a50163a );
 a50170a <=( A202  and  (not A201) );
 a50173a <=( A233  and  (not A232) );
 a50174a <=( a50173a  and  a50170a );
 a50175a <=( a50174a  and  a50167a );
 a50178a <=( (not A235)  and  (not A234) );
 a50181a <=( (not A265)  and  (not A236) );
 a50182a <=( a50181a  and  a50178a );
 a50185a <=( (not A267)  and  A266 );
 a50188a <=( (not A269)  and  (not A268) );
 a50189a <=( a50188a  and  a50185a );
 a50190a <=( a50189a  and  a50182a );
 a50193a <=( A168  and  A169 );
 a50196a <=( (not A166)  and  A167 );
 a50197a <=( a50196a  and  a50193a );
 a50200a <=( A202  and  (not A201) );
 a50203a <=( A233  and  (not A232) );
 a50204a <=( a50203a  and  a50200a );
 a50205a <=( a50204a  and  a50197a );
 a50208a <=( (not A235)  and  (not A234) );
 a50211a <=( A265  and  (not A236) );
 a50212a <=( a50211a  and  a50208a );
 a50215a <=( (not A267)  and  (not A266) );
 a50218a <=( (not A269)  and  (not A268) );
 a50219a <=( a50218a  and  a50215a );
 a50220a <=( a50219a  and  a50212a );
 a50223a <=( A168  and  A169 );
 a50226a <=( (not A166)  and  A167 );
 a50227a <=( a50226a  and  a50223a );
 a50230a <=( A202  and  (not A201) );
 a50233a <=( (not A233)  and  A232 );
 a50234a <=( a50233a  and  a50230a );
 a50235a <=( a50234a  and  a50227a );
 a50238a <=( (not A235)  and  (not A234) );
 a50241a <=( A298  and  (not A236) );
 a50242a <=( a50241a  and  a50238a );
 a50245a <=( (not A300)  and  (not A299) );
 a50248a <=( (not A302)  and  (not A301) );
 a50249a <=( a50248a  and  a50245a );
 a50250a <=( a50249a  and  a50242a );
 a50253a <=( A168  and  A169 );
 a50256a <=( (not A166)  and  A167 );
 a50257a <=( a50256a  and  a50253a );
 a50260a <=( A202  and  (not A201) );
 a50263a <=( (not A233)  and  A232 );
 a50264a <=( a50263a  and  a50260a );
 a50265a <=( a50264a  and  a50257a );
 a50268a <=( (not A235)  and  (not A234) );
 a50271a <=( (not A298)  and  (not A236) );
 a50272a <=( a50271a  and  a50268a );
 a50275a <=( (not A300)  and  A299 );
 a50278a <=( (not A302)  and  (not A301) );
 a50279a <=( a50278a  and  a50275a );
 a50280a <=( a50279a  and  a50272a );
 a50283a <=( A168  and  A169 );
 a50286a <=( (not A166)  and  A167 );
 a50287a <=( a50286a  and  a50283a );
 a50290a <=( A202  and  (not A201) );
 a50293a <=( (not A233)  and  A232 );
 a50294a <=( a50293a  and  a50290a );
 a50295a <=( a50294a  and  a50287a );
 a50298a <=( (not A235)  and  (not A234) );
 a50301a <=( (not A265)  and  (not A236) );
 a50302a <=( a50301a  and  a50298a );
 a50305a <=( (not A267)  and  A266 );
 a50308a <=( (not A269)  and  (not A268) );
 a50309a <=( a50308a  and  a50305a );
 a50310a <=( a50309a  and  a50302a );
 a50313a <=( A168  and  A169 );
 a50316a <=( (not A166)  and  A167 );
 a50317a <=( a50316a  and  a50313a );
 a50320a <=( A202  and  (not A201) );
 a50323a <=( (not A233)  and  A232 );
 a50324a <=( a50323a  and  a50320a );
 a50325a <=( a50324a  and  a50317a );
 a50328a <=( (not A235)  and  (not A234) );
 a50331a <=( A265  and  (not A236) );
 a50332a <=( a50331a  and  a50328a );
 a50335a <=( (not A267)  and  (not A266) );
 a50338a <=( (not A269)  and  (not A268) );
 a50339a <=( a50338a  and  a50335a );
 a50340a <=( a50339a  and  a50332a );
 a50343a <=( A168  and  A169 );
 a50346a <=( (not A166)  and  A167 );
 a50347a <=( a50346a  and  a50343a );
 a50350a <=( A203  and  (not A201) );
 a50353a <=( A233  and  (not A232) );
 a50354a <=( a50353a  and  a50350a );
 a50355a <=( a50354a  and  a50347a );
 a50358a <=( (not A235)  and  (not A234) );
 a50361a <=( A298  and  (not A236) );
 a50362a <=( a50361a  and  a50358a );
 a50365a <=( (not A300)  and  (not A299) );
 a50368a <=( (not A302)  and  (not A301) );
 a50369a <=( a50368a  and  a50365a );
 a50370a <=( a50369a  and  a50362a );
 a50373a <=( A168  and  A169 );
 a50376a <=( (not A166)  and  A167 );
 a50377a <=( a50376a  and  a50373a );
 a50380a <=( A203  and  (not A201) );
 a50383a <=( A233  and  (not A232) );
 a50384a <=( a50383a  and  a50380a );
 a50385a <=( a50384a  and  a50377a );
 a50388a <=( (not A235)  and  (not A234) );
 a50391a <=( (not A298)  and  (not A236) );
 a50392a <=( a50391a  and  a50388a );
 a50395a <=( (not A300)  and  A299 );
 a50398a <=( (not A302)  and  (not A301) );
 a50399a <=( a50398a  and  a50395a );
 a50400a <=( a50399a  and  a50392a );
 a50403a <=( A168  and  A169 );
 a50406a <=( (not A166)  and  A167 );
 a50407a <=( a50406a  and  a50403a );
 a50410a <=( A203  and  (not A201) );
 a50413a <=( A233  and  (not A232) );
 a50414a <=( a50413a  and  a50410a );
 a50415a <=( a50414a  and  a50407a );
 a50418a <=( (not A235)  and  (not A234) );
 a50421a <=( (not A265)  and  (not A236) );
 a50422a <=( a50421a  and  a50418a );
 a50425a <=( (not A267)  and  A266 );
 a50428a <=( (not A269)  and  (not A268) );
 a50429a <=( a50428a  and  a50425a );
 a50430a <=( a50429a  and  a50422a );
 a50433a <=( A168  and  A169 );
 a50436a <=( (not A166)  and  A167 );
 a50437a <=( a50436a  and  a50433a );
 a50440a <=( A203  and  (not A201) );
 a50443a <=( A233  and  (not A232) );
 a50444a <=( a50443a  and  a50440a );
 a50445a <=( a50444a  and  a50437a );
 a50448a <=( (not A235)  and  (not A234) );
 a50451a <=( A265  and  (not A236) );
 a50452a <=( a50451a  and  a50448a );
 a50455a <=( (not A267)  and  (not A266) );
 a50458a <=( (not A269)  and  (not A268) );
 a50459a <=( a50458a  and  a50455a );
 a50460a <=( a50459a  and  a50452a );
 a50463a <=( A168  and  A169 );
 a50466a <=( (not A166)  and  A167 );
 a50467a <=( a50466a  and  a50463a );
 a50470a <=( A203  and  (not A201) );
 a50473a <=( (not A233)  and  A232 );
 a50474a <=( a50473a  and  a50470a );
 a50475a <=( a50474a  and  a50467a );
 a50478a <=( (not A235)  and  (not A234) );
 a50481a <=( A298  and  (not A236) );
 a50482a <=( a50481a  and  a50478a );
 a50485a <=( (not A300)  and  (not A299) );
 a50488a <=( (not A302)  and  (not A301) );
 a50489a <=( a50488a  and  a50485a );
 a50490a <=( a50489a  and  a50482a );
 a50493a <=( A168  and  A169 );
 a50496a <=( (not A166)  and  A167 );
 a50497a <=( a50496a  and  a50493a );
 a50500a <=( A203  and  (not A201) );
 a50503a <=( (not A233)  and  A232 );
 a50504a <=( a50503a  and  a50500a );
 a50505a <=( a50504a  and  a50497a );
 a50508a <=( (not A235)  and  (not A234) );
 a50511a <=( (not A298)  and  (not A236) );
 a50512a <=( a50511a  and  a50508a );
 a50515a <=( (not A300)  and  A299 );
 a50518a <=( (not A302)  and  (not A301) );
 a50519a <=( a50518a  and  a50515a );
 a50520a <=( a50519a  and  a50512a );
 a50523a <=( A168  and  A169 );
 a50526a <=( (not A166)  and  A167 );
 a50527a <=( a50526a  and  a50523a );
 a50530a <=( A203  and  (not A201) );
 a50533a <=( (not A233)  and  A232 );
 a50534a <=( a50533a  and  a50530a );
 a50535a <=( a50534a  and  a50527a );
 a50538a <=( (not A235)  and  (not A234) );
 a50541a <=( (not A265)  and  (not A236) );
 a50542a <=( a50541a  and  a50538a );
 a50545a <=( (not A267)  and  A266 );
 a50548a <=( (not A269)  and  (not A268) );
 a50549a <=( a50548a  and  a50545a );
 a50550a <=( a50549a  and  a50542a );
 a50553a <=( A168  and  A169 );
 a50556a <=( (not A166)  and  A167 );
 a50557a <=( a50556a  and  a50553a );
 a50560a <=( A203  and  (not A201) );
 a50563a <=( (not A233)  and  A232 );
 a50564a <=( a50563a  and  a50560a );
 a50565a <=( a50564a  and  a50557a );
 a50568a <=( (not A235)  and  (not A234) );
 a50571a <=( A265  and  (not A236) );
 a50572a <=( a50571a  and  a50568a );
 a50575a <=( (not A267)  and  (not A266) );
 a50578a <=( (not A269)  and  (not A268) );
 a50579a <=( a50578a  and  a50575a );
 a50580a <=( a50579a  and  a50572a );
 a50583a <=( A168  and  A169 );
 a50586a <=( (not A166)  and  A167 );
 a50587a <=( a50586a  and  a50583a );
 a50590a <=( A200  and  A199 );
 a50593a <=( A233  and  (not A232) );
 a50594a <=( a50593a  and  a50590a );
 a50595a <=( a50594a  and  a50587a );
 a50598a <=( (not A235)  and  (not A234) );
 a50601a <=( A298  and  (not A236) );
 a50602a <=( a50601a  and  a50598a );
 a50605a <=( (not A300)  and  (not A299) );
 a50608a <=( (not A302)  and  (not A301) );
 a50609a <=( a50608a  and  a50605a );
 a50610a <=( a50609a  and  a50602a );
 a50613a <=( A168  and  A169 );
 a50616a <=( (not A166)  and  A167 );
 a50617a <=( a50616a  and  a50613a );
 a50620a <=( A200  and  A199 );
 a50623a <=( A233  and  (not A232) );
 a50624a <=( a50623a  and  a50620a );
 a50625a <=( a50624a  and  a50617a );
 a50628a <=( (not A235)  and  (not A234) );
 a50631a <=( (not A298)  and  (not A236) );
 a50632a <=( a50631a  and  a50628a );
 a50635a <=( (not A300)  and  A299 );
 a50638a <=( (not A302)  and  (not A301) );
 a50639a <=( a50638a  and  a50635a );
 a50640a <=( a50639a  and  a50632a );
 a50643a <=( A168  and  A169 );
 a50646a <=( (not A166)  and  A167 );
 a50647a <=( a50646a  and  a50643a );
 a50650a <=( A200  and  A199 );
 a50653a <=( A233  and  (not A232) );
 a50654a <=( a50653a  and  a50650a );
 a50655a <=( a50654a  and  a50647a );
 a50658a <=( (not A235)  and  (not A234) );
 a50661a <=( (not A265)  and  (not A236) );
 a50662a <=( a50661a  and  a50658a );
 a50665a <=( (not A267)  and  A266 );
 a50668a <=( (not A269)  and  (not A268) );
 a50669a <=( a50668a  and  a50665a );
 a50670a <=( a50669a  and  a50662a );
 a50673a <=( A168  and  A169 );
 a50676a <=( (not A166)  and  A167 );
 a50677a <=( a50676a  and  a50673a );
 a50680a <=( A200  and  A199 );
 a50683a <=( A233  and  (not A232) );
 a50684a <=( a50683a  and  a50680a );
 a50685a <=( a50684a  and  a50677a );
 a50688a <=( (not A235)  and  (not A234) );
 a50691a <=( A265  and  (not A236) );
 a50692a <=( a50691a  and  a50688a );
 a50695a <=( (not A267)  and  (not A266) );
 a50698a <=( (not A269)  and  (not A268) );
 a50699a <=( a50698a  and  a50695a );
 a50700a <=( a50699a  and  a50692a );
 a50703a <=( A168  and  A169 );
 a50706a <=( (not A166)  and  A167 );
 a50707a <=( a50706a  and  a50703a );
 a50710a <=( A200  and  A199 );
 a50713a <=( (not A233)  and  A232 );
 a50714a <=( a50713a  and  a50710a );
 a50715a <=( a50714a  and  a50707a );
 a50718a <=( (not A235)  and  (not A234) );
 a50721a <=( A298  and  (not A236) );
 a50722a <=( a50721a  and  a50718a );
 a50725a <=( (not A300)  and  (not A299) );
 a50728a <=( (not A302)  and  (not A301) );
 a50729a <=( a50728a  and  a50725a );
 a50730a <=( a50729a  and  a50722a );
 a50733a <=( A168  and  A169 );
 a50736a <=( (not A166)  and  A167 );
 a50737a <=( a50736a  and  a50733a );
 a50740a <=( A200  and  A199 );
 a50743a <=( (not A233)  and  A232 );
 a50744a <=( a50743a  and  a50740a );
 a50745a <=( a50744a  and  a50737a );
 a50748a <=( (not A235)  and  (not A234) );
 a50751a <=( (not A298)  and  (not A236) );
 a50752a <=( a50751a  and  a50748a );
 a50755a <=( (not A300)  and  A299 );
 a50758a <=( (not A302)  and  (not A301) );
 a50759a <=( a50758a  and  a50755a );
 a50760a <=( a50759a  and  a50752a );
 a50763a <=( A168  and  A169 );
 a50766a <=( (not A166)  and  A167 );
 a50767a <=( a50766a  and  a50763a );
 a50770a <=( A200  and  A199 );
 a50773a <=( (not A233)  and  A232 );
 a50774a <=( a50773a  and  a50770a );
 a50775a <=( a50774a  and  a50767a );
 a50778a <=( (not A235)  and  (not A234) );
 a50781a <=( (not A265)  and  (not A236) );
 a50782a <=( a50781a  and  a50778a );
 a50785a <=( (not A267)  and  A266 );
 a50788a <=( (not A269)  and  (not A268) );
 a50789a <=( a50788a  and  a50785a );
 a50790a <=( a50789a  and  a50782a );
 a50793a <=( A168  and  A169 );
 a50796a <=( (not A166)  and  A167 );
 a50797a <=( a50796a  and  a50793a );
 a50800a <=( A200  and  A199 );
 a50803a <=( (not A233)  and  A232 );
 a50804a <=( a50803a  and  a50800a );
 a50805a <=( a50804a  and  a50797a );
 a50808a <=( (not A235)  and  (not A234) );
 a50811a <=( A265  and  (not A236) );
 a50812a <=( a50811a  and  a50808a );
 a50815a <=( (not A267)  and  (not A266) );
 a50818a <=( (not A269)  and  (not A268) );
 a50819a <=( a50818a  and  a50815a );
 a50820a <=( a50819a  and  a50812a );
 a50823a <=( A168  and  A169 );
 a50826a <=( (not A166)  and  A167 );
 a50827a <=( a50826a  and  a50823a );
 a50830a <=( (not A200)  and  (not A199) );
 a50833a <=( A233  and  (not A232) );
 a50834a <=( a50833a  and  a50830a );
 a50835a <=( a50834a  and  a50827a );
 a50838a <=( (not A235)  and  (not A234) );
 a50841a <=( A298  and  (not A236) );
 a50842a <=( a50841a  and  a50838a );
 a50845a <=( (not A300)  and  (not A299) );
 a50848a <=( (not A302)  and  (not A301) );
 a50849a <=( a50848a  and  a50845a );
 a50850a <=( a50849a  and  a50842a );
 a50853a <=( A168  and  A169 );
 a50856a <=( (not A166)  and  A167 );
 a50857a <=( a50856a  and  a50853a );
 a50860a <=( (not A200)  and  (not A199) );
 a50863a <=( A233  and  (not A232) );
 a50864a <=( a50863a  and  a50860a );
 a50865a <=( a50864a  and  a50857a );
 a50868a <=( (not A235)  and  (not A234) );
 a50871a <=( (not A298)  and  (not A236) );
 a50872a <=( a50871a  and  a50868a );
 a50875a <=( (not A300)  and  A299 );
 a50878a <=( (not A302)  and  (not A301) );
 a50879a <=( a50878a  and  a50875a );
 a50880a <=( a50879a  and  a50872a );
 a50883a <=( A168  and  A169 );
 a50886a <=( (not A166)  and  A167 );
 a50887a <=( a50886a  and  a50883a );
 a50890a <=( (not A200)  and  (not A199) );
 a50893a <=( A233  and  (not A232) );
 a50894a <=( a50893a  and  a50890a );
 a50895a <=( a50894a  and  a50887a );
 a50898a <=( (not A235)  and  (not A234) );
 a50901a <=( (not A265)  and  (not A236) );
 a50902a <=( a50901a  and  a50898a );
 a50905a <=( (not A267)  and  A266 );
 a50908a <=( (not A269)  and  (not A268) );
 a50909a <=( a50908a  and  a50905a );
 a50910a <=( a50909a  and  a50902a );
 a50913a <=( A168  and  A169 );
 a50916a <=( (not A166)  and  A167 );
 a50917a <=( a50916a  and  a50913a );
 a50920a <=( (not A200)  and  (not A199) );
 a50923a <=( A233  and  (not A232) );
 a50924a <=( a50923a  and  a50920a );
 a50925a <=( a50924a  and  a50917a );
 a50928a <=( (not A235)  and  (not A234) );
 a50931a <=( A265  and  (not A236) );
 a50932a <=( a50931a  and  a50928a );
 a50935a <=( (not A267)  and  (not A266) );
 a50938a <=( (not A269)  and  (not A268) );
 a50939a <=( a50938a  and  a50935a );
 a50940a <=( a50939a  and  a50932a );
 a50943a <=( A168  and  A169 );
 a50946a <=( (not A166)  and  A167 );
 a50947a <=( a50946a  and  a50943a );
 a50950a <=( (not A200)  and  (not A199) );
 a50953a <=( (not A233)  and  A232 );
 a50954a <=( a50953a  and  a50950a );
 a50955a <=( a50954a  and  a50947a );
 a50958a <=( (not A235)  and  (not A234) );
 a50961a <=( A298  and  (not A236) );
 a50962a <=( a50961a  and  a50958a );
 a50965a <=( (not A300)  and  (not A299) );
 a50968a <=( (not A302)  and  (not A301) );
 a50969a <=( a50968a  and  a50965a );
 a50970a <=( a50969a  and  a50962a );
 a50973a <=( A168  and  A169 );
 a50976a <=( (not A166)  and  A167 );
 a50977a <=( a50976a  and  a50973a );
 a50980a <=( (not A200)  and  (not A199) );
 a50983a <=( (not A233)  and  A232 );
 a50984a <=( a50983a  and  a50980a );
 a50985a <=( a50984a  and  a50977a );
 a50988a <=( (not A235)  and  (not A234) );
 a50991a <=( (not A298)  and  (not A236) );
 a50992a <=( a50991a  and  a50988a );
 a50995a <=( (not A300)  and  A299 );
 a50998a <=( (not A302)  and  (not A301) );
 a50999a <=( a50998a  and  a50995a );
 a51000a <=( a50999a  and  a50992a );
 a51003a <=( A168  and  A169 );
 a51006a <=( (not A166)  and  A167 );
 a51007a <=( a51006a  and  a51003a );
 a51010a <=( (not A200)  and  (not A199) );
 a51013a <=( (not A233)  and  A232 );
 a51014a <=( a51013a  and  a51010a );
 a51015a <=( a51014a  and  a51007a );
 a51018a <=( (not A235)  and  (not A234) );
 a51021a <=( (not A265)  and  (not A236) );
 a51022a <=( a51021a  and  a51018a );
 a51025a <=( (not A267)  and  A266 );
 a51028a <=( (not A269)  and  (not A268) );
 a51029a <=( a51028a  and  a51025a );
 a51030a <=( a51029a  and  a51022a );
 a51033a <=( A168  and  A169 );
 a51036a <=( (not A166)  and  A167 );
 a51037a <=( a51036a  and  a51033a );
 a51040a <=( (not A200)  and  (not A199) );
 a51043a <=( (not A233)  and  A232 );
 a51044a <=( a51043a  and  a51040a );
 a51045a <=( a51044a  and  a51037a );
 a51048a <=( (not A235)  and  (not A234) );
 a51051a <=( A265  and  (not A236) );
 a51052a <=( a51051a  and  a51048a );
 a51055a <=( (not A267)  and  (not A266) );
 a51058a <=( (not A269)  and  (not A268) );
 a51059a <=( a51058a  and  a51055a );
 a51060a <=( a51059a  and  a51052a );
 a51063a <=( A168  and  A169 );
 a51066a <=( A166  and  (not A167) );
 a51067a <=( a51066a  and  a51063a );
 a51070a <=( (not A202)  and  A201 );
 a51073a <=( (not A232)  and  (not A203) );
 a51074a <=( a51073a  and  a51070a );
 a51075a <=( a51074a  and  a51067a );
 a51078a <=( A234  and  A233 );
 a51081a <=( A298  and  A235 );
 a51082a <=( a51081a  and  a51078a );
 a51085a <=( (not A300)  and  (not A299) );
 a51088a <=( (not A302)  and  (not A301) );
 a51089a <=( a51088a  and  a51085a );
 a51090a <=( a51089a  and  a51082a );
 a51093a <=( A168  and  A169 );
 a51096a <=( A166  and  (not A167) );
 a51097a <=( a51096a  and  a51093a );
 a51100a <=( (not A202)  and  A201 );
 a51103a <=( (not A232)  and  (not A203) );
 a51104a <=( a51103a  and  a51100a );
 a51105a <=( a51104a  and  a51097a );
 a51108a <=( A234  and  A233 );
 a51111a <=( (not A298)  and  A235 );
 a51112a <=( a51111a  and  a51108a );
 a51115a <=( (not A300)  and  A299 );
 a51118a <=( (not A302)  and  (not A301) );
 a51119a <=( a51118a  and  a51115a );
 a51120a <=( a51119a  and  a51112a );
 a51123a <=( A168  and  A169 );
 a51126a <=( A166  and  (not A167) );
 a51127a <=( a51126a  and  a51123a );
 a51130a <=( (not A202)  and  A201 );
 a51133a <=( (not A232)  and  (not A203) );
 a51134a <=( a51133a  and  a51130a );
 a51135a <=( a51134a  and  a51127a );
 a51138a <=( A234  and  A233 );
 a51141a <=( (not A265)  and  A235 );
 a51142a <=( a51141a  and  a51138a );
 a51145a <=( (not A267)  and  A266 );
 a51148a <=( (not A269)  and  (not A268) );
 a51149a <=( a51148a  and  a51145a );
 a51150a <=( a51149a  and  a51142a );
 a51153a <=( A168  and  A169 );
 a51156a <=( A166  and  (not A167) );
 a51157a <=( a51156a  and  a51153a );
 a51160a <=( (not A202)  and  A201 );
 a51163a <=( (not A232)  and  (not A203) );
 a51164a <=( a51163a  and  a51160a );
 a51165a <=( a51164a  and  a51157a );
 a51168a <=( A234  and  A233 );
 a51171a <=( A265  and  A235 );
 a51172a <=( a51171a  and  a51168a );
 a51175a <=( (not A267)  and  (not A266) );
 a51178a <=( (not A269)  and  (not A268) );
 a51179a <=( a51178a  and  a51175a );
 a51180a <=( a51179a  and  a51172a );
 a51183a <=( A168  and  A169 );
 a51186a <=( A166  and  (not A167) );
 a51187a <=( a51186a  and  a51183a );
 a51190a <=( (not A202)  and  A201 );
 a51193a <=( (not A232)  and  (not A203) );
 a51194a <=( a51193a  and  a51190a );
 a51195a <=( a51194a  and  a51187a );
 a51198a <=( A234  and  A233 );
 a51201a <=( A298  and  A236 );
 a51202a <=( a51201a  and  a51198a );
 a51205a <=( (not A300)  and  (not A299) );
 a51208a <=( (not A302)  and  (not A301) );
 a51209a <=( a51208a  and  a51205a );
 a51210a <=( a51209a  and  a51202a );
 a51213a <=( A168  and  A169 );
 a51216a <=( A166  and  (not A167) );
 a51217a <=( a51216a  and  a51213a );
 a51220a <=( (not A202)  and  A201 );
 a51223a <=( (not A232)  and  (not A203) );
 a51224a <=( a51223a  and  a51220a );
 a51225a <=( a51224a  and  a51217a );
 a51228a <=( A234  and  A233 );
 a51231a <=( (not A298)  and  A236 );
 a51232a <=( a51231a  and  a51228a );
 a51235a <=( (not A300)  and  A299 );
 a51238a <=( (not A302)  and  (not A301) );
 a51239a <=( a51238a  and  a51235a );
 a51240a <=( a51239a  and  a51232a );
 a51243a <=( A168  and  A169 );
 a51246a <=( A166  and  (not A167) );
 a51247a <=( a51246a  and  a51243a );
 a51250a <=( (not A202)  and  A201 );
 a51253a <=( (not A232)  and  (not A203) );
 a51254a <=( a51253a  and  a51250a );
 a51255a <=( a51254a  and  a51247a );
 a51258a <=( A234  and  A233 );
 a51261a <=( (not A265)  and  A236 );
 a51262a <=( a51261a  and  a51258a );
 a51265a <=( (not A267)  and  A266 );
 a51268a <=( (not A269)  and  (not A268) );
 a51269a <=( a51268a  and  a51265a );
 a51270a <=( a51269a  and  a51262a );
 a51273a <=( A168  and  A169 );
 a51276a <=( A166  and  (not A167) );
 a51277a <=( a51276a  and  a51273a );
 a51280a <=( (not A202)  and  A201 );
 a51283a <=( (not A232)  and  (not A203) );
 a51284a <=( a51283a  and  a51280a );
 a51285a <=( a51284a  and  a51277a );
 a51288a <=( A234  and  A233 );
 a51291a <=( A265  and  A236 );
 a51292a <=( a51291a  and  a51288a );
 a51295a <=( (not A267)  and  (not A266) );
 a51298a <=( (not A269)  and  (not A268) );
 a51299a <=( a51298a  and  a51295a );
 a51300a <=( a51299a  and  a51292a );
 a51303a <=( A168  and  A169 );
 a51306a <=( A166  and  (not A167) );
 a51307a <=( a51306a  and  a51303a );
 a51310a <=( (not A202)  and  A201 );
 a51313a <=( (not A232)  and  (not A203) );
 a51314a <=( a51313a  and  a51310a );
 a51315a <=( a51314a  and  a51307a );
 a51318a <=( (not A234)  and  A233 );
 a51321a <=( (not A236)  and  (not A235) );
 a51322a <=( a51321a  and  a51318a );
 a51325a <=( (not A299)  and  A298 );
 a51328a <=( A301  and  A300 );
 a51329a <=( a51328a  and  a51325a );
 a51330a <=( a51329a  and  a51322a );
 a51333a <=( A168  and  A169 );
 a51336a <=( A166  and  (not A167) );
 a51337a <=( a51336a  and  a51333a );
 a51340a <=( (not A202)  and  A201 );
 a51343a <=( (not A232)  and  (not A203) );
 a51344a <=( a51343a  and  a51340a );
 a51345a <=( a51344a  and  a51337a );
 a51348a <=( (not A234)  and  A233 );
 a51351a <=( (not A236)  and  (not A235) );
 a51352a <=( a51351a  and  a51348a );
 a51355a <=( (not A299)  and  A298 );
 a51358a <=( A302  and  A300 );
 a51359a <=( a51358a  and  a51355a );
 a51360a <=( a51359a  and  a51352a );
 a51363a <=( A168  and  A169 );
 a51366a <=( A166  and  (not A167) );
 a51367a <=( a51366a  and  a51363a );
 a51370a <=( (not A202)  and  A201 );
 a51373a <=( (not A232)  and  (not A203) );
 a51374a <=( a51373a  and  a51370a );
 a51375a <=( a51374a  and  a51367a );
 a51378a <=( (not A234)  and  A233 );
 a51381a <=( (not A236)  and  (not A235) );
 a51382a <=( a51381a  and  a51378a );
 a51385a <=( A299  and  (not A298) );
 a51388a <=( A301  and  A300 );
 a51389a <=( a51388a  and  a51385a );
 a51390a <=( a51389a  and  a51382a );
 a51393a <=( A168  and  A169 );
 a51396a <=( A166  and  (not A167) );
 a51397a <=( a51396a  and  a51393a );
 a51400a <=( (not A202)  and  A201 );
 a51403a <=( (not A232)  and  (not A203) );
 a51404a <=( a51403a  and  a51400a );
 a51405a <=( a51404a  and  a51397a );
 a51408a <=( (not A234)  and  A233 );
 a51411a <=( (not A236)  and  (not A235) );
 a51412a <=( a51411a  and  a51408a );
 a51415a <=( A299  and  (not A298) );
 a51418a <=( A302  and  A300 );
 a51419a <=( a51418a  and  a51415a );
 a51420a <=( a51419a  and  a51412a );
 a51423a <=( A168  and  A169 );
 a51426a <=( A166  and  (not A167) );
 a51427a <=( a51426a  and  a51423a );
 a51430a <=( (not A202)  and  A201 );
 a51433a <=( (not A232)  and  (not A203) );
 a51434a <=( a51433a  and  a51430a );
 a51435a <=( a51434a  and  a51427a );
 a51438a <=( (not A234)  and  A233 );
 a51441a <=( (not A236)  and  (not A235) );
 a51442a <=( a51441a  and  a51438a );
 a51445a <=( A266  and  (not A265) );
 a51448a <=( A268  and  A267 );
 a51449a <=( a51448a  and  a51445a );
 a51450a <=( a51449a  and  a51442a );
 a51453a <=( A168  and  A169 );
 a51456a <=( A166  and  (not A167) );
 a51457a <=( a51456a  and  a51453a );
 a51460a <=( (not A202)  and  A201 );
 a51463a <=( (not A232)  and  (not A203) );
 a51464a <=( a51463a  and  a51460a );
 a51465a <=( a51464a  and  a51457a );
 a51468a <=( (not A234)  and  A233 );
 a51471a <=( (not A236)  and  (not A235) );
 a51472a <=( a51471a  and  a51468a );
 a51475a <=( A266  and  (not A265) );
 a51478a <=( A269  and  A267 );
 a51479a <=( a51478a  and  a51475a );
 a51480a <=( a51479a  and  a51472a );
 a51483a <=( A168  and  A169 );
 a51486a <=( A166  and  (not A167) );
 a51487a <=( a51486a  and  a51483a );
 a51490a <=( (not A202)  and  A201 );
 a51493a <=( (not A232)  and  (not A203) );
 a51494a <=( a51493a  and  a51490a );
 a51495a <=( a51494a  and  a51487a );
 a51498a <=( (not A234)  and  A233 );
 a51501a <=( (not A236)  and  (not A235) );
 a51502a <=( a51501a  and  a51498a );
 a51505a <=( (not A266)  and  A265 );
 a51508a <=( A268  and  A267 );
 a51509a <=( a51508a  and  a51505a );
 a51510a <=( a51509a  and  a51502a );
 a51513a <=( A168  and  A169 );
 a51516a <=( A166  and  (not A167) );
 a51517a <=( a51516a  and  a51513a );
 a51520a <=( (not A202)  and  A201 );
 a51523a <=( (not A232)  and  (not A203) );
 a51524a <=( a51523a  and  a51520a );
 a51525a <=( a51524a  and  a51517a );
 a51528a <=( (not A234)  and  A233 );
 a51531a <=( (not A236)  and  (not A235) );
 a51532a <=( a51531a  and  a51528a );
 a51535a <=( (not A266)  and  A265 );
 a51538a <=( A269  and  A267 );
 a51539a <=( a51538a  and  a51535a );
 a51540a <=( a51539a  and  a51532a );
 a51543a <=( A168  and  A169 );
 a51546a <=( A166  and  (not A167) );
 a51547a <=( a51546a  and  a51543a );
 a51550a <=( (not A202)  and  A201 );
 a51553a <=( A232  and  (not A203) );
 a51554a <=( a51553a  and  a51550a );
 a51555a <=( a51554a  and  a51547a );
 a51558a <=( A234  and  (not A233) );
 a51561a <=( A298  and  A235 );
 a51562a <=( a51561a  and  a51558a );
 a51565a <=( (not A300)  and  (not A299) );
 a51568a <=( (not A302)  and  (not A301) );
 a51569a <=( a51568a  and  a51565a );
 a51570a <=( a51569a  and  a51562a );
 a51573a <=( A168  and  A169 );
 a51576a <=( A166  and  (not A167) );
 a51577a <=( a51576a  and  a51573a );
 a51580a <=( (not A202)  and  A201 );
 a51583a <=( A232  and  (not A203) );
 a51584a <=( a51583a  and  a51580a );
 a51585a <=( a51584a  and  a51577a );
 a51588a <=( A234  and  (not A233) );
 a51591a <=( (not A298)  and  A235 );
 a51592a <=( a51591a  and  a51588a );
 a51595a <=( (not A300)  and  A299 );
 a51598a <=( (not A302)  and  (not A301) );
 a51599a <=( a51598a  and  a51595a );
 a51600a <=( a51599a  and  a51592a );
 a51603a <=( A168  and  A169 );
 a51606a <=( A166  and  (not A167) );
 a51607a <=( a51606a  and  a51603a );
 a51610a <=( (not A202)  and  A201 );
 a51613a <=( A232  and  (not A203) );
 a51614a <=( a51613a  and  a51610a );
 a51615a <=( a51614a  and  a51607a );
 a51618a <=( A234  and  (not A233) );
 a51621a <=( (not A265)  and  A235 );
 a51622a <=( a51621a  and  a51618a );
 a51625a <=( (not A267)  and  A266 );
 a51628a <=( (not A269)  and  (not A268) );
 a51629a <=( a51628a  and  a51625a );
 a51630a <=( a51629a  and  a51622a );
 a51633a <=( A168  and  A169 );
 a51636a <=( A166  and  (not A167) );
 a51637a <=( a51636a  and  a51633a );
 a51640a <=( (not A202)  and  A201 );
 a51643a <=( A232  and  (not A203) );
 a51644a <=( a51643a  and  a51640a );
 a51645a <=( a51644a  and  a51637a );
 a51648a <=( A234  and  (not A233) );
 a51651a <=( A265  and  A235 );
 a51652a <=( a51651a  and  a51648a );
 a51655a <=( (not A267)  and  (not A266) );
 a51658a <=( (not A269)  and  (not A268) );
 a51659a <=( a51658a  and  a51655a );
 a51660a <=( a51659a  and  a51652a );
 a51663a <=( A168  and  A169 );
 a51666a <=( A166  and  (not A167) );
 a51667a <=( a51666a  and  a51663a );
 a51670a <=( (not A202)  and  A201 );
 a51673a <=( A232  and  (not A203) );
 a51674a <=( a51673a  and  a51670a );
 a51675a <=( a51674a  and  a51667a );
 a51678a <=( A234  and  (not A233) );
 a51681a <=( A298  and  A236 );
 a51682a <=( a51681a  and  a51678a );
 a51685a <=( (not A300)  and  (not A299) );
 a51688a <=( (not A302)  and  (not A301) );
 a51689a <=( a51688a  and  a51685a );
 a51690a <=( a51689a  and  a51682a );
 a51693a <=( A168  and  A169 );
 a51696a <=( A166  and  (not A167) );
 a51697a <=( a51696a  and  a51693a );
 a51700a <=( (not A202)  and  A201 );
 a51703a <=( A232  and  (not A203) );
 a51704a <=( a51703a  and  a51700a );
 a51705a <=( a51704a  and  a51697a );
 a51708a <=( A234  and  (not A233) );
 a51711a <=( (not A298)  and  A236 );
 a51712a <=( a51711a  and  a51708a );
 a51715a <=( (not A300)  and  A299 );
 a51718a <=( (not A302)  and  (not A301) );
 a51719a <=( a51718a  and  a51715a );
 a51720a <=( a51719a  and  a51712a );
 a51723a <=( A168  and  A169 );
 a51726a <=( A166  and  (not A167) );
 a51727a <=( a51726a  and  a51723a );
 a51730a <=( (not A202)  and  A201 );
 a51733a <=( A232  and  (not A203) );
 a51734a <=( a51733a  and  a51730a );
 a51735a <=( a51734a  and  a51727a );
 a51738a <=( A234  and  (not A233) );
 a51741a <=( (not A265)  and  A236 );
 a51742a <=( a51741a  and  a51738a );
 a51745a <=( (not A267)  and  A266 );
 a51748a <=( (not A269)  and  (not A268) );
 a51749a <=( a51748a  and  a51745a );
 a51750a <=( a51749a  and  a51742a );
 a51753a <=( A168  and  A169 );
 a51756a <=( A166  and  (not A167) );
 a51757a <=( a51756a  and  a51753a );
 a51760a <=( (not A202)  and  A201 );
 a51763a <=( A232  and  (not A203) );
 a51764a <=( a51763a  and  a51760a );
 a51765a <=( a51764a  and  a51757a );
 a51768a <=( A234  and  (not A233) );
 a51771a <=( A265  and  A236 );
 a51772a <=( a51771a  and  a51768a );
 a51775a <=( (not A267)  and  (not A266) );
 a51778a <=( (not A269)  and  (not A268) );
 a51779a <=( a51778a  and  a51775a );
 a51780a <=( a51779a  and  a51772a );
 a51783a <=( A168  and  A169 );
 a51786a <=( A166  and  (not A167) );
 a51787a <=( a51786a  and  a51783a );
 a51790a <=( (not A202)  and  A201 );
 a51793a <=( A232  and  (not A203) );
 a51794a <=( a51793a  and  a51790a );
 a51795a <=( a51794a  and  a51787a );
 a51798a <=( (not A234)  and  (not A233) );
 a51801a <=( (not A236)  and  (not A235) );
 a51802a <=( a51801a  and  a51798a );
 a51805a <=( (not A299)  and  A298 );
 a51808a <=( A301  and  A300 );
 a51809a <=( a51808a  and  a51805a );
 a51810a <=( a51809a  and  a51802a );
 a51813a <=( A168  and  A169 );
 a51816a <=( A166  and  (not A167) );
 a51817a <=( a51816a  and  a51813a );
 a51820a <=( (not A202)  and  A201 );
 a51823a <=( A232  and  (not A203) );
 a51824a <=( a51823a  and  a51820a );
 a51825a <=( a51824a  and  a51817a );
 a51828a <=( (not A234)  and  (not A233) );
 a51831a <=( (not A236)  and  (not A235) );
 a51832a <=( a51831a  and  a51828a );
 a51835a <=( (not A299)  and  A298 );
 a51838a <=( A302  and  A300 );
 a51839a <=( a51838a  and  a51835a );
 a51840a <=( a51839a  and  a51832a );
 a51843a <=( A168  and  A169 );
 a51846a <=( A166  and  (not A167) );
 a51847a <=( a51846a  and  a51843a );
 a51850a <=( (not A202)  and  A201 );
 a51853a <=( A232  and  (not A203) );
 a51854a <=( a51853a  and  a51850a );
 a51855a <=( a51854a  and  a51847a );
 a51858a <=( (not A234)  and  (not A233) );
 a51861a <=( (not A236)  and  (not A235) );
 a51862a <=( a51861a  and  a51858a );
 a51865a <=( A299  and  (not A298) );
 a51868a <=( A301  and  A300 );
 a51869a <=( a51868a  and  a51865a );
 a51870a <=( a51869a  and  a51862a );
 a51873a <=( A168  and  A169 );
 a51876a <=( A166  and  (not A167) );
 a51877a <=( a51876a  and  a51873a );
 a51880a <=( (not A202)  and  A201 );
 a51883a <=( A232  and  (not A203) );
 a51884a <=( a51883a  and  a51880a );
 a51885a <=( a51884a  and  a51877a );
 a51888a <=( (not A234)  and  (not A233) );
 a51891a <=( (not A236)  and  (not A235) );
 a51892a <=( a51891a  and  a51888a );
 a51895a <=( A299  and  (not A298) );
 a51898a <=( A302  and  A300 );
 a51899a <=( a51898a  and  a51895a );
 a51900a <=( a51899a  and  a51892a );
 a51903a <=( A168  and  A169 );
 a51906a <=( A166  and  (not A167) );
 a51907a <=( a51906a  and  a51903a );
 a51910a <=( (not A202)  and  A201 );
 a51913a <=( A232  and  (not A203) );
 a51914a <=( a51913a  and  a51910a );
 a51915a <=( a51914a  and  a51907a );
 a51918a <=( (not A234)  and  (not A233) );
 a51921a <=( (not A236)  and  (not A235) );
 a51922a <=( a51921a  and  a51918a );
 a51925a <=( A266  and  (not A265) );
 a51928a <=( A268  and  A267 );
 a51929a <=( a51928a  and  a51925a );
 a51930a <=( a51929a  and  a51922a );
 a51933a <=( A168  and  A169 );
 a51936a <=( A166  and  (not A167) );
 a51937a <=( a51936a  and  a51933a );
 a51940a <=( (not A202)  and  A201 );
 a51943a <=( A232  and  (not A203) );
 a51944a <=( a51943a  and  a51940a );
 a51945a <=( a51944a  and  a51937a );
 a51948a <=( (not A234)  and  (not A233) );
 a51951a <=( (not A236)  and  (not A235) );
 a51952a <=( a51951a  and  a51948a );
 a51955a <=( A266  and  (not A265) );
 a51958a <=( A269  and  A267 );
 a51959a <=( a51958a  and  a51955a );
 a51960a <=( a51959a  and  a51952a );
 a51963a <=( A168  and  A169 );
 a51966a <=( A166  and  (not A167) );
 a51967a <=( a51966a  and  a51963a );
 a51970a <=( (not A202)  and  A201 );
 a51973a <=( A232  and  (not A203) );
 a51974a <=( a51973a  and  a51970a );
 a51975a <=( a51974a  and  a51967a );
 a51978a <=( (not A234)  and  (not A233) );
 a51981a <=( (not A236)  and  (not A235) );
 a51982a <=( a51981a  and  a51978a );
 a51985a <=( (not A266)  and  A265 );
 a51988a <=( A268  and  A267 );
 a51989a <=( a51988a  and  a51985a );
 a51990a <=( a51989a  and  a51982a );
 a51993a <=( A168  and  A169 );
 a51996a <=( A166  and  (not A167) );
 a51997a <=( a51996a  and  a51993a );
 a52000a <=( (not A202)  and  A201 );
 a52003a <=( A232  and  (not A203) );
 a52004a <=( a52003a  and  a52000a );
 a52005a <=( a52004a  and  a51997a );
 a52008a <=( (not A234)  and  (not A233) );
 a52011a <=( (not A236)  and  (not A235) );
 a52012a <=( a52011a  and  a52008a );
 a52015a <=( (not A266)  and  A265 );
 a52018a <=( A269  and  A267 );
 a52019a <=( a52018a  and  a52015a );
 a52020a <=( a52019a  and  a52012a );
 a52023a <=( A168  and  A169 );
 a52026a <=( A166  and  (not A167) );
 a52027a <=( a52026a  and  a52023a );
 a52030a <=( A202  and  (not A201) );
 a52033a <=( A233  and  (not A232) );
 a52034a <=( a52033a  and  a52030a );
 a52035a <=( a52034a  and  a52027a );
 a52038a <=( (not A235)  and  (not A234) );
 a52041a <=( A298  and  (not A236) );
 a52042a <=( a52041a  and  a52038a );
 a52045a <=( (not A300)  and  (not A299) );
 a52048a <=( (not A302)  and  (not A301) );
 a52049a <=( a52048a  and  a52045a );
 a52050a <=( a52049a  and  a52042a );
 a52053a <=( A168  and  A169 );
 a52056a <=( A166  and  (not A167) );
 a52057a <=( a52056a  and  a52053a );
 a52060a <=( A202  and  (not A201) );
 a52063a <=( A233  and  (not A232) );
 a52064a <=( a52063a  and  a52060a );
 a52065a <=( a52064a  and  a52057a );
 a52068a <=( (not A235)  and  (not A234) );
 a52071a <=( (not A298)  and  (not A236) );
 a52072a <=( a52071a  and  a52068a );
 a52075a <=( (not A300)  and  A299 );
 a52078a <=( (not A302)  and  (not A301) );
 a52079a <=( a52078a  and  a52075a );
 a52080a <=( a52079a  and  a52072a );
 a52083a <=( A168  and  A169 );
 a52086a <=( A166  and  (not A167) );
 a52087a <=( a52086a  and  a52083a );
 a52090a <=( A202  and  (not A201) );
 a52093a <=( A233  and  (not A232) );
 a52094a <=( a52093a  and  a52090a );
 a52095a <=( a52094a  and  a52087a );
 a52098a <=( (not A235)  and  (not A234) );
 a52101a <=( (not A265)  and  (not A236) );
 a52102a <=( a52101a  and  a52098a );
 a52105a <=( (not A267)  and  A266 );
 a52108a <=( (not A269)  and  (not A268) );
 a52109a <=( a52108a  and  a52105a );
 a52110a <=( a52109a  and  a52102a );
 a52113a <=( A168  and  A169 );
 a52116a <=( A166  and  (not A167) );
 a52117a <=( a52116a  and  a52113a );
 a52120a <=( A202  and  (not A201) );
 a52123a <=( A233  and  (not A232) );
 a52124a <=( a52123a  and  a52120a );
 a52125a <=( a52124a  and  a52117a );
 a52128a <=( (not A235)  and  (not A234) );
 a52131a <=( A265  and  (not A236) );
 a52132a <=( a52131a  and  a52128a );
 a52135a <=( (not A267)  and  (not A266) );
 a52138a <=( (not A269)  and  (not A268) );
 a52139a <=( a52138a  and  a52135a );
 a52140a <=( a52139a  and  a52132a );
 a52143a <=( A168  and  A169 );
 a52146a <=( A166  and  (not A167) );
 a52147a <=( a52146a  and  a52143a );
 a52150a <=( A202  and  (not A201) );
 a52153a <=( (not A233)  and  A232 );
 a52154a <=( a52153a  and  a52150a );
 a52155a <=( a52154a  and  a52147a );
 a52158a <=( (not A235)  and  (not A234) );
 a52161a <=( A298  and  (not A236) );
 a52162a <=( a52161a  and  a52158a );
 a52165a <=( (not A300)  and  (not A299) );
 a52168a <=( (not A302)  and  (not A301) );
 a52169a <=( a52168a  and  a52165a );
 a52170a <=( a52169a  and  a52162a );
 a52173a <=( A168  and  A169 );
 a52176a <=( A166  and  (not A167) );
 a52177a <=( a52176a  and  a52173a );
 a52180a <=( A202  and  (not A201) );
 a52183a <=( (not A233)  and  A232 );
 a52184a <=( a52183a  and  a52180a );
 a52185a <=( a52184a  and  a52177a );
 a52188a <=( (not A235)  and  (not A234) );
 a52191a <=( (not A298)  and  (not A236) );
 a52192a <=( a52191a  and  a52188a );
 a52195a <=( (not A300)  and  A299 );
 a52198a <=( (not A302)  and  (not A301) );
 a52199a <=( a52198a  and  a52195a );
 a52200a <=( a52199a  and  a52192a );
 a52203a <=( A168  and  A169 );
 a52206a <=( A166  and  (not A167) );
 a52207a <=( a52206a  and  a52203a );
 a52210a <=( A202  and  (not A201) );
 a52213a <=( (not A233)  and  A232 );
 a52214a <=( a52213a  and  a52210a );
 a52215a <=( a52214a  and  a52207a );
 a52218a <=( (not A235)  and  (not A234) );
 a52221a <=( (not A265)  and  (not A236) );
 a52222a <=( a52221a  and  a52218a );
 a52225a <=( (not A267)  and  A266 );
 a52228a <=( (not A269)  and  (not A268) );
 a52229a <=( a52228a  and  a52225a );
 a52230a <=( a52229a  and  a52222a );
 a52233a <=( A168  and  A169 );
 a52236a <=( A166  and  (not A167) );
 a52237a <=( a52236a  and  a52233a );
 a52240a <=( A202  and  (not A201) );
 a52243a <=( (not A233)  and  A232 );
 a52244a <=( a52243a  and  a52240a );
 a52245a <=( a52244a  and  a52237a );
 a52248a <=( (not A235)  and  (not A234) );
 a52251a <=( A265  and  (not A236) );
 a52252a <=( a52251a  and  a52248a );
 a52255a <=( (not A267)  and  (not A266) );
 a52258a <=( (not A269)  and  (not A268) );
 a52259a <=( a52258a  and  a52255a );
 a52260a <=( a52259a  and  a52252a );
 a52263a <=( A168  and  A169 );
 a52266a <=( A166  and  (not A167) );
 a52267a <=( a52266a  and  a52263a );
 a52270a <=( A203  and  (not A201) );
 a52273a <=( A233  and  (not A232) );
 a52274a <=( a52273a  and  a52270a );
 a52275a <=( a52274a  and  a52267a );
 a52278a <=( (not A235)  and  (not A234) );
 a52281a <=( A298  and  (not A236) );
 a52282a <=( a52281a  and  a52278a );
 a52285a <=( (not A300)  and  (not A299) );
 a52288a <=( (not A302)  and  (not A301) );
 a52289a <=( a52288a  and  a52285a );
 a52290a <=( a52289a  and  a52282a );
 a52293a <=( A168  and  A169 );
 a52296a <=( A166  and  (not A167) );
 a52297a <=( a52296a  and  a52293a );
 a52300a <=( A203  and  (not A201) );
 a52303a <=( A233  and  (not A232) );
 a52304a <=( a52303a  and  a52300a );
 a52305a <=( a52304a  and  a52297a );
 a52308a <=( (not A235)  and  (not A234) );
 a52311a <=( (not A298)  and  (not A236) );
 a52312a <=( a52311a  and  a52308a );
 a52315a <=( (not A300)  and  A299 );
 a52318a <=( (not A302)  and  (not A301) );
 a52319a <=( a52318a  and  a52315a );
 a52320a <=( a52319a  and  a52312a );
 a52323a <=( A168  and  A169 );
 a52326a <=( A166  and  (not A167) );
 a52327a <=( a52326a  and  a52323a );
 a52330a <=( A203  and  (not A201) );
 a52333a <=( A233  and  (not A232) );
 a52334a <=( a52333a  and  a52330a );
 a52335a <=( a52334a  and  a52327a );
 a52338a <=( (not A235)  and  (not A234) );
 a52341a <=( (not A265)  and  (not A236) );
 a52342a <=( a52341a  and  a52338a );
 a52345a <=( (not A267)  and  A266 );
 a52348a <=( (not A269)  and  (not A268) );
 a52349a <=( a52348a  and  a52345a );
 a52350a <=( a52349a  and  a52342a );
 a52353a <=( A168  and  A169 );
 a52356a <=( A166  and  (not A167) );
 a52357a <=( a52356a  and  a52353a );
 a52360a <=( A203  and  (not A201) );
 a52363a <=( A233  and  (not A232) );
 a52364a <=( a52363a  and  a52360a );
 a52365a <=( a52364a  and  a52357a );
 a52368a <=( (not A235)  and  (not A234) );
 a52371a <=( A265  and  (not A236) );
 a52372a <=( a52371a  and  a52368a );
 a52375a <=( (not A267)  and  (not A266) );
 a52378a <=( (not A269)  and  (not A268) );
 a52379a <=( a52378a  and  a52375a );
 a52380a <=( a52379a  and  a52372a );
 a52383a <=( A168  and  A169 );
 a52386a <=( A166  and  (not A167) );
 a52387a <=( a52386a  and  a52383a );
 a52390a <=( A203  and  (not A201) );
 a52393a <=( (not A233)  and  A232 );
 a52394a <=( a52393a  and  a52390a );
 a52395a <=( a52394a  and  a52387a );
 a52398a <=( (not A235)  and  (not A234) );
 a52401a <=( A298  and  (not A236) );
 a52402a <=( a52401a  and  a52398a );
 a52405a <=( (not A300)  and  (not A299) );
 a52408a <=( (not A302)  and  (not A301) );
 a52409a <=( a52408a  and  a52405a );
 a52410a <=( a52409a  and  a52402a );
 a52413a <=( A168  and  A169 );
 a52416a <=( A166  and  (not A167) );
 a52417a <=( a52416a  and  a52413a );
 a52420a <=( A203  and  (not A201) );
 a52423a <=( (not A233)  and  A232 );
 a52424a <=( a52423a  and  a52420a );
 a52425a <=( a52424a  and  a52417a );
 a52428a <=( (not A235)  and  (not A234) );
 a52431a <=( (not A298)  and  (not A236) );
 a52432a <=( a52431a  and  a52428a );
 a52435a <=( (not A300)  and  A299 );
 a52438a <=( (not A302)  and  (not A301) );
 a52439a <=( a52438a  and  a52435a );
 a52440a <=( a52439a  and  a52432a );
 a52443a <=( A168  and  A169 );
 a52446a <=( A166  and  (not A167) );
 a52447a <=( a52446a  and  a52443a );
 a52450a <=( A203  and  (not A201) );
 a52453a <=( (not A233)  and  A232 );
 a52454a <=( a52453a  and  a52450a );
 a52455a <=( a52454a  and  a52447a );
 a52458a <=( (not A235)  and  (not A234) );
 a52461a <=( (not A265)  and  (not A236) );
 a52462a <=( a52461a  and  a52458a );
 a52465a <=( (not A267)  and  A266 );
 a52468a <=( (not A269)  and  (not A268) );
 a52469a <=( a52468a  and  a52465a );
 a52470a <=( a52469a  and  a52462a );
 a52473a <=( A168  and  A169 );
 a52476a <=( A166  and  (not A167) );
 a52477a <=( a52476a  and  a52473a );
 a52480a <=( A203  and  (not A201) );
 a52483a <=( (not A233)  and  A232 );
 a52484a <=( a52483a  and  a52480a );
 a52485a <=( a52484a  and  a52477a );
 a52488a <=( (not A235)  and  (not A234) );
 a52491a <=( A265  and  (not A236) );
 a52492a <=( a52491a  and  a52488a );
 a52495a <=( (not A267)  and  (not A266) );
 a52498a <=( (not A269)  and  (not A268) );
 a52499a <=( a52498a  and  a52495a );
 a52500a <=( a52499a  and  a52492a );
 a52503a <=( A168  and  A169 );
 a52506a <=( A166  and  (not A167) );
 a52507a <=( a52506a  and  a52503a );
 a52510a <=( A200  and  A199 );
 a52513a <=( A233  and  (not A232) );
 a52514a <=( a52513a  and  a52510a );
 a52515a <=( a52514a  and  a52507a );
 a52518a <=( (not A235)  and  (not A234) );
 a52521a <=( A298  and  (not A236) );
 a52522a <=( a52521a  and  a52518a );
 a52525a <=( (not A300)  and  (not A299) );
 a52528a <=( (not A302)  and  (not A301) );
 a52529a <=( a52528a  and  a52525a );
 a52530a <=( a52529a  and  a52522a );
 a52533a <=( A168  and  A169 );
 a52536a <=( A166  and  (not A167) );
 a52537a <=( a52536a  and  a52533a );
 a52540a <=( A200  and  A199 );
 a52543a <=( A233  and  (not A232) );
 a52544a <=( a52543a  and  a52540a );
 a52545a <=( a52544a  and  a52537a );
 a52548a <=( (not A235)  and  (not A234) );
 a52551a <=( (not A298)  and  (not A236) );
 a52552a <=( a52551a  and  a52548a );
 a52555a <=( (not A300)  and  A299 );
 a52558a <=( (not A302)  and  (not A301) );
 a52559a <=( a52558a  and  a52555a );
 a52560a <=( a52559a  and  a52552a );
 a52563a <=( A168  and  A169 );
 a52566a <=( A166  and  (not A167) );
 a52567a <=( a52566a  and  a52563a );
 a52570a <=( A200  and  A199 );
 a52573a <=( A233  and  (not A232) );
 a52574a <=( a52573a  and  a52570a );
 a52575a <=( a52574a  and  a52567a );
 a52578a <=( (not A235)  and  (not A234) );
 a52581a <=( (not A265)  and  (not A236) );
 a52582a <=( a52581a  and  a52578a );
 a52585a <=( (not A267)  and  A266 );
 a52588a <=( (not A269)  and  (not A268) );
 a52589a <=( a52588a  and  a52585a );
 a52590a <=( a52589a  and  a52582a );
 a52593a <=( A168  and  A169 );
 a52596a <=( A166  and  (not A167) );
 a52597a <=( a52596a  and  a52593a );
 a52600a <=( A200  and  A199 );
 a52603a <=( A233  and  (not A232) );
 a52604a <=( a52603a  and  a52600a );
 a52605a <=( a52604a  and  a52597a );
 a52608a <=( (not A235)  and  (not A234) );
 a52611a <=( A265  and  (not A236) );
 a52612a <=( a52611a  and  a52608a );
 a52615a <=( (not A267)  and  (not A266) );
 a52618a <=( (not A269)  and  (not A268) );
 a52619a <=( a52618a  and  a52615a );
 a52620a <=( a52619a  and  a52612a );
 a52623a <=( A168  and  A169 );
 a52626a <=( A166  and  (not A167) );
 a52627a <=( a52626a  and  a52623a );
 a52630a <=( A200  and  A199 );
 a52633a <=( (not A233)  and  A232 );
 a52634a <=( a52633a  and  a52630a );
 a52635a <=( a52634a  and  a52627a );
 a52638a <=( (not A235)  and  (not A234) );
 a52641a <=( A298  and  (not A236) );
 a52642a <=( a52641a  and  a52638a );
 a52645a <=( (not A300)  and  (not A299) );
 a52648a <=( (not A302)  and  (not A301) );
 a52649a <=( a52648a  and  a52645a );
 a52650a <=( a52649a  and  a52642a );
 a52653a <=( A168  and  A169 );
 a52656a <=( A166  and  (not A167) );
 a52657a <=( a52656a  and  a52653a );
 a52660a <=( A200  and  A199 );
 a52663a <=( (not A233)  and  A232 );
 a52664a <=( a52663a  and  a52660a );
 a52665a <=( a52664a  and  a52657a );
 a52668a <=( (not A235)  and  (not A234) );
 a52671a <=( (not A298)  and  (not A236) );
 a52672a <=( a52671a  and  a52668a );
 a52675a <=( (not A300)  and  A299 );
 a52678a <=( (not A302)  and  (not A301) );
 a52679a <=( a52678a  and  a52675a );
 a52680a <=( a52679a  and  a52672a );
 a52683a <=( A168  and  A169 );
 a52686a <=( A166  and  (not A167) );
 a52687a <=( a52686a  and  a52683a );
 a52690a <=( A200  and  A199 );
 a52693a <=( (not A233)  and  A232 );
 a52694a <=( a52693a  and  a52690a );
 a52695a <=( a52694a  and  a52687a );
 a52698a <=( (not A235)  and  (not A234) );
 a52701a <=( (not A265)  and  (not A236) );
 a52702a <=( a52701a  and  a52698a );
 a52705a <=( (not A267)  and  A266 );
 a52708a <=( (not A269)  and  (not A268) );
 a52709a <=( a52708a  and  a52705a );
 a52710a <=( a52709a  and  a52702a );
 a52713a <=( A168  and  A169 );
 a52716a <=( A166  and  (not A167) );
 a52717a <=( a52716a  and  a52713a );
 a52720a <=( A200  and  A199 );
 a52723a <=( (not A233)  and  A232 );
 a52724a <=( a52723a  and  a52720a );
 a52725a <=( a52724a  and  a52717a );
 a52728a <=( (not A235)  and  (not A234) );
 a52731a <=( A265  and  (not A236) );
 a52732a <=( a52731a  and  a52728a );
 a52735a <=( (not A267)  and  (not A266) );
 a52738a <=( (not A269)  and  (not A268) );
 a52739a <=( a52738a  and  a52735a );
 a52740a <=( a52739a  and  a52732a );
 a52743a <=( A168  and  A169 );
 a52746a <=( A166  and  (not A167) );
 a52747a <=( a52746a  and  a52743a );
 a52750a <=( (not A200)  and  (not A199) );
 a52753a <=( A233  and  (not A232) );
 a52754a <=( a52753a  and  a52750a );
 a52755a <=( a52754a  and  a52747a );
 a52758a <=( (not A235)  and  (not A234) );
 a52761a <=( A298  and  (not A236) );
 a52762a <=( a52761a  and  a52758a );
 a52765a <=( (not A300)  and  (not A299) );
 a52768a <=( (not A302)  and  (not A301) );
 a52769a <=( a52768a  and  a52765a );
 a52770a <=( a52769a  and  a52762a );
 a52773a <=( A168  and  A169 );
 a52776a <=( A166  and  (not A167) );
 a52777a <=( a52776a  and  a52773a );
 a52780a <=( (not A200)  and  (not A199) );
 a52783a <=( A233  and  (not A232) );
 a52784a <=( a52783a  and  a52780a );
 a52785a <=( a52784a  and  a52777a );
 a52788a <=( (not A235)  and  (not A234) );
 a52791a <=( (not A298)  and  (not A236) );
 a52792a <=( a52791a  and  a52788a );
 a52795a <=( (not A300)  and  A299 );
 a52798a <=( (not A302)  and  (not A301) );
 a52799a <=( a52798a  and  a52795a );
 a52800a <=( a52799a  and  a52792a );
 a52803a <=( A168  and  A169 );
 a52806a <=( A166  and  (not A167) );
 a52807a <=( a52806a  and  a52803a );
 a52810a <=( (not A200)  and  (not A199) );
 a52813a <=( A233  and  (not A232) );
 a52814a <=( a52813a  and  a52810a );
 a52815a <=( a52814a  and  a52807a );
 a52818a <=( (not A235)  and  (not A234) );
 a52821a <=( (not A265)  and  (not A236) );
 a52822a <=( a52821a  and  a52818a );
 a52825a <=( (not A267)  and  A266 );
 a52828a <=( (not A269)  and  (not A268) );
 a52829a <=( a52828a  and  a52825a );
 a52830a <=( a52829a  and  a52822a );
 a52833a <=( A168  and  A169 );
 a52836a <=( A166  and  (not A167) );
 a52837a <=( a52836a  and  a52833a );
 a52840a <=( (not A200)  and  (not A199) );
 a52843a <=( A233  and  (not A232) );
 a52844a <=( a52843a  and  a52840a );
 a52845a <=( a52844a  and  a52837a );
 a52848a <=( (not A235)  and  (not A234) );
 a52851a <=( A265  and  (not A236) );
 a52852a <=( a52851a  and  a52848a );
 a52855a <=( (not A267)  and  (not A266) );
 a52858a <=( (not A269)  and  (not A268) );
 a52859a <=( a52858a  and  a52855a );
 a52860a <=( a52859a  and  a52852a );
 a52863a <=( A168  and  A169 );
 a52866a <=( A166  and  (not A167) );
 a52867a <=( a52866a  and  a52863a );
 a52870a <=( (not A200)  and  (not A199) );
 a52873a <=( (not A233)  and  A232 );
 a52874a <=( a52873a  and  a52870a );
 a52875a <=( a52874a  and  a52867a );
 a52878a <=( (not A235)  and  (not A234) );
 a52881a <=( A298  and  (not A236) );
 a52882a <=( a52881a  and  a52878a );
 a52885a <=( (not A300)  and  (not A299) );
 a52888a <=( (not A302)  and  (not A301) );
 a52889a <=( a52888a  and  a52885a );
 a52890a <=( a52889a  and  a52882a );
 a52893a <=( A168  and  A169 );
 a52896a <=( A166  and  (not A167) );
 a52897a <=( a52896a  and  a52893a );
 a52900a <=( (not A200)  and  (not A199) );
 a52903a <=( (not A233)  and  A232 );
 a52904a <=( a52903a  and  a52900a );
 a52905a <=( a52904a  and  a52897a );
 a52908a <=( (not A235)  and  (not A234) );
 a52911a <=( (not A298)  and  (not A236) );
 a52912a <=( a52911a  and  a52908a );
 a52915a <=( (not A300)  and  A299 );
 a52918a <=( (not A302)  and  (not A301) );
 a52919a <=( a52918a  and  a52915a );
 a52920a <=( a52919a  and  a52912a );
 a52923a <=( A168  and  A169 );
 a52926a <=( A166  and  (not A167) );
 a52927a <=( a52926a  and  a52923a );
 a52930a <=( (not A200)  and  (not A199) );
 a52933a <=( (not A233)  and  A232 );
 a52934a <=( a52933a  and  a52930a );
 a52935a <=( a52934a  and  a52927a );
 a52938a <=( (not A235)  and  (not A234) );
 a52941a <=( (not A265)  and  (not A236) );
 a52942a <=( a52941a  and  a52938a );
 a52945a <=( (not A267)  and  A266 );
 a52948a <=( (not A269)  and  (not A268) );
 a52949a <=( a52948a  and  a52945a );
 a52950a <=( a52949a  and  a52942a );
 a52953a <=( A168  and  A169 );
 a52956a <=( A166  and  (not A167) );
 a52957a <=( a52956a  and  a52953a );
 a52960a <=( (not A200)  and  (not A199) );
 a52963a <=( (not A233)  and  A232 );
 a52964a <=( a52963a  and  a52960a );
 a52965a <=( a52964a  and  a52957a );
 a52968a <=( (not A235)  and  (not A234) );
 a52971a <=( A265  and  (not A236) );
 a52972a <=( a52971a  and  a52968a );
 a52975a <=( (not A267)  and  (not A266) );
 a52978a <=( (not A269)  and  (not A268) );
 a52979a <=( a52978a  and  a52975a );
 a52980a <=( a52979a  and  a52972a );
 a52983a <=( (not A169)  and  A170 );
 a52986a <=( A167  and  (not A168) );
 a52987a <=( a52986a  and  a52983a );
 a52990a <=( A201  and  (not A166) );
 a52993a <=( (not A203)  and  (not A202) );
 a52994a <=( a52993a  and  a52990a );
 a52995a <=( a52994a  and  a52987a );
 a52998a <=( A233  and  (not A232) );
 a53001a <=( A235  and  A234 );
 a53002a <=( a53001a  and  a52998a );
 a53005a <=( (not A299)  and  A298 );
 a53008a <=( A301  and  A300 );
 a53009a <=( a53008a  and  a53005a );
 a53010a <=( a53009a  and  a53002a );
 a53013a <=( (not A169)  and  A170 );
 a53016a <=( A167  and  (not A168) );
 a53017a <=( a53016a  and  a53013a );
 a53020a <=( A201  and  (not A166) );
 a53023a <=( (not A203)  and  (not A202) );
 a53024a <=( a53023a  and  a53020a );
 a53025a <=( a53024a  and  a53017a );
 a53028a <=( A233  and  (not A232) );
 a53031a <=( A235  and  A234 );
 a53032a <=( a53031a  and  a53028a );
 a53035a <=( (not A299)  and  A298 );
 a53038a <=( A302  and  A300 );
 a53039a <=( a53038a  and  a53035a );
 a53040a <=( a53039a  and  a53032a );
 a53043a <=( (not A169)  and  A170 );
 a53046a <=( A167  and  (not A168) );
 a53047a <=( a53046a  and  a53043a );
 a53050a <=( A201  and  (not A166) );
 a53053a <=( (not A203)  and  (not A202) );
 a53054a <=( a53053a  and  a53050a );
 a53055a <=( a53054a  and  a53047a );
 a53058a <=( A233  and  (not A232) );
 a53061a <=( A235  and  A234 );
 a53062a <=( a53061a  and  a53058a );
 a53065a <=( A299  and  (not A298) );
 a53068a <=( A301  and  A300 );
 a53069a <=( a53068a  and  a53065a );
 a53070a <=( a53069a  and  a53062a );
 a53073a <=( (not A169)  and  A170 );
 a53076a <=( A167  and  (not A168) );
 a53077a <=( a53076a  and  a53073a );
 a53080a <=( A201  and  (not A166) );
 a53083a <=( (not A203)  and  (not A202) );
 a53084a <=( a53083a  and  a53080a );
 a53085a <=( a53084a  and  a53077a );
 a53088a <=( A233  and  (not A232) );
 a53091a <=( A235  and  A234 );
 a53092a <=( a53091a  and  a53088a );
 a53095a <=( A299  and  (not A298) );
 a53098a <=( A302  and  A300 );
 a53099a <=( a53098a  and  a53095a );
 a53100a <=( a53099a  and  a53092a );
 a53103a <=( (not A169)  and  A170 );
 a53106a <=( A167  and  (not A168) );
 a53107a <=( a53106a  and  a53103a );
 a53110a <=( A201  and  (not A166) );
 a53113a <=( (not A203)  and  (not A202) );
 a53114a <=( a53113a  and  a53110a );
 a53115a <=( a53114a  and  a53107a );
 a53118a <=( A233  and  (not A232) );
 a53121a <=( A235  and  A234 );
 a53122a <=( a53121a  and  a53118a );
 a53125a <=( A266  and  (not A265) );
 a53128a <=( A268  and  A267 );
 a53129a <=( a53128a  and  a53125a );
 a53130a <=( a53129a  and  a53122a );
 a53133a <=( (not A169)  and  A170 );
 a53136a <=( A167  and  (not A168) );
 a53137a <=( a53136a  and  a53133a );
 a53140a <=( A201  and  (not A166) );
 a53143a <=( (not A203)  and  (not A202) );
 a53144a <=( a53143a  and  a53140a );
 a53145a <=( a53144a  and  a53137a );
 a53148a <=( A233  and  (not A232) );
 a53151a <=( A235  and  A234 );
 a53152a <=( a53151a  and  a53148a );
 a53155a <=( A266  and  (not A265) );
 a53158a <=( A269  and  A267 );
 a53159a <=( a53158a  and  a53155a );
 a53160a <=( a53159a  and  a53152a );
 a53163a <=( (not A169)  and  A170 );
 a53166a <=( A167  and  (not A168) );
 a53167a <=( a53166a  and  a53163a );
 a53170a <=( A201  and  (not A166) );
 a53173a <=( (not A203)  and  (not A202) );
 a53174a <=( a53173a  and  a53170a );
 a53175a <=( a53174a  and  a53167a );
 a53178a <=( A233  and  (not A232) );
 a53181a <=( A235  and  A234 );
 a53182a <=( a53181a  and  a53178a );
 a53185a <=( (not A266)  and  A265 );
 a53188a <=( A268  and  A267 );
 a53189a <=( a53188a  and  a53185a );
 a53190a <=( a53189a  and  a53182a );
 a53193a <=( (not A169)  and  A170 );
 a53196a <=( A167  and  (not A168) );
 a53197a <=( a53196a  and  a53193a );
 a53200a <=( A201  and  (not A166) );
 a53203a <=( (not A203)  and  (not A202) );
 a53204a <=( a53203a  and  a53200a );
 a53205a <=( a53204a  and  a53197a );
 a53208a <=( A233  and  (not A232) );
 a53211a <=( A235  and  A234 );
 a53212a <=( a53211a  and  a53208a );
 a53215a <=( (not A266)  and  A265 );
 a53218a <=( A269  and  A267 );
 a53219a <=( a53218a  and  a53215a );
 a53220a <=( a53219a  and  a53212a );
 a53223a <=( (not A169)  and  A170 );
 a53226a <=( A167  and  (not A168) );
 a53227a <=( a53226a  and  a53223a );
 a53230a <=( A201  and  (not A166) );
 a53233a <=( (not A203)  and  (not A202) );
 a53234a <=( a53233a  and  a53230a );
 a53235a <=( a53234a  and  a53227a );
 a53238a <=( A233  and  (not A232) );
 a53241a <=( A236  and  A234 );
 a53242a <=( a53241a  and  a53238a );
 a53245a <=( (not A299)  and  A298 );
 a53248a <=( A301  and  A300 );
 a53249a <=( a53248a  and  a53245a );
 a53250a <=( a53249a  and  a53242a );
 a53253a <=( (not A169)  and  A170 );
 a53256a <=( A167  and  (not A168) );
 a53257a <=( a53256a  and  a53253a );
 a53260a <=( A201  and  (not A166) );
 a53263a <=( (not A203)  and  (not A202) );
 a53264a <=( a53263a  and  a53260a );
 a53265a <=( a53264a  and  a53257a );
 a53268a <=( A233  and  (not A232) );
 a53271a <=( A236  and  A234 );
 a53272a <=( a53271a  and  a53268a );
 a53275a <=( (not A299)  and  A298 );
 a53278a <=( A302  and  A300 );
 a53279a <=( a53278a  and  a53275a );
 a53280a <=( a53279a  and  a53272a );
 a53283a <=( (not A169)  and  A170 );
 a53286a <=( A167  and  (not A168) );
 a53287a <=( a53286a  and  a53283a );
 a53290a <=( A201  and  (not A166) );
 a53293a <=( (not A203)  and  (not A202) );
 a53294a <=( a53293a  and  a53290a );
 a53295a <=( a53294a  and  a53287a );
 a53298a <=( A233  and  (not A232) );
 a53301a <=( A236  and  A234 );
 a53302a <=( a53301a  and  a53298a );
 a53305a <=( A299  and  (not A298) );
 a53308a <=( A301  and  A300 );
 a53309a <=( a53308a  and  a53305a );
 a53310a <=( a53309a  and  a53302a );
 a53313a <=( (not A169)  and  A170 );
 a53316a <=( A167  and  (not A168) );
 a53317a <=( a53316a  and  a53313a );
 a53320a <=( A201  and  (not A166) );
 a53323a <=( (not A203)  and  (not A202) );
 a53324a <=( a53323a  and  a53320a );
 a53325a <=( a53324a  and  a53317a );
 a53328a <=( A233  and  (not A232) );
 a53331a <=( A236  and  A234 );
 a53332a <=( a53331a  and  a53328a );
 a53335a <=( A299  and  (not A298) );
 a53338a <=( A302  and  A300 );
 a53339a <=( a53338a  and  a53335a );
 a53340a <=( a53339a  and  a53332a );
 a53343a <=( (not A169)  and  A170 );
 a53346a <=( A167  and  (not A168) );
 a53347a <=( a53346a  and  a53343a );
 a53350a <=( A201  and  (not A166) );
 a53353a <=( (not A203)  and  (not A202) );
 a53354a <=( a53353a  and  a53350a );
 a53355a <=( a53354a  and  a53347a );
 a53358a <=( A233  and  (not A232) );
 a53361a <=( A236  and  A234 );
 a53362a <=( a53361a  and  a53358a );
 a53365a <=( A266  and  (not A265) );
 a53368a <=( A268  and  A267 );
 a53369a <=( a53368a  and  a53365a );
 a53370a <=( a53369a  and  a53362a );
 a53373a <=( (not A169)  and  A170 );
 a53376a <=( A167  and  (not A168) );
 a53377a <=( a53376a  and  a53373a );
 a53380a <=( A201  and  (not A166) );
 a53383a <=( (not A203)  and  (not A202) );
 a53384a <=( a53383a  and  a53380a );
 a53385a <=( a53384a  and  a53377a );
 a53388a <=( A233  and  (not A232) );
 a53391a <=( A236  and  A234 );
 a53392a <=( a53391a  and  a53388a );
 a53395a <=( A266  and  (not A265) );
 a53398a <=( A269  and  A267 );
 a53399a <=( a53398a  and  a53395a );
 a53400a <=( a53399a  and  a53392a );
 a53403a <=( (not A169)  and  A170 );
 a53406a <=( A167  and  (not A168) );
 a53407a <=( a53406a  and  a53403a );
 a53410a <=( A201  and  (not A166) );
 a53413a <=( (not A203)  and  (not A202) );
 a53414a <=( a53413a  and  a53410a );
 a53415a <=( a53414a  and  a53407a );
 a53418a <=( A233  and  (not A232) );
 a53421a <=( A236  and  A234 );
 a53422a <=( a53421a  and  a53418a );
 a53425a <=( (not A266)  and  A265 );
 a53428a <=( A268  and  A267 );
 a53429a <=( a53428a  and  a53425a );
 a53430a <=( a53429a  and  a53422a );
 a53433a <=( (not A169)  and  A170 );
 a53436a <=( A167  and  (not A168) );
 a53437a <=( a53436a  and  a53433a );
 a53440a <=( A201  and  (not A166) );
 a53443a <=( (not A203)  and  (not A202) );
 a53444a <=( a53443a  and  a53440a );
 a53445a <=( a53444a  and  a53437a );
 a53448a <=( A233  and  (not A232) );
 a53451a <=( A236  and  A234 );
 a53452a <=( a53451a  and  a53448a );
 a53455a <=( (not A266)  and  A265 );
 a53458a <=( A269  and  A267 );
 a53459a <=( a53458a  and  a53455a );
 a53460a <=( a53459a  and  a53452a );
 a53463a <=( (not A169)  and  A170 );
 a53466a <=( A167  and  (not A168) );
 a53467a <=( a53466a  and  a53463a );
 a53470a <=( A201  and  (not A166) );
 a53473a <=( (not A203)  and  (not A202) );
 a53474a <=( a53473a  and  a53470a );
 a53475a <=( a53474a  and  a53467a );
 a53478a <=( (not A233)  and  A232 );
 a53481a <=( A235  and  A234 );
 a53482a <=( a53481a  and  a53478a );
 a53485a <=( (not A299)  and  A298 );
 a53488a <=( A301  and  A300 );
 a53489a <=( a53488a  and  a53485a );
 a53490a <=( a53489a  and  a53482a );
 a53493a <=( (not A169)  and  A170 );
 a53496a <=( A167  and  (not A168) );
 a53497a <=( a53496a  and  a53493a );
 a53500a <=( A201  and  (not A166) );
 a53503a <=( (not A203)  and  (not A202) );
 a53504a <=( a53503a  and  a53500a );
 a53505a <=( a53504a  and  a53497a );
 a53508a <=( (not A233)  and  A232 );
 a53511a <=( A235  and  A234 );
 a53512a <=( a53511a  and  a53508a );
 a53515a <=( (not A299)  and  A298 );
 a53518a <=( A302  and  A300 );
 a53519a <=( a53518a  and  a53515a );
 a53520a <=( a53519a  and  a53512a );
 a53523a <=( (not A169)  and  A170 );
 a53526a <=( A167  and  (not A168) );
 a53527a <=( a53526a  and  a53523a );
 a53530a <=( A201  and  (not A166) );
 a53533a <=( (not A203)  and  (not A202) );
 a53534a <=( a53533a  and  a53530a );
 a53535a <=( a53534a  and  a53527a );
 a53538a <=( (not A233)  and  A232 );
 a53541a <=( A235  and  A234 );
 a53542a <=( a53541a  and  a53538a );
 a53545a <=( A299  and  (not A298) );
 a53548a <=( A301  and  A300 );
 a53549a <=( a53548a  and  a53545a );
 a53550a <=( a53549a  and  a53542a );
 a53553a <=( (not A169)  and  A170 );
 a53556a <=( A167  and  (not A168) );
 a53557a <=( a53556a  and  a53553a );
 a53560a <=( A201  and  (not A166) );
 a53563a <=( (not A203)  and  (not A202) );
 a53564a <=( a53563a  and  a53560a );
 a53565a <=( a53564a  and  a53557a );
 a53568a <=( (not A233)  and  A232 );
 a53571a <=( A235  and  A234 );
 a53572a <=( a53571a  and  a53568a );
 a53575a <=( A299  and  (not A298) );
 a53578a <=( A302  and  A300 );
 a53579a <=( a53578a  and  a53575a );
 a53580a <=( a53579a  and  a53572a );
 a53583a <=( (not A169)  and  A170 );
 a53586a <=( A167  and  (not A168) );
 a53587a <=( a53586a  and  a53583a );
 a53590a <=( A201  and  (not A166) );
 a53593a <=( (not A203)  and  (not A202) );
 a53594a <=( a53593a  and  a53590a );
 a53595a <=( a53594a  and  a53587a );
 a53598a <=( (not A233)  and  A232 );
 a53601a <=( A235  and  A234 );
 a53602a <=( a53601a  and  a53598a );
 a53605a <=( A266  and  (not A265) );
 a53608a <=( A268  and  A267 );
 a53609a <=( a53608a  and  a53605a );
 a53610a <=( a53609a  and  a53602a );
 a53613a <=( (not A169)  and  A170 );
 a53616a <=( A167  and  (not A168) );
 a53617a <=( a53616a  and  a53613a );
 a53620a <=( A201  and  (not A166) );
 a53623a <=( (not A203)  and  (not A202) );
 a53624a <=( a53623a  and  a53620a );
 a53625a <=( a53624a  and  a53617a );
 a53628a <=( (not A233)  and  A232 );
 a53631a <=( A235  and  A234 );
 a53632a <=( a53631a  and  a53628a );
 a53635a <=( A266  and  (not A265) );
 a53638a <=( A269  and  A267 );
 a53639a <=( a53638a  and  a53635a );
 a53640a <=( a53639a  and  a53632a );
 a53643a <=( (not A169)  and  A170 );
 a53646a <=( A167  and  (not A168) );
 a53647a <=( a53646a  and  a53643a );
 a53650a <=( A201  and  (not A166) );
 a53653a <=( (not A203)  and  (not A202) );
 a53654a <=( a53653a  and  a53650a );
 a53655a <=( a53654a  and  a53647a );
 a53658a <=( (not A233)  and  A232 );
 a53661a <=( A235  and  A234 );
 a53662a <=( a53661a  and  a53658a );
 a53665a <=( (not A266)  and  A265 );
 a53668a <=( A268  and  A267 );
 a53669a <=( a53668a  and  a53665a );
 a53670a <=( a53669a  and  a53662a );
 a53673a <=( (not A169)  and  A170 );
 a53676a <=( A167  and  (not A168) );
 a53677a <=( a53676a  and  a53673a );
 a53680a <=( A201  and  (not A166) );
 a53683a <=( (not A203)  and  (not A202) );
 a53684a <=( a53683a  and  a53680a );
 a53685a <=( a53684a  and  a53677a );
 a53688a <=( (not A233)  and  A232 );
 a53691a <=( A235  and  A234 );
 a53692a <=( a53691a  and  a53688a );
 a53695a <=( (not A266)  and  A265 );
 a53698a <=( A269  and  A267 );
 a53699a <=( a53698a  and  a53695a );
 a53700a <=( a53699a  and  a53692a );
 a53703a <=( (not A169)  and  A170 );
 a53706a <=( A167  and  (not A168) );
 a53707a <=( a53706a  and  a53703a );
 a53710a <=( A201  and  (not A166) );
 a53713a <=( (not A203)  and  (not A202) );
 a53714a <=( a53713a  and  a53710a );
 a53715a <=( a53714a  and  a53707a );
 a53718a <=( (not A233)  and  A232 );
 a53721a <=( A236  and  A234 );
 a53722a <=( a53721a  and  a53718a );
 a53725a <=( (not A299)  and  A298 );
 a53728a <=( A301  and  A300 );
 a53729a <=( a53728a  and  a53725a );
 a53730a <=( a53729a  and  a53722a );
 a53733a <=( (not A169)  and  A170 );
 a53736a <=( A167  and  (not A168) );
 a53737a <=( a53736a  and  a53733a );
 a53740a <=( A201  and  (not A166) );
 a53743a <=( (not A203)  and  (not A202) );
 a53744a <=( a53743a  and  a53740a );
 a53745a <=( a53744a  and  a53737a );
 a53748a <=( (not A233)  and  A232 );
 a53751a <=( A236  and  A234 );
 a53752a <=( a53751a  and  a53748a );
 a53755a <=( (not A299)  and  A298 );
 a53758a <=( A302  and  A300 );
 a53759a <=( a53758a  and  a53755a );
 a53760a <=( a53759a  and  a53752a );
 a53763a <=( (not A169)  and  A170 );
 a53766a <=( A167  and  (not A168) );
 a53767a <=( a53766a  and  a53763a );
 a53770a <=( A201  and  (not A166) );
 a53773a <=( (not A203)  and  (not A202) );
 a53774a <=( a53773a  and  a53770a );
 a53775a <=( a53774a  and  a53767a );
 a53778a <=( (not A233)  and  A232 );
 a53781a <=( A236  and  A234 );
 a53782a <=( a53781a  and  a53778a );
 a53785a <=( A299  and  (not A298) );
 a53788a <=( A301  and  A300 );
 a53789a <=( a53788a  and  a53785a );
 a53790a <=( a53789a  and  a53782a );
 a53793a <=( (not A169)  and  A170 );
 a53796a <=( A167  and  (not A168) );
 a53797a <=( a53796a  and  a53793a );
 a53800a <=( A201  and  (not A166) );
 a53803a <=( (not A203)  and  (not A202) );
 a53804a <=( a53803a  and  a53800a );
 a53805a <=( a53804a  and  a53797a );
 a53808a <=( (not A233)  and  A232 );
 a53811a <=( A236  and  A234 );
 a53812a <=( a53811a  and  a53808a );
 a53815a <=( A299  and  (not A298) );
 a53818a <=( A302  and  A300 );
 a53819a <=( a53818a  and  a53815a );
 a53820a <=( a53819a  and  a53812a );
 a53823a <=( (not A169)  and  A170 );
 a53826a <=( A167  and  (not A168) );
 a53827a <=( a53826a  and  a53823a );
 a53830a <=( A201  and  (not A166) );
 a53833a <=( (not A203)  and  (not A202) );
 a53834a <=( a53833a  and  a53830a );
 a53835a <=( a53834a  and  a53827a );
 a53838a <=( (not A233)  and  A232 );
 a53841a <=( A236  and  A234 );
 a53842a <=( a53841a  and  a53838a );
 a53845a <=( A266  and  (not A265) );
 a53848a <=( A268  and  A267 );
 a53849a <=( a53848a  and  a53845a );
 a53850a <=( a53849a  and  a53842a );
 a53853a <=( (not A169)  and  A170 );
 a53856a <=( A167  and  (not A168) );
 a53857a <=( a53856a  and  a53853a );
 a53860a <=( A201  and  (not A166) );
 a53863a <=( (not A203)  and  (not A202) );
 a53864a <=( a53863a  and  a53860a );
 a53865a <=( a53864a  and  a53857a );
 a53868a <=( (not A233)  and  A232 );
 a53871a <=( A236  and  A234 );
 a53872a <=( a53871a  and  a53868a );
 a53875a <=( A266  and  (not A265) );
 a53878a <=( A269  and  A267 );
 a53879a <=( a53878a  and  a53875a );
 a53880a <=( a53879a  and  a53872a );
 a53883a <=( (not A169)  and  A170 );
 a53886a <=( A167  and  (not A168) );
 a53887a <=( a53886a  and  a53883a );
 a53890a <=( A201  and  (not A166) );
 a53893a <=( (not A203)  and  (not A202) );
 a53894a <=( a53893a  and  a53890a );
 a53895a <=( a53894a  and  a53887a );
 a53898a <=( (not A233)  and  A232 );
 a53901a <=( A236  and  A234 );
 a53902a <=( a53901a  and  a53898a );
 a53905a <=( (not A266)  and  A265 );
 a53908a <=( A268  and  A267 );
 a53909a <=( a53908a  and  a53905a );
 a53910a <=( a53909a  and  a53902a );
 a53913a <=( (not A169)  and  A170 );
 a53916a <=( A167  and  (not A168) );
 a53917a <=( a53916a  and  a53913a );
 a53920a <=( A201  and  (not A166) );
 a53923a <=( (not A203)  and  (not A202) );
 a53924a <=( a53923a  and  a53920a );
 a53925a <=( a53924a  and  a53917a );
 a53928a <=( (not A233)  and  A232 );
 a53931a <=( A236  and  A234 );
 a53932a <=( a53931a  and  a53928a );
 a53935a <=( (not A266)  and  A265 );
 a53938a <=( A269  and  A267 );
 a53939a <=( a53938a  and  a53935a );
 a53940a <=( a53939a  and  a53932a );
 a53943a <=( (not A169)  and  A170 );
 a53946a <=( A167  and  (not A168) );
 a53947a <=( a53946a  and  a53943a );
 a53950a <=( (not A201)  and  (not A166) );
 a53953a <=( (not A232)  and  A202 );
 a53954a <=( a53953a  and  a53950a );
 a53955a <=( a53954a  and  a53947a );
 a53958a <=( A234  and  A233 );
 a53961a <=( A298  and  A235 );
 a53962a <=( a53961a  and  a53958a );
 a53965a <=( (not A300)  and  (not A299) );
 a53968a <=( (not A302)  and  (not A301) );
 a53969a <=( a53968a  and  a53965a );
 a53970a <=( a53969a  and  a53962a );
 a53973a <=( (not A169)  and  A170 );
 a53976a <=( A167  and  (not A168) );
 a53977a <=( a53976a  and  a53973a );
 a53980a <=( (not A201)  and  (not A166) );
 a53983a <=( (not A232)  and  A202 );
 a53984a <=( a53983a  and  a53980a );
 a53985a <=( a53984a  and  a53977a );
 a53988a <=( A234  and  A233 );
 a53991a <=( (not A298)  and  A235 );
 a53992a <=( a53991a  and  a53988a );
 a53995a <=( (not A300)  and  A299 );
 a53998a <=( (not A302)  and  (not A301) );
 a53999a <=( a53998a  and  a53995a );
 a54000a <=( a53999a  and  a53992a );
 a54003a <=( (not A169)  and  A170 );
 a54006a <=( A167  and  (not A168) );
 a54007a <=( a54006a  and  a54003a );
 a54010a <=( (not A201)  and  (not A166) );
 a54013a <=( (not A232)  and  A202 );
 a54014a <=( a54013a  and  a54010a );
 a54015a <=( a54014a  and  a54007a );
 a54018a <=( A234  and  A233 );
 a54021a <=( (not A265)  and  A235 );
 a54022a <=( a54021a  and  a54018a );
 a54025a <=( (not A267)  and  A266 );
 a54028a <=( (not A269)  and  (not A268) );
 a54029a <=( a54028a  and  a54025a );
 a54030a <=( a54029a  and  a54022a );
 a54033a <=( (not A169)  and  A170 );
 a54036a <=( A167  and  (not A168) );
 a54037a <=( a54036a  and  a54033a );
 a54040a <=( (not A201)  and  (not A166) );
 a54043a <=( (not A232)  and  A202 );
 a54044a <=( a54043a  and  a54040a );
 a54045a <=( a54044a  and  a54037a );
 a54048a <=( A234  and  A233 );
 a54051a <=( A265  and  A235 );
 a54052a <=( a54051a  and  a54048a );
 a54055a <=( (not A267)  and  (not A266) );
 a54058a <=( (not A269)  and  (not A268) );
 a54059a <=( a54058a  and  a54055a );
 a54060a <=( a54059a  and  a54052a );
 a54063a <=( (not A169)  and  A170 );
 a54066a <=( A167  and  (not A168) );
 a54067a <=( a54066a  and  a54063a );
 a54070a <=( (not A201)  and  (not A166) );
 a54073a <=( (not A232)  and  A202 );
 a54074a <=( a54073a  and  a54070a );
 a54075a <=( a54074a  and  a54067a );
 a54078a <=( A234  and  A233 );
 a54081a <=( A298  and  A236 );
 a54082a <=( a54081a  and  a54078a );
 a54085a <=( (not A300)  and  (not A299) );
 a54088a <=( (not A302)  and  (not A301) );
 a54089a <=( a54088a  and  a54085a );
 a54090a <=( a54089a  and  a54082a );
 a54093a <=( (not A169)  and  A170 );
 a54096a <=( A167  and  (not A168) );
 a54097a <=( a54096a  and  a54093a );
 a54100a <=( (not A201)  and  (not A166) );
 a54103a <=( (not A232)  and  A202 );
 a54104a <=( a54103a  and  a54100a );
 a54105a <=( a54104a  and  a54097a );
 a54108a <=( A234  and  A233 );
 a54111a <=( (not A298)  and  A236 );
 a54112a <=( a54111a  and  a54108a );
 a54115a <=( (not A300)  and  A299 );
 a54118a <=( (not A302)  and  (not A301) );
 a54119a <=( a54118a  and  a54115a );
 a54120a <=( a54119a  and  a54112a );
 a54123a <=( (not A169)  and  A170 );
 a54126a <=( A167  and  (not A168) );
 a54127a <=( a54126a  and  a54123a );
 a54130a <=( (not A201)  and  (not A166) );
 a54133a <=( (not A232)  and  A202 );
 a54134a <=( a54133a  and  a54130a );
 a54135a <=( a54134a  and  a54127a );
 a54138a <=( A234  and  A233 );
 a54141a <=( (not A265)  and  A236 );
 a54142a <=( a54141a  and  a54138a );
 a54145a <=( (not A267)  and  A266 );
 a54148a <=( (not A269)  and  (not A268) );
 a54149a <=( a54148a  and  a54145a );
 a54150a <=( a54149a  and  a54142a );
 a54153a <=( (not A169)  and  A170 );
 a54156a <=( A167  and  (not A168) );
 a54157a <=( a54156a  and  a54153a );
 a54160a <=( (not A201)  and  (not A166) );
 a54163a <=( (not A232)  and  A202 );
 a54164a <=( a54163a  and  a54160a );
 a54165a <=( a54164a  and  a54157a );
 a54168a <=( A234  and  A233 );
 a54171a <=( A265  and  A236 );
 a54172a <=( a54171a  and  a54168a );
 a54175a <=( (not A267)  and  (not A266) );
 a54178a <=( (not A269)  and  (not A268) );
 a54179a <=( a54178a  and  a54175a );
 a54180a <=( a54179a  and  a54172a );
 a54183a <=( (not A169)  and  A170 );
 a54186a <=( A167  and  (not A168) );
 a54187a <=( a54186a  and  a54183a );
 a54190a <=( (not A201)  and  (not A166) );
 a54193a <=( (not A232)  and  A202 );
 a54194a <=( a54193a  and  a54190a );
 a54195a <=( a54194a  and  a54187a );
 a54198a <=( (not A234)  and  A233 );
 a54201a <=( (not A236)  and  (not A235) );
 a54202a <=( a54201a  and  a54198a );
 a54205a <=( (not A299)  and  A298 );
 a54208a <=( A301  and  A300 );
 a54209a <=( a54208a  and  a54205a );
 a54210a <=( a54209a  and  a54202a );
 a54213a <=( (not A169)  and  A170 );
 a54216a <=( A167  and  (not A168) );
 a54217a <=( a54216a  and  a54213a );
 a54220a <=( (not A201)  and  (not A166) );
 a54223a <=( (not A232)  and  A202 );
 a54224a <=( a54223a  and  a54220a );
 a54225a <=( a54224a  and  a54217a );
 a54228a <=( (not A234)  and  A233 );
 a54231a <=( (not A236)  and  (not A235) );
 a54232a <=( a54231a  and  a54228a );
 a54235a <=( (not A299)  and  A298 );
 a54238a <=( A302  and  A300 );
 a54239a <=( a54238a  and  a54235a );
 a54240a <=( a54239a  and  a54232a );
 a54243a <=( (not A169)  and  A170 );
 a54246a <=( A167  and  (not A168) );
 a54247a <=( a54246a  and  a54243a );
 a54250a <=( (not A201)  and  (not A166) );
 a54253a <=( (not A232)  and  A202 );
 a54254a <=( a54253a  and  a54250a );
 a54255a <=( a54254a  and  a54247a );
 a54258a <=( (not A234)  and  A233 );
 a54261a <=( (not A236)  and  (not A235) );
 a54262a <=( a54261a  and  a54258a );
 a54265a <=( A299  and  (not A298) );
 a54268a <=( A301  and  A300 );
 a54269a <=( a54268a  and  a54265a );
 a54270a <=( a54269a  and  a54262a );
 a54273a <=( (not A169)  and  A170 );
 a54276a <=( A167  and  (not A168) );
 a54277a <=( a54276a  and  a54273a );
 a54280a <=( (not A201)  and  (not A166) );
 a54283a <=( (not A232)  and  A202 );
 a54284a <=( a54283a  and  a54280a );
 a54285a <=( a54284a  and  a54277a );
 a54288a <=( (not A234)  and  A233 );
 a54291a <=( (not A236)  and  (not A235) );
 a54292a <=( a54291a  and  a54288a );
 a54295a <=( A299  and  (not A298) );
 a54298a <=( A302  and  A300 );
 a54299a <=( a54298a  and  a54295a );
 a54300a <=( a54299a  and  a54292a );
 a54303a <=( (not A169)  and  A170 );
 a54306a <=( A167  and  (not A168) );
 a54307a <=( a54306a  and  a54303a );
 a54310a <=( (not A201)  and  (not A166) );
 a54313a <=( (not A232)  and  A202 );
 a54314a <=( a54313a  and  a54310a );
 a54315a <=( a54314a  and  a54307a );
 a54318a <=( (not A234)  and  A233 );
 a54321a <=( (not A236)  and  (not A235) );
 a54322a <=( a54321a  and  a54318a );
 a54325a <=( A266  and  (not A265) );
 a54328a <=( A268  and  A267 );
 a54329a <=( a54328a  and  a54325a );
 a54330a <=( a54329a  and  a54322a );
 a54333a <=( (not A169)  and  A170 );
 a54336a <=( A167  and  (not A168) );
 a54337a <=( a54336a  and  a54333a );
 a54340a <=( (not A201)  and  (not A166) );
 a54343a <=( (not A232)  and  A202 );
 a54344a <=( a54343a  and  a54340a );
 a54345a <=( a54344a  and  a54337a );
 a54348a <=( (not A234)  and  A233 );
 a54351a <=( (not A236)  and  (not A235) );
 a54352a <=( a54351a  and  a54348a );
 a54355a <=( A266  and  (not A265) );
 a54358a <=( A269  and  A267 );
 a54359a <=( a54358a  and  a54355a );
 a54360a <=( a54359a  and  a54352a );
 a54363a <=( (not A169)  and  A170 );
 a54366a <=( A167  and  (not A168) );
 a54367a <=( a54366a  and  a54363a );
 a54370a <=( (not A201)  and  (not A166) );
 a54373a <=( (not A232)  and  A202 );
 a54374a <=( a54373a  and  a54370a );
 a54375a <=( a54374a  and  a54367a );
 a54378a <=( (not A234)  and  A233 );
 a54381a <=( (not A236)  and  (not A235) );
 a54382a <=( a54381a  and  a54378a );
 a54385a <=( (not A266)  and  A265 );
 a54388a <=( A268  and  A267 );
 a54389a <=( a54388a  and  a54385a );
 a54390a <=( a54389a  and  a54382a );
 a54393a <=( (not A169)  and  A170 );
 a54396a <=( A167  and  (not A168) );
 a54397a <=( a54396a  and  a54393a );
 a54400a <=( (not A201)  and  (not A166) );
 a54403a <=( (not A232)  and  A202 );
 a54404a <=( a54403a  and  a54400a );
 a54405a <=( a54404a  and  a54397a );
 a54408a <=( (not A234)  and  A233 );
 a54411a <=( (not A236)  and  (not A235) );
 a54412a <=( a54411a  and  a54408a );
 a54415a <=( (not A266)  and  A265 );
 a54418a <=( A269  and  A267 );
 a54419a <=( a54418a  and  a54415a );
 a54420a <=( a54419a  and  a54412a );
 a54423a <=( (not A169)  and  A170 );
 a54426a <=( A167  and  (not A168) );
 a54427a <=( a54426a  and  a54423a );
 a54430a <=( (not A201)  and  (not A166) );
 a54433a <=( A232  and  A202 );
 a54434a <=( a54433a  and  a54430a );
 a54435a <=( a54434a  and  a54427a );
 a54438a <=( A234  and  (not A233) );
 a54441a <=( A298  and  A235 );
 a54442a <=( a54441a  and  a54438a );
 a54445a <=( (not A300)  and  (not A299) );
 a54448a <=( (not A302)  and  (not A301) );
 a54449a <=( a54448a  and  a54445a );
 a54450a <=( a54449a  and  a54442a );
 a54453a <=( (not A169)  and  A170 );
 a54456a <=( A167  and  (not A168) );
 a54457a <=( a54456a  and  a54453a );
 a54460a <=( (not A201)  and  (not A166) );
 a54463a <=( A232  and  A202 );
 a54464a <=( a54463a  and  a54460a );
 a54465a <=( a54464a  and  a54457a );
 a54468a <=( A234  and  (not A233) );
 a54471a <=( (not A298)  and  A235 );
 a54472a <=( a54471a  and  a54468a );
 a54475a <=( (not A300)  and  A299 );
 a54478a <=( (not A302)  and  (not A301) );
 a54479a <=( a54478a  and  a54475a );
 a54480a <=( a54479a  and  a54472a );
 a54483a <=( (not A169)  and  A170 );
 a54486a <=( A167  and  (not A168) );
 a54487a <=( a54486a  and  a54483a );
 a54490a <=( (not A201)  and  (not A166) );
 a54493a <=( A232  and  A202 );
 a54494a <=( a54493a  and  a54490a );
 a54495a <=( a54494a  and  a54487a );
 a54498a <=( A234  and  (not A233) );
 a54501a <=( (not A265)  and  A235 );
 a54502a <=( a54501a  and  a54498a );
 a54505a <=( (not A267)  and  A266 );
 a54508a <=( (not A269)  and  (not A268) );
 a54509a <=( a54508a  and  a54505a );
 a54510a <=( a54509a  and  a54502a );
 a54513a <=( (not A169)  and  A170 );
 a54516a <=( A167  and  (not A168) );
 a54517a <=( a54516a  and  a54513a );
 a54520a <=( (not A201)  and  (not A166) );
 a54523a <=( A232  and  A202 );
 a54524a <=( a54523a  and  a54520a );
 a54525a <=( a54524a  and  a54517a );
 a54528a <=( A234  and  (not A233) );
 a54531a <=( A265  and  A235 );
 a54532a <=( a54531a  and  a54528a );
 a54535a <=( (not A267)  and  (not A266) );
 a54538a <=( (not A269)  and  (not A268) );
 a54539a <=( a54538a  and  a54535a );
 a54540a <=( a54539a  and  a54532a );
 a54543a <=( (not A169)  and  A170 );
 a54546a <=( A167  and  (not A168) );
 a54547a <=( a54546a  and  a54543a );
 a54550a <=( (not A201)  and  (not A166) );
 a54553a <=( A232  and  A202 );
 a54554a <=( a54553a  and  a54550a );
 a54555a <=( a54554a  and  a54547a );
 a54558a <=( A234  and  (not A233) );
 a54561a <=( A298  and  A236 );
 a54562a <=( a54561a  and  a54558a );
 a54565a <=( (not A300)  and  (not A299) );
 a54568a <=( (not A302)  and  (not A301) );
 a54569a <=( a54568a  and  a54565a );
 a54570a <=( a54569a  and  a54562a );
 a54573a <=( (not A169)  and  A170 );
 a54576a <=( A167  and  (not A168) );
 a54577a <=( a54576a  and  a54573a );
 a54580a <=( (not A201)  and  (not A166) );
 a54583a <=( A232  and  A202 );
 a54584a <=( a54583a  and  a54580a );
 a54585a <=( a54584a  and  a54577a );
 a54588a <=( A234  and  (not A233) );
 a54591a <=( (not A298)  and  A236 );
 a54592a <=( a54591a  and  a54588a );
 a54595a <=( (not A300)  and  A299 );
 a54598a <=( (not A302)  and  (not A301) );
 a54599a <=( a54598a  and  a54595a );
 a54600a <=( a54599a  and  a54592a );
 a54603a <=( (not A169)  and  A170 );
 a54606a <=( A167  and  (not A168) );
 a54607a <=( a54606a  and  a54603a );
 a54610a <=( (not A201)  and  (not A166) );
 a54613a <=( A232  and  A202 );
 a54614a <=( a54613a  and  a54610a );
 a54615a <=( a54614a  and  a54607a );
 a54618a <=( A234  and  (not A233) );
 a54621a <=( (not A265)  and  A236 );
 a54622a <=( a54621a  and  a54618a );
 a54625a <=( (not A267)  and  A266 );
 a54628a <=( (not A269)  and  (not A268) );
 a54629a <=( a54628a  and  a54625a );
 a54630a <=( a54629a  and  a54622a );
 a54633a <=( (not A169)  and  A170 );
 a54636a <=( A167  and  (not A168) );
 a54637a <=( a54636a  and  a54633a );
 a54640a <=( (not A201)  and  (not A166) );
 a54643a <=( A232  and  A202 );
 a54644a <=( a54643a  and  a54640a );
 a54645a <=( a54644a  and  a54637a );
 a54648a <=( A234  and  (not A233) );
 a54651a <=( A265  and  A236 );
 a54652a <=( a54651a  and  a54648a );
 a54655a <=( (not A267)  and  (not A266) );
 a54658a <=( (not A269)  and  (not A268) );
 a54659a <=( a54658a  and  a54655a );
 a54660a <=( a54659a  and  a54652a );
 a54663a <=( (not A169)  and  A170 );
 a54666a <=( A167  and  (not A168) );
 a54667a <=( a54666a  and  a54663a );
 a54670a <=( (not A201)  and  (not A166) );
 a54673a <=( A232  and  A202 );
 a54674a <=( a54673a  and  a54670a );
 a54675a <=( a54674a  and  a54667a );
 a54678a <=( (not A234)  and  (not A233) );
 a54681a <=( (not A236)  and  (not A235) );
 a54682a <=( a54681a  and  a54678a );
 a54685a <=( (not A299)  and  A298 );
 a54688a <=( A301  and  A300 );
 a54689a <=( a54688a  and  a54685a );
 a54690a <=( a54689a  and  a54682a );
 a54693a <=( (not A169)  and  A170 );
 a54696a <=( A167  and  (not A168) );
 a54697a <=( a54696a  and  a54693a );
 a54700a <=( (not A201)  and  (not A166) );
 a54703a <=( A232  and  A202 );
 a54704a <=( a54703a  and  a54700a );
 a54705a <=( a54704a  and  a54697a );
 a54708a <=( (not A234)  and  (not A233) );
 a54711a <=( (not A236)  and  (not A235) );
 a54712a <=( a54711a  and  a54708a );
 a54715a <=( (not A299)  and  A298 );
 a54718a <=( A302  and  A300 );
 a54719a <=( a54718a  and  a54715a );
 a54720a <=( a54719a  and  a54712a );
 a54723a <=( (not A169)  and  A170 );
 a54726a <=( A167  and  (not A168) );
 a54727a <=( a54726a  and  a54723a );
 a54730a <=( (not A201)  and  (not A166) );
 a54733a <=( A232  and  A202 );
 a54734a <=( a54733a  and  a54730a );
 a54735a <=( a54734a  and  a54727a );
 a54738a <=( (not A234)  and  (not A233) );
 a54741a <=( (not A236)  and  (not A235) );
 a54742a <=( a54741a  and  a54738a );
 a54745a <=( A299  and  (not A298) );
 a54748a <=( A301  and  A300 );
 a54749a <=( a54748a  and  a54745a );
 a54750a <=( a54749a  and  a54742a );
 a54753a <=( (not A169)  and  A170 );
 a54756a <=( A167  and  (not A168) );
 a54757a <=( a54756a  and  a54753a );
 a54760a <=( (not A201)  and  (not A166) );
 a54763a <=( A232  and  A202 );
 a54764a <=( a54763a  and  a54760a );
 a54765a <=( a54764a  and  a54757a );
 a54768a <=( (not A234)  and  (not A233) );
 a54771a <=( (not A236)  and  (not A235) );
 a54772a <=( a54771a  and  a54768a );
 a54775a <=( A299  and  (not A298) );
 a54778a <=( A302  and  A300 );
 a54779a <=( a54778a  and  a54775a );
 a54780a <=( a54779a  and  a54772a );
 a54783a <=( (not A169)  and  A170 );
 a54786a <=( A167  and  (not A168) );
 a54787a <=( a54786a  and  a54783a );
 a54790a <=( (not A201)  and  (not A166) );
 a54793a <=( A232  and  A202 );
 a54794a <=( a54793a  and  a54790a );
 a54795a <=( a54794a  and  a54787a );
 a54798a <=( (not A234)  and  (not A233) );
 a54801a <=( (not A236)  and  (not A235) );
 a54802a <=( a54801a  and  a54798a );
 a54805a <=( A266  and  (not A265) );
 a54808a <=( A268  and  A267 );
 a54809a <=( a54808a  and  a54805a );
 a54810a <=( a54809a  and  a54802a );
 a54813a <=( (not A169)  and  A170 );
 a54816a <=( A167  and  (not A168) );
 a54817a <=( a54816a  and  a54813a );
 a54820a <=( (not A201)  and  (not A166) );
 a54823a <=( A232  and  A202 );
 a54824a <=( a54823a  and  a54820a );
 a54825a <=( a54824a  and  a54817a );
 a54828a <=( (not A234)  and  (not A233) );
 a54831a <=( (not A236)  and  (not A235) );
 a54832a <=( a54831a  and  a54828a );
 a54835a <=( A266  and  (not A265) );
 a54838a <=( A269  and  A267 );
 a54839a <=( a54838a  and  a54835a );
 a54840a <=( a54839a  and  a54832a );
 a54843a <=( (not A169)  and  A170 );
 a54846a <=( A167  and  (not A168) );
 a54847a <=( a54846a  and  a54843a );
 a54850a <=( (not A201)  and  (not A166) );
 a54853a <=( A232  and  A202 );
 a54854a <=( a54853a  and  a54850a );
 a54855a <=( a54854a  and  a54847a );
 a54858a <=( (not A234)  and  (not A233) );
 a54861a <=( (not A236)  and  (not A235) );
 a54862a <=( a54861a  and  a54858a );
 a54865a <=( (not A266)  and  A265 );
 a54868a <=( A268  and  A267 );
 a54869a <=( a54868a  and  a54865a );
 a54870a <=( a54869a  and  a54862a );
 a54873a <=( (not A169)  and  A170 );
 a54876a <=( A167  and  (not A168) );
 a54877a <=( a54876a  and  a54873a );
 a54880a <=( (not A201)  and  (not A166) );
 a54883a <=( A232  and  A202 );
 a54884a <=( a54883a  and  a54880a );
 a54885a <=( a54884a  and  a54877a );
 a54888a <=( (not A234)  and  (not A233) );
 a54891a <=( (not A236)  and  (not A235) );
 a54892a <=( a54891a  and  a54888a );
 a54895a <=( (not A266)  and  A265 );
 a54898a <=( A269  and  A267 );
 a54899a <=( a54898a  and  a54895a );
 a54900a <=( a54899a  and  a54892a );
 a54903a <=( (not A169)  and  A170 );
 a54906a <=( A167  and  (not A168) );
 a54907a <=( a54906a  and  a54903a );
 a54910a <=( (not A201)  and  (not A166) );
 a54913a <=( (not A232)  and  A203 );
 a54914a <=( a54913a  and  a54910a );
 a54915a <=( a54914a  and  a54907a );
 a54918a <=( A234  and  A233 );
 a54921a <=( A298  and  A235 );
 a54922a <=( a54921a  and  a54918a );
 a54925a <=( (not A300)  and  (not A299) );
 a54928a <=( (not A302)  and  (not A301) );
 a54929a <=( a54928a  and  a54925a );
 a54930a <=( a54929a  and  a54922a );
 a54933a <=( (not A169)  and  A170 );
 a54936a <=( A167  and  (not A168) );
 a54937a <=( a54936a  and  a54933a );
 a54940a <=( (not A201)  and  (not A166) );
 a54943a <=( (not A232)  and  A203 );
 a54944a <=( a54943a  and  a54940a );
 a54945a <=( a54944a  and  a54937a );
 a54948a <=( A234  and  A233 );
 a54951a <=( (not A298)  and  A235 );
 a54952a <=( a54951a  and  a54948a );
 a54955a <=( (not A300)  and  A299 );
 a54958a <=( (not A302)  and  (not A301) );
 a54959a <=( a54958a  and  a54955a );
 a54960a <=( a54959a  and  a54952a );
 a54963a <=( (not A169)  and  A170 );
 a54966a <=( A167  and  (not A168) );
 a54967a <=( a54966a  and  a54963a );
 a54970a <=( (not A201)  and  (not A166) );
 a54973a <=( (not A232)  and  A203 );
 a54974a <=( a54973a  and  a54970a );
 a54975a <=( a54974a  and  a54967a );
 a54978a <=( A234  and  A233 );
 a54981a <=( (not A265)  and  A235 );
 a54982a <=( a54981a  and  a54978a );
 a54985a <=( (not A267)  and  A266 );
 a54988a <=( (not A269)  and  (not A268) );
 a54989a <=( a54988a  and  a54985a );
 a54990a <=( a54989a  and  a54982a );
 a54993a <=( (not A169)  and  A170 );
 a54996a <=( A167  and  (not A168) );
 a54997a <=( a54996a  and  a54993a );
 a55000a <=( (not A201)  and  (not A166) );
 a55003a <=( (not A232)  and  A203 );
 a55004a <=( a55003a  and  a55000a );
 a55005a <=( a55004a  and  a54997a );
 a55008a <=( A234  and  A233 );
 a55011a <=( A265  and  A235 );
 a55012a <=( a55011a  and  a55008a );
 a55015a <=( (not A267)  and  (not A266) );
 a55018a <=( (not A269)  and  (not A268) );
 a55019a <=( a55018a  and  a55015a );
 a55020a <=( a55019a  and  a55012a );
 a55023a <=( (not A169)  and  A170 );
 a55026a <=( A167  and  (not A168) );
 a55027a <=( a55026a  and  a55023a );
 a55030a <=( (not A201)  and  (not A166) );
 a55033a <=( (not A232)  and  A203 );
 a55034a <=( a55033a  and  a55030a );
 a55035a <=( a55034a  and  a55027a );
 a55038a <=( A234  and  A233 );
 a55041a <=( A298  and  A236 );
 a55042a <=( a55041a  and  a55038a );
 a55045a <=( (not A300)  and  (not A299) );
 a55048a <=( (not A302)  and  (not A301) );
 a55049a <=( a55048a  and  a55045a );
 a55050a <=( a55049a  and  a55042a );
 a55053a <=( (not A169)  and  A170 );
 a55056a <=( A167  and  (not A168) );
 a55057a <=( a55056a  and  a55053a );
 a55060a <=( (not A201)  and  (not A166) );
 a55063a <=( (not A232)  and  A203 );
 a55064a <=( a55063a  and  a55060a );
 a55065a <=( a55064a  and  a55057a );
 a55068a <=( A234  and  A233 );
 a55071a <=( (not A298)  and  A236 );
 a55072a <=( a55071a  and  a55068a );
 a55075a <=( (not A300)  and  A299 );
 a55078a <=( (not A302)  and  (not A301) );
 a55079a <=( a55078a  and  a55075a );
 a55080a <=( a55079a  and  a55072a );
 a55083a <=( (not A169)  and  A170 );
 a55086a <=( A167  and  (not A168) );
 a55087a <=( a55086a  and  a55083a );
 a55090a <=( (not A201)  and  (not A166) );
 a55093a <=( (not A232)  and  A203 );
 a55094a <=( a55093a  and  a55090a );
 a55095a <=( a55094a  and  a55087a );
 a55098a <=( A234  and  A233 );
 a55101a <=( (not A265)  and  A236 );
 a55102a <=( a55101a  and  a55098a );
 a55105a <=( (not A267)  and  A266 );
 a55108a <=( (not A269)  and  (not A268) );
 a55109a <=( a55108a  and  a55105a );
 a55110a <=( a55109a  and  a55102a );
 a55113a <=( (not A169)  and  A170 );
 a55116a <=( A167  and  (not A168) );
 a55117a <=( a55116a  and  a55113a );
 a55120a <=( (not A201)  and  (not A166) );
 a55123a <=( (not A232)  and  A203 );
 a55124a <=( a55123a  and  a55120a );
 a55125a <=( a55124a  and  a55117a );
 a55128a <=( A234  and  A233 );
 a55131a <=( A265  and  A236 );
 a55132a <=( a55131a  and  a55128a );
 a55135a <=( (not A267)  and  (not A266) );
 a55138a <=( (not A269)  and  (not A268) );
 a55139a <=( a55138a  and  a55135a );
 a55140a <=( a55139a  and  a55132a );
 a55143a <=( (not A169)  and  A170 );
 a55146a <=( A167  and  (not A168) );
 a55147a <=( a55146a  and  a55143a );
 a55150a <=( (not A201)  and  (not A166) );
 a55153a <=( (not A232)  and  A203 );
 a55154a <=( a55153a  and  a55150a );
 a55155a <=( a55154a  and  a55147a );
 a55158a <=( (not A234)  and  A233 );
 a55161a <=( (not A236)  and  (not A235) );
 a55162a <=( a55161a  and  a55158a );
 a55165a <=( (not A299)  and  A298 );
 a55168a <=( A301  and  A300 );
 a55169a <=( a55168a  and  a55165a );
 a55170a <=( a55169a  and  a55162a );
 a55173a <=( (not A169)  and  A170 );
 a55176a <=( A167  and  (not A168) );
 a55177a <=( a55176a  and  a55173a );
 a55180a <=( (not A201)  and  (not A166) );
 a55183a <=( (not A232)  and  A203 );
 a55184a <=( a55183a  and  a55180a );
 a55185a <=( a55184a  and  a55177a );
 a55188a <=( (not A234)  and  A233 );
 a55191a <=( (not A236)  and  (not A235) );
 a55192a <=( a55191a  and  a55188a );
 a55195a <=( (not A299)  and  A298 );
 a55198a <=( A302  and  A300 );
 a55199a <=( a55198a  and  a55195a );
 a55200a <=( a55199a  and  a55192a );
 a55203a <=( (not A169)  and  A170 );
 a55206a <=( A167  and  (not A168) );
 a55207a <=( a55206a  and  a55203a );
 a55210a <=( (not A201)  and  (not A166) );
 a55213a <=( (not A232)  and  A203 );
 a55214a <=( a55213a  and  a55210a );
 a55215a <=( a55214a  and  a55207a );
 a55218a <=( (not A234)  and  A233 );
 a55221a <=( (not A236)  and  (not A235) );
 a55222a <=( a55221a  and  a55218a );
 a55225a <=( A299  and  (not A298) );
 a55228a <=( A301  and  A300 );
 a55229a <=( a55228a  and  a55225a );
 a55230a <=( a55229a  and  a55222a );
 a55233a <=( (not A169)  and  A170 );
 a55236a <=( A167  and  (not A168) );
 a55237a <=( a55236a  and  a55233a );
 a55240a <=( (not A201)  and  (not A166) );
 a55243a <=( (not A232)  and  A203 );
 a55244a <=( a55243a  and  a55240a );
 a55245a <=( a55244a  and  a55237a );
 a55248a <=( (not A234)  and  A233 );
 a55251a <=( (not A236)  and  (not A235) );
 a55252a <=( a55251a  and  a55248a );
 a55255a <=( A299  and  (not A298) );
 a55258a <=( A302  and  A300 );
 a55259a <=( a55258a  and  a55255a );
 a55260a <=( a55259a  and  a55252a );
 a55263a <=( (not A169)  and  A170 );
 a55266a <=( A167  and  (not A168) );
 a55267a <=( a55266a  and  a55263a );
 a55270a <=( (not A201)  and  (not A166) );
 a55273a <=( (not A232)  and  A203 );
 a55274a <=( a55273a  and  a55270a );
 a55275a <=( a55274a  and  a55267a );
 a55278a <=( (not A234)  and  A233 );
 a55281a <=( (not A236)  and  (not A235) );
 a55282a <=( a55281a  and  a55278a );
 a55285a <=( A266  and  (not A265) );
 a55288a <=( A268  and  A267 );
 a55289a <=( a55288a  and  a55285a );
 a55290a <=( a55289a  and  a55282a );
 a55293a <=( (not A169)  and  A170 );
 a55296a <=( A167  and  (not A168) );
 a55297a <=( a55296a  and  a55293a );
 a55300a <=( (not A201)  and  (not A166) );
 a55303a <=( (not A232)  and  A203 );
 a55304a <=( a55303a  and  a55300a );
 a55305a <=( a55304a  and  a55297a );
 a55308a <=( (not A234)  and  A233 );
 a55311a <=( (not A236)  and  (not A235) );
 a55312a <=( a55311a  and  a55308a );
 a55315a <=( A266  and  (not A265) );
 a55318a <=( A269  and  A267 );
 a55319a <=( a55318a  and  a55315a );
 a55320a <=( a55319a  and  a55312a );
 a55323a <=( (not A169)  and  A170 );
 a55326a <=( A167  and  (not A168) );
 a55327a <=( a55326a  and  a55323a );
 a55330a <=( (not A201)  and  (not A166) );
 a55333a <=( (not A232)  and  A203 );
 a55334a <=( a55333a  and  a55330a );
 a55335a <=( a55334a  and  a55327a );
 a55338a <=( (not A234)  and  A233 );
 a55341a <=( (not A236)  and  (not A235) );
 a55342a <=( a55341a  and  a55338a );
 a55345a <=( (not A266)  and  A265 );
 a55348a <=( A268  and  A267 );
 a55349a <=( a55348a  and  a55345a );
 a55350a <=( a55349a  and  a55342a );
 a55353a <=( (not A169)  and  A170 );
 a55356a <=( A167  and  (not A168) );
 a55357a <=( a55356a  and  a55353a );
 a55360a <=( (not A201)  and  (not A166) );
 a55363a <=( (not A232)  and  A203 );
 a55364a <=( a55363a  and  a55360a );
 a55365a <=( a55364a  and  a55357a );
 a55368a <=( (not A234)  and  A233 );
 a55371a <=( (not A236)  and  (not A235) );
 a55372a <=( a55371a  and  a55368a );
 a55375a <=( (not A266)  and  A265 );
 a55378a <=( A269  and  A267 );
 a55379a <=( a55378a  and  a55375a );
 a55380a <=( a55379a  and  a55372a );
 a55383a <=( (not A169)  and  A170 );
 a55386a <=( A167  and  (not A168) );
 a55387a <=( a55386a  and  a55383a );
 a55390a <=( (not A201)  and  (not A166) );
 a55393a <=( A232  and  A203 );
 a55394a <=( a55393a  and  a55390a );
 a55395a <=( a55394a  and  a55387a );
 a55398a <=( A234  and  (not A233) );
 a55401a <=( A298  and  A235 );
 a55402a <=( a55401a  and  a55398a );
 a55405a <=( (not A300)  and  (not A299) );
 a55408a <=( (not A302)  and  (not A301) );
 a55409a <=( a55408a  and  a55405a );
 a55410a <=( a55409a  and  a55402a );
 a55413a <=( (not A169)  and  A170 );
 a55416a <=( A167  and  (not A168) );
 a55417a <=( a55416a  and  a55413a );
 a55420a <=( (not A201)  and  (not A166) );
 a55423a <=( A232  and  A203 );
 a55424a <=( a55423a  and  a55420a );
 a55425a <=( a55424a  and  a55417a );
 a55428a <=( A234  and  (not A233) );
 a55431a <=( (not A298)  and  A235 );
 a55432a <=( a55431a  and  a55428a );
 a55435a <=( (not A300)  and  A299 );
 a55438a <=( (not A302)  and  (not A301) );
 a55439a <=( a55438a  and  a55435a );
 a55440a <=( a55439a  and  a55432a );
 a55443a <=( (not A169)  and  A170 );
 a55446a <=( A167  and  (not A168) );
 a55447a <=( a55446a  and  a55443a );
 a55450a <=( (not A201)  and  (not A166) );
 a55453a <=( A232  and  A203 );
 a55454a <=( a55453a  and  a55450a );
 a55455a <=( a55454a  and  a55447a );
 a55458a <=( A234  and  (not A233) );
 a55461a <=( (not A265)  and  A235 );
 a55462a <=( a55461a  and  a55458a );
 a55465a <=( (not A267)  and  A266 );
 a55468a <=( (not A269)  and  (not A268) );
 a55469a <=( a55468a  and  a55465a );
 a55470a <=( a55469a  and  a55462a );
 a55473a <=( (not A169)  and  A170 );
 a55476a <=( A167  and  (not A168) );
 a55477a <=( a55476a  and  a55473a );
 a55480a <=( (not A201)  and  (not A166) );
 a55483a <=( A232  and  A203 );
 a55484a <=( a55483a  and  a55480a );
 a55485a <=( a55484a  and  a55477a );
 a55488a <=( A234  and  (not A233) );
 a55491a <=( A265  and  A235 );
 a55492a <=( a55491a  and  a55488a );
 a55495a <=( (not A267)  and  (not A266) );
 a55498a <=( (not A269)  and  (not A268) );
 a55499a <=( a55498a  and  a55495a );
 a55500a <=( a55499a  and  a55492a );
 a55503a <=( (not A169)  and  A170 );
 a55506a <=( A167  and  (not A168) );
 a55507a <=( a55506a  and  a55503a );
 a55510a <=( (not A201)  and  (not A166) );
 a55513a <=( A232  and  A203 );
 a55514a <=( a55513a  and  a55510a );
 a55515a <=( a55514a  and  a55507a );
 a55518a <=( A234  and  (not A233) );
 a55521a <=( A298  and  A236 );
 a55522a <=( a55521a  and  a55518a );
 a55525a <=( (not A300)  and  (not A299) );
 a55528a <=( (not A302)  and  (not A301) );
 a55529a <=( a55528a  and  a55525a );
 a55530a <=( a55529a  and  a55522a );
 a55533a <=( (not A169)  and  A170 );
 a55536a <=( A167  and  (not A168) );
 a55537a <=( a55536a  and  a55533a );
 a55540a <=( (not A201)  and  (not A166) );
 a55543a <=( A232  and  A203 );
 a55544a <=( a55543a  and  a55540a );
 a55545a <=( a55544a  and  a55537a );
 a55548a <=( A234  and  (not A233) );
 a55551a <=( (not A298)  and  A236 );
 a55552a <=( a55551a  and  a55548a );
 a55555a <=( (not A300)  and  A299 );
 a55558a <=( (not A302)  and  (not A301) );
 a55559a <=( a55558a  and  a55555a );
 a55560a <=( a55559a  and  a55552a );
 a55563a <=( (not A169)  and  A170 );
 a55566a <=( A167  and  (not A168) );
 a55567a <=( a55566a  and  a55563a );
 a55570a <=( (not A201)  and  (not A166) );
 a55573a <=( A232  and  A203 );
 a55574a <=( a55573a  and  a55570a );
 a55575a <=( a55574a  and  a55567a );
 a55578a <=( A234  and  (not A233) );
 a55581a <=( (not A265)  and  A236 );
 a55582a <=( a55581a  and  a55578a );
 a55585a <=( (not A267)  and  A266 );
 a55588a <=( (not A269)  and  (not A268) );
 a55589a <=( a55588a  and  a55585a );
 a55590a <=( a55589a  and  a55582a );
 a55593a <=( (not A169)  and  A170 );
 a55596a <=( A167  and  (not A168) );
 a55597a <=( a55596a  and  a55593a );
 a55600a <=( (not A201)  and  (not A166) );
 a55603a <=( A232  and  A203 );
 a55604a <=( a55603a  and  a55600a );
 a55605a <=( a55604a  and  a55597a );
 a55608a <=( A234  and  (not A233) );
 a55611a <=( A265  and  A236 );
 a55612a <=( a55611a  and  a55608a );
 a55615a <=( (not A267)  and  (not A266) );
 a55618a <=( (not A269)  and  (not A268) );
 a55619a <=( a55618a  and  a55615a );
 a55620a <=( a55619a  and  a55612a );
 a55623a <=( (not A169)  and  A170 );
 a55626a <=( A167  and  (not A168) );
 a55627a <=( a55626a  and  a55623a );
 a55630a <=( (not A201)  and  (not A166) );
 a55633a <=( A232  and  A203 );
 a55634a <=( a55633a  and  a55630a );
 a55635a <=( a55634a  and  a55627a );
 a55638a <=( (not A234)  and  (not A233) );
 a55641a <=( (not A236)  and  (not A235) );
 a55642a <=( a55641a  and  a55638a );
 a55645a <=( (not A299)  and  A298 );
 a55648a <=( A301  and  A300 );
 a55649a <=( a55648a  and  a55645a );
 a55650a <=( a55649a  and  a55642a );
 a55653a <=( (not A169)  and  A170 );
 a55656a <=( A167  and  (not A168) );
 a55657a <=( a55656a  and  a55653a );
 a55660a <=( (not A201)  and  (not A166) );
 a55663a <=( A232  and  A203 );
 a55664a <=( a55663a  and  a55660a );
 a55665a <=( a55664a  and  a55657a );
 a55668a <=( (not A234)  and  (not A233) );
 a55671a <=( (not A236)  and  (not A235) );
 a55672a <=( a55671a  and  a55668a );
 a55675a <=( (not A299)  and  A298 );
 a55678a <=( A302  and  A300 );
 a55679a <=( a55678a  and  a55675a );
 a55680a <=( a55679a  and  a55672a );
 a55683a <=( (not A169)  and  A170 );
 a55686a <=( A167  and  (not A168) );
 a55687a <=( a55686a  and  a55683a );
 a55690a <=( (not A201)  and  (not A166) );
 a55693a <=( A232  and  A203 );
 a55694a <=( a55693a  and  a55690a );
 a55695a <=( a55694a  and  a55687a );
 a55698a <=( (not A234)  and  (not A233) );
 a55701a <=( (not A236)  and  (not A235) );
 a55702a <=( a55701a  and  a55698a );
 a55705a <=( A299  and  (not A298) );
 a55708a <=( A301  and  A300 );
 a55709a <=( a55708a  and  a55705a );
 a55710a <=( a55709a  and  a55702a );
 a55713a <=( (not A169)  and  A170 );
 a55716a <=( A167  and  (not A168) );
 a55717a <=( a55716a  and  a55713a );
 a55720a <=( (not A201)  and  (not A166) );
 a55723a <=( A232  and  A203 );
 a55724a <=( a55723a  and  a55720a );
 a55725a <=( a55724a  and  a55717a );
 a55728a <=( (not A234)  and  (not A233) );
 a55731a <=( (not A236)  and  (not A235) );
 a55732a <=( a55731a  and  a55728a );
 a55735a <=( A299  and  (not A298) );
 a55738a <=( A302  and  A300 );
 a55739a <=( a55738a  and  a55735a );
 a55740a <=( a55739a  and  a55732a );
 a55743a <=( (not A169)  and  A170 );
 a55746a <=( A167  and  (not A168) );
 a55747a <=( a55746a  and  a55743a );
 a55750a <=( (not A201)  and  (not A166) );
 a55753a <=( A232  and  A203 );
 a55754a <=( a55753a  and  a55750a );
 a55755a <=( a55754a  and  a55747a );
 a55758a <=( (not A234)  and  (not A233) );
 a55761a <=( (not A236)  and  (not A235) );
 a55762a <=( a55761a  and  a55758a );
 a55765a <=( A266  and  (not A265) );
 a55768a <=( A268  and  A267 );
 a55769a <=( a55768a  and  a55765a );
 a55770a <=( a55769a  and  a55762a );
 a55773a <=( (not A169)  and  A170 );
 a55776a <=( A167  and  (not A168) );
 a55777a <=( a55776a  and  a55773a );
 a55780a <=( (not A201)  and  (not A166) );
 a55783a <=( A232  and  A203 );
 a55784a <=( a55783a  and  a55780a );
 a55785a <=( a55784a  and  a55777a );
 a55788a <=( (not A234)  and  (not A233) );
 a55791a <=( (not A236)  and  (not A235) );
 a55792a <=( a55791a  and  a55788a );
 a55795a <=( A266  and  (not A265) );
 a55798a <=( A269  and  A267 );
 a55799a <=( a55798a  and  a55795a );
 a55800a <=( a55799a  and  a55792a );
 a55803a <=( (not A169)  and  A170 );
 a55806a <=( A167  and  (not A168) );
 a55807a <=( a55806a  and  a55803a );
 a55810a <=( (not A201)  and  (not A166) );
 a55813a <=( A232  and  A203 );
 a55814a <=( a55813a  and  a55810a );
 a55815a <=( a55814a  and  a55807a );
 a55818a <=( (not A234)  and  (not A233) );
 a55821a <=( (not A236)  and  (not A235) );
 a55822a <=( a55821a  and  a55818a );
 a55825a <=( (not A266)  and  A265 );
 a55828a <=( A268  and  A267 );
 a55829a <=( a55828a  and  a55825a );
 a55830a <=( a55829a  and  a55822a );
 a55833a <=( (not A169)  and  A170 );
 a55836a <=( A167  and  (not A168) );
 a55837a <=( a55836a  and  a55833a );
 a55840a <=( (not A201)  and  (not A166) );
 a55843a <=( A232  and  A203 );
 a55844a <=( a55843a  and  a55840a );
 a55845a <=( a55844a  and  a55837a );
 a55848a <=( (not A234)  and  (not A233) );
 a55851a <=( (not A236)  and  (not A235) );
 a55852a <=( a55851a  and  a55848a );
 a55855a <=( (not A266)  and  A265 );
 a55858a <=( A269  and  A267 );
 a55859a <=( a55858a  and  a55855a );
 a55860a <=( a55859a  and  a55852a );
 a55863a <=( (not A169)  and  A170 );
 a55866a <=( A167  and  (not A168) );
 a55867a <=( a55866a  and  a55863a );
 a55870a <=( A199  and  (not A166) );
 a55873a <=( (not A232)  and  A200 );
 a55874a <=( a55873a  and  a55870a );
 a55875a <=( a55874a  and  a55867a );
 a55878a <=( A234  and  A233 );
 a55881a <=( A298  and  A235 );
 a55882a <=( a55881a  and  a55878a );
 a55885a <=( (not A300)  and  (not A299) );
 a55888a <=( (not A302)  and  (not A301) );
 a55889a <=( a55888a  and  a55885a );
 a55890a <=( a55889a  and  a55882a );
 a55893a <=( (not A169)  and  A170 );
 a55896a <=( A167  and  (not A168) );
 a55897a <=( a55896a  and  a55893a );
 a55900a <=( A199  and  (not A166) );
 a55903a <=( (not A232)  and  A200 );
 a55904a <=( a55903a  and  a55900a );
 a55905a <=( a55904a  and  a55897a );
 a55908a <=( A234  and  A233 );
 a55911a <=( (not A298)  and  A235 );
 a55912a <=( a55911a  and  a55908a );
 a55915a <=( (not A300)  and  A299 );
 a55918a <=( (not A302)  and  (not A301) );
 a55919a <=( a55918a  and  a55915a );
 a55920a <=( a55919a  and  a55912a );
 a55923a <=( (not A169)  and  A170 );
 a55926a <=( A167  and  (not A168) );
 a55927a <=( a55926a  and  a55923a );
 a55930a <=( A199  and  (not A166) );
 a55933a <=( (not A232)  and  A200 );
 a55934a <=( a55933a  and  a55930a );
 a55935a <=( a55934a  and  a55927a );
 a55938a <=( A234  and  A233 );
 a55941a <=( (not A265)  and  A235 );
 a55942a <=( a55941a  and  a55938a );
 a55945a <=( (not A267)  and  A266 );
 a55948a <=( (not A269)  and  (not A268) );
 a55949a <=( a55948a  and  a55945a );
 a55950a <=( a55949a  and  a55942a );
 a55953a <=( (not A169)  and  A170 );
 a55956a <=( A167  and  (not A168) );
 a55957a <=( a55956a  and  a55953a );
 a55960a <=( A199  and  (not A166) );
 a55963a <=( (not A232)  and  A200 );
 a55964a <=( a55963a  and  a55960a );
 a55965a <=( a55964a  and  a55957a );
 a55968a <=( A234  and  A233 );
 a55971a <=( A265  and  A235 );
 a55972a <=( a55971a  and  a55968a );
 a55975a <=( (not A267)  and  (not A266) );
 a55978a <=( (not A269)  and  (not A268) );
 a55979a <=( a55978a  and  a55975a );
 a55980a <=( a55979a  and  a55972a );
 a55983a <=( (not A169)  and  A170 );
 a55986a <=( A167  and  (not A168) );
 a55987a <=( a55986a  and  a55983a );
 a55990a <=( A199  and  (not A166) );
 a55993a <=( (not A232)  and  A200 );
 a55994a <=( a55993a  and  a55990a );
 a55995a <=( a55994a  and  a55987a );
 a55998a <=( A234  and  A233 );
 a56001a <=( A298  and  A236 );
 a56002a <=( a56001a  and  a55998a );
 a56005a <=( (not A300)  and  (not A299) );
 a56008a <=( (not A302)  and  (not A301) );
 a56009a <=( a56008a  and  a56005a );
 a56010a <=( a56009a  and  a56002a );
 a56013a <=( (not A169)  and  A170 );
 a56016a <=( A167  and  (not A168) );
 a56017a <=( a56016a  and  a56013a );
 a56020a <=( A199  and  (not A166) );
 a56023a <=( (not A232)  and  A200 );
 a56024a <=( a56023a  and  a56020a );
 a56025a <=( a56024a  and  a56017a );
 a56028a <=( A234  and  A233 );
 a56031a <=( (not A298)  and  A236 );
 a56032a <=( a56031a  and  a56028a );
 a56035a <=( (not A300)  and  A299 );
 a56038a <=( (not A302)  and  (not A301) );
 a56039a <=( a56038a  and  a56035a );
 a56040a <=( a56039a  and  a56032a );
 a56043a <=( (not A169)  and  A170 );
 a56046a <=( A167  and  (not A168) );
 a56047a <=( a56046a  and  a56043a );
 a56050a <=( A199  and  (not A166) );
 a56053a <=( (not A232)  and  A200 );
 a56054a <=( a56053a  and  a56050a );
 a56055a <=( a56054a  and  a56047a );
 a56058a <=( A234  and  A233 );
 a56061a <=( (not A265)  and  A236 );
 a56062a <=( a56061a  and  a56058a );
 a56065a <=( (not A267)  and  A266 );
 a56068a <=( (not A269)  and  (not A268) );
 a56069a <=( a56068a  and  a56065a );
 a56070a <=( a56069a  and  a56062a );
 a56073a <=( (not A169)  and  A170 );
 a56076a <=( A167  and  (not A168) );
 a56077a <=( a56076a  and  a56073a );
 a56080a <=( A199  and  (not A166) );
 a56083a <=( (not A232)  and  A200 );
 a56084a <=( a56083a  and  a56080a );
 a56085a <=( a56084a  and  a56077a );
 a56088a <=( A234  and  A233 );
 a56091a <=( A265  and  A236 );
 a56092a <=( a56091a  and  a56088a );
 a56095a <=( (not A267)  and  (not A266) );
 a56098a <=( (not A269)  and  (not A268) );
 a56099a <=( a56098a  and  a56095a );
 a56100a <=( a56099a  and  a56092a );
 a56103a <=( (not A169)  and  A170 );
 a56106a <=( A167  and  (not A168) );
 a56107a <=( a56106a  and  a56103a );
 a56110a <=( A199  and  (not A166) );
 a56113a <=( (not A232)  and  A200 );
 a56114a <=( a56113a  and  a56110a );
 a56115a <=( a56114a  and  a56107a );
 a56118a <=( (not A234)  and  A233 );
 a56121a <=( (not A236)  and  (not A235) );
 a56122a <=( a56121a  and  a56118a );
 a56125a <=( (not A299)  and  A298 );
 a56128a <=( A301  and  A300 );
 a56129a <=( a56128a  and  a56125a );
 a56130a <=( a56129a  and  a56122a );
 a56133a <=( (not A169)  and  A170 );
 a56136a <=( A167  and  (not A168) );
 a56137a <=( a56136a  and  a56133a );
 a56140a <=( A199  and  (not A166) );
 a56143a <=( (not A232)  and  A200 );
 a56144a <=( a56143a  and  a56140a );
 a56145a <=( a56144a  and  a56137a );
 a56148a <=( (not A234)  and  A233 );
 a56151a <=( (not A236)  and  (not A235) );
 a56152a <=( a56151a  and  a56148a );
 a56155a <=( (not A299)  and  A298 );
 a56158a <=( A302  and  A300 );
 a56159a <=( a56158a  and  a56155a );
 a56160a <=( a56159a  and  a56152a );
 a56163a <=( (not A169)  and  A170 );
 a56166a <=( A167  and  (not A168) );
 a56167a <=( a56166a  and  a56163a );
 a56170a <=( A199  and  (not A166) );
 a56173a <=( (not A232)  and  A200 );
 a56174a <=( a56173a  and  a56170a );
 a56175a <=( a56174a  and  a56167a );
 a56178a <=( (not A234)  and  A233 );
 a56181a <=( (not A236)  and  (not A235) );
 a56182a <=( a56181a  and  a56178a );
 a56185a <=( A299  and  (not A298) );
 a56188a <=( A301  and  A300 );
 a56189a <=( a56188a  and  a56185a );
 a56190a <=( a56189a  and  a56182a );
 a56193a <=( (not A169)  and  A170 );
 a56196a <=( A167  and  (not A168) );
 a56197a <=( a56196a  and  a56193a );
 a56200a <=( A199  and  (not A166) );
 a56203a <=( (not A232)  and  A200 );
 a56204a <=( a56203a  and  a56200a );
 a56205a <=( a56204a  and  a56197a );
 a56208a <=( (not A234)  and  A233 );
 a56211a <=( (not A236)  and  (not A235) );
 a56212a <=( a56211a  and  a56208a );
 a56215a <=( A299  and  (not A298) );
 a56218a <=( A302  and  A300 );
 a56219a <=( a56218a  and  a56215a );
 a56220a <=( a56219a  and  a56212a );
 a56223a <=( (not A169)  and  A170 );
 a56226a <=( A167  and  (not A168) );
 a56227a <=( a56226a  and  a56223a );
 a56230a <=( A199  and  (not A166) );
 a56233a <=( (not A232)  and  A200 );
 a56234a <=( a56233a  and  a56230a );
 a56235a <=( a56234a  and  a56227a );
 a56238a <=( (not A234)  and  A233 );
 a56241a <=( (not A236)  and  (not A235) );
 a56242a <=( a56241a  and  a56238a );
 a56245a <=( A266  and  (not A265) );
 a56248a <=( A268  and  A267 );
 a56249a <=( a56248a  and  a56245a );
 a56250a <=( a56249a  and  a56242a );
 a56253a <=( (not A169)  and  A170 );
 a56256a <=( A167  and  (not A168) );
 a56257a <=( a56256a  and  a56253a );
 a56260a <=( A199  and  (not A166) );
 a56263a <=( (not A232)  and  A200 );
 a56264a <=( a56263a  and  a56260a );
 a56265a <=( a56264a  and  a56257a );
 a56268a <=( (not A234)  and  A233 );
 a56271a <=( (not A236)  and  (not A235) );
 a56272a <=( a56271a  and  a56268a );
 a56275a <=( A266  and  (not A265) );
 a56278a <=( A269  and  A267 );
 a56279a <=( a56278a  and  a56275a );
 a56280a <=( a56279a  and  a56272a );
 a56283a <=( (not A169)  and  A170 );
 a56286a <=( A167  and  (not A168) );
 a56287a <=( a56286a  and  a56283a );
 a56290a <=( A199  and  (not A166) );
 a56293a <=( (not A232)  and  A200 );
 a56294a <=( a56293a  and  a56290a );
 a56295a <=( a56294a  and  a56287a );
 a56298a <=( (not A234)  and  A233 );
 a56301a <=( (not A236)  and  (not A235) );
 a56302a <=( a56301a  and  a56298a );
 a56305a <=( (not A266)  and  A265 );
 a56308a <=( A268  and  A267 );
 a56309a <=( a56308a  and  a56305a );
 a56310a <=( a56309a  and  a56302a );
 a56313a <=( (not A169)  and  A170 );
 a56316a <=( A167  and  (not A168) );
 a56317a <=( a56316a  and  a56313a );
 a56320a <=( A199  and  (not A166) );
 a56323a <=( (not A232)  and  A200 );
 a56324a <=( a56323a  and  a56320a );
 a56325a <=( a56324a  and  a56317a );
 a56328a <=( (not A234)  and  A233 );
 a56331a <=( (not A236)  and  (not A235) );
 a56332a <=( a56331a  and  a56328a );
 a56335a <=( (not A266)  and  A265 );
 a56338a <=( A269  and  A267 );
 a56339a <=( a56338a  and  a56335a );
 a56340a <=( a56339a  and  a56332a );
 a56343a <=( (not A169)  and  A170 );
 a56346a <=( A167  and  (not A168) );
 a56347a <=( a56346a  and  a56343a );
 a56350a <=( A199  and  (not A166) );
 a56353a <=( A232  and  A200 );
 a56354a <=( a56353a  and  a56350a );
 a56355a <=( a56354a  and  a56347a );
 a56358a <=( A234  and  (not A233) );
 a56361a <=( A298  and  A235 );
 a56362a <=( a56361a  and  a56358a );
 a56365a <=( (not A300)  and  (not A299) );
 a56368a <=( (not A302)  and  (not A301) );
 a56369a <=( a56368a  and  a56365a );
 a56370a <=( a56369a  and  a56362a );
 a56373a <=( (not A169)  and  A170 );
 a56376a <=( A167  and  (not A168) );
 a56377a <=( a56376a  and  a56373a );
 a56380a <=( A199  and  (not A166) );
 a56383a <=( A232  and  A200 );
 a56384a <=( a56383a  and  a56380a );
 a56385a <=( a56384a  and  a56377a );
 a56388a <=( A234  and  (not A233) );
 a56391a <=( (not A298)  and  A235 );
 a56392a <=( a56391a  and  a56388a );
 a56395a <=( (not A300)  and  A299 );
 a56398a <=( (not A302)  and  (not A301) );
 a56399a <=( a56398a  and  a56395a );
 a56400a <=( a56399a  and  a56392a );
 a56403a <=( (not A169)  and  A170 );
 a56406a <=( A167  and  (not A168) );
 a56407a <=( a56406a  and  a56403a );
 a56410a <=( A199  and  (not A166) );
 a56413a <=( A232  and  A200 );
 a56414a <=( a56413a  and  a56410a );
 a56415a <=( a56414a  and  a56407a );
 a56418a <=( A234  and  (not A233) );
 a56421a <=( (not A265)  and  A235 );
 a56422a <=( a56421a  and  a56418a );
 a56425a <=( (not A267)  and  A266 );
 a56428a <=( (not A269)  and  (not A268) );
 a56429a <=( a56428a  and  a56425a );
 a56430a <=( a56429a  and  a56422a );
 a56433a <=( (not A169)  and  A170 );
 a56436a <=( A167  and  (not A168) );
 a56437a <=( a56436a  and  a56433a );
 a56440a <=( A199  and  (not A166) );
 a56443a <=( A232  and  A200 );
 a56444a <=( a56443a  and  a56440a );
 a56445a <=( a56444a  and  a56437a );
 a56448a <=( A234  and  (not A233) );
 a56451a <=( A265  and  A235 );
 a56452a <=( a56451a  and  a56448a );
 a56455a <=( (not A267)  and  (not A266) );
 a56458a <=( (not A269)  and  (not A268) );
 a56459a <=( a56458a  and  a56455a );
 a56460a <=( a56459a  and  a56452a );
 a56463a <=( (not A169)  and  A170 );
 a56466a <=( A167  and  (not A168) );
 a56467a <=( a56466a  and  a56463a );
 a56470a <=( A199  and  (not A166) );
 a56473a <=( A232  and  A200 );
 a56474a <=( a56473a  and  a56470a );
 a56475a <=( a56474a  and  a56467a );
 a56478a <=( A234  and  (not A233) );
 a56481a <=( A298  and  A236 );
 a56482a <=( a56481a  and  a56478a );
 a56485a <=( (not A300)  and  (not A299) );
 a56488a <=( (not A302)  and  (not A301) );
 a56489a <=( a56488a  and  a56485a );
 a56490a <=( a56489a  and  a56482a );
 a56493a <=( (not A169)  and  A170 );
 a56496a <=( A167  and  (not A168) );
 a56497a <=( a56496a  and  a56493a );
 a56500a <=( A199  and  (not A166) );
 a56503a <=( A232  and  A200 );
 a56504a <=( a56503a  and  a56500a );
 a56505a <=( a56504a  and  a56497a );
 a56508a <=( A234  and  (not A233) );
 a56511a <=( (not A298)  and  A236 );
 a56512a <=( a56511a  and  a56508a );
 a56515a <=( (not A300)  and  A299 );
 a56518a <=( (not A302)  and  (not A301) );
 a56519a <=( a56518a  and  a56515a );
 a56520a <=( a56519a  and  a56512a );
 a56523a <=( (not A169)  and  A170 );
 a56526a <=( A167  and  (not A168) );
 a56527a <=( a56526a  and  a56523a );
 a56530a <=( A199  and  (not A166) );
 a56533a <=( A232  and  A200 );
 a56534a <=( a56533a  and  a56530a );
 a56535a <=( a56534a  and  a56527a );
 a56538a <=( A234  and  (not A233) );
 a56541a <=( (not A265)  and  A236 );
 a56542a <=( a56541a  and  a56538a );
 a56545a <=( (not A267)  and  A266 );
 a56548a <=( (not A269)  and  (not A268) );
 a56549a <=( a56548a  and  a56545a );
 a56550a <=( a56549a  and  a56542a );
 a56553a <=( (not A169)  and  A170 );
 a56556a <=( A167  and  (not A168) );
 a56557a <=( a56556a  and  a56553a );
 a56560a <=( A199  and  (not A166) );
 a56563a <=( A232  and  A200 );
 a56564a <=( a56563a  and  a56560a );
 a56565a <=( a56564a  and  a56557a );
 a56568a <=( A234  and  (not A233) );
 a56571a <=( A265  and  A236 );
 a56572a <=( a56571a  and  a56568a );
 a56575a <=( (not A267)  and  (not A266) );
 a56578a <=( (not A269)  and  (not A268) );
 a56579a <=( a56578a  and  a56575a );
 a56580a <=( a56579a  and  a56572a );
 a56583a <=( (not A169)  and  A170 );
 a56586a <=( A167  and  (not A168) );
 a56587a <=( a56586a  and  a56583a );
 a56590a <=( A199  and  (not A166) );
 a56593a <=( A232  and  A200 );
 a56594a <=( a56593a  and  a56590a );
 a56595a <=( a56594a  and  a56587a );
 a56598a <=( (not A234)  and  (not A233) );
 a56601a <=( (not A236)  and  (not A235) );
 a56602a <=( a56601a  and  a56598a );
 a56605a <=( (not A299)  and  A298 );
 a56608a <=( A301  and  A300 );
 a56609a <=( a56608a  and  a56605a );
 a56610a <=( a56609a  and  a56602a );
 a56613a <=( (not A169)  and  A170 );
 a56616a <=( A167  and  (not A168) );
 a56617a <=( a56616a  and  a56613a );
 a56620a <=( A199  and  (not A166) );
 a56623a <=( A232  and  A200 );
 a56624a <=( a56623a  and  a56620a );
 a56625a <=( a56624a  and  a56617a );
 a56628a <=( (not A234)  and  (not A233) );
 a56631a <=( (not A236)  and  (not A235) );
 a56632a <=( a56631a  and  a56628a );
 a56635a <=( (not A299)  and  A298 );
 a56638a <=( A302  and  A300 );
 a56639a <=( a56638a  and  a56635a );
 a56640a <=( a56639a  and  a56632a );
 a56643a <=( (not A169)  and  A170 );
 a56646a <=( A167  and  (not A168) );
 a56647a <=( a56646a  and  a56643a );
 a56650a <=( A199  and  (not A166) );
 a56653a <=( A232  and  A200 );
 a56654a <=( a56653a  and  a56650a );
 a56655a <=( a56654a  and  a56647a );
 a56658a <=( (not A234)  and  (not A233) );
 a56661a <=( (not A236)  and  (not A235) );
 a56662a <=( a56661a  and  a56658a );
 a56665a <=( A299  and  (not A298) );
 a56668a <=( A301  and  A300 );
 a56669a <=( a56668a  and  a56665a );
 a56670a <=( a56669a  and  a56662a );
 a56673a <=( (not A169)  and  A170 );
 a56676a <=( A167  and  (not A168) );
 a56677a <=( a56676a  and  a56673a );
 a56680a <=( A199  and  (not A166) );
 a56683a <=( A232  and  A200 );
 a56684a <=( a56683a  and  a56680a );
 a56685a <=( a56684a  and  a56677a );
 a56688a <=( (not A234)  and  (not A233) );
 a56691a <=( (not A236)  and  (not A235) );
 a56692a <=( a56691a  and  a56688a );
 a56695a <=( A299  and  (not A298) );
 a56698a <=( A302  and  A300 );
 a56699a <=( a56698a  and  a56695a );
 a56700a <=( a56699a  and  a56692a );
 a56703a <=( (not A169)  and  A170 );
 a56706a <=( A167  and  (not A168) );
 a56707a <=( a56706a  and  a56703a );
 a56710a <=( A199  and  (not A166) );
 a56713a <=( A232  and  A200 );
 a56714a <=( a56713a  and  a56710a );
 a56715a <=( a56714a  and  a56707a );
 a56718a <=( (not A234)  and  (not A233) );
 a56721a <=( (not A236)  and  (not A235) );
 a56722a <=( a56721a  and  a56718a );
 a56725a <=( A266  and  (not A265) );
 a56728a <=( A268  and  A267 );
 a56729a <=( a56728a  and  a56725a );
 a56730a <=( a56729a  and  a56722a );
 a56733a <=( (not A169)  and  A170 );
 a56736a <=( A167  and  (not A168) );
 a56737a <=( a56736a  and  a56733a );
 a56740a <=( A199  and  (not A166) );
 a56743a <=( A232  and  A200 );
 a56744a <=( a56743a  and  a56740a );
 a56745a <=( a56744a  and  a56737a );
 a56748a <=( (not A234)  and  (not A233) );
 a56751a <=( (not A236)  and  (not A235) );
 a56752a <=( a56751a  and  a56748a );
 a56755a <=( A266  and  (not A265) );
 a56758a <=( A269  and  A267 );
 a56759a <=( a56758a  and  a56755a );
 a56760a <=( a56759a  and  a56752a );
 a56763a <=( (not A169)  and  A170 );
 a56766a <=( A167  and  (not A168) );
 a56767a <=( a56766a  and  a56763a );
 a56770a <=( A199  and  (not A166) );
 a56773a <=( A232  and  A200 );
 a56774a <=( a56773a  and  a56770a );
 a56775a <=( a56774a  and  a56767a );
 a56778a <=( (not A234)  and  (not A233) );
 a56781a <=( (not A236)  and  (not A235) );
 a56782a <=( a56781a  and  a56778a );
 a56785a <=( (not A266)  and  A265 );
 a56788a <=( A268  and  A267 );
 a56789a <=( a56788a  and  a56785a );
 a56790a <=( a56789a  and  a56782a );
 a56793a <=( (not A169)  and  A170 );
 a56796a <=( A167  and  (not A168) );
 a56797a <=( a56796a  and  a56793a );
 a56800a <=( A199  and  (not A166) );
 a56803a <=( A232  and  A200 );
 a56804a <=( a56803a  and  a56800a );
 a56805a <=( a56804a  and  a56797a );
 a56808a <=( (not A234)  and  (not A233) );
 a56811a <=( (not A236)  and  (not A235) );
 a56812a <=( a56811a  and  a56808a );
 a56815a <=( (not A266)  and  A265 );
 a56818a <=( A269  and  A267 );
 a56819a <=( a56818a  and  a56815a );
 a56820a <=( a56819a  and  a56812a );
 a56823a <=( (not A169)  and  A170 );
 a56826a <=( A167  and  (not A168) );
 a56827a <=( a56826a  and  a56823a );
 a56830a <=( (not A199)  and  (not A166) );
 a56833a <=( (not A232)  and  (not A200) );
 a56834a <=( a56833a  and  a56830a );
 a56835a <=( a56834a  and  a56827a );
 a56838a <=( A234  and  A233 );
 a56841a <=( A298  and  A235 );
 a56842a <=( a56841a  and  a56838a );
 a56845a <=( (not A300)  and  (not A299) );
 a56848a <=( (not A302)  and  (not A301) );
 a56849a <=( a56848a  and  a56845a );
 a56850a <=( a56849a  and  a56842a );
 a56853a <=( (not A169)  and  A170 );
 a56856a <=( A167  and  (not A168) );
 a56857a <=( a56856a  and  a56853a );
 a56860a <=( (not A199)  and  (not A166) );
 a56863a <=( (not A232)  and  (not A200) );
 a56864a <=( a56863a  and  a56860a );
 a56865a <=( a56864a  and  a56857a );
 a56868a <=( A234  and  A233 );
 a56871a <=( (not A298)  and  A235 );
 a56872a <=( a56871a  and  a56868a );
 a56875a <=( (not A300)  and  A299 );
 a56878a <=( (not A302)  and  (not A301) );
 a56879a <=( a56878a  and  a56875a );
 a56880a <=( a56879a  and  a56872a );
 a56883a <=( (not A169)  and  A170 );
 a56886a <=( A167  and  (not A168) );
 a56887a <=( a56886a  and  a56883a );
 a56890a <=( (not A199)  and  (not A166) );
 a56893a <=( (not A232)  and  (not A200) );
 a56894a <=( a56893a  and  a56890a );
 a56895a <=( a56894a  and  a56887a );
 a56898a <=( A234  and  A233 );
 a56901a <=( (not A265)  and  A235 );
 a56902a <=( a56901a  and  a56898a );
 a56905a <=( (not A267)  and  A266 );
 a56908a <=( (not A269)  and  (not A268) );
 a56909a <=( a56908a  and  a56905a );
 a56910a <=( a56909a  and  a56902a );
 a56913a <=( (not A169)  and  A170 );
 a56916a <=( A167  and  (not A168) );
 a56917a <=( a56916a  and  a56913a );
 a56920a <=( (not A199)  and  (not A166) );
 a56923a <=( (not A232)  and  (not A200) );
 a56924a <=( a56923a  and  a56920a );
 a56925a <=( a56924a  and  a56917a );
 a56928a <=( A234  and  A233 );
 a56931a <=( A265  and  A235 );
 a56932a <=( a56931a  and  a56928a );
 a56935a <=( (not A267)  and  (not A266) );
 a56938a <=( (not A269)  and  (not A268) );
 a56939a <=( a56938a  and  a56935a );
 a56940a <=( a56939a  and  a56932a );
 a56943a <=( (not A169)  and  A170 );
 a56946a <=( A167  and  (not A168) );
 a56947a <=( a56946a  and  a56943a );
 a56950a <=( (not A199)  and  (not A166) );
 a56953a <=( (not A232)  and  (not A200) );
 a56954a <=( a56953a  and  a56950a );
 a56955a <=( a56954a  and  a56947a );
 a56958a <=( A234  and  A233 );
 a56961a <=( A298  and  A236 );
 a56962a <=( a56961a  and  a56958a );
 a56965a <=( (not A300)  and  (not A299) );
 a56968a <=( (not A302)  and  (not A301) );
 a56969a <=( a56968a  and  a56965a );
 a56970a <=( a56969a  and  a56962a );
 a56973a <=( (not A169)  and  A170 );
 a56976a <=( A167  and  (not A168) );
 a56977a <=( a56976a  and  a56973a );
 a56980a <=( (not A199)  and  (not A166) );
 a56983a <=( (not A232)  and  (not A200) );
 a56984a <=( a56983a  and  a56980a );
 a56985a <=( a56984a  and  a56977a );
 a56988a <=( A234  and  A233 );
 a56991a <=( (not A298)  and  A236 );
 a56992a <=( a56991a  and  a56988a );
 a56995a <=( (not A300)  and  A299 );
 a56998a <=( (not A302)  and  (not A301) );
 a56999a <=( a56998a  and  a56995a );
 a57000a <=( a56999a  and  a56992a );
 a57003a <=( (not A169)  and  A170 );
 a57006a <=( A167  and  (not A168) );
 a57007a <=( a57006a  and  a57003a );
 a57010a <=( (not A199)  and  (not A166) );
 a57013a <=( (not A232)  and  (not A200) );
 a57014a <=( a57013a  and  a57010a );
 a57015a <=( a57014a  and  a57007a );
 a57018a <=( A234  and  A233 );
 a57021a <=( (not A265)  and  A236 );
 a57022a <=( a57021a  and  a57018a );
 a57025a <=( (not A267)  and  A266 );
 a57028a <=( (not A269)  and  (not A268) );
 a57029a <=( a57028a  and  a57025a );
 a57030a <=( a57029a  and  a57022a );
 a57033a <=( (not A169)  and  A170 );
 a57036a <=( A167  and  (not A168) );
 a57037a <=( a57036a  and  a57033a );
 a57040a <=( (not A199)  and  (not A166) );
 a57043a <=( (not A232)  and  (not A200) );
 a57044a <=( a57043a  and  a57040a );
 a57045a <=( a57044a  and  a57037a );
 a57048a <=( A234  and  A233 );
 a57051a <=( A265  and  A236 );
 a57052a <=( a57051a  and  a57048a );
 a57055a <=( (not A267)  and  (not A266) );
 a57058a <=( (not A269)  and  (not A268) );
 a57059a <=( a57058a  and  a57055a );
 a57060a <=( a57059a  and  a57052a );
 a57063a <=( (not A169)  and  A170 );
 a57066a <=( A167  and  (not A168) );
 a57067a <=( a57066a  and  a57063a );
 a57070a <=( (not A199)  and  (not A166) );
 a57073a <=( (not A232)  and  (not A200) );
 a57074a <=( a57073a  and  a57070a );
 a57075a <=( a57074a  and  a57067a );
 a57078a <=( (not A234)  and  A233 );
 a57081a <=( (not A236)  and  (not A235) );
 a57082a <=( a57081a  and  a57078a );
 a57085a <=( (not A299)  and  A298 );
 a57088a <=( A301  and  A300 );
 a57089a <=( a57088a  and  a57085a );
 a57090a <=( a57089a  and  a57082a );
 a57093a <=( (not A169)  and  A170 );
 a57096a <=( A167  and  (not A168) );
 a57097a <=( a57096a  and  a57093a );
 a57100a <=( (not A199)  and  (not A166) );
 a57103a <=( (not A232)  and  (not A200) );
 a57104a <=( a57103a  and  a57100a );
 a57105a <=( a57104a  and  a57097a );
 a57108a <=( (not A234)  and  A233 );
 a57111a <=( (not A236)  and  (not A235) );
 a57112a <=( a57111a  and  a57108a );
 a57115a <=( (not A299)  and  A298 );
 a57118a <=( A302  and  A300 );
 a57119a <=( a57118a  and  a57115a );
 a57120a <=( a57119a  and  a57112a );
 a57123a <=( (not A169)  and  A170 );
 a57126a <=( A167  and  (not A168) );
 a57127a <=( a57126a  and  a57123a );
 a57130a <=( (not A199)  and  (not A166) );
 a57133a <=( (not A232)  and  (not A200) );
 a57134a <=( a57133a  and  a57130a );
 a57135a <=( a57134a  and  a57127a );
 a57138a <=( (not A234)  and  A233 );
 a57141a <=( (not A236)  and  (not A235) );
 a57142a <=( a57141a  and  a57138a );
 a57145a <=( A299  and  (not A298) );
 a57148a <=( A301  and  A300 );
 a57149a <=( a57148a  and  a57145a );
 a57150a <=( a57149a  and  a57142a );
 a57153a <=( (not A169)  and  A170 );
 a57156a <=( A167  and  (not A168) );
 a57157a <=( a57156a  and  a57153a );
 a57160a <=( (not A199)  and  (not A166) );
 a57163a <=( (not A232)  and  (not A200) );
 a57164a <=( a57163a  and  a57160a );
 a57165a <=( a57164a  and  a57157a );
 a57168a <=( (not A234)  and  A233 );
 a57171a <=( (not A236)  and  (not A235) );
 a57172a <=( a57171a  and  a57168a );
 a57175a <=( A299  and  (not A298) );
 a57178a <=( A302  and  A300 );
 a57179a <=( a57178a  and  a57175a );
 a57180a <=( a57179a  and  a57172a );
 a57183a <=( (not A169)  and  A170 );
 a57186a <=( A167  and  (not A168) );
 a57187a <=( a57186a  and  a57183a );
 a57190a <=( (not A199)  and  (not A166) );
 a57193a <=( (not A232)  and  (not A200) );
 a57194a <=( a57193a  and  a57190a );
 a57195a <=( a57194a  and  a57187a );
 a57198a <=( (not A234)  and  A233 );
 a57201a <=( (not A236)  and  (not A235) );
 a57202a <=( a57201a  and  a57198a );
 a57205a <=( A266  and  (not A265) );
 a57208a <=( A268  and  A267 );
 a57209a <=( a57208a  and  a57205a );
 a57210a <=( a57209a  and  a57202a );
 a57213a <=( (not A169)  and  A170 );
 a57216a <=( A167  and  (not A168) );
 a57217a <=( a57216a  and  a57213a );
 a57220a <=( (not A199)  and  (not A166) );
 a57223a <=( (not A232)  and  (not A200) );
 a57224a <=( a57223a  and  a57220a );
 a57225a <=( a57224a  and  a57217a );
 a57228a <=( (not A234)  and  A233 );
 a57231a <=( (not A236)  and  (not A235) );
 a57232a <=( a57231a  and  a57228a );
 a57235a <=( A266  and  (not A265) );
 a57238a <=( A269  and  A267 );
 a57239a <=( a57238a  and  a57235a );
 a57240a <=( a57239a  and  a57232a );
 a57243a <=( (not A169)  and  A170 );
 a57246a <=( A167  and  (not A168) );
 a57247a <=( a57246a  and  a57243a );
 a57250a <=( (not A199)  and  (not A166) );
 a57253a <=( (not A232)  and  (not A200) );
 a57254a <=( a57253a  and  a57250a );
 a57255a <=( a57254a  and  a57247a );
 a57258a <=( (not A234)  and  A233 );
 a57261a <=( (not A236)  and  (not A235) );
 a57262a <=( a57261a  and  a57258a );
 a57265a <=( (not A266)  and  A265 );
 a57268a <=( A268  and  A267 );
 a57269a <=( a57268a  and  a57265a );
 a57270a <=( a57269a  and  a57262a );
 a57273a <=( (not A169)  and  A170 );
 a57276a <=( A167  and  (not A168) );
 a57277a <=( a57276a  and  a57273a );
 a57280a <=( (not A199)  and  (not A166) );
 a57283a <=( (not A232)  and  (not A200) );
 a57284a <=( a57283a  and  a57280a );
 a57285a <=( a57284a  and  a57277a );
 a57288a <=( (not A234)  and  A233 );
 a57291a <=( (not A236)  and  (not A235) );
 a57292a <=( a57291a  and  a57288a );
 a57295a <=( (not A266)  and  A265 );
 a57298a <=( A269  and  A267 );
 a57299a <=( a57298a  and  a57295a );
 a57300a <=( a57299a  and  a57292a );
 a57303a <=( (not A169)  and  A170 );
 a57306a <=( A167  and  (not A168) );
 a57307a <=( a57306a  and  a57303a );
 a57310a <=( (not A199)  and  (not A166) );
 a57313a <=( A232  and  (not A200) );
 a57314a <=( a57313a  and  a57310a );
 a57315a <=( a57314a  and  a57307a );
 a57318a <=( A234  and  (not A233) );
 a57321a <=( A298  and  A235 );
 a57322a <=( a57321a  and  a57318a );
 a57325a <=( (not A300)  and  (not A299) );
 a57328a <=( (not A302)  and  (not A301) );
 a57329a <=( a57328a  and  a57325a );
 a57330a <=( a57329a  and  a57322a );
 a57333a <=( (not A169)  and  A170 );
 a57336a <=( A167  and  (not A168) );
 a57337a <=( a57336a  and  a57333a );
 a57340a <=( (not A199)  and  (not A166) );
 a57343a <=( A232  and  (not A200) );
 a57344a <=( a57343a  and  a57340a );
 a57345a <=( a57344a  and  a57337a );
 a57348a <=( A234  and  (not A233) );
 a57351a <=( (not A298)  and  A235 );
 a57352a <=( a57351a  and  a57348a );
 a57355a <=( (not A300)  and  A299 );
 a57358a <=( (not A302)  and  (not A301) );
 a57359a <=( a57358a  and  a57355a );
 a57360a <=( a57359a  and  a57352a );
 a57363a <=( (not A169)  and  A170 );
 a57366a <=( A167  and  (not A168) );
 a57367a <=( a57366a  and  a57363a );
 a57370a <=( (not A199)  and  (not A166) );
 a57373a <=( A232  and  (not A200) );
 a57374a <=( a57373a  and  a57370a );
 a57375a <=( a57374a  and  a57367a );
 a57378a <=( A234  and  (not A233) );
 a57381a <=( (not A265)  and  A235 );
 a57382a <=( a57381a  and  a57378a );
 a57385a <=( (not A267)  and  A266 );
 a57388a <=( (not A269)  and  (not A268) );
 a57389a <=( a57388a  and  a57385a );
 a57390a <=( a57389a  and  a57382a );
 a57393a <=( (not A169)  and  A170 );
 a57396a <=( A167  and  (not A168) );
 a57397a <=( a57396a  and  a57393a );
 a57400a <=( (not A199)  and  (not A166) );
 a57403a <=( A232  and  (not A200) );
 a57404a <=( a57403a  and  a57400a );
 a57405a <=( a57404a  and  a57397a );
 a57408a <=( A234  and  (not A233) );
 a57411a <=( A265  and  A235 );
 a57412a <=( a57411a  and  a57408a );
 a57415a <=( (not A267)  and  (not A266) );
 a57418a <=( (not A269)  and  (not A268) );
 a57419a <=( a57418a  and  a57415a );
 a57420a <=( a57419a  and  a57412a );
 a57423a <=( (not A169)  and  A170 );
 a57426a <=( A167  and  (not A168) );
 a57427a <=( a57426a  and  a57423a );
 a57430a <=( (not A199)  and  (not A166) );
 a57433a <=( A232  and  (not A200) );
 a57434a <=( a57433a  and  a57430a );
 a57435a <=( a57434a  and  a57427a );
 a57438a <=( A234  and  (not A233) );
 a57441a <=( A298  and  A236 );
 a57442a <=( a57441a  and  a57438a );
 a57445a <=( (not A300)  and  (not A299) );
 a57448a <=( (not A302)  and  (not A301) );
 a57449a <=( a57448a  and  a57445a );
 a57450a <=( a57449a  and  a57442a );
 a57453a <=( (not A169)  and  A170 );
 a57456a <=( A167  and  (not A168) );
 a57457a <=( a57456a  and  a57453a );
 a57460a <=( (not A199)  and  (not A166) );
 a57463a <=( A232  and  (not A200) );
 a57464a <=( a57463a  and  a57460a );
 a57465a <=( a57464a  and  a57457a );
 a57468a <=( A234  and  (not A233) );
 a57471a <=( (not A298)  and  A236 );
 a57472a <=( a57471a  and  a57468a );
 a57475a <=( (not A300)  and  A299 );
 a57478a <=( (not A302)  and  (not A301) );
 a57479a <=( a57478a  and  a57475a );
 a57480a <=( a57479a  and  a57472a );
 a57483a <=( (not A169)  and  A170 );
 a57486a <=( A167  and  (not A168) );
 a57487a <=( a57486a  and  a57483a );
 a57490a <=( (not A199)  and  (not A166) );
 a57493a <=( A232  and  (not A200) );
 a57494a <=( a57493a  and  a57490a );
 a57495a <=( a57494a  and  a57487a );
 a57498a <=( A234  and  (not A233) );
 a57501a <=( (not A265)  and  A236 );
 a57502a <=( a57501a  and  a57498a );
 a57505a <=( (not A267)  and  A266 );
 a57508a <=( (not A269)  and  (not A268) );
 a57509a <=( a57508a  and  a57505a );
 a57510a <=( a57509a  and  a57502a );
 a57513a <=( (not A169)  and  A170 );
 a57516a <=( A167  and  (not A168) );
 a57517a <=( a57516a  and  a57513a );
 a57520a <=( (not A199)  and  (not A166) );
 a57523a <=( A232  and  (not A200) );
 a57524a <=( a57523a  and  a57520a );
 a57525a <=( a57524a  and  a57517a );
 a57528a <=( A234  and  (not A233) );
 a57531a <=( A265  and  A236 );
 a57532a <=( a57531a  and  a57528a );
 a57535a <=( (not A267)  and  (not A266) );
 a57538a <=( (not A269)  and  (not A268) );
 a57539a <=( a57538a  and  a57535a );
 a57540a <=( a57539a  and  a57532a );
 a57543a <=( (not A169)  and  A170 );
 a57546a <=( A167  and  (not A168) );
 a57547a <=( a57546a  and  a57543a );
 a57550a <=( (not A199)  and  (not A166) );
 a57553a <=( A232  and  (not A200) );
 a57554a <=( a57553a  and  a57550a );
 a57555a <=( a57554a  and  a57547a );
 a57558a <=( (not A234)  and  (not A233) );
 a57561a <=( (not A236)  and  (not A235) );
 a57562a <=( a57561a  and  a57558a );
 a57565a <=( (not A299)  and  A298 );
 a57568a <=( A301  and  A300 );
 a57569a <=( a57568a  and  a57565a );
 a57570a <=( a57569a  and  a57562a );
 a57573a <=( (not A169)  and  A170 );
 a57576a <=( A167  and  (not A168) );
 a57577a <=( a57576a  and  a57573a );
 a57580a <=( (not A199)  and  (not A166) );
 a57583a <=( A232  and  (not A200) );
 a57584a <=( a57583a  and  a57580a );
 a57585a <=( a57584a  and  a57577a );
 a57588a <=( (not A234)  and  (not A233) );
 a57591a <=( (not A236)  and  (not A235) );
 a57592a <=( a57591a  and  a57588a );
 a57595a <=( (not A299)  and  A298 );
 a57598a <=( A302  and  A300 );
 a57599a <=( a57598a  and  a57595a );
 a57600a <=( a57599a  and  a57592a );
 a57603a <=( (not A169)  and  A170 );
 a57606a <=( A167  and  (not A168) );
 a57607a <=( a57606a  and  a57603a );
 a57610a <=( (not A199)  and  (not A166) );
 a57613a <=( A232  and  (not A200) );
 a57614a <=( a57613a  and  a57610a );
 a57615a <=( a57614a  and  a57607a );
 a57618a <=( (not A234)  and  (not A233) );
 a57621a <=( (not A236)  and  (not A235) );
 a57622a <=( a57621a  and  a57618a );
 a57625a <=( A299  and  (not A298) );
 a57628a <=( A301  and  A300 );
 a57629a <=( a57628a  and  a57625a );
 a57630a <=( a57629a  and  a57622a );
 a57633a <=( (not A169)  and  A170 );
 a57636a <=( A167  and  (not A168) );
 a57637a <=( a57636a  and  a57633a );
 a57640a <=( (not A199)  and  (not A166) );
 a57643a <=( A232  and  (not A200) );
 a57644a <=( a57643a  and  a57640a );
 a57645a <=( a57644a  and  a57637a );
 a57648a <=( (not A234)  and  (not A233) );
 a57651a <=( (not A236)  and  (not A235) );
 a57652a <=( a57651a  and  a57648a );
 a57655a <=( A299  and  (not A298) );
 a57658a <=( A302  and  A300 );
 a57659a <=( a57658a  and  a57655a );
 a57660a <=( a57659a  and  a57652a );
 a57663a <=( (not A169)  and  A170 );
 a57666a <=( A167  and  (not A168) );
 a57667a <=( a57666a  and  a57663a );
 a57670a <=( (not A199)  and  (not A166) );
 a57673a <=( A232  and  (not A200) );
 a57674a <=( a57673a  and  a57670a );
 a57675a <=( a57674a  and  a57667a );
 a57678a <=( (not A234)  and  (not A233) );
 a57681a <=( (not A236)  and  (not A235) );
 a57682a <=( a57681a  and  a57678a );
 a57685a <=( A266  and  (not A265) );
 a57688a <=( A268  and  A267 );
 a57689a <=( a57688a  and  a57685a );
 a57690a <=( a57689a  and  a57682a );
 a57693a <=( (not A169)  and  A170 );
 a57696a <=( A167  and  (not A168) );
 a57697a <=( a57696a  and  a57693a );
 a57700a <=( (not A199)  and  (not A166) );
 a57703a <=( A232  and  (not A200) );
 a57704a <=( a57703a  and  a57700a );
 a57705a <=( a57704a  and  a57697a );
 a57708a <=( (not A234)  and  (not A233) );
 a57711a <=( (not A236)  and  (not A235) );
 a57712a <=( a57711a  and  a57708a );
 a57715a <=( A266  and  (not A265) );
 a57718a <=( A269  and  A267 );
 a57719a <=( a57718a  and  a57715a );
 a57720a <=( a57719a  and  a57712a );
 a57723a <=( (not A169)  and  A170 );
 a57726a <=( A167  and  (not A168) );
 a57727a <=( a57726a  and  a57723a );
 a57730a <=( (not A199)  and  (not A166) );
 a57733a <=( A232  and  (not A200) );
 a57734a <=( a57733a  and  a57730a );
 a57735a <=( a57734a  and  a57727a );
 a57738a <=( (not A234)  and  (not A233) );
 a57741a <=( (not A236)  and  (not A235) );
 a57742a <=( a57741a  and  a57738a );
 a57745a <=( (not A266)  and  A265 );
 a57748a <=( A268  and  A267 );
 a57749a <=( a57748a  and  a57745a );
 a57750a <=( a57749a  and  a57742a );
 a57753a <=( (not A169)  and  A170 );
 a57756a <=( A167  and  (not A168) );
 a57757a <=( a57756a  and  a57753a );
 a57760a <=( (not A199)  and  (not A166) );
 a57763a <=( A232  and  (not A200) );
 a57764a <=( a57763a  and  a57760a );
 a57765a <=( a57764a  and  a57757a );
 a57768a <=( (not A234)  and  (not A233) );
 a57771a <=( (not A236)  and  (not A235) );
 a57772a <=( a57771a  and  a57768a );
 a57775a <=( (not A266)  and  A265 );
 a57778a <=( A269  and  A267 );
 a57779a <=( a57778a  and  a57775a );
 a57780a <=( a57779a  and  a57772a );
 a57783a <=( (not A169)  and  A170 );
 a57786a <=( (not A167)  and  (not A168) );
 a57787a <=( a57786a  and  a57783a );
 a57790a <=( A201  and  A166 );
 a57793a <=( (not A203)  and  (not A202) );
 a57794a <=( a57793a  and  a57790a );
 a57795a <=( a57794a  and  a57787a );
 a57798a <=( A233  and  (not A232) );
 a57801a <=( A235  and  A234 );
 a57802a <=( a57801a  and  a57798a );
 a57805a <=( (not A299)  and  A298 );
 a57808a <=( A301  and  A300 );
 a57809a <=( a57808a  and  a57805a );
 a57810a <=( a57809a  and  a57802a );
 a57813a <=( (not A169)  and  A170 );
 a57816a <=( (not A167)  and  (not A168) );
 a57817a <=( a57816a  and  a57813a );
 a57820a <=( A201  and  A166 );
 a57823a <=( (not A203)  and  (not A202) );
 a57824a <=( a57823a  and  a57820a );
 a57825a <=( a57824a  and  a57817a );
 a57828a <=( A233  and  (not A232) );
 a57831a <=( A235  and  A234 );
 a57832a <=( a57831a  and  a57828a );
 a57835a <=( (not A299)  and  A298 );
 a57838a <=( A302  and  A300 );
 a57839a <=( a57838a  and  a57835a );
 a57840a <=( a57839a  and  a57832a );
 a57843a <=( (not A169)  and  A170 );
 a57846a <=( (not A167)  and  (not A168) );
 a57847a <=( a57846a  and  a57843a );
 a57850a <=( A201  and  A166 );
 a57853a <=( (not A203)  and  (not A202) );
 a57854a <=( a57853a  and  a57850a );
 a57855a <=( a57854a  and  a57847a );
 a57858a <=( A233  and  (not A232) );
 a57861a <=( A235  and  A234 );
 a57862a <=( a57861a  and  a57858a );
 a57865a <=( A299  and  (not A298) );
 a57868a <=( A301  and  A300 );
 a57869a <=( a57868a  and  a57865a );
 a57870a <=( a57869a  and  a57862a );
 a57873a <=( (not A169)  and  A170 );
 a57876a <=( (not A167)  and  (not A168) );
 a57877a <=( a57876a  and  a57873a );
 a57880a <=( A201  and  A166 );
 a57883a <=( (not A203)  and  (not A202) );
 a57884a <=( a57883a  and  a57880a );
 a57885a <=( a57884a  and  a57877a );
 a57888a <=( A233  and  (not A232) );
 a57891a <=( A235  and  A234 );
 a57892a <=( a57891a  and  a57888a );
 a57895a <=( A299  and  (not A298) );
 a57898a <=( A302  and  A300 );
 a57899a <=( a57898a  and  a57895a );
 a57900a <=( a57899a  and  a57892a );
 a57903a <=( (not A169)  and  A170 );
 a57906a <=( (not A167)  and  (not A168) );
 a57907a <=( a57906a  and  a57903a );
 a57910a <=( A201  and  A166 );
 a57913a <=( (not A203)  and  (not A202) );
 a57914a <=( a57913a  and  a57910a );
 a57915a <=( a57914a  and  a57907a );
 a57918a <=( A233  and  (not A232) );
 a57921a <=( A235  and  A234 );
 a57922a <=( a57921a  and  a57918a );
 a57925a <=( A266  and  (not A265) );
 a57928a <=( A268  and  A267 );
 a57929a <=( a57928a  and  a57925a );
 a57930a <=( a57929a  and  a57922a );
 a57933a <=( (not A169)  and  A170 );
 a57936a <=( (not A167)  and  (not A168) );
 a57937a <=( a57936a  and  a57933a );
 a57940a <=( A201  and  A166 );
 a57943a <=( (not A203)  and  (not A202) );
 a57944a <=( a57943a  and  a57940a );
 a57945a <=( a57944a  and  a57937a );
 a57948a <=( A233  and  (not A232) );
 a57951a <=( A235  and  A234 );
 a57952a <=( a57951a  and  a57948a );
 a57955a <=( A266  and  (not A265) );
 a57958a <=( A269  and  A267 );
 a57959a <=( a57958a  and  a57955a );
 a57960a <=( a57959a  and  a57952a );
 a57963a <=( (not A169)  and  A170 );
 a57966a <=( (not A167)  and  (not A168) );
 a57967a <=( a57966a  and  a57963a );
 a57970a <=( A201  and  A166 );
 a57973a <=( (not A203)  and  (not A202) );
 a57974a <=( a57973a  and  a57970a );
 a57975a <=( a57974a  and  a57967a );
 a57978a <=( A233  and  (not A232) );
 a57981a <=( A235  and  A234 );
 a57982a <=( a57981a  and  a57978a );
 a57985a <=( (not A266)  and  A265 );
 a57988a <=( A268  and  A267 );
 a57989a <=( a57988a  and  a57985a );
 a57990a <=( a57989a  and  a57982a );
 a57993a <=( (not A169)  and  A170 );
 a57996a <=( (not A167)  and  (not A168) );
 a57997a <=( a57996a  and  a57993a );
 a58000a <=( A201  and  A166 );
 a58003a <=( (not A203)  and  (not A202) );
 a58004a <=( a58003a  and  a58000a );
 a58005a <=( a58004a  and  a57997a );
 a58008a <=( A233  and  (not A232) );
 a58011a <=( A235  and  A234 );
 a58012a <=( a58011a  and  a58008a );
 a58015a <=( (not A266)  and  A265 );
 a58018a <=( A269  and  A267 );
 a58019a <=( a58018a  and  a58015a );
 a58020a <=( a58019a  and  a58012a );
 a58023a <=( (not A169)  and  A170 );
 a58026a <=( (not A167)  and  (not A168) );
 a58027a <=( a58026a  and  a58023a );
 a58030a <=( A201  and  A166 );
 a58033a <=( (not A203)  and  (not A202) );
 a58034a <=( a58033a  and  a58030a );
 a58035a <=( a58034a  and  a58027a );
 a58038a <=( A233  and  (not A232) );
 a58041a <=( A236  and  A234 );
 a58042a <=( a58041a  and  a58038a );
 a58045a <=( (not A299)  and  A298 );
 a58048a <=( A301  and  A300 );
 a58049a <=( a58048a  and  a58045a );
 a58050a <=( a58049a  and  a58042a );
 a58053a <=( (not A169)  and  A170 );
 a58056a <=( (not A167)  and  (not A168) );
 a58057a <=( a58056a  and  a58053a );
 a58060a <=( A201  and  A166 );
 a58063a <=( (not A203)  and  (not A202) );
 a58064a <=( a58063a  and  a58060a );
 a58065a <=( a58064a  and  a58057a );
 a58068a <=( A233  and  (not A232) );
 a58071a <=( A236  and  A234 );
 a58072a <=( a58071a  and  a58068a );
 a58075a <=( (not A299)  and  A298 );
 a58078a <=( A302  and  A300 );
 a58079a <=( a58078a  and  a58075a );
 a58080a <=( a58079a  and  a58072a );
 a58083a <=( (not A169)  and  A170 );
 a58086a <=( (not A167)  and  (not A168) );
 a58087a <=( a58086a  and  a58083a );
 a58090a <=( A201  and  A166 );
 a58093a <=( (not A203)  and  (not A202) );
 a58094a <=( a58093a  and  a58090a );
 a58095a <=( a58094a  and  a58087a );
 a58098a <=( A233  and  (not A232) );
 a58101a <=( A236  and  A234 );
 a58102a <=( a58101a  and  a58098a );
 a58105a <=( A299  and  (not A298) );
 a58108a <=( A301  and  A300 );
 a58109a <=( a58108a  and  a58105a );
 a58110a <=( a58109a  and  a58102a );
 a58113a <=( (not A169)  and  A170 );
 a58116a <=( (not A167)  and  (not A168) );
 a58117a <=( a58116a  and  a58113a );
 a58120a <=( A201  and  A166 );
 a58123a <=( (not A203)  and  (not A202) );
 a58124a <=( a58123a  and  a58120a );
 a58125a <=( a58124a  and  a58117a );
 a58128a <=( A233  and  (not A232) );
 a58131a <=( A236  and  A234 );
 a58132a <=( a58131a  and  a58128a );
 a58135a <=( A299  and  (not A298) );
 a58138a <=( A302  and  A300 );
 a58139a <=( a58138a  and  a58135a );
 a58140a <=( a58139a  and  a58132a );
 a58143a <=( (not A169)  and  A170 );
 a58146a <=( (not A167)  and  (not A168) );
 a58147a <=( a58146a  and  a58143a );
 a58150a <=( A201  and  A166 );
 a58153a <=( (not A203)  and  (not A202) );
 a58154a <=( a58153a  and  a58150a );
 a58155a <=( a58154a  and  a58147a );
 a58158a <=( A233  and  (not A232) );
 a58161a <=( A236  and  A234 );
 a58162a <=( a58161a  and  a58158a );
 a58165a <=( A266  and  (not A265) );
 a58168a <=( A268  and  A267 );
 a58169a <=( a58168a  and  a58165a );
 a58170a <=( a58169a  and  a58162a );
 a58173a <=( (not A169)  and  A170 );
 a58176a <=( (not A167)  and  (not A168) );
 a58177a <=( a58176a  and  a58173a );
 a58180a <=( A201  and  A166 );
 a58183a <=( (not A203)  and  (not A202) );
 a58184a <=( a58183a  and  a58180a );
 a58185a <=( a58184a  and  a58177a );
 a58188a <=( A233  and  (not A232) );
 a58191a <=( A236  and  A234 );
 a58192a <=( a58191a  and  a58188a );
 a58195a <=( A266  and  (not A265) );
 a58198a <=( A269  and  A267 );
 a58199a <=( a58198a  and  a58195a );
 a58200a <=( a58199a  and  a58192a );
 a58203a <=( (not A169)  and  A170 );
 a58206a <=( (not A167)  and  (not A168) );
 a58207a <=( a58206a  and  a58203a );
 a58210a <=( A201  and  A166 );
 a58213a <=( (not A203)  and  (not A202) );
 a58214a <=( a58213a  and  a58210a );
 a58215a <=( a58214a  and  a58207a );
 a58218a <=( A233  and  (not A232) );
 a58221a <=( A236  and  A234 );
 a58222a <=( a58221a  and  a58218a );
 a58225a <=( (not A266)  and  A265 );
 a58228a <=( A268  and  A267 );
 a58229a <=( a58228a  and  a58225a );
 a58230a <=( a58229a  and  a58222a );
 a58233a <=( (not A169)  and  A170 );
 a58236a <=( (not A167)  and  (not A168) );
 a58237a <=( a58236a  and  a58233a );
 a58240a <=( A201  and  A166 );
 a58243a <=( (not A203)  and  (not A202) );
 a58244a <=( a58243a  and  a58240a );
 a58245a <=( a58244a  and  a58237a );
 a58248a <=( A233  and  (not A232) );
 a58251a <=( A236  and  A234 );
 a58252a <=( a58251a  and  a58248a );
 a58255a <=( (not A266)  and  A265 );
 a58258a <=( A269  and  A267 );
 a58259a <=( a58258a  and  a58255a );
 a58260a <=( a58259a  and  a58252a );
 a58263a <=( (not A169)  and  A170 );
 a58266a <=( (not A167)  and  (not A168) );
 a58267a <=( a58266a  and  a58263a );
 a58270a <=( A201  and  A166 );
 a58273a <=( (not A203)  and  (not A202) );
 a58274a <=( a58273a  and  a58270a );
 a58275a <=( a58274a  and  a58267a );
 a58278a <=( (not A233)  and  A232 );
 a58281a <=( A235  and  A234 );
 a58282a <=( a58281a  and  a58278a );
 a58285a <=( (not A299)  and  A298 );
 a58288a <=( A301  and  A300 );
 a58289a <=( a58288a  and  a58285a );
 a58290a <=( a58289a  and  a58282a );
 a58293a <=( (not A169)  and  A170 );
 a58296a <=( (not A167)  and  (not A168) );
 a58297a <=( a58296a  and  a58293a );
 a58300a <=( A201  and  A166 );
 a58303a <=( (not A203)  and  (not A202) );
 a58304a <=( a58303a  and  a58300a );
 a58305a <=( a58304a  and  a58297a );
 a58308a <=( (not A233)  and  A232 );
 a58311a <=( A235  and  A234 );
 a58312a <=( a58311a  and  a58308a );
 a58315a <=( (not A299)  and  A298 );
 a58318a <=( A302  and  A300 );
 a58319a <=( a58318a  and  a58315a );
 a58320a <=( a58319a  and  a58312a );
 a58323a <=( (not A169)  and  A170 );
 a58326a <=( (not A167)  and  (not A168) );
 a58327a <=( a58326a  and  a58323a );
 a58330a <=( A201  and  A166 );
 a58333a <=( (not A203)  and  (not A202) );
 a58334a <=( a58333a  and  a58330a );
 a58335a <=( a58334a  and  a58327a );
 a58338a <=( (not A233)  and  A232 );
 a58341a <=( A235  and  A234 );
 a58342a <=( a58341a  and  a58338a );
 a58345a <=( A299  and  (not A298) );
 a58348a <=( A301  and  A300 );
 a58349a <=( a58348a  and  a58345a );
 a58350a <=( a58349a  and  a58342a );
 a58353a <=( (not A169)  and  A170 );
 a58356a <=( (not A167)  and  (not A168) );
 a58357a <=( a58356a  and  a58353a );
 a58360a <=( A201  and  A166 );
 a58363a <=( (not A203)  and  (not A202) );
 a58364a <=( a58363a  and  a58360a );
 a58365a <=( a58364a  and  a58357a );
 a58368a <=( (not A233)  and  A232 );
 a58371a <=( A235  and  A234 );
 a58372a <=( a58371a  and  a58368a );
 a58375a <=( A299  and  (not A298) );
 a58378a <=( A302  and  A300 );
 a58379a <=( a58378a  and  a58375a );
 a58380a <=( a58379a  and  a58372a );
 a58383a <=( (not A169)  and  A170 );
 a58386a <=( (not A167)  and  (not A168) );
 a58387a <=( a58386a  and  a58383a );
 a58390a <=( A201  and  A166 );
 a58393a <=( (not A203)  and  (not A202) );
 a58394a <=( a58393a  and  a58390a );
 a58395a <=( a58394a  and  a58387a );
 a58398a <=( (not A233)  and  A232 );
 a58401a <=( A235  and  A234 );
 a58402a <=( a58401a  and  a58398a );
 a58405a <=( A266  and  (not A265) );
 a58408a <=( A268  and  A267 );
 a58409a <=( a58408a  and  a58405a );
 a58410a <=( a58409a  and  a58402a );
 a58413a <=( (not A169)  and  A170 );
 a58416a <=( (not A167)  and  (not A168) );
 a58417a <=( a58416a  and  a58413a );
 a58420a <=( A201  and  A166 );
 a58423a <=( (not A203)  and  (not A202) );
 a58424a <=( a58423a  and  a58420a );
 a58425a <=( a58424a  and  a58417a );
 a58428a <=( (not A233)  and  A232 );
 a58431a <=( A235  and  A234 );
 a58432a <=( a58431a  and  a58428a );
 a58435a <=( A266  and  (not A265) );
 a58438a <=( A269  and  A267 );
 a58439a <=( a58438a  and  a58435a );
 a58440a <=( a58439a  and  a58432a );
 a58443a <=( (not A169)  and  A170 );
 a58446a <=( (not A167)  and  (not A168) );
 a58447a <=( a58446a  and  a58443a );
 a58450a <=( A201  and  A166 );
 a58453a <=( (not A203)  and  (not A202) );
 a58454a <=( a58453a  and  a58450a );
 a58455a <=( a58454a  and  a58447a );
 a58458a <=( (not A233)  and  A232 );
 a58461a <=( A235  and  A234 );
 a58462a <=( a58461a  and  a58458a );
 a58465a <=( (not A266)  and  A265 );
 a58468a <=( A268  and  A267 );
 a58469a <=( a58468a  and  a58465a );
 a58470a <=( a58469a  and  a58462a );
 a58473a <=( (not A169)  and  A170 );
 a58476a <=( (not A167)  and  (not A168) );
 a58477a <=( a58476a  and  a58473a );
 a58480a <=( A201  and  A166 );
 a58483a <=( (not A203)  and  (not A202) );
 a58484a <=( a58483a  and  a58480a );
 a58485a <=( a58484a  and  a58477a );
 a58488a <=( (not A233)  and  A232 );
 a58491a <=( A235  and  A234 );
 a58492a <=( a58491a  and  a58488a );
 a58495a <=( (not A266)  and  A265 );
 a58498a <=( A269  and  A267 );
 a58499a <=( a58498a  and  a58495a );
 a58500a <=( a58499a  and  a58492a );
 a58503a <=( (not A169)  and  A170 );
 a58506a <=( (not A167)  and  (not A168) );
 a58507a <=( a58506a  and  a58503a );
 a58510a <=( A201  and  A166 );
 a58513a <=( (not A203)  and  (not A202) );
 a58514a <=( a58513a  and  a58510a );
 a58515a <=( a58514a  and  a58507a );
 a58518a <=( (not A233)  and  A232 );
 a58521a <=( A236  and  A234 );
 a58522a <=( a58521a  and  a58518a );
 a58525a <=( (not A299)  and  A298 );
 a58528a <=( A301  and  A300 );
 a58529a <=( a58528a  and  a58525a );
 a58530a <=( a58529a  and  a58522a );
 a58533a <=( (not A169)  and  A170 );
 a58536a <=( (not A167)  and  (not A168) );
 a58537a <=( a58536a  and  a58533a );
 a58540a <=( A201  and  A166 );
 a58543a <=( (not A203)  and  (not A202) );
 a58544a <=( a58543a  and  a58540a );
 a58545a <=( a58544a  and  a58537a );
 a58548a <=( (not A233)  and  A232 );
 a58551a <=( A236  and  A234 );
 a58552a <=( a58551a  and  a58548a );
 a58555a <=( (not A299)  and  A298 );
 a58558a <=( A302  and  A300 );
 a58559a <=( a58558a  and  a58555a );
 a58560a <=( a58559a  and  a58552a );
 a58563a <=( (not A169)  and  A170 );
 a58566a <=( (not A167)  and  (not A168) );
 a58567a <=( a58566a  and  a58563a );
 a58570a <=( A201  and  A166 );
 a58573a <=( (not A203)  and  (not A202) );
 a58574a <=( a58573a  and  a58570a );
 a58575a <=( a58574a  and  a58567a );
 a58578a <=( (not A233)  and  A232 );
 a58581a <=( A236  and  A234 );
 a58582a <=( a58581a  and  a58578a );
 a58585a <=( A299  and  (not A298) );
 a58588a <=( A301  and  A300 );
 a58589a <=( a58588a  and  a58585a );
 a58590a <=( a58589a  and  a58582a );
 a58593a <=( (not A169)  and  A170 );
 a58596a <=( (not A167)  and  (not A168) );
 a58597a <=( a58596a  and  a58593a );
 a58600a <=( A201  and  A166 );
 a58603a <=( (not A203)  and  (not A202) );
 a58604a <=( a58603a  and  a58600a );
 a58605a <=( a58604a  and  a58597a );
 a58608a <=( (not A233)  and  A232 );
 a58611a <=( A236  and  A234 );
 a58612a <=( a58611a  and  a58608a );
 a58615a <=( A299  and  (not A298) );
 a58618a <=( A302  and  A300 );
 a58619a <=( a58618a  and  a58615a );
 a58620a <=( a58619a  and  a58612a );
 a58623a <=( (not A169)  and  A170 );
 a58626a <=( (not A167)  and  (not A168) );
 a58627a <=( a58626a  and  a58623a );
 a58630a <=( A201  and  A166 );
 a58633a <=( (not A203)  and  (not A202) );
 a58634a <=( a58633a  and  a58630a );
 a58635a <=( a58634a  and  a58627a );
 a58638a <=( (not A233)  and  A232 );
 a58641a <=( A236  and  A234 );
 a58642a <=( a58641a  and  a58638a );
 a58645a <=( A266  and  (not A265) );
 a58648a <=( A268  and  A267 );
 a58649a <=( a58648a  and  a58645a );
 a58650a <=( a58649a  and  a58642a );
 a58653a <=( (not A169)  and  A170 );
 a58656a <=( (not A167)  and  (not A168) );
 a58657a <=( a58656a  and  a58653a );
 a58660a <=( A201  and  A166 );
 a58663a <=( (not A203)  and  (not A202) );
 a58664a <=( a58663a  and  a58660a );
 a58665a <=( a58664a  and  a58657a );
 a58668a <=( (not A233)  and  A232 );
 a58671a <=( A236  and  A234 );
 a58672a <=( a58671a  and  a58668a );
 a58675a <=( A266  and  (not A265) );
 a58678a <=( A269  and  A267 );
 a58679a <=( a58678a  and  a58675a );
 a58680a <=( a58679a  and  a58672a );
 a58683a <=( (not A169)  and  A170 );
 a58686a <=( (not A167)  and  (not A168) );
 a58687a <=( a58686a  and  a58683a );
 a58690a <=( A201  and  A166 );
 a58693a <=( (not A203)  and  (not A202) );
 a58694a <=( a58693a  and  a58690a );
 a58695a <=( a58694a  and  a58687a );
 a58698a <=( (not A233)  and  A232 );
 a58701a <=( A236  and  A234 );
 a58702a <=( a58701a  and  a58698a );
 a58705a <=( (not A266)  and  A265 );
 a58708a <=( A268  and  A267 );
 a58709a <=( a58708a  and  a58705a );
 a58710a <=( a58709a  and  a58702a );
 a58713a <=( (not A169)  and  A170 );
 a58716a <=( (not A167)  and  (not A168) );
 a58717a <=( a58716a  and  a58713a );
 a58720a <=( A201  and  A166 );
 a58723a <=( (not A203)  and  (not A202) );
 a58724a <=( a58723a  and  a58720a );
 a58725a <=( a58724a  and  a58717a );
 a58728a <=( (not A233)  and  A232 );
 a58731a <=( A236  and  A234 );
 a58732a <=( a58731a  and  a58728a );
 a58735a <=( (not A266)  and  A265 );
 a58738a <=( A269  and  A267 );
 a58739a <=( a58738a  and  a58735a );
 a58740a <=( a58739a  and  a58732a );
 a58743a <=( (not A169)  and  A170 );
 a58746a <=( (not A167)  and  (not A168) );
 a58747a <=( a58746a  and  a58743a );
 a58750a <=( (not A201)  and  A166 );
 a58753a <=( (not A232)  and  A202 );
 a58754a <=( a58753a  and  a58750a );
 a58755a <=( a58754a  and  a58747a );
 a58758a <=( A234  and  A233 );
 a58761a <=( A298  and  A235 );
 a58762a <=( a58761a  and  a58758a );
 a58765a <=( (not A300)  and  (not A299) );
 a58768a <=( (not A302)  and  (not A301) );
 a58769a <=( a58768a  and  a58765a );
 a58770a <=( a58769a  and  a58762a );
 a58773a <=( (not A169)  and  A170 );
 a58776a <=( (not A167)  and  (not A168) );
 a58777a <=( a58776a  and  a58773a );
 a58780a <=( (not A201)  and  A166 );
 a58783a <=( (not A232)  and  A202 );
 a58784a <=( a58783a  and  a58780a );
 a58785a <=( a58784a  and  a58777a );
 a58788a <=( A234  and  A233 );
 a58791a <=( (not A298)  and  A235 );
 a58792a <=( a58791a  and  a58788a );
 a58795a <=( (not A300)  and  A299 );
 a58798a <=( (not A302)  and  (not A301) );
 a58799a <=( a58798a  and  a58795a );
 a58800a <=( a58799a  and  a58792a );
 a58803a <=( (not A169)  and  A170 );
 a58806a <=( (not A167)  and  (not A168) );
 a58807a <=( a58806a  and  a58803a );
 a58810a <=( (not A201)  and  A166 );
 a58813a <=( (not A232)  and  A202 );
 a58814a <=( a58813a  and  a58810a );
 a58815a <=( a58814a  and  a58807a );
 a58818a <=( A234  and  A233 );
 a58821a <=( (not A265)  and  A235 );
 a58822a <=( a58821a  and  a58818a );
 a58825a <=( (not A267)  and  A266 );
 a58828a <=( (not A269)  and  (not A268) );
 a58829a <=( a58828a  and  a58825a );
 a58830a <=( a58829a  and  a58822a );
 a58833a <=( (not A169)  and  A170 );
 a58836a <=( (not A167)  and  (not A168) );
 a58837a <=( a58836a  and  a58833a );
 a58840a <=( (not A201)  and  A166 );
 a58843a <=( (not A232)  and  A202 );
 a58844a <=( a58843a  and  a58840a );
 a58845a <=( a58844a  and  a58837a );
 a58848a <=( A234  and  A233 );
 a58851a <=( A265  and  A235 );
 a58852a <=( a58851a  and  a58848a );
 a58855a <=( (not A267)  and  (not A266) );
 a58858a <=( (not A269)  and  (not A268) );
 a58859a <=( a58858a  and  a58855a );
 a58860a <=( a58859a  and  a58852a );
 a58863a <=( (not A169)  and  A170 );
 a58866a <=( (not A167)  and  (not A168) );
 a58867a <=( a58866a  and  a58863a );
 a58870a <=( (not A201)  and  A166 );
 a58873a <=( (not A232)  and  A202 );
 a58874a <=( a58873a  and  a58870a );
 a58875a <=( a58874a  and  a58867a );
 a58878a <=( A234  and  A233 );
 a58881a <=( A298  and  A236 );
 a58882a <=( a58881a  and  a58878a );
 a58885a <=( (not A300)  and  (not A299) );
 a58888a <=( (not A302)  and  (not A301) );
 a58889a <=( a58888a  and  a58885a );
 a58890a <=( a58889a  and  a58882a );
 a58893a <=( (not A169)  and  A170 );
 a58896a <=( (not A167)  and  (not A168) );
 a58897a <=( a58896a  and  a58893a );
 a58900a <=( (not A201)  and  A166 );
 a58903a <=( (not A232)  and  A202 );
 a58904a <=( a58903a  and  a58900a );
 a58905a <=( a58904a  and  a58897a );
 a58908a <=( A234  and  A233 );
 a58911a <=( (not A298)  and  A236 );
 a58912a <=( a58911a  and  a58908a );
 a58915a <=( (not A300)  and  A299 );
 a58918a <=( (not A302)  and  (not A301) );
 a58919a <=( a58918a  and  a58915a );
 a58920a <=( a58919a  and  a58912a );
 a58923a <=( (not A169)  and  A170 );
 a58926a <=( (not A167)  and  (not A168) );
 a58927a <=( a58926a  and  a58923a );
 a58930a <=( (not A201)  and  A166 );
 a58933a <=( (not A232)  and  A202 );
 a58934a <=( a58933a  and  a58930a );
 a58935a <=( a58934a  and  a58927a );
 a58938a <=( A234  and  A233 );
 a58941a <=( (not A265)  and  A236 );
 a58942a <=( a58941a  and  a58938a );
 a58945a <=( (not A267)  and  A266 );
 a58948a <=( (not A269)  and  (not A268) );
 a58949a <=( a58948a  and  a58945a );
 a58950a <=( a58949a  and  a58942a );
 a58953a <=( (not A169)  and  A170 );
 a58956a <=( (not A167)  and  (not A168) );
 a58957a <=( a58956a  and  a58953a );
 a58960a <=( (not A201)  and  A166 );
 a58963a <=( (not A232)  and  A202 );
 a58964a <=( a58963a  and  a58960a );
 a58965a <=( a58964a  and  a58957a );
 a58968a <=( A234  and  A233 );
 a58971a <=( A265  and  A236 );
 a58972a <=( a58971a  and  a58968a );
 a58975a <=( (not A267)  and  (not A266) );
 a58978a <=( (not A269)  and  (not A268) );
 a58979a <=( a58978a  and  a58975a );
 a58980a <=( a58979a  and  a58972a );
 a58983a <=( (not A169)  and  A170 );
 a58986a <=( (not A167)  and  (not A168) );
 a58987a <=( a58986a  and  a58983a );
 a58990a <=( (not A201)  and  A166 );
 a58993a <=( (not A232)  and  A202 );
 a58994a <=( a58993a  and  a58990a );
 a58995a <=( a58994a  and  a58987a );
 a58998a <=( (not A234)  and  A233 );
 a59001a <=( (not A236)  and  (not A235) );
 a59002a <=( a59001a  and  a58998a );
 a59005a <=( (not A299)  and  A298 );
 a59008a <=( A301  and  A300 );
 a59009a <=( a59008a  and  a59005a );
 a59010a <=( a59009a  and  a59002a );
 a59013a <=( (not A169)  and  A170 );
 a59016a <=( (not A167)  and  (not A168) );
 a59017a <=( a59016a  and  a59013a );
 a59020a <=( (not A201)  and  A166 );
 a59023a <=( (not A232)  and  A202 );
 a59024a <=( a59023a  and  a59020a );
 a59025a <=( a59024a  and  a59017a );
 a59028a <=( (not A234)  and  A233 );
 a59031a <=( (not A236)  and  (not A235) );
 a59032a <=( a59031a  and  a59028a );
 a59035a <=( (not A299)  and  A298 );
 a59038a <=( A302  and  A300 );
 a59039a <=( a59038a  and  a59035a );
 a59040a <=( a59039a  and  a59032a );
 a59043a <=( (not A169)  and  A170 );
 a59046a <=( (not A167)  and  (not A168) );
 a59047a <=( a59046a  and  a59043a );
 a59050a <=( (not A201)  and  A166 );
 a59053a <=( (not A232)  and  A202 );
 a59054a <=( a59053a  and  a59050a );
 a59055a <=( a59054a  and  a59047a );
 a59058a <=( (not A234)  and  A233 );
 a59061a <=( (not A236)  and  (not A235) );
 a59062a <=( a59061a  and  a59058a );
 a59065a <=( A299  and  (not A298) );
 a59068a <=( A301  and  A300 );
 a59069a <=( a59068a  and  a59065a );
 a59070a <=( a59069a  and  a59062a );
 a59073a <=( (not A169)  and  A170 );
 a59076a <=( (not A167)  and  (not A168) );
 a59077a <=( a59076a  and  a59073a );
 a59080a <=( (not A201)  and  A166 );
 a59083a <=( (not A232)  and  A202 );
 a59084a <=( a59083a  and  a59080a );
 a59085a <=( a59084a  and  a59077a );
 a59088a <=( (not A234)  and  A233 );
 a59091a <=( (not A236)  and  (not A235) );
 a59092a <=( a59091a  and  a59088a );
 a59095a <=( A299  and  (not A298) );
 a59098a <=( A302  and  A300 );
 a59099a <=( a59098a  and  a59095a );
 a59100a <=( a59099a  and  a59092a );
 a59103a <=( (not A169)  and  A170 );
 a59106a <=( (not A167)  and  (not A168) );
 a59107a <=( a59106a  and  a59103a );
 a59110a <=( (not A201)  and  A166 );
 a59113a <=( (not A232)  and  A202 );
 a59114a <=( a59113a  and  a59110a );
 a59115a <=( a59114a  and  a59107a );
 a59118a <=( (not A234)  and  A233 );
 a59121a <=( (not A236)  and  (not A235) );
 a59122a <=( a59121a  and  a59118a );
 a59125a <=( A266  and  (not A265) );
 a59128a <=( A268  and  A267 );
 a59129a <=( a59128a  and  a59125a );
 a59130a <=( a59129a  and  a59122a );
 a59133a <=( (not A169)  and  A170 );
 a59136a <=( (not A167)  and  (not A168) );
 a59137a <=( a59136a  and  a59133a );
 a59140a <=( (not A201)  and  A166 );
 a59143a <=( (not A232)  and  A202 );
 a59144a <=( a59143a  and  a59140a );
 a59145a <=( a59144a  and  a59137a );
 a59148a <=( (not A234)  and  A233 );
 a59151a <=( (not A236)  and  (not A235) );
 a59152a <=( a59151a  and  a59148a );
 a59155a <=( A266  and  (not A265) );
 a59158a <=( A269  and  A267 );
 a59159a <=( a59158a  and  a59155a );
 a59160a <=( a59159a  and  a59152a );
 a59163a <=( (not A169)  and  A170 );
 a59166a <=( (not A167)  and  (not A168) );
 a59167a <=( a59166a  and  a59163a );
 a59170a <=( (not A201)  and  A166 );
 a59173a <=( (not A232)  and  A202 );
 a59174a <=( a59173a  and  a59170a );
 a59175a <=( a59174a  and  a59167a );
 a59178a <=( (not A234)  and  A233 );
 a59181a <=( (not A236)  and  (not A235) );
 a59182a <=( a59181a  and  a59178a );
 a59185a <=( (not A266)  and  A265 );
 a59188a <=( A268  and  A267 );
 a59189a <=( a59188a  and  a59185a );
 a59190a <=( a59189a  and  a59182a );
 a59193a <=( (not A169)  and  A170 );
 a59196a <=( (not A167)  and  (not A168) );
 a59197a <=( a59196a  and  a59193a );
 a59200a <=( (not A201)  and  A166 );
 a59203a <=( (not A232)  and  A202 );
 a59204a <=( a59203a  and  a59200a );
 a59205a <=( a59204a  and  a59197a );
 a59208a <=( (not A234)  and  A233 );
 a59211a <=( (not A236)  and  (not A235) );
 a59212a <=( a59211a  and  a59208a );
 a59215a <=( (not A266)  and  A265 );
 a59218a <=( A269  and  A267 );
 a59219a <=( a59218a  and  a59215a );
 a59220a <=( a59219a  and  a59212a );
 a59223a <=( (not A169)  and  A170 );
 a59226a <=( (not A167)  and  (not A168) );
 a59227a <=( a59226a  and  a59223a );
 a59230a <=( (not A201)  and  A166 );
 a59233a <=( A232  and  A202 );
 a59234a <=( a59233a  and  a59230a );
 a59235a <=( a59234a  and  a59227a );
 a59238a <=( A234  and  (not A233) );
 a59241a <=( A298  and  A235 );
 a59242a <=( a59241a  and  a59238a );
 a59245a <=( (not A300)  and  (not A299) );
 a59248a <=( (not A302)  and  (not A301) );
 a59249a <=( a59248a  and  a59245a );
 a59250a <=( a59249a  and  a59242a );
 a59253a <=( (not A169)  and  A170 );
 a59256a <=( (not A167)  and  (not A168) );
 a59257a <=( a59256a  and  a59253a );
 a59260a <=( (not A201)  and  A166 );
 a59263a <=( A232  and  A202 );
 a59264a <=( a59263a  and  a59260a );
 a59265a <=( a59264a  and  a59257a );
 a59268a <=( A234  and  (not A233) );
 a59271a <=( (not A298)  and  A235 );
 a59272a <=( a59271a  and  a59268a );
 a59275a <=( (not A300)  and  A299 );
 a59278a <=( (not A302)  and  (not A301) );
 a59279a <=( a59278a  and  a59275a );
 a59280a <=( a59279a  and  a59272a );
 a59283a <=( (not A169)  and  A170 );
 a59286a <=( (not A167)  and  (not A168) );
 a59287a <=( a59286a  and  a59283a );
 a59290a <=( (not A201)  and  A166 );
 a59293a <=( A232  and  A202 );
 a59294a <=( a59293a  and  a59290a );
 a59295a <=( a59294a  and  a59287a );
 a59298a <=( A234  and  (not A233) );
 a59301a <=( (not A265)  and  A235 );
 a59302a <=( a59301a  and  a59298a );
 a59305a <=( (not A267)  and  A266 );
 a59308a <=( (not A269)  and  (not A268) );
 a59309a <=( a59308a  and  a59305a );
 a59310a <=( a59309a  and  a59302a );
 a59313a <=( (not A169)  and  A170 );
 a59316a <=( (not A167)  and  (not A168) );
 a59317a <=( a59316a  and  a59313a );
 a59320a <=( (not A201)  and  A166 );
 a59323a <=( A232  and  A202 );
 a59324a <=( a59323a  and  a59320a );
 a59325a <=( a59324a  and  a59317a );
 a59328a <=( A234  and  (not A233) );
 a59331a <=( A265  and  A235 );
 a59332a <=( a59331a  and  a59328a );
 a59335a <=( (not A267)  and  (not A266) );
 a59338a <=( (not A269)  and  (not A268) );
 a59339a <=( a59338a  and  a59335a );
 a59340a <=( a59339a  and  a59332a );
 a59343a <=( (not A169)  and  A170 );
 a59346a <=( (not A167)  and  (not A168) );
 a59347a <=( a59346a  and  a59343a );
 a59350a <=( (not A201)  and  A166 );
 a59353a <=( A232  and  A202 );
 a59354a <=( a59353a  and  a59350a );
 a59355a <=( a59354a  and  a59347a );
 a59358a <=( A234  and  (not A233) );
 a59361a <=( A298  and  A236 );
 a59362a <=( a59361a  and  a59358a );
 a59365a <=( (not A300)  and  (not A299) );
 a59368a <=( (not A302)  and  (not A301) );
 a59369a <=( a59368a  and  a59365a );
 a59370a <=( a59369a  and  a59362a );
 a59373a <=( (not A169)  and  A170 );
 a59376a <=( (not A167)  and  (not A168) );
 a59377a <=( a59376a  and  a59373a );
 a59380a <=( (not A201)  and  A166 );
 a59383a <=( A232  and  A202 );
 a59384a <=( a59383a  and  a59380a );
 a59385a <=( a59384a  and  a59377a );
 a59388a <=( A234  and  (not A233) );
 a59391a <=( (not A298)  and  A236 );
 a59392a <=( a59391a  and  a59388a );
 a59395a <=( (not A300)  and  A299 );
 a59398a <=( (not A302)  and  (not A301) );
 a59399a <=( a59398a  and  a59395a );
 a59400a <=( a59399a  and  a59392a );
 a59403a <=( (not A169)  and  A170 );
 a59406a <=( (not A167)  and  (not A168) );
 a59407a <=( a59406a  and  a59403a );
 a59410a <=( (not A201)  and  A166 );
 a59413a <=( A232  and  A202 );
 a59414a <=( a59413a  and  a59410a );
 a59415a <=( a59414a  and  a59407a );
 a59418a <=( A234  and  (not A233) );
 a59421a <=( (not A265)  and  A236 );
 a59422a <=( a59421a  and  a59418a );
 a59425a <=( (not A267)  and  A266 );
 a59428a <=( (not A269)  and  (not A268) );
 a59429a <=( a59428a  and  a59425a );
 a59430a <=( a59429a  and  a59422a );
 a59433a <=( (not A169)  and  A170 );
 a59436a <=( (not A167)  and  (not A168) );
 a59437a <=( a59436a  and  a59433a );
 a59440a <=( (not A201)  and  A166 );
 a59443a <=( A232  and  A202 );
 a59444a <=( a59443a  and  a59440a );
 a59445a <=( a59444a  and  a59437a );
 a59448a <=( A234  and  (not A233) );
 a59451a <=( A265  and  A236 );
 a59452a <=( a59451a  and  a59448a );
 a59455a <=( (not A267)  and  (not A266) );
 a59458a <=( (not A269)  and  (not A268) );
 a59459a <=( a59458a  and  a59455a );
 a59460a <=( a59459a  and  a59452a );
 a59463a <=( (not A169)  and  A170 );
 a59466a <=( (not A167)  and  (not A168) );
 a59467a <=( a59466a  and  a59463a );
 a59470a <=( (not A201)  and  A166 );
 a59473a <=( A232  and  A202 );
 a59474a <=( a59473a  and  a59470a );
 a59475a <=( a59474a  and  a59467a );
 a59478a <=( (not A234)  and  (not A233) );
 a59481a <=( (not A236)  and  (not A235) );
 a59482a <=( a59481a  and  a59478a );
 a59485a <=( (not A299)  and  A298 );
 a59488a <=( A301  and  A300 );
 a59489a <=( a59488a  and  a59485a );
 a59490a <=( a59489a  and  a59482a );
 a59493a <=( (not A169)  and  A170 );
 a59496a <=( (not A167)  and  (not A168) );
 a59497a <=( a59496a  and  a59493a );
 a59500a <=( (not A201)  and  A166 );
 a59503a <=( A232  and  A202 );
 a59504a <=( a59503a  and  a59500a );
 a59505a <=( a59504a  and  a59497a );
 a59508a <=( (not A234)  and  (not A233) );
 a59511a <=( (not A236)  and  (not A235) );
 a59512a <=( a59511a  and  a59508a );
 a59515a <=( (not A299)  and  A298 );
 a59518a <=( A302  and  A300 );
 a59519a <=( a59518a  and  a59515a );
 a59520a <=( a59519a  and  a59512a );
 a59523a <=( (not A169)  and  A170 );
 a59526a <=( (not A167)  and  (not A168) );
 a59527a <=( a59526a  and  a59523a );
 a59530a <=( (not A201)  and  A166 );
 a59533a <=( A232  and  A202 );
 a59534a <=( a59533a  and  a59530a );
 a59535a <=( a59534a  and  a59527a );
 a59538a <=( (not A234)  and  (not A233) );
 a59541a <=( (not A236)  and  (not A235) );
 a59542a <=( a59541a  and  a59538a );
 a59545a <=( A299  and  (not A298) );
 a59548a <=( A301  and  A300 );
 a59549a <=( a59548a  and  a59545a );
 a59550a <=( a59549a  and  a59542a );
 a59553a <=( (not A169)  and  A170 );
 a59556a <=( (not A167)  and  (not A168) );
 a59557a <=( a59556a  and  a59553a );
 a59560a <=( (not A201)  and  A166 );
 a59563a <=( A232  and  A202 );
 a59564a <=( a59563a  and  a59560a );
 a59565a <=( a59564a  and  a59557a );
 a59568a <=( (not A234)  and  (not A233) );
 a59571a <=( (not A236)  and  (not A235) );
 a59572a <=( a59571a  and  a59568a );
 a59575a <=( A299  and  (not A298) );
 a59578a <=( A302  and  A300 );
 a59579a <=( a59578a  and  a59575a );
 a59580a <=( a59579a  and  a59572a );
 a59583a <=( (not A169)  and  A170 );
 a59586a <=( (not A167)  and  (not A168) );
 a59587a <=( a59586a  and  a59583a );
 a59590a <=( (not A201)  and  A166 );
 a59593a <=( A232  and  A202 );
 a59594a <=( a59593a  and  a59590a );
 a59595a <=( a59594a  and  a59587a );
 a59598a <=( (not A234)  and  (not A233) );
 a59601a <=( (not A236)  and  (not A235) );
 a59602a <=( a59601a  and  a59598a );
 a59605a <=( A266  and  (not A265) );
 a59608a <=( A268  and  A267 );
 a59609a <=( a59608a  and  a59605a );
 a59610a <=( a59609a  and  a59602a );
 a59613a <=( (not A169)  and  A170 );
 a59616a <=( (not A167)  and  (not A168) );
 a59617a <=( a59616a  and  a59613a );
 a59620a <=( (not A201)  and  A166 );
 a59623a <=( A232  and  A202 );
 a59624a <=( a59623a  and  a59620a );
 a59625a <=( a59624a  and  a59617a );
 a59628a <=( (not A234)  and  (not A233) );
 a59631a <=( (not A236)  and  (not A235) );
 a59632a <=( a59631a  and  a59628a );
 a59635a <=( A266  and  (not A265) );
 a59638a <=( A269  and  A267 );
 a59639a <=( a59638a  and  a59635a );
 a59640a <=( a59639a  and  a59632a );
 a59643a <=( (not A169)  and  A170 );
 a59646a <=( (not A167)  and  (not A168) );
 a59647a <=( a59646a  and  a59643a );
 a59650a <=( (not A201)  and  A166 );
 a59653a <=( A232  and  A202 );
 a59654a <=( a59653a  and  a59650a );
 a59655a <=( a59654a  and  a59647a );
 a59658a <=( (not A234)  and  (not A233) );
 a59661a <=( (not A236)  and  (not A235) );
 a59662a <=( a59661a  and  a59658a );
 a59665a <=( (not A266)  and  A265 );
 a59668a <=( A268  and  A267 );
 a59669a <=( a59668a  and  a59665a );
 a59670a <=( a59669a  and  a59662a );
 a59673a <=( (not A169)  and  A170 );
 a59676a <=( (not A167)  and  (not A168) );
 a59677a <=( a59676a  and  a59673a );
 a59680a <=( (not A201)  and  A166 );
 a59683a <=( A232  and  A202 );
 a59684a <=( a59683a  and  a59680a );
 a59685a <=( a59684a  and  a59677a );
 a59688a <=( (not A234)  and  (not A233) );
 a59691a <=( (not A236)  and  (not A235) );
 a59692a <=( a59691a  and  a59688a );
 a59695a <=( (not A266)  and  A265 );
 a59698a <=( A269  and  A267 );
 a59699a <=( a59698a  and  a59695a );
 a59700a <=( a59699a  and  a59692a );
 a59703a <=( (not A169)  and  A170 );
 a59706a <=( (not A167)  and  (not A168) );
 a59707a <=( a59706a  and  a59703a );
 a59710a <=( (not A201)  and  A166 );
 a59713a <=( (not A232)  and  A203 );
 a59714a <=( a59713a  and  a59710a );
 a59715a <=( a59714a  and  a59707a );
 a59718a <=( A234  and  A233 );
 a59721a <=( A298  and  A235 );
 a59722a <=( a59721a  and  a59718a );
 a59725a <=( (not A300)  and  (not A299) );
 a59728a <=( (not A302)  and  (not A301) );
 a59729a <=( a59728a  and  a59725a );
 a59730a <=( a59729a  and  a59722a );
 a59733a <=( (not A169)  and  A170 );
 a59736a <=( (not A167)  and  (not A168) );
 a59737a <=( a59736a  and  a59733a );
 a59740a <=( (not A201)  and  A166 );
 a59743a <=( (not A232)  and  A203 );
 a59744a <=( a59743a  and  a59740a );
 a59745a <=( a59744a  and  a59737a );
 a59748a <=( A234  and  A233 );
 a59751a <=( (not A298)  and  A235 );
 a59752a <=( a59751a  and  a59748a );
 a59755a <=( (not A300)  and  A299 );
 a59758a <=( (not A302)  and  (not A301) );
 a59759a <=( a59758a  and  a59755a );
 a59760a <=( a59759a  and  a59752a );
 a59763a <=( (not A169)  and  A170 );
 a59766a <=( (not A167)  and  (not A168) );
 a59767a <=( a59766a  and  a59763a );
 a59770a <=( (not A201)  and  A166 );
 a59773a <=( (not A232)  and  A203 );
 a59774a <=( a59773a  and  a59770a );
 a59775a <=( a59774a  and  a59767a );
 a59778a <=( A234  and  A233 );
 a59781a <=( (not A265)  and  A235 );
 a59782a <=( a59781a  and  a59778a );
 a59785a <=( (not A267)  and  A266 );
 a59788a <=( (not A269)  and  (not A268) );
 a59789a <=( a59788a  and  a59785a );
 a59790a <=( a59789a  and  a59782a );
 a59793a <=( (not A169)  and  A170 );
 a59796a <=( (not A167)  and  (not A168) );
 a59797a <=( a59796a  and  a59793a );
 a59800a <=( (not A201)  and  A166 );
 a59803a <=( (not A232)  and  A203 );
 a59804a <=( a59803a  and  a59800a );
 a59805a <=( a59804a  and  a59797a );
 a59808a <=( A234  and  A233 );
 a59811a <=( A265  and  A235 );
 a59812a <=( a59811a  and  a59808a );
 a59815a <=( (not A267)  and  (not A266) );
 a59818a <=( (not A269)  and  (not A268) );
 a59819a <=( a59818a  and  a59815a );
 a59820a <=( a59819a  and  a59812a );
 a59823a <=( (not A169)  and  A170 );
 a59826a <=( (not A167)  and  (not A168) );
 a59827a <=( a59826a  and  a59823a );
 a59830a <=( (not A201)  and  A166 );
 a59833a <=( (not A232)  and  A203 );
 a59834a <=( a59833a  and  a59830a );
 a59835a <=( a59834a  and  a59827a );
 a59838a <=( A234  and  A233 );
 a59841a <=( A298  and  A236 );
 a59842a <=( a59841a  and  a59838a );
 a59845a <=( (not A300)  and  (not A299) );
 a59848a <=( (not A302)  and  (not A301) );
 a59849a <=( a59848a  and  a59845a );
 a59850a <=( a59849a  and  a59842a );
 a59853a <=( (not A169)  and  A170 );
 a59856a <=( (not A167)  and  (not A168) );
 a59857a <=( a59856a  and  a59853a );
 a59860a <=( (not A201)  and  A166 );
 a59863a <=( (not A232)  and  A203 );
 a59864a <=( a59863a  and  a59860a );
 a59865a <=( a59864a  and  a59857a );
 a59868a <=( A234  and  A233 );
 a59871a <=( (not A298)  and  A236 );
 a59872a <=( a59871a  and  a59868a );
 a59875a <=( (not A300)  and  A299 );
 a59878a <=( (not A302)  and  (not A301) );
 a59879a <=( a59878a  and  a59875a );
 a59880a <=( a59879a  and  a59872a );
 a59883a <=( (not A169)  and  A170 );
 a59886a <=( (not A167)  and  (not A168) );
 a59887a <=( a59886a  and  a59883a );
 a59890a <=( (not A201)  and  A166 );
 a59893a <=( (not A232)  and  A203 );
 a59894a <=( a59893a  and  a59890a );
 a59895a <=( a59894a  and  a59887a );
 a59898a <=( A234  and  A233 );
 a59901a <=( (not A265)  and  A236 );
 a59902a <=( a59901a  and  a59898a );
 a59905a <=( (not A267)  and  A266 );
 a59908a <=( (not A269)  and  (not A268) );
 a59909a <=( a59908a  and  a59905a );
 a59910a <=( a59909a  and  a59902a );
 a59913a <=( (not A169)  and  A170 );
 a59916a <=( (not A167)  and  (not A168) );
 a59917a <=( a59916a  and  a59913a );
 a59920a <=( (not A201)  and  A166 );
 a59923a <=( (not A232)  and  A203 );
 a59924a <=( a59923a  and  a59920a );
 a59925a <=( a59924a  and  a59917a );
 a59928a <=( A234  and  A233 );
 a59931a <=( A265  and  A236 );
 a59932a <=( a59931a  and  a59928a );
 a59935a <=( (not A267)  and  (not A266) );
 a59938a <=( (not A269)  and  (not A268) );
 a59939a <=( a59938a  and  a59935a );
 a59940a <=( a59939a  and  a59932a );
 a59943a <=( (not A169)  and  A170 );
 a59946a <=( (not A167)  and  (not A168) );
 a59947a <=( a59946a  and  a59943a );
 a59950a <=( (not A201)  and  A166 );
 a59953a <=( (not A232)  and  A203 );
 a59954a <=( a59953a  and  a59950a );
 a59955a <=( a59954a  and  a59947a );
 a59958a <=( (not A234)  and  A233 );
 a59961a <=( (not A236)  and  (not A235) );
 a59962a <=( a59961a  and  a59958a );
 a59965a <=( (not A299)  and  A298 );
 a59968a <=( A301  and  A300 );
 a59969a <=( a59968a  and  a59965a );
 a59970a <=( a59969a  and  a59962a );
 a59973a <=( (not A169)  and  A170 );
 a59976a <=( (not A167)  and  (not A168) );
 a59977a <=( a59976a  and  a59973a );
 a59980a <=( (not A201)  and  A166 );
 a59983a <=( (not A232)  and  A203 );
 a59984a <=( a59983a  and  a59980a );
 a59985a <=( a59984a  and  a59977a );
 a59988a <=( (not A234)  and  A233 );
 a59991a <=( (not A236)  and  (not A235) );
 a59992a <=( a59991a  and  a59988a );
 a59995a <=( (not A299)  and  A298 );
 a59998a <=( A302  and  A300 );
 a59999a <=( a59998a  and  a59995a );
 a60000a <=( a59999a  and  a59992a );
 a60003a <=( (not A169)  and  A170 );
 a60006a <=( (not A167)  and  (not A168) );
 a60007a <=( a60006a  and  a60003a );
 a60010a <=( (not A201)  and  A166 );
 a60013a <=( (not A232)  and  A203 );
 a60014a <=( a60013a  and  a60010a );
 a60015a <=( a60014a  and  a60007a );
 a60018a <=( (not A234)  and  A233 );
 a60021a <=( (not A236)  and  (not A235) );
 a60022a <=( a60021a  and  a60018a );
 a60025a <=( A299  and  (not A298) );
 a60028a <=( A301  and  A300 );
 a60029a <=( a60028a  and  a60025a );
 a60030a <=( a60029a  and  a60022a );
 a60033a <=( (not A169)  and  A170 );
 a60036a <=( (not A167)  and  (not A168) );
 a60037a <=( a60036a  and  a60033a );
 a60040a <=( (not A201)  and  A166 );
 a60043a <=( (not A232)  and  A203 );
 a60044a <=( a60043a  and  a60040a );
 a60045a <=( a60044a  and  a60037a );
 a60048a <=( (not A234)  and  A233 );
 a60051a <=( (not A236)  and  (not A235) );
 a60052a <=( a60051a  and  a60048a );
 a60055a <=( A299  and  (not A298) );
 a60058a <=( A302  and  A300 );
 a60059a <=( a60058a  and  a60055a );
 a60060a <=( a60059a  and  a60052a );
 a60063a <=( (not A169)  and  A170 );
 a60066a <=( (not A167)  and  (not A168) );
 a60067a <=( a60066a  and  a60063a );
 a60070a <=( (not A201)  and  A166 );
 a60073a <=( (not A232)  and  A203 );
 a60074a <=( a60073a  and  a60070a );
 a60075a <=( a60074a  and  a60067a );
 a60078a <=( (not A234)  and  A233 );
 a60081a <=( (not A236)  and  (not A235) );
 a60082a <=( a60081a  and  a60078a );
 a60085a <=( A266  and  (not A265) );
 a60088a <=( A268  and  A267 );
 a60089a <=( a60088a  and  a60085a );
 a60090a <=( a60089a  and  a60082a );
 a60093a <=( (not A169)  and  A170 );
 a60096a <=( (not A167)  and  (not A168) );
 a60097a <=( a60096a  and  a60093a );
 a60100a <=( (not A201)  and  A166 );
 a60103a <=( (not A232)  and  A203 );
 a60104a <=( a60103a  and  a60100a );
 a60105a <=( a60104a  and  a60097a );
 a60108a <=( (not A234)  and  A233 );
 a60111a <=( (not A236)  and  (not A235) );
 a60112a <=( a60111a  and  a60108a );
 a60115a <=( A266  and  (not A265) );
 a60118a <=( A269  and  A267 );
 a60119a <=( a60118a  and  a60115a );
 a60120a <=( a60119a  and  a60112a );
 a60123a <=( (not A169)  and  A170 );
 a60126a <=( (not A167)  and  (not A168) );
 a60127a <=( a60126a  and  a60123a );
 a60130a <=( (not A201)  and  A166 );
 a60133a <=( (not A232)  and  A203 );
 a60134a <=( a60133a  and  a60130a );
 a60135a <=( a60134a  and  a60127a );
 a60138a <=( (not A234)  and  A233 );
 a60141a <=( (not A236)  and  (not A235) );
 a60142a <=( a60141a  and  a60138a );
 a60145a <=( (not A266)  and  A265 );
 a60148a <=( A268  and  A267 );
 a60149a <=( a60148a  and  a60145a );
 a60150a <=( a60149a  and  a60142a );
 a60153a <=( (not A169)  and  A170 );
 a60156a <=( (not A167)  and  (not A168) );
 a60157a <=( a60156a  and  a60153a );
 a60160a <=( (not A201)  and  A166 );
 a60163a <=( (not A232)  and  A203 );
 a60164a <=( a60163a  and  a60160a );
 a60165a <=( a60164a  and  a60157a );
 a60168a <=( (not A234)  and  A233 );
 a60171a <=( (not A236)  and  (not A235) );
 a60172a <=( a60171a  and  a60168a );
 a60175a <=( (not A266)  and  A265 );
 a60178a <=( A269  and  A267 );
 a60179a <=( a60178a  and  a60175a );
 a60180a <=( a60179a  and  a60172a );
 a60183a <=( (not A169)  and  A170 );
 a60186a <=( (not A167)  and  (not A168) );
 a60187a <=( a60186a  and  a60183a );
 a60190a <=( (not A201)  and  A166 );
 a60193a <=( A232  and  A203 );
 a60194a <=( a60193a  and  a60190a );
 a60195a <=( a60194a  and  a60187a );
 a60198a <=( A234  and  (not A233) );
 a60201a <=( A298  and  A235 );
 a60202a <=( a60201a  and  a60198a );
 a60205a <=( (not A300)  and  (not A299) );
 a60208a <=( (not A302)  and  (not A301) );
 a60209a <=( a60208a  and  a60205a );
 a60210a <=( a60209a  and  a60202a );
 a60213a <=( (not A169)  and  A170 );
 a60216a <=( (not A167)  and  (not A168) );
 a60217a <=( a60216a  and  a60213a );
 a60220a <=( (not A201)  and  A166 );
 a60223a <=( A232  and  A203 );
 a60224a <=( a60223a  and  a60220a );
 a60225a <=( a60224a  and  a60217a );
 a60228a <=( A234  and  (not A233) );
 a60231a <=( (not A298)  and  A235 );
 a60232a <=( a60231a  and  a60228a );
 a60235a <=( (not A300)  and  A299 );
 a60238a <=( (not A302)  and  (not A301) );
 a60239a <=( a60238a  and  a60235a );
 a60240a <=( a60239a  and  a60232a );
 a60243a <=( (not A169)  and  A170 );
 a60246a <=( (not A167)  and  (not A168) );
 a60247a <=( a60246a  and  a60243a );
 a60250a <=( (not A201)  and  A166 );
 a60253a <=( A232  and  A203 );
 a60254a <=( a60253a  and  a60250a );
 a60255a <=( a60254a  and  a60247a );
 a60258a <=( A234  and  (not A233) );
 a60261a <=( (not A265)  and  A235 );
 a60262a <=( a60261a  and  a60258a );
 a60265a <=( (not A267)  and  A266 );
 a60268a <=( (not A269)  and  (not A268) );
 a60269a <=( a60268a  and  a60265a );
 a60270a <=( a60269a  and  a60262a );
 a60273a <=( (not A169)  and  A170 );
 a60276a <=( (not A167)  and  (not A168) );
 a60277a <=( a60276a  and  a60273a );
 a60280a <=( (not A201)  and  A166 );
 a60283a <=( A232  and  A203 );
 a60284a <=( a60283a  and  a60280a );
 a60285a <=( a60284a  and  a60277a );
 a60288a <=( A234  and  (not A233) );
 a60291a <=( A265  and  A235 );
 a60292a <=( a60291a  and  a60288a );
 a60295a <=( (not A267)  and  (not A266) );
 a60298a <=( (not A269)  and  (not A268) );
 a60299a <=( a60298a  and  a60295a );
 a60300a <=( a60299a  and  a60292a );
 a60303a <=( (not A169)  and  A170 );
 a60306a <=( (not A167)  and  (not A168) );
 a60307a <=( a60306a  and  a60303a );
 a60310a <=( (not A201)  and  A166 );
 a60313a <=( A232  and  A203 );
 a60314a <=( a60313a  and  a60310a );
 a60315a <=( a60314a  and  a60307a );
 a60318a <=( A234  and  (not A233) );
 a60321a <=( A298  and  A236 );
 a60322a <=( a60321a  and  a60318a );
 a60325a <=( (not A300)  and  (not A299) );
 a60328a <=( (not A302)  and  (not A301) );
 a60329a <=( a60328a  and  a60325a );
 a60330a <=( a60329a  and  a60322a );
 a60333a <=( (not A169)  and  A170 );
 a60336a <=( (not A167)  and  (not A168) );
 a60337a <=( a60336a  and  a60333a );
 a60340a <=( (not A201)  and  A166 );
 a60343a <=( A232  and  A203 );
 a60344a <=( a60343a  and  a60340a );
 a60345a <=( a60344a  and  a60337a );
 a60348a <=( A234  and  (not A233) );
 a60351a <=( (not A298)  and  A236 );
 a60352a <=( a60351a  and  a60348a );
 a60355a <=( (not A300)  and  A299 );
 a60358a <=( (not A302)  and  (not A301) );
 a60359a <=( a60358a  and  a60355a );
 a60360a <=( a60359a  and  a60352a );
 a60363a <=( (not A169)  and  A170 );
 a60366a <=( (not A167)  and  (not A168) );
 a60367a <=( a60366a  and  a60363a );
 a60370a <=( (not A201)  and  A166 );
 a60373a <=( A232  and  A203 );
 a60374a <=( a60373a  and  a60370a );
 a60375a <=( a60374a  and  a60367a );
 a60378a <=( A234  and  (not A233) );
 a60381a <=( (not A265)  and  A236 );
 a60382a <=( a60381a  and  a60378a );
 a60385a <=( (not A267)  and  A266 );
 a60388a <=( (not A269)  and  (not A268) );
 a60389a <=( a60388a  and  a60385a );
 a60390a <=( a60389a  and  a60382a );
 a60393a <=( (not A169)  and  A170 );
 a60396a <=( (not A167)  and  (not A168) );
 a60397a <=( a60396a  and  a60393a );
 a60400a <=( (not A201)  and  A166 );
 a60403a <=( A232  and  A203 );
 a60404a <=( a60403a  and  a60400a );
 a60405a <=( a60404a  and  a60397a );
 a60408a <=( A234  and  (not A233) );
 a60411a <=( A265  and  A236 );
 a60412a <=( a60411a  and  a60408a );
 a60415a <=( (not A267)  and  (not A266) );
 a60418a <=( (not A269)  and  (not A268) );
 a60419a <=( a60418a  and  a60415a );
 a60420a <=( a60419a  and  a60412a );
 a60423a <=( (not A169)  and  A170 );
 a60426a <=( (not A167)  and  (not A168) );
 a60427a <=( a60426a  and  a60423a );
 a60430a <=( (not A201)  and  A166 );
 a60433a <=( A232  and  A203 );
 a60434a <=( a60433a  and  a60430a );
 a60435a <=( a60434a  and  a60427a );
 a60438a <=( (not A234)  and  (not A233) );
 a60441a <=( (not A236)  and  (not A235) );
 a60442a <=( a60441a  and  a60438a );
 a60445a <=( (not A299)  and  A298 );
 a60448a <=( A301  and  A300 );
 a60449a <=( a60448a  and  a60445a );
 a60450a <=( a60449a  and  a60442a );
 a60453a <=( (not A169)  and  A170 );
 a60456a <=( (not A167)  and  (not A168) );
 a60457a <=( a60456a  and  a60453a );
 a60460a <=( (not A201)  and  A166 );
 a60463a <=( A232  and  A203 );
 a60464a <=( a60463a  and  a60460a );
 a60465a <=( a60464a  and  a60457a );
 a60468a <=( (not A234)  and  (not A233) );
 a60471a <=( (not A236)  and  (not A235) );
 a60472a <=( a60471a  and  a60468a );
 a60475a <=( (not A299)  and  A298 );
 a60478a <=( A302  and  A300 );
 a60479a <=( a60478a  and  a60475a );
 a60480a <=( a60479a  and  a60472a );
 a60483a <=( (not A169)  and  A170 );
 a60486a <=( (not A167)  and  (not A168) );
 a60487a <=( a60486a  and  a60483a );
 a60490a <=( (not A201)  and  A166 );
 a60493a <=( A232  and  A203 );
 a60494a <=( a60493a  and  a60490a );
 a60495a <=( a60494a  and  a60487a );
 a60498a <=( (not A234)  and  (not A233) );
 a60501a <=( (not A236)  and  (not A235) );
 a60502a <=( a60501a  and  a60498a );
 a60505a <=( A299  and  (not A298) );
 a60508a <=( A301  and  A300 );
 a60509a <=( a60508a  and  a60505a );
 a60510a <=( a60509a  and  a60502a );
 a60513a <=( (not A169)  and  A170 );
 a60516a <=( (not A167)  and  (not A168) );
 a60517a <=( a60516a  and  a60513a );
 a60520a <=( (not A201)  and  A166 );
 a60523a <=( A232  and  A203 );
 a60524a <=( a60523a  and  a60520a );
 a60525a <=( a60524a  and  a60517a );
 a60528a <=( (not A234)  and  (not A233) );
 a60531a <=( (not A236)  and  (not A235) );
 a60532a <=( a60531a  and  a60528a );
 a60535a <=( A299  and  (not A298) );
 a60538a <=( A302  and  A300 );
 a60539a <=( a60538a  and  a60535a );
 a60540a <=( a60539a  and  a60532a );
 a60543a <=( (not A169)  and  A170 );
 a60546a <=( (not A167)  and  (not A168) );
 a60547a <=( a60546a  and  a60543a );
 a60550a <=( (not A201)  and  A166 );
 a60553a <=( A232  and  A203 );
 a60554a <=( a60553a  and  a60550a );
 a60555a <=( a60554a  and  a60547a );
 a60558a <=( (not A234)  and  (not A233) );
 a60561a <=( (not A236)  and  (not A235) );
 a60562a <=( a60561a  and  a60558a );
 a60565a <=( A266  and  (not A265) );
 a60568a <=( A268  and  A267 );
 a60569a <=( a60568a  and  a60565a );
 a60570a <=( a60569a  and  a60562a );
 a60573a <=( (not A169)  and  A170 );
 a60576a <=( (not A167)  and  (not A168) );
 a60577a <=( a60576a  and  a60573a );
 a60580a <=( (not A201)  and  A166 );
 a60583a <=( A232  and  A203 );
 a60584a <=( a60583a  and  a60580a );
 a60585a <=( a60584a  and  a60577a );
 a60588a <=( (not A234)  and  (not A233) );
 a60591a <=( (not A236)  and  (not A235) );
 a60592a <=( a60591a  and  a60588a );
 a60595a <=( A266  and  (not A265) );
 a60598a <=( A269  and  A267 );
 a60599a <=( a60598a  and  a60595a );
 a60600a <=( a60599a  and  a60592a );
 a60603a <=( (not A169)  and  A170 );
 a60606a <=( (not A167)  and  (not A168) );
 a60607a <=( a60606a  and  a60603a );
 a60610a <=( (not A201)  and  A166 );
 a60613a <=( A232  and  A203 );
 a60614a <=( a60613a  and  a60610a );
 a60615a <=( a60614a  and  a60607a );
 a60618a <=( (not A234)  and  (not A233) );
 a60621a <=( (not A236)  and  (not A235) );
 a60622a <=( a60621a  and  a60618a );
 a60625a <=( (not A266)  and  A265 );
 a60628a <=( A268  and  A267 );
 a60629a <=( a60628a  and  a60625a );
 a60630a <=( a60629a  and  a60622a );
 a60633a <=( (not A169)  and  A170 );
 a60636a <=( (not A167)  and  (not A168) );
 a60637a <=( a60636a  and  a60633a );
 a60640a <=( (not A201)  and  A166 );
 a60643a <=( A232  and  A203 );
 a60644a <=( a60643a  and  a60640a );
 a60645a <=( a60644a  and  a60637a );
 a60648a <=( (not A234)  and  (not A233) );
 a60651a <=( (not A236)  and  (not A235) );
 a60652a <=( a60651a  and  a60648a );
 a60655a <=( (not A266)  and  A265 );
 a60658a <=( A269  and  A267 );
 a60659a <=( a60658a  and  a60655a );
 a60660a <=( a60659a  and  a60652a );
 a60663a <=( (not A169)  and  A170 );
 a60666a <=( (not A167)  and  (not A168) );
 a60667a <=( a60666a  and  a60663a );
 a60670a <=( A199  and  A166 );
 a60673a <=( (not A232)  and  A200 );
 a60674a <=( a60673a  and  a60670a );
 a60675a <=( a60674a  and  a60667a );
 a60678a <=( A234  and  A233 );
 a60681a <=( A298  and  A235 );
 a60682a <=( a60681a  and  a60678a );
 a60685a <=( (not A300)  and  (not A299) );
 a60688a <=( (not A302)  and  (not A301) );
 a60689a <=( a60688a  and  a60685a );
 a60690a <=( a60689a  and  a60682a );
 a60693a <=( (not A169)  and  A170 );
 a60696a <=( (not A167)  and  (not A168) );
 a60697a <=( a60696a  and  a60693a );
 a60700a <=( A199  and  A166 );
 a60703a <=( (not A232)  and  A200 );
 a60704a <=( a60703a  and  a60700a );
 a60705a <=( a60704a  and  a60697a );
 a60708a <=( A234  and  A233 );
 a60711a <=( (not A298)  and  A235 );
 a60712a <=( a60711a  and  a60708a );
 a60715a <=( (not A300)  and  A299 );
 a60718a <=( (not A302)  and  (not A301) );
 a60719a <=( a60718a  and  a60715a );
 a60720a <=( a60719a  and  a60712a );
 a60723a <=( (not A169)  and  A170 );
 a60726a <=( (not A167)  and  (not A168) );
 a60727a <=( a60726a  and  a60723a );
 a60730a <=( A199  and  A166 );
 a60733a <=( (not A232)  and  A200 );
 a60734a <=( a60733a  and  a60730a );
 a60735a <=( a60734a  and  a60727a );
 a60738a <=( A234  and  A233 );
 a60741a <=( (not A265)  and  A235 );
 a60742a <=( a60741a  and  a60738a );
 a60745a <=( (not A267)  and  A266 );
 a60748a <=( (not A269)  and  (not A268) );
 a60749a <=( a60748a  and  a60745a );
 a60750a <=( a60749a  and  a60742a );
 a60753a <=( (not A169)  and  A170 );
 a60756a <=( (not A167)  and  (not A168) );
 a60757a <=( a60756a  and  a60753a );
 a60760a <=( A199  and  A166 );
 a60763a <=( (not A232)  and  A200 );
 a60764a <=( a60763a  and  a60760a );
 a60765a <=( a60764a  and  a60757a );
 a60768a <=( A234  and  A233 );
 a60771a <=( A265  and  A235 );
 a60772a <=( a60771a  and  a60768a );
 a60775a <=( (not A267)  and  (not A266) );
 a60778a <=( (not A269)  and  (not A268) );
 a60779a <=( a60778a  and  a60775a );
 a60780a <=( a60779a  and  a60772a );
 a60783a <=( (not A169)  and  A170 );
 a60786a <=( (not A167)  and  (not A168) );
 a60787a <=( a60786a  and  a60783a );
 a60790a <=( A199  and  A166 );
 a60793a <=( (not A232)  and  A200 );
 a60794a <=( a60793a  and  a60790a );
 a60795a <=( a60794a  and  a60787a );
 a60798a <=( A234  and  A233 );
 a60801a <=( A298  and  A236 );
 a60802a <=( a60801a  and  a60798a );
 a60805a <=( (not A300)  and  (not A299) );
 a60808a <=( (not A302)  and  (not A301) );
 a60809a <=( a60808a  and  a60805a );
 a60810a <=( a60809a  and  a60802a );
 a60813a <=( (not A169)  and  A170 );
 a60816a <=( (not A167)  and  (not A168) );
 a60817a <=( a60816a  and  a60813a );
 a60820a <=( A199  and  A166 );
 a60823a <=( (not A232)  and  A200 );
 a60824a <=( a60823a  and  a60820a );
 a60825a <=( a60824a  and  a60817a );
 a60828a <=( A234  and  A233 );
 a60831a <=( (not A298)  and  A236 );
 a60832a <=( a60831a  and  a60828a );
 a60835a <=( (not A300)  and  A299 );
 a60838a <=( (not A302)  and  (not A301) );
 a60839a <=( a60838a  and  a60835a );
 a60840a <=( a60839a  and  a60832a );
 a60843a <=( (not A169)  and  A170 );
 a60846a <=( (not A167)  and  (not A168) );
 a60847a <=( a60846a  and  a60843a );
 a60850a <=( A199  and  A166 );
 a60853a <=( (not A232)  and  A200 );
 a60854a <=( a60853a  and  a60850a );
 a60855a <=( a60854a  and  a60847a );
 a60858a <=( A234  and  A233 );
 a60861a <=( (not A265)  and  A236 );
 a60862a <=( a60861a  and  a60858a );
 a60865a <=( (not A267)  and  A266 );
 a60868a <=( (not A269)  and  (not A268) );
 a60869a <=( a60868a  and  a60865a );
 a60870a <=( a60869a  and  a60862a );
 a60873a <=( (not A169)  and  A170 );
 a60876a <=( (not A167)  and  (not A168) );
 a60877a <=( a60876a  and  a60873a );
 a60880a <=( A199  and  A166 );
 a60883a <=( (not A232)  and  A200 );
 a60884a <=( a60883a  and  a60880a );
 a60885a <=( a60884a  and  a60877a );
 a60888a <=( A234  and  A233 );
 a60891a <=( A265  and  A236 );
 a60892a <=( a60891a  and  a60888a );
 a60895a <=( (not A267)  and  (not A266) );
 a60898a <=( (not A269)  and  (not A268) );
 a60899a <=( a60898a  and  a60895a );
 a60900a <=( a60899a  and  a60892a );
 a60903a <=( (not A169)  and  A170 );
 a60906a <=( (not A167)  and  (not A168) );
 a60907a <=( a60906a  and  a60903a );
 a60910a <=( A199  and  A166 );
 a60913a <=( (not A232)  and  A200 );
 a60914a <=( a60913a  and  a60910a );
 a60915a <=( a60914a  and  a60907a );
 a60918a <=( (not A234)  and  A233 );
 a60921a <=( (not A236)  and  (not A235) );
 a60922a <=( a60921a  and  a60918a );
 a60925a <=( (not A299)  and  A298 );
 a60928a <=( A301  and  A300 );
 a60929a <=( a60928a  and  a60925a );
 a60930a <=( a60929a  and  a60922a );
 a60933a <=( (not A169)  and  A170 );
 a60936a <=( (not A167)  and  (not A168) );
 a60937a <=( a60936a  and  a60933a );
 a60940a <=( A199  and  A166 );
 a60943a <=( (not A232)  and  A200 );
 a60944a <=( a60943a  and  a60940a );
 a60945a <=( a60944a  and  a60937a );
 a60948a <=( (not A234)  and  A233 );
 a60951a <=( (not A236)  and  (not A235) );
 a60952a <=( a60951a  and  a60948a );
 a60955a <=( (not A299)  and  A298 );
 a60958a <=( A302  and  A300 );
 a60959a <=( a60958a  and  a60955a );
 a60960a <=( a60959a  and  a60952a );
 a60963a <=( (not A169)  and  A170 );
 a60966a <=( (not A167)  and  (not A168) );
 a60967a <=( a60966a  and  a60963a );
 a60970a <=( A199  and  A166 );
 a60973a <=( (not A232)  and  A200 );
 a60974a <=( a60973a  and  a60970a );
 a60975a <=( a60974a  and  a60967a );
 a60978a <=( (not A234)  and  A233 );
 a60981a <=( (not A236)  and  (not A235) );
 a60982a <=( a60981a  and  a60978a );
 a60985a <=( A299  and  (not A298) );
 a60988a <=( A301  and  A300 );
 a60989a <=( a60988a  and  a60985a );
 a60990a <=( a60989a  and  a60982a );
 a60993a <=( (not A169)  and  A170 );
 a60996a <=( (not A167)  and  (not A168) );
 a60997a <=( a60996a  and  a60993a );
 a61000a <=( A199  and  A166 );
 a61003a <=( (not A232)  and  A200 );
 a61004a <=( a61003a  and  a61000a );
 a61005a <=( a61004a  and  a60997a );
 a61008a <=( (not A234)  and  A233 );
 a61011a <=( (not A236)  and  (not A235) );
 a61012a <=( a61011a  and  a61008a );
 a61015a <=( A299  and  (not A298) );
 a61018a <=( A302  and  A300 );
 a61019a <=( a61018a  and  a61015a );
 a61020a <=( a61019a  and  a61012a );
 a61023a <=( (not A169)  and  A170 );
 a61026a <=( (not A167)  and  (not A168) );
 a61027a <=( a61026a  and  a61023a );
 a61030a <=( A199  and  A166 );
 a61033a <=( (not A232)  and  A200 );
 a61034a <=( a61033a  and  a61030a );
 a61035a <=( a61034a  and  a61027a );
 a61038a <=( (not A234)  and  A233 );
 a61041a <=( (not A236)  and  (not A235) );
 a61042a <=( a61041a  and  a61038a );
 a61045a <=( A266  and  (not A265) );
 a61048a <=( A268  and  A267 );
 a61049a <=( a61048a  and  a61045a );
 a61050a <=( a61049a  and  a61042a );
 a61053a <=( (not A169)  and  A170 );
 a61056a <=( (not A167)  and  (not A168) );
 a61057a <=( a61056a  and  a61053a );
 a61060a <=( A199  and  A166 );
 a61063a <=( (not A232)  and  A200 );
 a61064a <=( a61063a  and  a61060a );
 a61065a <=( a61064a  and  a61057a );
 a61068a <=( (not A234)  and  A233 );
 a61071a <=( (not A236)  and  (not A235) );
 a61072a <=( a61071a  and  a61068a );
 a61075a <=( A266  and  (not A265) );
 a61078a <=( A269  and  A267 );
 a61079a <=( a61078a  and  a61075a );
 a61080a <=( a61079a  and  a61072a );
 a61083a <=( (not A169)  and  A170 );
 a61086a <=( (not A167)  and  (not A168) );
 a61087a <=( a61086a  and  a61083a );
 a61090a <=( A199  and  A166 );
 a61093a <=( (not A232)  and  A200 );
 a61094a <=( a61093a  and  a61090a );
 a61095a <=( a61094a  and  a61087a );
 a61098a <=( (not A234)  and  A233 );
 a61101a <=( (not A236)  and  (not A235) );
 a61102a <=( a61101a  and  a61098a );
 a61105a <=( (not A266)  and  A265 );
 a61108a <=( A268  and  A267 );
 a61109a <=( a61108a  and  a61105a );
 a61110a <=( a61109a  and  a61102a );
 a61113a <=( (not A169)  and  A170 );
 a61116a <=( (not A167)  and  (not A168) );
 a61117a <=( a61116a  and  a61113a );
 a61120a <=( A199  and  A166 );
 a61123a <=( (not A232)  and  A200 );
 a61124a <=( a61123a  and  a61120a );
 a61125a <=( a61124a  and  a61117a );
 a61128a <=( (not A234)  and  A233 );
 a61131a <=( (not A236)  and  (not A235) );
 a61132a <=( a61131a  and  a61128a );
 a61135a <=( (not A266)  and  A265 );
 a61138a <=( A269  and  A267 );
 a61139a <=( a61138a  and  a61135a );
 a61140a <=( a61139a  and  a61132a );
 a61143a <=( (not A169)  and  A170 );
 a61146a <=( (not A167)  and  (not A168) );
 a61147a <=( a61146a  and  a61143a );
 a61150a <=( A199  and  A166 );
 a61153a <=( A232  and  A200 );
 a61154a <=( a61153a  and  a61150a );
 a61155a <=( a61154a  and  a61147a );
 a61158a <=( A234  and  (not A233) );
 a61161a <=( A298  and  A235 );
 a61162a <=( a61161a  and  a61158a );
 a61165a <=( (not A300)  and  (not A299) );
 a61168a <=( (not A302)  and  (not A301) );
 a61169a <=( a61168a  and  a61165a );
 a61170a <=( a61169a  and  a61162a );
 a61173a <=( (not A169)  and  A170 );
 a61176a <=( (not A167)  and  (not A168) );
 a61177a <=( a61176a  and  a61173a );
 a61180a <=( A199  and  A166 );
 a61183a <=( A232  and  A200 );
 a61184a <=( a61183a  and  a61180a );
 a61185a <=( a61184a  and  a61177a );
 a61188a <=( A234  and  (not A233) );
 a61191a <=( (not A298)  and  A235 );
 a61192a <=( a61191a  and  a61188a );
 a61195a <=( (not A300)  and  A299 );
 a61198a <=( (not A302)  and  (not A301) );
 a61199a <=( a61198a  and  a61195a );
 a61200a <=( a61199a  and  a61192a );
 a61203a <=( (not A169)  and  A170 );
 a61206a <=( (not A167)  and  (not A168) );
 a61207a <=( a61206a  and  a61203a );
 a61210a <=( A199  and  A166 );
 a61213a <=( A232  and  A200 );
 a61214a <=( a61213a  and  a61210a );
 a61215a <=( a61214a  and  a61207a );
 a61218a <=( A234  and  (not A233) );
 a61221a <=( (not A265)  and  A235 );
 a61222a <=( a61221a  and  a61218a );
 a61225a <=( (not A267)  and  A266 );
 a61228a <=( (not A269)  and  (not A268) );
 a61229a <=( a61228a  and  a61225a );
 a61230a <=( a61229a  and  a61222a );
 a61233a <=( (not A169)  and  A170 );
 a61236a <=( (not A167)  and  (not A168) );
 a61237a <=( a61236a  and  a61233a );
 a61240a <=( A199  and  A166 );
 a61243a <=( A232  and  A200 );
 a61244a <=( a61243a  and  a61240a );
 a61245a <=( a61244a  and  a61237a );
 a61248a <=( A234  and  (not A233) );
 a61251a <=( A265  and  A235 );
 a61252a <=( a61251a  and  a61248a );
 a61255a <=( (not A267)  and  (not A266) );
 a61258a <=( (not A269)  and  (not A268) );
 a61259a <=( a61258a  and  a61255a );
 a61260a <=( a61259a  and  a61252a );
 a61263a <=( (not A169)  and  A170 );
 a61266a <=( (not A167)  and  (not A168) );
 a61267a <=( a61266a  and  a61263a );
 a61270a <=( A199  and  A166 );
 a61273a <=( A232  and  A200 );
 a61274a <=( a61273a  and  a61270a );
 a61275a <=( a61274a  and  a61267a );
 a61278a <=( A234  and  (not A233) );
 a61281a <=( A298  and  A236 );
 a61282a <=( a61281a  and  a61278a );
 a61285a <=( (not A300)  and  (not A299) );
 a61288a <=( (not A302)  and  (not A301) );
 a61289a <=( a61288a  and  a61285a );
 a61290a <=( a61289a  and  a61282a );
 a61293a <=( (not A169)  and  A170 );
 a61296a <=( (not A167)  and  (not A168) );
 a61297a <=( a61296a  and  a61293a );
 a61300a <=( A199  and  A166 );
 a61303a <=( A232  and  A200 );
 a61304a <=( a61303a  and  a61300a );
 a61305a <=( a61304a  and  a61297a );
 a61308a <=( A234  and  (not A233) );
 a61311a <=( (not A298)  and  A236 );
 a61312a <=( a61311a  and  a61308a );
 a61315a <=( (not A300)  and  A299 );
 a61318a <=( (not A302)  and  (not A301) );
 a61319a <=( a61318a  and  a61315a );
 a61320a <=( a61319a  and  a61312a );
 a61323a <=( (not A169)  and  A170 );
 a61326a <=( (not A167)  and  (not A168) );
 a61327a <=( a61326a  and  a61323a );
 a61330a <=( A199  and  A166 );
 a61333a <=( A232  and  A200 );
 a61334a <=( a61333a  and  a61330a );
 a61335a <=( a61334a  and  a61327a );
 a61338a <=( A234  and  (not A233) );
 a61341a <=( (not A265)  and  A236 );
 a61342a <=( a61341a  and  a61338a );
 a61345a <=( (not A267)  and  A266 );
 a61348a <=( (not A269)  and  (not A268) );
 a61349a <=( a61348a  and  a61345a );
 a61350a <=( a61349a  and  a61342a );
 a61353a <=( (not A169)  and  A170 );
 a61356a <=( (not A167)  and  (not A168) );
 a61357a <=( a61356a  and  a61353a );
 a61360a <=( A199  and  A166 );
 a61363a <=( A232  and  A200 );
 a61364a <=( a61363a  and  a61360a );
 a61365a <=( a61364a  and  a61357a );
 a61368a <=( A234  and  (not A233) );
 a61371a <=( A265  and  A236 );
 a61372a <=( a61371a  and  a61368a );
 a61375a <=( (not A267)  and  (not A266) );
 a61378a <=( (not A269)  and  (not A268) );
 a61379a <=( a61378a  and  a61375a );
 a61380a <=( a61379a  and  a61372a );
 a61383a <=( (not A169)  and  A170 );
 a61386a <=( (not A167)  and  (not A168) );
 a61387a <=( a61386a  and  a61383a );
 a61390a <=( A199  and  A166 );
 a61393a <=( A232  and  A200 );
 a61394a <=( a61393a  and  a61390a );
 a61395a <=( a61394a  and  a61387a );
 a61398a <=( (not A234)  and  (not A233) );
 a61401a <=( (not A236)  and  (not A235) );
 a61402a <=( a61401a  and  a61398a );
 a61405a <=( (not A299)  and  A298 );
 a61408a <=( A301  and  A300 );
 a61409a <=( a61408a  and  a61405a );
 a61410a <=( a61409a  and  a61402a );
 a61413a <=( (not A169)  and  A170 );
 a61416a <=( (not A167)  and  (not A168) );
 a61417a <=( a61416a  and  a61413a );
 a61420a <=( A199  and  A166 );
 a61423a <=( A232  and  A200 );
 a61424a <=( a61423a  and  a61420a );
 a61425a <=( a61424a  and  a61417a );
 a61428a <=( (not A234)  and  (not A233) );
 a61431a <=( (not A236)  and  (not A235) );
 a61432a <=( a61431a  and  a61428a );
 a61435a <=( (not A299)  and  A298 );
 a61438a <=( A302  and  A300 );
 a61439a <=( a61438a  and  a61435a );
 a61440a <=( a61439a  and  a61432a );
 a61443a <=( (not A169)  and  A170 );
 a61446a <=( (not A167)  and  (not A168) );
 a61447a <=( a61446a  and  a61443a );
 a61450a <=( A199  and  A166 );
 a61453a <=( A232  and  A200 );
 a61454a <=( a61453a  and  a61450a );
 a61455a <=( a61454a  and  a61447a );
 a61458a <=( (not A234)  and  (not A233) );
 a61461a <=( (not A236)  and  (not A235) );
 a61462a <=( a61461a  and  a61458a );
 a61465a <=( A299  and  (not A298) );
 a61468a <=( A301  and  A300 );
 a61469a <=( a61468a  and  a61465a );
 a61470a <=( a61469a  and  a61462a );
 a61473a <=( (not A169)  and  A170 );
 a61476a <=( (not A167)  and  (not A168) );
 a61477a <=( a61476a  and  a61473a );
 a61480a <=( A199  and  A166 );
 a61483a <=( A232  and  A200 );
 a61484a <=( a61483a  and  a61480a );
 a61485a <=( a61484a  and  a61477a );
 a61488a <=( (not A234)  and  (not A233) );
 a61491a <=( (not A236)  and  (not A235) );
 a61492a <=( a61491a  and  a61488a );
 a61495a <=( A299  and  (not A298) );
 a61498a <=( A302  and  A300 );
 a61499a <=( a61498a  and  a61495a );
 a61500a <=( a61499a  and  a61492a );
 a61503a <=( (not A169)  and  A170 );
 a61506a <=( (not A167)  and  (not A168) );
 a61507a <=( a61506a  and  a61503a );
 a61510a <=( A199  and  A166 );
 a61513a <=( A232  and  A200 );
 a61514a <=( a61513a  and  a61510a );
 a61515a <=( a61514a  and  a61507a );
 a61518a <=( (not A234)  and  (not A233) );
 a61521a <=( (not A236)  and  (not A235) );
 a61522a <=( a61521a  and  a61518a );
 a61525a <=( A266  and  (not A265) );
 a61528a <=( A268  and  A267 );
 a61529a <=( a61528a  and  a61525a );
 a61530a <=( a61529a  and  a61522a );
 a61533a <=( (not A169)  and  A170 );
 a61536a <=( (not A167)  and  (not A168) );
 a61537a <=( a61536a  and  a61533a );
 a61540a <=( A199  and  A166 );
 a61543a <=( A232  and  A200 );
 a61544a <=( a61543a  and  a61540a );
 a61545a <=( a61544a  and  a61537a );
 a61548a <=( (not A234)  and  (not A233) );
 a61551a <=( (not A236)  and  (not A235) );
 a61552a <=( a61551a  and  a61548a );
 a61555a <=( A266  and  (not A265) );
 a61558a <=( A269  and  A267 );
 a61559a <=( a61558a  and  a61555a );
 a61560a <=( a61559a  and  a61552a );
 a61563a <=( (not A169)  and  A170 );
 a61566a <=( (not A167)  and  (not A168) );
 a61567a <=( a61566a  and  a61563a );
 a61570a <=( A199  and  A166 );
 a61573a <=( A232  and  A200 );
 a61574a <=( a61573a  and  a61570a );
 a61575a <=( a61574a  and  a61567a );
 a61578a <=( (not A234)  and  (not A233) );
 a61581a <=( (not A236)  and  (not A235) );
 a61582a <=( a61581a  and  a61578a );
 a61585a <=( (not A266)  and  A265 );
 a61588a <=( A268  and  A267 );
 a61589a <=( a61588a  and  a61585a );
 a61590a <=( a61589a  and  a61582a );
 a61593a <=( (not A169)  and  A170 );
 a61596a <=( (not A167)  and  (not A168) );
 a61597a <=( a61596a  and  a61593a );
 a61600a <=( A199  and  A166 );
 a61603a <=( A232  and  A200 );
 a61604a <=( a61603a  and  a61600a );
 a61605a <=( a61604a  and  a61597a );
 a61608a <=( (not A234)  and  (not A233) );
 a61611a <=( (not A236)  and  (not A235) );
 a61612a <=( a61611a  and  a61608a );
 a61615a <=( (not A266)  and  A265 );
 a61618a <=( A269  and  A267 );
 a61619a <=( a61618a  and  a61615a );
 a61620a <=( a61619a  and  a61612a );
 a61623a <=( (not A169)  and  A170 );
 a61626a <=( (not A167)  and  (not A168) );
 a61627a <=( a61626a  and  a61623a );
 a61630a <=( (not A199)  and  A166 );
 a61633a <=( (not A232)  and  (not A200) );
 a61634a <=( a61633a  and  a61630a );
 a61635a <=( a61634a  and  a61627a );
 a61638a <=( A234  and  A233 );
 a61641a <=( A298  and  A235 );
 a61642a <=( a61641a  and  a61638a );
 a61645a <=( (not A300)  and  (not A299) );
 a61648a <=( (not A302)  and  (not A301) );
 a61649a <=( a61648a  and  a61645a );
 a61650a <=( a61649a  and  a61642a );
 a61653a <=( (not A169)  and  A170 );
 a61656a <=( (not A167)  and  (not A168) );
 a61657a <=( a61656a  and  a61653a );
 a61660a <=( (not A199)  and  A166 );
 a61663a <=( (not A232)  and  (not A200) );
 a61664a <=( a61663a  and  a61660a );
 a61665a <=( a61664a  and  a61657a );
 a61668a <=( A234  and  A233 );
 a61671a <=( (not A298)  and  A235 );
 a61672a <=( a61671a  and  a61668a );
 a61675a <=( (not A300)  and  A299 );
 a61678a <=( (not A302)  and  (not A301) );
 a61679a <=( a61678a  and  a61675a );
 a61680a <=( a61679a  and  a61672a );
 a61683a <=( (not A169)  and  A170 );
 a61686a <=( (not A167)  and  (not A168) );
 a61687a <=( a61686a  and  a61683a );
 a61690a <=( (not A199)  and  A166 );
 a61693a <=( (not A232)  and  (not A200) );
 a61694a <=( a61693a  and  a61690a );
 a61695a <=( a61694a  and  a61687a );
 a61698a <=( A234  and  A233 );
 a61701a <=( (not A265)  and  A235 );
 a61702a <=( a61701a  and  a61698a );
 a61705a <=( (not A267)  and  A266 );
 a61708a <=( (not A269)  and  (not A268) );
 a61709a <=( a61708a  and  a61705a );
 a61710a <=( a61709a  and  a61702a );
 a61713a <=( (not A169)  and  A170 );
 a61716a <=( (not A167)  and  (not A168) );
 a61717a <=( a61716a  and  a61713a );
 a61720a <=( (not A199)  and  A166 );
 a61723a <=( (not A232)  and  (not A200) );
 a61724a <=( a61723a  and  a61720a );
 a61725a <=( a61724a  and  a61717a );
 a61728a <=( A234  and  A233 );
 a61731a <=( A265  and  A235 );
 a61732a <=( a61731a  and  a61728a );
 a61735a <=( (not A267)  and  (not A266) );
 a61738a <=( (not A269)  and  (not A268) );
 a61739a <=( a61738a  and  a61735a );
 a61740a <=( a61739a  and  a61732a );
 a61743a <=( (not A169)  and  A170 );
 a61746a <=( (not A167)  and  (not A168) );
 a61747a <=( a61746a  and  a61743a );
 a61750a <=( (not A199)  and  A166 );
 a61753a <=( (not A232)  and  (not A200) );
 a61754a <=( a61753a  and  a61750a );
 a61755a <=( a61754a  and  a61747a );
 a61758a <=( A234  and  A233 );
 a61761a <=( A298  and  A236 );
 a61762a <=( a61761a  and  a61758a );
 a61765a <=( (not A300)  and  (not A299) );
 a61768a <=( (not A302)  and  (not A301) );
 a61769a <=( a61768a  and  a61765a );
 a61770a <=( a61769a  and  a61762a );
 a61773a <=( (not A169)  and  A170 );
 a61776a <=( (not A167)  and  (not A168) );
 a61777a <=( a61776a  and  a61773a );
 a61780a <=( (not A199)  and  A166 );
 a61783a <=( (not A232)  and  (not A200) );
 a61784a <=( a61783a  and  a61780a );
 a61785a <=( a61784a  and  a61777a );
 a61788a <=( A234  and  A233 );
 a61791a <=( (not A298)  and  A236 );
 a61792a <=( a61791a  and  a61788a );
 a61795a <=( (not A300)  and  A299 );
 a61798a <=( (not A302)  and  (not A301) );
 a61799a <=( a61798a  and  a61795a );
 a61800a <=( a61799a  and  a61792a );
 a61803a <=( (not A169)  and  A170 );
 a61806a <=( (not A167)  and  (not A168) );
 a61807a <=( a61806a  and  a61803a );
 a61810a <=( (not A199)  and  A166 );
 a61813a <=( (not A232)  and  (not A200) );
 a61814a <=( a61813a  and  a61810a );
 a61815a <=( a61814a  and  a61807a );
 a61818a <=( A234  and  A233 );
 a61821a <=( (not A265)  and  A236 );
 a61822a <=( a61821a  and  a61818a );
 a61825a <=( (not A267)  and  A266 );
 a61828a <=( (not A269)  and  (not A268) );
 a61829a <=( a61828a  and  a61825a );
 a61830a <=( a61829a  and  a61822a );
 a61833a <=( (not A169)  and  A170 );
 a61836a <=( (not A167)  and  (not A168) );
 a61837a <=( a61836a  and  a61833a );
 a61840a <=( (not A199)  and  A166 );
 a61843a <=( (not A232)  and  (not A200) );
 a61844a <=( a61843a  and  a61840a );
 a61845a <=( a61844a  and  a61837a );
 a61848a <=( A234  and  A233 );
 a61851a <=( A265  and  A236 );
 a61852a <=( a61851a  and  a61848a );
 a61855a <=( (not A267)  and  (not A266) );
 a61858a <=( (not A269)  and  (not A268) );
 a61859a <=( a61858a  and  a61855a );
 a61860a <=( a61859a  and  a61852a );
 a61863a <=( (not A169)  and  A170 );
 a61866a <=( (not A167)  and  (not A168) );
 a61867a <=( a61866a  and  a61863a );
 a61870a <=( (not A199)  and  A166 );
 a61873a <=( (not A232)  and  (not A200) );
 a61874a <=( a61873a  and  a61870a );
 a61875a <=( a61874a  and  a61867a );
 a61878a <=( (not A234)  and  A233 );
 a61881a <=( (not A236)  and  (not A235) );
 a61882a <=( a61881a  and  a61878a );
 a61885a <=( (not A299)  and  A298 );
 a61888a <=( A301  and  A300 );
 a61889a <=( a61888a  and  a61885a );
 a61890a <=( a61889a  and  a61882a );
 a61893a <=( (not A169)  and  A170 );
 a61896a <=( (not A167)  and  (not A168) );
 a61897a <=( a61896a  and  a61893a );
 a61900a <=( (not A199)  and  A166 );
 a61903a <=( (not A232)  and  (not A200) );
 a61904a <=( a61903a  and  a61900a );
 a61905a <=( a61904a  and  a61897a );
 a61908a <=( (not A234)  and  A233 );
 a61911a <=( (not A236)  and  (not A235) );
 a61912a <=( a61911a  and  a61908a );
 a61915a <=( (not A299)  and  A298 );
 a61918a <=( A302  and  A300 );
 a61919a <=( a61918a  and  a61915a );
 a61920a <=( a61919a  and  a61912a );
 a61923a <=( (not A169)  and  A170 );
 a61926a <=( (not A167)  and  (not A168) );
 a61927a <=( a61926a  and  a61923a );
 a61930a <=( (not A199)  and  A166 );
 a61933a <=( (not A232)  and  (not A200) );
 a61934a <=( a61933a  and  a61930a );
 a61935a <=( a61934a  and  a61927a );
 a61938a <=( (not A234)  and  A233 );
 a61941a <=( (not A236)  and  (not A235) );
 a61942a <=( a61941a  and  a61938a );
 a61945a <=( A299  and  (not A298) );
 a61948a <=( A301  and  A300 );
 a61949a <=( a61948a  and  a61945a );
 a61950a <=( a61949a  and  a61942a );
 a61953a <=( (not A169)  and  A170 );
 a61956a <=( (not A167)  and  (not A168) );
 a61957a <=( a61956a  and  a61953a );
 a61960a <=( (not A199)  and  A166 );
 a61963a <=( (not A232)  and  (not A200) );
 a61964a <=( a61963a  and  a61960a );
 a61965a <=( a61964a  and  a61957a );
 a61968a <=( (not A234)  and  A233 );
 a61971a <=( (not A236)  and  (not A235) );
 a61972a <=( a61971a  and  a61968a );
 a61975a <=( A299  and  (not A298) );
 a61978a <=( A302  and  A300 );
 a61979a <=( a61978a  and  a61975a );
 a61980a <=( a61979a  and  a61972a );
 a61983a <=( (not A169)  and  A170 );
 a61986a <=( (not A167)  and  (not A168) );
 a61987a <=( a61986a  and  a61983a );
 a61990a <=( (not A199)  and  A166 );
 a61993a <=( (not A232)  and  (not A200) );
 a61994a <=( a61993a  and  a61990a );
 a61995a <=( a61994a  and  a61987a );
 a61998a <=( (not A234)  and  A233 );
 a62001a <=( (not A236)  and  (not A235) );
 a62002a <=( a62001a  and  a61998a );
 a62005a <=( A266  and  (not A265) );
 a62008a <=( A268  and  A267 );
 a62009a <=( a62008a  and  a62005a );
 a62010a <=( a62009a  and  a62002a );
 a62013a <=( (not A169)  and  A170 );
 a62016a <=( (not A167)  and  (not A168) );
 a62017a <=( a62016a  and  a62013a );
 a62020a <=( (not A199)  and  A166 );
 a62023a <=( (not A232)  and  (not A200) );
 a62024a <=( a62023a  and  a62020a );
 a62025a <=( a62024a  and  a62017a );
 a62028a <=( (not A234)  and  A233 );
 a62031a <=( (not A236)  and  (not A235) );
 a62032a <=( a62031a  and  a62028a );
 a62035a <=( A266  and  (not A265) );
 a62038a <=( A269  and  A267 );
 a62039a <=( a62038a  and  a62035a );
 a62040a <=( a62039a  and  a62032a );
 a62043a <=( (not A169)  and  A170 );
 a62046a <=( (not A167)  and  (not A168) );
 a62047a <=( a62046a  and  a62043a );
 a62050a <=( (not A199)  and  A166 );
 a62053a <=( (not A232)  and  (not A200) );
 a62054a <=( a62053a  and  a62050a );
 a62055a <=( a62054a  and  a62047a );
 a62058a <=( (not A234)  and  A233 );
 a62061a <=( (not A236)  and  (not A235) );
 a62062a <=( a62061a  and  a62058a );
 a62065a <=( (not A266)  and  A265 );
 a62068a <=( A268  and  A267 );
 a62069a <=( a62068a  and  a62065a );
 a62070a <=( a62069a  and  a62062a );
 a62073a <=( (not A169)  and  A170 );
 a62076a <=( (not A167)  and  (not A168) );
 a62077a <=( a62076a  and  a62073a );
 a62080a <=( (not A199)  and  A166 );
 a62083a <=( (not A232)  and  (not A200) );
 a62084a <=( a62083a  and  a62080a );
 a62085a <=( a62084a  and  a62077a );
 a62088a <=( (not A234)  and  A233 );
 a62091a <=( (not A236)  and  (not A235) );
 a62092a <=( a62091a  and  a62088a );
 a62095a <=( (not A266)  and  A265 );
 a62098a <=( A269  and  A267 );
 a62099a <=( a62098a  and  a62095a );
 a62100a <=( a62099a  and  a62092a );
 a62103a <=( (not A169)  and  A170 );
 a62106a <=( (not A167)  and  (not A168) );
 a62107a <=( a62106a  and  a62103a );
 a62110a <=( (not A199)  and  A166 );
 a62113a <=( A232  and  (not A200) );
 a62114a <=( a62113a  and  a62110a );
 a62115a <=( a62114a  and  a62107a );
 a62118a <=( A234  and  (not A233) );
 a62121a <=( A298  and  A235 );
 a62122a <=( a62121a  and  a62118a );
 a62125a <=( (not A300)  and  (not A299) );
 a62128a <=( (not A302)  and  (not A301) );
 a62129a <=( a62128a  and  a62125a );
 a62130a <=( a62129a  and  a62122a );
 a62133a <=( (not A169)  and  A170 );
 a62136a <=( (not A167)  and  (not A168) );
 a62137a <=( a62136a  and  a62133a );
 a62140a <=( (not A199)  and  A166 );
 a62143a <=( A232  and  (not A200) );
 a62144a <=( a62143a  and  a62140a );
 a62145a <=( a62144a  and  a62137a );
 a62148a <=( A234  and  (not A233) );
 a62151a <=( (not A298)  and  A235 );
 a62152a <=( a62151a  and  a62148a );
 a62155a <=( (not A300)  and  A299 );
 a62158a <=( (not A302)  and  (not A301) );
 a62159a <=( a62158a  and  a62155a );
 a62160a <=( a62159a  and  a62152a );
 a62163a <=( (not A169)  and  A170 );
 a62166a <=( (not A167)  and  (not A168) );
 a62167a <=( a62166a  and  a62163a );
 a62170a <=( (not A199)  and  A166 );
 a62173a <=( A232  and  (not A200) );
 a62174a <=( a62173a  and  a62170a );
 a62175a <=( a62174a  and  a62167a );
 a62178a <=( A234  and  (not A233) );
 a62181a <=( (not A265)  and  A235 );
 a62182a <=( a62181a  and  a62178a );
 a62185a <=( (not A267)  and  A266 );
 a62188a <=( (not A269)  and  (not A268) );
 a62189a <=( a62188a  and  a62185a );
 a62190a <=( a62189a  and  a62182a );
 a62193a <=( (not A169)  and  A170 );
 a62196a <=( (not A167)  and  (not A168) );
 a62197a <=( a62196a  and  a62193a );
 a62200a <=( (not A199)  and  A166 );
 a62203a <=( A232  and  (not A200) );
 a62204a <=( a62203a  and  a62200a );
 a62205a <=( a62204a  and  a62197a );
 a62208a <=( A234  and  (not A233) );
 a62211a <=( A265  and  A235 );
 a62212a <=( a62211a  and  a62208a );
 a62215a <=( (not A267)  and  (not A266) );
 a62218a <=( (not A269)  and  (not A268) );
 a62219a <=( a62218a  and  a62215a );
 a62220a <=( a62219a  and  a62212a );
 a62223a <=( (not A169)  and  A170 );
 a62226a <=( (not A167)  and  (not A168) );
 a62227a <=( a62226a  and  a62223a );
 a62230a <=( (not A199)  and  A166 );
 a62233a <=( A232  and  (not A200) );
 a62234a <=( a62233a  and  a62230a );
 a62235a <=( a62234a  and  a62227a );
 a62238a <=( A234  and  (not A233) );
 a62241a <=( A298  and  A236 );
 a62242a <=( a62241a  and  a62238a );
 a62245a <=( (not A300)  and  (not A299) );
 a62248a <=( (not A302)  and  (not A301) );
 a62249a <=( a62248a  and  a62245a );
 a62250a <=( a62249a  and  a62242a );
 a62253a <=( (not A169)  and  A170 );
 a62256a <=( (not A167)  and  (not A168) );
 a62257a <=( a62256a  and  a62253a );
 a62260a <=( (not A199)  and  A166 );
 a62263a <=( A232  and  (not A200) );
 a62264a <=( a62263a  and  a62260a );
 a62265a <=( a62264a  and  a62257a );
 a62268a <=( A234  and  (not A233) );
 a62271a <=( (not A298)  and  A236 );
 a62272a <=( a62271a  and  a62268a );
 a62275a <=( (not A300)  and  A299 );
 a62278a <=( (not A302)  and  (not A301) );
 a62279a <=( a62278a  and  a62275a );
 a62280a <=( a62279a  and  a62272a );
 a62283a <=( (not A169)  and  A170 );
 a62286a <=( (not A167)  and  (not A168) );
 a62287a <=( a62286a  and  a62283a );
 a62290a <=( (not A199)  and  A166 );
 a62293a <=( A232  and  (not A200) );
 a62294a <=( a62293a  and  a62290a );
 a62295a <=( a62294a  and  a62287a );
 a62298a <=( A234  and  (not A233) );
 a62301a <=( (not A265)  and  A236 );
 a62302a <=( a62301a  and  a62298a );
 a62305a <=( (not A267)  and  A266 );
 a62308a <=( (not A269)  and  (not A268) );
 a62309a <=( a62308a  and  a62305a );
 a62310a <=( a62309a  and  a62302a );
 a62313a <=( (not A169)  and  A170 );
 a62316a <=( (not A167)  and  (not A168) );
 a62317a <=( a62316a  and  a62313a );
 a62320a <=( (not A199)  and  A166 );
 a62323a <=( A232  and  (not A200) );
 a62324a <=( a62323a  and  a62320a );
 a62325a <=( a62324a  and  a62317a );
 a62328a <=( A234  and  (not A233) );
 a62331a <=( A265  and  A236 );
 a62332a <=( a62331a  and  a62328a );
 a62335a <=( (not A267)  and  (not A266) );
 a62338a <=( (not A269)  and  (not A268) );
 a62339a <=( a62338a  and  a62335a );
 a62340a <=( a62339a  and  a62332a );
 a62343a <=( (not A169)  and  A170 );
 a62346a <=( (not A167)  and  (not A168) );
 a62347a <=( a62346a  and  a62343a );
 a62350a <=( (not A199)  and  A166 );
 a62353a <=( A232  and  (not A200) );
 a62354a <=( a62353a  and  a62350a );
 a62355a <=( a62354a  and  a62347a );
 a62358a <=( (not A234)  and  (not A233) );
 a62361a <=( (not A236)  and  (not A235) );
 a62362a <=( a62361a  and  a62358a );
 a62365a <=( (not A299)  and  A298 );
 a62368a <=( A301  and  A300 );
 a62369a <=( a62368a  and  a62365a );
 a62370a <=( a62369a  and  a62362a );
 a62373a <=( (not A169)  and  A170 );
 a62376a <=( (not A167)  and  (not A168) );
 a62377a <=( a62376a  and  a62373a );
 a62380a <=( (not A199)  and  A166 );
 a62383a <=( A232  and  (not A200) );
 a62384a <=( a62383a  and  a62380a );
 a62385a <=( a62384a  and  a62377a );
 a62388a <=( (not A234)  and  (not A233) );
 a62391a <=( (not A236)  and  (not A235) );
 a62392a <=( a62391a  and  a62388a );
 a62395a <=( (not A299)  and  A298 );
 a62398a <=( A302  and  A300 );
 a62399a <=( a62398a  and  a62395a );
 a62400a <=( a62399a  and  a62392a );
 a62403a <=( (not A169)  and  A170 );
 a62406a <=( (not A167)  and  (not A168) );
 a62407a <=( a62406a  and  a62403a );
 a62410a <=( (not A199)  and  A166 );
 a62413a <=( A232  and  (not A200) );
 a62414a <=( a62413a  and  a62410a );
 a62415a <=( a62414a  and  a62407a );
 a62418a <=( (not A234)  and  (not A233) );
 a62421a <=( (not A236)  and  (not A235) );
 a62422a <=( a62421a  and  a62418a );
 a62425a <=( A299  and  (not A298) );
 a62428a <=( A301  and  A300 );
 a62429a <=( a62428a  and  a62425a );
 a62430a <=( a62429a  and  a62422a );
 a62433a <=( (not A169)  and  A170 );
 a62436a <=( (not A167)  and  (not A168) );
 a62437a <=( a62436a  and  a62433a );
 a62440a <=( (not A199)  and  A166 );
 a62443a <=( A232  and  (not A200) );
 a62444a <=( a62443a  and  a62440a );
 a62445a <=( a62444a  and  a62437a );
 a62448a <=( (not A234)  and  (not A233) );
 a62451a <=( (not A236)  and  (not A235) );
 a62452a <=( a62451a  and  a62448a );
 a62455a <=( A299  and  (not A298) );
 a62458a <=( A302  and  A300 );
 a62459a <=( a62458a  and  a62455a );
 a62460a <=( a62459a  and  a62452a );
 a62463a <=( (not A169)  and  A170 );
 a62466a <=( (not A167)  and  (not A168) );
 a62467a <=( a62466a  and  a62463a );
 a62470a <=( (not A199)  and  A166 );
 a62473a <=( A232  and  (not A200) );
 a62474a <=( a62473a  and  a62470a );
 a62475a <=( a62474a  and  a62467a );
 a62478a <=( (not A234)  and  (not A233) );
 a62481a <=( (not A236)  and  (not A235) );
 a62482a <=( a62481a  and  a62478a );
 a62485a <=( A266  and  (not A265) );
 a62488a <=( A268  and  A267 );
 a62489a <=( a62488a  and  a62485a );
 a62490a <=( a62489a  and  a62482a );
 a62493a <=( (not A169)  and  A170 );
 a62496a <=( (not A167)  and  (not A168) );
 a62497a <=( a62496a  and  a62493a );
 a62500a <=( (not A199)  and  A166 );
 a62503a <=( A232  and  (not A200) );
 a62504a <=( a62503a  and  a62500a );
 a62505a <=( a62504a  and  a62497a );
 a62508a <=( (not A234)  and  (not A233) );
 a62511a <=( (not A236)  and  (not A235) );
 a62512a <=( a62511a  and  a62508a );
 a62515a <=( A266  and  (not A265) );
 a62518a <=( A269  and  A267 );
 a62519a <=( a62518a  and  a62515a );
 a62520a <=( a62519a  and  a62512a );
 a62523a <=( (not A169)  and  A170 );
 a62526a <=( (not A167)  and  (not A168) );
 a62527a <=( a62526a  and  a62523a );
 a62530a <=( (not A199)  and  A166 );
 a62533a <=( A232  and  (not A200) );
 a62534a <=( a62533a  and  a62530a );
 a62535a <=( a62534a  and  a62527a );
 a62538a <=( (not A234)  and  (not A233) );
 a62541a <=( (not A236)  and  (not A235) );
 a62542a <=( a62541a  and  a62538a );
 a62545a <=( (not A266)  and  A265 );
 a62548a <=( A268  and  A267 );
 a62549a <=( a62548a  and  a62545a );
 a62550a <=( a62549a  and  a62542a );
 a62553a <=( (not A169)  and  A170 );
 a62556a <=( (not A167)  and  (not A168) );
 a62557a <=( a62556a  and  a62553a );
 a62560a <=( (not A199)  and  A166 );
 a62563a <=( A232  and  (not A200) );
 a62564a <=( a62563a  and  a62560a );
 a62565a <=( a62564a  and  a62557a );
 a62568a <=( (not A234)  and  (not A233) );
 a62571a <=( (not A236)  and  (not A235) );
 a62572a <=( a62571a  and  a62568a );
 a62575a <=( (not A266)  and  A265 );
 a62578a <=( A269  and  A267 );
 a62579a <=( a62578a  and  a62575a );
 a62580a <=( a62579a  and  a62572a );
 a62583a <=( A168  and  (not A170) );
 a62586a <=( (not A166)  and  A167 );
 a62587a <=( a62586a  and  a62583a );
 a62590a <=( (not A202)  and  A201 );
 a62593a <=( (not A232)  and  (not A203) );
 a62594a <=( a62593a  and  a62590a );
 a62595a <=( a62594a  and  a62587a );
 a62598a <=( (not A234)  and  A233 );
 a62601a <=( (not A236)  and  (not A235) );
 a62602a <=( a62601a  and  a62598a );
 a62605a <=( (not A299)  and  A298 );
 a62609a <=( (not A302)  and  (not A301) );
 a62610a <=( (not A300)  and  a62609a );
 a62611a <=( a62610a  and  a62605a );
 a62612a <=( a62611a  and  a62602a );
 a62615a <=( A168  and  (not A170) );
 a62618a <=( (not A166)  and  A167 );
 a62619a <=( a62618a  and  a62615a );
 a62622a <=( (not A202)  and  A201 );
 a62625a <=( (not A232)  and  (not A203) );
 a62626a <=( a62625a  and  a62622a );
 a62627a <=( a62626a  and  a62619a );
 a62630a <=( (not A234)  and  A233 );
 a62633a <=( (not A236)  and  (not A235) );
 a62634a <=( a62633a  and  a62630a );
 a62637a <=( A299  and  (not A298) );
 a62641a <=( (not A302)  and  (not A301) );
 a62642a <=( (not A300)  and  a62641a );
 a62643a <=( a62642a  and  a62637a );
 a62644a <=( a62643a  and  a62634a );
 a62647a <=( A168  and  (not A170) );
 a62650a <=( (not A166)  and  A167 );
 a62651a <=( a62650a  and  a62647a );
 a62654a <=( (not A202)  and  A201 );
 a62657a <=( (not A232)  and  (not A203) );
 a62658a <=( a62657a  and  a62654a );
 a62659a <=( a62658a  and  a62651a );
 a62662a <=( (not A234)  and  A233 );
 a62665a <=( (not A236)  and  (not A235) );
 a62666a <=( a62665a  and  a62662a );
 a62669a <=( A266  and  (not A265) );
 a62673a <=( (not A269)  and  (not A268) );
 a62674a <=( (not A267)  and  a62673a );
 a62675a <=( a62674a  and  a62669a );
 a62676a <=( a62675a  and  a62666a );
 a62679a <=( A168  and  (not A170) );
 a62682a <=( (not A166)  and  A167 );
 a62683a <=( a62682a  and  a62679a );
 a62686a <=( (not A202)  and  A201 );
 a62689a <=( (not A232)  and  (not A203) );
 a62690a <=( a62689a  and  a62686a );
 a62691a <=( a62690a  and  a62683a );
 a62694a <=( (not A234)  and  A233 );
 a62697a <=( (not A236)  and  (not A235) );
 a62698a <=( a62697a  and  a62694a );
 a62701a <=( (not A266)  and  A265 );
 a62705a <=( (not A269)  and  (not A268) );
 a62706a <=( (not A267)  and  a62705a );
 a62707a <=( a62706a  and  a62701a );
 a62708a <=( a62707a  and  a62698a );
 a62711a <=( A168  and  (not A170) );
 a62714a <=( (not A166)  and  A167 );
 a62715a <=( a62714a  and  a62711a );
 a62718a <=( (not A202)  and  A201 );
 a62721a <=( A232  and  (not A203) );
 a62722a <=( a62721a  and  a62718a );
 a62723a <=( a62722a  and  a62715a );
 a62726a <=( (not A234)  and  (not A233) );
 a62729a <=( (not A236)  and  (not A235) );
 a62730a <=( a62729a  and  a62726a );
 a62733a <=( (not A299)  and  A298 );
 a62737a <=( (not A302)  and  (not A301) );
 a62738a <=( (not A300)  and  a62737a );
 a62739a <=( a62738a  and  a62733a );
 a62740a <=( a62739a  and  a62730a );
 a62743a <=( A168  and  (not A170) );
 a62746a <=( (not A166)  and  A167 );
 a62747a <=( a62746a  and  a62743a );
 a62750a <=( (not A202)  and  A201 );
 a62753a <=( A232  and  (not A203) );
 a62754a <=( a62753a  and  a62750a );
 a62755a <=( a62754a  and  a62747a );
 a62758a <=( (not A234)  and  (not A233) );
 a62761a <=( (not A236)  and  (not A235) );
 a62762a <=( a62761a  and  a62758a );
 a62765a <=( A299  and  (not A298) );
 a62769a <=( (not A302)  and  (not A301) );
 a62770a <=( (not A300)  and  a62769a );
 a62771a <=( a62770a  and  a62765a );
 a62772a <=( a62771a  and  a62762a );
 a62775a <=( A168  and  (not A170) );
 a62778a <=( (not A166)  and  A167 );
 a62779a <=( a62778a  and  a62775a );
 a62782a <=( (not A202)  and  A201 );
 a62785a <=( A232  and  (not A203) );
 a62786a <=( a62785a  and  a62782a );
 a62787a <=( a62786a  and  a62779a );
 a62790a <=( (not A234)  and  (not A233) );
 a62793a <=( (not A236)  and  (not A235) );
 a62794a <=( a62793a  and  a62790a );
 a62797a <=( A266  and  (not A265) );
 a62801a <=( (not A269)  and  (not A268) );
 a62802a <=( (not A267)  and  a62801a );
 a62803a <=( a62802a  and  a62797a );
 a62804a <=( a62803a  and  a62794a );
 a62807a <=( A168  and  (not A170) );
 a62810a <=( (not A166)  and  A167 );
 a62811a <=( a62810a  and  a62807a );
 a62814a <=( (not A202)  and  A201 );
 a62817a <=( A232  and  (not A203) );
 a62818a <=( a62817a  and  a62814a );
 a62819a <=( a62818a  and  a62811a );
 a62822a <=( (not A234)  and  (not A233) );
 a62825a <=( (not A236)  and  (not A235) );
 a62826a <=( a62825a  and  a62822a );
 a62829a <=( (not A266)  and  A265 );
 a62833a <=( (not A269)  and  (not A268) );
 a62834a <=( (not A267)  and  a62833a );
 a62835a <=( a62834a  and  a62829a );
 a62836a <=( a62835a  and  a62826a );
 a62839a <=( A168  and  (not A170) );
 a62842a <=( A166  and  (not A167) );
 a62843a <=( a62842a  and  a62839a );
 a62846a <=( (not A202)  and  A201 );
 a62849a <=( (not A232)  and  (not A203) );
 a62850a <=( a62849a  and  a62846a );
 a62851a <=( a62850a  and  a62843a );
 a62854a <=( (not A234)  and  A233 );
 a62857a <=( (not A236)  and  (not A235) );
 a62858a <=( a62857a  and  a62854a );
 a62861a <=( (not A299)  and  A298 );
 a62865a <=( (not A302)  and  (not A301) );
 a62866a <=( (not A300)  and  a62865a );
 a62867a <=( a62866a  and  a62861a );
 a62868a <=( a62867a  and  a62858a );
 a62871a <=( A168  and  (not A170) );
 a62874a <=( A166  and  (not A167) );
 a62875a <=( a62874a  and  a62871a );
 a62878a <=( (not A202)  and  A201 );
 a62881a <=( (not A232)  and  (not A203) );
 a62882a <=( a62881a  and  a62878a );
 a62883a <=( a62882a  and  a62875a );
 a62886a <=( (not A234)  and  A233 );
 a62889a <=( (not A236)  and  (not A235) );
 a62890a <=( a62889a  and  a62886a );
 a62893a <=( A299  and  (not A298) );
 a62897a <=( (not A302)  and  (not A301) );
 a62898a <=( (not A300)  and  a62897a );
 a62899a <=( a62898a  and  a62893a );
 a62900a <=( a62899a  and  a62890a );
 a62903a <=( A168  and  (not A170) );
 a62906a <=( A166  and  (not A167) );
 a62907a <=( a62906a  and  a62903a );
 a62910a <=( (not A202)  and  A201 );
 a62913a <=( (not A232)  and  (not A203) );
 a62914a <=( a62913a  and  a62910a );
 a62915a <=( a62914a  and  a62907a );
 a62918a <=( (not A234)  and  A233 );
 a62921a <=( (not A236)  and  (not A235) );
 a62922a <=( a62921a  and  a62918a );
 a62925a <=( A266  and  (not A265) );
 a62929a <=( (not A269)  and  (not A268) );
 a62930a <=( (not A267)  and  a62929a );
 a62931a <=( a62930a  and  a62925a );
 a62932a <=( a62931a  and  a62922a );
 a62935a <=( A168  and  (not A170) );
 a62938a <=( A166  and  (not A167) );
 a62939a <=( a62938a  and  a62935a );
 a62942a <=( (not A202)  and  A201 );
 a62945a <=( (not A232)  and  (not A203) );
 a62946a <=( a62945a  and  a62942a );
 a62947a <=( a62946a  and  a62939a );
 a62950a <=( (not A234)  and  A233 );
 a62953a <=( (not A236)  and  (not A235) );
 a62954a <=( a62953a  and  a62950a );
 a62957a <=( (not A266)  and  A265 );
 a62961a <=( (not A269)  and  (not A268) );
 a62962a <=( (not A267)  and  a62961a );
 a62963a <=( a62962a  and  a62957a );
 a62964a <=( a62963a  and  a62954a );
 a62967a <=( A168  and  (not A170) );
 a62970a <=( A166  and  (not A167) );
 a62971a <=( a62970a  and  a62967a );
 a62974a <=( (not A202)  and  A201 );
 a62977a <=( A232  and  (not A203) );
 a62978a <=( a62977a  and  a62974a );
 a62979a <=( a62978a  and  a62971a );
 a62982a <=( (not A234)  and  (not A233) );
 a62985a <=( (not A236)  and  (not A235) );
 a62986a <=( a62985a  and  a62982a );
 a62989a <=( (not A299)  and  A298 );
 a62993a <=( (not A302)  and  (not A301) );
 a62994a <=( (not A300)  and  a62993a );
 a62995a <=( a62994a  and  a62989a );
 a62996a <=( a62995a  and  a62986a );
 a62999a <=( A168  and  (not A170) );
 a63002a <=( A166  and  (not A167) );
 a63003a <=( a63002a  and  a62999a );
 a63006a <=( (not A202)  and  A201 );
 a63009a <=( A232  and  (not A203) );
 a63010a <=( a63009a  and  a63006a );
 a63011a <=( a63010a  and  a63003a );
 a63014a <=( (not A234)  and  (not A233) );
 a63017a <=( (not A236)  and  (not A235) );
 a63018a <=( a63017a  and  a63014a );
 a63021a <=( A299  and  (not A298) );
 a63025a <=( (not A302)  and  (not A301) );
 a63026a <=( (not A300)  and  a63025a );
 a63027a <=( a63026a  and  a63021a );
 a63028a <=( a63027a  and  a63018a );
 a63031a <=( A168  and  (not A170) );
 a63034a <=( A166  and  (not A167) );
 a63035a <=( a63034a  and  a63031a );
 a63038a <=( (not A202)  and  A201 );
 a63041a <=( A232  and  (not A203) );
 a63042a <=( a63041a  and  a63038a );
 a63043a <=( a63042a  and  a63035a );
 a63046a <=( (not A234)  and  (not A233) );
 a63049a <=( (not A236)  and  (not A235) );
 a63050a <=( a63049a  and  a63046a );
 a63053a <=( A266  and  (not A265) );
 a63057a <=( (not A269)  and  (not A268) );
 a63058a <=( (not A267)  and  a63057a );
 a63059a <=( a63058a  and  a63053a );
 a63060a <=( a63059a  and  a63050a );
 a63063a <=( A168  and  (not A170) );
 a63066a <=( A166  and  (not A167) );
 a63067a <=( a63066a  and  a63063a );
 a63070a <=( (not A202)  and  A201 );
 a63073a <=( A232  and  (not A203) );
 a63074a <=( a63073a  and  a63070a );
 a63075a <=( a63074a  and  a63067a );
 a63078a <=( (not A234)  and  (not A233) );
 a63081a <=( (not A236)  and  (not A235) );
 a63082a <=( a63081a  and  a63078a );
 a63085a <=( (not A266)  and  A265 );
 a63089a <=( (not A269)  and  (not A268) );
 a63090a <=( (not A267)  and  a63089a );
 a63091a <=( a63090a  and  a63085a );
 a63092a <=( a63091a  and  a63082a );
 a63095a <=( A168  and  A169 );
 a63098a <=( (not A166)  and  A167 );
 a63099a <=( a63098a  and  a63095a );
 a63102a <=( (not A202)  and  A201 );
 a63105a <=( (not A232)  and  (not A203) );
 a63106a <=( a63105a  and  a63102a );
 a63107a <=( a63106a  and  a63099a );
 a63110a <=( (not A234)  and  A233 );
 a63113a <=( (not A236)  and  (not A235) );
 a63114a <=( a63113a  and  a63110a );
 a63117a <=( (not A299)  and  A298 );
 a63121a <=( (not A302)  and  (not A301) );
 a63122a <=( (not A300)  and  a63121a );
 a63123a <=( a63122a  and  a63117a );
 a63124a <=( a63123a  and  a63114a );
 a63127a <=( A168  and  A169 );
 a63130a <=( (not A166)  and  A167 );
 a63131a <=( a63130a  and  a63127a );
 a63134a <=( (not A202)  and  A201 );
 a63137a <=( (not A232)  and  (not A203) );
 a63138a <=( a63137a  and  a63134a );
 a63139a <=( a63138a  and  a63131a );
 a63142a <=( (not A234)  and  A233 );
 a63145a <=( (not A236)  and  (not A235) );
 a63146a <=( a63145a  and  a63142a );
 a63149a <=( A299  and  (not A298) );
 a63153a <=( (not A302)  and  (not A301) );
 a63154a <=( (not A300)  and  a63153a );
 a63155a <=( a63154a  and  a63149a );
 a63156a <=( a63155a  and  a63146a );
 a63159a <=( A168  and  A169 );
 a63162a <=( (not A166)  and  A167 );
 a63163a <=( a63162a  and  a63159a );
 a63166a <=( (not A202)  and  A201 );
 a63169a <=( (not A232)  and  (not A203) );
 a63170a <=( a63169a  and  a63166a );
 a63171a <=( a63170a  and  a63163a );
 a63174a <=( (not A234)  and  A233 );
 a63177a <=( (not A236)  and  (not A235) );
 a63178a <=( a63177a  and  a63174a );
 a63181a <=( A266  and  (not A265) );
 a63185a <=( (not A269)  and  (not A268) );
 a63186a <=( (not A267)  and  a63185a );
 a63187a <=( a63186a  and  a63181a );
 a63188a <=( a63187a  and  a63178a );
 a63191a <=( A168  and  A169 );
 a63194a <=( (not A166)  and  A167 );
 a63195a <=( a63194a  and  a63191a );
 a63198a <=( (not A202)  and  A201 );
 a63201a <=( (not A232)  and  (not A203) );
 a63202a <=( a63201a  and  a63198a );
 a63203a <=( a63202a  and  a63195a );
 a63206a <=( (not A234)  and  A233 );
 a63209a <=( (not A236)  and  (not A235) );
 a63210a <=( a63209a  and  a63206a );
 a63213a <=( (not A266)  and  A265 );
 a63217a <=( (not A269)  and  (not A268) );
 a63218a <=( (not A267)  and  a63217a );
 a63219a <=( a63218a  and  a63213a );
 a63220a <=( a63219a  and  a63210a );
 a63223a <=( A168  and  A169 );
 a63226a <=( (not A166)  and  A167 );
 a63227a <=( a63226a  and  a63223a );
 a63230a <=( (not A202)  and  A201 );
 a63233a <=( A232  and  (not A203) );
 a63234a <=( a63233a  and  a63230a );
 a63235a <=( a63234a  and  a63227a );
 a63238a <=( (not A234)  and  (not A233) );
 a63241a <=( (not A236)  and  (not A235) );
 a63242a <=( a63241a  and  a63238a );
 a63245a <=( (not A299)  and  A298 );
 a63249a <=( (not A302)  and  (not A301) );
 a63250a <=( (not A300)  and  a63249a );
 a63251a <=( a63250a  and  a63245a );
 a63252a <=( a63251a  and  a63242a );
 a63255a <=( A168  and  A169 );
 a63258a <=( (not A166)  and  A167 );
 a63259a <=( a63258a  and  a63255a );
 a63262a <=( (not A202)  and  A201 );
 a63265a <=( A232  and  (not A203) );
 a63266a <=( a63265a  and  a63262a );
 a63267a <=( a63266a  and  a63259a );
 a63270a <=( (not A234)  and  (not A233) );
 a63273a <=( (not A236)  and  (not A235) );
 a63274a <=( a63273a  and  a63270a );
 a63277a <=( A299  and  (not A298) );
 a63281a <=( (not A302)  and  (not A301) );
 a63282a <=( (not A300)  and  a63281a );
 a63283a <=( a63282a  and  a63277a );
 a63284a <=( a63283a  and  a63274a );
 a63287a <=( A168  and  A169 );
 a63290a <=( (not A166)  and  A167 );
 a63291a <=( a63290a  and  a63287a );
 a63294a <=( (not A202)  and  A201 );
 a63297a <=( A232  and  (not A203) );
 a63298a <=( a63297a  and  a63294a );
 a63299a <=( a63298a  and  a63291a );
 a63302a <=( (not A234)  and  (not A233) );
 a63305a <=( (not A236)  and  (not A235) );
 a63306a <=( a63305a  and  a63302a );
 a63309a <=( A266  and  (not A265) );
 a63313a <=( (not A269)  and  (not A268) );
 a63314a <=( (not A267)  and  a63313a );
 a63315a <=( a63314a  and  a63309a );
 a63316a <=( a63315a  and  a63306a );
 a63319a <=( A168  and  A169 );
 a63322a <=( (not A166)  and  A167 );
 a63323a <=( a63322a  and  a63319a );
 a63326a <=( (not A202)  and  A201 );
 a63329a <=( A232  and  (not A203) );
 a63330a <=( a63329a  and  a63326a );
 a63331a <=( a63330a  and  a63323a );
 a63334a <=( (not A234)  and  (not A233) );
 a63337a <=( (not A236)  and  (not A235) );
 a63338a <=( a63337a  and  a63334a );
 a63341a <=( (not A266)  and  A265 );
 a63345a <=( (not A269)  and  (not A268) );
 a63346a <=( (not A267)  and  a63345a );
 a63347a <=( a63346a  and  a63341a );
 a63348a <=( a63347a  and  a63338a );
 a63351a <=( A168  and  A169 );
 a63354a <=( A166  and  (not A167) );
 a63355a <=( a63354a  and  a63351a );
 a63358a <=( (not A202)  and  A201 );
 a63361a <=( (not A232)  and  (not A203) );
 a63362a <=( a63361a  and  a63358a );
 a63363a <=( a63362a  and  a63355a );
 a63366a <=( (not A234)  and  A233 );
 a63369a <=( (not A236)  and  (not A235) );
 a63370a <=( a63369a  and  a63366a );
 a63373a <=( (not A299)  and  A298 );
 a63377a <=( (not A302)  and  (not A301) );
 a63378a <=( (not A300)  and  a63377a );
 a63379a <=( a63378a  and  a63373a );
 a63380a <=( a63379a  and  a63370a );
 a63383a <=( A168  and  A169 );
 a63386a <=( A166  and  (not A167) );
 a63387a <=( a63386a  and  a63383a );
 a63390a <=( (not A202)  and  A201 );
 a63393a <=( (not A232)  and  (not A203) );
 a63394a <=( a63393a  and  a63390a );
 a63395a <=( a63394a  and  a63387a );
 a63398a <=( (not A234)  and  A233 );
 a63401a <=( (not A236)  and  (not A235) );
 a63402a <=( a63401a  and  a63398a );
 a63405a <=( A299  and  (not A298) );
 a63409a <=( (not A302)  and  (not A301) );
 a63410a <=( (not A300)  and  a63409a );
 a63411a <=( a63410a  and  a63405a );
 a63412a <=( a63411a  and  a63402a );
 a63415a <=( A168  and  A169 );
 a63418a <=( A166  and  (not A167) );
 a63419a <=( a63418a  and  a63415a );
 a63422a <=( (not A202)  and  A201 );
 a63425a <=( (not A232)  and  (not A203) );
 a63426a <=( a63425a  and  a63422a );
 a63427a <=( a63426a  and  a63419a );
 a63430a <=( (not A234)  and  A233 );
 a63433a <=( (not A236)  and  (not A235) );
 a63434a <=( a63433a  and  a63430a );
 a63437a <=( A266  and  (not A265) );
 a63441a <=( (not A269)  and  (not A268) );
 a63442a <=( (not A267)  and  a63441a );
 a63443a <=( a63442a  and  a63437a );
 a63444a <=( a63443a  and  a63434a );
 a63447a <=( A168  and  A169 );
 a63450a <=( A166  and  (not A167) );
 a63451a <=( a63450a  and  a63447a );
 a63454a <=( (not A202)  and  A201 );
 a63457a <=( (not A232)  and  (not A203) );
 a63458a <=( a63457a  and  a63454a );
 a63459a <=( a63458a  and  a63451a );
 a63462a <=( (not A234)  and  A233 );
 a63465a <=( (not A236)  and  (not A235) );
 a63466a <=( a63465a  and  a63462a );
 a63469a <=( (not A266)  and  A265 );
 a63473a <=( (not A269)  and  (not A268) );
 a63474a <=( (not A267)  and  a63473a );
 a63475a <=( a63474a  and  a63469a );
 a63476a <=( a63475a  and  a63466a );
 a63479a <=( A168  and  A169 );
 a63482a <=( A166  and  (not A167) );
 a63483a <=( a63482a  and  a63479a );
 a63486a <=( (not A202)  and  A201 );
 a63489a <=( A232  and  (not A203) );
 a63490a <=( a63489a  and  a63486a );
 a63491a <=( a63490a  and  a63483a );
 a63494a <=( (not A234)  and  (not A233) );
 a63497a <=( (not A236)  and  (not A235) );
 a63498a <=( a63497a  and  a63494a );
 a63501a <=( (not A299)  and  A298 );
 a63505a <=( (not A302)  and  (not A301) );
 a63506a <=( (not A300)  and  a63505a );
 a63507a <=( a63506a  and  a63501a );
 a63508a <=( a63507a  and  a63498a );
 a63511a <=( A168  and  A169 );
 a63514a <=( A166  and  (not A167) );
 a63515a <=( a63514a  and  a63511a );
 a63518a <=( (not A202)  and  A201 );
 a63521a <=( A232  and  (not A203) );
 a63522a <=( a63521a  and  a63518a );
 a63523a <=( a63522a  and  a63515a );
 a63526a <=( (not A234)  and  (not A233) );
 a63529a <=( (not A236)  and  (not A235) );
 a63530a <=( a63529a  and  a63526a );
 a63533a <=( A299  and  (not A298) );
 a63537a <=( (not A302)  and  (not A301) );
 a63538a <=( (not A300)  and  a63537a );
 a63539a <=( a63538a  and  a63533a );
 a63540a <=( a63539a  and  a63530a );
 a63543a <=( A168  and  A169 );
 a63546a <=( A166  and  (not A167) );
 a63547a <=( a63546a  and  a63543a );
 a63550a <=( (not A202)  and  A201 );
 a63553a <=( A232  and  (not A203) );
 a63554a <=( a63553a  and  a63550a );
 a63555a <=( a63554a  and  a63547a );
 a63558a <=( (not A234)  and  (not A233) );
 a63561a <=( (not A236)  and  (not A235) );
 a63562a <=( a63561a  and  a63558a );
 a63565a <=( A266  and  (not A265) );
 a63569a <=( (not A269)  and  (not A268) );
 a63570a <=( (not A267)  and  a63569a );
 a63571a <=( a63570a  and  a63565a );
 a63572a <=( a63571a  and  a63562a );
 a63575a <=( A168  and  A169 );
 a63578a <=( A166  and  (not A167) );
 a63579a <=( a63578a  and  a63575a );
 a63582a <=( (not A202)  and  A201 );
 a63585a <=( A232  and  (not A203) );
 a63586a <=( a63585a  and  a63582a );
 a63587a <=( a63586a  and  a63579a );
 a63590a <=( (not A234)  and  (not A233) );
 a63593a <=( (not A236)  and  (not A235) );
 a63594a <=( a63593a  and  a63590a );
 a63597a <=( (not A266)  and  A265 );
 a63601a <=( (not A269)  and  (not A268) );
 a63602a <=( (not A267)  and  a63601a );
 a63603a <=( a63602a  and  a63597a );
 a63604a <=( a63603a  and  a63594a );
 a63607a <=( (not A169)  and  A170 );
 a63610a <=( A167  and  (not A168) );
 a63611a <=( a63610a  and  a63607a );
 a63614a <=( A201  and  (not A166) );
 a63617a <=( (not A203)  and  (not A202) );
 a63618a <=( a63617a  and  a63614a );
 a63619a <=( a63618a  and  a63611a );
 a63622a <=( A233  and  (not A232) );
 a63625a <=( A235  and  A234 );
 a63626a <=( a63625a  and  a63622a );
 a63629a <=( (not A299)  and  A298 );
 a63633a <=( (not A302)  and  (not A301) );
 a63634a <=( (not A300)  and  a63633a );
 a63635a <=( a63634a  and  a63629a );
 a63636a <=( a63635a  and  a63626a );
 a63639a <=( (not A169)  and  A170 );
 a63642a <=( A167  and  (not A168) );
 a63643a <=( a63642a  and  a63639a );
 a63646a <=( A201  and  (not A166) );
 a63649a <=( (not A203)  and  (not A202) );
 a63650a <=( a63649a  and  a63646a );
 a63651a <=( a63650a  and  a63643a );
 a63654a <=( A233  and  (not A232) );
 a63657a <=( A235  and  A234 );
 a63658a <=( a63657a  and  a63654a );
 a63661a <=( A299  and  (not A298) );
 a63665a <=( (not A302)  and  (not A301) );
 a63666a <=( (not A300)  and  a63665a );
 a63667a <=( a63666a  and  a63661a );
 a63668a <=( a63667a  and  a63658a );
 a63671a <=( (not A169)  and  A170 );
 a63674a <=( A167  and  (not A168) );
 a63675a <=( a63674a  and  a63671a );
 a63678a <=( A201  and  (not A166) );
 a63681a <=( (not A203)  and  (not A202) );
 a63682a <=( a63681a  and  a63678a );
 a63683a <=( a63682a  and  a63675a );
 a63686a <=( A233  and  (not A232) );
 a63689a <=( A235  and  A234 );
 a63690a <=( a63689a  and  a63686a );
 a63693a <=( A266  and  (not A265) );
 a63697a <=( (not A269)  and  (not A268) );
 a63698a <=( (not A267)  and  a63697a );
 a63699a <=( a63698a  and  a63693a );
 a63700a <=( a63699a  and  a63690a );
 a63703a <=( (not A169)  and  A170 );
 a63706a <=( A167  and  (not A168) );
 a63707a <=( a63706a  and  a63703a );
 a63710a <=( A201  and  (not A166) );
 a63713a <=( (not A203)  and  (not A202) );
 a63714a <=( a63713a  and  a63710a );
 a63715a <=( a63714a  and  a63707a );
 a63718a <=( A233  and  (not A232) );
 a63721a <=( A235  and  A234 );
 a63722a <=( a63721a  and  a63718a );
 a63725a <=( (not A266)  and  A265 );
 a63729a <=( (not A269)  and  (not A268) );
 a63730a <=( (not A267)  and  a63729a );
 a63731a <=( a63730a  and  a63725a );
 a63732a <=( a63731a  and  a63722a );
 a63735a <=( (not A169)  and  A170 );
 a63738a <=( A167  and  (not A168) );
 a63739a <=( a63738a  and  a63735a );
 a63742a <=( A201  and  (not A166) );
 a63745a <=( (not A203)  and  (not A202) );
 a63746a <=( a63745a  and  a63742a );
 a63747a <=( a63746a  and  a63739a );
 a63750a <=( A233  and  (not A232) );
 a63753a <=( A236  and  A234 );
 a63754a <=( a63753a  and  a63750a );
 a63757a <=( (not A299)  and  A298 );
 a63761a <=( (not A302)  and  (not A301) );
 a63762a <=( (not A300)  and  a63761a );
 a63763a <=( a63762a  and  a63757a );
 a63764a <=( a63763a  and  a63754a );
 a63767a <=( (not A169)  and  A170 );
 a63770a <=( A167  and  (not A168) );
 a63771a <=( a63770a  and  a63767a );
 a63774a <=( A201  and  (not A166) );
 a63777a <=( (not A203)  and  (not A202) );
 a63778a <=( a63777a  and  a63774a );
 a63779a <=( a63778a  and  a63771a );
 a63782a <=( A233  and  (not A232) );
 a63785a <=( A236  and  A234 );
 a63786a <=( a63785a  and  a63782a );
 a63789a <=( A299  and  (not A298) );
 a63793a <=( (not A302)  and  (not A301) );
 a63794a <=( (not A300)  and  a63793a );
 a63795a <=( a63794a  and  a63789a );
 a63796a <=( a63795a  and  a63786a );
 a63799a <=( (not A169)  and  A170 );
 a63802a <=( A167  and  (not A168) );
 a63803a <=( a63802a  and  a63799a );
 a63806a <=( A201  and  (not A166) );
 a63809a <=( (not A203)  and  (not A202) );
 a63810a <=( a63809a  and  a63806a );
 a63811a <=( a63810a  and  a63803a );
 a63814a <=( A233  and  (not A232) );
 a63817a <=( A236  and  A234 );
 a63818a <=( a63817a  and  a63814a );
 a63821a <=( A266  and  (not A265) );
 a63825a <=( (not A269)  and  (not A268) );
 a63826a <=( (not A267)  and  a63825a );
 a63827a <=( a63826a  and  a63821a );
 a63828a <=( a63827a  and  a63818a );
 a63831a <=( (not A169)  and  A170 );
 a63834a <=( A167  and  (not A168) );
 a63835a <=( a63834a  and  a63831a );
 a63838a <=( A201  and  (not A166) );
 a63841a <=( (not A203)  and  (not A202) );
 a63842a <=( a63841a  and  a63838a );
 a63843a <=( a63842a  and  a63835a );
 a63846a <=( A233  and  (not A232) );
 a63849a <=( A236  and  A234 );
 a63850a <=( a63849a  and  a63846a );
 a63853a <=( (not A266)  and  A265 );
 a63857a <=( (not A269)  and  (not A268) );
 a63858a <=( (not A267)  and  a63857a );
 a63859a <=( a63858a  and  a63853a );
 a63860a <=( a63859a  and  a63850a );
 a63863a <=( (not A169)  and  A170 );
 a63866a <=( A167  and  (not A168) );
 a63867a <=( a63866a  and  a63863a );
 a63870a <=( A201  and  (not A166) );
 a63873a <=( (not A203)  and  (not A202) );
 a63874a <=( a63873a  and  a63870a );
 a63875a <=( a63874a  and  a63867a );
 a63878a <=( A233  and  (not A232) );
 a63881a <=( (not A235)  and  (not A234) );
 a63882a <=( a63881a  and  a63878a );
 a63885a <=( A298  and  (not A236) );
 a63889a <=( A301  and  A300 );
 a63890a <=( (not A299)  and  a63889a );
 a63891a <=( a63890a  and  a63885a );
 a63892a <=( a63891a  and  a63882a );
 a63895a <=( (not A169)  and  A170 );
 a63898a <=( A167  and  (not A168) );
 a63899a <=( a63898a  and  a63895a );
 a63902a <=( A201  and  (not A166) );
 a63905a <=( (not A203)  and  (not A202) );
 a63906a <=( a63905a  and  a63902a );
 a63907a <=( a63906a  and  a63899a );
 a63910a <=( A233  and  (not A232) );
 a63913a <=( (not A235)  and  (not A234) );
 a63914a <=( a63913a  and  a63910a );
 a63917a <=( A298  and  (not A236) );
 a63921a <=( A302  and  A300 );
 a63922a <=( (not A299)  and  a63921a );
 a63923a <=( a63922a  and  a63917a );
 a63924a <=( a63923a  and  a63914a );
 a63927a <=( (not A169)  and  A170 );
 a63930a <=( A167  and  (not A168) );
 a63931a <=( a63930a  and  a63927a );
 a63934a <=( A201  and  (not A166) );
 a63937a <=( (not A203)  and  (not A202) );
 a63938a <=( a63937a  and  a63934a );
 a63939a <=( a63938a  and  a63931a );
 a63942a <=( A233  and  (not A232) );
 a63945a <=( (not A235)  and  (not A234) );
 a63946a <=( a63945a  and  a63942a );
 a63949a <=( (not A298)  and  (not A236) );
 a63953a <=( A301  and  A300 );
 a63954a <=( A299  and  a63953a );
 a63955a <=( a63954a  and  a63949a );
 a63956a <=( a63955a  and  a63946a );
 a63959a <=( (not A169)  and  A170 );
 a63962a <=( A167  and  (not A168) );
 a63963a <=( a63962a  and  a63959a );
 a63966a <=( A201  and  (not A166) );
 a63969a <=( (not A203)  and  (not A202) );
 a63970a <=( a63969a  and  a63966a );
 a63971a <=( a63970a  and  a63963a );
 a63974a <=( A233  and  (not A232) );
 a63977a <=( (not A235)  and  (not A234) );
 a63978a <=( a63977a  and  a63974a );
 a63981a <=( (not A298)  and  (not A236) );
 a63985a <=( A302  and  A300 );
 a63986a <=( A299  and  a63985a );
 a63987a <=( a63986a  and  a63981a );
 a63988a <=( a63987a  and  a63978a );
 a63991a <=( (not A169)  and  A170 );
 a63994a <=( A167  and  (not A168) );
 a63995a <=( a63994a  and  a63991a );
 a63998a <=( A201  and  (not A166) );
 a64001a <=( (not A203)  and  (not A202) );
 a64002a <=( a64001a  and  a63998a );
 a64003a <=( a64002a  and  a63995a );
 a64006a <=( A233  and  (not A232) );
 a64009a <=( (not A235)  and  (not A234) );
 a64010a <=( a64009a  and  a64006a );
 a64013a <=( (not A265)  and  (not A236) );
 a64017a <=( A268  and  A267 );
 a64018a <=( A266  and  a64017a );
 a64019a <=( a64018a  and  a64013a );
 a64020a <=( a64019a  and  a64010a );
 a64023a <=( (not A169)  and  A170 );
 a64026a <=( A167  and  (not A168) );
 a64027a <=( a64026a  and  a64023a );
 a64030a <=( A201  and  (not A166) );
 a64033a <=( (not A203)  and  (not A202) );
 a64034a <=( a64033a  and  a64030a );
 a64035a <=( a64034a  and  a64027a );
 a64038a <=( A233  and  (not A232) );
 a64041a <=( (not A235)  and  (not A234) );
 a64042a <=( a64041a  and  a64038a );
 a64045a <=( (not A265)  and  (not A236) );
 a64049a <=( A269  and  A267 );
 a64050a <=( A266  and  a64049a );
 a64051a <=( a64050a  and  a64045a );
 a64052a <=( a64051a  and  a64042a );
 a64055a <=( (not A169)  and  A170 );
 a64058a <=( A167  and  (not A168) );
 a64059a <=( a64058a  and  a64055a );
 a64062a <=( A201  and  (not A166) );
 a64065a <=( (not A203)  and  (not A202) );
 a64066a <=( a64065a  and  a64062a );
 a64067a <=( a64066a  and  a64059a );
 a64070a <=( A233  and  (not A232) );
 a64073a <=( (not A235)  and  (not A234) );
 a64074a <=( a64073a  and  a64070a );
 a64077a <=( A265  and  (not A236) );
 a64081a <=( A268  and  A267 );
 a64082a <=( (not A266)  and  a64081a );
 a64083a <=( a64082a  and  a64077a );
 a64084a <=( a64083a  and  a64074a );
 a64087a <=( (not A169)  and  A170 );
 a64090a <=( A167  and  (not A168) );
 a64091a <=( a64090a  and  a64087a );
 a64094a <=( A201  and  (not A166) );
 a64097a <=( (not A203)  and  (not A202) );
 a64098a <=( a64097a  and  a64094a );
 a64099a <=( a64098a  and  a64091a );
 a64102a <=( A233  and  (not A232) );
 a64105a <=( (not A235)  and  (not A234) );
 a64106a <=( a64105a  and  a64102a );
 a64109a <=( A265  and  (not A236) );
 a64113a <=( A269  and  A267 );
 a64114a <=( (not A266)  and  a64113a );
 a64115a <=( a64114a  and  a64109a );
 a64116a <=( a64115a  and  a64106a );
 a64119a <=( (not A169)  and  A170 );
 a64122a <=( A167  and  (not A168) );
 a64123a <=( a64122a  and  a64119a );
 a64126a <=( A201  and  (not A166) );
 a64129a <=( (not A203)  and  (not A202) );
 a64130a <=( a64129a  and  a64126a );
 a64131a <=( a64130a  and  a64123a );
 a64134a <=( (not A233)  and  A232 );
 a64137a <=( A235  and  A234 );
 a64138a <=( a64137a  and  a64134a );
 a64141a <=( (not A299)  and  A298 );
 a64145a <=( (not A302)  and  (not A301) );
 a64146a <=( (not A300)  and  a64145a );
 a64147a <=( a64146a  and  a64141a );
 a64148a <=( a64147a  and  a64138a );
 a64151a <=( (not A169)  and  A170 );
 a64154a <=( A167  and  (not A168) );
 a64155a <=( a64154a  and  a64151a );
 a64158a <=( A201  and  (not A166) );
 a64161a <=( (not A203)  and  (not A202) );
 a64162a <=( a64161a  and  a64158a );
 a64163a <=( a64162a  and  a64155a );
 a64166a <=( (not A233)  and  A232 );
 a64169a <=( A235  and  A234 );
 a64170a <=( a64169a  and  a64166a );
 a64173a <=( A299  and  (not A298) );
 a64177a <=( (not A302)  and  (not A301) );
 a64178a <=( (not A300)  and  a64177a );
 a64179a <=( a64178a  and  a64173a );
 a64180a <=( a64179a  and  a64170a );
 a64183a <=( (not A169)  and  A170 );
 a64186a <=( A167  and  (not A168) );
 a64187a <=( a64186a  and  a64183a );
 a64190a <=( A201  and  (not A166) );
 a64193a <=( (not A203)  and  (not A202) );
 a64194a <=( a64193a  and  a64190a );
 a64195a <=( a64194a  and  a64187a );
 a64198a <=( (not A233)  and  A232 );
 a64201a <=( A235  and  A234 );
 a64202a <=( a64201a  and  a64198a );
 a64205a <=( A266  and  (not A265) );
 a64209a <=( (not A269)  and  (not A268) );
 a64210a <=( (not A267)  and  a64209a );
 a64211a <=( a64210a  and  a64205a );
 a64212a <=( a64211a  and  a64202a );
 a64215a <=( (not A169)  and  A170 );
 a64218a <=( A167  and  (not A168) );
 a64219a <=( a64218a  and  a64215a );
 a64222a <=( A201  and  (not A166) );
 a64225a <=( (not A203)  and  (not A202) );
 a64226a <=( a64225a  and  a64222a );
 a64227a <=( a64226a  and  a64219a );
 a64230a <=( (not A233)  and  A232 );
 a64233a <=( A235  and  A234 );
 a64234a <=( a64233a  and  a64230a );
 a64237a <=( (not A266)  and  A265 );
 a64241a <=( (not A269)  and  (not A268) );
 a64242a <=( (not A267)  and  a64241a );
 a64243a <=( a64242a  and  a64237a );
 a64244a <=( a64243a  and  a64234a );
 a64247a <=( (not A169)  and  A170 );
 a64250a <=( A167  and  (not A168) );
 a64251a <=( a64250a  and  a64247a );
 a64254a <=( A201  and  (not A166) );
 a64257a <=( (not A203)  and  (not A202) );
 a64258a <=( a64257a  and  a64254a );
 a64259a <=( a64258a  and  a64251a );
 a64262a <=( (not A233)  and  A232 );
 a64265a <=( A236  and  A234 );
 a64266a <=( a64265a  and  a64262a );
 a64269a <=( (not A299)  and  A298 );
 a64273a <=( (not A302)  and  (not A301) );
 a64274a <=( (not A300)  and  a64273a );
 a64275a <=( a64274a  and  a64269a );
 a64276a <=( a64275a  and  a64266a );
 a64279a <=( (not A169)  and  A170 );
 a64282a <=( A167  and  (not A168) );
 a64283a <=( a64282a  and  a64279a );
 a64286a <=( A201  and  (not A166) );
 a64289a <=( (not A203)  and  (not A202) );
 a64290a <=( a64289a  and  a64286a );
 a64291a <=( a64290a  and  a64283a );
 a64294a <=( (not A233)  and  A232 );
 a64297a <=( A236  and  A234 );
 a64298a <=( a64297a  and  a64294a );
 a64301a <=( A299  and  (not A298) );
 a64305a <=( (not A302)  and  (not A301) );
 a64306a <=( (not A300)  and  a64305a );
 a64307a <=( a64306a  and  a64301a );
 a64308a <=( a64307a  and  a64298a );
 a64311a <=( (not A169)  and  A170 );
 a64314a <=( A167  and  (not A168) );
 a64315a <=( a64314a  and  a64311a );
 a64318a <=( A201  and  (not A166) );
 a64321a <=( (not A203)  and  (not A202) );
 a64322a <=( a64321a  and  a64318a );
 a64323a <=( a64322a  and  a64315a );
 a64326a <=( (not A233)  and  A232 );
 a64329a <=( A236  and  A234 );
 a64330a <=( a64329a  and  a64326a );
 a64333a <=( A266  and  (not A265) );
 a64337a <=( (not A269)  and  (not A268) );
 a64338a <=( (not A267)  and  a64337a );
 a64339a <=( a64338a  and  a64333a );
 a64340a <=( a64339a  and  a64330a );
 a64343a <=( (not A169)  and  A170 );
 a64346a <=( A167  and  (not A168) );
 a64347a <=( a64346a  and  a64343a );
 a64350a <=( A201  and  (not A166) );
 a64353a <=( (not A203)  and  (not A202) );
 a64354a <=( a64353a  and  a64350a );
 a64355a <=( a64354a  and  a64347a );
 a64358a <=( (not A233)  and  A232 );
 a64361a <=( A236  and  A234 );
 a64362a <=( a64361a  and  a64358a );
 a64365a <=( (not A266)  and  A265 );
 a64369a <=( (not A269)  and  (not A268) );
 a64370a <=( (not A267)  and  a64369a );
 a64371a <=( a64370a  and  a64365a );
 a64372a <=( a64371a  and  a64362a );
 a64375a <=( (not A169)  and  A170 );
 a64378a <=( A167  and  (not A168) );
 a64379a <=( a64378a  and  a64375a );
 a64382a <=( A201  and  (not A166) );
 a64385a <=( (not A203)  and  (not A202) );
 a64386a <=( a64385a  and  a64382a );
 a64387a <=( a64386a  and  a64379a );
 a64390a <=( (not A233)  and  A232 );
 a64393a <=( (not A235)  and  (not A234) );
 a64394a <=( a64393a  and  a64390a );
 a64397a <=( A298  and  (not A236) );
 a64401a <=( A301  and  A300 );
 a64402a <=( (not A299)  and  a64401a );
 a64403a <=( a64402a  and  a64397a );
 a64404a <=( a64403a  and  a64394a );
 a64407a <=( (not A169)  and  A170 );
 a64410a <=( A167  and  (not A168) );
 a64411a <=( a64410a  and  a64407a );
 a64414a <=( A201  and  (not A166) );
 a64417a <=( (not A203)  and  (not A202) );
 a64418a <=( a64417a  and  a64414a );
 a64419a <=( a64418a  and  a64411a );
 a64422a <=( (not A233)  and  A232 );
 a64425a <=( (not A235)  and  (not A234) );
 a64426a <=( a64425a  and  a64422a );
 a64429a <=( A298  and  (not A236) );
 a64433a <=( A302  and  A300 );
 a64434a <=( (not A299)  and  a64433a );
 a64435a <=( a64434a  and  a64429a );
 a64436a <=( a64435a  and  a64426a );
 a64439a <=( (not A169)  and  A170 );
 a64442a <=( A167  and  (not A168) );
 a64443a <=( a64442a  and  a64439a );
 a64446a <=( A201  and  (not A166) );
 a64449a <=( (not A203)  and  (not A202) );
 a64450a <=( a64449a  and  a64446a );
 a64451a <=( a64450a  and  a64443a );
 a64454a <=( (not A233)  and  A232 );
 a64457a <=( (not A235)  and  (not A234) );
 a64458a <=( a64457a  and  a64454a );
 a64461a <=( (not A298)  and  (not A236) );
 a64465a <=( A301  and  A300 );
 a64466a <=( A299  and  a64465a );
 a64467a <=( a64466a  and  a64461a );
 a64468a <=( a64467a  and  a64458a );
 a64471a <=( (not A169)  and  A170 );
 a64474a <=( A167  and  (not A168) );
 a64475a <=( a64474a  and  a64471a );
 a64478a <=( A201  and  (not A166) );
 a64481a <=( (not A203)  and  (not A202) );
 a64482a <=( a64481a  and  a64478a );
 a64483a <=( a64482a  and  a64475a );
 a64486a <=( (not A233)  and  A232 );
 a64489a <=( (not A235)  and  (not A234) );
 a64490a <=( a64489a  and  a64486a );
 a64493a <=( (not A298)  and  (not A236) );
 a64497a <=( A302  and  A300 );
 a64498a <=( A299  and  a64497a );
 a64499a <=( a64498a  and  a64493a );
 a64500a <=( a64499a  and  a64490a );
 a64503a <=( (not A169)  and  A170 );
 a64506a <=( A167  and  (not A168) );
 a64507a <=( a64506a  and  a64503a );
 a64510a <=( A201  and  (not A166) );
 a64513a <=( (not A203)  and  (not A202) );
 a64514a <=( a64513a  and  a64510a );
 a64515a <=( a64514a  and  a64507a );
 a64518a <=( (not A233)  and  A232 );
 a64521a <=( (not A235)  and  (not A234) );
 a64522a <=( a64521a  and  a64518a );
 a64525a <=( (not A265)  and  (not A236) );
 a64529a <=( A268  and  A267 );
 a64530a <=( A266  and  a64529a );
 a64531a <=( a64530a  and  a64525a );
 a64532a <=( a64531a  and  a64522a );
 a64535a <=( (not A169)  and  A170 );
 a64538a <=( A167  and  (not A168) );
 a64539a <=( a64538a  and  a64535a );
 a64542a <=( A201  and  (not A166) );
 a64545a <=( (not A203)  and  (not A202) );
 a64546a <=( a64545a  and  a64542a );
 a64547a <=( a64546a  and  a64539a );
 a64550a <=( (not A233)  and  A232 );
 a64553a <=( (not A235)  and  (not A234) );
 a64554a <=( a64553a  and  a64550a );
 a64557a <=( (not A265)  and  (not A236) );
 a64561a <=( A269  and  A267 );
 a64562a <=( A266  and  a64561a );
 a64563a <=( a64562a  and  a64557a );
 a64564a <=( a64563a  and  a64554a );
 a64567a <=( (not A169)  and  A170 );
 a64570a <=( A167  and  (not A168) );
 a64571a <=( a64570a  and  a64567a );
 a64574a <=( A201  and  (not A166) );
 a64577a <=( (not A203)  and  (not A202) );
 a64578a <=( a64577a  and  a64574a );
 a64579a <=( a64578a  and  a64571a );
 a64582a <=( (not A233)  and  A232 );
 a64585a <=( (not A235)  and  (not A234) );
 a64586a <=( a64585a  and  a64582a );
 a64589a <=( A265  and  (not A236) );
 a64593a <=( A268  and  A267 );
 a64594a <=( (not A266)  and  a64593a );
 a64595a <=( a64594a  and  a64589a );
 a64596a <=( a64595a  and  a64586a );
 a64599a <=( (not A169)  and  A170 );
 a64602a <=( A167  and  (not A168) );
 a64603a <=( a64602a  and  a64599a );
 a64606a <=( A201  and  (not A166) );
 a64609a <=( (not A203)  and  (not A202) );
 a64610a <=( a64609a  and  a64606a );
 a64611a <=( a64610a  and  a64603a );
 a64614a <=( (not A233)  and  A232 );
 a64617a <=( (not A235)  and  (not A234) );
 a64618a <=( a64617a  and  a64614a );
 a64621a <=( A265  and  (not A236) );
 a64625a <=( A269  and  A267 );
 a64626a <=( (not A266)  and  a64625a );
 a64627a <=( a64626a  and  a64621a );
 a64628a <=( a64627a  and  a64618a );
 a64631a <=( (not A169)  and  A170 );
 a64634a <=( A167  and  (not A168) );
 a64635a <=( a64634a  and  a64631a );
 a64638a <=( (not A201)  and  (not A166) );
 a64641a <=( (not A232)  and  A202 );
 a64642a <=( a64641a  and  a64638a );
 a64643a <=( a64642a  and  a64635a );
 a64646a <=( (not A234)  and  A233 );
 a64649a <=( (not A236)  and  (not A235) );
 a64650a <=( a64649a  and  a64646a );
 a64653a <=( (not A299)  and  A298 );
 a64657a <=( (not A302)  and  (not A301) );
 a64658a <=( (not A300)  and  a64657a );
 a64659a <=( a64658a  and  a64653a );
 a64660a <=( a64659a  and  a64650a );
 a64663a <=( (not A169)  and  A170 );
 a64666a <=( A167  and  (not A168) );
 a64667a <=( a64666a  and  a64663a );
 a64670a <=( (not A201)  and  (not A166) );
 a64673a <=( (not A232)  and  A202 );
 a64674a <=( a64673a  and  a64670a );
 a64675a <=( a64674a  and  a64667a );
 a64678a <=( (not A234)  and  A233 );
 a64681a <=( (not A236)  and  (not A235) );
 a64682a <=( a64681a  and  a64678a );
 a64685a <=( A299  and  (not A298) );
 a64689a <=( (not A302)  and  (not A301) );
 a64690a <=( (not A300)  and  a64689a );
 a64691a <=( a64690a  and  a64685a );
 a64692a <=( a64691a  and  a64682a );
 a64695a <=( (not A169)  and  A170 );
 a64698a <=( A167  and  (not A168) );
 a64699a <=( a64698a  and  a64695a );
 a64702a <=( (not A201)  and  (not A166) );
 a64705a <=( (not A232)  and  A202 );
 a64706a <=( a64705a  and  a64702a );
 a64707a <=( a64706a  and  a64699a );
 a64710a <=( (not A234)  and  A233 );
 a64713a <=( (not A236)  and  (not A235) );
 a64714a <=( a64713a  and  a64710a );
 a64717a <=( A266  and  (not A265) );
 a64721a <=( (not A269)  and  (not A268) );
 a64722a <=( (not A267)  and  a64721a );
 a64723a <=( a64722a  and  a64717a );
 a64724a <=( a64723a  and  a64714a );
 a64727a <=( (not A169)  and  A170 );
 a64730a <=( A167  and  (not A168) );
 a64731a <=( a64730a  and  a64727a );
 a64734a <=( (not A201)  and  (not A166) );
 a64737a <=( (not A232)  and  A202 );
 a64738a <=( a64737a  and  a64734a );
 a64739a <=( a64738a  and  a64731a );
 a64742a <=( (not A234)  and  A233 );
 a64745a <=( (not A236)  and  (not A235) );
 a64746a <=( a64745a  and  a64742a );
 a64749a <=( (not A266)  and  A265 );
 a64753a <=( (not A269)  and  (not A268) );
 a64754a <=( (not A267)  and  a64753a );
 a64755a <=( a64754a  and  a64749a );
 a64756a <=( a64755a  and  a64746a );
 a64759a <=( (not A169)  and  A170 );
 a64762a <=( A167  and  (not A168) );
 a64763a <=( a64762a  and  a64759a );
 a64766a <=( (not A201)  and  (not A166) );
 a64769a <=( A232  and  A202 );
 a64770a <=( a64769a  and  a64766a );
 a64771a <=( a64770a  and  a64763a );
 a64774a <=( (not A234)  and  (not A233) );
 a64777a <=( (not A236)  and  (not A235) );
 a64778a <=( a64777a  and  a64774a );
 a64781a <=( (not A299)  and  A298 );
 a64785a <=( (not A302)  and  (not A301) );
 a64786a <=( (not A300)  and  a64785a );
 a64787a <=( a64786a  and  a64781a );
 a64788a <=( a64787a  and  a64778a );
 a64791a <=( (not A169)  and  A170 );
 a64794a <=( A167  and  (not A168) );
 a64795a <=( a64794a  and  a64791a );
 a64798a <=( (not A201)  and  (not A166) );
 a64801a <=( A232  and  A202 );
 a64802a <=( a64801a  and  a64798a );
 a64803a <=( a64802a  and  a64795a );
 a64806a <=( (not A234)  and  (not A233) );
 a64809a <=( (not A236)  and  (not A235) );
 a64810a <=( a64809a  and  a64806a );
 a64813a <=( A299  and  (not A298) );
 a64817a <=( (not A302)  and  (not A301) );
 a64818a <=( (not A300)  and  a64817a );
 a64819a <=( a64818a  and  a64813a );
 a64820a <=( a64819a  and  a64810a );
 a64823a <=( (not A169)  and  A170 );
 a64826a <=( A167  and  (not A168) );
 a64827a <=( a64826a  and  a64823a );
 a64830a <=( (not A201)  and  (not A166) );
 a64833a <=( A232  and  A202 );
 a64834a <=( a64833a  and  a64830a );
 a64835a <=( a64834a  and  a64827a );
 a64838a <=( (not A234)  and  (not A233) );
 a64841a <=( (not A236)  and  (not A235) );
 a64842a <=( a64841a  and  a64838a );
 a64845a <=( A266  and  (not A265) );
 a64849a <=( (not A269)  and  (not A268) );
 a64850a <=( (not A267)  and  a64849a );
 a64851a <=( a64850a  and  a64845a );
 a64852a <=( a64851a  and  a64842a );
 a64855a <=( (not A169)  and  A170 );
 a64858a <=( A167  and  (not A168) );
 a64859a <=( a64858a  and  a64855a );
 a64862a <=( (not A201)  and  (not A166) );
 a64865a <=( A232  and  A202 );
 a64866a <=( a64865a  and  a64862a );
 a64867a <=( a64866a  and  a64859a );
 a64870a <=( (not A234)  and  (not A233) );
 a64873a <=( (not A236)  and  (not A235) );
 a64874a <=( a64873a  and  a64870a );
 a64877a <=( (not A266)  and  A265 );
 a64881a <=( (not A269)  and  (not A268) );
 a64882a <=( (not A267)  and  a64881a );
 a64883a <=( a64882a  and  a64877a );
 a64884a <=( a64883a  and  a64874a );
 a64887a <=( (not A169)  and  A170 );
 a64890a <=( A167  and  (not A168) );
 a64891a <=( a64890a  and  a64887a );
 a64894a <=( (not A201)  and  (not A166) );
 a64897a <=( (not A232)  and  A203 );
 a64898a <=( a64897a  and  a64894a );
 a64899a <=( a64898a  and  a64891a );
 a64902a <=( (not A234)  and  A233 );
 a64905a <=( (not A236)  and  (not A235) );
 a64906a <=( a64905a  and  a64902a );
 a64909a <=( (not A299)  and  A298 );
 a64913a <=( (not A302)  and  (not A301) );
 a64914a <=( (not A300)  and  a64913a );
 a64915a <=( a64914a  and  a64909a );
 a64916a <=( a64915a  and  a64906a );
 a64919a <=( (not A169)  and  A170 );
 a64922a <=( A167  and  (not A168) );
 a64923a <=( a64922a  and  a64919a );
 a64926a <=( (not A201)  and  (not A166) );
 a64929a <=( (not A232)  and  A203 );
 a64930a <=( a64929a  and  a64926a );
 a64931a <=( a64930a  and  a64923a );
 a64934a <=( (not A234)  and  A233 );
 a64937a <=( (not A236)  and  (not A235) );
 a64938a <=( a64937a  and  a64934a );
 a64941a <=( A299  and  (not A298) );
 a64945a <=( (not A302)  and  (not A301) );
 a64946a <=( (not A300)  and  a64945a );
 a64947a <=( a64946a  and  a64941a );
 a64948a <=( a64947a  and  a64938a );
 a64951a <=( (not A169)  and  A170 );
 a64954a <=( A167  and  (not A168) );
 a64955a <=( a64954a  and  a64951a );
 a64958a <=( (not A201)  and  (not A166) );
 a64961a <=( (not A232)  and  A203 );
 a64962a <=( a64961a  and  a64958a );
 a64963a <=( a64962a  and  a64955a );
 a64966a <=( (not A234)  and  A233 );
 a64969a <=( (not A236)  and  (not A235) );
 a64970a <=( a64969a  and  a64966a );
 a64973a <=( A266  and  (not A265) );
 a64977a <=( (not A269)  and  (not A268) );
 a64978a <=( (not A267)  and  a64977a );
 a64979a <=( a64978a  and  a64973a );
 a64980a <=( a64979a  and  a64970a );
 a64983a <=( (not A169)  and  A170 );
 a64986a <=( A167  and  (not A168) );
 a64987a <=( a64986a  and  a64983a );
 a64990a <=( (not A201)  and  (not A166) );
 a64993a <=( (not A232)  and  A203 );
 a64994a <=( a64993a  and  a64990a );
 a64995a <=( a64994a  and  a64987a );
 a64998a <=( (not A234)  and  A233 );
 a65001a <=( (not A236)  and  (not A235) );
 a65002a <=( a65001a  and  a64998a );
 a65005a <=( (not A266)  and  A265 );
 a65009a <=( (not A269)  and  (not A268) );
 a65010a <=( (not A267)  and  a65009a );
 a65011a <=( a65010a  and  a65005a );
 a65012a <=( a65011a  and  a65002a );
 a65015a <=( (not A169)  and  A170 );
 a65018a <=( A167  and  (not A168) );
 a65019a <=( a65018a  and  a65015a );
 a65022a <=( (not A201)  and  (not A166) );
 a65025a <=( A232  and  A203 );
 a65026a <=( a65025a  and  a65022a );
 a65027a <=( a65026a  and  a65019a );
 a65030a <=( (not A234)  and  (not A233) );
 a65033a <=( (not A236)  and  (not A235) );
 a65034a <=( a65033a  and  a65030a );
 a65037a <=( (not A299)  and  A298 );
 a65041a <=( (not A302)  and  (not A301) );
 a65042a <=( (not A300)  and  a65041a );
 a65043a <=( a65042a  and  a65037a );
 a65044a <=( a65043a  and  a65034a );
 a65047a <=( (not A169)  and  A170 );
 a65050a <=( A167  and  (not A168) );
 a65051a <=( a65050a  and  a65047a );
 a65054a <=( (not A201)  and  (not A166) );
 a65057a <=( A232  and  A203 );
 a65058a <=( a65057a  and  a65054a );
 a65059a <=( a65058a  and  a65051a );
 a65062a <=( (not A234)  and  (not A233) );
 a65065a <=( (not A236)  and  (not A235) );
 a65066a <=( a65065a  and  a65062a );
 a65069a <=( A299  and  (not A298) );
 a65073a <=( (not A302)  and  (not A301) );
 a65074a <=( (not A300)  and  a65073a );
 a65075a <=( a65074a  and  a65069a );
 a65076a <=( a65075a  and  a65066a );
 a65079a <=( (not A169)  and  A170 );
 a65082a <=( A167  and  (not A168) );
 a65083a <=( a65082a  and  a65079a );
 a65086a <=( (not A201)  and  (not A166) );
 a65089a <=( A232  and  A203 );
 a65090a <=( a65089a  and  a65086a );
 a65091a <=( a65090a  and  a65083a );
 a65094a <=( (not A234)  and  (not A233) );
 a65097a <=( (not A236)  and  (not A235) );
 a65098a <=( a65097a  and  a65094a );
 a65101a <=( A266  and  (not A265) );
 a65105a <=( (not A269)  and  (not A268) );
 a65106a <=( (not A267)  and  a65105a );
 a65107a <=( a65106a  and  a65101a );
 a65108a <=( a65107a  and  a65098a );
 a65111a <=( (not A169)  and  A170 );
 a65114a <=( A167  and  (not A168) );
 a65115a <=( a65114a  and  a65111a );
 a65118a <=( (not A201)  and  (not A166) );
 a65121a <=( A232  and  A203 );
 a65122a <=( a65121a  and  a65118a );
 a65123a <=( a65122a  and  a65115a );
 a65126a <=( (not A234)  and  (not A233) );
 a65129a <=( (not A236)  and  (not A235) );
 a65130a <=( a65129a  and  a65126a );
 a65133a <=( (not A266)  and  A265 );
 a65137a <=( (not A269)  and  (not A268) );
 a65138a <=( (not A267)  and  a65137a );
 a65139a <=( a65138a  and  a65133a );
 a65140a <=( a65139a  and  a65130a );
 a65143a <=( (not A169)  and  A170 );
 a65146a <=( A167  and  (not A168) );
 a65147a <=( a65146a  and  a65143a );
 a65150a <=( A199  and  (not A166) );
 a65153a <=( (not A232)  and  A200 );
 a65154a <=( a65153a  and  a65150a );
 a65155a <=( a65154a  and  a65147a );
 a65158a <=( (not A234)  and  A233 );
 a65161a <=( (not A236)  and  (not A235) );
 a65162a <=( a65161a  and  a65158a );
 a65165a <=( (not A299)  and  A298 );
 a65169a <=( (not A302)  and  (not A301) );
 a65170a <=( (not A300)  and  a65169a );
 a65171a <=( a65170a  and  a65165a );
 a65172a <=( a65171a  and  a65162a );
 a65175a <=( (not A169)  and  A170 );
 a65178a <=( A167  and  (not A168) );
 a65179a <=( a65178a  and  a65175a );
 a65182a <=( A199  and  (not A166) );
 a65185a <=( (not A232)  and  A200 );
 a65186a <=( a65185a  and  a65182a );
 a65187a <=( a65186a  and  a65179a );
 a65190a <=( (not A234)  and  A233 );
 a65193a <=( (not A236)  and  (not A235) );
 a65194a <=( a65193a  and  a65190a );
 a65197a <=( A299  and  (not A298) );
 a65201a <=( (not A302)  and  (not A301) );
 a65202a <=( (not A300)  and  a65201a );
 a65203a <=( a65202a  and  a65197a );
 a65204a <=( a65203a  and  a65194a );
 a65207a <=( (not A169)  and  A170 );
 a65210a <=( A167  and  (not A168) );
 a65211a <=( a65210a  and  a65207a );
 a65214a <=( A199  and  (not A166) );
 a65217a <=( (not A232)  and  A200 );
 a65218a <=( a65217a  and  a65214a );
 a65219a <=( a65218a  and  a65211a );
 a65222a <=( (not A234)  and  A233 );
 a65225a <=( (not A236)  and  (not A235) );
 a65226a <=( a65225a  and  a65222a );
 a65229a <=( A266  and  (not A265) );
 a65233a <=( (not A269)  and  (not A268) );
 a65234a <=( (not A267)  and  a65233a );
 a65235a <=( a65234a  and  a65229a );
 a65236a <=( a65235a  and  a65226a );
 a65239a <=( (not A169)  and  A170 );
 a65242a <=( A167  and  (not A168) );
 a65243a <=( a65242a  and  a65239a );
 a65246a <=( A199  and  (not A166) );
 a65249a <=( (not A232)  and  A200 );
 a65250a <=( a65249a  and  a65246a );
 a65251a <=( a65250a  and  a65243a );
 a65254a <=( (not A234)  and  A233 );
 a65257a <=( (not A236)  and  (not A235) );
 a65258a <=( a65257a  and  a65254a );
 a65261a <=( (not A266)  and  A265 );
 a65265a <=( (not A269)  and  (not A268) );
 a65266a <=( (not A267)  and  a65265a );
 a65267a <=( a65266a  and  a65261a );
 a65268a <=( a65267a  and  a65258a );
 a65271a <=( (not A169)  and  A170 );
 a65274a <=( A167  and  (not A168) );
 a65275a <=( a65274a  and  a65271a );
 a65278a <=( A199  and  (not A166) );
 a65281a <=( A232  and  A200 );
 a65282a <=( a65281a  and  a65278a );
 a65283a <=( a65282a  and  a65275a );
 a65286a <=( (not A234)  and  (not A233) );
 a65289a <=( (not A236)  and  (not A235) );
 a65290a <=( a65289a  and  a65286a );
 a65293a <=( (not A299)  and  A298 );
 a65297a <=( (not A302)  and  (not A301) );
 a65298a <=( (not A300)  and  a65297a );
 a65299a <=( a65298a  and  a65293a );
 a65300a <=( a65299a  and  a65290a );
 a65303a <=( (not A169)  and  A170 );
 a65306a <=( A167  and  (not A168) );
 a65307a <=( a65306a  and  a65303a );
 a65310a <=( A199  and  (not A166) );
 a65313a <=( A232  and  A200 );
 a65314a <=( a65313a  and  a65310a );
 a65315a <=( a65314a  and  a65307a );
 a65318a <=( (not A234)  and  (not A233) );
 a65321a <=( (not A236)  and  (not A235) );
 a65322a <=( a65321a  and  a65318a );
 a65325a <=( A299  and  (not A298) );
 a65329a <=( (not A302)  and  (not A301) );
 a65330a <=( (not A300)  and  a65329a );
 a65331a <=( a65330a  and  a65325a );
 a65332a <=( a65331a  and  a65322a );
 a65335a <=( (not A169)  and  A170 );
 a65338a <=( A167  and  (not A168) );
 a65339a <=( a65338a  and  a65335a );
 a65342a <=( A199  and  (not A166) );
 a65345a <=( A232  and  A200 );
 a65346a <=( a65345a  and  a65342a );
 a65347a <=( a65346a  and  a65339a );
 a65350a <=( (not A234)  and  (not A233) );
 a65353a <=( (not A236)  and  (not A235) );
 a65354a <=( a65353a  and  a65350a );
 a65357a <=( A266  and  (not A265) );
 a65361a <=( (not A269)  and  (not A268) );
 a65362a <=( (not A267)  and  a65361a );
 a65363a <=( a65362a  and  a65357a );
 a65364a <=( a65363a  and  a65354a );
 a65367a <=( (not A169)  and  A170 );
 a65370a <=( A167  and  (not A168) );
 a65371a <=( a65370a  and  a65367a );
 a65374a <=( A199  and  (not A166) );
 a65377a <=( A232  and  A200 );
 a65378a <=( a65377a  and  a65374a );
 a65379a <=( a65378a  and  a65371a );
 a65382a <=( (not A234)  and  (not A233) );
 a65385a <=( (not A236)  and  (not A235) );
 a65386a <=( a65385a  and  a65382a );
 a65389a <=( (not A266)  and  A265 );
 a65393a <=( (not A269)  and  (not A268) );
 a65394a <=( (not A267)  and  a65393a );
 a65395a <=( a65394a  and  a65389a );
 a65396a <=( a65395a  and  a65386a );
 a65399a <=( (not A169)  and  A170 );
 a65402a <=( A167  and  (not A168) );
 a65403a <=( a65402a  and  a65399a );
 a65406a <=( (not A199)  and  (not A166) );
 a65409a <=( (not A232)  and  (not A200) );
 a65410a <=( a65409a  and  a65406a );
 a65411a <=( a65410a  and  a65403a );
 a65414a <=( (not A234)  and  A233 );
 a65417a <=( (not A236)  and  (not A235) );
 a65418a <=( a65417a  and  a65414a );
 a65421a <=( (not A299)  and  A298 );
 a65425a <=( (not A302)  and  (not A301) );
 a65426a <=( (not A300)  and  a65425a );
 a65427a <=( a65426a  and  a65421a );
 a65428a <=( a65427a  and  a65418a );
 a65431a <=( (not A169)  and  A170 );
 a65434a <=( A167  and  (not A168) );
 a65435a <=( a65434a  and  a65431a );
 a65438a <=( (not A199)  and  (not A166) );
 a65441a <=( (not A232)  and  (not A200) );
 a65442a <=( a65441a  and  a65438a );
 a65443a <=( a65442a  and  a65435a );
 a65446a <=( (not A234)  and  A233 );
 a65449a <=( (not A236)  and  (not A235) );
 a65450a <=( a65449a  and  a65446a );
 a65453a <=( A299  and  (not A298) );
 a65457a <=( (not A302)  and  (not A301) );
 a65458a <=( (not A300)  and  a65457a );
 a65459a <=( a65458a  and  a65453a );
 a65460a <=( a65459a  and  a65450a );
 a65463a <=( (not A169)  and  A170 );
 a65466a <=( A167  and  (not A168) );
 a65467a <=( a65466a  and  a65463a );
 a65470a <=( (not A199)  and  (not A166) );
 a65473a <=( (not A232)  and  (not A200) );
 a65474a <=( a65473a  and  a65470a );
 a65475a <=( a65474a  and  a65467a );
 a65478a <=( (not A234)  and  A233 );
 a65481a <=( (not A236)  and  (not A235) );
 a65482a <=( a65481a  and  a65478a );
 a65485a <=( A266  and  (not A265) );
 a65489a <=( (not A269)  and  (not A268) );
 a65490a <=( (not A267)  and  a65489a );
 a65491a <=( a65490a  and  a65485a );
 a65492a <=( a65491a  and  a65482a );
 a65495a <=( (not A169)  and  A170 );
 a65498a <=( A167  and  (not A168) );
 a65499a <=( a65498a  and  a65495a );
 a65502a <=( (not A199)  and  (not A166) );
 a65505a <=( (not A232)  and  (not A200) );
 a65506a <=( a65505a  and  a65502a );
 a65507a <=( a65506a  and  a65499a );
 a65510a <=( (not A234)  and  A233 );
 a65513a <=( (not A236)  and  (not A235) );
 a65514a <=( a65513a  and  a65510a );
 a65517a <=( (not A266)  and  A265 );
 a65521a <=( (not A269)  and  (not A268) );
 a65522a <=( (not A267)  and  a65521a );
 a65523a <=( a65522a  and  a65517a );
 a65524a <=( a65523a  and  a65514a );
 a65527a <=( (not A169)  and  A170 );
 a65530a <=( A167  and  (not A168) );
 a65531a <=( a65530a  and  a65527a );
 a65534a <=( (not A199)  and  (not A166) );
 a65537a <=( A232  and  (not A200) );
 a65538a <=( a65537a  and  a65534a );
 a65539a <=( a65538a  and  a65531a );
 a65542a <=( (not A234)  and  (not A233) );
 a65545a <=( (not A236)  and  (not A235) );
 a65546a <=( a65545a  and  a65542a );
 a65549a <=( (not A299)  and  A298 );
 a65553a <=( (not A302)  and  (not A301) );
 a65554a <=( (not A300)  and  a65553a );
 a65555a <=( a65554a  and  a65549a );
 a65556a <=( a65555a  and  a65546a );
 a65559a <=( (not A169)  and  A170 );
 a65562a <=( A167  and  (not A168) );
 a65563a <=( a65562a  and  a65559a );
 a65566a <=( (not A199)  and  (not A166) );
 a65569a <=( A232  and  (not A200) );
 a65570a <=( a65569a  and  a65566a );
 a65571a <=( a65570a  and  a65563a );
 a65574a <=( (not A234)  and  (not A233) );
 a65577a <=( (not A236)  and  (not A235) );
 a65578a <=( a65577a  and  a65574a );
 a65581a <=( A299  and  (not A298) );
 a65585a <=( (not A302)  and  (not A301) );
 a65586a <=( (not A300)  and  a65585a );
 a65587a <=( a65586a  and  a65581a );
 a65588a <=( a65587a  and  a65578a );
 a65591a <=( (not A169)  and  A170 );
 a65594a <=( A167  and  (not A168) );
 a65595a <=( a65594a  and  a65591a );
 a65598a <=( (not A199)  and  (not A166) );
 a65601a <=( A232  and  (not A200) );
 a65602a <=( a65601a  and  a65598a );
 a65603a <=( a65602a  and  a65595a );
 a65606a <=( (not A234)  and  (not A233) );
 a65609a <=( (not A236)  and  (not A235) );
 a65610a <=( a65609a  and  a65606a );
 a65613a <=( A266  and  (not A265) );
 a65617a <=( (not A269)  and  (not A268) );
 a65618a <=( (not A267)  and  a65617a );
 a65619a <=( a65618a  and  a65613a );
 a65620a <=( a65619a  and  a65610a );
 a65623a <=( (not A169)  and  A170 );
 a65626a <=( A167  and  (not A168) );
 a65627a <=( a65626a  and  a65623a );
 a65630a <=( (not A199)  and  (not A166) );
 a65633a <=( A232  and  (not A200) );
 a65634a <=( a65633a  and  a65630a );
 a65635a <=( a65634a  and  a65627a );
 a65638a <=( (not A234)  and  (not A233) );
 a65641a <=( (not A236)  and  (not A235) );
 a65642a <=( a65641a  and  a65638a );
 a65645a <=( (not A266)  and  A265 );
 a65649a <=( (not A269)  and  (not A268) );
 a65650a <=( (not A267)  and  a65649a );
 a65651a <=( a65650a  and  a65645a );
 a65652a <=( a65651a  and  a65642a );
 a65655a <=( (not A169)  and  A170 );
 a65658a <=( (not A167)  and  (not A168) );
 a65659a <=( a65658a  and  a65655a );
 a65662a <=( A201  and  A166 );
 a65665a <=( (not A203)  and  (not A202) );
 a65666a <=( a65665a  and  a65662a );
 a65667a <=( a65666a  and  a65659a );
 a65670a <=( A233  and  (not A232) );
 a65673a <=( A235  and  A234 );
 a65674a <=( a65673a  and  a65670a );
 a65677a <=( (not A299)  and  A298 );
 a65681a <=( (not A302)  and  (not A301) );
 a65682a <=( (not A300)  and  a65681a );
 a65683a <=( a65682a  and  a65677a );
 a65684a <=( a65683a  and  a65674a );
 a65687a <=( (not A169)  and  A170 );
 a65690a <=( (not A167)  and  (not A168) );
 a65691a <=( a65690a  and  a65687a );
 a65694a <=( A201  and  A166 );
 a65697a <=( (not A203)  and  (not A202) );
 a65698a <=( a65697a  and  a65694a );
 a65699a <=( a65698a  and  a65691a );
 a65702a <=( A233  and  (not A232) );
 a65705a <=( A235  and  A234 );
 a65706a <=( a65705a  and  a65702a );
 a65709a <=( A299  and  (not A298) );
 a65713a <=( (not A302)  and  (not A301) );
 a65714a <=( (not A300)  and  a65713a );
 a65715a <=( a65714a  and  a65709a );
 a65716a <=( a65715a  and  a65706a );
 a65719a <=( (not A169)  and  A170 );
 a65722a <=( (not A167)  and  (not A168) );
 a65723a <=( a65722a  and  a65719a );
 a65726a <=( A201  and  A166 );
 a65729a <=( (not A203)  and  (not A202) );
 a65730a <=( a65729a  and  a65726a );
 a65731a <=( a65730a  and  a65723a );
 a65734a <=( A233  and  (not A232) );
 a65737a <=( A235  and  A234 );
 a65738a <=( a65737a  and  a65734a );
 a65741a <=( A266  and  (not A265) );
 a65745a <=( (not A269)  and  (not A268) );
 a65746a <=( (not A267)  and  a65745a );
 a65747a <=( a65746a  and  a65741a );
 a65748a <=( a65747a  and  a65738a );
 a65751a <=( (not A169)  and  A170 );
 a65754a <=( (not A167)  and  (not A168) );
 a65755a <=( a65754a  and  a65751a );
 a65758a <=( A201  and  A166 );
 a65761a <=( (not A203)  and  (not A202) );
 a65762a <=( a65761a  and  a65758a );
 a65763a <=( a65762a  and  a65755a );
 a65766a <=( A233  and  (not A232) );
 a65769a <=( A235  and  A234 );
 a65770a <=( a65769a  and  a65766a );
 a65773a <=( (not A266)  and  A265 );
 a65777a <=( (not A269)  and  (not A268) );
 a65778a <=( (not A267)  and  a65777a );
 a65779a <=( a65778a  and  a65773a );
 a65780a <=( a65779a  and  a65770a );
 a65783a <=( (not A169)  and  A170 );
 a65786a <=( (not A167)  and  (not A168) );
 a65787a <=( a65786a  and  a65783a );
 a65790a <=( A201  and  A166 );
 a65793a <=( (not A203)  and  (not A202) );
 a65794a <=( a65793a  and  a65790a );
 a65795a <=( a65794a  and  a65787a );
 a65798a <=( A233  and  (not A232) );
 a65801a <=( A236  and  A234 );
 a65802a <=( a65801a  and  a65798a );
 a65805a <=( (not A299)  and  A298 );
 a65809a <=( (not A302)  and  (not A301) );
 a65810a <=( (not A300)  and  a65809a );
 a65811a <=( a65810a  and  a65805a );
 a65812a <=( a65811a  and  a65802a );
 a65815a <=( (not A169)  and  A170 );
 a65818a <=( (not A167)  and  (not A168) );
 a65819a <=( a65818a  and  a65815a );
 a65822a <=( A201  and  A166 );
 a65825a <=( (not A203)  and  (not A202) );
 a65826a <=( a65825a  and  a65822a );
 a65827a <=( a65826a  and  a65819a );
 a65830a <=( A233  and  (not A232) );
 a65833a <=( A236  and  A234 );
 a65834a <=( a65833a  and  a65830a );
 a65837a <=( A299  and  (not A298) );
 a65841a <=( (not A302)  and  (not A301) );
 a65842a <=( (not A300)  and  a65841a );
 a65843a <=( a65842a  and  a65837a );
 a65844a <=( a65843a  and  a65834a );
 a65847a <=( (not A169)  and  A170 );
 a65850a <=( (not A167)  and  (not A168) );
 a65851a <=( a65850a  and  a65847a );
 a65854a <=( A201  and  A166 );
 a65857a <=( (not A203)  and  (not A202) );
 a65858a <=( a65857a  and  a65854a );
 a65859a <=( a65858a  and  a65851a );
 a65862a <=( A233  and  (not A232) );
 a65865a <=( A236  and  A234 );
 a65866a <=( a65865a  and  a65862a );
 a65869a <=( A266  and  (not A265) );
 a65873a <=( (not A269)  and  (not A268) );
 a65874a <=( (not A267)  and  a65873a );
 a65875a <=( a65874a  and  a65869a );
 a65876a <=( a65875a  and  a65866a );
 a65879a <=( (not A169)  and  A170 );
 a65882a <=( (not A167)  and  (not A168) );
 a65883a <=( a65882a  and  a65879a );
 a65886a <=( A201  and  A166 );
 a65889a <=( (not A203)  and  (not A202) );
 a65890a <=( a65889a  and  a65886a );
 a65891a <=( a65890a  and  a65883a );
 a65894a <=( A233  and  (not A232) );
 a65897a <=( A236  and  A234 );
 a65898a <=( a65897a  and  a65894a );
 a65901a <=( (not A266)  and  A265 );
 a65905a <=( (not A269)  and  (not A268) );
 a65906a <=( (not A267)  and  a65905a );
 a65907a <=( a65906a  and  a65901a );
 a65908a <=( a65907a  and  a65898a );
 a65911a <=( (not A169)  and  A170 );
 a65914a <=( (not A167)  and  (not A168) );
 a65915a <=( a65914a  and  a65911a );
 a65918a <=( A201  and  A166 );
 a65921a <=( (not A203)  and  (not A202) );
 a65922a <=( a65921a  and  a65918a );
 a65923a <=( a65922a  and  a65915a );
 a65926a <=( A233  and  (not A232) );
 a65929a <=( (not A235)  and  (not A234) );
 a65930a <=( a65929a  and  a65926a );
 a65933a <=( A298  and  (not A236) );
 a65937a <=( A301  and  A300 );
 a65938a <=( (not A299)  and  a65937a );
 a65939a <=( a65938a  and  a65933a );
 a65940a <=( a65939a  and  a65930a );
 a65943a <=( (not A169)  and  A170 );
 a65946a <=( (not A167)  and  (not A168) );
 a65947a <=( a65946a  and  a65943a );
 a65950a <=( A201  and  A166 );
 a65953a <=( (not A203)  and  (not A202) );
 a65954a <=( a65953a  and  a65950a );
 a65955a <=( a65954a  and  a65947a );
 a65958a <=( A233  and  (not A232) );
 a65961a <=( (not A235)  and  (not A234) );
 a65962a <=( a65961a  and  a65958a );
 a65965a <=( A298  and  (not A236) );
 a65969a <=( A302  and  A300 );
 a65970a <=( (not A299)  and  a65969a );
 a65971a <=( a65970a  and  a65965a );
 a65972a <=( a65971a  and  a65962a );
 a65975a <=( (not A169)  and  A170 );
 a65978a <=( (not A167)  and  (not A168) );
 a65979a <=( a65978a  and  a65975a );
 a65982a <=( A201  and  A166 );
 a65985a <=( (not A203)  and  (not A202) );
 a65986a <=( a65985a  and  a65982a );
 a65987a <=( a65986a  and  a65979a );
 a65990a <=( A233  and  (not A232) );
 a65993a <=( (not A235)  and  (not A234) );
 a65994a <=( a65993a  and  a65990a );
 a65997a <=( (not A298)  and  (not A236) );
 a66001a <=( A301  and  A300 );
 a66002a <=( A299  and  a66001a );
 a66003a <=( a66002a  and  a65997a );
 a66004a <=( a66003a  and  a65994a );
 a66007a <=( (not A169)  and  A170 );
 a66010a <=( (not A167)  and  (not A168) );
 a66011a <=( a66010a  and  a66007a );
 a66014a <=( A201  and  A166 );
 a66017a <=( (not A203)  and  (not A202) );
 a66018a <=( a66017a  and  a66014a );
 a66019a <=( a66018a  and  a66011a );
 a66022a <=( A233  and  (not A232) );
 a66025a <=( (not A235)  and  (not A234) );
 a66026a <=( a66025a  and  a66022a );
 a66029a <=( (not A298)  and  (not A236) );
 a66033a <=( A302  and  A300 );
 a66034a <=( A299  and  a66033a );
 a66035a <=( a66034a  and  a66029a );
 a66036a <=( a66035a  and  a66026a );
 a66039a <=( (not A169)  and  A170 );
 a66042a <=( (not A167)  and  (not A168) );
 a66043a <=( a66042a  and  a66039a );
 a66046a <=( A201  and  A166 );
 a66049a <=( (not A203)  and  (not A202) );
 a66050a <=( a66049a  and  a66046a );
 a66051a <=( a66050a  and  a66043a );
 a66054a <=( A233  and  (not A232) );
 a66057a <=( (not A235)  and  (not A234) );
 a66058a <=( a66057a  and  a66054a );
 a66061a <=( (not A265)  and  (not A236) );
 a66065a <=( A268  and  A267 );
 a66066a <=( A266  and  a66065a );
 a66067a <=( a66066a  and  a66061a );
 a66068a <=( a66067a  and  a66058a );
 a66071a <=( (not A169)  and  A170 );
 a66074a <=( (not A167)  and  (not A168) );
 a66075a <=( a66074a  and  a66071a );
 a66078a <=( A201  and  A166 );
 a66081a <=( (not A203)  and  (not A202) );
 a66082a <=( a66081a  and  a66078a );
 a66083a <=( a66082a  and  a66075a );
 a66086a <=( A233  and  (not A232) );
 a66089a <=( (not A235)  and  (not A234) );
 a66090a <=( a66089a  and  a66086a );
 a66093a <=( (not A265)  and  (not A236) );
 a66097a <=( A269  and  A267 );
 a66098a <=( A266  and  a66097a );
 a66099a <=( a66098a  and  a66093a );
 a66100a <=( a66099a  and  a66090a );
 a66103a <=( (not A169)  and  A170 );
 a66106a <=( (not A167)  and  (not A168) );
 a66107a <=( a66106a  and  a66103a );
 a66110a <=( A201  and  A166 );
 a66113a <=( (not A203)  and  (not A202) );
 a66114a <=( a66113a  and  a66110a );
 a66115a <=( a66114a  and  a66107a );
 a66118a <=( A233  and  (not A232) );
 a66121a <=( (not A235)  and  (not A234) );
 a66122a <=( a66121a  and  a66118a );
 a66125a <=( A265  and  (not A236) );
 a66129a <=( A268  and  A267 );
 a66130a <=( (not A266)  and  a66129a );
 a66131a <=( a66130a  and  a66125a );
 a66132a <=( a66131a  and  a66122a );
 a66135a <=( (not A169)  and  A170 );
 a66138a <=( (not A167)  and  (not A168) );
 a66139a <=( a66138a  and  a66135a );
 a66142a <=( A201  and  A166 );
 a66145a <=( (not A203)  and  (not A202) );
 a66146a <=( a66145a  and  a66142a );
 a66147a <=( a66146a  and  a66139a );
 a66150a <=( A233  and  (not A232) );
 a66153a <=( (not A235)  and  (not A234) );
 a66154a <=( a66153a  and  a66150a );
 a66157a <=( A265  and  (not A236) );
 a66161a <=( A269  and  A267 );
 a66162a <=( (not A266)  and  a66161a );
 a66163a <=( a66162a  and  a66157a );
 a66164a <=( a66163a  and  a66154a );
 a66167a <=( (not A169)  and  A170 );
 a66170a <=( (not A167)  and  (not A168) );
 a66171a <=( a66170a  and  a66167a );
 a66174a <=( A201  and  A166 );
 a66177a <=( (not A203)  and  (not A202) );
 a66178a <=( a66177a  and  a66174a );
 a66179a <=( a66178a  and  a66171a );
 a66182a <=( (not A233)  and  A232 );
 a66185a <=( A235  and  A234 );
 a66186a <=( a66185a  and  a66182a );
 a66189a <=( (not A299)  and  A298 );
 a66193a <=( (not A302)  and  (not A301) );
 a66194a <=( (not A300)  and  a66193a );
 a66195a <=( a66194a  and  a66189a );
 a66196a <=( a66195a  and  a66186a );
 a66199a <=( (not A169)  and  A170 );
 a66202a <=( (not A167)  and  (not A168) );
 a66203a <=( a66202a  and  a66199a );
 a66206a <=( A201  and  A166 );
 a66209a <=( (not A203)  and  (not A202) );
 a66210a <=( a66209a  and  a66206a );
 a66211a <=( a66210a  and  a66203a );
 a66214a <=( (not A233)  and  A232 );
 a66217a <=( A235  and  A234 );
 a66218a <=( a66217a  and  a66214a );
 a66221a <=( A299  and  (not A298) );
 a66225a <=( (not A302)  and  (not A301) );
 a66226a <=( (not A300)  and  a66225a );
 a66227a <=( a66226a  and  a66221a );
 a66228a <=( a66227a  and  a66218a );
 a66231a <=( (not A169)  and  A170 );
 a66234a <=( (not A167)  and  (not A168) );
 a66235a <=( a66234a  and  a66231a );
 a66238a <=( A201  and  A166 );
 a66241a <=( (not A203)  and  (not A202) );
 a66242a <=( a66241a  and  a66238a );
 a66243a <=( a66242a  and  a66235a );
 a66246a <=( (not A233)  and  A232 );
 a66249a <=( A235  and  A234 );
 a66250a <=( a66249a  and  a66246a );
 a66253a <=( A266  and  (not A265) );
 a66257a <=( (not A269)  and  (not A268) );
 a66258a <=( (not A267)  and  a66257a );
 a66259a <=( a66258a  and  a66253a );
 a66260a <=( a66259a  and  a66250a );
 a66263a <=( (not A169)  and  A170 );
 a66266a <=( (not A167)  and  (not A168) );
 a66267a <=( a66266a  and  a66263a );
 a66270a <=( A201  and  A166 );
 a66273a <=( (not A203)  and  (not A202) );
 a66274a <=( a66273a  and  a66270a );
 a66275a <=( a66274a  and  a66267a );
 a66278a <=( (not A233)  and  A232 );
 a66281a <=( A235  and  A234 );
 a66282a <=( a66281a  and  a66278a );
 a66285a <=( (not A266)  and  A265 );
 a66289a <=( (not A269)  and  (not A268) );
 a66290a <=( (not A267)  and  a66289a );
 a66291a <=( a66290a  and  a66285a );
 a66292a <=( a66291a  and  a66282a );
 a66295a <=( (not A169)  and  A170 );
 a66298a <=( (not A167)  and  (not A168) );
 a66299a <=( a66298a  and  a66295a );
 a66302a <=( A201  and  A166 );
 a66305a <=( (not A203)  and  (not A202) );
 a66306a <=( a66305a  and  a66302a );
 a66307a <=( a66306a  and  a66299a );
 a66310a <=( (not A233)  and  A232 );
 a66313a <=( A236  and  A234 );
 a66314a <=( a66313a  and  a66310a );
 a66317a <=( (not A299)  and  A298 );
 a66321a <=( (not A302)  and  (not A301) );
 a66322a <=( (not A300)  and  a66321a );
 a66323a <=( a66322a  and  a66317a );
 a66324a <=( a66323a  and  a66314a );
 a66327a <=( (not A169)  and  A170 );
 a66330a <=( (not A167)  and  (not A168) );
 a66331a <=( a66330a  and  a66327a );
 a66334a <=( A201  and  A166 );
 a66337a <=( (not A203)  and  (not A202) );
 a66338a <=( a66337a  and  a66334a );
 a66339a <=( a66338a  and  a66331a );
 a66342a <=( (not A233)  and  A232 );
 a66345a <=( A236  and  A234 );
 a66346a <=( a66345a  and  a66342a );
 a66349a <=( A299  and  (not A298) );
 a66353a <=( (not A302)  and  (not A301) );
 a66354a <=( (not A300)  and  a66353a );
 a66355a <=( a66354a  and  a66349a );
 a66356a <=( a66355a  and  a66346a );
 a66359a <=( (not A169)  and  A170 );
 a66362a <=( (not A167)  and  (not A168) );
 a66363a <=( a66362a  and  a66359a );
 a66366a <=( A201  and  A166 );
 a66369a <=( (not A203)  and  (not A202) );
 a66370a <=( a66369a  and  a66366a );
 a66371a <=( a66370a  and  a66363a );
 a66374a <=( (not A233)  and  A232 );
 a66377a <=( A236  and  A234 );
 a66378a <=( a66377a  and  a66374a );
 a66381a <=( A266  and  (not A265) );
 a66385a <=( (not A269)  and  (not A268) );
 a66386a <=( (not A267)  and  a66385a );
 a66387a <=( a66386a  and  a66381a );
 a66388a <=( a66387a  and  a66378a );
 a66391a <=( (not A169)  and  A170 );
 a66394a <=( (not A167)  and  (not A168) );
 a66395a <=( a66394a  and  a66391a );
 a66398a <=( A201  and  A166 );
 a66401a <=( (not A203)  and  (not A202) );
 a66402a <=( a66401a  and  a66398a );
 a66403a <=( a66402a  and  a66395a );
 a66406a <=( (not A233)  and  A232 );
 a66409a <=( A236  and  A234 );
 a66410a <=( a66409a  and  a66406a );
 a66413a <=( (not A266)  and  A265 );
 a66417a <=( (not A269)  and  (not A268) );
 a66418a <=( (not A267)  and  a66417a );
 a66419a <=( a66418a  and  a66413a );
 a66420a <=( a66419a  and  a66410a );
 a66423a <=( (not A169)  and  A170 );
 a66426a <=( (not A167)  and  (not A168) );
 a66427a <=( a66426a  and  a66423a );
 a66430a <=( A201  and  A166 );
 a66433a <=( (not A203)  and  (not A202) );
 a66434a <=( a66433a  and  a66430a );
 a66435a <=( a66434a  and  a66427a );
 a66438a <=( (not A233)  and  A232 );
 a66441a <=( (not A235)  and  (not A234) );
 a66442a <=( a66441a  and  a66438a );
 a66445a <=( A298  and  (not A236) );
 a66449a <=( A301  and  A300 );
 a66450a <=( (not A299)  and  a66449a );
 a66451a <=( a66450a  and  a66445a );
 a66452a <=( a66451a  and  a66442a );
 a66455a <=( (not A169)  and  A170 );
 a66458a <=( (not A167)  and  (not A168) );
 a66459a <=( a66458a  and  a66455a );
 a66462a <=( A201  and  A166 );
 a66465a <=( (not A203)  and  (not A202) );
 a66466a <=( a66465a  and  a66462a );
 a66467a <=( a66466a  and  a66459a );
 a66470a <=( (not A233)  and  A232 );
 a66473a <=( (not A235)  and  (not A234) );
 a66474a <=( a66473a  and  a66470a );
 a66477a <=( A298  and  (not A236) );
 a66481a <=( A302  and  A300 );
 a66482a <=( (not A299)  and  a66481a );
 a66483a <=( a66482a  and  a66477a );
 a66484a <=( a66483a  and  a66474a );
 a66487a <=( (not A169)  and  A170 );
 a66490a <=( (not A167)  and  (not A168) );
 a66491a <=( a66490a  and  a66487a );
 a66494a <=( A201  and  A166 );
 a66497a <=( (not A203)  and  (not A202) );
 a66498a <=( a66497a  and  a66494a );
 a66499a <=( a66498a  and  a66491a );
 a66502a <=( (not A233)  and  A232 );
 a66505a <=( (not A235)  and  (not A234) );
 a66506a <=( a66505a  and  a66502a );
 a66509a <=( (not A298)  and  (not A236) );
 a66513a <=( A301  and  A300 );
 a66514a <=( A299  and  a66513a );
 a66515a <=( a66514a  and  a66509a );
 a66516a <=( a66515a  and  a66506a );
 a66519a <=( (not A169)  and  A170 );
 a66522a <=( (not A167)  and  (not A168) );
 a66523a <=( a66522a  and  a66519a );
 a66526a <=( A201  and  A166 );
 a66529a <=( (not A203)  and  (not A202) );
 a66530a <=( a66529a  and  a66526a );
 a66531a <=( a66530a  and  a66523a );
 a66534a <=( (not A233)  and  A232 );
 a66537a <=( (not A235)  and  (not A234) );
 a66538a <=( a66537a  and  a66534a );
 a66541a <=( (not A298)  and  (not A236) );
 a66545a <=( A302  and  A300 );
 a66546a <=( A299  and  a66545a );
 a66547a <=( a66546a  and  a66541a );
 a66548a <=( a66547a  and  a66538a );
 a66551a <=( (not A169)  and  A170 );
 a66554a <=( (not A167)  and  (not A168) );
 a66555a <=( a66554a  and  a66551a );
 a66558a <=( A201  and  A166 );
 a66561a <=( (not A203)  and  (not A202) );
 a66562a <=( a66561a  and  a66558a );
 a66563a <=( a66562a  and  a66555a );
 a66566a <=( (not A233)  and  A232 );
 a66569a <=( (not A235)  and  (not A234) );
 a66570a <=( a66569a  and  a66566a );
 a66573a <=( (not A265)  and  (not A236) );
 a66577a <=( A268  and  A267 );
 a66578a <=( A266  and  a66577a );
 a66579a <=( a66578a  and  a66573a );
 a66580a <=( a66579a  and  a66570a );
 a66583a <=( (not A169)  and  A170 );
 a66586a <=( (not A167)  and  (not A168) );
 a66587a <=( a66586a  and  a66583a );
 a66590a <=( A201  and  A166 );
 a66593a <=( (not A203)  and  (not A202) );
 a66594a <=( a66593a  and  a66590a );
 a66595a <=( a66594a  and  a66587a );
 a66598a <=( (not A233)  and  A232 );
 a66601a <=( (not A235)  and  (not A234) );
 a66602a <=( a66601a  and  a66598a );
 a66605a <=( (not A265)  and  (not A236) );
 a66609a <=( A269  and  A267 );
 a66610a <=( A266  and  a66609a );
 a66611a <=( a66610a  and  a66605a );
 a66612a <=( a66611a  and  a66602a );
 a66615a <=( (not A169)  and  A170 );
 a66618a <=( (not A167)  and  (not A168) );
 a66619a <=( a66618a  and  a66615a );
 a66622a <=( A201  and  A166 );
 a66625a <=( (not A203)  and  (not A202) );
 a66626a <=( a66625a  and  a66622a );
 a66627a <=( a66626a  and  a66619a );
 a66630a <=( (not A233)  and  A232 );
 a66633a <=( (not A235)  and  (not A234) );
 a66634a <=( a66633a  and  a66630a );
 a66637a <=( A265  and  (not A236) );
 a66641a <=( A268  and  A267 );
 a66642a <=( (not A266)  and  a66641a );
 a66643a <=( a66642a  and  a66637a );
 a66644a <=( a66643a  and  a66634a );
 a66647a <=( (not A169)  and  A170 );
 a66650a <=( (not A167)  and  (not A168) );
 a66651a <=( a66650a  and  a66647a );
 a66654a <=( A201  and  A166 );
 a66657a <=( (not A203)  and  (not A202) );
 a66658a <=( a66657a  and  a66654a );
 a66659a <=( a66658a  and  a66651a );
 a66662a <=( (not A233)  and  A232 );
 a66665a <=( (not A235)  and  (not A234) );
 a66666a <=( a66665a  and  a66662a );
 a66669a <=( A265  and  (not A236) );
 a66673a <=( A269  and  A267 );
 a66674a <=( (not A266)  and  a66673a );
 a66675a <=( a66674a  and  a66669a );
 a66676a <=( a66675a  and  a66666a );
 a66679a <=( (not A169)  and  A170 );
 a66682a <=( (not A167)  and  (not A168) );
 a66683a <=( a66682a  and  a66679a );
 a66686a <=( (not A201)  and  A166 );
 a66689a <=( (not A232)  and  A202 );
 a66690a <=( a66689a  and  a66686a );
 a66691a <=( a66690a  and  a66683a );
 a66694a <=( (not A234)  and  A233 );
 a66697a <=( (not A236)  and  (not A235) );
 a66698a <=( a66697a  and  a66694a );
 a66701a <=( (not A299)  and  A298 );
 a66705a <=( (not A302)  and  (not A301) );
 a66706a <=( (not A300)  and  a66705a );
 a66707a <=( a66706a  and  a66701a );
 a66708a <=( a66707a  and  a66698a );
 a66711a <=( (not A169)  and  A170 );
 a66714a <=( (not A167)  and  (not A168) );
 a66715a <=( a66714a  and  a66711a );
 a66718a <=( (not A201)  and  A166 );
 a66721a <=( (not A232)  and  A202 );
 a66722a <=( a66721a  and  a66718a );
 a66723a <=( a66722a  and  a66715a );
 a66726a <=( (not A234)  and  A233 );
 a66729a <=( (not A236)  and  (not A235) );
 a66730a <=( a66729a  and  a66726a );
 a66733a <=( A299  and  (not A298) );
 a66737a <=( (not A302)  and  (not A301) );
 a66738a <=( (not A300)  and  a66737a );
 a66739a <=( a66738a  and  a66733a );
 a66740a <=( a66739a  and  a66730a );
 a66743a <=( (not A169)  and  A170 );
 a66746a <=( (not A167)  and  (not A168) );
 a66747a <=( a66746a  and  a66743a );
 a66750a <=( (not A201)  and  A166 );
 a66753a <=( (not A232)  and  A202 );
 a66754a <=( a66753a  and  a66750a );
 a66755a <=( a66754a  and  a66747a );
 a66758a <=( (not A234)  and  A233 );
 a66761a <=( (not A236)  and  (not A235) );
 a66762a <=( a66761a  and  a66758a );
 a66765a <=( A266  and  (not A265) );
 a66769a <=( (not A269)  and  (not A268) );
 a66770a <=( (not A267)  and  a66769a );
 a66771a <=( a66770a  and  a66765a );
 a66772a <=( a66771a  and  a66762a );
 a66775a <=( (not A169)  and  A170 );
 a66778a <=( (not A167)  and  (not A168) );
 a66779a <=( a66778a  and  a66775a );
 a66782a <=( (not A201)  and  A166 );
 a66785a <=( (not A232)  and  A202 );
 a66786a <=( a66785a  and  a66782a );
 a66787a <=( a66786a  and  a66779a );
 a66790a <=( (not A234)  and  A233 );
 a66793a <=( (not A236)  and  (not A235) );
 a66794a <=( a66793a  and  a66790a );
 a66797a <=( (not A266)  and  A265 );
 a66801a <=( (not A269)  and  (not A268) );
 a66802a <=( (not A267)  and  a66801a );
 a66803a <=( a66802a  and  a66797a );
 a66804a <=( a66803a  and  a66794a );
 a66807a <=( (not A169)  and  A170 );
 a66810a <=( (not A167)  and  (not A168) );
 a66811a <=( a66810a  and  a66807a );
 a66814a <=( (not A201)  and  A166 );
 a66817a <=( A232  and  A202 );
 a66818a <=( a66817a  and  a66814a );
 a66819a <=( a66818a  and  a66811a );
 a66822a <=( (not A234)  and  (not A233) );
 a66825a <=( (not A236)  and  (not A235) );
 a66826a <=( a66825a  and  a66822a );
 a66829a <=( (not A299)  and  A298 );
 a66833a <=( (not A302)  and  (not A301) );
 a66834a <=( (not A300)  and  a66833a );
 a66835a <=( a66834a  and  a66829a );
 a66836a <=( a66835a  and  a66826a );
 a66839a <=( (not A169)  and  A170 );
 a66842a <=( (not A167)  and  (not A168) );
 a66843a <=( a66842a  and  a66839a );
 a66846a <=( (not A201)  and  A166 );
 a66849a <=( A232  and  A202 );
 a66850a <=( a66849a  and  a66846a );
 a66851a <=( a66850a  and  a66843a );
 a66854a <=( (not A234)  and  (not A233) );
 a66857a <=( (not A236)  and  (not A235) );
 a66858a <=( a66857a  and  a66854a );
 a66861a <=( A299  and  (not A298) );
 a66865a <=( (not A302)  and  (not A301) );
 a66866a <=( (not A300)  and  a66865a );
 a66867a <=( a66866a  and  a66861a );
 a66868a <=( a66867a  and  a66858a );
 a66871a <=( (not A169)  and  A170 );
 a66874a <=( (not A167)  and  (not A168) );
 a66875a <=( a66874a  and  a66871a );
 a66878a <=( (not A201)  and  A166 );
 a66881a <=( A232  and  A202 );
 a66882a <=( a66881a  and  a66878a );
 a66883a <=( a66882a  and  a66875a );
 a66886a <=( (not A234)  and  (not A233) );
 a66889a <=( (not A236)  and  (not A235) );
 a66890a <=( a66889a  and  a66886a );
 a66893a <=( A266  and  (not A265) );
 a66897a <=( (not A269)  and  (not A268) );
 a66898a <=( (not A267)  and  a66897a );
 a66899a <=( a66898a  and  a66893a );
 a66900a <=( a66899a  and  a66890a );
 a66903a <=( (not A169)  and  A170 );
 a66906a <=( (not A167)  and  (not A168) );
 a66907a <=( a66906a  and  a66903a );
 a66910a <=( (not A201)  and  A166 );
 a66913a <=( A232  and  A202 );
 a66914a <=( a66913a  and  a66910a );
 a66915a <=( a66914a  and  a66907a );
 a66918a <=( (not A234)  and  (not A233) );
 a66921a <=( (not A236)  and  (not A235) );
 a66922a <=( a66921a  and  a66918a );
 a66925a <=( (not A266)  and  A265 );
 a66929a <=( (not A269)  and  (not A268) );
 a66930a <=( (not A267)  and  a66929a );
 a66931a <=( a66930a  and  a66925a );
 a66932a <=( a66931a  and  a66922a );
 a66935a <=( (not A169)  and  A170 );
 a66938a <=( (not A167)  and  (not A168) );
 a66939a <=( a66938a  and  a66935a );
 a66942a <=( (not A201)  and  A166 );
 a66945a <=( (not A232)  and  A203 );
 a66946a <=( a66945a  and  a66942a );
 a66947a <=( a66946a  and  a66939a );
 a66950a <=( (not A234)  and  A233 );
 a66953a <=( (not A236)  and  (not A235) );
 a66954a <=( a66953a  and  a66950a );
 a66957a <=( (not A299)  and  A298 );
 a66961a <=( (not A302)  and  (not A301) );
 a66962a <=( (not A300)  and  a66961a );
 a66963a <=( a66962a  and  a66957a );
 a66964a <=( a66963a  and  a66954a );
 a66967a <=( (not A169)  and  A170 );
 a66970a <=( (not A167)  and  (not A168) );
 a66971a <=( a66970a  and  a66967a );
 a66974a <=( (not A201)  and  A166 );
 a66977a <=( (not A232)  and  A203 );
 a66978a <=( a66977a  and  a66974a );
 a66979a <=( a66978a  and  a66971a );
 a66982a <=( (not A234)  and  A233 );
 a66985a <=( (not A236)  and  (not A235) );
 a66986a <=( a66985a  and  a66982a );
 a66989a <=( A299  and  (not A298) );
 a66993a <=( (not A302)  and  (not A301) );
 a66994a <=( (not A300)  and  a66993a );
 a66995a <=( a66994a  and  a66989a );
 a66996a <=( a66995a  and  a66986a );
 a66999a <=( (not A169)  and  A170 );
 a67002a <=( (not A167)  and  (not A168) );
 a67003a <=( a67002a  and  a66999a );
 a67006a <=( (not A201)  and  A166 );
 a67009a <=( (not A232)  and  A203 );
 a67010a <=( a67009a  and  a67006a );
 a67011a <=( a67010a  and  a67003a );
 a67014a <=( (not A234)  and  A233 );
 a67017a <=( (not A236)  and  (not A235) );
 a67018a <=( a67017a  and  a67014a );
 a67021a <=( A266  and  (not A265) );
 a67025a <=( (not A269)  and  (not A268) );
 a67026a <=( (not A267)  and  a67025a );
 a67027a <=( a67026a  and  a67021a );
 a67028a <=( a67027a  and  a67018a );
 a67031a <=( (not A169)  and  A170 );
 a67034a <=( (not A167)  and  (not A168) );
 a67035a <=( a67034a  and  a67031a );
 a67038a <=( (not A201)  and  A166 );
 a67041a <=( (not A232)  and  A203 );
 a67042a <=( a67041a  and  a67038a );
 a67043a <=( a67042a  and  a67035a );
 a67046a <=( (not A234)  and  A233 );
 a67049a <=( (not A236)  and  (not A235) );
 a67050a <=( a67049a  and  a67046a );
 a67053a <=( (not A266)  and  A265 );
 a67057a <=( (not A269)  and  (not A268) );
 a67058a <=( (not A267)  and  a67057a );
 a67059a <=( a67058a  and  a67053a );
 a67060a <=( a67059a  and  a67050a );
 a67063a <=( (not A169)  and  A170 );
 a67066a <=( (not A167)  and  (not A168) );
 a67067a <=( a67066a  and  a67063a );
 a67070a <=( (not A201)  and  A166 );
 a67073a <=( A232  and  A203 );
 a67074a <=( a67073a  and  a67070a );
 a67075a <=( a67074a  and  a67067a );
 a67078a <=( (not A234)  and  (not A233) );
 a67081a <=( (not A236)  and  (not A235) );
 a67082a <=( a67081a  and  a67078a );
 a67085a <=( (not A299)  and  A298 );
 a67089a <=( (not A302)  and  (not A301) );
 a67090a <=( (not A300)  and  a67089a );
 a67091a <=( a67090a  and  a67085a );
 a67092a <=( a67091a  and  a67082a );
 a67095a <=( (not A169)  and  A170 );
 a67098a <=( (not A167)  and  (not A168) );
 a67099a <=( a67098a  and  a67095a );
 a67102a <=( (not A201)  and  A166 );
 a67105a <=( A232  and  A203 );
 a67106a <=( a67105a  and  a67102a );
 a67107a <=( a67106a  and  a67099a );
 a67110a <=( (not A234)  and  (not A233) );
 a67113a <=( (not A236)  and  (not A235) );
 a67114a <=( a67113a  and  a67110a );
 a67117a <=( A299  and  (not A298) );
 a67121a <=( (not A302)  and  (not A301) );
 a67122a <=( (not A300)  and  a67121a );
 a67123a <=( a67122a  and  a67117a );
 a67124a <=( a67123a  and  a67114a );
 a67127a <=( (not A169)  and  A170 );
 a67130a <=( (not A167)  and  (not A168) );
 a67131a <=( a67130a  and  a67127a );
 a67134a <=( (not A201)  and  A166 );
 a67137a <=( A232  and  A203 );
 a67138a <=( a67137a  and  a67134a );
 a67139a <=( a67138a  and  a67131a );
 a67142a <=( (not A234)  and  (not A233) );
 a67145a <=( (not A236)  and  (not A235) );
 a67146a <=( a67145a  and  a67142a );
 a67149a <=( A266  and  (not A265) );
 a67153a <=( (not A269)  and  (not A268) );
 a67154a <=( (not A267)  and  a67153a );
 a67155a <=( a67154a  and  a67149a );
 a67156a <=( a67155a  and  a67146a );
 a67159a <=( (not A169)  and  A170 );
 a67162a <=( (not A167)  and  (not A168) );
 a67163a <=( a67162a  and  a67159a );
 a67166a <=( (not A201)  and  A166 );
 a67169a <=( A232  and  A203 );
 a67170a <=( a67169a  and  a67166a );
 a67171a <=( a67170a  and  a67163a );
 a67174a <=( (not A234)  and  (not A233) );
 a67177a <=( (not A236)  and  (not A235) );
 a67178a <=( a67177a  and  a67174a );
 a67181a <=( (not A266)  and  A265 );
 a67185a <=( (not A269)  and  (not A268) );
 a67186a <=( (not A267)  and  a67185a );
 a67187a <=( a67186a  and  a67181a );
 a67188a <=( a67187a  and  a67178a );
 a67191a <=( (not A169)  and  A170 );
 a67194a <=( (not A167)  and  (not A168) );
 a67195a <=( a67194a  and  a67191a );
 a67198a <=( A199  and  A166 );
 a67201a <=( (not A232)  and  A200 );
 a67202a <=( a67201a  and  a67198a );
 a67203a <=( a67202a  and  a67195a );
 a67206a <=( (not A234)  and  A233 );
 a67209a <=( (not A236)  and  (not A235) );
 a67210a <=( a67209a  and  a67206a );
 a67213a <=( (not A299)  and  A298 );
 a67217a <=( (not A302)  and  (not A301) );
 a67218a <=( (not A300)  and  a67217a );
 a67219a <=( a67218a  and  a67213a );
 a67220a <=( a67219a  and  a67210a );
 a67223a <=( (not A169)  and  A170 );
 a67226a <=( (not A167)  and  (not A168) );
 a67227a <=( a67226a  and  a67223a );
 a67230a <=( A199  and  A166 );
 a67233a <=( (not A232)  and  A200 );
 a67234a <=( a67233a  and  a67230a );
 a67235a <=( a67234a  and  a67227a );
 a67238a <=( (not A234)  and  A233 );
 a67241a <=( (not A236)  and  (not A235) );
 a67242a <=( a67241a  and  a67238a );
 a67245a <=( A299  and  (not A298) );
 a67249a <=( (not A302)  and  (not A301) );
 a67250a <=( (not A300)  and  a67249a );
 a67251a <=( a67250a  and  a67245a );
 a67252a <=( a67251a  and  a67242a );
 a67255a <=( (not A169)  and  A170 );
 a67258a <=( (not A167)  and  (not A168) );
 a67259a <=( a67258a  and  a67255a );
 a67262a <=( A199  and  A166 );
 a67265a <=( (not A232)  and  A200 );
 a67266a <=( a67265a  and  a67262a );
 a67267a <=( a67266a  and  a67259a );
 a67270a <=( (not A234)  and  A233 );
 a67273a <=( (not A236)  and  (not A235) );
 a67274a <=( a67273a  and  a67270a );
 a67277a <=( A266  and  (not A265) );
 a67281a <=( (not A269)  and  (not A268) );
 a67282a <=( (not A267)  and  a67281a );
 a67283a <=( a67282a  and  a67277a );
 a67284a <=( a67283a  and  a67274a );
 a67287a <=( (not A169)  and  A170 );
 a67290a <=( (not A167)  and  (not A168) );
 a67291a <=( a67290a  and  a67287a );
 a67294a <=( A199  and  A166 );
 a67297a <=( (not A232)  and  A200 );
 a67298a <=( a67297a  and  a67294a );
 a67299a <=( a67298a  and  a67291a );
 a67302a <=( (not A234)  and  A233 );
 a67305a <=( (not A236)  and  (not A235) );
 a67306a <=( a67305a  and  a67302a );
 a67309a <=( (not A266)  and  A265 );
 a67313a <=( (not A269)  and  (not A268) );
 a67314a <=( (not A267)  and  a67313a );
 a67315a <=( a67314a  and  a67309a );
 a67316a <=( a67315a  and  a67306a );
 a67319a <=( (not A169)  and  A170 );
 a67322a <=( (not A167)  and  (not A168) );
 a67323a <=( a67322a  and  a67319a );
 a67326a <=( A199  and  A166 );
 a67329a <=( A232  and  A200 );
 a67330a <=( a67329a  and  a67326a );
 a67331a <=( a67330a  and  a67323a );
 a67334a <=( (not A234)  and  (not A233) );
 a67337a <=( (not A236)  and  (not A235) );
 a67338a <=( a67337a  and  a67334a );
 a67341a <=( (not A299)  and  A298 );
 a67345a <=( (not A302)  and  (not A301) );
 a67346a <=( (not A300)  and  a67345a );
 a67347a <=( a67346a  and  a67341a );
 a67348a <=( a67347a  and  a67338a );
 a67351a <=( (not A169)  and  A170 );
 a67354a <=( (not A167)  and  (not A168) );
 a67355a <=( a67354a  and  a67351a );
 a67358a <=( A199  and  A166 );
 a67361a <=( A232  and  A200 );
 a67362a <=( a67361a  and  a67358a );
 a67363a <=( a67362a  and  a67355a );
 a67366a <=( (not A234)  and  (not A233) );
 a67369a <=( (not A236)  and  (not A235) );
 a67370a <=( a67369a  and  a67366a );
 a67373a <=( A299  and  (not A298) );
 a67377a <=( (not A302)  and  (not A301) );
 a67378a <=( (not A300)  and  a67377a );
 a67379a <=( a67378a  and  a67373a );
 a67380a <=( a67379a  and  a67370a );
 a67383a <=( (not A169)  and  A170 );
 a67386a <=( (not A167)  and  (not A168) );
 a67387a <=( a67386a  and  a67383a );
 a67390a <=( A199  and  A166 );
 a67393a <=( A232  and  A200 );
 a67394a <=( a67393a  and  a67390a );
 a67395a <=( a67394a  and  a67387a );
 a67398a <=( (not A234)  and  (not A233) );
 a67401a <=( (not A236)  and  (not A235) );
 a67402a <=( a67401a  and  a67398a );
 a67405a <=( A266  and  (not A265) );
 a67409a <=( (not A269)  and  (not A268) );
 a67410a <=( (not A267)  and  a67409a );
 a67411a <=( a67410a  and  a67405a );
 a67412a <=( a67411a  and  a67402a );
 a67415a <=( (not A169)  and  A170 );
 a67418a <=( (not A167)  and  (not A168) );
 a67419a <=( a67418a  and  a67415a );
 a67422a <=( A199  and  A166 );
 a67425a <=( A232  and  A200 );
 a67426a <=( a67425a  and  a67422a );
 a67427a <=( a67426a  and  a67419a );
 a67430a <=( (not A234)  and  (not A233) );
 a67433a <=( (not A236)  and  (not A235) );
 a67434a <=( a67433a  and  a67430a );
 a67437a <=( (not A266)  and  A265 );
 a67441a <=( (not A269)  and  (not A268) );
 a67442a <=( (not A267)  and  a67441a );
 a67443a <=( a67442a  and  a67437a );
 a67444a <=( a67443a  and  a67434a );
 a67447a <=( (not A169)  and  A170 );
 a67450a <=( (not A167)  and  (not A168) );
 a67451a <=( a67450a  and  a67447a );
 a67454a <=( (not A199)  and  A166 );
 a67457a <=( (not A232)  and  (not A200) );
 a67458a <=( a67457a  and  a67454a );
 a67459a <=( a67458a  and  a67451a );
 a67462a <=( (not A234)  and  A233 );
 a67465a <=( (not A236)  and  (not A235) );
 a67466a <=( a67465a  and  a67462a );
 a67469a <=( (not A299)  and  A298 );
 a67473a <=( (not A302)  and  (not A301) );
 a67474a <=( (not A300)  and  a67473a );
 a67475a <=( a67474a  and  a67469a );
 a67476a <=( a67475a  and  a67466a );
 a67479a <=( (not A169)  and  A170 );
 a67482a <=( (not A167)  and  (not A168) );
 a67483a <=( a67482a  and  a67479a );
 a67486a <=( (not A199)  and  A166 );
 a67489a <=( (not A232)  and  (not A200) );
 a67490a <=( a67489a  and  a67486a );
 a67491a <=( a67490a  and  a67483a );
 a67494a <=( (not A234)  and  A233 );
 a67497a <=( (not A236)  and  (not A235) );
 a67498a <=( a67497a  and  a67494a );
 a67501a <=( A299  and  (not A298) );
 a67505a <=( (not A302)  and  (not A301) );
 a67506a <=( (not A300)  and  a67505a );
 a67507a <=( a67506a  and  a67501a );
 a67508a <=( a67507a  and  a67498a );
 a67511a <=( (not A169)  and  A170 );
 a67514a <=( (not A167)  and  (not A168) );
 a67515a <=( a67514a  and  a67511a );
 a67518a <=( (not A199)  and  A166 );
 a67521a <=( (not A232)  and  (not A200) );
 a67522a <=( a67521a  and  a67518a );
 a67523a <=( a67522a  and  a67515a );
 a67526a <=( (not A234)  and  A233 );
 a67529a <=( (not A236)  and  (not A235) );
 a67530a <=( a67529a  and  a67526a );
 a67533a <=( A266  and  (not A265) );
 a67537a <=( (not A269)  and  (not A268) );
 a67538a <=( (not A267)  and  a67537a );
 a67539a <=( a67538a  and  a67533a );
 a67540a <=( a67539a  and  a67530a );
 a67543a <=( (not A169)  and  A170 );
 a67546a <=( (not A167)  and  (not A168) );
 a67547a <=( a67546a  and  a67543a );
 a67550a <=( (not A199)  and  A166 );
 a67553a <=( (not A232)  and  (not A200) );
 a67554a <=( a67553a  and  a67550a );
 a67555a <=( a67554a  and  a67547a );
 a67558a <=( (not A234)  and  A233 );
 a67561a <=( (not A236)  and  (not A235) );
 a67562a <=( a67561a  and  a67558a );
 a67565a <=( (not A266)  and  A265 );
 a67569a <=( (not A269)  and  (not A268) );
 a67570a <=( (not A267)  and  a67569a );
 a67571a <=( a67570a  and  a67565a );
 a67572a <=( a67571a  and  a67562a );
 a67575a <=( (not A169)  and  A170 );
 a67578a <=( (not A167)  and  (not A168) );
 a67579a <=( a67578a  and  a67575a );
 a67582a <=( (not A199)  and  A166 );
 a67585a <=( A232  and  (not A200) );
 a67586a <=( a67585a  and  a67582a );
 a67587a <=( a67586a  and  a67579a );
 a67590a <=( (not A234)  and  (not A233) );
 a67593a <=( (not A236)  and  (not A235) );
 a67594a <=( a67593a  and  a67590a );
 a67597a <=( (not A299)  and  A298 );
 a67601a <=( (not A302)  and  (not A301) );
 a67602a <=( (not A300)  and  a67601a );
 a67603a <=( a67602a  and  a67597a );
 a67604a <=( a67603a  and  a67594a );
 a67607a <=( (not A169)  and  A170 );
 a67610a <=( (not A167)  and  (not A168) );
 a67611a <=( a67610a  and  a67607a );
 a67614a <=( (not A199)  and  A166 );
 a67617a <=( A232  and  (not A200) );
 a67618a <=( a67617a  and  a67614a );
 a67619a <=( a67618a  and  a67611a );
 a67622a <=( (not A234)  and  (not A233) );
 a67625a <=( (not A236)  and  (not A235) );
 a67626a <=( a67625a  and  a67622a );
 a67629a <=( A299  and  (not A298) );
 a67633a <=( (not A302)  and  (not A301) );
 a67634a <=( (not A300)  and  a67633a );
 a67635a <=( a67634a  and  a67629a );
 a67636a <=( a67635a  and  a67626a );
 a67639a <=( (not A169)  and  A170 );
 a67642a <=( (not A167)  and  (not A168) );
 a67643a <=( a67642a  and  a67639a );
 a67646a <=( (not A199)  and  A166 );
 a67649a <=( A232  and  (not A200) );
 a67650a <=( a67649a  and  a67646a );
 a67651a <=( a67650a  and  a67643a );
 a67654a <=( (not A234)  and  (not A233) );
 a67657a <=( (not A236)  and  (not A235) );
 a67658a <=( a67657a  and  a67654a );
 a67661a <=( A266  and  (not A265) );
 a67665a <=( (not A269)  and  (not A268) );
 a67666a <=( (not A267)  and  a67665a );
 a67667a <=( a67666a  and  a67661a );
 a67668a <=( a67667a  and  a67658a );
 a67671a <=( (not A169)  and  A170 );
 a67674a <=( (not A167)  and  (not A168) );
 a67675a <=( a67674a  and  a67671a );
 a67678a <=( (not A199)  and  A166 );
 a67681a <=( A232  and  (not A200) );
 a67682a <=( a67681a  and  a67678a );
 a67683a <=( a67682a  and  a67675a );
 a67686a <=( (not A234)  and  (not A233) );
 a67689a <=( (not A236)  and  (not A235) );
 a67690a <=( a67689a  and  a67686a );
 a67693a <=( (not A266)  and  A265 );
 a67697a <=( (not A269)  and  (not A268) );
 a67698a <=( (not A267)  and  a67697a );
 a67699a <=( a67698a  and  a67693a );
 a67700a <=( a67699a  and  a67690a );
 a67703a <=( (not A169)  and  A170 );
 a67706a <=( A167  and  (not A168) );
 a67707a <=( a67706a  and  a67703a );
 a67710a <=( A201  and  (not A166) );
 a67714a <=( (not A232)  and  (not A203) );
 a67715a <=( (not A202)  and  a67714a );
 a67716a <=( a67715a  and  a67710a );
 a67717a <=( a67716a  and  a67707a );
 a67720a <=( (not A234)  and  A233 );
 a67723a <=( (not A236)  and  (not A235) );
 a67724a <=( a67723a  and  a67720a );
 a67727a <=( (not A299)  and  A298 );
 a67731a <=( (not A302)  and  (not A301) );
 a67732a <=( (not A300)  and  a67731a );
 a67733a <=( a67732a  and  a67727a );
 a67734a <=( a67733a  and  a67724a );
 a67737a <=( (not A169)  and  A170 );
 a67740a <=( A167  and  (not A168) );
 a67741a <=( a67740a  and  a67737a );
 a67744a <=( A201  and  (not A166) );
 a67748a <=( (not A232)  and  (not A203) );
 a67749a <=( (not A202)  and  a67748a );
 a67750a <=( a67749a  and  a67744a );
 a67751a <=( a67750a  and  a67741a );
 a67754a <=( (not A234)  and  A233 );
 a67757a <=( (not A236)  and  (not A235) );
 a67758a <=( a67757a  and  a67754a );
 a67761a <=( A299  and  (not A298) );
 a67765a <=( (not A302)  and  (not A301) );
 a67766a <=( (not A300)  and  a67765a );
 a67767a <=( a67766a  and  a67761a );
 a67768a <=( a67767a  and  a67758a );
 a67771a <=( (not A169)  and  A170 );
 a67774a <=( A167  and  (not A168) );
 a67775a <=( a67774a  and  a67771a );
 a67778a <=( A201  and  (not A166) );
 a67782a <=( (not A232)  and  (not A203) );
 a67783a <=( (not A202)  and  a67782a );
 a67784a <=( a67783a  and  a67778a );
 a67785a <=( a67784a  and  a67775a );
 a67788a <=( (not A234)  and  A233 );
 a67791a <=( (not A236)  and  (not A235) );
 a67792a <=( a67791a  and  a67788a );
 a67795a <=( A266  and  (not A265) );
 a67799a <=( (not A269)  and  (not A268) );
 a67800a <=( (not A267)  and  a67799a );
 a67801a <=( a67800a  and  a67795a );
 a67802a <=( a67801a  and  a67792a );
 a67805a <=( (not A169)  and  A170 );
 a67808a <=( A167  and  (not A168) );
 a67809a <=( a67808a  and  a67805a );
 a67812a <=( A201  and  (not A166) );
 a67816a <=( (not A232)  and  (not A203) );
 a67817a <=( (not A202)  and  a67816a );
 a67818a <=( a67817a  and  a67812a );
 a67819a <=( a67818a  and  a67809a );
 a67822a <=( (not A234)  and  A233 );
 a67825a <=( (not A236)  and  (not A235) );
 a67826a <=( a67825a  and  a67822a );
 a67829a <=( (not A266)  and  A265 );
 a67833a <=( (not A269)  and  (not A268) );
 a67834a <=( (not A267)  and  a67833a );
 a67835a <=( a67834a  and  a67829a );
 a67836a <=( a67835a  and  a67826a );
 a67839a <=( (not A169)  and  A170 );
 a67842a <=( A167  and  (not A168) );
 a67843a <=( a67842a  and  a67839a );
 a67846a <=( A201  and  (not A166) );
 a67850a <=( A232  and  (not A203) );
 a67851a <=( (not A202)  and  a67850a );
 a67852a <=( a67851a  and  a67846a );
 a67853a <=( a67852a  and  a67843a );
 a67856a <=( (not A234)  and  (not A233) );
 a67859a <=( (not A236)  and  (not A235) );
 a67860a <=( a67859a  and  a67856a );
 a67863a <=( (not A299)  and  A298 );
 a67867a <=( (not A302)  and  (not A301) );
 a67868a <=( (not A300)  and  a67867a );
 a67869a <=( a67868a  and  a67863a );
 a67870a <=( a67869a  and  a67860a );
 a67873a <=( (not A169)  and  A170 );
 a67876a <=( A167  and  (not A168) );
 a67877a <=( a67876a  and  a67873a );
 a67880a <=( A201  and  (not A166) );
 a67884a <=( A232  and  (not A203) );
 a67885a <=( (not A202)  and  a67884a );
 a67886a <=( a67885a  and  a67880a );
 a67887a <=( a67886a  and  a67877a );
 a67890a <=( (not A234)  and  (not A233) );
 a67893a <=( (not A236)  and  (not A235) );
 a67894a <=( a67893a  and  a67890a );
 a67897a <=( A299  and  (not A298) );
 a67901a <=( (not A302)  and  (not A301) );
 a67902a <=( (not A300)  and  a67901a );
 a67903a <=( a67902a  and  a67897a );
 a67904a <=( a67903a  and  a67894a );
 a67907a <=( (not A169)  and  A170 );
 a67910a <=( A167  and  (not A168) );
 a67911a <=( a67910a  and  a67907a );
 a67914a <=( A201  and  (not A166) );
 a67918a <=( A232  and  (not A203) );
 a67919a <=( (not A202)  and  a67918a );
 a67920a <=( a67919a  and  a67914a );
 a67921a <=( a67920a  and  a67911a );
 a67924a <=( (not A234)  and  (not A233) );
 a67927a <=( (not A236)  and  (not A235) );
 a67928a <=( a67927a  and  a67924a );
 a67931a <=( A266  and  (not A265) );
 a67935a <=( (not A269)  and  (not A268) );
 a67936a <=( (not A267)  and  a67935a );
 a67937a <=( a67936a  and  a67931a );
 a67938a <=( a67937a  and  a67928a );
 a67941a <=( (not A169)  and  A170 );
 a67944a <=( A167  and  (not A168) );
 a67945a <=( a67944a  and  a67941a );
 a67948a <=( A201  and  (not A166) );
 a67952a <=( A232  and  (not A203) );
 a67953a <=( (not A202)  and  a67952a );
 a67954a <=( a67953a  and  a67948a );
 a67955a <=( a67954a  and  a67945a );
 a67958a <=( (not A234)  and  (not A233) );
 a67961a <=( (not A236)  and  (not A235) );
 a67962a <=( a67961a  and  a67958a );
 a67965a <=( (not A266)  and  A265 );
 a67969a <=( (not A269)  and  (not A268) );
 a67970a <=( (not A267)  and  a67969a );
 a67971a <=( a67970a  and  a67965a );
 a67972a <=( a67971a  and  a67962a );
 a67975a <=( (not A169)  and  A170 );
 a67978a <=( (not A167)  and  (not A168) );
 a67979a <=( a67978a  and  a67975a );
 a67982a <=( A201  and  A166 );
 a67986a <=( (not A232)  and  (not A203) );
 a67987a <=( (not A202)  and  a67986a );
 a67988a <=( a67987a  and  a67982a );
 a67989a <=( a67988a  and  a67979a );
 a67992a <=( (not A234)  and  A233 );
 a67995a <=( (not A236)  and  (not A235) );
 a67996a <=( a67995a  and  a67992a );
 a67999a <=( (not A299)  and  A298 );
 a68003a <=( (not A302)  and  (not A301) );
 a68004a <=( (not A300)  and  a68003a );
 a68005a <=( a68004a  and  a67999a );
 a68006a <=( a68005a  and  a67996a );
 a68009a <=( (not A169)  and  A170 );
 a68012a <=( (not A167)  and  (not A168) );
 a68013a <=( a68012a  and  a68009a );
 a68016a <=( A201  and  A166 );
 a68020a <=( (not A232)  and  (not A203) );
 a68021a <=( (not A202)  and  a68020a );
 a68022a <=( a68021a  and  a68016a );
 a68023a <=( a68022a  and  a68013a );
 a68026a <=( (not A234)  and  A233 );
 a68029a <=( (not A236)  and  (not A235) );
 a68030a <=( a68029a  and  a68026a );
 a68033a <=( A299  and  (not A298) );
 a68037a <=( (not A302)  and  (not A301) );
 a68038a <=( (not A300)  and  a68037a );
 a68039a <=( a68038a  and  a68033a );
 a68040a <=( a68039a  and  a68030a );
 a68043a <=( (not A169)  and  A170 );
 a68046a <=( (not A167)  and  (not A168) );
 a68047a <=( a68046a  and  a68043a );
 a68050a <=( A201  and  A166 );
 a68054a <=( (not A232)  and  (not A203) );
 a68055a <=( (not A202)  and  a68054a );
 a68056a <=( a68055a  and  a68050a );
 a68057a <=( a68056a  and  a68047a );
 a68060a <=( (not A234)  and  A233 );
 a68063a <=( (not A236)  and  (not A235) );
 a68064a <=( a68063a  and  a68060a );
 a68067a <=( A266  and  (not A265) );
 a68071a <=( (not A269)  and  (not A268) );
 a68072a <=( (not A267)  and  a68071a );
 a68073a <=( a68072a  and  a68067a );
 a68074a <=( a68073a  and  a68064a );
 a68077a <=( (not A169)  and  A170 );
 a68080a <=( (not A167)  and  (not A168) );
 a68081a <=( a68080a  and  a68077a );
 a68084a <=( A201  and  A166 );
 a68088a <=( (not A232)  and  (not A203) );
 a68089a <=( (not A202)  and  a68088a );
 a68090a <=( a68089a  and  a68084a );
 a68091a <=( a68090a  and  a68081a );
 a68094a <=( (not A234)  and  A233 );
 a68097a <=( (not A236)  and  (not A235) );
 a68098a <=( a68097a  and  a68094a );
 a68101a <=( (not A266)  and  A265 );
 a68105a <=( (not A269)  and  (not A268) );
 a68106a <=( (not A267)  and  a68105a );
 a68107a <=( a68106a  and  a68101a );
 a68108a <=( a68107a  and  a68098a );
 a68111a <=( (not A169)  and  A170 );
 a68114a <=( (not A167)  and  (not A168) );
 a68115a <=( a68114a  and  a68111a );
 a68118a <=( A201  and  A166 );
 a68122a <=( A232  and  (not A203) );
 a68123a <=( (not A202)  and  a68122a );
 a68124a <=( a68123a  and  a68118a );
 a68125a <=( a68124a  and  a68115a );
 a68128a <=( (not A234)  and  (not A233) );
 a68131a <=( (not A236)  and  (not A235) );
 a68132a <=( a68131a  and  a68128a );
 a68135a <=( (not A299)  and  A298 );
 a68139a <=( (not A302)  and  (not A301) );
 a68140a <=( (not A300)  and  a68139a );
 a68141a <=( a68140a  and  a68135a );
 a68142a <=( a68141a  and  a68132a );
 a68145a <=( (not A169)  and  A170 );
 a68148a <=( (not A167)  and  (not A168) );
 a68149a <=( a68148a  and  a68145a );
 a68152a <=( A201  and  A166 );
 a68156a <=( A232  and  (not A203) );
 a68157a <=( (not A202)  and  a68156a );
 a68158a <=( a68157a  and  a68152a );
 a68159a <=( a68158a  and  a68149a );
 a68162a <=( (not A234)  and  (not A233) );
 a68165a <=( (not A236)  and  (not A235) );
 a68166a <=( a68165a  and  a68162a );
 a68169a <=( A299  and  (not A298) );
 a68173a <=( (not A302)  and  (not A301) );
 a68174a <=( (not A300)  and  a68173a );
 a68175a <=( a68174a  and  a68169a );
 a68176a <=( a68175a  and  a68166a );
 a68179a <=( (not A169)  and  A170 );
 a68182a <=( (not A167)  and  (not A168) );
 a68183a <=( a68182a  and  a68179a );
 a68186a <=( A201  and  A166 );
 a68190a <=( A232  and  (not A203) );
 a68191a <=( (not A202)  and  a68190a );
 a68192a <=( a68191a  and  a68186a );
 a68193a <=( a68192a  and  a68183a );
 a68196a <=( (not A234)  and  (not A233) );
 a68199a <=( (not A236)  and  (not A235) );
 a68200a <=( a68199a  and  a68196a );
 a68203a <=( A266  and  (not A265) );
 a68207a <=( (not A269)  and  (not A268) );
 a68208a <=( (not A267)  and  a68207a );
 a68209a <=( a68208a  and  a68203a );
 a68210a <=( a68209a  and  a68200a );
 a68213a <=( (not A169)  and  A170 );
 a68216a <=( (not A167)  and  (not A168) );
 a68217a <=( a68216a  and  a68213a );
 a68220a <=( A201  and  A166 );
 a68224a <=( A232  and  (not A203) );
 a68225a <=( (not A202)  and  a68224a );
 a68226a <=( a68225a  and  a68220a );
 a68227a <=( a68226a  and  a68217a );
 a68230a <=( (not A234)  and  (not A233) );
 a68233a <=( (not A236)  and  (not A235) );
 a68234a <=( a68233a  and  a68230a );
 a68237a <=( (not A266)  and  A265 );
 a68241a <=( (not A269)  and  (not A268) );
 a68242a <=( (not A267)  and  a68241a );
 a68243a <=( a68242a  and  a68237a );
 a68244a <=( a68243a  and  a68234a );


end x25_2x_behav;
