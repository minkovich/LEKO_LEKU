Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_6x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A109: buffer std_logic
);
end x25_6x;

architecture x25_6x_behav of x25_6x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2196a,a2197a,a2198a,a2199a,a2200a,a2201a,a2202a,a2203a,a2204a,a2205a,a2206a,a2207a,a2208a,a2209a,a2210a,a2211a,a2212a,a2213a,a2214a,a2215a,a2216a,a2217a,a2218a,a2219a,a2220a,a2221a,a2222a,a2223a,a2224a,a2225a,a2226a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2237a,a2238a,a2239a,a2240a,a2241a,a2242a,a2243a,a2244a,a2245a,a2246a,a2247a,a2248a,a2249a,a2250a,a2251a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2258a,a2259a,a2260a,a2261a,a2262a,a2263a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2271a,a2272a,a2273a,a2274a,a2275a,a2276a,a2277a,a2278a,a2279a,a2280a,a2281a,a2282a,a2283a,a2284a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2297a,a2298a,a2299a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2306a,a2307a,a2308a,a2309a,a2310a,a2311a,a2312a,a2313a,a2314a,a2315a,a2316a,a2317a,a2318a,a2319a,a2320a,a2321a,a2322a,a2323a,a2324a,a2325a,a2326a,a2327a,a2328a,a2329a,a2330a,a2331a,a2332a,a2333a,a2334a,a2335a,a2336a,a2337a,a2338a,a2339a,a2340a,a2341a,a2342a,a2343a,a2344a,a2345a,a2346a,a2347a,a2348a,a2349a,a2350a,a2351a,a2352a,a2353a,a2354a,a2355a,a2356a,a2357a,a2358a,a2359a,a2360a,a2361a,a2362a,a2363a,a2364a,a2365a,a2366a,a2367a,a2368a,a2369a,a2370a,a2371a,a2372a,a2373a,a2374a,a2375a,a2376a,a2377a,a2378a,a2379a,a2380a,a2381a,a2382a,a2383a,a2384a,a2385a,a2386a,a2387a,a2388a,a2389a,a2390a,a2391a,a2392a,a2393a,a2394a,a2395a,a2396a,a2397a,a2398a,a2399a,a2400a,a2401a,a2402a,a2403a,a2404a,a2405a,a2406a,a2407a,a2408a,a2409a,a2410a,a2411a,a2412a,a2413a,a2414a,a2415a,a2416a,a2417a,a2418a,a2419a,a2420a,a2421a,a2422a,a2423a,a2424a,a2425a,a2426a,a2427a,a2428a,a2429a,a2430a,a2431a,a2432a,a2433a,a2434a,a2435a,a2436a,a2437a,a2438a,a2439a,a2440a,a2441a,a2442a,a2443a,a2444a,a2445a,a2446a,a2447a,a2448a,a2449a,a2450a,a2451a,a2452a,a2453a,a2454a,a2455a,a2456a,a2457a,a2458a,a2459a,a2460a,a2461a,a2462a,a2463a,a2464a,a2465a,a2466a,a2467a,a2468a,a2469a,a2470a,a2471a,a2472a,a2473a,a2474a,a2475a,a2476a,a2477a,a2478a,a2479a,a2480a,a2481a,a2482a,a2483a,a2484a,a2485a,a2486a,a2487a,a2488a,a2489a,a2490a,a2491a,a2492a,a2493a,a2494a,a2495a,a2496a,a2497a,a2498a,a2499a,a2500a,a2501a,a2502a,a2503a,a2504a,a2505a,a2506a,a2507a,a2508a,a2509a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2516a,a2517a,a2518a,a2519a,a2520a,a2521a,a2522a,a2523a,a2524a,a2525a,a2526a,a2527a,a2528a,a2529a,a2530a,a2531a,a2532a,a2533a,a2534a,a2535a,a2536a,a2537a,a2538a,a2539a,a2540a,a2541a,a2542a,a2543a,a2544a,a2545a,a2546a,a2547a,a2548a,a2549a,a2550a,a2551a,a2552a,a2553a,a2554a,a2555a,a2556a,a2557a,a2558a,a2559a,a2560a,a2561a,a2562a,a2563a,a2564a,a2565a,a2566a,a2567a,a2568a,a2569a,a2570a,a2571a,a2572a,a2573a,a2574a,a2575a,a2576a,a2577a,a2578a,a2579a,a2580a,a2581a,a2582a,a2583a,a2584a,a2585a,a2586a,a2587a,a2588a,a2589a,a2590a,a2591a,a2592a,a2593a,a2594a,a2595a,a2596a,a2597a,a2598a,a2599a,a2600a,a2601a,a2602a,a2603a,a2604a,a2605a,a2606a,a2607a,a2608a,a2609a,a2610a,a2611a,a2612a,a2613a,a2614a,a2615a,a2616a,a2617a,a2618a,a2619a,a2620a,a2621a,a2622a,a2623a,a2624a,a2625a,a2626a,a2627a,a2628a,a2629a,a2630a,a2631a,a2632a,a2633a,a2634a,a2635a,a2636a,a2637a,a2638a,a2639a,a2640a,a2641a,a2642a,a2643a,a2644a,a2645a,a2646a,a2647a,a2648a,a2649a,a2650a,a2651a,a2652a,a2653a,a2654a,a2655a,a2656a,a2657a,a2658a,a2659a,a2660a,a2661a,a2662a,a2663a,a2664a,a2665a,a2666a,a2667a,a2668a,a2669a,a2670a,a2671a,a2672a,a2673a,a2674a,a2675a,a2676a,a2677a,a2678a,a2679a,a2680a,a2681a,a2682a,a2683a,a2684a,a2685a,a2686a,a2687a,a2688a,a2689a,a2690a,a2691a,a2692a,a2693a,a2694a,a2695a,a2696a,a2697a,a2698a,a2699a,a2700a,a2701a,a2702a,a2703a,a2704a,a2705a,a2706a,a2707a,a2708a,a2709a,a2710a,a2711a,a2712a,a2713a,a2714a,a2715a,a2716a,a2717a,a2718a,a2719a,a2720a,a2721a,a2722a,a2723a,a2724a,a2725a,a2726a,a2727a,a2728a,a2729a,a2730a,a2731a,a2732a,a2733a,a2734a,a2735a,a2736a,a2737a,a2738a,a2739a,a2740a,a2741a,a2742a,a2743a,a2744a,a2745a,a2746a,a2747a,a2748a,a2749a,a2750a,a2751a,a2752a,a2753a,a2754a,a2755a,a2756a,a2757a,a2758a,a2759a,a2760a,a2761a,a2762a,a2763a,a2764a,a2765a,a2766a,a2767a,a2768a,a2769a,a2770a,a2771a,a2772a,a2773a,a2774a,a2775a,a2776a,a2777a,a2778a,a2779a,a2780a,a2781a,a2782a,a2783a,a2784a,a2785a,a2786a,a2787a,a2788a,a2789a,a2790a,a2791a,a2792a,a2793a,a2794a,a2795a,a2796a,a2797a,a2798a,a2799a,a2800a,a2801a,a2802a,a2803a,a2804a,a2805a,a2806a,a2807a,a2808a,a2809a,a2810a,a2811a,a2812a,a2813a,a2814a,a2815a,a2816a,a2817a,a2818a,a2819a,a2820a,a2821a,a2822a,a2823a,a2824a,a2825a,a2826a,a2827a,a2828a,a2829a,a2830a,a2831a,a2832a,a2833a,a2834a,a2835a,a2836a,a2837a,a2838a,a2839a,a2840a,a2841a,a2842a,a2843a,a2844a,a2845a,a2846a,a2847a,a2848a,a2849a,a2850a,a2851a,a2852a,a2853a,a2854a,a2855a,a2856a,a2857a,a2858a,a2859a,a2860a,a2861a,a2862a,a2863a,a2864a,a2865a,a2866a,a2867a,a2868a,a2869a,a2870a,a2871a,a2872a,a2873a,a2874a,a2875a,a2876a,a2877a,a2878a,a2879a,a2880a,a2881a,a2882a,a2883a,a2884a,a2885a,a2886a,a2887a,a2888a,a2889a,a2890a,a2891a,a2892a,a2893a,a2894a,a2895a,a2896a,a2897a,a2898a,a2899a,a2900a,a2901a,a2902a,a2903a,a2904a,a2905a,a2906a,a2907a,a2908a,a2909a,a2910a,a2911a,a2912a,a2913a,a2914a,a2915a,a2916a,a2917a,a2918a,a2919a,a2920a,a2921a,a2922a,a2923a,a2924a,a2925a,a2926a,a2927a,a2928a,a2929a,a2930a,a2931a,a2932a,a2933a,a2934a,a2935a,a2936a,a2937a,a2938a,a2939a,a2940a,a2941a,a2942a,a2943a,a2944a,a2945a,a2946a,a2947a,a2948a,a2949a,a2950a,a2951a,a2952a,a2953a,a2954a,a2955a,a2956a,a2957a,a2958a,a2959a,a2960a,a2961a,a2962a,a2963a,a2964a,a2965a,a2966a,a2967a,a2968a,a2969a,a2970a,a2971a,a2972a,a2973a,a2974a,a2975a,a2976a,a2977a,a2978a,a2979a,a2980a,a2981a,a2982a,a2983a,a2984a,a2985a,a2986a,a2987a,a2988a,a2989a,a2990a,a2991a,a2992a,a2993a,a2994a,a2995a,a2996a,a2997a,a2998a,a2999a,a3000a,a3001a,a3002a,a3003a,a3004a,a3005a,a3006a,a3007a,a3008a,a3009a,a3010a,a3011a,a3012a,a3013a,a3014a,a3015a,a3016a,a3017a,a3018a,a3019a,a3020a,a3021a,a3022a,a3023a,a3024a,a3025a,a3026a,a3027a,a3028a,a3029a,a3030a,a3031a,a3032a,a3033a,a3034a,a3035a,a3036a,a3037a,a3038a,a3039a,a3040a,a3041a,a3042a,a3043a,a3044a,a3045a,a3046a,a3047a,a3048a,a3049a,a3050a,a3051a,a3052a,a3053a,a3054a,a3055a,a3056a,a3057a,a3058a,a3059a,a3060a,a3061a,a3062a,a3063a,a3064a,a3065a,a3066a,a3067a,a3068a,a3069a,a3070a,a3071a,a3072a,a3073a,a3074a,a3075a,a3076a,a3077a,a3078a,a3079a,a3080a,a3081a,a3082a,a3083a,a3084a,a3085a,a3086a,a3087a,a3088a,a3089a,a3090a,a3091a,a3092a,a3093a,a3094a,a3095a,a3096a,a3097a,a3098a,a3099a,a3100a,a3101a,a3102a,a3103a,a3104a,a3105a,a3106a,a3107a,a3108a,a3109a,a3110a,a3111a,a3112a,a3113a,a3114a,a3115a,a3116a,a3117a,a3118a,a3119a,a3120a,a3121a,a3122a,a3123a,a3124a,a3125a,a3126a,a3127a,a3128a,a3129a,a3130a,a3131a,a3132a,a3133a,a3134a,a3135a,a3136a,a3137a,a3138a,a3139a,a3140a,a3141a,a3142a,a3143a,a3144a,a3145a,a3146a,a3147a,a3148a,a3149a,a3150a,a3151a,a3152a,a3153a,a3154a,a3155a,a3156a,a3157a,a3158a,a3159a,a3160a,a3161a,a3162a,a3163a,a3164a,a3165a,a3166a,a3167a,a3168a,a3169a,a3170a,a3171a,a3172a,a3173a,a3174a,a3175a,a3176a,a3177a,a3178a,a3179a,a3180a,a3181a,a3182a,a3183a,a3184a,a3185a,a3186a,a3187a,a3188a,a3189a,a3190a,a3191a,a3192a,a3193a,a3194a,a3195a,a3196a,a3197a,a3198a,a3199a,a3200a,a3201a,a3202a,a3203a,a3204a,a3205a,a3206a,a3207a,a3208a,a3209a,a3210a,a3211a,a3212a,a3213a,a3214a,a3215a,a3216a,a3217a,a3218a,a3219a,a3220a,a3221a,a3222a,a3223a,a3224a,a3225a,a3226a,a3227a,a3228a,a3229a,a3230a,a3231a,a3232a,a3233a,a3234a,a3235a,a3236a,a3237a,a3238a,a3239a,a3240a,a3241a,a3242a,a3243a,a3244a,a3245a,a3246a,a3247a,a3248a,a3249a,a3250a,a3251a,a3252a,a3253a,a3254a,a3255a,a3256a,a3257a,a3258a,a3259a,a3260a,a3261a,a3262a,a3263a,a3264a,a3265a,a3266a,a3267a,a3268a,a3269a,a3270a,a3271a,a3272a,a3273a,a3274a,a3275a,a3276a,a3277a,a3278a,a3279a,a3280a,a3281a,a3282a,a3283a,a3284a,a3285a,a3286a,a3287a,a3288a,a3289a,a3290a,a3291a,a3292a,a3293a,a3294a,a3295a,a3296a,a3297a,a3298a,a3299a,a3300a,a3301a,a3302a,a3303a,a3304a,a3305a,a3306a,a3307a,a3308a,a3309a,a3310a,a3311a,a3312a,a3313a,a3314a,a3315a,a3316a,a3317a,a3318a,a3319a,a3320a,a3321a,a3322a,a3323a,a3324a,a3325a,a3326a,a3327a,a3328a,a3329a,a3330a,a3331a,a3332a,a3333a,a3334a,a3335a,a3336a,a3337a,a3338a,a3339a,a3340a,a3341a,a3342a,a3343a,a3344a,a3345a,a3346a,a3347a,a3348a,a3349a,a3350a,a3351a,a3352a,a3353a,a3354a,a3355a,a3356a,a3357a,a3358a,a3359a,a3360a,a3361a,a3362a,a3363a,a3364a,a3365a,a3366a,a3367a,a3368a,a3369a,a3370a,a3371a,a3372a,a3373a,a3374a,a3375a,a3376a,a3377a,a3378a,a3379a,a3380a,a3381a,a3382a,a3383a,a3384a,a3385a,a3386a,a3387a,a3388a,a3389a,a3390a,a3391a,a3392a,a3393a,a3394a,a3395a,a3396a,a3397a,a3398a,a3399a,a3400a,a3401a,a3402a,a3403a,a3404a,a3405a,a3406a,a3407a,a3408a,a3409a,a3410a,a3411a,a3412a,a3413a,a3414a,a3415a,a3416a,a3417a,a3418a,a3419a,a3420a,a3421a,a3422a,a3423a,a3424a,a3425a,a3426a,a3427a,a3428a,a3429a,a3430a,a3431a,a3432a,a3433a,a3434a,a3435a,a3436a,a3437a,a3438a,a3439a,a3440a,a3441a,a3442a,a3443a,a3444a,a3445a,a3446a,a3447a,a3448a,a3449a,a3450a,a3451a,a3452a,a3453a,a3454a,a3455a,a3456a,a3457a,a3458a,a3459a,a3460a,a3461a,a3462a,a3463a,a3464a,a3465a,a3466a,a3467a,a3468a,a3469a,a3470a,a3471a,a3472a,a3473a,a3474a,a3475a,a3476a,a3477a,a3478a,a3479a,a3480a,a3481a,a3482a,a3483a,a3484a,a3485a,a3486a,a3487a,a3488a,a3489a,a3490a,a3491a,a3492a,a3493a,a3494a,a3495a,a3496a,a3497a,a3498a,a3499a,a3500a,a3501a,a3502a,a3503a,a3504a,a3505a,a3506a,a3507a,a3508a,a3509a,a3510a,a3511a,a3512a,a3513a,a3514a,a3515a,a3516a,a3517a,a3518a,a3519a,a3520a,a3521a,a3522a,a3523a,a3524a,a3525a,a3526a,a3527a,a3528a,a3529a,a3530a,a3531a,a3532a,a3533a,a3534a,a3535a,a3536a,a3537a,a3538a,a3539a,a3540a,a3541a,a3542a,a3543a,a3544a,a3545a,a3546a,a3547a,a3548a,a3549a,a3550a,a3551a,a3552a,a3553a,a3554a,a3555a,a3556a,a3557a,a3558a,a3559a,a3560a,a3561a,a3562a,a3563a,a3564a,a3565a,a3566a,a3567a,a3568a,a3569a,a3570a,a3571a,a3572a,a3573a,a3574a,a3575a,a3576a,a3577a,a3578a,a3579a,a3580a,a3581a,a3582a,a3583a,a3584a,a3585a,a3586a,a3587a,a3588a,a3589a,a3590a,a3591a,a3592a,a3593a,a3594a,a3595a,a3596a,a3597a,a3598a,a3599a,a3600a,a3601a,a3602a,a3603a,a3604a,a3605a,a3606a,a3607a,a3608a,a3609a,a3610a,a3611a,a3612a,a3613a,a3614a,a3615a,a3616a,a3617a,a3618a,a3619a,a3620a,a3621a,a3622a,a3623a,a3624a,a3625a,a3626a,a3627a,a3628a,a3629a,a3630a,a3631a,a3632a,a3633a,a3634a,a3635a,a3636a,a3637a,a3638a,a3639a,a3640a,a3641a,a3642a,a3643a,a3644a,a3645a,a3646a,a3647a,a3648a,a3649a,a3650a,a3651a,a3652a,a3653a,a3654a,a3655a,a3656a,a3657a,a3658a,a3659a,a3660a,a3661a,a3662a,a3663a,a3664a,a3665a,a3666a,a3667a,a3668a,a3669a,a3670a,a3671a,a3672a,a3673a,a3674a,a3675a,a3676a,a3677a,a3678a,a3679a,a3680a,a3681a,a3682a,a3683a,a3684a,a3685a,a3686a,a3687a,a3688a,a3689a,a3690a,a3691a,a3692a,a3693a,a3694a,a3695a,a3696a,a3697a,a3698a,a3699a,a3700a,a3701a,a3702a,a3703a,a3704a,a3705a,a3706a,a3707a,a3708a,a3709a,a3710a,a3711a,a3712a,a3713a,a3714a,a3715a,a3716a,a3717a,a3718a,a3719a,a3720a,a3721a,a3722a,a3723a,a3724a,a3725a,a3726a,a3727a,a3728a,a3729a,a3730a,a3731a,a3732a,a3733a,a3734a,a3735a,a3736a,a3737a,a3738a,a3739a,a3740a,a3741a,a3742a,a3743a,a3744a,a3745a,a3746a,a3747a,a3748a,a3749a,a3750a,a3751a,a3752a,a3753a,a3754a,a3755a,a3756a,a3757a,a3758a,a3759a,a3760a,a3761a,a3762a,a3763a,a3764a,a3765a,a3766a,a3767a,a3768a,a3769a,a3770a,a3771a,a3772a,a3776a,a3777a,a3780a,a3783a,a3784a,a3785a,a3789a,a3790a,a3793a,a3796a,a3797a,a3798a,a3799a,a3803a,a3804a,a3807a,a3810a,a3811a,a3812a,a3815a,a3818a,a3819a,a3822a,a3825a,a3826a,a3827a,a3828a,a3829a,a3833a,a3834a,a3837a,a3840a,a3841a,a3842a,a3846a,a3847a,a3850a,a3853a,a3854a,a3855a,a3856a,a3860a,a3861a,a3864a,a3867a,a3868a,a3869a,a3872a,a3875a,a3876a,a3879a,a3882a,a3883a,a3884a,a3885a,a3886a,a3887a,a3891a,a3892a,a3895a,a3898a,a3899a,a3900a,a3904a,a3905a,a3908a,a3911a,a3912a,a3913a,a3914a,a3918a,a3919a,a3922a,a3925a,a3926a,a3927a,a3930a,a3933a,a3934a,a3937a,a3940a,a3941a,a3942a,a3943a,a3944a,a3948a,a3949a,a3952a,a3955a,a3956a,a3957a,a3960a,a3963a,a3964a,a3967a,a3970a,a3971a,a3972a,a3973a,a3977a,a3978a,a3981a,a3984a,a3985a,a3986a,a3989a,a3992a,a3993a,a3996a,a3999a,a4000a,a4001a,a4002a,a4003a,a4004a,a4005a,a4009a,a4010a,a4013a,a4016a,a4017a,a4018a,a4022a,a4023a,a4026a,a4029a,a4030a,a4031a,a4032a,a4036a,a4037a,a4040a,a4043a,a4044a,a4045a,a4048a,a4051a,a4052a,a4055a,a4058a,a4059a,a4060a,a4061a,a4062a,a4066a,a4067a,a4070a,a4073a,a4074a,a4075a,a4078a,a4081a,a4082a,a4085a,a4088a,a4089a,a4090a,a4091a,a4095a,a4096a,a4099a,a4102a,a4103a,a4104a,a4107a,a4110a,a4111a,a4114a,a4117a,a4118a,a4119a,a4120a,a4121a,a4122a,a4126a,a4127a,a4130a,a4133a,a4134a,a4135a,a4139a,a4140a,a4143a,a4146a,a4147a,a4148a,a4149a,a4153a,a4154a,a4157a,a4160a,a4161a,a4162a,a4165a,a4168a,a4169a,a4172a,a4175a,a4176a,a4177a,a4178a,a4179a,a4183a,a4184a,a4187a,a4190a,a4191a,a4192a,a4195a,a4198a,a4199a,a4202a,a4205a,a4206a,a4207a,a4208a,a4212a,a4213a,a4216a,a4219a,a4220a,a4221a,a4224a,a4227a,a4228a,a4231a,a4234a,a4235a,a4236a,a4237a,a4238a,a4239a,a4240a,a4241a,a4245a,a4246a,a4249a,a4252a,a4253a,a4254a,a4258a,a4259a,a4262a,a4265a,a4266a,a4267a,a4268a,a4272a,a4273a,a4276a,a4279a,a4280a,a4281a,a4284a,a4287a,a4288a,a4291a,a4294a,a4295a,a4296a,a4297a,a4298a,a4302a,a4303a,a4306a,a4309a,a4310a,a4311a,a4314a,a4317a,a4318a,a4321a,a4324a,a4325a,a4326a,a4327a,a4331a,a4332a,a4335a,a4338a,a4339a,a4340a,a4343a,a4346a,a4347a,a4350a,a4353a,a4354a,a4355a,a4356a,a4357a,a4358a,a4362a,a4363a,a4366a,a4369a,a4370a,a4371a,a4375a,a4376a,a4379a,a4382a,a4383a,a4384a,a4385a,a4389a,a4390a,a4393a,a4396a,a4397a,a4398a,a4401a,a4404a,a4405a,a4408a,a4411a,a4412a,a4413a,a4414a,a4415a,a4419a,a4420a,a4423a,a4426a,a4427a,a4428a,a4431a,a4434a,a4435a,a4438a,a4441a,a4442a,a4443a,a4444a,a4448a,a4449a,a4452a,a4455a,a4456a,a4457a,a4460a,a4463a,a4464a,a4467a,a4470a,a4471a,a4472a,a4473a,a4474a,a4475a,a4476a,a4480a,a4481a,a4484a,a4487a,a4488a,a4489a,a4493a,a4494a,a4497a,a4500a,a4501a,a4502a,a4503a,a4507a,a4508a,a4511a,a4514a,a4515a,a4516a,a4519a,a4522a,a4523a,a4526a,a4529a,a4530a,a4531a,a4532a,a4533a,a4537a,a4538a,a4541a,a4544a,a4545a,a4546a,a4549a,a4552a,a4553a,a4556a,a4559a,a4560a,a4561a,a4562a,a4566a,a4567a,a4570a,a4573a,a4574a,a4575a,a4578a,a4581a,a4582a,a4585a,a4588a,a4589a,a4590a,a4591a,a4592a,a4593a,a4597a,a4598a,a4601a,a4604a,a4605a,a4606a,a4610a,a4611a,a4614a,a4617a,a4618a,a4619a,a4620a,a4624a,a4625a,a4628a,a4631a,a4632a,a4633a,a4636a,a4639a,a4640a,a4643a,a4646a,a4647a,a4648a,a4649a,a4650a,a4654a,a4655a,a4658a,a4661a,a4662a,a4663a,a4666a,a4669a,a4670a,a4673a,a4676a,a4677a,a4678a,a4679a,a4683a,a4684a,a4687a,a4690a,a4691a,a4692a,a4695a,a4698a,a4699a,a4702a,a4705a,a4706a,a4707a,a4708a,a4709a,a4710a,a4711a,a4712a,a4713a,a4717a,a4718a,a4721a,a4724a,a4725a,a4726a,a4730a,a4731a,a4734a,a4737a,a4738a,a4739a,a4740a,a4744a,a4745a,a4748a,a4751a,a4752a,a4753a,a4756a,a4759a,a4760a,a4763a,a4766a,a4767a,a4768a,a4769a,a4770a,a4774a,a4775a,a4778a,a4781a,a4782a,a4783a,a4786a,a4789a,a4790a,a4793a,a4796a,a4797a,a4798a,a4799a,a4803a,a4804a,a4807a,a4810a,a4811a,a4812a,a4815a,a4818a,a4819a,a4822a,a4825a,a4826a,a4827a,a4828a,a4829a,a4830a,a4834a,a4835a,a4838a,a4841a,a4842a,a4843a,a4847a,a4848a,a4851a,a4854a,a4855a,a4856a,a4857a,a4861a,a4862a,a4865a,a4868a,a4869a,a4870a,a4873a,a4876a,a4877a,a4880a,a4883a,a4884a,a4885a,a4886a,a4887a,a4891a,a4892a,a4895a,a4898a,a4899a,a4900a,a4903a,a4906a,a4907a,a4910a,a4913a,a4914a,a4915a,a4916a,a4920a,a4921a,a4924a,a4927a,a4928a,a4929a,a4932a,a4935a,a4936a,a4939a,a4942a,a4943a,a4944a,a4945a,a4946a,a4947a,a4948a,a4952a,a4953a,a4956a,a4959a,a4960a,a4961a,a4965a,a4966a,a4969a,a4972a,a4973a,a4974a,a4975a,a4979a,a4980a,a4983a,a4986a,a4987a,a4988a,a4991a,a4994a,a4995a,a4998a,a5001a,a5002a,a5003a,a5004a,a5005a,a5009a,a5010a,a5013a,a5016a,a5017a,a5018a,a5021a,a5024a,a5025a,a5028a,a5031a,a5032a,a5033a,a5034a,a5038a,a5039a,a5042a,a5045a,a5046a,a5047a,a5050a,a5053a,a5054a,a5057a,a5060a,a5061a,a5062a,a5063a,a5064a,a5065a,a5069a,a5070a,a5073a,a5076a,a5077a,a5078a,a5082a,a5083a,a5086a,a5089a,a5090a,a5091a,a5092a,a5096a,a5097a,a5100a,a5103a,a5104a,a5105a,a5108a,a5111a,a5112a,a5115a,a5118a,a5119a,a5120a,a5121a,a5122a,a5126a,a5127a,a5130a,a5133a,a5134a,a5135a,a5138a,a5141a,a5142a,a5145a,a5148a,a5149a,a5150a,a5151a,a5155a,a5156a,a5159a,a5162a,a5163a,a5164a,a5167a,a5170a,a5171a,a5174a,a5177a,a5178a,a5179a,a5180a,a5181a,a5182a,a5183a,a5184a,a5188a,a5189a,a5192a,a5195a,a5196a,a5197a,a5201a,a5202a,a5205a,a5208a,a5209a,a5210a,a5211a,a5215a,a5216a,a5219a,a5222a,a5223a,a5224a,a5227a,a5230a,a5231a,a5234a,a5237a,a5238a,a5239a,a5240a,a5241a,a5245a,a5246a,a5249a,a5252a,a5253a,a5254a,a5257a,a5260a,a5261a,a5264a,a5267a,a5268a,a5269a,a5270a,a5274a,a5275a,a5278a,a5281a,a5282a,a5283a,a5286a,a5289a,a5290a,a5293a,a5296a,a5297a,a5298a,a5299a,a5300a,a5301a,a5305a,a5306a,a5309a,a5312a,a5313a,a5314a,a5318a,a5319a,a5322a,a5325a,a5326a,a5327a,a5328a,a5332a,a5333a,a5336a,a5339a,a5340a,a5341a,a5344a,a5347a,a5348a,a5351a,a5354a,a5355a,a5356a,a5357a,a5358a,a5362a,a5363a,a5366a,a5369a,a5370a,a5371a,a5374a,a5377a,a5378a,a5381a,a5384a,a5385a,a5386a,a5387a,a5391a,a5392a,a5395a,a5398a,a5399a,a5400a,a5403a,a5406a,a5407a,a5410a,a5413a,a5414a,a5415a,a5416a,a5417a,a5418a,a5419a,a5423a,a5424a,a5427a,a5430a,a5431a,a5432a,a5436a,a5437a,a5440a,a5443a,a5444a,a5445a,a5446a,a5450a,a5451a,a5454a,a5457a,a5458a,a5459a,a5462a,a5465a,a5466a,a5469a,a5472a,a5473a,a5474a,a5475a,a5476a,a5480a,a5481a,a5484a,a5487a,a5488a,a5489a,a5492a,a5495a,a5496a,a5499a,a5502a,a5503a,a5504a,a5505a,a5509a,a5510a,a5513a,a5516a,a5517a,a5518a,a5521a,a5524a,a5525a,a5528a,a5531a,a5532a,a5533a,a5534a,a5535a,a5536a,a5540a,a5541a,a5544a,a5547a,a5548a,a5549a,a5553a,a5554a,a5557a,a5560a,a5561a,a5562a,a5563a,a5567a,a5568a,a5571a,a5574a,a5575a,a5576a,a5579a,a5582a,a5583a,a5586a,a5589a,a5590a,a5591a,a5592a,a5593a,a5597a,a5598a,a5601a,a5604a,a5605a,a5606a,a5609a,a5612a,a5613a,a5616a,a5619a,a5620a,a5621a,a5622a,a5626a,a5627a,a5630a,a5633a,a5634a,a5635a,a5638a,a5641a,a5642a,a5645a,a5648a,a5649a,a5650a,a5651a,a5652a,a5653a,a5654a,a5655a,a5656a,a5657a,a5661a,a5662a,a5665a,a5668a,a5669a,a5670a,a5674a,a5675a,a5678a,a5681a,a5682a,a5683a,a5684a,a5688a,a5689a,a5692a,a5695a,a5696a,a5697a,a5700a,a5703a,a5704a,a5707a,a5710a,a5711a,a5712a,a5713a,a5714a,a5718a,a5719a,a5722a,a5725a,a5726a,a5727a,a5731a,a5732a,a5735a,a5738a,a5739a,a5740a,a5741a,a5745a,a5746a,a5749a,a5752a,a5753a,a5754a,a5757a,a5760a,a5761a,a5764a,a5767a,a5768a,a5769a,a5770a,a5771a,a5772a,a5776a,a5777a,a5780a,a5783a,a5784a,a5785a,a5789a,a5790a,a5793a,a5796a,a5797a,a5798a,a5799a,a5803a,a5804a,a5807a,a5810a,a5811a,a5812a,a5815a,a5818a,a5819a,a5822a,a5825a,a5826a,a5827a,a5828a,a5829a,a5833a,a5834a,a5837a,a5840a,a5841a,a5842a,a5845a,a5848a,a5849a,a5852a,a5855a,a5856a,a5857a,a5858a,a5862a,a5863a,a5866a,a5869a,a5870a,a5871a,a5874a,a5877a,a5878a,a5881a,a5884a,a5885a,a5886a,a5887a,a5888a,a5889a,a5890a,a5894a,a5895a,a5898a,a5901a,a5902a,a5903a,a5907a,a5908a,a5911a,a5914a,a5915a,a5916a,a5917a,a5921a,a5922a,a5925a,a5928a,a5929a,a5930a,a5933a,a5936a,a5937a,a5940a,a5943a,a5944a,a5945a,a5946a,a5947a,a5951a,a5952a,a5955a,a5958a,a5959a,a5960a,a5963a,a5966a,a5967a,a5970a,a5973a,a5974a,a5975a,a5976a,a5980a,a5981a,a5984a,a5987a,a5988a,a5989a,a5992a,a5995a,a5996a,a5999a,a6002a,a6003a,a6004a,a6005a,a6006a,a6007a,a6011a,a6012a,a6015a,a6018a,a6019a,a6020a,a6024a,a6025a,a6028a,a6031a,a6032a,a6033a,a6034a,a6038a,a6039a,a6042a,a6045a,a6046a,a6047a,a6050a,a6053a,a6054a,a6057a,a6060a,a6061a,a6062a,a6063a,a6064a,a6068a,a6069a,a6072a,a6075a,a6076a,a6077a,a6080a,a6083a,a6084a,a6087a,a6090a,a6091a,a6092a,a6093a,a6097a,a6098a,a6101a,a6104a,a6105a,a6106a,a6109a,a6112a,a6113a,a6116a,a6119a,a6120a,a6121a,a6122a,a6123a,a6124a,a6125a,a6126a,a6130a,a6131a,a6134a,a6137a,a6138a,a6139a,a6143a,a6144a,a6147a,a6150a,a6151a,a6152a,a6153a,a6157a,a6158a,a6161a,a6164a,a6165a,a6166a,a6169a,a6172a,a6173a,a6176a,a6179a,a6180a,a6181a,a6182a,a6183a,a6187a,a6188a,a6191a,a6194a,a6195a,a6196a,a6199a,a6202a,a6203a,a6206a,a6209a,a6210a,a6211a,a6212a,a6216a,a6217a,a6220a,a6223a,a6224a,a6225a,a6228a,a6231a,a6232a,a6235a,a6238a,a6239a,a6240a,a6241a,a6242a,a6243a,a6247a,a6248a,a6251a,a6254a,a6255a,a6256a,a6260a,a6261a,a6264a,a6267a,a6268a,a6269a,a6270a,a6274a,a6275a,a6278a,a6281a,a6282a,a6283a,a6286a,a6289a,a6290a,a6293a,a6296a,a6297a,a6298a,a6299a,a6300a,a6304a,a6305a,a6308a,a6311a,a6312a,a6313a,a6316a,a6319a,a6320a,a6323a,a6326a,a6327a,a6328a,a6329a,a6333a,a6334a,a6337a,a6340a,a6341a,a6342a,a6345a,a6348a,a6349a,a6352a,a6355a,a6356a,a6357a,a6358a,a6359a,a6360a,a6361a,a6365a,a6366a,a6369a,a6372a,a6373a,a6374a,a6378a,a6379a,a6382a,a6385a,a6386a,a6387a,a6388a,a6392a,a6393a,a6396a,a6399a,a6400a,a6401a,a6404a,a6407a,a6408a,a6411a,a6414a,a6415a,a6416a,a6417a,a6418a,a6422a,a6423a,a6426a,a6429a,a6430a,a6431a,a6434a,a6437a,a6438a,a6441a,a6444a,a6445a,a6446a,a6447a,a6451a,a6452a,a6455a,a6458a,a6459a,a6460a,a6463a,a6466a,a6467a,a6470a,a6473a,a6474a,a6475a,a6476a,a6477a,a6478a,a6482a,a6483a,a6486a,a6489a,a6490a,a6491a,a6495a,a6496a,a6499a,a6502a,a6503a,a6504a,a6505a,a6509a,a6510a,a6513a,a6516a,a6517a,a6518a,a6521a,a6524a,a6525a,a6528a,a6531a,a6532a,a6533a,a6534a,a6535a,a6539a,a6540a,a6543a,a6546a,a6547a,a6548a,a6551a,a6554a,a6555a,a6558a,a6561a,a6562a,a6563a,a6564a,a6568a,a6569a,a6572a,a6575a,a6576a,a6577a,a6580a,a6583a,a6584a,a6587a,a6590a,a6591a,a6592a,a6593a,a6594a,a6595a,a6596a,a6597a,a6598a,a6602a,a6603a,a6606a,a6609a,a6610a,a6611a,a6615a,a6616a,a6619a,a6622a,a6623a,a6624a,a6625a,a6629a,a6630a,a6633a,a6636a,a6637a,a6638a,a6641a,a6644a,a6645a,a6648a,a6651a,a6652a,a6653a,a6654a,a6655a,a6659a,a6660a,a6663a,a6666a,a6667a,a6668a,a6671a,a6674a,a6675a,a6678a,a6681a,a6682a,a6683a,a6684a,a6688a,a6689a,a6692a,a6695a,a6696a,a6697a,a6700a,a6703a,a6704a,a6707a,a6710a,a6711a,a6712a,a6713a,a6714a,a6715a,a6719a,a6720a,a6723a,a6726a,a6727a,a6728a,a6732a,a6733a,a6736a,a6739a,a6740a,a6741a,a6742a,a6746a,a6747a,a6750a,a6753a,a6754a,a6755a,a6758a,a6761a,a6762a,a6765a,a6768a,a6769a,a6770a,a6771a,a6772a,a6776a,a6777a,a6780a,a6783a,a6784a,a6785a,a6788a,a6791a,a6792a,a6795a,a6798a,a6799a,a6800a,a6801a,a6805a,a6806a,a6809a,a6812a,a6813a,a6814a,a6817a,a6820a,a6821a,a6824a,a6827a,a6828a,a6829a,a6830a,a6831a,a6832a,a6833a,a6837a,a6838a,a6841a,a6844a,a6845a,a6846a,a6850a,a6851a,a6854a,a6857a,a6858a,a6859a,a6860a,a6864a,a6865a,a6868a,a6871a,a6872a,a6873a,a6876a,a6879a,a6880a,a6883a,a6886a,a6887a,a6888a,a6889a,a6890a,a6894a,a6895a,a6898a,a6901a,a6902a,a6903a,a6906a,a6909a,a6910a,a6913a,a6916a,a6917a,a6918a,a6919a,a6923a,a6924a,a6927a,a6930a,a6931a,a6932a,a6935a,a6938a,a6939a,a6942a,a6945a,a6946a,a6947a,a6948a,a6949a,a6950a,a6954a,a6955a,a6958a,a6961a,a6962a,a6963a,a6967a,a6968a,a6971a,a6974a,a6975a,a6976a,a6977a,a6981a,a6982a,a6985a,a6988a,a6989a,a6990a,a6993a,a6996a,a6997a,a7000a,a7003a,a7004a,a7005a,a7006a,a7007a,a7011a,a7012a,a7015a,a7018a,a7019a,a7020a,a7023a,a7026a,a7027a,a7030a,a7033a,a7034a,a7035a,a7036a,a7040a,a7041a,a7044a,a7047a,a7048a,a7049a,a7052a,a7055a,a7056a,a7059a,a7062a,a7063a,a7064a,a7065a,a7066a,a7067a,a7068a,a7069a,a7073a,a7074a,a7077a,a7080a,a7081a,a7082a,a7086a,a7087a,a7090a,a7093a,a7094a,a7095a,a7096a,a7100a,a7101a,a7104a,a7107a,a7108a,a7109a,a7112a,a7115a,a7116a,a7119a,a7122a,a7123a,a7124a,a7125a,a7126a,a7130a,a7131a,a7134a,a7137a,a7138a,a7139a,a7142a,a7145a,a7146a,a7149a,a7152a,a7153a,a7154a,a7155a,a7159a,a7160a,a7163a,a7166a,a7167a,a7168a,a7171a,a7174a,a7175a,a7178a,a7181a,a7182a,a7183a,a7184a,a7185a,a7186a,a7190a,a7191a,a7194a,a7197a,a7198a,a7199a,a7203a,a7204a,a7207a,a7210a,a7211a,a7212a,a7213a,a7217a,a7218a,a7221a,a7224a,a7225a,a7226a,a7229a,a7232a,a7233a,a7236a,a7239a,a7240a,a7241a,a7242a,a7243a,a7247a,a7248a,a7251a,a7254a,a7255a,a7256a,a7259a,a7262a,a7263a,a7266a,a7269a,a7270a,a7271a,a7272a,a7276a,a7277a,a7280a,a7283a,a7284a,a7285a,a7288a,a7291a,a7292a,a7295a,a7298a,a7299a,a7300a,a7301a,a7302a,a7303a,a7304a,a7308a,a7309a,a7312a,a7315a,a7316a,a7317a,a7321a,a7322a,a7325a,a7328a,a7329a,a7330a,a7331a,a7335a,a7336a,a7339a,a7342a,a7343a,a7344a,a7347a,a7350a,a7351a,a7354a,a7357a,a7358a,a7359a,a7360a,a7361a,a7365a,a7366a,a7369a,a7372a,a7373a,a7374a,a7377a,a7380a,a7381a,a7384a,a7387a,a7388a,a7389a,a7390a,a7394a,a7395a,a7398a,a7401a,a7402a,a7403a,a7406a,a7409a,a7410a,a7413a,a7416a,a7417a,a7418a,a7419a,a7420a,a7421a,a7425a,a7426a,a7429a,a7432a,a7433a,a7434a,a7438a,a7439a,a7442a,a7445a,a7446a,a7447a,a7448a,a7452a,a7453a,a7456a,a7459a,a7460a,a7461a,a7464a,a7467a,a7468a,a7471a,a7474a,a7475a,a7476a,a7477a,a7478a,a7482a,a7483a,a7486a,a7489a,a7490a,a7491a,a7494a,a7497a,a7498a,a7501a,a7504a,a7505a,a7506a,a7507a,a7511a,a7512a,a7515a,a7518a,a7519a,a7520a,a7523a,a7526a,a7527a,a7530a,a7533a,a7534a,a7535a,a7536a,a7537a,a7538a,a7539a,a7540a,a7541a,a7542a,a7543a,a7547a,a7548a,a7551a,a7554a,a7555a,a7556a,a7560a,a7561a,a7564a,a7567a,a7568a,a7569a,a7570a,a7574a,a7575a,a7578a,a7581a,a7582a,a7583a,a7586a,a7589a,a7590a,a7593a,a7596a,a7597a,a7598a,a7599a,a7600a,a7604a,a7605a,a7608a,a7611a,a7612a,a7613a,a7617a,a7618a,a7621a,a7624a,a7625a,a7626a,a7627a,a7631a,a7632a,a7635a,a7638a,a7639a,a7640a,a7643a,a7646a,a7647a,a7650a,a7653a,a7654a,a7655a,a7656a,a7657a,a7658a,a7662a,a7663a,a7666a,a7669a,a7670a,a7671a,a7675a,a7676a,a7679a,a7682a,a7683a,a7684a,a7685a,a7689a,a7690a,a7693a,a7696a,a7697a,a7698a,a7701a,a7704a,a7705a,a7708a,a7711a,a7712a,a7713a,a7714a,a7715a,a7719a,a7720a,a7723a,a7726a,a7727a,a7728a,a7731a,a7734a,a7735a,a7738a,a7741a,a7742a,a7743a,a7744a,a7748a,a7749a,a7752a,a7755a,a7756a,a7757a,a7760a,a7763a,a7764a,a7767a,a7770a,a7771a,a7772a,a7773a,a7774a,a7775a,a7776a,a7780a,a7781a,a7784a,a7787a,a7788a,a7789a,a7793a,a7794a,a7797a,a7800a,a7801a,a7802a,a7803a,a7807a,a7808a,a7811a,a7814a,a7815a,a7816a,a7819a,a7822a,a7823a,a7826a,a7829a,a7830a,a7831a,a7832a,a7833a,a7837a,a7838a,a7841a,a7844a,a7845a,a7846a,a7849a,a7852a,a7853a,a7856a,a7859a,a7860a,a7861a,a7862a,a7866a,a7867a,a7870a,a7873a,a7874a,a7875a,a7878a,a7881a,a7882a,a7885a,a7888a,a7889a,a7890a,a7891a,a7892a,a7893a,a7897a,a7898a,a7901a,a7904a,a7905a,a7906a,a7910a,a7911a,a7914a,a7917a,a7918a,a7919a,a7920a,a7924a,a7925a,a7928a,a7931a,a7932a,a7933a,a7936a,a7939a,a7940a,a7943a,a7946a,a7947a,a7948a,a7949a,a7950a,a7954a,a7955a,a7958a,a7961a,a7962a,a7963a,a7966a,a7969a,a7970a,a7973a,a7976a,a7977a,a7978a,a7979a,a7983a,a7984a,a7987a,a7990a,a7991a,a7992a,a7995a,a7998a,a7999a,a8002a,a8005a,a8006a,a8007a,a8008a,a8009a,a8010a,a8011a,a8012a,a8016a,a8017a,a8020a,a8023a,a8024a,a8025a,a8029a,a8030a,a8033a,a8036a,a8037a,a8038a,a8039a,a8043a,a8044a,a8047a,a8050a,a8051a,a8052a,a8055a,a8058a,a8059a,a8062a,a8065a,a8066a,a8067a,a8068a,a8069a,a8073a,a8074a,a8077a,a8080a,a8081a,a8082a,a8085a,a8088a,a8089a,a8092a,a8095a,a8096a,a8097a,a8098a,a8102a,a8103a,a8106a,a8109a,a8110a,a8111a,a8114a,a8117a,a8118a,a8121a,a8124a,a8125a,a8126a,a8127a,a8128a,a8129a,a8133a,a8134a,a8137a,a8140a,a8141a,a8142a,a8146a,a8147a,a8150a,a8153a,a8154a,a8155a,a8156a,a8160a,a8161a,a8164a,a8167a,a8168a,a8169a,a8172a,a8175a,a8176a,a8179a,a8182a,a8183a,a8184a,a8185a,a8186a,a8190a,a8191a,a8194a,a8197a,a8198a,a8199a,a8202a,a8205a,a8206a,a8209a,a8212a,a8213a,a8214a,a8215a,a8219a,a8220a,a8223a,a8226a,a8227a,a8228a,a8231a,a8234a,a8235a,a8238a,a8241a,a8242a,a8243a,a8244a,a8245a,a8246a,a8247a,a8251a,a8252a,a8255a,a8258a,a8259a,a8260a,a8264a,a8265a,a8268a,a8271a,a8272a,a8273a,a8274a,a8278a,a8279a,a8282a,a8285a,a8286a,a8287a,a8290a,a8293a,a8294a,a8297a,a8300a,a8301a,a8302a,a8303a,a8304a,a8308a,a8309a,a8312a,a8315a,a8316a,a8317a,a8320a,a8323a,a8324a,a8327a,a8330a,a8331a,a8332a,a8333a,a8337a,a8338a,a8341a,a8344a,a8345a,a8346a,a8349a,a8352a,a8353a,a8356a,a8359a,a8360a,a8361a,a8362a,a8363a,a8364a,a8368a,a8369a,a8372a,a8375a,a8376a,a8377a,a8381a,a8382a,a8385a,a8388a,a8389a,a8390a,a8391a,a8395a,a8396a,a8399a,a8402a,a8403a,a8404a,a8407a,a8410a,a8411a,a8414a,a8417a,a8418a,a8419a,a8420a,a8421a,a8425a,a8426a,a8429a,a8432a,a8433a,a8434a,a8437a,a8440a,a8441a,a8444a,a8447a,a8448a,a8449a,a8450a,a8454a,a8455a,a8458a,a8461a,a8462a,a8463a,a8466a,a8469a,a8470a,a8473a,a8476a,a8477a,a8478a,a8479a,a8480a,a8481a,a8482a,a8483a,a8484a,a8488a,a8489a,a8492a,a8495a,a8496a,a8497a,a8501a,a8502a,a8505a,a8508a,a8509a,a8510a,a8511a,a8515a,a8516a,a8519a,a8522a,a8523a,a8524a,a8527a,a8530a,a8531a,a8534a,a8537a,a8538a,a8539a,a8540a,a8541a,a8545a,a8546a,a8549a,a8552a,a8553a,a8554a,a8557a,a8560a,a8561a,a8564a,a8567a,a8568a,a8569a,a8570a,a8574a,a8575a,a8578a,a8581a,a8582a,a8583a,a8586a,a8589a,a8590a,a8593a,a8596a,a8597a,a8598a,a8599a,a8600a,a8601a,a8605a,a8606a,a8609a,a8612a,a8613a,a8614a,a8618a,a8619a,a8622a,a8625a,a8626a,a8627a,a8628a,a8632a,a8633a,a8636a,a8639a,a8640a,a8641a,a8644a,a8647a,a8648a,a8651a,a8654a,a8655a,a8656a,a8657a,a8658a,a8662a,a8663a,a8666a,a8669a,a8670a,a8671a,a8674a,a8677a,a8678a,a8681a,a8684a,a8685a,a8686a,a8687a,a8691a,a8692a,a8695a,a8698a,a8699a,a8700a,a8703a,a8706a,a8707a,a8710a,a8713a,a8714a,a8715a,a8716a,a8717a,a8718a,a8719a,a8723a,a8724a,a8727a,a8730a,a8731a,a8732a,a8736a,a8737a,a8740a,a8743a,a8744a,a8745a,a8746a,a8750a,a8751a,a8754a,a8757a,a8758a,a8759a,a8762a,a8765a,a8766a,a8769a,a8772a,a8773a,a8774a,a8775a,a8776a,a8780a,a8781a,a8784a,a8787a,a8788a,a8789a,a8792a,a8795a,a8796a,a8799a,a8802a,a8803a,a8804a,a8805a,a8809a,a8810a,a8813a,a8816a,a8817a,a8818a,a8821a,a8824a,a8825a,a8828a,a8831a,a8832a,a8833a,a8834a,a8835a,a8836a,a8840a,a8841a,a8844a,a8847a,a8848a,a8849a,a8853a,a8854a,a8857a,a8860a,a8861a,a8862a,a8863a,a8867a,a8868a,a8871a,a8874a,a8875a,a8876a,a8879a,a8882a,a8883a,a8886a,a8889a,a8890a,a8891a,a8892a,a8893a,a8897a,a8898a,a8901a,a8904a,a8905a,a8906a,a8909a,a8912a,a8913a,a8916a,a8919a,a8920a,a8921a,a8922a,a8926a,a8927a,a8930a,a8933a,a8934a,a8935a,a8938a,a8941a,a8942a,a8945a,a8948a,a8949a,a8950a,a8951a,a8952a,a8953a,a8954a,a8955a,a8959a,a8960a,a8963a,a8966a,a8967a,a8968a,a8972a,a8973a,a8976a,a8979a,a8980a,a8981a,a8982a,a8986a,a8987a,a8990a,a8993a,a8994a,a8995a,a8998a,a9001a,a9002a,a9005a,a9008a,a9009a,a9010a,a9011a,a9012a,a9016a,a9017a,a9020a,a9023a,a9024a,a9025a,a9028a,a9031a,a9032a,a9035a,a9038a,a9039a,a9040a,a9041a,a9045a,a9046a,a9049a,a9052a,a9053a,a9054a,a9057a,a9060a,a9061a,a9064a,a9067a,a9068a,a9069a,a9070a,a9071a,a9072a,a9076a,a9077a,a9080a,a9083a,a9084a,a9085a,a9089a,a9090a,a9093a,a9096a,a9097a,a9098a,a9099a,a9103a,a9104a,a9107a,a9110a,a9111a,a9112a,a9115a,a9118a,a9119a,a9122a,a9125a,a9126a,a9127a,a9128a,a9129a,a9133a,a9134a,a9137a,a9140a,a9141a,a9142a,a9145a,a9148a,a9149a,a9152a,a9155a,a9156a,a9157a,a9158a,a9162a,a9163a,a9166a,a9169a,a9170a,a9171a,a9174a,a9177a,a9178a,a9181a,a9184a,a9185a,a9186a,a9187a,a9188a,a9189a,a9190a,a9194a,a9195a,a9198a,a9201a,a9202a,a9203a,a9207a,a9208a,a9211a,a9214a,a9215a,a9216a,a9217a,a9221a,a9222a,a9225a,a9228a,a9229a,a9230a,a9233a,a9236a,a9237a,a9240a,a9243a,a9244a,a9245a,a9246a,a9247a,a9251a,a9252a,a9255a,a9258a,a9259a,a9260a,a9263a,a9266a,a9267a,a9270a,a9273a,a9274a,a9275a,a9276a,a9280a,a9281a,a9284a,a9287a,a9288a,a9289a,a9292a,a9295a,a9296a,a9299a,a9302a,a9303a,a9304a,a9305a,a9306a,a9307a,a9311a,a9312a,a9315a,a9318a,a9319a,a9320a,a9324a,a9325a,a9328a,a9331a,a9332a,a9333a,a9334a,a9338a,a9339a,a9342a,a9345a,a9346a,a9347a,a9350a,a9353a,a9354a,a9357a,a9360a,a9361a,a9362a,a9363a,a9364a,a9368a,a9369a,a9372a,a9375a,a9376a,a9377a,a9380a,a9383a,a9384a,a9387a,a9390a,a9391a,a9392a,a9393a,a9397a,a9398a,a9401a,a9404a,a9405a,a9406a,a9409a,a9412a,a9413a,a9416a,a9419a,a9420a,a9421a,a9422a,a9423a,a9424a,a9425a,a9426a,a9427a,a9428a,a9432a,a9433a,a9436a,a9439a,a9440a,a9441a,a9445a,a9446a,a9449a,a9452a,a9453a,a9454a,a9455a,a9459a,a9460a,a9463a,a9466a,a9467a,a9468a,a9471a,a9474a,a9475a,a9478a,a9481a,a9482a,a9483a,a9484a,a9485a,a9489a,a9490a,a9493a,a9496a,a9497a,a9498a,a9502a,a9503a,a9506a,a9509a,a9510a,a9511a,a9512a,a9516a,a9517a,a9520a,a9523a,a9524a,a9525a,a9528a,a9531a,a9532a,a9535a,a9538a,a9539a,a9540a,a9541a,a9542a,a9543a,a9547a,a9548a,a9551a,a9554a,a9555a,a9556a,a9560a,a9561a,a9564a,a9567a,a9568a,a9569a,a9570a,a9574a,a9575a,a9578a,a9581a,a9582a,a9583a,a9586a,a9589a,a9590a,a9593a,a9596a,a9597a,a9598a,a9599a,a9600a,a9604a,a9605a,a9608a,a9611a,a9612a,a9613a,a9616a,a9619a,a9620a,a9623a,a9626a,a9627a,a9628a,a9629a,a9633a,a9634a,a9637a,a9640a,a9641a,a9642a,a9645a,a9648a,a9649a,a9652a,a9655a,a9656a,a9657a,a9658a,a9659a,a9660a,a9661a,a9665a,a9666a,a9669a,a9672a,a9673a,a9674a,a9678a,a9679a,a9682a,a9685a,a9686a,a9687a,a9688a,a9692a,a9693a,a9696a,a9699a,a9700a,a9701a,a9704a,a9707a,a9708a,a9711a,a9714a,a9715a,a9716a,a9717a,a9718a,a9722a,a9723a,a9726a,a9729a,a9730a,a9731a,a9734a,a9737a,a9738a,a9741a,a9744a,a9745a,a9746a,a9747a,a9751a,a9752a,a9755a,a9758a,a9759a,a9760a,a9763a,a9766a,a9767a,a9770a,a9773a,a9774a,a9775a,a9776a,a9777a,a9778a,a9782a,a9783a,a9786a,a9789a,a9790a,a9791a,a9795a,a9796a,a9799a,a9802a,a9803a,a9804a,a9805a,a9809a,a9810a,a9813a,a9816a,a9817a,a9818a,a9821a,a9824a,a9825a,a9828a,a9831a,a9832a,a9833a,a9834a,a9835a,a9839a,a9840a,a9843a,a9846a,a9847a,a9848a,a9851a,a9854a,a9855a,a9858a,a9861a,a9862a,a9863a,a9864a,a9868a,a9869a,a9872a,a9875a,a9876a,a9877a,a9880a,a9883a,a9884a,a9887a,a9890a,a9891a,a9892a,a9893a,a9894a,a9895a,a9896a,a9897a,a9901a,a9902a,a9905a,a9908a,a9909a,a9910a,a9914a,a9915a,a9918a,a9921a,a9922a,a9923a,a9924a,a9928a,a9929a,a9932a,a9935a,a9936a,a9937a,a9940a,a9943a,a9944a,a9947a,a9950a,a9951a,a9952a,a9953a,a9954a,a9958a,a9959a,a9962a,a9965a,a9966a,a9967a,a9970a,a9973a,a9974a,a9977a,a9980a,a9981a,a9982a,a9983a,a9987a,a9988a,a9991a,a9994a,a9995a,a9996a,a9999a,a10002a,a10003a,a10006a,a10009a,a10010a,a10011a,a10012a,a10013a,a10014a,a10018a,a10019a,a10022a,a10025a,a10026a,a10027a,a10031a,a10032a,a10035a,a10038a,a10039a,a10040a,a10041a,a10045a,a10046a,a10049a,a10052a,a10053a,a10054a,a10057a,a10060a,a10061a,a10064a,a10067a,a10068a,a10069a,a10070a,a10071a,a10075a,a10076a,a10079a,a10082a,a10083a,a10084a,a10087a,a10090a,a10091a,a10094a,a10097a,a10098a,a10099a,a10100a,a10104a,a10105a,a10108a,a10111a,a10112a,a10113a,a10116a,a10119a,a10120a,a10123a,a10126a,a10127a,a10128a,a10129a,a10130a,a10131a,a10132a,a10136a,a10137a,a10140a,a10143a,a10144a,a10145a,a10149a,a10150a,a10153a,a10156a,a10157a,a10158a,a10159a,a10163a,a10164a,a10167a,a10170a,a10171a,a10172a,a10175a,a10178a,a10179a,a10182a,a10185a,a10186a,a10187a,a10188a,a10189a,a10193a,a10194a,a10197a,a10200a,a10201a,a10202a,a10205a,a10208a,a10209a,a10212a,a10215a,a10216a,a10217a,a10218a,a10222a,a10223a,a10226a,a10229a,a10230a,a10231a,a10234a,a10237a,a10238a,a10241a,a10244a,a10245a,a10246a,a10247a,a10248a,a10249a,a10253a,a10254a,a10257a,a10260a,a10261a,a10262a,a10266a,a10267a,a10270a,a10273a,a10274a,a10275a,a10276a,a10280a,a10281a,a10284a,a10287a,a10288a,a10289a,a10292a,a10295a,a10296a,a10299a,a10302a,a10303a,a10304a,a10305a,a10306a,a10310a,a10311a,a10314a,a10317a,a10318a,a10319a,a10322a,a10325a,a10326a,a10329a,a10332a,a10333a,a10334a,a10335a,a10339a,a10340a,a10343a,a10346a,a10347a,a10348a,a10351a,a10354a,a10355a,a10358a,a10361a,a10362a,a10363a,a10364a,a10365a,a10366a,a10367a,a10368a,a10369a,a10373a,a10374a,a10377a,a10380a,a10381a,a10382a,a10386a,a10387a,a10390a,a10393a,a10394a,a10395a,a10396a,a10400a,a10401a,a10404a,a10407a,a10408a,a10409a,a10412a,a10415a,a10416a,a10419a,a10422a,a10423a,a10424a,a10425a,a10426a,a10430a,a10431a,a10434a,a10437a,a10438a,a10439a,a10442a,a10445a,a10446a,a10449a,a10452a,a10453a,a10454a,a10455a,a10459a,a10460a,a10463a,a10466a,a10467a,a10468a,a10471a,a10474a,a10475a,a10478a,a10481a,a10482a,a10483a,a10484a,a10485a,a10486a,a10490a,a10491a,a10494a,a10497a,a10498a,a10499a,a10503a,a10504a,a10507a,a10510a,a10511a,a10512a,a10513a,a10517a,a10518a,a10521a,a10524a,a10525a,a10526a,a10529a,a10532a,a10533a,a10536a,a10539a,a10540a,a10541a,a10542a,a10543a,a10547a,a10548a,a10551a,a10554a,a10555a,a10556a,a10559a,a10562a,a10563a,a10566a,a10569a,a10570a,a10571a,a10572a,a10576a,a10577a,a10580a,a10583a,a10584a,a10585a,a10588a,a10591a,a10592a,a10595a,a10598a,a10599a,a10600a,a10601a,a10602a,a10603a,a10604a,a10608a,a10609a,a10612a,a10615a,a10616a,a10617a,a10621a,a10622a,a10625a,a10628a,a10629a,a10630a,a10631a,a10635a,a10636a,a10639a,a10642a,a10643a,a10644a,a10647a,a10650a,a10651a,a10654a,a10657a,a10658a,a10659a,a10660a,a10661a,a10665a,a10666a,a10669a,a10672a,a10673a,a10674a,a10677a,a10680a,a10681a,a10684a,a10687a,a10688a,a10689a,a10690a,a10694a,a10695a,a10698a,a10701a,a10702a,a10703a,a10706a,a10709a,a10710a,a10713a,a10716a,a10717a,a10718a,a10719a,a10720a,a10721a,a10725a,a10726a,a10729a,a10732a,a10733a,a10734a,a10738a,a10739a,a10742a,a10745a,a10746a,a10747a,a10748a,a10752a,a10753a,a10756a,a10759a,a10760a,a10761a,a10764a,a10767a,a10768a,a10771a,a10774a,a10775a,a10776a,a10777a,a10778a,a10782a,a10783a,a10786a,a10789a,a10790a,a10791a,a10794a,a10797a,a10798a,a10801a,a10804a,a10805a,a10806a,a10807a,a10811a,a10812a,a10815a,a10818a,a10819a,a10820a,a10823a,a10826a,a10827a,a10830a,a10833a,a10834a,a10835a,a10836a,a10837a,a10838a,a10839a,a10840a,a10844a,a10845a,a10848a,a10851a,a10852a,a10853a,a10857a,a10858a,a10861a,a10864a,a10865a,a10866a,a10867a,a10871a,a10872a,a10875a,a10878a,a10879a,a10880a,a10883a,a10886a,a10887a,a10890a,a10893a,a10894a,a10895a,a10896a,a10897a,a10901a,a10902a,a10905a,a10908a,a10909a,a10910a,a10913a,a10916a,a10917a,a10920a,a10923a,a10924a,a10925a,a10926a,a10930a,a10931a,a10934a,a10937a,a10938a,a10939a,a10942a,a10945a,a10946a,a10949a,a10952a,a10953a,a10954a,a10955a,a10956a,a10957a,a10961a,a10962a,a10965a,a10968a,a10969a,a10970a,a10974a,a10975a,a10978a,a10981a,a10982a,a10983a,a10984a,a10988a,a10989a,a10992a,a10995a,a10996a,a10997a,a11000a,a11003a,a11004a,a11007a,a11010a,a11011a,a11012a,a11013a,a11014a,a11018a,a11019a,a11022a,a11025a,a11026a,a11027a,a11030a,a11033a,a11034a,a11037a,a11040a,a11041a,a11042a,a11043a,a11047a,a11048a,a11051a,a11054a,a11055a,a11056a,a11059a,a11062a,a11063a,a11066a,a11069a,a11070a,a11071a,a11072a,a11073a,a11074a,a11075a,a11079a,a11080a,a11083a,a11086a,a11087a,a11088a,a11092a,a11093a,a11096a,a11099a,a11100a,a11101a,a11102a,a11106a,a11107a,a11110a,a11113a,a11114a,a11115a,a11118a,a11121a,a11122a,a11125a,a11128a,a11129a,a11130a,a11131a,a11132a,a11136a,a11137a,a11140a,a11143a,a11144a,a11145a,a11148a,a11151a,a11152a,a11155a,a11158a,a11159a,a11160a,a11161a,a11165a,a11166a,a11169a,a11172a,a11173a,a11174a,a11177a,a11180a,a11181a,a11184a,a11187a,a11188a,a11189a,a11190a,a11191a,a11192a,a11196a,a11197a,a11200a,a11203a,a11204a,a11205a,a11209a,a11210a,a11213a,a11216a,a11217a,a11218a,a11219a,a11223a,a11224a,a11227a,a11230a,a11231a,a11232a,a11235a,a11238a,a11239a,a11242a,a11245a,a11246a,a11247a,a11248a,a11249a,a11253a,a11254a,a11257a,a11260a,a11261a,a11262a,a11265a,a11268a,a11269a,a11272a,a11275a,a11276a,a11277a,a11278a,a11282a,a11283a,a11286a,a11289a,a11290a,a11291a,a11294a,a11297a,a11298a,a11301a,a11304a,a11305a,a11306a,a11307a,a11308a,a11309a,a11310a,a11311a,a11312a,a11313a,a11314a,a11317a,a11320a,a11321a,a11324a,a11327a,a11328a,a11331a,a11334a,a11335a,a11338a,a11341a,a11342a,a11345a,a11348a,a11349a,a11352a,a11355a,a11356a,a11359a,a11362a,a11363a,a11366a,a11369a,a11370a,a11373a,a11376a,a11377a,a11380a,a11383a,a11384a,a11387a,a11390a,a11391a,a11394a,a11397a,a11398a,a11401a,a11404a,a11405a,a11408a,a11411a,a11412a,a11415a,a11418a,a11419a,a11422a,a11425a,a11426a,a11429a,a11432a,a11433a,a11436a,a11439a,a11440a,a11443a,a11446a,a11447a,a11450a,a11453a,a11454a,a11457a,a11460a,a11461a,a11464a,a11467a,a11468a,a11471a,a11474a,a11475a,a11478a,a11481a,a11482a,a11485a,a11488a,a11489a,a11492a,a11496a,a11497a,a11498a,a11501a,a11504a,a11505a,a11508a,a11512a,a11513a,a11514a,a11517a,a11520a,a11521a,a11524a,a11528a,a11529a,a11530a,a11533a,a11536a,a11537a,a11540a,a11544a,a11545a,a11546a,a11549a,a11552a,a11553a,a11556a,a11560a,a11561a,a11562a,a11565a,a11568a,a11569a,a11572a,a11576a,a11577a,a11578a,a11581a,a11584a,a11585a,a11588a,a11592a,a11593a,a11594a,a11597a,a11600a,a11601a,a11604a,a11608a,a11609a,a11610a,a11613a,a11617a,a11618a,a11619a,a11622a,a11626a,a11627a,a11628a,a11631a,a11635a,a11636a,a11637a,a11640a,a11644a,a11645a,a11646a,a11649a,a11653a,a11654a,a11655a,a11658a,a11662a,a11663a,a11664a,a11667a,a11671a,a11672a,a11673a,a11676a,a11680a,a11681a,a11682a,a11685a,a11689a,a11690a,a11691a,a11694a,a11698a,a11699a,a11700a,a11703a,a11707a,a11708a,a11709a,a11712a,a11716a,a11717a,a11718a,a11721a,a11725a,a11726a,a11727a,a11730a,a11734a,a11735a,a11736a,a11739a,a11743a,a11744a,a11745a,a11748a,a11752a,a11753a,a11754a,a11757a,a11761a,a11762a,a11763a,a11766a,a11770a,a11771a,a11772a,a11775a,a11779a,a11780a,a11781a,a11784a,a11788a,a11789a,a11790a,a11793a,a11797a,a11798a,a11799a,a11802a,a11806a,a11807a,a11808a,a11811a,a11815a,a11816a,a11817a,a11820a,a11824a,a11825a,a11826a,a11829a,a11833a,a11834a,a11835a,a11838a,a11842a,a11843a,a11844a,a11847a,a11851a,a11852a,a11853a,a11856a,a11860a,a11861a,a11862a,a11865a,a11869a,a11870a,a11871a,a11874a,a11878a,a11879a,a11880a,a11883a,a11887a,a11888a,a11889a,a11892a,a11896a,a11897a,a11898a,a11901a,a11905a,a11906a,a11907a,a11910a,a11914a,a11915a,a11916a,a11919a,a11923a,a11924a,a11925a,a11928a,a11932a,a11933a,a11934a,a11937a,a11941a,a11942a,a11943a,a11946a,a11950a,a11951a,a11952a,a11955a,a11959a,a11960a,a11961a,a11964a,a11968a,a11969a,a11970a,a11973a,a11977a,a11978a,a11979a,a11982a,a11986a,a11987a,a11988a,a11991a,a11995a,a11996a,a11997a,a12000a,a12004a,a12005a,a12006a,a12009a,a12013a,a12014a,a12015a,a12018a,a12022a,a12023a,a12024a,a12027a,a12031a,a12032a,a12033a,a12036a,a12040a,a12041a,a12042a,a12045a,a12049a,a12050a,a12051a,a12054a,a12058a,a12059a,a12060a,a12063a,a12067a,a12068a,a12069a,a12072a,a12076a,a12077a,a12078a,a12081a,a12085a,a12086a,a12087a,a12090a,a12094a,a12095a,a12096a,a12099a,a12103a,a12104a,a12105a,a12108a,a12112a,a12113a,a12114a,a12117a,a12121a,a12122a,a12123a,a12126a,a12130a,a12131a,a12132a,a12135a,a12139a,a12140a,a12141a,a12144a,a12148a,a12149a,a12150a,a12153a,a12157a,a12158a,a12159a,a12162a,a12166a,a12167a,a12168a,a12171a,a12175a,a12176a,a12177a,a12180a,a12184a,a12185a,a12186a,a12189a,a12193a,a12194a,a12195a,a12198a,a12202a,a12203a,a12204a,a12207a,a12211a,a12212a,a12213a,a12216a,a12220a,a12221a,a12222a,a12225a,a12229a,a12230a,a12231a,a12234a,a12238a,a12239a,a12240a,a12243a,a12247a,a12248a,a12249a,a12252a,a12256a,a12257a,a12258a,a12261a,a12265a,a12266a,a12267a,a12270a,a12274a,a12275a,a12276a,a12279a,a12283a,a12284a,a12285a,a12288a,a12292a,a12293a,a12294a,a12297a,a12301a,a12302a,a12303a,a12306a,a12310a,a12311a,a12312a,a12315a,a12319a,a12320a,a12321a,a12324a,a12328a,a12329a,a12330a,a12333a,a12337a,a12338a,a12339a,a12342a,a12346a,a12347a,a12348a,a12351a,a12355a,a12356a,a12357a,a12360a,a12364a,a12365a,a12366a,a12369a,a12373a,a12374a,a12375a,a12378a,a12382a,a12383a,a12384a,a12387a,a12391a,a12392a,a12393a,a12396a,a12400a,a12401a,a12402a,a12405a,a12409a,a12410a,a12411a,a12414a,a12418a,a12419a,a12420a,a12423a,a12427a,a12428a,a12429a,a12432a,a12436a,a12437a,a12438a,a12441a,a12445a,a12446a,a12447a,a12450a,a12454a,a12455a,a12456a,a12459a,a12463a,a12464a,a12465a,a12468a,a12472a,a12473a,a12474a,a12477a,a12481a,a12482a,a12483a,a12486a,a12490a,a12491a,a12492a,a12495a,a12499a,a12500a,a12501a,a12504a,a12508a,a12509a,a12510a,a12513a,a12517a,a12518a,a12519a,a12522a,a12526a,a12527a,a12528a,a12531a,a12535a,a12536a,a12537a,a12540a,a12544a,a12545a,a12546a,a12549a,a12553a,a12554a,a12555a,a12558a,a12562a,a12563a,a12564a,a12567a,a12571a,a12572a,a12573a,a12576a,a12580a,a12581a,a12582a,a12585a,a12589a,a12590a,a12591a,a12594a,a12598a,a12599a,a12600a,a12603a,a12607a,a12608a,a12609a,a12612a,a12616a,a12617a,a12618a,a12621a,a12625a,a12626a,a12627a,a12630a,a12634a,a12635a,a12636a,a12639a,a12643a,a12644a,a12645a,a12648a,a12652a,a12653a,a12654a,a12657a,a12661a,a12662a,a12663a,a12666a,a12670a,a12671a,a12672a,a12675a,a12679a,a12680a,a12681a,a12684a,a12688a,a12689a,a12690a,a12693a,a12697a,a12698a,a12699a,a12702a,a12706a,a12707a,a12708a,a12711a,a12715a,a12716a,a12717a,a12720a,a12724a,a12725a,a12726a,a12729a,a12733a,a12734a,a12735a,a12738a,a12742a,a12743a,a12744a,a12747a,a12751a,a12752a,a12753a,a12756a,a12760a,a12761a,a12762a,a12765a,a12769a,a12770a,a12771a,a12774a,a12778a,a12779a,a12780a,a12783a,a12787a,a12788a,a12789a,a12792a,a12796a,a12797a,a12798a,a12801a,a12805a,a12806a,a12807a,a12810a,a12814a,a12815a,a12816a,a12819a,a12823a,a12824a,a12825a,a12828a,a12832a,a12833a,a12834a,a12837a,a12841a,a12842a,a12843a,a12846a,a12850a,a12851a,a12852a,a12855a,a12859a,a12860a,a12861a,a12864a,a12868a,a12869a,a12870a,a12873a,a12877a,a12878a,a12879a,a12882a,a12886a,a12887a,a12888a,a12891a,a12895a,a12896a,a12897a,a12900a,a12904a,a12905a,a12906a,a12909a,a12913a,a12914a,a12915a,a12918a,a12922a,a12923a,a12924a,a12927a,a12931a,a12932a,a12933a,a12936a,a12940a,a12941a,a12942a,a12945a,a12949a,a12950a,a12951a,a12954a,a12958a,a12959a,a12960a,a12963a,a12967a,a12968a,a12969a,a12972a,a12976a,a12977a,a12978a,a12981a,a12985a,a12986a,a12987a,a12990a,a12994a,a12995a,a12996a,a12999a,a13003a,a13004a,a13005a,a13008a,a13012a,a13013a,a13014a,a13017a,a13021a,a13022a,a13023a,a13026a,a13030a,a13031a,a13032a,a13035a,a13039a,a13040a,a13041a,a13044a,a13048a,a13049a,a13050a,a13053a,a13057a,a13058a,a13059a,a13062a,a13066a,a13067a,a13068a,a13071a,a13075a,a13076a,a13077a,a13080a,a13084a,a13085a,a13086a,a13089a,a13093a,a13094a,a13095a,a13098a,a13102a,a13103a,a13104a,a13107a,a13111a,a13112a,a13113a,a13116a,a13120a,a13121a,a13122a,a13125a,a13129a,a13130a,a13131a,a13134a,a13138a,a13139a,a13140a,a13143a,a13147a,a13148a,a13149a,a13152a,a13156a,a13157a,a13158a,a13161a,a13165a,a13166a,a13167a,a13170a,a13174a,a13175a,a13176a,a13179a,a13183a,a13184a,a13185a,a13188a,a13192a,a13193a,a13194a,a13197a,a13201a,a13202a,a13203a,a13206a,a13210a,a13211a,a13212a,a13215a,a13219a,a13220a,a13221a,a13224a,a13228a,a13229a,a13230a,a13233a,a13237a,a13238a,a13239a,a13242a,a13246a,a13247a,a13248a,a13251a,a13255a,a13256a,a13257a,a13260a,a13264a,a13265a,a13266a,a13269a,a13273a,a13274a,a13275a,a13278a,a13282a,a13283a,a13284a,a13287a,a13291a,a13292a,a13293a,a13296a,a13300a,a13301a,a13302a,a13305a,a13309a,a13310a,a13311a,a13314a,a13318a,a13319a,a13320a,a13323a,a13327a,a13328a,a13329a,a13332a,a13336a,a13337a,a13338a,a13341a,a13345a,a13346a,a13347a,a13350a,a13354a,a13355a,a13356a,a13359a,a13363a,a13364a,a13365a,a13368a,a13372a,a13373a,a13374a,a13377a,a13381a,a13382a,a13383a,a13386a,a13390a,a13391a,a13392a,a13395a,a13399a,a13400a,a13401a,a13404a,a13408a,a13409a,a13410a,a13413a,a13417a,a13418a,a13419a,a13422a,a13426a,a13427a,a13428a,a13431a,a13435a,a13436a,a13437a,a13440a,a13444a,a13445a,a13446a,a13449a,a13453a,a13454a,a13455a,a13458a,a13462a,a13463a,a13464a,a13467a,a13471a,a13472a,a13473a,a13476a,a13480a,a13481a,a13482a,a13485a,a13489a,a13490a,a13491a,a13494a,a13498a,a13499a,a13500a,a13503a,a13507a,a13508a,a13509a,a13512a,a13516a,a13517a,a13518a,a13521a,a13525a,a13526a,a13527a,a13530a,a13534a,a13535a,a13536a,a13539a,a13543a,a13544a,a13545a,a13548a,a13552a,a13553a,a13554a,a13557a,a13561a,a13562a,a13563a,a13566a,a13570a,a13571a,a13572a,a13575a,a13579a,a13580a,a13581a,a13584a,a13588a,a13589a,a13590a,a13593a,a13597a,a13598a,a13599a,a13602a,a13606a,a13607a,a13608a,a13611a,a13615a,a13616a,a13617a,a13620a,a13624a,a13625a,a13626a,a13629a,a13633a,a13634a,a13635a,a13638a,a13642a,a13643a,a13644a,a13647a,a13651a,a13652a,a13653a,a13656a,a13660a,a13661a,a13662a,a13665a,a13669a,a13670a,a13671a,a13674a,a13678a,a13679a,a13680a,a13683a,a13687a,a13688a,a13689a,a13692a,a13696a,a13697a,a13698a,a13701a,a13705a,a13706a,a13707a,a13710a,a13714a,a13715a,a13716a,a13719a,a13723a,a13724a,a13725a,a13728a,a13732a,a13733a,a13734a,a13737a,a13741a,a13742a,a13743a,a13746a,a13750a,a13751a,a13752a,a13755a,a13759a,a13760a,a13761a,a13764a,a13768a,a13769a,a13770a,a13773a,a13777a,a13778a,a13779a,a13782a,a13786a,a13787a,a13788a,a13791a,a13795a,a13796a,a13797a,a13800a,a13804a,a13805a,a13806a,a13809a,a13813a,a13814a,a13815a,a13818a,a13822a,a13823a,a13824a,a13827a,a13831a,a13832a,a13833a,a13836a,a13840a,a13841a,a13842a,a13845a,a13849a,a13850a,a13851a,a13854a,a13858a,a13859a,a13860a,a13863a,a13867a,a13868a,a13869a,a13872a,a13876a,a13877a,a13878a,a13881a,a13885a,a13886a,a13887a,a13890a,a13894a,a13895a,a13896a,a13899a,a13903a,a13904a,a13905a,a13908a,a13912a,a13913a,a13914a,a13917a,a13921a,a13922a,a13923a,a13926a,a13930a,a13931a,a13932a,a13935a,a13939a,a13940a,a13941a,a13944a,a13948a,a13949a,a13950a,a13953a,a13957a,a13958a,a13959a,a13962a,a13966a,a13967a,a13968a,a13971a,a13975a,a13976a,a13977a,a13980a,a13984a,a13985a,a13986a,a13989a,a13993a,a13994a,a13995a,a13998a,a14002a,a14003a,a14004a,a14007a,a14011a,a14012a,a14013a,a14016a,a14020a,a14021a,a14022a,a14025a,a14029a,a14030a,a14031a,a14034a,a14038a,a14039a,a14040a,a14043a,a14047a,a14048a,a14049a,a14052a,a14056a,a14057a,a14058a,a14061a,a14065a,a14066a,a14067a,a14070a,a14074a,a14075a,a14076a,a14079a,a14083a,a14084a,a14085a,a14088a,a14092a,a14093a,a14094a,a14097a,a14101a,a14102a,a14103a,a14106a,a14110a,a14111a,a14112a,a14115a,a14119a,a14120a,a14121a,a14124a,a14128a,a14129a,a14130a,a14133a,a14137a,a14138a,a14139a,a14142a,a14146a,a14147a,a14148a,a14151a,a14155a,a14156a,a14157a,a14160a,a14164a,a14165a,a14166a,a14169a,a14173a,a14174a,a14175a,a14178a,a14182a,a14183a,a14184a,a14187a,a14191a,a14192a,a14193a,a14196a,a14200a,a14201a,a14202a,a14205a,a14209a,a14210a,a14211a,a14214a,a14218a,a14219a,a14220a,a14223a,a14227a,a14228a,a14229a,a14232a,a14236a,a14237a,a14238a,a14241a,a14245a,a14246a,a14247a,a14250a,a14254a,a14255a,a14256a,a14259a,a14263a,a14264a,a14265a,a14268a,a14272a,a14273a,a14274a,a14277a,a14281a,a14282a,a14283a,a14286a,a14290a,a14291a,a14292a,a14295a,a14299a,a14300a,a14301a,a14304a,a14308a,a14309a,a14310a,a14313a,a14317a,a14318a,a14319a,a14322a,a14326a,a14327a,a14328a,a14331a,a14335a,a14336a,a14337a,a14340a,a14344a,a14345a,a14346a,a14349a,a14353a,a14354a,a14355a,a14358a,a14362a,a14363a,a14364a,a14367a,a14371a,a14372a,a14373a,a14376a,a14380a,a14381a,a14382a,a14385a,a14389a,a14390a,a14391a,a14394a,a14398a,a14399a,a14400a,a14403a,a14407a,a14408a,a14409a,a14412a,a14416a,a14417a,a14418a,a14421a,a14425a,a14426a,a14427a,a14430a,a14434a,a14435a,a14436a,a14439a,a14443a,a14444a,a14445a,a14448a,a14452a,a14453a,a14454a,a14457a,a14461a,a14462a,a14463a,a14466a,a14470a,a14471a,a14472a,a14475a,a14479a,a14480a,a14481a,a14484a,a14488a,a14489a,a14490a,a14493a,a14497a,a14498a,a14499a,a14502a,a14506a,a14507a,a14508a,a14511a,a14515a,a14516a,a14517a,a14520a,a14524a,a14525a,a14526a,a14529a,a14533a,a14534a,a14535a,a14538a,a14542a,a14543a,a14544a,a14547a,a14551a,a14552a,a14553a,a14556a,a14560a,a14561a,a14562a,a14565a,a14569a,a14570a,a14571a,a14574a,a14578a,a14579a,a14580a,a14583a,a14587a,a14588a,a14589a,a14592a,a14596a,a14597a,a14598a,a14601a,a14605a,a14606a,a14607a,a14610a,a14614a,a14615a,a14616a,a14619a,a14623a,a14624a,a14625a,a14628a,a14632a,a14633a,a14634a,a14637a,a14641a,a14642a,a14643a,a14646a,a14650a,a14651a,a14652a,a14655a,a14659a,a14660a,a14661a,a14664a,a14668a,a14669a,a14670a,a14673a,a14677a,a14678a,a14679a,a14682a,a14686a,a14687a,a14688a,a14691a,a14695a,a14696a,a14697a,a14700a,a14704a,a14705a,a14706a,a14709a,a14713a,a14714a,a14715a,a14718a,a14722a,a14723a,a14724a,a14727a,a14731a,a14732a,a14733a,a14736a,a14740a,a14741a,a14742a,a14745a,a14749a,a14750a,a14751a,a14754a,a14758a,a14759a,a14760a,a14763a,a14767a,a14768a,a14769a,a14772a,a14776a,a14777a,a14778a,a14781a,a14785a,a14786a,a14787a,a14790a,a14794a,a14795a,a14796a,a14799a,a14803a,a14804a,a14805a,a14808a,a14812a,a14813a,a14814a,a14817a,a14821a,a14822a,a14823a,a14826a,a14830a,a14831a,a14832a,a14835a,a14839a,a14840a,a14841a,a14844a,a14848a,a14849a,a14850a,a14853a,a14857a,a14858a,a14859a,a14862a,a14866a,a14867a,a14868a,a14871a,a14875a,a14876a,a14877a,a14880a,a14884a,a14885a,a14886a,a14889a,a14893a,a14894a,a14895a,a14898a,a14902a,a14903a,a14904a,a14907a,a14911a,a14912a,a14913a,a14916a,a14920a,a14921a,a14922a,a14925a,a14929a,a14930a,a14931a,a14934a,a14938a,a14939a,a14940a,a14943a,a14947a,a14948a,a14949a,a14952a,a14956a,a14957a,a14958a,a14961a,a14965a,a14966a,a14967a,a14970a,a14974a,a14975a,a14976a,a14979a,a14983a,a14984a,a14985a,a14988a,a14992a,a14993a,a14994a,a14997a,a15001a,a15002a,a15003a,a15006a,a15010a,a15011a,a15012a,a15015a,a15019a,a15020a,a15021a,a15024a,a15028a,a15029a,a15030a,a15033a,a15037a,a15038a,a15039a,a15042a,a15046a,a15047a,a15048a,a15051a,a15055a,a15056a,a15057a,a15060a,a15064a,a15065a,a15066a,a15069a,a15073a,a15074a,a15075a,a15078a,a15082a,a15083a,a15084a,a15087a,a15091a,a15092a,a15093a,a15096a,a15100a,a15101a,a15102a,a15105a,a15109a,a15110a,a15111a,a15114a,a15118a,a15119a,a15120a,a15123a,a15127a,a15128a,a15129a,a15132a,a15136a,a15137a,a15138a,a15141a,a15145a,a15146a,a15147a,a15150a,a15154a,a15155a,a15156a,a15159a,a15163a,a15164a,a15165a,a15168a,a15172a,a15173a,a15174a,a15177a,a15181a,a15182a,a15183a,a15186a,a15190a,a15191a,a15192a,a15195a,a15199a,a15200a,a15201a,a15204a,a15208a,a15209a,a15210a,a15213a,a15217a,a15218a,a15219a,a15222a,a15226a,a15227a,a15228a,a15231a,a15235a,a15236a,a15237a,a15240a,a15244a,a15245a,a15246a,a15249a,a15253a,a15254a,a15255a,a15258a,a15262a,a15263a,a15264a,a15267a,a15271a,a15272a,a15273a,a15276a,a15280a,a15281a,a15282a,a15285a,a15289a,a15290a,a15291a,a15294a,a15298a,a15299a,a15300a,a15303a,a15307a,a15308a,a15309a,a15312a,a15316a,a15317a,a15318a,a15321a,a15325a,a15326a,a15327a,a15330a,a15334a,a15335a,a15336a,a15339a,a15343a,a15344a,a15345a,a15348a,a15352a,a15353a,a15354a,a15357a,a15361a,a15362a,a15363a,a15366a,a15370a,a15371a,a15372a,a15375a,a15379a,a15380a,a15381a,a15384a,a15388a,a15389a,a15390a,a15393a,a15397a,a15398a,a15399a,a15402a,a15406a,a15407a,a15408a,a15411a,a15415a,a15416a,a15417a,a15420a,a15424a,a15425a,a15426a,a15429a,a15433a,a15434a,a15435a,a15438a,a15442a,a15443a,a15444a,a15447a,a15451a,a15452a,a15453a,a15456a,a15460a,a15461a,a15462a,a15465a,a15469a,a15470a,a15471a,a15474a,a15478a,a15479a,a15480a,a15483a,a15487a,a15488a,a15489a,a15492a,a15496a,a15497a,a15498a,a15501a,a15505a,a15506a,a15507a,a15510a,a15514a,a15515a,a15516a,a15519a,a15523a,a15524a,a15525a,a15528a,a15532a,a15533a,a15534a,a15537a,a15541a,a15542a,a15543a,a15546a,a15550a,a15551a,a15552a,a15555a,a15559a,a15560a,a15561a,a15564a,a15568a,a15569a,a15570a,a15573a,a15577a,a15578a,a15579a,a15582a,a15586a,a15587a,a15588a,a15591a,a15595a,a15596a,a15597a,a15600a,a15604a,a15605a,a15606a,a15609a,a15613a,a15614a,a15615a,a15618a,a15622a,a15623a,a15624a,a15627a,a15631a,a15632a,a15633a,a15636a,a15640a,a15641a,a15642a,a15645a,a15649a,a15650a,a15651a,a15654a,a15658a,a15659a,a15660a,a15663a,a15667a,a15668a,a15669a,a15672a,a15676a,a15677a,a15678a,a15681a,a15685a,a15686a,a15687a,a15690a,a15694a,a15695a,a15696a,a15699a,a15703a,a15704a,a15705a,a15708a,a15712a,a15713a,a15714a,a15717a,a15721a,a15722a,a15723a,a15726a,a15730a,a15731a,a15732a,a15735a,a15739a,a15740a,a15741a,a15744a,a15748a,a15749a,a15750a,a15753a,a15757a,a15758a,a15759a,a15762a,a15766a,a15767a,a15768a,a15771a,a15775a,a15776a,a15777a,a15780a,a15784a,a15785a,a15786a,a15789a,a15793a,a15794a,a15795a,a15798a,a15802a,a15803a,a15804a,a15807a,a15811a,a15812a,a15813a,a15816a,a15820a,a15821a,a15822a,a15825a,a15829a,a15830a,a15831a,a15834a,a15838a,a15839a,a15840a,a15843a,a15847a,a15848a,a15849a,a15852a,a15856a,a15857a,a15858a,a15861a,a15865a,a15866a,a15867a,a15870a,a15874a,a15875a,a15876a,a15879a,a15883a,a15884a,a15885a,a15888a,a15892a,a15893a,a15894a,a15897a,a15901a,a15902a,a15903a,a15906a,a15910a,a15911a,a15912a,a15915a,a15919a,a15920a,a15921a,a15924a,a15928a,a15929a,a15930a,a15933a,a15937a,a15938a,a15939a,a15942a,a15946a,a15947a,a15948a,a15951a,a15955a,a15956a,a15957a,a15960a,a15964a,a15965a,a15966a,a15969a,a15973a,a15974a,a15975a,a15978a,a15982a,a15983a,a15984a,a15987a,a15991a,a15992a,a15993a,a15996a,a16000a,a16001a,a16002a,a16005a,a16009a,a16010a,a16011a,a16014a,a16018a,a16019a,a16020a,a16023a,a16027a,a16028a,a16029a,a16032a,a16036a,a16037a,a16038a,a16041a,a16045a,a16046a,a16047a,a16051a,a16052a,a16056a,a16057a,a16058a,a16061a,a16065a,a16066a,a16067a,a16071a,a16072a,a16076a,a16077a,a16078a,a16081a,a16085a,a16086a,a16087a,a16091a,a16092a,a16096a,a16097a,a16098a,a16101a,a16105a,a16106a,a16107a,a16111a,a16112a,a16116a,a16117a,a16118a,a16121a,a16125a,a16126a,a16127a,a16131a,a16132a,a16136a,a16137a,a16138a,a16141a,a16145a,a16146a,a16147a,a16151a,a16152a,a16156a,a16157a,a16158a,a16161a,a16165a,a16166a,a16167a,a16171a,a16172a,a16176a,a16177a,a16178a,a16181a,a16185a,a16186a,a16187a,a16191a,a16192a,a16196a,a16197a,a16198a,a16201a,a16205a,a16206a,a16207a,a16211a,a16212a,a16216a,a16217a,a16218a,a16221a,a16225a,a16226a,a16227a,a16231a,a16232a,a16236a,a16237a,a16238a,a16241a,a16245a,a16246a,a16247a,a16251a,a16252a,a16256a,a16257a,a16258a,a16261a,a16265a,a16266a,a16267a,a16271a,a16272a,a16276a,a16277a,a16278a,a16281a,a16285a,a16286a,a16287a,a16291a,a16292a,a16296a,a16297a,a16298a,a16301a,a16305a,a16306a,a16307a,a16311a,a16312a,a16316a,a16317a,a16318a,a16321a,a16325a,a16326a,a16327a,a16331a,a16332a,a16336a,a16337a,a16338a,a16341a,a16345a,a16346a,a16347a,a16351a,a16352a,a16356a,a16357a,a16358a,a16361a,a16365a,a16366a,a16367a,a16371a,a16372a,a16376a,a16377a,a16378a,a16381a,a16385a,a16386a,a16387a,a16391a,a16392a,a16396a,a16397a,a16398a,a16401a,a16405a,a16406a,a16407a,a16411a,a16412a,a16416a,a16417a,a16418a,a16421a,a16425a,a16426a,a16427a,a16431a,a16432a,a16436a,a16437a,a16438a,a16441a,a16445a,a16446a,a16447a,a16451a,a16452a,a16456a,a16457a,a16458a,a16461a,a16465a,a16466a,a16467a,a16471a,a16472a,a16476a,a16477a,a16478a,a16481a,a16485a,a16486a,a16487a,a16491a,a16492a,a16496a,a16497a,a16498a,a16501a,a16505a,a16506a,a16507a,a16511a,a16512a,a16516a,a16517a,a16518a,a16521a,a16525a,a16526a,a16527a,a16531a,a16532a,a16536a,a16537a,a16538a,a16541a,a16545a,a16546a,a16547a,a16551a,a16552a,a16556a,a16557a,a16558a,a16561a,a16565a,a16566a,a16567a,a16571a,a16572a,a16576a,a16577a,a16578a,a16581a,a16585a,a16586a,a16587a,a16591a,a16592a,a16596a,a16597a,a16598a,a16601a,a16605a,a16606a,a16607a,a16611a,a16612a,a16616a,a16617a,a16618a,a16621a,a16625a,a16626a,a16627a,a16631a,a16632a,a16636a,a16637a,a16638a,a16641a,a16645a,a16646a,a16647a,a16651a,a16652a,a16656a,a16657a,a16658a,a16661a,a16665a,a16666a,a16667a,a16671a,a16672a,a16676a,a16677a,a16678a,a16681a,a16685a,a16686a,a16687a,a16691a,a16692a,a16696a,a16697a,a16698a,a16701a,a16705a,a16706a,a16707a,a16711a,a16712a,a16716a,a16717a,a16718a,a16721a,a16725a,a16726a,a16727a,a16731a,a16732a,a16736a,a16737a,a16738a,a16741a,a16745a,a16746a,a16747a,a16751a,a16752a,a16756a,a16757a,a16758a,a16761a,a16765a,a16766a,a16767a,a16771a,a16772a,a16776a,a16777a,a16778a,a16781a,a16785a,a16786a,a16787a,a16791a,a16792a,a16796a,a16797a,a16798a,a16801a,a16805a,a16806a,a16807a,a16811a,a16812a,a16816a,a16817a,a16818a,a16821a,a16825a,a16826a,a16827a,a16831a,a16832a,a16836a,a16837a,a16838a,a16841a,a16845a,a16846a,a16847a,a16851a,a16852a,a16856a,a16857a,a16858a,a16861a,a16865a,a16866a,a16867a,a16871a,a16872a,a16876a,a16877a,a16878a,a16881a,a16885a,a16886a,a16887a,a16891a,a16892a,a16896a,a16897a,a16898a,a16901a,a16905a,a16906a,a16907a,a16911a,a16912a,a16916a,a16917a,a16918a,a16921a,a16925a,a16926a,a16927a,a16931a,a16932a,a16936a,a16937a,a16938a,a16941a,a16945a,a16946a,a16947a,a16951a,a16952a,a16956a,a16957a,a16958a,a16961a,a16965a,a16966a,a16967a,a16971a,a16972a,a16976a,a16977a,a16978a,a16981a,a16985a,a16986a,a16987a,a16991a,a16992a,a16996a,a16997a,a16998a,a17001a,a17005a,a17006a,a17007a,a17011a,a17012a,a17016a,a17017a,a17018a,a17021a,a17025a,a17026a,a17027a,a17031a,a17032a,a17036a,a17037a,a17038a,a17041a,a17045a,a17046a,a17047a,a17051a,a17052a,a17056a,a17057a,a17058a,a17061a,a17065a,a17066a,a17067a,a17071a,a17072a,a17076a,a17077a,a17078a,a17081a,a17085a,a17086a,a17087a,a17091a,a17092a,a17096a,a17097a,a17098a,a17101a,a17105a,a17106a,a17107a,a17111a,a17112a,a17116a,a17117a,a17118a,a17121a,a17125a,a17126a,a17127a,a17131a,a17132a,a17136a,a17137a,a17138a,a17141a,a17145a,a17146a,a17147a,a17151a,a17152a,a17156a,a17157a,a17158a,a17161a,a17165a,a17166a,a17167a,a17171a,a17172a,a17176a,a17177a,a17178a,a17181a,a17185a,a17186a,a17187a,a17191a,a17192a,a17196a,a17197a,a17198a,a17201a,a17205a,a17206a,a17207a,a17211a,a17212a,a17216a,a17217a,a17218a,a17221a,a17225a,a17226a,a17227a,a17231a,a17232a,a17236a,a17237a,a17238a,a17241a,a17245a,a17246a,a17247a,a17251a,a17252a,a17256a,a17257a,a17258a,a17261a,a17265a,a17266a,a17267a,a17271a,a17272a,a17276a,a17277a,a17278a,a17281a,a17285a,a17286a,a17287a,a17291a,a17292a,a17296a,a17297a,a17298a,a17301a,a17305a,a17306a,a17307a,a17311a,a17312a,a17316a,a17317a,a17318a,a17321a,a17325a,a17326a,a17327a,a17331a,a17332a,a17336a,a17337a,a17338a,a17341a,a17345a,a17346a,a17347a,a17351a,a17352a,a17356a,a17357a,a17358a,a17361a,a17365a,a17366a,a17367a,a17371a,a17372a,a17376a,a17377a,a17378a,a17381a,a17385a,a17386a,a17387a,a17391a,a17392a,a17396a,a17397a,a17398a,a17401a,a17405a,a17406a,a17407a,a17411a,a17412a,a17416a,a17417a,a17418a,a17421a,a17425a,a17426a,a17427a,a17431a,a17432a,a17436a,a17437a,a17438a,a17441a,a17445a,a17446a,a17447a,a17451a,a17452a,a17456a,a17457a,a17458a,a17461a,a17465a,a17466a,a17467a,a17471a,a17472a,a17476a,a17477a,a17478a,a17481a,a17485a,a17486a,a17487a,a17491a,a17492a,a17496a,a17497a,a17498a,a17501a,a17505a,a17506a,a17507a,a17511a,a17512a,a17516a,a17517a,a17518a,a17521a,a17525a,a17526a,a17527a,a17531a,a17532a,a17536a,a17537a,a17538a,a17541a,a17545a,a17546a,a17547a,a17551a,a17552a,a17556a,a17557a,a17558a,a17561a,a17565a,a17566a,a17567a,a17571a,a17572a,a17576a,a17577a,a17578a,a17581a,a17585a,a17586a,a17587a,a17591a,a17592a,a17596a,a17597a,a17598a,a17601a,a17605a,a17606a,a17607a,a17611a,a17612a,a17616a,a17617a,a17618a,a17621a,a17625a,a17626a,a17627a,a17631a,a17632a,a17636a,a17637a,a17638a,a17641a,a17645a,a17646a,a17647a,a17651a,a17652a,a17656a,a17657a,a17658a,a17661a,a17665a,a17666a,a17667a,a17671a,a17672a,a17676a,a17677a,a17678a,a17681a,a17685a,a17686a,a17687a,a17691a,a17692a,a17696a,a17697a,a17698a,a17701a,a17705a,a17706a,a17707a,a17711a,a17712a,a17716a,a17717a,a17718a,a17721a,a17725a,a17726a,a17727a,a17731a,a17732a,a17736a,a17737a,a17738a,a17741a,a17745a,a17746a,a17747a,a17751a,a17752a,a17756a,a17757a,a17758a,a17761a,a17765a,a17766a,a17767a,a17771a,a17772a,a17776a,a17777a,a17778a,a17781a,a17785a,a17786a,a17787a,a17791a,a17792a,a17796a,a17797a,a17798a,a17801a,a17805a,a17806a,a17807a,a17811a,a17812a,a17816a,a17817a,a17818a,a17821a,a17825a,a17826a,a17827a,a17831a,a17832a,a17836a,a17837a,a17838a,a17841a,a17845a,a17846a,a17847a,a17851a,a17852a,a17856a,a17857a,a17858a,a17861a,a17865a,a17866a,a17867a,a17871a,a17872a,a17876a,a17877a,a17878a,a17881a,a17885a,a17886a,a17887a,a17891a,a17892a,a17896a,a17897a,a17898a,a17901a,a17905a,a17906a,a17907a,a17911a,a17912a,a17916a,a17917a,a17918a,a17921a,a17925a,a17926a,a17927a,a17931a,a17932a,a17936a,a17937a,a17938a,a17941a,a17945a,a17946a,a17947a,a17951a,a17952a,a17956a,a17957a,a17958a,a17961a,a17965a,a17966a,a17967a,a17971a,a17972a,a17976a,a17977a,a17978a,a17981a,a17985a,a17986a,a17987a,a17991a,a17992a,a17996a,a17997a,a17998a,a18001a,a18005a,a18006a,a18007a,a18011a,a18012a,a18016a,a18017a,a18018a,a18021a,a18025a,a18026a,a18027a,a18031a,a18032a,a18036a,a18037a,a18038a,a18041a,a18045a,a18046a,a18047a,a18051a,a18052a,a18056a,a18057a,a18058a,a18061a,a18065a,a18066a,a18067a,a18071a,a18072a,a18076a,a18077a,a18078a,a18081a,a18085a,a18086a,a18087a,a18091a,a18092a,a18096a,a18097a,a18098a,a18101a,a18105a,a18106a,a18107a,a18111a,a18112a,a18116a,a18117a,a18118a,a18121a,a18125a,a18126a,a18127a,a18131a,a18132a,a18136a,a18137a,a18138a,a18141a,a18145a,a18146a,a18147a,a18151a,a18152a,a18156a,a18157a,a18158a,a18161a,a18165a,a18166a,a18167a,a18171a,a18172a,a18176a,a18177a,a18178a,a18181a,a18185a,a18186a,a18187a,a18191a,a18192a,a18196a,a18197a,a18198a,a18201a,a18205a,a18206a,a18207a,a18211a,a18212a,a18216a,a18217a,a18218a,a18221a,a18225a,a18226a,a18227a,a18231a,a18232a,a18236a,a18237a,a18238a,a18241a,a18245a,a18246a,a18247a,a18251a,a18252a,a18256a,a18257a,a18258a,a18261a,a18265a,a18266a,a18267a,a18271a,a18272a,a18276a,a18277a,a18278a,a18281a,a18285a,a18286a,a18287a,a18291a,a18292a,a18296a,a18297a,a18298a,a18301a,a18305a,a18306a,a18307a,a18311a,a18312a,a18316a,a18317a,a18318a,a18321a,a18325a,a18326a,a18327a,a18331a,a18332a,a18336a,a18337a,a18338a,a18341a,a18345a,a18346a,a18347a,a18351a,a18352a,a18356a,a18357a,a18358a,a18361a,a18365a,a18366a,a18367a,a18371a,a18372a,a18376a,a18377a,a18378a,a18381a,a18385a,a18386a,a18387a,a18391a,a18392a,a18396a,a18397a,a18398a,a18401a,a18405a,a18406a,a18407a,a18411a,a18412a,a18416a,a18417a,a18418a,a18421a,a18425a,a18426a,a18427a,a18431a,a18432a,a18436a,a18437a,a18438a,a18441a,a18445a,a18446a,a18447a,a18451a,a18452a,a18456a,a18457a,a18458a,a18461a,a18465a,a18466a,a18467a,a18471a,a18472a,a18476a,a18477a,a18478a,a18481a,a18485a,a18486a,a18487a,a18491a,a18492a,a18496a,a18497a,a18498a,a18501a,a18505a,a18506a,a18507a,a18511a,a18512a,a18516a,a18517a,a18518a,a18521a,a18525a,a18526a,a18527a,a18531a,a18532a,a18536a,a18537a,a18538a,a18541a,a18545a,a18546a,a18547a,a18551a,a18552a,a18556a,a18557a,a18558a,a18561a,a18565a,a18566a,a18567a,a18571a,a18572a,a18576a,a18577a,a18578a,a18581a,a18585a,a18586a,a18587a,a18591a,a18592a,a18596a,a18597a,a18598a,a18601a,a18605a,a18606a,a18607a,a18611a,a18612a,a18616a,a18617a,a18618a,a18621a,a18625a,a18626a,a18627a,a18631a,a18632a,a18636a,a18637a,a18638a,a18641a,a18645a,a18646a,a18647a,a18651a,a18652a,a18656a,a18657a,a18658a,a18661a,a18665a,a18666a,a18667a,a18671a,a18672a,a18676a,a18677a,a18678a,a18681a,a18685a,a18686a,a18687a,a18691a,a18692a,a18696a,a18697a,a18698a,a18701a,a18705a,a18706a,a18707a,a18711a,a18712a,a18716a,a18717a,a18718a,a18721a,a18725a,a18726a,a18727a,a18731a,a18732a,a18736a,a18737a,a18738a,a18741a,a18745a,a18746a,a18747a,a18751a,a18752a,a18756a,a18757a,a18758a,a18761a,a18765a,a18766a,a18767a,a18771a,a18772a,a18776a,a18777a,a18778a,a18781a,a18785a,a18786a,a18787a,a18791a,a18792a,a18796a,a18797a,a18798a,a18801a,a18805a,a18806a,a18807a,a18811a,a18812a,a18816a,a18817a,a18818a,a18821a,a18825a,a18826a,a18827a,a18831a,a18832a,a18836a,a18837a,a18838a,a18841a,a18845a,a18846a,a18847a,a18851a,a18852a,a18856a,a18857a,a18858a,a18861a,a18865a,a18866a,a18867a,a18871a,a18872a,a18876a,a18877a,a18878a,a18881a,a18885a,a18886a,a18887a,a18891a,a18892a,a18896a,a18897a,a18898a,a18901a,a18905a,a18906a,a18907a,a18911a,a18912a,a18916a,a18917a,a18918a,a18921a,a18925a,a18926a,a18927a,a18931a,a18932a,a18936a,a18937a,a18938a,a18941a,a18945a,a18946a,a18947a,a18951a,a18952a,a18956a,a18957a,a18958a,a18961a,a18965a,a18966a,a18967a,a18971a,a18972a,a18976a,a18977a,a18978a,a18981a,a18985a,a18986a,a18987a,a18991a,a18992a,a18996a,a18997a,a18998a,a19001a,a19005a,a19006a,a19007a,a19011a,a19012a,a19016a,a19017a,a19018a,a19021a,a19025a,a19026a,a19027a,a19031a,a19032a,a19036a,a19037a,a19038a,a19041a,a19045a,a19046a,a19047a,a19051a,a19052a,a19056a,a19057a,a19058a,a19061a,a19065a,a19066a,a19067a,a19071a,a19072a,a19076a,a19077a,a19078a,a19081a,a19085a,a19086a,a19087a,a19091a,a19092a,a19096a,a19097a,a19098a,a19101a,a19105a,a19106a,a19107a,a19111a,a19112a,a19116a,a19117a,a19118a,a19121a,a19125a,a19126a,a19127a,a19131a,a19132a,a19136a,a19137a,a19138a,a19141a,a19145a,a19146a,a19147a,a19151a,a19152a,a19156a,a19157a,a19158a,a19161a,a19165a,a19166a,a19167a,a19171a,a19172a,a19176a,a19177a,a19178a,a19181a,a19185a,a19186a,a19187a,a19191a,a19192a,a19196a,a19197a,a19198a,a19201a,a19205a,a19206a,a19207a,a19211a,a19212a,a19216a,a19217a,a19218a,a19221a,a19225a,a19226a,a19227a,a19231a,a19232a,a19236a,a19237a,a19238a,a19241a,a19245a,a19246a,a19247a,a19251a,a19252a,a19256a,a19257a,a19258a,a19261a,a19265a,a19266a,a19267a,a19271a,a19272a,a19276a,a19277a,a19278a,a19281a,a19285a,a19286a,a19287a,a19291a,a19292a,a19296a,a19297a,a19298a,a19301a,a19305a,a19306a,a19307a,a19311a,a19312a,a19316a,a19317a,a19318a,a19321a,a19325a,a19326a,a19327a,a19331a,a19332a,a19336a,a19337a,a19338a,a19341a,a19345a,a19346a,a19347a,a19351a,a19352a,a19356a,a19357a,a19358a,a19361a,a19365a,a19366a,a19367a,a19371a,a19372a,a19376a,a19377a,a19378a,a19381a,a19385a,a19386a,a19387a,a19391a,a19392a,a19396a,a19397a,a19398a,a19401a,a19405a,a19406a,a19407a,a19411a,a19412a,a19416a,a19417a,a19418a,a19421a,a19425a,a19426a,a19427a,a19431a,a19432a,a19436a,a19437a,a19438a,a19441a,a19445a,a19446a,a19447a,a19451a,a19452a,a19456a,a19457a,a19458a,a19461a,a19465a,a19466a,a19467a,a19471a,a19472a,a19476a,a19477a,a19478a,a19481a,a19485a,a19486a,a19487a,a19491a,a19492a,a19496a,a19497a,a19498a,a19501a,a19505a,a19506a,a19507a,a19511a,a19512a,a19516a,a19517a,a19518a,a19521a,a19525a,a19526a,a19527a,a19531a,a19532a,a19536a,a19537a,a19538a,a19541a,a19545a,a19546a,a19547a,a19551a,a19552a,a19556a,a19557a,a19558a,a19561a,a19565a,a19566a,a19567a,a19571a,a19572a,a19576a,a19577a,a19578a,a19581a,a19585a,a19586a,a19587a,a19591a,a19592a,a19596a,a19597a,a19598a,a19601a,a19605a,a19606a,a19607a,a19611a,a19612a,a19616a,a19617a,a19618a,a19621a,a19625a,a19626a,a19627a,a19631a,a19632a,a19636a,a19637a,a19638a,a19641a,a19645a,a19646a,a19647a,a19651a,a19652a,a19656a,a19657a,a19658a,a19661a,a19665a,a19666a,a19667a,a19671a,a19672a,a19676a,a19677a,a19678a,a19681a,a19685a,a19686a,a19687a,a19691a,a19692a,a19696a,a19697a,a19698a,a19701a,a19705a,a19706a,a19707a,a19711a,a19712a,a19716a,a19717a,a19718a,a19721a,a19725a,a19726a,a19727a,a19731a,a19732a,a19736a,a19737a,a19738a,a19741a,a19745a,a19746a,a19747a,a19751a,a19752a,a19756a,a19757a,a19758a,a19761a,a19765a,a19766a,a19767a,a19771a,a19772a,a19776a,a19777a,a19778a,a19781a,a19785a,a19786a,a19787a,a19791a,a19792a,a19796a,a19797a,a19798a,a19801a,a19805a,a19806a,a19807a,a19811a,a19812a,a19816a,a19817a,a19818a,a19821a,a19825a,a19826a,a19827a,a19831a,a19832a,a19836a,a19837a,a19838a,a19841a,a19845a,a19846a,a19847a,a19851a,a19852a,a19856a,a19857a,a19858a,a19861a,a19865a,a19866a,a19867a,a19871a,a19872a,a19876a,a19877a,a19878a,a19881a,a19885a,a19886a,a19887a,a19891a,a19892a,a19896a,a19897a,a19898a,a19901a,a19905a,a19906a,a19907a,a19911a,a19912a,a19916a,a19917a,a19918a,a19921a,a19925a,a19926a,a19927a,a19931a,a19932a,a19936a,a19937a,a19938a,a19941a,a19945a,a19946a,a19947a,a19951a,a19952a,a19956a,a19957a,a19958a,a19961a,a19965a,a19966a,a19967a,a19971a,a19972a,a19976a,a19977a,a19978a,a19981a,a19985a,a19986a,a19987a,a19991a,a19992a,a19996a,a19997a,a19998a,a20001a,a20005a,a20006a,a20007a,a20011a,a20012a,a20016a,a20017a,a20018a,a20021a,a20025a,a20026a,a20027a,a20031a,a20032a,a20036a,a20037a,a20038a,a20041a,a20045a,a20046a,a20047a,a20051a,a20052a,a20056a,a20057a,a20058a,a20061a,a20065a,a20066a,a20067a,a20071a,a20072a,a20076a,a20077a,a20078a,a20081a,a20085a,a20086a,a20087a,a20091a,a20092a,a20096a,a20097a,a20098a,a20101a,a20105a,a20106a,a20107a,a20111a,a20112a,a20116a,a20117a,a20118a,a20121a,a20125a,a20126a,a20127a,a20131a,a20132a,a20136a,a20137a,a20138a,a20141a,a20145a,a20146a,a20147a,a20151a,a20152a,a20156a,a20157a,a20158a,a20161a,a20165a,a20166a,a20167a,a20171a,a20172a,a20176a,a20177a,a20178a,a20181a,a20185a,a20186a,a20187a,a20191a,a20192a,a20196a,a20197a,a20198a,a20201a,a20205a,a20206a,a20207a,a20211a,a20212a,a20216a,a20217a,a20218a,a20221a,a20225a,a20226a,a20227a,a20231a,a20232a,a20236a,a20237a,a20238a,a20241a,a20245a,a20246a,a20247a,a20251a,a20252a,a20256a,a20257a,a20258a,a20261a,a20265a,a20266a,a20267a,a20271a,a20272a,a20276a,a20277a,a20278a,a20281a,a20285a,a20286a,a20287a,a20291a,a20292a,a20296a,a20297a,a20298a,a20301a,a20305a,a20306a,a20307a,a20311a,a20312a,a20316a,a20317a,a20318a,a20321a,a20325a,a20326a,a20327a,a20331a,a20332a,a20336a,a20337a,a20338a,a20341a,a20345a,a20346a,a20347a,a20351a,a20352a,a20356a,a20357a,a20358a,a20361a,a20365a,a20366a,a20367a,a20371a,a20372a,a20376a,a20377a,a20378a,a20381a,a20385a,a20386a,a20387a,a20391a,a20392a,a20396a,a20397a,a20398a,a20401a,a20405a,a20406a,a20407a,a20411a,a20412a,a20416a,a20417a,a20418a,a20421a,a20425a,a20426a,a20427a,a20431a,a20432a,a20436a,a20437a,a20438a,a20441a,a20445a,a20446a,a20447a,a20451a,a20452a,a20456a,a20457a,a20458a,a20461a,a20465a,a20466a,a20467a,a20471a,a20472a,a20476a,a20477a,a20478a,a20481a,a20485a,a20486a,a20487a,a20491a,a20492a,a20496a,a20497a,a20498a,a20501a,a20505a,a20506a,a20507a,a20511a,a20512a,a20516a,a20517a,a20518a,a20521a,a20525a,a20526a,a20527a,a20531a,a20532a,a20536a,a20537a,a20538a,a20541a,a20545a,a20546a,a20547a,a20551a,a20552a,a20556a,a20557a,a20558a,a20561a,a20565a,a20566a,a20567a,a20571a,a20572a,a20576a,a20577a,a20578a,a20581a,a20585a,a20586a,a20587a,a20591a,a20592a,a20596a,a20597a,a20598a,a20601a,a20605a,a20606a,a20607a,a20611a,a20612a,a20616a,a20617a,a20618a,a20621a,a20625a,a20626a,a20627a,a20631a,a20632a,a20636a,a20637a,a20638a,a20641a,a20645a,a20646a,a20647a,a20651a,a20652a,a20656a,a20657a,a20658a,a20661a,a20665a,a20666a,a20667a,a20671a,a20672a,a20676a,a20677a,a20678a,a20681a,a20685a,a20686a,a20687a,a20691a,a20692a,a20696a,a20697a,a20698a,a20701a,a20705a,a20706a,a20707a,a20711a,a20712a,a20716a,a20717a,a20718a,a20721a,a20725a,a20726a,a20727a,a20731a,a20732a,a20736a,a20737a,a20738a,a20741a,a20745a,a20746a,a20747a,a20751a,a20752a,a20756a,a20757a,a20758a,a20761a,a20765a,a20766a,a20767a,a20771a,a20772a,a20776a,a20777a,a20778a,a20781a,a20785a,a20786a,a20787a,a20791a,a20792a,a20796a,a20797a,a20798a,a20801a,a20805a,a20806a,a20807a,a20811a,a20812a,a20816a,a20817a,a20818a,a20821a,a20825a,a20826a,a20827a,a20831a,a20832a,a20836a,a20837a,a20838a,a20841a,a20845a,a20846a,a20847a,a20851a,a20852a,a20856a,a20857a,a20858a,a20861a,a20865a,a20866a,a20867a,a20871a,a20872a,a20876a,a20877a,a20878a,a20881a,a20885a,a20886a,a20887a,a20891a,a20892a,a20896a,a20897a,a20898a,a20901a,a20905a,a20906a,a20907a,a20911a,a20912a,a20916a,a20917a,a20918a,a20921a,a20925a,a20926a,a20927a,a20931a,a20932a,a20936a,a20937a,a20938a,a20941a,a20945a,a20946a,a20947a,a20951a,a20952a,a20956a,a20957a,a20958a,a20961a,a20965a,a20966a,a20967a,a20971a,a20972a,a20976a,a20977a,a20978a,a20981a,a20985a,a20986a,a20987a,a20991a,a20992a,a20996a,a20997a,a20998a,a21001a,a21005a,a21006a,a21007a,a21011a,a21012a,a21016a,a21017a,a21018a,a21021a,a21025a,a21026a,a21027a,a21031a,a21032a,a21036a,a21037a,a21038a,a21041a,a21045a,a21046a,a21047a,a21051a,a21052a,a21056a,a21057a,a21058a,a21061a,a21065a,a21066a,a21067a,a21071a,a21072a,a21076a,a21077a,a21078a,a21081a,a21085a,a21086a,a21087a,a21091a,a21092a,a21096a,a21097a,a21098a,a21101a,a21105a,a21106a,a21107a,a21111a,a21112a,a21116a,a21117a,a21118a,a21121a,a21125a,a21126a,a21127a,a21131a,a21132a,a21136a,a21137a,a21138a,a21141a,a21145a,a21146a,a21147a,a21151a,a21152a,a21156a,a21157a,a21158a,a21161a,a21165a,a21166a,a21167a,a21171a,a21172a,a21176a,a21177a,a21178a,a21181a,a21185a,a21186a,a21187a,a21191a,a21192a,a21196a,a21197a,a21198a,a21201a,a21205a,a21206a,a21207a,a21211a,a21212a,a21216a,a21217a,a21218a,a21221a,a21225a,a21226a,a21227a,a21231a,a21232a,a21236a,a21237a,a21238a,a21241a,a21245a,a21246a,a21247a,a21251a,a21252a,a21256a,a21257a,a21258a,a21261a,a21265a,a21266a,a21267a,a21271a,a21272a,a21276a,a21277a,a21278a,a21281a,a21285a,a21286a,a21287a,a21291a,a21292a,a21296a,a21297a,a21298a,a21301a,a21305a,a21306a,a21307a,a21311a,a21312a,a21316a,a21317a,a21318a,a21321a,a21325a,a21326a,a21327a,a21331a,a21332a,a21336a,a21337a,a21338a,a21341a,a21345a,a21346a,a21347a,a21351a,a21352a,a21356a,a21357a,a21358a,a21361a,a21365a,a21366a,a21367a,a21371a,a21372a,a21376a,a21377a,a21378a,a21381a,a21385a,a21386a,a21387a,a21391a,a21392a,a21396a,a21397a,a21398a,a21401a,a21405a,a21406a,a21407a,a21411a,a21412a,a21416a,a21417a,a21418a,a21421a,a21425a,a21426a,a21427a,a21431a,a21432a,a21436a,a21437a,a21438a,a21441a,a21445a,a21446a,a21447a,a21451a,a21452a,a21456a,a21457a,a21458a,a21461a,a21465a,a21466a,a21467a,a21471a,a21472a,a21476a,a21477a,a21478a,a21481a,a21485a,a21486a,a21487a,a21491a,a21492a,a21496a,a21497a,a21498a,a21501a,a21505a,a21506a,a21507a,a21511a,a21512a,a21516a,a21517a,a21518a,a21521a,a21525a,a21526a,a21527a,a21531a,a21532a,a21536a,a21537a,a21538a,a21541a,a21545a,a21546a,a21547a,a21551a,a21552a,a21556a,a21557a,a21558a,a21561a,a21565a,a21566a,a21567a,a21571a,a21572a,a21576a,a21577a,a21578a,a21581a,a21585a,a21586a,a21587a,a21591a,a21592a,a21596a,a21597a,a21598a,a21601a,a21605a,a21606a,a21607a,a21611a,a21612a,a21616a,a21617a,a21618a,a21621a,a21625a,a21626a,a21627a,a21631a,a21632a,a21636a,a21637a,a21638a,a21641a,a21645a,a21646a,a21647a,a21651a,a21652a,a21656a,a21657a,a21658a,a21661a,a21665a,a21666a,a21667a,a21671a,a21672a,a21676a,a21677a,a21678a,a21681a,a21685a,a21686a,a21687a,a21691a,a21692a,a21696a,a21697a,a21698a,a21701a,a21705a,a21706a,a21707a,a21711a,a21712a,a21716a,a21717a,a21718a,a21721a,a21725a,a21726a,a21727a,a21731a,a21732a,a21736a,a21737a,a21738a,a21741a,a21745a,a21746a,a21747a,a21751a,a21752a,a21756a,a21757a,a21758a,a21761a,a21765a,a21766a,a21767a,a21771a,a21772a,a21776a,a21777a,a21778a,a21781a,a21785a,a21786a,a21787a,a21791a,a21792a,a21796a,a21797a,a21798a,a21801a,a21805a,a21806a,a21807a,a21811a,a21812a,a21816a,a21817a,a21818a,a21821a,a21825a,a21826a,a21827a,a21831a,a21832a,a21836a,a21837a,a21838a,a21841a,a21845a,a21846a,a21847a,a21851a,a21852a,a21856a,a21857a,a21858a,a21861a,a21865a,a21866a,a21867a,a21871a,a21872a,a21876a,a21877a,a21878a,a21881a,a21885a,a21886a,a21887a,a21891a,a21892a,a21896a,a21897a,a21898a,a21901a,a21905a,a21906a,a21907a,a21911a,a21912a,a21916a,a21917a,a21918a,a21921a,a21925a,a21926a,a21927a,a21931a,a21932a,a21936a,a21937a,a21938a,a21941a,a21945a,a21946a,a21947a,a21951a,a21952a,a21956a,a21957a,a21958a,a21961a,a21965a,a21966a,a21967a,a21971a,a21972a,a21976a,a21977a,a21978a,a21981a,a21985a,a21986a,a21987a,a21991a,a21992a,a21996a,a21997a,a21998a,a22001a,a22005a,a22006a,a22007a,a22011a,a22012a,a22016a,a22017a,a22018a,a22021a,a22025a,a22026a,a22027a,a22031a,a22032a,a22036a,a22037a,a22038a,a22041a,a22045a,a22046a,a22047a,a22051a,a22052a,a22056a,a22057a,a22058a,a22061a,a22065a,a22066a,a22067a,a22071a,a22072a,a22076a,a22077a,a22078a,a22081a,a22085a,a22086a,a22087a,a22091a,a22092a,a22096a,a22097a,a22098a,a22101a,a22105a,a22106a,a22107a,a22111a,a22112a,a22116a,a22117a,a22118a,a22121a,a22125a,a22126a,a22127a,a22131a,a22132a,a22136a,a22137a,a22138a,a22141a,a22145a,a22146a,a22147a,a22151a,a22152a,a22156a,a22157a,a22158a,a22161a,a22165a,a22166a,a22167a,a22171a,a22172a,a22176a,a22177a,a22178a,a22181a,a22185a,a22186a,a22187a,a22191a,a22192a,a22196a,a22197a,a22198a,a22201a,a22205a,a22206a,a22207a,a22211a,a22212a,a22216a,a22217a,a22218a,a22221a,a22225a,a22226a,a22227a,a22231a,a22232a,a22236a,a22237a,a22238a,a22241a,a22245a,a22246a,a22247a,a22251a,a22252a,a22256a,a22257a,a22258a,a22261a,a22265a,a22266a,a22267a,a22271a,a22272a,a22276a,a22277a,a22278a,a22281a,a22285a,a22286a,a22287a,a22291a,a22292a,a22296a,a22297a,a22298a,a22301a,a22305a,a22306a,a22307a,a22311a,a22312a,a22316a,a22317a,a22318a,a22321a,a22325a,a22326a,a22327a,a22331a,a22332a,a22336a,a22337a,a22338a,a22341a,a22345a,a22346a,a22347a,a22351a,a22352a,a22356a,a22357a,a22358a,a22361a,a22365a,a22366a,a22367a,a22371a,a22372a,a22376a,a22377a,a22378a,a22381a,a22385a,a22386a,a22387a,a22391a,a22392a,a22396a,a22397a,a22398a,a22401a,a22405a,a22406a,a22407a,a22411a,a22412a,a22416a,a22417a,a22418a,a22421a,a22425a,a22426a,a22427a,a22431a,a22432a,a22436a,a22437a,a22438a,a22441a,a22445a,a22446a,a22447a,a22451a,a22452a,a22456a,a22457a,a22458a,a22461a,a22465a,a22466a,a22467a,a22471a,a22472a,a22476a,a22477a,a22478a,a22482a,a22483a,a22487a,a22488a,a22489a,a22493a,a22494a,a22498a,a22499a,a22500a,a22504a,a22505a,a22509a,a22510a,a22511a,a22515a,a22516a,a22520a,a22521a,a22522a,a22526a,a22527a,a22531a,a22532a,a22533a,a22537a,a22538a,a22542a,a22543a,a22544a,a22548a,a22549a,a22553a,a22554a,a22555a,a22559a,a22560a,a22564a,a22565a,a22566a,a22570a,a22571a,a22575a,a22576a,a22577a,a22581a,a22582a,a22586a,a22587a,a22588a,a22592a,a22593a,a22597a,a22598a,a22599a,a22603a,a22604a,a22608a,a22609a,a22610a,a22614a,a22615a,a22619a,a22620a,a22621a,a22625a,a22626a,a22630a,a22631a,a22632a,a22636a,a22637a,a22641a,a22642a,a22643a,a22647a,a22648a,a22652a,a22653a,a22654a,a22658a,a22659a,a22663a,a22664a,a22665a,a22669a,a22670a,a22674a,a22675a,a22676a,a22680a,a22681a,a22685a,a22686a,a22687a,a22691a,a22692a,a22696a,a22697a,a22698a,a22702a,a22703a,a22707a,a22708a,a22709a,a22713a,a22714a,a22718a,a22719a,a22720a,a22724a,a22725a,a22729a,a22730a,a22731a,a22735a,a22736a,a22740a,a22741a,a22742a,a22746a,a22747a,a22751a,a22752a,a22753a,a22757a,a22758a,a22762a,a22763a,a22764a,a22768a,a22769a,a22773a,a22774a,a22775a,a22779a,a22780a,a22784a,a22785a,a22786a,a22790a,a22791a,a22795a,a22796a,a22797a,a22801a,a22802a,a22806a,a22807a,a22808a,a22812a,a22813a,a22817a,a22818a,a22819a,a22823a,a22824a,a22828a,a22829a,a22830a,a22834a,a22835a,a22839a,a22840a,a22841a,a22845a,a22846a,a22850a,a22851a,a22852a,a22856a,a22857a,a22861a,a22862a,a22863a,a22867a,a22868a,a22872a,a22873a,a22874a,a22878a,a22879a,a22883a,a22884a,a22885a,a22889a,a22890a,a22894a,a22895a,a22896a,a22900a,a22901a,a22905a,a22906a,a22907a,a22911a,a22912a,a22916a,a22917a,a22918a,a22922a,a22923a,a22927a,a22928a,a22929a,a22933a,a22934a,a22938a,a22939a,a22940a,a22944a,a22945a,a22949a,a22950a,a22951a,a22955a,a22956a,a22960a,a22961a,a22962a,a22966a,a22967a,a22971a,a22972a,a22973a,a22977a,a22978a,a22982a,a22983a,a22984a,a22988a,a22989a,a22993a,a22994a,a22995a,a22999a,a23000a,a23004a,a23005a,a23006a,a23010a,a23011a,a23015a,a23016a,a23017a,a23021a,a23022a,a23026a,a23027a,a23028a,a23032a,a23033a,a23037a,a23038a,a23039a,a23043a,a23044a,a23048a,a23049a,a23050a,a23054a,a23055a,a23059a,a23060a,a23061a,a23065a,a23066a,a23070a,a23071a,a23072a,a23076a,a23077a,a23081a,a23082a,a23083a,a23087a,a23088a,a23092a,a23093a,a23094a,a23098a,a23099a,a23103a,a23104a,a23105a,a23109a,a23110a,a23114a,a23115a,a23116a,a23120a,a23121a,a23125a,a23126a,a23127a,a23131a,a23132a,a23136a,a23137a,a23138a,a23142a,a23143a,a23147a,a23148a,a23149a,a23153a,a23154a,a23158a,a23159a,a23160a,a23164a,a23165a,a23169a,a23170a,a23171a,a23175a,a23176a,a23180a,a23181a,a23182a,a23186a,a23187a,a23191a,a23192a,a23193a,a23197a,a23198a,a23202a,a23203a,a23204a,a23208a,a23209a,a23213a,a23214a,a23215a,a23219a,a23220a,a23224a,a23225a,a23226a,a23230a,a23231a,a23235a,a23236a,a23237a,a23241a,a23242a,a23246a,a23247a,a23248a,a23252a,a23253a,a23257a,a23258a,a23259a,a23263a,a23264a,a23268a,a23269a,a23270a,a23274a,a23275a,a23279a,a23280a,a23281a,a23285a,a23286a,a23290a,a23291a,a23292a,a23296a,a23297a,a23301a,a23302a,a23303a,a23307a,a23308a,a23312a,a23313a,a23314a,a23318a,a23319a,a23323a,a23324a,a23325a,a23329a,a23330a,a23334a,a23335a,a23336a,a23340a,a23341a,a23345a,a23346a,a23347a,a23351a,a23352a,a23356a,a23357a,a23358a,a23362a,a23363a,a23367a,a23368a,a23369a,a23373a,a23374a,a23378a,a23379a,a23380a,a23384a,a23385a,a23389a,a23390a,a23391a,a23395a,a23396a,a23400a,a23401a,a23402a,a23406a,a23407a,a23411a,a23412a,a23413a,a23417a,a23418a,a23422a,a23423a,a23424a,a23428a,a23429a,a23433a,a23434a,a23435a,a23439a,a23440a,a23444a,a23445a,a23446a,a23450a,a23451a,a23455a,a23456a,a23457a,a23461a,a23462a,a23466a,a23467a,a23468a,a23472a,a23473a,a23477a,a23478a,a23479a,a23483a,a23484a,a23488a,a23489a,a23490a,a23494a,a23495a,a23499a,a23500a,a23501a,a23505a,a23506a,a23510a,a23511a,a23512a,a23516a,a23517a,a23521a,a23522a,a23523a,a23527a,a23528a,a23532a,a23533a,a23534a,a23538a,a23539a,a23543a,a23544a,a23545a,a23549a,a23550a,a23554a,a23555a,a23556a,a23560a,a23561a,a23565a,a23566a,a23567a,a23571a,a23572a,a23576a,a23577a,a23578a,a23582a,a23583a,a23587a,a23588a,a23589a,a23593a,a23594a,a23598a,a23599a,a23600a,a23604a,a23605a,a23609a,a23610a,a23611a,a23615a,a23616a,a23620a,a23621a,a23622a,a23626a,a23627a,a23631a,a23632a,a23633a,a23637a,a23638a,a23642a,a23643a,a23644a,a23648a,a23649a,a23653a,a23654a,a23655a,a23659a,a23660a,a23664a,a23665a,a23666a,a23670a,a23671a,a23675a,a23676a,a23677a,a23681a,a23682a,a23686a,a23687a,a23688a,a23692a,a23693a,a23697a,a23698a,a23699a,a23703a,a23704a,a23708a,a23709a,a23710a,a23714a,a23715a,a23719a,a23720a,a23721a,a23725a,a23726a,a23730a,a23731a,a23732a,a23736a,a23737a,a23741a,a23742a,a23743a,a23747a,a23748a,a23752a,a23753a,a23754a,a23758a,a23759a,a23763a,a23764a,a23765a,a23769a,a23770a,a23774a,a23775a,a23776a,a23780a,a23781a,a23785a,a23786a,a23787a,a23791a,a23792a,a23796a,a23797a,a23798a,a23802a,a23803a,a23807a,a23808a,a23809a,a23813a,a23814a,a23818a,a23819a,a23820a,a23824a,a23825a,a23829a,a23830a,a23831a,a23835a,a23836a,a23840a,a23841a,a23842a,a23846a,a23847a,a23851a,a23852a,a23853a,a23857a,a23858a,a23862a,a23863a,a23864a,a23868a,a23869a,a23873a,a23874a,a23875a,a23879a,a23880a,a23884a,a23885a,a23886a,a23890a,a23891a,a23895a,a23896a,a23897a,a23901a,a23902a,a23906a,a23907a,a23908a,a23912a,a23913a,a23917a,a23918a,a23919a,a23923a,a23924a,a23928a,a23929a,a23930a,a23934a,a23935a,a23939a,a23940a,a23941a,a23945a,a23946a,a23950a,a23951a,a23952a,a23956a,a23957a,a23961a,a23962a,a23963a,a23967a,a23968a,a23972a,a23973a,a23974a,a23978a,a23979a,a23983a,a23984a,a23985a,a23989a,a23990a,a23994a,a23995a,a23996a,a24000a,a24001a,a24005a,a24006a,a24007a,a24011a,a24012a,a24016a,a24017a,a24018a,a24022a,a24023a,a24027a,a24028a,a24029a,a24033a,a24034a,a24038a,a24039a,a24040a,a24044a,a24045a,a24049a,a24050a,a24051a,a24055a,a24056a,a24060a,a24061a,a24062a,a24066a,a24067a,a24071a,a24072a,a24073a,a24077a,a24078a,a24082a,a24083a,a24084a,a24088a,a24089a,a24093a,a24094a,a24095a,a24099a,a24100a,a24104a,a24105a,a24106a,a24110a,a24111a,a24115a,a24116a,a24117a,a24121a,a24122a,a24126a,a24127a,a24128a,a24132a,a24133a,a24137a,a24138a,a24139a,a24143a,a24144a,a24148a,a24149a,a24150a,a24154a,a24155a,a24159a,a24160a,a24161a,a24165a,a24166a,a24170a,a24171a,a24172a,a24176a,a24177a,a24181a,a24182a,a24183a,a24187a,a24188a,a24192a,a24193a,a24194a,a24198a,a24199a,a24203a,a24204a,a24205a,a24209a,a24210a,a24214a,a24215a,a24216a,a24220a,a24221a,a24225a,a24226a,a24227a,a24231a,a24232a,a24236a,a24237a,a24238a,a24242a,a24243a,a24247a,a24248a,a24249a,a24253a,a24254a,a24258a,a24259a,a24260a,a24264a,a24265a,a24269a,a24270a,a24271a,a24275a,a24276a,a24280a,a24281a,a24282a,a24286a,a24287a,a24291a,a24292a,a24293a,a24297a,a24298a,a24302a,a24303a,a24304a,a24308a,a24309a,a24313a,a24314a,a24315a,a24319a,a24320a,a24324a,a24325a,a24326a,a24330a,a24331a,a24335a,a24336a,a24337a,a24341a,a24342a,a24346a,a24347a,a24348a,a24352a,a24353a,a24357a,a24358a,a24359a,a24363a,a24364a,a24368a,a24369a,a24370a,a24374a,a24375a,a24379a,a24380a,a24381a,a24385a,a24386a,a24390a,a24391a,a24392a,a24396a,a24397a,a24401a,a24402a,a24403a,a24407a,a24408a,a24412a,a24413a,a24414a,a24418a,a24419a,a24423a,a24424a,a24425a,a24429a,a24430a,a24434a,a24435a,a24436a,a24440a,a24441a,a24445a,a24446a,a24447a,a24451a,a24452a,a24456a,a24457a,a24458a,a24462a,a24463a,a24467a,a24468a,a24469a,a24473a,a24474a,a24478a,a24479a,a24480a,a24484a,a24485a,a24489a,a24490a,a24491a,a24495a,a24496a,a24500a,a24501a,a24502a,a24506a,a24507a,a24511a,a24512a,a24513a,a24517a,a24518a,a24522a,a24523a,a24524a,a24528a,a24529a,a24533a,a24534a,a24535a,a24539a,a24540a,a24544a,a24545a,a24546a,a24550a,a24551a,a24555a,a24556a,a24557a,a24561a,a24562a,a24566a,a24567a,a24568a,a24572a,a24573a,a24577a,a24578a,a24579a,a24583a,a24584a,a24588a,a24589a,a24590a,a24594a,a24595a,a24599a,a24600a,a24601a,a24605a,a24606a,a24610a,a24611a,a24612a,a24616a,a24617a,a24621a,a24622a,a24623a,a24627a,a24628a,a24632a,a24633a,a24634a,a24638a,a24639a,a24643a,a24644a,a24645a,a24649a,a24650a,a24654a,a24655a,a24656a,a24660a,a24661a,a24665a,a24666a,a24667a,a24671a,a24672a,a24676a,a24677a,a24678a,a24682a,a24683a,a24687a,a24688a,a24689a,a24693a,a24694a,a24698a,a24699a,a24700a,a24704a,a24705a,a24709a,a24710a,a24711a,a24715a,a24716a,a24720a,a24721a,a24722a,a24726a,a24727a,a24731a,a24732a,a24733a,a24737a,a24738a,a24742a,a24743a,a24744a,a24748a,a24749a,a24753a,a24754a,a24755a,a24759a,a24760a,a24764a,a24765a,a24766a,a24770a,a24771a,a24775a,a24776a,a24777a,a24781a,a24782a,a24786a,a24787a,a24788a,a24792a,a24793a,a24797a,a24798a,a24799a,a24803a,a24804a,a24808a,a24809a,a24810a,a24814a,a24815a,a24819a,a24820a,a24821a,a24825a,a24826a,a24830a,a24831a,a24832a,a24836a,a24837a,a24841a,a24842a,a24843a,a24847a,a24848a,a24852a,a24853a,a24854a,a24858a,a24859a,a24863a,a24864a,a24865a,a24869a,a24870a,a24874a,a24875a,a24876a,a24880a,a24881a,a24885a,a24886a,a24887a,a24891a,a24892a,a24896a,a24897a,a24898a,a24902a,a24903a,a24907a,a24908a,a24909a,a24913a,a24914a,a24918a,a24919a,a24920a,a24924a,a24925a,a24929a,a24930a,a24931a,a24935a,a24936a,a24940a,a24941a,a24942a,a24946a,a24947a,a24951a,a24952a,a24953a,a24957a,a24958a,a24962a,a24963a,a24964a,a24968a,a24969a,a24973a,a24974a,a24975a,a24979a,a24980a,a24984a,a24985a,a24986a,a24990a,a24991a,a24995a,a24996a,a24997a,a25001a,a25002a,a25006a,a25007a,a25008a,a25012a,a25013a,a25017a,a25018a,a25019a,a25023a,a25024a,a25028a,a25029a,a25030a,a25034a,a25035a,a25039a,a25040a,a25041a,a25045a,a25046a,a25050a,a25051a,a25052a,a25056a,a25057a,a25061a,a25062a,a25063a,a25067a,a25068a,a25072a,a25073a,a25074a,a25078a,a25079a,a25083a,a25084a,a25085a,a25089a,a25090a,a25094a,a25095a,a25096a,a25100a,a25101a,a25105a,a25106a,a25107a,a25111a,a25112a,a25116a,a25117a,a25118a,a25122a,a25123a,a25127a,a25128a,a25129a,a25133a,a25134a,a25138a,a25139a,a25140a,a25144a,a25145a,a25149a,a25150a,a25151a,a25155a,a25156a,a25160a,a25161a,a25162a,a25166a,a25167a,a25171a,a25172a,a25173a,a25177a,a25178a,a25182a,a25183a,a25184a,a25188a,a25189a,a25193a,a25194a,a25195a,a25199a,a25200a,a25204a,a25205a,a25206a,a25210a,a25211a,a25215a,a25216a,a25217a,a25221a,a25222a,a25226a,a25227a,a25228a,a25232a,a25233a,a25237a,a25238a,a25239a,a25243a,a25244a,a25248a,a25249a,a25250a,a25254a,a25255a,a25259a,a25260a,a25261a,a25265a,a25266a,a25270a,a25271a,a25272a,a25276a,a25277a,a25281a,a25282a,a25283a,a25287a,a25288a,a25292a,a25293a,a25294a,a25298a,a25299a,a25303a,a25304a,a25305a,a25309a,a25310a,a25314a,a25315a,a25316a,a25320a,a25321a,a25325a,a25326a,a25327a,a25331a,a25332a,a25336a,a25337a,a25338a,a25342a,a25343a,a25347a,a25348a,a25349a,a25353a,a25354a,a25358a,a25359a,a25360a,a25364a,a25365a,a25369a,a25370a,a25371a,a25375a,a25376a,a25380a,a25381a,a25382a,a25386a,a25387a,a25391a,a25392a,a25393a,a25397a,a25398a,a25402a,a25403a,a25404a,a25408a,a25409a,a25413a,a25414a,a25415a,a25419a,a25420a,a25424a,a25425a,a25426a,a25430a,a25431a,a25435a,a25436a,a25437a,a25441a,a25442a,a25446a,a25447a,a25448a,a25452a,a25453a,a25457a,a25458a,a25459a,a25463a,a25464a,a25468a,a25469a,a25470a,a25474a,a25475a,a25479a,a25480a,a25481a,a25485a,a25486a,a25490a,a25491a,a25492a,a25496a,a25497a,a25501a,a25502a,a25503a,a25507a,a25508a,a25512a,a25513a,a25514a,a25518a,a25519a,a25523a,a25524a,a25525a,a25529a,a25530a,a25534a,a25535a,a25536a,a25540a,a25541a,a25545a,a25546a,a25547a,a25551a,a25552a,a25556a,a25557a,a25558a,a25562a,a25563a,a25567a,a25568a,a25569a,a25573a,a25574a,a25578a,a25579a,a25580a,a25584a,a25585a,a25589a,a25590a,a25591a,a25595a,a25596a,a25600a,a25601a,a25602a,a25606a,a25607a,a25611a,a25612a,a25613a,a25617a,a25618a,a25622a,a25623a,a25624a,a25628a,a25629a,a25633a,a25634a,a25635a,a25639a,a25640a,a25644a,a25645a,a25646a,a25650a,a25651a,a25655a,a25656a,a25657a,a25661a,a25662a,a25666a,a25667a,a25668a,a25672a,a25673a,a25677a,a25678a,a25679a,a25683a,a25684a,a25688a,a25689a,a25690a,a25694a,a25695a,a25699a,a25700a,a25701a,a25705a,a25706a,a25710a,a25711a,a25712a,a25716a,a25717a,a25721a,a25722a,a25723a,a25727a,a25728a,a25732a,a25733a,a25734a,a25738a,a25739a,a25743a,a25744a,a25745a,a25749a,a25750a,a25754a,a25755a,a25756a,a25760a,a25761a,a25765a,a25766a,a25767a,a25771a,a25772a,a25776a,a25777a,a25778a,a25782a,a25783a,a25787a,a25788a,a25789a,a25793a,a25794a,a25798a,a25799a,a25800a,a25804a,a25805a,a25809a,a25810a,a25811a,a25815a,a25816a,a25820a,a25821a,a25822a,a25826a,a25827a,a25831a,a25832a,a25833a,a25837a,a25838a,a25842a,a25843a,a25844a,a25848a,a25849a,a25853a,a25854a,a25855a,a25859a,a25860a,a25864a,a25865a,a25866a,a25870a,a25871a,a25875a,a25876a,a25877a,a25881a,a25882a,a25886a,a25887a,a25888a,a25892a,a25893a,a25897a,a25898a,a25899a,a25903a,a25904a,a25908a,a25909a,a25910a,a25914a,a25915a,a25919a,a25920a,a25921a,a25925a,a25926a,a25930a,a25931a,a25932a,a25936a,a25937a,a25941a,a25942a,a25943a,a25947a,a25948a,a25952a,a25953a,a25954a,a25958a,a25959a,a25963a,a25964a,a25965a,a25969a,a25970a,a25974a,a25975a,a25976a,a25980a,a25981a,a25985a,a25986a,a25987a,a25991a,a25992a,a25996a,a25997a,a25998a,a26002a,a26003a,a26007a,a26008a,a26009a,a26013a,a26014a,a26018a,a26019a,a26020a,a26024a,a26025a,a26029a,a26030a,a26031a,a26035a,a26036a,a26040a,a26041a,a26042a,a26046a,a26047a,a26051a,a26052a,a26053a,a26057a,a26058a,a26062a,a26063a,a26064a,a26068a,a26069a,a26073a,a26074a,a26075a,a26079a,a26080a,a26084a,a26085a,a26086a,a26090a,a26091a,a26095a,a26096a,a26097a,a26101a,a26102a,a26106a,a26107a,a26108a,a26112a,a26113a,a26117a,a26118a,a26119a,a26123a,a26124a,a26128a,a26129a,a26130a,a26134a,a26135a,a26139a,a26140a,a26141a,a26145a,a26146a,a26150a,a26151a,a26152a,a26156a,a26157a,a26161a,a26162a,a26163a,a26167a,a26168a,a26172a,a26173a,a26174a,a26178a,a26179a,a26183a,a26184a,a26185a,a26189a,a26190a,a26194a,a26195a,a26196a,a26200a,a26201a,a26205a,a26206a,a26207a,a26211a,a26212a,a26216a,a26217a,a26218a,a26222a,a26223a,a26227a,a26228a,a26229a,a26233a,a26234a,a26238a,a26239a,a26240a,a26244a,a26245a,a26249a,a26250a,a26251a,a26255a,a26256a,a26260a,a26261a,a26262a,a26266a,a26267a,a26271a,a26272a,a26273a,a26277a,a26278a,a26282a,a26283a,a26284a,a26288a,a26289a,a26293a,a26294a,a26295a,a26299a,a26300a,a26304a,a26305a,a26306a,a26310a,a26311a,a26315a,a26316a,a26317a,a26321a,a26322a,a26326a,a26327a,a26328a,a26332a,a26333a,a26337a,a26338a,a26339a,a26343a,a26344a,a26348a,a26349a,a26350a,a26354a,a26355a,a26359a,a26360a,a26361a,a26365a,a26366a,a26370a,a26371a,a26372a,a26376a,a26377a,a26381a,a26382a,a26383a,a26387a,a26388a,a26392a,a26393a,a26394a,a26398a,a26399a,a26403a,a26404a,a26405a,a26409a,a26410a,a26414a,a26415a,a26416a,a26420a,a26421a,a26425a,a26426a,a26427a,a26431a,a26432a,a26436a,a26437a,a26438a,a26442a,a26443a,a26447a,a26448a,a26449a,a26453a,a26454a,a26458a,a26459a,a26460a,a26464a,a26465a,a26469a,a26470a,a26471a,a26475a,a26476a,a26480a,a26481a,a26482a,a26486a,a26487a,a26491a,a26492a,a26493a,a26497a,a26498a,a26502a,a26503a,a26504a,a26508a,a26509a,a26513a,a26514a,a26515a,a26519a,a26520a,a26524a,a26525a,a26526a,a26530a,a26531a,a26535a,a26536a,a26537a,a26541a,a26542a,a26546a,a26547a,a26548a,a26552a,a26553a,a26557a,a26558a,a26559a,a26563a,a26564a,a26568a,a26569a,a26570a,a26574a,a26575a,a26579a,a26580a,a26581a,a26585a,a26586a,a26590a,a26591a,a26592a,a26596a,a26597a,a26601a,a26602a,a26603a,a26607a,a26608a,a26612a,a26613a,a26614a,a26618a,a26619a,a26623a,a26624a,a26625a,a26629a,a26630a,a26634a,a26635a,a26636a,a26640a,a26641a,a26645a,a26646a,a26647a,a26651a,a26652a,a26656a,a26657a,a26658a,a26662a,a26663a,a26667a,a26668a,a26669a,a26673a,a26674a,a26678a,a26679a,a26680a,a26684a,a26685a,a26689a,a26690a,a26691a,a26695a,a26696a,a26700a,a26701a,a26702a,a26706a,a26707a,a26711a,a26712a,a26713a,a26717a,a26718a,a26722a,a26723a,a26724a,a26728a,a26729a,a26733a,a26734a,a26735a,a26739a,a26740a,a26744a,a26745a,a26746a,a26750a,a26751a,a26755a,a26756a,a26757a,a26761a,a26762a,a26766a,a26767a,a26768a,a26772a,a26773a,a26777a,a26778a,a26779a,a26783a,a26784a,a26788a,a26789a,a26790a,a26794a,a26795a,a26799a,a26800a,a26801a,a26805a,a26806a,a26810a,a26811a,a26812a,a26816a,a26817a,a26821a,a26822a,a26823a,a26827a,a26828a,a26832a,a26833a,a26834a,a26838a,a26839a,a26843a,a26844a,a26845a,a26849a,a26850a,a26854a,a26855a,a26856a,a26860a,a26861a,a26865a,a26866a,a26867a,a26871a,a26872a,a26876a,a26877a,a26878a,a26882a,a26883a,a26887a,a26888a,a26889a,a26893a,a26894a,a26898a,a26899a,a26900a,a26904a,a26905a,a26909a,a26910a,a26911a,a26915a,a26916a,a26920a,a26921a,a26922a,a26926a,a26927a,a26931a,a26932a,a26933a,a26937a,a26938a,a26942a,a26943a,a26944a,a26948a,a26949a,a26953a,a26954a,a26955a,a26959a,a26960a,a26964a,a26965a,a26966a,a26970a,a26971a,a26975a,a26976a,a26977a,a26981a,a26982a,a26986a,a26987a,a26988a,a26992a,a26993a,a26997a,a26998a,a26999a,a27003a,a27004a,a27008a,a27009a,a27010a,a27014a,a27015a,a27019a,a27020a,a27021a,a27025a,a27026a,a27030a,a27031a,a27032a,a27036a,a27037a,a27041a,a27042a,a27043a,a27047a,a27048a,a27052a,a27053a,a27054a,a27058a,a27059a,a27063a,a27064a,a27065a,a27069a,a27070a,a27074a,a27075a,a27076a,a27080a,a27081a,a27085a,a27086a,a27087a,a27091a,a27092a,a27096a,a27097a,a27098a,a27102a,a27103a,a27107a,a27108a,a27109a,a27113a,a27114a,a27118a,a27119a,a27120a,a27124a,a27125a,a27129a,a27130a,a27131a,a27135a,a27136a,a27140a,a27141a,a27142a,a27146a,a27147a,a27151a,a27152a,a27153a,a27157a,a27158a,a27162a,a27163a,a27164a,a27168a,a27169a,a27173a,a27174a,a27175a,a27179a,a27180a,a27184a,a27185a,a27186a,a27190a,a27191a,a27195a,a27196a,a27197a,a27201a,a27202a,a27206a,a27207a,a27208a,a27212a,a27213a,a27217a,a27218a,a27219a,a27223a,a27224a,a27228a,a27229a,a27230a,a27234a,a27235a,a27239a,a27240a,a27241a,a27245a,a27246a,a27250a,a27251a,a27252a,a27256a,a27257a,a27261a,a27262a,a27263a,a27267a,a27268a,a27272a,a27273a,a27274a,a27278a,a27279a,a27283a,a27284a,a27285a,a27289a,a27290a,a27294a,a27295a,a27296a,a27300a,a27301a,a27305a,a27306a,a27307a,a27311a,a27312a,a27316a,a27317a,a27318a,a27322a,a27323a,a27327a,a27328a,a27329a,a27333a,a27334a,a27338a,a27339a,a27340a,a27344a,a27345a,a27349a,a27350a,a27351a,a27355a,a27356a,a27360a,a27361a,a27362a,a27366a,a27367a,a27371a,a27372a,a27373a,a27377a,a27378a,a27382a,a27383a,a27384a,a27388a,a27389a,a27393a,a27394a,a27395a,a27399a,a27400a,a27404a,a27405a,a27406a,a27410a,a27411a,a27415a,a27416a,a27417a,a27421a,a27422a,a27426a,a27427a,a27428a,a27432a,a27433a,a27437a,a27438a,a27439a,a27443a,a27444a,a27448a,a27449a,a27450a,a27454a,a27455a,a27459a,a27460a,a27461a,a27465a,a27466a,a27470a,a27471a,a27472a,a27476a,a27477a,a27481a,a27482a,a27483a,a27487a,a27488a,a27492a,a27493a,a27494a,a27498a,a27499a,a27503a,a27504a,a27505a,a27509a,a27510a,a27514a,a27515a,a27516a,a27520a,a27521a,a27525a,a27526a,a27527a,a27531a,a27532a,a27536a,a27537a,a27538a,a27542a,a27543a,a27547a,a27548a,a27549a,a27553a,a27554a,a27558a,a27559a,a27560a,a27564a,a27565a,a27569a,a27570a,a27571a,a27575a,a27576a,a27580a,a27581a,a27582a,a27586a,a27587a,a27591a,a27592a,a27593a,a27597a,a27598a,a27602a,a27603a,a27604a,a27608a,a27609a,a27613a,a27614a,a27615a,a27619a,a27620a,a27624a,a27625a,a27626a,a27630a,a27631a,a27635a,a27636a,a27637a,a27641a,a27642a,a27646a,a27647a,a27648a,a27652a,a27653a,a27657a,a27658a,a27659a,a27663a,a27664a,a27668a,a27669a,a27670a,a27674a,a27675a,a27679a,a27680a,a27681a,a27685a,a27686a,a27690a,a27691a,a27692a,a27696a,a27697a,a27701a,a27702a,a27703a,a27707a,a27708a,a27712a,a27713a,a27714a,a27718a,a27719a,a27723a,a27724a,a27725a,a27729a,a27730a,a27734a,a27735a,a27736a,a27740a,a27741a,a27745a,a27746a,a27747a,a27751a,a27752a,a27756a,a27757a,a27758a,a27762a,a27763a,a27767a,a27768a,a27769a,a27773a,a27774a,a27778a,a27779a,a27780a,a27784a,a27785a,a27789a,a27790a,a27791a,a27795a,a27796a,a27800a,a27801a,a27802a,a27806a,a27807a,a27811a,a27812a,a27813a,a27817a,a27818a,a27822a,a27823a,a27824a,a27828a,a27829a,a27833a,a27834a,a27835a,a27839a,a27840a,a27844a,a27845a,a27846a,a27850a,a27851a,a27855a,a27856a,a27857a,a27861a,a27862a,a27866a,a27867a,a27868a,a27872a,a27873a,a27877a,a27878a,a27879a,a27883a,a27884a,a27888a,a27889a,a27890a,a27894a,a27895a,a27899a,a27900a,a27901a,a27905a,a27906a,a27910a,a27911a,a27912a,a27916a,a27917a,a27921a,a27922a,a27923a,a27927a,a27928a,a27932a,a27933a,a27934a,a27938a,a27939a,a27943a,a27944a,a27945a,a27949a,a27950a,a27954a,a27955a,a27956a,a27960a,a27961a,a27965a,a27966a,a27967a,a27971a,a27972a,a27976a,a27977a,a27978a,a27982a,a27983a,a27987a,a27988a,a27989a,a27993a,a27994a,a27998a,a27999a,a28000a,a28004a,a28005a,a28009a,a28010a,a28011a,a28015a,a28016a,a28020a,a28021a,a28022a,a28026a,a28027a,a28031a,a28032a,a28033a,a28037a,a28038a,a28042a,a28043a,a28044a,a28048a,a28049a,a28053a,a28054a,a28055a,a28059a,a28060a,a28064a,a28065a,a28066a,a28070a,a28071a,a28075a,a28076a,a28077a,a28081a,a28082a,a28086a,a28087a,a28088a,a28092a,a28093a,a28097a,a28098a,a28099a,a28103a,a28104a,a28108a,a28109a,a28110a,a28114a,a28115a,a28119a,a28120a,a28121a,a28125a,a28126a,a28130a,a28131a,a28132a,a28136a,a28137a,a28141a,a28142a,a28143a,a28147a,a28148a,a28152a,a28153a,a28154a,a28158a,a28159a,a28163a,a28164a,a28165a,a28169a,a28170a,a28174a,a28175a,a28176a,a28180a,a28181a,a28185a,a28186a,a28187a,a28191a,a28192a,a28196a,a28197a,a28198a,a28202a,a28203a,a28207a,a28208a,a28209a,a28213a,a28214a,a28218a,a28219a,a28220a,a28224a,a28225a,a28229a,a28230a,a28231a,a28235a,a28236a,a28240a,a28241a,a28242a,a28246a,a28247a,a28251a,a28252a,a28253a,a28257a,a28258a,a28262a,a28263a,a28264a,a28268a,a28269a,a28273a,a28274a,a28275a,a28279a,a28280a,a28284a,a28285a,a28286a,a28290a,a28291a,a28295a,a28296a,a28297a,a28301a,a28302a,a28306a,a28307a,a28308a,a28312a,a28313a,a28317a,a28318a,a28319a,a28323a,a28324a,a28328a,a28329a,a28330a,a28334a,a28335a,a28339a,a28340a,a28341a,a28345a,a28346a,a28350a,a28351a,a28352a,a28356a,a28357a,a28361a,a28362a,a28363a,a28367a,a28368a,a28372a,a28373a,a28374a,a28378a,a28379a,a28383a,a28384a,a28385a,a28389a,a28390a,a28394a,a28395a,a28396a,a28400a,a28401a,a28405a,a28406a,a28407a,a28411a,a28412a,a28416a,a28417a,a28418a,a28422a,a28423a,a28427a,a28428a,a28429a,a28433a,a28434a,a28438a,a28439a,a28440a,a28444a,a28445a,a28449a,a28450a,a28451a,a28455a,a28456a,a28460a,a28461a,a28462a,a28466a,a28467a,a28471a,a28472a,a28473a,a28477a,a28478a,a28482a,a28483a,a28484a,a28488a,a28489a,a28493a,a28494a,a28495a,a28499a,a28500a,a28504a,a28505a,a28506a,a28510a,a28511a,a28515a,a28516a,a28517a,a28521a,a28522a,a28526a,a28527a,a28528a,a28532a,a28533a,a28537a,a28538a,a28539a,a28543a,a28544a,a28548a,a28549a,a28550a,a28554a,a28555a,a28559a,a28560a,a28561a,a28565a,a28566a,a28570a,a28571a,a28572a,a28576a,a28577a,a28581a,a28582a,a28583a,a28587a,a28588a,a28592a,a28593a,a28594a,a28598a,a28599a,a28603a,a28604a,a28605a,a28609a,a28610a,a28614a,a28615a,a28616a,a28620a,a28621a,a28625a,a28626a,a28627a,a28631a,a28632a,a28636a,a28637a,a28638a,a28642a,a28643a,a28647a,a28648a,a28649a,a28653a,a28654a,a28658a,a28659a,a28660a,a28664a,a28665a,a28669a,a28670a,a28671a,a28675a,a28676a,a28680a,a28681a,a28682a,a28686a,a28687a,a28691a,a28692a,a28693a,a28697a,a28698a,a28702a,a28703a,a28704a,a28708a,a28709a,a28713a,a28714a,a28715a,a28719a,a28720a,a28724a,a28725a,a28726a,a28730a,a28731a,a28735a,a28736a,a28737a,a28741a,a28742a,a28746a,a28747a,a28748a,a28752a,a28753a,a28757a,a28758a,a28759a,a28763a,a28764a,a28768a,a28769a,a28770a,a28774a,a28775a,a28779a,a28780a,a28781a,a28785a,a28786a,a28790a,a28791a,a28792a,a28796a,a28797a,a28801a,a28802a,a28803a,a28807a,a28808a,a28812a,a28813a,a28814a,a28818a,a28819a,a28823a,a28824a,a28825a,a28829a,a28830a,a28834a,a28835a,a28836a,a28840a,a28841a,a28845a,a28846a,a28847a,a28851a,a28852a,a28856a,a28857a,a28858a,a28862a,a28863a,a28867a,a28868a,a28869a,a28873a,a28874a,a28878a,a28879a,a28880a,a28884a,a28885a,a28889a,a28890a,a28891a,a28895a,a28896a,a28900a,a28901a,a28902a,a28906a,a28907a,a28911a,a28912a,a28913a,a28917a,a28918a,a28922a,a28923a,a28924a,a28928a,a28929a,a28933a,a28934a,a28935a,a28939a,a28940a,a28944a,a28945a,a28946a,a28950a,a28951a,a28955a,a28956a,a28957a,a28961a,a28962a,a28966a,a28967a,a28968a,a28972a,a28973a,a28977a,a28978a,a28979a,a28983a,a28984a,a28988a,a28989a,a28990a,a28994a,a28995a,a28999a,a29000a,a29001a,a29005a,a29006a,a29010a,a29011a,a29012a,a29016a,a29017a,a29021a,a29022a,a29023a,a29027a,a29028a,a29032a,a29033a,a29034a,a29038a,a29039a,a29043a,a29044a,a29045a,a29049a,a29050a,a29054a,a29055a,a29056a,a29060a,a29061a,a29065a,a29066a,a29067a,a29071a,a29072a,a29076a,a29077a,a29078a,a29082a,a29083a,a29087a,a29088a,a29089a,a29093a,a29094a,a29098a,a29099a,a29100a,a29104a,a29105a,a29109a,a29110a,a29111a,a29115a,a29116a,a29120a,a29121a,a29122a,a29126a,a29127a,a29131a,a29132a,a29133a,a29137a,a29138a,a29142a,a29143a,a29144a,a29148a,a29149a,a29153a,a29154a,a29155a,a29159a,a29160a,a29164a,a29165a,a29166a,a29170a,a29171a,a29175a,a29176a,a29177a,a29181a,a29182a,a29186a,a29187a,a29188a,a29192a,a29193a,a29197a,a29198a,a29199a,a29203a,a29204a,a29208a,a29209a,a29210a,a29214a,a29215a,a29219a,a29220a,a29221a,a29225a,a29226a,a29230a,a29231a,a29232a,a29236a,a29237a,a29241a,a29242a,a29243a,a29247a,a29248a,a29252a,a29253a,a29254a,a29258a,a29259a,a29263a,a29264a,a29265a,a29269a,a29270a,a29274a,a29275a,a29276a,a29280a,a29281a,a29285a,a29286a,a29287a,a29291a,a29292a,a29296a,a29297a,a29298a,a29302a,a29303a,a29307a,a29308a,a29309a,a29313a,a29314a,a29318a,a29319a,a29320a,a29324a,a29325a,a29329a,a29330a,a29331a,a29335a,a29336a,a29340a,a29341a,a29342a,a29346a,a29347a,a29351a,a29352a,a29353a,a29357a,a29358a,a29362a,a29363a,a29364a,a29368a,a29369a,a29373a,a29374a,a29375a,a29379a,a29380a,a29384a,a29385a,a29386a,a29390a,a29391a,a29395a,a29396a,a29397a,a29401a,a29402a,a29406a,a29407a,a29408a,a29412a,a29413a,a29417a,a29418a,a29419a,a29423a,a29424a,a29428a,a29429a,a29430a,a29434a,a29435a,a29439a,a29440a,a29441a,a29445a,a29446a,a29450a,a29451a,a29452a,a29456a,a29457a,a29461a,a29462a,a29463a,a29467a,a29468a,a29472a,a29473a,a29474a,a29478a,a29479a,a29483a,a29484a,a29485a,a29489a,a29490a,a29494a,a29495a,a29496a,a29500a,a29501a,a29505a,a29506a,a29507a,a29511a,a29512a,a29516a,a29517a,a29518a,a29522a,a29523a,a29527a,a29528a,a29529a,a29533a,a29534a,a29538a,a29539a,a29540a,a29544a,a29545a,a29549a,a29550a,a29551a,a29555a,a29556a,a29560a,a29561a,a29562a,a29566a,a29567a,a29571a,a29572a,a29573a,a29577a,a29578a,a29582a,a29583a,a29584a,a29588a,a29589a,a29593a,a29594a,a29595a,a29599a,a29600a,a29604a,a29605a,a29606a,a29610a,a29611a,a29615a,a29616a,a29617a,a29621a,a29622a,a29626a,a29627a,a29628a,a29632a,a29633a,a29637a,a29638a,a29639a,a29643a,a29644a,a29648a,a29649a,a29650a,a29654a,a29655a,a29659a,a29660a,a29661a,a29665a,a29666a,a29670a,a29671a,a29672a,a29676a,a29677a,a29681a,a29682a,a29683a,a29687a,a29688a,a29692a,a29693a,a29694a,a29698a,a29699a,a29703a,a29704a,a29705a,a29709a,a29710a,a29714a,a29715a,a29716a,a29720a,a29721a,a29725a,a29726a,a29727a,a29731a,a29732a,a29736a,a29737a,a29738a,a29742a,a29743a,a29747a,a29748a,a29749a,a29753a,a29754a,a29758a,a29759a,a29760a,a29764a,a29765a,a29769a,a29770a,a29771a,a29775a,a29776a,a29780a,a29781a,a29782a,a29786a,a29787a,a29791a,a29792a,a29793a,a29797a,a29798a,a29802a,a29803a,a29804a,a29808a,a29809a,a29813a,a29814a,a29815a,a29819a,a29820a,a29824a,a29825a,a29826a,a29830a,a29831a,a29835a,a29836a,a29837a,a29841a,a29842a,a29846a,a29847a,a29848a,a29852a,a29853a,a29857a,a29858a,a29859a,a29863a,a29864a,a29868a,a29869a,a29870a,a29874a,a29875a,a29879a,a29880a,a29881a,a29885a,a29886a,a29890a,a29891a,a29892a,a29896a,a29897a,a29901a,a29902a,a29903a,a29907a,a29908a,a29912a,a29913a,a29914a,a29918a,a29919a,a29923a,a29924a,a29925a,a29929a,a29930a,a29934a,a29935a,a29936a,a29940a,a29941a,a29945a,a29946a,a29947a,a29951a,a29952a,a29956a,a29957a,a29958a,a29962a,a29963a,a29967a,a29968a,a29969a,a29973a,a29974a,a29978a,a29979a,a29980a,a29984a,a29985a,a29989a,a29990a,a29991a,a29995a,a29996a,a30000a,a30001a,a30002a,a30006a,a30007a,a30011a,a30012a,a30013a,a30017a,a30018a,a30022a,a30023a,a30024a,a30028a,a30029a,a30033a,a30034a,a30035a,a30039a,a30040a,a30044a,a30045a,a30046a,a30050a,a30051a,a30055a,a30056a,a30057a,a30061a,a30062a,a30066a,a30067a,a30068a,a30072a,a30073a,a30077a,a30078a,a30079a,a30083a,a30084a,a30088a,a30089a,a30090a,a30094a,a30095a,a30099a,a30100a,a30101a,a30105a,a30106a,a30110a,a30111a,a30112a,a30116a,a30117a,a30121a,a30122a,a30123a,a30127a,a30128a,a30132a,a30133a,a30134a,a30138a,a30139a,a30143a,a30144a,a30145a,a30149a,a30150a,a30154a,a30155a,a30156a,a30160a,a30161a,a30165a,a30166a,a30167a,a30171a,a30172a,a30176a,a30177a,a30178a,a30182a,a30183a,a30187a,a30188a,a30189a,a30193a,a30194a,a30198a,a30199a,a30200a,a30204a,a30205a,a30209a,a30210a,a30211a,a30215a,a30216a,a30220a,a30221a,a30222a,a30226a,a30227a,a30231a,a30232a,a30233a,a30237a,a30238a,a30242a,a30243a,a30244a,a30248a,a30249a,a30253a,a30254a,a30255a,a30259a,a30260a,a30264a,a30265a,a30266a,a30270a,a30271a,a30275a,a30276a,a30277a,a30281a,a30282a,a30286a,a30287a,a30288a,a30292a,a30293a,a30297a,a30298a,a30299a,a30303a,a30304a,a30308a,a30309a,a30310a,a30314a,a30315a,a30319a,a30320a,a30321a,a30325a,a30326a,a30330a,a30331a,a30332a,a30336a,a30337a,a30341a,a30342a,a30343a,a30347a,a30348a,a30352a,a30353a,a30354a,a30358a,a30359a,a30363a,a30364a,a30365a,a30369a,a30370a,a30374a,a30375a,a30376a,a30380a,a30381a,a30385a,a30386a,a30387a,a30391a,a30392a,a30396a,a30397a,a30398a,a30402a,a30403a,a30407a,a30408a,a30409a,a30413a,a30414a,a30418a,a30419a,a30420a,a30424a,a30425a,a30429a,a30430a,a30431a,a30435a,a30436a,a30440a,a30441a,a30442a,a30446a,a30447a,a30451a,a30452a,a30453a,a30457a,a30458a,a30462a,a30463a,a30464a,a30468a,a30469a,a30473a,a30474a,a30475a,a30479a,a30480a,a30484a,a30485a,a30486a,a30490a,a30491a,a30495a,a30496a,a30497a,a30501a,a30502a,a30506a,a30507a,a30508a,a30512a,a30513a,a30517a,a30518a,a30519a,a30523a,a30524a,a30528a,a30529a,a30530a,a30534a,a30535a,a30539a,a30540a,a30541a,a30545a,a30546a,a30550a,a30551a,a30552a,a30556a,a30557a,a30561a,a30562a,a30563a,a30567a,a30568a,a30572a,a30573a,a30574a,a30578a,a30579a,a30583a,a30584a,a30585a,a30589a,a30590a,a30594a,a30595a,a30596a,a30600a,a30601a,a30605a,a30606a,a30607a,a30611a,a30612a,a30616a,a30617a,a30618a,a30622a,a30623a,a30627a,a30628a,a30629a,a30633a,a30634a,a30638a,a30639a,a30640a,a30644a,a30645a,a30649a,a30650a,a30651a,a30655a,a30656a,a30660a,a30661a,a30662a,a30666a,a30667a,a30671a,a30672a,a30673a,a30677a,a30678a,a30682a,a30683a,a30684a,a30688a,a30689a,a30693a,a30694a,a30695a,a30699a,a30700a,a30704a,a30705a,a30706a,a30710a,a30711a,a30715a,a30716a,a30717a,a30721a,a30722a,a30726a,a30727a,a30728a,a30732a,a30733a,a30737a,a30738a,a30739a,a30743a,a30744a,a30748a,a30749a,a30750a,a30754a,a30755a,a30759a,a30760a,a30761a,a30765a,a30766a,a30770a,a30771a,a30772a,a30776a,a30777a,a30781a,a30782a,a30783a,a30787a,a30788a,a30792a,a30793a,a30794a,a30798a,a30799a,a30803a,a30804a,a30805a,a30809a,a30810a,a30814a,a30815a,a30816a,a30820a,a30821a,a30825a,a30826a,a30827a,a30831a,a30832a,a30836a,a30837a,a30838a,a30842a,a30843a,a30847a,a30848a,a30849a,a30853a,a30854a,a30858a,a30859a,a30860a,a30864a,a30865a,a30869a,a30870a,a30871a,a30875a,a30876a,a30880a,a30881a,a30882a,a30886a,a30887a,a30891a,a30892a,a30893a,a30897a,a30898a,a30902a,a30903a,a30904a,a30908a,a30909a,a30913a,a30914a,a30915a,a30919a,a30920a,a30924a,a30925a,a30926a,a30930a,a30931a,a30935a,a30936a,a30937a,a30941a,a30942a,a30946a,a30947a,a30948a,a30952a,a30953a,a30957a,a30958a,a30959a,a30963a,a30964a,a30968a,a30969a,a30970a,a30974a,a30975a,a30979a,a30980a,a30981a,a30985a,a30986a,a30990a,a30991a,a30992a,a30996a,a30997a,a31001a,a31002a,a31003a,a31007a,a31008a,a31012a,a31013a,a31014a,a31018a,a31019a,a31023a,a31024a,a31025a,a31029a,a31030a,a31034a,a31035a,a31036a,a31040a,a31041a,a31045a,a31046a,a31047a,a31051a,a31052a,a31056a,a31057a,a31058a,a31062a,a31063a,a31067a,a31068a,a31069a,a31073a,a31074a,a31078a,a31079a,a31080a,a31084a,a31085a,a31089a,a31090a,a31091a,a31095a,a31096a,a31100a,a31101a,a31102a,a31106a,a31107a,a31111a,a31112a,a31113a,a31117a,a31118a,a31122a,a31123a,a31124a,a31128a,a31129a,a31133a,a31134a,a31135a,a31139a,a31140a,a31144a,a31145a,a31146a,a31150a,a31151a,a31155a,a31156a,a31157a,a31161a,a31162a,a31166a,a31167a,a31168a,a31172a,a31173a,a31177a,a31178a,a31179a,a31183a,a31184a,a31188a,a31189a,a31190a,a31194a,a31195a,a31199a,a31200a,a31201a,a31205a,a31206a,a31210a,a31211a,a31212a,a31216a,a31217a,a31221a,a31222a,a31223a,a31227a,a31228a,a31232a,a31233a,a31234a,a31238a,a31239a,a31243a,a31244a,a31245a,a31249a,a31250a,a31254a,a31255a,a31256a,a31260a,a31261a,a31265a,a31266a,a31267a,a31271a,a31272a,a31276a,a31277a,a31278a,a31282a,a31283a,a31287a,a31288a,a31289a,a31293a,a31294a,a31298a,a31299a,a31300a,a31304a,a31305a,a31309a,a31310a,a31311a,a31315a,a31316a,a31320a,a31321a,a31322a,a31326a,a31327a,a31331a,a31332a,a31333a,a31337a,a31338a,a31342a,a31343a,a31344a,a31348a,a31349a,a31353a,a31354a,a31355a,a31359a,a31360a,a31364a,a31365a,a31366a,a31370a,a31371a,a31375a,a31376a,a31377a,a31381a,a31382a,a31386a,a31387a,a31388a,a31392a,a31393a,a31397a,a31398a,a31399a,a31403a,a31404a,a31408a,a31409a,a31410a,a31414a,a31415a,a31419a,a31420a,a31421a,a31425a,a31426a,a31430a,a31431a,a31432a,a31436a,a31437a,a31441a,a31442a,a31443a,a31447a,a31448a,a31452a,a31453a,a31454a,a31458a,a31459a,a31463a,a31464a,a31465a,a31469a,a31470a,a31474a,a31475a,a31476a,a31480a,a31481a,a31485a,a31486a,a31487a,a31491a,a31492a,a31496a,a31497a,a31498a,a31502a,a31503a,a31507a,a31508a,a31509a,a31513a,a31514a,a31518a,a31519a,a31520a,a31524a,a31525a,a31529a,a31530a,a31531a,a31535a,a31536a,a31540a,a31541a,a31542a,a31546a,a31547a,a31551a,a31552a,a31553a,a31557a,a31558a,a31562a,a31563a,a31564a,a31568a,a31569a,a31573a,a31574a,a31575a,a31579a,a31580a,a31584a,a31585a,a31586a,a31590a,a31591a,a31595a,a31596a,a31597a,a31601a,a31602a,a31606a,a31607a,a31608a,a31612a,a31613a,a31617a,a31618a,a31619a,a31623a,a31624a,a31628a,a31629a,a31630a,a31634a,a31635a,a31639a,a31640a,a31641a,a31645a,a31646a,a31650a,a31651a,a31652a,a31656a,a31657a,a31661a,a31662a,a31663a,a31667a,a31668a,a31672a,a31673a,a31674a,a31678a,a31679a,a31683a,a31684a,a31685a,a31689a,a31690a,a31694a,a31695a,a31696a,a31700a,a31701a,a31705a,a31706a,a31707a,a31711a,a31712a,a31716a,a31717a,a31718a,a31722a,a31723a,a31727a,a31728a,a31729a,a31733a,a31734a,a31738a,a31739a,a31740a,a31744a,a31745a,a31749a,a31750a,a31751a,a31755a,a31756a,a31760a,a31761a,a31762a,a31766a,a31767a,a31771a,a31772a,a31773a,a31777a,a31778a,a31782a,a31783a,a31784a,a31788a,a31789a,a31793a,a31794a,a31795a,a31799a,a31800a,a31804a,a31805a,a31806a,a31810a,a31811a,a31815a,a31816a,a31817a,a31821a,a31822a,a31826a,a31827a,a31828a,a31832a,a31833a,a31837a,a31838a,a31839a,a31843a,a31844a,a31848a,a31849a,a31850a,a31854a,a31855a,a31859a,a31860a,a31861a,a31865a,a31866a,a31870a,a31871a,a31872a,a31876a,a31877a,a31881a,a31882a,a31883a,a31887a,a31888a,a31892a,a31893a,a31894a,a31898a,a31899a,a31903a,a31904a,a31905a,a31909a,a31910a,a31914a,a31915a,a31916a,a31920a,a31921a,a31925a,a31926a,a31927a,a31931a,a31932a,a31936a,a31937a,a31938a,a31942a,a31943a,a31947a,a31948a,a31949a,a31953a,a31954a,a31958a,a31959a,a31960a,a31964a,a31965a,a31969a,a31970a,a31971a,a31975a,a31976a,a31980a,a31981a,a31982a,a31986a,a31987a,a31991a,a31992a,a31993a,a31997a,a31998a,a32002a,a32003a,a32004a,a32008a,a32009a,a32013a,a32014a,a32015a,a32019a,a32020a,a32024a,a32025a,a32026a,a32030a,a32031a,a32035a,a32036a,a32037a,a32041a,a32042a,a32046a,a32047a,a32048a,a32052a,a32053a,a32057a,a32058a,a32059a,a32063a,a32064a,a32068a,a32069a,a32070a,a32074a,a32075a,a32079a,a32080a,a32081a,a32085a,a32086a,a32090a,a32091a,a32092a,a32096a,a32097a,a32101a,a32102a,a32103a,a32107a,a32108a,a32112a,a32113a,a32114a,a32118a,a32119a,a32123a,a32124a,a32125a,a32129a,a32130a,a32134a,a32135a,a32136a,a32140a,a32141a,a32145a,a32146a,a32147a,a32151a,a32152a,a32156a,a32157a,a32158a,a32162a,a32163a,a32167a,a32168a,a32169a,a32173a,a32174a,a32178a,a32179a,a32180a,a32184a,a32185a,a32189a,a32190a,a32191a,a32195a,a32196a,a32200a,a32201a,a32202a,a32206a,a32207a,a32211a,a32212a,a32213a,a32217a,a32218a,a32222a,a32223a,a32224a,a32228a,a32229a,a32233a,a32234a,a32235a,a32239a,a32240a,a32244a,a32245a,a32246a,a32250a,a32251a,a32255a,a32256a,a32257a,a32261a,a32262a,a32266a,a32267a,a32268a,a32272a,a32273a,a32277a,a32278a,a32279a,a32283a,a32284a,a32288a,a32289a,a32290a,a32294a,a32295a,a32299a,a32300a,a32301a,a32305a,a32306a,a32310a,a32311a,a32312a,a32316a,a32317a,a32321a,a32322a,a32323a,a32327a,a32328a,a32332a,a32333a,a32334a,a32338a,a32339a,a32343a,a32344a,a32345a,a32349a,a32350a,a32354a,a32355a,a32356a,a32360a,a32361a,a32365a,a32366a,a32367a,a32371a,a32372a,a32376a,a32377a,a32378a,a32382a,a32383a,a32387a,a32388a,a32389a,a32393a,a32394a,a32398a,a32399a,a32400a,a32404a,a32405a,a32409a,a32410a,a32411a,a32415a,a32416a,a32420a,a32421a,a32422a,a32426a,a32427a,a32431a,a32432a,a32433a,a32437a,a32438a,a32442a,a32443a,a32444a,a32448a,a32449a,a32453a,a32454a,a32455a,a32459a,a32460a,a32464a,a32465a,a32466a,a32470a,a32471a,a32475a,a32476a,a32477a,a32481a,a32482a,a32486a,a32487a,a32488a,a32492a,a32493a,a32497a,a32498a,a32499a,a32503a,a32504a,a32508a,a32509a,a32510a,a32514a,a32515a,a32519a,a32520a,a32521a,a32525a,a32526a,a32530a,a32531a,a32532a,a32536a,a32537a,a32541a,a32542a,a32543a,a32547a,a32548a,a32552a,a32553a,a32554a,a32558a,a32559a,a32563a,a32564a,a32565a,a32569a,a32570a,a32574a,a32575a,a32576a,a32580a,a32581a,a32585a,a32586a,a32587a,a32591a,a32592a,a32596a,a32597a,a32598a,a32602a,a32603a,a32607a,a32608a,a32609a,a32613a,a32614a,a32618a,a32619a,a32620a,a32624a,a32625a,a32629a,a32630a,a32631a,a32635a,a32636a,a32640a,a32641a,a32642a,a32646a,a32647a,a32651a,a32652a,a32653a,a32657a,a32658a,a32662a,a32663a,a32664a,a32668a,a32669a,a32673a,a32674a,a32675a,a32679a,a32680a,a32684a,a32685a,a32686a,a32690a,a32691a,a32695a,a32696a,a32697a,a32701a,a32702a,a32706a,a32707a,a32708a,a32712a,a32713a,a32717a,a32718a,a32719a,a32723a,a32724a,a32728a,a32729a,a32730a,a32734a,a32735a,a32739a,a32740a,a32741a,a32745a,a32746a,a32750a,a32751a,a32752a,a32756a,a32757a,a32761a,a32762a,a32763a,a32767a,a32768a,a32772a,a32773a,a32774a,a32778a,a32779a,a32783a,a32784a,a32785a,a32789a,a32790a,a32794a,a32795a,a32796a,a32800a,a32801a,a32805a,a32806a,a32807a,a32811a,a32812a,a32816a,a32817a,a32818a,a32822a,a32823a,a32827a,a32828a,a32829a,a32833a,a32834a,a32838a,a32839a,a32840a,a32844a,a32845a,a32849a,a32850a,a32851a,a32855a,a32856a,a32860a,a32861a,a32862a,a32866a,a32867a,a32871a,a32872a,a32873a,a32877a,a32878a,a32882a,a32883a,a32884a,a32888a,a32889a,a32893a,a32894a,a32895a,a32899a,a32900a,a32904a,a32905a,a32906a,a32910a,a32911a,a32915a,a32916a,a32917a,a32921a,a32922a,a32926a,a32927a,a32928a,a32932a,a32933a,a32937a,a32938a,a32939a,a32943a,a32944a,a32948a,a32949a,a32950a,a32954a,a32955a,a32959a,a32960a,a32961a,a32965a,a32966a,a32970a,a32971a,a32972a,a32976a,a32977a,a32981a,a32982a,a32983a,a32987a,a32988a,a32992a,a32993a,a32994a,a32998a,a32999a,a33003a,a33004a,a33005a,a33009a,a33010a,a33014a,a33015a,a33016a,a33020a,a33021a,a33025a,a33026a,a33027a,a33031a,a33032a,a33036a,a33037a,a33038a,a33042a,a33043a,a33047a,a33048a,a33049a,a33053a,a33054a,a33058a,a33059a,a33060a,a33064a,a33065a,a33069a,a33070a,a33071a,a33075a,a33076a,a33080a,a33081a,a33082a,a33086a,a33087a,a33091a,a33092a,a33093a,a33097a,a33098a,a33102a,a33103a,a33104a,a33108a,a33109a,a33113a,a33114a,a33115a,a33119a,a33120a,a33124a,a33125a,a33126a,a33130a,a33131a,a33135a,a33136a,a33137a,a33141a,a33142a,a33146a,a33147a,a33148a,a33152a,a33153a,a33157a,a33158a,a33159a,a33163a,a33164a,a33168a,a33169a,a33170a,a33174a,a33175a,a33179a,a33180a,a33181a,a33185a,a33186a,a33190a,a33191a,a33192a,a33196a,a33197a,a33201a,a33202a,a33203a,a33207a,a33208a,a33212a,a33213a,a33214a,a33218a,a33219a,a33223a,a33224a,a33225a,a33229a,a33230a,a33234a,a33235a,a33236a,a33240a,a33241a,a33245a,a33246a,a33247a,a33251a,a33252a,a33256a,a33257a,a33258a,a33262a,a33263a,a33267a,a33268a,a33269a,a33273a,a33274a,a33278a,a33279a,a33280a,a33284a,a33285a,a33289a,a33290a,a33291a,a33295a,a33296a,a33300a,a33301a,a33302a,a33306a,a33307a,a33311a,a33312a,a33313a,a33317a,a33318a,a33322a,a33323a,a33324a,a33328a,a33329a,a33333a,a33334a,a33335a,a33339a,a33340a,a33344a,a33345a,a33346a,a33350a,a33351a,a33355a,a33356a,a33357a,a33361a,a33362a,a33366a,a33367a,a33368a,a33372a,a33373a,a33377a,a33378a,a33379a,a33383a,a33384a,a33388a,a33389a,a33390a,a33394a,a33395a,a33399a,a33400a,a33401a,a33405a,a33406a,a33410a,a33411a,a33412a,a33416a,a33417a,a33421a,a33422a,a33423a,a33427a,a33428a,a33432a,a33433a,a33434a,a33438a,a33439a,a33443a,a33444a,a33445a,a33449a,a33450a,a33454a,a33455a,a33456a,a33460a,a33461a,a33465a,a33466a,a33467a,a33471a,a33472a,a33476a,a33477a,a33478a,a33482a,a33483a,a33487a,a33488a,a33489a,a33493a,a33494a,a33498a,a33499a,a33500a,a33504a,a33505a,a33509a,a33510a,a33511a,a33515a,a33516a,a33520a,a33521a,a33522a,a33526a,a33527a,a33531a,a33532a,a33533a,a33537a,a33538a,a33542a,a33543a,a33544a,a33548a,a33549a,a33553a,a33554a,a33555a,a33559a,a33560a,a33564a,a33565a,a33566a,a33570a,a33571a,a33575a,a33576a,a33577a,a33581a,a33582a,a33586a,a33587a,a33588a,a33592a,a33593a,a33597a,a33598a,a33599a,a33603a,a33604a,a33608a,a33609a,a33610a,a33614a,a33615a,a33619a,a33620a,a33621a,a33625a,a33626a,a33630a,a33631a,a33632a,a33636a,a33637a,a33641a,a33642a,a33643a,a33647a,a33648a,a33652a,a33653a,a33654a,a33658a,a33659a,a33663a,a33664a,a33665a,a33669a,a33670a,a33674a,a33675a,a33676a,a33680a,a33681a,a33685a,a33686a,a33687a,a33691a,a33692a,a33696a,a33697a,a33698a,a33702a,a33703a,a33707a,a33708a,a33709a,a33713a,a33714a,a33718a,a33719a,a33720a,a33724a,a33725a,a33729a,a33730a,a33731a,a33735a,a33736a,a33740a,a33741a,a33742a,a33746a,a33747a,a33751a,a33752a,a33753a,a33757a,a33758a,a33762a,a33763a,a33764a,a33768a,a33769a,a33773a,a33774a,a33775a,a33779a,a33780a,a33784a,a33785a,a33786a,a33790a,a33791a,a33795a,a33796a,a33797a,a33801a,a33802a,a33806a,a33807a,a33808a,a33812a,a33813a,a33817a,a33818a,a33819a,a33823a,a33824a,a33828a,a33829a,a33830a,a33834a,a33835a,a33839a,a33840a,a33841a,a33845a,a33846a,a33850a,a33851a,a33852a,a33856a,a33857a,a33861a,a33862a,a33863a,a33867a,a33868a,a33872a,a33873a,a33874a,a33878a,a33879a,a33883a,a33884a,a33885a,a33889a,a33890a,a33894a,a33895a,a33896a,a33900a,a33901a,a33905a,a33906a,a33907a,a33911a,a33912a,a33916a,a33917a,a33918a,a33922a,a33923a,a33927a,a33928a,a33929a,a33933a,a33934a,a33938a,a33939a,a33940a,a33944a,a33945a,a33949a,a33950a,a33951a,a33955a,a33956a,a33960a,a33961a,a33962a,a33966a,a33967a,a33971a,a33972a,a33973a,a33977a,a33978a,a33982a,a33983a,a33984a,a33988a,a33989a,a33993a,a33994a,a33995a,a33999a,a34000a,a34004a,a34005a,a34006a,a34010a,a34011a,a34015a,a34016a,a34017a,a34021a,a34022a,a34026a,a34027a,a34028a,a34032a,a34033a,a34037a,a34038a,a34039a,a34043a,a34044a,a34048a,a34049a,a34050a,a34054a,a34055a,a34059a,a34060a,a34061a,a34065a,a34066a,a34070a,a34071a,a34072a,a34076a,a34077a,a34081a,a34082a,a34083a,a34087a,a34088a,a34092a,a34093a,a34094a,a34098a,a34099a,a34103a,a34104a,a34105a,a34109a,a34110a,a34114a,a34115a,a34116a,a34120a,a34121a,a34125a,a34126a,a34127a,a34131a,a34132a,a34136a,a34137a,a34138a,a34142a,a34143a,a34147a,a34148a,a34149a,a34153a,a34154a,a34158a,a34159a,a34160a,a34164a,a34165a,a34169a,a34170a,a34171a,a34175a,a34176a,a34180a,a34181a,a34182a,a34186a,a34187a,a34191a,a34192a,a34193a,a34197a,a34198a,a34202a,a34203a,a34204a,a34208a,a34209a,a34213a,a34214a,a34215a,a34219a,a34220a,a34224a,a34225a,a34226a,a34230a,a34231a,a34235a,a34236a,a34237a,a34241a,a34242a,a34246a,a34247a,a34248a,a34252a,a34253a,a34257a,a34258a,a34259a,a34263a,a34264a,a34268a,a34269a,a34270a,a34274a,a34275a,a34279a,a34280a,a34281a,a34285a,a34286a,a34290a,a34291a,a34292a,a34296a,a34297a,a34301a,a34302a,a34303a,a34307a,a34308a,a34312a,a34313a,a34314a,a34318a,a34319a,a34323a,a34324a,a34325a,a34329a,a34330a,a34334a,a34335a,a34336a,a34340a,a34341a,a34345a,a34346a,a34347a,a34351a,a34352a,a34356a,a34357a,a34358a,a34362a,a34363a,a34367a,a34368a,a34369a,a34373a,a34374a,a34378a,a34379a,a34380a,a34384a,a34385a,a34389a,a34390a,a34391a,a34395a,a34396a,a34400a,a34401a,a34402a,a34406a,a34407a,a34411a,a34412a,a34413a,a34417a,a34418a,a34422a,a34423a,a34424a,a34428a,a34429a,a34433a,a34434a,a34435a,a34439a,a34440a,a34444a,a34445a,a34446a,a34450a,a34451a,a34455a,a34456a,a34457a,a34461a,a34462a,a34466a,a34467a,a34468a,a34472a,a34473a,a34477a,a34478a,a34479a,a34483a,a34484a,a34488a,a34489a,a34490a,a34494a,a34495a,a34499a,a34500a,a34501a,a34505a,a34506a,a34510a,a34511a,a34512a,a34516a,a34517a,a34521a,a34522a,a34523a,a34527a,a34528a,a34532a,a34533a,a34534a,a34538a,a34539a,a34543a,a34544a,a34545a,a34549a,a34550a,a34554a,a34555a,a34556a,a34560a,a34561a,a34565a,a34566a,a34567a,a34571a,a34572a,a34576a,a34577a,a34578a,a34582a,a34583a,a34587a,a34588a,a34589a,a34593a,a34594a,a34598a,a34599a,a34600a,a34604a,a34605a,a34609a,a34610a,a34611a,a34615a,a34616a,a34620a,a34621a,a34622a,a34626a,a34627a,a34631a,a34632a,a34633a,a34637a,a34638a,a34642a,a34643a,a34644a,a34648a,a34649a,a34653a,a34654a,a34655a,a34659a,a34660a,a34664a,a34665a,a34666a,a34670a,a34671a,a34675a,a34676a,a34677a,a34681a,a34682a,a34686a,a34687a,a34688a,a34692a,a34693a,a34697a,a34698a,a34699a,a34703a,a34704a,a34708a,a34709a,a34710a,a34714a,a34715a,a34719a,a34720a,a34721a,a34725a,a34726a,a34730a,a34731a,a34732a,a34736a,a34737a,a34741a,a34742a,a34743a,a34747a,a34748a,a34752a,a34753a,a34754a,a34758a,a34759a,a34763a,a34764a,a34765a,a34769a,a34770a,a34774a,a34775a,a34776a,a34780a,a34781a,a34785a,a34786a,a34787a,a34791a,a34792a,a34796a,a34797a,a34798a,a34802a,a34803a,a34807a,a34808a,a34809a,a34813a,a34814a,a34818a,a34819a,a34820a,a34824a,a34825a,a34829a,a34830a,a34831a,a34835a,a34836a,a34840a,a34841a,a34842a,a34846a,a34847a,a34851a,a34852a,a34853a,a34857a,a34858a,a34862a,a34863a,a34864a,a34868a,a34869a,a34873a,a34874a,a34875a,a34879a,a34880a,a34884a,a34885a,a34886a,a34890a,a34891a,a34895a,a34896a,a34897a,a34901a,a34902a,a34906a,a34907a,a34908a,a34912a,a34913a,a34917a,a34918a,a34919a,a34923a,a34924a,a34928a,a34929a,a34930a,a34934a,a34935a,a34939a,a34940a,a34941a,a34945a,a34946a,a34950a,a34951a,a34952a,a34956a,a34957a,a34961a,a34962a,a34963a,a34967a,a34968a,a34972a,a34973a,a34974a,a34978a,a34979a,a34983a,a34984a,a34985a,a34989a,a34990a,a34994a,a34995a,a34996a,a35000a,a35001a,a35005a,a35006a,a35007a,a35011a,a35012a,a35016a,a35017a,a35018a,a35022a,a35023a,a35027a,a35028a,a35029a,a35033a,a35034a,a35038a,a35039a,a35040a,a35044a,a35045a,a35049a,a35050a,a35051a,a35055a,a35056a,a35060a,a35061a,a35062a,a35066a,a35067a,a35071a,a35072a,a35073a,a35077a,a35078a,a35082a,a35083a,a35084a,a35088a,a35089a,a35093a,a35094a,a35095a,a35099a,a35100a,a35104a,a35105a,a35106a,a35110a,a35111a,a35115a,a35116a,a35117a,a35121a,a35122a,a35126a,a35127a,a35128a,a35132a,a35133a,a35137a,a35138a,a35139a,a35143a,a35144a,a35148a,a35149a,a35150a,a35154a,a35155a,a35159a,a35160a,a35161a,a35165a,a35166a,a35170a,a35171a,a35172a,a35176a,a35177a,a35181a,a35182a,a35183a,a35187a,a35188a,a35192a,a35193a,a35194a,a35198a,a35199a,a35203a,a35204a,a35205a,a35209a,a35210a,a35214a,a35215a,a35216a,a35220a,a35221a,a35225a,a35226a,a35227a,a35231a,a35232a,a35236a,a35237a,a35238a,a35242a,a35243a,a35247a,a35248a,a35249a,a35253a,a35254a,a35258a,a35259a,a35260a,a35264a,a35265a,a35269a,a35270a,a35271a,a35275a,a35276a,a35280a,a35281a,a35282a,a35286a,a35287a,a35291a,a35292a,a35293a,a35297a,a35298a,a35302a,a35303a,a35304a,a35308a,a35309a,a35313a,a35314a,a35315a,a35319a,a35320a,a35324a,a35325a,a35326a,a35330a,a35331a,a35335a,a35336a,a35337a,a35341a,a35342a,a35346a,a35347a,a35348a,a35352a,a35353a,a35357a,a35358a,a35359a,a35363a,a35364a,a35368a,a35369a,a35370a,a35374a,a35375a,a35379a,a35380a,a35381a,a35385a,a35386a,a35390a,a35391a,a35392a,a35396a,a35397a,a35401a,a35402a,a35403a,a35407a,a35408a,a35412a,a35413a,a35414a,a35418a,a35419a,a35423a,a35424a,a35425a,a35429a,a35430a,a35434a,a35435a,a35436a,a35440a,a35441a,a35445a,a35446a,a35447a,a35451a,a35452a,a35456a,a35457a,a35458a,a35462a,a35463a,a35467a,a35468a,a35469a,a35473a,a35474a,a35478a,a35479a,a35480a,a35484a,a35485a,a35489a,a35490a,a35491a,a35495a,a35496a,a35500a,a35501a,a35502a,a35506a,a35507a,a35511a,a35512a,a35513a,a35517a,a35518a,a35522a,a35523a,a35524a,a35528a,a35529a,a35533a,a35534a,a35535a,a35539a,a35540a,a35544a,a35545a,a35546a,a35550a,a35551a,a35555a,a35556a,a35557a,a35561a,a35562a,a35566a,a35567a,a35568a,a35572a,a35573a,a35577a,a35578a,a35579a,a35583a,a35584a,a35588a,a35589a,a35590a,a35594a,a35595a,a35599a,a35600a,a35601a,a35605a,a35606a,a35610a,a35611a,a35612a,a35616a,a35617a,a35621a,a35622a,a35623a,a35627a,a35628a,a35632a,a35633a,a35634a,a35638a,a35639a,a35643a,a35644a,a35645a,a35649a,a35650a,a35654a,a35655a,a35656a,a35660a,a35661a,a35665a,a35666a,a35667a,a35671a,a35672a,a35676a,a35677a,a35678a,a35682a,a35683a,a35687a,a35688a,a35689a,a35693a,a35694a,a35698a,a35699a,a35700a,a35704a,a35705a,a35709a,a35710a,a35711a,a35715a,a35716a,a35720a,a35721a,a35722a,a35726a,a35727a,a35731a,a35732a,a35733a,a35737a,a35738a,a35742a,a35743a,a35744a,a35748a,a35749a,a35753a,a35754a,a35755a,a35759a,a35760a,a35764a,a35765a,a35766a,a35770a,a35771a,a35775a,a35776a,a35777a,a35781a,a35782a,a35786a,a35787a,a35788a,a35792a,a35793a,a35797a,a35798a,a35799a,a35803a,a35804a,a35808a,a35809a,a35810a,a35814a,a35815a,a35819a,a35820a,a35821a,a35825a,a35826a,a35830a,a35831a,a35832a,a35836a,a35837a,a35841a,a35842a,a35843a,a35847a,a35848a,a35852a,a35853a,a35854a,a35858a,a35859a,a35863a,a35864a,a35865a,a35869a,a35870a,a35874a,a35875a,a35876a,a35880a,a35881a,a35885a,a35886a,a35887a,a35891a,a35892a,a35896a,a35897a,a35898a,a35902a,a35903a,a35907a,a35908a,a35909a,a35913a,a35914a,a35918a,a35919a,a35920a,a35924a,a35925a,a35929a,a35930a,a35931a,a35935a,a35936a,a35940a,a35941a,a35942a,a35946a,a35947a,a35951a,a35952a,a35953a,a35957a,a35958a,a35962a,a35963a,a35964a,a35968a,a35969a,a35973a,a35974a,a35975a,a35979a,a35980a,a35984a,a35985a,a35986a,a35990a,a35991a,a35995a,a35996a,a35997a,a36001a,a36002a,a36006a,a36007a,a36008a,a36012a,a36013a,a36017a,a36018a,a36019a,a36023a,a36024a,a36028a,a36029a,a36030a,a36034a,a36035a,a36039a,a36040a,a36041a,a36045a,a36046a,a36050a,a36051a,a36052a,a36056a,a36057a,a36061a,a36062a,a36063a,a36067a,a36068a,a36072a,a36073a,a36074a,a36078a,a36079a,a36083a,a36084a,a36085a,a36089a,a36090a,a36094a,a36095a,a36096a,a36100a,a36101a,a36105a,a36106a,a36107a,a36111a,a36112a,a36116a,a36117a,a36118a,a36122a,a36123a,a36127a,a36128a,a36129a,a36133a,a36134a,a36138a,a36139a,a36140a,a36144a,a36145a,a36149a,a36150a,a36151a,a36155a,a36156a,a36160a,a36161a,a36162a,a36166a,a36167a,a36171a,a36172a,a36173a,a36177a,a36178a,a36182a,a36183a,a36184a,a36188a,a36189a,a36193a,a36194a,a36195a,a36199a,a36200a,a36204a,a36205a,a36206a,a36210a,a36211a,a36215a,a36216a,a36217a,a36221a,a36222a,a36226a,a36227a,a36228a,a36232a,a36233a,a36237a,a36238a,a36239a,a36243a,a36244a,a36248a,a36249a,a36250a,a36254a,a36255a,a36259a,a36260a,a36261a,a36265a,a36266a,a36270a,a36271a,a36272a,a36276a,a36277a,a36281a,a36282a,a36283a,a36287a,a36288a,a36292a,a36293a,a36294a,a36298a,a36299a,a36303a,a36304a,a36305a,a36309a,a36310a,a36314a,a36315a,a36316a,a36320a,a36321a,a36325a,a36326a,a36327a,a36331a,a36332a,a36336a,a36337a,a36338a,a36342a,a36343a,a36347a,a36348a,a36349a,a36353a,a36354a,a36358a,a36359a,a36360a,a36364a,a36365a,a36369a,a36370a,a36371a,a36375a,a36376a,a36380a,a36381a,a36382a,a36386a,a36387a,a36391a,a36392a,a36393a,a36397a,a36398a,a36402a,a36403a,a36404a,a36408a,a36409a,a36413a,a36414a,a36415a,a36419a,a36420a,a36424a,a36425a,a36426a,a36430a,a36431a,a36435a,a36436a,a36437a,a36441a,a36442a,a36446a,a36447a,a36448a,a36452a,a36453a,a36457a,a36458a,a36459a,a36463a,a36464a,a36468a,a36469a,a36470a,a36474a,a36475a,a36479a,a36480a,a36481a,a36485a,a36486a,a36490a,a36491a,a36492a,a36496a,a36497a,a36501a,a36502a,a36503a,a36507a,a36508a,a36512a,a36513a,a36514a,a36518a,a36519a,a36523a,a36524a,a36525a,a36529a,a36530a,a36534a,a36535a,a36536a,a36540a,a36541a,a36545a,a36546a,a36547a,a36551a,a36552a,a36556a,a36557a,a36558a,a36562a,a36563a,a36567a,a36568a,a36569a,a36573a,a36574a,a36578a,a36579a,a36580a,a36584a,a36585a,a36589a,a36590a,a36591a,a36595a,a36596a,a36600a,a36601a,a36602a,a36606a,a36607a,a36611a,a36612a,a36613a,a36617a,a36618a,a36622a,a36623a,a36624a,a36628a,a36629a,a36633a,a36634a,a36635a,a36639a,a36640a,a36644a,a36645a,a36646a,a36650a,a36651a,a36655a,a36656a,a36657a,a36661a,a36662a,a36666a,a36667a,a36668a,a36672a,a36673a,a36677a,a36678a,a36679a,a36683a,a36684a,a36688a,a36689a,a36690a,a36694a,a36695a,a36699a,a36700a,a36701a,a36705a,a36706a,a36710a,a36711a,a36712a,a36716a,a36717a,a36721a,a36722a,a36723a,a36727a,a36728a,a36732a,a36733a,a36734a,a36738a,a36739a,a36743a,a36744a,a36745a,a36749a,a36750a,a36754a,a36755a,a36756a,a36760a,a36761a,a36765a,a36766a,a36767a,a36771a,a36772a,a36776a,a36777a,a36778a,a36782a,a36783a,a36787a,a36788a,a36789a,a36793a,a36794a,a36798a,a36799a,a36800a,a36804a,a36805a,a36809a,a36810a,a36811a,a36815a,a36816a,a36820a,a36821a,a36822a,a36826a,a36827a,a36831a,a36832a,a36833a,a36837a,a36838a,a36842a,a36843a,a36844a,a36848a,a36849a,a36853a,a36854a,a36855a,a36859a,a36860a,a36864a,a36865a,a36866a,a36870a,a36871a,a36875a,a36876a,a36877a,a36881a,a36882a,a36886a,a36887a,a36888a,a36892a,a36893a,a36897a,a36898a,a36899a,a36903a,a36904a,a36908a,a36909a,a36910a,a36914a,a36915a,a36919a,a36920a,a36921a,a36925a,a36926a,a36930a,a36931a,a36932a,a36936a,a36937a,a36941a,a36942a,a36943a,a36947a,a36948a,a36952a,a36953a,a36954a,a36958a,a36959a,a36963a,a36964a,a36965a,a36969a,a36970a,a36974a,a36975a,a36976a,a36980a,a36981a,a36985a,a36986a,a36987a,a36991a,a36992a,a36996a,a36997a,a36998a,a37002a,a37003a,a37007a,a37008a,a37009a,a37013a,a37014a,a37018a,a37019a,a37020a,a37024a,a37025a,a37029a,a37030a,a37031a,a37035a,a37036a,a37040a,a37041a,a37042a,a37046a,a37047a,a37051a,a37052a,a37053a,a37057a,a37058a,a37062a,a37063a,a37064a,a37068a,a37069a,a37073a,a37074a,a37075a,a37079a,a37080a,a37084a,a37085a,a37086a,a37090a,a37091a,a37095a,a37096a,a37097a,a37101a,a37102a,a37106a,a37107a,a37108a,a37112a,a37113a,a37117a,a37118a,a37119a,a37123a,a37124a,a37128a,a37129a,a37130a,a37134a,a37135a,a37139a,a37140a,a37141a,a37145a,a37146a,a37150a,a37151a,a37152a,a37156a,a37157a,a37161a,a37162a,a37163a,a37167a,a37168a,a37172a,a37173a,a37174a,a37178a,a37179a,a37183a,a37184a,a37185a,a37189a,a37190a,a37194a,a37195a,a37196a,a37200a,a37201a,a37205a,a37206a,a37207a,a37211a,a37212a,a37216a,a37217a,a37218a,a37222a,a37223a,a37227a,a37228a,a37229a,a37233a,a37234a,a37238a,a37239a,a37240a,a37244a,a37245a,a37249a,a37250a,a37251a,a37255a,a37256a,a37260a,a37261a,a37262a,a37266a,a37267a,a37271a,a37272a,a37273a,a37277a,a37278a,a37282a,a37283a,a37284a,a37288a,a37289a,a37293a,a37294a,a37295a,a37299a,a37300a,a37304a,a37305a,a37306a,a37310a,a37311a,a37315a,a37316a,a37317a,a37321a,a37322a,a37326a,a37327a,a37328a,a37332a,a37333a,a37337a,a37338a,a37339a,a37343a,a37344a,a37348a,a37349a,a37350a,a37354a,a37355a,a37359a,a37360a,a37361a,a37365a,a37366a,a37370a,a37371a,a37372a,a37376a,a37377a,a37381a,a37382a,a37383a,a37387a,a37388a,a37392a,a37393a,a37394a,a37398a,a37399a,a37403a,a37404a,a37405a,a37409a,a37410a,a37414a,a37415a,a37416a,a37420a,a37421a,a37425a,a37426a,a37427a,a37431a,a37432a,a37436a,a37437a,a37438a,a37442a,a37443a,a37447a,a37448a,a37449a,a37453a,a37454a,a37458a,a37459a,a37460a,a37464a,a37465a,a37469a,a37470a,a37471a,a37475a,a37476a,a37480a,a37481a,a37482a,a37486a,a37487a,a37491a,a37492a,a37493a,a37497a,a37498a,a37502a,a37503a,a37504a,a37508a,a37509a,a37513a,a37514a,a37515a,a37519a,a37520a,a37524a,a37525a,a37526a,a37530a,a37531a,a37535a,a37536a,a37537a,a37541a,a37542a,a37546a,a37547a,a37548a,a37552a,a37553a,a37557a,a37558a,a37559a,a37563a,a37564a,a37568a,a37569a,a37570a,a37574a,a37575a,a37579a,a37580a,a37581a,a37585a,a37586a,a37590a,a37591a,a37592a,a37596a,a37597a,a37601a,a37602a,a37603a,a37607a,a37608a,a37612a,a37613a,a37614a,a37618a,a37619a,a37623a,a37624a,a37625a,a37629a,a37630a,a37634a,a37635a,a37636a,a37640a,a37641a,a37645a,a37646a,a37647a,a37651a,a37652a,a37656a,a37657a,a37658a,a37662a,a37663a,a37667a,a37668a,a37669a,a37673a,a37674a,a37678a,a37679a,a37680a,a37684a,a37685a,a37689a,a37690a,a37691a,a37695a,a37696a,a37700a,a37701a,a37702a,a37706a,a37707a,a37711a,a37712a,a37713a,a37717a,a37718a,a37722a,a37723a,a37724a,a37728a,a37729a,a37733a,a37734a,a37735a,a37739a,a37740a,a37744a,a37745a,a37746a,a37750a,a37751a,a37755a,a37756a,a37757a,a37761a,a37762a,a37766a,a37767a,a37768a,a37772a,a37773a,a37777a,a37778a,a37779a,a37783a,a37784a,a37788a,a37789a,a37790a,a37794a,a37795a,a37799a,a37800a,a37801a,a37805a,a37806a,a37810a,a37811a,a37812a,a37816a,a37817a,a37821a,a37822a,a37823a,a37827a,a37828a,a37832a,a37833a,a37834a,a37838a,a37839a,a37843a,a37844a,a37845a,a37849a,a37850a,a37854a,a37855a,a37856a,a37860a,a37861a,a37865a,a37866a,a37867a,a37871a,a37872a,a37876a,a37877a,a37878a,a37882a,a37883a,a37887a,a37888a,a37889a,a37893a,a37894a,a37898a,a37899a,a37900a,a37904a,a37905a,a37909a,a37910a,a37911a,a37915a,a37916a,a37920a,a37921a,a37922a,a37926a,a37927a,a37931a,a37932a,a37933a,a37937a,a37938a,a37942a,a37943a,a37944a,a37948a,a37949a,a37953a,a37954a,a37955a,a37959a,a37960a,a37964a,a37965a,a37966a,a37970a,a37971a,a37975a,a37976a,a37977a,a37981a,a37982a,a37986a,a37987a,a37988a,a37992a,a37993a,a37997a,a37998a,a37999a,a38003a,a38004a,a38008a,a38009a,a38010a,a38014a,a38015a,a38019a,a38020a,a38021a,a38025a,a38026a,a38030a,a38031a,a38032a,a38036a,a38037a,a38041a,a38042a,a38043a,a38047a,a38048a,a38052a,a38053a,a38054a,a38058a,a38059a,a38063a,a38064a,a38065a,a38069a,a38070a,a38074a,a38075a,a38076a,a38080a,a38081a,a38085a,a38086a,a38087a,a38091a,a38092a,a38096a,a38097a,a38098a,a38102a,a38103a,a38107a,a38108a,a38109a,a38113a,a38114a,a38118a,a38119a,a38120a,a38124a,a38125a,a38129a,a38130a,a38131a,a38135a,a38136a,a38140a,a38141a,a38142a,a38146a,a38147a,a38151a,a38152a,a38153a,a38157a,a38158a,a38162a,a38163a,a38164a,a38168a,a38169a,a38173a,a38174a,a38175a,a38179a,a38180a,a38184a,a38185a,a38186a,a38190a,a38191a,a38195a,a38196a,a38197a,a38201a,a38202a,a38206a,a38207a,a38208a,a38212a,a38213a,a38217a,a38218a,a38219a,a38223a,a38224a,a38228a,a38229a,a38230a,a38234a,a38235a,a38239a,a38240a,a38241a,a38245a,a38246a,a38250a,a38251a,a38252a,a38256a,a38257a,a38261a,a38262a,a38263a,a38267a,a38268a,a38272a,a38273a,a38274a,a38278a,a38279a,a38283a,a38284a,a38285a,a38289a,a38290a,a38294a,a38295a,a38296a,a38300a,a38301a,a38305a,a38306a,a38307a,a38311a,a38312a,a38316a,a38317a,a38318a,a38322a,a38323a,a38327a,a38328a,a38329a,a38333a,a38334a,a38338a,a38339a,a38340a,a38344a,a38345a,a38349a,a38350a,a38351a,a38355a,a38356a,a38360a,a38361a,a38362a,a38366a,a38367a,a38371a,a38372a,a38373a,a38377a,a38378a,a38382a,a38383a,a38384a,a38388a,a38389a,a38393a,a38394a,a38395a,a38399a,a38400a,a38404a,a38405a,a38406a,a38410a,a38411a,a38415a,a38416a,a38417a,a38421a,a38422a,a38426a,a38427a,a38428a,a38432a,a38433a,a38437a,a38438a,a38439a,a38443a,a38444a,a38448a,a38449a,a38450a,a38454a,a38455a,a38459a,a38460a,a38461a,a38465a,a38466a,a38470a,a38471a,a38472a,a38476a,a38477a,a38481a,a38482a,a38483a,a38487a,a38488a,a38492a,a38493a,a38494a,a38498a,a38499a,a38503a,a38504a,a38505a,a38509a,a38510a,a38514a,a38515a,a38516a,a38520a,a38521a,a38525a,a38526a,a38527a,a38531a,a38532a,a38536a,a38537a,a38538a,a38542a,a38543a,a38547a,a38548a,a38549a,a38553a,a38554a,a38558a,a38559a,a38560a,a38564a,a38565a,a38569a,a38570a,a38571a,a38575a,a38576a,a38580a,a38581a,a38582a,a38586a,a38587a,a38591a,a38592a,a38593a,a38597a,a38598a,a38602a,a38603a,a38604a,a38608a,a38609a,a38613a,a38614a,a38615a,a38619a,a38620a,a38624a,a38625a,a38626a,a38630a,a38631a,a38635a,a38636a,a38637a,a38641a,a38642a,a38646a,a38647a,a38648a,a38652a,a38653a,a38657a,a38658a,a38659a,a38663a,a38664a,a38668a,a38669a,a38670a,a38674a,a38675a,a38679a,a38680a,a38681a,a38685a,a38686a,a38690a,a38691a,a38692a,a38696a,a38697a,a38701a,a38702a,a38703a,a38707a,a38708a,a38712a,a38713a,a38714a,a38718a,a38719a,a38723a,a38724a,a38725a,a38729a,a38730a,a38734a,a38735a,a38736a,a38740a,a38741a,a38745a,a38746a,a38747a,a38751a,a38752a,a38756a,a38757a,a38758a,a38762a,a38763a,a38767a,a38768a,a38769a,a38773a,a38774a,a38778a,a38779a,a38780a,a38784a,a38785a,a38789a,a38790a,a38791a,a38795a,a38796a,a38800a,a38801a,a38802a,a38806a,a38807a,a38811a,a38812a,a38813a,a38817a,a38818a,a38822a,a38823a,a38824a,a38828a,a38829a,a38833a,a38834a,a38835a,a38839a,a38840a,a38844a,a38845a,a38846a,a38850a,a38851a,a38855a,a38856a,a38857a,a38861a,a38862a,a38866a,a38867a,a38868a,a38872a,a38873a,a38877a,a38878a,a38879a,a38883a,a38884a,a38888a,a38889a,a38890a,a38894a,a38895a,a38899a,a38900a,a38901a,a38905a,a38906a,a38910a,a38911a,a38912a,a38916a,a38917a,a38921a,a38922a,a38923a,a38927a,a38928a,a38932a,a38933a,a38934a,a38938a,a38939a,a38943a,a38944a,a38945a,a38949a,a38950a,a38954a,a38955a,a38956a,a38960a,a38961a,a38965a,a38966a,a38967a,a38971a,a38972a,a38976a,a38977a,a38978a,a38982a,a38983a,a38987a,a38988a,a38989a,a38993a,a38994a,a38998a,a38999a,a39000a,a39004a,a39005a,a39009a,a39010a,a39011a,a39015a,a39016a,a39020a,a39021a,a39022a,a39026a,a39027a,a39031a,a39032a,a39033a,a39037a,a39038a,a39042a,a39043a,a39044a,a39048a,a39049a,a39053a,a39054a,a39055a,a39059a,a39060a,a39064a,a39065a,a39066a,a39070a,a39071a,a39075a,a39076a,a39077a,a39081a,a39082a,a39086a,a39087a,a39088a,a39092a,a39093a,a39097a,a39098a,a39099a,a39103a,a39104a,a39108a,a39109a,a39110a,a39114a,a39115a,a39119a,a39120a,a39121a,a39125a,a39126a,a39130a,a39131a,a39132a,a39136a,a39137a,a39141a,a39142a,a39143a,a39147a,a39148a,a39152a,a39153a,a39154a,a39158a,a39159a,a39163a,a39164a,a39165a,a39169a,a39170a,a39174a,a39175a,a39176a,a39180a,a39181a,a39185a,a39186a,a39187a,a39191a,a39192a,a39196a,a39197a,a39198a,a39202a,a39203a,a39207a,a39208a,a39209a,a39213a,a39214a,a39218a,a39219a,a39220a,a39224a,a39225a,a39229a,a39230a,a39231a,a39235a,a39236a,a39240a,a39241a,a39242a,a39246a,a39247a,a39251a,a39252a,a39253a,a39257a,a39258a,a39262a,a39263a,a39264a,a39268a,a39269a,a39273a,a39274a,a39275a,a39279a,a39280a,a39284a,a39285a,a39286a,a39290a,a39291a,a39295a,a39296a,a39297a,a39301a,a39302a,a39306a,a39307a,a39308a,a39312a,a39313a,a39317a,a39318a,a39319a,a39323a,a39324a,a39328a,a39329a,a39330a,a39334a,a39335a,a39339a,a39340a,a39341a,a39345a,a39346a,a39350a,a39351a,a39352a,a39356a,a39357a,a39361a,a39362a,a39363a,a39367a,a39368a,a39372a,a39373a,a39374a,a39378a,a39379a,a39383a,a39384a,a39385a,a39389a,a39390a,a39394a,a39395a,a39396a,a39400a,a39401a,a39405a,a39406a,a39407a,a39411a,a39412a,a39416a,a39417a,a39418a,a39422a,a39423a,a39427a,a39428a,a39429a,a39433a,a39434a,a39438a,a39439a,a39440a,a39444a,a39445a,a39449a,a39450a,a39451a,a39455a,a39456a,a39460a,a39461a,a39462a,a39466a,a39467a,a39471a,a39472a,a39473a,a39477a,a39478a,a39482a,a39483a,a39484a,a39488a,a39489a,a39493a,a39494a,a39495a,a39499a,a39500a,a39504a,a39505a,a39506a,a39510a,a39511a,a39515a,a39516a,a39517a,a39521a,a39522a,a39526a,a39527a,a39528a,a39532a,a39533a,a39537a,a39538a,a39539a,a39543a,a39544a,a39548a,a39549a,a39550a,a39554a,a39555a,a39559a,a39560a,a39561a,a39565a,a39566a,a39570a,a39571a,a39572a,a39576a,a39577a,a39581a,a39582a,a39583a,a39587a,a39588a,a39592a,a39593a,a39594a,a39598a,a39599a,a39603a,a39604a,a39605a,a39609a,a39610a,a39614a,a39615a,a39616a,a39620a,a39621a,a39625a,a39626a,a39627a,a39631a,a39632a,a39636a,a39637a,a39638a,a39642a,a39643a,a39647a,a39648a,a39649a,a39653a,a39654a,a39658a,a39659a,a39660a,a39664a,a39665a,a39669a,a39670a,a39671a,a39675a,a39676a,a39680a,a39681a,a39682a,a39686a,a39687a,a39691a,a39692a,a39693a,a39697a,a39698a,a39702a,a39703a,a39704a,a39708a,a39709a,a39713a,a39714a,a39715a,a39719a,a39720a,a39724a,a39725a,a39726a,a39730a,a39731a,a39735a,a39736a,a39737a,a39741a,a39742a,a39746a,a39747a,a39748a,a39752a,a39753a,a39757a,a39758a,a39759a,a39763a,a39764a,a39768a,a39769a,a39770a,a39774a,a39775a,a39779a,a39780a,a39781a,a39785a,a39786a,a39790a,a39791a,a39792a,a39796a,a39797a,a39801a,a39802a,a39803a,a39807a,a39808a,a39812a,a39813a,a39814a,a39818a,a39819a,a39823a,a39824a,a39825a,a39829a,a39830a,a39834a,a39835a,a39836a,a39840a,a39841a,a39845a,a39846a,a39847a,a39851a,a39852a,a39856a,a39857a,a39858a,a39862a,a39863a,a39867a,a39868a,a39869a,a39873a,a39874a,a39878a,a39879a,a39880a,a39884a,a39885a,a39889a,a39890a,a39891a,a39895a,a39896a,a39900a,a39901a,a39902a,a39906a,a39907a,a39911a,a39912a,a39913a,a39917a,a39918a,a39922a,a39923a,a39924a,a39928a,a39929a,a39933a,a39934a,a39935a,a39939a,a39940a,a39944a,a39945a,a39946a,a39950a,a39951a,a39955a,a39956a,a39957a,a39961a,a39962a,a39966a,a39967a,a39968a,a39972a,a39973a,a39977a,a39978a,a39979a,a39983a,a39984a,a39988a,a39989a,a39990a,a39994a,a39995a,a39999a,a40000a,a40001a,a40005a,a40006a,a40010a,a40011a,a40012a,a40016a,a40017a,a40021a,a40022a,a40023a,a40027a,a40028a,a40032a,a40033a,a40034a,a40038a,a40039a,a40043a,a40044a,a40045a,a40049a,a40050a,a40054a,a40055a,a40056a,a40060a,a40061a,a40065a,a40066a,a40067a,a40071a,a40072a,a40076a,a40077a,a40078a,a40082a,a40083a,a40087a,a40088a,a40089a,a40093a,a40094a,a40098a,a40099a,a40100a,a40104a,a40105a,a40109a,a40110a,a40111a,a40115a,a40116a,a40120a,a40121a,a40122a,a40126a,a40127a,a40131a,a40132a,a40133a,a40137a,a40138a,a40142a,a40143a,a40144a,a40148a,a40149a,a40153a,a40154a,a40155a,a40159a,a40160a,a40164a,a40165a,a40166a,a40170a,a40171a,a40175a,a40176a,a40177a,a40181a,a40182a,a40186a,a40187a,a40188a,a40192a,a40193a,a40197a,a40198a,a40199a,a40203a,a40204a,a40208a,a40209a,a40210a,a40214a,a40215a,a40219a,a40220a,a40221a,a40225a,a40226a,a40230a,a40231a,a40232a,a40236a,a40237a,a40241a,a40242a,a40243a,a40247a,a40248a,a40252a,a40253a,a40254a,a40258a,a40259a,a40263a,a40264a,a40265a,a40269a,a40270a,a40274a,a40275a,a40276a,a40280a,a40281a,a40285a,a40286a,a40287a,a40291a,a40292a,a40296a,a40297a,a40298a,a40302a,a40303a,a40307a,a40308a,a40309a,a40313a,a40314a,a40318a,a40319a,a40320a,a40324a,a40325a,a40329a,a40330a,a40331a,a40335a,a40336a,a40340a,a40341a,a40342a,a40346a,a40347a,a40351a,a40352a,a40353a,a40357a,a40358a,a40362a,a40363a,a40364a,a40368a,a40369a,a40373a,a40374a,a40375a,a40379a,a40380a,a40384a,a40385a,a40386a,a40390a,a40391a,a40395a,a40396a,a40397a,a40401a,a40402a,a40406a,a40407a,a40408a,a40412a,a40413a,a40417a,a40418a,a40419a,a40423a,a40424a,a40428a,a40429a,a40430a,a40434a,a40435a,a40439a,a40440a,a40441a,a40445a,a40446a,a40450a,a40451a,a40452a,a40456a,a40457a,a40461a,a40462a,a40463a,a40467a,a40468a,a40472a,a40473a,a40474a,a40478a,a40479a,a40483a,a40484a,a40485a,a40489a,a40490a,a40494a,a40495a,a40496a,a40500a,a40501a,a40505a,a40506a,a40507a,a40511a,a40512a,a40516a,a40517a,a40518a,a40522a,a40523a,a40527a,a40528a,a40529a,a40533a,a40534a,a40538a,a40539a,a40540a,a40544a,a40545a,a40549a,a40550a,a40551a,a40555a,a40556a,a40560a,a40561a,a40562a,a40566a,a40567a,a40571a,a40572a,a40573a,a40577a,a40578a,a40582a,a40583a,a40584a,a40588a,a40589a,a40593a,a40594a,a40595a,a40599a,a40600a,a40604a,a40605a,a40606a,a40610a,a40611a,a40615a,a40616a,a40617a,a40621a,a40622a,a40626a,a40627a,a40628a,a40632a,a40633a,a40637a,a40638a,a40639a,a40643a,a40644a,a40648a,a40649a,a40650a,a40654a,a40655a,a40659a,a40660a,a40661a,a40665a,a40666a,a40670a,a40671a,a40672a,a40676a,a40677a,a40681a,a40682a,a40683a,a40687a,a40688a,a40692a,a40693a,a40694a,a40698a,a40699a,a40703a,a40704a,a40705a,a40709a,a40710a,a40714a,a40715a,a40716a,a40720a,a40721a,a40725a,a40726a,a40727a,a40731a,a40732a,a40736a,a40737a,a40738a,a40742a,a40743a,a40747a,a40748a,a40749a,a40753a,a40754a,a40758a,a40759a,a40760a,a40764a,a40765a,a40769a,a40770a,a40771a,a40775a,a40776a,a40780a,a40781a,a40782a,a40786a,a40787a,a40791a,a40792a,a40793a,a40797a,a40798a,a40802a,a40803a,a40804a,a40808a,a40809a,a40813a,a40814a,a40815a,a40819a,a40820a,a40824a,a40825a,a40826a,a40830a,a40831a,a40835a,a40836a,a40837a,a40841a,a40842a,a40846a,a40847a,a40848a,a40852a,a40853a,a40857a,a40858a,a40859a,a40863a,a40864a,a40868a,a40869a,a40870a,a40874a,a40875a,a40879a,a40880a,a40881a,a40885a,a40886a,a40890a,a40891a,a40892a,a40896a,a40897a,a40901a,a40902a,a40903a,a40907a,a40908a,a40912a,a40913a,a40914a,a40918a,a40919a,a40923a,a40924a,a40925a,a40929a,a40930a,a40934a,a40935a,a40936a,a40940a,a40941a,a40945a,a40946a,a40947a,a40951a,a40952a,a40956a,a40957a,a40958a,a40962a,a40963a,a40967a,a40968a,a40969a,a40973a,a40974a,a40978a,a40979a,a40980a,a40984a,a40985a,a40989a,a40990a,a40991a,a40995a,a40996a,a41000a,a41001a,a41002a,a41006a,a41007a,a41011a,a41012a,a41013a,a41017a,a41018a,a41022a,a41023a,a41024a,a41028a,a41029a,a41033a,a41034a,a41035a,a41039a,a41040a,a41044a,a41045a,a41046a,a41050a,a41051a,a41055a,a41056a,a41057a,a41061a,a41062a,a41066a,a41067a,a41068a,a41072a,a41073a,a41077a,a41078a,a41079a,a41083a,a41084a,a41088a,a41089a,a41090a,a41094a,a41095a,a41099a,a41100a,a41101a,a41105a,a41106a,a41110a,a41111a,a41112a,a41116a,a41117a,a41121a,a41122a,a41123a,a41127a,a41128a,a41132a,a41133a,a41134a,a41138a,a41139a,a41143a,a41144a,a41145a,a41149a,a41150a,a41154a,a41155a,a41156a,a41160a,a41161a,a41165a,a41166a,a41167a,a41171a,a41172a,a41176a,a41177a,a41178a,a41182a,a41183a,a41187a,a41188a,a41189a,a41193a,a41194a,a41198a,a41199a,a41200a,a41204a,a41205a,a41209a,a41210a,a41211a,a41215a,a41216a,a41220a,a41221a,a41222a,a41226a,a41227a,a41231a,a41232a,a41233a,a41237a,a41238a,a41242a,a41243a,a41244a,a41248a,a41249a,a41253a,a41254a,a41255a,a41259a,a41260a,a41264a,a41265a,a41266a,a41270a,a41271a,a41275a,a41276a,a41277a,a41281a,a41282a,a41286a,a41287a,a41288a,a41292a,a41293a,a41297a,a41298a,a41299a,a41303a,a41304a,a41308a,a41309a,a41310a,a41314a,a41315a,a41319a,a41320a,a41321a,a41325a,a41326a,a41329a,a41332a,a41333a,a41334a,a41338a,a41339a,a41343a,a41344a,a41345a,a41349a,a41350a,a41353a,a41356a,a41357a,a41358a,a41362a,a41363a,a41367a,a41368a,a41369a,a41373a,a41374a,a41377a,a41380a,a41381a,a41382a,a41386a,a41387a,a41391a,a41392a,a41393a,a41397a,a41398a,a41401a,a41404a,a41405a,a41406a,a41410a,a41411a,a41415a,a41416a,a41417a,a41421a,a41422a,a41425a,a41428a,a41429a,a41430a,a41434a,a41435a,a41439a,a41440a,a41441a,a41445a,a41446a,a41449a,a41452a,a41453a,a41454a,a41458a,a41459a,a41463a,a41464a,a41465a,a41469a,a41470a,a41473a,a41476a,a41477a,a41478a,a41482a,a41483a,a41487a,a41488a,a41489a,a41493a,a41494a,a41497a,a41500a,a41501a,a41502a,a41506a,a41507a,a41511a,a41512a,a41513a,a41517a,a41518a,a41521a,a41524a,a41525a,a41526a,a41530a,a41531a,a41535a,a41536a,a41537a,a41541a,a41542a,a41545a,a41548a,a41549a,a41550a,a41554a,a41555a,a41559a,a41560a,a41561a,a41565a,a41566a,a41569a,a41572a,a41573a,a41574a,a41578a,a41579a,a41583a,a41584a,a41585a,a41589a,a41590a,a41593a,a41596a,a41597a,a41598a,a41602a,a41603a,a41607a,a41608a,a41609a,a41613a,a41614a,a41617a,a41620a,a41621a,a41622a,a41626a,a41627a,a41631a,a41632a,a41633a,a41637a,a41638a,a41641a,a41644a,a41645a,a41646a,a41650a,a41651a,a41655a,a41656a,a41657a,a41661a,a41662a,a41665a,a41668a,a41669a,a41670a,a41674a,a41675a,a41679a,a41680a,a41681a,a41685a,a41686a,a41689a,a41692a,a41693a,a41694a,a41698a,a41699a,a41703a,a41704a,a41705a,a41709a,a41710a,a41713a,a41716a,a41717a,a41718a,a41722a,a41723a,a41727a,a41728a,a41729a,a41733a,a41734a,a41737a,a41740a,a41741a,a41742a,a41746a,a41747a,a41751a,a41752a,a41753a,a41757a,a41758a,a41761a,a41764a,a41765a,a41766a,a41770a,a41771a,a41775a,a41776a,a41777a,a41781a,a41782a,a41785a,a41788a,a41789a,a41790a,a41794a,a41795a,a41799a,a41800a,a41801a,a41805a,a41806a,a41809a,a41812a,a41813a,a41814a,a41818a,a41819a,a41823a,a41824a,a41825a,a41829a,a41830a,a41833a,a41836a,a41837a,a41838a,a41842a,a41843a,a41847a,a41848a,a41849a,a41853a,a41854a,a41857a,a41860a,a41861a,a41862a,a41866a,a41867a,a41871a,a41872a,a41873a,a41877a,a41878a,a41881a,a41884a,a41885a,a41886a,a41890a,a41891a,a41895a,a41896a,a41897a,a41901a,a41902a,a41905a,a41908a,a41909a,a41910a,a41914a,a41915a,a41919a,a41920a,a41921a,a41925a,a41926a,a41929a,a41932a,a41933a,a41934a,a41938a,a41939a,a41943a,a41944a,a41945a,a41949a,a41950a,a41953a,a41956a,a41957a,a41958a,a41962a,a41963a,a41967a,a41968a,a41969a,a41973a,a41974a,a41977a,a41980a,a41981a,a41982a,a41986a,a41987a,a41991a,a41992a,a41993a,a41997a,a41998a,a42001a,a42004a,a42005a,a42006a,a42010a,a42011a,a42015a,a42016a,a42017a,a42021a,a42022a,a42025a,a42028a,a42029a,a42030a,a42034a,a42035a,a42039a,a42040a,a42041a,a42045a,a42046a,a42049a,a42052a,a42053a,a42054a,a42058a,a42059a,a42063a,a42064a,a42065a,a42069a,a42070a,a42073a,a42076a,a42077a,a42078a,a42082a,a42083a,a42087a,a42088a,a42089a,a42093a,a42094a,a42097a,a42100a,a42101a,a42102a,a42106a,a42107a,a42111a,a42112a,a42113a,a42117a,a42118a,a42121a,a42124a,a42125a,a42126a,a42130a,a42131a,a42135a,a42136a,a42137a,a42141a,a42142a,a42145a,a42148a,a42149a,a42150a,a42154a,a42155a,a42159a,a42160a,a42161a,a42165a,a42166a,a42169a,a42172a,a42173a,a42174a,a42178a,a42179a,a42183a,a42184a,a42185a,a42189a,a42190a,a42193a,a42196a,a42197a,a42198a,a42202a,a42203a,a42207a,a42208a,a42209a,a42213a,a42214a,a42217a,a42220a,a42221a,a42222a,a42226a,a42227a,a42231a,a42232a,a42233a,a42237a,a42238a,a42241a,a42244a,a42245a,a42246a,a42250a,a42251a,a42255a,a42256a,a42257a,a42261a,a42262a,a42265a,a42268a,a42269a,a42270a,a42274a,a42275a,a42279a,a42280a,a42281a,a42285a,a42286a,a42289a,a42292a,a42293a,a42294a,a42298a,a42299a,a42303a,a42304a,a42305a,a42309a,a42310a,a42313a,a42316a,a42317a,a42318a,a42322a,a42323a,a42327a,a42328a,a42329a,a42333a,a42334a,a42337a,a42340a,a42341a,a42342a,a42346a,a42347a,a42351a,a42352a,a42353a,a42357a,a42358a,a42361a,a42364a,a42365a,a42366a,a42370a,a42371a,a42375a,a42376a,a42377a,a42381a,a42382a,a42385a,a42388a,a42389a,a42390a,a42394a,a42395a,a42399a,a42400a,a42401a,a42405a,a42406a,a42409a,a42412a,a42413a,a42414a,a42418a,a42419a,a42423a,a42424a,a42425a,a42429a,a42430a,a42433a,a42436a,a42437a,a42438a,a42442a,a42443a,a42447a,a42448a,a42449a,a42453a,a42454a,a42457a,a42460a,a42461a,a42462a,a42466a,a42467a,a42471a,a42472a,a42473a,a42477a,a42478a,a42481a,a42484a,a42485a,a42486a,a42490a,a42491a,a42495a,a42496a,a42497a,a42501a,a42502a,a42505a,a42508a,a42509a,a42510a,a42514a,a42515a,a42519a,a42520a,a42521a,a42525a,a42526a,a42529a,a42532a,a42533a,a42534a,a42538a,a42539a,a42543a,a42544a,a42545a,a42549a,a42550a,a42553a,a42556a,a42557a,a42558a,a42562a,a42563a,a42567a,a42568a,a42569a,a42573a,a42574a,a42577a,a42580a,a42581a,a42582a,a42586a,a42587a,a42591a,a42592a,a42593a,a42597a,a42598a,a42601a,a42604a,a42605a,a42606a,a42610a,a42611a,a42615a,a42616a,a42617a,a42621a,a42622a,a42625a,a42628a,a42629a,a42630a,a42634a,a42635a,a42639a,a42640a,a42641a,a42645a,a42646a,a42649a,a42652a,a42653a,a42654a,a42658a,a42659a,a42663a,a42664a,a42665a,a42669a,a42670a,a42673a,a42676a,a42677a,a42678a,a42682a,a42683a,a42687a,a42688a,a42689a,a42693a,a42694a,a42697a,a42700a,a42701a,a42702a,a42706a,a42707a,a42711a,a42712a,a42713a,a42717a,a42718a,a42721a,a42724a,a42725a,a42726a,a42730a,a42731a,a42735a,a42736a,a42737a,a42741a,a42742a,a42745a,a42748a,a42749a,a42750a,a42754a,a42755a,a42759a,a42760a,a42761a,a42765a,a42766a,a42769a,a42772a,a42773a,a42774a,a42778a,a42779a,a42783a,a42784a,a42785a,a42789a,a42790a,a42793a,a42796a,a42797a,a42798a,a42802a,a42803a,a42807a,a42808a,a42809a,a42813a,a42814a,a42817a,a42820a,a42821a,a42822a,a42826a,a42827a,a42831a,a42832a,a42833a,a42837a,a42838a,a42841a,a42844a,a42845a,a42846a,a42850a,a42851a,a42855a,a42856a,a42857a,a42861a,a42862a,a42865a,a42868a,a42869a,a42870a,a42874a,a42875a,a42879a,a42880a,a42881a,a42885a,a42886a,a42889a,a42892a,a42893a,a42894a,a42898a,a42899a,a42903a,a42904a,a42905a,a42909a,a42910a,a42913a,a42916a,a42917a,a42918a,a42922a,a42923a,a42927a,a42928a,a42929a,a42933a,a42934a,a42937a,a42940a,a42941a,a42942a,a42946a,a42947a,a42951a,a42952a,a42953a,a42957a,a42958a,a42961a,a42964a,a42965a,a42966a,a42970a,a42971a,a42975a,a42976a,a42977a,a42981a,a42982a,a42985a,a42988a,a42989a,a42990a,a42994a,a42995a,a42999a,a43000a,a43001a,a43005a,a43006a,a43009a,a43012a,a43013a,a43014a,a43018a,a43019a,a43023a,a43024a,a43025a,a43029a,a43030a,a43033a,a43036a,a43037a,a43038a,a43042a,a43043a,a43047a,a43048a,a43049a,a43053a,a43054a,a43057a,a43060a,a43061a,a43062a,a43066a,a43067a,a43071a,a43072a,a43073a,a43077a,a43078a,a43081a,a43084a,a43085a,a43086a,a43090a,a43091a,a43095a,a43096a,a43097a,a43101a,a43102a,a43105a,a43108a,a43109a,a43110a,a43114a,a43115a,a43119a,a43120a,a43121a,a43125a,a43126a,a43129a,a43132a,a43133a,a43134a,a43138a,a43139a,a43143a,a43144a,a43145a,a43149a,a43150a,a43153a,a43156a,a43157a,a43158a,a43162a,a43163a,a43167a,a43168a,a43169a,a43173a,a43174a,a43177a,a43180a,a43181a,a43182a,a43186a,a43187a,a43191a,a43192a,a43193a,a43197a,a43198a,a43201a,a43204a,a43205a,a43206a,a43210a,a43211a,a43215a,a43216a,a43217a,a43221a,a43222a,a43225a,a43228a,a43229a,a43230a,a43234a,a43235a,a43239a,a43240a,a43241a,a43245a,a43246a,a43249a,a43252a,a43253a,a43254a,a43258a,a43259a,a43263a,a43264a,a43265a,a43269a,a43270a,a43273a,a43276a,a43277a,a43278a,a43282a,a43283a,a43287a,a43288a,a43289a,a43293a,a43294a,a43297a,a43300a,a43301a,a43302a,a43306a,a43307a,a43311a,a43312a,a43313a,a43317a,a43318a,a43321a,a43324a,a43325a,a43326a,a43330a,a43331a,a43335a,a43336a,a43337a,a43341a,a43342a,a43345a,a43348a,a43349a,a43350a,a43354a,a43355a,a43359a,a43360a,a43361a,a43365a,a43366a,a43369a,a43372a,a43373a,a43374a,a43378a,a43379a,a43383a,a43384a,a43385a,a43389a,a43390a,a43393a,a43396a,a43397a,a43398a,a43402a,a43403a,a43407a,a43408a,a43409a,a43413a,a43414a,a43417a,a43420a,a43421a,a43422a,a43426a,a43427a,a43431a,a43432a,a43433a,a43437a,a43438a,a43441a,a43444a,a43445a,a43446a,a43450a,a43451a,a43455a,a43456a,a43457a,a43461a,a43462a,a43465a,a43468a,a43469a,a43470a,a43474a,a43475a,a43479a,a43480a,a43481a,a43485a,a43486a,a43489a,a43492a,a43493a,a43494a,a43498a,a43499a,a43503a,a43504a,a43505a,a43509a,a43510a,a43513a,a43516a,a43517a,a43518a,a43522a,a43523a,a43527a,a43528a,a43529a,a43533a,a43534a,a43537a,a43540a,a43541a,a43542a,a43546a,a43547a,a43551a,a43552a,a43553a,a43557a,a43558a,a43561a,a43564a,a43565a,a43566a,a43570a,a43571a,a43575a,a43576a,a43577a,a43581a,a43582a,a43585a,a43588a,a43589a,a43590a,a43594a,a43595a,a43599a,a43600a,a43601a,a43605a,a43606a,a43609a,a43612a,a43613a,a43614a,a43618a,a43619a,a43623a,a43624a,a43625a,a43629a,a43630a,a43633a,a43636a,a43637a,a43638a,a43642a,a43643a,a43647a,a43648a,a43649a,a43653a,a43654a,a43657a,a43660a,a43661a,a43662a,a43666a,a43667a,a43671a,a43672a,a43673a,a43677a,a43678a,a43681a,a43684a,a43685a,a43686a,a43690a,a43691a,a43695a,a43696a,a43697a,a43701a,a43702a,a43705a,a43708a,a43709a,a43710a,a43714a,a43715a,a43719a,a43720a,a43721a,a43725a,a43726a,a43729a,a43732a,a43733a,a43734a,a43738a,a43739a,a43743a,a43744a,a43745a,a43749a,a43750a,a43753a,a43756a,a43757a,a43758a,a43762a,a43763a,a43767a,a43768a,a43769a,a43773a,a43774a,a43777a,a43780a,a43781a,a43782a,a43786a,a43787a,a43791a,a43792a,a43793a,a43797a,a43798a,a43801a,a43804a,a43805a,a43806a,a43810a,a43811a,a43815a,a43816a,a43817a,a43821a,a43822a,a43825a,a43828a,a43829a,a43830a,a43834a,a43835a,a43839a,a43840a,a43841a,a43845a,a43846a,a43849a,a43852a,a43853a,a43854a,a43858a,a43859a,a43863a,a43864a,a43865a,a43869a,a43870a,a43873a,a43876a,a43877a,a43878a,a43882a,a43883a,a43887a,a43888a,a43889a,a43893a,a43894a,a43897a,a43900a,a43901a,a43902a,a43906a,a43907a,a43911a,a43912a,a43913a,a43917a,a43918a,a43921a,a43924a,a43925a,a43926a,a43930a,a43931a,a43935a,a43936a,a43937a,a43941a,a43942a,a43945a,a43948a,a43949a,a43950a,a43954a,a43955a,a43959a,a43960a,a43961a,a43965a,a43966a,a43969a,a43972a,a43973a,a43974a,a43978a,a43979a,a43983a,a43984a,a43985a,a43989a,a43990a,a43993a,a43996a,a43997a,a43998a,a44002a,a44003a,a44007a,a44008a,a44009a,a44013a,a44014a,a44017a,a44020a,a44021a,a44022a,a44026a,a44027a,a44031a,a44032a,a44033a,a44037a,a44038a,a44041a,a44044a,a44045a,a44046a,a44050a,a44051a,a44055a,a44056a,a44057a,a44061a,a44062a,a44065a,a44068a,a44069a,a44070a,a44074a,a44075a,a44079a,a44080a,a44081a,a44085a,a44086a,a44089a,a44092a,a44093a,a44094a,a44098a,a44099a,a44103a,a44104a,a44105a,a44109a,a44110a,a44113a,a44116a,a44117a,a44118a,a44122a,a44123a,a44127a,a44128a,a44129a,a44133a,a44134a,a44137a,a44140a,a44141a,a44142a,a44146a,a44147a,a44151a,a44152a,a44153a,a44157a,a44158a,a44161a,a44164a,a44165a,a44166a,a44170a,a44171a,a44175a,a44176a,a44177a,a44181a,a44182a,a44185a,a44188a,a44189a,a44190a,a44194a,a44195a,a44199a,a44200a,a44201a,a44205a,a44206a,a44209a,a44212a,a44213a,a44214a,a44218a,a44219a,a44223a,a44224a,a44225a,a44229a,a44230a,a44233a,a44236a,a44237a,a44238a,a44242a,a44243a,a44247a,a44248a,a44249a,a44253a,a44254a,a44257a,a44260a,a44261a,a44262a,a44266a,a44267a,a44271a,a44272a,a44273a,a44277a,a44278a,a44281a,a44284a,a44285a,a44286a,a44290a,a44291a,a44295a,a44296a,a44297a,a44301a,a44302a,a44305a,a44308a,a44309a,a44310a,a44314a,a44315a,a44319a,a44320a,a44321a,a44325a,a44326a,a44329a,a44332a,a44333a,a44334a,a44338a,a44339a,a44343a,a44344a,a44345a,a44349a,a44350a,a44353a,a44356a,a44357a,a44358a,a44362a,a44363a,a44367a,a44368a,a44369a,a44373a,a44374a,a44377a,a44380a,a44381a,a44382a,a44386a,a44387a,a44391a,a44392a,a44393a,a44397a,a44398a,a44401a,a44404a,a44405a,a44406a,a44410a,a44411a,a44415a,a44416a,a44417a,a44421a,a44422a,a44425a,a44428a,a44429a,a44430a,a44434a,a44435a,a44439a,a44440a,a44441a,a44445a,a44446a,a44449a,a44452a,a44453a,a44454a,a44458a,a44459a,a44463a,a44464a,a44465a,a44469a,a44470a,a44473a,a44476a,a44477a,a44478a,a44482a,a44483a,a44487a,a44488a,a44489a,a44493a,a44494a,a44497a,a44500a,a44501a,a44502a,a44506a,a44507a,a44511a,a44512a,a44513a,a44517a,a44518a,a44521a,a44524a,a44525a,a44526a,a44530a,a44531a,a44535a,a44536a,a44537a,a44541a,a44542a,a44545a,a44548a,a44549a,a44550a,a44554a,a44555a,a44559a,a44560a,a44561a,a44565a,a44566a,a44569a,a44572a,a44573a,a44574a,a44578a,a44579a,a44583a,a44584a,a44585a,a44589a,a44590a,a44593a,a44596a,a44597a,a44598a,a44602a,a44603a,a44607a,a44608a,a44609a,a44613a,a44614a,a44617a,a44620a,a44621a,a44622a,a44626a,a44627a,a44631a,a44632a,a44633a,a44637a,a44638a,a44641a,a44644a,a44645a,a44646a,a44650a,a44651a,a44655a,a44656a,a44657a,a44661a,a44662a,a44665a,a44668a,a44669a,a44670a,a44674a,a44675a,a44679a,a44680a,a44681a,a44685a,a44686a,a44689a,a44692a,a44693a,a44694a,a44698a,a44699a,a44703a,a44704a,a44705a,a44709a,a44710a,a44713a,a44716a,a44717a,a44718a,a44722a,a44723a,a44727a,a44728a,a44729a,a44733a,a44734a,a44737a,a44740a,a44741a,a44742a,a44746a,a44747a,a44751a,a44752a,a44753a,a44757a,a44758a,a44761a,a44764a,a44765a,a44766a,a44770a,a44771a,a44775a,a44776a,a44777a,a44781a,a44782a,a44785a,a44788a,a44789a,a44790a,a44794a,a44795a,a44799a,a44800a,a44801a,a44805a,a44806a,a44809a,a44812a,a44813a,a44814a,a44818a,a44819a,a44823a,a44824a,a44825a,a44829a,a44830a,a44833a,a44836a,a44837a,a44838a,a44842a,a44843a,a44847a,a44848a,a44849a,a44853a,a44854a,a44857a,a44860a,a44861a,a44862a,a44866a,a44867a,a44871a,a44872a,a44873a,a44877a,a44878a,a44881a,a44884a,a44885a,a44886a,a44890a,a44891a,a44895a,a44896a,a44897a,a44901a,a44902a,a44905a,a44908a,a44909a,a44910a,a44914a,a44915a,a44919a,a44920a,a44921a,a44925a,a44926a,a44929a,a44932a,a44933a,a44934a,a44938a,a44939a,a44943a,a44944a,a44945a,a44949a,a44950a,a44953a,a44956a,a44957a,a44958a,a44962a,a44963a,a44967a,a44968a,a44969a,a44973a,a44974a,a44977a,a44980a,a44981a,a44982a,a44986a,a44987a,a44991a,a44992a,a44993a,a44997a,a44998a,a45001a,a45004a,a45005a,a45006a,a45010a,a45011a,a45015a,a45016a,a45017a,a45021a,a45022a,a45025a,a45028a,a45029a,a45030a,a45034a,a45035a,a45039a,a45040a,a45041a,a45045a,a45046a,a45049a,a45052a,a45053a,a45054a,a45058a,a45059a,a45063a,a45064a,a45065a,a45069a,a45070a,a45073a,a45076a,a45077a,a45078a,a45082a,a45083a,a45087a,a45088a,a45089a,a45093a,a45094a,a45097a,a45100a,a45101a,a45102a,a45106a,a45107a,a45111a,a45112a,a45113a,a45117a,a45118a,a45121a,a45124a,a45125a,a45126a,a45130a,a45131a,a45135a,a45136a,a45137a,a45141a,a45142a,a45145a,a45148a,a45149a,a45150a,a45154a,a45155a,a45159a,a45160a,a45161a,a45165a,a45166a,a45169a,a45172a,a45173a,a45174a,a45178a,a45179a,a45183a,a45184a,a45185a,a45189a,a45190a,a45193a,a45196a,a45197a,a45198a,a45202a,a45203a,a45207a,a45208a,a45209a,a45213a,a45214a,a45217a,a45220a,a45221a,a45222a,a45226a,a45227a,a45231a,a45232a,a45233a,a45237a,a45238a,a45241a,a45244a,a45245a,a45246a,a45250a,a45251a,a45255a,a45256a,a45257a,a45261a,a45262a,a45265a,a45268a,a45269a,a45270a,a45274a,a45275a,a45279a,a45280a,a45281a,a45285a,a45286a,a45289a,a45292a,a45293a,a45294a,a45298a,a45299a,a45303a,a45304a,a45305a,a45309a,a45310a,a45313a,a45316a,a45317a,a45318a,a45322a,a45323a,a45327a,a45328a,a45329a,a45333a,a45334a,a45337a,a45340a,a45341a,a45342a,a45346a,a45347a,a45351a,a45352a,a45353a,a45357a,a45358a,a45361a,a45364a,a45365a,a45366a,a45370a,a45371a,a45375a,a45376a,a45377a,a45381a,a45382a,a45385a,a45388a,a45389a,a45390a,a45394a,a45395a,a45399a,a45400a,a45401a,a45405a,a45406a,a45409a,a45412a,a45413a,a45414a,a45418a,a45419a,a45423a,a45424a,a45425a,a45429a,a45430a,a45433a,a45436a,a45437a,a45438a,a45442a,a45443a,a45447a,a45448a,a45449a,a45453a,a45454a,a45457a,a45460a,a45461a,a45462a,a45466a,a45467a,a45471a,a45472a,a45473a,a45477a,a45478a,a45481a,a45484a,a45485a,a45486a,a45490a,a45491a,a45495a,a45496a,a45497a,a45501a,a45502a,a45505a,a45508a,a45509a,a45510a,a45514a,a45515a,a45519a,a45520a,a45521a,a45525a,a45526a,a45529a,a45532a,a45533a,a45534a,a45538a,a45539a,a45543a,a45544a,a45545a,a45549a,a45550a,a45553a,a45556a,a45557a,a45558a,a45562a,a45563a,a45567a,a45568a,a45569a,a45573a,a45574a,a45577a,a45580a,a45581a,a45582a,a45586a,a45587a,a45591a,a45592a,a45593a,a45597a,a45598a,a45601a,a45604a,a45605a,a45606a,a45610a,a45611a,a45615a,a45616a,a45617a,a45621a,a45622a,a45625a,a45628a,a45629a,a45630a,a45634a,a45635a,a45639a,a45640a,a45641a,a45645a,a45646a,a45649a,a45652a,a45653a,a45654a,a45658a,a45659a,a45663a,a45664a,a45665a,a45669a,a45670a,a45673a,a45676a,a45677a,a45678a,a45682a,a45683a,a45687a,a45688a,a45689a,a45693a,a45694a,a45697a,a45700a,a45701a,a45702a,a45706a,a45707a,a45711a,a45712a,a45713a,a45717a,a45718a,a45721a,a45724a,a45725a,a45726a,a45730a,a45731a,a45735a,a45736a,a45737a,a45741a,a45742a,a45745a,a45748a,a45749a,a45750a,a45754a,a45755a,a45759a,a45760a,a45761a,a45765a,a45766a,a45769a,a45772a,a45773a,a45774a,a45778a,a45779a,a45783a,a45784a,a45785a,a45789a,a45790a,a45793a,a45796a,a45797a,a45798a,a45802a,a45803a,a45807a,a45808a,a45809a,a45813a,a45814a,a45817a,a45820a,a45821a,a45822a,a45826a,a45827a,a45831a,a45832a,a45833a,a45837a,a45838a,a45841a,a45844a,a45845a,a45846a,a45850a,a45851a,a45855a,a45856a,a45857a,a45861a,a45862a,a45865a,a45868a,a45869a,a45870a,a45874a,a45875a,a45879a,a45880a,a45881a,a45885a,a45886a,a45889a,a45892a,a45893a,a45894a,a45898a,a45899a,a45903a,a45904a,a45905a,a45909a,a45910a,a45913a,a45916a,a45917a,a45918a,a45922a,a45923a,a45927a,a45928a,a45929a,a45933a,a45934a,a45937a,a45940a,a45941a,a45942a,a45946a,a45947a,a45951a,a45952a,a45953a,a45957a,a45958a,a45961a,a45964a,a45965a,a45966a,a45970a,a45971a,a45975a,a45976a,a45977a,a45981a,a45982a,a45985a,a45988a,a45989a,a45990a,a45994a,a45995a,a45999a,a46000a,a46001a,a46005a,a46006a,a46009a,a46012a,a46013a,a46014a,a46018a,a46019a,a46023a,a46024a,a46025a,a46029a,a46030a,a46033a,a46036a,a46037a,a46038a,a46042a,a46043a,a46047a,a46048a,a46049a,a46053a,a46054a,a46057a,a46060a,a46061a,a46062a,a46066a,a46067a,a46071a,a46072a,a46073a,a46077a,a46078a,a46081a,a46084a,a46085a,a46086a,a46090a,a46091a,a46095a,a46096a,a46097a,a46101a,a46102a,a46105a,a46108a,a46109a,a46110a,a46114a,a46115a,a46119a,a46120a,a46121a,a46125a,a46126a,a46129a,a46132a,a46133a,a46134a,a46138a,a46139a,a46143a,a46144a,a46145a,a46149a,a46150a,a46153a,a46156a,a46157a,a46158a,a46162a,a46163a,a46167a,a46168a,a46169a,a46173a,a46174a,a46177a,a46180a,a46181a,a46182a,a46186a,a46187a,a46191a,a46192a,a46193a,a46197a,a46198a,a46201a,a46204a,a46205a,a46206a,a46210a,a46211a,a46215a,a46216a,a46217a,a46221a,a46222a,a46225a,a46228a,a46229a,a46230a,a46234a,a46235a,a46239a,a46240a,a46241a,a46245a,a46246a,a46249a,a46252a,a46253a,a46254a,a46258a,a46259a,a46263a,a46264a,a46265a,a46269a,a46270a,a46273a,a46276a,a46277a,a46278a,a46282a,a46283a,a46287a,a46288a,a46289a,a46293a,a46294a,a46297a,a46300a,a46301a,a46302a,a46306a,a46307a,a46311a,a46312a,a46313a,a46317a,a46318a,a46321a,a46324a,a46325a,a46326a,a46330a,a46331a,a46335a,a46336a,a46337a,a46341a,a46342a,a46345a,a46348a,a46349a,a46350a,a46354a,a46355a,a46359a,a46360a,a46361a,a46365a,a46366a,a46369a,a46372a,a46373a,a46374a,a46378a,a46379a,a46383a,a46384a,a46385a,a46389a,a46390a,a46393a,a46396a,a46397a,a46398a,a46402a,a46403a,a46407a,a46408a,a46409a,a46413a,a46414a,a46417a,a46420a,a46421a,a46422a,a46426a,a46427a,a46431a,a46432a,a46433a,a46437a,a46438a,a46441a,a46444a,a46445a,a46446a,a46450a,a46451a,a46455a,a46456a,a46457a,a46461a,a46462a,a46465a,a46468a,a46469a,a46470a,a46474a,a46475a,a46479a,a46480a,a46481a,a46485a,a46486a,a46489a,a46492a,a46493a,a46494a,a46498a,a46499a,a46503a,a46504a,a46505a,a46509a,a46510a,a46513a,a46516a,a46517a,a46518a,a46522a,a46523a,a46527a,a46528a,a46529a,a46533a,a46534a,a46537a,a46540a,a46541a,a46542a,a46546a,a46547a,a46551a,a46552a,a46553a,a46557a,a46558a,a46561a,a46564a,a46565a,a46566a,a46570a,a46571a,a46575a,a46576a,a46577a,a46581a,a46582a,a46585a,a46588a,a46589a,a46590a,a46594a,a46595a,a46599a,a46600a,a46601a,a46605a,a46606a,a46609a,a46612a,a46613a,a46614a,a46618a,a46619a,a46623a,a46624a,a46625a,a46629a,a46630a,a46633a,a46636a,a46637a,a46638a,a46642a,a46643a,a46647a,a46648a,a46649a,a46653a,a46654a,a46657a,a46660a,a46661a,a46662a,a46666a,a46667a,a46671a,a46672a,a46673a,a46677a,a46678a,a46681a,a46684a,a46685a,a46686a,a46690a,a46691a,a46695a,a46696a,a46697a,a46701a,a46702a,a46705a,a46708a,a46709a,a46710a,a46714a,a46715a,a46719a,a46720a,a46721a,a46725a,a46726a,a46729a,a46732a,a46733a,a46734a,a46738a,a46739a,a46743a,a46744a,a46745a,a46749a,a46750a,a46753a,a46756a,a46757a,a46758a,a46762a,a46763a,a46767a,a46768a,a46769a,a46773a,a46774a,a46777a,a46780a,a46781a,a46782a,a46786a,a46787a,a46791a,a46792a,a46793a,a46797a,a46798a,a46801a,a46804a,a46805a,a46806a,a46810a,a46811a,a46815a,a46816a,a46817a,a46821a,a46822a,a46825a,a46828a,a46829a,a46830a,a46834a,a46835a,a46839a,a46840a,a46841a,a46845a,a46846a,a46849a,a46852a,a46853a,a46854a,a46858a,a46859a,a46863a,a46864a,a46865a,a46869a,a46870a,a46873a,a46876a,a46877a,a46878a,a46882a,a46883a,a46887a,a46888a,a46889a,a46893a,a46894a,a46897a,a46900a,a46901a,a46902a,a46906a,a46907a,a46911a,a46912a,a46913a,a46917a,a46918a,a46921a,a46924a,a46925a,a46926a,a46930a,a46931a,a46935a,a46936a,a46937a,a46941a,a46942a,a46945a,a46948a,a46949a,a46950a,a46954a,a46955a,a46959a,a46960a,a46961a,a46965a,a46966a,a46969a,a46972a,a46973a,a46974a,a46978a,a46979a,a46983a,a46984a,a46985a,a46989a,a46990a,a46993a,a46996a,a46997a,a46998a,a47002a,a47003a,a47007a,a47008a,a47009a,a47013a,a47014a,a47017a,a47020a,a47021a,a47022a,a47026a,a47027a,a47031a,a47032a,a47033a,a47037a,a47038a,a47041a,a47044a,a47045a,a47046a,a47050a,a47051a,a47055a,a47056a,a47057a,a47061a,a47062a,a47065a,a47068a,a47069a,a47070a,a47074a,a47075a,a47079a,a47080a,a47081a,a47085a,a47086a,a47089a,a47092a,a47093a,a47094a,a47098a,a47099a,a47103a,a47104a,a47105a,a47109a,a47110a,a47113a,a47116a,a47117a,a47118a,a47122a,a47123a,a47127a,a47128a,a47129a,a47133a,a47134a,a47137a,a47140a,a47141a,a47142a,a47146a,a47147a,a47151a,a47152a,a47153a,a47157a,a47158a,a47161a,a47164a,a47165a,a47166a,a47170a,a47171a,a47175a,a47176a,a47177a,a47181a,a47182a,a47185a,a47188a,a47189a,a47190a,a47194a,a47195a,a47199a,a47200a,a47201a,a47205a,a47206a,a47209a,a47212a,a47213a,a47214a,a47218a,a47219a,a47223a,a47224a,a47225a,a47229a,a47230a,a47233a,a47236a,a47237a,a47238a,a47242a,a47243a,a47247a,a47248a,a47249a,a47253a,a47254a,a47257a,a47260a,a47261a,a47262a,a47266a,a47267a,a47271a,a47272a,a47273a,a47277a,a47278a,a47281a,a47284a,a47285a,a47286a,a47290a,a47291a,a47295a,a47296a,a47297a,a47301a,a47302a,a47305a,a47308a,a47309a,a47310a,a47314a,a47315a,a47319a,a47320a,a47321a,a47325a,a47326a,a47329a,a47332a,a47333a,a47334a,a47338a,a47339a,a47343a,a47344a,a47345a,a47349a,a47350a,a47353a,a47356a,a47357a,a47358a,a47362a,a47363a,a47367a,a47368a,a47369a,a47373a,a47374a,a47377a,a47380a,a47381a,a47382a,a47386a,a47387a,a47391a,a47392a,a47393a,a47397a,a47398a,a47401a,a47404a,a47405a,a47406a,a47410a,a47411a,a47415a,a47416a,a47417a,a47421a,a47422a,a47425a,a47428a,a47429a,a47430a,a47434a,a47435a,a47439a,a47440a,a47441a,a47445a,a47446a,a47449a,a47452a,a47453a,a47454a,a47458a,a47459a,a47463a,a47464a,a47465a,a47469a,a47470a,a47473a,a47476a,a47477a,a47478a,a47482a,a47483a,a47487a,a47488a,a47489a,a47493a,a47494a,a47497a,a47500a,a47501a,a47502a,a47506a,a47507a,a47511a,a47512a,a47513a,a47517a,a47518a,a47521a,a47524a,a47525a,a47526a,a47530a,a47531a,a47535a,a47536a,a47537a,a47541a,a47542a,a47545a,a47548a,a47549a,a47550a,a47554a,a47555a,a47559a,a47560a,a47561a,a47565a,a47566a,a47569a,a47572a,a47573a,a47574a,a47578a,a47579a,a47583a,a47584a,a47585a,a47589a,a47590a,a47593a,a47596a,a47597a,a47598a,a47602a,a47603a,a47607a,a47608a,a47609a,a47613a,a47614a,a47617a,a47620a,a47621a,a47622a,a47626a,a47627a,a47631a,a47632a,a47633a,a47637a,a47638a,a47641a,a47644a,a47645a,a47646a,a47650a,a47651a,a47655a,a47656a,a47657a,a47661a,a47662a,a47665a,a47668a,a47669a,a47670a,a47674a,a47675a,a47679a,a47680a,a47681a,a47685a,a47686a,a47689a,a47692a,a47693a,a47694a,a47698a,a47699a,a47703a,a47704a,a47705a,a47709a,a47710a,a47713a,a47716a,a47717a,a47718a,a47722a,a47723a,a47727a,a47728a,a47729a,a47733a,a47734a,a47737a,a47740a,a47741a,a47742a,a47746a,a47747a,a47751a,a47752a,a47753a,a47757a,a47758a,a47761a,a47764a,a47765a,a47766a,a47770a,a47771a,a47775a,a47776a,a47777a,a47781a,a47782a,a47785a,a47788a,a47789a,a47790a,a47794a,a47795a,a47799a,a47800a,a47801a,a47805a,a47806a,a47809a,a47812a,a47813a,a47814a,a47818a,a47819a,a47823a,a47824a,a47825a,a47829a,a47830a,a47833a,a47836a,a47837a,a47838a,a47842a,a47843a,a47847a,a47848a,a47849a,a47853a,a47854a,a47857a,a47860a,a47861a,a47862a,a47866a,a47867a,a47871a,a47872a,a47873a,a47877a,a47878a,a47881a,a47884a,a47885a,a47886a,a47890a,a47891a,a47895a,a47896a,a47897a,a47901a,a47902a,a47905a,a47908a,a47909a,a47910a,a47914a,a47915a,a47919a,a47920a,a47921a,a47925a,a47926a,a47929a,a47932a,a47933a,a47934a,a47938a,a47939a,a47943a,a47944a,a47945a,a47949a,a47950a,a47953a,a47956a,a47957a,a47958a,a47962a,a47963a,a47967a,a47968a,a47969a,a47973a,a47974a,a47977a,a47980a,a47981a,a47982a,a47986a,a47987a,a47991a,a47992a,a47993a,a47997a,a47998a,a48001a,a48004a,a48005a,a48006a,a48010a,a48011a,a48015a,a48016a,a48017a,a48021a,a48022a,a48025a,a48028a,a48029a,a48030a,a48034a,a48035a,a48039a,a48040a,a48041a,a48045a,a48046a,a48049a,a48052a,a48053a,a48054a,a48058a,a48059a,a48063a,a48064a,a48065a,a48069a,a48070a,a48073a,a48076a,a48077a,a48078a,a48082a,a48083a,a48087a,a48088a,a48089a,a48093a,a48094a,a48097a,a48100a,a48101a,a48102a,a48106a,a48107a,a48111a,a48112a,a48113a,a48117a,a48118a,a48121a,a48124a,a48125a,a48126a,a48130a,a48131a,a48135a,a48136a,a48137a,a48141a,a48142a,a48145a,a48148a,a48149a,a48150a,a48154a,a48155a,a48159a,a48160a,a48161a,a48165a,a48166a,a48169a,a48172a,a48173a,a48174a,a48178a,a48179a,a48183a,a48184a,a48185a,a48189a,a48190a,a48193a,a48196a,a48197a,a48198a,a48202a,a48203a,a48207a,a48208a,a48209a,a48213a,a48214a,a48217a,a48220a,a48221a,a48222a,a48226a,a48227a,a48231a,a48232a,a48233a,a48237a,a48238a,a48241a,a48244a,a48245a,a48246a,a48250a,a48251a,a48255a,a48256a,a48257a,a48261a,a48262a,a48265a,a48268a,a48269a,a48270a,a48274a,a48275a,a48279a,a48280a,a48281a,a48285a,a48286a,a48289a,a48292a,a48293a,a48294a,a48298a,a48299a,a48303a,a48304a,a48305a,a48309a,a48310a,a48313a,a48316a,a48317a,a48318a,a48322a,a48323a,a48327a,a48328a,a48329a,a48333a,a48334a,a48337a,a48340a,a48341a,a48342a,a48346a,a48347a,a48351a,a48352a,a48353a,a48357a,a48358a,a48361a,a48364a,a48365a,a48366a,a48370a,a48371a,a48375a,a48376a,a48377a,a48381a,a48382a,a48385a,a48388a,a48389a,a48390a,a48394a,a48395a,a48399a,a48400a,a48401a,a48405a,a48406a,a48409a,a48412a,a48413a,a48414a,a48418a,a48419a,a48423a,a48424a,a48425a,a48429a,a48430a,a48433a,a48436a,a48437a,a48438a,a48442a,a48443a,a48447a,a48448a,a48449a,a48453a,a48454a,a48457a,a48460a,a48461a,a48462a,a48466a,a48467a,a48471a,a48472a,a48473a,a48477a,a48478a,a48481a,a48484a,a48485a,a48486a,a48490a,a48491a,a48495a,a48496a,a48497a,a48501a,a48502a,a48505a,a48508a,a48509a,a48510a,a48514a,a48515a,a48519a,a48520a,a48521a,a48525a,a48526a,a48529a,a48532a,a48533a,a48534a,a48538a,a48539a,a48543a,a48544a,a48545a,a48549a,a48550a,a48553a,a48556a,a48557a,a48558a,a48562a,a48563a,a48567a,a48568a,a48569a,a48573a,a48574a,a48577a,a48580a,a48581a,a48582a,a48586a,a48587a,a48591a,a48592a,a48593a,a48597a,a48598a,a48601a,a48604a,a48605a,a48606a,a48610a,a48611a,a48615a,a48616a,a48617a,a48621a,a48622a,a48625a,a48628a,a48629a,a48630a,a48634a,a48635a,a48639a,a48640a,a48641a,a48645a,a48646a,a48649a,a48652a,a48653a,a48654a,a48658a,a48659a,a48663a,a48664a,a48665a,a48669a,a48670a,a48673a,a48676a,a48677a,a48678a,a48682a,a48683a,a48687a,a48688a,a48689a,a48693a,a48694a,a48697a,a48700a,a48701a,a48702a,a48706a,a48707a,a48711a,a48712a,a48713a,a48717a,a48718a,a48721a,a48724a,a48725a,a48726a,a48730a,a48731a,a48735a,a48736a,a48737a,a48741a,a48742a,a48745a,a48748a,a48749a,a48750a,a48754a,a48755a,a48759a,a48760a,a48761a,a48765a,a48766a,a48769a,a48772a,a48773a,a48774a,a48778a,a48779a,a48783a,a48784a,a48785a,a48789a,a48790a,a48793a,a48796a,a48797a,a48798a,a48802a,a48803a,a48807a,a48808a,a48809a,a48813a,a48814a,a48817a,a48820a,a48821a,a48822a,a48826a,a48827a,a48831a,a48832a,a48833a,a48837a,a48838a,a48841a,a48844a,a48845a,a48846a,a48850a,a48851a,a48855a,a48856a,a48857a,a48861a,a48862a,a48865a,a48868a,a48869a,a48870a,a48874a,a48875a,a48879a,a48880a,a48881a,a48885a,a48886a,a48889a,a48892a,a48893a,a48894a,a48898a,a48899a,a48903a,a48904a,a48905a,a48909a,a48910a,a48913a,a48916a,a48917a,a48918a,a48922a,a48923a,a48927a,a48928a,a48929a,a48933a,a48934a,a48937a,a48940a,a48941a,a48942a,a48946a,a48947a,a48951a,a48952a,a48953a,a48957a,a48958a,a48961a,a48964a,a48965a,a48966a,a48970a,a48971a,a48975a,a48976a,a48977a,a48981a,a48982a,a48985a,a48988a,a48989a,a48990a,a48994a,a48995a,a48999a,a49000a,a49001a,a49005a,a49006a,a49009a,a49012a,a49013a,a49014a,a49018a,a49019a,a49023a,a49024a,a49025a,a49029a,a49030a,a49033a,a49036a,a49037a,a49038a,a49042a,a49043a,a49047a,a49048a,a49049a,a49053a,a49054a,a49057a,a49060a,a49061a,a49062a,a49066a,a49067a,a49071a,a49072a,a49073a,a49077a,a49078a,a49081a,a49084a,a49085a,a49086a,a49090a,a49091a,a49095a,a49096a,a49097a,a49101a,a49102a,a49105a,a49108a,a49109a,a49110a,a49114a,a49115a,a49119a,a49120a,a49121a,a49125a,a49126a,a49129a,a49132a,a49133a,a49134a,a49138a,a49139a,a49143a,a49144a,a49145a,a49149a,a49150a,a49153a,a49156a,a49157a,a49158a,a49162a,a49163a,a49167a,a49168a,a49169a,a49173a,a49174a,a49177a,a49180a,a49181a,a49182a,a49186a,a49187a,a49191a,a49192a,a49193a,a49197a,a49198a,a49201a,a49204a,a49205a,a49206a,a49210a,a49211a,a49215a,a49216a,a49217a,a49221a,a49222a,a49225a,a49228a,a49229a,a49230a,a49234a,a49235a,a49239a,a49240a,a49241a,a49245a,a49246a,a49249a,a49252a,a49253a,a49254a,a49258a,a49259a,a49263a,a49264a,a49265a,a49269a,a49270a,a49273a,a49276a,a49277a,a49278a,a49282a,a49283a,a49287a,a49288a,a49289a,a49293a,a49294a,a49297a,a49300a,a49301a,a49302a,a49306a,a49307a,a49311a,a49312a,a49313a,a49317a,a49318a,a49321a,a49324a,a49325a,a49326a,a49330a,a49331a,a49335a,a49336a,a49337a,a49341a,a49342a,a49345a,a49348a,a49349a,a49350a,a49354a,a49355a,a49359a,a49360a,a49361a,a49365a,a49366a,a49369a,a49372a,a49373a,a49374a,a49378a,a49379a,a49383a,a49384a,a49385a,a49389a,a49390a,a49393a,a49396a,a49397a,a49398a,a49402a,a49403a,a49407a,a49408a,a49409a,a49413a,a49414a,a49417a,a49420a,a49421a,a49422a,a49426a,a49427a,a49431a,a49432a,a49433a,a49437a,a49438a,a49441a,a49444a,a49445a,a49446a,a49450a,a49451a,a49455a,a49456a,a49457a,a49461a,a49462a,a49465a,a49468a,a49469a,a49470a,a49474a,a49475a,a49479a,a49480a,a49481a,a49485a,a49486a,a49489a,a49492a,a49493a,a49494a,a49498a,a49499a,a49503a,a49504a,a49505a,a49509a,a49510a,a49513a,a49516a,a49517a,a49518a,a49522a,a49523a,a49527a,a49528a,a49529a,a49533a,a49534a,a49537a,a49540a,a49541a,a49542a,a49546a,a49547a,a49551a,a49552a,a49553a,a49557a,a49558a,a49561a,a49564a,a49565a,a49566a,a49570a,a49571a,a49575a,a49576a,a49577a,a49581a,a49582a,a49585a,a49588a,a49589a,a49590a,a49594a,a49595a,a49599a,a49600a,a49601a,a49605a,a49606a,a49609a,a49612a,a49613a,a49614a,a49618a,a49619a,a49623a,a49624a,a49625a,a49629a,a49630a,a49633a,a49636a,a49637a,a49638a,a49642a,a49643a,a49647a,a49648a,a49649a,a49653a,a49654a,a49657a,a49660a,a49661a,a49662a,a49666a,a49667a,a49671a,a49672a,a49673a,a49677a,a49678a,a49681a,a49684a,a49685a,a49686a,a49690a,a49691a,a49695a,a49696a,a49697a,a49701a,a49702a,a49705a,a49708a,a49709a,a49710a,a49714a,a49715a,a49719a,a49720a,a49721a,a49725a,a49726a,a49729a,a49732a,a49733a,a49734a,a49738a,a49739a,a49743a,a49744a,a49745a,a49749a,a49750a,a49753a,a49756a,a49757a,a49758a,a49762a,a49763a,a49767a,a49768a,a49769a,a49773a,a49774a,a49777a,a49780a,a49781a,a49782a,a49786a,a49787a,a49791a,a49792a,a49793a,a49797a,a49798a,a49801a,a49804a,a49805a,a49806a,a49810a,a49811a,a49815a,a49816a,a49817a,a49821a,a49822a,a49825a,a49828a,a49829a,a49830a,a49834a,a49835a,a49839a,a49840a,a49841a,a49845a,a49846a,a49849a,a49852a,a49853a,a49854a,a49858a,a49859a,a49863a,a49864a,a49865a,a49869a,a49870a,a49873a,a49876a,a49877a,a49878a,a49882a,a49883a,a49887a,a49888a,a49889a,a49893a,a49894a,a49897a,a49900a,a49901a,a49902a,a49906a,a49907a,a49911a,a49912a,a49913a,a49917a,a49918a,a49921a,a49924a,a49925a,a49926a,a49930a,a49931a,a49935a,a49936a,a49937a,a49941a,a49942a,a49945a,a49948a,a49949a,a49950a,a49954a,a49955a,a49959a,a49960a,a49961a,a49965a,a49966a,a49969a,a49972a,a49973a,a49974a,a49978a,a49979a,a49983a,a49984a,a49985a,a49989a,a49990a,a49993a,a49996a,a49997a,a49998a,a50002a,a50003a,a50007a,a50008a,a50009a,a50013a,a50014a,a50017a,a50020a,a50021a,a50022a,a50026a,a50027a,a50031a,a50032a,a50033a,a50037a,a50038a,a50041a,a50044a,a50045a,a50046a,a50050a,a50051a,a50055a,a50056a,a50057a,a50061a,a50062a,a50065a,a50068a,a50069a,a50070a,a50074a,a50075a,a50079a,a50080a,a50081a,a50085a,a50086a,a50089a,a50092a,a50093a,a50094a,a50098a,a50099a,a50103a,a50104a,a50105a,a50109a,a50110a,a50113a,a50116a,a50117a,a50118a,a50122a,a50123a,a50127a,a50128a,a50129a,a50133a,a50134a,a50137a,a50140a,a50141a,a50142a,a50146a,a50147a,a50151a,a50152a,a50153a,a50157a,a50158a,a50161a,a50164a,a50165a,a50166a,a50170a,a50171a,a50175a,a50176a,a50177a,a50181a,a50182a,a50185a,a50188a,a50189a,a50190a,a50194a,a50195a,a50199a,a50200a,a50201a,a50205a,a50206a,a50209a,a50212a,a50213a,a50214a,a50218a,a50219a,a50223a,a50224a,a50225a,a50229a,a50230a,a50233a,a50236a,a50237a,a50238a,a50242a,a50243a,a50247a,a50248a,a50249a,a50253a,a50254a,a50257a,a50260a,a50261a,a50262a,a50266a,a50267a,a50271a,a50272a,a50273a,a50277a,a50278a,a50281a,a50284a,a50285a,a50286a,a50290a,a50291a,a50295a,a50296a,a50297a,a50301a,a50302a,a50305a,a50308a,a50309a,a50310a,a50314a,a50315a,a50319a,a50320a,a50321a,a50325a,a50326a,a50329a,a50332a,a50333a,a50334a,a50338a,a50339a,a50343a,a50344a,a50345a,a50349a,a50350a,a50353a,a50356a,a50357a,a50358a,a50362a,a50363a,a50367a,a50368a,a50369a,a50373a,a50374a,a50377a,a50380a,a50381a,a50382a,a50386a,a50387a,a50391a,a50392a,a50393a,a50397a,a50398a,a50401a,a50404a,a50405a,a50406a,a50410a,a50411a,a50415a,a50416a,a50417a,a50421a,a50422a,a50425a,a50428a,a50429a,a50430a,a50434a,a50435a,a50439a,a50440a,a50441a,a50445a,a50446a,a50449a,a50452a,a50453a,a50454a,a50458a,a50459a,a50463a,a50464a,a50465a,a50469a,a50470a,a50473a,a50476a,a50477a,a50478a,a50482a,a50483a,a50487a,a50488a,a50489a,a50493a,a50494a,a50497a,a50500a,a50501a,a50502a,a50506a,a50507a,a50511a,a50512a,a50513a,a50517a,a50518a,a50521a,a50524a,a50525a,a50526a,a50530a,a50531a,a50535a,a50536a,a50537a,a50541a,a50542a,a50545a,a50548a,a50549a,a50550a,a50554a,a50555a,a50559a,a50560a,a50561a,a50565a,a50566a,a50569a,a50572a,a50573a,a50574a,a50578a,a50579a,a50583a,a50584a,a50585a,a50589a,a50590a,a50593a,a50596a,a50597a,a50598a,a50602a,a50603a,a50607a,a50608a,a50609a,a50613a,a50614a,a50617a,a50620a,a50621a,a50622a,a50626a,a50627a,a50631a,a50632a,a50633a,a50637a,a50638a,a50641a,a50644a,a50645a,a50646a,a50650a,a50651a,a50655a,a50656a,a50657a,a50661a,a50662a,a50665a,a50668a,a50669a,a50670a,a50674a,a50675a,a50679a,a50680a,a50681a,a50685a,a50686a,a50689a,a50692a,a50693a,a50694a,a50698a,a50699a,a50703a,a50704a,a50705a,a50709a,a50710a,a50713a,a50716a,a50717a,a50718a,a50722a,a50723a,a50727a,a50728a,a50729a,a50733a,a50734a,a50737a,a50740a,a50741a,a50742a,a50746a,a50747a,a50751a,a50752a,a50753a,a50757a,a50758a,a50761a,a50764a,a50765a,a50766a,a50770a,a50771a,a50775a,a50776a,a50777a,a50781a,a50782a,a50785a,a50788a,a50789a,a50790a,a50794a,a50795a,a50799a,a50800a,a50801a,a50805a,a50806a,a50809a,a50812a,a50813a,a50814a,a50818a,a50819a,a50823a,a50824a,a50825a,a50829a,a50830a,a50833a,a50836a,a50837a,a50838a,a50842a,a50843a,a50847a,a50848a,a50849a,a50853a,a50854a,a50857a,a50860a,a50861a,a50862a,a50866a,a50867a,a50871a,a50872a,a50873a,a50877a,a50878a,a50881a,a50884a,a50885a,a50886a,a50890a,a50891a,a50895a,a50896a,a50897a,a50901a,a50902a,a50905a,a50908a,a50909a,a50910a,a50914a,a50915a,a50919a,a50920a,a50921a,a50925a,a50926a,a50929a,a50932a,a50933a,a50934a,a50938a,a50939a,a50943a,a50944a,a50945a,a50949a,a50950a,a50953a,a50956a,a50957a,a50958a,a50962a,a50963a,a50967a,a50968a,a50969a,a50973a,a50974a,a50977a,a50980a,a50981a,a50982a,a50986a,a50987a,a50991a,a50992a,a50993a,a50997a,a50998a,a51001a,a51004a,a51005a,a51006a,a51010a,a51011a,a51015a,a51016a,a51017a,a51021a,a51022a,a51025a,a51028a,a51029a,a51030a,a51034a,a51035a,a51039a,a51040a,a51041a,a51045a,a51046a,a51049a,a51052a,a51053a,a51054a,a51058a,a51059a,a51063a,a51064a,a51065a,a51069a,a51070a,a51073a,a51076a,a51077a,a51078a,a51082a,a51083a,a51087a,a51088a,a51089a,a51093a,a51094a,a51097a,a51100a,a51101a,a51102a,a51106a,a51107a,a51111a,a51112a,a51113a,a51117a,a51118a,a51121a,a51124a,a51125a,a51126a,a51130a,a51131a,a51135a,a51136a,a51137a,a51141a,a51142a,a51145a,a51148a,a51149a,a51150a,a51154a,a51155a,a51159a,a51160a,a51161a,a51165a,a51166a,a51169a,a51172a,a51173a,a51174a,a51178a,a51179a,a51183a,a51184a,a51185a,a51189a,a51190a,a51193a,a51196a,a51197a,a51198a,a51202a,a51203a,a51207a,a51208a,a51209a,a51213a,a51214a,a51217a,a51220a,a51221a,a51222a,a51226a,a51227a,a51231a,a51232a,a51233a,a51237a,a51238a,a51241a,a51244a,a51245a,a51246a,a51250a,a51251a,a51255a,a51256a,a51257a,a51261a,a51262a,a51265a,a51268a,a51269a,a51270a,a51274a,a51275a,a51279a,a51280a,a51281a,a51285a,a51286a,a51289a,a51292a,a51293a,a51294a,a51298a,a51299a,a51303a,a51304a,a51305a,a51309a,a51310a,a51313a,a51316a,a51317a,a51318a,a51322a,a51323a,a51327a,a51328a,a51329a,a51333a,a51334a,a51337a,a51340a,a51341a,a51342a,a51346a,a51347a,a51351a,a51352a,a51353a,a51357a,a51358a,a51361a,a51364a,a51365a,a51366a,a51370a,a51371a,a51375a,a51376a,a51377a,a51381a,a51382a,a51385a,a51388a,a51389a,a51390a,a51394a,a51395a,a51399a,a51400a,a51401a,a51405a,a51406a,a51409a,a51412a,a51413a,a51414a,a51418a,a51419a,a51423a,a51424a,a51425a,a51429a,a51430a,a51433a,a51436a,a51437a,a51438a,a51442a,a51443a,a51447a,a51448a,a51449a,a51453a,a51454a,a51457a,a51460a,a51461a,a51462a,a51466a,a51467a,a51471a,a51472a,a51473a,a51477a,a51478a,a51481a,a51484a,a51485a,a51486a,a51490a,a51491a,a51495a,a51496a,a51497a,a51501a,a51502a,a51505a,a51508a,a51509a,a51510a,a51514a,a51515a,a51519a,a51520a,a51521a,a51525a,a51526a,a51529a,a51532a,a51533a,a51534a,a51538a,a51539a,a51543a,a51544a,a51545a,a51549a,a51550a,a51553a,a51556a,a51557a,a51558a,a51562a,a51563a,a51567a,a51568a,a51569a,a51573a,a51574a,a51577a,a51580a,a51581a,a51582a,a51586a,a51587a,a51591a,a51592a,a51593a,a51597a,a51598a,a51601a,a51604a,a51605a,a51606a,a51610a,a51611a,a51615a,a51616a,a51617a,a51621a,a51622a,a51625a,a51628a,a51629a,a51630a,a51634a,a51635a,a51639a,a51640a,a51641a,a51645a,a51646a,a51649a,a51652a,a51653a,a51654a,a51658a,a51659a,a51663a,a51664a,a51665a,a51669a,a51670a,a51673a,a51676a,a51677a,a51678a,a51682a,a51683a,a51687a,a51688a,a51689a,a51693a,a51694a,a51697a,a51700a,a51701a,a51702a,a51706a,a51707a,a51711a,a51712a,a51713a,a51717a,a51718a,a51721a,a51724a,a51725a,a51726a,a51730a,a51731a,a51735a,a51736a,a51737a,a51741a,a51742a,a51745a,a51748a,a51749a,a51750a,a51754a,a51755a,a51759a,a51760a,a51761a,a51765a,a51766a,a51769a,a51772a,a51773a,a51774a,a51778a,a51779a,a51783a,a51784a,a51785a,a51789a,a51790a,a51793a,a51796a,a51797a,a51798a,a51802a,a51803a,a51807a,a51808a,a51809a,a51813a,a51814a,a51817a,a51820a,a51821a,a51822a,a51826a,a51827a,a51831a,a51832a,a51833a,a51837a,a51838a,a51841a,a51844a,a51845a,a51846a,a51850a,a51851a,a51855a,a51856a,a51857a,a51861a,a51862a,a51865a,a51868a,a51869a,a51870a,a51874a,a51875a,a51879a,a51880a,a51881a,a51885a,a51886a,a51889a,a51892a,a51893a,a51894a,a51898a,a51899a,a51903a,a51904a,a51905a,a51909a,a51910a,a51913a,a51916a,a51917a,a51918a,a51922a,a51923a,a51927a,a51928a,a51929a,a51933a,a51934a,a51937a,a51940a,a51941a,a51942a,a51946a,a51947a,a51951a,a51952a,a51953a,a51957a,a51958a,a51961a,a51964a,a51965a,a51966a,a51970a,a51971a,a51975a,a51976a,a51977a,a51981a,a51982a,a51985a,a51988a,a51989a,a51990a,a51994a,a51995a,a51999a,a52000a,a52001a,a52005a,a52006a,a52009a,a52012a,a52013a,a52014a,a52018a,a52019a,a52023a,a52024a,a52025a,a52029a,a52030a,a52033a,a52036a,a52037a,a52038a,a52042a,a52043a,a52047a,a52048a,a52049a,a52053a,a52054a,a52057a,a52060a,a52061a,a52062a,a52066a,a52067a,a52071a,a52072a,a52073a,a52077a,a52078a,a52081a,a52084a,a52085a,a52086a,a52090a,a52091a,a52095a,a52096a,a52097a,a52101a,a52102a,a52105a,a52108a,a52109a,a52110a,a52114a,a52115a,a52119a,a52120a,a52121a,a52125a,a52126a,a52129a,a52132a,a52133a,a52134a,a52138a,a52139a,a52143a,a52144a,a52145a,a52149a,a52150a,a52153a,a52156a,a52157a,a52158a,a52162a,a52163a,a52167a,a52168a,a52169a,a52173a,a52174a,a52177a,a52180a,a52181a,a52182a,a52186a,a52187a,a52191a,a52192a,a52193a,a52197a,a52198a,a52201a,a52204a,a52205a,a52206a,a52210a,a52211a,a52215a,a52216a,a52217a,a52221a,a52222a,a52225a,a52228a,a52229a,a52230a,a52234a,a52235a,a52239a,a52240a,a52241a,a52245a,a52246a,a52249a,a52252a,a52253a,a52254a,a52258a,a52259a,a52263a,a52264a,a52265a,a52269a,a52270a,a52273a,a52276a,a52277a,a52278a,a52282a,a52283a,a52287a,a52288a,a52289a,a52293a,a52294a,a52297a,a52300a,a52301a,a52302a,a52306a,a52307a,a52311a,a52312a,a52313a,a52317a,a52318a,a52321a,a52324a,a52325a,a52326a,a52330a,a52331a,a52335a,a52336a,a52337a,a52341a,a52342a,a52345a,a52348a,a52349a,a52350a,a52354a,a52355a,a52359a,a52360a,a52361a,a52365a,a52366a,a52369a,a52372a,a52373a,a52374a,a52378a,a52379a,a52383a,a52384a,a52385a,a52389a,a52390a,a52393a,a52396a,a52397a,a52398a,a52402a,a52403a,a52407a,a52408a,a52409a,a52413a,a52414a,a52417a,a52420a,a52421a,a52422a,a52426a,a52427a,a52431a,a52432a,a52433a,a52437a,a52438a,a52441a,a52444a,a52445a,a52446a,a52450a,a52451a,a52455a,a52456a,a52457a,a52461a,a52462a,a52465a,a52468a,a52469a,a52470a,a52474a,a52475a,a52479a,a52480a,a52481a,a52485a,a52486a,a52489a,a52492a,a52493a,a52494a,a52498a,a52499a,a52503a,a52504a,a52505a,a52509a,a52510a,a52513a,a52516a,a52517a,a52518a,a52522a,a52523a,a52527a,a52528a,a52529a,a52533a,a52534a,a52537a,a52540a,a52541a,a52542a,a52546a,a52547a,a52551a,a52552a,a52553a,a52557a,a52558a,a52561a,a52564a,a52565a,a52566a,a52570a,a52571a,a52575a,a52576a,a52577a,a52581a,a52582a,a52585a,a52588a,a52589a,a52590a,a52594a,a52595a,a52599a,a52600a,a52601a,a52605a,a52606a,a52609a,a52612a,a52613a,a52614a,a52618a,a52619a,a52623a,a52624a,a52625a,a52629a,a52630a,a52633a,a52636a,a52637a,a52638a,a52642a,a52643a,a52647a,a52648a,a52649a,a52653a,a52654a,a52657a,a52660a,a52661a,a52662a,a52666a,a52667a,a52671a,a52672a,a52673a,a52677a,a52678a,a52681a,a52684a,a52685a,a52686a,a52690a,a52691a,a52695a,a52696a,a52697a,a52701a,a52702a,a52705a,a52708a,a52709a,a52710a,a52714a,a52715a,a52719a,a52720a,a52721a,a52725a,a52726a,a52729a,a52732a,a52733a,a52734a,a52738a,a52739a,a52743a,a52744a,a52745a,a52749a,a52750a,a52753a,a52756a,a52757a,a52758a,a52762a,a52763a,a52767a,a52768a,a52769a,a52773a,a52774a,a52777a,a52780a,a52781a,a52782a,a52786a,a52787a,a52791a,a52792a,a52793a,a52797a,a52798a,a52801a,a52804a,a52805a,a52806a,a52810a,a52811a,a52815a,a52816a,a52817a,a52821a,a52822a,a52825a,a52828a,a52829a,a52830a,a52834a,a52835a,a52839a,a52840a,a52841a,a52845a,a52846a,a52849a,a52852a,a52853a,a52854a,a52858a,a52859a,a52863a,a52864a,a52865a,a52869a,a52870a,a52873a,a52876a,a52877a,a52878a,a52882a,a52883a,a52887a,a52888a,a52889a,a52893a,a52894a,a52897a,a52900a,a52901a,a52902a,a52906a,a52907a,a52911a,a52912a,a52913a,a52917a,a52918a,a52921a,a52924a,a52925a,a52926a,a52930a,a52931a,a52935a,a52936a,a52937a,a52941a,a52942a,a52945a,a52948a,a52949a,a52950a,a52954a,a52955a,a52959a,a52960a,a52961a,a52965a,a52966a,a52969a,a52972a,a52973a,a52974a,a52978a,a52979a,a52983a,a52984a,a52985a,a52989a,a52990a,a52993a,a52996a,a52997a,a52998a,a53002a,a53003a,a53007a,a53008a,a53009a,a53013a,a53014a,a53017a,a53020a,a53021a,a53022a,a53026a,a53027a,a53031a,a53032a,a53033a,a53037a,a53038a,a53041a,a53044a,a53045a,a53046a,a53050a,a53051a,a53055a,a53056a,a53057a,a53061a,a53062a,a53065a,a53068a,a53069a,a53070a,a53074a,a53075a,a53079a,a53080a,a53081a,a53085a,a53086a,a53089a,a53092a,a53093a,a53094a,a53098a,a53099a,a53103a,a53104a,a53105a,a53109a,a53110a,a53113a,a53116a,a53117a,a53118a,a53122a,a53123a,a53127a,a53128a,a53129a,a53133a,a53134a,a53137a,a53140a,a53141a,a53142a,a53146a,a53147a,a53151a,a53152a,a53153a,a53157a,a53158a,a53161a,a53164a,a53165a,a53166a,a53170a,a53171a,a53175a,a53176a,a53177a,a53181a,a53182a,a53185a,a53188a,a53189a,a53190a,a53194a,a53195a,a53199a,a53200a,a53201a,a53205a,a53206a,a53209a,a53212a,a53213a,a53214a,a53218a,a53219a,a53223a,a53224a,a53225a,a53229a,a53230a,a53233a,a53236a,a53237a,a53238a,a53242a,a53243a,a53247a,a53248a,a53249a,a53253a,a53254a,a53257a,a53260a,a53261a,a53262a,a53266a,a53267a,a53271a,a53272a,a53273a,a53277a,a53278a,a53281a,a53284a,a53285a,a53286a,a53290a,a53291a,a53295a,a53296a,a53297a,a53301a,a53302a,a53305a,a53308a,a53309a,a53310a,a53314a,a53315a,a53319a,a53320a,a53321a,a53325a,a53326a,a53329a,a53332a,a53333a,a53334a,a53338a,a53339a,a53343a,a53344a,a53345a,a53349a,a53350a,a53353a,a53356a,a53357a,a53358a,a53362a,a53363a,a53367a,a53368a,a53369a,a53373a,a53374a,a53377a,a53380a,a53381a,a53382a,a53386a,a53387a,a53391a,a53392a,a53393a,a53397a,a53398a,a53401a,a53404a,a53405a,a53406a,a53410a,a53411a,a53415a,a53416a,a53417a,a53421a,a53422a,a53425a,a53428a,a53429a,a53430a,a53434a,a53435a,a53439a,a53440a,a53441a,a53445a,a53446a,a53449a,a53452a,a53453a,a53454a,a53458a,a53459a,a53463a,a53464a,a53465a,a53469a,a53470a,a53473a,a53476a,a53477a,a53478a,a53482a,a53483a,a53487a,a53488a,a53489a,a53493a,a53494a,a53497a,a53500a,a53501a,a53502a,a53506a,a53507a,a53511a,a53512a,a53513a,a53517a,a53518a,a53521a,a53524a,a53525a,a53526a,a53530a,a53531a,a53535a,a53536a,a53537a,a53541a,a53542a,a53545a,a53548a,a53549a,a53550a,a53554a,a53555a,a53559a,a53560a,a53561a,a53565a,a53566a,a53569a,a53572a,a53573a,a53574a,a53578a,a53579a,a53583a,a53584a,a53585a,a53589a,a53590a,a53593a,a53596a,a53597a,a53598a,a53602a,a53603a,a53607a,a53608a,a53609a,a53613a,a53614a,a53617a,a53620a,a53621a,a53622a,a53626a,a53627a,a53631a,a53632a,a53633a,a53637a,a53638a,a53641a,a53644a,a53645a,a53646a,a53650a,a53651a,a53655a,a53656a,a53657a,a53661a,a53662a,a53665a,a53668a,a53669a,a53670a,a53674a,a53675a,a53679a,a53680a,a53681a,a53685a,a53686a,a53689a,a53692a,a53693a,a53694a,a53698a,a53699a,a53703a,a53704a,a53705a,a53709a,a53710a,a53713a,a53716a,a53717a,a53718a,a53722a,a53723a,a53727a,a53728a,a53729a,a53733a,a53734a,a53737a,a53740a,a53741a,a53742a,a53746a,a53747a,a53751a,a53752a,a53753a,a53757a,a53758a,a53761a,a53764a,a53765a,a53766a,a53770a,a53771a,a53775a,a53776a,a53777a,a53781a,a53782a,a53785a,a53788a,a53789a,a53790a,a53794a,a53795a,a53799a,a53800a,a53801a,a53805a,a53806a,a53809a,a53812a,a53813a,a53814a,a53818a,a53819a,a53823a,a53824a,a53825a,a53829a,a53830a,a53833a,a53836a,a53837a,a53838a,a53842a,a53843a,a53847a,a53848a,a53849a,a53853a,a53854a,a53857a,a53860a,a53861a,a53862a,a53866a,a53867a,a53871a,a53872a,a53873a,a53877a,a53878a,a53881a,a53884a,a53885a,a53886a,a53890a,a53891a,a53895a,a53896a,a53897a,a53901a,a53902a,a53905a,a53908a,a53909a,a53910a,a53914a,a53915a,a53919a,a53920a,a53921a,a53925a,a53926a,a53929a,a53932a,a53933a,a53934a,a53938a,a53939a,a53943a,a53944a,a53945a,a53949a,a53950a,a53953a,a53956a,a53957a,a53958a,a53962a,a53963a,a53967a,a53968a,a53969a,a53973a,a53974a,a53977a,a53980a,a53981a,a53982a,a53986a,a53987a,a53991a,a53992a,a53993a,a53997a,a53998a,a54001a,a54004a,a54005a,a54006a,a54010a,a54011a,a54015a,a54016a,a54017a,a54021a,a54022a,a54025a,a54028a,a54029a,a54030a,a54034a,a54035a,a54039a,a54040a,a54041a,a54045a,a54046a,a54049a,a54052a,a54053a,a54054a,a54058a,a54059a,a54063a,a54064a,a54065a,a54069a,a54070a,a54073a,a54076a,a54077a,a54078a,a54082a,a54083a,a54087a,a54088a,a54089a,a54093a,a54094a,a54097a,a54100a,a54101a,a54102a,a54106a,a54107a,a54111a,a54112a,a54113a,a54117a,a54118a,a54121a,a54124a,a54125a,a54126a,a54130a,a54131a,a54135a,a54136a,a54137a,a54141a,a54142a,a54145a,a54148a,a54149a,a54150a,a54154a,a54155a,a54159a,a54160a,a54161a,a54165a,a54166a,a54169a,a54172a,a54173a,a54174a,a54178a,a54179a,a54183a,a54184a,a54185a,a54189a,a54190a,a54193a,a54196a,a54197a,a54198a,a54202a,a54203a,a54207a,a54208a,a54209a,a54213a,a54214a,a54217a,a54220a,a54221a,a54222a,a54226a,a54227a,a54231a,a54232a,a54233a,a54237a,a54238a,a54241a,a54244a,a54245a,a54246a,a54250a,a54251a,a54255a,a54256a,a54257a,a54261a,a54262a,a54265a,a54268a,a54269a,a54270a,a54274a,a54275a,a54279a,a54280a,a54281a,a54285a,a54286a,a54289a,a54292a,a54293a,a54294a,a54298a,a54299a,a54303a,a54304a,a54305a,a54309a,a54310a,a54313a,a54316a,a54317a,a54318a,a54322a,a54323a,a54327a,a54328a,a54329a,a54333a,a54334a,a54337a,a54340a,a54341a,a54342a,a54346a,a54347a,a54351a,a54352a,a54353a,a54357a,a54358a,a54361a,a54364a,a54365a,a54366a,a54370a,a54371a,a54375a,a54376a,a54377a,a54381a,a54382a,a54385a,a54388a,a54389a,a54390a,a54394a,a54395a,a54399a,a54400a,a54401a,a54405a,a54406a,a54409a,a54412a,a54413a,a54414a,a54418a,a54419a,a54423a,a54424a,a54425a,a54429a,a54430a,a54433a,a54436a,a54437a,a54438a,a54442a,a54443a,a54447a,a54448a,a54449a,a54453a,a54454a,a54457a,a54460a,a54461a,a54462a,a54466a,a54467a,a54471a,a54472a,a54473a,a54477a,a54478a,a54481a,a54484a,a54485a,a54486a,a54490a,a54491a,a54495a,a54496a,a54497a,a54501a,a54502a,a54505a,a54508a,a54509a,a54510a,a54514a,a54515a,a54519a,a54520a,a54521a,a54525a,a54526a,a54529a,a54532a,a54533a,a54534a,a54538a,a54539a,a54543a,a54544a,a54545a,a54549a,a54550a,a54553a,a54556a,a54557a,a54558a,a54562a,a54563a,a54567a,a54568a,a54569a,a54573a,a54574a,a54577a,a54580a,a54581a,a54582a,a54586a,a54587a,a54591a,a54592a,a54593a,a54597a,a54598a,a54601a,a54604a,a54605a,a54606a,a54610a,a54611a,a54615a,a54616a,a54617a,a54621a,a54622a,a54625a,a54628a,a54629a,a54630a,a54634a,a54635a,a54639a,a54640a,a54641a,a54645a,a54646a,a54649a,a54652a,a54653a,a54654a,a54658a,a54659a,a54663a,a54664a,a54665a,a54669a,a54670a,a54673a,a54676a,a54677a,a54678a,a54682a,a54683a,a54687a,a54688a,a54689a,a54693a,a54694a,a54697a,a54700a,a54701a,a54702a,a54706a,a54707a,a54711a,a54712a,a54713a,a54717a,a54718a,a54721a,a54724a,a54725a,a54726a,a54730a,a54731a,a54735a,a54736a,a54737a,a54741a,a54742a,a54745a,a54748a,a54749a,a54750a,a54754a,a54755a,a54759a,a54760a,a54761a,a54765a,a54766a,a54769a,a54772a,a54773a,a54774a,a54778a,a54779a,a54783a,a54784a,a54785a,a54789a,a54790a,a54793a,a54796a,a54797a,a54798a,a54802a,a54803a,a54807a,a54808a,a54809a,a54813a,a54814a,a54817a,a54820a,a54821a,a54822a,a54826a,a54827a,a54831a,a54832a,a54833a,a54837a,a54838a,a54841a,a54844a,a54845a,a54846a,a54850a,a54851a,a54855a,a54856a,a54857a,a54861a,a54862a,a54865a,a54868a,a54869a,a54870a,a54874a,a54875a,a54879a,a54880a,a54881a,a54885a,a54886a,a54889a,a54892a,a54893a,a54894a,a54898a,a54899a,a54903a,a54904a,a54905a,a54909a,a54910a,a54913a,a54916a,a54917a,a54918a,a54922a,a54923a,a54927a,a54928a,a54929a,a54933a,a54934a,a54937a,a54940a,a54941a,a54942a,a54946a,a54947a,a54951a,a54952a,a54953a,a54957a,a54958a,a54961a,a54964a,a54965a,a54966a,a54970a,a54971a,a54975a,a54976a,a54977a,a54981a,a54982a,a54985a,a54988a,a54989a,a54990a,a54994a,a54995a,a54999a,a55000a,a55001a,a55005a,a55006a,a55009a,a55012a,a55013a,a55014a,a55018a,a55019a,a55023a,a55024a,a55025a,a55029a,a55030a,a55033a,a55036a,a55037a,a55038a,a55042a,a55043a,a55047a,a55048a,a55049a,a55053a,a55054a,a55057a,a55060a,a55061a,a55062a,a55066a,a55067a,a55071a,a55072a,a55073a,a55077a,a55078a,a55081a,a55084a,a55085a,a55086a,a55090a,a55091a,a55095a,a55096a,a55097a,a55101a,a55102a,a55105a,a55108a,a55109a,a55110a,a55114a,a55115a,a55119a,a55120a,a55121a,a55125a,a55126a,a55129a,a55132a,a55133a,a55134a,a55138a,a55139a,a55143a,a55144a,a55145a,a55149a,a55150a,a55153a,a55156a,a55157a,a55158a,a55162a,a55163a,a55167a,a55168a,a55169a,a55173a,a55174a,a55177a,a55180a,a55181a,a55182a,a55186a,a55187a,a55191a,a55192a,a55193a,a55197a,a55198a,a55201a,a55204a,a55205a,a55206a,a55210a,a55211a,a55215a,a55216a,a55217a,a55221a,a55222a,a55225a,a55228a,a55229a,a55230a,a55234a,a55235a,a55239a,a55240a,a55241a,a55245a,a55246a,a55249a,a55252a,a55253a,a55254a,a55258a,a55259a,a55263a,a55264a,a55265a,a55269a,a55270a,a55273a,a55276a,a55277a,a55278a,a55282a,a55283a,a55287a,a55288a,a55289a,a55293a,a55294a,a55297a,a55300a,a55301a,a55302a,a55306a,a55307a,a55311a,a55312a,a55313a,a55317a,a55318a,a55321a,a55324a,a55325a,a55326a,a55330a,a55331a,a55335a,a55336a,a55337a,a55341a,a55342a,a55345a,a55348a,a55349a,a55350a,a55354a,a55355a,a55359a,a55360a,a55361a,a55365a,a55366a,a55369a,a55372a,a55373a,a55374a,a55378a,a55379a,a55383a,a55384a,a55385a,a55389a,a55390a,a55393a,a55396a,a55397a,a55398a,a55402a,a55403a,a55407a,a55408a,a55409a,a55413a,a55414a,a55417a,a55420a,a55421a,a55422a,a55426a,a55427a,a55431a,a55432a,a55433a,a55437a,a55438a,a55441a,a55444a,a55445a,a55446a,a55450a,a55451a,a55455a,a55456a,a55457a,a55461a,a55462a,a55465a,a55468a,a55469a,a55470a,a55474a,a55475a,a55479a,a55480a,a55481a,a55485a,a55486a,a55489a,a55492a,a55493a,a55494a,a55498a,a55499a,a55503a,a55504a,a55505a,a55509a,a55510a,a55513a,a55516a,a55517a,a55518a,a55522a,a55523a,a55527a,a55528a,a55529a,a55533a,a55534a,a55537a,a55540a,a55541a,a55542a,a55546a,a55547a,a55551a,a55552a,a55553a,a55557a,a55558a,a55561a,a55564a,a55565a,a55566a,a55570a,a55571a,a55575a,a55576a,a55577a,a55581a,a55582a,a55585a,a55588a,a55589a,a55590a,a55594a,a55595a,a55599a,a55600a,a55601a,a55605a,a55606a,a55609a,a55612a,a55613a,a55614a,a55618a,a55619a,a55623a,a55624a,a55625a,a55629a,a55630a,a55633a,a55636a,a55637a,a55638a,a55642a,a55643a,a55647a,a55648a,a55649a,a55653a,a55654a,a55657a,a55660a,a55661a,a55662a,a55666a,a55667a,a55671a,a55672a,a55673a,a55677a,a55678a,a55681a,a55684a,a55685a,a55686a,a55690a,a55691a,a55695a,a55696a,a55697a,a55701a,a55702a,a55705a,a55708a,a55709a,a55710a,a55714a,a55715a,a55719a,a55720a,a55721a,a55725a,a55726a,a55729a,a55732a,a55733a,a55734a,a55738a,a55739a,a55743a,a55744a,a55745a,a55749a,a55750a,a55753a,a55756a,a55757a,a55758a,a55762a,a55763a,a55767a,a55768a,a55769a,a55773a,a55774a,a55777a,a55780a,a55781a,a55782a,a55786a,a55787a,a55791a,a55792a,a55793a,a55797a,a55798a,a55801a,a55804a,a55805a,a55806a,a55810a,a55811a,a55815a,a55816a,a55817a,a55821a,a55822a,a55825a,a55828a,a55829a,a55830a,a55834a,a55835a,a55839a,a55840a,a55841a,a55845a,a55846a,a55849a,a55852a,a55853a,a55854a,a55858a,a55859a,a55863a,a55864a,a55865a,a55869a,a55870a,a55873a,a55876a,a55877a,a55878a,a55882a,a55883a,a55887a,a55888a,a55889a,a55893a,a55894a,a55897a,a55900a,a55901a,a55902a,a55906a,a55907a,a55911a,a55912a,a55913a,a55917a,a55918a,a55921a,a55924a,a55925a,a55926a,a55930a,a55931a,a55935a,a55936a,a55937a,a55941a,a55942a,a55945a,a55948a,a55949a,a55950a,a55954a,a55955a,a55959a,a55960a,a55961a,a55965a,a55966a,a55969a,a55972a,a55973a,a55974a,a55978a,a55979a,a55983a,a55984a,a55985a,a55989a,a55990a,a55993a,a55996a,a55997a,a55998a,a56002a,a56003a,a56007a,a56008a,a56009a,a56013a,a56014a,a56017a,a56020a,a56021a,a56022a,a56026a,a56027a,a56031a,a56032a,a56033a,a56037a,a56038a,a56041a,a56044a,a56045a,a56046a,a56050a,a56051a,a56055a,a56056a,a56057a,a56061a,a56062a,a56065a,a56068a,a56069a,a56070a,a56074a,a56075a,a56079a,a56080a,a56081a,a56085a,a56086a,a56089a,a56092a,a56093a,a56094a,a56098a,a56099a,a56103a,a56104a,a56105a,a56109a,a56110a,a56113a,a56116a,a56117a,a56118a,a56122a,a56123a,a56127a,a56128a,a56129a,a56133a,a56134a,a56137a,a56140a,a56141a,a56142a,a56146a,a56147a,a56151a,a56152a,a56153a,a56157a,a56158a,a56161a,a56164a,a56165a,a56166a,a56170a,a56171a,a56175a,a56176a,a56177a,a56181a,a56182a,a56185a,a56188a,a56189a,a56190a,a56194a,a56195a,a56199a,a56200a,a56201a,a56205a,a56206a,a56209a,a56212a,a56213a,a56214a,a56218a,a56219a,a56223a,a56224a,a56225a,a56229a,a56230a,a56233a,a56236a,a56237a,a56238a,a56242a,a56243a,a56247a,a56248a,a56249a,a56253a,a56254a,a56257a,a56260a,a56261a,a56262a,a56266a,a56267a,a56271a,a56272a,a56273a,a56277a,a56278a,a56281a,a56284a,a56285a,a56286a,a56290a,a56291a,a56295a,a56296a,a56297a,a56301a,a56302a,a56305a,a56308a,a56309a,a56310a,a56314a,a56315a,a56319a,a56320a,a56321a,a56325a,a56326a,a56329a,a56332a,a56333a,a56334a,a56338a,a56339a,a56343a,a56344a,a56345a,a56349a,a56350a,a56353a,a56356a,a56357a,a56358a,a56362a,a56363a,a56367a,a56368a,a56369a,a56373a,a56374a,a56377a,a56380a,a56381a,a56382a,a56386a,a56387a,a56391a,a56392a,a56393a,a56397a,a56398a,a56401a,a56404a,a56405a,a56406a,a56410a,a56411a,a56415a,a56416a,a56417a,a56421a,a56422a,a56425a,a56428a,a56429a,a56430a,a56434a,a56435a,a56439a,a56440a,a56441a,a56445a,a56446a,a56449a,a56452a,a56453a,a56454a,a56458a,a56459a,a56463a,a56464a,a56465a,a56469a,a56470a,a56473a,a56476a,a56477a,a56478a,a56482a,a56483a,a56487a,a56488a,a56489a,a56493a,a56494a,a56497a,a56500a,a56501a,a56502a,a56506a,a56507a,a56511a,a56512a,a56513a,a56517a,a56518a,a56521a,a56524a,a56525a,a56526a,a56530a,a56531a,a56535a,a56536a,a56537a,a56541a,a56542a,a56545a,a56548a,a56549a,a56550a,a56554a,a56555a,a56559a,a56560a,a56561a,a56565a,a56566a,a56569a,a56572a,a56573a,a56574a,a56578a,a56579a,a56583a,a56584a,a56585a,a56589a,a56590a,a56593a,a56596a,a56597a,a56598a,a56602a,a56603a,a56607a,a56608a,a56609a,a56613a,a56614a,a56617a,a56620a,a56621a,a56622a,a56626a,a56627a,a56631a,a56632a,a56633a,a56637a,a56638a,a56641a,a56644a,a56645a,a56646a,a56650a,a56651a,a56655a,a56656a,a56657a,a56661a,a56662a,a56665a,a56668a,a56669a,a56670a,a56674a,a56675a,a56679a,a56680a,a56681a,a56685a,a56686a,a56689a,a56692a,a56693a,a56694a,a56698a,a56699a,a56703a,a56704a,a56705a,a56709a,a56710a,a56713a,a56716a,a56717a,a56718a,a56722a,a56723a,a56727a,a56728a,a56729a,a56733a,a56734a,a56737a,a56740a,a56741a,a56742a,a56746a,a56747a,a56751a,a56752a,a56753a,a56757a,a56758a,a56761a,a56764a,a56765a,a56766a,a56770a,a56771a,a56775a,a56776a,a56777a,a56781a,a56782a,a56785a,a56788a,a56789a,a56790a,a56794a,a56795a,a56799a,a56800a,a56801a,a56805a,a56806a,a56809a,a56812a,a56813a,a56814a,a56818a,a56819a,a56823a,a56824a,a56825a,a56829a,a56830a,a56833a,a56836a,a56837a,a56838a,a56842a,a56843a,a56847a,a56848a,a56849a,a56853a,a56854a,a56857a,a56860a,a56861a,a56862a,a56866a,a56867a,a56871a,a56872a,a56873a,a56877a,a56878a,a56881a,a56884a,a56885a,a56886a,a56890a,a56891a,a56895a,a56896a,a56897a,a56901a,a56902a,a56905a,a56908a,a56909a,a56910a,a56914a,a56915a,a56919a,a56920a,a56921a,a56925a,a56926a,a56929a,a56932a,a56933a,a56934a,a56938a,a56939a,a56943a,a56944a,a56945a,a56949a,a56950a,a56953a,a56956a,a56957a,a56958a,a56962a,a56963a,a56967a,a56968a,a56969a,a56973a,a56974a,a56977a,a56980a,a56981a,a56982a,a56986a,a56987a,a56991a,a56992a,a56993a,a56997a,a56998a,a57001a,a57004a,a57005a,a57006a,a57010a,a57011a,a57015a,a57016a,a57017a,a57021a,a57022a,a57025a,a57028a,a57029a,a57030a,a57034a,a57035a,a57039a,a57040a,a57041a,a57045a,a57046a,a57049a,a57052a,a57053a,a57054a,a57058a,a57059a,a57063a,a57064a,a57065a,a57069a,a57070a,a57073a,a57076a,a57077a,a57078a,a57082a,a57083a,a57087a,a57088a,a57089a,a57093a,a57094a,a57097a,a57100a,a57101a,a57102a,a57106a,a57107a,a57111a,a57112a,a57113a,a57117a,a57118a,a57121a,a57124a,a57125a,a57126a,a57130a,a57131a,a57135a,a57136a,a57137a,a57141a,a57142a,a57145a,a57148a,a57149a,a57150a,a57154a,a57155a,a57159a,a57160a,a57161a,a57165a,a57166a,a57169a,a57172a,a57173a,a57174a,a57178a,a57179a,a57183a,a57184a,a57185a,a57189a,a57190a,a57193a,a57196a,a57197a,a57198a,a57202a,a57203a,a57207a,a57208a,a57209a,a57213a,a57214a,a57217a,a57220a,a57221a,a57222a,a57226a,a57227a,a57231a,a57232a,a57233a,a57237a,a57238a,a57241a,a57244a,a57245a,a57246a,a57250a,a57251a,a57255a,a57256a,a57257a,a57261a,a57262a,a57265a,a57268a,a57269a,a57270a,a57274a,a57275a,a57279a,a57280a,a57281a,a57285a,a57286a,a57289a,a57292a,a57293a,a57294a,a57298a,a57299a,a57303a,a57304a,a57305a,a57309a,a57310a,a57313a,a57316a,a57317a,a57318a,a57322a,a57323a,a57327a,a57328a,a57329a,a57333a,a57334a,a57337a,a57340a,a57341a,a57342a,a57346a,a57347a,a57351a,a57352a,a57353a,a57357a,a57358a,a57361a,a57364a,a57365a,a57366a,a57370a,a57371a,a57375a,a57376a,a57377a,a57381a,a57382a,a57385a,a57388a,a57389a,a57390a,a57394a,a57395a,a57399a,a57400a,a57401a,a57405a,a57406a,a57409a,a57412a,a57413a,a57414a,a57418a,a57419a,a57423a,a57424a,a57425a,a57429a,a57430a,a57433a,a57436a,a57437a,a57438a,a57442a,a57443a,a57447a,a57448a,a57449a,a57453a,a57454a,a57457a,a57460a,a57461a,a57462a,a57466a,a57467a,a57471a,a57472a,a57473a,a57477a,a57478a,a57481a,a57484a,a57485a,a57486a,a57490a,a57491a,a57495a,a57496a,a57497a,a57501a,a57502a,a57505a,a57508a,a57509a,a57510a,a57514a,a57515a,a57519a,a57520a,a57521a,a57525a,a57526a,a57529a,a57532a,a57533a,a57534a,a57538a,a57539a,a57543a,a57544a,a57545a,a57549a,a57550a,a57553a,a57556a,a57557a,a57558a,a57562a,a57563a,a57567a,a57568a,a57569a,a57573a,a57574a,a57577a,a57580a,a57581a,a57582a,a57586a,a57587a,a57591a,a57592a,a57593a,a57597a,a57598a,a57601a,a57604a,a57605a,a57606a,a57610a,a57611a,a57615a,a57616a,a57617a,a57621a,a57622a,a57625a,a57628a,a57629a,a57630a,a57634a,a57635a,a57639a,a57640a,a57641a,a57645a,a57646a,a57649a,a57652a,a57653a,a57654a,a57658a,a57659a,a57663a,a57664a,a57665a,a57669a,a57670a,a57673a,a57676a,a57677a,a57678a,a57682a,a57683a,a57687a,a57688a,a57689a,a57693a,a57694a,a57697a,a57700a,a57701a,a57702a,a57706a,a57707a,a57711a,a57712a,a57713a,a57717a,a57718a,a57721a,a57724a,a57725a,a57726a,a57730a,a57731a,a57735a,a57736a,a57737a,a57741a,a57742a,a57745a,a57748a,a57749a,a57750a,a57754a,a57755a,a57759a,a57760a,a57761a,a57765a,a57766a,a57769a,a57772a,a57773a,a57774a,a57778a,a57779a,a57783a,a57784a,a57785a,a57789a,a57790a,a57793a,a57796a,a57797a,a57798a,a57802a,a57803a,a57807a,a57808a,a57809a,a57813a,a57814a,a57817a,a57820a,a57821a,a57822a,a57826a,a57827a,a57831a,a57832a,a57833a,a57837a,a57838a,a57841a,a57844a,a57845a,a57846a,a57850a,a57851a,a57855a,a57856a,a57857a,a57861a,a57862a,a57865a,a57868a,a57869a,a57870a,a57874a,a57875a,a57879a,a57880a,a57881a,a57885a,a57886a,a57889a,a57892a,a57893a,a57894a,a57898a,a57899a,a57903a,a57904a,a57905a,a57909a,a57910a,a57913a,a57916a,a57917a,a57918a,a57922a,a57923a,a57927a,a57928a,a57929a,a57933a,a57934a,a57937a,a57940a,a57941a,a57942a,a57946a,a57947a,a57951a,a57952a,a57953a,a57957a,a57958a,a57961a,a57964a,a57965a,a57966a,a57970a,a57971a,a57975a,a57976a,a57977a,a57981a,a57982a,a57985a,a57988a,a57989a,a57990a,a57994a,a57995a,a57999a,a58000a,a58001a,a58005a,a58006a,a58009a,a58012a,a58013a,a58014a,a58018a,a58019a,a58023a,a58024a,a58025a,a58029a,a58030a,a58033a,a58036a,a58037a,a58038a,a58042a,a58043a,a58047a,a58048a,a58049a,a58053a,a58054a,a58057a,a58060a,a58061a,a58062a,a58066a,a58067a,a58071a,a58072a,a58073a,a58077a,a58078a,a58081a,a58084a,a58085a,a58086a,a58090a,a58091a,a58095a,a58096a,a58097a,a58101a,a58102a,a58105a,a58108a,a58109a,a58110a,a58114a,a58115a,a58119a,a58120a,a58121a,a58125a,a58126a,a58129a,a58132a,a58133a,a58134a,a58138a,a58139a,a58143a,a58144a,a58145a,a58149a,a58150a,a58153a,a58156a,a58157a,a58158a,a58162a,a58163a,a58167a,a58168a,a58169a,a58173a,a58174a,a58177a,a58180a,a58181a,a58182a,a58186a,a58187a,a58191a,a58192a,a58193a,a58197a,a58198a,a58201a,a58204a,a58205a,a58206a,a58210a,a58211a,a58215a,a58216a,a58217a,a58221a,a58222a,a58225a,a58228a,a58229a,a58230a,a58234a,a58235a,a58239a,a58240a,a58241a,a58245a,a58246a,a58249a,a58252a,a58253a,a58254a,a58258a,a58259a,a58263a,a58264a,a58265a,a58269a,a58270a,a58273a,a58276a,a58277a,a58278a,a58282a,a58283a,a58287a,a58288a,a58289a,a58293a,a58294a,a58297a,a58300a,a58301a,a58302a,a58306a,a58307a,a58311a,a58312a,a58313a,a58317a,a58318a,a58321a,a58324a,a58325a,a58326a,a58330a,a58331a,a58335a,a58336a,a58337a,a58341a,a58342a,a58345a,a58348a,a58349a,a58350a,a58354a,a58355a,a58359a,a58360a,a58361a,a58365a,a58366a,a58369a,a58372a,a58373a,a58374a,a58378a,a58379a,a58383a,a58384a,a58385a,a58389a,a58390a,a58393a,a58396a,a58397a,a58398a,a58402a,a58403a,a58407a,a58408a,a58409a,a58413a,a58414a,a58417a,a58420a,a58421a,a58422a,a58426a,a58427a,a58431a,a58432a,a58433a,a58437a,a58438a,a58441a,a58444a,a58445a,a58446a,a58450a,a58451a,a58455a,a58456a,a58457a,a58461a,a58462a,a58465a,a58468a,a58469a,a58470a,a58474a,a58475a,a58479a,a58480a,a58481a,a58485a,a58486a,a58489a,a58492a,a58493a,a58494a,a58498a,a58499a,a58503a,a58504a,a58505a,a58509a,a58510a,a58513a,a58516a,a58517a,a58518a,a58522a,a58523a,a58527a,a58528a,a58529a,a58533a,a58534a,a58537a,a58540a,a58541a,a58542a,a58546a,a58547a,a58551a,a58552a,a58553a,a58557a,a58558a,a58561a,a58564a,a58565a,a58566a,a58570a,a58571a,a58575a,a58576a,a58577a,a58581a,a58582a,a58585a,a58588a,a58589a,a58590a,a58594a,a58595a,a58599a,a58600a,a58601a,a58605a,a58606a,a58609a,a58612a,a58613a,a58614a,a58618a,a58619a,a58623a,a58624a,a58625a,a58629a,a58630a,a58633a,a58636a,a58637a,a58638a,a58642a,a58643a,a58647a,a58648a,a58649a,a58653a,a58654a,a58657a,a58660a,a58661a,a58662a,a58666a,a58667a,a58671a,a58672a,a58673a,a58677a,a58678a,a58681a,a58684a,a58685a,a58686a,a58690a,a58691a,a58695a,a58696a,a58697a,a58701a,a58702a,a58705a,a58708a,a58709a,a58710a,a58714a,a58715a,a58719a,a58720a,a58721a,a58725a,a58726a,a58729a,a58732a,a58733a,a58734a,a58738a,a58739a,a58743a,a58744a,a58745a,a58749a,a58750a,a58753a,a58756a,a58757a,a58758a,a58762a,a58763a,a58767a,a58768a,a58769a,a58773a,a58774a,a58777a,a58780a,a58781a,a58782a,a58786a,a58787a,a58791a,a58792a,a58793a,a58797a,a58798a,a58801a,a58804a,a58805a,a58806a,a58810a,a58811a,a58815a,a58816a,a58817a,a58821a,a58822a,a58825a,a58828a,a58829a,a58830a,a58834a,a58835a,a58839a,a58840a,a58841a,a58845a,a58846a,a58849a,a58852a,a58853a,a58854a,a58858a,a58859a,a58863a,a58864a,a58865a,a58869a,a58870a,a58873a,a58876a,a58877a,a58878a,a58882a,a58883a,a58887a,a58888a,a58889a,a58893a,a58894a,a58897a,a58900a,a58901a,a58902a,a58906a,a58907a,a58911a,a58912a,a58913a,a58917a,a58918a,a58921a,a58924a,a58925a,a58926a,a58930a,a58931a,a58935a,a58936a,a58937a,a58941a,a58942a,a58945a,a58948a,a58949a,a58950a,a58954a,a58955a,a58959a,a58960a,a58961a,a58965a,a58966a,a58969a,a58972a,a58973a,a58974a,a58978a,a58979a,a58983a,a58984a,a58985a,a58989a,a58990a,a58993a,a58996a,a58997a,a58998a,a59002a,a59003a,a59007a,a59008a,a59009a,a59013a,a59014a,a59017a,a59020a,a59021a,a59022a,a59026a,a59027a,a59031a,a59032a,a59033a,a59037a,a59038a,a59041a,a59044a,a59045a,a59046a,a59050a,a59051a,a59055a,a59056a,a59057a,a59061a,a59062a,a59065a,a59068a,a59069a,a59070a,a59074a,a59075a,a59079a,a59080a,a59081a,a59085a,a59086a,a59089a,a59092a,a59093a,a59094a,a59098a,a59099a,a59103a,a59104a,a59105a,a59109a,a59110a,a59113a,a59116a,a59117a,a59118a,a59122a,a59123a,a59127a,a59128a,a59129a,a59133a,a59134a,a59137a,a59140a,a59141a,a59142a,a59146a,a59147a,a59151a,a59152a,a59153a,a59157a,a59158a,a59161a,a59164a,a59165a,a59166a,a59170a,a59171a,a59175a,a59176a,a59177a,a59181a,a59182a,a59185a,a59188a,a59189a,a59190a,a59194a,a59195a,a59199a,a59200a,a59201a,a59205a,a59206a,a59209a,a59212a,a59213a,a59214a,a59218a,a59219a,a59223a,a59224a,a59225a,a59229a,a59230a,a59233a,a59236a,a59237a,a59238a,a59242a,a59243a,a59247a,a59248a,a59249a,a59253a,a59254a,a59257a,a59260a,a59261a,a59262a,a59266a,a59267a,a59271a,a59272a,a59273a,a59277a,a59278a,a59281a,a59284a,a59285a,a59286a,a59290a,a59291a,a59295a,a59296a,a59297a,a59301a,a59302a,a59305a,a59308a,a59309a,a59310a,a59314a,a59315a,a59319a,a59320a,a59321a,a59325a,a59326a,a59329a,a59332a,a59333a,a59334a,a59338a,a59339a,a59343a,a59344a,a59345a,a59349a,a59350a,a59353a,a59356a,a59357a,a59358a,a59362a,a59363a,a59367a,a59368a,a59369a,a59373a,a59374a,a59377a,a59380a,a59381a,a59382a,a59386a,a59387a,a59391a,a59392a,a59393a,a59397a,a59398a,a59401a,a59404a,a59405a,a59406a,a59410a,a59411a,a59415a,a59416a,a59417a,a59421a,a59422a,a59425a,a59428a,a59429a,a59430a,a59434a,a59435a,a59439a,a59440a,a59441a,a59445a,a59446a,a59449a,a59452a,a59453a,a59454a,a59458a,a59459a,a59463a,a59464a,a59465a,a59469a,a59470a,a59473a,a59476a,a59477a,a59478a,a59482a,a59483a,a59487a,a59488a,a59489a,a59493a,a59494a,a59497a,a59500a,a59501a,a59502a,a59506a,a59507a,a59511a,a59512a,a59513a,a59517a,a59518a,a59521a,a59524a,a59525a,a59526a,a59530a,a59531a,a59535a,a59536a,a59537a,a59541a,a59542a,a59545a,a59548a,a59549a,a59550a,a59554a,a59555a,a59559a,a59560a,a59561a,a59565a,a59566a,a59569a,a59572a,a59573a,a59574a,a59578a,a59579a,a59583a,a59584a,a59585a,a59589a,a59590a,a59593a,a59596a,a59597a,a59598a,a59602a,a59603a,a59607a,a59608a,a59609a,a59613a,a59614a,a59617a,a59620a,a59621a,a59622a,a59626a,a59627a,a59631a,a59632a,a59633a,a59637a,a59638a,a59641a,a59644a,a59645a,a59646a,a59650a,a59651a,a59655a,a59656a,a59657a,a59661a,a59662a,a59665a,a59668a,a59669a,a59670a,a59674a,a59675a,a59679a,a59680a,a59681a,a59685a,a59686a,a59689a,a59692a,a59693a,a59694a,a59698a,a59699a,a59703a,a59704a,a59705a,a59709a,a59710a,a59713a,a59716a,a59717a,a59718a,a59722a,a59723a,a59727a,a59728a,a59729a,a59733a,a59734a,a59737a,a59740a,a59741a,a59742a,a59746a,a59747a,a59751a,a59752a,a59753a,a59757a,a59758a,a59761a,a59764a,a59765a,a59766a,a59770a,a59771a,a59775a,a59776a,a59777a,a59781a,a59782a,a59785a,a59788a,a59789a,a59790a,a59794a,a59795a,a59799a,a59800a,a59801a,a59805a,a59806a,a59809a,a59812a,a59813a,a59814a,a59818a,a59819a,a59823a,a59824a,a59825a,a59829a,a59830a,a59833a,a59836a,a59837a,a59838a,a59842a,a59843a,a59847a,a59848a,a59849a,a59853a,a59854a,a59857a,a59860a,a59861a,a59862a,a59866a,a59867a,a59871a,a59872a,a59873a,a59877a,a59878a,a59881a,a59884a,a59885a,a59886a,a59890a,a59891a,a59895a,a59896a,a59897a,a59901a,a59902a,a59905a,a59908a,a59909a,a59910a,a59914a,a59915a,a59919a,a59920a,a59921a,a59925a,a59926a,a59929a,a59932a,a59933a,a59934a,a59938a,a59939a,a59943a,a59944a,a59945a,a59949a,a59950a,a59953a,a59956a,a59957a,a59958a,a59962a,a59963a,a59967a,a59968a,a59969a,a59973a,a59974a,a59977a,a59980a,a59981a,a59982a,a59986a,a59987a,a59991a,a59992a,a59993a,a59997a,a59998a,a60001a,a60004a,a60005a,a60006a,a60010a,a60011a,a60015a,a60016a,a60017a,a60021a,a60022a,a60025a,a60028a,a60029a,a60030a,a60034a,a60035a,a60039a,a60040a,a60041a,a60045a,a60046a,a60049a,a60052a,a60053a,a60054a,a60058a,a60059a,a60063a,a60064a,a60065a,a60069a,a60070a,a60073a,a60076a,a60077a,a60078a,a60082a,a60083a,a60087a,a60088a,a60089a,a60093a,a60094a,a60097a,a60100a,a60101a,a60102a,a60106a,a60107a,a60111a,a60112a,a60113a,a60117a,a60118a,a60121a,a60124a,a60125a,a60126a,a60130a,a60131a,a60135a,a60136a,a60137a,a60141a,a60142a,a60145a,a60148a,a60149a,a60150a,a60154a,a60155a,a60159a,a60160a,a60161a,a60165a,a60166a,a60169a,a60172a,a60173a,a60174a,a60178a,a60179a,a60183a,a60184a,a60185a,a60189a,a60190a,a60193a,a60196a,a60197a,a60198a,a60202a,a60203a,a60207a,a60208a,a60209a,a60213a,a60214a,a60217a,a60220a,a60221a,a60222a,a60226a,a60227a,a60231a,a60232a,a60233a,a60237a,a60238a,a60241a,a60244a,a60245a,a60246a,a60250a,a60251a,a60255a,a60256a,a60257a,a60261a,a60262a,a60265a,a60268a,a60269a,a60270a,a60274a,a60275a,a60279a,a60280a,a60281a,a60285a,a60286a,a60289a,a60292a,a60293a,a60294a,a60298a,a60299a,a60303a,a60304a,a60305a,a60309a,a60310a,a60313a,a60316a,a60317a,a60318a,a60322a,a60323a,a60327a,a60328a,a60329a,a60333a,a60334a,a60337a,a60340a,a60341a,a60342a,a60346a,a60347a,a60351a,a60352a,a60353a,a60357a,a60358a,a60361a,a60364a,a60365a,a60366a,a60370a,a60371a,a60375a,a60376a,a60377a,a60381a,a60382a,a60385a,a60388a,a60389a,a60390a,a60394a,a60395a,a60399a,a60400a,a60401a,a60405a,a60406a,a60409a,a60412a,a60413a,a60414a,a60418a,a60419a,a60423a,a60424a,a60425a,a60429a,a60430a,a60433a,a60436a,a60437a,a60438a,a60442a,a60443a,a60447a,a60448a,a60449a,a60453a,a60454a,a60457a,a60460a,a60461a,a60462a,a60466a,a60467a,a60471a,a60472a,a60473a,a60477a,a60478a,a60481a,a60484a,a60485a,a60486a,a60490a,a60491a,a60495a,a60496a,a60497a,a60501a,a60502a,a60505a,a60508a,a60509a,a60510a,a60514a,a60515a,a60519a,a60520a,a60521a,a60525a,a60526a,a60529a,a60532a,a60533a,a60534a,a60538a,a60539a,a60543a,a60544a,a60545a,a60549a,a60550a,a60553a,a60556a,a60557a,a60558a,a60562a,a60563a,a60567a,a60568a,a60569a,a60573a,a60574a,a60577a,a60580a,a60581a,a60582a,a60586a,a60587a,a60591a,a60592a,a60593a,a60597a,a60598a,a60601a,a60604a,a60605a,a60606a,a60610a,a60611a,a60615a,a60616a,a60617a,a60621a,a60622a,a60625a,a60628a,a60629a,a60630a,a60634a,a60635a,a60639a,a60640a,a60641a,a60645a,a60646a,a60649a,a60652a,a60653a,a60654a,a60658a,a60659a,a60663a,a60664a,a60665a,a60669a,a60670a,a60673a,a60676a,a60677a,a60678a,a60682a,a60683a,a60687a,a60688a,a60689a,a60693a,a60694a,a60697a,a60700a,a60701a,a60702a,a60706a,a60707a,a60711a,a60712a,a60713a,a60717a,a60718a,a60721a,a60724a,a60725a,a60726a,a60730a,a60731a,a60735a,a60736a,a60737a,a60741a,a60742a,a60745a,a60748a,a60749a,a60750a,a60754a,a60755a,a60759a,a60760a,a60761a,a60765a,a60766a,a60769a,a60772a,a60773a,a60774a,a60778a,a60779a,a60783a,a60784a,a60785a,a60789a,a60790a,a60793a,a60796a,a60797a,a60798a,a60802a,a60803a,a60807a,a60808a,a60809a,a60813a,a60814a,a60817a,a60820a,a60821a,a60822a,a60826a,a60827a,a60831a,a60832a,a60833a,a60837a,a60838a,a60841a,a60844a,a60845a,a60846a,a60850a,a60851a,a60855a,a60856a,a60857a,a60861a,a60862a,a60865a,a60868a,a60869a,a60870a,a60874a,a60875a,a60879a,a60880a,a60881a,a60885a,a60886a,a60889a,a60892a,a60893a,a60894a,a60898a,a60899a,a60903a,a60904a,a60905a,a60909a,a60910a,a60913a,a60916a,a60917a,a60918a,a60922a,a60923a,a60927a,a60928a,a60929a,a60933a,a60934a,a60937a,a60940a,a60941a,a60942a,a60946a,a60947a,a60951a,a60952a,a60953a,a60957a,a60958a,a60961a,a60964a,a60965a,a60966a,a60970a,a60971a,a60975a,a60976a,a60977a,a60981a,a60982a,a60985a,a60988a,a60989a,a60990a,a60994a,a60995a,a60999a,a61000a,a61001a,a61005a,a61006a,a61009a,a61012a,a61013a,a61014a,a61018a,a61019a,a61023a,a61024a,a61025a,a61029a,a61030a,a61033a,a61036a,a61037a,a61038a,a61042a,a61043a,a61047a,a61048a,a61049a,a61053a,a61054a,a61057a,a61060a,a61061a,a61062a,a61066a,a61067a,a61071a,a61072a,a61073a,a61077a,a61078a,a61081a,a61084a,a61085a,a61086a,a61090a,a61091a,a61095a,a61096a,a61097a,a61101a,a61102a,a61105a,a61108a,a61109a,a61110a,a61114a,a61115a,a61119a,a61120a,a61121a,a61125a,a61126a,a61129a,a61132a,a61133a,a61134a,a61138a,a61139a,a61143a,a61144a,a61145a,a61149a,a61150a,a61153a,a61156a,a61157a,a61158a,a61162a,a61163a,a61167a,a61168a,a61169a,a61173a,a61174a,a61177a,a61180a,a61181a,a61182a,a61186a,a61187a,a61191a,a61192a,a61193a,a61197a,a61198a,a61201a,a61204a,a61205a,a61206a,a61210a,a61211a,a61215a,a61216a,a61217a,a61221a,a61222a,a61225a,a61228a,a61229a,a61230a,a61234a,a61235a,a61239a,a61240a,a61241a,a61245a,a61246a,a61249a,a61252a,a61253a,a61254a,a61258a,a61259a,a61263a,a61264a,a61265a,a61269a,a61270a,a61273a,a61276a,a61277a,a61278a,a61282a,a61283a,a61287a,a61288a,a61289a,a61293a,a61294a,a61297a,a61300a,a61301a,a61302a,a61306a,a61307a,a61311a,a61312a,a61313a,a61317a,a61318a,a61321a,a61324a,a61325a,a61326a,a61330a,a61331a,a61335a,a61336a,a61337a,a61341a,a61342a,a61345a,a61348a,a61349a,a61350a,a61354a,a61355a,a61359a,a61360a,a61361a,a61365a,a61366a,a61369a,a61372a,a61373a,a61374a,a61378a,a61379a,a61383a,a61384a,a61385a,a61389a,a61390a,a61393a,a61396a,a61397a,a61398a,a61402a,a61403a,a61407a,a61408a,a61409a,a61413a,a61414a,a61417a,a61420a,a61421a,a61422a,a61426a,a61427a,a61431a,a61432a,a61433a,a61437a,a61438a,a61441a,a61444a,a61445a,a61446a,a61450a,a61451a,a61455a,a61456a,a61457a,a61461a,a61462a,a61465a,a61468a,a61469a,a61470a,a61474a,a61475a,a61479a,a61480a,a61481a,a61485a,a61486a,a61489a,a61492a,a61493a,a61494a,a61498a,a61499a,a61503a,a61504a,a61505a,a61509a,a61510a,a61513a,a61516a,a61517a,a61518a,a61522a,a61523a,a61527a,a61528a,a61529a,a61533a,a61534a,a61537a,a61540a,a61541a,a61542a,a61546a,a61547a,a61551a,a61552a,a61553a,a61557a,a61558a,a61561a,a61564a,a61565a,a61566a,a61570a,a61571a,a61575a,a61576a,a61577a,a61581a,a61582a,a61585a,a61588a,a61589a,a61590a,a61594a,a61595a,a61599a,a61600a,a61601a,a61605a,a61606a,a61609a,a61612a,a61613a,a61614a,a61618a,a61619a,a61623a,a61624a,a61625a,a61629a,a61630a,a61633a,a61636a,a61637a,a61638a,a61642a,a61643a,a61647a,a61648a,a61649a,a61653a,a61654a,a61657a,a61660a,a61661a,a61662a,a61666a,a61667a,a61671a,a61672a,a61673a,a61677a,a61678a,a61681a,a61684a,a61685a,a61686a,a61690a,a61691a,a61695a,a61696a,a61697a,a61701a,a61702a,a61705a,a61708a,a61709a,a61710a,a61714a,a61715a,a61719a,a61720a,a61721a,a61725a,a61726a,a61729a,a61732a,a61733a,a61734a,a61738a,a61739a,a61743a,a61744a,a61745a,a61749a,a61750a,a61753a,a61756a,a61757a,a61758a,a61762a,a61763a,a61767a,a61768a,a61769a,a61773a,a61774a,a61777a,a61780a,a61781a,a61782a,a61786a,a61787a,a61791a,a61792a,a61793a,a61797a,a61798a,a61801a,a61804a,a61805a,a61806a,a61810a,a61811a,a61815a,a61816a,a61817a,a61821a,a61822a,a61825a,a61828a,a61829a,a61830a,a61834a,a61835a,a61839a,a61840a,a61841a,a61845a,a61846a,a61849a,a61852a,a61853a,a61854a,a61858a,a61859a,a61863a,a61864a,a61865a,a61869a,a61870a,a61873a,a61876a,a61877a,a61878a,a61882a,a61883a,a61887a,a61888a,a61889a,a61893a,a61894a,a61897a,a61900a,a61901a,a61902a,a61906a,a61907a,a61911a,a61912a,a61913a,a61917a,a61918a,a61921a,a61924a,a61925a,a61926a,a61930a,a61931a,a61935a,a61936a,a61937a,a61941a,a61942a,a61945a,a61948a,a61949a,a61950a,a61954a,a61955a,a61959a,a61960a,a61961a,a61965a,a61966a,a61969a,a61972a,a61973a,a61974a,a61978a,a61979a,a61983a,a61984a,a61985a,a61989a,a61990a,a61993a,a61996a,a61997a,a61998a,a62002a,a62003a,a62007a,a62008a,a62009a,a62013a,a62014a,a62017a,a62020a,a62021a,a62022a,a62026a,a62027a,a62031a,a62032a,a62033a,a62037a,a62038a,a62041a,a62044a,a62045a,a62046a,a62050a,a62051a,a62055a,a62056a,a62057a,a62061a,a62062a,a62065a,a62068a,a62069a,a62070a,a62074a,a62075a,a62079a,a62080a,a62081a,a62085a,a62086a,a62089a,a62092a,a62093a,a62094a,a62098a,a62099a,a62103a,a62104a,a62105a,a62109a,a62110a,a62113a,a62116a,a62117a,a62118a,a62122a,a62123a,a62127a,a62128a,a62129a,a62133a,a62134a,a62137a,a62140a,a62141a,a62142a,a62146a,a62147a,a62151a,a62152a,a62153a,a62157a,a62158a,a62161a,a62164a,a62165a,a62166a,a62170a,a62171a,a62175a,a62176a,a62177a,a62181a,a62182a,a62185a,a62188a,a62189a,a62190a,a62194a,a62195a,a62199a,a62200a,a62201a,a62205a,a62206a,a62209a,a62212a,a62213a,a62214a,a62218a,a62219a,a62223a,a62224a,a62225a,a62229a,a62230a,a62233a,a62236a,a62237a,a62238a,a62242a,a62243a,a62247a,a62248a,a62249a,a62253a,a62254a,a62257a,a62260a,a62261a,a62262a,a62266a,a62267a,a62271a,a62272a,a62273a,a62277a,a62278a,a62281a,a62284a,a62285a,a62286a,a62290a,a62291a,a62295a,a62296a,a62297a,a62301a,a62302a,a62305a,a62308a,a62309a,a62310a,a62314a,a62315a,a62319a,a62320a,a62321a,a62325a,a62326a,a62329a,a62332a,a62333a,a62334a,a62338a,a62339a,a62343a,a62344a,a62345a,a62349a,a62350a,a62353a,a62356a,a62357a,a62358a,a62362a,a62363a,a62367a,a62368a,a62369a,a62373a,a62374a,a62377a,a62380a,a62381a,a62382a,a62386a,a62387a,a62391a,a62392a,a62393a,a62397a,a62398a,a62401a,a62404a,a62405a,a62406a,a62410a,a62411a,a62415a,a62416a,a62417a,a62421a,a62422a,a62425a,a62428a,a62429a,a62430a,a62434a,a62435a,a62439a,a62440a,a62441a,a62445a,a62446a,a62449a,a62452a,a62453a,a62454a,a62458a,a62459a,a62463a,a62464a,a62465a,a62469a,a62470a,a62473a,a62476a,a62477a,a62478a,a62482a,a62483a,a62487a,a62488a,a62489a,a62493a,a62494a,a62497a,a62500a,a62501a,a62502a,a62506a,a62507a,a62511a,a62512a,a62513a,a62517a,a62518a,a62521a,a62524a,a62525a,a62526a,a62530a,a62531a,a62535a,a62536a,a62537a,a62541a,a62542a,a62545a,a62548a,a62549a,a62550a,a62554a,a62555a,a62559a,a62560a,a62561a,a62565a,a62566a,a62569a,a62572a,a62573a,a62574a,a62578a,a62579a,a62583a,a62584a,a62585a,a62589a,a62590a,a62593a,a62596a,a62597a,a62598a,a62602a,a62603a,a62607a,a62608a,a62609a,a62613a,a62614a,a62617a,a62620a,a62621a,a62622a,a62626a,a62627a,a62631a,a62632a,a62633a,a62637a,a62638a,a62641a,a62644a,a62645a,a62646a,a62650a,a62651a,a62655a,a62656a,a62657a,a62661a,a62662a,a62665a,a62668a,a62669a,a62670a,a62674a,a62675a,a62679a,a62680a,a62681a,a62685a,a62686a,a62689a,a62692a,a62693a,a62694a,a62698a,a62699a,a62703a,a62704a,a62705a,a62709a,a62710a,a62713a,a62716a,a62717a,a62718a,a62722a,a62723a,a62727a,a62728a,a62729a,a62733a,a62734a,a62737a,a62740a,a62741a,a62742a,a62746a,a62747a,a62751a,a62752a,a62753a,a62757a,a62758a,a62761a,a62764a,a62765a,a62766a,a62770a,a62771a,a62775a,a62776a,a62777a,a62781a,a62782a,a62785a,a62788a,a62789a,a62790a,a62794a,a62795a,a62799a,a62800a,a62801a,a62805a,a62806a,a62809a,a62812a,a62813a,a62814a,a62818a,a62819a,a62823a,a62824a,a62825a,a62829a,a62830a,a62833a,a62836a,a62837a,a62838a,a62842a,a62843a,a62847a,a62848a,a62849a,a62853a,a62854a,a62857a,a62860a,a62861a,a62862a,a62866a,a62867a,a62871a,a62872a,a62873a,a62877a,a62878a,a62881a,a62884a,a62885a,a62886a,a62890a,a62891a,a62895a,a62896a,a62897a,a62901a,a62902a,a62905a,a62908a,a62909a,a62910a,a62914a,a62915a,a62919a,a62920a,a62921a,a62925a,a62926a,a62929a,a62932a,a62933a,a62934a,a62938a,a62939a,a62943a,a62944a,a62945a,a62949a,a62950a,a62953a,a62956a,a62957a,a62958a,a62962a,a62963a,a62967a,a62968a,a62969a,a62973a,a62974a,a62977a,a62980a,a62981a,a62982a,a62986a,a62987a,a62991a,a62992a,a62993a,a62997a,a62998a,a63001a,a63004a,a63005a,a63006a,a63010a,a63011a,a63015a,a63016a,a63017a,a63021a,a63022a,a63025a,a63028a,a63029a,a63030a,a63034a,a63035a,a63039a,a63040a,a63041a,a63045a,a63046a,a63049a,a63052a,a63053a,a63054a,a63058a,a63059a,a63063a,a63064a,a63065a,a63069a,a63070a,a63073a,a63076a,a63077a,a63078a,a63082a,a63083a,a63087a,a63088a,a63089a,a63093a,a63094a,a63097a,a63100a,a63101a,a63102a,a63106a,a63107a,a63111a,a63112a,a63113a,a63117a,a63118a,a63121a,a63124a,a63125a,a63126a,a63130a,a63131a,a63135a,a63136a,a63137a,a63141a,a63142a,a63145a,a63148a,a63149a,a63150a,a63154a,a63155a,a63159a,a63160a,a63161a,a63165a,a63166a,a63169a,a63172a,a63173a,a63174a,a63178a,a63179a,a63183a,a63184a,a63185a,a63189a,a63190a,a63193a,a63196a,a63197a,a63198a,a63202a,a63203a,a63207a,a63208a,a63209a,a63213a,a63214a,a63217a,a63220a,a63221a,a63222a,a63226a,a63227a,a63231a,a63232a,a63233a,a63237a,a63238a,a63241a,a63244a,a63245a,a63246a,a63250a,a63251a,a63255a,a63256a,a63257a,a63261a,a63262a,a63265a,a63268a,a63269a,a63270a,a63274a,a63275a,a63279a,a63280a,a63281a,a63285a,a63286a,a63289a,a63292a,a63293a,a63294a,a63298a,a63299a,a63303a,a63304a,a63305a,a63309a,a63310a,a63313a,a63316a,a63317a,a63318a,a63322a,a63323a,a63327a,a63328a,a63329a,a63333a,a63334a,a63337a,a63340a,a63341a,a63342a,a63346a,a63347a,a63351a,a63352a,a63353a,a63357a,a63358a,a63361a,a63364a,a63365a,a63366a,a63370a,a63371a,a63375a,a63376a,a63377a,a63381a,a63382a,a63385a,a63388a,a63389a,a63390a,a63394a,a63395a,a63399a,a63400a,a63401a,a63405a,a63406a,a63409a,a63412a,a63413a,a63414a,a63418a,a63419a,a63423a,a63424a,a63425a,a63429a,a63430a,a63433a,a63436a,a63437a,a63438a,a63442a,a63443a,a63447a,a63448a,a63449a,a63453a,a63454a,a63457a,a63460a,a63461a,a63462a,a63466a,a63467a,a63471a,a63472a,a63473a,a63477a,a63478a,a63481a,a63484a,a63485a,a63486a,a63490a,a63491a,a63495a,a63496a,a63497a,a63501a,a63502a,a63505a,a63508a,a63509a,a63510a,a63514a,a63515a,a63519a,a63520a,a63521a,a63525a,a63526a,a63529a,a63532a,a63533a,a63534a,a63538a,a63539a,a63543a,a63544a,a63545a,a63549a,a63550a,a63553a,a63556a,a63557a,a63558a,a63562a,a63563a,a63567a,a63568a,a63569a,a63573a,a63574a,a63577a,a63580a,a63581a,a63582a,a63586a,a63587a,a63591a,a63592a,a63593a,a63597a,a63598a,a63601a,a63604a,a63605a,a63606a,a63610a,a63611a,a63615a,a63616a,a63617a,a63621a,a63622a,a63625a,a63628a,a63629a,a63630a,a63634a,a63635a,a63639a,a63640a,a63641a,a63645a,a63646a,a63649a,a63652a,a63653a,a63654a,a63658a,a63659a,a63663a,a63664a,a63665a,a63669a,a63670a,a63673a,a63676a,a63677a,a63678a,a63682a,a63683a,a63687a,a63688a,a63689a,a63693a,a63694a,a63697a,a63700a,a63701a,a63702a,a63706a,a63707a,a63711a,a63712a,a63713a,a63717a,a63718a,a63721a,a63724a,a63725a,a63726a,a63730a,a63731a,a63735a,a63736a,a63737a,a63741a,a63742a,a63745a,a63748a,a63749a,a63750a,a63754a,a63755a,a63759a,a63760a,a63761a,a63765a,a63766a,a63769a,a63772a,a63773a,a63774a,a63778a,a63779a,a63783a,a63784a,a63785a,a63789a,a63790a,a63793a,a63796a,a63797a,a63798a,a63802a,a63803a,a63807a,a63808a,a63809a,a63813a,a63814a,a63817a,a63820a,a63821a,a63822a,a63826a,a63827a,a63831a,a63832a,a63833a,a63837a,a63838a,a63841a,a63844a,a63845a,a63846a,a63850a,a63851a,a63855a,a63856a,a63857a,a63861a,a63862a,a63865a,a63868a,a63869a,a63870a,a63874a,a63875a,a63879a,a63880a,a63881a,a63885a,a63886a,a63889a,a63892a,a63893a,a63894a,a63898a,a63899a,a63903a,a63904a,a63905a,a63909a,a63910a,a63913a,a63916a,a63917a,a63918a,a63922a,a63923a,a63927a,a63928a,a63929a,a63933a,a63934a,a63937a,a63940a,a63941a,a63942a,a63946a,a63947a,a63951a,a63952a,a63953a,a63957a,a63958a,a63961a,a63964a,a63965a,a63966a,a63970a,a63971a,a63975a,a63976a,a63977a,a63981a,a63982a,a63985a,a63988a,a63989a,a63990a,a63994a,a63995a,a63999a,a64000a,a64001a,a64005a,a64006a,a64009a,a64012a,a64013a,a64014a,a64018a,a64019a,a64023a,a64024a,a64025a,a64029a,a64030a,a64033a,a64036a,a64037a,a64038a,a64042a,a64043a,a64047a,a64048a,a64049a,a64053a,a64054a,a64057a,a64060a,a64061a,a64062a,a64066a,a64067a,a64071a,a64072a,a64073a,a64077a,a64078a,a64081a,a64084a,a64085a,a64086a,a64090a,a64091a,a64095a,a64096a,a64097a,a64101a,a64102a,a64105a,a64108a,a64109a,a64110a,a64114a,a64115a,a64119a,a64120a,a64121a,a64125a,a64126a,a64129a,a64132a,a64133a,a64134a,a64138a,a64139a,a64143a,a64144a,a64145a,a64149a,a64150a,a64153a,a64156a,a64157a,a64158a,a64162a,a64163a,a64167a,a64168a,a64169a,a64173a,a64174a,a64177a,a64180a,a64181a,a64182a,a64186a,a64187a,a64191a,a64192a,a64193a,a64197a,a64198a,a64201a,a64204a,a64205a,a64206a,a64210a,a64211a,a64215a,a64216a,a64217a,a64221a,a64222a,a64225a,a64228a,a64229a,a64230a,a64234a,a64235a,a64239a,a64240a,a64241a,a64245a,a64246a,a64249a,a64252a,a64253a,a64254a,a64258a,a64259a,a64263a,a64264a,a64265a,a64269a,a64270a,a64273a,a64276a,a64277a,a64278a,a64282a,a64283a,a64287a,a64288a,a64289a,a64293a,a64294a,a64297a,a64300a,a64301a,a64302a,a64306a,a64307a,a64311a,a64312a,a64313a,a64317a,a64318a,a64321a,a64324a,a64325a,a64326a,a64330a,a64331a,a64335a,a64336a,a64337a,a64341a,a64342a,a64345a,a64348a,a64349a,a64350a,a64354a,a64355a,a64359a,a64360a,a64361a,a64365a,a64366a,a64369a,a64372a,a64373a,a64374a,a64378a,a64379a,a64383a,a64384a,a64385a,a64389a,a64390a,a64393a,a64396a,a64397a,a64398a,a64402a,a64403a,a64407a,a64408a,a64409a,a64413a,a64414a,a64417a,a64420a,a64421a,a64422a,a64426a,a64427a,a64431a,a64432a,a64433a,a64437a,a64438a,a64441a,a64444a,a64445a,a64446a,a64450a,a64451a,a64455a,a64456a,a64457a,a64461a,a64462a,a64465a,a64468a,a64469a,a64470a,a64474a,a64475a,a64479a,a64480a,a64481a,a64485a,a64486a,a64489a,a64492a,a64493a,a64494a,a64498a,a64499a,a64503a,a64504a,a64505a,a64509a,a64510a,a64513a,a64516a,a64517a,a64518a,a64522a,a64523a,a64527a,a64528a,a64529a,a64533a,a64534a,a64537a,a64540a,a64541a,a64542a,a64546a,a64547a,a64551a,a64552a,a64553a,a64557a,a64558a,a64561a,a64564a,a64565a,a64566a,a64570a,a64571a,a64575a,a64576a,a64577a,a64581a,a64582a,a64585a,a64588a,a64589a,a64590a,a64594a,a64595a,a64599a,a64600a,a64601a,a64605a,a64606a,a64609a,a64612a,a64613a,a64614a,a64618a,a64619a,a64623a,a64624a,a64625a,a64629a,a64630a,a64633a,a64636a,a64637a,a64638a,a64642a,a64643a,a64646a,a64649a,a64650a,a64651a,a64655a,a64656a,a64659a,a64662a,a64663a,a64664a,a64668a,a64669a,a64672a,a64675a,a64676a,a64677a,a64681a,a64682a,a64685a,a64688a,a64689a,a64690a,a64694a,a64695a,a64698a,a64701a,a64702a,a64703a,a64707a,a64708a,a64711a,a64714a,a64715a,a64716a,a64720a,a64721a,a64724a,a64727a,a64728a,a64729a,a64733a,a64734a,a64737a,a64740a,a64741a,a64742a,a64746a,a64747a,a64750a,a64753a,a64754a,a64755a,a64759a,a64760a,a64763a,a64766a,a64767a,a64768a,a64772a,a64773a,a64776a,a64779a,a64780a,a64781a,a64785a,a64786a,a64789a,a64792a,a64793a,a64794a,a64798a,a64799a,a64802a,a64805a,a64806a,a64807a,a64811a,a64812a,a64815a,a64818a,a64819a,a64820a,a64824a,a64825a,a64828a,a64831a,a64832a,a64833a,a64837a,a64838a,a64841a,a64844a,a64845a,a64846a,a64850a,a64851a,a64854a,a64857a,a64858a,a64859a,a64863a,a64864a,a64867a,a64870a,a64871a,a64872a,a64876a,a64877a,a64880a,a64883a,a64884a,a64885a,a64889a,a64890a,a64893a,a64896a,a64897a,a64898a,a64902a,a64903a,a64906a,a64909a,a64910a,a64911a,a64915a,a64916a,a64919a,a64922a,a64923a,a64924a,a64928a,a64929a,a64932a,a64935a,a64936a,a64937a,a64941a,a64942a,a64945a,a64948a,a64949a,a64950a,a64954a,a64955a,a64958a,a64961a,a64962a,a64963a,a64967a,a64968a,a64971a,a64974a,a64975a,a64976a,a64980a,a64981a,a64984a,a64987a,a64988a,a64989a,a64993a,a64994a,a64997a,a65000a,a65001a,a65002a,a65006a,a65007a,a65010a,a65013a,a65014a,a65015a,a65019a,a65020a,a65023a,a65026a,a65027a,a65028a,a65032a,a65033a,a65036a,a65039a,a65040a,a65041a,a65045a,a65046a,a65049a,a65052a,a65053a,a65054a,a65058a,a65059a,a65062a,a65065a,a65066a,a65067a,a65071a,a65072a,a65075a,a65078a,a65079a,a65080a,a65084a,a65085a,a65088a,a65091a,a65092a,a65093a,a65097a,a65098a,a65101a,a65104a,a65105a,a65106a,a65110a,a65111a,a65114a,a65117a,a65118a,a65119a,a65123a,a65124a,a65127a,a65130a,a65131a,a65132a,a65136a,a65137a,a65140a,a65143a,a65144a,a65145a,a65149a,a65150a,a65153a,a65156a,a65157a,a65158a,a65162a,a65163a,a65166a,a65169a,a65170a,a65171a,a65175a,a65176a,a65179a,a65182a,a65183a,a65184a,a65188a,a65189a,a65192a,a65195a,a65196a,a65197a,a65201a,a65202a,a65205a,a65208a,a65209a,a65210a,a65214a,a65215a,a65218a,a65221a,a65222a,a65223a,a65227a,a65228a,a65231a,a65234a,a65235a,a65236a,a65240a,a65241a,a65244a,a65247a,a65248a,a65249a,a65253a,a65254a,a65257a,a65260a,a65261a,a65262a,a65266a,a65267a,a65270a,a65273a,a65274a,a65275a,a65279a,a65280a,a65283a,a65286a,a65287a,a65288a,a65292a,a65293a,a65296a,a65299a,a65300a,a65301a,a65305a,a65306a,a65309a,a65312a,a65313a,a65314a,a65318a,a65319a,a65322a,a65325a,a65326a,a65327a,a65331a,a65332a,a65335a,a65338a,a65339a,a65340a,a65344a,a65345a,a65348a,a65351a,a65352a,a65353a,a65357a,a65358a,a65361a,a65364a,a65365a,a65366a,a65370a,a65371a,a65374a,a65377a,a65378a,a65379a,a65383a,a65384a,a65387a,a65390a,a65391a,a65392a,a65396a,a65397a,a65400a,a65403a,a65404a,a65405a,a65409a,a65410a,a65413a,a65416a,a65417a,a65418a,a65422a,a65423a,a65426a,a65429a,a65430a,a65431a,a65435a,a65436a,a65439a,a65442a,a65443a,a65444a,a65448a,a65449a,a65452a,a65455a,a65456a,a65457a,a65461a,a65462a,a65465a,a65468a,a65469a,a65470a,a65474a,a65475a,a65478a,a65481a,a65482a,a65483a,a65487a,a65488a,a65491a,a65494a,a65495a,a65496a,a65500a,a65501a,a65504a,a65507a,a65508a,a65509a,a65513a,a65514a,a65517a,a65520a,a65521a,a65522a,a65526a,a65527a,a65530a,a65533a,a65534a,a65535a,a65539a,a65540a,a65543a,a65546a,a65547a,a65548a,a65552a,a65553a,a65556a,a65559a,a65560a,a65561a,a65565a,a65566a,a65569a,a65572a,a65573a,a65574a,a65578a,a65579a,a65582a,a65585a,a65586a,a65587a,a65591a,a65592a,a65595a,a65598a,a65599a,a65600a,a65604a,a65605a,a65608a,a65611a,a65612a,a65613a,a65617a,a65618a,a65621a,a65624a,a65625a,a65626a,a65630a,a65631a,a65634a,a65637a,a65638a,a65639a,a65643a,a65644a,a65647a,a65650a,a65651a,a65652a,a65656a,a65657a,a65660a,a65663a,a65664a,a65665a,a65669a,a65670a,a65673a,a65676a,a65677a,a65678a,a65682a,a65683a,a65686a,a65689a,a65690a,a65691a,a65695a,a65696a,a65699a,a65702a,a65703a,a65704a,a65708a,a65709a,a65712a,a65715a,a65716a,a65717a,a65721a,a65722a,a65725a,a65728a,a65729a,a65730a,a65734a,a65735a,a65738a,a65741a,a65742a,a65743a,a65747a,a65748a,a65751a,a65754a,a65755a,a65756a,a65760a,a65761a,a65764a,a65767a,a65768a,a65769a,a65773a,a65774a,a65777a,a65780a,a65781a,a65782a,a65786a,a65787a,a65790a,a65793a,a65794a,a65795a,a65799a,a65800a,a65803a,a65806a,a65807a,a65808a,a65812a,a65813a,a65816a,a65819a,a65820a,a65821a,a65825a,a65826a,a65829a,a65832a,a65833a,a65834a,a65838a,a65839a,a65842a,a65845a,a65846a,a65847a,a65851a,a65852a,a65855a,a65858a,a65859a,a65860a,a65864a,a65865a,a65868a,a65871a,a65872a,a65873a,a65877a,a65878a,a65881a,a65884a,a65885a,a65886a,a65890a,a65891a,a65894a,a65897a,a65898a,a65899a,a65903a,a65904a,a65907a,a65910a,a65911a,a65912a,a65916a,a65917a,a65920a,a65923a,a65924a,a65925a,a65929a,a65930a,a65933a,a65936a,a65937a,a65938a,a65942a,a65943a,a65946a,a65949a,a65950a,a65951a,a65955a,a65956a,a65959a,a65962a,a65963a,a65964a,a65968a,a65969a,a65972a,a65975a,a65976a,a65977a,a65981a,a65982a,a65985a,a65988a,a65989a,a65990a,a65994a,a65995a,a65998a,a66001a,a66002a,a66003a,a66007a,a66008a,a66011a,a66014a,a66015a,a66016a,a66020a,a66021a,a66024a,a66027a,a66028a,a66029a,a66033a,a66034a,a66037a,a66040a,a66041a,a66042a,a66046a,a66047a,a66050a,a66053a,a66054a,a66055a,a66059a,a66060a,a66063a,a66066a,a66067a,a66068a,a66072a,a66073a,a66076a,a66079a,a66080a,a66081a,a66085a,a66086a,a66089a,a66092a,a66093a,a66094a,a66098a,a66099a,a66102a,a66105a,a66106a,a66107a,a66111a,a66112a,a66115a,a66118a,a66119a,a66120a,a66124a,a66125a,a66128a,a66131a,a66132a,a66133a,a66137a,a66138a,a66141a,a66144a,a66145a,a66146a,a66150a,a66151a,a66154a,a66157a,a66158a,a66159a,a66163a,a66164a,a66167a,a66170a,a66171a,a66172a,a66176a,a66177a,a66180a,a66183a,a66184a,a66185a,a66189a,a66190a,a66193a,a66196a,a66197a,a66198a,a66202a,a66203a,a66206a,a66209a,a66210a,a66211a,a66215a,a66216a,a66219a,a66222a,a66223a,a66224a,a66228a,a66229a,a66232a,a66235a,a66236a,a66237a,a66241a,a66242a,a66245a,a66248a,a66249a,a66250a,a66254a,a66255a,a66258a,a66261a,a66262a,a66263a,a66267a,a66268a,a66271a,a66274a,a66275a,a66276a,a66280a,a66281a,a66284a,a66287a,a66288a,a66289a,a66293a,a66294a,a66297a,a66300a,a66301a,a66302a,a66306a,a66307a,a66310a,a66313a,a66314a,a66315a,a66319a,a66320a,a66323a,a66326a,a66327a,a66328a,a66332a,a66333a,a66336a,a66339a,a66340a,a66341a,a66345a,a66346a,a66349a,a66352a,a66353a,a66354a,a66358a,a66359a,a66362a,a66365a,a66366a,a66367a,a66371a,a66372a,a66375a,a66378a,a66379a,a66380a,a66384a,a66385a,a66388a,a66391a,a66392a,a66393a,a66397a,a66398a,a66401a,a66404a,a66405a,a66406a,a66410a,a66411a,a66414a,a66417a,a66418a,a66419a,a66423a,a66424a,a66427a,a66430a,a66431a,a66432a,a66436a,a66437a,a66440a,a66443a,a66444a,a66445a,a66449a,a66450a,a66453a,a66456a,a66457a,a66458a,a66462a,a66463a,a66466a,a66469a,a66470a,a66471a,a66475a,a66476a,a66479a,a66482a,a66483a,a66484a,a66488a,a66489a,a66492a,a66495a,a66496a,a66497a,a66501a,a66502a,a66505a,a66508a,a66509a,a66510a,a66514a,a66515a,a66518a,a66521a,a66522a,a66523a,a66527a,a66528a,a66531a,a66534a,a66535a,a66536a,a66540a,a66541a,a66544a,a66547a,a66548a,a66549a,a66553a,a66554a,a66557a,a66560a,a66561a,a66562a,a66566a,a66567a,a66570a,a66573a,a66574a,a66575a,a66579a,a66580a,a66583a,a66586a,a66587a,a66588a,a66592a,a66593a,a66596a,a66599a,a66600a,a66601a,a66605a,a66606a,a66609a,a66612a,a66613a,a66614a,a66618a,a66619a,a66622a,a66625a,a66626a,a66627a,a66631a,a66632a,a66635a,a66638a,a66639a,a66640a,a66644a,a66645a,a66648a,a66651a,a66652a,a66653a,a66657a,a66658a,a66661a,a66664a,a66665a,a66666a,a66670a,a66671a,a66674a,a66677a,a66678a,a66679a,a66683a,a66684a,a66687a,a66690a,a66691a,a66692a,a66696a,a66697a,a66700a,a66703a,a66704a,a66705a,a66709a,a66710a,a66713a,a66716a,a66717a,a66718a,a66722a,a66723a,a66726a,a66729a,a66730a,a66731a,a66735a,a66736a,a66739a,a66742a,a66743a,a66744a,a66748a,a66749a,a66752a,a66755a,a66756a,a66757a,a66761a,a66762a,a66765a,a66768a,a66769a,a66770a,a66774a,a66775a,a66778a,a66781a,a66782a,a66783a,a66787a,a66788a,a66791a,a66794a,a66795a,a66796a,a66800a,a66801a,a66804a,a66807a,a66808a,a66809a,a66813a,a66814a,a66817a,a66820a,a66821a,a66822a,a66826a,a66827a,a66830a,a66833a,a66834a,a66835a,a66839a,a66840a,a66843a,a66846a,a66847a,a66848a,a66852a,a66853a,a66856a,a66859a,a66860a,a66861a,a66865a,a66866a,a66869a,a66872a,a66873a,a66874a,a66878a,a66879a,a66882a,a66885a,a66886a,a66887a,a66891a,a66892a,a66895a,a66898a,a66899a,a66900a,a66904a,a66905a,a66908a,a66911a,a66912a,a66913a,a66917a,a66918a,a66921a,a66924a,a66925a,a66926a,a66930a,a66931a,a66934a,a66937a,a66938a,a66939a,a66943a,a66944a,a66947a,a66950a,a66951a,a66952a,a66956a,a66957a,a66960a,a66963a,a66964a,a66965a,a66969a,a66970a,a66973a,a66976a,a66977a,a66978a,a66982a,a66983a,a66986a,a66989a,a66990a,a66991a,a66995a,a66996a,a66999a,a67002a,a67003a,a67004a,a67008a,a67009a,a67012a,a67015a,a67016a,a67017a,a67021a,a67022a,a67025a,a67028a,a67029a,a67030a,a67034a,a67035a,a67038a,a67041a,a67042a,a67043a,a67047a,a67048a,a67051a,a67054a,a67055a,a67056a,a67060a,a67061a,a67064a,a67067a,a67068a,a67069a,a67073a,a67074a,a67077a,a67080a,a67081a,a67082a,a67086a,a67087a,a67090a,a67093a,a67094a,a67095a,a67099a,a67100a,a67103a,a67106a,a67107a,a67108a,a67112a,a67113a,a67116a,a67119a,a67120a,a67121a,a67125a,a67126a,a67129a,a67132a,a67133a,a67134a,a67138a,a67139a,a67142a,a67145a,a67146a,a67147a,a67151a,a67152a,a67155a,a67158a,a67159a,a67160a,a67164a,a67165a,a67168a,a67171a,a67172a,a67173a,a67177a,a67178a,a67181a,a67184a,a67185a,a67186a,a67190a,a67191a,a67194a,a67197a,a67198a,a67199a,a67203a,a67204a,a67207a,a67210a,a67211a,a67212a,a67216a,a67217a,a67220a,a67223a,a67224a,a67225a,a67229a,a67230a,a67233a,a67236a,a67237a,a67238a,a67242a,a67243a,a67246a,a67249a,a67250a,a67251a,a67255a,a67256a,a67259a,a67262a,a67263a,a67264a,a67268a,a67269a,a67272a,a67275a,a67276a,a67277a,a67281a,a67282a,a67285a,a67288a,a67289a,a67290a,a67294a,a67295a,a67298a,a67301a,a67302a,a67303a,a67307a,a67308a,a67311a,a67314a,a67315a,a67316a,a67320a,a67321a,a67324a,a67327a,a67328a,a67329a,a67333a,a67334a,a67337a,a67340a,a67341a,a67342a,a67346a,a67347a,a67350a,a67353a,a67354a,a67355a,a67359a,a67360a,a67363a,a67366a,a67367a,a67368a,a67372a,a67373a,a67376a,a67379a,a67380a,a67381a,a67385a,a67386a,a67389a,a67392a,a67393a,a67394a,a67398a,a67399a,a67402a,a67405a,a67406a,a67407a,a67411a,a67412a,a67415a,a67418a,a67419a,a67420a,a67424a,a67425a,a67428a,a67431a,a67432a,a67433a,a67437a,a67438a,a67441a,a67444a,a67445a,a67446a,a67450a,a67451a,a67454a,a67457a,a67458a,a67459a,a67463a,a67464a,a67467a,a67470a,a67471a,a67472a,a67476a,a67477a,a67480a,a67483a,a67484a,a67485a,a67489a,a67490a,a67493a,a67496a,a67497a,a67498a,a67502a,a67503a,a67506a,a67509a,a67510a,a67511a,a67515a,a67516a,a67519a,a67522a,a67523a,a67524a,a67528a,a67529a,a67532a,a67535a,a67536a,a67537a,a67541a,a67542a,a67545a,a67548a,a67549a,a67550a,a67554a,a67555a,a67558a,a67561a,a67562a,a67563a,a67567a,a67568a,a67571a,a67574a,a67575a,a67576a,a67580a,a67581a,a67584a,a67587a,a67588a,a67589a,a67593a,a67594a,a67597a,a67600a,a67601a,a67602a,a67606a,a67607a,a67610a,a67613a,a67614a,a67615a,a67619a,a67620a,a67623a,a67626a,a67627a,a67628a,a67632a,a67633a,a67636a,a67639a,a67640a,a67641a,a67645a,a67646a,a67649a,a67652a,a67653a,a67654a,a67658a,a67659a,a67662a,a67665a,a67666a,a67667a,a67671a,a67672a,a67675a,a67678a,a67679a,a67680a,a67684a,a67685a,a67688a,a67691a,a67692a,a67693a,a67697a,a67698a,a67701a,a67704a,a67705a,a67706a,a67710a,a67711a,a67714a,a67717a,a67718a,a67719a,a67723a,a67724a,a67727a,a67730a,a67731a,a67732a,a67736a,a67737a,a67740a,a67743a,a67744a,a67745a,a67749a,a67750a,a67753a,a67756a,a67757a,a67758a,a67762a,a67763a,a67766a,a67769a,a67770a,a67771a,a67775a,a67776a,a67779a,a67782a,a67783a,a67784a,a67788a,a67789a,a67792a,a67795a,a67796a,a67797a,a67801a,a67802a,a67805a,a67808a,a67809a,a67810a,a67814a,a67815a,a67818a,a67821a,a67822a,a67823a,a67827a,a67828a,a67831a,a67834a,a67835a,a67836a,a67840a,a67841a,a67844a,a67847a,a67848a,a67849a,a67853a,a67854a,a67857a,a67860a,a67861a,a67862a,a67866a,a67867a,a67870a,a67873a,a67874a,a67875a,a67879a,a67880a,a67883a,a67886a,a67887a,a67888a,a67892a,a67893a,a67896a,a67899a,a67900a,a67901a,a67905a,a67906a,a67909a,a67912a,a67913a,a67914a,a67918a,a67919a,a67922a,a67925a,a67926a,a67927a,a67931a,a67932a,a67935a,a67938a,a67939a,a67940a,a67944a,a67945a,a67948a,a67951a,a67952a,a67953a,a67957a,a67958a,a67961a,a67964a,a67965a,a67966a,a67970a,a67971a,a67974a,a67977a,a67978a,a67979a,a67983a,a67984a,a67987a,a67990a,a67991a,a67992a,a67996a,a67997a,a68000a,a68003a,a68004a,a68005a,a68009a,a68010a,a68013a,a68016a,a68017a,a68018a,a68022a,a68023a,a68026a,a68029a,a68030a,a68031a,a68035a,a68036a,a68039a,a68042a,a68043a,a68044a,a68048a,a68049a,a68052a,a68055a,a68056a,a68057a,a68061a,a68062a,a68065a,a68068a,a68069a,a68070a,a68074a,a68075a,a68078a,a68081a,a68082a,a68083a,a68087a,a68088a,a68091a,a68094a,a68095a,a68096a,a68100a,a68101a,a68104a,a68107a,a68108a,a68109a,a68113a,a68114a,a68117a,a68120a,a68121a,a68122a,a68126a,a68127a,a68130a,a68133a,a68134a,a68135a,a68139a,a68140a,a68143a,a68146a,a68147a,a68148a,a68152a,a68153a,a68156a,a68159a,a68160a,a68161a,a68165a,a68166a,a68169a,a68172a,a68173a,a68174a,a68178a,a68179a,a68182a,a68185a,a68186a,a68187a,a68191a,a68192a,a68195a,a68198a,a68199a,a68200a,a68204a,a68205a,a68208a,a68211a,a68212a,a68213a,a68217a,a68218a,a68221a,a68224a,a68225a,a68226a,a68230a,a68231a,a68234a,a68237a,a68238a,a68239a,a68243a,a68244a,a68247a,a68250a,a68251a,a68252a,a68256a,a68257a,a68260a,a68263a,a68264a,a68265a,a68269a,a68270a,a68273a,a68276a,a68277a,a68278a,a68282a,a68283a,a68286a,a68289a,a68290a,a68291a,a68295a,a68296a,a68299a,a68302a,a68303a,a68304a,a68308a,a68309a,a68312a,a68315a,a68316a,a68317a,a68321a,a68322a,a68325a,a68328a,a68329a,a68330a,a68334a,a68335a,a68338a,a68341a,a68342a,a68343a,a68347a,a68348a,a68351a,a68354a,a68355a,a68356a,a68360a,a68361a,a68364a,a68367a,a68368a,a68369a,a68373a,a68374a,a68377a,a68380a,a68381a,a68382a,a68386a,a68387a,a68390a,a68393a,a68394a,a68395a,a68399a,a68400a,a68403a,a68406a,a68407a,a68408a,a68412a,a68413a,a68416a,a68419a,a68420a,a68421a,a68425a,a68426a,a68429a,a68432a,a68433a,a68434a,a68438a,a68439a,a68442a,a68445a,a68446a,a68447a,a68451a,a68452a,a68455a,a68458a,a68459a,a68460a,a68464a,a68465a,a68468a,a68471a,a68472a,a68473a,a68477a,a68478a,a68481a,a68484a,a68485a,a68486a,a68490a,a68491a,a68494a,a68497a,a68498a,a68499a,a68503a,a68504a,a68507a,a68510a,a68511a,a68512a,a68516a,a68517a,a68520a,a68523a,a68524a,a68525a,a68529a,a68530a,a68533a,a68536a,a68537a,a68538a,a68542a,a68543a,a68546a,a68549a,a68550a,a68551a,a68555a,a68556a,a68559a,a68562a,a68563a,a68564a,a68568a,a68569a,a68572a,a68575a,a68576a,a68577a,a68581a,a68582a,a68585a,a68588a,a68589a,a68590a,a68594a,a68595a,a68598a,a68601a,a68602a,a68603a,a68607a,a68608a,a68611a,a68614a,a68615a,a68616a,a68620a,a68621a,a68624a,a68627a,a68628a,a68629a,a68633a,a68634a,a68637a,a68640a,a68641a,a68642a,a68646a,a68647a,a68650a,a68653a,a68654a,a68655a,a68659a,a68660a,a68663a,a68666a,a68667a,a68668a,a68672a,a68673a,a68676a,a68679a,a68680a,a68681a,a68685a,a68686a,a68689a,a68692a,a68693a,a68694a,a68698a,a68699a,a68702a,a68705a,a68706a,a68707a,a68711a,a68712a,a68715a,a68718a,a68719a,a68720a,a68724a,a68725a,a68728a,a68731a,a68732a,a68733a,a68737a,a68738a,a68741a,a68744a,a68745a,a68746a,a68750a,a68751a,a68754a,a68757a,a68758a,a68759a,a68763a,a68764a,a68767a,a68770a,a68771a,a68772a,a68776a,a68777a,a68780a,a68783a,a68784a,a68785a,a68789a,a68790a,a68793a,a68796a,a68797a,a68798a,a68802a,a68803a,a68806a,a68809a,a68810a,a68811a,a68815a,a68816a,a68819a,a68822a,a68823a,a68824a,a68828a,a68829a,a68832a,a68835a,a68836a,a68837a,a68841a,a68842a,a68845a,a68848a,a68849a,a68850a,a68854a,a68855a,a68858a,a68861a,a68862a,a68863a,a68867a,a68868a,a68871a,a68874a,a68875a,a68876a,a68880a,a68881a,a68884a,a68887a,a68888a,a68889a,a68893a,a68894a,a68897a,a68900a,a68901a,a68902a,a68906a,a68907a,a68910a,a68913a,a68914a,a68915a,a68919a,a68920a,a68923a,a68926a,a68927a,a68928a,a68932a,a68933a,a68936a,a68939a,a68940a,a68941a,a68945a,a68946a,a68949a,a68952a,a68953a,a68954a,a68958a,a68959a,a68962a,a68965a,a68966a,a68967a,a68971a,a68972a,a68975a,a68978a,a68979a,a68980a,a68984a,a68985a,a68988a,a68991a,a68992a,a68993a,a68997a,a68998a,a69001a,a69004a,a69005a,a69006a,a69010a,a69011a,a69014a,a69017a,a69018a,a69019a,a69023a,a69024a,a69027a,a69030a,a69031a,a69032a,a69036a,a69037a,a69040a,a69043a,a69044a,a69045a,a69049a,a69050a,a69053a,a69056a,a69057a,a69058a,a69062a,a69063a,a69066a,a69069a,a69070a,a69071a,a69075a,a69076a,a69079a,a69082a,a69083a,a69084a,a69088a,a69089a,a69092a,a69095a,a69096a,a69097a,a69101a,a69102a,a69105a,a69108a,a69109a,a69110a,a69114a,a69115a,a69118a,a69121a,a69122a,a69123a,a69127a,a69128a,a69131a,a69134a,a69135a,a69136a,a69140a,a69141a,a69144a,a69147a,a69148a,a69149a,a69153a,a69154a,a69157a,a69160a,a69161a,a69162a,a69166a,a69167a,a69170a,a69173a,a69174a,a69175a,a69179a,a69180a,a69183a,a69186a,a69187a,a69188a,a69192a,a69193a,a69196a,a69199a,a69200a,a69201a,a69205a,a69206a,a69209a,a69212a,a69213a,a69214a,a69218a,a69219a,a69222a,a69225a,a69226a,a69227a,a69231a,a69232a,a69235a,a69238a,a69239a,a69240a,a69244a,a69245a,a69248a,a69251a,a69252a,a69253a,a69257a,a69258a,a69261a,a69264a,a69265a,a69266a,a69270a,a69271a,a69274a,a69277a,a69278a,a69279a,a69283a,a69284a,a69287a,a69290a,a69291a,a69292a,a69296a,a69297a,a69300a,a69303a,a69304a,a69305a,a69309a,a69310a,a69313a,a69316a,a69317a,a69318a,a69322a,a69323a,a69326a,a69329a,a69330a,a69331a,a69335a,a69336a,a69339a,a69342a,a69343a,a69344a,a69348a,a69349a,a69352a,a69355a,a69356a,a69357a,a69361a,a69362a,a69365a,a69368a,a69369a,a69370a,a69374a,a69375a,a69378a,a69381a,a69382a,a69383a,a69387a,a69388a,a69391a,a69394a,a69395a,a69396a,a69400a,a69401a,a69404a,a69407a,a69408a,a69409a,a69413a,a69414a,a69417a,a69420a,a69421a,a69422a,a69426a,a69427a,a69430a,a69433a,a69434a,a69435a,a69439a,a69440a,a69443a,a69446a,a69447a,a69448a,a69452a,a69453a,a69456a,a69459a,a69460a,a69461a,a69465a,a69466a,a69469a,a69472a,a69473a,a69474a,a69478a,a69479a,a69482a,a69485a,a69486a,a69487a,a69491a,a69492a,a69495a,a69498a,a69499a,a69500a,a69504a,a69505a,a69508a,a69511a,a69512a,a69513a,a69517a,a69518a,a69521a,a69524a,a69525a,a69526a,a69530a,a69531a,a69534a,a69537a,a69538a,a69539a,a69543a,a69544a,a69547a,a69550a,a69551a,a69552a,a69556a,a69557a,a69560a,a69563a,a69564a,a69565a,a69569a,a69570a,a69573a,a69576a,a69577a,a69578a,a69582a,a69583a,a69586a,a69589a,a69590a,a69591a,a69595a,a69596a,a69599a,a69602a,a69603a,a69604a,a69608a,a69609a,a69612a,a69615a,a69616a,a69617a,a69621a,a69622a,a69625a,a69628a,a69629a,a69630a,a69634a,a69635a,a69638a,a69641a,a69642a,a69643a,a69647a,a69648a,a69651a,a69654a,a69655a,a69656a,a69660a,a69661a,a69664a,a69667a,a69668a,a69669a,a69673a,a69674a,a69677a,a69680a,a69681a,a69682a,a69686a,a69687a,a69690a,a69693a,a69694a,a69695a,a69699a,a69700a,a69703a,a69706a,a69707a,a69708a,a69712a,a69713a,a69716a,a69719a,a69720a,a69721a,a69725a,a69726a,a69729a,a69732a,a69733a,a69734a,a69738a,a69739a,a69742a,a69745a,a69746a,a69747a,a69751a,a69752a,a69755a,a69758a,a69759a,a69760a,a69764a,a69765a,a69768a,a69771a,a69772a,a69773a,a69777a,a69778a,a69781a,a69784a,a69785a,a69786a,a69790a,a69791a,a69794a,a69797a,a69798a,a69799a,a69803a,a69804a,a69807a,a69810a,a69811a,a69812a,a69816a,a69817a,a69820a,a69823a,a69824a,a69825a,a69829a,a69830a,a69833a,a69836a,a69837a,a69838a,a69842a,a69843a,a69846a,a69849a,a69850a,a69851a,a69855a,a69856a,a69859a,a69862a,a69863a,a69864a,a69868a,a69869a,a69872a,a69875a,a69876a,a69877a,a69881a,a69882a,a69885a,a69888a,a69889a,a69890a,a69894a,a69895a,a69898a,a69901a,a69902a,a69903a,a69907a,a69908a,a69911a,a69914a,a69915a,a69916a,a69920a,a69921a,a69924a,a69927a,a69928a,a69929a,a69933a,a69934a,a69937a,a69940a,a69941a,a69942a,a69946a,a69947a,a69950a,a69953a,a69954a,a69955a,a69959a,a69960a,a69963a,a69966a,a69967a,a69968a,a69972a,a69973a,a69976a,a69979a,a69980a,a69981a,a69985a,a69986a,a69989a,a69992a,a69993a,a69994a,a69998a,a69999a,a70002a,a70005a,a70006a,a70007a,a70011a,a70012a,a70015a,a70018a,a70019a,a70020a,a70024a,a70025a,a70028a,a70031a,a70032a,a70033a,a70037a,a70038a,a70041a,a70044a,a70045a,a70046a,a70050a,a70051a,a70054a,a70057a,a70058a,a70059a,a70063a,a70064a,a70067a,a70070a,a70071a,a70072a,a70076a,a70077a,a70080a,a70083a,a70084a,a70085a,a70089a,a70090a,a70093a,a70096a,a70097a,a70098a,a70102a,a70103a,a70106a,a70109a,a70110a,a70111a,a70115a,a70116a,a70119a,a70122a,a70123a,a70124a,a70128a,a70129a,a70132a,a70135a,a70136a,a70137a,a70141a,a70142a,a70145a,a70148a,a70149a,a70150a,a70154a,a70155a,a70158a,a70161a,a70162a,a70163a,a70167a,a70168a,a70171a,a70174a,a70175a,a70176a,a70180a,a70181a,a70184a,a70187a,a70188a,a70189a,a70193a,a70194a,a70197a,a70200a,a70201a,a70202a,a70206a,a70207a,a70210a,a70213a,a70214a,a70215a,a70219a,a70220a,a70223a,a70226a,a70227a,a70228a,a70232a,a70233a,a70236a,a70239a,a70240a,a70241a,a70245a,a70246a,a70249a,a70252a,a70253a,a70254a,a70258a,a70259a,a70262a,a70265a,a70266a,a70267a,a70271a,a70272a,a70275a,a70278a,a70279a,a70280a,a70284a,a70285a,a70288a,a70291a,a70292a,a70293a,a70297a,a70298a,a70301a,a70304a,a70305a,a70306a,a70310a,a70311a,a70314a,a70317a,a70318a,a70319a,a70323a,a70324a,a70327a,a70330a,a70331a,a70332a,a70336a,a70337a,a70340a,a70343a,a70344a,a70345a,a70349a,a70350a,a70353a,a70356a,a70357a,a70358a,a70362a,a70363a,a70366a,a70369a,a70370a,a70371a,a70375a,a70376a,a70379a,a70382a,a70383a,a70384a,a70388a,a70389a,a70392a,a70395a,a70396a,a70397a,a70401a,a70402a,a70405a,a70408a,a70409a,a70410a,a70414a,a70415a,a70418a,a70421a,a70422a,a70423a,a70427a,a70428a,a70431a,a70434a,a70435a,a70436a,a70440a,a70441a,a70444a,a70447a,a70448a,a70449a,a70453a,a70454a,a70457a,a70460a,a70461a,a70462a,a70466a,a70467a,a70470a,a70473a,a70474a,a70475a,a70479a,a70480a,a70483a,a70486a,a70487a,a70488a,a70492a,a70493a,a70496a,a70499a,a70500a,a70501a,a70505a,a70506a,a70509a,a70512a,a70513a,a70514a,a70518a,a70519a,a70522a,a70525a,a70526a,a70527a,a70531a,a70532a,a70535a,a70538a,a70539a,a70540a,a70544a,a70545a,a70548a,a70551a,a70552a,a70553a,a70557a,a70558a,a70561a,a70564a,a70565a,a70566a,a70570a,a70571a,a70574a,a70577a,a70578a,a70579a,a70583a,a70584a,a70587a,a70590a,a70591a,a70592a,a70596a,a70597a,a70600a,a70603a,a70604a,a70605a,a70609a,a70610a,a70613a,a70616a,a70617a,a70618a,a70622a,a70623a,a70626a,a70629a,a70630a,a70631a,a70635a,a70636a,a70639a,a70642a,a70643a,a70644a,a70648a,a70649a,a70652a,a70655a,a70656a,a70657a,a70661a,a70662a,a70665a,a70668a,a70669a,a70670a,a70674a,a70675a,a70678a,a70681a,a70682a,a70683a,a70687a,a70688a,a70691a,a70694a,a70695a,a70696a,a70700a,a70701a,a70704a,a70707a,a70708a,a70709a,a70713a,a70714a,a70717a,a70720a,a70721a,a70722a,a70726a,a70727a,a70730a,a70733a,a70734a,a70735a,a70739a,a70740a,a70743a,a70746a,a70747a,a70748a,a70752a,a70753a,a70756a,a70759a,a70760a,a70761a,a70765a,a70766a,a70769a,a70772a,a70773a,a70774a,a70778a,a70779a,a70782a,a70785a,a70786a,a70787a,a70791a,a70792a,a70795a,a70798a,a70799a,a70800a,a70804a,a70805a,a70808a,a70811a,a70812a,a70813a,a70817a,a70818a,a70821a,a70824a,a70825a,a70826a,a70830a,a70831a,a70834a,a70837a,a70838a,a70839a,a70843a,a70844a,a70847a,a70850a,a70851a,a70852a,a70856a,a70857a,a70860a,a70863a,a70864a,a70865a,a70869a,a70870a,a70873a,a70876a,a70877a,a70878a,a70882a,a70883a,a70886a,a70889a,a70890a,a70891a,a70895a,a70896a,a70899a,a70902a,a70903a,a70904a,a70908a,a70909a,a70912a,a70915a,a70916a,a70917a,a70921a,a70922a,a70925a,a70928a,a70929a,a70930a,a70934a,a70935a,a70938a,a70941a,a70942a,a70943a,a70947a,a70948a,a70951a,a70954a,a70955a,a70956a,a70960a,a70961a,a70964a,a70967a,a70968a,a70969a,a70973a,a70974a,a70977a,a70980a,a70981a,a70982a,a70986a,a70987a,a70990a,a70993a,a70994a,a70995a,a70999a,a71000a,a71003a,a71006a,a71007a,a71008a,a71012a,a71013a,a71016a,a71019a,a71020a,a71021a,a71025a,a71026a,a71029a,a71032a,a71033a,a71034a,a71038a,a71039a,a71042a,a71045a,a71046a,a71047a,a71051a,a71052a,a71055a,a71058a,a71059a,a71060a,a71064a,a71065a,a71068a,a71071a,a71072a,a71073a,a71077a,a71078a,a71081a,a71084a,a71085a,a71086a,a71090a,a71091a,a71094a,a71097a,a71098a,a71099a,a71103a,a71104a,a71107a,a71110a,a71111a,a71112a,a71116a,a71117a,a71120a,a71123a,a71124a,a71125a,a71129a,a71130a,a71133a,a71136a,a71137a,a71138a,a71142a,a71143a,a71146a,a71149a,a71150a,a71151a,a71155a,a71156a,a71159a,a71162a,a71163a,a71164a,a71168a,a71169a,a71172a,a71175a,a71176a,a71177a,a71181a,a71182a,a71185a,a71188a,a71189a,a71190a,a71194a,a71195a,a71198a,a71201a,a71202a,a71203a,a71207a,a71208a,a71211a,a71214a,a71215a,a71216a,a71220a,a71221a,a71224a,a71227a,a71228a,a71229a,a71233a,a71234a,a71237a,a71240a,a71241a,a71242a,a71246a,a71247a,a71250a,a71253a,a71254a,a71255a,a71259a,a71260a,a71263a,a71266a,a71267a,a71268a,a71272a,a71273a,a71276a,a71279a,a71280a,a71281a,a71285a,a71286a,a71289a,a71292a,a71293a,a71294a,a71298a,a71299a,a71302a,a71305a,a71306a,a71307a,a71311a,a71312a,a71315a,a71318a,a71319a,a71320a,a71324a,a71325a,a71328a,a71331a,a71332a,a71333a,a71337a,a71338a,a71341a,a71344a,a71345a,a71346a,a71350a,a71351a,a71354a,a71357a,a71358a,a71359a,a71363a,a71364a,a71367a,a71370a,a71371a,a71372a,a71376a,a71377a,a71380a,a71383a,a71384a,a71385a,a71389a,a71390a,a71393a,a71396a,a71397a,a71398a,a71402a,a71403a,a71406a,a71409a,a71410a,a71411a,a71415a,a71416a,a71419a,a71422a,a71423a,a71424a,a71428a,a71429a,a71432a,a71435a,a71436a,a71437a,a71441a,a71442a,a71445a,a71448a,a71449a,a71450a,a71454a,a71455a,a71458a,a71461a,a71462a,a71463a,a71467a,a71468a,a71471a,a71474a,a71475a,a71476a,a71480a,a71481a,a71484a,a71487a,a71488a,a71489a,a71493a,a71494a,a71497a,a71500a,a71501a,a71502a,a71506a,a71507a,a71510a,a71513a,a71514a,a71515a,a71519a,a71520a,a71523a,a71526a,a71527a,a71528a,a71532a,a71533a,a71536a,a71539a,a71540a,a71541a,a71545a,a71546a,a71549a,a71552a,a71553a,a71554a,a71558a,a71559a,a71562a,a71565a,a71566a,a71567a,a71571a,a71572a,a71575a,a71578a,a71579a,a71580a,a71584a,a71585a,a71588a,a71591a,a71592a,a71593a,a71597a,a71598a,a71601a,a71604a,a71605a,a71606a,a71610a,a71611a,a71614a,a71617a,a71618a,a71619a,a71623a,a71624a,a71627a,a71630a,a71631a,a71632a,a71636a,a71637a,a71640a,a71643a,a71644a,a71645a,a71649a,a71650a,a71653a,a71656a,a71657a,a71658a,a71662a,a71663a,a71666a,a71669a,a71670a,a71671a,a71675a,a71676a,a71679a,a71682a,a71683a,a71684a,a71688a,a71689a,a71692a,a71695a,a71696a,a71697a,a71701a,a71702a,a71705a,a71708a,a71709a,a71710a,a71714a,a71715a,a71718a,a71721a,a71722a,a71723a,a71727a,a71728a,a71731a,a71734a,a71735a,a71736a,a71740a,a71741a,a71744a,a71747a,a71748a,a71749a,a71753a,a71754a,a71757a,a71760a,a71761a,a71762a,a71766a,a71767a,a71770a,a71773a,a71774a,a71775a,a71779a,a71780a,a71783a,a71786a,a71787a,a71788a,a71792a,a71793a,a71796a,a71799a,a71800a,a71801a,a71805a,a71806a,a71809a,a71812a,a71813a,a71814a,a71818a,a71819a,a71822a,a71825a,a71826a,a71827a,a71831a,a71832a,a71835a,a71838a,a71839a,a71840a,a71844a,a71845a,a71848a,a71851a,a71852a,a71853a,a71857a,a71858a,a71861a,a71864a,a71865a,a71866a,a71870a,a71871a,a71874a,a71877a,a71878a,a71879a,a71883a,a71884a,a71887a,a71890a,a71891a,a71892a,a71896a,a71897a,a71900a,a71903a,a71904a,a71905a,a71909a,a71910a,a71913a,a71916a,a71917a,a71918a,a71922a,a71923a,a71926a,a71929a,a71930a,a71931a,a71935a,a71936a,a71939a,a71942a,a71943a,a71944a,a71948a,a71949a,a71952a,a71955a,a71956a,a71957a,a71961a,a71962a,a71965a,a71968a,a71969a,a71970a,a71974a,a71975a,a71978a,a71981a,a71982a,a71983a,a71987a,a71988a,a71991a,a71994a,a71995a,a71996a,a72000a,a72001a,a72004a,a72007a,a72008a,a72009a,a72013a,a72014a,a72017a,a72020a,a72021a,a72022a,a72026a,a72027a,a72030a,a72033a,a72034a,a72035a,a72039a,a72040a,a72043a,a72046a,a72047a,a72048a,a72052a,a72053a,a72056a,a72059a,a72060a,a72061a,a72065a,a72066a,a72069a,a72072a,a72073a,a72074a,a72078a,a72079a,a72082a,a72085a,a72086a,a72087a,a72091a,a72092a,a72095a,a72098a,a72099a,a72100a,a72104a,a72105a,a72108a,a72111a,a72112a,a72113a,a72117a,a72118a,a72121a,a72124a,a72125a,a72126a,a72130a,a72131a,a72134a,a72137a,a72138a,a72139a,a72143a,a72144a,a72147a,a72150a,a72151a,a72152a,a72156a,a72157a,a72160a,a72163a,a72164a,a72165a,a72169a,a72170a,a72173a,a72176a,a72177a,a72178a,a72182a,a72183a,a72186a,a72189a,a72190a,a72191a,a72195a,a72196a,a72199a,a72202a,a72203a,a72204a,a72208a,a72209a,a72212a,a72215a,a72216a,a72217a,a72221a,a72222a,a72225a,a72228a,a72229a,a72230a,a72234a,a72235a,a72238a,a72241a,a72242a,a72243a,a72247a,a72248a,a72251a,a72254a,a72255a,a72256a,a72260a,a72261a,a72264a,a72267a,a72268a,a72269a,a72273a,a72274a,a72277a,a72280a,a72281a,a72282a,a72286a,a72287a,a72290a,a72293a,a72294a,a72295a,a72299a,a72300a,a72303a,a72306a,a72307a,a72308a,a72312a,a72313a,a72316a,a72319a,a72320a,a72321a,a72325a,a72326a,a72329a,a72332a,a72333a,a72334a,a72338a,a72339a,a72342a,a72345a,a72346a,a72347a,a72351a,a72352a,a72355a,a72358a,a72359a,a72360a,a72364a,a72365a,a72368a,a72371a,a72372a,a72373a,a72377a,a72378a,a72381a,a72384a,a72385a,a72386a,a72390a,a72391a,a72394a,a72397a,a72398a,a72399a,a72403a,a72404a,a72407a,a72410a,a72411a,a72412a,a72416a,a72417a,a72420a,a72423a,a72424a,a72425a,a72429a,a72430a,a72433a,a72436a,a72437a,a72438a,a72442a,a72443a,a72446a,a72449a,a72450a,a72451a,a72455a,a72456a,a72459a,a72462a,a72463a,a72464a,a72468a,a72469a,a72472a,a72475a,a72476a,a72477a,a72481a,a72482a,a72485a,a72488a,a72489a,a72490a,a72494a,a72495a,a72498a,a72501a,a72502a,a72503a,a72507a,a72508a,a72511a,a72514a,a72515a,a72516a,a72520a,a72521a,a72524a,a72527a,a72528a,a72529a,a72533a,a72534a,a72537a,a72540a,a72541a,a72542a,a72546a,a72547a,a72550a,a72553a,a72554a,a72555a,a72559a,a72560a,a72563a,a72566a,a72567a,a72568a,a72572a,a72573a,a72576a,a72579a,a72580a,a72581a,a72585a,a72586a,a72589a,a72592a,a72593a,a72594a,a72598a,a72599a,a72602a,a72605a,a72606a,a72607a,a72611a,a72612a,a72615a,a72618a,a72619a,a72620a,a72624a,a72625a,a72628a,a72631a,a72632a,a72633a,a72637a,a72638a,a72641a,a72644a,a72645a,a72646a,a72650a,a72651a,a72654a,a72657a,a72658a,a72659a,a72663a,a72664a,a72667a,a72670a,a72671a,a72672a,a72676a,a72677a,a72680a,a72683a,a72684a,a72685a,a72689a,a72690a,a72693a,a72696a,a72697a,a72698a,a72702a,a72703a,a72706a,a72709a,a72710a,a72711a,a72715a,a72716a,a72719a,a72722a,a72723a,a72724a,a72728a,a72729a,a72732a,a72735a,a72736a,a72737a,a72741a,a72742a,a72745a,a72748a,a72749a,a72750a,a72754a,a72755a,a72758a,a72761a,a72762a,a72763a,a72767a,a72768a,a72771a,a72774a,a72775a,a72776a,a72780a,a72781a,a72784a,a72787a,a72788a,a72789a,a72793a,a72794a,a72797a,a72800a,a72801a,a72802a,a72806a,a72807a,a72810a,a72813a,a72814a,a72815a,a72819a,a72820a,a72823a,a72826a,a72827a,a72828a,a72832a,a72833a,a72836a,a72839a,a72840a,a72841a,a72845a,a72846a,a72849a,a72852a,a72853a,a72854a,a72858a,a72859a,a72862a,a72865a,a72866a,a72867a,a72871a,a72872a,a72875a,a72878a,a72879a,a72880a,a72884a,a72885a,a72888a,a72891a,a72892a,a72893a,a72897a,a72898a,a72901a,a72904a,a72905a,a72906a,a72910a,a72911a,a72914a,a72917a,a72918a,a72919a,a72923a,a72924a,a72927a,a72930a,a72931a,a72932a,a72936a,a72937a,a72940a,a72943a,a72944a,a72945a,a72949a,a72950a,a72953a,a72956a,a72957a,a72958a,a72962a,a72963a,a72966a,a72969a,a72970a,a72971a,a72975a,a72976a,a72979a,a72982a,a72983a,a72984a,a72988a,a72989a,a72992a,a72995a,a72996a,a72997a,a73001a,a73002a,a73005a,a73008a,a73009a,a73010a,a73014a,a73015a,a73018a,a73021a,a73022a,a73023a,a73027a,a73028a,a73031a,a73034a,a73035a,a73036a,a73040a,a73041a,a73044a,a73047a,a73048a,a73049a,a73053a,a73054a,a73057a,a73060a,a73061a,a73062a,a73066a,a73067a,a73070a,a73073a,a73074a,a73075a,a73079a,a73080a,a73083a,a73086a,a73087a,a73088a,a73092a,a73093a,a73096a,a73099a,a73100a,a73101a,a73105a,a73106a,a73109a,a73112a,a73113a,a73114a,a73118a,a73119a,a73122a,a73125a,a73126a,a73127a,a73131a,a73132a,a73135a,a73138a,a73139a,a73140a,a73144a,a73145a,a73148a,a73151a,a73152a,a73153a,a73157a,a73158a,a73161a,a73164a,a73165a,a73166a,a73170a,a73171a,a73174a,a73177a,a73178a,a73179a,a73183a,a73184a,a73187a,a73190a,a73191a,a73192a,a73196a,a73197a,a73200a,a73203a,a73204a,a73205a,a73209a,a73210a,a73213a,a73216a,a73217a,a73218a,a73222a,a73223a,a73226a,a73229a,a73230a,a73231a,a73235a,a73236a,a73239a,a73242a,a73243a,a73244a,a73248a,a73249a,a73252a,a73255a,a73256a,a73257a,a73261a,a73262a,a73265a,a73268a,a73269a,a73270a,a73274a,a73275a,a73278a,a73281a,a73282a,a73283a,a73287a,a73288a,a73291a,a73294a,a73295a,a73296a,a73300a,a73301a,a73304a,a73307a,a73308a,a73309a,a73313a,a73314a,a73317a,a73320a,a73321a,a73322a,a73326a,a73327a,a73330a,a73333a,a73334a,a73335a,a73339a,a73340a,a73343a,a73346a,a73347a,a73348a,a73352a,a73353a,a73356a,a73359a,a73360a,a73361a,a73365a,a73366a,a73369a,a73372a,a73373a,a73374a,a73378a,a73379a,a73382a,a73385a,a73386a,a73387a,a73391a,a73392a,a73395a,a73398a,a73399a,a73400a,a73404a,a73405a,a73408a,a73411a,a73412a,a73413a,a73417a,a73418a,a73421a,a73424a,a73425a,a73426a,a73430a,a73431a,a73434a,a73437a,a73438a,a73439a,a73443a,a73444a,a73447a,a73450a,a73451a,a73452a,a73456a,a73457a,a73460a,a73463a,a73464a,a73465a,a73469a,a73470a,a73473a,a73476a,a73477a,a73478a,a73482a,a73483a,a73486a,a73489a,a73490a,a73491a,a73495a,a73496a,a73499a,a73502a,a73503a,a73504a,a73508a,a73509a,a73512a,a73515a,a73516a,a73517a,a73521a,a73522a,a73525a,a73528a,a73529a,a73530a,a73534a,a73535a,a73538a,a73541a,a73542a,a73543a,a73547a,a73548a,a73551a,a73554a,a73555a,a73556a,a73560a,a73561a,a73564a,a73567a,a73568a,a73569a,a73573a,a73574a,a73577a,a73580a,a73581a,a73582a,a73586a,a73587a,a73590a,a73593a,a73594a,a73595a,a73599a,a73600a,a73603a,a73606a,a73607a,a73608a,a73612a,a73613a,a73616a,a73619a,a73620a,a73621a,a73625a,a73626a,a73629a,a73632a,a73633a,a73634a,a73638a,a73639a,a73642a,a73645a,a73646a,a73647a,a73651a,a73652a,a73655a,a73658a,a73659a,a73660a,a73664a,a73665a,a73668a,a73671a,a73672a,a73673a,a73677a,a73678a,a73681a,a73684a,a73685a,a73686a,a73690a,a73691a,a73694a,a73697a,a73698a,a73699a,a73703a,a73704a,a73707a,a73710a,a73711a,a73712a,a73716a,a73717a,a73720a,a73723a,a73724a,a73725a,a73729a,a73730a,a73733a,a73736a,a73737a,a73738a,a73742a,a73743a,a73746a,a73749a,a73750a,a73751a,a73755a,a73756a,a73759a,a73762a,a73763a,a73764a,a73768a,a73769a,a73772a,a73775a,a73776a,a73777a,a73781a,a73782a,a73785a,a73788a,a73789a,a73790a,a73794a,a73795a,a73798a,a73801a,a73802a,a73803a,a73807a,a73808a,a73811a,a73814a,a73815a,a73816a,a73820a,a73821a,a73824a,a73827a,a73828a,a73829a,a73833a,a73834a,a73837a,a73840a,a73841a,a73842a,a73846a,a73847a,a73850a,a73853a,a73854a,a73855a,a73859a,a73860a,a73863a,a73866a,a73867a,a73868a,a73872a,a73873a,a73876a,a73879a,a73880a,a73881a,a73885a,a73886a,a73889a,a73892a,a73893a,a73894a,a73898a,a73899a,a73902a,a73905a,a73906a,a73907a,a73911a,a73912a,a73915a,a73918a,a73919a,a73920a,a73924a,a73925a,a73928a,a73931a,a73932a,a73933a,a73937a,a73938a,a73941a,a73944a,a73945a,a73946a,a73950a,a73951a,a73954a,a73957a,a73958a,a73959a,a73963a,a73964a,a73967a,a73970a,a73971a,a73972a,a73976a,a73977a,a73980a,a73983a,a73984a,a73985a,a73989a,a73990a,a73993a,a73996a,a73997a,a73998a,a74002a,a74003a,a74006a,a74009a,a74010a,a74011a,a74015a,a74016a,a74019a,a74022a,a74023a,a74024a,a74028a,a74029a,a74032a,a74035a,a74036a,a74037a,a74041a,a74042a,a74045a,a74048a,a74049a,a74050a,a74054a,a74055a,a74058a,a74061a,a74062a,a74063a,a74067a,a74068a,a74071a,a74074a,a74075a,a74076a,a74080a,a74081a,a74084a,a74087a,a74088a,a74089a,a74093a,a74094a,a74097a,a74100a,a74101a,a74102a,a74106a,a74107a,a74110a,a74113a,a74114a,a74115a,a74119a,a74120a,a74123a,a74126a,a74127a,a74128a,a74132a,a74133a,a74136a,a74139a,a74140a,a74141a,a74145a,a74146a,a74149a,a74152a,a74153a,a74154a,a74158a,a74159a,a74162a,a74165a,a74166a,a74167a,a74171a,a74172a,a74175a,a74178a,a74179a,a74180a,a74184a,a74185a,a74188a,a74191a,a74192a,a74193a,a74197a,a74198a,a74201a,a74204a,a74205a,a74206a,a74210a,a74211a,a74214a,a74217a,a74218a,a74219a,a74223a,a74224a,a74227a,a74230a,a74231a,a74232a,a74236a,a74237a,a74240a,a74243a,a74244a,a74245a,a74249a,a74250a,a74253a,a74256a,a74257a,a74258a,a74262a,a74263a,a74266a,a74269a,a74270a,a74271a,a74275a,a74276a,a74279a,a74282a,a74283a,a74284a,a74288a,a74289a,a74292a,a74295a,a74296a,a74297a,a74301a,a74302a,a74305a,a74308a,a74309a,a74310a,a74314a,a74315a,a74318a,a74321a,a74322a,a74323a,a74327a,a74328a,a74331a,a74334a,a74335a,a74336a,a74340a,a74341a,a74344a,a74347a,a74348a,a74349a,a74353a,a74354a,a74357a,a74360a,a74361a,a74362a,a74366a,a74367a,a74370a,a74373a,a74374a,a74375a,a74379a,a74380a,a74383a,a74386a,a74387a,a74388a,a74392a,a74393a,a74396a,a74399a,a74400a,a74401a,a74405a,a74406a,a74409a,a74412a,a74413a,a74414a,a74418a,a74419a,a74422a,a74425a,a74426a,a74427a,a74431a,a74432a,a74435a,a74438a,a74439a,a74440a,a74444a,a74445a,a74448a,a74451a,a74452a,a74453a,a74457a,a74458a,a74461a,a74464a,a74465a,a74466a,a74470a,a74471a,a74474a,a74477a,a74478a,a74479a,a74483a,a74484a,a74487a,a74490a,a74491a,a74492a,a74496a,a74497a,a74500a,a74503a,a74504a,a74505a,a74509a,a74510a,a74513a,a74516a,a74517a,a74518a,a74522a,a74523a,a74526a,a74529a,a74530a,a74531a,a74535a,a74536a,a74539a,a74542a,a74543a,a74544a,a74548a,a74549a,a74552a,a74555a,a74556a,a74557a,a74561a,a74562a,a74565a,a74568a,a74569a,a74570a,a74574a,a74575a,a74578a,a74581a,a74582a,a74583a,a74587a,a74588a,a74591a,a74594a,a74595a,a74596a,a74600a,a74601a,a74604a,a74607a,a74608a,a74609a,a74613a,a74614a,a74617a,a74620a,a74621a,a74622a,a74626a,a74627a,a74630a,a74633a,a74634a,a74635a,a74639a,a74640a,a74643a,a74646a,a74647a,a74648a,a74652a,a74653a,a74656a,a74659a,a74660a,a74661a,a74665a,a74666a,a74669a,a74672a,a74673a,a74674a,a74678a,a74679a,a74682a,a74685a,a74686a,a74687a,a74691a,a74692a,a74695a,a74698a,a74699a,a74700a,a74704a,a74705a,a74708a,a74711a,a74712a,a74713a,a74717a,a74718a,a74721a,a74724a,a74725a,a74726a,a74730a,a74731a,a74734a,a74737a,a74738a,a74739a,a74743a,a74744a,a74747a,a74750a,a74751a,a74752a,a74756a,a74757a,a74760a,a74763a,a74764a,a74765a,a74769a,a74770a,a74773a,a74776a,a74777a,a74778a,a74782a,a74783a,a74786a,a74789a,a74790a,a74791a,a74795a,a74796a,a74799a,a74802a,a74803a,a74804a,a74808a,a74809a,a74812a,a74815a,a74816a,a74817a,a74821a,a74822a,a74825a,a74828a,a74829a,a74830a,a74834a,a74835a,a74838a,a74841a,a74842a,a74843a,a74847a,a74848a,a74851a,a74854a,a74855a,a74856a,a74860a,a74861a,a74864a,a74867a,a74868a,a74869a,a74873a,a74874a,a74877a,a74880a,a74881a,a74882a,a74886a,a74887a,a74890a,a74893a,a74894a,a74895a,a74899a,a74900a,a74903a,a74906a,a74907a,a74908a,a74912a,a74913a,a74916a,a74919a,a74920a,a74921a,a74925a,a74926a,a74929a,a74932a,a74933a,a74934a,a74938a,a74939a,a74942a,a74945a,a74946a,a74947a,a74951a,a74952a,a74955a,a74958a,a74959a,a74960a,a74964a,a74965a,a74968a,a74971a,a74972a,a74973a,a74977a,a74978a,a74981a,a74984a,a74985a,a74986a,a74990a,a74991a,a74994a,a74997a,a74998a,a74999a,a75003a,a75004a,a75007a,a75010a,a75011a,a75012a,a75016a,a75017a,a75020a,a75023a,a75024a,a75025a,a75029a,a75030a,a75033a,a75036a,a75037a,a75038a,a75042a,a75043a,a75046a,a75049a,a75050a,a75051a,a75055a,a75056a,a75059a,a75062a,a75063a,a75064a,a75068a,a75069a,a75072a,a75075a,a75076a,a75077a,a75081a,a75082a,a75085a,a75088a,a75089a,a75090a,a75094a,a75095a,a75098a,a75101a,a75102a,a75103a,a75107a,a75108a,a75111a,a75114a,a75115a,a75116a,a75120a,a75121a,a75124a,a75127a,a75128a,a75129a,a75133a,a75134a,a75137a,a75140a,a75141a,a75142a,a75146a,a75147a,a75150a,a75153a,a75154a,a75155a,a75159a,a75160a,a75163a,a75166a,a75167a,a75168a,a75172a,a75173a,a75176a,a75179a,a75180a,a75181a,a75185a,a75186a,a75189a,a75192a,a75193a,a75194a,a75198a,a75199a,a75202a,a75205a,a75206a,a75207a,a75211a,a75212a,a75215a,a75218a,a75219a,a75220a,a75224a,a75225a,a75228a,a75231a,a75232a,a75233a,a75237a,a75238a,a75241a,a75244a,a75245a,a75246a,a75250a,a75251a,a75254a,a75257a,a75258a,a75259a,a75263a,a75264a,a75267a,a75270a,a75271a,a75272a,a75276a,a75277a,a75280a,a75283a,a75284a,a75285a,a75289a,a75290a,a75293a,a75296a,a75297a,a75298a,a75302a,a75303a,a75306a,a75309a,a75310a,a75311a,a75315a,a75316a,a75319a,a75322a,a75323a,a75324a,a75328a,a75329a,a75332a,a75335a,a75336a,a75337a,a75341a,a75342a,a75345a,a75348a,a75349a,a75350a,a75354a,a75355a,a75358a,a75361a,a75362a,a75363a,a75367a,a75368a,a75371a,a75374a,a75375a,a75376a,a75380a,a75381a,a75384a,a75387a,a75388a,a75389a,a75393a,a75394a,a75397a,a75400a,a75401a,a75402a,a75406a,a75407a,a75410a,a75413a,a75414a,a75415a,a75419a,a75420a,a75423a,a75426a,a75427a,a75428a,a75432a,a75433a,a75436a,a75439a,a75440a,a75441a,a75445a,a75446a,a75449a,a75452a,a75453a,a75454a,a75458a,a75459a,a75462a,a75465a,a75466a,a75467a,a75471a,a75472a,a75475a,a75478a,a75479a,a75480a,a75484a,a75485a,a75488a,a75491a,a75492a,a75493a,a75497a,a75498a,a75501a,a75504a,a75505a,a75506a,a75510a,a75511a,a75514a,a75517a,a75518a,a75519a,a75523a,a75524a,a75527a,a75530a,a75531a,a75532a,a75536a,a75537a,a75540a,a75543a,a75544a,a75545a,a75549a,a75550a,a75553a,a75556a,a75557a,a75558a,a75562a,a75563a,a75566a,a75569a,a75570a,a75571a,a75575a,a75576a,a75579a,a75582a,a75583a,a75584a,a75588a,a75589a,a75592a,a75595a,a75596a,a75597a,a75601a,a75602a,a75605a,a75608a,a75609a,a75610a,a75614a,a75615a,a75618a,a75621a,a75622a,a75623a,a75627a,a75628a,a75631a,a75634a,a75635a,a75636a,a75640a,a75641a,a75644a,a75647a,a75648a,a75649a,a75653a,a75654a,a75657a,a75660a,a75661a,a75662a,a75666a,a75667a,a75670a,a75673a,a75674a,a75675a,a75679a,a75680a,a75683a,a75686a,a75687a,a75688a,a75692a,a75693a,a75696a,a75699a,a75700a,a75701a,a75705a,a75706a,a75709a,a75712a,a75713a,a75714a,a75718a,a75719a,a75722a,a75725a,a75726a,a75727a,a75731a,a75732a,a75735a,a75738a,a75739a,a75740a,a75744a,a75745a,a75748a,a75751a,a75752a,a75753a,a75757a,a75758a,a75761a,a75764a,a75765a,a75766a,a75770a,a75771a,a75774a,a75777a,a75778a,a75779a,a75783a,a75784a,a75787a,a75790a,a75791a,a75792a,a75796a,a75797a,a75800a,a75803a,a75804a,a75805a,a75809a,a75810a,a75813a,a75816a,a75817a,a75818a,a75822a,a75823a,a75826a,a75829a,a75830a,a75831a,a75835a,a75836a,a75839a,a75842a,a75843a,a75844a,a75848a,a75849a,a75852a,a75855a,a75856a,a75857a,a75861a,a75862a,a75865a,a75868a,a75869a,a75870a,a75874a,a75875a,a75878a,a75881a,a75882a,a75883a,a75887a,a75888a,a75891a,a75894a,a75895a,a75896a,a75900a,a75901a,a75904a,a75907a,a75908a,a75909a,a75913a,a75914a,a75917a,a75920a,a75921a,a75922a,a75926a,a75927a,a75930a,a75933a,a75934a,a75935a,a75939a,a75940a,a75943a,a75946a,a75947a,a75948a,a75952a,a75953a,a75956a,a75959a,a75960a,a75961a,a75965a,a75966a,a75969a,a75972a,a75973a,a75974a,a75978a,a75979a,a75982a,a75985a,a75986a,a75987a,a75991a,a75992a,a75995a,a75998a,a75999a,a76000a,a76004a,a76005a,a76008a,a76011a,a76012a,a76013a,a76017a,a76018a,a76021a,a76024a,a76025a,a76026a,a76030a,a76031a,a76034a,a76037a,a76038a,a76039a,a76043a,a76044a,a76047a,a76050a,a76051a,a76052a,a76056a,a76057a,a76060a,a76063a,a76064a,a76065a,a76069a,a76070a,a76073a,a76076a,a76077a,a76078a,a76082a,a76083a,a76086a,a76089a,a76090a,a76091a,a76095a,a76096a,a76099a,a76102a,a76103a,a76104a,a76108a,a76109a,a76112a,a76115a,a76116a,a76117a,a76121a,a76122a,a76125a,a76128a,a76129a,a76130a,a76134a,a76135a,a76138a,a76141a,a76142a,a76143a,a76147a,a76148a,a76151a,a76154a,a76155a,a76156a,a76160a,a76161a,a76164a,a76167a,a76168a,a76169a,a76173a,a76174a,a76177a,a76180a,a76181a,a76182a,a76186a,a76187a,a76190a,a76193a,a76194a,a76195a,a76199a,a76200a,a76203a,a76206a,a76207a,a76208a,a76212a,a76213a,a76216a,a76219a,a76220a,a76221a,a76225a,a76226a,a76229a,a76232a,a76233a,a76234a,a76238a,a76239a,a76242a,a76245a,a76246a,a76247a,a76251a,a76252a,a76255a,a76258a,a76259a,a76260a,a76264a,a76265a,a76268a,a76271a,a76272a,a76273a,a76277a,a76278a,a76281a,a76284a,a76285a,a76286a,a76290a,a76291a,a76294a,a76297a,a76298a,a76299a,a76303a,a76304a,a76307a,a76310a,a76311a,a76312a,a76316a,a76317a,a76320a,a76323a,a76324a,a76325a,a76329a,a76330a,a76333a,a76336a,a76337a,a76338a,a76342a,a76343a,a76346a,a76349a,a76350a,a76351a,a76355a,a76356a,a76359a,a76362a,a76363a,a76364a,a76368a,a76369a,a76372a,a76375a,a76376a,a76377a,a76381a,a76382a,a76385a,a76388a,a76389a,a76390a,a76394a,a76395a,a76398a,a76401a,a76402a,a76403a,a76407a,a76408a,a76411a,a76414a,a76415a,a76416a,a76420a,a76421a,a76424a,a76427a,a76428a,a76429a,a76433a,a76434a,a76437a,a76440a,a76441a,a76442a,a76446a,a76447a,a76450a,a76453a,a76454a,a76455a,a76459a,a76460a,a76463a,a76466a,a76467a,a76468a,a76472a,a76473a,a76476a,a76479a,a76480a,a76481a,a76485a,a76486a,a76489a,a76492a,a76493a,a76494a,a76498a,a76499a,a76502a,a76505a,a76506a,a76507a,a76511a,a76512a,a76515a,a76518a,a76519a,a76520a,a76524a,a76525a,a76528a,a76531a,a76532a,a76533a,a76537a,a76538a,a76541a,a76544a,a76545a,a76546a,a76550a,a76551a,a76554a,a76557a,a76558a,a76559a,a76563a,a76564a,a76567a,a76570a,a76571a,a76572a,a76576a,a76577a,a76580a,a76583a,a76584a,a76585a,a76589a,a76590a,a76593a,a76596a,a76597a,a76598a,a76602a,a76603a,a76606a,a76609a,a76610a,a76611a,a76615a,a76616a,a76619a,a76622a,a76623a,a76624a,a76628a,a76629a,a76632a,a76635a,a76636a,a76637a,a76641a,a76642a,a76645a,a76648a,a76649a,a76650a,a76654a,a76655a,a76658a,a76661a,a76662a,a76663a,a76667a,a76668a,a76671a,a76674a,a76675a,a76676a,a76680a,a76681a,a76684a,a76687a,a76688a,a76689a,a76693a,a76694a,a76697a,a76700a,a76701a,a76702a,a76706a,a76707a,a76710a,a76713a,a76714a,a76715a,a76719a,a76720a,a76723a,a76726a,a76727a,a76728a,a76732a,a76733a,a76736a,a76739a,a76740a,a76741a,a76745a,a76746a,a76749a,a76752a,a76753a,a76754a,a76758a,a76759a,a76762a,a76765a,a76766a,a76767a,a76771a,a76772a,a76775a,a76778a,a76779a,a76780a,a76784a,a76785a,a76788a,a76791a,a76792a,a76793a,a76797a,a76798a,a76801a,a76804a,a76805a,a76806a,a76810a,a76811a,a76814a,a76817a,a76818a,a76819a,a76823a,a76824a,a76827a,a76830a,a76831a,a76832a,a76836a,a76837a,a76840a,a76843a,a76844a,a76845a,a76849a,a76850a,a76853a,a76856a,a76857a,a76858a,a76862a,a76863a,a76866a,a76869a,a76870a,a76871a,a76875a,a76876a,a76879a,a76882a,a76883a,a76884a,a76888a,a76889a,a76892a,a76895a,a76896a,a76897a,a76901a,a76902a,a76905a,a76908a,a76909a,a76910a,a76914a,a76915a,a76918a,a76921a,a76922a,a76923a,a76927a,a76928a,a76931a,a76934a,a76935a,a76936a,a76940a,a76941a,a76944a,a76947a,a76948a,a76949a,a76953a,a76954a,a76957a,a76960a,a76961a,a76962a,a76966a,a76967a,a76970a,a76973a,a76974a,a76975a,a76979a,a76980a,a76983a,a76986a,a76987a,a76988a,a76992a,a76993a,a76996a,a76999a,a77000a,a77001a,a77005a,a77006a,a77009a,a77012a,a77013a,a77014a,a77018a,a77019a,a77022a,a77025a,a77026a,a77027a,a77031a,a77032a,a77035a,a77038a,a77039a,a77040a,a77044a,a77045a,a77048a,a77051a,a77052a,a77053a,a77057a,a77058a,a77061a,a77064a,a77065a,a77066a,a77070a,a77071a,a77074a,a77077a,a77078a,a77079a,a77083a,a77084a,a77087a,a77090a,a77091a,a77092a,a77096a,a77097a,a77100a,a77103a,a77104a,a77105a,a77109a,a77110a,a77113a,a77116a,a77117a,a77118a,a77122a,a77123a,a77126a,a77129a,a77130a,a77131a,a77135a,a77136a,a77139a,a77142a,a77143a,a77144a,a77148a,a77149a,a77152a,a77155a,a77156a,a77157a,a77161a,a77162a,a77165a,a77168a,a77169a,a77170a,a77174a,a77175a,a77178a,a77181a,a77182a,a77183a,a77187a,a77188a,a77191a,a77194a,a77195a,a77196a,a77200a,a77201a,a77204a,a77207a,a77208a,a77209a,a77213a,a77214a,a77217a,a77220a,a77221a,a77222a,a77226a,a77227a,a77230a,a77233a,a77234a,a77235a,a77239a,a77240a,a77243a,a77246a,a77247a,a77248a,a77252a,a77253a,a77256a,a77259a,a77260a,a77261a,a77265a,a77266a,a77269a,a77272a,a77273a,a77274a,a77278a,a77279a,a77282a,a77285a,a77286a,a77287a,a77291a,a77292a,a77295a,a77298a,a77299a,a77300a,a77304a,a77305a,a77308a,a77311a,a77312a,a77313a,a77317a,a77318a,a77321a,a77324a,a77325a,a77326a,a77330a,a77331a,a77334a,a77337a,a77338a,a77339a,a77343a,a77344a,a77347a,a77350a,a77351a,a77352a,a77356a,a77357a,a77360a,a77363a,a77364a,a77365a,a77369a,a77370a,a77373a,a77376a,a77377a,a77378a,a77382a,a77383a,a77386a,a77389a,a77390a,a77391a,a77395a,a77396a,a77399a,a77402a,a77403a,a77404a,a77408a,a77409a,a77412a,a77415a,a77416a,a77417a,a77421a,a77422a,a77425a,a77428a,a77429a,a77430a,a77434a,a77435a,a77438a,a77441a,a77442a,a77443a,a77447a,a77448a,a77451a,a77454a,a77455a,a77456a,a77460a,a77461a,a77464a,a77467a,a77468a,a77469a,a77473a,a77474a,a77477a,a77480a,a77481a,a77482a,a77486a,a77487a,a77490a,a77493a,a77494a,a77495a,a77499a,a77500a,a77503a,a77506a,a77507a,a77508a,a77512a,a77513a,a77516a,a77519a,a77520a,a77521a,a77525a,a77526a,a77529a,a77532a,a77533a,a77534a,a77538a,a77539a,a77542a,a77545a,a77546a,a77547a,a77551a,a77552a,a77555a,a77558a,a77559a,a77560a,a77564a,a77565a,a77568a,a77571a,a77572a,a77573a,a77577a,a77578a,a77581a,a77584a,a77585a,a77586a,a77590a,a77591a,a77594a,a77597a,a77598a,a77599a,a77603a,a77604a,a77607a,a77610a,a77611a,a77612a,a77616a,a77617a,a77620a,a77623a,a77624a,a77625a,a77629a,a77630a,a77633a,a77636a,a77637a,a77638a,a77642a,a77643a,a77646a,a77649a,a77650a,a77651a,a77655a,a77656a,a77659a,a77662a,a77663a,a77664a,a77668a,a77669a,a77672a,a77675a,a77676a,a77677a,a77681a,a77682a,a77685a,a77688a,a77689a,a77690a,a77694a,a77695a,a77698a,a77701a,a77702a,a77703a,a77707a,a77708a,a77711a,a77714a,a77715a,a77716a,a77720a,a77721a,a77724a,a77727a,a77728a,a77729a,a77733a,a77734a,a77737a,a77740a,a77741a,a77742a,a77746a,a77747a,a77750a,a77753a,a77754a,a77755a,a77759a,a77760a,a77763a,a77766a,a77767a,a77768a,a77772a,a77773a,a77776a,a77779a,a77780a,a77781a,a77785a,a77786a,a77789a,a77792a,a77793a,a77794a,a77798a,a77799a,a77802a,a77805a,a77806a,a77807a,a77811a,a77812a,a77815a,a77818a,a77819a,a77820a,a77824a,a77825a,a77828a,a77831a,a77832a,a77833a,a77837a,a77838a,a77841a,a77844a,a77845a,a77846a,a77850a,a77851a,a77854a,a77857a,a77858a,a77859a,a77863a,a77864a,a77867a,a77870a,a77871a,a77872a,a77876a,a77877a,a77880a,a77883a,a77884a,a77885a,a77889a,a77890a,a77893a,a77896a,a77897a,a77898a,a77902a,a77903a,a77906a,a77909a,a77910a,a77911a,a77915a,a77916a,a77919a,a77922a,a77923a,a77924a,a77928a,a77929a,a77932a,a77935a,a77936a,a77937a,a77941a,a77942a,a77945a,a77948a,a77949a,a77950a,a77954a,a77955a,a77958a,a77961a,a77962a,a77963a,a77967a,a77968a,a77971a,a77974a,a77975a,a77976a,a77980a,a77981a,a77984a,a77987a,a77988a,a77989a,a77993a,a77994a,a77997a,a78000a,a78001a,a78002a,a78006a,a78007a,a78010a,a78013a,a78014a,a78015a,a78019a,a78020a,a78023a,a78026a,a78027a,a78028a,a78032a,a78033a,a78036a,a78039a,a78040a,a78041a,a78045a,a78046a,a78049a,a78052a,a78053a,a78054a,a78058a,a78059a,a78062a,a78065a,a78066a,a78067a,a78071a,a78072a,a78075a,a78078a,a78079a,a78080a,a78084a,a78085a,a78088a,a78091a,a78092a,a78093a,a78097a,a78098a,a78101a,a78104a,a78105a,a78106a,a78110a,a78111a,a78114a,a78117a,a78118a,a78119a,a78123a,a78124a,a78127a,a78130a,a78131a,a78132a,a78136a,a78137a,a78140a,a78143a,a78144a,a78145a,a78149a,a78150a,a78153a,a78156a,a78157a,a78158a,a78162a,a78163a,a78166a,a78169a,a78170a,a78171a,a78175a,a78176a,a78179a,a78182a,a78183a,a78184a,a78188a,a78189a,a78192a,a78195a,a78196a,a78197a,a78201a,a78202a,a78205a,a78208a,a78209a,a78210a,a78214a,a78215a,a78218a,a78221a,a78222a,a78223a,a78227a,a78228a,a78231a,a78234a,a78235a,a78236a,a78240a,a78241a,a78244a,a78247a,a78248a,a78249a,a78253a,a78254a,a78257a,a78260a,a78261a,a78262a,a78266a,a78267a,a78270a,a78273a,a78274a,a78275a,a78279a,a78280a,a78283a,a78286a,a78287a,a78288a,a78292a,a78293a,a78296a,a78299a,a78300a,a78301a,a78305a,a78306a,a78309a,a78312a,a78313a,a78314a,a78318a,a78319a,a78322a,a78325a,a78326a,a78327a,a78331a,a78332a,a78335a,a78338a,a78339a,a78340a,a78344a,a78345a,a78348a,a78351a,a78352a,a78353a,a78357a,a78358a,a78361a,a78364a,a78365a,a78366a,a78370a,a78371a,a78374a,a78377a,a78378a,a78379a,a78383a,a78384a,a78387a,a78390a,a78391a,a78392a,a78396a,a78397a,a78400a,a78403a,a78404a,a78405a,a78409a,a78410a,a78413a,a78416a,a78417a,a78418a,a78422a,a78423a,a78426a,a78429a,a78430a,a78431a,a78435a,a78436a,a78439a,a78442a,a78443a,a78444a,a78448a,a78449a,a78452a,a78455a,a78456a,a78457a,a78461a,a78462a,a78465a,a78468a,a78469a,a78470a,a78474a,a78475a,a78478a,a78481a,a78482a,a78483a,a78487a,a78488a,a78491a,a78494a,a78495a,a78496a,a78500a,a78501a,a78504a,a78507a,a78508a,a78509a,a78513a,a78514a,a78517a,a78520a,a78521a,a78522a,a78526a,a78527a,a78530a,a78533a,a78534a,a78535a,a78539a,a78540a,a78543a,a78546a,a78547a,a78548a,a78552a,a78553a,a78556a,a78559a,a78560a,a78561a,a78565a,a78566a,a78569a,a78572a,a78573a,a78574a,a78578a,a78579a,a78582a,a78585a,a78586a,a78587a,a78591a,a78592a,a78595a,a78598a,a78599a,a78600a,a78604a,a78605a,a78608a,a78611a,a78612a,a78613a,a78617a,a78618a,a78621a,a78624a,a78625a,a78626a,a78630a,a78631a,a78634a,a78637a,a78638a,a78639a,a78643a,a78644a,a78647a,a78650a,a78651a,a78652a,a78656a,a78657a,a78660a,a78663a,a78664a,a78665a,a78669a,a78670a,a78673a,a78676a,a78677a,a78678a,a78682a,a78683a,a78686a,a78689a,a78690a,a78691a,a78695a,a78696a,a78699a,a78702a,a78703a,a78704a,a78708a,a78709a,a78712a,a78715a,a78716a,a78717a,a78721a,a78722a,a78725a,a78728a,a78729a,a78730a,a78734a,a78735a,a78738a,a78741a,a78742a,a78743a,a78747a,a78748a,a78751a,a78754a,a78755a,a78756a,a78760a,a78761a,a78764a,a78767a,a78768a,a78769a,a78773a,a78774a,a78777a,a78780a,a78781a,a78782a,a78786a,a78787a,a78790a,a78793a,a78794a,a78795a,a78799a,a78800a,a78803a,a78806a,a78807a,a78808a,a78812a,a78813a,a78816a,a78819a,a78820a,a78821a,a78825a,a78826a,a78829a,a78832a,a78833a,a78834a,a78838a,a78839a,a78842a,a78845a,a78846a,a78847a,a78851a,a78852a,a78855a,a78858a,a78859a,a78860a,a78864a,a78865a,a78868a,a78871a,a78872a,a78873a,a78877a,a78878a,a78881a,a78884a,a78885a,a78886a,a78890a,a78891a,a78894a,a78897a,a78898a,a78899a,a78903a,a78904a,a78907a,a78910a,a78911a,a78912a,a78916a,a78917a,a78920a,a78923a,a78924a,a78925a,a78929a,a78930a,a78933a,a78936a,a78937a,a78938a,a78942a,a78943a,a78946a,a78949a,a78950a,a78951a,a78955a,a78956a,a78959a,a78962a,a78963a,a78964a,a78968a,a78969a,a78972a,a78975a,a78976a,a78977a,a78981a,a78982a,a78985a,a78988a,a78989a,a78990a,a78994a,a78995a,a78998a,a79001a,a79002a,a79003a,a79007a,a79008a,a79011a,a79014a,a79015a,a79016a,a79020a,a79021a,a79024a,a79027a,a79028a,a79029a,a79033a,a79034a,a79037a,a79040a,a79041a,a79042a,a79046a,a79047a,a79050a,a79053a,a79054a,a79055a,a79059a,a79060a,a79063a,a79066a,a79067a,a79068a,a79072a,a79073a,a79076a,a79079a,a79080a,a79081a,a79085a,a79086a,a79089a,a79092a,a79093a,a79094a,a79098a,a79099a,a79102a,a79105a,a79106a,a79107a,a79111a,a79112a,a79115a,a79118a,a79119a,a79120a,a79124a,a79125a,a79128a,a79131a,a79132a,a79133a,a79137a,a79138a,a79141a,a79144a,a79145a,a79146a,a79150a,a79151a,a79154a,a79157a,a79158a,a79159a,a79163a,a79164a,a79167a,a79170a,a79171a,a79172a,a79176a,a79177a,a79180a,a79183a,a79184a,a79185a,a79189a,a79190a,a79193a,a79196a,a79197a,a79198a,a79202a,a79203a,a79206a,a79209a,a79210a,a79211a,a79215a,a79216a,a79219a,a79222a,a79223a,a79224a,a79228a,a79229a,a79232a,a79235a,a79236a,a79237a,a79241a,a79242a,a79245a,a79248a,a79249a,a79250a,a79254a,a79255a,a79258a,a79261a,a79262a,a79263a,a79267a,a79268a,a79271a,a79274a,a79275a,a79276a,a79280a,a79281a,a79284a,a79287a,a79288a,a79289a,a79293a,a79294a,a79297a,a79300a,a79301a,a79302a,a79306a,a79307a,a79310a,a79313a,a79314a,a79315a,a79319a,a79320a,a79323a,a79326a,a79327a,a79328a,a79332a,a79333a,a79336a,a79339a,a79340a,a79341a,a79345a,a79346a,a79349a,a79352a,a79353a,a79354a,a79358a,a79359a,a79362a,a79365a,a79366a,a79367a,a79371a,a79372a,a79375a,a79378a,a79379a,a79380a,a79384a,a79385a,a79388a,a79391a,a79392a,a79393a,a79397a,a79398a,a79401a,a79404a,a79405a,a79406a,a79410a,a79411a,a79414a,a79417a,a79418a,a79419a,a79423a,a79424a,a79427a,a79430a,a79431a,a79432a,a79436a,a79437a,a79440a,a79443a,a79444a,a79445a,a79449a,a79450a,a79453a,a79456a,a79457a,a79458a,a79462a,a79463a,a79466a,a79469a,a79470a,a79471a,a79475a,a79476a,a79479a,a79482a,a79483a,a79484a,a79488a,a79489a,a79492a,a79495a,a79496a,a79497a,a79501a,a79502a,a79505a,a79508a,a79509a,a79510a,a79514a,a79515a,a79518a,a79521a,a79522a,a79523a,a79527a,a79528a,a79531a,a79534a,a79535a,a79536a,a79540a,a79541a,a79544a,a79547a,a79548a,a79549a,a79553a,a79554a,a79557a,a79560a,a79561a,a79562a,a79566a,a79567a,a79570a,a79573a,a79574a,a79575a,a79579a,a79580a,a79583a,a79586a,a79587a,a79588a,a79592a,a79593a,a79596a,a79599a,a79600a,a79601a,a79605a,a79606a,a79609a,a79612a,a79613a,a79614a,a79618a,a79619a,a79622a,a79625a,a79626a,a79627a,a79631a,a79632a,a79635a,a79638a,a79639a,a79640a,a79644a,a79645a,a79648a,a79651a,a79652a,a79653a,a79657a,a79658a,a79661a,a79664a,a79665a,a79666a,a79670a,a79671a,a79674a,a79677a,a79678a,a79679a,a79683a,a79684a,a79687a,a79690a,a79691a,a79692a,a79696a,a79697a,a79700a,a79703a,a79704a,a79705a,a79709a,a79710a,a79713a,a79716a,a79717a,a79718a,a79722a,a79723a,a79726a,a79729a,a79730a,a79731a,a79735a,a79736a,a79739a,a79742a,a79743a,a79744a,a79748a,a79749a,a79752a,a79755a,a79756a,a79757a,a79761a,a79762a,a79765a,a79768a,a79769a,a79770a,a79774a,a79775a,a79778a,a79781a,a79782a,a79783a,a79787a,a79788a,a79791a,a79794a,a79795a,a79796a,a79800a,a79801a,a79804a,a79807a,a79808a,a79809a,a79813a,a79814a,a79817a,a79820a,a79821a,a79822a,a79826a,a79827a,a79830a,a79833a,a79834a,a79835a,a79839a,a79840a,a79843a,a79846a,a79847a,a79848a,a79852a,a79853a,a79856a,a79859a,a79860a,a79861a,a79865a,a79866a,a79869a,a79872a,a79873a,a79874a,a79878a,a79879a,a79882a,a79885a,a79886a,a79887a,a79891a,a79892a,a79895a,a79898a,a79899a,a79900a,a79904a,a79905a,a79908a,a79911a,a79912a,a79913a,a79917a,a79918a,a79921a,a79924a,a79925a,a79926a,a79930a,a79931a,a79934a,a79937a,a79938a,a79939a,a79943a,a79944a,a79947a,a79950a,a79951a,a79952a,a79956a,a79957a,a79960a,a79963a,a79964a,a79965a,a79969a,a79970a,a79973a,a79976a,a79977a,a79978a,a79982a,a79983a,a79986a,a79989a,a79990a,a79991a,a79995a,a79996a,a79999a,a80002a,a80003a,a80004a,a80008a,a80009a,a80012a,a80015a,a80016a,a80017a,a80021a,a80022a,a80025a,a80028a,a80029a,a80030a,a80034a,a80035a,a80038a,a80041a,a80042a,a80043a,a80047a,a80048a,a80051a,a80054a,a80055a,a80056a,a80060a,a80061a,a80064a,a80067a,a80068a,a80069a,a80073a,a80074a,a80077a,a80080a,a80081a,a80082a,a80086a,a80087a,a80090a,a80093a,a80094a,a80095a,a80099a,a80100a,a80103a,a80106a,a80107a,a80108a,a80112a,a80113a,a80116a,a80119a,a80120a,a80121a,a80125a,a80126a,a80129a,a80132a,a80133a,a80134a,a80138a,a80139a,a80142a,a80145a,a80146a,a80147a,a80151a,a80152a,a80155a,a80158a,a80159a,a80160a,a80164a,a80165a,a80168a,a80171a,a80172a,a80173a,a80177a,a80178a,a80181a,a80184a,a80185a,a80186a,a80190a,a80191a,a80194a,a80197a,a80198a,a80199a,a80203a,a80204a,a80207a,a80210a,a80211a,a80212a,a80216a,a80217a,a80220a,a80223a,a80224a,a80225a,a80229a,a80230a,a80233a,a80236a,a80237a,a80238a,a80242a,a80243a,a80246a,a80249a,a80250a,a80251a,a80255a,a80256a,a80259a,a80262a,a80263a,a80264a,a80268a,a80269a,a80272a,a80275a,a80276a,a80277a,a80281a,a80282a,a80285a,a80288a,a80289a,a80290a,a80294a,a80295a,a80298a,a80301a,a80302a,a80303a,a80307a,a80308a,a80311a,a80314a,a80315a,a80316a,a80320a,a80321a,a80324a,a80327a,a80328a,a80329a,a80333a,a80334a,a80337a,a80340a,a80341a,a80342a,a80346a,a80347a,a80350a,a80353a,a80354a,a80355a,a80359a,a80360a,a80363a,a80366a,a80367a,a80368a,a80372a,a80373a,a80376a,a80379a,a80380a,a80381a,a80385a,a80386a,a80389a,a80392a,a80393a,a80394a,a80398a,a80399a,a80402a,a80405a,a80406a,a80407a,a80411a,a80412a,a80415a,a80418a,a80419a,a80420a,a80424a,a80425a,a80428a,a80431a,a80432a,a80433a,a80437a,a80438a,a80441a,a80444a,a80445a,a80446a,a80450a,a80451a,a80454a,a80457a,a80458a,a80459a,a80463a,a80464a,a80467a,a80470a,a80471a,a80472a,a80476a,a80477a,a80480a,a80483a,a80484a,a80485a,a80489a,a80490a,a80493a,a80496a,a80497a,a80498a,a80502a,a80503a,a80506a,a80509a,a80510a,a80511a,a80515a,a80516a,a80519a,a80522a,a80523a,a80524a,a80528a,a80529a,a80532a,a80535a,a80536a,a80537a,a80541a,a80542a,a80545a,a80548a,a80549a,a80550a,a80554a,a80555a,a80558a,a80561a,a80562a,a80563a,a80567a,a80568a,a80571a,a80574a,a80575a,a80576a,a80580a,a80581a,a80584a,a80587a,a80588a,a80589a,a80593a,a80594a,a80597a,a80600a,a80601a,a80602a,a80606a,a80607a,a80610a,a80613a,a80614a,a80615a,a80619a,a80620a,a80623a,a80626a,a80627a,a80628a,a80632a,a80633a,a80636a,a80639a,a80640a,a80641a,a80645a,a80646a,a80649a,a80652a,a80653a,a80654a,a80658a,a80659a,a80662a,a80665a,a80666a,a80667a,a80671a,a80672a,a80675a,a80678a,a80679a,a80680a,a80684a,a80685a,a80688a,a80691a,a80692a,a80693a,a80697a,a80698a,a80701a,a80704a,a80705a,a80706a,a80710a,a80711a,a80714a,a80717a,a80718a,a80719a,a80723a,a80724a,a80727a,a80730a,a80731a,a80732a,a80736a,a80737a,a80740a,a80743a,a80744a,a80745a,a80749a,a80750a,a80753a,a80756a,a80757a,a80758a,a80762a,a80763a,a80766a,a80769a,a80770a,a80771a,a80775a,a80776a,a80779a,a80782a,a80783a,a80784a,a80788a,a80789a,a80792a,a80795a,a80796a,a80797a,a80801a,a80802a,a80805a,a80808a,a80809a,a80810a,a80814a,a80815a,a80818a,a80821a,a80822a,a80823a,a80827a,a80828a,a80831a,a80834a,a80835a,a80836a,a80840a,a80841a,a80844a,a80847a,a80848a,a80849a,a80853a,a80854a,a80857a,a80860a,a80861a,a80862a,a80866a,a80867a,a80870a,a80873a,a80874a,a80875a,a80879a,a80880a,a80883a,a80886a,a80887a,a80888a,a80892a,a80893a,a80896a,a80899a,a80900a,a80901a,a80905a,a80906a,a80909a,a80912a,a80913a,a80914a,a80918a,a80919a,a80922a,a80925a,a80926a,a80927a,a80931a,a80932a,a80935a,a80938a,a80939a,a80940a,a80944a,a80945a,a80948a,a80951a,a80952a,a80953a,a80957a,a80958a,a80961a,a80964a,a80965a,a80966a,a80970a,a80971a,a80974a,a80977a,a80978a,a80979a,a80983a,a80984a,a80987a,a80990a,a80991a,a80992a,a80996a,a80997a,a81000a,a81003a,a81004a,a81005a,a81009a,a81010a,a81013a,a81016a,a81017a,a81018a,a81022a,a81023a,a81026a,a81029a,a81030a,a81031a,a81035a,a81036a,a81039a,a81042a,a81043a,a81044a,a81048a,a81049a,a81052a,a81055a,a81056a,a81057a,a81061a,a81062a,a81065a,a81068a,a81069a,a81070a,a81074a,a81075a,a81078a,a81081a,a81082a,a81083a,a81087a,a81088a,a81091a,a81094a,a81095a,a81096a,a81100a,a81101a,a81104a,a81107a,a81108a,a81109a,a81113a,a81114a,a81117a,a81120a,a81121a,a81122a,a81126a,a81127a,a81130a,a81133a,a81134a,a81135a,a81139a,a81140a,a81143a,a81146a,a81147a,a81148a,a81152a,a81153a,a81156a,a81159a,a81160a,a81161a,a81165a,a81166a,a81169a,a81172a,a81173a,a81174a,a81178a,a81179a,a81182a,a81185a,a81186a,a81187a,a81191a,a81192a,a81195a,a81198a,a81199a,a81200a,a81204a,a81205a,a81208a,a81211a,a81212a,a81213a,a81217a,a81218a,a81221a,a81224a,a81225a,a81226a,a81230a,a81231a,a81234a,a81237a,a81238a,a81239a,a81243a,a81244a,a81247a,a81250a,a81251a,a81252a,a81256a,a81257a,a81260a,a81263a,a81264a,a81265a,a81269a,a81270a,a81273a,a81276a,a81277a,a81278a,a81282a,a81283a,a81286a,a81289a,a81290a,a81291a,a81295a,a81296a,a81299a,a81302a,a81303a,a81304a,a81308a,a81309a,a81312a,a81315a,a81316a,a81317a,a81321a,a81322a,a81325a,a81328a,a81329a,a81330a,a81334a,a81335a,a81338a,a81341a,a81342a,a81343a,a81347a,a81348a,a81351a,a81354a,a81355a,a81356a,a81360a,a81361a,a81364a,a81367a,a81368a,a81369a,a81373a,a81374a,a81377a,a81380a,a81381a,a81382a,a81386a,a81387a,a81390a,a81393a,a81394a,a81395a,a81399a,a81400a,a81403a,a81406a,a81407a,a81408a,a81412a,a81413a,a81416a,a81419a,a81420a,a81421a,a81425a,a81426a,a81429a,a81432a,a81433a,a81434a,a81438a,a81439a,a81442a,a81445a,a81446a,a81447a,a81451a,a81452a,a81455a,a81458a,a81459a,a81460a,a81464a,a81465a,a81468a,a81471a,a81472a,a81473a,a81477a,a81478a,a81481a,a81484a,a81485a,a81486a,a81490a,a81491a,a81494a,a81497a,a81498a,a81499a,a81503a,a81504a,a81507a,a81510a,a81511a,a81512a,a81516a,a81517a,a81520a,a81523a,a81524a,a81525a,a81529a,a81530a,a81533a,a81536a,a81537a,a81538a,a81542a,a81543a,a81546a,a81549a,a81550a,a81551a,a81555a,a81556a,a81559a,a81562a,a81563a,a81564a,a81568a,a81569a,a81572a,a81575a,a81576a,a81577a,a81581a,a81582a,a81585a,a81588a,a81589a,a81590a,a81594a,a81595a,a81598a,a81601a,a81602a,a81603a,a81607a,a81608a,a81611a,a81614a,a81615a,a81616a,a81620a,a81621a,a81624a,a81627a,a81628a,a81629a,a81633a,a81634a,a81637a,a81640a,a81641a,a81642a,a81646a,a81647a,a81650a,a81653a,a81654a,a81655a,a81659a,a81660a,a81663a,a81666a,a81667a,a81668a,a81672a,a81673a,a81676a,a81679a,a81680a,a81681a,a81685a,a81686a,a81689a,a81692a,a81693a,a81694a,a81698a,a81699a,a81702a,a81705a,a81706a,a81707a,a81711a,a81712a,a81715a,a81718a,a81719a,a81720a,a81724a,a81725a,a81728a,a81731a,a81732a,a81733a,a81737a,a81738a,a81741a,a81744a,a81745a,a81746a,a81750a,a81751a,a81754a,a81757a,a81758a,a81759a,a81763a,a81764a,a81767a,a81770a,a81771a,a81772a,a81776a,a81777a,a81780a,a81783a,a81784a,a81785a,a81789a,a81790a,a81793a,a81796a,a81797a,a81798a,a81802a,a81803a,a81806a,a81809a,a81810a,a81811a,a81815a,a81816a,a81819a,a81822a,a81823a,a81824a,a81828a,a81829a,a81832a,a81835a,a81836a,a81837a,a81841a,a81842a,a81845a,a81848a,a81849a,a81850a,a81854a,a81855a,a81858a,a81861a,a81862a,a81863a,a81867a,a81868a,a81871a,a81874a,a81875a,a81876a,a81880a,a81881a,a81884a,a81887a,a81888a,a81889a,a81893a,a81894a,a81897a,a81900a,a81901a,a81902a,a81906a,a81907a,a81910a,a81913a,a81914a,a81915a,a81919a,a81920a,a81923a,a81926a,a81927a,a81928a,a81932a,a81933a,a81936a,a81939a,a81940a,a81941a,a81945a,a81946a,a81949a,a81952a,a81953a,a81954a,a81958a,a81959a,a81962a,a81965a,a81966a,a81967a,a81971a,a81972a,a81975a,a81978a,a81979a,a81980a,a81984a,a81985a,a81988a,a81991a,a81992a,a81993a,a81997a,a81998a,a82001a,a82004a,a82005a,a82006a,a82010a,a82011a,a82014a,a82017a,a82018a,a82019a,a82023a,a82024a,a82027a,a82030a,a82031a,a82032a,a82036a,a82037a,a82040a,a82043a,a82044a,a82045a,a82049a,a82050a,a82053a,a82056a,a82057a,a82058a,a82062a,a82063a,a82066a,a82069a,a82070a,a82071a,a82075a,a82076a,a82079a,a82082a,a82083a,a82084a,a82088a,a82089a,a82092a,a82095a,a82096a,a82097a,a82101a,a82102a,a82105a,a82108a,a82109a,a82110a,a82114a,a82115a,a82118a,a82121a,a82122a,a82123a,a82127a,a82128a,a82131a,a82134a,a82135a,a82136a,a82140a,a82141a,a82144a,a82147a,a82148a,a82149a,a82153a,a82154a,a82157a,a82160a,a82161a,a82162a,a82166a,a82167a,a82170a,a82173a,a82174a,a82175a,a82179a,a82180a,a82183a,a82186a,a82187a,a82188a,a82192a,a82193a,a82196a,a82199a,a82200a,a82201a,a82205a,a82206a,a82209a,a82212a,a82213a,a82214a,a82218a,a82219a,a82222a,a82225a,a82226a,a82227a,a82231a,a82232a,a82235a,a82238a,a82239a,a82240a,a82244a,a82245a,a82248a,a82251a,a82252a,a82253a,a82257a,a82258a,a82261a,a82264a,a82265a,a82266a,a82270a,a82271a,a82274a,a82277a,a82278a,a82279a,a82283a,a82284a,a82287a,a82290a,a82291a,a82292a,a82296a,a82297a,a82300a,a82303a,a82304a,a82305a,a82309a,a82310a,a82313a,a82316a,a82317a,a82318a,a82322a,a82323a,a82326a,a82329a,a82330a,a82331a,a82335a,a82336a,a82339a,a82342a,a82343a,a82344a,a82348a,a82349a,a82352a,a82355a,a82356a,a82357a,a82361a,a82362a,a82365a,a82368a,a82369a,a82370a,a82374a,a82375a,a82378a,a82381a,a82382a,a82383a,a82387a,a82388a,a82391a,a82394a,a82395a,a82396a,a82400a,a82401a,a82404a,a82407a,a82408a,a82409a,a82413a,a82414a,a82417a,a82420a,a82421a,a82422a,a82426a,a82427a,a82430a,a82433a,a82434a,a82435a,a82439a,a82440a,a82443a,a82446a,a82447a,a82448a,a82452a,a82453a,a82456a,a82459a,a82460a,a82461a,a82465a,a82466a,a82469a,a82472a,a82473a,a82474a,a82478a,a82479a,a82482a,a82485a,a82486a,a82487a,a82491a,a82492a,a82495a,a82498a,a82499a,a82500a,a82504a,a82505a,a82508a,a82511a,a82512a,a82513a,a82517a,a82518a,a82521a,a82524a,a82525a,a82526a,a82530a,a82531a,a82534a,a82537a,a82538a,a82539a,a82543a,a82544a,a82547a,a82550a,a82551a,a82552a,a82556a,a82557a,a82560a,a82563a,a82564a,a82565a,a82569a,a82570a,a82573a,a82576a,a82577a,a82578a,a82582a,a82583a,a82586a,a82589a,a82590a,a82591a,a82595a,a82596a,a82599a,a82602a,a82603a,a82604a,a82608a,a82609a,a82612a,a82615a,a82616a,a82617a,a82621a,a82622a,a82625a,a82628a,a82629a,a82630a,a82634a,a82635a,a82638a,a82641a,a82642a,a82643a,a82647a,a82648a,a82651a,a82654a,a82655a,a82656a,a82660a,a82661a,a82664a,a82667a,a82668a,a82669a,a82673a,a82674a,a82677a,a82680a,a82681a,a82682a,a82686a,a82687a,a82690a,a82693a,a82694a,a82695a,a82699a,a82700a,a82703a,a82706a,a82707a,a82708a,a82712a,a82713a,a82716a,a82719a,a82720a,a82721a,a82725a,a82726a,a82729a,a82732a,a82733a,a82734a,a82738a,a82739a,a82742a,a82745a,a82746a,a82747a,a82751a,a82752a,a82755a,a82758a,a82759a,a82760a,a82764a,a82765a,a82768a,a82771a,a82772a,a82773a,a82777a,a82778a,a82781a,a82784a,a82785a,a82786a,a82790a,a82791a,a82794a,a82797a,a82798a,a82799a,a82803a,a82804a,a82807a,a82810a,a82811a,a82812a,a82816a,a82817a,a82820a,a82823a,a82824a,a82825a,a82829a,a82830a,a82833a,a82836a,a82837a,a82838a,a82842a,a82843a,a82846a,a82849a,a82850a,a82851a,a82855a,a82856a,a82859a,a82862a,a82863a,a82864a,a82868a,a82869a,a82872a,a82875a,a82876a,a82877a,a82881a,a82882a,a82885a,a82888a,a82889a,a82890a,a82894a,a82895a,a82898a,a82901a,a82902a,a82903a,a82907a,a82908a,a82911a,a82914a,a82915a,a82916a,a82920a,a82921a,a82924a,a82927a,a82928a,a82929a,a82933a,a82934a,a82937a,a82940a,a82941a,a82942a,a82946a,a82947a,a82950a,a82953a,a82954a,a82955a,a82959a,a82960a,a82963a,a82966a,a82967a,a82968a,a82972a,a82973a,a82976a,a82979a,a82980a,a82981a,a82985a,a82986a,a82989a,a82992a,a82993a,a82994a,a82998a,a82999a,a83002a,a83005a,a83006a,a83007a,a83011a,a83012a,a83015a,a83018a,a83019a,a83020a,a83024a,a83025a,a83028a,a83031a,a83032a,a83033a,a83037a,a83038a,a83041a,a83044a,a83045a,a83046a,a83050a,a83051a,a83054a,a83057a,a83058a,a83059a,a83063a,a83064a,a83067a,a83070a,a83071a,a83072a,a83076a,a83077a,a83080a,a83083a,a83084a,a83085a,a83089a,a83090a,a83093a,a83096a,a83097a,a83098a,a83102a,a83103a,a83106a,a83109a,a83110a,a83111a,a83115a,a83116a,a83119a,a83122a,a83123a,a83124a,a83128a,a83129a,a83132a,a83135a,a83136a,a83137a,a83141a,a83142a,a83145a,a83148a,a83149a,a83150a,a83154a,a83155a,a83158a,a83161a,a83162a,a83163a,a83167a,a83168a,a83171a,a83174a,a83175a,a83176a,a83180a,a83181a,a83184a,a83187a,a83188a,a83189a,a83193a,a83194a,a83197a,a83200a,a83201a,a83202a,a83206a,a83207a,a83210a,a83213a,a83214a,a83215a,a83219a,a83220a,a83223a,a83226a,a83227a,a83228a,a83232a,a83233a,a83236a,a83239a,a83240a,a83241a,a83245a,a83246a,a83249a,a83252a,a83253a,a83254a,a83258a,a83259a,a83262a,a83265a,a83266a,a83267a,a83271a,a83272a,a83275a,a83278a,a83279a,a83280a,a83284a,a83285a,a83288a,a83291a,a83292a,a83293a,a83297a,a83298a,a83301a,a83304a,a83305a,a83306a,a83310a,a83311a,a83314a,a83317a,a83318a,a83319a,a83323a,a83324a,a83327a,a83330a,a83331a,a83332a,a83336a,a83337a,a83340a,a83343a,a83344a,a83345a,a83349a,a83350a,a83353a,a83356a,a83357a,a83358a,a83362a,a83363a,a83366a,a83369a,a83370a,a83371a,a83375a,a83376a,a83379a,a83382a,a83383a,a83384a,a83388a,a83389a,a83392a,a83395a,a83396a,a83397a,a83401a,a83402a,a83405a,a83408a,a83409a,a83410a,a83414a,a83415a,a83418a,a83421a,a83422a,a83423a,a83427a,a83428a,a83431a,a83434a,a83435a,a83436a,a83440a,a83441a,a83444a,a83447a,a83448a,a83449a,a83453a,a83454a,a83457a,a83460a,a83461a,a83462a,a83466a,a83467a,a83470a,a83473a,a83474a,a83475a,a83479a,a83480a,a83483a,a83486a,a83487a,a83488a,a83492a,a83493a,a83496a,a83499a,a83500a,a83501a,a83505a,a83506a,a83509a,a83512a,a83513a,a83514a,a83518a,a83519a,a83522a,a83525a,a83526a,a83527a,a83531a,a83532a,a83535a,a83538a,a83539a,a83540a,a83544a,a83545a,a83548a,a83551a,a83552a,a83553a,a83557a,a83558a,a83561a,a83564a,a83565a,a83566a,a83570a,a83571a,a83574a,a83577a,a83578a,a83579a,a83583a,a83584a,a83587a,a83590a,a83591a,a83592a,a83596a,a83597a,a83600a,a83603a,a83604a,a83605a,a83609a,a83610a,a83613a,a83616a,a83617a,a83618a,a83622a,a83623a,a83626a,a83629a,a83630a,a83631a,a83635a,a83636a,a83639a,a83642a,a83643a,a83644a,a83648a,a83649a,a83652a,a83655a,a83656a,a83657a,a83661a,a83662a,a83665a,a83668a,a83669a,a83670a,a83674a,a83675a,a83678a,a83681a,a83682a,a83683a,a83687a,a83688a,a83691a,a83694a,a83695a,a83696a,a83700a,a83701a,a83704a,a83707a,a83708a,a83709a,a83713a,a83714a,a83717a,a83720a,a83721a,a83722a,a83726a,a83727a,a83730a,a83733a,a83734a,a83735a,a83739a,a83740a,a83743a,a83746a,a83747a,a83748a,a83752a,a83753a,a83756a,a83759a,a83760a,a83761a,a83765a,a83766a,a83769a,a83772a,a83773a,a83774a,a83778a,a83779a,a83782a,a83785a,a83786a,a83787a,a83791a,a83792a,a83795a,a83798a,a83799a,a83800a,a83804a,a83805a,a83808a,a83811a,a83812a,a83813a,a83817a,a83818a,a83821a,a83824a,a83825a,a83826a,a83830a,a83831a,a83834a,a83837a,a83838a,a83839a,a83843a,a83844a,a83847a,a83850a,a83851a,a83852a,a83856a,a83857a,a83860a,a83863a,a83864a,a83865a,a83869a,a83870a,a83873a,a83876a,a83877a,a83878a,a83882a,a83883a,a83886a,a83889a,a83890a,a83891a,a83895a,a83896a,a83899a,a83902a,a83903a,a83904a,a83908a,a83909a,a83912a,a83915a,a83916a,a83917a,a83921a,a83922a,a83925a,a83928a,a83929a,a83930a,a83934a,a83935a,a83938a,a83941a,a83942a,a83943a,a83947a,a83948a,a83951a,a83954a,a83955a,a83956a,a83960a,a83961a,a83964a,a83967a,a83968a,a83969a,a83973a,a83974a,a83977a,a83980a,a83981a,a83982a,a83986a,a83987a,a83990a,a83993a,a83994a,a83995a,a83999a,a84000a,a84003a,a84006a,a84007a,a84008a,a84012a,a84013a,a84016a,a84019a,a84020a,a84021a,a84025a,a84026a,a84029a,a84032a,a84033a,a84034a,a84038a,a84039a,a84042a,a84045a,a84046a,a84047a,a84051a,a84052a,a84055a,a84058a,a84059a,a84060a,a84064a,a84065a,a84068a,a84071a,a84072a,a84073a,a84077a,a84078a,a84081a,a84084a,a84085a,a84086a,a84090a,a84091a,a84094a,a84097a,a84098a,a84099a,a84103a,a84104a,a84107a,a84110a,a84111a,a84112a,a84116a,a84117a,a84120a,a84123a,a84124a,a84125a,a84129a,a84130a,a84133a,a84136a,a84137a,a84138a,a84142a,a84143a,a84146a,a84149a,a84150a,a84151a,a84155a,a84156a,a84159a,a84162a,a84163a,a84164a,a84168a,a84169a,a84172a,a84175a,a84176a,a84177a,a84181a,a84182a,a84185a,a84188a,a84189a,a84190a,a84194a,a84195a,a84198a,a84201a,a84202a,a84203a,a84207a,a84208a,a84211a,a84214a,a84215a,a84216a,a84220a,a84221a,a84224a,a84227a,a84228a,a84229a,a84233a,a84234a,a84237a,a84240a,a84241a,a84242a,a84246a,a84247a,a84250a,a84253a,a84254a,a84255a,a84259a,a84260a,a84263a,a84266a,a84267a,a84268a,a84272a,a84273a,a84276a,a84279a,a84280a,a84281a,a84285a,a84286a,a84289a,a84292a,a84293a,a84294a,a84298a,a84299a,a84302a,a84305a,a84306a,a84307a,a84311a,a84312a,a84315a,a84318a,a84319a,a84320a,a84324a,a84325a,a84328a,a84331a,a84332a,a84333a,a84337a,a84338a,a84341a,a84344a,a84345a,a84346a,a84350a,a84351a,a84354a,a84357a,a84358a,a84359a,a84363a,a84364a,a84367a,a84370a,a84371a,a84372a,a84376a,a84377a,a84380a,a84383a,a84384a,a84385a,a84389a,a84390a,a84393a,a84396a,a84397a,a84398a,a84402a,a84403a,a84406a,a84409a,a84410a,a84411a,a84415a,a84416a,a84419a,a84422a,a84423a,a84424a,a84428a,a84429a,a84432a,a84435a,a84436a,a84437a,a84441a,a84442a,a84445a,a84448a,a84449a,a84450a,a84454a,a84455a,a84458a,a84461a,a84462a,a84463a,a84467a,a84468a,a84471a,a84474a,a84475a,a84476a,a84480a,a84481a,a84484a,a84487a,a84488a,a84489a,a84493a,a84494a,a84497a,a84500a,a84501a,a84502a,a84506a,a84507a,a84510a,a84513a,a84514a,a84515a,a84519a,a84520a,a84523a,a84526a,a84527a,a84528a,a84532a,a84533a,a84536a,a84539a,a84540a,a84541a,a84545a,a84546a,a84549a,a84552a,a84553a,a84554a,a84558a,a84559a,a84562a,a84565a,a84566a,a84567a,a84571a,a84572a,a84575a,a84578a,a84579a,a84580a,a84584a,a84585a,a84588a,a84591a,a84592a,a84593a,a84597a,a84598a,a84601a,a84604a,a84605a,a84606a,a84610a,a84611a,a84614a,a84617a,a84618a,a84619a,a84623a,a84624a,a84627a,a84630a,a84631a,a84632a,a84636a,a84637a,a84640a,a84643a,a84644a,a84645a,a84649a,a84650a,a84653a,a84656a,a84657a,a84658a,a84662a,a84663a,a84666a,a84669a,a84670a,a84671a,a84675a,a84676a,a84679a,a84682a,a84683a,a84684a,a84688a,a84689a,a84692a,a84695a,a84696a,a84697a,a84701a,a84702a,a84705a,a84708a,a84709a,a84710a,a84714a,a84715a,a84718a,a84721a,a84722a,a84723a,a84727a,a84728a,a84731a,a84734a,a84735a,a84736a,a84740a,a84741a,a84744a,a84747a,a84748a,a84749a,a84753a,a84754a,a84757a,a84760a,a84761a,a84762a,a84766a,a84767a,a84770a,a84773a,a84774a,a84775a,a84779a,a84780a,a84783a,a84786a,a84787a,a84788a,a84792a,a84793a,a84796a,a84799a,a84800a,a84801a,a84805a,a84806a,a84809a,a84812a,a84813a,a84814a,a84818a,a84819a,a84822a,a84825a,a84826a,a84827a,a84831a,a84832a,a84835a,a84838a,a84839a,a84840a,a84844a,a84845a,a84848a,a84851a,a84852a,a84853a,a84857a,a84858a,a84861a,a84864a,a84865a,a84866a,a84870a,a84871a,a84874a,a84877a,a84878a,a84879a,a84883a,a84884a,a84887a,a84890a,a84891a,a84892a,a84896a,a84897a,a84900a,a84903a,a84904a,a84905a,a84909a,a84910a,a84913a,a84916a,a84917a,a84918a,a84922a,a84923a,a84926a,a84929a,a84930a,a84931a,a84935a,a84936a,a84939a,a84942a,a84943a,a84944a,a84948a,a84949a,a84952a,a84955a,a84956a,a84957a,a84961a,a84962a,a84965a,a84968a,a84969a,a84970a,a84974a,a84975a,a84978a,a84981a,a84982a,a84983a,a84987a,a84988a,a84991a,a84994a,a84995a,a84996a,a85000a,a85001a,a85004a,a85007a,a85008a,a85009a,a85013a,a85014a,a85017a,a85020a,a85021a,a85022a,a85026a,a85027a,a85030a,a85033a,a85034a,a85035a,a85039a,a85040a,a85043a,a85046a,a85047a,a85048a,a85052a,a85053a,a85056a,a85059a,a85060a,a85061a,a85065a,a85066a,a85069a,a85072a,a85073a,a85074a,a85078a,a85079a,a85082a,a85085a,a85086a,a85087a,a85091a,a85092a,a85095a,a85098a,a85099a,a85100a,a85104a,a85105a,a85108a,a85111a,a85112a,a85113a,a85117a,a85118a,a85121a,a85124a,a85125a,a85126a,a85130a,a85131a,a85134a,a85137a,a85138a,a85139a,a85143a,a85144a,a85147a,a85150a,a85151a,a85152a,a85156a,a85157a,a85160a,a85163a,a85164a,a85165a,a85169a,a85170a,a85173a,a85176a,a85177a,a85178a,a85182a,a85183a,a85186a,a85189a,a85190a,a85191a,a85195a,a85196a,a85199a,a85202a,a85203a,a85204a,a85208a,a85209a,a85212a,a85215a,a85216a,a85217a,a85221a,a85222a,a85225a,a85228a,a85229a,a85230a,a85234a,a85235a,a85238a,a85241a,a85242a,a85243a,a85247a,a85248a,a85251a,a85254a,a85255a,a85256a,a85260a,a85261a,a85264a,a85267a,a85268a,a85269a,a85273a,a85274a,a85277a,a85280a,a85281a,a85282a,a85286a,a85287a,a85290a,a85293a,a85294a,a85295a,a85299a,a85300a,a85303a,a85306a,a85307a,a85308a,a85312a,a85313a,a85316a,a85319a,a85320a,a85321a,a85325a,a85326a,a85329a,a85332a,a85333a,a85334a,a85338a,a85339a,a85342a,a85345a,a85346a,a85347a,a85351a,a85352a,a85355a,a85358a,a85359a,a85360a,a85364a,a85365a,a85368a,a85371a,a85372a,a85373a,a85377a,a85378a,a85381a,a85384a,a85385a,a85386a,a85390a,a85391a,a85394a,a85397a,a85398a,a85399a,a85403a,a85404a,a85407a,a85410a,a85411a,a85412a,a85416a,a85417a,a85420a,a85423a,a85424a,a85425a,a85429a,a85430a,a85433a,a85436a,a85437a,a85438a,a85442a,a85443a,a85446a,a85449a,a85450a,a85451a,a85455a,a85456a,a85459a,a85462a,a85463a,a85464a,a85468a,a85469a,a85472a,a85475a,a85476a,a85477a,a85481a,a85482a,a85485a,a85488a,a85489a,a85490a,a85494a,a85495a,a85498a,a85501a,a85502a,a85503a,a85507a,a85508a,a85511a,a85514a,a85515a,a85516a,a85520a,a85521a,a85524a,a85527a,a85528a,a85529a,a85533a,a85534a,a85537a,a85540a,a85541a,a85542a,a85546a,a85547a,a85550a,a85553a,a85554a,a85555a,a85559a,a85560a,a85563a,a85566a,a85567a,a85568a,a85572a,a85573a,a85576a,a85579a,a85580a,a85581a,a85585a,a85586a,a85589a,a85592a,a85593a,a85594a,a85598a,a85599a,a85602a,a85605a,a85606a,a85607a,a85611a,a85612a,a85615a,a85618a,a85619a,a85620a,a85624a,a85625a,a85628a,a85631a,a85632a,a85633a,a85637a,a85638a,a85641a,a85644a,a85645a,a85646a,a85650a,a85651a,a85654a,a85657a,a85658a,a85659a,a85663a,a85664a,a85667a,a85670a,a85671a,a85672a,a85676a,a85677a,a85680a,a85683a,a85684a,a85685a,a85689a,a85690a,a85693a,a85696a,a85697a,a85698a,a85702a,a85703a,a85706a,a85709a,a85710a,a85711a,a85715a,a85716a,a85719a,a85722a,a85723a,a85724a,a85728a,a85729a,a85732a,a85735a,a85736a,a85737a,a85741a,a85742a,a85745a,a85748a,a85749a,a85750a,a85754a,a85755a,a85758a,a85761a,a85762a,a85763a,a85767a,a85768a,a85771a,a85774a,a85775a,a85776a,a85780a,a85781a,a85784a,a85787a,a85788a,a85789a,a85793a,a85794a,a85797a,a85800a,a85801a,a85802a,a85806a,a85807a,a85810a,a85813a,a85814a,a85815a,a85819a,a85820a,a85823a,a85826a,a85827a,a85828a,a85832a,a85833a,a85836a,a85839a,a85840a,a85841a,a85845a,a85846a,a85849a,a85852a,a85853a,a85854a,a85858a,a85859a,a85862a,a85865a,a85866a,a85867a,a85871a,a85872a,a85875a,a85878a,a85879a,a85880a,a85884a,a85885a,a85888a,a85891a,a85892a,a85893a,a85897a,a85898a,a85901a,a85904a,a85905a,a85906a,a85910a,a85911a,a85914a,a85917a,a85918a,a85919a,a85923a,a85924a,a85927a,a85930a,a85931a,a85932a,a85936a,a85937a,a85940a,a85943a,a85944a,a85945a,a85949a,a85950a,a85953a,a85956a,a85957a,a85958a,a85962a,a85963a,a85966a,a85969a,a85970a,a85971a,a85975a,a85976a,a85979a,a85982a,a85983a,a85984a,a85988a,a85989a,a85992a,a85995a,a85996a,a85997a,a86001a,a86002a,a86005a,a86008a,a86009a,a86010a,a86014a,a86015a,a86018a,a86021a,a86022a,a86023a,a86027a,a86028a,a86031a,a86034a,a86035a,a86036a,a86040a,a86041a,a86044a,a86047a,a86048a,a86049a,a86053a,a86054a,a86057a,a86060a,a86061a,a86062a,a86066a,a86067a,a86070a,a86073a,a86074a,a86075a,a86079a,a86080a,a86083a,a86086a,a86087a,a86088a,a86092a,a86093a,a86096a,a86099a,a86100a,a86101a,a86105a,a86106a,a86109a,a86112a,a86113a,a86114a,a86118a,a86119a,a86122a,a86125a,a86126a,a86127a,a86131a,a86132a,a86135a,a86138a,a86139a,a86140a,a86144a,a86145a,a86148a,a86151a,a86152a,a86153a,a86157a,a86158a,a86161a,a86164a,a86165a,a86166a,a86170a,a86171a,a86174a,a86177a,a86178a,a86179a,a86183a,a86184a,a86187a,a86190a,a86191a,a86192a,a86196a,a86197a,a86200a,a86203a,a86204a,a86205a,a86209a,a86210a,a86213a,a86216a,a86217a,a86218a,a86222a,a86223a,a86226a,a86229a,a86230a,a86231a,a86235a,a86236a,a86239a,a86242a,a86243a,a86244a,a86248a,a86249a,a86252a,a86255a,a86256a,a86257a,a86261a,a86262a,a86265a,a86268a,a86269a,a86270a,a86274a,a86275a,a86278a,a86281a,a86282a,a86283a,a86287a,a86288a,a86291a,a86294a,a86295a,a86296a,a86300a,a86301a,a86304a,a86307a,a86308a,a86309a,a86313a,a86314a,a86317a,a86320a,a86321a,a86322a,a86326a,a86327a,a86330a,a86333a,a86334a,a86335a,a86339a,a86340a,a86343a,a86346a,a86347a,a86348a,a86352a,a86353a,a86356a,a86359a,a86360a,a86361a,a86365a,a86366a,a86369a,a86372a,a86373a,a86374a,a86378a,a86379a,a86382a,a86385a,a86386a,a86387a,a86391a,a86392a,a86395a,a86398a,a86399a,a86400a,a86404a,a86405a,a86408a,a86411a,a86412a,a86413a,a86417a,a86418a,a86421a,a86424a,a86425a,a86426a,a86430a,a86431a,a86434a,a86437a,a86438a,a86439a,a86443a,a86444a,a86447a,a86450a,a86451a,a86452a,a86456a,a86457a,a86460a,a86463a,a86464a,a86465a,a86469a,a86470a,a86473a,a86476a,a86477a,a86478a,a86482a,a86483a,a86486a,a86489a,a86490a,a86491a,a86495a,a86496a,a86499a,a86502a,a86503a,a86504a,a86508a,a86509a,a86512a,a86515a,a86516a,a86517a,a86521a,a86522a,a86525a,a86528a,a86529a,a86530a,a86534a,a86535a,a86538a,a86541a,a86542a,a86543a,a86547a,a86548a,a86551a,a86554a,a86555a,a86556a,a86560a,a86561a,a86564a,a86567a,a86568a,a86569a,a86573a,a86574a,a86577a,a86580a,a86581a,a86582a,a86586a,a86587a,a86590a,a86593a,a86594a,a86595a,a86599a,a86600a,a86603a,a86606a,a86607a,a86608a,a86612a,a86613a,a86616a,a86619a,a86620a,a86621a,a86625a,a86626a,a86629a,a86632a,a86633a,a86634a,a86638a,a86639a,a86642a,a86645a,a86646a,a86647a,a86651a,a86652a,a86655a,a86658a,a86659a,a86660a,a86664a,a86665a,a86668a,a86671a,a86672a,a86673a,a86677a,a86678a,a86681a,a86684a,a86685a,a86686a,a86690a,a86691a,a86694a,a86697a,a86698a,a86699a,a86703a,a86704a,a86707a,a86710a,a86711a,a86712a,a86716a,a86717a,a86720a,a86723a,a86724a,a86725a,a86729a,a86730a,a86733a,a86736a,a86737a,a86738a,a86742a,a86743a,a86746a,a86749a,a86750a,a86751a,a86755a,a86756a,a86759a,a86762a,a86763a,a86764a,a86768a,a86769a,a86772a,a86775a,a86776a,a86777a,a86781a,a86782a,a86785a,a86788a,a86789a,a86790a,a86794a,a86795a,a86798a,a86801a,a86802a,a86803a,a86806a,a86809a,a86810a,a86813a,a86816a,a86817a,a86818a,a86822a,a86823a,a86826a,a86829a,a86830a,a86831a,a86834a,a86837a,a86838a,a86841a,a86844a,a86845a,a86846a,a86850a,a86851a,a86854a,a86857a,a86858a,a86859a,a86862a,a86865a,a86866a,a86869a,a86872a,a86873a,a86874a,a86878a,a86879a,a86882a,a86885a,a86886a,a86887a,a86890a,a86893a,a86894a,a86897a,a86900a,a86901a,a86902a,a86906a,a86907a,a86910a,a86913a,a86914a,a86915a,a86918a,a86921a,a86922a,a86925a,a86928a,a86929a,a86930a,a86934a,a86935a,a86938a,a86941a,a86942a,a86943a,a86946a,a86949a,a86950a,a86953a,a86956a,a86957a,a86958a,a86962a,a86963a,a86966a,a86969a,a86970a,a86971a,a86974a,a86977a,a86978a,a86981a,a86984a,a86985a,a86986a,a86990a,a86991a,a86994a,a86997a,a86998a,a86999a,a87002a,a87005a,a87006a,a87009a,a87012a,a87013a,a87014a,a87018a,a87019a,a87022a,a87025a,a87026a,a87027a,a87030a,a87033a,a87034a,a87037a,a87040a,a87041a,a87042a,a87046a,a87047a,a87050a,a87053a,a87054a,a87055a,a87058a,a87061a,a87062a,a87065a,a87068a,a87069a,a87070a,a87074a,a87075a,a87078a,a87081a,a87082a,a87083a,a87086a,a87089a,a87090a,a87093a,a87096a,a87097a,a87098a,a87102a,a87103a,a87106a,a87109a,a87110a,a87111a,a87114a,a87117a,a87118a,a87121a,a87124a,a87125a,a87126a,a87130a,a87131a,a87134a,a87137a,a87138a,a87139a,a87142a,a87145a,a87146a,a87149a,a87152a,a87153a,a87154a,a87158a,a87159a,a87162a,a87165a,a87166a,a87167a,a87170a,a87173a,a87174a,a87177a,a87180a,a87181a,a87182a,a87186a,a87187a,a87190a,a87193a,a87194a,a87195a,a87198a,a87201a,a87202a,a87205a,a87208a,a87209a,a87210a,a87214a,a87215a,a87218a,a87221a,a87222a,a87223a,a87226a,a87229a,a87230a,a87233a,a87236a,a87237a,a87238a,a87242a,a87243a,a87246a,a87249a,a87250a,a87251a,a87254a,a87257a,a87258a,a87261a,a87264a,a87265a,a87266a,a87270a,a87271a,a87274a,a87277a,a87278a,a87279a,a87282a,a87285a,a87286a,a87289a,a87292a,a87293a,a87294a,a87298a,a87299a,a87302a,a87305a,a87306a,a87307a,a87310a,a87313a,a87314a,a87317a,a87320a,a87321a,a87322a,a87326a,a87327a,a87330a,a87333a,a87334a,a87335a,a87338a,a87341a,a87342a,a87345a,a87348a,a87349a,a87350a,a87354a,a87355a,a87358a,a87361a,a87362a,a87363a,a87366a,a87369a,a87370a,a87373a,a87376a,a87377a,a87378a,a87382a,a87383a,a87386a,a87389a,a87390a,a87391a,a87394a,a87397a,a87398a,a87401a,a87404a,a87405a,a87406a,a87410a,a87411a,a87414a,a87417a,a87418a,a87419a,a87422a,a87425a,a87426a,a87429a,a87432a,a87433a,a87434a,a87438a,a87439a,a87442a,a87445a,a87446a,a87447a,a87450a,a87453a,a87454a,a87457a,a87460a,a87461a,a87462a,a87466a,a87467a,a87470a,a87473a,a87474a,a87475a,a87478a,a87481a,a87482a,a87485a,a87488a,a87489a,a87490a,a87494a,a87495a,a87498a,a87501a,a87502a,a87503a,a87506a,a87509a,a87510a,a87513a,a87516a,a87517a,a87518a,a87522a,a87523a,a87526a,a87529a,a87530a,a87531a,a87534a,a87537a,a87538a,a87541a,a87544a,a87545a,a87546a,a87550a,a87551a,a87554a,a87557a,a87558a,a87559a,a87562a,a87565a,a87566a,a87569a,a87572a,a87573a,a87574a,a87578a,a87579a,a87582a,a87585a,a87586a,a87587a,a87590a,a87593a,a87594a,a87597a,a87600a,a87601a,a87602a,a87606a,a87607a,a87610a,a87613a,a87614a,a87615a,a87618a,a87621a,a87622a,a87625a,a87628a,a87629a,a87630a,a87634a,a87635a,a87638a,a87641a,a87642a,a87643a,a87646a,a87649a,a87650a,a87653a,a87656a,a87657a,a87658a,a87662a,a87663a,a87666a,a87669a,a87670a,a87671a,a87674a,a87677a,a87678a,a87681a,a87684a,a87685a,a87686a,a87690a,a87691a,a87694a,a87697a,a87698a,a87699a,a87702a,a87705a,a87706a,a87709a,a87712a,a87713a,a87714a,a87718a,a87719a,a87722a,a87725a,a87726a,a87727a,a87730a,a87733a,a87734a,a87737a,a87740a,a87741a,a87742a,a87746a,a87747a,a87750a,a87753a,a87754a,a87755a,a87758a,a87761a,a87762a,a87765a,a87768a,a87769a,a87770a,a87774a,a87775a,a87778a,a87781a,a87782a,a87783a,a87786a,a87789a,a87790a,a87793a,a87796a,a87797a,a87798a,a87802a,a87803a,a87806a,a87809a,a87810a,a87811a,a87814a,a87817a,a87818a,a87821a,a87824a,a87825a,a87826a,a87830a,a87831a,a87834a,a87837a,a87838a,a87839a,a87842a,a87845a,a87846a,a87849a,a87852a,a87853a,a87854a,a87858a,a87859a,a87862a,a87865a,a87866a,a87867a,a87870a,a87873a,a87874a,a87877a,a87880a,a87881a,a87882a,a87886a,a87887a,a87890a,a87893a,a87894a,a87895a,a87898a,a87901a,a87902a,a87905a,a87908a,a87909a,a87910a,a87914a,a87915a,a87918a,a87921a,a87922a,a87923a,a87926a,a87929a,a87930a,a87933a,a87936a,a87937a,a87938a,a87942a,a87943a,a87946a,a87949a,a87950a,a87951a,a87954a,a87957a,a87958a,a87961a,a87964a,a87965a,a87966a,a87970a,a87971a,a87974a,a87977a,a87978a,a87979a,a87982a,a87985a,a87986a,a87989a,a87992a,a87993a,a87994a,a87998a,a87999a,a88002a,a88005a,a88006a,a88007a,a88010a,a88013a,a88014a,a88017a,a88020a,a88021a,a88022a,a88026a,a88027a,a88030a,a88033a,a88034a,a88035a,a88038a,a88041a,a88042a,a88045a,a88048a,a88049a,a88050a,a88054a,a88055a,a88058a,a88061a,a88062a,a88063a,a88066a,a88069a,a88070a,a88073a,a88076a,a88077a,a88078a,a88082a,a88083a,a88086a,a88089a,a88090a,a88091a,a88094a,a88097a,a88098a,a88101a,a88104a,a88105a,a88106a,a88110a,a88111a,a88114a,a88117a,a88118a,a88119a,a88122a,a88125a,a88126a,a88129a,a88132a,a88133a,a88134a,a88138a,a88139a,a88142a,a88145a,a88146a,a88147a,a88150a,a88153a,a88154a,a88157a,a88160a,a88161a,a88162a,a88166a,a88167a,a88170a,a88173a,a88174a,a88175a,a88178a,a88181a,a88182a,a88185a,a88188a,a88189a,a88190a,a88194a,a88195a,a88198a,a88201a,a88202a,a88203a,a88206a,a88209a,a88210a,a88213a,a88216a,a88217a,a88218a,a88222a,a88223a,a88226a,a88229a,a88230a,a88231a,a88234a,a88237a,a88238a,a88241a,a88244a,a88245a,a88246a,a88250a,a88251a,a88254a,a88257a,a88258a,a88259a,a88262a,a88265a,a88266a,a88269a,a88272a,a88273a,a88274a,a88278a,a88279a,a88282a,a88285a,a88286a,a88287a,a88290a,a88293a,a88294a,a88297a,a88300a,a88301a,a88302a,a88306a,a88307a,a88310a,a88313a,a88314a,a88315a,a88318a,a88321a,a88322a,a88325a,a88328a,a88329a,a88330a,a88334a,a88335a,a88338a,a88341a,a88342a,a88343a,a88346a,a88349a,a88350a,a88353a,a88356a,a88357a,a88358a,a88362a,a88363a,a88366a,a88369a,a88370a,a88371a,a88374a,a88377a,a88378a,a88381a,a88384a,a88385a,a88386a,a88390a,a88391a,a88394a,a88397a,a88398a,a88399a,a88402a,a88405a,a88406a,a88409a,a88412a,a88413a,a88414a,a88418a,a88419a,a88422a,a88425a,a88426a,a88427a,a88430a,a88433a,a88434a,a88437a,a88440a,a88441a,a88442a,a88446a,a88447a,a88450a,a88453a,a88454a,a88455a,a88458a,a88461a,a88462a,a88465a,a88468a,a88469a,a88470a,a88474a,a88475a,a88478a,a88481a,a88482a,a88483a,a88486a,a88489a,a88490a,a88493a,a88496a,a88497a,a88498a,a88502a,a88503a,a88506a,a88509a,a88510a,a88511a,a88514a,a88517a,a88518a,a88521a,a88524a,a88525a,a88526a,a88530a,a88531a,a88534a,a88537a,a88538a,a88539a,a88542a,a88545a,a88546a,a88549a,a88552a,a88553a,a88554a,a88558a,a88559a,a88562a,a88565a,a88566a,a88567a,a88570a,a88573a,a88574a,a88577a,a88580a,a88581a,a88582a,a88586a,a88587a,a88590a,a88593a,a88594a,a88595a,a88598a,a88601a,a88602a,a88605a,a88608a,a88609a,a88610a,a88614a,a88615a,a88618a,a88621a,a88622a,a88623a,a88626a,a88629a,a88630a,a88633a,a88636a,a88637a,a88638a,a88642a,a88643a,a88646a,a88649a,a88650a,a88651a,a88654a,a88657a,a88658a,a88661a,a88664a,a88665a,a88666a,a88670a,a88671a,a88674a,a88677a,a88678a,a88679a,a88682a,a88685a,a88686a,a88689a,a88692a,a88693a,a88694a,a88698a,a88699a,a88702a,a88705a,a88706a,a88707a,a88710a,a88713a,a88714a,a88717a,a88720a,a88721a,a88722a,a88726a,a88727a,a88730a,a88733a,a88734a,a88735a,a88738a,a88741a,a88742a,a88745a,a88748a,a88749a,a88750a,a88754a,a88755a,a88758a,a88761a,a88762a,a88763a,a88766a,a88769a,a88770a,a88773a,a88776a,a88777a,a88778a,a88782a,a88783a,a88786a,a88789a,a88790a,a88791a,a88794a,a88797a,a88798a,a88801a,a88804a,a88805a,a88806a,a88810a,a88811a,a88814a,a88817a,a88818a,a88819a,a88822a,a88825a,a88826a,a88829a,a88832a,a88833a,a88834a,a88838a,a88839a,a88842a,a88845a,a88846a,a88847a,a88850a,a88853a,a88854a,a88857a,a88860a,a88861a,a88862a,a88866a,a88867a,a88870a,a88873a,a88874a,a88875a,a88878a,a88881a,a88882a,a88885a,a88888a,a88889a,a88890a,a88894a,a88895a,a88898a,a88901a,a88902a,a88903a,a88906a,a88909a,a88910a,a88913a,a88916a,a88917a,a88918a,a88922a,a88923a,a88926a,a88929a,a88930a,a88931a,a88934a,a88937a,a88938a,a88941a,a88944a,a88945a,a88946a,a88950a,a88951a,a88954a,a88957a,a88958a,a88959a,a88962a,a88965a,a88966a,a88969a,a88972a,a88973a,a88974a,a88978a,a88979a,a88982a,a88985a,a88986a,a88987a,a88990a,a88993a,a88994a,a88997a,a89000a,a89001a,a89002a,a89006a,a89007a,a89010a,a89013a,a89014a,a89015a,a89018a,a89021a,a89022a,a89025a,a89028a,a89029a,a89030a,a89034a,a89035a,a89038a,a89041a,a89042a,a89043a,a89046a,a89049a,a89050a,a89053a,a89056a,a89057a,a89058a,a89062a,a89063a,a89066a,a89069a,a89070a,a89071a,a89074a,a89077a,a89078a,a89081a,a89084a,a89085a,a89086a,a89090a,a89091a,a89094a,a89097a,a89098a,a89099a,a89102a,a89105a,a89106a,a89109a,a89112a,a89113a,a89114a,a89118a,a89119a,a89122a,a89125a,a89126a,a89127a,a89130a,a89133a,a89134a,a89137a,a89140a,a89141a,a89142a,a89146a,a89147a,a89150a,a89153a,a89154a,a89155a,a89158a,a89161a,a89162a,a89165a,a89168a,a89169a,a89170a,a89174a,a89175a,a89178a,a89181a,a89182a,a89183a,a89186a,a89189a,a89190a,a89193a,a89196a,a89197a,a89198a,a89202a,a89203a,a89206a,a89209a,a89210a,a89211a,a89214a,a89217a,a89218a,a89221a,a89224a,a89225a,a89226a,a89230a,a89231a,a89234a,a89237a,a89238a,a89239a,a89242a,a89245a,a89246a,a89249a,a89252a,a89253a,a89254a,a89258a,a89259a,a89262a,a89265a,a89266a,a89267a,a89270a,a89273a,a89274a,a89277a,a89280a,a89281a,a89282a,a89286a,a89287a,a89290a,a89293a,a89294a,a89295a,a89298a,a89301a,a89302a,a89305a,a89308a,a89309a,a89310a,a89314a,a89315a,a89318a,a89321a,a89322a,a89323a,a89326a,a89329a,a89330a,a89333a,a89336a,a89337a,a89338a,a89342a,a89343a,a89346a,a89349a,a89350a,a89351a,a89354a,a89357a,a89358a,a89361a,a89364a,a89365a,a89366a,a89370a,a89371a,a89374a,a89377a,a89378a,a89379a,a89382a,a89385a,a89386a,a89389a,a89392a,a89393a,a89394a,a89398a,a89399a,a89402a,a89405a,a89406a,a89407a,a89410a,a89413a,a89414a,a89417a,a89420a,a89421a,a89422a,a89426a,a89427a,a89430a,a89433a,a89434a,a89435a,a89438a,a89441a,a89442a,a89445a,a89448a,a89449a,a89450a,a89454a,a89455a,a89458a,a89461a,a89462a,a89463a,a89466a,a89469a,a89470a,a89473a,a89476a,a89477a,a89478a,a89482a,a89483a,a89486a,a89489a,a89490a,a89491a,a89494a,a89497a,a89498a,a89501a,a89504a,a89505a,a89506a,a89510a,a89511a,a89514a,a89517a,a89518a,a89519a,a89522a,a89525a,a89526a,a89529a,a89532a,a89533a,a89534a,a89538a,a89539a,a89542a,a89545a,a89546a,a89547a,a89550a,a89553a,a89554a,a89557a,a89560a,a89561a,a89562a,a89566a,a89567a,a89570a,a89573a,a89574a,a89575a,a89578a,a89581a,a89582a,a89585a,a89588a,a89589a,a89590a,a89594a,a89595a,a89598a,a89601a,a89602a,a89603a,a89606a,a89609a,a89610a,a89613a,a89616a,a89617a,a89618a,a89622a,a89623a,a89626a,a89629a,a89630a,a89631a,a89634a,a89637a,a89638a,a89641a,a89644a,a89645a,a89646a,a89650a,a89651a,a89654a,a89657a,a89658a,a89659a,a89662a,a89665a,a89666a,a89669a,a89672a,a89673a,a89674a,a89678a,a89679a,a89682a,a89685a,a89686a,a89687a,a89690a,a89693a,a89694a,a89697a,a89700a,a89701a,a89702a,a89706a,a89707a,a89710a,a89713a,a89714a,a89715a,a89718a,a89721a,a89722a,a89725a,a89728a,a89729a,a89730a,a89734a,a89735a,a89738a,a89741a,a89742a,a89743a,a89746a,a89749a,a89750a,a89753a,a89756a,a89757a,a89758a,a89762a,a89763a,a89766a,a89769a,a89770a,a89771a,a89774a,a89777a,a89778a,a89781a,a89784a,a89785a,a89786a,a89790a,a89791a,a89794a,a89797a,a89798a,a89799a,a89802a,a89805a,a89806a,a89809a,a89812a,a89813a,a89814a,a89818a,a89819a,a89822a,a89825a,a89826a,a89827a,a89830a,a89833a,a89834a,a89837a,a89840a,a89841a,a89842a,a89846a,a89847a,a89850a,a89853a,a89854a,a89855a,a89858a,a89861a,a89862a,a89865a,a89868a,a89869a,a89870a,a89874a,a89875a,a89878a,a89881a,a89882a,a89883a,a89886a,a89889a,a89890a,a89893a,a89896a,a89897a,a89898a,a89902a,a89903a,a89906a,a89909a,a89910a,a89911a,a89914a,a89917a,a89918a,a89921a,a89924a,a89925a,a89926a,a89930a,a89931a,a89934a,a89937a,a89938a,a89939a,a89942a,a89945a,a89946a,a89949a,a89952a,a89953a,a89954a,a89958a,a89959a,a89962a,a89965a,a89966a,a89967a,a89970a,a89973a,a89974a,a89977a,a89980a,a89981a,a89982a,a89986a,a89987a,a89990a,a89993a,a89994a,a89995a,a89998a,a90001a,a90002a,a90005a,a90008a,a90009a,a90010a,a90014a,a90015a,a90018a,a90021a,a90022a,a90023a,a90026a,a90029a,a90030a,a90033a,a90036a,a90037a,a90038a,a90042a,a90043a,a90046a,a90049a,a90050a,a90051a,a90054a,a90057a,a90058a,a90061a,a90064a,a90065a,a90066a,a90070a,a90071a,a90074a,a90077a,a90078a,a90079a,a90082a,a90085a,a90086a,a90089a,a90092a,a90093a,a90094a,a90098a,a90099a,a90102a,a90105a,a90106a,a90107a,a90110a,a90113a,a90114a,a90117a,a90120a,a90121a,a90122a,a90126a,a90127a,a90130a,a90133a,a90134a,a90135a,a90138a,a90141a,a90142a,a90145a,a90148a,a90149a,a90150a,a90154a,a90155a,a90158a,a90161a,a90162a,a90163a,a90166a,a90169a,a90170a,a90173a,a90176a,a90177a,a90178a,a90182a,a90183a,a90186a,a90189a,a90190a,a90191a,a90194a,a90197a,a90198a,a90201a,a90204a,a90205a,a90206a,a90210a,a90211a,a90214a,a90217a,a90218a,a90219a,a90222a,a90225a,a90226a,a90229a,a90232a,a90233a,a90234a,a90238a,a90239a,a90242a,a90245a,a90246a,a90247a,a90250a,a90253a,a90254a,a90257a,a90260a,a90261a,a90262a,a90266a,a90267a,a90270a,a90273a,a90274a,a90275a,a90278a,a90281a,a90282a,a90285a,a90288a,a90289a,a90290a,a90294a,a90295a,a90298a,a90301a,a90302a,a90303a,a90306a,a90309a,a90310a,a90313a,a90316a,a90317a,a90318a,a90322a,a90323a,a90326a,a90329a,a90330a,a90331a,a90334a,a90337a,a90338a,a90341a,a90344a,a90345a,a90346a,a90350a,a90351a,a90354a,a90357a,a90358a,a90359a,a90362a,a90365a,a90366a,a90369a,a90372a,a90373a,a90374a,a90378a,a90379a,a90382a,a90385a,a90386a,a90387a,a90390a,a90393a,a90394a,a90397a,a90400a,a90401a,a90402a,a90406a,a90407a,a90410a,a90413a,a90414a,a90415a,a90418a,a90421a,a90422a,a90425a,a90428a,a90429a,a90430a,a90434a,a90435a,a90438a,a90441a,a90442a,a90443a,a90446a,a90449a,a90450a,a90453a,a90456a,a90457a,a90458a,a90462a,a90463a,a90466a,a90469a,a90470a,a90471a,a90474a,a90477a,a90478a,a90481a,a90484a,a90485a,a90486a,a90490a,a90491a,a90494a,a90497a,a90498a,a90499a,a90502a,a90505a,a90506a,a90509a,a90512a,a90513a,a90514a,a90518a,a90519a,a90522a,a90525a,a90526a,a90527a,a90530a,a90533a,a90534a,a90537a,a90540a,a90541a,a90542a,a90546a,a90547a,a90550a,a90553a,a90554a,a90555a,a90558a,a90561a,a90562a,a90565a,a90568a,a90569a,a90570a,a90574a,a90575a,a90578a,a90581a,a90582a,a90583a,a90586a,a90589a,a90590a,a90593a,a90596a,a90597a,a90598a,a90602a,a90603a,a90606a,a90609a,a90610a,a90611a,a90614a,a90617a,a90618a,a90621a,a90624a,a90625a,a90626a,a90630a,a90631a,a90634a,a90637a,a90638a,a90639a,a90642a,a90645a,a90646a,a90649a,a90652a,a90653a,a90654a,a90658a,a90659a,a90662a,a90665a,a90666a,a90667a,a90670a,a90673a,a90674a,a90677a,a90680a,a90681a,a90682a,a90686a,a90687a,a90690a,a90693a,a90694a,a90695a,a90698a,a90701a,a90702a,a90705a,a90708a,a90709a,a90710a,a90714a,a90715a,a90718a,a90721a,a90722a,a90723a,a90726a,a90729a,a90730a,a90733a,a90736a,a90737a,a90738a,a90742a,a90743a,a90746a,a90749a,a90750a,a90751a,a90754a,a90757a,a90758a,a90761a,a90764a,a90765a,a90766a,a90770a,a90771a,a90774a,a90777a,a90778a,a90779a,a90782a,a90785a,a90786a,a90789a,a90792a,a90793a,a90794a,a90798a,a90799a,a90802a,a90805a,a90806a,a90807a,a90810a,a90813a,a90814a,a90817a,a90820a,a90821a,a90822a,a90826a,a90827a,a90830a,a90833a,a90834a,a90835a,a90838a,a90841a,a90842a,a90845a,a90848a,a90849a,a90850a,a90854a,a90855a,a90858a,a90861a,a90862a,a90863a,a90866a,a90869a,a90870a,a90873a,a90876a,a90877a,a90878a,a90882a,a90883a,a90886a,a90889a,a90890a,a90891a,a90894a,a90897a,a90898a,a90901a,a90904a,a90905a,a90906a,a90910a,a90911a,a90914a,a90917a,a90918a,a90919a,a90922a,a90925a,a90926a,a90929a,a90932a,a90933a,a90934a,a90938a,a90939a,a90942a,a90945a,a90946a,a90947a,a90950a,a90953a,a90954a,a90957a,a90960a,a90961a,a90962a,a90966a,a90967a,a90970a,a90973a,a90974a,a90975a,a90978a,a90981a,a90982a,a90985a,a90988a,a90989a,a90990a,a90994a,a90995a,a90998a,a91001a,a91002a,a91003a,a91006a,a91009a,a91010a,a91013a,a91016a,a91017a,a91018a,a91022a,a91023a,a91026a,a91029a,a91030a,a91031a,a91034a,a91037a,a91038a,a91041a,a91044a,a91045a,a91046a,a91050a,a91051a,a91054a,a91057a,a91058a,a91059a,a91062a,a91065a,a91066a,a91069a,a91072a,a91073a,a91074a,a91078a,a91079a,a91082a,a91085a,a91086a,a91087a,a91090a,a91093a,a91094a,a91097a,a91100a,a91101a,a91102a,a91106a,a91107a,a91110a,a91113a,a91114a,a91115a,a91118a,a91121a,a91122a,a91125a,a91128a,a91129a,a91130a,a91134a,a91135a,a91138a,a91141a,a91142a,a91143a,a91146a,a91149a,a91150a,a91153a,a91156a,a91157a,a91158a,a91162a,a91163a,a91166a,a91169a,a91170a,a91171a,a91174a,a91177a,a91178a,a91181a,a91184a,a91185a,a91186a,a91190a,a91191a,a91194a,a91197a,a91198a,a91199a,a91202a,a91205a,a91206a,a91209a,a91212a,a91213a,a91214a,a91218a,a91219a,a91222a,a91225a,a91226a,a91227a,a91230a,a91233a,a91234a,a91237a,a91240a,a91241a,a91242a,a91246a,a91247a,a91250a,a91253a,a91254a,a91255a,a91258a,a91261a,a91262a,a91265a,a91268a,a91269a,a91270a,a91274a,a91275a,a91278a,a91281a,a91282a,a91283a,a91286a,a91289a,a91290a,a91293a,a91296a,a91297a,a91298a,a91302a,a91303a,a91306a,a91309a,a91310a,a91311a,a91314a,a91317a,a91318a,a91321a,a91324a,a91325a,a91326a,a91330a,a91331a,a91334a,a91337a,a91338a,a91339a,a91342a,a91345a,a91346a,a91349a,a91352a,a91353a,a91354a,a91358a,a91359a,a91362a,a91365a,a91366a,a91367a,a91370a,a91373a,a91374a,a91377a,a91380a,a91381a,a91382a,a91386a,a91387a,a91390a,a91393a,a91394a,a91395a,a91398a,a91401a,a91402a,a91405a,a91408a,a91409a,a91410a,a91414a,a91415a,a91418a,a91421a,a91422a,a91423a,a91426a,a91429a,a91430a,a91433a,a91436a,a91437a,a91438a,a91442a,a91443a,a91446a,a91449a,a91450a,a91451a,a91454a,a91457a,a91458a,a91461a,a91464a,a91465a,a91466a,a91470a,a91471a,a91474a,a91477a,a91478a,a91479a,a91482a,a91485a,a91486a,a91489a,a91492a,a91493a,a91494a,a91498a,a91499a,a91502a,a91505a,a91506a,a91507a,a91510a,a91513a,a91514a,a91517a,a91520a,a91521a,a91522a,a91526a,a91527a,a91530a,a91533a,a91534a,a91535a,a91538a,a91541a,a91542a,a91545a,a91548a,a91549a,a91550a,a91554a,a91555a,a91558a,a91561a,a91562a,a91563a,a91566a,a91569a,a91570a,a91573a,a91576a,a91577a,a91578a,a91582a,a91583a,a91586a,a91589a,a91590a,a91591a,a91594a,a91597a,a91598a,a91601a,a91604a,a91605a,a91606a,a91610a,a91611a,a91614a,a91617a,a91618a,a91619a,a91622a,a91625a,a91626a,a91629a,a91632a,a91633a,a91634a,a91638a,a91639a,a91642a,a91645a,a91646a,a91647a,a91650a,a91653a,a91654a,a91657a,a91660a,a91661a,a91662a,a91666a,a91667a,a91670a,a91673a,a91674a,a91675a,a91678a,a91681a,a91682a,a91685a,a91688a,a91689a,a91690a,a91694a,a91695a,a91698a,a91701a,a91702a,a91703a,a91706a,a91709a,a91710a,a91713a,a91716a,a91717a,a91718a,a91722a,a91723a,a91726a,a91729a,a91730a,a91731a,a91734a,a91737a,a91738a,a91741a,a91744a,a91745a,a91746a,a91750a,a91751a,a91754a,a91757a,a91758a,a91759a,a91762a,a91765a,a91766a,a91769a,a91772a,a91773a,a91774a,a91778a,a91779a,a91782a,a91785a,a91786a,a91787a,a91790a,a91793a,a91794a,a91797a,a91800a,a91801a,a91802a,a91806a,a91807a,a91810a,a91813a,a91814a,a91815a,a91818a,a91821a,a91822a,a91825a,a91828a,a91829a,a91830a,a91834a,a91835a,a91838a,a91841a,a91842a,a91843a,a91846a,a91849a,a91850a,a91853a,a91856a,a91857a,a91858a,a91862a,a91863a,a91866a,a91869a,a91870a,a91871a,a91874a,a91877a,a91878a,a91881a,a91884a,a91885a,a91886a,a91890a,a91891a,a91894a,a91897a,a91898a,a91899a,a91902a,a91905a,a91906a,a91909a,a91912a,a91913a,a91914a,a91918a,a91919a,a91922a,a91925a,a91926a,a91927a,a91930a,a91933a,a91934a,a91937a,a91940a,a91941a,a91942a,a91946a,a91947a,a91950a,a91953a,a91954a,a91955a,a91958a,a91961a,a91962a,a91965a,a91968a,a91969a,a91970a,a91974a,a91975a,a91978a,a91981a,a91982a,a91983a,a91986a,a91989a,a91990a,a91993a,a91996a,a91997a,a91998a,a92002a,a92003a,a92006a,a92009a,a92010a,a92011a,a92014a,a92017a,a92018a,a92021a,a92024a,a92025a,a92026a,a92030a,a92031a,a92034a,a92037a,a92038a,a92039a,a92042a,a92045a,a92046a,a92049a,a92052a,a92053a,a92054a,a92058a,a92059a,a92062a,a92065a,a92066a,a92067a,a92070a,a92073a,a92074a,a92077a,a92080a,a92081a,a92082a,a92086a,a92087a,a92090a,a92093a,a92094a,a92095a,a92098a,a92101a,a92102a,a92105a,a92108a,a92109a,a92110a,a92114a,a92115a,a92118a,a92121a,a92122a,a92123a,a92126a,a92129a,a92130a,a92133a,a92136a,a92137a,a92138a,a92142a,a92143a,a92146a,a92149a,a92150a,a92151a,a92154a,a92157a,a92158a,a92161a,a92164a,a92165a,a92166a,a92170a,a92171a,a92174a,a92177a,a92178a,a92179a,a92182a,a92185a,a92186a,a92189a,a92192a,a92193a,a92194a,a92198a,a92199a,a92202a,a92205a,a92206a,a92207a,a92210a,a92213a,a92214a,a92217a,a92220a,a92221a,a92222a,a92226a,a92227a,a92230a,a92233a,a92234a,a92235a,a92238a,a92241a,a92242a,a92245a,a92248a,a92249a,a92250a,a92254a,a92255a,a92258a,a92261a,a92262a,a92263a,a92266a,a92269a,a92270a,a92273a,a92276a,a92277a,a92278a,a92282a,a92283a,a92286a,a92289a,a92290a,a92291a,a92294a,a92297a,a92298a,a92301a,a92304a,a92305a,a92306a,a92310a,a92311a,a92314a,a92317a,a92318a,a92319a,a92322a,a92325a,a92326a,a92329a,a92332a,a92333a,a92334a,a92338a,a92339a,a92342a,a92345a,a92346a,a92347a,a92350a,a92353a,a92354a,a92357a,a92360a,a92361a,a92362a,a92366a,a92367a,a92370a,a92373a,a92374a,a92375a,a92378a,a92381a,a92382a,a92385a,a92388a,a92389a,a92390a,a92394a,a92395a,a92398a,a92401a,a92402a,a92403a,a92406a,a92409a,a92410a,a92413a,a92416a,a92417a,a92418a,a92422a,a92423a,a92426a,a92429a,a92430a,a92431a,a92434a,a92437a,a92438a,a92441a,a92444a,a92445a,a92446a,a92450a,a92451a,a92454a,a92457a,a92458a,a92459a,a92462a,a92465a,a92466a,a92469a,a92472a,a92473a,a92474a,a92478a,a92479a,a92482a,a92485a,a92486a,a92487a,a92490a,a92493a,a92494a,a92497a,a92500a,a92501a,a92502a,a92506a,a92507a,a92510a,a92513a,a92514a,a92515a,a92518a,a92521a,a92522a,a92525a,a92528a,a92529a,a92530a,a92534a,a92535a,a92538a,a92541a,a92542a,a92543a,a92546a,a92549a,a92550a,a92553a,a92556a,a92557a,a92558a,a92562a,a92563a,a92566a,a92569a,a92570a,a92571a,a92574a,a92577a,a92578a,a92581a,a92584a,a92585a,a92586a,a92590a,a92591a,a92594a,a92597a,a92598a,a92599a,a92602a,a92605a,a92606a,a92609a,a92612a,a92613a,a92614a,a92618a,a92619a,a92622a,a92625a,a92626a,a92627a,a92630a,a92633a,a92634a,a92637a,a92640a,a92641a,a92642a,a92646a,a92647a,a92650a,a92653a,a92654a,a92655a,a92658a,a92661a,a92662a,a92665a,a92668a,a92669a,a92670a,a92674a,a92675a,a92678a,a92681a,a92682a,a92683a,a92686a,a92689a,a92690a,a92693a,a92696a,a92697a,a92698a,a92702a,a92703a,a92706a,a92709a,a92710a,a92711a,a92714a,a92717a,a92718a,a92721a,a92724a,a92725a,a92726a,a92730a,a92731a,a92734a,a92737a,a92738a,a92739a,a92742a,a92745a,a92746a,a92749a,a92752a,a92753a,a92754a,a92758a,a92759a,a92762a,a92765a,a92766a,a92767a,a92770a,a92773a,a92774a,a92777a,a92780a,a92781a,a92782a,a92786a,a92787a,a92790a,a92793a,a92794a,a92795a,a92798a,a92801a,a92802a,a92805a,a92808a,a92809a,a92810a,a92814a,a92815a,a92818a,a92821a,a92822a,a92823a,a92826a,a92829a,a92830a,a92833a,a92836a,a92837a,a92838a,a92842a,a92843a,a92846a,a92849a,a92850a,a92851a,a92854a,a92857a,a92858a,a92861a,a92864a,a92865a,a92866a,a92870a,a92871a,a92874a,a92877a,a92878a,a92879a,a92882a,a92885a,a92886a,a92889a,a92892a,a92893a,a92894a,a92898a,a92899a,a92902a,a92905a,a92906a,a92907a,a92910a,a92913a,a92914a,a92917a,a92920a,a92921a,a92922a,a92926a,a92927a,a92930a,a92933a,a92934a,a92935a,a92938a,a92941a,a92942a,a92945a,a92948a,a92949a,a92950a,a92954a,a92955a,a92958a,a92961a,a92962a,a92963a,a92966a,a92969a,a92970a,a92973a,a92976a,a92977a,a92978a,a92982a,a92983a,a92986a,a92989a,a92990a,a92991a,a92994a,a92997a,a92998a,a93001a,a93004a,a93005a,a93006a,a93010a,a93011a,a93014a,a93017a,a93018a,a93019a,a93022a,a93025a,a93026a,a93029a,a93032a,a93033a,a93034a,a93038a,a93039a,a93042a,a93045a,a93046a,a93047a,a93050a,a93053a,a93054a,a93057a,a93060a,a93061a,a93062a,a93066a,a93067a,a93070a,a93073a,a93074a,a93075a,a93078a,a93081a,a93082a,a93085a,a93088a,a93089a,a93090a,a93094a,a93095a,a93098a,a93101a,a93102a,a93103a,a93106a,a93109a,a93110a,a93113a,a93116a,a93117a,a93118a,a93122a,a93123a,a93126a,a93129a,a93130a,a93131a,a93134a,a93137a,a93138a,a93141a,a93144a,a93145a,a93146a,a93150a,a93151a,a93154a,a93157a,a93158a,a93159a,a93162a,a93165a,a93166a,a93169a,a93172a,a93173a,a93174a,a93178a,a93179a,a93182a,a93185a,a93186a,a93187a,a93190a,a93193a,a93194a,a93197a,a93200a,a93201a,a93202a,a93206a,a93207a,a93210a,a93213a,a93214a,a93215a,a93218a,a93221a,a93222a,a93225a,a93228a,a93229a,a93230a,a93234a,a93235a,a93238a,a93241a,a93242a,a93243a,a93246a,a93249a,a93250a,a93253a,a93256a,a93257a,a93258a,a93262a,a93263a,a93266a,a93269a,a93270a,a93271a,a93274a,a93277a,a93278a,a93281a,a93284a,a93285a,a93286a,a93290a,a93291a,a93294a,a93297a,a93298a,a93299a,a93302a,a93305a,a93306a,a93309a,a93312a,a93313a,a93314a,a93318a,a93319a,a93322a,a93325a,a93326a,a93327a,a93330a,a93333a,a93334a,a93337a,a93340a,a93341a,a93342a,a93346a,a93347a,a93350a,a93353a,a93354a,a93355a,a93358a,a93361a,a93362a,a93365a,a93368a,a93369a,a93370a,a93374a,a93375a,a93378a,a93381a,a93382a,a93383a,a93386a,a93389a,a93390a,a93393a,a93396a,a93397a,a93398a,a93402a,a93403a,a93406a,a93409a,a93410a,a93411a,a93414a,a93417a,a93418a,a93421a,a93424a,a93425a,a93426a,a93430a,a93431a,a93434a,a93437a,a93438a,a93439a,a93442a,a93445a,a93446a,a93449a,a93452a,a93453a,a93454a,a93458a,a93459a,a93462a,a93465a,a93466a,a93467a,a93470a,a93473a,a93474a,a93477a,a93480a,a93481a,a93482a,a93486a,a93487a,a93490a,a93493a,a93494a,a93495a,a93498a,a93501a,a93502a,a93505a,a93508a,a93509a,a93510a,a93514a,a93515a,a93518a,a93521a,a93522a,a93523a,a93526a,a93529a,a93530a,a93533a,a93536a,a93537a,a93538a,a93542a,a93543a,a93546a,a93549a,a93550a,a93551a,a93554a,a93557a,a93558a,a93561a,a93564a,a93565a,a93566a,a93570a,a93571a,a93574a,a93577a,a93578a,a93579a,a93582a,a93585a,a93586a,a93589a,a93592a,a93593a,a93594a,a93598a,a93599a,a93602a,a93605a,a93606a,a93607a,a93610a,a93613a,a93614a,a93617a,a93620a,a93621a,a93622a,a93626a,a93627a,a93630a,a93633a,a93634a,a93635a,a93638a,a93641a,a93642a,a93645a,a93648a,a93649a,a93650a,a93654a,a93655a,a93658a,a93661a,a93662a,a93663a,a93666a,a93669a,a93670a,a93673a,a93676a,a93677a,a93678a,a93682a,a93683a,a93686a,a93689a,a93690a,a93691a,a93694a,a93697a,a93698a,a93701a,a93704a,a93705a,a93706a,a93710a,a93711a,a93714a,a93717a,a93718a,a93719a,a93722a,a93725a,a93726a,a93729a,a93732a,a93733a,a93734a,a93738a,a93739a,a93742a,a93745a,a93746a,a93747a,a93750a,a93753a,a93754a,a93757a,a93760a,a93761a,a93762a,a93766a,a93767a,a93770a,a93773a,a93774a,a93775a,a93778a,a93781a,a93782a,a93785a,a93788a,a93789a,a93790a,a93794a,a93795a,a93798a,a93801a,a93802a,a93803a,a93806a,a93809a,a93810a,a93813a,a93816a,a93817a,a93818a,a93822a,a93823a,a93826a,a93829a,a93830a,a93831a,a93834a,a93837a,a93838a,a93841a,a93844a,a93845a,a93846a,a93850a,a93851a,a93854a,a93857a,a93858a,a93859a,a93862a,a93865a,a93866a,a93869a,a93872a,a93873a,a93874a,a93878a,a93879a,a93882a,a93885a,a93886a,a93887a,a93890a,a93893a,a93894a,a93897a,a93900a,a93901a,a93902a,a93906a,a93907a,a93910a,a93913a,a93914a,a93915a,a93918a,a93921a,a93922a,a93925a,a93928a,a93929a,a93930a,a93934a,a93935a,a93938a,a93941a,a93942a,a93943a,a93946a,a93949a,a93950a,a93953a,a93956a,a93957a,a93958a,a93962a,a93963a,a93966a,a93969a,a93970a,a93971a,a93974a,a93977a,a93978a,a93981a,a93984a,a93985a,a93986a,a93990a,a93991a,a93994a,a93997a,a93998a,a93999a,a94002a,a94005a,a94006a,a94009a,a94012a,a94013a,a94014a,a94018a,a94019a,a94022a,a94025a,a94026a,a94027a,a94030a,a94033a,a94034a,a94037a,a94040a,a94041a,a94042a,a94046a,a94047a,a94050a,a94053a,a94054a,a94055a,a94058a,a94061a,a94062a,a94065a,a94068a,a94069a,a94070a,a94074a,a94075a,a94078a,a94081a,a94082a,a94083a,a94086a,a94089a,a94090a,a94093a,a94096a,a94097a,a94098a,a94102a,a94103a,a94106a,a94109a,a94110a,a94111a,a94114a,a94117a,a94118a,a94121a,a94124a,a94125a,a94126a,a94130a,a94131a,a94134a,a94137a,a94138a,a94139a,a94142a,a94145a,a94146a,a94149a,a94152a,a94153a,a94154a,a94158a,a94159a,a94162a,a94165a,a94166a,a94167a,a94170a,a94173a,a94174a,a94177a,a94180a,a94181a,a94182a,a94186a,a94187a,a94190a,a94193a,a94194a,a94195a,a94198a,a94201a,a94202a,a94205a,a94208a,a94209a,a94210a,a94214a,a94215a,a94218a,a94221a,a94222a,a94223a,a94226a,a94229a,a94230a,a94233a,a94236a,a94237a,a94238a,a94242a,a94243a,a94246a,a94249a,a94250a,a94251a,a94254a,a94257a,a94258a,a94261a,a94264a,a94265a,a94266a,a94270a,a94271a,a94274a,a94277a,a94278a,a94279a,a94282a,a94285a,a94286a,a94289a,a94292a,a94293a,a94294a,a94298a,a94299a,a94302a,a94305a,a94306a,a94307a,a94310a,a94313a,a94314a,a94317a,a94320a,a94321a,a94322a,a94326a,a94327a,a94330a,a94333a,a94334a,a94335a,a94338a,a94341a,a94342a,a94345a,a94348a,a94349a,a94350a,a94354a,a94355a,a94358a,a94361a,a94362a,a94363a,a94366a,a94369a,a94370a,a94373a,a94376a,a94377a,a94378a,a94382a,a94383a,a94386a,a94389a,a94390a,a94391a,a94394a,a94397a,a94398a,a94401a,a94404a,a94405a,a94406a,a94410a,a94411a,a94414a,a94417a,a94418a,a94419a,a94422a,a94425a,a94426a,a94429a,a94432a,a94433a,a94434a,a94438a,a94439a,a94442a,a94445a,a94446a,a94447a,a94450a,a94453a,a94454a,a94457a,a94460a,a94461a,a94462a,a94466a,a94467a,a94470a,a94473a,a94474a,a94475a,a94478a,a94481a,a94482a,a94485a,a94488a,a94489a,a94490a,a94494a,a94495a,a94498a,a94501a,a94502a,a94503a,a94506a,a94509a,a94510a,a94513a,a94516a,a94517a,a94518a,a94522a,a94523a,a94526a,a94529a,a94530a,a94531a,a94534a,a94537a,a94538a,a94541a,a94544a,a94545a,a94546a,a94550a,a94551a,a94554a,a94557a,a94558a,a94559a,a94562a,a94565a,a94566a,a94569a,a94572a,a94573a,a94574a,a94578a,a94579a,a94582a,a94585a,a94586a,a94587a,a94590a,a94593a,a94594a,a94597a,a94600a,a94601a,a94602a,a94606a,a94607a,a94610a,a94613a,a94614a,a94615a,a94618a,a94621a,a94622a,a94625a,a94628a,a94629a,a94630a,a94634a,a94635a,a94638a,a94641a,a94642a,a94643a,a94646a,a94649a,a94650a,a94653a,a94656a,a94657a,a94658a,a94662a,a94663a,a94666a,a94669a,a94670a,a94671a,a94674a,a94677a,a94678a,a94681a,a94684a,a94685a,a94686a,a94690a,a94691a,a94694a,a94697a,a94698a,a94699a,a94702a,a94705a,a94706a,a94709a,a94712a,a94713a,a94714a,a94718a,a94719a,a94722a,a94725a,a94726a,a94727a,a94730a,a94733a,a94734a,a94737a,a94740a,a94741a,a94742a,a94746a,a94747a,a94750a,a94753a,a94754a,a94755a,a94758a,a94761a,a94762a,a94765a,a94768a,a94769a,a94770a,a94774a,a94775a,a94778a,a94781a,a94782a,a94783a,a94786a,a94789a,a94790a,a94793a,a94796a,a94797a,a94798a,a94802a,a94803a,a94806a,a94809a,a94810a,a94811a,a94814a,a94817a,a94818a,a94821a,a94824a,a94825a,a94826a,a94830a,a94831a,a94834a,a94837a,a94838a,a94839a,a94842a,a94845a,a94846a,a94849a,a94852a,a94853a,a94854a,a94858a,a94859a,a94862a,a94865a,a94866a,a94867a,a94870a,a94873a,a94874a,a94877a,a94880a,a94881a,a94882a,a94886a,a94887a,a94890a,a94893a,a94894a,a94895a,a94898a,a94901a,a94902a,a94905a,a94908a,a94909a,a94910a,a94914a,a94915a,a94918a,a94921a,a94922a,a94923a,a94926a,a94929a,a94930a,a94933a,a94936a,a94937a,a94938a,a94942a,a94943a,a94946a,a94949a,a94950a,a94951a,a94954a,a94957a,a94958a,a94961a,a94964a,a94965a,a94966a,a94970a,a94971a,a94974a,a94977a,a94978a,a94979a,a94982a,a94985a,a94986a,a94989a,a94992a,a94993a,a94994a,a94998a,a94999a,a95002a,a95005a,a95006a,a95007a,a95010a,a95013a,a95014a,a95017a,a95020a,a95021a,a95022a,a95026a,a95027a,a95030a,a95033a,a95034a,a95035a,a95038a,a95041a,a95042a,a95045a,a95048a,a95049a,a95050a,a95054a,a95055a,a95058a,a95061a,a95062a,a95063a,a95066a,a95069a,a95070a,a95073a,a95076a,a95077a,a95078a,a95082a,a95083a,a95086a,a95089a,a95090a,a95091a,a95094a,a95097a,a95098a,a95101a,a95104a,a95105a,a95106a,a95110a,a95111a,a95114a,a95117a,a95118a,a95119a,a95122a,a95125a,a95126a,a95129a,a95132a,a95133a,a95134a,a95138a,a95139a,a95142a,a95145a,a95146a,a95147a,a95150a,a95153a,a95154a,a95157a,a95160a,a95161a,a95162a,a95166a,a95167a,a95170a,a95173a,a95174a,a95175a,a95178a,a95181a,a95182a,a95185a,a95188a,a95189a,a95190a,a95194a,a95195a,a95198a,a95201a,a95202a,a95203a,a95206a,a95209a,a95210a,a95213a,a95216a,a95217a,a95218a,a95222a,a95223a,a95226a,a95229a,a95230a,a95231a,a95234a,a95237a,a95238a,a95241a,a95244a,a95245a,a95246a,a95250a,a95251a,a95254a,a95257a,a95258a,a95259a,a95262a,a95265a,a95266a,a95269a,a95272a,a95273a,a95274a,a95278a,a95279a,a95282a,a95285a,a95286a,a95287a,a95290a,a95293a,a95294a,a95297a,a95300a,a95301a,a95302a,a95306a,a95307a,a95310a,a95313a,a95314a,a95315a,a95318a,a95321a,a95322a,a95325a,a95328a,a95329a,a95330a,a95334a,a95335a,a95338a,a95341a,a95342a,a95343a,a95346a,a95349a,a95350a,a95353a,a95356a,a95357a,a95358a,a95362a,a95363a,a95366a,a95369a,a95370a,a95371a,a95374a,a95377a,a95378a,a95381a,a95384a,a95385a,a95386a,a95390a,a95391a,a95394a,a95397a,a95398a,a95399a,a95402a,a95405a,a95406a,a95409a,a95412a,a95413a,a95414a,a95418a,a95419a,a95422a,a95425a,a95426a,a95427a,a95430a,a95433a,a95434a,a95437a,a95440a,a95441a,a95442a,a95446a,a95447a,a95450a,a95453a,a95454a,a95455a,a95458a,a95461a,a95462a,a95465a,a95468a,a95469a,a95470a,a95474a,a95475a,a95478a,a95481a,a95482a,a95483a,a95486a,a95489a,a95490a,a95493a,a95496a,a95497a,a95498a,a95502a,a95503a,a95506a,a95509a,a95510a,a95511a,a95514a,a95517a,a95518a,a95521a,a95524a,a95525a,a95526a,a95530a,a95531a,a95534a,a95537a,a95538a,a95539a,a95542a,a95545a,a95546a,a95549a,a95552a,a95553a,a95554a,a95558a,a95559a,a95562a,a95565a,a95566a,a95567a,a95570a,a95573a,a95574a,a95577a,a95580a,a95581a,a95582a,a95586a,a95587a,a95590a,a95593a,a95594a,a95595a,a95598a,a95601a,a95602a,a95605a,a95608a,a95609a,a95610a,a95614a,a95615a,a95618a,a95621a,a95622a,a95623a,a95626a,a95629a,a95630a,a95633a,a95636a,a95637a,a95638a,a95642a,a95643a,a95646a,a95649a,a95650a,a95651a,a95654a,a95657a,a95658a,a95661a,a95664a,a95665a,a95666a,a95670a,a95671a,a95674a,a95677a,a95678a,a95679a,a95682a,a95685a,a95686a,a95689a,a95692a,a95693a,a95694a,a95698a,a95699a,a95702a,a95705a,a95706a,a95707a,a95710a,a95713a,a95714a,a95717a,a95720a,a95721a,a95722a,a95726a,a95727a,a95730a,a95733a,a95734a,a95735a,a95738a,a95741a,a95742a,a95745a,a95748a,a95749a,a95750a,a95754a,a95755a,a95758a,a95761a,a95762a,a95763a,a95766a,a95769a,a95770a,a95773a,a95776a,a95777a,a95778a,a95782a,a95783a,a95786a,a95789a,a95790a,a95791a,a95794a,a95797a,a95798a,a95801a,a95804a,a95805a,a95806a,a95810a,a95811a,a95814a,a95817a,a95818a,a95819a,a95822a,a95825a,a95826a,a95829a,a95832a,a95833a,a95834a,a95838a,a95839a,a95842a,a95845a,a95846a,a95847a,a95850a,a95853a,a95854a,a95857a,a95860a,a95861a,a95862a,a95866a,a95867a,a95870a,a95873a,a95874a,a95875a,a95878a,a95881a,a95882a,a95885a,a95888a,a95889a,a95890a,a95894a,a95895a,a95898a,a95901a,a95902a,a95903a,a95906a,a95909a,a95910a,a95913a,a95916a,a95917a,a95918a,a95922a,a95923a,a95926a,a95929a,a95930a,a95931a,a95934a,a95937a,a95938a,a95941a,a95944a,a95945a,a95946a,a95950a,a95951a,a95954a,a95957a,a95958a,a95959a,a95962a,a95965a,a95966a,a95969a,a95972a,a95973a,a95974a,a95978a,a95979a,a95982a,a95985a,a95986a,a95987a,a95990a,a95993a,a95994a,a95997a,a96000a,a96001a,a96002a,a96006a,a96007a,a96010a,a96013a,a96014a,a96015a,a96018a,a96021a,a96022a,a96025a,a96028a,a96029a,a96030a,a96034a,a96035a,a96038a,a96041a,a96042a,a96043a,a96046a,a96049a,a96050a,a96053a,a96056a,a96057a,a96058a,a96062a,a96063a,a96066a,a96069a,a96070a,a96071a,a96074a,a96077a,a96078a,a96081a,a96084a,a96085a,a96086a,a96090a,a96091a,a96094a,a96097a,a96098a,a96099a,a96102a,a96105a,a96106a,a96109a,a96112a,a96113a,a96114a,a96118a,a96119a,a96122a,a96125a,a96126a,a96127a,a96130a,a96133a,a96134a,a96137a,a96140a,a96141a,a96142a,a96146a,a96147a,a96150a,a96153a,a96154a,a96155a,a96158a,a96161a,a96162a,a96165a,a96168a,a96169a,a96170a,a96174a,a96175a,a96178a,a96181a,a96182a,a96183a,a96186a,a96189a,a96190a,a96193a,a96196a,a96197a,a96198a,a96202a,a96203a,a96206a,a96209a,a96210a,a96211a,a96214a,a96217a,a96218a,a96221a,a96224a,a96225a,a96226a,a96230a,a96231a,a96234a,a96237a,a96238a,a96239a,a96242a,a96245a,a96246a,a96249a,a96252a,a96253a,a96254a,a96258a,a96259a,a96262a,a96265a,a96266a,a96267a,a96270a,a96273a,a96274a,a96277a,a96280a,a96281a,a96282a,a96286a,a96287a,a96290a,a96293a,a96294a,a96295a,a96298a,a96301a,a96302a,a96305a,a96308a,a96309a,a96310a,a96314a,a96315a,a96318a,a96321a,a96322a,a96323a,a96326a,a96329a,a96330a,a96333a,a96336a,a96337a,a96338a,a96342a,a96343a,a96346a,a96349a,a96350a,a96351a,a96354a,a96357a,a96358a,a96361a,a96364a,a96365a,a96366a,a96370a,a96371a,a96374a,a96377a,a96378a,a96379a,a96382a,a96385a,a96386a,a96389a,a96392a,a96393a,a96394a,a96398a,a96399a,a96402a,a96405a,a96406a,a96407a,a96410a,a96413a,a96414a,a96417a,a96420a,a96421a,a96422a,a96426a,a96427a,a96430a,a96433a,a96434a,a96435a,a96438a,a96441a,a96442a,a96445a,a96448a,a96449a,a96450a,a96454a,a96455a,a96458a,a96461a,a96462a,a96463a,a96466a,a96469a,a96470a,a96473a,a96476a,a96477a,a96478a,a96482a,a96483a,a96486a,a96489a,a96490a,a96491a,a96494a,a96497a,a96498a,a96501a,a96504a,a96505a,a96506a,a96510a,a96511a,a96514a,a96517a,a96518a,a96519a,a96522a,a96525a,a96526a,a96529a,a96532a,a96533a,a96534a,a96538a,a96539a,a96542a,a96545a,a96546a,a96547a,a96550a,a96553a,a96554a,a96557a,a96560a,a96561a,a96562a,a96566a,a96567a,a96570a,a96573a,a96574a,a96575a,a96578a,a96581a,a96582a,a96585a,a96588a,a96589a,a96590a,a96594a,a96595a,a96598a,a96601a,a96602a,a96603a,a96606a,a96609a,a96610a,a96613a,a96616a,a96617a,a96618a,a96622a,a96623a,a96626a,a96629a,a96630a,a96631a,a96634a,a96637a,a96638a,a96641a,a96644a,a96645a,a96646a,a96650a,a96651a,a96654a,a96657a,a96658a,a96659a,a96662a,a96665a,a96666a,a96669a,a96672a,a96673a,a96674a,a96678a,a96679a,a96682a,a96685a,a96686a,a96687a,a96690a,a96693a,a96694a,a96697a,a96700a,a96701a,a96702a,a96706a,a96707a,a96710a,a96713a,a96714a,a96715a,a96718a,a96721a,a96722a,a96725a,a96728a,a96729a,a96730a,a96734a,a96735a,a96738a,a96741a,a96742a,a96743a,a96746a,a96749a,a96750a,a96753a,a96756a,a96757a,a96758a,a96762a,a96763a,a96766a,a96769a,a96770a,a96771a,a96774a,a96777a,a96778a,a96781a,a96784a,a96785a,a96786a,a96790a,a96791a,a96794a,a96797a,a96798a,a96799a,a96802a,a96805a,a96806a,a96809a,a96812a,a96813a,a96814a,a96818a,a96819a,a96822a,a96825a,a96826a,a96827a,a96830a,a96833a,a96834a,a96837a,a96840a,a96841a,a96842a,a96846a,a96847a,a96850a,a96853a,a96854a,a96855a,a96858a,a96861a,a96862a,a96865a,a96868a,a96869a,a96870a,a96874a,a96875a,a96878a,a96881a,a96882a,a96883a,a96886a,a96889a,a96890a,a96893a,a96896a,a96897a,a96898a,a96902a,a96903a,a96906a,a96909a,a96910a,a96911a,a96914a,a96917a,a96918a,a96921a,a96924a,a96925a,a96926a,a96930a,a96931a,a96934a,a96937a,a96938a,a96939a,a96942a,a96945a,a96946a,a96949a,a96952a,a96953a,a96954a,a96958a,a96959a,a96962a,a96965a,a96966a,a96967a,a96970a,a96973a,a96974a,a96977a,a96980a,a96981a,a96982a,a96986a,a96987a,a96990a,a96993a,a96994a,a96995a,a96998a,a97001a,a97002a,a97005a,a97008a,a97009a,a97010a,a97014a,a97015a,a97018a,a97021a,a97022a,a97023a,a97026a,a97029a,a97030a,a97033a,a97036a,a97037a,a97038a,a97042a,a97043a,a97046a,a97049a,a97050a,a97051a,a97054a,a97057a,a97058a,a97061a,a97064a,a97065a,a97066a,a97070a,a97071a,a97074a,a97077a,a97078a,a97079a,a97082a,a97085a,a97086a,a97089a,a97092a,a97093a,a97094a,a97098a,a97099a,a97102a,a97105a,a97106a,a97107a,a97110a,a97113a,a97114a,a97117a,a97120a,a97121a,a97122a,a97126a,a97127a,a97130a,a97133a,a97134a,a97135a,a97138a,a97141a,a97142a,a97145a,a97148a,a97149a,a97150a,a97154a,a97155a,a97158a,a97161a,a97162a,a97163a,a97166a,a97169a,a97170a,a97173a,a97176a,a97177a,a97178a,a97182a,a97183a,a97186a,a97189a,a97190a,a97191a,a97194a,a97197a,a97198a,a97201a,a97204a,a97205a,a97206a,a97210a,a97211a,a97214a,a97217a,a97218a,a97219a,a97222a,a97225a,a97226a,a97229a,a97232a,a97233a,a97234a,a97238a,a97239a,a97242a,a97245a,a97246a,a97247a,a97250a,a97253a,a97254a,a97257a,a97260a,a97261a,a97262a,a97266a,a97267a,a97270a,a97273a,a97274a,a97275a,a97278a,a97281a,a97282a,a97285a,a97288a,a97289a,a97290a,a97294a,a97295a,a97298a,a97301a,a97302a,a97303a,a97306a,a97309a,a97310a,a97313a,a97316a,a97317a,a97318a,a97322a,a97323a,a97326a,a97329a,a97330a,a97331a,a97334a,a97337a,a97338a,a97341a,a97344a,a97345a,a97346a,a97350a,a97351a,a97354a,a97357a,a97358a,a97359a,a97362a,a97365a,a97366a,a97369a,a97372a,a97373a,a97374a,a97378a,a97379a,a97382a,a97385a,a97386a,a97387a,a97390a,a97393a,a97394a,a97397a,a97400a,a97401a,a97402a,a97406a,a97407a,a97410a,a97413a,a97414a,a97415a,a97418a,a97421a,a97422a,a97425a,a97428a,a97429a,a97430a,a97434a,a97435a,a97438a,a97441a,a97442a,a97443a,a97446a,a97449a,a97450a,a97453a,a97456a,a97457a,a97458a,a97462a,a97463a,a97466a,a97469a,a97470a,a97471a,a97474a,a97477a,a97478a,a97481a,a97484a,a97485a,a97486a,a97490a,a97491a,a97494a,a97497a,a97498a,a97499a,a97502a,a97505a,a97506a,a97509a,a97512a,a97513a,a97514a,a97518a,a97519a,a97522a,a97525a,a97526a,a97527a,a97530a,a97533a,a97534a,a97537a,a97540a,a97541a,a97542a,a97545a,a97548a,a97549a,a97552a,a97555a,a97556a,a97557a,a97560a,a97563a,a97564a,a97567a,a97570a,a97571a,a97572a,a97575a,a97578a,a97579a,a97582a,a97585a,a97586a,a97587a,a97590a,a97593a,a97594a,a97597a,a97600a,a97601a,a97602a,a97605a,a97608a,a97609a,a97612a,a97615a,a97616a,a97617a,a97620a,a97623a,a97624a,a97627a,a97630a,a97631a,a97632a,a97635a,a97638a,a97639a,a97642a,a97645a,a97646a,a97647a,a97650a,a97653a,a97654a,a97657a,a97660a,a97661a,a97662a,a97665a,a97668a,a97669a,a97672a,a97675a,a97676a,a97677a,a97680a,a97683a,a97684a,a97687a,a97690a,a97691a,a97692a,a97695a,a97698a,a97699a,a97702a,a97705a,a97706a,a97707a,a97710a,a97713a,a97714a,a97717a,a97720a,a97721a,a97722a,a97725a,a97728a,a97729a,a97732a,a97735a,a97736a,a97737a,a97740a,a97743a,a97744a,a97747a,a97750a,a97751a,a97752a,a97755a,a97758a,a97759a,a97762a,a97765a,a97766a,a97767a,a97770a,a97773a,a97774a,a97777a,a97780a,a97781a,a97782a,a97785a,a97788a,a97789a,a97792a,a97795a,a97796a,a97797a,a97800a,a97803a,a97804a,a97807a,a97810a,a97811a,a97812a,a97815a,a97818a,a97819a,a97822a,a97825a,a97826a,a97827a,a97830a,a97833a,a97834a,a97837a,a97840a,a97841a,a97842a,a97845a,a97848a,a97849a,a97852a,a97855a,a97856a,a97857a,a97860a,a97863a,a97864a,a97867a,a97870a,a97871a,a97872a,a97875a,a97878a,a97879a,a97882a,a97885a,a97886a,a97887a,a97890a,a97893a,a97894a,a97897a,a97900a,a97901a,a97902a,a97905a,a97908a,a97909a,a97912a,a97915a,a97916a,a97917a,a97920a,a97923a,a97924a,a97927a,a97930a,a97931a,a97932a,a97935a,a97938a,a97939a,a97942a,a97945a,a97946a,a97947a,a97950a,a97953a,a97954a,a97957a,a97960a,a97961a,a97962a,a97965a,a97968a,a97969a,a97972a,a97975a,a97976a,a97977a,a97980a,a97983a,a97984a,a97987a,a97990a,a97991a,a97992a,a97995a,a97998a,a97999a,a98002a,a98005a,a98006a,a98007a,a98010a,a98013a,a98014a,a98017a,a98020a,a98021a,a98022a,a98025a,a98028a,a98029a,a98032a,a98035a,a98036a,a98037a,a98040a,a98043a,a98044a,a98047a,a98050a,a98051a,a98052a,a98055a,a98058a,a98059a,a98062a,a98065a,a98066a,a98067a,a98070a,a98073a,a98074a,a98077a,a98080a,a98081a,a98082a,a98085a,a98088a,a98089a,a98092a,a98095a,a98096a,a98097a,a98100a,a98103a,a98104a,a98107a,a98110a,a98111a,a98112a,a98115a,a98118a,a98119a,a98122a,a98125a,a98126a,a98127a,a98130a,a98133a,a98134a,a98137a,a98140a,a98141a,a98142a,a98145a,a98148a,a98149a,a98152a,a98155a,a98156a,a98157a,a98160a,a98163a,a98164a,a98167a,a98170a,a98171a,a98172a,a98175a,a98178a,a98179a,a98182a,a98185a,a98186a,a98187a,a98190a,a98193a,a98194a,a98197a,a98200a,a98201a,a98202a,a98205a,a98208a,a98209a,a98212a,a98215a,a98216a,a98217a,a98220a,a98223a,a98224a,a98227a,a98230a,a98231a,a98232a,a98235a,a98238a,a98239a,a98242a,a98245a,a98246a,a98247a,a98250a,a98253a,a98254a,a98257a,a98260a,a98261a,a98262a,a98265a,a98268a,a98269a,a98272a,a98275a,a98276a,a98277a,a98280a,a98283a,a98284a,a98287a,a98290a,a98291a,a98292a,a98295a,a98298a,a98299a,a98302a,a98305a,a98306a,a98307a,a98310a,a98313a,a98314a,a98317a,a98320a,a98321a,a98322a,a98325a,a98328a,a98329a,a98332a,a98335a,a98336a,a98337a,a98340a,a98343a,a98344a,a98347a,a98350a,a98351a,a98352a,a98355a,a98358a,a98359a,a98362a,a98365a,a98366a,a98367a,a98370a,a98373a,a98374a,a98377a,a98380a,a98381a,a98382a,a98385a,a98388a,a98389a,a98392a,a98395a,a98396a,a98397a,a98400a,a98403a,a98404a,a98407a,a98410a,a98411a,a98412a,a98415a,a98418a,a98419a,a98422a,a98425a,a98426a,a98427a,a98430a,a98433a,a98434a,a98437a,a98440a,a98441a,a98442a,a98445a,a98448a,a98449a,a98452a,a98455a,a98456a,a98457a,a98460a,a98463a,a98464a,a98467a,a98470a,a98471a,a98472a,a98475a,a98478a,a98479a,a98482a,a98485a,a98486a,a98487a,a98490a,a98493a,a98494a,a98497a,a98500a,a98501a,a98502a,a98505a,a98508a,a98509a,a98512a,a98515a,a98516a,a98517a,a98520a,a98523a,a98524a,a98527a,a98530a,a98531a,a98532a,a98535a,a98538a,a98539a,a98542a,a98545a,a98546a,a98547a,a98550a,a98553a,a98554a,a98557a,a98560a,a98561a,a98562a,a98565a,a98568a,a98569a,a98572a,a98575a,a98576a,a98577a,a98580a,a98583a,a98584a,a98587a,a98590a,a98591a,a98592a,a98595a,a98598a,a98599a,a98602a,a98605a,a98606a,a98607a,a98610a,a98613a,a98614a,a98617a,a98620a,a98621a,a98622a,a98625a,a98628a,a98629a,a98632a,a98635a,a98636a,a98637a,a98640a,a98643a,a98644a,a98647a,a98650a,a98651a,a98652a,a98655a,a98658a,a98659a,a98662a,a98665a,a98666a,a98667a,a98670a,a98673a,a98674a,a98677a,a98680a,a98681a,a98682a,a98685a,a98688a,a98689a,a98692a,a98695a,a98696a,a98697a,a98700a,a98703a,a98704a,a98707a,a98710a,a98711a,a98712a,a98715a,a98718a,a98719a,a98722a,a98725a,a98726a,a98727a,a98730a,a98733a,a98734a,a98737a,a98740a,a98741a,a98742a,a98745a,a98748a,a98749a,a98752a,a98755a,a98756a,a98757a,a98760a,a98763a,a98764a,a98767a,a98770a,a98771a,a98772a,a98775a,a98778a,a98779a,a98782a,a98785a,a98786a,a98787a,a98790a,a98793a,a98794a,a98797a,a98800a,a98801a,a98802a,a98805a,a98808a,a98809a,a98812a,a98815a,a98816a,a98817a,a98820a,a98823a,a98824a,a98827a,a98830a,a98831a,a98832a,a98835a,a98838a,a98839a,a98842a,a98845a,a98846a,a98847a,a98850a,a98853a,a98854a,a98857a,a98860a,a98861a,a98862a,a98865a,a98868a,a98869a,a98872a,a98875a,a98876a,a98877a,a98880a,a98883a,a98884a,a98887a,a98890a,a98891a,a98892a,a98895a,a98898a,a98899a,a98902a,a98905a,a98906a,a98907a,a98910a,a98913a,a98914a,a98917a,a98920a,a98921a,a98922a,a98925a,a98928a,a98929a,a98932a,a98935a,a98936a,a98937a,a98940a,a98943a,a98944a,a98947a,a98950a,a98951a,a98952a,a98955a,a98958a,a98959a,a98962a,a98965a,a98966a,a98967a,a98970a,a98973a,a98974a,a98977a,a98980a,a98981a,a98982a,a98985a,a98988a,a98989a,a98992a,a98995a,a98996a,a98997a,a99000a,a99003a,a99004a,a99007a,a99010a,a99011a,a99012a,a99015a,a99018a,a99019a,a99022a,a99025a,a99026a,a99027a,a99030a,a99033a,a99034a,a99037a,a99040a,a99041a,a99042a,a99045a,a99048a,a99049a,a99052a,a99055a,a99056a,a99057a,a99060a,a99063a,a99064a,a99067a,a99070a,a99071a,a99072a,a99075a,a99078a,a99079a,a99082a,a99085a,a99086a,a99087a,a99090a,a99093a,a99094a,a99097a,a99100a,a99101a,a99102a,a99105a,a99108a,a99109a,a99112a,a99115a,a99116a,a99117a,a99120a,a99123a,a99124a,a99127a,a99130a,a99131a,a99132a,a99135a,a99138a,a99139a,a99142a,a99145a,a99146a,a99147a,a99150a,a99153a,a99154a,a99157a,a99160a,a99161a,a99162a,a99165a,a99168a,a99169a,a99172a,a99175a,a99176a,a99177a,a99180a,a99183a,a99184a,a99187a,a99190a,a99191a,a99192a,a99195a,a99198a,a99199a,a99202a,a99205a,a99206a,a99207a,a99210a,a99213a,a99214a,a99217a,a99220a,a99221a,a99222a,a99225a,a99228a,a99229a,a99232a,a99235a,a99236a,a99237a,a99240a,a99243a,a99244a,a99247a,a99250a,a99251a,a99252a,a99255a,a99258a,a99259a,a99262a,a99265a,a99266a,a99267a,a99270a,a99273a,a99274a,a99277a,a99280a,a99281a,a99282a,a99285a,a99288a,a99289a,a99292a,a99295a,a99296a,a99297a,a99300a,a99303a,a99304a,a99307a,a99310a,a99311a,a99312a,a99315a,a99318a,a99319a,a99322a,a99325a,a99326a,a99327a,a99330a,a99333a,a99334a,a99337a,a99340a,a99341a,a99342a,a99345a,a99348a,a99349a,a99352a,a99355a,a99356a,a99357a,a99360a,a99363a,a99364a,a99367a,a99370a,a99371a,a99372a,a99375a,a99378a,a99379a,a99382a,a99385a,a99386a,a99387a,a99390a,a99393a,a99394a,a99397a,a99400a,a99401a,a99402a,a99405a,a99408a,a99409a,a99412a,a99415a,a99416a,a99417a,a99420a,a99423a,a99424a,a99427a,a99430a,a99431a,a99432a,a99435a,a99438a,a99439a,a99442a,a99445a,a99446a,a99447a,a99450a,a99453a,a99454a,a99457a,a99460a,a99461a,a99462a,a99465a,a99468a,a99469a,a99472a,a99475a,a99476a,a99477a,a99480a,a99483a,a99484a,a99487a,a99490a,a99491a,a99492a,a99495a,a99498a,a99499a,a99502a,a99505a,a99506a,a99507a,a99510a,a99513a,a99514a,a99517a,a99520a,a99521a,a99522a,a99525a,a99528a,a99529a,a99532a,a99535a,a99536a,a99537a,a99540a,a99543a,a99544a,a99547a,a99550a,a99551a,a99552a,a99555a,a99558a,a99559a,a99562a,a99565a,a99566a,a99567a,a99570a,a99573a,a99574a,a99577a,a99580a,a99581a,a99582a,a99585a,a99588a,a99589a,a99592a,a99595a,a99596a,a99597a,a99600a,a99603a,a99604a,a99607a,a99610a,a99611a,a99612a,a99615a,a99618a,a99619a,a99622a,a99625a,a99626a,a99627a,a99630a,a99633a,a99634a,a99637a,a99640a,a99641a,a99642a,a99645a,a99648a,a99649a,a99652a,a99655a,a99656a,a99657a,a99660a,a99663a,a99664a,a99667a,a99670a,a99671a,a99672a,a99675a,a99678a,a99679a,a99682a,a99685a,a99686a,a99687a,a99690a,a99693a,a99694a,a99697a,a99700a,a99701a,a99702a,a99705a,a99708a,a99709a,a99712a,a99715a,a99716a,a99717a,a99720a,a99723a,a99724a,a99727a,a99730a,a99731a,a99732a,a99735a,a99738a,a99739a,a99742a,a99745a,a99746a,a99747a,a99750a,a99753a,a99754a,a99757a,a99760a,a99761a,a99762a,a99765a,a99768a,a99769a,a99772a,a99775a,a99776a,a99777a,a99780a,a99783a,a99784a,a99787a,a99790a,a99791a,a99792a,a99795a,a99798a,a99799a,a99802a,a99805a,a99806a,a99807a,a99810a,a99813a,a99814a,a99817a,a99820a,a99821a,a99822a,a99825a,a99828a,a99829a,a99832a,a99835a,a99836a,a99837a,a99840a,a99843a,a99844a,a99847a,a99850a,a99851a,a99852a,a99855a,a99858a,a99859a,a99862a,a99865a,a99866a,a99867a,a99870a,a99873a,a99874a,a99877a,a99880a,a99881a,a99882a,a99885a,a99888a,a99889a,a99892a,a99895a,a99896a,a99897a,a99900a,a99903a,a99904a,a99907a,a99910a,a99911a,a99912a,a99915a,a99918a,a99919a,a99922a,a99925a,a99926a,a99927a,a99930a,a99933a,a99934a,a99937a,a99940a,a99941a,a99942a,a99945a,a99948a,a99949a,a99952a,a99955a,a99956a,a99957a,a99960a,a99963a,a99964a,a99967a,a99970a,a99971a,a99972a,a99975a,a99978a,a99979a,a99982a,a99985a,a99986a,a99987a,a99990a,a99993a,a99994a,a99997a,a100000a,a100001a,a100002a,a100005a,a100008a,a100009a,a100012a,a100015a,a100016a,a100017a,a100020a,a100023a,a100024a,a100027a,a100030a,a100031a,a100032a,a100035a,a100038a,a100039a,a100042a,a100045a,a100046a,a100047a,a100050a,a100053a,a100054a,a100057a,a100060a,a100061a,a100062a,a100065a,a100068a,a100069a,a100072a,a100075a,a100076a,a100077a,a100080a,a100083a,a100084a,a100087a,a100090a,a100091a,a100092a,a100095a,a100098a,a100099a,a100102a,a100105a,a100106a,a100107a,a100110a,a100113a,a100114a,a100117a,a100120a,a100121a,a100122a,a100125a,a100128a,a100129a,a100132a,a100135a,a100136a,a100137a,a100140a,a100143a,a100144a,a100147a,a100150a,a100151a,a100152a,a100155a,a100158a,a100159a,a100162a,a100165a,a100166a,a100167a,a100170a,a100173a,a100174a,a100177a,a100180a,a100181a,a100182a,a100185a,a100188a,a100189a,a100192a,a100195a,a100196a,a100197a,a100200a,a100203a,a100204a,a100207a,a100210a,a100211a,a100212a,a100215a,a100218a,a100219a,a100222a,a100225a,a100226a,a100227a,a100230a,a100233a,a100234a,a100237a,a100240a,a100241a,a100242a,a100245a,a100248a,a100249a,a100252a,a100255a,a100256a,a100257a,a100260a,a100263a,a100264a,a100267a,a100270a,a100271a,a100272a,a100275a,a100278a,a100279a,a100282a,a100285a,a100286a,a100287a,a100290a,a100293a,a100294a,a100297a,a100300a,a100301a,a100302a,a100305a,a100308a,a100309a,a100312a,a100315a,a100316a,a100317a,a100320a,a100323a,a100324a,a100327a,a100330a,a100331a,a100332a,a100335a,a100338a,a100339a,a100342a,a100345a,a100346a,a100347a,a100350a,a100353a,a100354a,a100357a,a100360a,a100361a,a100362a,a100365a,a100368a,a100369a,a100372a,a100375a,a100376a,a100377a,a100380a,a100383a,a100384a,a100387a,a100390a,a100391a,a100392a,a100395a,a100398a,a100399a,a100402a,a100405a,a100406a,a100407a,a100410a,a100413a,a100414a,a100417a,a100420a,a100421a,a100422a,a100425a,a100428a,a100429a,a100432a,a100435a,a100436a,a100437a,a100440a,a100443a,a100444a,a100447a,a100450a,a100451a,a100452a,a100455a,a100458a,a100459a,a100462a,a100465a,a100466a,a100467a,a100470a,a100473a,a100474a,a100477a,a100480a,a100481a,a100482a,a100485a,a100488a,a100489a,a100492a,a100495a,a100496a,a100497a,a100500a,a100503a,a100504a,a100507a,a100510a,a100511a,a100512a,a100515a,a100518a,a100519a,a100522a,a100525a,a100526a,a100527a,a100530a,a100533a,a100534a,a100537a,a100540a,a100541a,a100542a,a100545a,a100548a,a100549a,a100552a,a100555a,a100556a,a100557a,a100560a,a100563a,a100564a,a100567a,a100570a,a100571a,a100572a,a100575a,a100578a,a100579a,a100582a,a100585a,a100586a,a100587a,a100590a,a100593a,a100594a,a100597a,a100600a,a100601a,a100602a,a100605a,a100608a,a100609a,a100612a,a100615a,a100616a,a100617a,a100620a,a100623a,a100624a,a100627a,a100630a,a100631a,a100632a,a100635a,a100638a,a100639a,a100642a,a100645a,a100646a,a100647a,a100650a,a100653a,a100654a,a100657a,a100660a,a100661a,a100662a,a100665a,a100668a,a100669a,a100672a,a100675a,a100676a,a100677a,a100680a,a100683a,a100684a,a100687a,a100690a,a100691a,a100692a,a100695a,a100698a,a100699a,a100702a,a100705a,a100706a,a100707a,a100710a,a100713a,a100714a,a100717a,a100720a,a100721a,a100722a,a100725a,a100728a,a100729a,a100732a,a100735a,a100736a,a100737a,a100740a,a100743a,a100744a,a100747a,a100750a,a100751a,a100752a,a100755a,a100758a,a100759a,a100762a,a100765a,a100766a,a100767a,a100770a,a100773a,a100774a,a100777a,a100780a,a100781a,a100782a,a100785a,a100788a,a100789a,a100792a,a100795a,a100796a,a100797a,a100800a,a100803a,a100804a,a100807a,a100810a,a100811a,a100812a,a100815a,a100818a,a100819a,a100822a,a100825a,a100826a,a100827a,a100830a,a100833a,a100834a,a100837a,a100840a,a100841a,a100842a,a100845a,a100848a,a100849a,a100852a,a100855a,a100856a,a100857a,a100860a,a100863a,a100864a,a100867a,a100870a,a100871a,a100872a,a100875a,a100878a,a100879a,a100882a,a100885a,a100886a,a100887a,a100890a,a100893a,a100894a,a100897a,a100900a,a100901a,a100902a,a100905a,a100908a,a100909a,a100912a,a100915a,a100916a,a100917a,a100920a,a100923a,a100924a,a100927a,a100930a,a100931a,a100932a,a100935a,a100938a,a100939a,a100942a,a100945a,a100946a,a100947a,a100950a,a100953a,a100954a,a100957a,a100960a,a100961a,a100962a,a100965a,a100968a,a100969a,a100972a,a100975a,a100976a,a100977a,a100980a,a100983a,a100984a,a100987a,a100991a,a100992a,a100993a,a100994a,a100997a,a101000a,a101001a,a101004a,a101007a,a101008a,a101009a,a101012a,a101015a,a101016a,a101019a,a101023a,a101024a,a101025a,a101026a,a101029a,a101032a,a101033a,a101036a,a101039a,a101040a,a101041a,a101044a,a101047a,a101048a,a101051a,a101055a,a101056a,a101057a,a101058a,a101061a,a101064a,a101065a,a101068a,a101071a,a101072a,a101073a,a101076a,a101079a,a101080a,a101083a,a101087a,a101088a,a101089a,a101090a,a101093a,a101096a,a101097a,a101100a,a101103a,a101104a,a101105a,a101108a,a101111a,a101112a,a101115a,a101119a,a101120a,a101121a,a101122a,a101125a,a101128a,a101129a,a101132a,a101135a,a101136a,a101137a,a101140a,a101143a,a101144a,a101147a,a101151a,a101152a,a101153a,a101154a: std_logic;
begin

A109 <=( a11314a ) or ( a7543a );
 a1a <=( a101154a  and  a101137a );
 a2a <=( a101122a  and  a101105a );
 a3a <=( a101090a  and  a101073a );
 a4a <=( a101058a  and  a101041a );
 a5a <=( a101026a  and  a101009a );
 a6a <=( a100994a  and  a100977a );
 a7a <=( a100962a  and  a100947a );
 a8a <=( a100932a  and  a100917a );
 a9a <=( a100902a  and  a100887a );
 a10a <=( a100872a  and  a100857a );
 a11a <=( a100842a  and  a100827a );
 a12a <=( a100812a  and  a100797a );
 a13a <=( a100782a  and  a100767a );
 a14a <=( a100752a  and  a100737a );
 a15a <=( a100722a  and  a100707a );
 a16a <=( a100692a  and  a100677a );
 a17a <=( a100662a  and  a100647a );
 a18a <=( a100632a  and  a100617a );
 a19a <=( a100602a  and  a100587a );
 a20a <=( a100572a  and  a100557a );
 a21a <=( a100542a  and  a100527a );
 a22a <=( a100512a  and  a100497a );
 a23a <=( a100482a  and  a100467a );
 a24a <=( a100452a  and  a100437a );
 a25a <=( a100422a  and  a100407a );
 a26a <=( a100392a  and  a100377a );
 a27a <=( a100362a  and  a100347a );
 a28a <=( a100332a  and  a100317a );
 a29a <=( a100302a  and  a100287a );
 a30a <=( a100272a  and  a100257a );
 a31a <=( a100242a  and  a100227a );
 a32a <=( a100212a  and  a100197a );
 a33a <=( a100182a  and  a100167a );
 a34a <=( a100152a  and  a100137a );
 a35a <=( a100122a  and  a100107a );
 a36a <=( a100092a  and  a100077a );
 a37a <=( a100062a  and  a100047a );
 a38a <=( a100032a  and  a100017a );
 a39a <=( a100002a  and  a99987a );
 a40a <=( a99972a  and  a99957a );
 a41a <=( a99942a  and  a99927a );
 a42a <=( a99912a  and  a99897a );
 a43a <=( a99882a  and  a99867a );
 a44a <=( a99852a  and  a99837a );
 a45a <=( a99822a  and  a99807a );
 a46a <=( a99792a  and  a99777a );
 a47a <=( a99762a  and  a99747a );
 a48a <=( a99732a  and  a99717a );
 a49a <=( a99702a  and  a99687a );
 a50a <=( a99672a  and  a99657a );
 a51a <=( a99642a  and  a99627a );
 a52a <=( a99612a  and  a99597a );
 a53a <=( a99582a  and  a99567a );
 a54a <=( a99552a  and  a99537a );
 a55a <=( a99522a  and  a99507a );
 a56a <=( a99492a  and  a99477a );
 a57a <=( a99462a  and  a99447a );
 a58a <=( a99432a  and  a99417a );
 a59a <=( a99402a  and  a99387a );
 a60a <=( a99372a  and  a99357a );
 a61a <=( a99342a  and  a99327a );
 a62a <=( a99312a  and  a99297a );
 a63a <=( a99282a  and  a99267a );
 a64a <=( a99252a  and  a99237a );
 a65a <=( a99222a  and  a99207a );
 a66a <=( a99192a  and  a99177a );
 a67a <=( a99162a  and  a99147a );
 a68a <=( a99132a  and  a99117a );
 a69a <=( a99102a  and  a99087a );
 a70a <=( a99072a  and  a99057a );
 a71a <=( a99042a  and  a99027a );
 a72a <=( a99012a  and  a98997a );
 a73a <=( a98982a  and  a98967a );
 a74a <=( a98952a  and  a98937a );
 a75a <=( a98922a  and  a98907a );
 a76a <=( a98892a  and  a98877a );
 a77a <=( a98862a  and  a98847a );
 a78a <=( a98832a  and  a98817a );
 a79a <=( a98802a  and  a98787a );
 a80a <=( a98772a  and  a98757a );
 a81a <=( a98742a  and  a98727a );
 a82a <=( a98712a  and  a98697a );
 a83a <=( a98682a  and  a98667a );
 a84a <=( a98652a  and  a98637a );
 a85a <=( a98622a  and  a98607a );
 a86a <=( a98592a  and  a98577a );
 a87a <=( a98562a  and  a98547a );
 a88a <=( a98532a  and  a98517a );
 a89a <=( a98502a  and  a98487a );
 a90a <=( a98472a  and  a98457a );
 a91a <=( a98442a  and  a98427a );
 a92a <=( a98412a  and  a98397a );
 a93a <=( a98382a  and  a98367a );
 a94a <=( a98352a  and  a98337a );
 a95a <=( a98322a  and  a98307a );
 a96a <=( a98292a  and  a98277a );
 a97a <=( a98262a  and  a98247a );
 a98a <=( a98232a  and  a98217a );
 a99a <=( a98202a  and  a98187a );
 a100a <=( a98172a  and  a98157a );
 a101a <=( a98142a  and  a98127a );
 a102a <=( a98112a  and  a98097a );
 a103a <=( a98082a  and  a98067a );
 a104a <=( a98052a  and  a98037a );
 a105a <=( a98022a  and  a98007a );
 a106a <=( a97992a  and  a97977a );
 a107a <=( a97962a  and  a97947a );
 a108a <=( a97932a  and  a97917a );
 a109a <=( a97902a  and  a97887a );
 a110a <=( a97872a  and  a97857a );
 a111a <=( a97842a  and  a97827a );
 a112a <=( a97812a  and  a97797a );
 a113a <=( a97782a  and  a97767a );
 a114a <=( a97752a  and  a97737a );
 a115a <=( a97722a  and  a97707a );
 a116a <=( a97692a  and  a97677a );
 a117a <=( a97662a  and  a97647a );
 a118a <=( a97632a  and  a97617a );
 a119a <=( a97602a  and  a97587a );
 a120a <=( a97572a  and  a97557a );
 a121a <=( a97542a  and  a97527a );
 a122a <=( a97514a  and  a97499a );
 a123a <=( a97486a  and  a97471a );
 a124a <=( a97458a  and  a97443a );
 a125a <=( a97430a  and  a97415a );
 a126a <=( a97402a  and  a97387a );
 a127a <=( a97374a  and  a97359a );
 a128a <=( a97346a  and  a97331a );
 a129a <=( a97318a  and  a97303a );
 a130a <=( a97290a  and  a97275a );
 a131a <=( a97262a  and  a97247a );
 a132a <=( a97234a  and  a97219a );
 a133a <=( a97206a  and  a97191a );
 a134a <=( a97178a  and  a97163a );
 a135a <=( a97150a  and  a97135a );
 a136a <=( a97122a  and  a97107a );
 a137a <=( a97094a  and  a97079a );
 a138a <=( a97066a  and  a97051a );
 a139a <=( a97038a  and  a97023a );
 a140a <=( a97010a  and  a96995a );
 a141a <=( a96982a  and  a96967a );
 a142a <=( a96954a  and  a96939a );
 a143a <=( a96926a  and  a96911a );
 a144a <=( a96898a  and  a96883a );
 a145a <=( a96870a  and  a96855a );
 a146a <=( a96842a  and  a96827a );
 a147a <=( a96814a  and  a96799a );
 a148a <=( a96786a  and  a96771a );
 a149a <=( a96758a  and  a96743a );
 a150a <=( a96730a  and  a96715a );
 a151a <=( a96702a  and  a96687a );
 a152a <=( a96674a  and  a96659a );
 a153a <=( a96646a  and  a96631a );
 a154a <=( a96618a  and  a96603a );
 a155a <=( a96590a  and  a96575a );
 a156a <=( a96562a  and  a96547a );
 a157a <=( a96534a  and  a96519a );
 a158a <=( a96506a  and  a96491a );
 a159a <=( a96478a  and  a96463a );
 a160a <=( a96450a  and  a96435a );
 a161a <=( a96422a  and  a96407a );
 a162a <=( a96394a  and  a96379a );
 a163a <=( a96366a  and  a96351a );
 a164a <=( a96338a  and  a96323a );
 a165a <=( a96310a  and  a96295a );
 a166a <=( a96282a  and  a96267a );
 a167a <=( a96254a  and  a96239a );
 a168a <=( a96226a  and  a96211a );
 a169a <=( a96198a  and  a96183a );
 a170a <=( a96170a  and  a96155a );
 a171a <=( a96142a  and  a96127a );
 a172a <=( a96114a  and  a96099a );
 a173a <=( a96086a  and  a96071a );
 a174a <=( a96058a  and  a96043a );
 a175a <=( a96030a  and  a96015a );
 a176a <=( a96002a  and  a95987a );
 a177a <=( a95974a  and  a95959a );
 a178a <=( a95946a  and  a95931a );
 a179a <=( a95918a  and  a95903a );
 a180a <=( a95890a  and  a95875a );
 a181a <=( a95862a  and  a95847a );
 a182a <=( a95834a  and  a95819a );
 a183a <=( a95806a  and  a95791a );
 a184a <=( a95778a  and  a95763a );
 a185a <=( a95750a  and  a95735a );
 a186a <=( a95722a  and  a95707a );
 a187a <=( a95694a  and  a95679a );
 a188a <=( a95666a  and  a95651a );
 a189a <=( a95638a  and  a95623a );
 a190a <=( a95610a  and  a95595a );
 a191a <=( a95582a  and  a95567a );
 a192a <=( a95554a  and  a95539a );
 a193a <=( a95526a  and  a95511a );
 a194a <=( a95498a  and  a95483a );
 a195a <=( a95470a  and  a95455a );
 a196a <=( a95442a  and  a95427a );
 a197a <=( a95414a  and  a95399a );
 a198a <=( a95386a  and  a95371a );
 a199a <=( a95358a  and  a95343a );
 a200a <=( a95330a  and  a95315a );
 a201a <=( a95302a  and  a95287a );
 a202a <=( a95274a  and  a95259a );
 a203a <=( a95246a  and  a95231a );
 a204a <=( a95218a  and  a95203a );
 a205a <=( a95190a  and  a95175a );
 a206a <=( a95162a  and  a95147a );
 a207a <=( a95134a  and  a95119a );
 a208a <=( a95106a  and  a95091a );
 a209a <=( a95078a  and  a95063a );
 a210a <=( a95050a  and  a95035a );
 a211a <=( a95022a  and  a95007a );
 a212a <=( a94994a  and  a94979a );
 a213a <=( a94966a  and  a94951a );
 a214a <=( a94938a  and  a94923a );
 a215a <=( a94910a  and  a94895a );
 a216a <=( a94882a  and  a94867a );
 a217a <=( a94854a  and  a94839a );
 a218a <=( a94826a  and  a94811a );
 a219a <=( a94798a  and  a94783a );
 a220a <=( a94770a  and  a94755a );
 a221a <=( a94742a  and  a94727a );
 a222a <=( a94714a  and  a94699a );
 a223a <=( a94686a  and  a94671a );
 a224a <=( a94658a  and  a94643a );
 a225a <=( a94630a  and  a94615a );
 a226a <=( a94602a  and  a94587a );
 a227a <=( a94574a  and  a94559a );
 a228a <=( a94546a  and  a94531a );
 a229a <=( a94518a  and  a94503a );
 a230a <=( a94490a  and  a94475a );
 a231a <=( a94462a  and  a94447a );
 a232a <=( a94434a  and  a94419a );
 a233a <=( a94406a  and  a94391a );
 a234a <=( a94378a  and  a94363a );
 a235a <=( a94350a  and  a94335a );
 a236a <=( a94322a  and  a94307a );
 a237a <=( a94294a  and  a94279a );
 a238a <=( a94266a  and  a94251a );
 a239a <=( a94238a  and  a94223a );
 a240a <=( a94210a  and  a94195a );
 a241a <=( a94182a  and  a94167a );
 a242a <=( a94154a  and  a94139a );
 a243a <=( a94126a  and  a94111a );
 a244a <=( a94098a  and  a94083a );
 a245a <=( a94070a  and  a94055a );
 a246a <=( a94042a  and  a94027a );
 a247a <=( a94014a  and  a93999a );
 a248a <=( a93986a  and  a93971a );
 a249a <=( a93958a  and  a93943a );
 a250a <=( a93930a  and  a93915a );
 a251a <=( a93902a  and  a93887a );
 a252a <=( a93874a  and  a93859a );
 a253a <=( a93846a  and  a93831a );
 a254a <=( a93818a  and  a93803a );
 a255a <=( a93790a  and  a93775a );
 a256a <=( a93762a  and  a93747a );
 a257a <=( a93734a  and  a93719a );
 a258a <=( a93706a  and  a93691a );
 a259a <=( a93678a  and  a93663a );
 a260a <=( a93650a  and  a93635a );
 a261a <=( a93622a  and  a93607a );
 a262a <=( a93594a  and  a93579a );
 a263a <=( a93566a  and  a93551a );
 a264a <=( a93538a  and  a93523a );
 a265a <=( a93510a  and  a93495a );
 a266a <=( a93482a  and  a93467a );
 a267a <=( a93454a  and  a93439a );
 a268a <=( a93426a  and  a93411a );
 a269a <=( a93398a  and  a93383a );
 a270a <=( a93370a  and  a93355a );
 a271a <=( a93342a  and  a93327a );
 a272a <=( a93314a  and  a93299a );
 a273a <=( a93286a  and  a93271a );
 a274a <=( a93258a  and  a93243a );
 a275a <=( a93230a  and  a93215a );
 a276a <=( a93202a  and  a93187a );
 a277a <=( a93174a  and  a93159a );
 a278a <=( a93146a  and  a93131a );
 a279a <=( a93118a  and  a93103a );
 a280a <=( a93090a  and  a93075a );
 a281a <=( a93062a  and  a93047a );
 a282a <=( a93034a  and  a93019a );
 a283a <=( a93006a  and  a92991a );
 a284a <=( a92978a  and  a92963a );
 a285a <=( a92950a  and  a92935a );
 a286a <=( a92922a  and  a92907a );
 a287a <=( a92894a  and  a92879a );
 a288a <=( a92866a  and  a92851a );
 a289a <=( a92838a  and  a92823a );
 a290a <=( a92810a  and  a92795a );
 a291a <=( a92782a  and  a92767a );
 a292a <=( a92754a  and  a92739a );
 a293a <=( a92726a  and  a92711a );
 a294a <=( a92698a  and  a92683a );
 a295a <=( a92670a  and  a92655a );
 a296a <=( a92642a  and  a92627a );
 a297a <=( a92614a  and  a92599a );
 a298a <=( a92586a  and  a92571a );
 a299a <=( a92558a  and  a92543a );
 a300a <=( a92530a  and  a92515a );
 a301a <=( a92502a  and  a92487a );
 a302a <=( a92474a  and  a92459a );
 a303a <=( a92446a  and  a92431a );
 a304a <=( a92418a  and  a92403a );
 a305a <=( a92390a  and  a92375a );
 a306a <=( a92362a  and  a92347a );
 a307a <=( a92334a  and  a92319a );
 a308a <=( a92306a  and  a92291a );
 a309a <=( a92278a  and  a92263a );
 a310a <=( a92250a  and  a92235a );
 a311a <=( a92222a  and  a92207a );
 a312a <=( a92194a  and  a92179a );
 a313a <=( a92166a  and  a92151a );
 a314a <=( a92138a  and  a92123a );
 a315a <=( a92110a  and  a92095a );
 a316a <=( a92082a  and  a92067a );
 a317a <=( a92054a  and  a92039a );
 a318a <=( a92026a  and  a92011a );
 a319a <=( a91998a  and  a91983a );
 a320a <=( a91970a  and  a91955a );
 a321a <=( a91942a  and  a91927a );
 a322a <=( a91914a  and  a91899a );
 a323a <=( a91886a  and  a91871a );
 a324a <=( a91858a  and  a91843a );
 a325a <=( a91830a  and  a91815a );
 a326a <=( a91802a  and  a91787a );
 a327a <=( a91774a  and  a91759a );
 a328a <=( a91746a  and  a91731a );
 a329a <=( a91718a  and  a91703a );
 a330a <=( a91690a  and  a91675a );
 a331a <=( a91662a  and  a91647a );
 a332a <=( a91634a  and  a91619a );
 a333a <=( a91606a  and  a91591a );
 a334a <=( a91578a  and  a91563a );
 a335a <=( a91550a  and  a91535a );
 a336a <=( a91522a  and  a91507a );
 a337a <=( a91494a  and  a91479a );
 a338a <=( a91466a  and  a91451a );
 a339a <=( a91438a  and  a91423a );
 a340a <=( a91410a  and  a91395a );
 a341a <=( a91382a  and  a91367a );
 a342a <=( a91354a  and  a91339a );
 a343a <=( a91326a  and  a91311a );
 a344a <=( a91298a  and  a91283a );
 a345a <=( a91270a  and  a91255a );
 a346a <=( a91242a  and  a91227a );
 a347a <=( a91214a  and  a91199a );
 a348a <=( a91186a  and  a91171a );
 a349a <=( a91158a  and  a91143a );
 a350a <=( a91130a  and  a91115a );
 a351a <=( a91102a  and  a91087a );
 a352a <=( a91074a  and  a91059a );
 a353a <=( a91046a  and  a91031a );
 a354a <=( a91018a  and  a91003a );
 a355a <=( a90990a  and  a90975a );
 a356a <=( a90962a  and  a90947a );
 a357a <=( a90934a  and  a90919a );
 a358a <=( a90906a  and  a90891a );
 a359a <=( a90878a  and  a90863a );
 a360a <=( a90850a  and  a90835a );
 a361a <=( a90822a  and  a90807a );
 a362a <=( a90794a  and  a90779a );
 a363a <=( a90766a  and  a90751a );
 a364a <=( a90738a  and  a90723a );
 a365a <=( a90710a  and  a90695a );
 a366a <=( a90682a  and  a90667a );
 a367a <=( a90654a  and  a90639a );
 a368a <=( a90626a  and  a90611a );
 a369a <=( a90598a  and  a90583a );
 a370a <=( a90570a  and  a90555a );
 a371a <=( a90542a  and  a90527a );
 a372a <=( a90514a  and  a90499a );
 a373a <=( a90486a  and  a90471a );
 a374a <=( a90458a  and  a90443a );
 a375a <=( a90430a  and  a90415a );
 a376a <=( a90402a  and  a90387a );
 a377a <=( a90374a  and  a90359a );
 a378a <=( a90346a  and  a90331a );
 a379a <=( a90318a  and  a90303a );
 a380a <=( a90290a  and  a90275a );
 a381a <=( a90262a  and  a90247a );
 a382a <=( a90234a  and  a90219a );
 a383a <=( a90206a  and  a90191a );
 a384a <=( a90178a  and  a90163a );
 a385a <=( a90150a  and  a90135a );
 a386a <=( a90122a  and  a90107a );
 a387a <=( a90094a  and  a90079a );
 a388a <=( a90066a  and  a90051a );
 a389a <=( a90038a  and  a90023a );
 a390a <=( a90010a  and  a89995a );
 a391a <=( a89982a  and  a89967a );
 a392a <=( a89954a  and  a89939a );
 a393a <=( a89926a  and  a89911a );
 a394a <=( a89898a  and  a89883a );
 a395a <=( a89870a  and  a89855a );
 a396a <=( a89842a  and  a89827a );
 a397a <=( a89814a  and  a89799a );
 a398a <=( a89786a  and  a89771a );
 a399a <=( a89758a  and  a89743a );
 a400a <=( a89730a  and  a89715a );
 a401a <=( a89702a  and  a89687a );
 a402a <=( a89674a  and  a89659a );
 a403a <=( a89646a  and  a89631a );
 a404a <=( a89618a  and  a89603a );
 a405a <=( a89590a  and  a89575a );
 a406a <=( a89562a  and  a89547a );
 a407a <=( a89534a  and  a89519a );
 a408a <=( a89506a  and  a89491a );
 a409a <=( a89478a  and  a89463a );
 a410a <=( a89450a  and  a89435a );
 a411a <=( a89422a  and  a89407a );
 a412a <=( a89394a  and  a89379a );
 a413a <=( a89366a  and  a89351a );
 a414a <=( a89338a  and  a89323a );
 a415a <=( a89310a  and  a89295a );
 a416a <=( a89282a  and  a89267a );
 a417a <=( a89254a  and  a89239a );
 a418a <=( a89226a  and  a89211a );
 a419a <=( a89198a  and  a89183a );
 a420a <=( a89170a  and  a89155a );
 a421a <=( a89142a  and  a89127a );
 a422a <=( a89114a  and  a89099a );
 a423a <=( a89086a  and  a89071a );
 a424a <=( a89058a  and  a89043a );
 a425a <=( a89030a  and  a89015a );
 a426a <=( a89002a  and  a88987a );
 a427a <=( a88974a  and  a88959a );
 a428a <=( a88946a  and  a88931a );
 a429a <=( a88918a  and  a88903a );
 a430a <=( a88890a  and  a88875a );
 a431a <=( a88862a  and  a88847a );
 a432a <=( a88834a  and  a88819a );
 a433a <=( a88806a  and  a88791a );
 a434a <=( a88778a  and  a88763a );
 a435a <=( a88750a  and  a88735a );
 a436a <=( a88722a  and  a88707a );
 a437a <=( a88694a  and  a88679a );
 a438a <=( a88666a  and  a88651a );
 a439a <=( a88638a  and  a88623a );
 a440a <=( a88610a  and  a88595a );
 a441a <=( a88582a  and  a88567a );
 a442a <=( a88554a  and  a88539a );
 a443a <=( a88526a  and  a88511a );
 a444a <=( a88498a  and  a88483a );
 a445a <=( a88470a  and  a88455a );
 a446a <=( a88442a  and  a88427a );
 a447a <=( a88414a  and  a88399a );
 a448a <=( a88386a  and  a88371a );
 a449a <=( a88358a  and  a88343a );
 a450a <=( a88330a  and  a88315a );
 a451a <=( a88302a  and  a88287a );
 a452a <=( a88274a  and  a88259a );
 a453a <=( a88246a  and  a88231a );
 a454a <=( a88218a  and  a88203a );
 a455a <=( a88190a  and  a88175a );
 a456a <=( a88162a  and  a88147a );
 a457a <=( a88134a  and  a88119a );
 a458a <=( a88106a  and  a88091a );
 a459a <=( a88078a  and  a88063a );
 a460a <=( a88050a  and  a88035a );
 a461a <=( a88022a  and  a88007a );
 a462a <=( a87994a  and  a87979a );
 a463a <=( a87966a  and  a87951a );
 a464a <=( a87938a  and  a87923a );
 a465a <=( a87910a  and  a87895a );
 a466a <=( a87882a  and  a87867a );
 a467a <=( a87854a  and  a87839a );
 a468a <=( a87826a  and  a87811a );
 a469a <=( a87798a  and  a87783a );
 a470a <=( a87770a  and  a87755a );
 a471a <=( a87742a  and  a87727a );
 a472a <=( a87714a  and  a87699a );
 a473a <=( a87686a  and  a87671a );
 a474a <=( a87658a  and  a87643a );
 a475a <=( a87630a  and  a87615a );
 a476a <=( a87602a  and  a87587a );
 a477a <=( a87574a  and  a87559a );
 a478a <=( a87546a  and  a87531a );
 a479a <=( a87518a  and  a87503a );
 a480a <=( a87490a  and  a87475a );
 a481a <=( a87462a  and  a87447a );
 a482a <=( a87434a  and  a87419a );
 a483a <=( a87406a  and  a87391a );
 a484a <=( a87378a  and  a87363a );
 a485a <=( a87350a  and  a87335a );
 a486a <=( a87322a  and  a87307a );
 a487a <=( a87294a  and  a87279a );
 a488a <=( a87266a  and  a87251a );
 a489a <=( a87238a  and  a87223a );
 a490a <=( a87210a  and  a87195a );
 a491a <=( a87182a  and  a87167a );
 a492a <=( a87154a  and  a87139a );
 a493a <=( a87126a  and  a87111a );
 a494a <=( a87098a  and  a87083a );
 a495a <=( a87070a  and  a87055a );
 a496a <=( a87042a  and  a87027a );
 a497a <=( a87014a  and  a86999a );
 a498a <=( a86986a  and  a86971a );
 a499a <=( a86958a  and  a86943a );
 a500a <=( a86930a  and  a86915a );
 a501a <=( a86902a  and  a86887a );
 a502a <=( a86874a  and  a86859a );
 a503a <=( a86846a  and  a86831a );
 a504a <=( a86818a  and  a86803a );
 a505a <=( a86790a  and  a86777a );
 a506a <=( a86764a  and  a86751a );
 a507a <=( a86738a  and  a86725a );
 a508a <=( a86712a  and  a86699a );
 a509a <=( a86686a  and  a86673a );
 a510a <=( a86660a  and  a86647a );
 a511a <=( a86634a  and  a86621a );
 a512a <=( a86608a  and  a86595a );
 a513a <=( a86582a  and  a86569a );
 a514a <=( a86556a  and  a86543a );
 a515a <=( a86530a  and  a86517a );
 a516a <=( a86504a  and  a86491a );
 a517a <=( a86478a  and  a86465a );
 a518a <=( a86452a  and  a86439a );
 a519a <=( a86426a  and  a86413a );
 a520a <=( a86400a  and  a86387a );
 a521a <=( a86374a  and  a86361a );
 a522a <=( a86348a  and  a86335a );
 a523a <=( a86322a  and  a86309a );
 a524a <=( a86296a  and  a86283a );
 a525a <=( a86270a  and  a86257a );
 a526a <=( a86244a  and  a86231a );
 a527a <=( a86218a  and  a86205a );
 a528a <=( a86192a  and  a86179a );
 a529a <=( a86166a  and  a86153a );
 a530a <=( a86140a  and  a86127a );
 a531a <=( a86114a  and  a86101a );
 a532a <=( a86088a  and  a86075a );
 a533a <=( a86062a  and  a86049a );
 a534a <=( a86036a  and  a86023a );
 a535a <=( a86010a  and  a85997a );
 a536a <=( a85984a  and  a85971a );
 a537a <=( a85958a  and  a85945a );
 a538a <=( a85932a  and  a85919a );
 a539a <=( a85906a  and  a85893a );
 a540a <=( a85880a  and  a85867a );
 a541a <=( a85854a  and  a85841a );
 a542a <=( a85828a  and  a85815a );
 a543a <=( a85802a  and  a85789a );
 a544a <=( a85776a  and  a85763a );
 a545a <=( a85750a  and  a85737a );
 a546a <=( a85724a  and  a85711a );
 a547a <=( a85698a  and  a85685a );
 a548a <=( a85672a  and  a85659a );
 a549a <=( a85646a  and  a85633a );
 a550a <=( a85620a  and  a85607a );
 a551a <=( a85594a  and  a85581a );
 a552a <=( a85568a  and  a85555a );
 a553a <=( a85542a  and  a85529a );
 a554a <=( a85516a  and  a85503a );
 a555a <=( a85490a  and  a85477a );
 a556a <=( a85464a  and  a85451a );
 a557a <=( a85438a  and  a85425a );
 a558a <=( a85412a  and  a85399a );
 a559a <=( a85386a  and  a85373a );
 a560a <=( a85360a  and  a85347a );
 a561a <=( a85334a  and  a85321a );
 a562a <=( a85308a  and  a85295a );
 a563a <=( a85282a  and  a85269a );
 a564a <=( a85256a  and  a85243a );
 a565a <=( a85230a  and  a85217a );
 a566a <=( a85204a  and  a85191a );
 a567a <=( a85178a  and  a85165a );
 a568a <=( a85152a  and  a85139a );
 a569a <=( a85126a  and  a85113a );
 a570a <=( a85100a  and  a85087a );
 a571a <=( a85074a  and  a85061a );
 a572a <=( a85048a  and  a85035a );
 a573a <=( a85022a  and  a85009a );
 a574a <=( a84996a  and  a84983a );
 a575a <=( a84970a  and  a84957a );
 a576a <=( a84944a  and  a84931a );
 a577a <=( a84918a  and  a84905a );
 a578a <=( a84892a  and  a84879a );
 a579a <=( a84866a  and  a84853a );
 a580a <=( a84840a  and  a84827a );
 a581a <=( a84814a  and  a84801a );
 a582a <=( a84788a  and  a84775a );
 a583a <=( a84762a  and  a84749a );
 a584a <=( a84736a  and  a84723a );
 a585a <=( a84710a  and  a84697a );
 a586a <=( a84684a  and  a84671a );
 a587a <=( a84658a  and  a84645a );
 a588a <=( a84632a  and  a84619a );
 a589a <=( a84606a  and  a84593a );
 a590a <=( a84580a  and  a84567a );
 a591a <=( a84554a  and  a84541a );
 a592a <=( a84528a  and  a84515a );
 a593a <=( a84502a  and  a84489a );
 a594a <=( a84476a  and  a84463a );
 a595a <=( a84450a  and  a84437a );
 a596a <=( a84424a  and  a84411a );
 a597a <=( a84398a  and  a84385a );
 a598a <=( a84372a  and  a84359a );
 a599a <=( a84346a  and  a84333a );
 a600a <=( a84320a  and  a84307a );
 a601a <=( a84294a  and  a84281a );
 a602a <=( a84268a  and  a84255a );
 a603a <=( a84242a  and  a84229a );
 a604a <=( a84216a  and  a84203a );
 a605a <=( a84190a  and  a84177a );
 a606a <=( a84164a  and  a84151a );
 a607a <=( a84138a  and  a84125a );
 a608a <=( a84112a  and  a84099a );
 a609a <=( a84086a  and  a84073a );
 a610a <=( a84060a  and  a84047a );
 a611a <=( a84034a  and  a84021a );
 a612a <=( a84008a  and  a83995a );
 a613a <=( a83982a  and  a83969a );
 a614a <=( a83956a  and  a83943a );
 a615a <=( a83930a  and  a83917a );
 a616a <=( a83904a  and  a83891a );
 a617a <=( a83878a  and  a83865a );
 a618a <=( a83852a  and  a83839a );
 a619a <=( a83826a  and  a83813a );
 a620a <=( a83800a  and  a83787a );
 a621a <=( a83774a  and  a83761a );
 a622a <=( a83748a  and  a83735a );
 a623a <=( a83722a  and  a83709a );
 a624a <=( a83696a  and  a83683a );
 a625a <=( a83670a  and  a83657a );
 a626a <=( a83644a  and  a83631a );
 a627a <=( a83618a  and  a83605a );
 a628a <=( a83592a  and  a83579a );
 a629a <=( a83566a  and  a83553a );
 a630a <=( a83540a  and  a83527a );
 a631a <=( a83514a  and  a83501a );
 a632a <=( a83488a  and  a83475a );
 a633a <=( a83462a  and  a83449a );
 a634a <=( a83436a  and  a83423a );
 a635a <=( a83410a  and  a83397a );
 a636a <=( a83384a  and  a83371a );
 a637a <=( a83358a  and  a83345a );
 a638a <=( a83332a  and  a83319a );
 a639a <=( a83306a  and  a83293a );
 a640a <=( a83280a  and  a83267a );
 a641a <=( a83254a  and  a83241a );
 a642a <=( a83228a  and  a83215a );
 a643a <=( a83202a  and  a83189a );
 a644a <=( a83176a  and  a83163a );
 a645a <=( a83150a  and  a83137a );
 a646a <=( a83124a  and  a83111a );
 a647a <=( a83098a  and  a83085a );
 a648a <=( a83072a  and  a83059a );
 a649a <=( a83046a  and  a83033a );
 a650a <=( a83020a  and  a83007a );
 a651a <=( a82994a  and  a82981a );
 a652a <=( a82968a  and  a82955a );
 a653a <=( a82942a  and  a82929a );
 a654a <=( a82916a  and  a82903a );
 a655a <=( a82890a  and  a82877a );
 a656a <=( a82864a  and  a82851a );
 a657a <=( a82838a  and  a82825a );
 a658a <=( a82812a  and  a82799a );
 a659a <=( a82786a  and  a82773a );
 a660a <=( a82760a  and  a82747a );
 a661a <=( a82734a  and  a82721a );
 a662a <=( a82708a  and  a82695a );
 a663a <=( a82682a  and  a82669a );
 a664a <=( a82656a  and  a82643a );
 a665a <=( a82630a  and  a82617a );
 a666a <=( a82604a  and  a82591a );
 a667a <=( a82578a  and  a82565a );
 a668a <=( a82552a  and  a82539a );
 a669a <=( a82526a  and  a82513a );
 a670a <=( a82500a  and  a82487a );
 a671a <=( a82474a  and  a82461a );
 a672a <=( a82448a  and  a82435a );
 a673a <=( a82422a  and  a82409a );
 a674a <=( a82396a  and  a82383a );
 a675a <=( a82370a  and  a82357a );
 a676a <=( a82344a  and  a82331a );
 a677a <=( a82318a  and  a82305a );
 a678a <=( a82292a  and  a82279a );
 a679a <=( a82266a  and  a82253a );
 a680a <=( a82240a  and  a82227a );
 a681a <=( a82214a  and  a82201a );
 a682a <=( a82188a  and  a82175a );
 a683a <=( a82162a  and  a82149a );
 a684a <=( a82136a  and  a82123a );
 a685a <=( a82110a  and  a82097a );
 a686a <=( a82084a  and  a82071a );
 a687a <=( a82058a  and  a82045a );
 a688a <=( a82032a  and  a82019a );
 a689a <=( a82006a  and  a81993a );
 a690a <=( a81980a  and  a81967a );
 a691a <=( a81954a  and  a81941a );
 a692a <=( a81928a  and  a81915a );
 a693a <=( a81902a  and  a81889a );
 a694a <=( a81876a  and  a81863a );
 a695a <=( a81850a  and  a81837a );
 a696a <=( a81824a  and  a81811a );
 a697a <=( a81798a  and  a81785a );
 a698a <=( a81772a  and  a81759a );
 a699a <=( a81746a  and  a81733a );
 a700a <=( a81720a  and  a81707a );
 a701a <=( a81694a  and  a81681a );
 a702a <=( a81668a  and  a81655a );
 a703a <=( a81642a  and  a81629a );
 a704a <=( a81616a  and  a81603a );
 a705a <=( a81590a  and  a81577a );
 a706a <=( a81564a  and  a81551a );
 a707a <=( a81538a  and  a81525a );
 a708a <=( a81512a  and  a81499a );
 a709a <=( a81486a  and  a81473a );
 a710a <=( a81460a  and  a81447a );
 a711a <=( a81434a  and  a81421a );
 a712a <=( a81408a  and  a81395a );
 a713a <=( a81382a  and  a81369a );
 a714a <=( a81356a  and  a81343a );
 a715a <=( a81330a  and  a81317a );
 a716a <=( a81304a  and  a81291a );
 a717a <=( a81278a  and  a81265a );
 a718a <=( a81252a  and  a81239a );
 a719a <=( a81226a  and  a81213a );
 a720a <=( a81200a  and  a81187a );
 a721a <=( a81174a  and  a81161a );
 a722a <=( a81148a  and  a81135a );
 a723a <=( a81122a  and  a81109a );
 a724a <=( a81096a  and  a81083a );
 a725a <=( a81070a  and  a81057a );
 a726a <=( a81044a  and  a81031a );
 a727a <=( a81018a  and  a81005a );
 a728a <=( a80992a  and  a80979a );
 a729a <=( a80966a  and  a80953a );
 a730a <=( a80940a  and  a80927a );
 a731a <=( a80914a  and  a80901a );
 a732a <=( a80888a  and  a80875a );
 a733a <=( a80862a  and  a80849a );
 a734a <=( a80836a  and  a80823a );
 a735a <=( a80810a  and  a80797a );
 a736a <=( a80784a  and  a80771a );
 a737a <=( a80758a  and  a80745a );
 a738a <=( a80732a  and  a80719a );
 a739a <=( a80706a  and  a80693a );
 a740a <=( a80680a  and  a80667a );
 a741a <=( a80654a  and  a80641a );
 a742a <=( a80628a  and  a80615a );
 a743a <=( a80602a  and  a80589a );
 a744a <=( a80576a  and  a80563a );
 a745a <=( a80550a  and  a80537a );
 a746a <=( a80524a  and  a80511a );
 a747a <=( a80498a  and  a80485a );
 a748a <=( a80472a  and  a80459a );
 a749a <=( a80446a  and  a80433a );
 a750a <=( a80420a  and  a80407a );
 a751a <=( a80394a  and  a80381a );
 a752a <=( a80368a  and  a80355a );
 a753a <=( a80342a  and  a80329a );
 a754a <=( a80316a  and  a80303a );
 a755a <=( a80290a  and  a80277a );
 a756a <=( a80264a  and  a80251a );
 a757a <=( a80238a  and  a80225a );
 a758a <=( a80212a  and  a80199a );
 a759a <=( a80186a  and  a80173a );
 a760a <=( a80160a  and  a80147a );
 a761a <=( a80134a  and  a80121a );
 a762a <=( a80108a  and  a80095a );
 a763a <=( a80082a  and  a80069a );
 a764a <=( a80056a  and  a80043a );
 a765a <=( a80030a  and  a80017a );
 a766a <=( a80004a  and  a79991a );
 a767a <=( a79978a  and  a79965a );
 a768a <=( a79952a  and  a79939a );
 a769a <=( a79926a  and  a79913a );
 a770a <=( a79900a  and  a79887a );
 a771a <=( a79874a  and  a79861a );
 a772a <=( a79848a  and  a79835a );
 a773a <=( a79822a  and  a79809a );
 a774a <=( a79796a  and  a79783a );
 a775a <=( a79770a  and  a79757a );
 a776a <=( a79744a  and  a79731a );
 a777a <=( a79718a  and  a79705a );
 a778a <=( a79692a  and  a79679a );
 a779a <=( a79666a  and  a79653a );
 a780a <=( a79640a  and  a79627a );
 a781a <=( a79614a  and  a79601a );
 a782a <=( a79588a  and  a79575a );
 a783a <=( a79562a  and  a79549a );
 a784a <=( a79536a  and  a79523a );
 a785a <=( a79510a  and  a79497a );
 a786a <=( a79484a  and  a79471a );
 a787a <=( a79458a  and  a79445a );
 a788a <=( a79432a  and  a79419a );
 a789a <=( a79406a  and  a79393a );
 a790a <=( a79380a  and  a79367a );
 a791a <=( a79354a  and  a79341a );
 a792a <=( a79328a  and  a79315a );
 a793a <=( a79302a  and  a79289a );
 a794a <=( a79276a  and  a79263a );
 a795a <=( a79250a  and  a79237a );
 a796a <=( a79224a  and  a79211a );
 a797a <=( a79198a  and  a79185a );
 a798a <=( a79172a  and  a79159a );
 a799a <=( a79146a  and  a79133a );
 a800a <=( a79120a  and  a79107a );
 a801a <=( a79094a  and  a79081a );
 a802a <=( a79068a  and  a79055a );
 a803a <=( a79042a  and  a79029a );
 a804a <=( a79016a  and  a79003a );
 a805a <=( a78990a  and  a78977a );
 a806a <=( a78964a  and  a78951a );
 a807a <=( a78938a  and  a78925a );
 a808a <=( a78912a  and  a78899a );
 a809a <=( a78886a  and  a78873a );
 a810a <=( a78860a  and  a78847a );
 a811a <=( a78834a  and  a78821a );
 a812a <=( a78808a  and  a78795a );
 a813a <=( a78782a  and  a78769a );
 a814a <=( a78756a  and  a78743a );
 a815a <=( a78730a  and  a78717a );
 a816a <=( a78704a  and  a78691a );
 a817a <=( a78678a  and  a78665a );
 a818a <=( a78652a  and  a78639a );
 a819a <=( a78626a  and  a78613a );
 a820a <=( a78600a  and  a78587a );
 a821a <=( a78574a  and  a78561a );
 a822a <=( a78548a  and  a78535a );
 a823a <=( a78522a  and  a78509a );
 a824a <=( a78496a  and  a78483a );
 a825a <=( a78470a  and  a78457a );
 a826a <=( a78444a  and  a78431a );
 a827a <=( a78418a  and  a78405a );
 a828a <=( a78392a  and  a78379a );
 a829a <=( a78366a  and  a78353a );
 a830a <=( a78340a  and  a78327a );
 a831a <=( a78314a  and  a78301a );
 a832a <=( a78288a  and  a78275a );
 a833a <=( a78262a  and  a78249a );
 a834a <=( a78236a  and  a78223a );
 a835a <=( a78210a  and  a78197a );
 a836a <=( a78184a  and  a78171a );
 a837a <=( a78158a  and  a78145a );
 a838a <=( a78132a  and  a78119a );
 a839a <=( a78106a  and  a78093a );
 a840a <=( a78080a  and  a78067a );
 a841a <=( a78054a  and  a78041a );
 a842a <=( a78028a  and  a78015a );
 a843a <=( a78002a  and  a77989a );
 a844a <=( a77976a  and  a77963a );
 a845a <=( a77950a  and  a77937a );
 a846a <=( a77924a  and  a77911a );
 a847a <=( a77898a  and  a77885a );
 a848a <=( a77872a  and  a77859a );
 a849a <=( a77846a  and  a77833a );
 a850a <=( a77820a  and  a77807a );
 a851a <=( a77794a  and  a77781a );
 a852a <=( a77768a  and  a77755a );
 a853a <=( a77742a  and  a77729a );
 a854a <=( a77716a  and  a77703a );
 a855a <=( a77690a  and  a77677a );
 a856a <=( a77664a  and  a77651a );
 a857a <=( a77638a  and  a77625a );
 a858a <=( a77612a  and  a77599a );
 a859a <=( a77586a  and  a77573a );
 a860a <=( a77560a  and  a77547a );
 a861a <=( a77534a  and  a77521a );
 a862a <=( a77508a  and  a77495a );
 a863a <=( a77482a  and  a77469a );
 a864a <=( a77456a  and  a77443a );
 a865a <=( a77430a  and  a77417a );
 a866a <=( a77404a  and  a77391a );
 a867a <=( a77378a  and  a77365a );
 a868a <=( a77352a  and  a77339a );
 a869a <=( a77326a  and  a77313a );
 a870a <=( a77300a  and  a77287a );
 a871a <=( a77274a  and  a77261a );
 a872a <=( a77248a  and  a77235a );
 a873a <=( a77222a  and  a77209a );
 a874a <=( a77196a  and  a77183a );
 a875a <=( a77170a  and  a77157a );
 a876a <=( a77144a  and  a77131a );
 a877a <=( a77118a  and  a77105a );
 a878a <=( a77092a  and  a77079a );
 a879a <=( a77066a  and  a77053a );
 a880a <=( a77040a  and  a77027a );
 a881a <=( a77014a  and  a77001a );
 a882a <=( a76988a  and  a76975a );
 a883a <=( a76962a  and  a76949a );
 a884a <=( a76936a  and  a76923a );
 a885a <=( a76910a  and  a76897a );
 a886a <=( a76884a  and  a76871a );
 a887a <=( a76858a  and  a76845a );
 a888a <=( a76832a  and  a76819a );
 a889a <=( a76806a  and  a76793a );
 a890a <=( a76780a  and  a76767a );
 a891a <=( a76754a  and  a76741a );
 a892a <=( a76728a  and  a76715a );
 a893a <=( a76702a  and  a76689a );
 a894a <=( a76676a  and  a76663a );
 a895a <=( a76650a  and  a76637a );
 a896a <=( a76624a  and  a76611a );
 a897a <=( a76598a  and  a76585a );
 a898a <=( a76572a  and  a76559a );
 a899a <=( a76546a  and  a76533a );
 a900a <=( a76520a  and  a76507a );
 a901a <=( a76494a  and  a76481a );
 a902a <=( a76468a  and  a76455a );
 a903a <=( a76442a  and  a76429a );
 a904a <=( a76416a  and  a76403a );
 a905a <=( a76390a  and  a76377a );
 a906a <=( a76364a  and  a76351a );
 a907a <=( a76338a  and  a76325a );
 a908a <=( a76312a  and  a76299a );
 a909a <=( a76286a  and  a76273a );
 a910a <=( a76260a  and  a76247a );
 a911a <=( a76234a  and  a76221a );
 a912a <=( a76208a  and  a76195a );
 a913a <=( a76182a  and  a76169a );
 a914a <=( a76156a  and  a76143a );
 a915a <=( a76130a  and  a76117a );
 a916a <=( a76104a  and  a76091a );
 a917a <=( a76078a  and  a76065a );
 a918a <=( a76052a  and  a76039a );
 a919a <=( a76026a  and  a76013a );
 a920a <=( a76000a  and  a75987a );
 a921a <=( a75974a  and  a75961a );
 a922a <=( a75948a  and  a75935a );
 a923a <=( a75922a  and  a75909a );
 a924a <=( a75896a  and  a75883a );
 a925a <=( a75870a  and  a75857a );
 a926a <=( a75844a  and  a75831a );
 a927a <=( a75818a  and  a75805a );
 a928a <=( a75792a  and  a75779a );
 a929a <=( a75766a  and  a75753a );
 a930a <=( a75740a  and  a75727a );
 a931a <=( a75714a  and  a75701a );
 a932a <=( a75688a  and  a75675a );
 a933a <=( a75662a  and  a75649a );
 a934a <=( a75636a  and  a75623a );
 a935a <=( a75610a  and  a75597a );
 a936a <=( a75584a  and  a75571a );
 a937a <=( a75558a  and  a75545a );
 a938a <=( a75532a  and  a75519a );
 a939a <=( a75506a  and  a75493a );
 a940a <=( a75480a  and  a75467a );
 a941a <=( a75454a  and  a75441a );
 a942a <=( a75428a  and  a75415a );
 a943a <=( a75402a  and  a75389a );
 a944a <=( a75376a  and  a75363a );
 a945a <=( a75350a  and  a75337a );
 a946a <=( a75324a  and  a75311a );
 a947a <=( a75298a  and  a75285a );
 a948a <=( a75272a  and  a75259a );
 a949a <=( a75246a  and  a75233a );
 a950a <=( a75220a  and  a75207a );
 a951a <=( a75194a  and  a75181a );
 a952a <=( a75168a  and  a75155a );
 a953a <=( a75142a  and  a75129a );
 a954a <=( a75116a  and  a75103a );
 a955a <=( a75090a  and  a75077a );
 a956a <=( a75064a  and  a75051a );
 a957a <=( a75038a  and  a75025a );
 a958a <=( a75012a  and  a74999a );
 a959a <=( a74986a  and  a74973a );
 a960a <=( a74960a  and  a74947a );
 a961a <=( a74934a  and  a74921a );
 a962a <=( a74908a  and  a74895a );
 a963a <=( a74882a  and  a74869a );
 a964a <=( a74856a  and  a74843a );
 a965a <=( a74830a  and  a74817a );
 a966a <=( a74804a  and  a74791a );
 a967a <=( a74778a  and  a74765a );
 a968a <=( a74752a  and  a74739a );
 a969a <=( a74726a  and  a74713a );
 a970a <=( a74700a  and  a74687a );
 a971a <=( a74674a  and  a74661a );
 a972a <=( a74648a  and  a74635a );
 a973a <=( a74622a  and  a74609a );
 a974a <=( a74596a  and  a74583a );
 a975a <=( a74570a  and  a74557a );
 a976a <=( a74544a  and  a74531a );
 a977a <=( a74518a  and  a74505a );
 a978a <=( a74492a  and  a74479a );
 a979a <=( a74466a  and  a74453a );
 a980a <=( a74440a  and  a74427a );
 a981a <=( a74414a  and  a74401a );
 a982a <=( a74388a  and  a74375a );
 a983a <=( a74362a  and  a74349a );
 a984a <=( a74336a  and  a74323a );
 a985a <=( a74310a  and  a74297a );
 a986a <=( a74284a  and  a74271a );
 a987a <=( a74258a  and  a74245a );
 a988a <=( a74232a  and  a74219a );
 a989a <=( a74206a  and  a74193a );
 a990a <=( a74180a  and  a74167a );
 a991a <=( a74154a  and  a74141a );
 a992a <=( a74128a  and  a74115a );
 a993a <=( a74102a  and  a74089a );
 a994a <=( a74076a  and  a74063a );
 a995a <=( a74050a  and  a74037a );
 a996a <=( a74024a  and  a74011a );
 a997a <=( a73998a  and  a73985a );
 a998a <=( a73972a  and  a73959a );
 a999a <=( a73946a  and  a73933a );
 a1000a <=( a73920a  and  a73907a );
 a1001a <=( a73894a  and  a73881a );
 a1002a <=( a73868a  and  a73855a );
 a1003a <=( a73842a  and  a73829a );
 a1004a <=( a73816a  and  a73803a );
 a1005a <=( a73790a  and  a73777a );
 a1006a <=( a73764a  and  a73751a );
 a1007a <=( a73738a  and  a73725a );
 a1008a <=( a73712a  and  a73699a );
 a1009a <=( a73686a  and  a73673a );
 a1010a <=( a73660a  and  a73647a );
 a1011a <=( a73634a  and  a73621a );
 a1012a <=( a73608a  and  a73595a );
 a1013a <=( a73582a  and  a73569a );
 a1014a <=( a73556a  and  a73543a );
 a1015a <=( a73530a  and  a73517a );
 a1016a <=( a73504a  and  a73491a );
 a1017a <=( a73478a  and  a73465a );
 a1018a <=( a73452a  and  a73439a );
 a1019a <=( a73426a  and  a73413a );
 a1020a <=( a73400a  and  a73387a );
 a1021a <=( a73374a  and  a73361a );
 a1022a <=( a73348a  and  a73335a );
 a1023a <=( a73322a  and  a73309a );
 a1024a <=( a73296a  and  a73283a );
 a1025a <=( a73270a  and  a73257a );
 a1026a <=( a73244a  and  a73231a );
 a1027a <=( a73218a  and  a73205a );
 a1028a <=( a73192a  and  a73179a );
 a1029a <=( a73166a  and  a73153a );
 a1030a <=( a73140a  and  a73127a );
 a1031a <=( a73114a  and  a73101a );
 a1032a <=( a73088a  and  a73075a );
 a1033a <=( a73062a  and  a73049a );
 a1034a <=( a73036a  and  a73023a );
 a1035a <=( a73010a  and  a72997a );
 a1036a <=( a72984a  and  a72971a );
 a1037a <=( a72958a  and  a72945a );
 a1038a <=( a72932a  and  a72919a );
 a1039a <=( a72906a  and  a72893a );
 a1040a <=( a72880a  and  a72867a );
 a1041a <=( a72854a  and  a72841a );
 a1042a <=( a72828a  and  a72815a );
 a1043a <=( a72802a  and  a72789a );
 a1044a <=( a72776a  and  a72763a );
 a1045a <=( a72750a  and  a72737a );
 a1046a <=( a72724a  and  a72711a );
 a1047a <=( a72698a  and  a72685a );
 a1048a <=( a72672a  and  a72659a );
 a1049a <=( a72646a  and  a72633a );
 a1050a <=( a72620a  and  a72607a );
 a1051a <=( a72594a  and  a72581a );
 a1052a <=( a72568a  and  a72555a );
 a1053a <=( a72542a  and  a72529a );
 a1054a <=( a72516a  and  a72503a );
 a1055a <=( a72490a  and  a72477a );
 a1056a <=( a72464a  and  a72451a );
 a1057a <=( a72438a  and  a72425a );
 a1058a <=( a72412a  and  a72399a );
 a1059a <=( a72386a  and  a72373a );
 a1060a <=( a72360a  and  a72347a );
 a1061a <=( a72334a  and  a72321a );
 a1062a <=( a72308a  and  a72295a );
 a1063a <=( a72282a  and  a72269a );
 a1064a <=( a72256a  and  a72243a );
 a1065a <=( a72230a  and  a72217a );
 a1066a <=( a72204a  and  a72191a );
 a1067a <=( a72178a  and  a72165a );
 a1068a <=( a72152a  and  a72139a );
 a1069a <=( a72126a  and  a72113a );
 a1070a <=( a72100a  and  a72087a );
 a1071a <=( a72074a  and  a72061a );
 a1072a <=( a72048a  and  a72035a );
 a1073a <=( a72022a  and  a72009a );
 a1074a <=( a71996a  and  a71983a );
 a1075a <=( a71970a  and  a71957a );
 a1076a <=( a71944a  and  a71931a );
 a1077a <=( a71918a  and  a71905a );
 a1078a <=( a71892a  and  a71879a );
 a1079a <=( a71866a  and  a71853a );
 a1080a <=( a71840a  and  a71827a );
 a1081a <=( a71814a  and  a71801a );
 a1082a <=( a71788a  and  a71775a );
 a1083a <=( a71762a  and  a71749a );
 a1084a <=( a71736a  and  a71723a );
 a1085a <=( a71710a  and  a71697a );
 a1086a <=( a71684a  and  a71671a );
 a1087a <=( a71658a  and  a71645a );
 a1088a <=( a71632a  and  a71619a );
 a1089a <=( a71606a  and  a71593a );
 a1090a <=( a71580a  and  a71567a );
 a1091a <=( a71554a  and  a71541a );
 a1092a <=( a71528a  and  a71515a );
 a1093a <=( a71502a  and  a71489a );
 a1094a <=( a71476a  and  a71463a );
 a1095a <=( a71450a  and  a71437a );
 a1096a <=( a71424a  and  a71411a );
 a1097a <=( a71398a  and  a71385a );
 a1098a <=( a71372a  and  a71359a );
 a1099a <=( a71346a  and  a71333a );
 a1100a <=( a71320a  and  a71307a );
 a1101a <=( a71294a  and  a71281a );
 a1102a <=( a71268a  and  a71255a );
 a1103a <=( a71242a  and  a71229a );
 a1104a <=( a71216a  and  a71203a );
 a1105a <=( a71190a  and  a71177a );
 a1106a <=( a71164a  and  a71151a );
 a1107a <=( a71138a  and  a71125a );
 a1108a <=( a71112a  and  a71099a );
 a1109a <=( a71086a  and  a71073a );
 a1110a <=( a71060a  and  a71047a );
 a1111a <=( a71034a  and  a71021a );
 a1112a <=( a71008a  and  a70995a );
 a1113a <=( a70982a  and  a70969a );
 a1114a <=( a70956a  and  a70943a );
 a1115a <=( a70930a  and  a70917a );
 a1116a <=( a70904a  and  a70891a );
 a1117a <=( a70878a  and  a70865a );
 a1118a <=( a70852a  and  a70839a );
 a1119a <=( a70826a  and  a70813a );
 a1120a <=( a70800a  and  a70787a );
 a1121a <=( a70774a  and  a70761a );
 a1122a <=( a70748a  and  a70735a );
 a1123a <=( a70722a  and  a70709a );
 a1124a <=( a70696a  and  a70683a );
 a1125a <=( a70670a  and  a70657a );
 a1126a <=( a70644a  and  a70631a );
 a1127a <=( a70618a  and  a70605a );
 a1128a <=( a70592a  and  a70579a );
 a1129a <=( a70566a  and  a70553a );
 a1130a <=( a70540a  and  a70527a );
 a1131a <=( a70514a  and  a70501a );
 a1132a <=( a70488a  and  a70475a );
 a1133a <=( a70462a  and  a70449a );
 a1134a <=( a70436a  and  a70423a );
 a1135a <=( a70410a  and  a70397a );
 a1136a <=( a70384a  and  a70371a );
 a1137a <=( a70358a  and  a70345a );
 a1138a <=( a70332a  and  a70319a );
 a1139a <=( a70306a  and  a70293a );
 a1140a <=( a70280a  and  a70267a );
 a1141a <=( a70254a  and  a70241a );
 a1142a <=( a70228a  and  a70215a );
 a1143a <=( a70202a  and  a70189a );
 a1144a <=( a70176a  and  a70163a );
 a1145a <=( a70150a  and  a70137a );
 a1146a <=( a70124a  and  a70111a );
 a1147a <=( a70098a  and  a70085a );
 a1148a <=( a70072a  and  a70059a );
 a1149a <=( a70046a  and  a70033a );
 a1150a <=( a70020a  and  a70007a );
 a1151a <=( a69994a  and  a69981a );
 a1152a <=( a69968a  and  a69955a );
 a1153a <=( a69942a  and  a69929a );
 a1154a <=( a69916a  and  a69903a );
 a1155a <=( a69890a  and  a69877a );
 a1156a <=( a69864a  and  a69851a );
 a1157a <=( a69838a  and  a69825a );
 a1158a <=( a69812a  and  a69799a );
 a1159a <=( a69786a  and  a69773a );
 a1160a <=( a69760a  and  a69747a );
 a1161a <=( a69734a  and  a69721a );
 a1162a <=( a69708a  and  a69695a );
 a1163a <=( a69682a  and  a69669a );
 a1164a <=( a69656a  and  a69643a );
 a1165a <=( a69630a  and  a69617a );
 a1166a <=( a69604a  and  a69591a );
 a1167a <=( a69578a  and  a69565a );
 a1168a <=( a69552a  and  a69539a );
 a1169a <=( a69526a  and  a69513a );
 a1170a <=( a69500a  and  a69487a );
 a1171a <=( a69474a  and  a69461a );
 a1172a <=( a69448a  and  a69435a );
 a1173a <=( a69422a  and  a69409a );
 a1174a <=( a69396a  and  a69383a );
 a1175a <=( a69370a  and  a69357a );
 a1176a <=( a69344a  and  a69331a );
 a1177a <=( a69318a  and  a69305a );
 a1178a <=( a69292a  and  a69279a );
 a1179a <=( a69266a  and  a69253a );
 a1180a <=( a69240a  and  a69227a );
 a1181a <=( a69214a  and  a69201a );
 a1182a <=( a69188a  and  a69175a );
 a1183a <=( a69162a  and  a69149a );
 a1184a <=( a69136a  and  a69123a );
 a1185a <=( a69110a  and  a69097a );
 a1186a <=( a69084a  and  a69071a );
 a1187a <=( a69058a  and  a69045a );
 a1188a <=( a69032a  and  a69019a );
 a1189a <=( a69006a  and  a68993a );
 a1190a <=( a68980a  and  a68967a );
 a1191a <=( a68954a  and  a68941a );
 a1192a <=( a68928a  and  a68915a );
 a1193a <=( a68902a  and  a68889a );
 a1194a <=( a68876a  and  a68863a );
 a1195a <=( a68850a  and  a68837a );
 a1196a <=( a68824a  and  a68811a );
 a1197a <=( a68798a  and  a68785a );
 a1198a <=( a68772a  and  a68759a );
 a1199a <=( a68746a  and  a68733a );
 a1200a <=( a68720a  and  a68707a );
 a1201a <=( a68694a  and  a68681a );
 a1202a <=( a68668a  and  a68655a );
 a1203a <=( a68642a  and  a68629a );
 a1204a <=( a68616a  and  a68603a );
 a1205a <=( a68590a  and  a68577a );
 a1206a <=( a68564a  and  a68551a );
 a1207a <=( a68538a  and  a68525a );
 a1208a <=( a68512a  and  a68499a );
 a1209a <=( a68486a  and  a68473a );
 a1210a <=( a68460a  and  a68447a );
 a1211a <=( a68434a  and  a68421a );
 a1212a <=( a68408a  and  a68395a );
 a1213a <=( a68382a  and  a68369a );
 a1214a <=( a68356a  and  a68343a );
 a1215a <=( a68330a  and  a68317a );
 a1216a <=( a68304a  and  a68291a );
 a1217a <=( a68278a  and  a68265a );
 a1218a <=( a68252a  and  a68239a );
 a1219a <=( a68226a  and  a68213a );
 a1220a <=( a68200a  and  a68187a );
 a1221a <=( a68174a  and  a68161a );
 a1222a <=( a68148a  and  a68135a );
 a1223a <=( a68122a  and  a68109a );
 a1224a <=( a68096a  and  a68083a );
 a1225a <=( a68070a  and  a68057a );
 a1226a <=( a68044a  and  a68031a );
 a1227a <=( a68018a  and  a68005a );
 a1228a <=( a67992a  and  a67979a );
 a1229a <=( a67966a  and  a67953a );
 a1230a <=( a67940a  and  a67927a );
 a1231a <=( a67914a  and  a67901a );
 a1232a <=( a67888a  and  a67875a );
 a1233a <=( a67862a  and  a67849a );
 a1234a <=( a67836a  and  a67823a );
 a1235a <=( a67810a  and  a67797a );
 a1236a <=( a67784a  and  a67771a );
 a1237a <=( a67758a  and  a67745a );
 a1238a <=( a67732a  and  a67719a );
 a1239a <=( a67706a  and  a67693a );
 a1240a <=( a67680a  and  a67667a );
 a1241a <=( a67654a  and  a67641a );
 a1242a <=( a67628a  and  a67615a );
 a1243a <=( a67602a  and  a67589a );
 a1244a <=( a67576a  and  a67563a );
 a1245a <=( a67550a  and  a67537a );
 a1246a <=( a67524a  and  a67511a );
 a1247a <=( a67498a  and  a67485a );
 a1248a <=( a67472a  and  a67459a );
 a1249a <=( a67446a  and  a67433a );
 a1250a <=( a67420a  and  a67407a );
 a1251a <=( a67394a  and  a67381a );
 a1252a <=( a67368a  and  a67355a );
 a1253a <=( a67342a  and  a67329a );
 a1254a <=( a67316a  and  a67303a );
 a1255a <=( a67290a  and  a67277a );
 a1256a <=( a67264a  and  a67251a );
 a1257a <=( a67238a  and  a67225a );
 a1258a <=( a67212a  and  a67199a );
 a1259a <=( a67186a  and  a67173a );
 a1260a <=( a67160a  and  a67147a );
 a1261a <=( a67134a  and  a67121a );
 a1262a <=( a67108a  and  a67095a );
 a1263a <=( a67082a  and  a67069a );
 a1264a <=( a67056a  and  a67043a );
 a1265a <=( a67030a  and  a67017a );
 a1266a <=( a67004a  and  a66991a );
 a1267a <=( a66978a  and  a66965a );
 a1268a <=( a66952a  and  a66939a );
 a1269a <=( a66926a  and  a66913a );
 a1270a <=( a66900a  and  a66887a );
 a1271a <=( a66874a  and  a66861a );
 a1272a <=( a66848a  and  a66835a );
 a1273a <=( a66822a  and  a66809a );
 a1274a <=( a66796a  and  a66783a );
 a1275a <=( a66770a  and  a66757a );
 a1276a <=( a66744a  and  a66731a );
 a1277a <=( a66718a  and  a66705a );
 a1278a <=( a66692a  and  a66679a );
 a1279a <=( a66666a  and  a66653a );
 a1280a <=( a66640a  and  a66627a );
 a1281a <=( a66614a  and  a66601a );
 a1282a <=( a66588a  and  a66575a );
 a1283a <=( a66562a  and  a66549a );
 a1284a <=( a66536a  and  a66523a );
 a1285a <=( a66510a  and  a66497a );
 a1286a <=( a66484a  and  a66471a );
 a1287a <=( a66458a  and  a66445a );
 a1288a <=( a66432a  and  a66419a );
 a1289a <=( a66406a  and  a66393a );
 a1290a <=( a66380a  and  a66367a );
 a1291a <=( a66354a  and  a66341a );
 a1292a <=( a66328a  and  a66315a );
 a1293a <=( a66302a  and  a66289a );
 a1294a <=( a66276a  and  a66263a );
 a1295a <=( a66250a  and  a66237a );
 a1296a <=( a66224a  and  a66211a );
 a1297a <=( a66198a  and  a66185a );
 a1298a <=( a66172a  and  a66159a );
 a1299a <=( a66146a  and  a66133a );
 a1300a <=( a66120a  and  a66107a );
 a1301a <=( a66094a  and  a66081a );
 a1302a <=( a66068a  and  a66055a );
 a1303a <=( a66042a  and  a66029a );
 a1304a <=( a66016a  and  a66003a );
 a1305a <=( a65990a  and  a65977a );
 a1306a <=( a65964a  and  a65951a );
 a1307a <=( a65938a  and  a65925a );
 a1308a <=( a65912a  and  a65899a );
 a1309a <=( a65886a  and  a65873a );
 a1310a <=( a65860a  and  a65847a );
 a1311a <=( a65834a  and  a65821a );
 a1312a <=( a65808a  and  a65795a );
 a1313a <=( a65782a  and  a65769a );
 a1314a <=( a65756a  and  a65743a );
 a1315a <=( a65730a  and  a65717a );
 a1316a <=( a65704a  and  a65691a );
 a1317a <=( a65678a  and  a65665a );
 a1318a <=( a65652a  and  a65639a );
 a1319a <=( a65626a  and  a65613a );
 a1320a <=( a65600a  and  a65587a );
 a1321a <=( a65574a  and  a65561a );
 a1322a <=( a65548a  and  a65535a );
 a1323a <=( a65522a  and  a65509a );
 a1324a <=( a65496a  and  a65483a );
 a1325a <=( a65470a  and  a65457a );
 a1326a <=( a65444a  and  a65431a );
 a1327a <=( a65418a  and  a65405a );
 a1328a <=( a65392a  and  a65379a );
 a1329a <=( a65366a  and  a65353a );
 a1330a <=( a65340a  and  a65327a );
 a1331a <=( a65314a  and  a65301a );
 a1332a <=( a65288a  and  a65275a );
 a1333a <=( a65262a  and  a65249a );
 a1334a <=( a65236a  and  a65223a );
 a1335a <=( a65210a  and  a65197a );
 a1336a <=( a65184a  and  a65171a );
 a1337a <=( a65158a  and  a65145a );
 a1338a <=( a65132a  and  a65119a );
 a1339a <=( a65106a  and  a65093a );
 a1340a <=( a65080a  and  a65067a );
 a1341a <=( a65054a  and  a65041a );
 a1342a <=( a65028a  and  a65015a );
 a1343a <=( a65002a  and  a64989a );
 a1344a <=( a64976a  and  a64963a );
 a1345a <=( a64950a  and  a64937a );
 a1346a <=( a64924a  and  a64911a );
 a1347a <=( a64898a  and  a64885a );
 a1348a <=( a64872a  and  a64859a );
 a1349a <=( a64846a  and  a64833a );
 a1350a <=( a64820a  and  a64807a );
 a1351a <=( a64794a  and  a64781a );
 a1352a <=( a64768a  and  a64755a );
 a1353a <=( a64742a  and  a64729a );
 a1354a <=( a64716a  and  a64703a );
 a1355a <=( a64690a  and  a64677a );
 a1356a <=( a64664a  and  a64651a );
 a1357a <=( a64638a  and  a64625a );
 a1358a <=( a64614a  and  a64601a );
 a1359a <=( a64590a  and  a64577a );
 a1360a <=( a64566a  and  a64553a );
 a1361a <=( a64542a  and  a64529a );
 a1362a <=( a64518a  and  a64505a );
 a1363a <=( a64494a  and  a64481a );
 a1364a <=( a64470a  and  a64457a );
 a1365a <=( a64446a  and  a64433a );
 a1366a <=( a64422a  and  a64409a );
 a1367a <=( a64398a  and  a64385a );
 a1368a <=( a64374a  and  a64361a );
 a1369a <=( a64350a  and  a64337a );
 a1370a <=( a64326a  and  a64313a );
 a1371a <=( a64302a  and  a64289a );
 a1372a <=( a64278a  and  a64265a );
 a1373a <=( a64254a  and  a64241a );
 a1374a <=( a64230a  and  a64217a );
 a1375a <=( a64206a  and  a64193a );
 a1376a <=( a64182a  and  a64169a );
 a1377a <=( a64158a  and  a64145a );
 a1378a <=( a64134a  and  a64121a );
 a1379a <=( a64110a  and  a64097a );
 a1380a <=( a64086a  and  a64073a );
 a1381a <=( a64062a  and  a64049a );
 a1382a <=( a64038a  and  a64025a );
 a1383a <=( a64014a  and  a64001a );
 a1384a <=( a63990a  and  a63977a );
 a1385a <=( a63966a  and  a63953a );
 a1386a <=( a63942a  and  a63929a );
 a1387a <=( a63918a  and  a63905a );
 a1388a <=( a63894a  and  a63881a );
 a1389a <=( a63870a  and  a63857a );
 a1390a <=( a63846a  and  a63833a );
 a1391a <=( a63822a  and  a63809a );
 a1392a <=( a63798a  and  a63785a );
 a1393a <=( a63774a  and  a63761a );
 a1394a <=( a63750a  and  a63737a );
 a1395a <=( a63726a  and  a63713a );
 a1396a <=( a63702a  and  a63689a );
 a1397a <=( a63678a  and  a63665a );
 a1398a <=( a63654a  and  a63641a );
 a1399a <=( a63630a  and  a63617a );
 a1400a <=( a63606a  and  a63593a );
 a1401a <=( a63582a  and  a63569a );
 a1402a <=( a63558a  and  a63545a );
 a1403a <=( a63534a  and  a63521a );
 a1404a <=( a63510a  and  a63497a );
 a1405a <=( a63486a  and  a63473a );
 a1406a <=( a63462a  and  a63449a );
 a1407a <=( a63438a  and  a63425a );
 a1408a <=( a63414a  and  a63401a );
 a1409a <=( a63390a  and  a63377a );
 a1410a <=( a63366a  and  a63353a );
 a1411a <=( a63342a  and  a63329a );
 a1412a <=( a63318a  and  a63305a );
 a1413a <=( a63294a  and  a63281a );
 a1414a <=( a63270a  and  a63257a );
 a1415a <=( a63246a  and  a63233a );
 a1416a <=( a63222a  and  a63209a );
 a1417a <=( a63198a  and  a63185a );
 a1418a <=( a63174a  and  a63161a );
 a1419a <=( a63150a  and  a63137a );
 a1420a <=( a63126a  and  a63113a );
 a1421a <=( a63102a  and  a63089a );
 a1422a <=( a63078a  and  a63065a );
 a1423a <=( a63054a  and  a63041a );
 a1424a <=( a63030a  and  a63017a );
 a1425a <=( a63006a  and  a62993a );
 a1426a <=( a62982a  and  a62969a );
 a1427a <=( a62958a  and  a62945a );
 a1428a <=( a62934a  and  a62921a );
 a1429a <=( a62910a  and  a62897a );
 a1430a <=( a62886a  and  a62873a );
 a1431a <=( a62862a  and  a62849a );
 a1432a <=( a62838a  and  a62825a );
 a1433a <=( a62814a  and  a62801a );
 a1434a <=( a62790a  and  a62777a );
 a1435a <=( a62766a  and  a62753a );
 a1436a <=( a62742a  and  a62729a );
 a1437a <=( a62718a  and  a62705a );
 a1438a <=( a62694a  and  a62681a );
 a1439a <=( a62670a  and  a62657a );
 a1440a <=( a62646a  and  a62633a );
 a1441a <=( a62622a  and  a62609a );
 a1442a <=( a62598a  and  a62585a );
 a1443a <=( a62574a  and  a62561a );
 a1444a <=( a62550a  and  a62537a );
 a1445a <=( a62526a  and  a62513a );
 a1446a <=( a62502a  and  a62489a );
 a1447a <=( a62478a  and  a62465a );
 a1448a <=( a62454a  and  a62441a );
 a1449a <=( a62430a  and  a62417a );
 a1450a <=( a62406a  and  a62393a );
 a1451a <=( a62382a  and  a62369a );
 a1452a <=( a62358a  and  a62345a );
 a1453a <=( a62334a  and  a62321a );
 a1454a <=( a62310a  and  a62297a );
 a1455a <=( a62286a  and  a62273a );
 a1456a <=( a62262a  and  a62249a );
 a1457a <=( a62238a  and  a62225a );
 a1458a <=( a62214a  and  a62201a );
 a1459a <=( a62190a  and  a62177a );
 a1460a <=( a62166a  and  a62153a );
 a1461a <=( a62142a  and  a62129a );
 a1462a <=( a62118a  and  a62105a );
 a1463a <=( a62094a  and  a62081a );
 a1464a <=( a62070a  and  a62057a );
 a1465a <=( a62046a  and  a62033a );
 a1466a <=( a62022a  and  a62009a );
 a1467a <=( a61998a  and  a61985a );
 a1468a <=( a61974a  and  a61961a );
 a1469a <=( a61950a  and  a61937a );
 a1470a <=( a61926a  and  a61913a );
 a1471a <=( a61902a  and  a61889a );
 a1472a <=( a61878a  and  a61865a );
 a1473a <=( a61854a  and  a61841a );
 a1474a <=( a61830a  and  a61817a );
 a1475a <=( a61806a  and  a61793a );
 a1476a <=( a61782a  and  a61769a );
 a1477a <=( a61758a  and  a61745a );
 a1478a <=( a61734a  and  a61721a );
 a1479a <=( a61710a  and  a61697a );
 a1480a <=( a61686a  and  a61673a );
 a1481a <=( a61662a  and  a61649a );
 a1482a <=( a61638a  and  a61625a );
 a1483a <=( a61614a  and  a61601a );
 a1484a <=( a61590a  and  a61577a );
 a1485a <=( a61566a  and  a61553a );
 a1486a <=( a61542a  and  a61529a );
 a1487a <=( a61518a  and  a61505a );
 a1488a <=( a61494a  and  a61481a );
 a1489a <=( a61470a  and  a61457a );
 a1490a <=( a61446a  and  a61433a );
 a1491a <=( a61422a  and  a61409a );
 a1492a <=( a61398a  and  a61385a );
 a1493a <=( a61374a  and  a61361a );
 a1494a <=( a61350a  and  a61337a );
 a1495a <=( a61326a  and  a61313a );
 a1496a <=( a61302a  and  a61289a );
 a1497a <=( a61278a  and  a61265a );
 a1498a <=( a61254a  and  a61241a );
 a1499a <=( a61230a  and  a61217a );
 a1500a <=( a61206a  and  a61193a );
 a1501a <=( a61182a  and  a61169a );
 a1502a <=( a61158a  and  a61145a );
 a1503a <=( a61134a  and  a61121a );
 a1504a <=( a61110a  and  a61097a );
 a1505a <=( a61086a  and  a61073a );
 a1506a <=( a61062a  and  a61049a );
 a1507a <=( a61038a  and  a61025a );
 a1508a <=( a61014a  and  a61001a );
 a1509a <=( a60990a  and  a60977a );
 a1510a <=( a60966a  and  a60953a );
 a1511a <=( a60942a  and  a60929a );
 a1512a <=( a60918a  and  a60905a );
 a1513a <=( a60894a  and  a60881a );
 a1514a <=( a60870a  and  a60857a );
 a1515a <=( a60846a  and  a60833a );
 a1516a <=( a60822a  and  a60809a );
 a1517a <=( a60798a  and  a60785a );
 a1518a <=( a60774a  and  a60761a );
 a1519a <=( a60750a  and  a60737a );
 a1520a <=( a60726a  and  a60713a );
 a1521a <=( a60702a  and  a60689a );
 a1522a <=( a60678a  and  a60665a );
 a1523a <=( a60654a  and  a60641a );
 a1524a <=( a60630a  and  a60617a );
 a1525a <=( a60606a  and  a60593a );
 a1526a <=( a60582a  and  a60569a );
 a1527a <=( a60558a  and  a60545a );
 a1528a <=( a60534a  and  a60521a );
 a1529a <=( a60510a  and  a60497a );
 a1530a <=( a60486a  and  a60473a );
 a1531a <=( a60462a  and  a60449a );
 a1532a <=( a60438a  and  a60425a );
 a1533a <=( a60414a  and  a60401a );
 a1534a <=( a60390a  and  a60377a );
 a1535a <=( a60366a  and  a60353a );
 a1536a <=( a60342a  and  a60329a );
 a1537a <=( a60318a  and  a60305a );
 a1538a <=( a60294a  and  a60281a );
 a1539a <=( a60270a  and  a60257a );
 a1540a <=( a60246a  and  a60233a );
 a1541a <=( a60222a  and  a60209a );
 a1542a <=( a60198a  and  a60185a );
 a1543a <=( a60174a  and  a60161a );
 a1544a <=( a60150a  and  a60137a );
 a1545a <=( a60126a  and  a60113a );
 a1546a <=( a60102a  and  a60089a );
 a1547a <=( a60078a  and  a60065a );
 a1548a <=( a60054a  and  a60041a );
 a1549a <=( a60030a  and  a60017a );
 a1550a <=( a60006a  and  a59993a );
 a1551a <=( a59982a  and  a59969a );
 a1552a <=( a59958a  and  a59945a );
 a1553a <=( a59934a  and  a59921a );
 a1554a <=( a59910a  and  a59897a );
 a1555a <=( a59886a  and  a59873a );
 a1556a <=( a59862a  and  a59849a );
 a1557a <=( a59838a  and  a59825a );
 a1558a <=( a59814a  and  a59801a );
 a1559a <=( a59790a  and  a59777a );
 a1560a <=( a59766a  and  a59753a );
 a1561a <=( a59742a  and  a59729a );
 a1562a <=( a59718a  and  a59705a );
 a1563a <=( a59694a  and  a59681a );
 a1564a <=( a59670a  and  a59657a );
 a1565a <=( a59646a  and  a59633a );
 a1566a <=( a59622a  and  a59609a );
 a1567a <=( a59598a  and  a59585a );
 a1568a <=( a59574a  and  a59561a );
 a1569a <=( a59550a  and  a59537a );
 a1570a <=( a59526a  and  a59513a );
 a1571a <=( a59502a  and  a59489a );
 a1572a <=( a59478a  and  a59465a );
 a1573a <=( a59454a  and  a59441a );
 a1574a <=( a59430a  and  a59417a );
 a1575a <=( a59406a  and  a59393a );
 a1576a <=( a59382a  and  a59369a );
 a1577a <=( a59358a  and  a59345a );
 a1578a <=( a59334a  and  a59321a );
 a1579a <=( a59310a  and  a59297a );
 a1580a <=( a59286a  and  a59273a );
 a1581a <=( a59262a  and  a59249a );
 a1582a <=( a59238a  and  a59225a );
 a1583a <=( a59214a  and  a59201a );
 a1584a <=( a59190a  and  a59177a );
 a1585a <=( a59166a  and  a59153a );
 a1586a <=( a59142a  and  a59129a );
 a1587a <=( a59118a  and  a59105a );
 a1588a <=( a59094a  and  a59081a );
 a1589a <=( a59070a  and  a59057a );
 a1590a <=( a59046a  and  a59033a );
 a1591a <=( a59022a  and  a59009a );
 a1592a <=( a58998a  and  a58985a );
 a1593a <=( a58974a  and  a58961a );
 a1594a <=( a58950a  and  a58937a );
 a1595a <=( a58926a  and  a58913a );
 a1596a <=( a58902a  and  a58889a );
 a1597a <=( a58878a  and  a58865a );
 a1598a <=( a58854a  and  a58841a );
 a1599a <=( a58830a  and  a58817a );
 a1600a <=( a58806a  and  a58793a );
 a1601a <=( a58782a  and  a58769a );
 a1602a <=( a58758a  and  a58745a );
 a1603a <=( a58734a  and  a58721a );
 a1604a <=( a58710a  and  a58697a );
 a1605a <=( a58686a  and  a58673a );
 a1606a <=( a58662a  and  a58649a );
 a1607a <=( a58638a  and  a58625a );
 a1608a <=( a58614a  and  a58601a );
 a1609a <=( a58590a  and  a58577a );
 a1610a <=( a58566a  and  a58553a );
 a1611a <=( a58542a  and  a58529a );
 a1612a <=( a58518a  and  a58505a );
 a1613a <=( a58494a  and  a58481a );
 a1614a <=( a58470a  and  a58457a );
 a1615a <=( a58446a  and  a58433a );
 a1616a <=( a58422a  and  a58409a );
 a1617a <=( a58398a  and  a58385a );
 a1618a <=( a58374a  and  a58361a );
 a1619a <=( a58350a  and  a58337a );
 a1620a <=( a58326a  and  a58313a );
 a1621a <=( a58302a  and  a58289a );
 a1622a <=( a58278a  and  a58265a );
 a1623a <=( a58254a  and  a58241a );
 a1624a <=( a58230a  and  a58217a );
 a1625a <=( a58206a  and  a58193a );
 a1626a <=( a58182a  and  a58169a );
 a1627a <=( a58158a  and  a58145a );
 a1628a <=( a58134a  and  a58121a );
 a1629a <=( a58110a  and  a58097a );
 a1630a <=( a58086a  and  a58073a );
 a1631a <=( a58062a  and  a58049a );
 a1632a <=( a58038a  and  a58025a );
 a1633a <=( a58014a  and  a58001a );
 a1634a <=( a57990a  and  a57977a );
 a1635a <=( a57966a  and  a57953a );
 a1636a <=( a57942a  and  a57929a );
 a1637a <=( a57918a  and  a57905a );
 a1638a <=( a57894a  and  a57881a );
 a1639a <=( a57870a  and  a57857a );
 a1640a <=( a57846a  and  a57833a );
 a1641a <=( a57822a  and  a57809a );
 a1642a <=( a57798a  and  a57785a );
 a1643a <=( a57774a  and  a57761a );
 a1644a <=( a57750a  and  a57737a );
 a1645a <=( a57726a  and  a57713a );
 a1646a <=( a57702a  and  a57689a );
 a1647a <=( a57678a  and  a57665a );
 a1648a <=( a57654a  and  a57641a );
 a1649a <=( a57630a  and  a57617a );
 a1650a <=( a57606a  and  a57593a );
 a1651a <=( a57582a  and  a57569a );
 a1652a <=( a57558a  and  a57545a );
 a1653a <=( a57534a  and  a57521a );
 a1654a <=( a57510a  and  a57497a );
 a1655a <=( a57486a  and  a57473a );
 a1656a <=( a57462a  and  a57449a );
 a1657a <=( a57438a  and  a57425a );
 a1658a <=( a57414a  and  a57401a );
 a1659a <=( a57390a  and  a57377a );
 a1660a <=( a57366a  and  a57353a );
 a1661a <=( a57342a  and  a57329a );
 a1662a <=( a57318a  and  a57305a );
 a1663a <=( a57294a  and  a57281a );
 a1664a <=( a57270a  and  a57257a );
 a1665a <=( a57246a  and  a57233a );
 a1666a <=( a57222a  and  a57209a );
 a1667a <=( a57198a  and  a57185a );
 a1668a <=( a57174a  and  a57161a );
 a1669a <=( a57150a  and  a57137a );
 a1670a <=( a57126a  and  a57113a );
 a1671a <=( a57102a  and  a57089a );
 a1672a <=( a57078a  and  a57065a );
 a1673a <=( a57054a  and  a57041a );
 a1674a <=( a57030a  and  a57017a );
 a1675a <=( a57006a  and  a56993a );
 a1676a <=( a56982a  and  a56969a );
 a1677a <=( a56958a  and  a56945a );
 a1678a <=( a56934a  and  a56921a );
 a1679a <=( a56910a  and  a56897a );
 a1680a <=( a56886a  and  a56873a );
 a1681a <=( a56862a  and  a56849a );
 a1682a <=( a56838a  and  a56825a );
 a1683a <=( a56814a  and  a56801a );
 a1684a <=( a56790a  and  a56777a );
 a1685a <=( a56766a  and  a56753a );
 a1686a <=( a56742a  and  a56729a );
 a1687a <=( a56718a  and  a56705a );
 a1688a <=( a56694a  and  a56681a );
 a1689a <=( a56670a  and  a56657a );
 a1690a <=( a56646a  and  a56633a );
 a1691a <=( a56622a  and  a56609a );
 a1692a <=( a56598a  and  a56585a );
 a1693a <=( a56574a  and  a56561a );
 a1694a <=( a56550a  and  a56537a );
 a1695a <=( a56526a  and  a56513a );
 a1696a <=( a56502a  and  a56489a );
 a1697a <=( a56478a  and  a56465a );
 a1698a <=( a56454a  and  a56441a );
 a1699a <=( a56430a  and  a56417a );
 a1700a <=( a56406a  and  a56393a );
 a1701a <=( a56382a  and  a56369a );
 a1702a <=( a56358a  and  a56345a );
 a1703a <=( a56334a  and  a56321a );
 a1704a <=( a56310a  and  a56297a );
 a1705a <=( a56286a  and  a56273a );
 a1706a <=( a56262a  and  a56249a );
 a1707a <=( a56238a  and  a56225a );
 a1708a <=( a56214a  and  a56201a );
 a1709a <=( a56190a  and  a56177a );
 a1710a <=( a56166a  and  a56153a );
 a1711a <=( a56142a  and  a56129a );
 a1712a <=( a56118a  and  a56105a );
 a1713a <=( a56094a  and  a56081a );
 a1714a <=( a56070a  and  a56057a );
 a1715a <=( a56046a  and  a56033a );
 a1716a <=( a56022a  and  a56009a );
 a1717a <=( a55998a  and  a55985a );
 a1718a <=( a55974a  and  a55961a );
 a1719a <=( a55950a  and  a55937a );
 a1720a <=( a55926a  and  a55913a );
 a1721a <=( a55902a  and  a55889a );
 a1722a <=( a55878a  and  a55865a );
 a1723a <=( a55854a  and  a55841a );
 a1724a <=( a55830a  and  a55817a );
 a1725a <=( a55806a  and  a55793a );
 a1726a <=( a55782a  and  a55769a );
 a1727a <=( a55758a  and  a55745a );
 a1728a <=( a55734a  and  a55721a );
 a1729a <=( a55710a  and  a55697a );
 a1730a <=( a55686a  and  a55673a );
 a1731a <=( a55662a  and  a55649a );
 a1732a <=( a55638a  and  a55625a );
 a1733a <=( a55614a  and  a55601a );
 a1734a <=( a55590a  and  a55577a );
 a1735a <=( a55566a  and  a55553a );
 a1736a <=( a55542a  and  a55529a );
 a1737a <=( a55518a  and  a55505a );
 a1738a <=( a55494a  and  a55481a );
 a1739a <=( a55470a  and  a55457a );
 a1740a <=( a55446a  and  a55433a );
 a1741a <=( a55422a  and  a55409a );
 a1742a <=( a55398a  and  a55385a );
 a1743a <=( a55374a  and  a55361a );
 a1744a <=( a55350a  and  a55337a );
 a1745a <=( a55326a  and  a55313a );
 a1746a <=( a55302a  and  a55289a );
 a1747a <=( a55278a  and  a55265a );
 a1748a <=( a55254a  and  a55241a );
 a1749a <=( a55230a  and  a55217a );
 a1750a <=( a55206a  and  a55193a );
 a1751a <=( a55182a  and  a55169a );
 a1752a <=( a55158a  and  a55145a );
 a1753a <=( a55134a  and  a55121a );
 a1754a <=( a55110a  and  a55097a );
 a1755a <=( a55086a  and  a55073a );
 a1756a <=( a55062a  and  a55049a );
 a1757a <=( a55038a  and  a55025a );
 a1758a <=( a55014a  and  a55001a );
 a1759a <=( a54990a  and  a54977a );
 a1760a <=( a54966a  and  a54953a );
 a1761a <=( a54942a  and  a54929a );
 a1762a <=( a54918a  and  a54905a );
 a1763a <=( a54894a  and  a54881a );
 a1764a <=( a54870a  and  a54857a );
 a1765a <=( a54846a  and  a54833a );
 a1766a <=( a54822a  and  a54809a );
 a1767a <=( a54798a  and  a54785a );
 a1768a <=( a54774a  and  a54761a );
 a1769a <=( a54750a  and  a54737a );
 a1770a <=( a54726a  and  a54713a );
 a1771a <=( a54702a  and  a54689a );
 a1772a <=( a54678a  and  a54665a );
 a1773a <=( a54654a  and  a54641a );
 a1774a <=( a54630a  and  a54617a );
 a1775a <=( a54606a  and  a54593a );
 a1776a <=( a54582a  and  a54569a );
 a1777a <=( a54558a  and  a54545a );
 a1778a <=( a54534a  and  a54521a );
 a1779a <=( a54510a  and  a54497a );
 a1780a <=( a54486a  and  a54473a );
 a1781a <=( a54462a  and  a54449a );
 a1782a <=( a54438a  and  a54425a );
 a1783a <=( a54414a  and  a54401a );
 a1784a <=( a54390a  and  a54377a );
 a1785a <=( a54366a  and  a54353a );
 a1786a <=( a54342a  and  a54329a );
 a1787a <=( a54318a  and  a54305a );
 a1788a <=( a54294a  and  a54281a );
 a1789a <=( a54270a  and  a54257a );
 a1790a <=( a54246a  and  a54233a );
 a1791a <=( a54222a  and  a54209a );
 a1792a <=( a54198a  and  a54185a );
 a1793a <=( a54174a  and  a54161a );
 a1794a <=( a54150a  and  a54137a );
 a1795a <=( a54126a  and  a54113a );
 a1796a <=( a54102a  and  a54089a );
 a1797a <=( a54078a  and  a54065a );
 a1798a <=( a54054a  and  a54041a );
 a1799a <=( a54030a  and  a54017a );
 a1800a <=( a54006a  and  a53993a );
 a1801a <=( a53982a  and  a53969a );
 a1802a <=( a53958a  and  a53945a );
 a1803a <=( a53934a  and  a53921a );
 a1804a <=( a53910a  and  a53897a );
 a1805a <=( a53886a  and  a53873a );
 a1806a <=( a53862a  and  a53849a );
 a1807a <=( a53838a  and  a53825a );
 a1808a <=( a53814a  and  a53801a );
 a1809a <=( a53790a  and  a53777a );
 a1810a <=( a53766a  and  a53753a );
 a1811a <=( a53742a  and  a53729a );
 a1812a <=( a53718a  and  a53705a );
 a1813a <=( a53694a  and  a53681a );
 a1814a <=( a53670a  and  a53657a );
 a1815a <=( a53646a  and  a53633a );
 a1816a <=( a53622a  and  a53609a );
 a1817a <=( a53598a  and  a53585a );
 a1818a <=( a53574a  and  a53561a );
 a1819a <=( a53550a  and  a53537a );
 a1820a <=( a53526a  and  a53513a );
 a1821a <=( a53502a  and  a53489a );
 a1822a <=( a53478a  and  a53465a );
 a1823a <=( a53454a  and  a53441a );
 a1824a <=( a53430a  and  a53417a );
 a1825a <=( a53406a  and  a53393a );
 a1826a <=( a53382a  and  a53369a );
 a1827a <=( a53358a  and  a53345a );
 a1828a <=( a53334a  and  a53321a );
 a1829a <=( a53310a  and  a53297a );
 a1830a <=( a53286a  and  a53273a );
 a1831a <=( a53262a  and  a53249a );
 a1832a <=( a53238a  and  a53225a );
 a1833a <=( a53214a  and  a53201a );
 a1834a <=( a53190a  and  a53177a );
 a1835a <=( a53166a  and  a53153a );
 a1836a <=( a53142a  and  a53129a );
 a1837a <=( a53118a  and  a53105a );
 a1838a <=( a53094a  and  a53081a );
 a1839a <=( a53070a  and  a53057a );
 a1840a <=( a53046a  and  a53033a );
 a1841a <=( a53022a  and  a53009a );
 a1842a <=( a52998a  and  a52985a );
 a1843a <=( a52974a  and  a52961a );
 a1844a <=( a52950a  and  a52937a );
 a1845a <=( a52926a  and  a52913a );
 a1846a <=( a52902a  and  a52889a );
 a1847a <=( a52878a  and  a52865a );
 a1848a <=( a52854a  and  a52841a );
 a1849a <=( a52830a  and  a52817a );
 a1850a <=( a52806a  and  a52793a );
 a1851a <=( a52782a  and  a52769a );
 a1852a <=( a52758a  and  a52745a );
 a1853a <=( a52734a  and  a52721a );
 a1854a <=( a52710a  and  a52697a );
 a1855a <=( a52686a  and  a52673a );
 a1856a <=( a52662a  and  a52649a );
 a1857a <=( a52638a  and  a52625a );
 a1858a <=( a52614a  and  a52601a );
 a1859a <=( a52590a  and  a52577a );
 a1860a <=( a52566a  and  a52553a );
 a1861a <=( a52542a  and  a52529a );
 a1862a <=( a52518a  and  a52505a );
 a1863a <=( a52494a  and  a52481a );
 a1864a <=( a52470a  and  a52457a );
 a1865a <=( a52446a  and  a52433a );
 a1866a <=( a52422a  and  a52409a );
 a1867a <=( a52398a  and  a52385a );
 a1868a <=( a52374a  and  a52361a );
 a1869a <=( a52350a  and  a52337a );
 a1870a <=( a52326a  and  a52313a );
 a1871a <=( a52302a  and  a52289a );
 a1872a <=( a52278a  and  a52265a );
 a1873a <=( a52254a  and  a52241a );
 a1874a <=( a52230a  and  a52217a );
 a1875a <=( a52206a  and  a52193a );
 a1876a <=( a52182a  and  a52169a );
 a1877a <=( a52158a  and  a52145a );
 a1878a <=( a52134a  and  a52121a );
 a1879a <=( a52110a  and  a52097a );
 a1880a <=( a52086a  and  a52073a );
 a1881a <=( a52062a  and  a52049a );
 a1882a <=( a52038a  and  a52025a );
 a1883a <=( a52014a  and  a52001a );
 a1884a <=( a51990a  and  a51977a );
 a1885a <=( a51966a  and  a51953a );
 a1886a <=( a51942a  and  a51929a );
 a1887a <=( a51918a  and  a51905a );
 a1888a <=( a51894a  and  a51881a );
 a1889a <=( a51870a  and  a51857a );
 a1890a <=( a51846a  and  a51833a );
 a1891a <=( a51822a  and  a51809a );
 a1892a <=( a51798a  and  a51785a );
 a1893a <=( a51774a  and  a51761a );
 a1894a <=( a51750a  and  a51737a );
 a1895a <=( a51726a  and  a51713a );
 a1896a <=( a51702a  and  a51689a );
 a1897a <=( a51678a  and  a51665a );
 a1898a <=( a51654a  and  a51641a );
 a1899a <=( a51630a  and  a51617a );
 a1900a <=( a51606a  and  a51593a );
 a1901a <=( a51582a  and  a51569a );
 a1902a <=( a51558a  and  a51545a );
 a1903a <=( a51534a  and  a51521a );
 a1904a <=( a51510a  and  a51497a );
 a1905a <=( a51486a  and  a51473a );
 a1906a <=( a51462a  and  a51449a );
 a1907a <=( a51438a  and  a51425a );
 a1908a <=( a51414a  and  a51401a );
 a1909a <=( a51390a  and  a51377a );
 a1910a <=( a51366a  and  a51353a );
 a1911a <=( a51342a  and  a51329a );
 a1912a <=( a51318a  and  a51305a );
 a1913a <=( a51294a  and  a51281a );
 a1914a <=( a51270a  and  a51257a );
 a1915a <=( a51246a  and  a51233a );
 a1916a <=( a51222a  and  a51209a );
 a1917a <=( a51198a  and  a51185a );
 a1918a <=( a51174a  and  a51161a );
 a1919a <=( a51150a  and  a51137a );
 a1920a <=( a51126a  and  a51113a );
 a1921a <=( a51102a  and  a51089a );
 a1922a <=( a51078a  and  a51065a );
 a1923a <=( a51054a  and  a51041a );
 a1924a <=( a51030a  and  a51017a );
 a1925a <=( a51006a  and  a50993a );
 a1926a <=( a50982a  and  a50969a );
 a1927a <=( a50958a  and  a50945a );
 a1928a <=( a50934a  and  a50921a );
 a1929a <=( a50910a  and  a50897a );
 a1930a <=( a50886a  and  a50873a );
 a1931a <=( a50862a  and  a50849a );
 a1932a <=( a50838a  and  a50825a );
 a1933a <=( a50814a  and  a50801a );
 a1934a <=( a50790a  and  a50777a );
 a1935a <=( a50766a  and  a50753a );
 a1936a <=( a50742a  and  a50729a );
 a1937a <=( a50718a  and  a50705a );
 a1938a <=( a50694a  and  a50681a );
 a1939a <=( a50670a  and  a50657a );
 a1940a <=( a50646a  and  a50633a );
 a1941a <=( a50622a  and  a50609a );
 a1942a <=( a50598a  and  a50585a );
 a1943a <=( a50574a  and  a50561a );
 a1944a <=( a50550a  and  a50537a );
 a1945a <=( a50526a  and  a50513a );
 a1946a <=( a50502a  and  a50489a );
 a1947a <=( a50478a  and  a50465a );
 a1948a <=( a50454a  and  a50441a );
 a1949a <=( a50430a  and  a50417a );
 a1950a <=( a50406a  and  a50393a );
 a1951a <=( a50382a  and  a50369a );
 a1952a <=( a50358a  and  a50345a );
 a1953a <=( a50334a  and  a50321a );
 a1954a <=( a50310a  and  a50297a );
 a1955a <=( a50286a  and  a50273a );
 a1956a <=( a50262a  and  a50249a );
 a1957a <=( a50238a  and  a50225a );
 a1958a <=( a50214a  and  a50201a );
 a1959a <=( a50190a  and  a50177a );
 a1960a <=( a50166a  and  a50153a );
 a1961a <=( a50142a  and  a50129a );
 a1962a <=( a50118a  and  a50105a );
 a1963a <=( a50094a  and  a50081a );
 a1964a <=( a50070a  and  a50057a );
 a1965a <=( a50046a  and  a50033a );
 a1966a <=( a50022a  and  a50009a );
 a1967a <=( a49998a  and  a49985a );
 a1968a <=( a49974a  and  a49961a );
 a1969a <=( a49950a  and  a49937a );
 a1970a <=( a49926a  and  a49913a );
 a1971a <=( a49902a  and  a49889a );
 a1972a <=( a49878a  and  a49865a );
 a1973a <=( a49854a  and  a49841a );
 a1974a <=( a49830a  and  a49817a );
 a1975a <=( a49806a  and  a49793a );
 a1976a <=( a49782a  and  a49769a );
 a1977a <=( a49758a  and  a49745a );
 a1978a <=( a49734a  and  a49721a );
 a1979a <=( a49710a  and  a49697a );
 a1980a <=( a49686a  and  a49673a );
 a1981a <=( a49662a  and  a49649a );
 a1982a <=( a49638a  and  a49625a );
 a1983a <=( a49614a  and  a49601a );
 a1984a <=( a49590a  and  a49577a );
 a1985a <=( a49566a  and  a49553a );
 a1986a <=( a49542a  and  a49529a );
 a1987a <=( a49518a  and  a49505a );
 a1988a <=( a49494a  and  a49481a );
 a1989a <=( a49470a  and  a49457a );
 a1990a <=( a49446a  and  a49433a );
 a1991a <=( a49422a  and  a49409a );
 a1992a <=( a49398a  and  a49385a );
 a1993a <=( a49374a  and  a49361a );
 a1994a <=( a49350a  and  a49337a );
 a1995a <=( a49326a  and  a49313a );
 a1996a <=( a49302a  and  a49289a );
 a1997a <=( a49278a  and  a49265a );
 a1998a <=( a49254a  and  a49241a );
 a1999a <=( a49230a  and  a49217a );
 a2000a <=( a49206a  and  a49193a );
 a2001a <=( a49182a  and  a49169a );
 a2002a <=( a49158a  and  a49145a );
 a2003a <=( a49134a  and  a49121a );
 a2004a <=( a49110a  and  a49097a );
 a2005a <=( a49086a  and  a49073a );
 a2006a <=( a49062a  and  a49049a );
 a2007a <=( a49038a  and  a49025a );
 a2008a <=( a49014a  and  a49001a );
 a2009a <=( a48990a  and  a48977a );
 a2010a <=( a48966a  and  a48953a );
 a2011a <=( a48942a  and  a48929a );
 a2012a <=( a48918a  and  a48905a );
 a2013a <=( a48894a  and  a48881a );
 a2014a <=( a48870a  and  a48857a );
 a2015a <=( a48846a  and  a48833a );
 a2016a <=( a48822a  and  a48809a );
 a2017a <=( a48798a  and  a48785a );
 a2018a <=( a48774a  and  a48761a );
 a2019a <=( a48750a  and  a48737a );
 a2020a <=( a48726a  and  a48713a );
 a2021a <=( a48702a  and  a48689a );
 a2022a <=( a48678a  and  a48665a );
 a2023a <=( a48654a  and  a48641a );
 a2024a <=( a48630a  and  a48617a );
 a2025a <=( a48606a  and  a48593a );
 a2026a <=( a48582a  and  a48569a );
 a2027a <=( a48558a  and  a48545a );
 a2028a <=( a48534a  and  a48521a );
 a2029a <=( a48510a  and  a48497a );
 a2030a <=( a48486a  and  a48473a );
 a2031a <=( a48462a  and  a48449a );
 a2032a <=( a48438a  and  a48425a );
 a2033a <=( a48414a  and  a48401a );
 a2034a <=( a48390a  and  a48377a );
 a2035a <=( a48366a  and  a48353a );
 a2036a <=( a48342a  and  a48329a );
 a2037a <=( a48318a  and  a48305a );
 a2038a <=( a48294a  and  a48281a );
 a2039a <=( a48270a  and  a48257a );
 a2040a <=( a48246a  and  a48233a );
 a2041a <=( a48222a  and  a48209a );
 a2042a <=( a48198a  and  a48185a );
 a2043a <=( a48174a  and  a48161a );
 a2044a <=( a48150a  and  a48137a );
 a2045a <=( a48126a  and  a48113a );
 a2046a <=( a48102a  and  a48089a );
 a2047a <=( a48078a  and  a48065a );
 a2048a <=( a48054a  and  a48041a );
 a2049a <=( a48030a  and  a48017a );
 a2050a <=( a48006a  and  a47993a );
 a2051a <=( a47982a  and  a47969a );
 a2052a <=( a47958a  and  a47945a );
 a2053a <=( a47934a  and  a47921a );
 a2054a <=( a47910a  and  a47897a );
 a2055a <=( a47886a  and  a47873a );
 a2056a <=( a47862a  and  a47849a );
 a2057a <=( a47838a  and  a47825a );
 a2058a <=( a47814a  and  a47801a );
 a2059a <=( a47790a  and  a47777a );
 a2060a <=( a47766a  and  a47753a );
 a2061a <=( a47742a  and  a47729a );
 a2062a <=( a47718a  and  a47705a );
 a2063a <=( a47694a  and  a47681a );
 a2064a <=( a47670a  and  a47657a );
 a2065a <=( a47646a  and  a47633a );
 a2066a <=( a47622a  and  a47609a );
 a2067a <=( a47598a  and  a47585a );
 a2068a <=( a47574a  and  a47561a );
 a2069a <=( a47550a  and  a47537a );
 a2070a <=( a47526a  and  a47513a );
 a2071a <=( a47502a  and  a47489a );
 a2072a <=( a47478a  and  a47465a );
 a2073a <=( a47454a  and  a47441a );
 a2074a <=( a47430a  and  a47417a );
 a2075a <=( a47406a  and  a47393a );
 a2076a <=( a47382a  and  a47369a );
 a2077a <=( a47358a  and  a47345a );
 a2078a <=( a47334a  and  a47321a );
 a2079a <=( a47310a  and  a47297a );
 a2080a <=( a47286a  and  a47273a );
 a2081a <=( a47262a  and  a47249a );
 a2082a <=( a47238a  and  a47225a );
 a2083a <=( a47214a  and  a47201a );
 a2084a <=( a47190a  and  a47177a );
 a2085a <=( a47166a  and  a47153a );
 a2086a <=( a47142a  and  a47129a );
 a2087a <=( a47118a  and  a47105a );
 a2088a <=( a47094a  and  a47081a );
 a2089a <=( a47070a  and  a47057a );
 a2090a <=( a47046a  and  a47033a );
 a2091a <=( a47022a  and  a47009a );
 a2092a <=( a46998a  and  a46985a );
 a2093a <=( a46974a  and  a46961a );
 a2094a <=( a46950a  and  a46937a );
 a2095a <=( a46926a  and  a46913a );
 a2096a <=( a46902a  and  a46889a );
 a2097a <=( a46878a  and  a46865a );
 a2098a <=( a46854a  and  a46841a );
 a2099a <=( a46830a  and  a46817a );
 a2100a <=( a46806a  and  a46793a );
 a2101a <=( a46782a  and  a46769a );
 a2102a <=( a46758a  and  a46745a );
 a2103a <=( a46734a  and  a46721a );
 a2104a <=( a46710a  and  a46697a );
 a2105a <=( a46686a  and  a46673a );
 a2106a <=( a46662a  and  a46649a );
 a2107a <=( a46638a  and  a46625a );
 a2108a <=( a46614a  and  a46601a );
 a2109a <=( a46590a  and  a46577a );
 a2110a <=( a46566a  and  a46553a );
 a2111a <=( a46542a  and  a46529a );
 a2112a <=( a46518a  and  a46505a );
 a2113a <=( a46494a  and  a46481a );
 a2114a <=( a46470a  and  a46457a );
 a2115a <=( a46446a  and  a46433a );
 a2116a <=( a46422a  and  a46409a );
 a2117a <=( a46398a  and  a46385a );
 a2118a <=( a46374a  and  a46361a );
 a2119a <=( a46350a  and  a46337a );
 a2120a <=( a46326a  and  a46313a );
 a2121a <=( a46302a  and  a46289a );
 a2122a <=( a46278a  and  a46265a );
 a2123a <=( a46254a  and  a46241a );
 a2124a <=( a46230a  and  a46217a );
 a2125a <=( a46206a  and  a46193a );
 a2126a <=( a46182a  and  a46169a );
 a2127a <=( a46158a  and  a46145a );
 a2128a <=( a46134a  and  a46121a );
 a2129a <=( a46110a  and  a46097a );
 a2130a <=( a46086a  and  a46073a );
 a2131a <=( a46062a  and  a46049a );
 a2132a <=( a46038a  and  a46025a );
 a2133a <=( a46014a  and  a46001a );
 a2134a <=( a45990a  and  a45977a );
 a2135a <=( a45966a  and  a45953a );
 a2136a <=( a45942a  and  a45929a );
 a2137a <=( a45918a  and  a45905a );
 a2138a <=( a45894a  and  a45881a );
 a2139a <=( a45870a  and  a45857a );
 a2140a <=( a45846a  and  a45833a );
 a2141a <=( a45822a  and  a45809a );
 a2142a <=( a45798a  and  a45785a );
 a2143a <=( a45774a  and  a45761a );
 a2144a <=( a45750a  and  a45737a );
 a2145a <=( a45726a  and  a45713a );
 a2146a <=( a45702a  and  a45689a );
 a2147a <=( a45678a  and  a45665a );
 a2148a <=( a45654a  and  a45641a );
 a2149a <=( a45630a  and  a45617a );
 a2150a <=( a45606a  and  a45593a );
 a2151a <=( a45582a  and  a45569a );
 a2152a <=( a45558a  and  a45545a );
 a2153a <=( a45534a  and  a45521a );
 a2154a <=( a45510a  and  a45497a );
 a2155a <=( a45486a  and  a45473a );
 a2156a <=( a45462a  and  a45449a );
 a2157a <=( a45438a  and  a45425a );
 a2158a <=( a45414a  and  a45401a );
 a2159a <=( a45390a  and  a45377a );
 a2160a <=( a45366a  and  a45353a );
 a2161a <=( a45342a  and  a45329a );
 a2162a <=( a45318a  and  a45305a );
 a2163a <=( a45294a  and  a45281a );
 a2164a <=( a45270a  and  a45257a );
 a2165a <=( a45246a  and  a45233a );
 a2166a <=( a45222a  and  a45209a );
 a2167a <=( a45198a  and  a45185a );
 a2168a <=( a45174a  and  a45161a );
 a2169a <=( a45150a  and  a45137a );
 a2170a <=( a45126a  and  a45113a );
 a2171a <=( a45102a  and  a45089a );
 a2172a <=( a45078a  and  a45065a );
 a2173a <=( a45054a  and  a45041a );
 a2174a <=( a45030a  and  a45017a );
 a2175a <=( a45006a  and  a44993a );
 a2176a <=( a44982a  and  a44969a );
 a2177a <=( a44958a  and  a44945a );
 a2178a <=( a44934a  and  a44921a );
 a2179a <=( a44910a  and  a44897a );
 a2180a <=( a44886a  and  a44873a );
 a2181a <=( a44862a  and  a44849a );
 a2182a <=( a44838a  and  a44825a );
 a2183a <=( a44814a  and  a44801a );
 a2184a <=( a44790a  and  a44777a );
 a2185a <=( a44766a  and  a44753a );
 a2186a <=( a44742a  and  a44729a );
 a2187a <=( a44718a  and  a44705a );
 a2188a <=( a44694a  and  a44681a );
 a2189a <=( a44670a  and  a44657a );
 a2190a <=( a44646a  and  a44633a );
 a2191a <=( a44622a  and  a44609a );
 a2192a <=( a44598a  and  a44585a );
 a2193a <=( a44574a  and  a44561a );
 a2194a <=( a44550a  and  a44537a );
 a2195a <=( a44526a  and  a44513a );
 a2196a <=( a44502a  and  a44489a );
 a2197a <=( a44478a  and  a44465a );
 a2198a <=( a44454a  and  a44441a );
 a2199a <=( a44430a  and  a44417a );
 a2200a <=( a44406a  and  a44393a );
 a2201a <=( a44382a  and  a44369a );
 a2202a <=( a44358a  and  a44345a );
 a2203a <=( a44334a  and  a44321a );
 a2204a <=( a44310a  and  a44297a );
 a2205a <=( a44286a  and  a44273a );
 a2206a <=( a44262a  and  a44249a );
 a2207a <=( a44238a  and  a44225a );
 a2208a <=( a44214a  and  a44201a );
 a2209a <=( a44190a  and  a44177a );
 a2210a <=( a44166a  and  a44153a );
 a2211a <=( a44142a  and  a44129a );
 a2212a <=( a44118a  and  a44105a );
 a2213a <=( a44094a  and  a44081a );
 a2214a <=( a44070a  and  a44057a );
 a2215a <=( a44046a  and  a44033a );
 a2216a <=( a44022a  and  a44009a );
 a2217a <=( a43998a  and  a43985a );
 a2218a <=( a43974a  and  a43961a );
 a2219a <=( a43950a  and  a43937a );
 a2220a <=( a43926a  and  a43913a );
 a2221a <=( a43902a  and  a43889a );
 a2222a <=( a43878a  and  a43865a );
 a2223a <=( a43854a  and  a43841a );
 a2224a <=( a43830a  and  a43817a );
 a2225a <=( a43806a  and  a43793a );
 a2226a <=( a43782a  and  a43769a );
 a2227a <=( a43758a  and  a43745a );
 a2228a <=( a43734a  and  a43721a );
 a2229a <=( a43710a  and  a43697a );
 a2230a <=( a43686a  and  a43673a );
 a2231a <=( a43662a  and  a43649a );
 a2232a <=( a43638a  and  a43625a );
 a2233a <=( a43614a  and  a43601a );
 a2234a <=( a43590a  and  a43577a );
 a2235a <=( a43566a  and  a43553a );
 a2236a <=( a43542a  and  a43529a );
 a2237a <=( a43518a  and  a43505a );
 a2238a <=( a43494a  and  a43481a );
 a2239a <=( a43470a  and  a43457a );
 a2240a <=( a43446a  and  a43433a );
 a2241a <=( a43422a  and  a43409a );
 a2242a <=( a43398a  and  a43385a );
 a2243a <=( a43374a  and  a43361a );
 a2244a <=( a43350a  and  a43337a );
 a2245a <=( a43326a  and  a43313a );
 a2246a <=( a43302a  and  a43289a );
 a2247a <=( a43278a  and  a43265a );
 a2248a <=( a43254a  and  a43241a );
 a2249a <=( a43230a  and  a43217a );
 a2250a <=( a43206a  and  a43193a );
 a2251a <=( a43182a  and  a43169a );
 a2252a <=( a43158a  and  a43145a );
 a2253a <=( a43134a  and  a43121a );
 a2254a <=( a43110a  and  a43097a );
 a2255a <=( a43086a  and  a43073a );
 a2256a <=( a43062a  and  a43049a );
 a2257a <=( a43038a  and  a43025a );
 a2258a <=( a43014a  and  a43001a );
 a2259a <=( a42990a  and  a42977a );
 a2260a <=( a42966a  and  a42953a );
 a2261a <=( a42942a  and  a42929a );
 a2262a <=( a42918a  and  a42905a );
 a2263a <=( a42894a  and  a42881a );
 a2264a <=( a42870a  and  a42857a );
 a2265a <=( a42846a  and  a42833a );
 a2266a <=( a42822a  and  a42809a );
 a2267a <=( a42798a  and  a42785a );
 a2268a <=( a42774a  and  a42761a );
 a2269a <=( a42750a  and  a42737a );
 a2270a <=( a42726a  and  a42713a );
 a2271a <=( a42702a  and  a42689a );
 a2272a <=( a42678a  and  a42665a );
 a2273a <=( a42654a  and  a42641a );
 a2274a <=( a42630a  and  a42617a );
 a2275a <=( a42606a  and  a42593a );
 a2276a <=( a42582a  and  a42569a );
 a2277a <=( a42558a  and  a42545a );
 a2278a <=( a42534a  and  a42521a );
 a2279a <=( a42510a  and  a42497a );
 a2280a <=( a42486a  and  a42473a );
 a2281a <=( a42462a  and  a42449a );
 a2282a <=( a42438a  and  a42425a );
 a2283a <=( a42414a  and  a42401a );
 a2284a <=( a42390a  and  a42377a );
 a2285a <=( a42366a  and  a42353a );
 a2286a <=( a42342a  and  a42329a );
 a2287a <=( a42318a  and  a42305a );
 a2288a <=( a42294a  and  a42281a );
 a2289a <=( a42270a  and  a42257a );
 a2290a <=( a42246a  and  a42233a );
 a2291a <=( a42222a  and  a42209a );
 a2292a <=( a42198a  and  a42185a );
 a2293a <=( a42174a  and  a42161a );
 a2294a <=( a42150a  and  a42137a );
 a2295a <=( a42126a  and  a42113a );
 a2296a <=( a42102a  and  a42089a );
 a2297a <=( a42078a  and  a42065a );
 a2298a <=( a42054a  and  a42041a );
 a2299a <=( a42030a  and  a42017a );
 a2300a <=( a42006a  and  a41993a );
 a2301a <=( a41982a  and  a41969a );
 a2302a <=( a41958a  and  a41945a );
 a2303a <=( a41934a  and  a41921a );
 a2304a <=( a41910a  and  a41897a );
 a2305a <=( a41886a  and  a41873a );
 a2306a <=( a41862a  and  a41849a );
 a2307a <=( a41838a  and  a41825a );
 a2308a <=( a41814a  and  a41801a );
 a2309a <=( a41790a  and  a41777a );
 a2310a <=( a41766a  and  a41753a );
 a2311a <=( a41742a  and  a41729a );
 a2312a <=( a41718a  and  a41705a );
 a2313a <=( a41694a  and  a41681a );
 a2314a <=( a41670a  and  a41657a );
 a2315a <=( a41646a  and  a41633a );
 a2316a <=( a41622a  and  a41609a );
 a2317a <=( a41598a  and  a41585a );
 a2318a <=( a41574a  and  a41561a );
 a2319a <=( a41550a  and  a41537a );
 a2320a <=( a41526a  and  a41513a );
 a2321a <=( a41502a  and  a41489a );
 a2322a <=( a41478a  and  a41465a );
 a2323a <=( a41454a  and  a41441a );
 a2324a <=( a41430a  and  a41417a );
 a2325a <=( a41406a  and  a41393a );
 a2326a <=( a41382a  and  a41369a );
 a2327a <=( a41358a  and  a41345a );
 a2328a <=( a41334a  and  a41321a );
 a2329a <=( a41310a  and  a41299a );
 a2330a <=( a41288a  and  a41277a );
 a2331a <=( a41266a  and  a41255a );
 a2332a <=( a41244a  and  a41233a );
 a2333a <=( a41222a  and  a41211a );
 a2334a <=( a41200a  and  a41189a );
 a2335a <=( a41178a  and  a41167a );
 a2336a <=( a41156a  and  a41145a );
 a2337a <=( a41134a  and  a41123a );
 a2338a <=( a41112a  and  a41101a );
 a2339a <=( a41090a  and  a41079a );
 a2340a <=( a41068a  and  a41057a );
 a2341a <=( a41046a  and  a41035a );
 a2342a <=( a41024a  and  a41013a );
 a2343a <=( a41002a  and  a40991a );
 a2344a <=( a40980a  and  a40969a );
 a2345a <=( a40958a  and  a40947a );
 a2346a <=( a40936a  and  a40925a );
 a2347a <=( a40914a  and  a40903a );
 a2348a <=( a40892a  and  a40881a );
 a2349a <=( a40870a  and  a40859a );
 a2350a <=( a40848a  and  a40837a );
 a2351a <=( a40826a  and  a40815a );
 a2352a <=( a40804a  and  a40793a );
 a2353a <=( a40782a  and  a40771a );
 a2354a <=( a40760a  and  a40749a );
 a2355a <=( a40738a  and  a40727a );
 a2356a <=( a40716a  and  a40705a );
 a2357a <=( a40694a  and  a40683a );
 a2358a <=( a40672a  and  a40661a );
 a2359a <=( a40650a  and  a40639a );
 a2360a <=( a40628a  and  a40617a );
 a2361a <=( a40606a  and  a40595a );
 a2362a <=( a40584a  and  a40573a );
 a2363a <=( a40562a  and  a40551a );
 a2364a <=( a40540a  and  a40529a );
 a2365a <=( a40518a  and  a40507a );
 a2366a <=( a40496a  and  a40485a );
 a2367a <=( a40474a  and  a40463a );
 a2368a <=( a40452a  and  a40441a );
 a2369a <=( a40430a  and  a40419a );
 a2370a <=( a40408a  and  a40397a );
 a2371a <=( a40386a  and  a40375a );
 a2372a <=( a40364a  and  a40353a );
 a2373a <=( a40342a  and  a40331a );
 a2374a <=( a40320a  and  a40309a );
 a2375a <=( a40298a  and  a40287a );
 a2376a <=( a40276a  and  a40265a );
 a2377a <=( a40254a  and  a40243a );
 a2378a <=( a40232a  and  a40221a );
 a2379a <=( a40210a  and  a40199a );
 a2380a <=( a40188a  and  a40177a );
 a2381a <=( a40166a  and  a40155a );
 a2382a <=( a40144a  and  a40133a );
 a2383a <=( a40122a  and  a40111a );
 a2384a <=( a40100a  and  a40089a );
 a2385a <=( a40078a  and  a40067a );
 a2386a <=( a40056a  and  a40045a );
 a2387a <=( a40034a  and  a40023a );
 a2388a <=( a40012a  and  a40001a );
 a2389a <=( a39990a  and  a39979a );
 a2390a <=( a39968a  and  a39957a );
 a2391a <=( a39946a  and  a39935a );
 a2392a <=( a39924a  and  a39913a );
 a2393a <=( a39902a  and  a39891a );
 a2394a <=( a39880a  and  a39869a );
 a2395a <=( a39858a  and  a39847a );
 a2396a <=( a39836a  and  a39825a );
 a2397a <=( a39814a  and  a39803a );
 a2398a <=( a39792a  and  a39781a );
 a2399a <=( a39770a  and  a39759a );
 a2400a <=( a39748a  and  a39737a );
 a2401a <=( a39726a  and  a39715a );
 a2402a <=( a39704a  and  a39693a );
 a2403a <=( a39682a  and  a39671a );
 a2404a <=( a39660a  and  a39649a );
 a2405a <=( a39638a  and  a39627a );
 a2406a <=( a39616a  and  a39605a );
 a2407a <=( a39594a  and  a39583a );
 a2408a <=( a39572a  and  a39561a );
 a2409a <=( a39550a  and  a39539a );
 a2410a <=( a39528a  and  a39517a );
 a2411a <=( a39506a  and  a39495a );
 a2412a <=( a39484a  and  a39473a );
 a2413a <=( a39462a  and  a39451a );
 a2414a <=( a39440a  and  a39429a );
 a2415a <=( a39418a  and  a39407a );
 a2416a <=( a39396a  and  a39385a );
 a2417a <=( a39374a  and  a39363a );
 a2418a <=( a39352a  and  a39341a );
 a2419a <=( a39330a  and  a39319a );
 a2420a <=( a39308a  and  a39297a );
 a2421a <=( a39286a  and  a39275a );
 a2422a <=( a39264a  and  a39253a );
 a2423a <=( a39242a  and  a39231a );
 a2424a <=( a39220a  and  a39209a );
 a2425a <=( a39198a  and  a39187a );
 a2426a <=( a39176a  and  a39165a );
 a2427a <=( a39154a  and  a39143a );
 a2428a <=( a39132a  and  a39121a );
 a2429a <=( a39110a  and  a39099a );
 a2430a <=( a39088a  and  a39077a );
 a2431a <=( a39066a  and  a39055a );
 a2432a <=( a39044a  and  a39033a );
 a2433a <=( a39022a  and  a39011a );
 a2434a <=( a39000a  and  a38989a );
 a2435a <=( a38978a  and  a38967a );
 a2436a <=( a38956a  and  a38945a );
 a2437a <=( a38934a  and  a38923a );
 a2438a <=( a38912a  and  a38901a );
 a2439a <=( a38890a  and  a38879a );
 a2440a <=( a38868a  and  a38857a );
 a2441a <=( a38846a  and  a38835a );
 a2442a <=( a38824a  and  a38813a );
 a2443a <=( a38802a  and  a38791a );
 a2444a <=( a38780a  and  a38769a );
 a2445a <=( a38758a  and  a38747a );
 a2446a <=( a38736a  and  a38725a );
 a2447a <=( a38714a  and  a38703a );
 a2448a <=( a38692a  and  a38681a );
 a2449a <=( a38670a  and  a38659a );
 a2450a <=( a38648a  and  a38637a );
 a2451a <=( a38626a  and  a38615a );
 a2452a <=( a38604a  and  a38593a );
 a2453a <=( a38582a  and  a38571a );
 a2454a <=( a38560a  and  a38549a );
 a2455a <=( a38538a  and  a38527a );
 a2456a <=( a38516a  and  a38505a );
 a2457a <=( a38494a  and  a38483a );
 a2458a <=( a38472a  and  a38461a );
 a2459a <=( a38450a  and  a38439a );
 a2460a <=( a38428a  and  a38417a );
 a2461a <=( a38406a  and  a38395a );
 a2462a <=( a38384a  and  a38373a );
 a2463a <=( a38362a  and  a38351a );
 a2464a <=( a38340a  and  a38329a );
 a2465a <=( a38318a  and  a38307a );
 a2466a <=( a38296a  and  a38285a );
 a2467a <=( a38274a  and  a38263a );
 a2468a <=( a38252a  and  a38241a );
 a2469a <=( a38230a  and  a38219a );
 a2470a <=( a38208a  and  a38197a );
 a2471a <=( a38186a  and  a38175a );
 a2472a <=( a38164a  and  a38153a );
 a2473a <=( a38142a  and  a38131a );
 a2474a <=( a38120a  and  a38109a );
 a2475a <=( a38098a  and  a38087a );
 a2476a <=( a38076a  and  a38065a );
 a2477a <=( a38054a  and  a38043a );
 a2478a <=( a38032a  and  a38021a );
 a2479a <=( a38010a  and  a37999a );
 a2480a <=( a37988a  and  a37977a );
 a2481a <=( a37966a  and  a37955a );
 a2482a <=( a37944a  and  a37933a );
 a2483a <=( a37922a  and  a37911a );
 a2484a <=( a37900a  and  a37889a );
 a2485a <=( a37878a  and  a37867a );
 a2486a <=( a37856a  and  a37845a );
 a2487a <=( a37834a  and  a37823a );
 a2488a <=( a37812a  and  a37801a );
 a2489a <=( a37790a  and  a37779a );
 a2490a <=( a37768a  and  a37757a );
 a2491a <=( a37746a  and  a37735a );
 a2492a <=( a37724a  and  a37713a );
 a2493a <=( a37702a  and  a37691a );
 a2494a <=( a37680a  and  a37669a );
 a2495a <=( a37658a  and  a37647a );
 a2496a <=( a37636a  and  a37625a );
 a2497a <=( a37614a  and  a37603a );
 a2498a <=( a37592a  and  a37581a );
 a2499a <=( a37570a  and  a37559a );
 a2500a <=( a37548a  and  a37537a );
 a2501a <=( a37526a  and  a37515a );
 a2502a <=( a37504a  and  a37493a );
 a2503a <=( a37482a  and  a37471a );
 a2504a <=( a37460a  and  a37449a );
 a2505a <=( a37438a  and  a37427a );
 a2506a <=( a37416a  and  a37405a );
 a2507a <=( a37394a  and  a37383a );
 a2508a <=( a37372a  and  a37361a );
 a2509a <=( a37350a  and  a37339a );
 a2510a <=( a37328a  and  a37317a );
 a2511a <=( a37306a  and  a37295a );
 a2512a <=( a37284a  and  a37273a );
 a2513a <=( a37262a  and  a37251a );
 a2514a <=( a37240a  and  a37229a );
 a2515a <=( a37218a  and  a37207a );
 a2516a <=( a37196a  and  a37185a );
 a2517a <=( a37174a  and  a37163a );
 a2518a <=( a37152a  and  a37141a );
 a2519a <=( a37130a  and  a37119a );
 a2520a <=( a37108a  and  a37097a );
 a2521a <=( a37086a  and  a37075a );
 a2522a <=( a37064a  and  a37053a );
 a2523a <=( a37042a  and  a37031a );
 a2524a <=( a37020a  and  a37009a );
 a2525a <=( a36998a  and  a36987a );
 a2526a <=( a36976a  and  a36965a );
 a2527a <=( a36954a  and  a36943a );
 a2528a <=( a36932a  and  a36921a );
 a2529a <=( a36910a  and  a36899a );
 a2530a <=( a36888a  and  a36877a );
 a2531a <=( a36866a  and  a36855a );
 a2532a <=( a36844a  and  a36833a );
 a2533a <=( a36822a  and  a36811a );
 a2534a <=( a36800a  and  a36789a );
 a2535a <=( a36778a  and  a36767a );
 a2536a <=( a36756a  and  a36745a );
 a2537a <=( a36734a  and  a36723a );
 a2538a <=( a36712a  and  a36701a );
 a2539a <=( a36690a  and  a36679a );
 a2540a <=( a36668a  and  a36657a );
 a2541a <=( a36646a  and  a36635a );
 a2542a <=( a36624a  and  a36613a );
 a2543a <=( a36602a  and  a36591a );
 a2544a <=( a36580a  and  a36569a );
 a2545a <=( a36558a  and  a36547a );
 a2546a <=( a36536a  and  a36525a );
 a2547a <=( a36514a  and  a36503a );
 a2548a <=( a36492a  and  a36481a );
 a2549a <=( a36470a  and  a36459a );
 a2550a <=( a36448a  and  a36437a );
 a2551a <=( a36426a  and  a36415a );
 a2552a <=( a36404a  and  a36393a );
 a2553a <=( a36382a  and  a36371a );
 a2554a <=( a36360a  and  a36349a );
 a2555a <=( a36338a  and  a36327a );
 a2556a <=( a36316a  and  a36305a );
 a2557a <=( a36294a  and  a36283a );
 a2558a <=( a36272a  and  a36261a );
 a2559a <=( a36250a  and  a36239a );
 a2560a <=( a36228a  and  a36217a );
 a2561a <=( a36206a  and  a36195a );
 a2562a <=( a36184a  and  a36173a );
 a2563a <=( a36162a  and  a36151a );
 a2564a <=( a36140a  and  a36129a );
 a2565a <=( a36118a  and  a36107a );
 a2566a <=( a36096a  and  a36085a );
 a2567a <=( a36074a  and  a36063a );
 a2568a <=( a36052a  and  a36041a );
 a2569a <=( a36030a  and  a36019a );
 a2570a <=( a36008a  and  a35997a );
 a2571a <=( a35986a  and  a35975a );
 a2572a <=( a35964a  and  a35953a );
 a2573a <=( a35942a  and  a35931a );
 a2574a <=( a35920a  and  a35909a );
 a2575a <=( a35898a  and  a35887a );
 a2576a <=( a35876a  and  a35865a );
 a2577a <=( a35854a  and  a35843a );
 a2578a <=( a35832a  and  a35821a );
 a2579a <=( a35810a  and  a35799a );
 a2580a <=( a35788a  and  a35777a );
 a2581a <=( a35766a  and  a35755a );
 a2582a <=( a35744a  and  a35733a );
 a2583a <=( a35722a  and  a35711a );
 a2584a <=( a35700a  and  a35689a );
 a2585a <=( a35678a  and  a35667a );
 a2586a <=( a35656a  and  a35645a );
 a2587a <=( a35634a  and  a35623a );
 a2588a <=( a35612a  and  a35601a );
 a2589a <=( a35590a  and  a35579a );
 a2590a <=( a35568a  and  a35557a );
 a2591a <=( a35546a  and  a35535a );
 a2592a <=( a35524a  and  a35513a );
 a2593a <=( a35502a  and  a35491a );
 a2594a <=( a35480a  and  a35469a );
 a2595a <=( a35458a  and  a35447a );
 a2596a <=( a35436a  and  a35425a );
 a2597a <=( a35414a  and  a35403a );
 a2598a <=( a35392a  and  a35381a );
 a2599a <=( a35370a  and  a35359a );
 a2600a <=( a35348a  and  a35337a );
 a2601a <=( a35326a  and  a35315a );
 a2602a <=( a35304a  and  a35293a );
 a2603a <=( a35282a  and  a35271a );
 a2604a <=( a35260a  and  a35249a );
 a2605a <=( a35238a  and  a35227a );
 a2606a <=( a35216a  and  a35205a );
 a2607a <=( a35194a  and  a35183a );
 a2608a <=( a35172a  and  a35161a );
 a2609a <=( a35150a  and  a35139a );
 a2610a <=( a35128a  and  a35117a );
 a2611a <=( a35106a  and  a35095a );
 a2612a <=( a35084a  and  a35073a );
 a2613a <=( a35062a  and  a35051a );
 a2614a <=( a35040a  and  a35029a );
 a2615a <=( a35018a  and  a35007a );
 a2616a <=( a34996a  and  a34985a );
 a2617a <=( a34974a  and  a34963a );
 a2618a <=( a34952a  and  a34941a );
 a2619a <=( a34930a  and  a34919a );
 a2620a <=( a34908a  and  a34897a );
 a2621a <=( a34886a  and  a34875a );
 a2622a <=( a34864a  and  a34853a );
 a2623a <=( a34842a  and  a34831a );
 a2624a <=( a34820a  and  a34809a );
 a2625a <=( a34798a  and  a34787a );
 a2626a <=( a34776a  and  a34765a );
 a2627a <=( a34754a  and  a34743a );
 a2628a <=( a34732a  and  a34721a );
 a2629a <=( a34710a  and  a34699a );
 a2630a <=( a34688a  and  a34677a );
 a2631a <=( a34666a  and  a34655a );
 a2632a <=( a34644a  and  a34633a );
 a2633a <=( a34622a  and  a34611a );
 a2634a <=( a34600a  and  a34589a );
 a2635a <=( a34578a  and  a34567a );
 a2636a <=( a34556a  and  a34545a );
 a2637a <=( a34534a  and  a34523a );
 a2638a <=( a34512a  and  a34501a );
 a2639a <=( a34490a  and  a34479a );
 a2640a <=( a34468a  and  a34457a );
 a2641a <=( a34446a  and  a34435a );
 a2642a <=( a34424a  and  a34413a );
 a2643a <=( a34402a  and  a34391a );
 a2644a <=( a34380a  and  a34369a );
 a2645a <=( a34358a  and  a34347a );
 a2646a <=( a34336a  and  a34325a );
 a2647a <=( a34314a  and  a34303a );
 a2648a <=( a34292a  and  a34281a );
 a2649a <=( a34270a  and  a34259a );
 a2650a <=( a34248a  and  a34237a );
 a2651a <=( a34226a  and  a34215a );
 a2652a <=( a34204a  and  a34193a );
 a2653a <=( a34182a  and  a34171a );
 a2654a <=( a34160a  and  a34149a );
 a2655a <=( a34138a  and  a34127a );
 a2656a <=( a34116a  and  a34105a );
 a2657a <=( a34094a  and  a34083a );
 a2658a <=( a34072a  and  a34061a );
 a2659a <=( a34050a  and  a34039a );
 a2660a <=( a34028a  and  a34017a );
 a2661a <=( a34006a  and  a33995a );
 a2662a <=( a33984a  and  a33973a );
 a2663a <=( a33962a  and  a33951a );
 a2664a <=( a33940a  and  a33929a );
 a2665a <=( a33918a  and  a33907a );
 a2666a <=( a33896a  and  a33885a );
 a2667a <=( a33874a  and  a33863a );
 a2668a <=( a33852a  and  a33841a );
 a2669a <=( a33830a  and  a33819a );
 a2670a <=( a33808a  and  a33797a );
 a2671a <=( a33786a  and  a33775a );
 a2672a <=( a33764a  and  a33753a );
 a2673a <=( a33742a  and  a33731a );
 a2674a <=( a33720a  and  a33709a );
 a2675a <=( a33698a  and  a33687a );
 a2676a <=( a33676a  and  a33665a );
 a2677a <=( a33654a  and  a33643a );
 a2678a <=( a33632a  and  a33621a );
 a2679a <=( a33610a  and  a33599a );
 a2680a <=( a33588a  and  a33577a );
 a2681a <=( a33566a  and  a33555a );
 a2682a <=( a33544a  and  a33533a );
 a2683a <=( a33522a  and  a33511a );
 a2684a <=( a33500a  and  a33489a );
 a2685a <=( a33478a  and  a33467a );
 a2686a <=( a33456a  and  a33445a );
 a2687a <=( a33434a  and  a33423a );
 a2688a <=( a33412a  and  a33401a );
 a2689a <=( a33390a  and  a33379a );
 a2690a <=( a33368a  and  a33357a );
 a2691a <=( a33346a  and  a33335a );
 a2692a <=( a33324a  and  a33313a );
 a2693a <=( a33302a  and  a33291a );
 a2694a <=( a33280a  and  a33269a );
 a2695a <=( a33258a  and  a33247a );
 a2696a <=( a33236a  and  a33225a );
 a2697a <=( a33214a  and  a33203a );
 a2698a <=( a33192a  and  a33181a );
 a2699a <=( a33170a  and  a33159a );
 a2700a <=( a33148a  and  a33137a );
 a2701a <=( a33126a  and  a33115a );
 a2702a <=( a33104a  and  a33093a );
 a2703a <=( a33082a  and  a33071a );
 a2704a <=( a33060a  and  a33049a );
 a2705a <=( a33038a  and  a33027a );
 a2706a <=( a33016a  and  a33005a );
 a2707a <=( a32994a  and  a32983a );
 a2708a <=( a32972a  and  a32961a );
 a2709a <=( a32950a  and  a32939a );
 a2710a <=( a32928a  and  a32917a );
 a2711a <=( a32906a  and  a32895a );
 a2712a <=( a32884a  and  a32873a );
 a2713a <=( a32862a  and  a32851a );
 a2714a <=( a32840a  and  a32829a );
 a2715a <=( a32818a  and  a32807a );
 a2716a <=( a32796a  and  a32785a );
 a2717a <=( a32774a  and  a32763a );
 a2718a <=( a32752a  and  a32741a );
 a2719a <=( a32730a  and  a32719a );
 a2720a <=( a32708a  and  a32697a );
 a2721a <=( a32686a  and  a32675a );
 a2722a <=( a32664a  and  a32653a );
 a2723a <=( a32642a  and  a32631a );
 a2724a <=( a32620a  and  a32609a );
 a2725a <=( a32598a  and  a32587a );
 a2726a <=( a32576a  and  a32565a );
 a2727a <=( a32554a  and  a32543a );
 a2728a <=( a32532a  and  a32521a );
 a2729a <=( a32510a  and  a32499a );
 a2730a <=( a32488a  and  a32477a );
 a2731a <=( a32466a  and  a32455a );
 a2732a <=( a32444a  and  a32433a );
 a2733a <=( a32422a  and  a32411a );
 a2734a <=( a32400a  and  a32389a );
 a2735a <=( a32378a  and  a32367a );
 a2736a <=( a32356a  and  a32345a );
 a2737a <=( a32334a  and  a32323a );
 a2738a <=( a32312a  and  a32301a );
 a2739a <=( a32290a  and  a32279a );
 a2740a <=( a32268a  and  a32257a );
 a2741a <=( a32246a  and  a32235a );
 a2742a <=( a32224a  and  a32213a );
 a2743a <=( a32202a  and  a32191a );
 a2744a <=( a32180a  and  a32169a );
 a2745a <=( a32158a  and  a32147a );
 a2746a <=( a32136a  and  a32125a );
 a2747a <=( a32114a  and  a32103a );
 a2748a <=( a32092a  and  a32081a );
 a2749a <=( a32070a  and  a32059a );
 a2750a <=( a32048a  and  a32037a );
 a2751a <=( a32026a  and  a32015a );
 a2752a <=( a32004a  and  a31993a );
 a2753a <=( a31982a  and  a31971a );
 a2754a <=( a31960a  and  a31949a );
 a2755a <=( a31938a  and  a31927a );
 a2756a <=( a31916a  and  a31905a );
 a2757a <=( a31894a  and  a31883a );
 a2758a <=( a31872a  and  a31861a );
 a2759a <=( a31850a  and  a31839a );
 a2760a <=( a31828a  and  a31817a );
 a2761a <=( a31806a  and  a31795a );
 a2762a <=( a31784a  and  a31773a );
 a2763a <=( a31762a  and  a31751a );
 a2764a <=( a31740a  and  a31729a );
 a2765a <=( a31718a  and  a31707a );
 a2766a <=( a31696a  and  a31685a );
 a2767a <=( a31674a  and  a31663a );
 a2768a <=( a31652a  and  a31641a );
 a2769a <=( a31630a  and  a31619a );
 a2770a <=( a31608a  and  a31597a );
 a2771a <=( a31586a  and  a31575a );
 a2772a <=( a31564a  and  a31553a );
 a2773a <=( a31542a  and  a31531a );
 a2774a <=( a31520a  and  a31509a );
 a2775a <=( a31498a  and  a31487a );
 a2776a <=( a31476a  and  a31465a );
 a2777a <=( a31454a  and  a31443a );
 a2778a <=( a31432a  and  a31421a );
 a2779a <=( a31410a  and  a31399a );
 a2780a <=( a31388a  and  a31377a );
 a2781a <=( a31366a  and  a31355a );
 a2782a <=( a31344a  and  a31333a );
 a2783a <=( a31322a  and  a31311a );
 a2784a <=( a31300a  and  a31289a );
 a2785a <=( a31278a  and  a31267a );
 a2786a <=( a31256a  and  a31245a );
 a2787a <=( a31234a  and  a31223a );
 a2788a <=( a31212a  and  a31201a );
 a2789a <=( a31190a  and  a31179a );
 a2790a <=( a31168a  and  a31157a );
 a2791a <=( a31146a  and  a31135a );
 a2792a <=( a31124a  and  a31113a );
 a2793a <=( a31102a  and  a31091a );
 a2794a <=( a31080a  and  a31069a );
 a2795a <=( a31058a  and  a31047a );
 a2796a <=( a31036a  and  a31025a );
 a2797a <=( a31014a  and  a31003a );
 a2798a <=( a30992a  and  a30981a );
 a2799a <=( a30970a  and  a30959a );
 a2800a <=( a30948a  and  a30937a );
 a2801a <=( a30926a  and  a30915a );
 a2802a <=( a30904a  and  a30893a );
 a2803a <=( a30882a  and  a30871a );
 a2804a <=( a30860a  and  a30849a );
 a2805a <=( a30838a  and  a30827a );
 a2806a <=( a30816a  and  a30805a );
 a2807a <=( a30794a  and  a30783a );
 a2808a <=( a30772a  and  a30761a );
 a2809a <=( a30750a  and  a30739a );
 a2810a <=( a30728a  and  a30717a );
 a2811a <=( a30706a  and  a30695a );
 a2812a <=( a30684a  and  a30673a );
 a2813a <=( a30662a  and  a30651a );
 a2814a <=( a30640a  and  a30629a );
 a2815a <=( a30618a  and  a30607a );
 a2816a <=( a30596a  and  a30585a );
 a2817a <=( a30574a  and  a30563a );
 a2818a <=( a30552a  and  a30541a );
 a2819a <=( a30530a  and  a30519a );
 a2820a <=( a30508a  and  a30497a );
 a2821a <=( a30486a  and  a30475a );
 a2822a <=( a30464a  and  a30453a );
 a2823a <=( a30442a  and  a30431a );
 a2824a <=( a30420a  and  a30409a );
 a2825a <=( a30398a  and  a30387a );
 a2826a <=( a30376a  and  a30365a );
 a2827a <=( a30354a  and  a30343a );
 a2828a <=( a30332a  and  a30321a );
 a2829a <=( a30310a  and  a30299a );
 a2830a <=( a30288a  and  a30277a );
 a2831a <=( a30266a  and  a30255a );
 a2832a <=( a30244a  and  a30233a );
 a2833a <=( a30222a  and  a30211a );
 a2834a <=( a30200a  and  a30189a );
 a2835a <=( a30178a  and  a30167a );
 a2836a <=( a30156a  and  a30145a );
 a2837a <=( a30134a  and  a30123a );
 a2838a <=( a30112a  and  a30101a );
 a2839a <=( a30090a  and  a30079a );
 a2840a <=( a30068a  and  a30057a );
 a2841a <=( a30046a  and  a30035a );
 a2842a <=( a30024a  and  a30013a );
 a2843a <=( a30002a  and  a29991a );
 a2844a <=( a29980a  and  a29969a );
 a2845a <=( a29958a  and  a29947a );
 a2846a <=( a29936a  and  a29925a );
 a2847a <=( a29914a  and  a29903a );
 a2848a <=( a29892a  and  a29881a );
 a2849a <=( a29870a  and  a29859a );
 a2850a <=( a29848a  and  a29837a );
 a2851a <=( a29826a  and  a29815a );
 a2852a <=( a29804a  and  a29793a );
 a2853a <=( a29782a  and  a29771a );
 a2854a <=( a29760a  and  a29749a );
 a2855a <=( a29738a  and  a29727a );
 a2856a <=( a29716a  and  a29705a );
 a2857a <=( a29694a  and  a29683a );
 a2858a <=( a29672a  and  a29661a );
 a2859a <=( a29650a  and  a29639a );
 a2860a <=( a29628a  and  a29617a );
 a2861a <=( a29606a  and  a29595a );
 a2862a <=( a29584a  and  a29573a );
 a2863a <=( a29562a  and  a29551a );
 a2864a <=( a29540a  and  a29529a );
 a2865a <=( a29518a  and  a29507a );
 a2866a <=( a29496a  and  a29485a );
 a2867a <=( a29474a  and  a29463a );
 a2868a <=( a29452a  and  a29441a );
 a2869a <=( a29430a  and  a29419a );
 a2870a <=( a29408a  and  a29397a );
 a2871a <=( a29386a  and  a29375a );
 a2872a <=( a29364a  and  a29353a );
 a2873a <=( a29342a  and  a29331a );
 a2874a <=( a29320a  and  a29309a );
 a2875a <=( a29298a  and  a29287a );
 a2876a <=( a29276a  and  a29265a );
 a2877a <=( a29254a  and  a29243a );
 a2878a <=( a29232a  and  a29221a );
 a2879a <=( a29210a  and  a29199a );
 a2880a <=( a29188a  and  a29177a );
 a2881a <=( a29166a  and  a29155a );
 a2882a <=( a29144a  and  a29133a );
 a2883a <=( a29122a  and  a29111a );
 a2884a <=( a29100a  and  a29089a );
 a2885a <=( a29078a  and  a29067a );
 a2886a <=( a29056a  and  a29045a );
 a2887a <=( a29034a  and  a29023a );
 a2888a <=( a29012a  and  a29001a );
 a2889a <=( a28990a  and  a28979a );
 a2890a <=( a28968a  and  a28957a );
 a2891a <=( a28946a  and  a28935a );
 a2892a <=( a28924a  and  a28913a );
 a2893a <=( a28902a  and  a28891a );
 a2894a <=( a28880a  and  a28869a );
 a2895a <=( a28858a  and  a28847a );
 a2896a <=( a28836a  and  a28825a );
 a2897a <=( a28814a  and  a28803a );
 a2898a <=( a28792a  and  a28781a );
 a2899a <=( a28770a  and  a28759a );
 a2900a <=( a28748a  and  a28737a );
 a2901a <=( a28726a  and  a28715a );
 a2902a <=( a28704a  and  a28693a );
 a2903a <=( a28682a  and  a28671a );
 a2904a <=( a28660a  and  a28649a );
 a2905a <=( a28638a  and  a28627a );
 a2906a <=( a28616a  and  a28605a );
 a2907a <=( a28594a  and  a28583a );
 a2908a <=( a28572a  and  a28561a );
 a2909a <=( a28550a  and  a28539a );
 a2910a <=( a28528a  and  a28517a );
 a2911a <=( a28506a  and  a28495a );
 a2912a <=( a28484a  and  a28473a );
 a2913a <=( a28462a  and  a28451a );
 a2914a <=( a28440a  and  a28429a );
 a2915a <=( a28418a  and  a28407a );
 a2916a <=( a28396a  and  a28385a );
 a2917a <=( a28374a  and  a28363a );
 a2918a <=( a28352a  and  a28341a );
 a2919a <=( a28330a  and  a28319a );
 a2920a <=( a28308a  and  a28297a );
 a2921a <=( a28286a  and  a28275a );
 a2922a <=( a28264a  and  a28253a );
 a2923a <=( a28242a  and  a28231a );
 a2924a <=( a28220a  and  a28209a );
 a2925a <=( a28198a  and  a28187a );
 a2926a <=( a28176a  and  a28165a );
 a2927a <=( a28154a  and  a28143a );
 a2928a <=( a28132a  and  a28121a );
 a2929a <=( a28110a  and  a28099a );
 a2930a <=( a28088a  and  a28077a );
 a2931a <=( a28066a  and  a28055a );
 a2932a <=( a28044a  and  a28033a );
 a2933a <=( a28022a  and  a28011a );
 a2934a <=( a28000a  and  a27989a );
 a2935a <=( a27978a  and  a27967a );
 a2936a <=( a27956a  and  a27945a );
 a2937a <=( a27934a  and  a27923a );
 a2938a <=( a27912a  and  a27901a );
 a2939a <=( a27890a  and  a27879a );
 a2940a <=( a27868a  and  a27857a );
 a2941a <=( a27846a  and  a27835a );
 a2942a <=( a27824a  and  a27813a );
 a2943a <=( a27802a  and  a27791a );
 a2944a <=( a27780a  and  a27769a );
 a2945a <=( a27758a  and  a27747a );
 a2946a <=( a27736a  and  a27725a );
 a2947a <=( a27714a  and  a27703a );
 a2948a <=( a27692a  and  a27681a );
 a2949a <=( a27670a  and  a27659a );
 a2950a <=( a27648a  and  a27637a );
 a2951a <=( a27626a  and  a27615a );
 a2952a <=( a27604a  and  a27593a );
 a2953a <=( a27582a  and  a27571a );
 a2954a <=( a27560a  and  a27549a );
 a2955a <=( a27538a  and  a27527a );
 a2956a <=( a27516a  and  a27505a );
 a2957a <=( a27494a  and  a27483a );
 a2958a <=( a27472a  and  a27461a );
 a2959a <=( a27450a  and  a27439a );
 a2960a <=( a27428a  and  a27417a );
 a2961a <=( a27406a  and  a27395a );
 a2962a <=( a27384a  and  a27373a );
 a2963a <=( a27362a  and  a27351a );
 a2964a <=( a27340a  and  a27329a );
 a2965a <=( a27318a  and  a27307a );
 a2966a <=( a27296a  and  a27285a );
 a2967a <=( a27274a  and  a27263a );
 a2968a <=( a27252a  and  a27241a );
 a2969a <=( a27230a  and  a27219a );
 a2970a <=( a27208a  and  a27197a );
 a2971a <=( a27186a  and  a27175a );
 a2972a <=( a27164a  and  a27153a );
 a2973a <=( a27142a  and  a27131a );
 a2974a <=( a27120a  and  a27109a );
 a2975a <=( a27098a  and  a27087a );
 a2976a <=( a27076a  and  a27065a );
 a2977a <=( a27054a  and  a27043a );
 a2978a <=( a27032a  and  a27021a );
 a2979a <=( a27010a  and  a26999a );
 a2980a <=( a26988a  and  a26977a );
 a2981a <=( a26966a  and  a26955a );
 a2982a <=( a26944a  and  a26933a );
 a2983a <=( a26922a  and  a26911a );
 a2984a <=( a26900a  and  a26889a );
 a2985a <=( a26878a  and  a26867a );
 a2986a <=( a26856a  and  a26845a );
 a2987a <=( a26834a  and  a26823a );
 a2988a <=( a26812a  and  a26801a );
 a2989a <=( a26790a  and  a26779a );
 a2990a <=( a26768a  and  a26757a );
 a2991a <=( a26746a  and  a26735a );
 a2992a <=( a26724a  and  a26713a );
 a2993a <=( a26702a  and  a26691a );
 a2994a <=( a26680a  and  a26669a );
 a2995a <=( a26658a  and  a26647a );
 a2996a <=( a26636a  and  a26625a );
 a2997a <=( a26614a  and  a26603a );
 a2998a <=( a26592a  and  a26581a );
 a2999a <=( a26570a  and  a26559a );
 a3000a <=( a26548a  and  a26537a );
 a3001a <=( a26526a  and  a26515a );
 a3002a <=( a26504a  and  a26493a );
 a3003a <=( a26482a  and  a26471a );
 a3004a <=( a26460a  and  a26449a );
 a3005a <=( a26438a  and  a26427a );
 a3006a <=( a26416a  and  a26405a );
 a3007a <=( a26394a  and  a26383a );
 a3008a <=( a26372a  and  a26361a );
 a3009a <=( a26350a  and  a26339a );
 a3010a <=( a26328a  and  a26317a );
 a3011a <=( a26306a  and  a26295a );
 a3012a <=( a26284a  and  a26273a );
 a3013a <=( a26262a  and  a26251a );
 a3014a <=( a26240a  and  a26229a );
 a3015a <=( a26218a  and  a26207a );
 a3016a <=( a26196a  and  a26185a );
 a3017a <=( a26174a  and  a26163a );
 a3018a <=( a26152a  and  a26141a );
 a3019a <=( a26130a  and  a26119a );
 a3020a <=( a26108a  and  a26097a );
 a3021a <=( a26086a  and  a26075a );
 a3022a <=( a26064a  and  a26053a );
 a3023a <=( a26042a  and  a26031a );
 a3024a <=( a26020a  and  a26009a );
 a3025a <=( a25998a  and  a25987a );
 a3026a <=( a25976a  and  a25965a );
 a3027a <=( a25954a  and  a25943a );
 a3028a <=( a25932a  and  a25921a );
 a3029a <=( a25910a  and  a25899a );
 a3030a <=( a25888a  and  a25877a );
 a3031a <=( a25866a  and  a25855a );
 a3032a <=( a25844a  and  a25833a );
 a3033a <=( a25822a  and  a25811a );
 a3034a <=( a25800a  and  a25789a );
 a3035a <=( a25778a  and  a25767a );
 a3036a <=( a25756a  and  a25745a );
 a3037a <=( a25734a  and  a25723a );
 a3038a <=( a25712a  and  a25701a );
 a3039a <=( a25690a  and  a25679a );
 a3040a <=( a25668a  and  a25657a );
 a3041a <=( a25646a  and  a25635a );
 a3042a <=( a25624a  and  a25613a );
 a3043a <=( a25602a  and  a25591a );
 a3044a <=( a25580a  and  a25569a );
 a3045a <=( a25558a  and  a25547a );
 a3046a <=( a25536a  and  a25525a );
 a3047a <=( a25514a  and  a25503a );
 a3048a <=( a25492a  and  a25481a );
 a3049a <=( a25470a  and  a25459a );
 a3050a <=( a25448a  and  a25437a );
 a3051a <=( a25426a  and  a25415a );
 a3052a <=( a25404a  and  a25393a );
 a3053a <=( a25382a  and  a25371a );
 a3054a <=( a25360a  and  a25349a );
 a3055a <=( a25338a  and  a25327a );
 a3056a <=( a25316a  and  a25305a );
 a3057a <=( a25294a  and  a25283a );
 a3058a <=( a25272a  and  a25261a );
 a3059a <=( a25250a  and  a25239a );
 a3060a <=( a25228a  and  a25217a );
 a3061a <=( a25206a  and  a25195a );
 a3062a <=( a25184a  and  a25173a );
 a3063a <=( a25162a  and  a25151a );
 a3064a <=( a25140a  and  a25129a );
 a3065a <=( a25118a  and  a25107a );
 a3066a <=( a25096a  and  a25085a );
 a3067a <=( a25074a  and  a25063a );
 a3068a <=( a25052a  and  a25041a );
 a3069a <=( a25030a  and  a25019a );
 a3070a <=( a25008a  and  a24997a );
 a3071a <=( a24986a  and  a24975a );
 a3072a <=( a24964a  and  a24953a );
 a3073a <=( a24942a  and  a24931a );
 a3074a <=( a24920a  and  a24909a );
 a3075a <=( a24898a  and  a24887a );
 a3076a <=( a24876a  and  a24865a );
 a3077a <=( a24854a  and  a24843a );
 a3078a <=( a24832a  and  a24821a );
 a3079a <=( a24810a  and  a24799a );
 a3080a <=( a24788a  and  a24777a );
 a3081a <=( a24766a  and  a24755a );
 a3082a <=( a24744a  and  a24733a );
 a3083a <=( a24722a  and  a24711a );
 a3084a <=( a24700a  and  a24689a );
 a3085a <=( a24678a  and  a24667a );
 a3086a <=( a24656a  and  a24645a );
 a3087a <=( a24634a  and  a24623a );
 a3088a <=( a24612a  and  a24601a );
 a3089a <=( a24590a  and  a24579a );
 a3090a <=( a24568a  and  a24557a );
 a3091a <=( a24546a  and  a24535a );
 a3092a <=( a24524a  and  a24513a );
 a3093a <=( a24502a  and  a24491a );
 a3094a <=( a24480a  and  a24469a );
 a3095a <=( a24458a  and  a24447a );
 a3096a <=( a24436a  and  a24425a );
 a3097a <=( a24414a  and  a24403a );
 a3098a <=( a24392a  and  a24381a );
 a3099a <=( a24370a  and  a24359a );
 a3100a <=( a24348a  and  a24337a );
 a3101a <=( a24326a  and  a24315a );
 a3102a <=( a24304a  and  a24293a );
 a3103a <=( a24282a  and  a24271a );
 a3104a <=( a24260a  and  a24249a );
 a3105a <=( a24238a  and  a24227a );
 a3106a <=( a24216a  and  a24205a );
 a3107a <=( a24194a  and  a24183a );
 a3108a <=( a24172a  and  a24161a );
 a3109a <=( a24150a  and  a24139a );
 a3110a <=( a24128a  and  a24117a );
 a3111a <=( a24106a  and  a24095a );
 a3112a <=( a24084a  and  a24073a );
 a3113a <=( a24062a  and  a24051a );
 a3114a <=( a24040a  and  a24029a );
 a3115a <=( a24018a  and  a24007a );
 a3116a <=( a23996a  and  a23985a );
 a3117a <=( a23974a  and  a23963a );
 a3118a <=( a23952a  and  a23941a );
 a3119a <=( a23930a  and  a23919a );
 a3120a <=( a23908a  and  a23897a );
 a3121a <=( a23886a  and  a23875a );
 a3122a <=( a23864a  and  a23853a );
 a3123a <=( a23842a  and  a23831a );
 a3124a <=( a23820a  and  a23809a );
 a3125a <=( a23798a  and  a23787a );
 a3126a <=( a23776a  and  a23765a );
 a3127a <=( a23754a  and  a23743a );
 a3128a <=( a23732a  and  a23721a );
 a3129a <=( a23710a  and  a23699a );
 a3130a <=( a23688a  and  a23677a );
 a3131a <=( a23666a  and  a23655a );
 a3132a <=( a23644a  and  a23633a );
 a3133a <=( a23622a  and  a23611a );
 a3134a <=( a23600a  and  a23589a );
 a3135a <=( a23578a  and  a23567a );
 a3136a <=( a23556a  and  a23545a );
 a3137a <=( a23534a  and  a23523a );
 a3138a <=( a23512a  and  a23501a );
 a3139a <=( a23490a  and  a23479a );
 a3140a <=( a23468a  and  a23457a );
 a3141a <=( a23446a  and  a23435a );
 a3142a <=( a23424a  and  a23413a );
 a3143a <=( a23402a  and  a23391a );
 a3144a <=( a23380a  and  a23369a );
 a3145a <=( a23358a  and  a23347a );
 a3146a <=( a23336a  and  a23325a );
 a3147a <=( a23314a  and  a23303a );
 a3148a <=( a23292a  and  a23281a );
 a3149a <=( a23270a  and  a23259a );
 a3150a <=( a23248a  and  a23237a );
 a3151a <=( a23226a  and  a23215a );
 a3152a <=( a23204a  and  a23193a );
 a3153a <=( a23182a  and  a23171a );
 a3154a <=( a23160a  and  a23149a );
 a3155a <=( a23138a  and  a23127a );
 a3156a <=( a23116a  and  a23105a );
 a3157a <=( a23094a  and  a23083a );
 a3158a <=( a23072a  and  a23061a );
 a3159a <=( a23050a  and  a23039a );
 a3160a <=( a23028a  and  a23017a );
 a3161a <=( a23006a  and  a22995a );
 a3162a <=( a22984a  and  a22973a );
 a3163a <=( a22962a  and  a22951a );
 a3164a <=( a22940a  and  a22929a );
 a3165a <=( a22918a  and  a22907a );
 a3166a <=( a22896a  and  a22885a );
 a3167a <=( a22874a  and  a22863a );
 a3168a <=( a22852a  and  a22841a );
 a3169a <=( a22830a  and  a22819a );
 a3170a <=( a22808a  and  a22797a );
 a3171a <=( a22786a  and  a22775a );
 a3172a <=( a22764a  and  a22753a );
 a3173a <=( a22742a  and  a22731a );
 a3174a <=( a22720a  and  a22709a );
 a3175a <=( a22698a  and  a22687a );
 a3176a <=( a22676a  and  a22665a );
 a3177a <=( a22654a  and  a22643a );
 a3178a <=( a22632a  and  a22621a );
 a3179a <=( a22610a  and  a22599a );
 a3180a <=( a22588a  and  a22577a );
 a3181a <=( a22566a  and  a22555a );
 a3182a <=( a22544a  and  a22533a );
 a3183a <=( a22522a  and  a22511a );
 a3184a <=( a22500a  and  a22489a );
 a3185a <=( a22478a  and  a22467a );
 a3186a <=( a22458a  and  a22447a );
 a3187a <=( a22438a  and  a22427a );
 a3188a <=( a22418a  and  a22407a );
 a3189a <=( a22398a  and  a22387a );
 a3190a <=( a22378a  and  a22367a );
 a3191a <=( a22358a  and  a22347a );
 a3192a <=( a22338a  and  a22327a );
 a3193a <=( a22318a  and  a22307a );
 a3194a <=( a22298a  and  a22287a );
 a3195a <=( a22278a  and  a22267a );
 a3196a <=( a22258a  and  a22247a );
 a3197a <=( a22238a  and  a22227a );
 a3198a <=( a22218a  and  a22207a );
 a3199a <=( a22198a  and  a22187a );
 a3200a <=( a22178a  and  a22167a );
 a3201a <=( a22158a  and  a22147a );
 a3202a <=( a22138a  and  a22127a );
 a3203a <=( a22118a  and  a22107a );
 a3204a <=( a22098a  and  a22087a );
 a3205a <=( a22078a  and  a22067a );
 a3206a <=( a22058a  and  a22047a );
 a3207a <=( a22038a  and  a22027a );
 a3208a <=( a22018a  and  a22007a );
 a3209a <=( a21998a  and  a21987a );
 a3210a <=( a21978a  and  a21967a );
 a3211a <=( a21958a  and  a21947a );
 a3212a <=( a21938a  and  a21927a );
 a3213a <=( a21918a  and  a21907a );
 a3214a <=( a21898a  and  a21887a );
 a3215a <=( a21878a  and  a21867a );
 a3216a <=( a21858a  and  a21847a );
 a3217a <=( a21838a  and  a21827a );
 a3218a <=( a21818a  and  a21807a );
 a3219a <=( a21798a  and  a21787a );
 a3220a <=( a21778a  and  a21767a );
 a3221a <=( a21758a  and  a21747a );
 a3222a <=( a21738a  and  a21727a );
 a3223a <=( a21718a  and  a21707a );
 a3224a <=( a21698a  and  a21687a );
 a3225a <=( a21678a  and  a21667a );
 a3226a <=( a21658a  and  a21647a );
 a3227a <=( a21638a  and  a21627a );
 a3228a <=( a21618a  and  a21607a );
 a3229a <=( a21598a  and  a21587a );
 a3230a <=( a21578a  and  a21567a );
 a3231a <=( a21558a  and  a21547a );
 a3232a <=( a21538a  and  a21527a );
 a3233a <=( a21518a  and  a21507a );
 a3234a <=( a21498a  and  a21487a );
 a3235a <=( a21478a  and  a21467a );
 a3236a <=( a21458a  and  a21447a );
 a3237a <=( a21438a  and  a21427a );
 a3238a <=( a21418a  and  a21407a );
 a3239a <=( a21398a  and  a21387a );
 a3240a <=( a21378a  and  a21367a );
 a3241a <=( a21358a  and  a21347a );
 a3242a <=( a21338a  and  a21327a );
 a3243a <=( a21318a  and  a21307a );
 a3244a <=( a21298a  and  a21287a );
 a3245a <=( a21278a  and  a21267a );
 a3246a <=( a21258a  and  a21247a );
 a3247a <=( a21238a  and  a21227a );
 a3248a <=( a21218a  and  a21207a );
 a3249a <=( a21198a  and  a21187a );
 a3250a <=( a21178a  and  a21167a );
 a3251a <=( a21158a  and  a21147a );
 a3252a <=( a21138a  and  a21127a );
 a3253a <=( a21118a  and  a21107a );
 a3254a <=( a21098a  and  a21087a );
 a3255a <=( a21078a  and  a21067a );
 a3256a <=( a21058a  and  a21047a );
 a3257a <=( a21038a  and  a21027a );
 a3258a <=( a21018a  and  a21007a );
 a3259a <=( a20998a  and  a20987a );
 a3260a <=( a20978a  and  a20967a );
 a3261a <=( a20958a  and  a20947a );
 a3262a <=( a20938a  and  a20927a );
 a3263a <=( a20918a  and  a20907a );
 a3264a <=( a20898a  and  a20887a );
 a3265a <=( a20878a  and  a20867a );
 a3266a <=( a20858a  and  a20847a );
 a3267a <=( a20838a  and  a20827a );
 a3268a <=( a20818a  and  a20807a );
 a3269a <=( a20798a  and  a20787a );
 a3270a <=( a20778a  and  a20767a );
 a3271a <=( a20758a  and  a20747a );
 a3272a <=( a20738a  and  a20727a );
 a3273a <=( a20718a  and  a20707a );
 a3274a <=( a20698a  and  a20687a );
 a3275a <=( a20678a  and  a20667a );
 a3276a <=( a20658a  and  a20647a );
 a3277a <=( a20638a  and  a20627a );
 a3278a <=( a20618a  and  a20607a );
 a3279a <=( a20598a  and  a20587a );
 a3280a <=( a20578a  and  a20567a );
 a3281a <=( a20558a  and  a20547a );
 a3282a <=( a20538a  and  a20527a );
 a3283a <=( a20518a  and  a20507a );
 a3284a <=( a20498a  and  a20487a );
 a3285a <=( a20478a  and  a20467a );
 a3286a <=( a20458a  and  a20447a );
 a3287a <=( a20438a  and  a20427a );
 a3288a <=( a20418a  and  a20407a );
 a3289a <=( a20398a  and  a20387a );
 a3290a <=( a20378a  and  a20367a );
 a3291a <=( a20358a  and  a20347a );
 a3292a <=( a20338a  and  a20327a );
 a3293a <=( a20318a  and  a20307a );
 a3294a <=( a20298a  and  a20287a );
 a3295a <=( a20278a  and  a20267a );
 a3296a <=( a20258a  and  a20247a );
 a3297a <=( a20238a  and  a20227a );
 a3298a <=( a20218a  and  a20207a );
 a3299a <=( a20198a  and  a20187a );
 a3300a <=( a20178a  and  a20167a );
 a3301a <=( a20158a  and  a20147a );
 a3302a <=( a20138a  and  a20127a );
 a3303a <=( a20118a  and  a20107a );
 a3304a <=( a20098a  and  a20087a );
 a3305a <=( a20078a  and  a20067a );
 a3306a <=( a20058a  and  a20047a );
 a3307a <=( a20038a  and  a20027a );
 a3308a <=( a20018a  and  a20007a );
 a3309a <=( a19998a  and  a19987a );
 a3310a <=( a19978a  and  a19967a );
 a3311a <=( a19958a  and  a19947a );
 a3312a <=( a19938a  and  a19927a );
 a3313a <=( a19918a  and  a19907a );
 a3314a <=( a19898a  and  a19887a );
 a3315a <=( a19878a  and  a19867a );
 a3316a <=( a19858a  and  a19847a );
 a3317a <=( a19838a  and  a19827a );
 a3318a <=( a19818a  and  a19807a );
 a3319a <=( a19798a  and  a19787a );
 a3320a <=( a19778a  and  a19767a );
 a3321a <=( a19758a  and  a19747a );
 a3322a <=( a19738a  and  a19727a );
 a3323a <=( a19718a  and  a19707a );
 a3324a <=( a19698a  and  a19687a );
 a3325a <=( a19678a  and  a19667a );
 a3326a <=( a19658a  and  a19647a );
 a3327a <=( a19638a  and  a19627a );
 a3328a <=( a19618a  and  a19607a );
 a3329a <=( a19598a  and  a19587a );
 a3330a <=( a19578a  and  a19567a );
 a3331a <=( a19558a  and  a19547a );
 a3332a <=( a19538a  and  a19527a );
 a3333a <=( a19518a  and  a19507a );
 a3334a <=( a19498a  and  a19487a );
 a3335a <=( a19478a  and  a19467a );
 a3336a <=( a19458a  and  a19447a );
 a3337a <=( a19438a  and  a19427a );
 a3338a <=( a19418a  and  a19407a );
 a3339a <=( a19398a  and  a19387a );
 a3340a <=( a19378a  and  a19367a );
 a3341a <=( a19358a  and  a19347a );
 a3342a <=( a19338a  and  a19327a );
 a3343a <=( a19318a  and  a19307a );
 a3344a <=( a19298a  and  a19287a );
 a3345a <=( a19278a  and  a19267a );
 a3346a <=( a19258a  and  a19247a );
 a3347a <=( a19238a  and  a19227a );
 a3348a <=( a19218a  and  a19207a );
 a3349a <=( a19198a  and  a19187a );
 a3350a <=( a19178a  and  a19167a );
 a3351a <=( a19158a  and  a19147a );
 a3352a <=( a19138a  and  a19127a );
 a3353a <=( a19118a  and  a19107a );
 a3354a <=( a19098a  and  a19087a );
 a3355a <=( a19078a  and  a19067a );
 a3356a <=( a19058a  and  a19047a );
 a3357a <=( a19038a  and  a19027a );
 a3358a <=( a19018a  and  a19007a );
 a3359a <=( a18998a  and  a18987a );
 a3360a <=( a18978a  and  a18967a );
 a3361a <=( a18958a  and  a18947a );
 a3362a <=( a18938a  and  a18927a );
 a3363a <=( a18918a  and  a18907a );
 a3364a <=( a18898a  and  a18887a );
 a3365a <=( a18878a  and  a18867a );
 a3366a <=( a18858a  and  a18847a );
 a3367a <=( a18838a  and  a18827a );
 a3368a <=( a18818a  and  a18807a );
 a3369a <=( a18798a  and  a18787a );
 a3370a <=( a18778a  and  a18767a );
 a3371a <=( a18758a  and  a18747a );
 a3372a <=( a18738a  and  a18727a );
 a3373a <=( a18718a  and  a18707a );
 a3374a <=( a18698a  and  a18687a );
 a3375a <=( a18678a  and  a18667a );
 a3376a <=( a18658a  and  a18647a );
 a3377a <=( a18638a  and  a18627a );
 a3378a <=( a18618a  and  a18607a );
 a3379a <=( a18598a  and  a18587a );
 a3380a <=( a18578a  and  a18567a );
 a3381a <=( a18558a  and  a18547a );
 a3382a <=( a18538a  and  a18527a );
 a3383a <=( a18518a  and  a18507a );
 a3384a <=( a18498a  and  a18487a );
 a3385a <=( a18478a  and  a18467a );
 a3386a <=( a18458a  and  a18447a );
 a3387a <=( a18438a  and  a18427a );
 a3388a <=( a18418a  and  a18407a );
 a3389a <=( a18398a  and  a18387a );
 a3390a <=( a18378a  and  a18367a );
 a3391a <=( a18358a  and  a18347a );
 a3392a <=( a18338a  and  a18327a );
 a3393a <=( a18318a  and  a18307a );
 a3394a <=( a18298a  and  a18287a );
 a3395a <=( a18278a  and  a18267a );
 a3396a <=( a18258a  and  a18247a );
 a3397a <=( a18238a  and  a18227a );
 a3398a <=( a18218a  and  a18207a );
 a3399a <=( a18198a  and  a18187a );
 a3400a <=( a18178a  and  a18167a );
 a3401a <=( a18158a  and  a18147a );
 a3402a <=( a18138a  and  a18127a );
 a3403a <=( a18118a  and  a18107a );
 a3404a <=( a18098a  and  a18087a );
 a3405a <=( a18078a  and  a18067a );
 a3406a <=( a18058a  and  a18047a );
 a3407a <=( a18038a  and  a18027a );
 a3408a <=( a18018a  and  a18007a );
 a3409a <=( a17998a  and  a17987a );
 a3410a <=( a17978a  and  a17967a );
 a3411a <=( a17958a  and  a17947a );
 a3412a <=( a17938a  and  a17927a );
 a3413a <=( a17918a  and  a17907a );
 a3414a <=( a17898a  and  a17887a );
 a3415a <=( a17878a  and  a17867a );
 a3416a <=( a17858a  and  a17847a );
 a3417a <=( a17838a  and  a17827a );
 a3418a <=( a17818a  and  a17807a );
 a3419a <=( a17798a  and  a17787a );
 a3420a <=( a17778a  and  a17767a );
 a3421a <=( a17758a  and  a17747a );
 a3422a <=( a17738a  and  a17727a );
 a3423a <=( a17718a  and  a17707a );
 a3424a <=( a17698a  and  a17687a );
 a3425a <=( a17678a  and  a17667a );
 a3426a <=( a17658a  and  a17647a );
 a3427a <=( a17638a  and  a17627a );
 a3428a <=( a17618a  and  a17607a );
 a3429a <=( a17598a  and  a17587a );
 a3430a <=( a17578a  and  a17567a );
 a3431a <=( a17558a  and  a17547a );
 a3432a <=( a17538a  and  a17527a );
 a3433a <=( a17518a  and  a17507a );
 a3434a <=( a17498a  and  a17487a );
 a3435a <=( a17478a  and  a17467a );
 a3436a <=( a17458a  and  a17447a );
 a3437a <=( a17438a  and  a17427a );
 a3438a <=( a17418a  and  a17407a );
 a3439a <=( a17398a  and  a17387a );
 a3440a <=( a17378a  and  a17367a );
 a3441a <=( a17358a  and  a17347a );
 a3442a <=( a17338a  and  a17327a );
 a3443a <=( a17318a  and  a17307a );
 a3444a <=( a17298a  and  a17287a );
 a3445a <=( a17278a  and  a17267a );
 a3446a <=( a17258a  and  a17247a );
 a3447a <=( a17238a  and  a17227a );
 a3448a <=( a17218a  and  a17207a );
 a3449a <=( a17198a  and  a17187a );
 a3450a <=( a17178a  and  a17167a );
 a3451a <=( a17158a  and  a17147a );
 a3452a <=( a17138a  and  a17127a );
 a3453a <=( a17118a  and  a17107a );
 a3454a <=( a17098a  and  a17087a );
 a3455a <=( a17078a  and  a17067a );
 a3456a <=( a17058a  and  a17047a );
 a3457a <=( a17038a  and  a17027a );
 a3458a <=( a17018a  and  a17007a );
 a3459a <=( a16998a  and  a16987a );
 a3460a <=( a16978a  and  a16967a );
 a3461a <=( a16958a  and  a16947a );
 a3462a <=( a16938a  and  a16927a );
 a3463a <=( a16918a  and  a16907a );
 a3464a <=( a16898a  and  a16887a );
 a3465a <=( a16878a  and  a16867a );
 a3466a <=( a16858a  and  a16847a );
 a3467a <=( a16838a  and  a16827a );
 a3468a <=( a16818a  and  a16807a );
 a3469a <=( a16798a  and  a16787a );
 a3470a <=( a16778a  and  a16767a );
 a3471a <=( a16758a  and  a16747a );
 a3472a <=( a16738a  and  a16727a );
 a3473a <=( a16718a  and  a16707a );
 a3474a <=( a16698a  and  a16687a );
 a3475a <=( a16678a  and  a16667a );
 a3476a <=( a16658a  and  a16647a );
 a3477a <=( a16638a  and  a16627a );
 a3478a <=( a16618a  and  a16607a );
 a3479a <=( a16598a  and  a16587a );
 a3480a <=( a16578a  and  a16567a );
 a3481a <=( a16558a  and  a16547a );
 a3482a <=( a16538a  and  a16527a );
 a3483a <=( a16518a  and  a16507a );
 a3484a <=( a16498a  and  a16487a );
 a3485a <=( a16478a  and  a16467a );
 a3486a <=( a16458a  and  a16447a );
 a3487a <=( a16438a  and  a16427a );
 a3488a <=( a16418a  and  a16407a );
 a3489a <=( a16398a  and  a16387a );
 a3490a <=( a16378a  and  a16367a );
 a3491a <=( a16358a  and  a16347a );
 a3492a <=( a16338a  and  a16327a );
 a3493a <=( a16318a  and  a16307a );
 a3494a <=( a16298a  and  a16287a );
 a3495a <=( a16278a  and  a16267a );
 a3496a <=( a16258a  and  a16247a );
 a3497a <=( a16238a  and  a16227a );
 a3498a <=( a16218a  and  a16207a );
 a3499a <=( a16198a  and  a16187a );
 a3500a <=( a16178a  and  a16167a );
 a3501a <=( a16158a  and  a16147a );
 a3502a <=( a16138a  and  a16127a );
 a3503a <=( a16118a  and  a16107a );
 a3504a <=( a16098a  and  a16087a );
 a3505a <=( a16078a  and  a16067a );
 a3506a <=( a16058a  and  a16047a );
 a3507a <=( a16038a  and  a16029a );
 a3508a <=( a16020a  and  a16011a );
 a3509a <=( a16002a  and  a15993a );
 a3510a <=( a15984a  and  a15975a );
 a3511a <=( a15966a  and  a15957a );
 a3512a <=( a15948a  and  a15939a );
 a3513a <=( a15930a  and  a15921a );
 a3514a <=( a15912a  and  a15903a );
 a3515a <=( a15894a  and  a15885a );
 a3516a <=( a15876a  and  a15867a );
 a3517a <=( a15858a  and  a15849a );
 a3518a <=( a15840a  and  a15831a );
 a3519a <=( a15822a  and  a15813a );
 a3520a <=( a15804a  and  a15795a );
 a3521a <=( a15786a  and  a15777a );
 a3522a <=( a15768a  and  a15759a );
 a3523a <=( a15750a  and  a15741a );
 a3524a <=( a15732a  and  a15723a );
 a3525a <=( a15714a  and  a15705a );
 a3526a <=( a15696a  and  a15687a );
 a3527a <=( a15678a  and  a15669a );
 a3528a <=( a15660a  and  a15651a );
 a3529a <=( a15642a  and  a15633a );
 a3530a <=( a15624a  and  a15615a );
 a3531a <=( a15606a  and  a15597a );
 a3532a <=( a15588a  and  a15579a );
 a3533a <=( a15570a  and  a15561a );
 a3534a <=( a15552a  and  a15543a );
 a3535a <=( a15534a  and  a15525a );
 a3536a <=( a15516a  and  a15507a );
 a3537a <=( a15498a  and  a15489a );
 a3538a <=( a15480a  and  a15471a );
 a3539a <=( a15462a  and  a15453a );
 a3540a <=( a15444a  and  a15435a );
 a3541a <=( a15426a  and  a15417a );
 a3542a <=( a15408a  and  a15399a );
 a3543a <=( a15390a  and  a15381a );
 a3544a <=( a15372a  and  a15363a );
 a3545a <=( a15354a  and  a15345a );
 a3546a <=( a15336a  and  a15327a );
 a3547a <=( a15318a  and  a15309a );
 a3548a <=( a15300a  and  a15291a );
 a3549a <=( a15282a  and  a15273a );
 a3550a <=( a15264a  and  a15255a );
 a3551a <=( a15246a  and  a15237a );
 a3552a <=( a15228a  and  a15219a );
 a3553a <=( a15210a  and  a15201a );
 a3554a <=( a15192a  and  a15183a );
 a3555a <=( a15174a  and  a15165a );
 a3556a <=( a15156a  and  a15147a );
 a3557a <=( a15138a  and  a15129a );
 a3558a <=( a15120a  and  a15111a );
 a3559a <=( a15102a  and  a15093a );
 a3560a <=( a15084a  and  a15075a );
 a3561a <=( a15066a  and  a15057a );
 a3562a <=( a15048a  and  a15039a );
 a3563a <=( a15030a  and  a15021a );
 a3564a <=( a15012a  and  a15003a );
 a3565a <=( a14994a  and  a14985a );
 a3566a <=( a14976a  and  a14967a );
 a3567a <=( a14958a  and  a14949a );
 a3568a <=( a14940a  and  a14931a );
 a3569a <=( a14922a  and  a14913a );
 a3570a <=( a14904a  and  a14895a );
 a3571a <=( a14886a  and  a14877a );
 a3572a <=( a14868a  and  a14859a );
 a3573a <=( a14850a  and  a14841a );
 a3574a <=( a14832a  and  a14823a );
 a3575a <=( a14814a  and  a14805a );
 a3576a <=( a14796a  and  a14787a );
 a3577a <=( a14778a  and  a14769a );
 a3578a <=( a14760a  and  a14751a );
 a3579a <=( a14742a  and  a14733a );
 a3580a <=( a14724a  and  a14715a );
 a3581a <=( a14706a  and  a14697a );
 a3582a <=( a14688a  and  a14679a );
 a3583a <=( a14670a  and  a14661a );
 a3584a <=( a14652a  and  a14643a );
 a3585a <=( a14634a  and  a14625a );
 a3586a <=( a14616a  and  a14607a );
 a3587a <=( a14598a  and  a14589a );
 a3588a <=( a14580a  and  a14571a );
 a3589a <=( a14562a  and  a14553a );
 a3590a <=( a14544a  and  a14535a );
 a3591a <=( a14526a  and  a14517a );
 a3592a <=( a14508a  and  a14499a );
 a3593a <=( a14490a  and  a14481a );
 a3594a <=( a14472a  and  a14463a );
 a3595a <=( a14454a  and  a14445a );
 a3596a <=( a14436a  and  a14427a );
 a3597a <=( a14418a  and  a14409a );
 a3598a <=( a14400a  and  a14391a );
 a3599a <=( a14382a  and  a14373a );
 a3600a <=( a14364a  and  a14355a );
 a3601a <=( a14346a  and  a14337a );
 a3602a <=( a14328a  and  a14319a );
 a3603a <=( a14310a  and  a14301a );
 a3604a <=( a14292a  and  a14283a );
 a3605a <=( a14274a  and  a14265a );
 a3606a <=( a14256a  and  a14247a );
 a3607a <=( a14238a  and  a14229a );
 a3608a <=( a14220a  and  a14211a );
 a3609a <=( a14202a  and  a14193a );
 a3610a <=( a14184a  and  a14175a );
 a3611a <=( a14166a  and  a14157a );
 a3612a <=( a14148a  and  a14139a );
 a3613a <=( a14130a  and  a14121a );
 a3614a <=( a14112a  and  a14103a );
 a3615a <=( a14094a  and  a14085a );
 a3616a <=( a14076a  and  a14067a );
 a3617a <=( a14058a  and  a14049a );
 a3618a <=( a14040a  and  a14031a );
 a3619a <=( a14022a  and  a14013a );
 a3620a <=( a14004a  and  a13995a );
 a3621a <=( a13986a  and  a13977a );
 a3622a <=( a13968a  and  a13959a );
 a3623a <=( a13950a  and  a13941a );
 a3624a <=( a13932a  and  a13923a );
 a3625a <=( a13914a  and  a13905a );
 a3626a <=( a13896a  and  a13887a );
 a3627a <=( a13878a  and  a13869a );
 a3628a <=( a13860a  and  a13851a );
 a3629a <=( a13842a  and  a13833a );
 a3630a <=( a13824a  and  a13815a );
 a3631a <=( a13806a  and  a13797a );
 a3632a <=( a13788a  and  a13779a );
 a3633a <=( a13770a  and  a13761a );
 a3634a <=( a13752a  and  a13743a );
 a3635a <=( a13734a  and  a13725a );
 a3636a <=( a13716a  and  a13707a );
 a3637a <=( a13698a  and  a13689a );
 a3638a <=( a13680a  and  a13671a );
 a3639a <=( a13662a  and  a13653a );
 a3640a <=( a13644a  and  a13635a );
 a3641a <=( a13626a  and  a13617a );
 a3642a <=( a13608a  and  a13599a );
 a3643a <=( a13590a  and  a13581a );
 a3644a <=( a13572a  and  a13563a );
 a3645a <=( a13554a  and  a13545a );
 a3646a <=( a13536a  and  a13527a );
 a3647a <=( a13518a  and  a13509a );
 a3648a <=( a13500a  and  a13491a );
 a3649a <=( a13482a  and  a13473a );
 a3650a <=( a13464a  and  a13455a );
 a3651a <=( a13446a  and  a13437a );
 a3652a <=( a13428a  and  a13419a );
 a3653a <=( a13410a  and  a13401a );
 a3654a <=( a13392a  and  a13383a );
 a3655a <=( a13374a  and  a13365a );
 a3656a <=( a13356a  and  a13347a );
 a3657a <=( a13338a  and  a13329a );
 a3658a <=( a13320a  and  a13311a );
 a3659a <=( a13302a  and  a13293a );
 a3660a <=( a13284a  and  a13275a );
 a3661a <=( a13266a  and  a13257a );
 a3662a <=( a13248a  and  a13239a );
 a3663a <=( a13230a  and  a13221a );
 a3664a <=( a13212a  and  a13203a );
 a3665a <=( a13194a  and  a13185a );
 a3666a <=( a13176a  and  a13167a );
 a3667a <=( a13158a  and  a13149a );
 a3668a <=( a13140a  and  a13131a );
 a3669a <=( a13122a  and  a13113a );
 a3670a <=( a13104a  and  a13095a );
 a3671a <=( a13086a  and  a13077a );
 a3672a <=( a13068a  and  a13059a );
 a3673a <=( a13050a  and  a13041a );
 a3674a <=( a13032a  and  a13023a );
 a3675a <=( a13014a  and  a13005a );
 a3676a <=( a12996a  and  a12987a );
 a3677a <=( a12978a  and  a12969a );
 a3678a <=( a12960a  and  a12951a );
 a3679a <=( a12942a  and  a12933a );
 a3680a <=( a12924a  and  a12915a );
 a3681a <=( a12906a  and  a12897a );
 a3682a <=( a12888a  and  a12879a );
 a3683a <=( a12870a  and  a12861a );
 a3684a <=( a12852a  and  a12843a );
 a3685a <=( a12834a  and  a12825a );
 a3686a <=( a12816a  and  a12807a );
 a3687a <=( a12798a  and  a12789a );
 a3688a <=( a12780a  and  a12771a );
 a3689a <=( a12762a  and  a12753a );
 a3690a <=( a12744a  and  a12735a );
 a3691a <=( a12726a  and  a12717a );
 a3692a <=( a12708a  and  a12699a );
 a3693a <=( a12690a  and  a12681a );
 a3694a <=( a12672a  and  a12663a );
 a3695a <=( a12654a  and  a12645a );
 a3696a <=( a12636a  and  a12627a );
 a3697a <=( a12618a  and  a12609a );
 a3698a <=( a12600a  and  a12591a );
 a3699a <=( a12582a  and  a12573a );
 a3700a <=( a12564a  and  a12555a );
 a3701a <=( a12546a  and  a12537a );
 a3702a <=( a12528a  and  a12519a );
 a3703a <=( a12510a  and  a12501a );
 a3704a <=( a12492a  and  a12483a );
 a3705a <=( a12474a  and  a12465a );
 a3706a <=( a12456a  and  a12447a );
 a3707a <=( a12438a  and  a12429a );
 a3708a <=( a12420a  and  a12411a );
 a3709a <=( a12402a  and  a12393a );
 a3710a <=( a12384a  and  a12375a );
 a3711a <=( a12366a  and  a12357a );
 a3712a <=( a12348a  and  a12339a );
 a3713a <=( a12330a  and  a12321a );
 a3714a <=( a12312a  and  a12303a );
 a3715a <=( a12294a  and  a12285a );
 a3716a <=( a12276a  and  a12267a );
 a3717a <=( a12258a  and  a12249a );
 a3718a <=( a12240a  and  a12231a );
 a3719a <=( a12222a  and  a12213a );
 a3720a <=( a12204a  and  a12195a );
 a3721a <=( a12186a  and  a12177a );
 a3722a <=( a12168a  and  a12159a );
 a3723a <=( a12150a  and  a12141a );
 a3724a <=( a12132a  and  a12123a );
 a3725a <=( a12114a  and  a12105a );
 a3726a <=( a12096a  and  a12087a );
 a3727a <=( a12078a  and  a12069a );
 a3728a <=( a12060a  and  a12051a );
 a3729a <=( a12042a  and  a12033a );
 a3730a <=( a12024a  and  a12015a );
 a3731a <=( a12006a  and  a11997a );
 a3732a <=( a11988a  and  a11979a );
 a3733a <=( a11970a  and  a11961a );
 a3734a <=( a11952a  and  a11943a );
 a3735a <=( a11934a  and  a11925a );
 a3736a <=( a11916a  and  a11907a );
 a3737a <=( a11898a  and  a11889a );
 a3738a <=( a11880a  and  a11871a );
 a3739a <=( a11862a  and  a11853a );
 a3740a <=( a11844a  and  a11835a );
 a3741a <=( a11826a  and  a11817a );
 a3742a <=( a11808a  and  a11799a );
 a3743a <=( a11790a  and  a11781a );
 a3744a <=( a11772a  and  a11763a );
 a3745a <=( a11754a  and  a11745a );
 a3746a <=( a11736a  and  a11727a );
 a3747a <=( a11718a  and  a11709a );
 a3748a <=( a11700a  and  a11691a );
 a3749a <=( a11682a  and  a11673a );
 a3750a <=( a11664a  and  a11655a );
 a3751a <=( a11646a  and  a11637a );
 a3752a <=( a11628a  and  a11619a );
 a3753a <=( a11610a  and  a11601a );
 a3754a <=( a11594a  and  a11585a );
 a3755a <=( a11578a  and  a11569a );
 a3756a <=( a11562a  and  a11553a );
 a3757a <=( a11546a  and  a11537a );
 a3758a <=( a11530a  and  a11521a );
 a3759a <=( a11514a  and  a11505a );
 a3760a <=( a11498a  and  a11489a );
 a3761a <=( a11482a  and  a11475a );
 a3762a <=( a11468a  and  a11461a );
 a3763a <=( a11454a  and  a11447a );
 a3764a <=( a11440a  and  a11433a );
 a3765a <=( a11426a  and  a11419a );
 a3766a <=( a11412a  and  a11405a );
 a3767a <=( a11398a  and  a11391a );
 a3768a <=( a11384a  and  a11377a );
 a3769a <=( a11370a  and  a11363a );
 a3770a <=( a11356a  and  a11349a );
 a3771a <=( a11342a  and  a11335a );
 a3772a <=( a11328a  and  a11321a );
 a3776a <=( a3770a ) or ( a3771a );
 a3777a <=( a3772a ) or ( a3776a );
 a3780a <=( a3768a ) or ( a3769a );
 a3783a <=( a3766a ) or ( a3767a );
 a3784a <=( a3783a ) or ( a3780a );
 a3785a <=( a3784a ) or ( a3777a );
 a3789a <=( a3763a ) or ( a3764a );
 a3790a <=( a3765a ) or ( a3789a );
 a3793a <=( a3761a ) or ( a3762a );
 a3796a <=( a3759a ) or ( a3760a );
 a3797a <=( a3796a ) or ( a3793a );
 a3798a <=( a3797a ) or ( a3790a );
 a3799a <=( a3798a ) or ( a3785a );
 a3803a <=( a3756a ) or ( a3757a );
 a3804a <=( a3758a ) or ( a3803a );
 a3807a <=( a3754a ) or ( a3755a );
 a3810a <=( a3752a ) or ( a3753a );
 a3811a <=( a3810a ) or ( a3807a );
 a3812a <=( a3811a ) or ( a3804a );
 a3815a <=( a3750a ) or ( a3751a );
 a3818a <=( a3748a ) or ( a3749a );
 a3819a <=( a3818a ) or ( a3815a );
 a3822a <=( a3746a ) or ( a3747a );
 a3825a <=( a3744a ) or ( a3745a );
 a3826a <=( a3825a ) or ( a3822a );
 a3827a <=( a3826a ) or ( a3819a );
 a3828a <=( a3827a ) or ( a3812a );
 a3829a <=( a3828a ) or ( a3799a );
 a3833a <=( a3741a ) or ( a3742a );
 a3834a <=( a3743a ) or ( a3833a );
 a3837a <=( a3739a ) or ( a3740a );
 a3840a <=( a3737a ) or ( a3738a );
 a3841a <=( a3840a ) or ( a3837a );
 a3842a <=( a3841a ) or ( a3834a );
 a3846a <=( a3734a ) or ( a3735a );
 a3847a <=( a3736a ) or ( a3846a );
 a3850a <=( a3732a ) or ( a3733a );
 a3853a <=( a3730a ) or ( a3731a );
 a3854a <=( a3853a ) or ( a3850a );
 a3855a <=( a3854a ) or ( a3847a );
 a3856a <=( a3855a ) or ( a3842a );
 a3860a <=( a3727a ) or ( a3728a );
 a3861a <=( a3729a ) or ( a3860a );
 a3864a <=( a3725a ) or ( a3726a );
 a3867a <=( a3723a ) or ( a3724a );
 a3868a <=( a3867a ) or ( a3864a );
 a3869a <=( a3868a ) or ( a3861a );
 a3872a <=( a3721a ) or ( a3722a );
 a3875a <=( a3719a ) or ( a3720a );
 a3876a <=( a3875a ) or ( a3872a );
 a3879a <=( a3717a ) or ( a3718a );
 a3882a <=( a3715a ) or ( a3716a );
 a3883a <=( a3882a ) or ( a3879a );
 a3884a <=( a3883a ) or ( a3876a );
 a3885a <=( a3884a ) or ( a3869a );
 a3886a <=( a3885a ) or ( a3856a );
 a3887a <=( a3886a ) or ( a3829a );
 a3891a <=( a3712a ) or ( a3713a );
 a3892a <=( a3714a ) or ( a3891a );
 a3895a <=( a3710a ) or ( a3711a );
 a3898a <=( a3708a ) or ( a3709a );
 a3899a <=( a3898a ) or ( a3895a );
 a3900a <=( a3899a ) or ( a3892a );
 a3904a <=( a3705a ) or ( a3706a );
 a3905a <=( a3707a ) or ( a3904a );
 a3908a <=( a3703a ) or ( a3704a );
 a3911a <=( a3701a ) or ( a3702a );
 a3912a <=( a3911a ) or ( a3908a );
 a3913a <=( a3912a ) or ( a3905a );
 a3914a <=( a3913a ) or ( a3900a );
 a3918a <=( a3698a ) or ( a3699a );
 a3919a <=( a3700a ) or ( a3918a );
 a3922a <=( a3696a ) or ( a3697a );
 a3925a <=( a3694a ) or ( a3695a );
 a3926a <=( a3925a ) or ( a3922a );
 a3927a <=( a3926a ) or ( a3919a );
 a3930a <=( a3692a ) or ( a3693a );
 a3933a <=( a3690a ) or ( a3691a );
 a3934a <=( a3933a ) or ( a3930a );
 a3937a <=( a3688a ) or ( a3689a );
 a3940a <=( a3686a ) or ( a3687a );
 a3941a <=( a3940a ) or ( a3937a );
 a3942a <=( a3941a ) or ( a3934a );
 a3943a <=( a3942a ) or ( a3927a );
 a3944a <=( a3943a ) or ( a3914a );
 a3948a <=( a3683a ) or ( a3684a );
 a3949a <=( a3685a ) or ( a3948a );
 a3952a <=( a3681a ) or ( a3682a );
 a3955a <=( a3679a ) or ( a3680a );
 a3956a <=( a3955a ) or ( a3952a );
 a3957a <=( a3956a ) or ( a3949a );
 a3960a <=( a3677a ) or ( a3678a );
 a3963a <=( a3675a ) or ( a3676a );
 a3964a <=( a3963a ) or ( a3960a );
 a3967a <=( a3673a ) or ( a3674a );
 a3970a <=( a3671a ) or ( a3672a );
 a3971a <=( a3970a ) or ( a3967a );
 a3972a <=( a3971a ) or ( a3964a );
 a3973a <=( a3972a ) or ( a3957a );
 a3977a <=( a3668a ) or ( a3669a );
 a3978a <=( a3670a ) or ( a3977a );
 a3981a <=( a3666a ) or ( a3667a );
 a3984a <=( a3664a ) or ( a3665a );
 a3985a <=( a3984a ) or ( a3981a );
 a3986a <=( a3985a ) or ( a3978a );
 a3989a <=( a3662a ) or ( a3663a );
 a3992a <=( a3660a ) or ( a3661a );
 a3993a <=( a3992a ) or ( a3989a );
 a3996a <=( a3658a ) or ( a3659a );
 a3999a <=( a3656a ) or ( a3657a );
 a4000a <=( a3999a ) or ( a3996a );
 a4001a <=( a4000a ) or ( a3993a );
 a4002a <=( a4001a ) or ( a3986a );
 a4003a <=( a4002a ) or ( a3973a );
 a4004a <=( a4003a ) or ( a3944a );
 a4005a <=( a4004a ) or ( a3887a );
 a4009a <=( a3653a ) or ( a3654a );
 a4010a <=( a3655a ) or ( a4009a );
 a4013a <=( a3651a ) or ( a3652a );
 a4016a <=( a3649a ) or ( a3650a );
 a4017a <=( a4016a ) or ( a4013a );
 a4018a <=( a4017a ) or ( a4010a );
 a4022a <=( a3646a ) or ( a3647a );
 a4023a <=( a3648a ) or ( a4022a );
 a4026a <=( a3644a ) or ( a3645a );
 a4029a <=( a3642a ) or ( a3643a );
 a4030a <=( a4029a ) or ( a4026a );
 a4031a <=( a4030a ) or ( a4023a );
 a4032a <=( a4031a ) or ( a4018a );
 a4036a <=( a3639a ) or ( a3640a );
 a4037a <=( a3641a ) or ( a4036a );
 a4040a <=( a3637a ) or ( a3638a );
 a4043a <=( a3635a ) or ( a3636a );
 a4044a <=( a4043a ) or ( a4040a );
 a4045a <=( a4044a ) or ( a4037a );
 a4048a <=( a3633a ) or ( a3634a );
 a4051a <=( a3631a ) or ( a3632a );
 a4052a <=( a4051a ) or ( a4048a );
 a4055a <=( a3629a ) or ( a3630a );
 a4058a <=( a3627a ) or ( a3628a );
 a4059a <=( a4058a ) or ( a4055a );
 a4060a <=( a4059a ) or ( a4052a );
 a4061a <=( a4060a ) or ( a4045a );
 a4062a <=( a4061a ) or ( a4032a );
 a4066a <=( a3624a ) or ( a3625a );
 a4067a <=( a3626a ) or ( a4066a );
 a4070a <=( a3622a ) or ( a3623a );
 a4073a <=( a3620a ) or ( a3621a );
 a4074a <=( a4073a ) or ( a4070a );
 a4075a <=( a4074a ) or ( a4067a );
 a4078a <=( a3618a ) or ( a3619a );
 a4081a <=( a3616a ) or ( a3617a );
 a4082a <=( a4081a ) or ( a4078a );
 a4085a <=( a3614a ) or ( a3615a );
 a4088a <=( a3612a ) or ( a3613a );
 a4089a <=( a4088a ) or ( a4085a );
 a4090a <=( a4089a ) or ( a4082a );
 a4091a <=( a4090a ) or ( a4075a );
 a4095a <=( a3609a ) or ( a3610a );
 a4096a <=( a3611a ) or ( a4095a );
 a4099a <=( a3607a ) or ( a3608a );
 a4102a <=( a3605a ) or ( a3606a );
 a4103a <=( a4102a ) or ( a4099a );
 a4104a <=( a4103a ) or ( a4096a );
 a4107a <=( a3603a ) or ( a3604a );
 a4110a <=( a3601a ) or ( a3602a );
 a4111a <=( a4110a ) or ( a4107a );
 a4114a <=( a3599a ) or ( a3600a );
 a4117a <=( a3597a ) or ( a3598a );
 a4118a <=( a4117a ) or ( a4114a );
 a4119a <=( a4118a ) or ( a4111a );
 a4120a <=( a4119a ) or ( a4104a );
 a4121a <=( a4120a ) or ( a4091a );
 a4122a <=( a4121a ) or ( a4062a );
 a4126a <=( a3594a ) or ( a3595a );
 a4127a <=( a3596a ) or ( a4126a );
 a4130a <=( a3592a ) or ( a3593a );
 a4133a <=( a3590a ) or ( a3591a );
 a4134a <=( a4133a ) or ( a4130a );
 a4135a <=( a4134a ) or ( a4127a );
 a4139a <=( a3587a ) or ( a3588a );
 a4140a <=( a3589a ) or ( a4139a );
 a4143a <=( a3585a ) or ( a3586a );
 a4146a <=( a3583a ) or ( a3584a );
 a4147a <=( a4146a ) or ( a4143a );
 a4148a <=( a4147a ) or ( a4140a );
 a4149a <=( a4148a ) or ( a4135a );
 a4153a <=( a3580a ) or ( a3581a );
 a4154a <=( a3582a ) or ( a4153a );
 a4157a <=( a3578a ) or ( a3579a );
 a4160a <=( a3576a ) or ( a3577a );
 a4161a <=( a4160a ) or ( a4157a );
 a4162a <=( a4161a ) or ( a4154a );
 a4165a <=( a3574a ) or ( a3575a );
 a4168a <=( a3572a ) or ( a3573a );
 a4169a <=( a4168a ) or ( a4165a );
 a4172a <=( a3570a ) or ( a3571a );
 a4175a <=( a3568a ) or ( a3569a );
 a4176a <=( a4175a ) or ( a4172a );
 a4177a <=( a4176a ) or ( a4169a );
 a4178a <=( a4177a ) or ( a4162a );
 a4179a <=( a4178a ) or ( a4149a );
 a4183a <=( a3565a ) or ( a3566a );
 a4184a <=( a3567a ) or ( a4183a );
 a4187a <=( a3563a ) or ( a3564a );
 a4190a <=( a3561a ) or ( a3562a );
 a4191a <=( a4190a ) or ( a4187a );
 a4192a <=( a4191a ) or ( a4184a );
 a4195a <=( a3559a ) or ( a3560a );
 a4198a <=( a3557a ) or ( a3558a );
 a4199a <=( a4198a ) or ( a4195a );
 a4202a <=( a3555a ) or ( a3556a );
 a4205a <=( a3553a ) or ( a3554a );
 a4206a <=( a4205a ) or ( a4202a );
 a4207a <=( a4206a ) or ( a4199a );
 a4208a <=( a4207a ) or ( a4192a );
 a4212a <=( a3550a ) or ( a3551a );
 a4213a <=( a3552a ) or ( a4212a );
 a4216a <=( a3548a ) or ( a3549a );
 a4219a <=( a3546a ) or ( a3547a );
 a4220a <=( a4219a ) or ( a4216a );
 a4221a <=( a4220a ) or ( a4213a );
 a4224a <=( a3544a ) or ( a3545a );
 a4227a <=( a3542a ) or ( a3543a );
 a4228a <=( a4227a ) or ( a4224a );
 a4231a <=( a3540a ) or ( a3541a );
 a4234a <=( a3538a ) or ( a3539a );
 a4235a <=( a4234a ) or ( a4231a );
 a4236a <=( a4235a ) or ( a4228a );
 a4237a <=( a4236a ) or ( a4221a );
 a4238a <=( a4237a ) or ( a4208a );
 a4239a <=( a4238a ) or ( a4179a );
 a4240a <=( a4239a ) or ( a4122a );
 a4241a <=( a4240a ) or ( a4005a );
 a4245a <=( a3535a ) or ( a3536a );
 a4246a <=( a3537a ) or ( a4245a );
 a4249a <=( a3533a ) or ( a3534a );
 a4252a <=( a3531a ) or ( a3532a );
 a4253a <=( a4252a ) or ( a4249a );
 a4254a <=( a4253a ) or ( a4246a );
 a4258a <=( a3528a ) or ( a3529a );
 a4259a <=( a3530a ) or ( a4258a );
 a4262a <=( a3526a ) or ( a3527a );
 a4265a <=( a3524a ) or ( a3525a );
 a4266a <=( a4265a ) or ( a4262a );
 a4267a <=( a4266a ) or ( a4259a );
 a4268a <=( a4267a ) or ( a4254a );
 a4272a <=( a3521a ) or ( a3522a );
 a4273a <=( a3523a ) or ( a4272a );
 a4276a <=( a3519a ) or ( a3520a );
 a4279a <=( a3517a ) or ( a3518a );
 a4280a <=( a4279a ) or ( a4276a );
 a4281a <=( a4280a ) or ( a4273a );
 a4284a <=( a3515a ) or ( a3516a );
 a4287a <=( a3513a ) or ( a3514a );
 a4288a <=( a4287a ) or ( a4284a );
 a4291a <=( a3511a ) or ( a3512a );
 a4294a <=( a3509a ) or ( a3510a );
 a4295a <=( a4294a ) or ( a4291a );
 a4296a <=( a4295a ) or ( a4288a );
 a4297a <=( a4296a ) or ( a4281a );
 a4298a <=( a4297a ) or ( a4268a );
 a4302a <=( a3506a ) or ( a3507a );
 a4303a <=( a3508a ) or ( a4302a );
 a4306a <=( a3504a ) or ( a3505a );
 a4309a <=( a3502a ) or ( a3503a );
 a4310a <=( a4309a ) or ( a4306a );
 a4311a <=( a4310a ) or ( a4303a );
 a4314a <=( a3500a ) or ( a3501a );
 a4317a <=( a3498a ) or ( a3499a );
 a4318a <=( a4317a ) or ( a4314a );
 a4321a <=( a3496a ) or ( a3497a );
 a4324a <=( a3494a ) or ( a3495a );
 a4325a <=( a4324a ) or ( a4321a );
 a4326a <=( a4325a ) or ( a4318a );
 a4327a <=( a4326a ) or ( a4311a );
 a4331a <=( a3491a ) or ( a3492a );
 a4332a <=( a3493a ) or ( a4331a );
 a4335a <=( a3489a ) or ( a3490a );
 a4338a <=( a3487a ) or ( a3488a );
 a4339a <=( a4338a ) or ( a4335a );
 a4340a <=( a4339a ) or ( a4332a );
 a4343a <=( a3485a ) or ( a3486a );
 a4346a <=( a3483a ) or ( a3484a );
 a4347a <=( a4346a ) or ( a4343a );
 a4350a <=( a3481a ) or ( a3482a );
 a4353a <=( a3479a ) or ( a3480a );
 a4354a <=( a4353a ) or ( a4350a );
 a4355a <=( a4354a ) or ( a4347a );
 a4356a <=( a4355a ) or ( a4340a );
 a4357a <=( a4356a ) or ( a4327a );
 a4358a <=( a4357a ) or ( a4298a );
 a4362a <=( a3476a ) or ( a3477a );
 a4363a <=( a3478a ) or ( a4362a );
 a4366a <=( a3474a ) or ( a3475a );
 a4369a <=( a3472a ) or ( a3473a );
 a4370a <=( a4369a ) or ( a4366a );
 a4371a <=( a4370a ) or ( a4363a );
 a4375a <=( a3469a ) or ( a3470a );
 a4376a <=( a3471a ) or ( a4375a );
 a4379a <=( a3467a ) or ( a3468a );
 a4382a <=( a3465a ) or ( a3466a );
 a4383a <=( a4382a ) or ( a4379a );
 a4384a <=( a4383a ) or ( a4376a );
 a4385a <=( a4384a ) or ( a4371a );
 a4389a <=( a3462a ) or ( a3463a );
 a4390a <=( a3464a ) or ( a4389a );
 a4393a <=( a3460a ) or ( a3461a );
 a4396a <=( a3458a ) or ( a3459a );
 a4397a <=( a4396a ) or ( a4393a );
 a4398a <=( a4397a ) or ( a4390a );
 a4401a <=( a3456a ) or ( a3457a );
 a4404a <=( a3454a ) or ( a3455a );
 a4405a <=( a4404a ) or ( a4401a );
 a4408a <=( a3452a ) or ( a3453a );
 a4411a <=( a3450a ) or ( a3451a );
 a4412a <=( a4411a ) or ( a4408a );
 a4413a <=( a4412a ) or ( a4405a );
 a4414a <=( a4413a ) or ( a4398a );
 a4415a <=( a4414a ) or ( a4385a );
 a4419a <=( a3447a ) or ( a3448a );
 a4420a <=( a3449a ) or ( a4419a );
 a4423a <=( a3445a ) or ( a3446a );
 a4426a <=( a3443a ) or ( a3444a );
 a4427a <=( a4426a ) or ( a4423a );
 a4428a <=( a4427a ) or ( a4420a );
 a4431a <=( a3441a ) or ( a3442a );
 a4434a <=( a3439a ) or ( a3440a );
 a4435a <=( a4434a ) or ( a4431a );
 a4438a <=( a3437a ) or ( a3438a );
 a4441a <=( a3435a ) or ( a3436a );
 a4442a <=( a4441a ) or ( a4438a );
 a4443a <=( a4442a ) or ( a4435a );
 a4444a <=( a4443a ) or ( a4428a );
 a4448a <=( a3432a ) or ( a3433a );
 a4449a <=( a3434a ) or ( a4448a );
 a4452a <=( a3430a ) or ( a3431a );
 a4455a <=( a3428a ) or ( a3429a );
 a4456a <=( a4455a ) or ( a4452a );
 a4457a <=( a4456a ) or ( a4449a );
 a4460a <=( a3426a ) or ( a3427a );
 a4463a <=( a3424a ) or ( a3425a );
 a4464a <=( a4463a ) or ( a4460a );
 a4467a <=( a3422a ) or ( a3423a );
 a4470a <=( a3420a ) or ( a3421a );
 a4471a <=( a4470a ) or ( a4467a );
 a4472a <=( a4471a ) or ( a4464a );
 a4473a <=( a4472a ) or ( a4457a );
 a4474a <=( a4473a ) or ( a4444a );
 a4475a <=( a4474a ) or ( a4415a );
 a4476a <=( a4475a ) or ( a4358a );
 a4480a <=( a3417a ) or ( a3418a );
 a4481a <=( a3419a ) or ( a4480a );
 a4484a <=( a3415a ) or ( a3416a );
 a4487a <=( a3413a ) or ( a3414a );
 a4488a <=( a4487a ) or ( a4484a );
 a4489a <=( a4488a ) or ( a4481a );
 a4493a <=( a3410a ) or ( a3411a );
 a4494a <=( a3412a ) or ( a4493a );
 a4497a <=( a3408a ) or ( a3409a );
 a4500a <=( a3406a ) or ( a3407a );
 a4501a <=( a4500a ) or ( a4497a );
 a4502a <=( a4501a ) or ( a4494a );
 a4503a <=( a4502a ) or ( a4489a );
 a4507a <=( a3403a ) or ( a3404a );
 a4508a <=( a3405a ) or ( a4507a );
 a4511a <=( a3401a ) or ( a3402a );
 a4514a <=( a3399a ) or ( a3400a );
 a4515a <=( a4514a ) or ( a4511a );
 a4516a <=( a4515a ) or ( a4508a );
 a4519a <=( a3397a ) or ( a3398a );
 a4522a <=( a3395a ) or ( a3396a );
 a4523a <=( a4522a ) or ( a4519a );
 a4526a <=( a3393a ) or ( a3394a );
 a4529a <=( a3391a ) or ( a3392a );
 a4530a <=( a4529a ) or ( a4526a );
 a4531a <=( a4530a ) or ( a4523a );
 a4532a <=( a4531a ) or ( a4516a );
 a4533a <=( a4532a ) or ( a4503a );
 a4537a <=( a3388a ) or ( a3389a );
 a4538a <=( a3390a ) or ( a4537a );
 a4541a <=( a3386a ) or ( a3387a );
 a4544a <=( a3384a ) or ( a3385a );
 a4545a <=( a4544a ) or ( a4541a );
 a4546a <=( a4545a ) or ( a4538a );
 a4549a <=( a3382a ) or ( a3383a );
 a4552a <=( a3380a ) or ( a3381a );
 a4553a <=( a4552a ) or ( a4549a );
 a4556a <=( a3378a ) or ( a3379a );
 a4559a <=( a3376a ) or ( a3377a );
 a4560a <=( a4559a ) or ( a4556a );
 a4561a <=( a4560a ) or ( a4553a );
 a4562a <=( a4561a ) or ( a4546a );
 a4566a <=( a3373a ) or ( a3374a );
 a4567a <=( a3375a ) or ( a4566a );
 a4570a <=( a3371a ) or ( a3372a );
 a4573a <=( a3369a ) or ( a3370a );
 a4574a <=( a4573a ) or ( a4570a );
 a4575a <=( a4574a ) or ( a4567a );
 a4578a <=( a3367a ) or ( a3368a );
 a4581a <=( a3365a ) or ( a3366a );
 a4582a <=( a4581a ) or ( a4578a );
 a4585a <=( a3363a ) or ( a3364a );
 a4588a <=( a3361a ) or ( a3362a );
 a4589a <=( a4588a ) or ( a4585a );
 a4590a <=( a4589a ) or ( a4582a );
 a4591a <=( a4590a ) or ( a4575a );
 a4592a <=( a4591a ) or ( a4562a );
 a4593a <=( a4592a ) or ( a4533a );
 a4597a <=( a3358a ) or ( a3359a );
 a4598a <=( a3360a ) or ( a4597a );
 a4601a <=( a3356a ) or ( a3357a );
 a4604a <=( a3354a ) or ( a3355a );
 a4605a <=( a4604a ) or ( a4601a );
 a4606a <=( a4605a ) or ( a4598a );
 a4610a <=( a3351a ) or ( a3352a );
 a4611a <=( a3353a ) or ( a4610a );
 a4614a <=( a3349a ) or ( a3350a );
 a4617a <=( a3347a ) or ( a3348a );
 a4618a <=( a4617a ) or ( a4614a );
 a4619a <=( a4618a ) or ( a4611a );
 a4620a <=( a4619a ) or ( a4606a );
 a4624a <=( a3344a ) or ( a3345a );
 a4625a <=( a3346a ) or ( a4624a );
 a4628a <=( a3342a ) or ( a3343a );
 a4631a <=( a3340a ) or ( a3341a );
 a4632a <=( a4631a ) or ( a4628a );
 a4633a <=( a4632a ) or ( a4625a );
 a4636a <=( a3338a ) or ( a3339a );
 a4639a <=( a3336a ) or ( a3337a );
 a4640a <=( a4639a ) or ( a4636a );
 a4643a <=( a3334a ) or ( a3335a );
 a4646a <=( a3332a ) or ( a3333a );
 a4647a <=( a4646a ) or ( a4643a );
 a4648a <=( a4647a ) or ( a4640a );
 a4649a <=( a4648a ) or ( a4633a );
 a4650a <=( a4649a ) or ( a4620a );
 a4654a <=( a3329a ) or ( a3330a );
 a4655a <=( a3331a ) or ( a4654a );
 a4658a <=( a3327a ) or ( a3328a );
 a4661a <=( a3325a ) or ( a3326a );
 a4662a <=( a4661a ) or ( a4658a );
 a4663a <=( a4662a ) or ( a4655a );
 a4666a <=( a3323a ) or ( a3324a );
 a4669a <=( a3321a ) or ( a3322a );
 a4670a <=( a4669a ) or ( a4666a );
 a4673a <=( a3319a ) or ( a3320a );
 a4676a <=( a3317a ) or ( a3318a );
 a4677a <=( a4676a ) or ( a4673a );
 a4678a <=( a4677a ) or ( a4670a );
 a4679a <=( a4678a ) or ( a4663a );
 a4683a <=( a3314a ) or ( a3315a );
 a4684a <=( a3316a ) or ( a4683a );
 a4687a <=( a3312a ) or ( a3313a );
 a4690a <=( a3310a ) or ( a3311a );
 a4691a <=( a4690a ) or ( a4687a );
 a4692a <=( a4691a ) or ( a4684a );
 a4695a <=( a3308a ) or ( a3309a );
 a4698a <=( a3306a ) or ( a3307a );
 a4699a <=( a4698a ) or ( a4695a );
 a4702a <=( a3304a ) or ( a3305a );
 a4705a <=( a3302a ) or ( a3303a );
 a4706a <=( a4705a ) or ( a4702a );
 a4707a <=( a4706a ) or ( a4699a );
 a4708a <=( a4707a ) or ( a4692a );
 a4709a <=( a4708a ) or ( a4679a );
 a4710a <=( a4709a ) or ( a4650a );
 a4711a <=( a4710a ) or ( a4593a );
 a4712a <=( a4711a ) or ( a4476a );
 a4713a <=( a4712a ) or ( a4241a );
 a4717a <=( a3299a ) or ( a3300a );
 a4718a <=( a3301a ) or ( a4717a );
 a4721a <=( a3297a ) or ( a3298a );
 a4724a <=( a3295a ) or ( a3296a );
 a4725a <=( a4724a ) or ( a4721a );
 a4726a <=( a4725a ) or ( a4718a );
 a4730a <=( a3292a ) or ( a3293a );
 a4731a <=( a3294a ) or ( a4730a );
 a4734a <=( a3290a ) or ( a3291a );
 a4737a <=( a3288a ) or ( a3289a );
 a4738a <=( a4737a ) or ( a4734a );
 a4739a <=( a4738a ) or ( a4731a );
 a4740a <=( a4739a ) or ( a4726a );
 a4744a <=( a3285a ) or ( a3286a );
 a4745a <=( a3287a ) or ( a4744a );
 a4748a <=( a3283a ) or ( a3284a );
 a4751a <=( a3281a ) or ( a3282a );
 a4752a <=( a4751a ) or ( a4748a );
 a4753a <=( a4752a ) or ( a4745a );
 a4756a <=( a3279a ) or ( a3280a );
 a4759a <=( a3277a ) or ( a3278a );
 a4760a <=( a4759a ) or ( a4756a );
 a4763a <=( a3275a ) or ( a3276a );
 a4766a <=( a3273a ) or ( a3274a );
 a4767a <=( a4766a ) or ( a4763a );
 a4768a <=( a4767a ) or ( a4760a );
 a4769a <=( a4768a ) or ( a4753a );
 a4770a <=( a4769a ) or ( a4740a );
 a4774a <=( a3270a ) or ( a3271a );
 a4775a <=( a3272a ) or ( a4774a );
 a4778a <=( a3268a ) or ( a3269a );
 a4781a <=( a3266a ) or ( a3267a );
 a4782a <=( a4781a ) or ( a4778a );
 a4783a <=( a4782a ) or ( a4775a );
 a4786a <=( a3264a ) or ( a3265a );
 a4789a <=( a3262a ) or ( a3263a );
 a4790a <=( a4789a ) or ( a4786a );
 a4793a <=( a3260a ) or ( a3261a );
 a4796a <=( a3258a ) or ( a3259a );
 a4797a <=( a4796a ) or ( a4793a );
 a4798a <=( a4797a ) or ( a4790a );
 a4799a <=( a4798a ) or ( a4783a );
 a4803a <=( a3255a ) or ( a3256a );
 a4804a <=( a3257a ) or ( a4803a );
 a4807a <=( a3253a ) or ( a3254a );
 a4810a <=( a3251a ) or ( a3252a );
 a4811a <=( a4810a ) or ( a4807a );
 a4812a <=( a4811a ) or ( a4804a );
 a4815a <=( a3249a ) or ( a3250a );
 a4818a <=( a3247a ) or ( a3248a );
 a4819a <=( a4818a ) or ( a4815a );
 a4822a <=( a3245a ) or ( a3246a );
 a4825a <=( a3243a ) or ( a3244a );
 a4826a <=( a4825a ) or ( a4822a );
 a4827a <=( a4826a ) or ( a4819a );
 a4828a <=( a4827a ) or ( a4812a );
 a4829a <=( a4828a ) or ( a4799a );
 a4830a <=( a4829a ) or ( a4770a );
 a4834a <=( a3240a ) or ( a3241a );
 a4835a <=( a3242a ) or ( a4834a );
 a4838a <=( a3238a ) or ( a3239a );
 a4841a <=( a3236a ) or ( a3237a );
 a4842a <=( a4841a ) or ( a4838a );
 a4843a <=( a4842a ) or ( a4835a );
 a4847a <=( a3233a ) or ( a3234a );
 a4848a <=( a3235a ) or ( a4847a );
 a4851a <=( a3231a ) or ( a3232a );
 a4854a <=( a3229a ) or ( a3230a );
 a4855a <=( a4854a ) or ( a4851a );
 a4856a <=( a4855a ) or ( a4848a );
 a4857a <=( a4856a ) or ( a4843a );
 a4861a <=( a3226a ) or ( a3227a );
 a4862a <=( a3228a ) or ( a4861a );
 a4865a <=( a3224a ) or ( a3225a );
 a4868a <=( a3222a ) or ( a3223a );
 a4869a <=( a4868a ) or ( a4865a );
 a4870a <=( a4869a ) or ( a4862a );
 a4873a <=( a3220a ) or ( a3221a );
 a4876a <=( a3218a ) or ( a3219a );
 a4877a <=( a4876a ) or ( a4873a );
 a4880a <=( a3216a ) or ( a3217a );
 a4883a <=( a3214a ) or ( a3215a );
 a4884a <=( a4883a ) or ( a4880a );
 a4885a <=( a4884a ) or ( a4877a );
 a4886a <=( a4885a ) or ( a4870a );
 a4887a <=( a4886a ) or ( a4857a );
 a4891a <=( a3211a ) or ( a3212a );
 a4892a <=( a3213a ) or ( a4891a );
 a4895a <=( a3209a ) or ( a3210a );
 a4898a <=( a3207a ) or ( a3208a );
 a4899a <=( a4898a ) or ( a4895a );
 a4900a <=( a4899a ) or ( a4892a );
 a4903a <=( a3205a ) or ( a3206a );
 a4906a <=( a3203a ) or ( a3204a );
 a4907a <=( a4906a ) or ( a4903a );
 a4910a <=( a3201a ) or ( a3202a );
 a4913a <=( a3199a ) or ( a3200a );
 a4914a <=( a4913a ) or ( a4910a );
 a4915a <=( a4914a ) or ( a4907a );
 a4916a <=( a4915a ) or ( a4900a );
 a4920a <=( a3196a ) or ( a3197a );
 a4921a <=( a3198a ) or ( a4920a );
 a4924a <=( a3194a ) or ( a3195a );
 a4927a <=( a3192a ) or ( a3193a );
 a4928a <=( a4927a ) or ( a4924a );
 a4929a <=( a4928a ) or ( a4921a );
 a4932a <=( a3190a ) or ( a3191a );
 a4935a <=( a3188a ) or ( a3189a );
 a4936a <=( a4935a ) or ( a4932a );
 a4939a <=( a3186a ) or ( a3187a );
 a4942a <=( a3184a ) or ( a3185a );
 a4943a <=( a4942a ) or ( a4939a );
 a4944a <=( a4943a ) or ( a4936a );
 a4945a <=( a4944a ) or ( a4929a );
 a4946a <=( a4945a ) or ( a4916a );
 a4947a <=( a4946a ) or ( a4887a );
 a4948a <=( a4947a ) or ( a4830a );
 a4952a <=( a3181a ) or ( a3182a );
 a4953a <=( a3183a ) or ( a4952a );
 a4956a <=( a3179a ) or ( a3180a );
 a4959a <=( a3177a ) or ( a3178a );
 a4960a <=( a4959a ) or ( a4956a );
 a4961a <=( a4960a ) or ( a4953a );
 a4965a <=( a3174a ) or ( a3175a );
 a4966a <=( a3176a ) or ( a4965a );
 a4969a <=( a3172a ) or ( a3173a );
 a4972a <=( a3170a ) or ( a3171a );
 a4973a <=( a4972a ) or ( a4969a );
 a4974a <=( a4973a ) or ( a4966a );
 a4975a <=( a4974a ) or ( a4961a );
 a4979a <=( a3167a ) or ( a3168a );
 a4980a <=( a3169a ) or ( a4979a );
 a4983a <=( a3165a ) or ( a3166a );
 a4986a <=( a3163a ) or ( a3164a );
 a4987a <=( a4986a ) or ( a4983a );
 a4988a <=( a4987a ) or ( a4980a );
 a4991a <=( a3161a ) or ( a3162a );
 a4994a <=( a3159a ) or ( a3160a );
 a4995a <=( a4994a ) or ( a4991a );
 a4998a <=( a3157a ) or ( a3158a );
 a5001a <=( a3155a ) or ( a3156a );
 a5002a <=( a5001a ) or ( a4998a );
 a5003a <=( a5002a ) or ( a4995a );
 a5004a <=( a5003a ) or ( a4988a );
 a5005a <=( a5004a ) or ( a4975a );
 a5009a <=( a3152a ) or ( a3153a );
 a5010a <=( a3154a ) or ( a5009a );
 a5013a <=( a3150a ) or ( a3151a );
 a5016a <=( a3148a ) or ( a3149a );
 a5017a <=( a5016a ) or ( a5013a );
 a5018a <=( a5017a ) or ( a5010a );
 a5021a <=( a3146a ) or ( a3147a );
 a5024a <=( a3144a ) or ( a3145a );
 a5025a <=( a5024a ) or ( a5021a );
 a5028a <=( a3142a ) or ( a3143a );
 a5031a <=( a3140a ) or ( a3141a );
 a5032a <=( a5031a ) or ( a5028a );
 a5033a <=( a5032a ) or ( a5025a );
 a5034a <=( a5033a ) or ( a5018a );
 a5038a <=( a3137a ) or ( a3138a );
 a5039a <=( a3139a ) or ( a5038a );
 a5042a <=( a3135a ) or ( a3136a );
 a5045a <=( a3133a ) or ( a3134a );
 a5046a <=( a5045a ) or ( a5042a );
 a5047a <=( a5046a ) or ( a5039a );
 a5050a <=( a3131a ) or ( a3132a );
 a5053a <=( a3129a ) or ( a3130a );
 a5054a <=( a5053a ) or ( a5050a );
 a5057a <=( a3127a ) or ( a3128a );
 a5060a <=( a3125a ) or ( a3126a );
 a5061a <=( a5060a ) or ( a5057a );
 a5062a <=( a5061a ) or ( a5054a );
 a5063a <=( a5062a ) or ( a5047a );
 a5064a <=( a5063a ) or ( a5034a );
 a5065a <=( a5064a ) or ( a5005a );
 a5069a <=( a3122a ) or ( a3123a );
 a5070a <=( a3124a ) or ( a5069a );
 a5073a <=( a3120a ) or ( a3121a );
 a5076a <=( a3118a ) or ( a3119a );
 a5077a <=( a5076a ) or ( a5073a );
 a5078a <=( a5077a ) or ( a5070a );
 a5082a <=( a3115a ) or ( a3116a );
 a5083a <=( a3117a ) or ( a5082a );
 a5086a <=( a3113a ) or ( a3114a );
 a5089a <=( a3111a ) or ( a3112a );
 a5090a <=( a5089a ) or ( a5086a );
 a5091a <=( a5090a ) or ( a5083a );
 a5092a <=( a5091a ) or ( a5078a );
 a5096a <=( a3108a ) or ( a3109a );
 a5097a <=( a3110a ) or ( a5096a );
 a5100a <=( a3106a ) or ( a3107a );
 a5103a <=( a3104a ) or ( a3105a );
 a5104a <=( a5103a ) or ( a5100a );
 a5105a <=( a5104a ) or ( a5097a );
 a5108a <=( a3102a ) or ( a3103a );
 a5111a <=( a3100a ) or ( a3101a );
 a5112a <=( a5111a ) or ( a5108a );
 a5115a <=( a3098a ) or ( a3099a );
 a5118a <=( a3096a ) or ( a3097a );
 a5119a <=( a5118a ) or ( a5115a );
 a5120a <=( a5119a ) or ( a5112a );
 a5121a <=( a5120a ) or ( a5105a );
 a5122a <=( a5121a ) or ( a5092a );
 a5126a <=( a3093a ) or ( a3094a );
 a5127a <=( a3095a ) or ( a5126a );
 a5130a <=( a3091a ) or ( a3092a );
 a5133a <=( a3089a ) or ( a3090a );
 a5134a <=( a5133a ) or ( a5130a );
 a5135a <=( a5134a ) or ( a5127a );
 a5138a <=( a3087a ) or ( a3088a );
 a5141a <=( a3085a ) or ( a3086a );
 a5142a <=( a5141a ) or ( a5138a );
 a5145a <=( a3083a ) or ( a3084a );
 a5148a <=( a3081a ) or ( a3082a );
 a5149a <=( a5148a ) or ( a5145a );
 a5150a <=( a5149a ) or ( a5142a );
 a5151a <=( a5150a ) or ( a5135a );
 a5155a <=( a3078a ) or ( a3079a );
 a5156a <=( a3080a ) or ( a5155a );
 a5159a <=( a3076a ) or ( a3077a );
 a5162a <=( a3074a ) or ( a3075a );
 a5163a <=( a5162a ) or ( a5159a );
 a5164a <=( a5163a ) or ( a5156a );
 a5167a <=( a3072a ) or ( a3073a );
 a5170a <=( a3070a ) or ( a3071a );
 a5171a <=( a5170a ) or ( a5167a );
 a5174a <=( a3068a ) or ( a3069a );
 a5177a <=( a3066a ) or ( a3067a );
 a5178a <=( a5177a ) or ( a5174a );
 a5179a <=( a5178a ) or ( a5171a );
 a5180a <=( a5179a ) or ( a5164a );
 a5181a <=( a5180a ) or ( a5151a );
 a5182a <=( a5181a ) or ( a5122a );
 a5183a <=( a5182a ) or ( a5065a );
 a5184a <=( a5183a ) or ( a4948a );
 a5188a <=( a3063a ) or ( a3064a );
 a5189a <=( a3065a ) or ( a5188a );
 a5192a <=( a3061a ) or ( a3062a );
 a5195a <=( a3059a ) or ( a3060a );
 a5196a <=( a5195a ) or ( a5192a );
 a5197a <=( a5196a ) or ( a5189a );
 a5201a <=( a3056a ) or ( a3057a );
 a5202a <=( a3058a ) or ( a5201a );
 a5205a <=( a3054a ) or ( a3055a );
 a5208a <=( a3052a ) or ( a3053a );
 a5209a <=( a5208a ) or ( a5205a );
 a5210a <=( a5209a ) or ( a5202a );
 a5211a <=( a5210a ) or ( a5197a );
 a5215a <=( a3049a ) or ( a3050a );
 a5216a <=( a3051a ) or ( a5215a );
 a5219a <=( a3047a ) or ( a3048a );
 a5222a <=( a3045a ) or ( a3046a );
 a5223a <=( a5222a ) or ( a5219a );
 a5224a <=( a5223a ) or ( a5216a );
 a5227a <=( a3043a ) or ( a3044a );
 a5230a <=( a3041a ) or ( a3042a );
 a5231a <=( a5230a ) or ( a5227a );
 a5234a <=( a3039a ) or ( a3040a );
 a5237a <=( a3037a ) or ( a3038a );
 a5238a <=( a5237a ) or ( a5234a );
 a5239a <=( a5238a ) or ( a5231a );
 a5240a <=( a5239a ) or ( a5224a );
 a5241a <=( a5240a ) or ( a5211a );
 a5245a <=( a3034a ) or ( a3035a );
 a5246a <=( a3036a ) or ( a5245a );
 a5249a <=( a3032a ) or ( a3033a );
 a5252a <=( a3030a ) or ( a3031a );
 a5253a <=( a5252a ) or ( a5249a );
 a5254a <=( a5253a ) or ( a5246a );
 a5257a <=( a3028a ) or ( a3029a );
 a5260a <=( a3026a ) or ( a3027a );
 a5261a <=( a5260a ) or ( a5257a );
 a5264a <=( a3024a ) or ( a3025a );
 a5267a <=( a3022a ) or ( a3023a );
 a5268a <=( a5267a ) or ( a5264a );
 a5269a <=( a5268a ) or ( a5261a );
 a5270a <=( a5269a ) or ( a5254a );
 a5274a <=( a3019a ) or ( a3020a );
 a5275a <=( a3021a ) or ( a5274a );
 a5278a <=( a3017a ) or ( a3018a );
 a5281a <=( a3015a ) or ( a3016a );
 a5282a <=( a5281a ) or ( a5278a );
 a5283a <=( a5282a ) or ( a5275a );
 a5286a <=( a3013a ) or ( a3014a );
 a5289a <=( a3011a ) or ( a3012a );
 a5290a <=( a5289a ) or ( a5286a );
 a5293a <=( a3009a ) or ( a3010a );
 a5296a <=( a3007a ) or ( a3008a );
 a5297a <=( a5296a ) or ( a5293a );
 a5298a <=( a5297a ) or ( a5290a );
 a5299a <=( a5298a ) or ( a5283a );
 a5300a <=( a5299a ) or ( a5270a );
 a5301a <=( a5300a ) or ( a5241a );
 a5305a <=( a3004a ) or ( a3005a );
 a5306a <=( a3006a ) or ( a5305a );
 a5309a <=( a3002a ) or ( a3003a );
 a5312a <=( a3000a ) or ( a3001a );
 a5313a <=( a5312a ) or ( a5309a );
 a5314a <=( a5313a ) or ( a5306a );
 a5318a <=( a2997a ) or ( a2998a );
 a5319a <=( a2999a ) or ( a5318a );
 a5322a <=( a2995a ) or ( a2996a );
 a5325a <=( a2993a ) or ( a2994a );
 a5326a <=( a5325a ) or ( a5322a );
 a5327a <=( a5326a ) or ( a5319a );
 a5328a <=( a5327a ) or ( a5314a );
 a5332a <=( a2990a ) or ( a2991a );
 a5333a <=( a2992a ) or ( a5332a );
 a5336a <=( a2988a ) or ( a2989a );
 a5339a <=( a2986a ) or ( a2987a );
 a5340a <=( a5339a ) or ( a5336a );
 a5341a <=( a5340a ) or ( a5333a );
 a5344a <=( a2984a ) or ( a2985a );
 a5347a <=( a2982a ) or ( a2983a );
 a5348a <=( a5347a ) or ( a5344a );
 a5351a <=( a2980a ) or ( a2981a );
 a5354a <=( a2978a ) or ( a2979a );
 a5355a <=( a5354a ) or ( a5351a );
 a5356a <=( a5355a ) or ( a5348a );
 a5357a <=( a5356a ) or ( a5341a );
 a5358a <=( a5357a ) or ( a5328a );
 a5362a <=( a2975a ) or ( a2976a );
 a5363a <=( a2977a ) or ( a5362a );
 a5366a <=( a2973a ) or ( a2974a );
 a5369a <=( a2971a ) or ( a2972a );
 a5370a <=( a5369a ) or ( a5366a );
 a5371a <=( a5370a ) or ( a5363a );
 a5374a <=( a2969a ) or ( a2970a );
 a5377a <=( a2967a ) or ( a2968a );
 a5378a <=( a5377a ) or ( a5374a );
 a5381a <=( a2965a ) or ( a2966a );
 a5384a <=( a2963a ) or ( a2964a );
 a5385a <=( a5384a ) or ( a5381a );
 a5386a <=( a5385a ) or ( a5378a );
 a5387a <=( a5386a ) or ( a5371a );
 a5391a <=( a2960a ) or ( a2961a );
 a5392a <=( a2962a ) or ( a5391a );
 a5395a <=( a2958a ) or ( a2959a );
 a5398a <=( a2956a ) or ( a2957a );
 a5399a <=( a5398a ) or ( a5395a );
 a5400a <=( a5399a ) or ( a5392a );
 a5403a <=( a2954a ) or ( a2955a );
 a5406a <=( a2952a ) or ( a2953a );
 a5407a <=( a5406a ) or ( a5403a );
 a5410a <=( a2950a ) or ( a2951a );
 a5413a <=( a2948a ) or ( a2949a );
 a5414a <=( a5413a ) or ( a5410a );
 a5415a <=( a5414a ) or ( a5407a );
 a5416a <=( a5415a ) or ( a5400a );
 a5417a <=( a5416a ) or ( a5387a );
 a5418a <=( a5417a ) or ( a5358a );
 a5419a <=( a5418a ) or ( a5301a );
 a5423a <=( a2945a ) or ( a2946a );
 a5424a <=( a2947a ) or ( a5423a );
 a5427a <=( a2943a ) or ( a2944a );
 a5430a <=( a2941a ) or ( a2942a );
 a5431a <=( a5430a ) or ( a5427a );
 a5432a <=( a5431a ) or ( a5424a );
 a5436a <=( a2938a ) or ( a2939a );
 a5437a <=( a2940a ) or ( a5436a );
 a5440a <=( a2936a ) or ( a2937a );
 a5443a <=( a2934a ) or ( a2935a );
 a5444a <=( a5443a ) or ( a5440a );
 a5445a <=( a5444a ) or ( a5437a );
 a5446a <=( a5445a ) or ( a5432a );
 a5450a <=( a2931a ) or ( a2932a );
 a5451a <=( a2933a ) or ( a5450a );
 a5454a <=( a2929a ) or ( a2930a );
 a5457a <=( a2927a ) or ( a2928a );
 a5458a <=( a5457a ) or ( a5454a );
 a5459a <=( a5458a ) or ( a5451a );
 a5462a <=( a2925a ) or ( a2926a );
 a5465a <=( a2923a ) or ( a2924a );
 a5466a <=( a5465a ) or ( a5462a );
 a5469a <=( a2921a ) or ( a2922a );
 a5472a <=( a2919a ) or ( a2920a );
 a5473a <=( a5472a ) or ( a5469a );
 a5474a <=( a5473a ) or ( a5466a );
 a5475a <=( a5474a ) or ( a5459a );
 a5476a <=( a5475a ) or ( a5446a );
 a5480a <=( a2916a ) or ( a2917a );
 a5481a <=( a2918a ) or ( a5480a );
 a5484a <=( a2914a ) or ( a2915a );
 a5487a <=( a2912a ) or ( a2913a );
 a5488a <=( a5487a ) or ( a5484a );
 a5489a <=( a5488a ) or ( a5481a );
 a5492a <=( a2910a ) or ( a2911a );
 a5495a <=( a2908a ) or ( a2909a );
 a5496a <=( a5495a ) or ( a5492a );
 a5499a <=( a2906a ) or ( a2907a );
 a5502a <=( a2904a ) or ( a2905a );
 a5503a <=( a5502a ) or ( a5499a );
 a5504a <=( a5503a ) or ( a5496a );
 a5505a <=( a5504a ) or ( a5489a );
 a5509a <=( a2901a ) or ( a2902a );
 a5510a <=( a2903a ) or ( a5509a );
 a5513a <=( a2899a ) or ( a2900a );
 a5516a <=( a2897a ) or ( a2898a );
 a5517a <=( a5516a ) or ( a5513a );
 a5518a <=( a5517a ) or ( a5510a );
 a5521a <=( a2895a ) or ( a2896a );
 a5524a <=( a2893a ) or ( a2894a );
 a5525a <=( a5524a ) or ( a5521a );
 a5528a <=( a2891a ) or ( a2892a );
 a5531a <=( a2889a ) or ( a2890a );
 a5532a <=( a5531a ) or ( a5528a );
 a5533a <=( a5532a ) or ( a5525a );
 a5534a <=( a5533a ) or ( a5518a );
 a5535a <=( a5534a ) or ( a5505a );
 a5536a <=( a5535a ) or ( a5476a );
 a5540a <=( a2886a ) or ( a2887a );
 a5541a <=( a2888a ) or ( a5540a );
 a5544a <=( a2884a ) or ( a2885a );
 a5547a <=( a2882a ) or ( a2883a );
 a5548a <=( a5547a ) or ( a5544a );
 a5549a <=( a5548a ) or ( a5541a );
 a5553a <=( a2879a ) or ( a2880a );
 a5554a <=( a2881a ) or ( a5553a );
 a5557a <=( a2877a ) or ( a2878a );
 a5560a <=( a2875a ) or ( a2876a );
 a5561a <=( a5560a ) or ( a5557a );
 a5562a <=( a5561a ) or ( a5554a );
 a5563a <=( a5562a ) or ( a5549a );
 a5567a <=( a2872a ) or ( a2873a );
 a5568a <=( a2874a ) or ( a5567a );
 a5571a <=( a2870a ) or ( a2871a );
 a5574a <=( a2868a ) or ( a2869a );
 a5575a <=( a5574a ) or ( a5571a );
 a5576a <=( a5575a ) or ( a5568a );
 a5579a <=( a2866a ) or ( a2867a );
 a5582a <=( a2864a ) or ( a2865a );
 a5583a <=( a5582a ) or ( a5579a );
 a5586a <=( a2862a ) or ( a2863a );
 a5589a <=( a2860a ) or ( a2861a );
 a5590a <=( a5589a ) or ( a5586a );
 a5591a <=( a5590a ) or ( a5583a );
 a5592a <=( a5591a ) or ( a5576a );
 a5593a <=( a5592a ) or ( a5563a );
 a5597a <=( a2857a ) or ( a2858a );
 a5598a <=( a2859a ) or ( a5597a );
 a5601a <=( a2855a ) or ( a2856a );
 a5604a <=( a2853a ) or ( a2854a );
 a5605a <=( a5604a ) or ( a5601a );
 a5606a <=( a5605a ) or ( a5598a );
 a5609a <=( a2851a ) or ( a2852a );
 a5612a <=( a2849a ) or ( a2850a );
 a5613a <=( a5612a ) or ( a5609a );
 a5616a <=( a2847a ) or ( a2848a );
 a5619a <=( a2845a ) or ( a2846a );
 a5620a <=( a5619a ) or ( a5616a );
 a5621a <=( a5620a ) or ( a5613a );
 a5622a <=( a5621a ) or ( a5606a );
 a5626a <=( a2842a ) or ( a2843a );
 a5627a <=( a2844a ) or ( a5626a );
 a5630a <=( a2840a ) or ( a2841a );
 a5633a <=( a2838a ) or ( a2839a );
 a5634a <=( a5633a ) or ( a5630a );
 a5635a <=( a5634a ) or ( a5627a );
 a5638a <=( a2836a ) or ( a2837a );
 a5641a <=( a2834a ) or ( a2835a );
 a5642a <=( a5641a ) or ( a5638a );
 a5645a <=( a2832a ) or ( a2833a );
 a5648a <=( a2830a ) or ( a2831a );
 a5649a <=( a5648a ) or ( a5645a );
 a5650a <=( a5649a ) or ( a5642a );
 a5651a <=( a5650a ) or ( a5635a );
 a5652a <=( a5651a ) or ( a5622a );
 a5653a <=( a5652a ) or ( a5593a );
 a5654a <=( a5653a ) or ( a5536a );
 a5655a <=( a5654a ) or ( a5419a );
 a5656a <=( a5655a ) or ( a5184a );
 a5657a <=( a5656a ) or ( a4713a );
 a5661a <=( a2827a ) or ( a2828a );
 a5662a <=( a2829a ) or ( a5661a );
 a5665a <=( a2825a ) or ( a2826a );
 a5668a <=( a2823a ) or ( a2824a );
 a5669a <=( a5668a ) or ( a5665a );
 a5670a <=( a5669a ) or ( a5662a );
 a5674a <=( a2820a ) or ( a2821a );
 a5675a <=( a2822a ) or ( a5674a );
 a5678a <=( a2818a ) or ( a2819a );
 a5681a <=( a2816a ) or ( a2817a );
 a5682a <=( a5681a ) or ( a5678a );
 a5683a <=( a5682a ) or ( a5675a );
 a5684a <=( a5683a ) or ( a5670a );
 a5688a <=( a2813a ) or ( a2814a );
 a5689a <=( a2815a ) or ( a5688a );
 a5692a <=( a2811a ) or ( a2812a );
 a5695a <=( a2809a ) or ( a2810a );
 a5696a <=( a5695a ) or ( a5692a );
 a5697a <=( a5696a ) or ( a5689a );
 a5700a <=( a2807a ) or ( a2808a );
 a5703a <=( a2805a ) or ( a2806a );
 a5704a <=( a5703a ) or ( a5700a );
 a5707a <=( a2803a ) or ( a2804a );
 a5710a <=( a2801a ) or ( a2802a );
 a5711a <=( a5710a ) or ( a5707a );
 a5712a <=( a5711a ) or ( a5704a );
 a5713a <=( a5712a ) or ( a5697a );
 a5714a <=( a5713a ) or ( a5684a );
 a5718a <=( a2798a ) or ( a2799a );
 a5719a <=( a2800a ) or ( a5718a );
 a5722a <=( a2796a ) or ( a2797a );
 a5725a <=( a2794a ) or ( a2795a );
 a5726a <=( a5725a ) or ( a5722a );
 a5727a <=( a5726a ) or ( a5719a );
 a5731a <=( a2791a ) or ( a2792a );
 a5732a <=( a2793a ) or ( a5731a );
 a5735a <=( a2789a ) or ( a2790a );
 a5738a <=( a2787a ) or ( a2788a );
 a5739a <=( a5738a ) or ( a5735a );
 a5740a <=( a5739a ) or ( a5732a );
 a5741a <=( a5740a ) or ( a5727a );
 a5745a <=( a2784a ) or ( a2785a );
 a5746a <=( a2786a ) or ( a5745a );
 a5749a <=( a2782a ) or ( a2783a );
 a5752a <=( a2780a ) or ( a2781a );
 a5753a <=( a5752a ) or ( a5749a );
 a5754a <=( a5753a ) or ( a5746a );
 a5757a <=( a2778a ) or ( a2779a );
 a5760a <=( a2776a ) or ( a2777a );
 a5761a <=( a5760a ) or ( a5757a );
 a5764a <=( a2774a ) or ( a2775a );
 a5767a <=( a2772a ) or ( a2773a );
 a5768a <=( a5767a ) or ( a5764a );
 a5769a <=( a5768a ) or ( a5761a );
 a5770a <=( a5769a ) or ( a5754a );
 a5771a <=( a5770a ) or ( a5741a );
 a5772a <=( a5771a ) or ( a5714a );
 a5776a <=( a2769a ) or ( a2770a );
 a5777a <=( a2771a ) or ( a5776a );
 a5780a <=( a2767a ) or ( a2768a );
 a5783a <=( a2765a ) or ( a2766a );
 a5784a <=( a5783a ) or ( a5780a );
 a5785a <=( a5784a ) or ( a5777a );
 a5789a <=( a2762a ) or ( a2763a );
 a5790a <=( a2764a ) or ( a5789a );
 a5793a <=( a2760a ) or ( a2761a );
 a5796a <=( a2758a ) or ( a2759a );
 a5797a <=( a5796a ) or ( a5793a );
 a5798a <=( a5797a ) or ( a5790a );
 a5799a <=( a5798a ) or ( a5785a );
 a5803a <=( a2755a ) or ( a2756a );
 a5804a <=( a2757a ) or ( a5803a );
 a5807a <=( a2753a ) or ( a2754a );
 a5810a <=( a2751a ) or ( a2752a );
 a5811a <=( a5810a ) or ( a5807a );
 a5812a <=( a5811a ) or ( a5804a );
 a5815a <=( a2749a ) or ( a2750a );
 a5818a <=( a2747a ) or ( a2748a );
 a5819a <=( a5818a ) or ( a5815a );
 a5822a <=( a2745a ) or ( a2746a );
 a5825a <=( a2743a ) or ( a2744a );
 a5826a <=( a5825a ) or ( a5822a );
 a5827a <=( a5826a ) or ( a5819a );
 a5828a <=( a5827a ) or ( a5812a );
 a5829a <=( a5828a ) or ( a5799a );
 a5833a <=( a2740a ) or ( a2741a );
 a5834a <=( a2742a ) or ( a5833a );
 a5837a <=( a2738a ) or ( a2739a );
 a5840a <=( a2736a ) or ( a2737a );
 a5841a <=( a5840a ) or ( a5837a );
 a5842a <=( a5841a ) or ( a5834a );
 a5845a <=( a2734a ) or ( a2735a );
 a5848a <=( a2732a ) or ( a2733a );
 a5849a <=( a5848a ) or ( a5845a );
 a5852a <=( a2730a ) or ( a2731a );
 a5855a <=( a2728a ) or ( a2729a );
 a5856a <=( a5855a ) or ( a5852a );
 a5857a <=( a5856a ) or ( a5849a );
 a5858a <=( a5857a ) or ( a5842a );
 a5862a <=( a2725a ) or ( a2726a );
 a5863a <=( a2727a ) or ( a5862a );
 a5866a <=( a2723a ) or ( a2724a );
 a5869a <=( a2721a ) or ( a2722a );
 a5870a <=( a5869a ) or ( a5866a );
 a5871a <=( a5870a ) or ( a5863a );
 a5874a <=( a2719a ) or ( a2720a );
 a5877a <=( a2717a ) or ( a2718a );
 a5878a <=( a5877a ) or ( a5874a );
 a5881a <=( a2715a ) or ( a2716a );
 a5884a <=( a2713a ) or ( a2714a );
 a5885a <=( a5884a ) or ( a5881a );
 a5886a <=( a5885a ) or ( a5878a );
 a5887a <=( a5886a ) or ( a5871a );
 a5888a <=( a5887a ) or ( a5858a );
 a5889a <=( a5888a ) or ( a5829a );
 a5890a <=( a5889a ) or ( a5772a );
 a5894a <=( a2710a ) or ( a2711a );
 a5895a <=( a2712a ) or ( a5894a );
 a5898a <=( a2708a ) or ( a2709a );
 a5901a <=( a2706a ) or ( a2707a );
 a5902a <=( a5901a ) or ( a5898a );
 a5903a <=( a5902a ) or ( a5895a );
 a5907a <=( a2703a ) or ( a2704a );
 a5908a <=( a2705a ) or ( a5907a );
 a5911a <=( a2701a ) or ( a2702a );
 a5914a <=( a2699a ) or ( a2700a );
 a5915a <=( a5914a ) or ( a5911a );
 a5916a <=( a5915a ) or ( a5908a );
 a5917a <=( a5916a ) or ( a5903a );
 a5921a <=( a2696a ) or ( a2697a );
 a5922a <=( a2698a ) or ( a5921a );
 a5925a <=( a2694a ) or ( a2695a );
 a5928a <=( a2692a ) or ( a2693a );
 a5929a <=( a5928a ) or ( a5925a );
 a5930a <=( a5929a ) or ( a5922a );
 a5933a <=( a2690a ) or ( a2691a );
 a5936a <=( a2688a ) or ( a2689a );
 a5937a <=( a5936a ) or ( a5933a );
 a5940a <=( a2686a ) or ( a2687a );
 a5943a <=( a2684a ) or ( a2685a );
 a5944a <=( a5943a ) or ( a5940a );
 a5945a <=( a5944a ) or ( a5937a );
 a5946a <=( a5945a ) or ( a5930a );
 a5947a <=( a5946a ) or ( a5917a );
 a5951a <=( a2681a ) or ( a2682a );
 a5952a <=( a2683a ) or ( a5951a );
 a5955a <=( a2679a ) or ( a2680a );
 a5958a <=( a2677a ) or ( a2678a );
 a5959a <=( a5958a ) or ( a5955a );
 a5960a <=( a5959a ) or ( a5952a );
 a5963a <=( a2675a ) or ( a2676a );
 a5966a <=( a2673a ) or ( a2674a );
 a5967a <=( a5966a ) or ( a5963a );
 a5970a <=( a2671a ) or ( a2672a );
 a5973a <=( a2669a ) or ( a2670a );
 a5974a <=( a5973a ) or ( a5970a );
 a5975a <=( a5974a ) or ( a5967a );
 a5976a <=( a5975a ) or ( a5960a );
 a5980a <=( a2666a ) or ( a2667a );
 a5981a <=( a2668a ) or ( a5980a );
 a5984a <=( a2664a ) or ( a2665a );
 a5987a <=( a2662a ) or ( a2663a );
 a5988a <=( a5987a ) or ( a5984a );
 a5989a <=( a5988a ) or ( a5981a );
 a5992a <=( a2660a ) or ( a2661a );
 a5995a <=( a2658a ) or ( a2659a );
 a5996a <=( a5995a ) or ( a5992a );
 a5999a <=( a2656a ) or ( a2657a );
 a6002a <=( a2654a ) or ( a2655a );
 a6003a <=( a6002a ) or ( a5999a );
 a6004a <=( a6003a ) or ( a5996a );
 a6005a <=( a6004a ) or ( a5989a );
 a6006a <=( a6005a ) or ( a5976a );
 a6007a <=( a6006a ) or ( a5947a );
 a6011a <=( a2651a ) or ( a2652a );
 a6012a <=( a2653a ) or ( a6011a );
 a6015a <=( a2649a ) or ( a2650a );
 a6018a <=( a2647a ) or ( a2648a );
 a6019a <=( a6018a ) or ( a6015a );
 a6020a <=( a6019a ) or ( a6012a );
 a6024a <=( a2644a ) or ( a2645a );
 a6025a <=( a2646a ) or ( a6024a );
 a6028a <=( a2642a ) or ( a2643a );
 a6031a <=( a2640a ) or ( a2641a );
 a6032a <=( a6031a ) or ( a6028a );
 a6033a <=( a6032a ) or ( a6025a );
 a6034a <=( a6033a ) or ( a6020a );
 a6038a <=( a2637a ) or ( a2638a );
 a6039a <=( a2639a ) or ( a6038a );
 a6042a <=( a2635a ) or ( a2636a );
 a6045a <=( a2633a ) or ( a2634a );
 a6046a <=( a6045a ) or ( a6042a );
 a6047a <=( a6046a ) or ( a6039a );
 a6050a <=( a2631a ) or ( a2632a );
 a6053a <=( a2629a ) or ( a2630a );
 a6054a <=( a6053a ) or ( a6050a );
 a6057a <=( a2627a ) or ( a2628a );
 a6060a <=( a2625a ) or ( a2626a );
 a6061a <=( a6060a ) or ( a6057a );
 a6062a <=( a6061a ) or ( a6054a );
 a6063a <=( a6062a ) or ( a6047a );
 a6064a <=( a6063a ) or ( a6034a );
 a6068a <=( a2622a ) or ( a2623a );
 a6069a <=( a2624a ) or ( a6068a );
 a6072a <=( a2620a ) or ( a2621a );
 a6075a <=( a2618a ) or ( a2619a );
 a6076a <=( a6075a ) or ( a6072a );
 a6077a <=( a6076a ) or ( a6069a );
 a6080a <=( a2616a ) or ( a2617a );
 a6083a <=( a2614a ) or ( a2615a );
 a6084a <=( a6083a ) or ( a6080a );
 a6087a <=( a2612a ) or ( a2613a );
 a6090a <=( a2610a ) or ( a2611a );
 a6091a <=( a6090a ) or ( a6087a );
 a6092a <=( a6091a ) or ( a6084a );
 a6093a <=( a6092a ) or ( a6077a );
 a6097a <=( a2607a ) or ( a2608a );
 a6098a <=( a2609a ) or ( a6097a );
 a6101a <=( a2605a ) or ( a2606a );
 a6104a <=( a2603a ) or ( a2604a );
 a6105a <=( a6104a ) or ( a6101a );
 a6106a <=( a6105a ) or ( a6098a );
 a6109a <=( a2601a ) or ( a2602a );
 a6112a <=( a2599a ) or ( a2600a );
 a6113a <=( a6112a ) or ( a6109a );
 a6116a <=( a2597a ) or ( a2598a );
 a6119a <=( a2595a ) or ( a2596a );
 a6120a <=( a6119a ) or ( a6116a );
 a6121a <=( a6120a ) or ( a6113a );
 a6122a <=( a6121a ) or ( a6106a );
 a6123a <=( a6122a ) or ( a6093a );
 a6124a <=( a6123a ) or ( a6064a );
 a6125a <=( a6124a ) or ( a6007a );
 a6126a <=( a6125a ) or ( a5890a );
 a6130a <=( a2592a ) or ( a2593a );
 a6131a <=( a2594a ) or ( a6130a );
 a6134a <=( a2590a ) or ( a2591a );
 a6137a <=( a2588a ) or ( a2589a );
 a6138a <=( a6137a ) or ( a6134a );
 a6139a <=( a6138a ) or ( a6131a );
 a6143a <=( a2585a ) or ( a2586a );
 a6144a <=( a2587a ) or ( a6143a );
 a6147a <=( a2583a ) or ( a2584a );
 a6150a <=( a2581a ) or ( a2582a );
 a6151a <=( a6150a ) or ( a6147a );
 a6152a <=( a6151a ) or ( a6144a );
 a6153a <=( a6152a ) or ( a6139a );
 a6157a <=( a2578a ) or ( a2579a );
 a6158a <=( a2580a ) or ( a6157a );
 a6161a <=( a2576a ) or ( a2577a );
 a6164a <=( a2574a ) or ( a2575a );
 a6165a <=( a6164a ) or ( a6161a );
 a6166a <=( a6165a ) or ( a6158a );
 a6169a <=( a2572a ) or ( a2573a );
 a6172a <=( a2570a ) or ( a2571a );
 a6173a <=( a6172a ) or ( a6169a );
 a6176a <=( a2568a ) or ( a2569a );
 a6179a <=( a2566a ) or ( a2567a );
 a6180a <=( a6179a ) or ( a6176a );
 a6181a <=( a6180a ) or ( a6173a );
 a6182a <=( a6181a ) or ( a6166a );
 a6183a <=( a6182a ) or ( a6153a );
 a6187a <=( a2563a ) or ( a2564a );
 a6188a <=( a2565a ) or ( a6187a );
 a6191a <=( a2561a ) or ( a2562a );
 a6194a <=( a2559a ) or ( a2560a );
 a6195a <=( a6194a ) or ( a6191a );
 a6196a <=( a6195a ) or ( a6188a );
 a6199a <=( a2557a ) or ( a2558a );
 a6202a <=( a2555a ) or ( a2556a );
 a6203a <=( a6202a ) or ( a6199a );
 a6206a <=( a2553a ) or ( a2554a );
 a6209a <=( a2551a ) or ( a2552a );
 a6210a <=( a6209a ) or ( a6206a );
 a6211a <=( a6210a ) or ( a6203a );
 a6212a <=( a6211a ) or ( a6196a );
 a6216a <=( a2548a ) or ( a2549a );
 a6217a <=( a2550a ) or ( a6216a );
 a6220a <=( a2546a ) or ( a2547a );
 a6223a <=( a2544a ) or ( a2545a );
 a6224a <=( a6223a ) or ( a6220a );
 a6225a <=( a6224a ) or ( a6217a );
 a6228a <=( a2542a ) or ( a2543a );
 a6231a <=( a2540a ) or ( a2541a );
 a6232a <=( a6231a ) or ( a6228a );
 a6235a <=( a2538a ) or ( a2539a );
 a6238a <=( a2536a ) or ( a2537a );
 a6239a <=( a6238a ) or ( a6235a );
 a6240a <=( a6239a ) or ( a6232a );
 a6241a <=( a6240a ) or ( a6225a );
 a6242a <=( a6241a ) or ( a6212a );
 a6243a <=( a6242a ) or ( a6183a );
 a6247a <=( a2533a ) or ( a2534a );
 a6248a <=( a2535a ) or ( a6247a );
 a6251a <=( a2531a ) or ( a2532a );
 a6254a <=( a2529a ) or ( a2530a );
 a6255a <=( a6254a ) or ( a6251a );
 a6256a <=( a6255a ) or ( a6248a );
 a6260a <=( a2526a ) or ( a2527a );
 a6261a <=( a2528a ) or ( a6260a );
 a6264a <=( a2524a ) or ( a2525a );
 a6267a <=( a2522a ) or ( a2523a );
 a6268a <=( a6267a ) or ( a6264a );
 a6269a <=( a6268a ) or ( a6261a );
 a6270a <=( a6269a ) or ( a6256a );
 a6274a <=( a2519a ) or ( a2520a );
 a6275a <=( a2521a ) or ( a6274a );
 a6278a <=( a2517a ) or ( a2518a );
 a6281a <=( a2515a ) or ( a2516a );
 a6282a <=( a6281a ) or ( a6278a );
 a6283a <=( a6282a ) or ( a6275a );
 a6286a <=( a2513a ) or ( a2514a );
 a6289a <=( a2511a ) or ( a2512a );
 a6290a <=( a6289a ) or ( a6286a );
 a6293a <=( a2509a ) or ( a2510a );
 a6296a <=( a2507a ) or ( a2508a );
 a6297a <=( a6296a ) or ( a6293a );
 a6298a <=( a6297a ) or ( a6290a );
 a6299a <=( a6298a ) or ( a6283a );
 a6300a <=( a6299a ) or ( a6270a );
 a6304a <=( a2504a ) or ( a2505a );
 a6305a <=( a2506a ) or ( a6304a );
 a6308a <=( a2502a ) or ( a2503a );
 a6311a <=( a2500a ) or ( a2501a );
 a6312a <=( a6311a ) or ( a6308a );
 a6313a <=( a6312a ) or ( a6305a );
 a6316a <=( a2498a ) or ( a2499a );
 a6319a <=( a2496a ) or ( a2497a );
 a6320a <=( a6319a ) or ( a6316a );
 a6323a <=( a2494a ) or ( a2495a );
 a6326a <=( a2492a ) or ( a2493a );
 a6327a <=( a6326a ) or ( a6323a );
 a6328a <=( a6327a ) or ( a6320a );
 a6329a <=( a6328a ) or ( a6313a );
 a6333a <=( a2489a ) or ( a2490a );
 a6334a <=( a2491a ) or ( a6333a );
 a6337a <=( a2487a ) or ( a2488a );
 a6340a <=( a2485a ) or ( a2486a );
 a6341a <=( a6340a ) or ( a6337a );
 a6342a <=( a6341a ) or ( a6334a );
 a6345a <=( a2483a ) or ( a2484a );
 a6348a <=( a2481a ) or ( a2482a );
 a6349a <=( a6348a ) or ( a6345a );
 a6352a <=( a2479a ) or ( a2480a );
 a6355a <=( a2477a ) or ( a2478a );
 a6356a <=( a6355a ) or ( a6352a );
 a6357a <=( a6356a ) or ( a6349a );
 a6358a <=( a6357a ) or ( a6342a );
 a6359a <=( a6358a ) or ( a6329a );
 a6360a <=( a6359a ) or ( a6300a );
 a6361a <=( a6360a ) or ( a6243a );
 a6365a <=( a2474a ) or ( a2475a );
 a6366a <=( a2476a ) or ( a6365a );
 a6369a <=( a2472a ) or ( a2473a );
 a6372a <=( a2470a ) or ( a2471a );
 a6373a <=( a6372a ) or ( a6369a );
 a6374a <=( a6373a ) or ( a6366a );
 a6378a <=( a2467a ) or ( a2468a );
 a6379a <=( a2469a ) or ( a6378a );
 a6382a <=( a2465a ) or ( a2466a );
 a6385a <=( a2463a ) or ( a2464a );
 a6386a <=( a6385a ) or ( a6382a );
 a6387a <=( a6386a ) or ( a6379a );
 a6388a <=( a6387a ) or ( a6374a );
 a6392a <=( a2460a ) or ( a2461a );
 a6393a <=( a2462a ) or ( a6392a );
 a6396a <=( a2458a ) or ( a2459a );
 a6399a <=( a2456a ) or ( a2457a );
 a6400a <=( a6399a ) or ( a6396a );
 a6401a <=( a6400a ) or ( a6393a );
 a6404a <=( a2454a ) or ( a2455a );
 a6407a <=( a2452a ) or ( a2453a );
 a6408a <=( a6407a ) or ( a6404a );
 a6411a <=( a2450a ) or ( a2451a );
 a6414a <=( a2448a ) or ( a2449a );
 a6415a <=( a6414a ) or ( a6411a );
 a6416a <=( a6415a ) or ( a6408a );
 a6417a <=( a6416a ) or ( a6401a );
 a6418a <=( a6417a ) or ( a6388a );
 a6422a <=( a2445a ) or ( a2446a );
 a6423a <=( a2447a ) or ( a6422a );
 a6426a <=( a2443a ) or ( a2444a );
 a6429a <=( a2441a ) or ( a2442a );
 a6430a <=( a6429a ) or ( a6426a );
 a6431a <=( a6430a ) or ( a6423a );
 a6434a <=( a2439a ) or ( a2440a );
 a6437a <=( a2437a ) or ( a2438a );
 a6438a <=( a6437a ) or ( a6434a );
 a6441a <=( a2435a ) or ( a2436a );
 a6444a <=( a2433a ) or ( a2434a );
 a6445a <=( a6444a ) or ( a6441a );
 a6446a <=( a6445a ) or ( a6438a );
 a6447a <=( a6446a ) or ( a6431a );
 a6451a <=( a2430a ) or ( a2431a );
 a6452a <=( a2432a ) or ( a6451a );
 a6455a <=( a2428a ) or ( a2429a );
 a6458a <=( a2426a ) or ( a2427a );
 a6459a <=( a6458a ) or ( a6455a );
 a6460a <=( a6459a ) or ( a6452a );
 a6463a <=( a2424a ) or ( a2425a );
 a6466a <=( a2422a ) or ( a2423a );
 a6467a <=( a6466a ) or ( a6463a );
 a6470a <=( a2420a ) or ( a2421a );
 a6473a <=( a2418a ) or ( a2419a );
 a6474a <=( a6473a ) or ( a6470a );
 a6475a <=( a6474a ) or ( a6467a );
 a6476a <=( a6475a ) or ( a6460a );
 a6477a <=( a6476a ) or ( a6447a );
 a6478a <=( a6477a ) or ( a6418a );
 a6482a <=( a2415a ) or ( a2416a );
 a6483a <=( a2417a ) or ( a6482a );
 a6486a <=( a2413a ) or ( a2414a );
 a6489a <=( a2411a ) or ( a2412a );
 a6490a <=( a6489a ) or ( a6486a );
 a6491a <=( a6490a ) or ( a6483a );
 a6495a <=( a2408a ) or ( a2409a );
 a6496a <=( a2410a ) or ( a6495a );
 a6499a <=( a2406a ) or ( a2407a );
 a6502a <=( a2404a ) or ( a2405a );
 a6503a <=( a6502a ) or ( a6499a );
 a6504a <=( a6503a ) or ( a6496a );
 a6505a <=( a6504a ) or ( a6491a );
 a6509a <=( a2401a ) or ( a2402a );
 a6510a <=( a2403a ) or ( a6509a );
 a6513a <=( a2399a ) or ( a2400a );
 a6516a <=( a2397a ) or ( a2398a );
 a6517a <=( a6516a ) or ( a6513a );
 a6518a <=( a6517a ) or ( a6510a );
 a6521a <=( a2395a ) or ( a2396a );
 a6524a <=( a2393a ) or ( a2394a );
 a6525a <=( a6524a ) or ( a6521a );
 a6528a <=( a2391a ) or ( a2392a );
 a6531a <=( a2389a ) or ( a2390a );
 a6532a <=( a6531a ) or ( a6528a );
 a6533a <=( a6532a ) or ( a6525a );
 a6534a <=( a6533a ) or ( a6518a );
 a6535a <=( a6534a ) or ( a6505a );
 a6539a <=( a2386a ) or ( a2387a );
 a6540a <=( a2388a ) or ( a6539a );
 a6543a <=( a2384a ) or ( a2385a );
 a6546a <=( a2382a ) or ( a2383a );
 a6547a <=( a6546a ) or ( a6543a );
 a6548a <=( a6547a ) or ( a6540a );
 a6551a <=( a2380a ) or ( a2381a );
 a6554a <=( a2378a ) or ( a2379a );
 a6555a <=( a6554a ) or ( a6551a );
 a6558a <=( a2376a ) or ( a2377a );
 a6561a <=( a2374a ) or ( a2375a );
 a6562a <=( a6561a ) or ( a6558a );
 a6563a <=( a6562a ) or ( a6555a );
 a6564a <=( a6563a ) or ( a6548a );
 a6568a <=( a2371a ) or ( a2372a );
 a6569a <=( a2373a ) or ( a6568a );
 a6572a <=( a2369a ) or ( a2370a );
 a6575a <=( a2367a ) or ( a2368a );
 a6576a <=( a6575a ) or ( a6572a );
 a6577a <=( a6576a ) or ( a6569a );
 a6580a <=( a2365a ) or ( a2366a );
 a6583a <=( a2363a ) or ( a2364a );
 a6584a <=( a6583a ) or ( a6580a );
 a6587a <=( a2361a ) or ( a2362a );
 a6590a <=( a2359a ) or ( a2360a );
 a6591a <=( a6590a ) or ( a6587a );
 a6592a <=( a6591a ) or ( a6584a );
 a6593a <=( a6592a ) or ( a6577a );
 a6594a <=( a6593a ) or ( a6564a );
 a6595a <=( a6594a ) or ( a6535a );
 a6596a <=( a6595a ) or ( a6478a );
 a6597a <=( a6596a ) or ( a6361a );
 a6598a <=( a6597a ) or ( a6126a );
 a6602a <=( a2356a ) or ( a2357a );
 a6603a <=( a2358a ) or ( a6602a );
 a6606a <=( a2354a ) or ( a2355a );
 a6609a <=( a2352a ) or ( a2353a );
 a6610a <=( a6609a ) or ( a6606a );
 a6611a <=( a6610a ) or ( a6603a );
 a6615a <=( a2349a ) or ( a2350a );
 a6616a <=( a2351a ) or ( a6615a );
 a6619a <=( a2347a ) or ( a2348a );
 a6622a <=( a2345a ) or ( a2346a );
 a6623a <=( a6622a ) or ( a6619a );
 a6624a <=( a6623a ) or ( a6616a );
 a6625a <=( a6624a ) or ( a6611a );
 a6629a <=( a2342a ) or ( a2343a );
 a6630a <=( a2344a ) or ( a6629a );
 a6633a <=( a2340a ) or ( a2341a );
 a6636a <=( a2338a ) or ( a2339a );
 a6637a <=( a6636a ) or ( a6633a );
 a6638a <=( a6637a ) or ( a6630a );
 a6641a <=( a2336a ) or ( a2337a );
 a6644a <=( a2334a ) or ( a2335a );
 a6645a <=( a6644a ) or ( a6641a );
 a6648a <=( a2332a ) or ( a2333a );
 a6651a <=( a2330a ) or ( a2331a );
 a6652a <=( a6651a ) or ( a6648a );
 a6653a <=( a6652a ) or ( a6645a );
 a6654a <=( a6653a ) or ( a6638a );
 a6655a <=( a6654a ) or ( a6625a );
 a6659a <=( a2327a ) or ( a2328a );
 a6660a <=( a2329a ) or ( a6659a );
 a6663a <=( a2325a ) or ( a2326a );
 a6666a <=( a2323a ) or ( a2324a );
 a6667a <=( a6666a ) or ( a6663a );
 a6668a <=( a6667a ) or ( a6660a );
 a6671a <=( a2321a ) or ( a2322a );
 a6674a <=( a2319a ) or ( a2320a );
 a6675a <=( a6674a ) or ( a6671a );
 a6678a <=( a2317a ) or ( a2318a );
 a6681a <=( a2315a ) or ( a2316a );
 a6682a <=( a6681a ) or ( a6678a );
 a6683a <=( a6682a ) or ( a6675a );
 a6684a <=( a6683a ) or ( a6668a );
 a6688a <=( a2312a ) or ( a2313a );
 a6689a <=( a2314a ) or ( a6688a );
 a6692a <=( a2310a ) or ( a2311a );
 a6695a <=( a2308a ) or ( a2309a );
 a6696a <=( a6695a ) or ( a6692a );
 a6697a <=( a6696a ) or ( a6689a );
 a6700a <=( a2306a ) or ( a2307a );
 a6703a <=( a2304a ) or ( a2305a );
 a6704a <=( a6703a ) or ( a6700a );
 a6707a <=( a2302a ) or ( a2303a );
 a6710a <=( a2300a ) or ( a2301a );
 a6711a <=( a6710a ) or ( a6707a );
 a6712a <=( a6711a ) or ( a6704a );
 a6713a <=( a6712a ) or ( a6697a );
 a6714a <=( a6713a ) or ( a6684a );
 a6715a <=( a6714a ) or ( a6655a );
 a6719a <=( a2297a ) or ( a2298a );
 a6720a <=( a2299a ) or ( a6719a );
 a6723a <=( a2295a ) or ( a2296a );
 a6726a <=( a2293a ) or ( a2294a );
 a6727a <=( a6726a ) or ( a6723a );
 a6728a <=( a6727a ) or ( a6720a );
 a6732a <=( a2290a ) or ( a2291a );
 a6733a <=( a2292a ) or ( a6732a );
 a6736a <=( a2288a ) or ( a2289a );
 a6739a <=( a2286a ) or ( a2287a );
 a6740a <=( a6739a ) or ( a6736a );
 a6741a <=( a6740a ) or ( a6733a );
 a6742a <=( a6741a ) or ( a6728a );
 a6746a <=( a2283a ) or ( a2284a );
 a6747a <=( a2285a ) or ( a6746a );
 a6750a <=( a2281a ) or ( a2282a );
 a6753a <=( a2279a ) or ( a2280a );
 a6754a <=( a6753a ) or ( a6750a );
 a6755a <=( a6754a ) or ( a6747a );
 a6758a <=( a2277a ) or ( a2278a );
 a6761a <=( a2275a ) or ( a2276a );
 a6762a <=( a6761a ) or ( a6758a );
 a6765a <=( a2273a ) or ( a2274a );
 a6768a <=( a2271a ) or ( a2272a );
 a6769a <=( a6768a ) or ( a6765a );
 a6770a <=( a6769a ) or ( a6762a );
 a6771a <=( a6770a ) or ( a6755a );
 a6772a <=( a6771a ) or ( a6742a );
 a6776a <=( a2268a ) or ( a2269a );
 a6777a <=( a2270a ) or ( a6776a );
 a6780a <=( a2266a ) or ( a2267a );
 a6783a <=( a2264a ) or ( a2265a );
 a6784a <=( a6783a ) or ( a6780a );
 a6785a <=( a6784a ) or ( a6777a );
 a6788a <=( a2262a ) or ( a2263a );
 a6791a <=( a2260a ) or ( a2261a );
 a6792a <=( a6791a ) or ( a6788a );
 a6795a <=( a2258a ) or ( a2259a );
 a6798a <=( a2256a ) or ( a2257a );
 a6799a <=( a6798a ) or ( a6795a );
 a6800a <=( a6799a ) or ( a6792a );
 a6801a <=( a6800a ) or ( a6785a );
 a6805a <=( a2253a ) or ( a2254a );
 a6806a <=( a2255a ) or ( a6805a );
 a6809a <=( a2251a ) or ( a2252a );
 a6812a <=( a2249a ) or ( a2250a );
 a6813a <=( a6812a ) or ( a6809a );
 a6814a <=( a6813a ) or ( a6806a );
 a6817a <=( a2247a ) or ( a2248a );
 a6820a <=( a2245a ) or ( a2246a );
 a6821a <=( a6820a ) or ( a6817a );
 a6824a <=( a2243a ) or ( a2244a );
 a6827a <=( a2241a ) or ( a2242a );
 a6828a <=( a6827a ) or ( a6824a );
 a6829a <=( a6828a ) or ( a6821a );
 a6830a <=( a6829a ) or ( a6814a );
 a6831a <=( a6830a ) or ( a6801a );
 a6832a <=( a6831a ) or ( a6772a );
 a6833a <=( a6832a ) or ( a6715a );
 a6837a <=( a2238a ) or ( a2239a );
 a6838a <=( a2240a ) or ( a6837a );
 a6841a <=( a2236a ) or ( a2237a );
 a6844a <=( a2234a ) or ( a2235a );
 a6845a <=( a6844a ) or ( a6841a );
 a6846a <=( a6845a ) or ( a6838a );
 a6850a <=( a2231a ) or ( a2232a );
 a6851a <=( a2233a ) or ( a6850a );
 a6854a <=( a2229a ) or ( a2230a );
 a6857a <=( a2227a ) or ( a2228a );
 a6858a <=( a6857a ) or ( a6854a );
 a6859a <=( a6858a ) or ( a6851a );
 a6860a <=( a6859a ) or ( a6846a );
 a6864a <=( a2224a ) or ( a2225a );
 a6865a <=( a2226a ) or ( a6864a );
 a6868a <=( a2222a ) or ( a2223a );
 a6871a <=( a2220a ) or ( a2221a );
 a6872a <=( a6871a ) or ( a6868a );
 a6873a <=( a6872a ) or ( a6865a );
 a6876a <=( a2218a ) or ( a2219a );
 a6879a <=( a2216a ) or ( a2217a );
 a6880a <=( a6879a ) or ( a6876a );
 a6883a <=( a2214a ) or ( a2215a );
 a6886a <=( a2212a ) or ( a2213a );
 a6887a <=( a6886a ) or ( a6883a );
 a6888a <=( a6887a ) or ( a6880a );
 a6889a <=( a6888a ) or ( a6873a );
 a6890a <=( a6889a ) or ( a6860a );
 a6894a <=( a2209a ) or ( a2210a );
 a6895a <=( a2211a ) or ( a6894a );
 a6898a <=( a2207a ) or ( a2208a );
 a6901a <=( a2205a ) or ( a2206a );
 a6902a <=( a6901a ) or ( a6898a );
 a6903a <=( a6902a ) or ( a6895a );
 a6906a <=( a2203a ) or ( a2204a );
 a6909a <=( a2201a ) or ( a2202a );
 a6910a <=( a6909a ) or ( a6906a );
 a6913a <=( a2199a ) or ( a2200a );
 a6916a <=( a2197a ) or ( a2198a );
 a6917a <=( a6916a ) or ( a6913a );
 a6918a <=( a6917a ) or ( a6910a );
 a6919a <=( a6918a ) or ( a6903a );
 a6923a <=( a2194a ) or ( a2195a );
 a6924a <=( a2196a ) or ( a6923a );
 a6927a <=( a2192a ) or ( a2193a );
 a6930a <=( a2190a ) or ( a2191a );
 a6931a <=( a6930a ) or ( a6927a );
 a6932a <=( a6931a ) or ( a6924a );
 a6935a <=( a2188a ) or ( a2189a );
 a6938a <=( a2186a ) or ( a2187a );
 a6939a <=( a6938a ) or ( a6935a );
 a6942a <=( a2184a ) or ( a2185a );
 a6945a <=( a2182a ) or ( a2183a );
 a6946a <=( a6945a ) or ( a6942a );
 a6947a <=( a6946a ) or ( a6939a );
 a6948a <=( a6947a ) or ( a6932a );
 a6949a <=( a6948a ) or ( a6919a );
 a6950a <=( a6949a ) or ( a6890a );
 a6954a <=( a2179a ) or ( a2180a );
 a6955a <=( a2181a ) or ( a6954a );
 a6958a <=( a2177a ) or ( a2178a );
 a6961a <=( a2175a ) or ( a2176a );
 a6962a <=( a6961a ) or ( a6958a );
 a6963a <=( a6962a ) or ( a6955a );
 a6967a <=( a2172a ) or ( a2173a );
 a6968a <=( a2174a ) or ( a6967a );
 a6971a <=( a2170a ) or ( a2171a );
 a6974a <=( a2168a ) or ( a2169a );
 a6975a <=( a6974a ) or ( a6971a );
 a6976a <=( a6975a ) or ( a6968a );
 a6977a <=( a6976a ) or ( a6963a );
 a6981a <=( a2165a ) or ( a2166a );
 a6982a <=( a2167a ) or ( a6981a );
 a6985a <=( a2163a ) or ( a2164a );
 a6988a <=( a2161a ) or ( a2162a );
 a6989a <=( a6988a ) or ( a6985a );
 a6990a <=( a6989a ) or ( a6982a );
 a6993a <=( a2159a ) or ( a2160a );
 a6996a <=( a2157a ) or ( a2158a );
 a6997a <=( a6996a ) or ( a6993a );
 a7000a <=( a2155a ) or ( a2156a );
 a7003a <=( a2153a ) or ( a2154a );
 a7004a <=( a7003a ) or ( a7000a );
 a7005a <=( a7004a ) or ( a6997a );
 a7006a <=( a7005a ) or ( a6990a );
 a7007a <=( a7006a ) or ( a6977a );
 a7011a <=( a2150a ) or ( a2151a );
 a7012a <=( a2152a ) or ( a7011a );
 a7015a <=( a2148a ) or ( a2149a );
 a7018a <=( a2146a ) or ( a2147a );
 a7019a <=( a7018a ) or ( a7015a );
 a7020a <=( a7019a ) or ( a7012a );
 a7023a <=( a2144a ) or ( a2145a );
 a7026a <=( a2142a ) or ( a2143a );
 a7027a <=( a7026a ) or ( a7023a );
 a7030a <=( a2140a ) or ( a2141a );
 a7033a <=( a2138a ) or ( a2139a );
 a7034a <=( a7033a ) or ( a7030a );
 a7035a <=( a7034a ) or ( a7027a );
 a7036a <=( a7035a ) or ( a7020a );
 a7040a <=( a2135a ) or ( a2136a );
 a7041a <=( a2137a ) or ( a7040a );
 a7044a <=( a2133a ) or ( a2134a );
 a7047a <=( a2131a ) or ( a2132a );
 a7048a <=( a7047a ) or ( a7044a );
 a7049a <=( a7048a ) or ( a7041a );
 a7052a <=( a2129a ) or ( a2130a );
 a7055a <=( a2127a ) or ( a2128a );
 a7056a <=( a7055a ) or ( a7052a );
 a7059a <=( a2125a ) or ( a2126a );
 a7062a <=( a2123a ) or ( a2124a );
 a7063a <=( a7062a ) or ( a7059a );
 a7064a <=( a7063a ) or ( a7056a );
 a7065a <=( a7064a ) or ( a7049a );
 a7066a <=( a7065a ) or ( a7036a );
 a7067a <=( a7066a ) or ( a7007a );
 a7068a <=( a7067a ) or ( a6950a );
 a7069a <=( a7068a ) or ( a6833a );
 a7073a <=( a2120a ) or ( a2121a );
 a7074a <=( a2122a ) or ( a7073a );
 a7077a <=( a2118a ) or ( a2119a );
 a7080a <=( a2116a ) or ( a2117a );
 a7081a <=( a7080a ) or ( a7077a );
 a7082a <=( a7081a ) or ( a7074a );
 a7086a <=( a2113a ) or ( a2114a );
 a7087a <=( a2115a ) or ( a7086a );
 a7090a <=( a2111a ) or ( a2112a );
 a7093a <=( a2109a ) or ( a2110a );
 a7094a <=( a7093a ) or ( a7090a );
 a7095a <=( a7094a ) or ( a7087a );
 a7096a <=( a7095a ) or ( a7082a );
 a7100a <=( a2106a ) or ( a2107a );
 a7101a <=( a2108a ) or ( a7100a );
 a7104a <=( a2104a ) or ( a2105a );
 a7107a <=( a2102a ) or ( a2103a );
 a7108a <=( a7107a ) or ( a7104a );
 a7109a <=( a7108a ) or ( a7101a );
 a7112a <=( a2100a ) or ( a2101a );
 a7115a <=( a2098a ) or ( a2099a );
 a7116a <=( a7115a ) or ( a7112a );
 a7119a <=( a2096a ) or ( a2097a );
 a7122a <=( a2094a ) or ( a2095a );
 a7123a <=( a7122a ) or ( a7119a );
 a7124a <=( a7123a ) or ( a7116a );
 a7125a <=( a7124a ) or ( a7109a );
 a7126a <=( a7125a ) or ( a7096a );
 a7130a <=( a2091a ) or ( a2092a );
 a7131a <=( a2093a ) or ( a7130a );
 a7134a <=( a2089a ) or ( a2090a );
 a7137a <=( a2087a ) or ( a2088a );
 a7138a <=( a7137a ) or ( a7134a );
 a7139a <=( a7138a ) or ( a7131a );
 a7142a <=( a2085a ) or ( a2086a );
 a7145a <=( a2083a ) or ( a2084a );
 a7146a <=( a7145a ) or ( a7142a );
 a7149a <=( a2081a ) or ( a2082a );
 a7152a <=( a2079a ) or ( a2080a );
 a7153a <=( a7152a ) or ( a7149a );
 a7154a <=( a7153a ) or ( a7146a );
 a7155a <=( a7154a ) or ( a7139a );
 a7159a <=( a2076a ) or ( a2077a );
 a7160a <=( a2078a ) or ( a7159a );
 a7163a <=( a2074a ) or ( a2075a );
 a7166a <=( a2072a ) or ( a2073a );
 a7167a <=( a7166a ) or ( a7163a );
 a7168a <=( a7167a ) or ( a7160a );
 a7171a <=( a2070a ) or ( a2071a );
 a7174a <=( a2068a ) or ( a2069a );
 a7175a <=( a7174a ) or ( a7171a );
 a7178a <=( a2066a ) or ( a2067a );
 a7181a <=( a2064a ) or ( a2065a );
 a7182a <=( a7181a ) or ( a7178a );
 a7183a <=( a7182a ) or ( a7175a );
 a7184a <=( a7183a ) or ( a7168a );
 a7185a <=( a7184a ) or ( a7155a );
 a7186a <=( a7185a ) or ( a7126a );
 a7190a <=( a2061a ) or ( a2062a );
 a7191a <=( a2063a ) or ( a7190a );
 a7194a <=( a2059a ) or ( a2060a );
 a7197a <=( a2057a ) or ( a2058a );
 a7198a <=( a7197a ) or ( a7194a );
 a7199a <=( a7198a ) or ( a7191a );
 a7203a <=( a2054a ) or ( a2055a );
 a7204a <=( a2056a ) or ( a7203a );
 a7207a <=( a2052a ) or ( a2053a );
 a7210a <=( a2050a ) or ( a2051a );
 a7211a <=( a7210a ) or ( a7207a );
 a7212a <=( a7211a ) or ( a7204a );
 a7213a <=( a7212a ) or ( a7199a );
 a7217a <=( a2047a ) or ( a2048a );
 a7218a <=( a2049a ) or ( a7217a );
 a7221a <=( a2045a ) or ( a2046a );
 a7224a <=( a2043a ) or ( a2044a );
 a7225a <=( a7224a ) or ( a7221a );
 a7226a <=( a7225a ) or ( a7218a );
 a7229a <=( a2041a ) or ( a2042a );
 a7232a <=( a2039a ) or ( a2040a );
 a7233a <=( a7232a ) or ( a7229a );
 a7236a <=( a2037a ) or ( a2038a );
 a7239a <=( a2035a ) or ( a2036a );
 a7240a <=( a7239a ) or ( a7236a );
 a7241a <=( a7240a ) or ( a7233a );
 a7242a <=( a7241a ) or ( a7226a );
 a7243a <=( a7242a ) or ( a7213a );
 a7247a <=( a2032a ) or ( a2033a );
 a7248a <=( a2034a ) or ( a7247a );
 a7251a <=( a2030a ) or ( a2031a );
 a7254a <=( a2028a ) or ( a2029a );
 a7255a <=( a7254a ) or ( a7251a );
 a7256a <=( a7255a ) or ( a7248a );
 a7259a <=( a2026a ) or ( a2027a );
 a7262a <=( a2024a ) or ( a2025a );
 a7263a <=( a7262a ) or ( a7259a );
 a7266a <=( a2022a ) or ( a2023a );
 a7269a <=( a2020a ) or ( a2021a );
 a7270a <=( a7269a ) or ( a7266a );
 a7271a <=( a7270a ) or ( a7263a );
 a7272a <=( a7271a ) or ( a7256a );
 a7276a <=( a2017a ) or ( a2018a );
 a7277a <=( a2019a ) or ( a7276a );
 a7280a <=( a2015a ) or ( a2016a );
 a7283a <=( a2013a ) or ( a2014a );
 a7284a <=( a7283a ) or ( a7280a );
 a7285a <=( a7284a ) or ( a7277a );
 a7288a <=( a2011a ) or ( a2012a );
 a7291a <=( a2009a ) or ( a2010a );
 a7292a <=( a7291a ) or ( a7288a );
 a7295a <=( a2007a ) or ( a2008a );
 a7298a <=( a2005a ) or ( a2006a );
 a7299a <=( a7298a ) or ( a7295a );
 a7300a <=( a7299a ) or ( a7292a );
 a7301a <=( a7300a ) or ( a7285a );
 a7302a <=( a7301a ) or ( a7272a );
 a7303a <=( a7302a ) or ( a7243a );
 a7304a <=( a7303a ) or ( a7186a );
 a7308a <=( a2002a ) or ( a2003a );
 a7309a <=( a2004a ) or ( a7308a );
 a7312a <=( a2000a ) or ( a2001a );
 a7315a <=( a1998a ) or ( a1999a );
 a7316a <=( a7315a ) or ( a7312a );
 a7317a <=( a7316a ) or ( a7309a );
 a7321a <=( a1995a ) or ( a1996a );
 a7322a <=( a1997a ) or ( a7321a );
 a7325a <=( a1993a ) or ( a1994a );
 a7328a <=( a1991a ) or ( a1992a );
 a7329a <=( a7328a ) or ( a7325a );
 a7330a <=( a7329a ) or ( a7322a );
 a7331a <=( a7330a ) or ( a7317a );
 a7335a <=( a1988a ) or ( a1989a );
 a7336a <=( a1990a ) or ( a7335a );
 a7339a <=( a1986a ) or ( a1987a );
 a7342a <=( a1984a ) or ( a1985a );
 a7343a <=( a7342a ) or ( a7339a );
 a7344a <=( a7343a ) or ( a7336a );
 a7347a <=( a1982a ) or ( a1983a );
 a7350a <=( a1980a ) or ( a1981a );
 a7351a <=( a7350a ) or ( a7347a );
 a7354a <=( a1978a ) or ( a1979a );
 a7357a <=( a1976a ) or ( a1977a );
 a7358a <=( a7357a ) or ( a7354a );
 a7359a <=( a7358a ) or ( a7351a );
 a7360a <=( a7359a ) or ( a7344a );
 a7361a <=( a7360a ) or ( a7331a );
 a7365a <=( a1973a ) or ( a1974a );
 a7366a <=( a1975a ) or ( a7365a );
 a7369a <=( a1971a ) or ( a1972a );
 a7372a <=( a1969a ) or ( a1970a );
 a7373a <=( a7372a ) or ( a7369a );
 a7374a <=( a7373a ) or ( a7366a );
 a7377a <=( a1967a ) or ( a1968a );
 a7380a <=( a1965a ) or ( a1966a );
 a7381a <=( a7380a ) or ( a7377a );
 a7384a <=( a1963a ) or ( a1964a );
 a7387a <=( a1961a ) or ( a1962a );
 a7388a <=( a7387a ) or ( a7384a );
 a7389a <=( a7388a ) or ( a7381a );
 a7390a <=( a7389a ) or ( a7374a );
 a7394a <=( a1958a ) or ( a1959a );
 a7395a <=( a1960a ) or ( a7394a );
 a7398a <=( a1956a ) or ( a1957a );
 a7401a <=( a1954a ) or ( a1955a );
 a7402a <=( a7401a ) or ( a7398a );
 a7403a <=( a7402a ) or ( a7395a );
 a7406a <=( a1952a ) or ( a1953a );
 a7409a <=( a1950a ) or ( a1951a );
 a7410a <=( a7409a ) or ( a7406a );
 a7413a <=( a1948a ) or ( a1949a );
 a7416a <=( a1946a ) or ( a1947a );
 a7417a <=( a7416a ) or ( a7413a );
 a7418a <=( a7417a ) or ( a7410a );
 a7419a <=( a7418a ) or ( a7403a );
 a7420a <=( a7419a ) or ( a7390a );
 a7421a <=( a7420a ) or ( a7361a );
 a7425a <=( a1943a ) or ( a1944a );
 a7426a <=( a1945a ) or ( a7425a );
 a7429a <=( a1941a ) or ( a1942a );
 a7432a <=( a1939a ) or ( a1940a );
 a7433a <=( a7432a ) or ( a7429a );
 a7434a <=( a7433a ) or ( a7426a );
 a7438a <=( a1936a ) or ( a1937a );
 a7439a <=( a1938a ) or ( a7438a );
 a7442a <=( a1934a ) or ( a1935a );
 a7445a <=( a1932a ) or ( a1933a );
 a7446a <=( a7445a ) or ( a7442a );
 a7447a <=( a7446a ) or ( a7439a );
 a7448a <=( a7447a ) or ( a7434a );
 a7452a <=( a1929a ) or ( a1930a );
 a7453a <=( a1931a ) or ( a7452a );
 a7456a <=( a1927a ) or ( a1928a );
 a7459a <=( a1925a ) or ( a1926a );
 a7460a <=( a7459a ) or ( a7456a );
 a7461a <=( a7460a ) or ( a7453a );
 a7464a <=( a1923a ) or ( a1924a );
 a7467a <=( a1921a ) or ( a1922a );
 a7468a <=( a7467a ) or ( a7464a );
 a7471a <=( a1919a ) or ( a1920a );
 a7474a <=( a1917a ) or ( a1918a );
 a7475a <=( a7474a ) or ( a7471a );
 a7476a <=( a7475a ) or ( a7468a );
 a7477a <=( a7476a ) or ( a7461a );
 a7478a <=( a7477a ) or ( a7448a );
 a7482a <=( a1914a ) or ( a1915a );
 a7483a <=( a1916a ) or ( a7482a );
 a7486a <=( a1912a ) or ( a1913a );
 a7489a <=( a1910a ) or ( a1911a );
 a7490a <=( a7489a ) or ( a7486a );
 a7491a <=( a7490a ) or ( a7483a );
 a7494a <=( a1908a ) or ( a1909a );
 a7497a <=( a1906a ) or ( a1907a );
 a7498a <=( a7497a ) or ( a7494a );
 a7501a <=( a1904a ) or ( a1905a );
 a7504a <=( a1902a ) or ( a1903a );
 a7505a <=( a7504a ) or ( a7501a );
 a7506a <=( a7505a ) or ( a7498a );
 a7507a <=( a7506a ) or ( a7491a );
 a7511a <=( a1899a ) or ( a1900a );
 a7512a <=( a1901a ) or ( a7511a );
 a7515a <=( a1897a ) or ( a1898a );
 a7518a <=( a1895a ) or ( a1896a );
 a7519a <=( a7518a ) or ( a7515a );
 a7520a <=( a7519a ) or ( a7512a );
 a7523a <=( a1893a ) or ( a1894a );
 a7526a <=( a1891a ) or ( a1892a );
 a7527a <=( a7526a ) or ( a7523a );
 a7530a <=( a1889a ) or ( a1890a );
 a7533a <=( a1887a ) or ( a1888a );
 a7534a <=( a7533a ) or ( a7530a );
 a7535a <=( a7534a ) or ( a7527a );
 a7536a <=( a7535a ) or ( a7520a );
 a7537a <=( a7536a ) or ( a7507a );
 a7538a <=( a7537a ) or ( a7478a );
 a7539a <=( a7538a ) or ( a7421a );
 a7540a <=( a7539a ) or ( a7304a );
 a7541a <=( a7540a ) or ( a7069a );
 a7542a <=( a7541a ) or ( a6598a );
 a7543a <=( a7542a ) or ( a5657a );
 a7547a <=( a1884a ) or ( a1885a );
 a7548a <=( a1886a ) or ( a7547a );
 a7551a <=( a1882a ) or ( a1883a );
 a7554a <=( a1880a ) or ( a1881a );
 a7555a <=( a7554a ) or ( a7551a );
 a7556a <=( a7555a ) or ( a7548a );
 a7560a <=( a1877a ) or ( a1878a );
 a7561a <=( a1879a ) or ( a7560a );
 a7564a <=( a1875a ) or ( a1876a );
 a7567a <=( a1873a ) or ( a1874a );
 a7568a <=( a7567a ) or ( a7564a );
 a7569a <=( a7568a ) or ( a7561a );
 a7570a <=( a7569a ) or ( a7556a );
 a7574a <=( a1870a ) or ( a1871a );
 a7575a <=( a1872a ) or ( a7574a );
 a7578a <=( a1868a ) or ( a1869a );
 a7581a <=( a1866a ) or ( a1867a );
 a7582a <=( a7581a ) or ( a7578a );
 a7583a <=( a7582a ) or ( a7575a );
 a7586a <=( a1864a ) or ( a1865a );
 a7589a <=( a1862a ) or ( a1863a );
 a7590a <=( a7589a ) or ( a7586a );
 a7593a <=( a1860a ) or ( a1861a );
 a7596a <=( a1858a ) or ( a1859a );
 a7597a <=( a7596a ) or ( a7593a );
 a7598a <=( a7597a ) or ( a7590a );
 a7599a <=( a7598a ) or ( a7583a );
 a7600a <=( a7599a ) or ( a7570a );
 a7604a <=( a1855a ) or ( a1856a );
 a7605a <=( a1857a ) or ( a7604a );
 a7608a <=( a1853a ) or ( a1854a );
 a7611a <=( a1851a ) or ( a1852a );
 a7612a <=( a7611a ) or ( a7608a );
 a7613a <=( a7612a ) or ( a7605a );
 a7617a <=( a1848a ) or ( a1849a );
 a7618a <=( a1850a ) or ( a7617a );
 a7621a <=( a1846a ) or ( a1847a );
 a7624a <=( a1844a ) or ( a1845a );
 a7625a <=( a7624a ) or ( a7621a );
 a7626a <=( a7625a ) or ( a7618a );
 a7627a <=( a7626a ) or ( a7613a );
 a7631a <=( a1841a ) or ( a1842a );
 a7632a <=( a1843a ) or ( a7631a );
 a7635a <=( a1839a ) or ( a1840a );
 a7638a <=( a1837a ) or ( a1838a );
 a7639a <=( a7638a ) or ( a7635a );
 a7640a <=( a7639a ) or ( a7632a );
 a7643a <=( a1835a ) or ( a1836a );
 a7646a <=( a1833a ) or ( a1834a );
 a7647a <=( a7646a ) or ( a7643a );
 a7650a <=( a1831a ) or ( a1832a );
 a7653a <=( a1829a ) or ( a1830a );
 a7654a <=( a7653a ) or ( a7650a );
 a7655a <=( a7654a ) or ( a7647a );
 a7656a <=( a7655a ) or ( a7640a );
 a7657a <=( a7656a ) or ( a7627a );
 a7658a <=( a7657a ) or ( a7600a );
 a7662a <=( a1826a ) or ( a1827a );
 a7663a <=( a1828a ) or ( a7662a );
 a7666a <=( a1824a ) or ( a1825a );
 a7669a <=( a1822a ) or ( a1823a );
 a7670a <=( a7669a ) or ( a7666a );
 a7671a <=( a7670a ) or ( a7663a );
 a7675a <=( a1819a ) or ( a1820a );
 a7676a <=( a1821a ) or ( a7675a );
 a7679a <=( a1817a ) or ( a1818a );
 a7682a <=( a1815a ) or ( a1816a );
 a7683a <=( a7682a ) or ( a7679a );
 a7684a <=( a7683a ) or ( a7676a );
 a7685a <=( a7684a ) or ( a7671a );
 a7689a <=( a1812a ) or ( a1813a );
 a7690a <=( a1814a ) or ( a7689a );
 a7693a <=( a1810a ) or ( a1811a );
 a7696a <=( a1808a ) or ( a1809a );
 a7697a <=( a7696a ) or ( a7693a );
 a7698a <=( a7697a ) or ( a7690a );
 a7701a <=( a1806a ) or ( a1807a );
 a7704a <=( a1804a ) or ( a1805a );
 a7705a <=( a7704a ) or ( a7701a );
 a7708a <=( a1802a ) or ( a1803a );
 a7711a <=( a1800a ) or ( a1801a );
 a7712a <=( a7711a ) or ( a7708a );
 a7713a <=( a7712a ) or ( a7705a );
 a7714a <=( a7713a ) or ( a7698a );
 a7715a <=( a7714a ) or ( a7685a );
 a7719a <=( a1797a ) or ( a1798a );
 a7720a <=( a1799a ) or ( a7719a );
 a7723a <=( a1795a ) or ( a1796a );
 a7726a <=( a1793a ) or ( a1794a );
 a7727a <=( a7726a ) or ( a7723a );
 a7728a <=( a7727a ) or ( a7720a );
 a7731a <=( a1791a ) or ( a1792a );
 a7734a <=( a1789a ) or ( a1790a );
 a7735a <=( a7734a ) or ( a7731a );
 a7738a <=( a1787a ) or ( a1788a );
 a7741a <=( a1785a ) or ( a1786a );
 a7742a <=( a7741a ) or ( a7738a );
 a7743a <=( a7742a ) or ( a7735a );
 a7744a <=( a7743a ) or ( a7728a );
 a7748a <=( a1782a ) or ( a1783a );
 a7749a <=( a1784a ) or ( a7748a );
 a7752a <=( a1780a ) or ( a1781a );
 a7755a <=( a1778a ) or ( a1779a );
 a7756a <=( a7755a ) or ( a7752a );
 a7757a <=( a7756a ) or ( a7749a );
 a7760a <=( a1776a ) or ( a1777a );
 a7763a <=( a1774a ) or ( a1775a );
 a7764a <=( a7763a ) or ( a7760a );
 a7767a <=( a1772a ) or ( a1773a );
 a7770a <=( a1770a ) or ( a1771a );
 a7771a <=( a7770a ) or ( a7767a );
 a7772a <=( a7771a ) or ( a7764a );
 a7773a <=( a7772a ) or ( a7757a );
 a7774a <=( a7773a ) or ( a7744a );
 a7775a <=( a7774a ) or ( a7715a );
 a7776a <=( a7775a ) or ( a7658a );
 a7780a <=( a1767a ) or ( a1768a );
 a7781a <=( a1769a ) or ( a7780a );
 a7784a <=( a1765a ) or ( a1766a );
 a7787a <=( a1763a ) or ( a1764a );
 a7788a <=( a7787a ) or ( a7784a );
 a7789a <=( a7788a ) or ( a7781a );
 a7793a <=( a1760a ) or ( a1761a );
 a7794a <=( a1762a ) or ( a7793a );
 a7797a <=( a1758a ) or ( a1759a );
 a7800a <=( a1756a ) or ( a1757a );
 a7801a <=( a7800a ) or ( a7797a );
 a7802a <=( a7801a ) or ( a7794a );
 a7803a <=( a7802a ) or ( a7789a );
 a7807a <=( a1753a ) or ( a1754a );
 a7808a <=( a1755a ) or ( a7807a );
 a7811a <=( a1751a ) or ( a1752a );
 a7814a <=( a1749a ) or ( a1750a );
 a7815a <=( a7814a ) or ( a7811a );
 a7816a <=( a7815a ) or ( a7808a );
 a7819a <=( a1747a ) or ( a1748a );
 a7822a <=( a1745a ) or ( a1746a );
 a7823a <=( a7822a ) or ( a7819a );
 a7826a <=( a1743a ) or ( a1744a );
 a7829a <=( a1741a ) or ( a1742a );
 a7830a <=( a7829a ) or ( a7826a );
 a7831a <=( a7830a ) or ( a7823a );
 a7832a <=( a7831a ) or ( a7816a );
 a7833a <=( a7832a ) or ( a7803a );
 a7837a <=( a1738a ) or ( a1739a );
 a7838a <=( a1740a ) or ( a7837a );
 a7841a <=( a1736a ) or ( a1737a );
 a7844a <=( a1734a ) or ( a1735a );
 a7845a <=( a7844a ) or ( a7841a );
 a7846a <=( a7845a ) or ( a7838a );
 a7849a <=( a1732a ) or ( a1733a );
 a7852a <=( a1730a ) or ( a1731a );
 a7853a <=( a7852a ) or ( a7849a );
 a7856a <=( a1728a ) or ( a1729a );
 a7859a <=( a1726a ) or ( a1727a );
 a7860a <=( a7859a ) or ( a7856a );
 a7861a <=( a7860a ) or ( a7853a );
 a7862a <=( a7861a ) or ( a7846a );
 a7866a <=( a1723a ) or ( a1724a );
 a7867a <=( a1725a ) or ( a7866a );
 a7870a <=( a1721a ) or ( a1722a );
 a7873a <=( a1719a ) or ( a1720a );
 a7874a <=( a7873a ) or ( a7870a );
 a7875a <=( a7874a ) or ( a7867a );
 a7878a <=( a1717a ) or ( a1718a );
 a7881a <=( a1715a ) or ( a1716a );
 a7882a <=( a7881a ) or ( a7878a );
 a7885a <=( a1713a ) or ( a1714a );
 a7888a <=( a1711a ) or ( a1712a );
 a7889a <=( a7888a ) or ( a7885a );
 a7890a <=( a7889a ) or ( a7882a );
 a7891a <=( a7890a ) or ( a7875a );
 a7892a <=( a7891a ) or ( a7862a );
 a7893a <=( a7892a ) or ( a7833a );
 a7897a <=( a1708a ) or ( a1709a );
 a7898a <=( a1710a ) or ( a7897a );
 a7901a <=( a1706a ) or ( a1707a );
 a7904a <=( a1704a ) or ( a1705a );
 a7905a <=( a7904a ) or ( a7901a );
 a7906a <=( a7905a ) or ( a7898a );
 a7910a <=( a1701a ) or ( a1702a );
 a7911a <=( a1703a ) or ( a7910a );
 a7914a <=( a1699a ) or ( a1700a );
 a7917a <=( a1697a ) or ( a1698a );
 a7918a <=( a7917a ) or ( a7914a );
 a7919a <=( a7918a ) or ( a7911a );
 a7920a <=( a7919a ) or ( a7906a );
 a7924a <=( a1694a ) or ( a1695a );
 a7925a <=( a1696a ) or ( a7924a );
 a7928a <=( a1692a ) or ( a1693a );
 a7931a <=( a1690a ) or ( a1691a );
 a7932a <=( a7931a ) or ( a7928a );
 a7933a <=( a7932a ) or ( a7925a );
 a7936a <=( a1688a ) or ( a1689a );
 a7939a <=( a1686a ) or ( a1687a );
 a7940a <=( a7939a ) or ( a7936a );
 a7943a <=( a1684a ) or ( a1685a );
 a7946a <=( a1682a ) or ( a1683a );
 a7947a <=( a7946a ) or ( a7943a );
 a7948a <=( a7947a ) or ( a7940a );
 a7949a <=( a7948a ) or ( a7933a );
 a7950a <=( a7949a ) or ( a7920a );
 a7954a <=( a1679a ) or ( a1680a );
 a7955a <=( a1681a ) or ( a7954a );
 a7958a <=( a1677a ) or ( a1678a );
 a7961a <=( a1675a ) or ( a1676a );
 a7962a <=( a7961a ) or ( a7958a );
 a7963a <=( a7962a ) or ( a7955a );
 a7966a <=( a1673a ) or ( a1674a );
 a7969a <=( a1671a ) or ( a1672a );
 a7970a <=( a7969a ) or ( a7966a );
 a7973a <=( a1669a ) or ( a1670a );
 a7976a <=( a1667a ) or ( a1668a );
 a7977a <=( a7976a ) or ( a7973a );
 a7978a <=( a7977a ) or ( a7970a );
 a7979a <=( a7978a ) or ( a7963a );
 a7983a <=( a1664a ) or ( a1665a );
 a7984a <=( a1666a ) or ( a7983a );
 a7987a <=( a1662a ) or ( a1663a );
 a7990a <=( a1660a ) or ( a1661a );
 a7991a <=( a7990a ) or ( a7987a );
 a7992a <=( a7991a ) or ( a7984a );
 a7995a <=( a1658a ) or ( a1659a );
 a7998a <=( a1656a ) or ( a1657a );
 a7999a <=( a7998a ) or ( a7995a );
 a8002a <=( a1654a ) or ( a1655a );
 a8005a <=( a1652a ) or ( a1653a );
 a8006a <=( a8005a ) or ( a8002a );
 a8007a <=( a8006a ) or ( a7999a );
 a8008a <=( a8007a ) or ( a7992a );
 a8009a <=( a8008a ) or ( a7979a );
 a8010a <=( a8009a ) or ( a7950a );
 a8011a <=( a8010a ) or ( a7893a );
 a8012a <=( a8011a ) or ( a7776a );
 a8016a <=( a1649a ) or ( a1650a );
 a8017a <=( a1651a ) or ( a8016a );
 a8020a <=( a1647a ) or ( a1648a );
 a8023a <=( a1645a ) or ( a1646a );
 a8024a <=( a8023a ) or ( a8020a );
 a8025a <=( a8024a ) or ( a8017a );
 a8029a <=( a1642a ) or ( a1643a );
 a8030a <=( a1644a ) or ( a8029a );
 a8033a <=( a1640a ) or ( a1641a );
 a8036a <=( a1638a ) or ( a1639a );
 a8037a <=( a8036a ) or ( a8033a );
 a8038a <=( a8037a ) or ( a8030a );
 a8039a <=( a8038a ) or ( a8025a );
 a8043a <=( a1635a ) or ( a1636a );
 a8044a <=( a1637a ) or ( a8043a );
 a8047a <=( a1633a ) or ( a1634a );
 a8050a <=( a1631a ) or ( a1632a );
 a8051a <=( a8050a ) or ( a8047a );
 a8052a <=( a8051a ) or ( a8044a );
 a8055a <=( a1629a ) or ( a1630a );
 a8058a <=( a1627a ) or ( a1628a );
 a8059a <=( a8058a ) or ( a8055a );
 a8062a <=( a1625a ) or ( a1626a );
 a8065a <=( a1623a ) or ( a1624a );
 a8066a <=( a8065a ) or ( a8062a );
 a8067a <=( a8066a ) or ( a8059a );
 a8068a <=( a8067a ) or ( a8052a );
 a8069a <=( a8068a ) or ( a8039a );
 a8073a <=( a1620a ) or ( a1621a );
 a8074a <=( a1622a ) or ( a8073a );
 a8077a <=( a1618a ) or ( a1619a );
 a8080a <=( a1616a ) or ( a1617a );
 a8081a <=( a8080a ) or ( a8077a );
 a8082a <=( a8081a ) or ( a8074a );
 a8085a <=( a1614a ) or ( a1615a );
 a8088a <=( a1612a ) or ( a1613a );
 a8089a <=( a8088a ) or ( a8085a );
 a8092a <=( a1610a ) or ( a1611a );
 a8095a <=( a1608a ) or ( a1609a );
 a8096a <=( a8095a ) or ( a8092a );
 a8097a <=( a8096a ) or ( a8089a );
 a8098a <=( a8097a ) or ( a8082a );
 a8102a <=( a1605a ) or ( a1606a );
 a8103a <=( a1607a ) or ( a8102a );
 a8106a <=( a1603a ) or ( a1604a );
 a8109a <=( a1601a ) or ( a1602a );
 a8110a <=( a8109a ) or ( a8106a );
 a8111a <=( a8110a ) or ( a8103a );
 a8114a <=( a1599a ) or ( a1600a );
 a8117a <=( a1597a ) or ( a1598a );
 a8118a <=( a8117a ) or ( a8114a );
 a8121a <=( a1595a ) or ( a1596a );
 a8124a <=( a1593a ) or ( a1594a );
 a8125a <=( a8124a ) or ( a8121a );
 a8126a <=( a8125a ) or ( a8118a );
 a8127a <=( a8126a ) or ( a8111a );
 a8128a <=( a8127a ) or ( a8098a );
 a8129a <=( a8128a ) or ( a8069a );
 a8133a <=( a1590a ) or ( a1591a );
 a8134a <=( a1592a ) or ( a8133a );
 a8137a <=( a1588a ) or ( a1589a );
 a8140a <=( a1586a ) or ( a1587a );
 a8141a <=( a8140a ) or ( a8137a );
 a8142a <=( a8141a ) or ( a8134a );
 a8146a <=( a1583a ) or ( a1584a );
 a8147a <=( a1585a ) or ( a8146a );
 a8150a <=( a1581a ) or ( a1582a );
 a8153a <=( a1579a ) or ( a1580a );
 a8154a <=( a8153a ) or ( a8150a );
 a8155a <=( a8154a ) or ( a8147a );
 a8156a <=( a8155a ) or ( a8142a );
 a8160a <=( a1576a ) or ( a1577a );
 a8161a <=( a1578a ) or ( a8160a );
 a8164a <=( a1574a ) or ( a1575a );
 a8167a <=( a1572a ) or ( a1573a );
 a8168a <=( a8167a ) or ( a8164a );
 a8169a <=( a8168a ) or ( a8161a );
 a8172a <=( a1570a ) or ( a1571a );
 a8175a <=( a1568a ) or ( a1569a );
 a8176a <=( a8175a ) or ( a8172a );
 a8179a <=( a1566a ) or ( a1567a );
 a8182a <=( a1564a ) or ( a1565a );
 a8183a <=( a8182a ) or ( a8179a );
 a8184a <=( a8183a ) or ( a8176a );
 a8185a <=( a8184a ) or ( a8169a );
 a8186a <=( a8185a ) or ( a8156a );
 a8190a <=( a1561a ) or ( a1562a );
 a8191a <=( a1563a ) or ( a8190a );
 a8194a <=( a1559a ) or ( a1560a );
 a8197a <=( a1557a ) or ( a1558a );
 a8198a <=( a8197a ) or ( a8194a );
 a8199a <=( a8198a ) or ( a8191a );
 a8202a <=( a1555a ) or ( a1556a );
 a8205a <=( a1553a ) or ( a1554a );
 a8206a <=( a8205a ) or ( a8202a );
 a8209a <=( a1551a ) or ( a1552a );
 a8212a <=( a1549a ) or ( a1550a );
 a8213a <=( a8212a ) or ( a8209a );
 a8214a <=( a8213a ) or ( a8206a );
 a8215a <=( a8214a ) or ( a8199a );
 a8219a <=( a1546a ) or ( a1547a );
 a8220a <=( a1548a ) or ( a8219a );
 a8223a <=( a1544a ) or ( a1545a );
 a8226a <=( a1542a ) or ( a1543a );
 a8227a <=( a8226a ) or ( a8223a );
 a8228a <=( a8227a ) or ( a8220a );
 a8231a <=( a1540a ) or ( a1541a );
 a8234a <=( a1538a ) or ( a1539a );
 a8235a <=( a8234a ) or ( a8231a );
 a8238a <=( a1536a ) or ( a1537a );
 a8241a <=( a1534a ) or ( a1535a );
 a8242a <=( a8241a ) or ( a8238a );
 a8243a <=( a8242a ) or ( a8235a );
 a8244a <=( a8243a ) or ( a8228a );
 a8245a <=( a8244a ) or ( a8215a );
 a8246a <=( a8245a ) or ( a8186a );
 a8247a <=( a8246a ) or ( a8129a );
 a8251a <=( a1531a ) or ( a1532a );
 a8252a <=( a1533a ) or ( a8251a );
 a8255a <=( a1529a ) or ( a1530a );
 a8258a <=( a1527a ) or ( a1528a );
 a8259a <=( a8258a ) or ( a8255a );
 a8260a <=( a8259a ) or ( a8252a );
 a8264a <=( a1524a ) or ( a1525a );
 a8265a <=( a1526a ) or ( a8264a );
 a8268a <=( a1522a ) or ( a1523a );
 a8271a <=( a1520a ) or ( a1521a );
 a8272a <=( a8271a ) or ( a8268a );
 a8273a <=( a8272a ) or ( a8265a );
 a8274a <=( a8273a ) or ( a8260a );
 a8278a <=( a1517a ) or ( a1518a );
 a8279a <=( a1519a ) or ( a8278a );
 a8282a <=( a1515a ) or ( a1516a );
 a8285a <=( a1513a ) or ( a1514a );
 a8286a <=( a8285a ) or ( a8282a );
 a8287a <=( a8286a ) or ( a8279a );
 a8290a <=( a1511a ) or ( a1512a );
 a8293a <=( a1509a ) or ( a1510a );
 a8294a <=( a8293a ) or ( a8290a );
 a8297a <=( a1507a ) or ( a1508a );
 a8300a <=( a1505a ) or ( a1506a );
 a8301a <=( a8300a ) or ( a8297a );
 a8302a <=( a8301a ) or ( a8294a );
 a8303a <=( a8302a ) or ( a8287a );
 a8304a <=( a8303a ) or ( a8274a );
 a8308a <=( a1502a ) or ( a1503a );
 a8309a <=( a1504a ) or ( a8308a );
 a8312a <=( a1500a ) or ( a1501a );
 a8315a <=( a1498a ) or ( a1499a );
 a8316a <=( a8315a ) or ( a8312a );
 a8317a <=( a8316a ) or ( a8309a );
 a8320a <=( a1496a ) or ( a1497a );
 a8323a <=( a1494a ) or ( a1495a );
 a8324a <=( a8323a ) or ( a8320a );
 a8327a <=( a1492a ) or ( a1493a );
 a8330a <=( a1490a ) or ( a1491a );
 a8331a <=( a8330a ) or ( a8327a );
 a8332a <=( a8331a ) or ( a8324a );
 a8333a <=( a8332a ) or ( a8317a );
 a8337a <=( a1487a ) or ( a1488a );
 a8338a <=( a1489a ) or ( a8337a );
 a8341a <=( a1485a ) or ( a1486a );
 a8344a <=( a1483a ) or ( a1484a );
 a8345a <=( a8344a ) or ( a8341a );
 a8346a <=( a8345a ) or ( a8338a );
 a8349a <=( a1481a ) or ( a1482a );
 a8352a <=( a1479a ) or ( a1480a );
 a8353a <=( a8352a ) or ( a8349a );
 a8356a <=( a1477a ) or ( a1478a );
 a8359a <=( a1475a ) or ( a1476a );
 a8360a <=( a8359a ) or ( a8356a );
 a8361a <=( a8360a ) or ( a8353a );
 a8362a <=( a8361a ) or ( a8346a );
 a8363a <=( a8362a ) or ( a8333a );
 a8364a <=( a8363a ) or ( a8304a );
 a8368a <=( a1472a ) or ( a1473a );
 a8369a <=( a1474a ) or ( a8368a );
 a8372a <=( a1470a ) or ( a1471a );
 a8375a <=( a1468a ) or ( a1469a );
 a8376a <=( a8375a ) or ( a8372a );
 a8377a <=( a8376a ) or ( a8369a );
 a8381a <=( a1465a ) or ( a1466a );
 a8382a <=( a1467a ) or ( a8381a );
 a8385a <=( a1463a ) or ( a1464a );
 a8388a <=( a1461a ) or ( a1462a );
 a8389a <=( a8388a ) or ( a8385a );
 a8390a <=( a8389a ) or ( a8382a );
 a8391a <=( a8390a ) or ( a8377a );
 a8395a <=( a1458a ) or ( a1459a );
 a8396a <=( a1460a ) or ( a8395a );
 a8399a <=( a1456a ) or ( a1457a );
 a8402a <=( a1454a ) or ( a1455a );
 a8403a <=( a8402a ) or ( a8399a );
 a8404a <=( a8403a ) or ( a8396a );
 a8407a <=( a1452a ) or ( a1453a );
 a8410a <=( a1450a ) or ( a1451a );
 a8411a <=( a8410a ) or ( a8407a );
 a8414a <=( a1448a ) or ( a1449a );
 a8417a <=( a1446a ) or ( a1447a );
 a8418a <=( a8417a ) or ( a8414a );
 a8419a <=( a8418a ) or ( a8411a );
 a8420a <=( a8419a ) or ( a8404a );
 a8421a <=( a8420a ) or ( a8391a );
 a8425a <=( a1443a ) or ( a1444a );
 a8426a <=( a1445a ) or ( a8425a );
 a8429a <=( a1441a ) or ( a1442a );
 a8432a <=( a1439a ) or ( a1440a );
 a8433a <=( a8432a ) or ( a8429a );
 a8434a <=( a8433a ) or ( a8426a );
 a8437a <=( a1437a ) or ( a1438a );
 a8440a <=( a1435a ) or ( a1436a );
 a8441a <=( a8440a ) or ( a8437a );
 a8444a <=( a1433a ) or ( a1434a );
 a8447a <=( a1431a ) or ( a1432a );
 a8448a <=( a8447a ) or ( a8444a );
 a8449a <=( a8448a ) or ( a8441a );
 a8450a <=( a8449a ) or ( a8434a );
 a8454a <=( a1428a ) or ( a1429a );
 a8455a <=( a1430a ) or ( a8454a );
 a8458a <=( a1426a ) or ( a1427a );
 a8461a <=( a1424a ) or ( a1425a );
 a8462a <=( a8461a ) or ( a8458a );
 a8463a <=( a8462a ) or ( a8455a );
 a8466a <=( a1422a ) or ( a1423a );
 a8469a <=( a1420a ) or ( a1421a );
 a8470a <=( a8469a ) or ( a8466a );
 a8473a <=( a1418a ) or ( a1419a );
 a8476a <=( a1416a ) or ( a1417a );
 a8477a <=( a8476a ) or ( a8473a );
 a8478a <=( a8477a ) or ( a8470a );
 a8479a <=( a8478a ) or ( a8463a );
 a8480a <=( a8479a ) or ( a8450a );
 a8481a <=( a8480a ) or ( a8421a );
 a8482a <=( a8481a ) or ( a8364a );
 a8483a <=( a8482a ) or ( a8247a );
 a8484a <=( a8483a ) or ( a8012a );
 a8488a <=( a1413a ) or ( a1414a );
 a8489a <=( a1415a ) or ( a8488a );
 a8492a <=( a1411a ) or ( a1412a );
 a8495a <=( a1409a ) or ( a1410a );
 a8496a <=( a8495a ) or ( a8492a );
 a8497a <=( a8496a ) or ( a8489a );
 a8501a <=( a1406a ) or ( a1407a );
 a8502a <=( a1408a ) or ( a8501a );
 a8505a <=( a1404a ) or ( a1405a );
 a8508a <=( a1402a ) or ( a1403a );
 a8509a <=( a8508a ) or ( a8505a );
 a8510a <=( a8509a ) or ( a8502a );
 a8511a <=( a8510a ) or ( a8497a );
 a8515a <=( a1399a ) or ( a1400a );
 a8516a <=( a1401a ) or ( a8515a );
 a8519a <=( a1397a ) or ( a1398a );
 a8522a <=( a1395a ) or ( a1396a );
 a8523a <=( a8522a ) or ( a8519a );
 a8524a <=( a8523a ) or ( a8516a );
 a8527a <=( a1393a ) or ( a1394a );
 a8530a <=( a1391a ) or ( a1392a );
 a8531a <=( a8530a ) or ( a8527a );
 a8534a <=( a1389a ) or ( a1390a );
 a8537a <=( a1387a ) or ( a1388a );
 a8538a <=( a8537a ) or ( a8534a );
 a8539a <=( a8538a ) or ( a8531a );
 a8540a <=( a8539a ) or ( a8524a );
 a8541a <=( a8540a ) or ( a8511a );
 a8545a <=( a1384a ) or ( a1385a );
 a8546a <=( a1386a ) or ( a8545a );
 a8549a <=( a1382a ) or ( a1383a );
 a8552a <=( a1380a ) or ( a1381a );
 a8553a <=( a8552a ) or ( a8549a );
 a8554a <=( a8553a ) or ( a8546a );
 a8557a <=( a1378a ) or ( a1379a );
 a8560a <=( a1376a ) or ( a1377a );
 a8561a <=( a8560a ) or ( a8557a );
 a8564a <=( a1374a ) or ( a1375a );
 a8567a <=( a1372a ) or ( a1373a );
 a8568a <=( a8567a ) or ( a8564a );
 a8569a <=( a8568a ) or ( a8561a );
 a8570a <=( a8569a ) or ( a8554a );
 a8574a <=( a1369a ) or ( a1370a );
 a8575a <=( a1371a ) or ( a8574a );
 a8578a <=( a1367a ) or ( a1368a );
 a8581a <=( a1365a ) or ( a1366a );
 a8582a <=( a8581a ) or ( a8578a );
 a8583a <=( a8582a ) or ( a8575a );
 a8586a <=( a1363a ) or ( a1364a );
 a8589a <=( a1361a ) or ( a1362a );
 a8590a <=( a8589a ) or ( a8586a );
 a8593a <=( a1359a ) or ( a1360a );
 a8596a <=( a1357a ) or ( a1358a );
 a8597a <=( a8596a ) or ( a8593a );
 a8598a <=( a8597a ) or ( a8590a );
 a8599a <=( a8598a ) or ( a8583a );
 a8600a <=( a8599a ) or ( a8570a );
 a8601a <=( a8600a ) or ( a8541a );
 a8605a <=( a1354a ) or ( a1355a );
 a8606a <=( a1356a ) or ( a8605a );
 a8609a <=( a1352a ) or ( a1353a );
 a8612a <=( a1350a ) or ( a1351a );
 a8613a <=( a8612a ) or ( a8609a );
 a8614a <=( a8613a ) or ( a8606a );
 a8618a <=( a1347a ) or ( a1348a );
 a8619a <=( a1349a ) or ( a8618a );
 a8622a <=( a1345a ) or ( a1346a );
 a8625a <=( a1343a ) or ( a1344a );
 a8626a <=( a8625a ) or ( a8622a );
 a8627a <=( a8626a ) or ( a8619a );
 a8628a <=( a8627a ) or ( a8614a );
 a8632a <=( a1340a ) or ( a1341a );
 a8633a <=( a1342a ) or ( a8632a );
 a8636a <=( a1338a ) or ( a1339a );
 a8639a <=( a1336a ) or ( a1337a );
 a8640a <=( a8639a ) or ( a8636a );
 a8641a <=( a8640a ) or ( a8633a );
 a8644a <=( a1334a ) or ( a1335a );
 a8647a <=( a1332a ) or ( a1333a );
 a8648a <=( a8647a ) or ( a8644a );
 a8651a <=( a1330a ) or ( a1331a );
 a8654a <=( a1328a ) or ( a1329a );
 a8655a <=( a8654a ) or ( a8651a );
 a8656a <=( a8655a ) or ( a8648a );
 a8657a <=( a8656a ) or ( a8641a );
 a8658a <=( a8657a ) or ( a8628a );
 a8662a <=( a1325a ) or ( a1326a );
 a8663a <=( a1327a ) or ( a8662a );
 a8666a <=( a1323a ) or ( a1324a );
 a8669a <=( a1321a ) or ( a1322a );
 a8670a <=( a8669a ) or ( a8666a );
 a8671a <=( a8670a ) or ( a8663a );
 a8674a <=( a1319a ) or ( a1320a );
 a8677a <=( a1317a ) or ( a1318a );
 a8678a <=( a8677a ) or ( a8674a );
 a8681a <=( a1315a ) or ( a1316a );
 a8684a <=( a1313a ) or ( a1314a );
 a8685a <=( a8684a ) or ( a8681a );
 a8686a <=( a8685a ) or ( a8678a );
 a8687a <=( a8686a ) or ( a8671a );
 a8691a <=( a1310a ) or ( a1311a );
 a8692a <=( a1312a ) or ( a8691a );
 a8695a <=( a1308a ) or ( a1309a );
 a8698a <=( a1306a ) or ( a1307a );
 a8699a <=( a8698a ) or ( a8695a );
 a8700a <=( a8699a ) or ( a8692a );
 a8703a <=( a1304a ) or ( a1305a );
 a8706a <=( a1302a ) or ( a1303a );
 a8707a <=( a8706a ) or ( a8703a );
 a8710a <=( a1300a ) or ( a1301a );
 a8713a <=( a1298a ) or ( a1299a );
 a8714a <=( a8713a ) or ( a8710a );
 a8715a <=( a8714a ) or ( a8707a );
 a8716a <=( a8715a ) or ( a8700a );
 a8717a <=( a8716a ) or ( a8687a );
 a8718a <=( a8717a ) or ( a8658a );
 a8719a <=( a8718a ) or ( a8601a );
 a8723a <=( a1295a ) or ( a1296a );
 a8724a <=( a1297a ) or ( a8723a );
 a8727a <=( a1293a ) or ( a1294a );
 a8730a <=( a1291a ) or ( a1292a );
 a8731a <=( a8730a ) or ( a8727a );
 a8732a <=( a8731a ) or ( a8724a );
 a8736a <=( a1288a ) or ( a1289a );
 a8737a <=( a1290a ) or ( a8736a );
 a8740a <=( a1286a ) or ( a1287a );
 a8743a <=( a1284a ) or ( a1285a );
 a8744a <=( a8743a ) or ( a8740a );
 a8745a <=( a8744a ) or ( a8737a );
 a8746a <=( a8745a ) or ( a8732a );
 a8750a <=( a1281a ) or ( a1282a );
 a8751a <=( a1283a ) or ( a8750a );
 a8754a <=( a1279a ) or ( a1280a );
 a8757a <=( a1277a ) or ( a1278a );
 a8758a <=( a8757a ) or ( a8754a );
 a8759a <=( a8758a ) or ( a8751a );
 a8762a <=( a1275a ) or ( a1276a );
 a8765a <=( a1273a ) or ( a1274a );
 a8766a <=( a8765a ) or ( a8762a );
 a8769a <=( a1271a ) or ( a1272a );
 a8772a <=( a1269a ) or ( a1270a );
 a8773a <=( a8772a ) or ( a8769a );
 a8774a <=( a8773a ) or ( a8766a );
 a8775a <=( a8774a ) or ( a8759a );
 a8776a <=( a8775a ) or ( a8746a );
 a8780a <=( a1266a ) or ( a1267a );
 a8781a <=( a1268a ) or ( a8780a );
 a8784a <=( a1264a ) or ( a1265a );
 a8787a <=( a1262a ) or ( a1263a );
 a8788a <=( a8787a ) or ( a8784a );
 a8789a <=( a8788a ) or ( a8781a );
 a8792a <=( a1260a ) or ( a1261a );
 a8795a <=( a1258a ) or ( a1259a );
 a8796a <=( a8795a ) or ( a8792a );
 a8799a <=( a1256a ) or ( a1257a );
 a8802a <=( a1254a ) or ( a1255a );
 a8803a <=( a8802a ) or ( a8799a );
 a8804a <=( a8803a ) or ( a8796a );
 a8805a <=( a8804a ) or ( a8789a );
 a8809a <=( a1251a ) or ( a1252a );
 a8810a <=( a1253a ) or ( a8809a );
 a8813a <=( a1249a ) or ( a1250a );
 a8816a <=( a1247a ) or ( a1248a );
 a8817a <=( a8816a ) or ( a8813a );
 a8818a <=( a8817a ) or ( a8810a );
 a8821a <=( a1245a ) or ( a1246a );
 a8824a <=( a1243a ) or ( a1244a );
 a8825a <=( a8824a ) or ( a8821a );
 a8828a <=( a1241a ) or ( a1242a );
 a8831a <=( a1239a ) or ( a1240a );
 a8832a <=( a8831a ) or ( a8828a );
 a8833a <=( a8832a ) or ( a8825a );
 a8834a <=( a8833a ) or ( a8818a );
 a8835a <=( a8834a ) or ( a8805a );
 a8836a <=( a8835a ) or ( a8776a );
 a8840a <=( a1236a ) or ( a1237a );
 a8841a <=( a1238a ) or ( a8840a );
 a8844a <=( a1234a ) or ( a1235a );
 a8847a <=( a1232a ) or ( a1233a );
 a8848a <=( a8847a ) or ( a8844a );
 a8849a <=( a8848a ) or ( a8841a );
 a8853a <=( a1229a ) or ( a1230a );
 a8854a <=( a1231a ) or ( a8853a );
 a8857a <=( a1227a ) or ( a1228a );
 a8860a <=( a1225a ) or ( a1226a );
 a8861a <=( a8860a ) or ( a8857a );
 a8862a <=( a8861a ) or ( a8854a );
 a8863a <=( a8862a ) or ( a8849a );
 a8867a <=( a1222a ) or ( a1223a );
 a8868a <=( a1224a ) or ( a8867a );
 a8871a <=( a1220a ) or ( a1221a );
 a8874a <=( a1218a ) or ( a1219a );
 a8875a <=( a8874a ) or ( a8871a );
 a8876a <=( a8875a ) or ( a8868a );
 a8879a <=( a1216a ) or ( a1217a );
 a8882a <=( a1214a ) or ( a1215a );
 a8883a <=( a8882a ) or ( a8879a );
 a8886a <=( a1212a ) or ( a1213a );
 a8889a <=( a1210a ) or ( a1211a );
 a8890a <=( a8889a ) or ( a8886a );
 a8891a <=( a8890a ) or ( a8883a );
 a8892a <=( a8891a ) or ( a8876a );
 a8893a <=( a8892a ) or ( a8863a );
 a8897a <=( a1207a ) or ( a1208a );
 a8898a <=( a1209a ) or ( a8897a );
 a8901a <=( a1205a ) or ( a1206a );
 a8904a <=( a1203a ) or ( a1204a );
 a8905a <=( a8904a ) or ( a8901a );
 a8906a <=( a8905a ) or ( a8898a );
 a8909a <=( a1201a ) or ( a1202a );
 a8912a <=( a1199a ) or ( a1200a );
 a8913a <=( a8912a ) or ( a8909a );
 a8916a <=( a1197a ) or ( a1198a );
 a8919a <=( a1195a ) or ( a1196a );
 a8920a <=( a8919a ) or ( a8916a );
 a8921a <=( a8920a ) or ( a8913a );
 a8922a <=( a8921a ) or ( a8906a );
 a8926a <=( a1192a ) or ( a1193a );
 a8927a <=( a1194a ) or ( a8926a );
 a8930a <=( a1190a ) or ( a1191a );
 a8933a <=( a1188a ) or ( a1189a );
 a8934a <=( a8933a ) or ( a8930a );
 a8935a <=( a8934a ) or ( a8927a );
 a8938a <=( a1186a ) or ( a1187a );
 a8941a <=( a1184a ) or ( a1185a );
 a8942a <=( a8941a ) or ( a8938a );
 a8945a <=( a1182a ) or ( a1183a );
 a8948a <=( a1180a ) or ( a1181a );
 a8949a <=( a8948a ) or ( a8945a );
 a8950a <=( a8949a ) or ( a8942a );
 a8951a <=( a8950a ) or ( a8935a );
 a8952a <=( a8951a ) or ( a8922a );
 a8953a <=( a8952a ) or ( a8893a );
 a8954a <=( a8953a ) or ( a8836a );
 a8955a <=( a8954a ) or ( a8719a );
 a8959a <=( a1177a ) or ( a1178a );
 a8960a <=( a1179a ) or ( a8959a );
 a8963a <=( a1175a ) or ( a1176a );
 a8966a <=( a1173a ) or ( a1174a );
 a8967a <=( a8966a ) or ( a8963a );
 a8968a <=( a8967a ) or ( a8960a );
 a8972a <=( a1170a ) or ( a1171a );
 a8973a <=( a1172a ) or ( a8972a );
 a8976a <=( a1168a ) or ( a1169a );
 a8979a <=( a1166a ) or ( a1167a );
 a8980a <=( a8979a ) or ( a8976a );
 a8981a <=( a8980a ) or ( a8973a );
 a8982a <=( a8981a ) or ( a8968a );
 a8986a <=( a1163a ) or ( a1164a );
 a8987a <=( a1165a ) or ( a8986a );
 a8990a <=( a1161a ) or ( a1162a );
 a8993a <=( a1159a ) or ( a1160a );
 a8994a <=( a8993a ) or ( a8990a );
 a8995a <=( a8994a ) or ( a8987a );
 a8998a <=( a1157a ) or ( a1158a );
 a9001a <=( a1155a ) or ( a1156a );
 a9002a <=( a9001a ) or ( a8998a );
 a9005a <=( a1153a ) or ( a1154a );
 a9008a <=( a1151a ) or ( a1152a );
 a9009a <=( a9008a ) or ( a9005a );
 a9010a <=( a9009a ) or ( a9002a );
 a9011a <=( a9010a ) or ( a8995a );
 a9012a <=( a9011a ) or ( a8982a );
 a9016a <=( a1148a ) or ( a1149a );
 a9017a <=( a1150a ) or ( a9016a );
 a9020a <=( a1146a ) or ( a1147a );
 a9023a <=( a1144a ) or ( a1145a );
 a9024a <=( a9023a ) or ( a9020a );
 a9025a <=( a9024a ) or ( a9017a );
 a9028a <=( a1142a ) or ( a1143a );
 a9031a <=( a1140a ) or ( a1141a );
 a9032a <=( a9031a ) or ( a9028a );
 a9035a <=( a1138a ) or ( a1139a );
 a9038a <=( a1136a ) or ( a1137a );
 a9039a <=( a9038a ) or ( a9035a );
 a9040a <=( a9039a ) or ( a9032a );
 a9041a <=( a9040a ) or ( a9025a );
 a9045a <=( a1133a ) or ( a1134a );
 a9046a <=( a1135a ) or ( a9045a );
 a9049a <=( a1131a ) or ( a1132a );
 a9052a <=( a1129a ) or ( a1130a );
 a9053a <=( a9052a ) or ( a9049a );
 a9054a <=( a9053a ) or ( a9046a );
 a9057a <=( a1127a ) or ( a1128a );
 a9060a <=( a1125a ) or ( a1126a );
 a9061a <=( a9060a ) or ( a9057a );
 a9064a <=( a1123a ) or ( a1124a );
 a9067a <=( a1121a ) or ( a1122a );
 a9068a <=( a9067a ) or ( a9064a );
 a9069a <=( a9068a ) or ( a9061a );
 a9070a <=( a9069a ) or ( a9054a );
 a9071a <=( a9070a ) or ( a9041a );
 a9072a <=( a9071a ) or ( a9012a );
 a9076a <=( a1118a ) or ( a1119a );
 a9077a <=( a1120a ) or ( a9076a );
 a9080a <=( a1116a ) or ( a1117a );
 a9083a <=( a1114a ) or ( a1115a );
 a9084a <=( a9083a ) or ( a9080a );
 a9085a <=( a9084a ) or ( a9077a );
 a9089a <=( a1111a ) or ( a1112a );
 a9090a <=( a1113a ) or ( a9089a );
 a9093a <=( a1109a ) or ( a1110a );
 a9096a <=( a1107a ) or ( a1108a );
 a9097a <=( a9096a ) or ( a9093a );
 a9098a <=( a9097a ) or ( a9090a );
 a9099a <=( a9098a ) or ( a9085a );
 a9103a <=( a1104a ) or ( a1105a );
 a9104a <=( a1106a ) or ( a9103a );
 a9107a <=( a1102a ) or ( a1103a );
 a9110a <=( a1100a ) or ( a1101a );
 a9111a <=( a9110a ) or ( a9107a );
 a9112a <=( a9111a ) or ( a9104a );
 a9115a <=( a1098a ) or ( a1099a );
 a9118a <=( a1096a ) or ( a1097a );
 a9119a <=( a9118a ) or ( a9115a );
 a9122a <=( a1094a ) or ( a1095a );
 a9125a <=( a1092a ) or ( a1093a );
 a9126a <=( a9125a ) or ( a9122a );
 a9127a <=( a9126a ) or ( a9119a );
 a9128a <=( a9127a ) or ( a9112a );
 a9129a <=( a9128a ) or ( a9099a );
 a9133a <=( a1089a ) or ( a1090a );
 a9134a <=( a1091a ) or ( a9133a );
 a9137a <=( a1087a ) or ( a1088a );
 a9140a <=( a1085a ) or ( a1086a );
 a9141a <=( a9140a ) or ( a9137a );
 a9142a <=( a9141a ) or ( a9134a );
 a9145a <=( a1083a ) or ( a1084a );
 a9148a <=( a1081a ) or ( a1082a );
 a9149a <=( a9148a ) or ( a9145a );
 a9152a <=( a1079a ) or ( a1080a );
 a9155a <=( a1077a ) or ( a1078a );
 a9156a <=( a9155a ) or ( a9152a );
 a9157a <=( a9156a ) or ( a9149a );
 a9158a <=( a9157a ) or ( a9142a );
 a9162a <=( a1074a ) or ( a1075a );
 a9163a <=( a1076a ) or ( a9162a );
 a9166a <=( a1072a ) or ( a1073a );
 a9169a <=( a1070a ) or ( a1071a );
 a9170a <=( a9169a ) or ( a9166a );
 a9171a <=( a9170a ) or ( a9163a );
 a9174a <=( a1068a ) or ( a1069a );
 a9177a <=( a1066a ) or ( a1067a );
 a9178a <=( a9177a ) or ( a9174a );
 a9181a <=( a1064a ) or ( a1065a );
 a9184a <=( a1062a ) or ( a1063a );
 a9185a <=( a9184a ) or ( a9181a );
 a9186a <=( a9185a ) or ( a9178a );
 a9187a <=( a9186a ) or ( a9171a );
 a9188a <=( a9187a ) or ( a9158a );
 a9189a <=( a9188a ) or ( a9129a );
 a9190a <=( a9189a ) or ( a9072a );
 a9194a <=( a1059a ) or ( a1060a );
 a9195a <=( a1061a ) or ( a9194a );
 a9198a <=( a1057a ) or ( a1058a );
 a9201a <=( a1055a ) or ( a1056a );
 a9202a <=( a9201a ) or ( a9198a );
 a9203a <=( a9202a ) or ( a9195a );
 a9207a <=( a1052a ) or ( a1053a );
 a9208a <=( a1054a ) or ( a9207a );
 a9211a <=( a1050a ) or ( a1051a );
 a9214a <=( a1048a ) or ( a1049a );
 a9215a <=( a9214a ) or ( a9211a );
 a9216a <=( a9215a ) or ( a9208a );
 a9217a <=( a9216a ) or ( a9203a );
 a9221a <=( a1045a ) or ( a1046a );
 a9222a <=( a1047a ) or ( a9221a );
 a9225a <=( a1043a ) or ( a1044a );
 a9228a <=( a1041a ) or ( a1042a );
 a9229a <=( a9228a ) or ( a9225a );
 a9230a <=( a9229a ) or ( a9222a );
 a9233a <=( a1039a ) or ( a1040a );
 a9236a <=( a1037a ) or ( a1038a );
 a9237a <=( a9236a ) or ( a9233a );
 a9240a <=( a1035a ) or ( a1036a );
 a9243a <=( a1033a ) or ( a1034a );
 a9244a <=( a9243a ) or ( a9240a );
 a9245a <=( a9244a ) or ( a9237a );
 a9246a <=( a9245a ) or ( a9230a );
 a9247a <=( a9246a ) or ( a9217a );
 a9251a <=( a1030a ) or ( a1031a );
 a9252a <=( a1032a ) or ( a9251a );
 a9255a <=( a1028a ) or ( a1029a );
 a9258a <=( a1026a ) or ( a1027a );
 a9259a <=( a9258a ) or ( a9255a );
 a9260a <=( a9259a ) or ( a9252a );
 a9263a <=( a1024a ) or ( a1025a );
 a9266a <=( a1022a ) or ( a1023a );
 a9267a <=( a9266a ) or ( a9263a );
 a9270a <=( a1020a ) or ( a1021a );
 a9273a <=( a1018a ) or ( a1019a );
 a9274a <=( a9273a ) or ( a9270a );
 a9275a <=( a9274a ) or ( a9267a );
 a9276a <=( a9275a ) or ( a9260a );
 a9280a <=( a1015a ) or ( a1016a );
 a9281a <=( a1017a ) or ( a9280a );
 a9284a <=( a1013a ) or ( a1014a );
 a9287a <=( a1011a ) or ( a1012a );
 a9288a <=( a9287a ) or ( a9284a );
 a9289a <=( a9288a ) or ( a9281a );
 a9292a <=( a1009a ) or ( a1010a );
 a9295a <=( a1007a ) or ( a1008a );
 a9296a <=( a9295a ) or ( a9292a );
 a9299a <=( a1005a ) or ( a1006a );
 a9302a <=( a1003a ) or ( a1004a );
 a9303a <=( a9302a ) or ( a9299a );
 a9304a <=( a9303a ) or ( a9296a );
 a9305a <=( a9304a ) or ( a9289a );
 a9306a <=( a9305a ) or ( a9276a );
 a9307a <=( a9306a ) or ( a9247a );
 a9311a <=( a1000a ) or ( a1001a );
 a9312a <=( a1002a ) or ( a9311a );
 a9315a <=( a998a ) or ( a999a );
 a9318a <=( a996a ) or ( a997a );
 a9319a <=( a9318a ) or ( a9315a );
 a9320a <=( a9319a ) or ( a9312a );
 a9324a <=( a993a ) or ( a994a );
 a9325a <=( a995a ) or ( a9324a );
 a9328a <=( a991a ) or ( a992a );
 a9331a <=( a989a ) or ( a990a );
 a9332a <=( a9331a ) or ( a9328a );
 a9333a <=( a9332a ) or ( a9325a );
 a9334a <=( a9333a ) or ( a9320a );
 a9338a <=( a986a ) or ( a987a );
 a9339a <=( a988a ) or ( a9338a );
 a9342a <=( a984a ) or ( a985a );
 a9345a <=( a982a ) or ( a983a );
 a9346a <=( a9345a ) or ( a9342a );
 a9347a <=( a9346a ) or ( a9339a );
 a9350a <=( a980a ) or ( a981a );
 a9353a <=( a978a ) or ( a979a );
 a9354a <=( a9353a ) or ( a9350a );
 a9357a <=( a976a ) or ( a977a );
 a9360a <=( a974a ) or ( a975a );
 a9361a <=( a9360a ) or ( a9357a );
 a9362a <=( a9361a ) or ( a9354a );
 a9363a <=( a9362a ) or ( a9347a );
 a9364a <=( a9363a ) or ( a9334a );
 a9368a <=( a971a ) or ( a972a );
 a9369a <=( a973a ) or ( a9368a );
 a9372a <=( a969a ) or ( a970a );
 a9375a <=( a967a ) or ( a968a );
 a9376a <=( a9375a ) or ( a9372a );
 a9377a <=( a9376a ) or ( a9369a );
 a9380a <=( a965a ) or ( a966a );
 a9383a <=( a963a ) or ( a964a );
 a9384a <=( a9383a ) or ( a9380a );
 a9387a <=( a961a ) or ( a962a );
 a9390a <=( a959a ) or ( a960a );
 a9391a <=( a9390a ) or ( a9387a );
 a9392a <=( a9391a ) or ( a9384a );
 a9393a <=( a9392a ) or ( a9377a );
 a9397a <=( a956a ) or ( a957a );
 a9398a <=( a958a ) or ( a9397a );
 a9401a <=( a954a ) or ( a955a );
 a9404a <=( a952a ) or ( a953a );
 a9405a <=( a9404a ) or ( a9401a );
 a9406a <=( a9405a ) or ( a9398a );
 a9409a <=( a950a ) or ( a951a );
 a9412a <=( a948a ) or ( a949a );
 a9413a <=( a9412a ) or ( a9409a );
 a9416a <=( a946a ) or ( a947a );
 a9419a <=( a944a ) or ( a945a );
 a9420a <=( a9419a ) or ( a9416a );
 a9421a <=( a9420a ) or ( a9413a );
 a9422a <=( a9421a ) or ( a9406a );
 a9423a <=( a9422a ) or ( a9393a );
 a9424a <=( a9423a ) or ( a9364a );
 a9425a <=( a9424a ) or ( a9307a );
 a9426a <=( a9425a ) or ( a9190a );
 a9427a <=( a9426a ) or ( a8955a );
 a9428a <=( a9427a ) or ( a8484a );
 a9432a <=( a941a ) or ( a942a );
 a9433a <=( a943a ) or ( a9432a );
 a9436a <=( a939a ) or ( a940a );
 a9439a <=( a937a ) or ( a938a );
 a9440a <=( a9439a ) or ( a9436a );
 a9441a <=( a9440a ) or ( a9433a );
 a9445a <=( a934a ) or ( a935a );
 a9446a <=( a936a ) or ( a9445a );
 a9449a <=( a932a ) or ( a933a );
 a9452a <=( a930a ) or ( a931a );
 a9453a <=( a9452a ) or ( a9449a );
 a9454a <=( a9453a ) or ( a9446a );
 a9455a <=( a9454a ) or ( a9441a );
 a9459a <=( a927a ) or ( a928a );
 a9460a <=( a929a ) or ( a9459a );
 a9463a <=( a925a ) or ( a926a );
 a9466a <=( a923a ) or ( a924a );
 a9467a <=( a9466a ) or ( a9463a );
 a9468a <=( a9467a ) or ( a9460a );
 a9471a <=( a921a ) or ( a922a );
 a9474a <=( a919a ) or ( a920a );
 a9475a <=( a9474a ) or ( a9471a );
 a9478a <=( a917a ) or ( a918a );
 a9481a <=( a915a ) or ( a916a );
 a9482a <=( a9481a ) or ( a9478a );
 a9483a <=( a9482a ) or ( a9475a );
 a9484a <=( a9483a ) or ( a9468a );
 a9485a <=( a9484a ) or ( a9455a );
 a9489a <=( a912a ) or ( a913a );
 a9490a <=( a914a ) or ( a9489a );
 a9493a <=( a910a ) or ( a911a );
 a9496a <=( a908a ) or ( a909a );
 a9497a <=( a9496a ) or ( a9493a );
 a9498a <=( a9497a ) or ( a9490a );
 a9502a <=( a905a ) or ( a906a );
 a9503a <=( a907a ) or ( a9502a );
 a9506a <=( a903a ) or ( a904a );
 a9509a <=( a901a ) or ( a902a );
 a9510a <=( a9509a ) or ( a9506a );
 a9511a <=( a9510a ) or ( a9503a );
 a9512a <=( a9511a ) or ( a9498a );
 a9516a <=( a898a ) or ( a899a );
 a9517a <=( a900a ) or ( a9516a );
 a9520a <=( a896a ) or ( a897a );
 a9523a <=( a894a ) or ( a895a );
 a9524a <=( a9523a ) or ( a9520a );
 a9525a <=( a9524a ) or ( a9517a );
 a9528a <=( a892a ) or ( a893a );
 a9531a <=( a890a ) or ( a891a );
 a9532a <=( a9531a ) or ( a9528a );
 a9535a <=( a888a ) or ( a889a );
 a9538a <=( a886a ) or ( a887a );
 a9539a <=( a9538a ) or ( a9535a );
 a9540a <=( a9539a ) or ( a9532a );
 a9541a <=( a9540a ) or ( a9525a );
 a9542a <=( a9541a ) or ( a9512a );
 a9543a <=( a9542a ) or ( a9485a );
 a9547a <=( a883a ) or ( a884a );
 a9548a <=( a885a ) or ( a9547a );
 a9551a <=( a881a ) or ( a882a );
 a9554a <=( a879a ) or ( a880a );
 a9555a <=( a9554a ) or ( a9551a );
 a9556a <=( a9555a ) or ( a9548a );
 a9560a <=( a876a ) or ( a877a );
 a9561a <=( a878a ) or ( a9560a );
 a9564a <=( a874a ) or ( a875a );
 a9567a <=( a872a ) or ( a873a );
 a9568a <=( a9567a ) or ( a9564a );
 a9569a <=( a9568a ) or ( a9561a );
 a9570a <=( a9569a ) or ( a9556a );
 a9574a <=( a869a ) or ( a870a );
 a9575a <=( a871a ) or ( a9574a );
 a9578a <=( a867a ) or ( a868a );
 a9581a <=( a865a ) or ( a866a );
 a9582a <=( a9581a ) or ( a9578a );
 a9583a <=( a9582a ) or ( a9575a );
 a9586a <=( a863a ) or ( a864a );
 a9589a <=( a861a ) or ( a862a );
 a9590a <=( a9589a ) or ( a9586a );
 a9593a <=( a859a ) or ( a860a );
 a9596a <=( a857a ) or ( a858a );
 a9597a <=( a9596a ) or ( a9593a );
 a9598a <=( a9597a ) or ( a9590a );
 a9599a <=( a9598a ) or ( a9583a );
 a9600a <=( a9599a ) or ( a9570a );
 a9604a <=( a854a ) or ( a855a );
 a9605a <=( a856a ) or ( a9604a );
 a9608a <=( a852a ) or ( a853a );
 a9611a <=( a850a ) or ( a851a );
 a9612a <=( a9611a ) or ( a9608a );
 a9613a <=( a9612a ) or ( a9605a );
 a9616a <=( a848a ) or ( a849a );
 a9619a <=( a846a ) or ( a847a );
 a9620a <=( a9619a ) or ( a9616a );
 a9623a <=( a844a ) or ( a845a );
 a9626a <=( a842a ) or ( a843a );
 a9627a <=( a9626a ) or ( a9623a );
 a9628a <=( a9627a ) or ( a9620a );
 a9629a <=( a9628a ) or ( a9613a );
 a9633a <=( a839a ) or ( a840a );
 a9634a <=( a841a ) or ( a9633a );
 a9637a <=( a837a ) or ( a838a );
 a9640a <=( a835a ) or ( a836a );
 a9641a <=( a9640a ) or ( a9637a );
 a9642a <=( a9641a ) or ( a9634a );
 a9645a <=( a833a ) or ( a834a );
 a9648a <=( a831a ) or ( a832a );
 a9649a <=( a9648a ) or ( a9645a );
 a9652a <=( a829a ) or ( a830a );
 a9655a <=( a827a ) or ( a828a );
 a9656a <=( a9655a ) or ( a9652a );
 a9657a <=( a9656a ) or ( a9649a );
 a9658a <=( a9657a ) or ( a9642a );
 a9659a <=( a9658a ) or ( a9629a );
 a9660a <=( a9659a ) or ( a9600a );
 a9661a <=( a9660a ) or ( a9543a );
 a9665a <=( a824a ) or ( a825a );
 a9666a <=( a826a ) or ( a9665a );
 a9669a <=( a822a ) or ( a823a );
 a9672a <=( a820a ) or ( a821a );
 a9673a <=( a9672a ) or ( a9669a );
 a9674a <=( a9673a ) or ( a9666a );
 a9678a <=( a817a ) or ( a818a );
 a9679a <=( a819a ) or ( a9678a );
 a9682a <=( a815a ) or ( a816a );
 a9685a <=( a813a ) or ( a814a );
 a9686a <=( a9685a ) or ( a9682a );
 a9687a <=( a9686a ) or ( a9679a );
 a9688a <=( a9687a ) or ( a9674a );
 a9692a <=( a810a ) or ( a811a );
 a9693a <=( a812a ) or ( a9692a );
 a9696a <=( a808a ) or ( a809a );
 a9699a <=( a806a ) or ( a807a );
 a9700a <=( a9699a ) or ( a9696a );
 a9701a <=( a9700a ) or ( a9693a );
 a9704a <=( a804a ) or ( a805a );
 a9707a <=( a802a ) or ( a803a );
 a9708a <=( a9707a ) or ( a9704a );
 a9711a <=( a800a ) or ( a801a );
 a9714a <=( a798a ) or ( a799a );
 a9715a <=( a9714a ) or ( a9711a );
 a9716a <=( a9715a ) or ( a9708a );
 a9717a <=( a9716a ) or ( a9701a );
 a9718a <=( a9717a ) or ( a9688a );
 a9722a <=( a795a ) or ( a796a );
 a9723a <=( a797a ) or ( a9722a );
 a9726a <=( a793a ) or ( a794a );
 a9729a <=( a791a ) or ( a792a );
 a9730a <=( a9729a ) or ( a9726a );
 a9731a <=( a9730a ) or ( a9723a );
 a9734a <=( a789a ) or ( a790a );
 a9737a <=( a787a ) or ( a788a );
 a9738a <=( a9737a ) or ( a9734a );
 a9741a <=( a785a ) or ( a786a );
 a9744a <=( a783a ) or ( a784a );
 a9745a <=( a9744a ) or ( a9741a );
 a9746a <=( a9745a ) or ( a9738a );
 a9747a <=( a9746a ) or ( a9731a );
 a9751a <=( a780a ) or ( a781a );
 a9752a <=( a782a ) or ( a9751a );
 a9755a <=( a778a ) or ( a779a );
 a9758a <=( a776a ) or ( a777a );
 a9759a <=( a9758a ) or ( a9755a );
 a9760a <=( a9759a ) or ( a9752a );
 a9763a <=( a774a ) or ( a775a );
 a9766a <=( a772a ) or ( a773a );
 a9767a <=( a9766a ) or ( a9763a );
 a9770a <=( a770a ) or ( a771a );
 a9773a <=( a768a ) or ( a769a );
 a9774a <=( a9773a ) or ( a9770a );
 a9775a <=( a9774a ) or ( a9767a );
 a9776a <=( a9775a ) or ( a9760a );
 a9777a <=( a9776a ) or ( a9747a );
 a9778a <=( a9777a ) or ( a9718a );
 a9782a <=( a765a ) or ( a766a );
 a9783a <=( a767a ) or ( a9782a );
 a9786a <=( a763a ) or ( a764a );
 a9789a <=( a761a ) or ( a762a );
 a9790a <=( a9789a ) or ( a9786a );
 a9791a <=( a9790a ) or ( a9783a );
 a9795a <=( a758a ) or ( a759a );
 a9796a <=( a760a ) or ( a9795a );
 a9799a <=( a756a ) or ( a757a );
 a9802a <=( a754a ) or ( a755a );
 a9803a <=( a9802a ) or ( a9799a );
 a9804a <=( a9803a ) or ( a9796a );
 a9805a <=( a9804a ) or ( a9791a );
 a9809a <=( a751a ) or ( a752a );
 a9810a <=( a753a ) or ( a9809a );
 a9813a <=( a749a ) or ( a750a );
 a9816a <=( a747a ) or ( a748a );
 a9817a <=( a9816a ) or ( a9813a );
 a9818a <=( a9817a ) or ( a9810a );
 a9821a <=( a745a ) or ( a746a );
 a9824a <=( a743a ) or ( a744a );
 a9825a <=( a9824a ) or ( a9821a );
 a9828a <=( a741a ) or ( a742a );
 a9831a <=( a739a ) or ( a740a );
 a9832a <=( a9831a ) or ( a9828a );
 a9833a <=( a9832a ) or ( a9825a );
 a9834a <=( a9833a ) or ( a9818a );
 a9835a <=( a9834a ) or ( a9805a );
 a9839a <=( a736a ) or ( a737a );
 a9840a <=( a738a ) or ( a9839a );
 a9843a <=( a734a ) or ( a735a );
 a9846a <=( a732a ) or ( a733a );
 a9847a <=( a9846a ) or ( a9843a );
 a9848a <=( a9847a ) or ( a9840a );
 a9851a <=( a730a ) or ( a731a );
 a9854a <=( a728a ) or ( a729a );
 a9855a <=( a9854a ) or ( a9851a );
 a9858a <=( a726a ) or ( a727a );
 a9861a <=( a724a ) or ( a725a );
 a9862a <=( a9861a ) or ( a9858a );
 a9863a <=( a9862a ) or ( a9855a );
 a9864a <=( a9863a ) or ( a9848a );
 a9868a <=( a721a ) or ( a722a );
 a9869a <=( a723a ) or ( a9868a );
 a9872a <=( a719a ) or ( a720a );
 a9875a <=( a717a ) or ( a718a );
 a9876a <=( a9875a ) or ( a9872a );
 a9877a <=( a9876a ) or ( a9869a );
 a9880a <=( a715a ) or ( a716a );
 a9883a <=( a713a ) or ( a714a );
 a9884a <=( a9883a ) or ( a9880a );
 a9887a <=( a711a ) or ( a712a );
 a9890a <=( a709a ) or ( a710a );
 a9891a <=( a9890a ) or ( a9887a );
 a9892a <=( a9891a ) or ( a9884a );
 a9893a <=( a9892a ) or ( a9877a );
 a9894a <=( a9893a ) or ( a9864a );
 a9895a <=( a9894a ) or ( a9835a );
 a9896a <=( a9895a ) or ( a9778a );
 a9897a <=( a9896a ) or ( a9661a );
 a9901a <=( a706a ) or ( a707a );
 a9902a <=( a708a ) or ( a9901a );
 a9905a <=( a704a ) or ( a705a );
 a9908a <=( a702a ) or ( a703a );
 a9909a <=( a9908a ) or ( a9905a );
 a9910a <=( a9909a ) or ( a9902a );
 a9914a <=( a699a ) or ( a700a );
 a9915a <=( a701a ) or ( a9914a );
 a9918a <=( a697a ) or ( a698a );
 a9921a <=( a695a ) or ( a696a );
 a9922a <=( a9921a ) or ( a9918a );
 a9923a <=( a9922a ) or ( a9915a );
 a9924a <=( a9923a ) or ( a9910a );
 a9928a <=( a692a ) or ( a693a );
 a9929a <=( a694a ) or ( a9928a );
 a9932a <=( a690a ) or ( a691a );
 a9935a <=( a688a ) or ( a689a );
 a9936a <=( a9935a ) or ( a9932a );
 a9937a <=( a9936a ) or ( a9929a );
 a9940a <=( a686a ) or ( a687a );
 a9943a <=( a684a ) or ( a685a );
 a9944a <=( a9943a ) or ( a9940a );
 a9947a <=( a682a ) or ( a683a );
 a9950a <=( a680a ) or ( a681a );
 a9951a <=( a9950a ) or ( a9947a );
 a9952a <=( a9951a ) or ( a9944a );
 a9953a <=( a9952a ) or ( a9937a );
 a9954a <=( a9953a ) or ( a9924a );
 a9958a <=( a677a ) or ( a678a );
 a9959a <=( a679a ) or ( a9958a );
 a9962a <=( a675a ) or ( a676a );
 a9965a <=( a673a ) or ( a674a );
 a9966a <=( a9965a ) or ( a9962a );
 a9967a <=( a9966a ) or ( a9959a );
 a9970a <=( a671a ) or ( a672a );
 a9973a <=( a669a ) or ( a670a );
 a9974a <=( a9973a ) or ( a9970a );
 a9977a <=( a667a ) or ( a668a );
 a9980a <=( a665a ) or ( a666a );
 a9981a <=( a9980a ) or ( a9977a );
 a9982a <=( a9981a ) or ( a9974a );
 a9983a <=( a9982a ) or ( a9967a );
 a9987a <=( a662a ) or ( a663a );
 a9988a <=( a664a ) or ( a9987a );
 a9991a <=( a660a ) or ( a661a );
 a9994a <=( a658a ) or ( a659a );
 a9995a <=( a9994a ) or ( a9991a );
 a9996a <=( a9995a ) or ( a9988a );
 a9999a <=( a656a ) or ( a657a );
 a10002a <=( a654a ) or ( a655a );
 a10003a <=( a10002a ) or ( a9999a );
 a10006a <=( a652a ) or ( a653a );
 a10009a <=( a650a ) or ( a651a );
 a10010a <=( a10009a ) or ( a10006a );
 a10011a <=( a10010a ) or ( a10003a );
 a10012a <=( a10011a ) or ( a9996a );
 a10013a <=( a10012a ) or ( a9983a );
 a10014a <=( a10013a ) or ( a9954a );
 a10018a <=( a647a ) or ( a648a );
 a10019a <=( a649a ) or ( a10018a );
 a10022a <=( a645a ) or ( a646a );
 a10025a <=( a643a ) or ( a644a );
 a10026a <=( a10025a ) or ( a10022a );
 a10027a <=( a10026a ) or ( a10019a );
 a10031a <=( a640a ) or ( a641a );
 a10032a <=( a642a ) or ( a10031a );
 a10035a <=( a638a ) or ( a639a );
 a10038a <=( a636a ) or ( a637a );
 a10039a <=( a10038a ) or ( a10035a );
 a10040a <=( a10039a ) or ( a10032a );
 a10041a <=( a10040a ) or ( a10027a );
 a10045a <=( a633a ) or ( a634a );
 a10046a <=( a635a ) or ( a10045a );
 a10049a <=( a631a ) or ( a632a );
 a10052a <=( a629a ) or ( a630a );
 a10053a <=( a10052a ) or ( a10049a );
 a10054a <=( a10053a ) or ( a10046a );
 a10057a <=( a627a ) or ( a628a );
 a10060a <=( a625a ) or ( a626a );
 a10061a <=( a10060a ) or ( a10057a );
 a10064a <=( a623a ) or ( a624a );
 a10067a <=( a621a ) or ( a622a );
 a10068a <=( a10067a ) or ( a10064a );
 a10069a <=( a10068a ) or ( a10061a );
 a10070a <=( a10069a ) or ( a10054a );
 a10071a <=( a10070a ) or ( a10041a );
 a10075a <=( a618a ) or ( a619a );
 a10076a <=( a620a ) or ( a10075a );
 a10079a <=( a616a ) or ( a617a );
 a10082a <=( a614a ) or ( a615a );
 a10083a <=( a10082a ) or ( a10079a );
 a10084a <=( a10083a ) or ( a10076a );
 a10087a <=( a612a ) or ( a613a );
 a10090a <=( a610a ) or ( a611a );
 a10091a <=( a10090a ) or ( a10087a );
 a10094a <=( a608a ) or ( a609a );
 a10097a <=( a606a ) or ( a607a );
 a10098a <=( a10097a ) or ( a10094a );
 a10099a <=( a10098a ) or ( a10091a );
 a10100a <=( a10099a ) or ( a10084a );
 a10104a <=( a603a ) or ( a604a );
 a10105a <=( a605a ) or ( a10104a );
 a10108a <=( a601a ) or ( a602a );
 a10111a <=( a599a ) or ( a600a );
 a10112a <=( a10111a ) or ( a10108a );
 a10113a <=( a10112a ) or ( a10105a );
 a10116a <=( a597a ) or ( a598a );
 a10119a <=( a595a ) or ( a596a );
 a10120a <=( a10119a ) or ( a10116a );
 a10123a <=( a593a ) or ( a594a );
 a10126a <=( a591a ) or ( a592a );
 a10127a <=( a10126a ) or ( a10123a );
 a10128a <=( a10127a ) or ( a10120a );
 a10129a <=( a10128a ) or ( a10113a );
 a10130a <=( a10129a ) or ( a10100a );
 a10131a <=( a10130a ) or ( a10071a );
 a10132a <=( a10131a ) or ( a10014a );
 a10136a <=( a588a ) or ( a589a );
 a10137a <=( a590a ) or ( a10136a );
 a10140a <=( a586a ) or ( a587a );
 a10143a <=( a584a ) or ( a585a );
 a10144a <=( a10143a ) or ( a10140a );
 a10145a <=( a10144a ) or ( a10137a );
 a10149a <=( a581a ) or ( a582a );
 a10150a <=( a583a ) or ( a10149a );
 a10153a <=( a579a ) or ( a580a );
 a10156a <=( a577a ) or ( a578a );
 a10157a <=( a10156a ) or ( a10153a );
 a10158a <=( a10157a ) or ( a10150a );
 a10159a <=( a10158a ) or ( a10145a );
 a10163a <=( a574a ) or ( a575a );
 a10164a <=( a576a ) or ( a10163a );
 a10167a <=( a572a ) or ( a573a );
 a10170a <=( a570a ) or ( a571a );
 a10171a <=( a10170a ) or ( a10167a );
 a10172a <=( a10171a ) or ( a10164a );
 a10175a <=( a568a ) or ( a569a );
 a10178a <=( a566a ) or ( a567a );
 a10179a <=( a10178a ) or ( a10175a );
 a10182a <=( a564a ) or ( a565a );
 a10185a <=( a562a ) or ( a563a );
 a10186a <=( a10185a ) or ( a10182a );
 a10187a <=( a10186a ) or ( a10179a );
 a10188a <=( a10187a ) or ( a10172a );
 a10189a <=( a10188a ) or ( a10159a );
 a10193a <=( a559a ) or ( a560a );
 a10194a <=( a561a ) or ( a10193a );
 a10197a <=( a557a ) or ( a558a );
 a10200a <=( a555a ) or ( a556a );
 a10201a <=( a10200a ) or ( a10197a );
 a10202a <=( a10201a ) or ( a10194a );
 a10205a <=( a553a ) or ( a554a );
 a10208a <=( a551a ) or ( a552a );
 a10209a <=( a10208a ) or ( a10205a );
 a10212a <=( a549a ) or ( a550a );
 a10215a <=( a547a ) or ( a548a );
 a10216a <=( a10215a ) or ( a10212a );
 a10217a <=( a10216a ) or ( a10209a );
 a10218a <=( a10217a ) or ( a10202a );
 a10222a <=( a544a ) or ( a545a );
 a10223a <=( a546a ) or ( a10222a );
 a10226a <=( a542a ) or ( a543a );
 a10229a <=( a540a ) or ( a541a );
 a10230a <=( a10229a ) or ( a10226a );
 a10231a <=( a10230a ) or ( a10223a );
 a10234a <=( a538a ) or ( a539a );
 a10237a <=( a536a ) or ( a537a );
 a10238a <=( a10237a ) or ( a10234a );
 a10241a <=( a534a ) or ( a535a );
 a10244a <=( a532a ) or ( a533a );
 a10245a <=( a10244a ) or ( a10241a );
 a10246a <=( a10245a ) or ( a10238a );
 a10247a <=( a10246a ) or ( a10231a );
 a10248a <=( a10247a ) or ( a10218a );
 a10249a <=( a10248a ) or ( a10189a );
 a10253a <=( a529a ) or ( a530a );
 a10254a <=( a531a ) or ( a10253a );
 a10257a <=( a527a ) or ( a528a );
 a10260a <=( a525a ) or ( a526a );
 a10261a <=( a10260a ) or ( a10257a );
 a10262a <=( a10261a ) or ( a10254a );
 a10266a <=( a522a ) or ( a523a );
 a10267a <=( a524a ) or ( a10266a );
 a10270a <=( a520a ) or ( a521a );
 a10273a <=( a518a ) or ( a519a );
 a10274a <=( a10273a ) or ( a10270a );
 a10275a <=( a10274a ) or ( a10267a );
 a10276a <=( a10275a ) or ( a10262a );
 a10280a <=( a515a ) or ( a516a );
 a10281a <=( a517a ) or ( a10280a );
 a10284a <=( a513a ) or ( a514a );
 a10287a <=( a511a ) or ( a512a );
 a10288a <=( a10287a ) or ( a10284a );
 a10289a <=( a10288a ) or ( a10281a );
 a10292a <=( a509a ) or ( a510a );
 a10295a <=( a507a ) or ( a508a );
 a10296a <=( a10295a ) or ( a10292a );
 a10299a <=( a505a ) or ( a506a );
 a10302a <=( a503a ) or ( a504a );
 a10303a <=( a10302a ) or ( a10299a );
 a10304a <=( a10303a ) or ( a10296a );
 a10305a <=( a10304a ) or ( a10289a );
 a10306a <=( a10305a ) or ( a10276a );
 a10310a <=( a500a ) or ( a501a );
 a10311a <=( a502a ) or ( a10310a );
 a10314a <=( a498a ) or ( a499a );
 a10317a <=( a496a ) or ( a497a );
 a10318a <=( a10317a ) or ( a10314a );
 a10319a <=( a10318a ) or ( a10311a );
 a10322a <=( a494a ) or ( a495a );
 a10325a <=( a492a ) or ( a493a );
 a10326a <=( a10325a ) or ( a10322a );
 a10329a <=( a490a ) or ( a491a );
 a10332a <=( a488a ) or ( a489a );
 a10333a <=( a10332a ) or ( a10329a );
 a10334a <=( a10333a ) or ( a10326a );
 a10335a <=( a10334a ) or ( a10319a );
 a10339a <=( a485a ) or ( a486a );
 a10340a <=( a487a ) or ( a10339a );
 a10343a <=( a483a ) or ( a484a );
 a10346a <=( a481a ) or ( a482a );
 a10347a <=( a10346a ) or ( a10343a );
 a10348a <=( a10347a ) or ( a10340a );
 a10351a <=( a479a ) or ( a480a );
 a10354a <=( a477a ) or ( a478a );
 a10355a <=( a10354a ) or ( a10351a );
 a10358a <=( a475a ) or ( a476a );
 a10361a <=( a473a ) or ( a474a );
 a10362a <=( a10361a ) or ( a10358a );
 a10363a <=( a10362a ) or ( a10355a );
 a10364a <=( a10363a ) or ( a10348a );
 a10365a <=( a10364a ) or ( a10335a );
 a10366a <=( a10365a ) or ( a10306a );
 a10367a <=( a10366a ) or ( a10249a );
 a10368a <=( a10367a ) or ( a10132a );
 a10369a <=( a10368a ) or ( a9897a );
 a10373a <=( a470a ) or ( a471a );
 a10374a <=( a472a ) or ( a10373a );
 a10377a <=( a468a ) or ( a469a );
 a10380a <=( a466a ) or ( a467a );
 a10381a <=( a10380a ) or ( a10377a );
 a10382a <=( a10381a ) or ( a10374a );
 a10386a <=( a463a ) or ( a464a );
 a10387a <=( a465a ) or ( a10386a );
 a10390a <=( a461a ) or ( a462a );
 a10393a <=( a459a ) or ( a460a );
 a10394a <=( a10393a ) or ( a10390a );
 a10395a <=( a10394a ) or ( a10387a );
 a10396a <=( a10395a ) or ( a10382a );
 a10400a <=( a456a ) or ( a457a );
 a10401a <=( a458a ) or ( a10400a );
 a10404a <=( a454a ) or ( a455a );
 a10407a <=( a452a ) or ( a453a );
 a10408a <=( a10407a ) or ( a10404a );
 a10409a <=( a10408a ) or ( a10401a );
 a10412a <=( a450a ) or ( a451a );
 a10415a <=( a448a ) or ( a449a );
 a10416a <=( a10415a ) or ( a10412a );
 a10419a <=( a446a ) or ( a447a );
 a10422a <=( a444a ) or ( a445a );
 a10423a <=( a10422a ) or ( a10419a );
 a10424a <=( a10423a ) or ( a10416a );
 a10425a <=( a10424a ) or ( a10409a );
 a10426a <=( a10425a ) or ( a10396a );
 a10430a <=( a441a ) or ( a442a );
 a10431a <=( a443a ) or ( a10430a );
 a10434a <=( a439a ) or ( a440a );
 a10437a <=( a437a ) or ( a438a );
 a10438a <=( a10437a ) or ( a10434a );
 a10439a <=( a10438a ) or ( a10431a );
 a10442a <=( a435a ) or ( a436a );
 a10445a <=( a433a ) or ( a434a );
 a10446a <=( a10445a ) or ( a10442a );
 a10449a <=( a431a ) or ( a432a );
 a10452a <=( a429a ) or ( a430a );
 a10453a <=( a10452a ) or ( a10449a );
 a10454a <=( a10453a ) or ( a10446a );
 a10455a <=( a10454a ) or ( a10439a );
 a10459a <=( a426a ) or ( a427a );
 a10460a <=( a428a ) or ( a10459a );
 a10463a <=( a424a ) or ( a425a );
 a10466a <=( a422a ) or ( a423a );
 a10467a <=( a10466a ) or ( a10463a );
 a10468a <=( a10467a ) or ( a10460a );
 a10471a <=( a420a ) or ( a421a );
 a10474a <=( a418a ) or ( a419a );
 a10475a <=( a10474a ) or ( a10471a );
 a10478a <=( a416a ) or ( a417a );
 a10481a <=( a414a ) or ( a415a );
 a10482a <=( a10481a ) or ( a10478a );
 a10483a <=( a10482a ) or ( a10475a );
 a10484a <=( a10483a ) or ( a10468a );
 a10485a <=( a10484a ) or ( a10455a );
 a10486a <=( a10485a ) or ( a10426a );
 a10490a <=( a411a ) or ( a412a );
 a10491a <=( a413a ) or ( a10490a );
 a10494a <=( a409a ) or ( a410a );
 a10497a <=( a407a ) or ( a408a );
 a10498a <=( a10497a ) or ( a10494a );
 a10499a <=( a10498a ) or ( a10491a );
 a10503a <=( a404a ) or ( a405a );
 a10504a <=( a406a ) or ( a10503a );
 a10507a <=( a402a ) or ( a403a );
 a10510a <=( a400a ) or ( a401a );
 a10511a <=( a10510a ) or ( a10507a );
 a10512a <=( a10511a ) or ( a10504a );
 a10513a <=( a10512a ) or ( a10499a );
 a10517a <=( a397a ) or ( a398a );
 a10518a <=( a399a ) or ( a10517a );
 a10521a <=( a395a ) or ( a396a );
 a10524a <=( a393a ) or ( a394a );
 a10525a <=( a10524a ) or ( a10521a );
 a10526a <=( a10525a ) or ( a10518a );
 a10529a <=( a391a ) or ( a392a );
 a10532a <=( a389a ) or ( a390a );
 a10533a <=( a10532a ) or ( a10529a );
 a10536a <=( a387a ) or ( a388a );
 a10539a <=( a385a ) or ( a386a );
 a10540a <=( a10539a ) or ( a10536a );
 a10541a <=( a10540a ) or ( a10533a );
 a10542a <=( a10541a ) or ( a10526a );
 a10543a <=( a10542a ) or ( a10513a );
 a10547a <=( a382a ) or ( a383a );
 a10548a <=( a384a ) or ( a10547a );
 a10551a <=( a380a ) or ( a381a );
 a10554a <=( a378a ) or ( a379a );
 a10555a <=( a10554a ) or ( a10551a );
 a10556a <=( a10555a ) or ( a10548a );
 a10559a <=( a376a ) or ( a377a );
 a10562a <=( a374a ) or ( a375a );
 a10563a <=( a10562a ) or ( a10559a );
 a10566a <=( a372a ) or ( a373a );
 a10569a <=( a370a ) or ( a371a );
 a10570a <=( a10569a ) or ( a10566a );
 a10571a <=( a10570a ) or ( a10563a );
 a10572a <=( a10571a ) or ( a10556a );
 a10576a <=( a367a ) or ( a368a );
 a10577a <=( a369a ) or ( a10576a );
 a10580a <=( a365a ) or ( a366a );
 a10583a <=( a363a ) or ( a364a );
 a10584a <=( a10583a ) or ( a10580a );
 a10585a <=( a10584a ) or ( a10577a );
 a10588a <=( a361a ) or ( a362a );
 a10591a <=( a359a ) or ( a360a );
 a10592a <=( a10591a ) or ( a10588a );
 a10595a <=( a357a ) or ( a358a );
 a10598a <=( a355a ) or ( a356a );
 a10599a <=( a10598a ) or ( a10595a );
 a10600a <=( a10599a ) or ( a10592a );
 a10601a <=( a10600a ) or ( a10585a );
 a10602a <=( a10601a ) or ( a10572a );
 a10603a <=( a10602a ) or ( a10543a );
 a10604a <=( a10603a ) or ( a10486a );
 a10608a <=( a352a ) or ( a353a );
 a10609a <=( a354a ) or ( a10608a );
 a10612a <=( a350a ) or ( a351a );
 a10615a <=( a348a ) or ( a349a );
 a10616a <=( a10615a ) or ( a10612a );
 a10617a <=( a10616a ) or ( a10609a );
 a10621a <=( a345a ) or ( a346a );
 a10622a <=( a347a ) or ( a10621a );
 a10625a <=( a343a ) or ( a344a );
 a10628a <=( a341a ) or ( a342a );
 a10629a <=( a10628a ) or ( a10625a );
 a10630a <=( a10629a ) or ( a10622a );
 a10631a <=( a10630a ) or ( a10617a );
 a10635a <=( a338a ) or ( a339a );
 a10636a <=( a340a ) or ( a10635a );
 a10639a <=( a336a ) or ( a337a );
 a10642a <=( a334a ) or ( a335a );
 a10643a <=( a10642a ) or ( a10639a );
 a10644a <=( a10643a ) or ( a10636a );
 a10647a <=( a332a ) or ( a333a );
 a10650a <=( a330a ) or ( a331a );
 a10651a <=( a10650a ) or ( a10647a );
 a10654a <=( a328a ) or ( a329a );
 a10657a <=( a326a ) or ( a327a );
 a10658a <=( a10657a ) or ( a10654a );
 a10659a <=( a10658a ) or ( a10651a );
 a10660a <=( a10659a ) or ( a10644a );
 a10661a <=( a10660a ) or ( a10631a );
 a10665a <=( a323a ) or ( a324a );
 a10666a <=( a325a ) or ( a10665a );
 a10669a <=( a321a ) or ( a322a );
 a10672a <=( a319a ) or ( a320a );
 a10673a <=( a10672a ) or ( a10669a );
 a10674a <=( a10673a ) or ( a10666a );
 a10677a <=( a317a ) or ( a318a );
 a10680a <=( a315a ) or ( a316a );
 a10681a <=( a10680a ) or ( a10677a );
 a10684a <=( a313a ) or ( a314a );
 a10687a <=( a311a ) or ( a312a );
 a10688a <=( a10687a ) or ( a10684a );
 a10689a <=( a10688a ) or ( a10681a );
 a10690a <=( a10689a ) or ( a10674a );
 a10694a <=( a308a ) or ( a309a );
 a10695a <=( a310a ) or ( a10694a );
 a10698a <=( a306a ) or ( a307a );
 a10701a <=( a304a ) or ( a305a );
 a10702a <=( a10701a ) or ( a10698a );
 a10703a <=( a10702a ) or ( a10695a );
 a10706a <=( a302a ) or ( a303a );
 a10709a <=( a300a ) or ( a301a );
 a10710a <=( a10709a ) or ( a10706a );
 a10713a <=( a298a ) or ( a299a );
 a10716a <=( a296a ) or ( a297a );
 a10717a <=( a10716a ) or ( a10713a );
 a10718a <=( a10717a ) or ( a10710a );
 a10719a <=( a10718a ) or ( a10703a );
 a10720a <=( a10719a ) or ( a10690a );
 a10721a <=( a10720a ) or ( a10661a );
 a10725a <=( a293a ) or ( a294a );
 a10726a <=( a295a ) or ( a10725a );
 a10729a <=( a291a ) or ( a292a );
 a10732a <=( a289a ) or ( a290a );
 a10733a <=( a10732a ) or ( a10729a );
 a10734a <=( a10733a ) or ( a10726a );
 a10738a <=( a286a ) or ( a287a );
 a10739a <=( a288a ) or ( a10738a );
 a10742a <=( a284a ) or ( a285a );
 a10745a <=( a282a ) or ( a283a );
 a10746a <=( a10745a ) or ( a10742a );
 a10747a <=( a10746a ) or ( a10739a );
 a10748a <=( a10747a ) or ( a10734a );
 a10752a <=( a279a ) or ( a280a );
 a10753a <=( a281a ) or ( a10752a );
 a10756a <=( a277a ) or ( a278a );
 a10759a <=( a275a ) or ( a276a );
 a10760a <=( a10759a ) or ( a10756a );
 a10761a <=( a10760a ) or ( a10753a );
 a10764a <=( a273a ) or ( a274a );
 a10767a <=( a271a ) or ( a272a );
 a10768a <=( a10767a ) or ( a10764a );
 a10771a <=( a269a ) or ( a270a );
 a10774a <=( a267a ) or ( a268a );
 a10775a <=( a10774a ) or ( a10771a );
 a10776a <=( a10775a ) or ( a10768a );
 a10777a <=( a10776a ) or ( a10761a );
 a10778a <=( a10777a ) or ( a10748a );
 a10782a <=( a264a ) or ( a265a );
 a10783a <=( a266a ) or ( a10782a );
 a10786a <=( a262a ) or ( a263a );
 a10789a <=( a260a ) or ( a261a );
 a10790a <=( a10789a ) or ( a10786a );
 a10791a <=( a10790a ) or ( a10783a );
 a10794a <=( a258a ) or ( a259a );
 a10797a <=( a256a ) or ( a257a );
 a10798a <=( a10797a ) or ( a10794a );
 a10801a <=( a254a ) or ( a255a );
 a10804a <=( a252a ) or ( a253a );
 a10805a <=( a10804a ) or ( a10801a );
 a10806a <=( a10805a ) or ( a10798a );
 a10807a <=( a10806a ) or ( a10791a );
 a10811a <=( a249a ) or ( a250a );
 a10812a <=( a251a ) or ( a10811a );
 a10815a <=( a247a ) or ( a248a );
 a10818a <=( a245a ) or ( a246a );
 a10819a <=( a10818a ) or ( a10815a );
 a10820a <=( a10819a ) or ( a10812a );
 a10823a <=( a243a ) or ( a244a );
 a10826a <=( a241a ) or ( a242a );
 a10827a <=( a10826a ) or ( a10823a );
 a10830a <=( a239a ) or ( a240a );
 a10833a <=( a237a ) or ( a238a );
 a10834a <=( a10833a ) or ( a10830a );
 a10835a <=( a10834a ) or ( a10827a );
 a10836a <=( a10835a ) or ( a10820a );
 a10837a <=( a10836a ) or ( a10807a );
 a10838a <=( a10837a ) or ( a10778a );
 a10839a <=( a10838a ) or ( a10721a );
 a10840a <=( a10839a ) or ( a10604a );
 a10844a <=( a234a ) or ( a235a );
 a10845a <=( a236a ) or ( a10844a );
 a10848a <=( a232a ) or ( a233a );
 a10851a <=( a230a ) or ( a231a );
 a10852a <=( a10851a ) or ( a10848a );
 a10853a <=( a10852a ) or ( a10845a );
 a10857a <=( a227a ) or ( a228a );
 a10858a <=( a229a ) or ( a10857a );
 a10861a <=( a225a ) or ( a226a );
 a10864a <=( a223a ) or ( a224a );
 a10865a <=( a10864a ) or ( a10861a );
 a10866a <=( a10865a ) or ( a10858a );
 a10867a <=( a10866a ) or ( a10853a );
 a10871a <=( a220a ) or ( a221a );
 a10872a <=( a222a ) or ( a10871a );
 a10875a <=( a218a ) or ( a219a );
 a10878a <=( a216a ) or ( a217a );
 a10879a <=( a10878a ) or ( a10875a );
 a10880a <=( a10879a ) or ( a10872a );
 a10883a <=( a214a ) or ( a215a );
 a10886a <=( a212a ) or ( a213a );
 a10887a <=( a10886a ) or ( a10883a );
 a10890a <=( a210a ) or ( a211a );
 a10893a <=( a208a ) or ( a209a );
 a10894a <=( a10893a ) or ( a10890a );
 a10895a <=( a10894a ) or ( a10887a );
 a10896a <=( a10895a ) or ( a10880a );
 a10897a <=( a10896a ) or ( a10867a );
 a10901a <=( a205a ) or ( a206a );
 a10902a <=( a207a ) or ( a10901a );
 a10905a <=( a203a ) or ( a204a );
 a10908a <=( a201a ) or ( a202a );
 a10909a <=( a10908a ) or ( a10905a );
 a10910a <=( a10909a ) or ( a10902a );
 a10913a <=( a199a ) or ( a200a );
 a10916a <=( a197a ) or ( a198a );
 a10917a <=( a10916a ) or ( a10913a );
 a10920a <=( a195a ) or ( a196a );
 a10923a <=( a193a ) or ( a194a );
 a10924a <=( a10923a ) or ( a10920a );
 a10925a <=( a10924a ) or ( a10917a );
 a10926a <=( a10925a ) or ( a10910a );
 a10930a <=( a190a ) or ( a191a );
 a10931a <=( a192a ) or ( a10930a );
 a10934a <=( a188a ) or ( a189a );
 a10937a <=( a186a ) or ( a187a );
 a10938a <=( a10937a ) or ( a10934a );
 a10939a <=( a10938a ) or ( a10931a );
 a10942a <=( a184a ) or ( a185a );
 a10945a <=( a182a ) or ( a183a );
 a10946a <=( a10945a ) or ( a10942a );
 a10949a <=( a180a ) or ( a181a );
 a10952a <=( a178a ) or ( a179a );
 a10953a <=( a10952a ) or ( a10949a );
 a10954a <=( a10953a ) or ( a10946a );
 a10955a <=( a10954a ) or ( a10939a );
 a10956a <=( a10955a ) or ( a10926a );
 a10957a <=( a10956a ) or ( a10897a );
 a10961a <=( a175a ) or ( a176a );
 a10962a <=( a177a ) or ( a10961a );
 a10965a <=( a173a ) or ( a174a );
 a10968a <=( a171a ) or ( a172a );
 a10969a <=( a10968a ) or ( a10965a );
 a10970a <=( a10969a ) or ( a10962a );
 a10974a <=( a168a ) or ( a169a );
 a10975a <=( a170a ) or ( a10974a );
 a10978a <=( a166a ) or ( a167a );
 a10981a <=( a164a ) or ( a165a );
 a10982a <=( a10981a ) or ( a10978a );
 a10983a <=( a10982a ) or ( a10975a );
 a10984a <=( a10983a ) or ( a10970a );
 a10988a <=( a161a ) or ( a162a );
 a10989a <=( a163a ) or ( a10988a );
 a10992a <=( a159a ) or ( a160a );
 a10995a <=( a157a ) or ( a158a );
 a10996a <=( a10995a ) or ( a10992a );
 a10997a <=( a10996a ) or ( a10989a );
 a11000a <=( a155a ) or ( a156a );
 a11003a <=( a153a ) or ( a154a );
 a11004a <=( a11003a ) or ( a11000a );
 a11007a <=( a151a ) or ( a152a );
 a11010a <=( a149a ) or ( a150a );
 a11011a <=( a11010a ) or ( a11007a );
 a11012a <=( a11011a ) or ( a11004a );
 a11013a <=( a11012a ) or ( a10997a );
 a11014a <=( a11013a ) or ( a10984a );
 a11018a <=( a146a ) or ( a147a );
 a11019a <=( a148a ) or ( a11018a );
 a11022a <=( a144a ) or ( a145a );
 a11025a <=( a142a ) or ( a143a );
 a11026a <=( a11025a ) or ( a11022a );
 a11027a <=( a11026a ) or ( a11019a );
 a11030a <=( a140a ) or ( a141a );
 a11033a <=( a138a ) or ( a139a );
 a11034a <=( a11033a ) or ( a11030a );
 a11037a <=( a136a ) or ( a137a );
 a11040a <=( a134a ) or ( a135a );
 a11041a <=( a11040a ) or ( a11037a );
 a11042a <=( a11041a ) or ( a11034a );
 a11043a <=( a11042a ) or ( a11027a );
 a11047a <=( a131a ) or ( a132a );
 a11048a <=( a133a ) or ( a11047a );
 a11051a <=( a129a ) or ( a130a );
 a11054a <=( a127a ) or ( a128a );
 a11055a <=( a11054a ) or ( a11051a );
 a11056a <=( a11055a ) or ( a11048a );
 a11059a <=( a125a ) or ( a126a );
 a11062a <=( a123a ) or ( a124a );
 a11063a <=( a11062a ) or ( a11059a );
 a11066a <=( a121a ) or ( a122a );
 a11069a <=( a119a ) or ( a120a );
 a11070a <=( a11069a ) or ( a11066a );
 a11071a <=( a11070a ) or ( a11063a );
 a11072a <=( a11071a ) or ( a11056a );
 a11073a <=( a11072a ) or ( a11043a );
 a11074a <=( a11073a ) or ( a11014a );
 a11075a <=( a11074a ) or ( a10957a );
 a11079a <=( a116a ) or ( a117a );
 a11080a <=( a118a ) or ( a11079a );
 a11083a <=( a114a ) or ( a115a );
 a11086a <=( a112a ) or ( a113a );
 a11087a <=( a11086a ) or ( a11083a );
 a11088a <=( a11087a ) or ( a11080a );
 a11092a <=( a109a ) or ( a110a );
 a11093a <=( a111a ) or ( a11092a );
 a11096a <=( a107a ) or ( a108a );
 a11099a <=( a105a ) or ( a106a );
 a11100a <=( a11099a ) or ( a11096a );
 a11101a <=( a11100a ) or ( a11093a );
 a11102a <=( a11101a ) or ( a11088a );
 a11106a <=( a102a ) or ( a103a );
 a11107a <=( a104a ) or ( a11106a );
 a11110a <=( a100a ) or ( a101a );
 a11113a <=( a98a ) or ( a99a );
 a11114a <=( a11113a ) or ( a11110a );
 a11115a <=( a11114a ) or ( a11107a );
 a11118a <=( a96a ) or ( a97a );
 a11121a <=( a94a ) or ( a95a );
 a11122a <=( a11121a ) or ( a11118a );
 a11125a <=( a92a ) or ( a93a );
 a11128a <=( a90a ) or ( a91a );
 a11129a <=( a11128a ) or ( a11125a );
 a11130a <=( a11129a ) or ( a11122a );
 a11131a <=( a11130a ) or ( a11115a );
 a11132a <=( a11131a ) or ( a11102a );
 a11136a <=( a87a ) or ( a88a );
 a11137a <=( a89a ) or ( a11136a );
 a11140a <=( a85a ) or ( a86a );
 a11143a <=( a83a ) or ( a84a );
 a11144a <=( a11143a ) or ( a11140a );
 a11145a <=( a11144a ) or ( a11137a );
 a11148a <=( a81a ) or ( a82a );
 a11151a <=( a79a ) or ( a80a );
 a11152a <=( a11151a ) or ( a11148a );
 a11155a <=( a77a ) or ( a78a );
 a11158a <=( a75a ) or ( a76a );
 a11159a <=( a11158a ) or ( a11155a );
 a11160a <=( a11159a ) or ( a11152a );
 a11161a <=( a11160a ) or ( a11145a );
 a11165a <=( a72a ) or ( a73a );
 a11166a <=( a74a ) or ( a11165a );
 a11169a <=( a70a ) or ( a71a );
 a11172a <=( a68a ) or ( a69a );
 a11173a <=( a11172a ) or ( a11169a );
 a11174a <=( a11173a ) or ( a11166a );
 a11177a <=( a66a ) or ( a67a );
 a11180a <=( a64a ) or ( a65a );
 a11181a <=( a11180a ) or ( a11177a );
 a11184a <=( a62a ) or ( a63a );
 a11187a <=( a60a ) or ( a61a );
 a11188a <=( a11187a ) or ( a11184a );
 a11189a <=( a11188a ) or ( a11181a );
 a11190a <=( a11189a ) or ( a11174a );
 a11191a <=( a11190a ) or ( a11161a );
 a11192a <=( a11191a ) or ( a11132a );
 a11196a <=( a57a ) or ( a58a );
 a11197a <=( a59a ) or ( a11196a );
 a11200a <=( a55a ) or ( a56a );
 a11203a <=( a53a ) or ( a54a );
 a11204a <=( a11203a ) or ( a11200a );
 a11205a <=( a11204a ) or ( a11197a );
 a11209a <=( a50a ) or ( a51a );
 a11210a <=( a52a ) or ( a11209a );
 a11213a <=( a48a ) or ( a49a );
 a11216a <=( a46a ) or ( a47a );
 a11217a <=( a11216a ) or ( a11213a );
 a11218a <=( a11217a ) or ( a11210a );
 a11219a <=( a11218a ) or ( a11205a );
 a11223a <=( a43a ) or ( a44a );
 a11224a <=( a45a ) or ( a11223a );
 a11227a <=( a41a ) or ( a42a );
 a11230a <=( a39a ) or ( a40a );
 a11231a <=( a11230a ) or ( a11227a );
 a11232a <=( a11231a ) or ( a11224a );
 a11235a <=( a37a ) or ( a38a );
 a11238a <=( a35a ) or ( a36a );
 a11239a <=( a11238a ) or ( a11235a );
 a11242a <=( a33a ) or ( a34a );
 a11245a <=( a31a ) or ( a32a );
 a11246a <=( a11245a ) or ( a11242a );
 a11247a <=( a11246a ) or ( a11239a );
 a11248a <=( a11247a ) or ( a11232a );
 a11249a <=( a11248a ) or ( a11219a );
 a11253a <=( a28a ) or ( a29a );
 a11254a <=( a30a ) or ( a11253a );
 a11257a <=( a26a ) or ( a27a );
 a11260a <=( a24a ) or ( a25a );
 a11261a <=( a11260a ) or ( a11257a );
 a11262a <=( a11261a ) or ( a11254a );
 a11265a <=( a22a ) or ( a23a );
 a11268a <=( a20a ) or ( a21a );
 a11269a <=( a11268a ) or ( a11265a );
 a11272a <=( a18a ) or ( a19a );
 a11275a <=( a16a ) or ( a17a );
 a11276a <=( a11275a ) or ( a11272a );
 a11277a <=( a11276a ) or ( a11269a );
 a11278a <=( a11277a ) or ( a11262a );
 a11282a <=( a13a ) or ( a14a );
 a11283a <=( a15a ) or ( a11282a );
 a11286a <=( a11a ) or ( a12a );
 a11289a <=( a9a ) or ( a10a );
 a11290a <=( a11289a ) or ( a11286a );
 a11291a <=( a11290a ) or ( a11283a );
 a11294a <=( a7a ) or ( a8a );
 a11297a <=( a5a ) or ( a6a );
 a11298a <=( a11297a ) or ( a11294a );
 a11301a <=( a3a ) or ( a4a );
 a11304a <=( a1a ) or ( a2a );
 a11305a <=( a11304a ) or ( a11301a );
 a11306a <=( a11305a ) or ( a11298a );
 a11307a <=( a11306a ) or ( a11291a );
 a11308a <=( a11307a ) or ( a11278a );
 a11309a <=( a11308a ) or ( a11249a );
 a11310a <=( a11309a ) or ( a11192a );
 a11311a <=( a11310a ) or ( a11075a );
 a11312a <=( a11311a ) or ( a10840a );
 a11313a <=( a11312a ) or ( a10369a );
 a11314a <=( a11313a ) or ( a9428a );
 a11317a <=( A166  and  A168 );
 a11320a <=( A200  and  A199 );
 a11321a <=( a11320a  and  a11317a );
 a11324a <=( A233  and  (not A232) );
 a11327a <=( A299  and  (not A298) );
 a11328a <=( a11327a  and  a11324a );
 a11331a <=( A166  and  A168 );
 a11334a <=( A200  and  A199 );
 a11335a <=( a11334a  and  a11331a );
 a11338a <=( A233  and  (not A232) );
 a11341a <=( A266  and  (not A265) );
 a11342a <=( a11341a  and  a11338a );
 a11345a <=( A166  and  A168 );
 a11348a <=( (not A201)  and  (not A200) );
 a11349a <=( a11348a  and  a11345a );
 a11352a <=( A233  and  (not A232) );
 a11355a <=( A299  and  (not A298) );
 a11356a <=( a11355a  and  a11352a );
 a11359a <=( A166  and  A168 );
 a11362a <=( (not A201)  and  (not A200) );
 a11363a <=( a11362a  and  a11359a );
 a11366a <=( A233  and  (not A232) );
 a11369a <=( A266  and  (not A265) );
 a11370a <=( a11369a  and  a11366a );
 a11373a <=( A166  and  A168 );
 a11376a <=( (not A200)  and  (not A199) );
 a11377a <=( a11376a  and  a11373a );
 a11380a <=( A233  and  (not A232) );
 a11383a <=( A299  and  (not A298) );
 a11384a <=( a11383a  and  a11380a );
 a11387a <=( A166  and  A168 );
 a11390a <=( (not A200)  and  (not A199) );
 a11391a <=( a11390a  and  a11387a );
 a11394a <=( A233  and  (not A232) );
 a11397a <=( A266  and  (not A265) );
 a11398a <=( a11397a  and  a11394a );
 a11401a <=( A167  and  A168 );
 a11404a <=( A200  and  A199 );
 a11405a <=( a11404a  and  a11401a );
 a11408a <=( A233  and  (not A232) );
 a11411a <=( A299  and  (not A298) );
 a11412a <=( a11411a  and  a11408a );
 a11415a <=( A167  and  A168 );
 a11418a <=( A200  and  A199 );
 a11419a <=( a11418a  and  a11415a );
 a11422a <=( A233  and  (not A232) );
 a11425a <=( A266  and  (not A265) );
 a11426a <=( a11425a  and  a11422a );
 a11429a <=( A167  and  A168 );
 a11432a <=( (not A201)  and  (not A200) );
 a11433a <=( a11432a  and  a11429a );
 a11436a <=( A233  and  (not A232) );
 a11439a <=( A299  and  (not A298) );
 a11440a <=( a11439a  and  a11436a );
 a11443a <=( A167  and  A168 );
 a11446a <=( (not A201)  and  (not A200) );
 a11447a <=( a11446a  and  a11443a );
 a11450a <=( A233  and  (not A232) );
 a11453a <=( A266  and  (not A265) );
 a11454a <=( a11453a  and  a11450a );
 a11457a <=( A167  and  A168 );
 a11460a <=( (not A200)  and  (not A199) );
 a11461a <=( a11460a  and  a11457a );
 a11464a <=( A233  and  (not A232) );
 a11467a <=( A299  and  (not A298) );
 a11468a <=( a11467a  and  a11464a );
 a11471a <=( A167  and  A168 );
 a11474a <=( (not A200)  and  (not A199) );
 a11475a <=( a11474a  and  a11471a );
 a11478a <=( A233  and  (not A232) );
 a11481a <=( A266  and  (not A265) );
 a11482a <=( a11481a  and  a11478a );
 a11485a <=( A166  and  A168 );
 a11488a <=( (not A202)  and  (not A200) );
 a11489a <=( a11488a  and  a11485a );
 a11492a <=( (not A232)  and  (not A203) );
 a11496a <=( A299  and  (not A298) );
 a11497a <=( A233  and  a11496a );
 a11498a <=( a11497a  and  a11492a );
 a11501a <=( A166  and  A168 );
 a11504a <=( (not A202)  and  (not A200) );
 a11505a <=( a11504a  and  a11501a );
 a11508a <=( (not A232)  and  (not A203) );
 a11512a <=( A266  and  (not A265) );
 a11513a <=( A233  and  a11512a );
 a11514a <=( a11513a  and  a11508a );
 a11517a <=( A167  and  A168 );
 a11520a <=( (not A202)  and  (not A200) );
 a11521a <=( a11520a  and  a11517a );
 a11524a <=( (not A232)  and  (not A203) );
 a11528a <=( A299  and  (not A298) );
 a11529a <=( A233  and  a11528a );
 a11530a <=( a11529a  and  a11524a );
 a11533a <=( A167  and  A168 );
 a11536a <=( (not A202)  and  (not A200) );
 a11537a <=( a11536a  and  a11533a );
 a11540a <=( (not A232)  and  (not A203) );
 a11544a <=( A266  and  (not A265) );
 a11545a <=( A233  and  a11544a );
 a11546a <=( a11545a  and  a11540a );
 a11549a <=( (not A167)  and  A170 );
 a11552a <=( (not A199)  and  (not A166) );
 a11553a <=( a11552a  and  a11549a );
 a11556a <=( (not A232)  and  A200 );
 a11560a <=( A299  and  (not A298) );
 a11561a <=( A233  and  a11560a );
 a11562a <=( a11561a  and  a11556a );
 a11565a <=( (not A167)  and  A170 );
 a11568a <=( (not A199)  and  (not A166) );
 a11569a <=( a11568a  and  a11565a );
 a11572a <=( (not A232)  and  A200 );
 a11576a <=( A266  and  (not A265) );
 a11577a <=( A233  and  a11576a );
 a11578a <=( a11577a  and  a11572a );
 a11581a <=( (not A167)  and  (not A169) );
 a11584a <=( (not A199)  and  (not A166) );
 a11585a <=( a11584a  and  a11581a );
 a11588a <=( (not A232)  and  A200 );
 a11592a <=( A299  and  (not A298) );
 a11593a <=( A233  and  a11592a );
 a11594a <=( a11593a  and  a11588a );
 a11597a <=( (not A167)  and  (not A169) );
 a11600a <=( (not A199)  and  (not A166) );
 a11601a <=( a11600a  and  a11597a );
 a11604a <=( (not A232)  and  A200 );
 a11608a <=( A266  and  (not A265) );
 a11609a <=( A233  and  a11608a );
 a11610a <=( a11609a  and  a11604a );
 a11613a <=( A166  and  A168 );
 a11617a <=( A232  and  A200 );
 a11618a <=( A199  and  a11617a );
 a11619a <=( a11618a  and  a11613a );
 a11622a <=( A265  and  A233 );
 a11626a <=( (not A300)  and  (not A299) );
 a11627a <=( (not A267)  and  a11626a );
 a11628a <=( a11627a  and  a11622a );
 a11631a <=( A166  and  A168 );
 a11635a <=( A232  and  A200 );
 a11636a <=( A199  and  a11635a );
 a11637a <=( a11636a  and  a11631a );
 a11640a <=( A265  and  A233 );
 a11644a <=( A299  and  A298 );
 a11645a <=( (not A267)  and  a11644a );
 a11646a <=( a11645a  and  a11640a );
 a11649a <=( A166  and  A168 );
 a11653a <=( A232  and  A200 );
 a11654a <=( A199  and  a11653a );
 a11655a <=( a11654a  and  a11649a );
 a11658a <=( A265  and  A233 );
 a11662a <=( (not A299)  and  (not A298) );
 a11663a <=( (not A267)  and  a11662a );
 a11664a <=( a11663a  and  a11658a );
 a11667a <=( A166  and  A168 );
 a11671a <=( A232  and  A200 );
 a11672a <=( A199  and  a11671a );
 a11673a <=( a11672a  and  a11667a );
 a11676a <=( A265  and  A233 );
 a11680a <=( (not A300)  and  (not A299) );
 a11681a <=( A266  and  a11680a );
 a11682a <=( a11681a  and  a11676a );
 a11685a <=( A166  and  A168 );
 a11689a <=( A232  and  A200 );
 a11690a <=( A199  and  a11689a );
 a11691a <=( a11690a  and  a11685a );
 a11694a <=( A265  and  A233 );
 a11698a <=( A299  and  A298 );
 a11699a <=( A266  and  a11698a );
 a11700a <=( a11699a  and  a11694a );
 a11703a <=( A166  and  A168 );
 a11707a <=( A232  and  A200 );
 a11708a <=( A199  and  a11707a );
 a11709a <=( a11708a  and  a11703a );
 a11712a <=( A265  and  A233 );
 a11716a <=( (not A299)  and  (not A298) );
 a11717a <=( A266  and  a11716a );
 a11718a <=( a11717a  and  a11712a );
 a11721a <=( A166  and  A168 );
 a11725a <=( A232  and  A200 );
 a11726a <=( A199  and  a11725a );
 a11727a <=( a11726a  and  a11721a );
 a11730a <=( (not A265)  and  A233 );
 a11734a <=( (not A300)  and  (not A299) );
 a11735a <=( (not A266)  and  a11734a );
 a11736a <=( a11735a  and  a11730a );
 a11739a <=( A166  and  A168 );
 a11743a <=( A232  and  A200 );
 a11744a <=( A199  and  a11743a );
 a11745a <=( a11744a  and  a11739a );
 a11748a <=( (not A265)  and  A233 );
 a11752a <=( A299  and  A298 );
 a11753a <=( (not A266)  and  a11752a );
 a11754a <=( a11753a  and  a11748a );
 a11757a <=( A166  and  A168 );
 a11761a <=( A232  and  A200 );
 a11762a <=( A199  and  a11761a );
 a11763a <=( a11762a  and  a11757a );
 a11766a <=( (not A265)  and  A233 );
 a11770a <=( (not A299)  and  (not A298) );
 a11771a <=( (not A266)  and  a11770a );
 a11772a <=( a11771a  and  a11766a );
 a11775a <=( A166  and  A168 );
 a11779a <=( (not A232)  and  A200 );
 a11780a <=( A199  and  a11779a );
 a11781a <=( a11780a  and  a11775a );
 a11784a <=( A298  and  A233 );
 a11788a <=( A301  and  A300 );
 a11789a <=( (not A299)  and  a11788a );
 a11790a <=( a11789a  and  a11784a );
 a11793a <=( A166  and  A168 );
 a11797a <=( (not A232)  and  A200 );
 a11798a <=( A199  and  a11797a );
 a11799a <=( a11798a  and  a11793a );
 a11802a <=( A298  and  A233 );
 a11806a <=( A302  and  A300 );
 a11807a <=( (not A299)  and  a11806a );
 a11808a <=( a11807a  and  a11802a );
 a11811a <=( A166  and  A168 );
 a11815a <=( (not A232)  and  A200 );
 a11816a <=( A199  and  a11815a );
 a11817a <=( a11816a  and  a11811a );
 a11820a <=( A265  and  A233 );
 a11824a <=( A268  and  A267 );
 a11825a <=( (not A266)  and  a11824a );
 a11826a <=( a11825a  and  a11820a );
 a11829a <=( A166  and  A168 );
 a11833a <=( (not A232)  and  A200 );
 a11834a <=( A199  and  a11833a );
 a11835a <=( a11834a  and  a11829a );
 a11838a <=( A265  and  A233 );
 a11842a <=( A269  and  A267 );
 a11843a <=( (not A266)  and  a11842a );
 a11844a <=( a11843a  and  a11838a );
 a11847a <=( A166  and  A168 );
 a11851a <=( (not A233)  and  A200 );
 a11852a <=( A199  and  a11851a );
 a11853a <=( a11852a  and  a11847a );
 a11856a <=( A265  and  (not A234) );
 a11860a <=( (not A300)  and  A298 );
 a11861a <=( A266  and  a11860a );
 a11862a <=( a11861a  and  a11856a );
 a11865a <=( A166  and  A168 );
 a11869a <=( (not A233)  and  A200 );
 a11870a <=( A199  and  a11869a );
 a11871a <=( a11870a  and  a11865a );
 a11874a <=( A265  and  (not A234) );
 a11878a <=( A299  and  A298 );
 a11879a <=( A266  and  a11878a );
 a11880a <=( a11879a  and  a11874a );
 a11883a <=( A166  and  A168 );
 a11887a <=( (not A233)  and  A200 );
 a11888a <=( A199  and  a11887a );
 a11889a <=( a11888a  and  a11883a );
 a11892a <=( A265  and  (not A234) );
 a11896a <=( (not A299)  and  (not A298) );
 a11897a <=( A266  and  a11896a );
 a11898a <=( a11897a  and  a11892a );
 a11901a <=( A166  and  A168 );
 a11905a <=( (not A233)  and  A200 );
 a11906a <=( A199  and  a11905a );
 a11907a <=( a11906a  and  a11901a );
 a11910a <=( (not A266)  and  (not A234) );
 a11914a <=( (not A300)  and  A298 );
 a11915a <=( (not A267)  and  a11914a );
 a11916a <=( a11915a  and  a11910a );
 a11919a <=( A166  and  A168 );
 a11923a <=( (not A233)  and  A200 );
 a11924a <=( A199  and  a11923a );
 a11925a <=( a11924a  and  a11919a );
 a11928a <=( (not A266)  and  (not A234) );
 a11932a <=( A299  and  A298 );
 a11933a <=( (not A267)  and  a11932a );
 a11934a <=( a11933a  and  a11928a );
 a11937a <=( A166  and  A168 );
 a11941a <=( (not A233)  and  A200 );
 a11942a <=( A199  and  a11941a );
 a11943a <=( a11942a  and  a11937a );
 a11946a <=( (not A266)  and  (not A234) );
 a11950a <=( (not A299)  and  (not A298) );
 a11951a <=( (not A267)  and  a11950a );
 a11952a <=( a11951a  and  a11946a );
 a11955a <=( A166  and  A168 );
 a11959a <=( (not A233)  and  A200 );
 a11960a <=( A199  and  a11959a );
 a11961a <=( a11960a  and  a11955a );
 a11964a <=( (not A265)  and  (not A234) );
 a11968a <=( (not A300)  and  A298 );
 a11969a <=( (not A266)  and  a11968a );
 a11970a <=( a11969a  and  a11964a );
 a11973a <=( A166  and  A168 );
 a11977a <=( (not A233)  and  A200 );
 a11978a <=( A199  and  a11977a );
 a11979a <=( a11978a  and  a11973a );
 a11982a <=( (not A265)  and  (not A234) );
 a11986a <=( A299  and  A298 );
 a11987a <=( (not A266)  and  a11986a );
 a11988a <=( a11987a  and  a11982a );
 a11991a <=( A166  and  A168 );
 a11995a <=( (not A233)  and  A200 );
 a11996a <=( A199  and  a11995a );
 a11997a <=( a11996a  and  a11991a );
 a12000a <=( (not A265)  and  (not A234) );
 a12004a <=( (not A299)  and  (not A298) );
 a12005a <=( (not A266)  and  a12004a );
 a12006a <=( a12005a  and  a12000a );
 a12009a <=( A166  and  A168 );
 a12013a <=( A232  and  A200 );
 a12014a <=( A199  and  a12013a );
 a12015a <=( a12014a  and  a12009a );
 a12018a <=( A234  and  (not A233) );
 a12022a <=( A299  and  (not A298) );
 a12023a <=( A235  and  a12022a );
 a12024a <=( a12023a  and  a12018a );
 a12027a <=( A166  and  A168 );
 a12031a <=( A232  and  A200 );
 a12032a <=( A199  and  a12031a );
 a12033a <=( a12032a  and  a12027a );
 a12036a <=( A234  and  (not A233) );
 a12040a <=( A266  and  (not A265) );
 a12041a <=( A235  and  a12040a );
 a12042a <=( a12041a  and  a12036a );
 a12045a <=( A166  and  A168 );
 a12049a <=( A232  and  A200 );
 a12050a <=( A199  and  a12049a );
 a12051a <=( a12050a  and  a12045a );
 a12054a <=( A234  and  (not A233) );
 a12058a <=( A299  and  (not A298) );
 a12059a <=( A236  and  a12058a );
 a12060a <=( a12059a  and  a12054a );
 a12063a <=( A166  and  A168 );
 a12067a <=( A232  and  A200 );
 a12068a <=( A199  and  a12067a );
 a12069a <=( a12068a  and  a12063a );
 a12072a <=( A234  and  (not A233) );
 a12076a <=( A266  and  (not A265) );
 a12077a <=( A236  and  a12076a );
 a12078a <=( a12077a  and  a12072a );
 a12081a <=( A166  and  A168 );
 a12085a <=( (not A232)  and  A200 );
 a12086a <=( A199  and  a12085a );
 a12087a <=( a12086a  and  a12081a );
 a12090a <=( A265  and  (not A233) );
 a12094a <=( (not A300)  and  A298 );
 a12095a <=( A266  and  a12094a );
 a12096a <=( a12095a  and  a12090a );
 a12099a <=( A166  and  A168 );
 a12103a <=( (not A232)  and  A200 );
 a12104a <=( A199  and  a12103a );
 a12105a <=( a12104a  and  a12099a );
 a12108a <=( A265  and  (not A233) );
 a12112a <=( A299  and  A298 );
 a12113a <=( A266  and  a12112a );
 a12114a <=( a12113a  and  a12108a );
 a12117a <=( A166  and  A168 );
 a12121a <=( (not A232)  and  A200 );
 a12122a <=( A199  and  a12121a );
 a12123a <=( a12122a  and  a12117a );
 a12126a <=( A265  and  (not A233) );
 a12130a <=( (not A299)  and  (not A298) );
 a12131a <=( A266  and  a12130a );
 a12132a <=( a12131a  and  a12126a );
 a12135a <=( A166  and  A168 );
 a12139a <=( (not A232)  and  A200 );
 a12140a <=( A199  and  a12139a );
 a12141a <=( a12140a  and  a12135a );
 a12144a <=( (not A266)  and  (not A233) );
 a12148a <=( (not A300)  and  A298 );
 a12149a <=( (not A267)  and  a12148a );
 a12150a <=( a12149a  and  a12144a );
 a12153a <=( A166  and  A168 );
 a12157a <=( (not A232)  and  A200 );
 a12158a <=( A199  and  a12157a );
 a12159a <=( a12158a  and  a12153a );
 a12162a <=( (not A266)  and  (not A233) );
 a12166a <=( A299  and  A298 );
 a12167a <=( (not A267)  and  a12166a );
 a12168a <=( a12167a  and  a12162a );
 a12171a <=( A166  and  A168 );
 a12175a <=( (not A232)  and  A200 );
 a12176a <=( A199  and  a12175a );
 a12177a <=( a12176a  and  a12171a );
 a12180a <=( (not A266)  and  (not A233) );
 a12184a <=( (not A299)  and  (not A298) );
 a12185a <=( (not A267)  and  a12184a );
 a12186a <=( a12185a  and  a12180a );
 a12189a <=( A166  and  A168 );
 a12193a <=( (not A232)  and  A200 );
 a12194a <=( A199  and  a12193a );
 a12195a <=( a12194a  and  a12189a );
 a12198a <=( (not A265)  and  (not A233) );
 a12202a <=( (not A300)  and  A298 );
 a12203a <=( (not A266)  and  a12202a );
 a12204a <=( a12203a  and  a12198a );
 a12207a <=( A166  and  A168 );
 a12211a <=( (not A232)  and  A200 );
 a12212a <=( A199  and  a12211a );
 a12213a <=( a12212a  and  a12207a );
 a12216a <=( (not A265)  and  (not A233) );
 a12220a <=( A299  and  A298 );
 a12221a <=( (not A266)  and  a12220a );
 a12222a <=( a12221a  and  a12216a );
 a12225a <=( A166  and  A168 );
 a12229a <=( (not A232)  and  A200 );
 a12230a <=( A199  and  a12229a );
 a12231a <=( a12230a  and  a12225a );
 a12234a <=( (not A265)  and  (not A233) );
 a12238a <=( (not A299)  and  (not A298) );
 a12239a <=( (not A266)  and  a12238a );
 a12240a <=( a12239a  and  a12234a );
 a12243a <=( A166  and  A168 );
 a12247a <=( A232  and  (not A201) );
 a12248a <=( (not A200)  and  a12247a );
 a12249a <=( a12248a  and  a12243a );
 a12252a <=( A265  and  A233 );
 a12256a <=( (not A300)  and  (not A299) );
 a12257a <=( (not A267)  and  a12256a );
 a12258a <=( a12257a  and  a12252a );
 a12261a <=( A166  and  A168 );
 a12265a <=( A232  and  (not A201) );
 a12266a <=( (not A200)  and  a12265a );
 a12267a <=( a12266a  and  a12261a );
 a12270a <=( A265  and  A233 );
 a12274a <=( A299  and  A298 );
 a12275a <=( (not A267)  and  a12274a );
 a12276a <=( a12275a  and  a12270a );
 a12279a <=( A166  and  A168 );
 a12283a <=( A232  and  (not A201) );
 a12284a <=( (not A200)  and  a12283a );
 a12285a <=( a12284a  and  a12279a );
 a12288a <=( A265  and  A233 );
 a12292a <=( (not A299)  and  (not A298) );
 a12293a <=( (not A267)  and  a12292a );
 a12294a <=( a12293a  and  a12288a );
 a12297a <=( A166  and  A168 );
 a12301a <=( A232  and  (not A201) );
 a12302a <=( (not A200)  and  a12301a );
 a12303a <=( a12302a  and  a12297a );
 a12306a <=( A265  and  A233 );
 a12310a <=( (not A300)  and  (not A299) );
 a12311a <=( A266  and  a12310a );
 a12312a <=( a12311a  and  a12306a );
 a12315a <=( A166  and  A168 );
 a12319a <=( A232  and  (not A201) );
 a12320a <=( (not A200)  and  a12319a );
 a12321a <=( a12320a  and  a12315a );
 a12324a <=( A265  and  A233 );
 a12328a <=( A299  and  A298 );
 a12329a <=( A266  and  a12328a );
 a12330a <=( a12329a  and  a12324a );
 a12333a <=( A166  and  A168 );
 a12337a <=( A232  and  (not A201) );
 a12338a <=( (not A200)  and  a12337a );
 a12339a <=( a12338a  and  a12333a );
 a12342a <=( A265  and  A233 );
 a12346a <=( (not A299)  and  (not A298) );
 a12347a <=( A266  and  a12346a );
 a12348a <=( a12347a  and  a12342a );
 a12351a <=( A166  and  A168 );
 a12355a <=( A232  and  (not A201) );
 a12356a <=( (not A200)  and  a12355a );
 a12357a <=( a12356a  and  a12351a );
 a12360a <=( (not A265)  and  A233 );
 a12364a <=( (not A300)  and  (not A299) );
 a12365a <=( (not A266)  and  a12364a );
 a12366a <=( a12365a  and  a12360a );
 a12369a <=( A166  and  A168 );
 a12373a <=( A232  and  (not A201) );
 a12374a <=( (not A200)  and  a12373a );
 a12375a <=( a12374a  and  a12369a );
 a12378a <=( (not A265)  and  A233 );
 a12382a <=( A299  and  A298 );
 a12383a <=( (not A266)  and  a12382a );
 a12384a <=( a12383a  and  a12378a );
 a12387a <=( A166  and  A168 );
 a12391a <=( A232  and  (not A201) );
 a12392a <=( (not A200)  and  a12391a );
 a12393a <=( a12392a  and  a12387a );
 a12396a <=( (not A265)  and  A233 );
 a12400a <=( (not A299)  and  (not A298) );
 a12401a <=( (not A266)  and  a12400a );
 a12402a <=( a12401a  and  a12396a );
 a12405a <=( A166  and  A168 );
 a12409a <=( (not A232)  and  (not A201) );
 a12410a <=( (not A200)  and  a12409a );
 a12411a <=( a12410a  and  a12405a );
 a12414a <=( A298  and  A233 );
 a12418a <=( A301  and  A300 );
 a12419a <=( (not A299)  and  a12418a );
 a12420a <=( a12419a  and  a12414a );
 a12423a <=( A166  and  A168 );
 a12427a <=( (not A232)  and  (not A201) );
 a12428a <=( (not A200)  and  a12427a );
 a12429a <=( a12428a  and  a12423a );
 a12432a <=( A298  and  A233 );
 a12436a <=( A302  and  A300 );
 a12437a <=( (not A299)  and  a12436a );
 a12438a <=( a12437a  and  a12432a );
 a12441a <=( A166  and  A168 );
 a12445a <=( (not A232)  and  (not A201) );
 a12446a <=( (not A200)  and  a12445a );
 a12447a <=( a12446a  and  a12441a );
 a12450a <=( A265  and  A233 );
 a12454a <=( A268  and  A267 );
 a12455a <=( (not A266)  and  a12454a );
 a12456a <=( a12455a  and  a12450a );
 a12459a <=( A166  and  A168 );
 a12463a <=( (not A232)  and  (not A201) );
 a12464a <=( (not A200)  and  a12463a );
 a12465a <=( a12464a  and  a12459a );
 a12468a <=( A265  and  A233 );
 a12472a <=( A269  and  A267 );
 a12473a <=( (not A266)  and  a12472a );
 a12474a <=( a12473a  and  a12468a );
 a12477a <=( A166  and  A168 );
 a12481a <=( (not A233)  and  (not A201) );
 a12482a <=( (not A200)  and  a12481a );
 a12483a <=( a12482a  and  a12477a );
 a12486a <=( A265  and  (not A234) );
 a12490a <=( (not A300)  and  A298 );
 a12491a <=( A266  and  a12490a );
 a12492a <=( a12491a  and  a12486a );
 a12495a <=( A166  and  A168 );
 a12499a <=( (not A233)  and  (not A201) );
 a12500a <=( (not A200)  and  a12499a );
 a12501a <=( a12500a  and  a12495a );
 a12504a <=( A265  and  (not A234) );
 a12508a <=( A299  and  A298 );
 a12509a <=( A266  and  a12508a );
 a12510a <=( a12509a  and  a12504a );
 a12513a <=( A166  and  A168 );
 a12517a <=( (not A233)  and  (not A201) );
 a12518a <=( (not A200)  and  a12517a );
 a12519a <=( a12518a  and  a12513a );
 a12522a <=( A265  and  (not A234) );
 a12526a <=( (not A299)  and  (not A298) );
 a12527a <=( A266  and  a12526a );
 a12528a <=( a12527a  and  a12522a );
 a12531a <=( A166  and  A168 );
 a12535a <=( (not A233)  and  (not A201) );
 a12536a <=( (not A200)  and  a12535a );
 a12537a <=( a12536a  and  a12531a );
 a12540a <=( (not A266)  and  (not A234) );
 a12544a <=( (not A300)  and  A298 );
 a12545a <=( (not A267)  and  a12544a );
 a12546a <=( a12545a  and  a12540a );
 a12549a <=( A166  and  A168 );
 a12553a <=( (not A233)  and  (not A201) );
 a12554a <=( (not A200)  and  a12553a );
 a12555a <=( a12554a  and  a12549a );
 a12558a <=( (not A266)  and  (not A234) );
 a12562a <=( A299  and  A298 );
 a12563a <=( (not A267)  and  a12562a );
 a12564a <=( a12563a  and  a12558a );
 a12567a <=( A166  and  A168 );
 a12571a <=( (not A233)  and  (not A201) );
 a12572a <=( (not A200)  and  a12571a );
 a12573a <=( a12572a  and  a12567a );
 a12576a <=( (not A266)  and  (not A234) );
 a12580a <=( (not A299)  and  (not A298) );
 a12581a <=( (not A267)  and  a12580a );
 a12582a <=( a12581a  and  a12576a );
 a12585a <=( A166  and  A168 );
 a12589a <=( (not A233)  and  (not A201) );
 a12590a <=( (not A200)  and  a12589a );
 a12591a <=( a12590a  and  a12585a );
 a12594a <=( (not A265)  and  (not A234) );
 a12598a <=( (not A300)  and  A298 );
 a12599a <=( (not A266)  and  a12598a );
 a12600a <=( a12599a  and  a12594a );
 a12603a <=( A166  and  A168 );
 a12607a <=( (not A233)  and  (not A201) );
 a12608a <=( (not A200)  and  a12607a );
 a12609a <=( a12608a  and  a12603a );
 a12612a <=( (not A265)  and  (not A234) );
 a12616a <=( A299  and  A298 );
 a12617a <=( (not A266)  and  a12616a );
 a12618a <=( a12617a  and  a12612a );
 a12621a <=( A166  and  A168 );
 a12625a <=( (not A233)  and  (not A201) );
 a12626a <=( (not A200)  and  a12625a );
 a12627a <=( a12626a  and  a12621a );
 a12630a <=( (not A265)  and  (not A234) );
 a12634a <=( (not A299)  and  (not A298) );
 a12635a <=( (not A266)  and  a12634a );
 a12636a <=( a12635a  and  a12630a );
 a12639a <=( A166  and  A168 );
 a12643a <=( A232  and  (not A201) );
 a12644a <=( (not A200)  and  a12643a );
 a12645a <=( a12644a  and  a12639a );
 a12648a <=( A234  and  (not A233) );
 a12652a <=( A299  and  (not A298) );
 a12653a <=( A235  and  a12652a );
 a12654a <=( a12653a  and  a12648a );
 a12657a <=( A166  and  A168 );
 a12661a <=( A232  and  (not A201) );
 a12662a <=( (not A200)  and  a12661a );
 a12663a <=( a12662a  and  a12657a );
 a12666a <=( A234  and  (not A233) );
 a12670a <=( A266  and  (not A265) );
 a12671a <=( A235  and  a12670a );
 a12672a <=( a12671a  and  a12666a );
 a12675a <=( A166  and  A168 );
 a12679a <=( A232  and  (not A201) );
 a12680a <=( (not A200)  and  a12679a );
 a12681a <=( a12680a  and  a12675a );
 a12684a <=( A234  and  (not A233) );
 a12688a <=( A299  and  (not A298) );
 a12689a <=( A236  and  a12688a );
 a12690a <=( a12689a  and  a12684a );
 a12693a <=( A166  and  A168 );
 a12697a <=( A232  and  (not A201) );
 a12698a <=( (not A200)  and  a12697a );
 a12699a <=( a12698a  and  a12693a );
 a12702a <=( A234  and  (not A233) );
 a12706a <=( A266  and  (not A265) );
 a12707a <=( A236  and  a12706a );
 a12708a <=( a12707a  and  a12702a );
 a12711a <=( A166  and  A168 );
 a12715a <=( (not A232)  and  (not A201) );
 a12716a <=( (not A200)  and  a12715a );
 a12717a <=( a12716a  and  a12711a );
 a12720a <=( A265  and  (not A233) );
 a12724a <=( (not A300)  and  A298 );
 a12725a <=( A266  and  a12724a );
 a12726a <=( a12725a  and  a12720a );
 a12729a <=( A166  and  A168 );
 a12733a <=( (not A232)  and  (not A201) );
 a12734a <=( (not A200)  and  a12733a );
 a12735a <=( a12734a  and  a12729a );
 a12738a <=( A265  and  (not A233) );
 a12742a <=( A299  and  A298 );
 a12743a <=( A266  and  a12742a );
 a12744a <=( a12743a  and  a12738a );
 a12747a <=( A166  and  A168 );
 a12751a <=( (not A232)  and  (not A201) );
 a12752a <=( (not A200)  and  a12751a );
 a12753a <=( a12752a  and  a12747a );
 a12756a <=( A265  and  (not A233) );
 a12760a <=( (not A299)  and  (not A298) );
 a12761a <=( A266  and  a12760a );
 a12762a <=( a12761a  and  a12756a );
 a12765a <=( A166  and  A168 );
 a12769a <=( (not A232)  and  (not A201) );
 a12770a <=( (not A200)  and  a12769a );
 a12771a <=( a12770a  and  a12765a );
 a12774a <=( (not A266)  and  (not A233) );
 a12778a <=( (not A300)  and  A298 );
 a12779a <=( (not A267)  and  a12778a );
 a12780a <=( a12779a  and  a12774a );
 a12783a <=( A166  and  A168 );
 a12787a <=( (not A232)  and  (not A201) );
 a12788a <=( (not A200)  and  a12787a );
 a12789a <=( a12788a  and  a12783a );
 a12792a <=( (not A266)  and  (not A233) );
 a12796a <=( A299  and  A298 );
 a12797a <=( (not A267)  and  a12796a );
 a12798a <=( a12797a  and  a12792a );
 a12801a <=( A166  and  A168 );
 a12805a <=( (not A232)  and  (not A201) );
 a12806a <=( (not A200)  and  a12805a );
 a12807a <=( a12806a  and  a12801a );
 a12810a <=( (not A266)  and  (not A233) );
 a12814a <=( (not A299)  and  (not A298) );
 a12815a <=( (not A267)  and  a12814a );
 a12816a <=( a12815a  and  a12810a );
 a12819a <=( A166  and  A168 );
 a12823a <=( (not A232)  and  (not A201) );
 a12824a <=( (not A200)  and  a12823a );
 a12825a <=( a12824a  and  a12819a );
 a12828a <=( (not A265)  and  (not A233) );
 a12832a <=( (not A300)  and  A298 );
 a12833a <=( (not A266)  and  a12832a );
 a12834a <=( a12833a  and  a12828a );
 a12837a <=( A166  and  A168 );
 a12841a <=( (not A232)  and  (not A201) );
 a12842a <=( (not A200)  and  a12841a );
 a12843a <=( a12842a  and  a12837a );
 a12846a <=( (not A265)  and  (not A233) );
 a12850a <=( A299  and  A298 );
 a12851a <=( (not A266)  and  a12850a );
 a12852a <=( a12851a  and  a12846a );
 a12855a <=( A166  and  A168 );
 a12859a <=( (not A232)  and  (not A201) );
 a12860a <=( (not A200)  and  a12859a );
 a12861a <=( a12860a  and  a12855a );
 a12864a <=( (not A265)  and  (not A233) );
 a12868a <=( (not A299)  and  (not A298) );
 a12869a <=( (not A266)  and  a12868a );
 a12870a <=( a12869a  and  a12864a );
 a12873a <=( A166  and  A168 );
 a12877a <=( A232  and  (not A200) );
 a12878a <=( (not A199)  and  a12877a );
 a12879a <=( a12878a  and  a12873a );
 a12882a <=( A265  and  A233 );
 a12886a <=( (not A300)  and  (not A299) );
 a12887a <=( (not A267)  and  a12886a );
 a12888a <=( a12887a  and  a12882a );
 a12891a <=( A166  and  A168 );
 a12895a <=( A232  and  (not A200) );
 a12896a <=( (not A199)  and  a12895a );
 a12897a <=( a12896a  and  a12891a );
 a12900a <=( A265  and  A233 );
 a12904a <=( A299  and  A298 );
 a12905a <=( (not A267)  and  a12904a );
 a12906a <=( a12905a  and  a12900a );
 a12909a <=( A166  and  A168 );
 a12913a <=( A232  and  (not A200) );
 a12914a <=( (not A199)  and  a12913a );
 a12915a <=( a12914a  and  a12909a );
 a12918a <=( A265  and  A233 );
 a12922a <=( (not A299)  and  (not A298) );
 a12923a <=( (not A267)  and  a12922a );
 a12924a <=( a12923a  and  a12918a );
 a12927a <=( A166  and  A168 );
 a12931a <=( A232  and  (not A200) );
 a12932a <=( (not A199)  and  a12931a );
 a12933a <=( a12932a  and  a12927a );
 a12936a <=( A265  and  A233 );
 a12940a <=( (not A300)  and  (not A299) );
 a12941a <=( A266  and  a12940a );
 a12942a <=( a12941a  and  a12936a );
 a12945a <=( A166  and  A168 );
 a12949a <=( A232  and  (not A200) );
 a12950a <=( (not A199)  and  a12949a );
 a12951a <=( a12950a  and  a12945a );
 a12954a <=( A265  and  A233 );
 a12958a <=( A299  and  A298 );
 a12959a <=( A266  and  a12958a );
 a12960a <=( a12959a  and  a12954a );
 a12963a <=( A166  and  A168 );
 a12967a <=( A232  and  (not A200) );
 a12968a <=( (not A199)  and  a12967a );
 a12969a <=( a12968a  and  a12963a );
 a12972a <=( A265  and  A233 );
 a12976a <=( (not A299)  and  (not A298) );
 a12977a <=( A266  and  a12976a );
 a12978a <=( a12977a  and  a12972a );
 a12981a <=( A166  and  A168 );
 a12985a <=( A232  and  (not A200) );
 a12986a <=( (not A199)  and  a12985a );
 a12987a <=( a12986a  and  a12981a );
 a12990a <=( (not A265)  and  A233 );
 a12994a <=( (not A300)  and  (not A299) );
 a12995a <=( (not A266)  and  a12994a );
 a12996a <=( a12995a  and  a12990a );
 a12999a <=( A166  and  A168 );
 a13003a <=( A232  and  (not A200) );
 a13004a <=( (not A199)  and  a13003a );
 a13005a <=( a13004a  and  a12999a );
 a13008a <=( (not A265)  and  A233 );
 a13012a <=( A299  and  A298 );
 a13013a <=( (not A266)  and  a13012a );
 a13014a <=( a13013a  and  a13008a );
 a13017a <=( A166  and  A168 );
 a13021a <=( A232  and  (not A200) );
 a13022a <=( (not A199)  and  a13021a );
 a13023a <=( a13022a  and  a13017a );
 a13026a <=( (not A265)  and  A233 );
 a13030a <=( (not A299)  and  (not A298) );
 a13031a <=( (not A266)  and  a13030a );
 a13032a <=( a13031a  and  a13026a );
 a13035a <=( A166  and  A168 );
 a13039a <=( (not A232)  and  (not A200) );
 a13040a <=( (not A199)  and  a13039a );
 a13041a <=( a13040a  and  a13035a );
 a13044a <=( A298  and  A233 );
 a13048a <=( A301  and  A300 );
 a13049a <=( (not A299)  and  a13048a );
 a13050a <=( a13049a  and  a13044a );
 a13053a <=( A166  and  A168 );
 a13057a <=( (not A232)  and  (not A200) );
 a13058a <=( (not A199)  and  a13057a );
 a13059a <=( a13058a  and  a13053a );
 a13062a <=( A298  and  A233 );
 a13066a <=( A302  and  A300 );
 a13067a <=( (not A299)  and  a13066a );
 a13068a <=( a13067a  and  a13062a );
 a13071a <=( A166  and  A168 );
 a13075a <=( (not A232)  and  (not A200) );
 a13076a <=( (not A199)  and  a13075a );
 a13077a <=( a13076a  and  a13071a );
 a13080a <=( A265  and  A233 );
 a13084a <=( A268  and  A267 );
 a13085a <=( (not A266)  and  a13084a );
 a13086a <=( a13085a  and  a13080a );
 a13089a <=( A166  and  A168 );
 a13093a <=( (not A232)  and  (not A200) );
 a13094a <=( (not A199)  and  a13093a );
 a13095a <=( a13094a  and  a13089a );
 a13098a <=( A265  and  A233 );
 a13102a <=( A269  and  A267 );
 a13103a <=( (not A266)  and  a13102a );
 a13104a <=( a13103a  and  a13098a );
 a13107a <=( A166  and  A168 );
 a13111a <=( (not A233)  and  (not A200) );
 a13112a <=( (not A199)  and  a13111a );
 a13113a <=( a13112a  and  a13107a );
 a13116a <=( A265  and  (not A234) );
 a13120a <=( (not A300)  and  A298 );
 a13121a <=( A266  and  a13120a );
 a13122a <=( a13121a  and  a13116a );
 a13125a <=( A166  and  A168 );
 a13129a <=( (not A233)  and  (not A200) );
 a13130a <=( (not A199)  and  a13129a );
 a13131a <=( a13130a  and  a13125a );
 a13134a <=( A265  and  (not A234) );
 a13138a <=( A299  and  A298 );
 a13139a <=( A266  and  a13138a );
 a13140a <=( a13139a  and  a13134a );
 a13143a <=( A166  and  A168 );
 a13147a <=( (not A233)  and  (not A200) );
 a13148a <=( (not A199)  and  a13147a );
 a13149a <=( a13148a  and  a13143a );
 a13152a <=( A265  and  (not A234) );
 a13156a <=( (not A299)  and  (not A298) );
 a13157a <=( A266  and  a13156a );
 a13158a <=( a13157a  and  a13152a );
 a13161a <=( A166  and  A168 );
 a13165a <=( (not A233)  and  (not A200) );
 a13166a <=( (not A199)  and  a13165a );
 a13167a <=( a13166a  and  a13161a );
 a13170a <=( (not A266)  and  (not A234) );
 a13174a <=( (not A300)  and  A298 );
 a13175a <=( (not A267)  and  a13174a );
 a13176a <=( a13175a  and  a13170a );
 a13179a <=( A166  and  A168 );
 a13183a <=( (not A233)  and  (not A200) );
 a13184a <=( (not A199)  and  a13183a );
 a13185a <=( a13184a  and  a13179a );
 a13188a <=( (not A266)  and  (not A234) );
 a13192a <=( A299  and  A298 );
 a13193a <=( (not A267)  and  a13192a );
 a13194a <=( a13193a  and  a13188a );
 a13197a <=( A166  and  A168 );
 a13201a <=( (not A233)  and  (not A200) );
 a13202a <=( (not A199)  and  a13201a );
 a13203a <=( a13202a  and  a13197a );
 a13206a <=( (not A266)  and  (not A234) );
 a13210a <=( (not A299)  and  (not A298) );
 a13211a <=( (not A267)  and  a13210a );
 a13212a <=( a13211a  and  a13206a );
 a13215a <=( A166  and  A168 );
 a13219a <=( (not A233)  and  (not A200) );
 a13220a <=( (not A199)  and  a13219a );
 a13221a <=( a13220a  and  a13215a );
 a13224a <=( (not A265)  and  (not A234) );
 a13228a <=( (not A300)  and  A298 );
 a13229a <=( (not A266)  and  a13228a );
 a13230a <=( a13229a  and  a13224a );
 a13233a <=( A166  and  A168 );
 a13237a <=( (not A233)  and  (not A200) );
 a13238a <=( (not A199)  and  a13237a );
 a13239a <=( a13238a  and  a13233a );
 a13242a <=( (not A265)  and  (not A234) );
 a13246a <=( A299  and  A298 );
 a13247a <=( (not A266)  and  a13246a );
 a13248a <=( a13247a  and  a13242a );
 a13251a <=( A166  and  A168 );
 a13255a <=( (not A233)  and  (not A200) );
 a13256a <=( (not A199)  and  a13255a );
 a13257a <=( a13256a  and  a13251a );
 a13260a <=( (not A265)  and  (not A234) );
 a13264a <=( (not A299)  and  (not A298) );
 a13265a <=( (not A266)  and  a13264a );
 a13266a <=( a13265a  and  a13260a );
 a13269a <=( A166  and  A168 );
 a13273a <=( A232  and  (not A200) );
 a13274a <=( (not A199)  and  a13273a );
 a13275a <=( a13274a  and  a13269a );
 a13278a <=( A234  and  (not A233) );
 a13282a <=( A299  and  (not A298) );
 a13283a <=( A235  and  a13282a );
 a13284a <=( a13283a  and  a13278a );
 a13287a <=( A166  and  A168 );
 a13291a <=( A232  and  (not A200) );
 a13292a <=( (not A199)  and  a13291a );
 a13293a <=( a13292a  and  a13287a );
 a13296a <=( A234  and  (not A233) );
 a13300a <=( A266  and  (not A265) );
 a13301a <=( A235  and  a13300a );
 a13302a <=( a13301a  and  a13296a );
 a13305a <=( A166  and  A168 );
 a13309a <=( A232  and  (not A200) );
 a13310a <=( (not A199)  and  a13309a );
 a13311a <=( a13310a  and  a13305a );
 a13314a <=( A234  and  (not A233) );
 a13318a <=( A299  and  (not A298) );
 a13319a <=( A236  and  a13318a );
 a13320a <=( a13319a  and  a13314a );
 a13323a <=( A166  and  A168 );
 a13327a <=( A232  and  (not A200) );
 a13328a <=( (not A199)  and  a13327a );
 a13329a <=( a13328a  and  a13323a );
 a13332a <=( A234  and  (not A233) );
 a13336a <=( A266  and  (not A265) );
 a13337a <=( A236  and  a13336a );
 a13338a <=( a13337a  and  a13332a );
 a13341a <=( A166  and  A168 );
 a13345a <=( (not A232)  and  (not A200) );
 a13346a <=( (not A199)  and  a13345a );
 a13347a <=( a13346a  and  a13341a );
 a13350a <=( A265  and  (not A233) );
 a13354a <=( (not A300)  and  A298 );
 a13355a <=( A266  and  a13354a );
 a13356a <=( a13355a  and  a13350a );
 a13359a <=( A166  and  A168 );
 a13363a <=( (not A232)  and  (not A200) );
 a13364a <=( (not A199)  and  a13363a );
 a13365a <=( a13364a  and  a13359a );
 a13368a <=( A265  and  (not A233) );
 a13372a <=( A299  and  A298 );
 a13373a <=( A266  and  a13372a );
 a13374a <=( a13373a  and  a13368a );
 a13377a <=( A166  and  A168 );
 a13381a <=( (not A232)  and  (not A200) );
 a13382a <=( (not A199)  and  a13381a );
 a13383a <=( a13382a  and  a13377a );
 a13386a <=( A265  and  (not A233) );
 a13390a <=( (not A299)  and  (not A298) );
 a13391a <=( A266  and  a13390a );
 a13392a <=( a13391a  and  a13386a );
 a13395a <=( A166  and  A168 );
 a13399a <=( (not A232)  and  (not A200) );
 a13400a <=( (not A199)  and  a13399a );
 a13401a <=( a13400a  and  a13395a );
 a13404a <=( (not A266)  and  (not A233) );
 a13408a <=( (not A300)  and  A298 );
 a13409a <=( (not A267)  and  a13408a );
 a13410a <=( a13409a  and  a13404a );
 a13413a <=( A166  and  A168 );
 a13417a <=( (not A232)  and  (not A200) );
 a13418a <=( (not A199)  and  a13417a );
 a13419a <=( a13418a  and  a13413a );
 a13422a <=( (not A266)  and  (not A233) );
 a13426a <=( A299  and  A298 );
 a13427a <=( (not A267)  and  a13426a );
 a13428a <=( a13427a  and  a13422a );
 a13431a <=( A166  and  A168 );
 a13435a <=( (not A232)  and  (not A200) );
 a13436a <=( (not A199)  and  a13435a );
 a13437a <=( a13436a  and  a13431a );
 a13440a <=( (not A266)  and  (not A233) );
 a13444a <=( (not A299)  and  (not A298) );
 a13445a <=( (not A267)  and  a13444a );
 a13446a <=( a13445a  and  a13440a );
 a13449a <=( A166  and  A168 );
 a13453a <=( (not A232)  and  (not A200) );
 a13454a <=( (not A199)  and  a13453a );
 a13455a <=( a13454a  and  a13449a );
 a13458a <=( (not A265)  and  (not A233) );
 a13462a <=( (not A300)  and  A298 );
 a13463a <=( (not A266)  and  a13462a );
 a13464a <=( a13463a  and  a13458a );
 a13467a <=( A166  and  A168 );
 a13471a <=( (not A232)  and  (not A200) );
 a13472a <=( (not A199)  and  a13471a );
 a13473a <=( a13472a  and  a13467a );
 a13476a <=( (not A265)  and  (not A233) );
 a13480a <=( A299  and  A298 );
 a13481a <=( (not A266)  and  a13480a );
 a13482a <=( a13481a  and  a13476a );
 a13485a <=( A166  and  A168 );
 a13489a <=( (not A232)  and  (not A200) );
 a13490a <=( (not A199)  and  a13489a );
 a13491a <=( a13490a  and  a13485a );
 a13494a <=( (not A265)  and  (not A233) );
 a13498a <=( (not A299)  and  (not A298) );
 a13499a <=( (not A266)  and  a13498a );
 a13500a <=( a13499a  and  a13494a );
 a13503a <=( A167  and  A168 );
 a13507a <=( A232  and  A200 );
 a13508a <=( A199  and  a13507a );
 a13509a <=( a13508a  and  a13503a );
 a13512a <=( A265  and  A233 );
 a13516a <=( (not A300)  and  (not A299) );
 a13517a <=( (not A267)  and  a13516a );
 a13518a <=( a13517a  and  a13512a );
 a13521a <=( A167  and  A168 );
 a13525a <=( A232  and  A200 );
 a13526a <=( A199  and  a13525a );
 a13527a <=( a13526a  and  a13521a );
 a13530a <=( A265  and  A233 );
 a13534a <=( A299  and  A298 );
 a13535a <=( (not A267)  and  a13534a );
 a13536a <=( a13535a  and  a13530a );
 a13539a <=( A167  and  A168 );
 a13543a <=( A232  and  A200 );
 a13544a <=( A199  and  a13543a );
 a13545a <=( a13544a  and  a13539a );
 a13548a <=( A265  and  A233 );
 a13552a <=( (not A299)  and  (not A298) );
 a13553a <=( (not A267)  and  a13552a );
 a13554a <=( a13553a  and  a13548a );
 a13557a <=( A167  and  A168 );
 a13561a <=( A232  and  A200 );
 a13562a <=( A199  and  a13561a );
 a13563a <=( a13562a  and  a13557a );
 a13566a <=( A265  and  A233 );
 a13570a <=( (not A300)  and  (not A299) );
 a13571a <=( A266  and  a13570a );
 a13572a <=( a13571a  and  a13566a );
 a13575a <=( A167  and  A168 );
 a13579a <=( A232  and  A200 );
 a13580a <=( A199  and  a13579a );
 a13581a <=( a13580a  and  a13575a );
 a13584a <=( A265  and  A233 );
 a13588a <=( A299  and  A298 );
 a13589a <=( A266  and  a13588a );
 a13590a <=( a13589a  and  a13584a );
 a13593a <=( A167  and  A168 );
 a13597a <=( A232  and  A200 );
 a13598a <=( A199  and  a13597a );
 a13599a <=( a13598a  and  a13593a );
 a13602a <=( A265  and  A233 );
 a13606a <=( (not A299)  and  (not A298) );
 a13607a <=( A266  and  a13606a );
 a13608a <=( a13607a  and  a13602a );
 a13611a <=( A167  and  A168 );
 a13615a <=( A232  and  A200 );
 a13616a <=( A199  and  a13615a );
 a13617a <=( a13616a  and  a13611a );
 a13620a <=( (not A265)  and  A233 );
 a13624a <=( (not A300)  and  (not A299) );
 a13625a <=( (not A266)  and  a13624a );
 a13626a <=( a13625a  and  a13620a );
 a13629a <=( A167  and  A168 );
 a13633a <=( A232  and  A200 );
 a13634a <=( A199  and  a13633a );
 a13635a <=( a13634a  and  a13629a );
 a13638a <=( (not A265)  and  A233 );
 a13642a <=( A299  and  A298 );
 a13643a <=( (not A266)  and  a13642a );
 a13644a <=( a13643a  and  a13638a );
 a13647a <=( A167  and  A168 );
 a13651a <=( A232  and  A200 );
 a13652a <=( A199  and  a13651a );
 a13653a <=( a13652a  and  a13647a );
 a13656a <=( (not A265)  and  A233 );
 a13660a <=( (not A299)  and  (not A298) );
 a13661a <=( (not A266)  and  a13660a );
 a13662a <=( a13661a  and  a13656a );
 a13665a <=( A167  and  A168 );
 a13669a <=( (not A232)  and  A200 );
 a13670a <=( A199  and  a13669a );
 a13671a <=( a13670a  and  a13665a );
 a13674a <=( A298  and  A233 );
 a13678a <=( A301  and  A300 );
 a13679a <=( (not A299)  and  a13678a );
 a13680a <=( a13679a  and  a13674a );
 a13683a <=( A167  and  A168 );
 a13687a <=( (not A232)  and  A200 );
 a13688a <=( A199  and  a13687a );
 a13689a <=( a13688a  and  a13683a );
 a13692a <=( A298  and  A233 );
 a13696a <=( A302  and  A300 );
 a13697a <=( (not A299)  and  a13696a );
 a13698a <=( a13697a  and  a13692a );
 a13701a <=( A167  and  A168 );
 a13705a <=( (not A232)  and  A200 );
 a13706a <=( A199  and  a13705a );
 a13707a <=( a13706a  and  a13701a );
 a13710a <=( A265  and  A233 );
 a13714a <=( A268  and  A267 );
 a13715a <=( (not A266)  and  a13714a );
 a13716a <=( a13715a  and  a13710a );
 a13719a <=( A167  and  A168 );
 a13723a <=( (not A232)  and  A200 );
 a13724a <=( A199  and  a13723a );
 a13725a <=( a13724a  and  a13719a );
 a13728a <=( A265  and  A233 );
 a13732a <=( A269  and  A267 );
 a13733a <=( (not A266)  and  a13732a );
 a13734a <=( a13733a  and  a13728a );
 a13737a <=( A167  and  A168 );
 a13741a <=( (not A233)  and  A200 );
 a13742a <=( A199  and  a13741a );
 a13743a <=( a13742a  and  a13737a );
 a13746a <=( A265  and  (not A234) );
 a13750a <=( (not A300)  and  A298 );
 a13751a <=( A266  and  a13750a );
 a13752a <=( a13751a  and  a13746a );
 a13755a <=( A167  and  A168 );
 a13759a <=( (not A233)  and  A200 );
 a13760a <=( A199  and  a13759a );
 a13761a <=( a13760a  and  a13755a );
 a13764a <=( A265  and  (not A234) );
 a13768a <=( A299  and  A298 );
 a13769a <=( A266  and  a13768a );
 a13770a <=( a13769a  and  a13764a );
 a13773a <=( A167  and  A168 );
 a13777a <=( (not A233)  and  A200 );
 a13778a <=( A199  and  a13777a );
 a13779a <=( a13778a  and  a13773a );
 a13782a <=( A265  and  (not A234) );
 a13786a <=( (not A299)  and  (not A298) );
 a13787a <=( A266  and  a13786a );
 a13788a <=( a13787a  and  a13782a );
 a13791a <=( A167  and  A168 );
 a13795a <=( (not A233)  and  A200 );
 a13796a <=( A199  and  a13795a );
 a13797a <=( a13796a  and  a13791a );
 a13800a <=( (not A266)  and  (not A234) );
 a13804a <=( (not A300)  and  A298 );
 a13805a <=( (not A267)  and  a13804a );
 a13806a <=( a13805a  and  a13800a );
 a13809a <=( A167  and  A168 );
 a13813a <=( (not A233)  and  A200 );
 a13814a <=( A199  and  a13813a );
 a13815a <=( a13814a  and  a13809a );
 a13818a <=( (not A266)  and  (not A234) );
 a13822a <=( A299  and  A298 );
 a13823a <=( (not A267)  and  a13822a );
 a13824a <=( a13823a  and  a13818a );
 a13827a <=( A167  and  A168 );
 a13831a <=( (not A233)  and  A200 );
 a13832a <=( A199  and  a13831a );
 a13833a <=( a13832a  and  a13827a );
 a13836a <=( (not A266)  and  (not A234) );
 a13840a <=( (not A299)  and  (not A298) );
 a13841a <=( (not A267)  and  a13840a );
 a13842a <=( a13841a  and  a13836a );
 a13845a <=( A167  and  A168 );
 a13849a <=( (not A233)  and  A200 );
 a13850a <=( A199  and  a13849a );
 a13851a <=( a13850a  and  a13845a );
 a13854a <=( (not A265)  and  (not A234) );
 a13858a <=( (not A300)  and  A298 );
 a13859a <=( (not A266)  and  a13858a );
 a13860a <=( a13859a  and  a13854a );
 a13863a <=( A167  and  A168 );
 a13867a <=( (not A233)  and  A200 );
 a13868a <=( A199  and  a13867a );
 a13869a <=( a13868a  and  a13863a );
 a13872a <=( (not A265)  and  (not A234) );
 a13876a <=( A299  and  A298 );
 a13877a <=( (not A266)  and  a13876a );
 a13878a <=( a13877a  and  a13872a );
 a13881a <=( A167  and  A168 );
 a13885a <=( (not A233)  and  A200 );
 a13886a <=( A199  and  a13885a );
 a13887a <=( a13886a  and  a13881a );
 a13890a <=( (not A265)  and  (not A234) );
 a13894a <=( (not A299)  and  (not A298) );
 a13895a <=( (not A266)  and  a13894a );
 a13896a <=( a13895a  and  a13890a );
 a13899a <=( A167  and  A168 );
 a13903a <=( A232  and  A200 );
 a13904a <=( A199  and  a13903a );
 a13905a <=( a13904a  and  a13899a );
 a13908a <=( A234  and  (not A233) );
 a13912a <=( A299  and  (not A298) );
 a13913a <=( A235  and  a13912a );
 a13914a <=( a13913a  and  a13908a );
 a13917a <=( A167  and  A168 );
 a13921a <=( A232  and  A200 );
 a13922a <=( A199  and  a13921a );
 a13923a <=( a13922a  and  a13917a );
 a13926a <=( A234  and  (not A233) );
 a13930a <=( A266  and  (not A265) );
 a13931a <=( A235  and  a13930a );
 a13932a <=( a13931a  and  a13926a );
 a13935a <=( A167  and  A168 );
 a13939a <=( A232  and  A200 );
 a13940a <=( A199  and  a13939a );
 a13941a <=( a13940a  and  a13935a );
 a13944a <=( A234  and  (not A233) );
 a13948a <=( A299  and  (not A298) );
 a13949a <=( A236  and  a13948a );
 a13950a <=( a13949a  and  a13944a );
 a13953a <=( A167  and  A168 );
 a13957a <=( A232  and  A200 );
 a13958a <=( A199  and  a13957a );
 a13959a <=( a13958a  and  a13953a );
 a13962a <=( A234  and  (not A233) );
 a13966a <=( A266  and  (not A265) );
 a13967a <=( A236  and  a13966a );
 a13968a <=( a13967a  and  a13962a );
 a13971a <=( A167  and  A168 );
 a13975a <=( (not A232)  and  A200 );
 a13976a <=( A199  and  a13975a );
 a13977a <=( a13976a  and  a13971a );
 a13980a <=( A265  and  (not A233) );
 a13984a <=( (not A300)  and  A298 );
 a13985a <=( A266  and  a13984a );
 a13986a <=( a13985a  and  a13980a );
 a13989a <=( A167  and  A168 );
 a13993a <=( (not A232)  and  A200 );
 a13994a <=( A199  and  a13993a );
 a13995a <=( a13994a  and  a13989a );
 a13998a <=( A265  and  (not A233) );
 a14002a <=( A299  and  A298 );
 a14003a <=( A266  and  a14002a );
 a14004a <=( a14003a  and  a13998a );
 a14007a <=( A167  and  A168 );
 a14011a <=( (not A232)  and  A200 );
 a14012a <=( A199  and  a14011a );
 a14013a <=( a14012a  and  a14007a );
 a14016a <=( A265  and  (not A233) );
 a14020a <=( (not A299)  and  (not A298) );
 a14021a <=( A266  and  a14020a );
 a14022a <=( a14021a  and  a14016a );
 a14025a <=( A167  and  A168 );
 a14029a <=( (not A232)  and  A200 );
 a14030a <=( A199  and  a14029a );
 a14031a <=( a14030a  and  a14025a );
 a14034a <=( (not A266)  and  (not A233) );
 a14038a <=( (not A300)  and  A298 );
 a14039a <=( (not A267)  and  a14038a );
 a14040a <=( a14039a  and  a14034a );
 a14043a <=( A167  and  A168 );
 a14047a <=( (not A232)  and  A200 );
 a14048a <=( A199  and  a14047a );
 a14049a <=( a14048a  and  a14043a );
 a14052a <=( (not A266)  and  (not A233) );
 a14056a <=( A299  and  A298 );
 a14057a <=( (not A267)  and  a14056a );
 a14058a <=( a14057a  and  a14052a );
 a14061a <=( A167  and  A168 );
 a14065a <=( (not A232)  and  A200 );
 a14066a <=( A199  and  a14065a );
 a14067a <=( a14066a  and  a14061a );
 a14070a <=( (not A266)  and  (not A233) );
 a14074a <=( (not A299)  and  (not A298) );
 a14075a <=( (not A267)  and  a14074a );
 a14076a <=( a14075a  and  a14070a );
 a14079a <=( A167  and  A168 );
 a14083a <=( (not A232)  and  A200 );
 a14084a <=( A199  and  a14083a );
 a14085a <=( a14084a  and  a14079a );
 a14088a <=( (not A265)  and  (not A233) );
 a14092a <=( (not A300)  and  A298 );
 a14093a <=( (not A266)  and  a14092a );
 a14094a <=( a14093a  and  a14088a );
 a14097a <=( A167  and  A168 );
 a14101a <=( (not A232)  and  A200 );
 a14102a <=( A199  and  a14101a );
 a14103a <=( a14102a  and  a14097a );
 a14106a <=( (not A265)  and  (not A233) );
 a14110a <=( A299  and  A298 );
 a14111a <=( (not A266)  and  a14110a );
 a14112a <=( a14111a  and  a14106a );
 a14115a <=( A167  and  A168 );
 a14119a <=( (not A232)  and  A200 );
 a14120a <=( A199  and  a14119a );
 a14121a <=( a14120a  and  a14115a );
 a14124a <=( (not A265)  and  (not A233) );
 a14128a <=( (not A299)  and  (not A298) );
 a14129a <=( (not A266)  and  a14128a );
 a14130a <=( a14129a  and  a14124a );
 a14133a <=( A167  and  A168 );
 a14137a <=( A232  and  (not A201) );
 a14138a <=( (not A200)  and  a14137a );
 a14139a <=( a14138a  and  a14133a );
 a14142a <=( A265  and  A233 );
 a14146a <=( (not A300)  and  (not A299) );
 a14147a <=( (not A267)  and  a14146a );
 a14148a <=( a14147a  and  a14142a );
 a14151a <=( A167  and  A168 );
 a14155a <=( A232  and  (not A201) );
 a14156a <=( (not A200)  and  a14155a );
 a14157a <=( a14156a  and  a14151a );
 a14160a <=( A265  and  A233 );
 a14164a <=( A299  and  A298 );
 a14165a <=( (not A267)  and  a14164a );
 a14166a <=( a14165a  and  a14160a );
 a14169a <=( A167  and  A168 );
 a14173a <=( A232  and  (not A201) );
 a14174a <=( (not A200)  and  a14173a );
 a14175a <=( a14174a  and  a14169a );
 a14178a <=( A265  and  A233 );
 a14182a <=( (not A299)  and  (not A298) );
 a14183a <=( (not A267)  and  a14182a );
 a14184a <=( a14183a  and  a14178a );
 a14187a <=( A167  and  A168 );
 a14191a <=( A232  and  (not A201) );
 a14192a <=( (not A200)  and  a14191a );
 a14193a <=( a14192a  and  a14187a );
 a14196a <=( A265  and  A233 );
 a14200a <=( (not A300)  and  (not A299) );
 a14201a <=( A266  and  a14200a );
 a14202a <=( a14201a  and  a14196a );
 a14205a <=( A167  and  A168 );
 a14209a <=( A232  and  (not A201) );
 a14210a <=( (not A200)  and  a14209a );
 a14211a <=( a14210a  and  a14205a );
 a14214a <=( A265  and  A233 );
 a14218a <=( A299  and  A298 );
 a14219a <=( A266  and  a14218a );
 a14220a <=( a14219a  and  a14214a );
 a14223a <=( A167  and  A168 );
 a14227a <=( A232  and  (not A201) );
 a14228a <=( (not A200)  and  a14227a );
 a14229a <=( a14228a  and  a14223a );
 a14232a <=( A265  and  A233 );
 a14236a <=( (not A299)  and  (not A298) );
 a14237a <=( A266  and  a14236a );
 a14238a <=( a14237a  and  a14232a );
 a14241a <=( A167  and  A168 );
 a14245a <=( A232  and  (not A201) );
 a14246a <=( (not A200)  and  a14245a );
 a14247a <=( a14246a  and  a14241a );
 a14250a <=( (not A265)  and  A233 );
 a14254a <=( (not A300)  and  (not A299) );
 a14255a <=( (not A266)  and  a14254a );
 a14256a <=( a14255a  and  a14250a );
 a14259a <=( A167  and  A168 );
 a14263a <=( A232  and  (not A201) );
 a14264a <=( (not A200)  and  a14263a );
 a14265a <=( a14264a  and  a14259a );
 a14268a <=( (not A265)  and  A233 );
 a14272a <=( A299  and  A298 );
 a14273a <=( (not A266)  and  a14272a );
 a14274a <=( a14273a  and  a14268a );
 a14277a <=( A167  and  A168 );
 a14281a <=( A232  and  (not A201) );
 a14282a <=( (not A200)  and  a14281a );
 a14283a <=( a14282a  and  a14277a );
 a14286a <=( (not A265)  and  A233 );
 a14290a <=( (not A299)  and  (not A298) );
 a14291a <=( (not A266)  and  a14290a );
 a14292a <=( a14291a  and  a14286a );
 a14295a <=( A167  and  A168 );
 a14299a <=( (not A232)  and  (not A201) );
 a14300a <=( (not A200)  and  a14299a );
 a14301a <=( a14300a  and  a14295a );
 a14304a <=( A298  and  A233 );
 a14308a <=( A301  and  A300 );
 a14309a <=( (not A299)  and  a14308a );
 a14310a <=( a14309a  and  a14304a );
 a14313a <=( A167  and  A168 );
 a14317a <=( (not A232)  and  (not A201) );
 a14318a <=( (not A200)  and  a14317a );
 a14319a <=( a14318a  and  a14313a );
 a14322a <=( A298  and  A233 );
 a14326a <=( A302  and  A300 );
 a14327a <=( (not A299)  and  a14326a );
 a14328a <=( a14327a  and  a14322a );
 a14331a <=( A167  and  A168 );
 a14335a <=( (not A232)  and  (not A201) );
 a14336a <=( (not A200)  and  a14335a );
 a14337a <=( a14336a  and  a14331a );
 a14340a <=( A265  and  A233 );
 a14344a <=( A268  and  A267 );
 a14345a <=( (not A266)  and  a14344a );
 a14346a <=( a14345a  and  a14340a );
 a14349a <=( A167  and  A168 );
 a14353a <=( (not A232)  and  (not A201) );
 a14354a <=( (not A200)  and  a14353a );
 a14355a <=( a14354a  and  a14349a );
 a14358a <=( A265  and  A233 );
 a14362a <=( A269  and  A267 );
 a14363a <=( (not A266)  and  a14362a );
 a14364a <=( a14363a  and  a14358a );
 a14367a <=( A167  and  A168 );
 a14371a <=( (not A233)  and  (not A201) );
 a14372a <=( (not A200)  and  a14371a );
 a14373a <=( a14372a  and  a14367a );
 a14376a <=( A265  and  (not A234) );
 a14380a <=( (not A300)  and  A298 );
 a14381a <=( A266  and  a14380a );
 a14382a <=( a14381a  and  a14376a );
 a14385a <=( A167  and  A168 );
 a14389a <=( (not A233)  and  (not A201) );
 a14390a <=( (not A200)  and  a14389a );
 a14391a <=( a14390a  and  a14385a );
 a14394a <=( A265  and  (not A234) );
 a14398a <=( A299  and  A298 );
 a14399a <=( A266  and  a14398a );
 a14400a <=( a14399a  and  a14394a );
 a14403a <=( A167  and  A168 );
 a14407a <=( (not A233)  and  (not A201) );
 a14408a <=( (not A200)  and  a14407a );
 a14409a <=( a14408a  and  a14403a );
 a14412a <=( A265  and  (not A234) );
 a14416a <=( (not A299)  and  (not A298) );
 a14417a <=( A266  and  a14416a );
 a14418a <=( a14417a  and  a14412a );
 a14421a <=( A167  and  A168 );
 a14425a <=( (not A233)  and  (not A201) );
 a14426a <=( (not A200)  and  a14425a );
 a14427a <=( a14426a  and  a14421a );
 a14430a <=( (not A266)  and  (not A234) );
 a14434a <=( (not A300)  and  A298 );
 a14435a <=( (not A267)  and  a14434a );
 a14436a <=( a14435a  and  a14430a );
 a14439a <=( A167  and  A168 );
 a14443a <=( (not A233)  and  (not A201) );
 a14444a <=( (not A200)  and  a14443a );
 a14445a <=( a14444a  and  a14439a );
 a14448a <=( (not A266)  and  (not A234) );
 a14452a <=( A299  and  A298 );
 a14453a <=( (not A267)  and  a14452a );
 a14454a <=( a14453a  and  a14448a );
 a14457a <=( A167  and  A168 );
 a14461a <=( (not A233)  and  (not A201) );
 a14462a <=( (not A200)  and  a14461a );
 a14463a <=( a14462a  and  a14457a );
 a14466a <=( (not A266)  and  (not A234) );
 a14470a <=( (not A299)  and  (not A298) );
 a14471a <=( (not A267)  and  a14470a );
 a14472a <=( a14471a  and  a14466a );
 a14475a <=( A167  and  A168 );
 a14479a <=( (not A233)  and  (not A201) );
 a14480a <=( (not A200)  and  a14479a );
 a14481a <=( a14480a  and  a14475a );
 a14484a <=( (not A265)  and  (not A234) );
 a14488a <=( (not A300)  and  A298 );
 a14489a <=( (not A266)  and  a14488a );
 a14490a <=( a14489a  and  a14484a );
 a14493a <=( A167  and  A168 );
 a14497a <=( (not A233)  and  (not A201) );
 a14498a <=( (not A200)  and  a14497a );
 a14499a <=( a14498a  and  a14493a );
 a14502a <=( (not A265)  and  (not A234) );
 a14506a <=( A299  and  A298 );
 a14507a <=( (not A266)  and  a14506a );
 a14508a <=( a14507a  and  a14502a );
 a14511a <=( A167  and  A168 );
 a14515a <=( (not A233)  and  (not A201) );
 a14516a <=( (not A200)  and  a14515a );
 a14517a <=( a14516a  and  a14511a );
 a14520a <=( (not A265)  and  (not A234) );
 a14524a <=( (not A299)  and  (not A298) );
 a14525a <=( (not A266)  and  a14524a );
 a14526a <=( a14525a  and  a14520a );
 a14529a <=( A167  and  A168 );
 a14533a <=( A232  and  (not A201) );
 a14534a <=( (not A200)  and  a14533a );
 a14535a <=( a14534a  and  a14529a );
 a14538a <=( A234  and  (not A233) );
 a14542a <=( A299  and  (not A298) );
 a14543a <=( A235  and  a14542a );
 a14544a <=( a14543a  and  a14538a );
 a14547a <=( A167  and  A168 );
 a14551a <=( A232  and  (not A201) );
 a14552a <=( (not A200)  and  a14551a );
 a14553a <=( a14552a  and  a14547a );
 a14556a <=( A234  and  (not A233) );
 a14560a <=( A266  and  (not A265) );
 a14561a <=( A235  and  a14560a );
 a14562a <=( a14561a  and  a14556a );
 a14565a <=( A167  and  A168 );
 a14569a <=( A232  and  (not A201) );
 a14570a <=( (not A200)  and  a14569a );
 a14571a <=( a14570a  and  a14565a );
 a14574a <=( A234  and  (not A233) );
 a14578a <=( A299  and  (not A298) );
 a14579a <=( A236  and  a14578a );
 a14580a <=( a14579a  and  a14574a );
 a14583a <=( A167  and  A168 );
 a14587a <=( A232  and  (not A201) );
 a14588a <=( (not A200)  and  a14587a );
 a14589a <=( a14588a  and  a14583a );
 a14592a <=( A234  and  (not A233) );
 a14596a <=( A266  and  (not A265) );
 a14597a <=( A236  and  a14596a );
 a14598a <=( a14597a  and  a14592a );
 a14601a <=( A167  and  A168 );
 a14605a <=( (not A232)  and  (not A201) );
 a14606a <=( (not A200)  and  a14605a );
 a14607a <=( a14606a  and  a14601a );
 a14610a <=( A265  and  (not A233) );
 a14614a <=( (not A300)  and  A298 );
 a14615a <=( A266  and  a14614a );
 a14616a <=( a14615a  and  a14610a );
 a14619a <=( A167  and  A168 );
 a14623a <=( (not A232)  and  (not A201) );
 a14624a <=( (not A200)  and  a14623a );
 a14625a <=( a14624a  and  a14619a );
 a14628a <=( A265  and  (not A233) );
 a14632a <=( A299  and  A298 );
 a14633a <=( A266  and  a14632a );
 a14634a <=( a14633a  and  a14628a );
 a14637a <=( A167  and  A168 );
 a14641a <=( (not A232)  and  (not A201) );
 a14642a <=( (not A200)  and  a14641a );
 a14643a <=( a14642a  and  a14637a );
 a14646a <=( A265  and  (not A233) );
 a14650a <=( (not A299)  and  (not A298) );
 a14651a <=( A266  and  a14650a );
 a14652a <=( a14651a  and  a14646a );
 a14655a <=( A167  and  A168 );
 a14659a <=( (not A232)  and  (not A201) );
 a14660a <=( (not A200)  and  a14659a );
 a14661a <=( a14660a  and  a14655a );
 a14664a <=( (not A266)  and  (not A233) );
 a14668a <=( (not A300)  and  A298 );
 a14669a <=( (not A267)  and  a14668a );
 a14670a <=( a14669a  and  a14664a );
 a14673a <=( A167  and  A168 );
 a14677a <=( (not A232)  and  (not A201) );
 a14678a <=( (not A200)  and  a14677a );
 a14679a <=( a14678a  and  a14673a );
 a14682a <=( (not A266)  and  (not A233) );
 a14686a <=( A299  and  A298 );
 a14687a <=( (not A267)  and  a14686a );
 a14688a <=( a14687a  and  a14682a );
 a14691a <=( A167  and  A168 );
 a14695a <=( (not A232)  and  (not A201) );
 a14696a <=( (not A200)  and  a14695a );
 a14697a <=( a14696a  and  a14691a );
 a14700a <=( (not A266)  and  (not A233) );
 a14704a <=( (not A299)  and  (not A298) );
 a14705a <=( (not A267)  and  a14704a );
 a14706a <=( a14705a  and  a14700a );
 a14709a <=( A167  and  A168 );
 a14713a <=( (not A232)  and  (not A201) );
 a14714a <=( (not A200)  and  a14713a );
 a14715a <=( a14714a  and  a14709a );
 a14718a <=( (not A265)  and  (not A233) );
 a14722a <=( (not A300)  and  A298 );
 a14723a <=( (not A266)  and  a14722a );
 a14724a <=( a14723a  and  a14718a );
 a14727a <=( A167  and  A168 );
 a14731a <=( (not A232)  and  (not A201) );
 a14732a <=( (not A200)  and  a14731a );
 a14733a <=( a14732a  and  a14727a );
 a14736a <=( (not A265)  and  (not A233) );
 a14740a <=( A299  and  A298 );
 a14741a <=( (not A266)  and  a14740a );
 a14742a <=( a14741a  and  a14736a );
 a14745a <=( A167  and  A168 );
 a14749a <=( (not A232)  and  (not A201) );
 a14750a <=( (not A200)  and  a14749a );
 a14751a <=( a14750a  and  a14745a );
 a14754a <=( (not A265)  and  (not A233) );
 a14758a <=( (not A299)  and  (not A298) );
 a14759a <=( (not A266)  and  a14758a );
 a14760a <=( a14759a  and  a14754a );
 a14763a <=( A167  and  A168 );
 a14767a <=( A232  and  (not A200) );
 a14768a <=( (not A199)  and  a14767a );
 a14769a <=( a14768a  and  a14763a );
 a14772a <=( A265  and  A233 );
 a14776a <=( (not A300)  and  (not A299) );
 a14777a <=( (not A267)  and  a14776a );
 a14778a <=( a14777a  and  a14772a );
 a14781a <=( A167  and  A168 );
 a14785a <=( A232  and  (not A200) );
 a14786a <=( (not A199)  and  a14785a );
 a14787a <=( a14786a  and  a14781a );
 a14790a <=( A265  and  A233 );
 a14794a <=( A299  and  A298 );
 a14795a <=( (not A267)  and  a14794a );
 a14796a <=( a14795a  and  a14790a );
 a14799a <=( A167  and  A168 );
 a14803a <=( A232  and  (not A200) );
 a14804a <=( (not A199)  and  a14803a );
 a14805a <=( a14804a  and  a14799a );
 a14808a <=( A265  and  A233 );
 a14812a <=( (not A299)  and  (not A298) );
 a14813a <=( (not A267)  and  a14812a );
 a14814a <=( a14813a  and  a14808a );
 a14817a <=( A167  and  A168 );
 a14821a <=( A232  and  (not A200) );
 a14822a <=( (not A199)  and  a14821a );
 a14823a <=( a14822a  and  a14817a );
 a14826a <=( A265  and  A233 );
 a14830a <=( (not A300)  and  (not A299) );
 a14831a <=( A266  and  a14830a );
 a14832a <=( a14831a  and  a14826a );
 a14835a <=( A167  and  A168 );
 a14839a <=( A232  and  (not A200) );
 a14840a <=( (not A199)  and  a14839a );
 a14841a <=( a14840a  and  a14835a );
 a14844a <=( A265  and  A233 );
 a14848a <=( A299  and  A298 );
 a14849a <=( A266  and  a14848a );
 a14850a <=( a14849a  and  a14844a );
 a14853a <=( A167  and  A168 );
 a14857a <=( A232  and  (not A200) );
 a14858a <=( (not A199)  and  a14857a );
 a14859a <=( a14858a  and  a14853a );
 a14862a <=( A265  and  A233 );
 a14866a <=( (not A299)  and  (not A298) );
 a14867a <=( A266  and  a14866a );
 a14868a <=( a14867a  and  a14862a );
 a14871a <=( A167  and  A168 );
 a14875a <=( A232  and  (not A200) );
 a14876a <=( (not A199)  and  a14875a );
 a14877a <=( a14876a  and  a14871a );
 a14880a <=( (not A265)  and  A233 );
 a14884a <=( (not A300)  and  (not A299) );
 a14885a <=( (not A266)  and  a14884a );
 a14886a <=( a14885a  and  a14880a );
 a14889a <=( A167  and  A168 );
 a14893a <=( A232  and  (not A200) );
 a14894a <=( (not A199)  and  a14893a );
 a14895a <=( a14894a  and  a14889a );
 a14898a <=( (not A265)  and  A233 );
 a14902a <=( A299  and  A298 );
 a14903a <=( (not A266)  and  a14902a );
 a14904a <=( a14903a  and  a14898a );
 a14907a <=( A167  and  A168 );
 a14911a <=( A232  and  (not A200) );
 a14912a <=( (not A199)  and  a14911a );
 a14913a <=( a14912a  and  a14907a );
 a14916a <=( (not A265)  and  A233 );
 a14920a <=( (not A299)  and  (not A298) );
 a14921a <=( (not A266)  and  a14920a );
 a14922a <=( a14921a  and  a14916a );
 a14925a <=( A167  and  A168 );
 a14929a <=( (not A232)  and  (not A200) );
 a14930a <=( (not A199)  and  a14929a );
 a14931a <=( a14930a  and  a14925a );
 a14934a <=( A298  and  A233 );
 a14938a <=( A301  and  A300 );
 a14939a <=( (not A299)  and  a14938a );
 a14940a <=( a14939a  and  a14934a );
 a14943a <=( A167  and  A168 );
 a14947a <=( (not A232)  and  (not A200) );
 a14948a <=( (not A199)  and  a14947a );
 a14949a <=( a14948a  and  a14943a );
 a14952a <=( A298  and  A233 );
 a14956a <=( A302  and  A300 );
 a14957a <=( (not A299)  and  a14956a );
 a14958a <=( a14957a  and  a14952a );
 a14961a <=( A167  and  A168 );
 a14965a <=( (not A232)  and  (not A200) );
 a14966a <=( (not A199)  and  a14965a );
 a14967a <=( a14966a  and  a14961a );
 a14970a <=( A265  and  A233 );
 a14974a <=( A268  and  A267 );
 a14975a <=( (not A266)  and  a14974a );
 a14976a <=( a14975a  and  a14970a );
 a14979a <=( A167  and  A168 );
 a14983a <=( (not A232)  and  (not A200) );
 a14984a <=( (not A199)  and  a14983a );
 a14985a <=( a14984a  and  a14979a );
 a14988a <=( A265  and  A233 );
 a14992a <=( A269  and  A267 );
 a14993a <=( (not A266)  and  a14992a );
 a14994a <=( a14993a  and  a14988a );
 a14997a <=( A167  and  A168 );
 a15001a <=( (not A233)  and  (not A200) );
 a15002a <=( (not A199)  and  a15001a );
 a15003a <=( a15002a  and  a14997a );
 a15006a <=( A265  and  (not A234) );
 a15010a <=( (not A300)  and  A298 );
 a15011a <=( A266  and  a15010a );
 a15012a <=( a15011a  and  a15006a );
 a15015a <=( A167  and  A168 );
 a15019a <=( (not A233)  and  (not A200) );
 a15020a <=( (not A199)  and  a15019a );
 a15021a <=( a15020a  and  a15015a );
 a15024a <=( A265  and  (not A234) );
 a15028a <=( A299  and  A298 );
 a15029a <=( A266  and  a15028a );
 a15030a <=( a15029a  and  a15024a );
 a15033a <=( A167  and  A168 );
 a15037a <=( (not A233)  and  (not A200) );
 a15038a <=( (not A199)  and  a15037a );
 a15039a <=( a15038a  and  a15033a );
 a15042a <=( A265  and  (not A234) );
 a15046a <=( (not A299)  and  (not A298) );
 a15047a <=( A266  and  a15046a );
 a15048a <=( a15047a  and  a15042a );
 a15051a <=( A167  and  A168 );
 a15055a <=( (not A233)  and  (not A200) );
 a15056a <=( (not A199)  and  a15055a );
 a15057a <=( a15056a  and  a15051a );
 a15060a <=( (not A266)  and  (not A234) );
 a15064a <=( (not A300)  and  A298 );
 a15065a <=( (not A267)  and  a15064a );
 a15066a <=( a15065a  and  a15060a );
 a15069a <=( A167  and  A168 );
 a15073a <=( (not A233)  and  (not A200) );
 a15074a <=( (not A199)  and  a15073a );
 a15075a <=( a15074a  and  a15069a );
 a15078a <=( (not A266)  and  (not A234) );
 a15082a <=( A299  and  A298 );
 a15083a <=( (not A267)  and  a15082a );
 a15084a <=( a15083a  and  a15078a );
 a15087a <=( A167  and  A168 );
 a15091a <=( (not A233)  and  (not A200) );
 a15092a <=( (not A199)  and  a15091a );
 a15093a <=( a15092a  and  a15087a );
 a15096a <=( (not A266)  and  (not A234) );
 a15100a <=( (not A299)  and  (not A298) );
 a15101a <=( (not A267)  and  a15100a );
 a15102a <=( a15101a  and  a15096a );
 a15105a <=( A167  and  A168 );
 a15109a <=( (not A233)  and  (not A200) );
 a15110a <=( (not A199)  and  a15109a );
 a15111a <=( a15110a  and  a15105a );
 a15114a <=( (not A265)  and  (not A234) );
 a15118a <=( (not A300)  and  A298 );
 a15119a <=( (not A266)  and  a15118a );
 a15120a <=( a15119a  and  a15114a );
 a15123a <=( A167  and  A168 );
 a15127a <=( (not A233)  and  (not A200) );
 a15128a <=( (not A199)  and  a15127a );
 a15129a <=( a15128a  and  a15123a );
 a15132a <=( (not A265)  and  (not A234) );
 a15136a <=( A299  and  A298 );
 a15137a <=( (not A266)  and  a15136a );
 a15138a <=( a15137a  and  a15132a );
 a15141a <=( A167  and  A168 );
 a15145a <=( (not A233)  and  (not A200) );
 a15146a <=( (not A199)  and  a15145a );
 a15147a <=( a15146a  and  a15141a );
 a15150a <=( (not A265)  and  (not A234) );
 a15154a <=( (not A299)  and  (not A298) );
 a15155a <=( (not A266)  and  a15154a );
 a15156a <=( a15155a  and  a15150a );
 a15159a <=( A167  and  A168 );
 a15163a <=( A232  and  (not A200) );
 a15164a <=( (not A199)  and  a15163a );
 a15165a <=( a15164a  and  a15159a );
 a15168a <=( A234  and  (not A233) );
 a15172a <=( A299  and  (not A298) );
 a15173a <=( A235  and  a15172a );
 a15174a <=( a15173a  and  a15168a );
 a15177a <=( A167  and  A168 );
 a15181a <=( A232  and  (not A200) );
 a15182a <=( (not A199)  and  a15181a );
 a15183a <=( a15182a  and  a15177a );
 a15186a <=( A234  and  (not A233) );
 a15190a <=( A266  and  (not A265) );
 a15191a <=( A235  and  a15190a );
 a15192a <=( a15191a  and  a15186a );
 a15195a <=( A167  and  A168 );
 a15199a <=( A232  and  (not A200) );
 a15200a <=( (not A199)  and  a15199a );
 a15201a <=( a15200a  and  a15195a );
 a15204a <=( A234  and  (not A233) );
 a15208a <=( A299  and  (not A298) );
 a15209a <=( A236  and  a15208a );
 a15210a <=( a15209a  and  a15204a );
 a15213a <=( A167  and  A168 );
 a15217a <=( A232  and  (not A200) );
 a15218a <=( (not A199)  and  a15217a );
 a15219a <=( a15218a  and  a15213a );
 a15222a <=( A234  and  (not A233) );
 a15226a <=( A266  and  (not A265) );
 a15227a <=( A236  and  a15226a );
 a15228a <=( a15227a  and  a15222a );
 a15231a <=( A167  and  A168 );
 a15235a <=( (not A232)  and  (not A200) );
 a15236a <=( (not A199)  and  a15235a );
 a15237a <=( a15236a  and  a15231a );
 a15240a <=( A265  and  (not A233) );
 a15244a <=( (not A300)  and  A298 );
 a15245a <=( A266  and  a15244a );
 a15246a <=( a15245a  and  a15240a );
 a15249a <=( A167  and  A168 );
 a15253a <=( (not A232)  and  (not A200) );
 a15254a <=( (not A199)  and  a15253a );
 a15255a <=( a15254a  and  a15249a );
 a15258a <=( A265  and  (not A233) );
 a15262a <=( A299  and  A298 );
 a15263a <=( A266  and  a15262a );
 a15264a <=( a15263a  and  a15258a );
 a15267a <=( A167  and  A168 );
 a15271a <=( (not A232)  and  (not A200) );
 a15272a <=( (not A199)  and  a15271a );
 a15273a <=( a15272a  and  a15267a );
 a15276a <=( A265  and  (not A233) );
 a15280a <=( (not A299)  and  (not A298) );
 a15281a <=( A266  and  a15280a );
 a15282a <=( a15281a  and  a15276a );
 a15285a <=( A167  and  A168 );
 a15289a <=( (not A232)  and  (not A200) );
 a15290a <=( (not A199)  and  a15289a );
 a15291a <=( a15290a  and  a15285a );
 a15294a <=( (not A266)  and  (not A233) );
 a15298a <=( (not A300)  and  A298 );
 a15299a <=( (not A267)  and  a15298a );
 a15300a <=( a15299a  and  a15294a );
 a15303a <=( A167  and  A168 );
 a15307a <=( (not A232)  and  (not A200) );
 a15308a <=( (not A199)  and  a15307a );
 a15309a <=( a15308a  and  a15303a );
 a15312a <=( (not A266)  and  (not A233) );
 a15316a <=( A299  and  A298 );
 a15317a <=( (not A267)  and  a15316a );
 a15318a <=( a15317a  and  a15312a );
 a15321a <=( A167  and  A168 );
 a15325a <=( (not A232)  and  (not A200) );
 a15326a <=( (not A199)  and  a15325a );
 a15327a <=( a15326a  and  a15321a );
 a15330a <=( (not A266)  and  (not A233) );
 a15334a <=( (not A299)  and  (not A298) );
 a15335a <=( (not A267)  and  a15334a );
 a15336a <=( a15335a  and  a15330a );
 a15339a <=( A167  and  A168 );
 a15343a <=( (not A232)  and  (not A200) );
 a15344a <=( (not A199)  and  a15343a );
 a15345a <=( a15344a  and  a15339a );
 a15348a <=( (not A265)  and  (not A233) );
 a15352a <=( (not A300)  and  A298 );
 a15353a <=( (not A266)  and  a15352a );
 a15354a <=( a15353a  and  a15348a );
 a15357a <=( A167  and  A168 );
 a15361a <=( (not A232)  and  (not A200) );
 a15362a <=( (not A199)  and  a15361a );
 a15363a <=( a15362a  and  a15357a );
 a15366a <=( (not A265)  and  (not A233) );
 a15370a <=( A299  and  A298 );
 a15371a <=( (not A266)  and  a15370a );
 a15372a <=( a15371a  and  a15366a );
 a15375a <=( A167  and  A168 );
 a15379a <=( (not A232)  and  (not A200) );
 a15380a <=( (not A199)  and  a15379a );
 a15381a <=( a15380a  and  a15375a );
 a15384a <=( (not A265)  and  (not A233) );
 a15388a <=( (not A299)  and  (not A298) );
 a15389a <=( (not A266)  and  a15388a );
 a15390a <=( a15389a  and  a15384a );
 a15393a <=( (not A168)  and  A170 );
 a15397a <=( (not A199)  and  A166 );
 a15398a <=( A167  and  a15397a );
 a15399a <=( a15398a  and  a15393a );
 a15402a <=( (not A232)  and  A200 );
 a15406a <=( A299  and  (not A298) );
 a15407a <=( A233  and  a15406a );
 a15408a <=( a15407a  and  a15402a );
 a15411a <=( (not A168)  and  A170 );
 a15415a <=( (not A199)  and  A166 );
 a15416a <=( A167  and  a15415a );
 a15417a <=( a15416a  and  a15411a );
 a15420a <=( (not A232)  and  A200 );
 a15424a <=( A266  and  (not A265) );
 a15425a <=( A233  and  a15424a );
 a15426a <=( a15425a  and  a15420a );
 a15429a <=( (not A168)  and  (not A170) );
 a15433a <=( (not A199)  and  (not A166) );
 a15434a <=( A167  and  a15433a );
 a15435a <=( a15434a  and  a15429a );
 a15438a <=( (not A232)  and  A200 );
 a15442a <=( A299  and  (not A298) );
 a15443a <=( A233  and  a15442a );
 a15444a <=( a15443a  and  a15438a );
 a15447a <=( (not A168)  and  (not A170) );
 a15451a <=( (not A199)  and  (not A166) );
 a15452a <=( A167  and  a15451a );
 a15453a <=( a15452a  and  a15447a );
 a15456a <=( (not A232)  and  A200 );
 a15460a <=( A266  and  (not A265) );
 a15461a <=( A233  and  a15460a );
 a15462a <=( a15461a  and  a15456a );
 a15465a <=( (not A168)  and  (not A170) );
 a15469a <=( (not A199)  and  A166 );
 a15470a <=( (not A167)  and  a15469a );
 a15471a <=( a15470a  and  a15465a );
 a15474a <=( (not A232)  and  A200 );
 a15478a <=( A299  and  (not A298) );
 a15479a <=( A233  and  a15478a );
 a15480a <=( a15479a  and  a15474a );
 a15483a <=( (not A168)  and  (not A170) );
 a15487a <=( (not A199)  and  A166 );
 a15488a <=( (not A167)  and  a15487a );
 a15489a <=( a15488a  and  a15483a );
 a15492a <=( (not A232)  and  A200 );
 a15496a <=( A266  and  (not A265) );
 a15497a <=( A233  and  a15496a );
 a15498a <=( a15497a  and  a15492a );
 a15501a <=( (not A168)  and  A169 );
 a15505a <=( (not A199)  and  (not A166) );
 a15506a <=( A167  and  a15505a );
 a15507a <=( a15506a  and  a15501a );
 a15510a <=( (not A232)  and  A200 );
 a15514a <=( A299  and  (not A298) );
 a15515a <=( A233  and  a15514a );
 a15516a <=( a15515a  and  a15510a );
 a15519a <=( (not A168)  and  A169 );
 a15523a <=( (not A199)  and  (not A166) );
 a15524a <=( A167  and  a15523a );
 a15525a <=( a15524a  and  a15519a );
 a15528a <=( (not A232)  and  A200 );
 a15532a <=( A266  and  (not A265) );
 a15533a <=( A233  and  a15532a );
 a15534a <=( a15533a  and  a15528a );
 a15537a <=( (not A168)  and  A169 );
 a15541a <=( (not A199)  and  A166 );
 a15542a <=( (not A167)  and  a15541a );
 a15543a <=( a15542a  and  a15537a );
 a15546a <=( (not A232)  and  A200 );
 a15550a <=( A299  and  (not A298) );
 a15551a <=( A233  and  a15550a );
 a15552a <=( a15551a  and  a15546a );
 a15555a <=( (not A168)  and  A169 );
 a15559a <=( (not A199)  and  A166 );
 a15560a <=( (not A167)  and  a15559a );
 a15561a <=( a15560a  and  a15555a );
 a15564a <=( (not A232)  and  A200 );
 a15568a <=( A266  and  (not A265) );
 a15569a <=( A233  and  a15568a );
 a15570a <=( a15569a  and  a15564a );
 a15573a <=( A169  and  (not A170) );
 a15577a <=( A199  and  A166 );
 a15578a <=( A167  and  a15577a );
 a15579a <=( a15578a  and  a15573a );
 a15582a <=( (not A232)  and  A200 );
 a15586a <=( A299  and  (not A298) );
 a15587a <=( A233  and  a15586a );
 a15588a <=( a15587a  and  a15582a );
 a15591a <=( A169  and  (not A170) );
 a15595a <=( A199  and  A166 );
 a15596a <=( A167  and  a15595a );
 a15597a <=( a15596a  and  a15591a );
 a15600a <=( (not A232)  and  A200 );
 a15604a <=( A266  and  (not A265) );
 a15605a <=( A233  and  a15604a );
 a15606a <=( a15605a  and  a15600a );
 a15609a <=( A169  and  (not A170) );
 a15613a <=( (not A200)  and  A166 );
 a15614a <=( A167  and  a15613a );
 a15615a <=( a15614a  and  a15609a );
 a15618a <=( (not A232)  and  (not A201) );
 a15622a <=( A299  and  (not A298) );
 a15623a <=( A233  and  a15622a );
 a15624a <=( a15623a  and  a15618a );
 a15627a <=( A169  and  (not A170) );
 a15631a <=( (not A200)  and  A166 );
 a15632a <=( A167  and  a15631a );
 a15633a <=( a15632a  and  a15627a );
 a15636a <=( (not A232)  and  (not A201) );
 a15640a <=( A266  and  (not A265) );
 a15641a <=( A233  and  a15640a );
 a15642a <=( a15641a  and  a15636a );
 a15645a <=( A169  and  (not A170) );
 a15649a <=( (not A199)  and  A166 );
 a15650a <=( A167  and  a15649a );
 a15651a <=( a15650a  and  a15645a );
 a15654a <=( (not A232)  and  (not A200) );
 a15658a <=( A299  and  (not A298) );
 a15659a <=( A233  and  a15658a );
 a15660a <=( a15659a  and  a15654a );
 a15663a <=( A169  and  (not A170) );
 a15667a <=( (not A199)  and  A166 );
 a15668a <=( A167  and  a15667a );
 a15669a <=( a15668a  and  a15663a );
 a15672a <=( (not A232)  and  (not A200) );
 a15676a <=( A266  and  (not A265) );
 a15677a <=( A233  and  a15676a );
 a15678a <=( a15677a  and  a15672a );
 a15681a <=( A169  and  (not A170) );
 a15685a <=( A199  and  (not A166) );
 a15686a <=( (not A167)  and  a15685a );
 a15687a <=( a15686a  and  a15681a );
 a15690a <=( (not A232)  and  A200 );
 a15694a <=( A299  and  (not A298) );
 a15695a <=( A233  and  a15694a );
 a15696a <=( a15695a  and  a15690a );
 a15699a <=( A169  and  (not A170) );
 a15703a <=( A199  and  (not A166) );
 a15704a <=( (not A167)  and  a15703a );
 a15705a <=( a15704a  and  a15699a );
 a15708a <=( (not A232)  and  A200 );
 a15712a <=( A266  and  (not A265) );
 a15713a <=( A233  and  a15712a );
 a15714a <=( a15713a  and  a15708a );
 a15717a <=( A169  and  (not A170) );
 a15721a <=( (not A200)  and  (not A166) );
 a15722a <=( (not A167)  and  a15721a );
 a15723a <=( a15722a  and  a15717a );
 a15726a <=( (not A232)  and  (not A201) );
 a15730a <=( A299  and  (not A298) );
 a15731a <=( A233  and  a15730a );
 a15732a <=( a15731a  and  a15726a );
 a15735a <=( A169  and  (not A170) );
 a15739a <=( (not A200)  and  (not A166) );
 a15740a <=( (not A167)  and  a15739a );
 a15741a <=( a15740a  and  a15735a );
 a15744a <=( (not A232)  and  (not A201) );
 a15748a <=( A266  and  (not A265) );
 a15749a <=( A233  and  a15748a );
 a15750a <=( a15749a  and  a15744a );
 a15753a <=( A169  and  (not A170) );
 a15757a <=( (not A199)  and  (not A166) );
 a15758a <=( (not A167)  and  a15757a );
 a15759a <=( a15758a  and  a15753a );
 a15762a <=( (not A232)  and  (not A200) );
 a15766a <=( A299  and  (not A298) );
 a15767a <=( A233  and  a15766a );
 a15768a <=( a15767a  and  a15762a );
 a15771a <=( A169  and  (not A170) );
 a15775a <=( (not A199)  and  (not A166) );
 a15776a <=( (not A167)  and  a15775a );
 a15777a <=( a15776a  and  a15771a );
 a15780a <=( (not A232)  and  (not A200) );
 a15784a <=( A266  and  (not A265) );
 a15785a <=( A233  and  a15784a );
 a15786a <=( a15785a  and  a15780a );
 a15789a <=( (not A168)  and  (not A169) );
 a15793a <=( (not A199)  and  A166 );
 a15794a <=( A167  and  a15793a );
 a15795a <=( a15794a  and  a15789a );
 a15798a <=( (not A232)  and  A200 );
 a15802a <=( A299  and  (not A298) );
 a15803a <=( A233  and  a15802a );
 a15804a <=( a15803a  and  a15798a );
 a15807a <=( (not A168)  and  (not A169) );
 a15811a <=( (not A199)  and  A166 );
 a15812a <=( A167  and  a15811a );
 a15813a <=( a15812a  and  a15807a );
 a15816a <=( (not A232)  and  A200 );
 a15820a <=( A266  and  (not A265) );
 a15821a <=( A233  and  a15820a );
 a15822a <=( a15821a  and  a15816a );
 a15825a <=( (not A169)  and  A170 );
 a15829a <=( A199  and  (not A166) );
 a15830a <=( A167  and  a15829a );
 a15831a <=( a15830a  and  a15825a );
 a15834a <=( (not A232)  and  A200 );
 a15838a <=( A299  and  (not A298) );
 a15839a <=( A233  and  a15838a );
 a15840a <=( a15839a  and  a15834a );
 a15843a <=( (not A169)  and  A170 );
 a15847a <=( A199  and  (not A166) );
 a15848a <=( A167  and  a15847a );
 a15849a <=( a15848a  and  a15843a );
 a15852a <=( (not A232)  and  A200 );
 a15856a <=( A266  and  (not A265) );
 a15857a <=( A233  and  a15856a );
 a15858a <=( a15857a  and  a15852a );
 a15861a <=( (not A169)  and  A170 );
 a15865a <=( (not A200)  and  (not A166) );
 a15866a <=( A167  and  a15865a );
 a15867a <=( a15866a  and  a15861a );
 a15870a <=( (not A232)  and  (not A201) );
 a15874a <=( A299  and  (not A298) );
 a15875a <=( A233  and  a15874a );
 a15876a <=( a15875a  and  a15870a );
 a15879a <=( (not A169)  and  A170 );
 a15883a <=( (not A200)  and  (not A166) );
 a15884a <=( A167  and  a15883a );
 a15885a <=( a15884a  and  a15879a );
 a15888a <=( (not A232)  and  (not A201) );
 a15892a <=( A266  and  (not A265) );
 a15893a <=( A233  and  a15892a );
 a15894a <=( a15893a  and  a15888a );
 a15897a <=( (not A169)  and  A170 );
 a15901a <=( (not A199)  and  (not A166) );
 a15902a <=( A167  and  a15901a );
 a15903a <=( a15902a  and  a15897a );
 a15906a <=( (not A232)  and  (not A200) );
 a15910a <=( A299  and  (not A298) );
 a15911a <=( A233  and  a15910a );
 a15912a <=( a15911a  and  a15906a );
 a15915a <=( (not A169)  and  A170 );
 a15919a <=( (not A199)  and  (not A166) );
 a15920a <=( A167  and  a15919a );
 a15921a <=( a15920a  and  a15915a );
 a15924a <=( (not A232)  and  (not A200) );
 a15928a <=( A266  and  (not A265) );
 a15929a <=( A233  and  a15928a );
 a15930a <=( a15929a  and  a15924a );
 a15933a <=( (not A169)  and  A170 );
 a15937a <=( A199  and  A166 );
 a15938a <=( (not A167)  and  a15937a );
 a15939a <=( a15938a  and  a15933a );
 a15942a <=( (not A232)  and  A200 );
 a15946a <=( A299  and  (not A298) );
 a15947a <=( A233  and  a15946a );
 a15948a <=( a15947a  and  a15942a );
 a15951a <=( (not A169)  and  A170 );
 a15955a <=( A199  and  A166 );
 a15956a <=( (not A167)  and  a15955a );
 a15957a <=( a15956a  and  a15951a );
 a15960a <=( (not A232)  and  A200 );
 a15964a <=( A266  and  (not A265) );
 a15965a <=( A233  and  a15964a );
 a15966a <=( a15965a  and  a15960a );
 a15969a <=( (not A169)  and  A170 );
 a15973a <=( (not A200)  and  A166 );
 a15974a <=( (not A167)  and  a15973a );
 a15975a <=( a15974a  and  a15969a );
 a15978a <=( (not A232)  and  (not A201) );
 a15982a <=( A299  and  (not A298) );
 a15983a <=( A233  and  a15982a );
 a15984a <=( a15983a  and  a15978a );
 a15987a <=( (not A169)  and  A170 );
 a15991a <=( (not A200)  and  A166 );
 a15992a <=( (not A167)  and  a15991a );
 a15993a <=( a15992a  and  a15987a );
 a15996a <=( (not A232)  and  (not A201) );
 a16000a <=( A266  and  (not A265) );
 a16001a <=( A233  and  a16000a );
 a16002a <=( a16001a  and  a15996a );
 a16005a <=( (not A169)  and  A170 );
 a16009a <=( (not A199)  and  A166 );
 a16010a <=( (not A167)  and  a16009a );
 a16011a <=( a16010a  and  a16005a );
 a16014a <=( (not A232)  and  (not A200) );
 a16018a <=( A299  and  (not A298) );
 a16019a <=( A233  and  a16018a );
 a16020a <=( a16019a  and  a16014a );
 a16023a <=( (not A169)  and  A170 );
 a16027a <=( (not A199)  and  A166 );
 a16028a <=( (not A167)  and  a16027a );
 a16029a <=( a16028a  and  a16023a );
 a16032a <=( (not A232)  and  (not A200) );
 a16036a <=( A266  and  (not A265) );
 a16037a <=( A233  and  a16036a );
 a16038a <=( a16037a  and  a16032a );
 a16041a <=( A166  and  A168 );
 a16045a <=( A232  and  A200 );
 a16046a <=( A199  and  a16045a );
 a16047a <=( a16046a  and  a16041a );
 a16051a <=( (not A268)  and  A265 );
 a16052a <=( A233  and  a16051a );
 a16056a <=( (not A300)  and  (not A299) );
 a16057a <=( (not A269)  and  a16056a );
 a16058a <=( a16057a  and  a16052a );
 a16061a <=( A166  and  A168 );
 a16065a <=( A232  and  A200 );
 a16066a <=( A199  and  a16065a );
 a16067a <=( a16066a  and  a16061a );
 a16071a <=( (not A268)  and  A265 );
 a16072a <=( A233  and  a16071a );
 a16076a <=( A299  and  A298 );
 a16077a <=( (not A269)  and  a16076a );
 a16078a <=( a16077a  and  a16072a );
 a16081a <=( A166  and  A168 );
 a16085a <=( A232  and  A200 );
 a16086a <=( A199  and  a16085a );
 a16087a <=( a16086a  and  a16081a );
 a16091a <=( (not A268)  and  A265 );
 a16092a <=( A233  and  a16091a );
 a16096a <=( (not A299)  and  (not A298) );
 a16097a <=( (not A269)  and  a16096a );
 a16098a <=( a16097a  and  a16092a );
 a16101a <=( A166  and  A168 );
 a16105a <=( A232  and  A200 );
 a16106a <=( A199  and  a16105a );
 a16107a <=( a16106a  and  a16101a );
 a16111a <=( (not A267)  and  A265 );
 a16112a <=( A233  and  a16111a );
 a16116a <=( (not A302)  and  (not A301) );
 a16117a <=( (not A299)  and  a16116a );
 a16118a <=( a16117a  and  a16112a );
 a16121a <=( A166  and  A168 );
 a16125a <=( A232  and  A200 );
 a16126a <=( A199  and  a16125a );
 a16127a <=( a16126a  and  a16121a );
 a16131a <=( A266  and  A265 );
 a16132a <=( A233  and  a16131a );
 a16136a <=( (not A302)  and  (not A301) );
 a16137a <=( (not A299)  and  a16136a );
 a16138a <=( a16137a  and  a16132a );
 a16141a <=( A166  and  A168 );
 a16145a <=( A232  and  A200 );
 a16146a <=( A199  and  a16145a );
 a16147a <=( a16146a  and  a16141a );
 a16151a <=( (not A266)  and  (not A265) );
 a16152a <=( A233  and  a16151a );
 a16156a <=( (not A302)  and  (not A301) );
 a16157a <=( (not A299)  and  a16156a );
 a16158a <=( a16157a  and  a16152a );
 a16161a <=( A166  and  A168 );
 a16165a <=( (not A233)  and  A200 );
 a16166a <=( A199  and  a16165a );
 a16167a <=( a16166a  and  a16161a );
 a16171a <=( A265  and  (not A236) );
 a16172a <=( (not A235)  and  a16171a );
 a16176a <=( (not A300)  and  A298 );
 a16177a <=( A266  and  a16176a );
 a16178a <=( a16177a  and  a16172a );
 a16181a <=( A166  and  A168 );
 a16185a <=( (not A233)  and  A200 );
 a16186a <=( A199  and  a16185a );
 a16187a <=( a16186a  and  a16181a );
 a16191a <=( A265  and  (not A236) );
 a16192a <=( (not A235)  and  a16191a );
 a16196a <=( A299  and  A298 );
 a16197a <=( A266  and  a16196a );
 a16198a <=( a16197a  and  a16192a );
 a16201a <=( A166  and  A168 );
 a16205a <=( (not A233)  and  A200 );
 a16206a <=( A199  and  a16205a );
 a16207a <=( a16206a  and  a16201a );
 a16211a <=( A265  and  (not A236) );
 a16212a <=( (not A235)  and  a16211a );
 a16216a <=( (not A299)  and  (not A298) );
 a16217a <=( A266  and  a16216a );
 a16218a <=( a16217a  and  a16212a );
 a16221a <=( A166  and  A168 );
 a16225a <=( (not A233)  and  A200 );
 a16226a <=( A199  and  a16225a );
 a16227a <=( a16226a  and  a16221a );
 a16231a <=( (not A266)  and  (not A236) );
 a16232a <=( (not A235)  and  a16231a );
 a16236a <=( (not A300)  and  A298 );
 a16237a <=( (not A267)  and  a16236a );
 a16238a <=( a16237a  and  a16232a );
 a16241a <=( A166  and  A168 );
 a16245a <=( (not A233)  and  A200 );
 a16246a <=( A199  and  a16245a );
 a16247a <=( a16246a  and  a16241a );
 a16251a <=( (not A266)  and  (not A236) );
 a16252a <=( (not A235)  and  a16251a );
 a16256a <=( A299  and  A298 );
 a16257a <=( (not A267)  and  a16256a );
 a16258a <=( a16257a  and  a16252a );
 a16261a <=( A166  and  A168 );
 a16265a <=( (not A233)  and  A200 );
 a16266a <=( A199  and  a16265a );
 a16267a <=( a16266a  and  a16261a );
 a16271a <=( (not A266)  and  (not A236) );
 a16272a <=( (not A235)  and  a16271a );
 a16276a <=( (not A299)  and  (not A298) );
 a16277a <=( (not A267)  and  a16276a );
 a16278a <=( a16277a  and  a16272a );
 a16281a <=( A166  and  A168 );
 a16285a <=( (not A233)  and  A200 );
 a16286a <=( A199  and  a16285a );
 a16287a <=( a16286a  and  a16281a );
 a16291a <=( (not A265)  and  (not A236) );
 a16292a <=( (not A235)  and  a16291a );
 a16296a <=( (not A300)  and  A298 );
 a16297a <=( (not A266)  and  a16296a );
 a16298a <=( a16297a  and  a16292a );
 a16301a <=( A166  and  A168 );
 a16305a <=( (not A233)  and  A200 );
 a16306a <=( A199  and  a16305a );
 a16307a <=( a16306a  and  a16301a );
 a16311a <=( (not A265)  and  (not A236) );
 a16312a <=( (not A235)  and  a16311a );
 a16316a <=( A299  and  A298 );
 a16317a <=( (not A266)  and  a16316a );
 a16318a <=( a16317a  and  a16312a );
 a16321a <=( A166  and  A168 );
 a16325a <=( (not A233)  and  A200 );
 a16326a <=( A199  and  a16325a );
 a16327a <=( a16326a  and  a16321a );
 a16331a <=( (not A265)  and  (not A236) );
 a16332a <=( (not A235)  and  a16331a );
 a16336a <=( (not A299)  and  (not A298) );
 a16337a <=( (not A266)  and  a16336a );
 a16338a <=( a16337a  and  a16332a );
 a16341a <=( A166  and  A168 );
 a16345a <=( (not A233)  and  A200 );
 a16346a <=( A199  and  a16345a );
 a16347a <=( a16346a  and  a16341a );
 a16351a <=( A266  and  A265 );
 a16352a <=( (not A234)  and  a16351a );
 a16356a <=( (not A302)  and  (not A301) );
 a16357a <=( A298  and  a16356a );
 a16358a <=( a16357a  and  a16352a );
 a16361a <=( A166  and  A168 );
 a16365a <=( (not A233)  and  A200 );
 a16366a <=( A199  and  a16365a );
 a16367a <=( a16366a  and  a16361a );
 a16371a <=( (not A268)  and  (not A266) );
 a16372a <=( (not A234)  and  a16371a );
 a16376a <=( (not A300)  and  A298 );
 a16377a <=( (not A269)  and  a16376a );
 a16378a <=( a16377a  and  a16372a );
 a16381a <=( A166  and  A168 );
 a16385a <=( (not A233)  and  A200 );
 a16386a <=( A199  and  a16385a );
 a16387a <=( a16386a  and  a16381a );
 a16391a <=( (not A268)  and  (not A266) );
 a16392a <=( (not A234)  and  a16391a );
 a16396a <=( A299  and  A298 );
 a16397a <=( (not A269)  and  a16396a );
 a16398a <=( a16397a  and  a16392a );
 a16401a <=( A166  and  A168 );
 a16405a <=( (not A233)  and  A200 );
 a16406a <=( A199  and  a16405a );
 a16407a <=( a16406a  and  a16401a );
 a16411a <=( (not A268)  and  (not A266) );
 a16412a <=( (not A234)  and  a16411a );
 a16416a <=( (not A299)  and  (not A298) );
 a16417a <=( (not A269)  and  a16416a );
 a16418a <=( a16417a  and  a16412a );
 a16421a <=( A166  and  A168 );
 a16425a <=( (not A233)  and  A200 );
 a16426a <=( A199  and  a16425a );
 a16427a <=( a16426a  and  a16421a );
 a16431a <=( (not A267)  and  (not A266) );
 a16432a <=( (not A234)  and  a16431a );
 a16436a <=( (not A302)  and  (not A301) );
 a16437a <=( A298  and  a16436a );
 a16438a <=( a16437a  and  a16432a );
 a16441a <=( A166  and  A168 );
 a16445a <=( (not A233)  and  A200 );
 a16446a <=( A199  and  a16445a );
 a16447a <=( a16446a  and  a16441a );
 a16451a <=( (not A266)  and  (not A265) );
 a16452a <=( (not A234)  and  a16451a );
 a16456a <=( (not A302)  and  (not A301) );
 a16457a <=( A298  and  a16456a );
 a16458a <=( a16457a  and  a16452a );
 a16461a <=( A166  and  A168 );
 a16465a <=( (not A232)  and  A200 );
 a16466a <=( A199  and  a16465a );
 a16467a <=( a16466a  and  a16461a );
 a16471a <=( A266  and  A265 );
 a16472a <=( (not A233)  and  a16471a );
 a16476a <=( (not A302)  and  (not A301) );
 a16477a <=( A298  and  a16476a );
 a16478a <=( a16477a  and  a16472a );
 a16481a <=( A166  and  A168 );
 a16485a <=( (not A232)  and  A200 );
 a16486a <=( A199  and  a16485a );
 a16487a <=( a16486a  and  a16481a );
 a16491a <=( (not A268)  and  (not A266) );
 a16492a <=( (not A233)  and  a16491a );
 a16496a <=( (not A300)  and  A298 );
 a16497a <=( (not A269)  and  a16496a );
 a16498a <=( a16497a  and  a16492a );
 a16501a <=( A166  and  A168 );
 a16505a <=( (not A232)  and  A200 );
 a16506a <=( A199  and  a16505a );
 a16507a <=( a16506a  and  a16501a );
 a16511a <=( (not A268)  and  (not A266) );
 a16512a <=( (not A233)  and  a16511a );
 a16516a <=( A299  and  A298 );
 a16517a <=( (not A269)  and  a16516a );
 a16518a <=( a16517a  and  a16512a );
 a16521a <=( A166  and  A168 );
 a16525a <=( (not A232)  and  A200 );
 a16526a <=( A199  and  a16525a );
 a16527a <=( a16526a  and  a16521a );
 a16531a <=( (not A268)  and  (not A266) );
 a16532a <=( (not A233)  and  a16531a );
 a16536a <=( (not A299)  and  (not A298) );
 a16537a <=( (not A269)  and  a16536a );
 a16538a <=( a16537a  and  a16532a );
 a16541a <=( A166  and  A168 );
 a16545a <=( (not A232)  and  A200 );
 a16546a <=( A199  and  a16545a );
 a16547a <=( a16546a  and  a16541a );
 a16551a <=( (not A267)  and  (not A266) );
 a16552a <=( (not A233)  and  a16551a );
 a16556a <=( (not A302)  and  (not A301) );
 a16557a <=( A298  and  a16556a );
 a16558a <=( a16557a  and  a16552a );
 a16561a <=( A166  and  A168 );
 a16565a <=( (not A232)  and  A200 );
 a16566a <=( A199  and  a16565a );
 a16567a <=( a16566a  and  a16561a );
 a16571a <=( (not A266)  and  (not A265) );
 a16572a <=( (not A233)  and  a16571a );
 a16576a <=( (not A302)  and  (not A301) );
 a16577a <=( A298  and  a16576a );
 a16578a <=( a16577a  and  a16572a );
 a16581a <=( A166  and  A168 );
 a16585a <=( (not A203)  and  (not A202) );
 a16586a <=( (not A200)  and  a16585a );
 a16587a <=( a16586a  and  a16581a );
 a16591a <=( A265  and  A233 );
 a16592a <=( A232  and  a16591a );
 a16596a <=( (not A300)  and  (not A299) );
 a16597a <=( (not A267)  and  a16596a );
 a16598a <=( a16597a  and  a16592a );
 a16601a <=( A166  and  A168 );
 a16605a <=( (not A203)  and  (not A202) );
 a16606a <=( (not A200)  and  a16605a );
 a16607a <=( a16606a  and  a16601a );
 a16611a <=( A265  and  A233 );
 a16612a <=( A232  and  a16611a );
 a16616a <=( A299  and  A298 );
 a16617a <=( (not A267)  and  a16616a );
 a16618a <=( a16617a  and  a16612a );
 a16621a <=( A166  and  A168 );
 a16625a <=( (not A203)  and  (not A202) );
 a16626a <=( (not A200)  and  a16625a );
 a16627a <=( a16626a  and  a16621a );
 a16631a <=( A265  and  A233 );
 a16632a <=( A232  and  a16631a );
 a16636a <=( (not A299)  and  (not A298) );
 a16637a <=( (not A267)  and  a16636a );
 a16638a <=( a16637a  and  a16632a );
 a16641a <=( A166  and  A168 );
 a16645a <=( (not A203)  and  (not A202) );
 a16646a <=( (not A200)  and  a16645a );
 a16647a <=( a16646a  and  a16641a );
 a16651a <=( A265  and  A233 );
 a16652a <=( A232  and  a16651a );
 a16656a <=( (not A300)  and  (not A299) );
 a16657a <=( A266  and  a16656a );
 a16658a <=( a16657a  and  a16652a );
 a16661a <=( A166  and  A168 );
 a16665a <=( (not A203)  and  (not A202) );
 a16666a <=( (not A200)  and  a16665a );
 a16667a <=( a16666a  and  a16661a );
 a16671a <=( A265  and  A233 );
 a16672a <=( A232  and  a16671a );
 a16676a <=( A299  and  A298 );
 a16677a <=( A266  and  a16676a );
 a16678a <=( a16677a  and  a16672a );
 a16681a <=( A166  and  A168 );
 a16685a <=( (not A203)  and  (not A202) );
 a16686a <=( (not A200)  and  a16685a );
 a16687a <=( a16686a  and  a16681a );
 a16691a <=( A265  and  A233 );
 a16692a <=( A232  and  a16691a );
 a16696a <=( (not A299)  and  (not A298) );
 a16697a <=( A266  and  a16696a );
 a16698a <=( a16697a  and  a16692a );
 a16701a <=( A166  and  A168 );
 a16705a <=( (not A203)  and  (not A202) );
 a16706a <=( (not A200)  and  a16705a );
 a16707a <=( a16706a  and  a16701a );
 a16711a <=( (not A265)  and  A233 );
 a16712a <=( A232  and  a16711a );
 a16716a <=( (not A300)  and  (not A299) );
 a16717a <=( (not A266)  and  a16716a );
 a16718a <=( a16717a  and  a16712a );
 a16721a <=( A166  and  A168 );
 a16725a <=( (not A203)  and  (not A202) );
 a16726a <=( (not A200)  and  a16725a );
 a16727a <=( a16726a  and  a16721a );
 a16731a <=( (not A265)  and  A233 );
 a16732a <=( A232  and  a16731a );
 a16736a <=( A299  and  A298 );
 a16737a <=( (not A266)  and  a16736a );
 a16738a <=( a16737a  and  a16732a );
 a16741a <=( A166  and  A168 );
 a16745a <=( (not A203)  and  (not A202) );
 a16746a <=( (not A200)  and  a16745a );
 a16747a <=( a16746a  and  a16741a );
 a16751a <=( (not A265)  and  A233 );
 a16752a <=( A232  and  a16751a );
 a16756a <=( (not A299)  and  (not A298) );
 a16757a <=( (not A266)  and  a16756a );
 a16758a <=( a16757a  and  a16752a );
 a16761a <=( A166  and  A168 );
 a16765a <=( (not A203)  and  (not A202) );
 a16766a <=( (not A200)  and  a16765a );
 a16767a <=( a16766a  and  a16761a );
 a16771a <=( A298  and  A233 );
 a16772a <=( (not A232)  and  a16771a );
 a16776a <=( A301  and  A300 );
 a16777a <=( (not A299)  and  a16776a );
 a16778a <=( a16777a  and  a16772a );
 a16781a <=( A166  and  A168 );
 a16785a <=( (not A203)  and  (not A202) );
 a16786a <=( (not A200)  and  a16785a );
 a16787a <=( a16786a  and  a16781a );
 a16791a <=( A298  and  A233 );
 a16792a <=( (not A232)  and  a16791a );
 a16796a <=( A302  and  A300 );
 a16797a <=( (not A299)  and  a16796a );
 a16798a <=( a16797a  and  a16792a );
 a16801a <=( A166  and  A168 );
 a16805a <=( (not A203)  and  (not A202) );
 a16806a <=( (not A200)  and  a16805a );
 a16807a <=( a16806a  and  a16801a );
 a16811a <=( A265  and  A233 );
 a16812a <=( (not A232)  and  a16811a );
 a16816a <=( A268  and  A267 );
 a16817a <=( (not A266)  and  a16816a );
 a16818a <=( a16817a  and  a16812a );
 a16821a <=( A166  and  A168 );
 a16825a <=( (not A203)  and  (not A202) );
 a16826a <=( (not A200)  and  a16825a );
 a16827a <=( a16826a  and  a16821a );
 a16831a <=( A265  and  A233 );
 a16832a <=( (not A232)  and  a16831a );
 a16836a <=( A269  and  A267 );
 a16837a <=( (not A266)  and  a16836a );
 a16838a <=( a16837a  and  a16832a );
 a16841a <=( A166  and  A168 );
 a16845a <=( (not A203)  and  (not A202) );
 a16846a <=( (not A200)  and  a16845a );
 a16847a <=( a16846a  and  a16841a );
 a16851a <=( A265  and  (not A234) );
 a16852a <=( (not A233)  and  a16851a );
 a16856a <=( (not A300)  and  A298 );
 a16857a <=( A266  and  a16856a );
 a16858a <=( a16857a  and  a16852a );
 a16861a <=( A166  and  A168 );
 a16865a <=( (not A203)  and  (not A202) );
 a16866a <=( (not A200)  and  a16865a );
 a16867a <=( a16866a  and  a16861a );
 a16871a <=( A265  and  (not A234) );
 a16872a <=( (not A233)  and  a16871a );
 a16876a <=( A299  and  A298 );
 a16877a <=( A266  and  a16876a );
 a16878a <=( a16877a  and  a16872a );
 a16881a <=( A166  and  A168 );
 a16885a <=( (not A203)  and  (not A202) );
 a16886a <=( (not A200)  and  a16885a );
 a16887a <=( a16886a  and  a16881a );
 a16891a <=( A265  and  (not A234) );
 a16892a <=( (not A233)  and  a16891a );
 a16896a <=( (not A299)  and  (not A298) );
 a16897a <=( A266  and  a16896a );
 a16898a <=( a16897a  and  a16892a );
 a16901a <=( A166  and  A168 );
 a16905a <=( (not A203)  and  (not A202) );
 a16906a <=( (not A200)  and  a16905a );
 a16907a <=( a16906a  and  a16901a );
 a16911a <=( (not A266)  and  (not A234) );
 a16912a <=( (not A233)  and  a16911a );
 a16916a <=( (not A300)  and  A298 );
 a16917a <=( (not A267)  and  a16916a );
 a16918a <=( a16917a  and  a16912a );
 a16921a <=( A166  and  A168 );
 a16925a <=( (not A203)  and  (not A202) );
 a16926a <=( (not A200)  and  a16925a );
 a16927a <=( a16926a  and  a16921a );
 a16931a <=( (not A266)  and  (not A234) );
 a16932a <=( (not A233)  and  a16931a );
 a16936a <=( A299  and  A298 );
 a16937a <=( (not A267)  and  a16936a );
 a16938a <=( a16937a  and  a16932a );
 a16941a <=( A166  and  A168 );
 a16945a <=( (not A203)  and  (not A202) );
 a16946a <=( (not A200)  and  a16945a );
 a16947a <=( a16946a  and  a16941a );
 a16951a <=( (not A266)  and  (not A234) );
 a16952a <=( (not A233)  and  a16951a );
 a16956a <=( (not A299)  and  (not A298) );
 a16957a <=( (not A267)  and  a16956a );
 a16958a <=( a16957a  and  a16952a );
 a16961a <=( A166  and  A168 );
 a16965a <=( (not A203)  and  (not A202) );
 a16966a <=( (not A200)  and  a16965a );
 a16967a <=( a16966a  and  a16961a );
 a16971a <=( (not A265)  and  (not A234) );
 a16972a <=( (not A233)  and  a16971a );
 a16976a <=( (not A300)  and  A298 );
 a16977a <=( (not A266)  and  a16976a );
 a16978a <=( a16977a  and  a16972a );
 a16981a <=( A166  and  A168 );
 a16985a <=( (not A203)  and  (not A202) );
 a16986a <=( (not A200)  and  a16985a );
 a16987a <=( a16986a  and  a16981a );
 a16991a <=( (not A265)  and  (not A234) );
 a16992a <=( (not A233)  and  a16991a );
 a16996a <=( A299  and  A298 );
 a16997a <=( (not A266)  and  a16996a );
 a16998a <=( a16997a  and  a16992a );
 a17001a <=( A166  and  A168 );
 a17005a <=( (not A203)  and  (not A202) );
 a17006a <=( (not A200)  and  a17005a );
 a17007a <=( a17006a  and  a17001a );
 a17011a <=( (not A265)  and  (not A234) );
 a17012a <=( (not A233)  and  a17011a );
 a17016a <=( (not A299)  and  (not A298) );
 a17017a <=( (not A266)  and  a17016a );
 a17018a <=( a17017a  and  a17012a );
 a17021a <=( A166  and  A168 );
 a17025a <=( (not A203)  and  (not A202) );
 a17026a <=( (not A200)  and  a17025a );
 a17027a <=( a17026a  and  a17021a );
 a17031a <=( A234  and  (not A233) );
 a17032a <=( A232  and  a17031a );
 a17036a <=( A299  and  (not A298) );
 a17037a <=( A235  and  a17036a );
 a17038a <=( a17037a  and  a17032a );
 a17041a <=( A166  and  A168 );
 a17045a <=( (not A203)  and  (not A202) );
 a17046a <=( (not A200)  and  a17045a );
 a17047a <=( a17046a  and  a17041a );
 a17051a <=( A234  and  (not A233) );
 a17052a <=( A232  and  a17051a );
 a17056a <=( A266  and  (not A265) );
 a17057a <=( A235  and  a17056a );
 a17058a <=( a17057a  and  a17052a );
 a17061a <=( A166  and  A168 );
 a17065a <=( (not A203)  and  (not A202) );
 a17066a <=( (not A200)  and  a17065a );
 a17067a <=( a17066a  and  a17061a );
 a17071a <=( A234  and  (not A233) );
 a17072a <=( A232  and  a17071a );
 a17076a <=( A299  and  (not A298) );
 a17077a <=( A236  and  a17076a );
 a17078a <=( a17077a  and  a17072a );
 a17081a <=( A166  and  A168 );
 a17085a <=( (not A203)  and  (not A202) );
 a17086a <=( (not A200)  and  a17085a );
 a17087a <=( a17086a  and  a17081a );
 a17091a <=( A234  and  (not A233) );
 a17092a <=( A232  and  a17091a );
 a17096a <=( A266  and  (not A265) );
 a17097a <=( A236  and  a17096a );
 a17098a <=( a17097a  and  a17092a );
 a17101a <=( A166  and  A168 );
 a17105a <=( (not A203)  and  (not A202) );
 a17106a <=( (not A200)  and  a17105a );
 a17107a <=( a17106a  and  a17101a );
 a17111a <=( A265  and  (not A233) );
 a17112a <=( (not A232)  and  a17111a );
 a17116a <=( (not A300)  and  A298 );
 a17117a <=( A266  and  a17116a );
 a17118a <=( a17117a  and  a17112a );
 a17121a <=( A166  and  A168 );
 a17125a <=( (not A203)  and  (not A202) );
 a17126a <=( (not A200)  and  a17125a );
 a17127a <=( a17126a  and  a17121a );
 a17131a <=( A265  and  (not A233) );
 a17132a <=( (not A232)  and  a17131a );
 a17136a <=( A299  and  A298 );
 a17137a <=( A266  and  a17136a );
 a17138a <=( a17137a  and  a17132a );
 a17141a <=( A166  and  A168 );
 a17145a <=( (not A203)  and  (not A202) );
 a17146a <=( (not A200)  and  a17145a );
 a17147a <=( a17146a  and  a17141a );
 a17151a <=( A265  and  (not A233) );
 a17152a <=( (not A232)  and  a17151a );
 a17156a <=( (not A299)  and  (not A298) );
 a17157a <=( A266  and  a17156a );
 a17158a <=( a17157a  and  a17152a );
 a17161a <=( A166  and  A168 );
 a17165a <=( (not A203)  and  (not A202) );
 a17166a <=( (not A200)  and  a17165a );
 a17167a <=( a17166a  and  a17161a );
 a17171a <=( (not A266)  and  (not A233) );
 a17172a <=( (not A232)  and  a17171a );
 a17176a <=( (not A300)  and  A298 );
 a17177a <=( (not A267)  and  a17176a );
 a17178a <=( a17177a  and  a17172a );
 a17181a <=( A166  and  A168 );
 a17185a <=( (not A203)  and  (not A202) );
 a17186a <=( (not A200)  and  a17185a );
 a17187a <=( a17186a  and  a17181a );
 a17191a <=( (not A266)  and  (not A233) );
 a17192a <=( (not A232)  and  a17191a );
 a17196a <=( A299  and  A298 );
 a17197a <=( (not A267)  and  a17196a );
 a17198a <=( a17197a  and  a17192a );
 a17201a <=( A166  and  A168 );
 a17205a <=( (not A203)  and  (not A202) );
 a17206a <=( (not A200)  and  a17205a );
 a17207a <=( a17206a  and  a17201a );
 a17211a <=( (not A266)  and  (not A233) );
 a17212a <=( (not A232)  and  a17211a );
 a17216a <=( (not A299)  and  (not A298) );
 a17217a <=( (not A267)  and  a17216a );
 a17218a <=( a17217a  and  a17212a );
 a17221a <=( A166  and  A168 );
 a17225a <=( (not A203)  and  (not A202) );
 a17226a <=( (not A200)  and  a17225a );
 a17227a <=( a17226a  and  a17221a );
 a17231a <=( (not A265)  and  (not A233) );
 a17232a <=( (not A232)  and  a17231a );
 a17236a <=( (not A300)  and  A298 );
 a17237a <=( (not A266)  and  a17236a );
 a17238a <=( a17237a  and  a17232a );
 a17241a <=( A166  and  A168 );
 a17245a <=( (not A203)  and  (not A202) );
 a17246a <=( (not A200)  and  a17245a );
 a17247a <=( a17246a  and  a17241a );
 a17251a <=( (not A265)  and  (not A233) );
 a17252a <=( (not A232)  and  a17251a );
 a17256a <=( A299  and  A298 );
 a17257a <=( (not A266)  and  a17256a );
 a17258a <=( a17257a  and  a17252a );
 a17261a <=( A166  and  A168 );
 a17265a <=( (not A203)  and  (not A202) );
 a17266a <=( (not A200)  and  a17265a );
 a17267a <=( a17266a  and  a17261a );
 a17271a <=( (not A265)  and  (not A233) );
 a17272a <=( (not A232)  and  a17271a );
 a17276a <=( (not A299)  and  (not A298) );
 a17277a <=( (not A266)  and  a17276a );
 a17278a <=( a17277a  and  a17272a );
 a17281a <=( A166  and  A168 );
 a17285a <=( A232  and  (not A201) );
 a17286a <=( (not A200)  and  a17285a );
 a17287a <=( a17286a  and  a17281a );
 a17291a <=( (not A268)  and  A265 );
 a17292a <=( A233  and  a17291a );
 a17296a <=( (not A300)  and  (not A299) );
 a17297a <=( (not A269)  and  a17296a );
 a17298a <=( a17297a  and  a17292a );
 a17301a <=( A166  and  A168 );
 a17305a <=( A232  and  (not A201) );
 a17306a <=( (not A200)  and  a17305a );
 a17307a <=( a17306a  and  a17301a );
 a17311a <=( (not A268)  and  A265 );
 a17312a <=( A233  and  a17311a );
 a17316a <=( A299  and  A298 );
 a17317a <=( (not A269)  and  a17316a );
 a17318a <=( a17317a  and  a17312a );
 a17321a <=( A166  and  A168 );
 a17325a <=( A232  and  (not A201) );
 a17326a <=( (not A200)  and  a17325a );
 a17327a <=( a17326a  and  a17321a );
 a17331a <=( (not A268)  and  A265 );
 a17332a <=( A233  and  a17331a );
 a17336a <=( (not A299)  and  (not A298) );
 a17337a <=( (not A269)  and  a17336a );
 a17338a <=( a17337a  and  a17332a );
 a17341a <=( A166  and  A168 );
 a17345a <=( A232  and  (not A201) );
 a17346a <=( (not A200)  and  a17345a );
 a17347a <=( a17346a  and  a17341a );
 a17351a <=( (not A267)  and  A265 );
 a17352a <=( A233  and  a17351a );
 a17356a <=( (not A302)  and  (not A301) );
 a17357a <=( (not A299)  and  a17356a );
 a17358a <=( a17357a  and  a17352a );
 a17361a <=( A166  and  A168 );
 a17365a <=( A232  and  (not A201) );
 a17366a <=( (not A200)  and  a17365a );
 a17367a <=( a17366a  and  a17361a );
 a17371a <=( A266  and  A265 );
 a17372a <=( A233  and  a17371a );
 a17376a <=( (not A302)  and  (not A301) );
 a17377a <=( (not A299)  and  a17376a );
 a17378a <=( a17377a  and  a17372a );
 a17381a <=( A166  and  A168 );
 a17385a <=( A232  and  (not A201) );
 a17386a <=( (not A200)  and  a17385a );
 a17387a <=( a17386a  and  a17381a );
 a17391a <=( (not A266)  and  (not A265) );
 a17392a <=( A233  and  a17391a );
 a17396a <=( (not A302)  and  (not A301) );
 a17397a <=( (not A299)  and  a17396a );
 a17398a <=( a17397a  and  a17392a );
 a17401a <=( A166  and  A168 );
 a17405a <=( (not A233)  and  (not A201) );
 a17406a <=( (not A200)  and  a17405a );
 a17407a <=( a17406a  and  a17401a );
 a17411a <=( A265  and  (not A236) );
 a17412a <=( (not A235)  and  a17411a );
 a17416a <=( (not A300)  and  A298 );
 a17417a <=( A266  and  a17416a );
 a17418a <=( a17417a  and  a17412a );
 a17421a <=( A166  and  A168 );
 a17425a <=( (not A233)  and  (not A201) );
 a17426a <=( (not A200)  and  a17425a );
 a17427a <=( a17426a  and  a17421a );
 a17431a <=( A265  and  (not A236) );
 a17432a <=( (not A235)  and  a17431a );
 a17436a <=( A299  and  A298 );
 a17437a <=( A266  and  a17436a );
 a17438a <=( a17437a  and  a17432a );
 a17441a <=( A166  and  A168 );
 a17445a <=( (not A233)  and  (not A201) );
 a17446a <=( (not A200)  and  a17445a );
 a17447a <=( a17446a  and  a17441a );
 a17451a <=( A265  and  (not A236) );
 a17452a <=( (not A235)  and  a17451a );
 a17456a <=( (not A299)  and  (not A298) );
 a17457a <=( A266  and  a17456a );
 a17458a <=( a17457a  and  a17452a );
 a17461a <=( A166  and  A168 );
 a17465a <=( (not A233)  and  (not A201) );
 a17466a <=( (not A200)  and  a17465a );
 a17467a <=( a17466a  and  a17461a );
 a17471a <=( (not A266)  and  (not A236) );
 a17472a <=( (not A235)  and  a17471a );
 a17476a <=( (not A300)  and  A298 );
 a17477a <=( (not A267)  and  a17476a );
 a17478a <=( a17477a  and  a17472a );
 a17481a <=( A166  and  A168 );
 a17485a <=( (not A233)  and  (not A201) );
 a17486a <=( (not A200)  and  a17485a );
 a17487a <=( a17486a  and  a17481a );
 a17491a <=( (not A266)  and  (not A236) );
 a17492a <=( (not A235)  and  a17491a );
 a17496a <=( A299  and  A298 );
 a17497a <=( (not A267)  and  a17496a );
 a17498a <=( a17497a  and  a17492a );
 a17501a <=( A166  and  A168 );
 a17505a <=( (not A233)  and  (not A201) );
 a17506a <=( (not A200)  and  a17505a );
 a17507a <=( a17506a  and  a17501a );
 a17511a <=( (not A266)  and  (not A236) );
 a17512a <=( (not A235)  and  a17511a );
 a17516a <=( (not A299)  and  (not A298) );
 a17517a <=( (not A267)  and  a17516a );
 a17518a <=( a17517a  and  a17512a );
 a17521a <=( A166  and  A168 );
 a17525a <=( (not A233)  and  (not A201) );
 a17526a <=( (not A200)  and  a17525a );
 a17527a <=( a17526a  and  a17521a );
 a17531a <=( (not A265)  and  (not A236) );
 a17532a <=( (not A235)  and  a17531a );
 a17536a <=( (not A300)  and  A298 );
 a17537a <=( (not A266)  and  a17536a );
 a17538a <=( a17537a  and  a17532a );
 a17541a <=( A166  and  A168 );
 a17545a <=( (not A233)  and  (not A201) );
 a17546a <=( (not A200)  and  a17545a );
 a17547a <=( a17546a  and  a17541a );
 a17551a <=( (not A265)  and  (not A236) );
 a17552a <=( (not A235)  and  a17551a );
 a17556a <=( A299  and  A298 );
 a17557a <=( (not A266)  and  a17556a );
 a17558a <=( a17557a  and  a17552a );
 a17561a <=( A166  and  A168 );
 a17565a <=( (not A233)  and  (not A201) );
 a17566a <=( (not A200)  and  a17565a );
 a17567a <=( a17566a  and  a17561a );
 a17571a <=( (not A265)  and  (not A236) );
 a17572a <=( (not A235)  and  a17571a );
 a17576a <=( (not A299)  and  (not A298) );
 a17577a <=( (not A266)  and  a17576a );
 a17578a <=( a17577a  and  a17572a );
 a17581a <=( A166  and  A168 );
 a17585a <=( (not A233)  and  (not A201) );
 a17586a <=( (not A200)  and  a17585a );
 a17587a <=( a17586a  and  a17581a );
 a17591a <=( A266  and  A265 );
 a17592a <=( (not A234)  and  a17591a );
 a17596a <=( (not A302)  and  (not A301) );
 a17597a <=( A298  and  a17596a );
 a17598a <=( a17597a  and  a17592a );
 a17601a <=( A166  and  A168 );
 a17605a <=( (not A233)  and  (not A201) );
 a17606a <=( (not A200)  and  a17605a );
 a17607a <=( a17606a  and  a17601a );
 a17611a <=( (not A268)  and  (not A266) );
 a17612a <=( (not A234)  and  a17611a );
 a17616a <=( (not A300)  and  A298 );
 a17617a <=( (not A269)  and  a17616a );
 a17618a <=( a17617a  and  a17612a );
 a17621a <=( A166  and  A168 );
 a17625a <=( (not A233)  and  (not A201) );
 a17626a <=( (not A200)  and  a17625a );
 a17627a <=( a17626a  and  a17621a );
 a17631a <=( (not A268)  and  (not A266) );
 a17632a <=( (not A234)  and  a17631a );
 a17636a <=( A299  and  A298 );
 a17637a <=( (not A269)  and  a17636a );
 a17638a <=( a17637a  and  a17632a );
 a17641a <=( A166  and  A168 );
 a17645a <=( (not A233)  and  (not A201) );
 a17646a <=( (not A200)  and  a17645a );
 a17647a <=( a17646a  and  a17641a );
 a17651a <=( (not A268)  and  (not A266) );
 a17652a <=( (not A234)  and  a17651a );
 a17656a <=( (not A299)  and  (not A298) );
 a17657a <=( (not A269)  and  a17656a );
 a17658a <=( a17657a  and  a17652a );
 a17661a <=( A166  and  A168 );
 a17665a <=( (not A233)  and  (not A201) );
 a17666a <=( (not A200)  and  a17665a );
 a17667a <=( a17666a  and  a17661a );
 a17671a <=( (not A267)  and  (not A266) );
 a17672a <=( (not A234)  and  a17671a );
 a17676a <=( (not A302)  and  (not A301) );
 a17677a <=( A298  and  a17676a );
 a17678a <=( a17677a  and  a17672a );
 a17681a <=( A166  and  A168 );
 a17685a <=( (not A233)  and  (not A201) );
 a17686a <=( (not A200)  and  a17685a );
 a17687a <=( a17686a  and  a17681a );
 a17691a <=( (not A266)  and  (not A265) );
 a17692a <=( (not A234)  and  a17691a );
 a17696a <=( (not A302)  and  (not A301) );
 a17697a <=( A298  and  a17696a );
 a17698a <=( a17697a  and  a17692a );
 a17701a <=( A166  and  A168 );
 a17705a <=( (not A232)  and  (not A201) );
 a17706a <=( (not A200)  and  a17705a );
 a17707a <=( a17706a  and  a17701a );
 a17711a <=( A266  and  A265 );
 a17712a <=( (not A233)  and  a17711a );
 a17716a <=( (not A302)  and  (not A301) );
 a17717a <=( A298  and  a17716a );
 a17718a <=( a17717a  and  a17712a );
 a17721a <=( A166  and  A168 );
 a17725a <=( (not A232)  and  (not A201) );
 a17726a <=( (not A200)  and  a17725a );
 a17727a <=( a17726a  and  a17721a );
 a17731a <=( (not A268)  and  (not A266) );
 a17732a <=( (not A233)  and  a17731a );
 a17736a <=( (not A300)  and  A298 );
 a17737a <=( (not A269)  and  a17736a );
 a17738a <=( a17737a  and  a17732a );
 a17741a <=( A166  and  A168 );
 a17745a <=( (not A232)  and  (not A201) );
 a17746a <=( (not A200)  and  a17745a );
 a17747a <=( a17746a  and  a17741a );
 a17751a <=( (not A268)  and  (not A266) );
 a17752a <=( (not A233)  and  a17751a );
 a17756a <=( A299  and  A298 );
 a17757a <=( (not A269)  and  a17756a );
 a17758a <=( a17757a  and  a17752a );
 a17761a <=( A166  and  A168 );
 a17765a <=( (not A232)  and  (not A201) );
 a17766a <=( (not A200)  and  a17765a );
 a17767a <=( a17766a  and  a17761a );
 a17771a <=( (not A268)  and  (not A266) );
 a17772a <=( (not A233)  and  a17771a );
 a17776a <=( (not A299)  and  (not A298) );
 a17777a <=( (not A269)  and  a17776a );
 a17778a <=( a17777a  and  a17772a );
 a17781a <=( A166  and  A168 );
 a17785a <=( (not A232)  and  (not A201) );
 a17786a <=( (not A200)  and  a17785a );
 a17787a <=( a17786a  and  a17781a );
 a17791a <=( (not A267)  and  (not A266) );
 a17792a <=( (not A233)  and  a17791a );
 a17796a <=( (not A302)  and  (not A301) );
 a17797a <=( A298  and  a17796a );
 a17798a <=( a17797a  and  a17792a );
 a17801a <=( A166  and  A168 );
 a17805a <=( (not A232)  and  (not A201) );
 a17806a <=( (not A200)  and  a17805a );
 a17807a <=( a17806a  and  a17801a );
 a17811a <=( (not A266)  and  (not A265) );
 a17812a <=( (not A233)  and  a17811a );
 a17816a <=( (not A302)  and  (not A301) );
 a17817a <=( A298  and  a17816a );
 a17818a <=( a17817a  and  a17812a );
 a17821a <=( A166  and  A168 );
 a17825a <=( A232  and  (not A200) );
 a17826a <=( (not A199)  and  a17825a );
 a17827a <=( a17826a  and  a17821a );
 a17831a <=( (not A268)  and  A265 );
 a17832a <=( A233  and  a17831a );
 a17836a <=( (not A300)  and  (not A299) );
 a17837a <=( (not A269)  and  a17836a );
 a17838a <=( a17837a  and  a17832a );
 a17841a <=( A166  and  A168 );
 a17845a <=( A232  and  (not A200) );
 a17846a <=( (not A199)  and  a17845a );
 a17847a <=( a17846a  and  a17841a );
 a17851a <=( (not A268)  and  A265 );
 a17852a <=( A233  and  a17851a );
 a17856a <=( A299  and  A298 );
 a17857a <=( (not A269)  and  a17856a );
 a17858a <=( a17857a  and  a17852a );
 a17861a <=( A166  and  A168 );
 a17865a <=( A232  and  (not A200) );
 a17866a <=( (not A199)  and  a17865a );
 a17867a <=( a17866a  and  a17861a );
 a17871a <=( (not A268)  and  A265 );
 a17872a <=( A233  and  a17871a );
 a17876a <=( (not A299)  and  (not A298) );
 a17877a <=( (not A269)  and  a17876a );
 a17878a <=( a17877a  and  a17872a );
 a17881a <=( A166  and  A168 );
 a17885a <=( A232  and  (not A200) );
 a17886a <=( (not A199)  and  a17885a );
 a17887a <=( a17886a  and  a17881a );
 a17891a <=( (not A267)  and  A265 );
 a17892a <=( A233  and  a17891a );
 a17896a <=( (not A302)  and  (not A301) );
 a17897a <=( (not A299)  and  a17896a );
 a17898a <=( a17897a  and  a17892a );
 a17901a <=( A166  and  A168 );
 a17905a <=( A232  and  (not A200) );
 a17906a <=( (not A199)  and  a17905a );
 a17907a <=( a17906a  and  a17901a );
 a17911a <=( A266  and  A265 );
 a17912a <=( A233  and  a17911a );
 a17916a <=( (not A302)  and  (not A301) );
 a17917a <=( (not A299)  and  a17916a );
 a17918a <=( a17917a  and  a17912a );
 a17921a <=( A166  and  A168 );
 a17925a <=( A232  and  (not A200) );
 a17926a <=( (not A199)  and  a17925a );
 a17927a <=( a17926a  and  a17921a );
 a17931a <=( (not A266)  and  (not A265) );
 a17932a <=( A233  and  a17931a );
 a17936a <=( (not A302)  and  (not A301) );
 a17937a <=( (not A299)  and  a17936a );
 a17938a <=( a17937a  and  a17932a );
 a17941a <=( A166  and  A168 );
 a17945a <=( (not A233)  and  (not A200) );
 a17946a <=( (not A199)  and  a17945a );
 a17947a <=( a17946a  and  a17941a );
 a17951a <=( A265  and  (not A236) );
 a17952a <=( (not A235)  and  a17951a );
 a17956a <=( (not A300)  and  A298 );
 a17957a <=( A266  and  a17956a );
 a17958a <=( a17957a  and  a17952a );
 a17961a <=( A166  and  A168 );
 a17965a <=( (not A233)  and  (not A200) );
 a17966a <=( (not A199)  and  a17965a );
 a17967a <=( a17966a  and  a17961a );
 a17971a <=( A265  and  (not A236) );
 a17972a <=( (not A235)  and  a17971a );
 a17976a <=( A299  and  A298 );
 a17977a <=( A266  and  a17976a );
 a17978a <=( a17977a  and  a17972a );
 a17981a <=( A166  and  A168 );
 a17985a <=( (not A233)  and  (not A200) );
 a17986a <=( (not A199)  and  a17985a );
 a17987a <=( a17986a  and  a17981a );
 a17991a <=( A265  and  (not A236) );
 a17992a <=( (not A235)  and  a17991a );
 a17996a <=( (not A299)  and  (not A298) );
 a17997a <=( A266  and  a17996a );
 a17998a <=( a17997a  and  a17992a );
 a18001a <=( A166  and  A168 );
 a18005a <=( (not A233)  and  (not A200) );
 a18006a <=( (not A199)  and  a18005a );
 a18007a <=( a18006a  and  a18001a );
 a18011a <=( (not A266)  and  (not A236) );
 a18012a <=( (not A235)  and  a18011a );
 a18016a <=( (not A300)  and  A298 );
 a18017a <=( (not A267)  and  a18016a );
 a18018a <=( a18017a  and  a18012a );
 a18021a <=( A166  and  A168 );
 a18025a <=( (not A233)  and  (not A200) );
 a18026a <=( (not A199)  and  a18025a );
 a18027a <=( a18026a  and  a18021a );
 a18031a <=( (not A266)  and  (not A236) );
 a18032a <=( (not A235)  and  a18031a );
 a18036a <=( A299  and  A298 );
 a18037a <=( (not A267)  and  a18036a );
 a18038a <=( a18037a  and  a18032a );
 a18041a <=( A166  and  A168 );
 a18045a <=( (not A233)  and  (not A200) );
 a18046a <=( (not A199)  and  a18045a );
 a18047a <=( a18046a  and  a18041a );
 a18051a <=( (not A266)  and  (not A236) );
 a18052a <=( (not A235)  and  a18051a );
 a18056a <=( (not A299)  and  (not A298) );
 a18057a <=( (not A267)  and  a18056a );
 a18058a <=( a18057a  and  a18052a );
 a18061a <=( A166  and  A168 );
 a18065a <=( (not A233)  and  (not A200) );
 a18066a <=( (not A199)  and  a18065a );
 a18067a <=( a18066a  and  a18061a );
 a18071a <=( (not A265)  and  (not A236) );
 a18072a <=( (not A235)  and  a18071a );
 a18076a <=( (not A300)  and  A298 );
 a18077a <=( (not A266)  and  a18076a );
 a18078a <=( a18077a  and  a18072a );
 a18081a <=( A166  and  A168 );
 a18085a <=( (not A233)  and  (not A200) );
 a18086a <=( (not A199)  and  a18085a );
 a18087a <=( a18086a  and  a18081a );
 a18091a <=( (not A265)  and  (not A236) );
 a18092a <=( (not A235)  and  a18091a );
 a18096a <=( A299  and  A298 );
 a18097a <=( (not A266)  and  a18096a );
 a18098a <=( a18097a  and  a18092a );
 a18101a <=( A166  and  A168 );
 a18105a <=( (not A233)  and  (not A200) );
 a18106a <=( (not A199)  and  a18105a );
 a18107a <=( a18106a  and  a18101a );
 a18111a <=( (not A265)  and  (not A236) );
 a18112a <=( (not A235)  and  a18111a );
 a18116a <=( (not A299)  and  (not A298) );
 a18117a <=( (not A266)  and  a18116a );
 a18118a <=( a18117a  and  a18112a );
 a18121a <=( A166  and  A168 );
 a18125a <=( (not A233)  and  (not A200) );
 a18126a <=( (not A199)  and  a18125a );
 a18127a <=( a18126a  and  a18121a );
 a18131a <=( A266  and  A265 );
 a18132a <=( (not A234)  and  a18131a );
 a18136a <=( (not A302)  and  (not A301) );
 a18137a <=( A298  and  a18136a );
 a18138a <=( a18137a  and  a18132a );
 a18141a <=( A166  and  A168 );
 a18145a <=( (not A233)  and  (not A200) );
 a18146a <=( (not A199)  and  a18145a );
 a18147a <=( a18146a  and  a18141a );
 a18151a <=( (not A268)  and  (not A266) );
 a18152a <=( (not A234)  and  a18151a );
 a18156a <=( (not A300)  and  A298 );
 a18157a <=( (not A269)  and  a18156a );
 a18158a <=( a18157a  and  a18152a );
 a18161a <=( A166  and  A168 );
 a18165a <=( (not A233)  and  (not A200) );
 a18166a <=( (not A199)  and  a18165a );
 a18167a <=( a18166a  and  a18161a );
 a18171a <=( (not A268)  and  (not A266) );
 a18172a <=( (not A234)  and  a18171a );
 a18176a <=( A299  and  A298 );
 a18177a <=( (not A269)  and  a18176a );
 a18178a <=( a18177a  and  a18172a );
 a18181a <=( A166  and  A168 );
 a18185a <=( (not A233)  and  (not A200) );
 a18186a <=( (not A199)  and  a18185a );
 a18187a <=( a18186a  and  a18181a );
 a18191a <=( (not A268)  and  (not A266) );
 a18192a <=( (not A234)  and  a18191a );
 a18196a <=( (not A299)  and  (not A298) );
 a18197a <=( (not A269)  and  a18196a );
 a18198a <=( a18197a  and  a18192a );
 a18201a <=( A166  and  A168 );
 a18205a <=( (not A233)  and  (not A200) );
 a18206a <=( (not A199)  and  a18205a );
 a18207a <=( a18206a  and  a18201a );
 a18211a <=( (not A267)  and  (not A266) );
 a18212a <=( (not A234)  and  a18211a );
 a18216a <=( (not A302)  and  (not A301) );
 a18217a <=( A298  and  a18216a );
 a18218a <=( a18217a  and  a18212a );
 a18221a <=( A166  and  A168 );
 a18225a <=( (not A233)  and  (not A200) );
 a18226a <=( (not A199)  and  a18225a );
 a18227a <=( a18226a  and  a18221a );
 a18231a <=( (not A266)  and  (not A265) );
 a18232a <=( (not A234)  and  a18231a );
 a18236a <=( (not A302)  and  (not A301) );
 a18237a <=( A298  and  a18236a );
 a18238a <=( a18237a  and  a18232a );
 a18241a <=( A166  and  A168 );
 a18245a <=( (not A232)  and  (not A200) );
 a18246a <=( (not A199)  and  a18245a );
 a18247a <=( a18246a  and  a18241a );
 a18251a <=( A266  and  A265 );
 a18252a <=( (not A233)  and  a18251a );
 a18256a <=( (not A302)  and  (not A301) );
 a18257a <=( A298  and  a18256a );
 a18258a <=( a18257a  and  a18252a );
 a18261a <=( A166  and  A168 );
 a18265a <=( (not A232)  and  (not A200) );
 a18266a <=( (not A199)  and  a18265a );
 a18267a <=( a18266a  and  a18261a );
 a18271a <=( (not A268)  and  (not A266) );
 a18272a <=( (not A233)  and  a18271a );
 a18276a <=( (not A300)  and  A298 );
 a18277a <=( (not A269)  and  a18276a );
 a18278a <=( a18277a  and  a18272a );
 a18281a <=( A166  and  A168 );
 a18285a <=( (not A232)  and  (not A200) );
 a18286a <=( (not A199)  and  a18285a );
 a18287a <=( a18286a  and  a18281a );
 a18291a <=( (not A268)  and  (not A266) );
 a18292a <=( (not A233)  and  a18291a );
 a18296a <=( A299  and  A298 );
 a18297a <=( (not A269)  and  a18296a );
 a18298a <=( a18297a  and  a18292a );
 a18301a <=( A166  and  A168 );
 a18305a <=( (not A232)  and  (not A200) );
 a18306a <=( (not A199)  and  a18305a );
 a18307a <=( a18306a  and  a18301a );
 a18311a <=( (not A268)  and  (not A266) );
 a18312a <=( (not A233)  and  a18311a );
 a18316a <=( (not A299)  and  (not A298) );
 a18317a <=( (not A269)  and  a18316a );
 a18318a <=( a18317a  and  a18312a );
 a18321a <=( A166  and  A168 );
 a18325a <=( (not A232)  and  (not A200) );
 a18326a <=( (not A199)  and  a18325a );
 a18327a <=( a18326a  and  a18321a );
 a18331a <=( (not A267)  and  (not A266) );
 a18332a <=( (not A233)  and  a18331a );
 a18336a <=( (not A302)  and  (not A301) );
 a18337a <=( A298  and  a18336a );
 a18338a <=( a18337a  and  a18332a );
 a18341a <=( A166  and  A168 );
 a18345a <=( (not A232)  and  (not A200) );
 a18346a <=( (not A199)  and  a18345a );
 a18347a <=( a18346a  and  a18341a );
 a18351a <=( (not A266)  and  (not A265) );
 a18352a <=( (not A233)  and  a18351a );
 a18356a <=( (not A302)  and  (not A301) );
 a18357a <=( A298  and  a18356a );
 a18358a <=( a18357a  and  a18352a );
 a18361a <=( A167  and  A168 );
 a18365a <=( A232  and  A200 );
 a18366a <=( A199  and  a18365a );
 a18367a <=( a18366a  and  a18361a );
 a18371a <=( (not A268)  and  A265 );
 a18372a <=( A233  and  a18371a );
 a18376a <=( (not A300)  and  (not A299) );
 a18377a <=( (not A269)  and  a18376a );
 a18378a <=( a18377a  and  a18372a );
 a18381a <=( A167  and  A168 );
 a18385a <=( A232  and  A200 );
 a18386a <=( A199  and  a18385a );
 a18387a <=( a18386a  and  a18381a );
 a18391a <=( (not A268)  and  A265 );
 a18392a <=( A233  and  a18391a );
 a18396a <=( A299  and  A298 );
 a18397a <=( (not A269)  and  a18396a );
 a18398a <=( a18397a  and  a18392a );
 a18401a <=( A167  and  A168 );
 a18405a <=( A232  and  A200 );
 a18406a <=( A199  and  a18405a );
 a18407a <=( a18406a  and  a18401a );
 a18411a <=( (not A268)  and  A265 );
 a18412a <=( A233  and  a18411a );
 a18416a <=( (not A299)  and  (not A298) );
 a18417a <=( (not A269)  and  a18416a );
 a18418a <=( a18417a  and  a18412a );
 a18421a <=( A167  and  A168 );
 a18425a <=( A232  and  A200 );
 a18426a <=( A199  and  a18425a );
 a18427a <=( a18426a  and  a18421a );
 a18431a <=( (not A267)  and  A265 );
 a18432a <=( A233  and  a18431a );
 a18436a <=( (not A302)  and  (not A301) );
 a18437a <=( (not A299)  and  a18436a );
 a18438a <=( a18437a  and  a18432a );
 a18441a <=( A167  and  A168 );
 a18445a <=( A232  and  A200 );
 a18446a <=( A199  and  a18445a );
 a18447a <=( a18446a  and  a18441a );
 a18451a <=( A266  and  A265 );
 a18452a <=( A233  and  a18451a );
 a18456a <=( (not A302)  and  (not A301) );
 a18457a <=( (not A299)  and  a18456a );
 a18458a <=( a18457a  and  a18452a );
 a18461a <=( A167  and  A168 );
 a18465a <=( A232  and  A200 );
 a18466a <=( A199  and  a18465a );
 a18467a <=( a18466a  and  a18461a );
 a18471a <=( (not A266)  and  (not A265) );
 a18472a <=( A233  and  a18471a );
 a18476a <=( (not A302)  and  (not A301) );
 a18477a <=( (not A299)  and  a18476a );
 a18478a <=( a18477a  and  a18472a );
 a18481a <=( A167  and  A168 );
 a18485a <=( (not A233)  and  A200 );
 a18486a <=( A199  and  a18485a );
 a18487a <=( a18486a  and  a18481a );
 a18491a <=( A265  and  (not A236) );
 a18492a <=( (not A235)  and  a18491a );
 a18496a <=( (not A300)  and  A298 );
 a18497a <=( A266  and  a18496a );
 a18498a <=( a18497a  and  a18492a );
 a18501a <=( A167  and  A168 );
 a18505a <=( (not A233)  and  A200 );
 a18506a <=( A199  and  a18505a );
 a18507a <=( a18506a  and  a18501a );
 a18511a <=( A265  and  (not A236) );
 a18512a <=( (not A235)  and  a18511a );
 a18516a <=( A299  and  A298 );
 a18517a <=( A266  and  a18516a );
 a18518a <=( a18517a  and  a18512a );
 a18521a <=( A167  and  A168 );
 a18525a <=( (not A233)  and  A200 );
 a18526a <=( A199  and  a18525a );
 a18527a <=( a18526a  and  a18521a );
 a18531a <=( A265  and  (not A236) );
 a18532a <=( (not A235)  and  a18531a );
 a18536a <=( (not A299)  and  (not A298) );
 a18537a <=( A266  and  a18536a );
 a18538a <=( a18537a  and  a18532a );
 a18541a <=( A167  and  A168 );
 a18545a <=( (not A233)  and  A200 );
 a18546a <=( A199  and  a18545a );
 a18547a <=( a18546a  and  a18541a );
 a18551a <=( (not A266)  and  (not A236) );
 a18552a <=( (not A235)  and  a18551a );
 a18556a <=( (not A300)  and  A298 );
 a18557a <=( (not A267)  and  a18556a );
 a18558a <=( a18557a  and  a18552a );
 a18561a <=( A167  and  A168 );
 a18565a <=( (not A233)  and  A200 );
 a18566a <=( A199  and  a18565a );
 a18567a <=( a18566a  and  a18561a );
 a18571a <=( (not A266)  and  (not A236) );
 a18572a <=( (not A235)  and  a18571a );
 a18576a <=( A299  and  A298 );
 a18577a <=( (not A267)  and  a18576a );
 a18578a <=( a18577a  and  a18572a );
 a18581a <=( A167  and  A168 );
 a18585a <=( (not A233)  and  A200 );
 a18586a <=( A199  and  a18585a );
 a18587a <=( a18586a  and  a18581a );
 a18591a <=( (not A266)  and  (not A236) );
 a18592a <=( (not A235)  and  a18591a );
 a18596a <=( (not A299)  and  (not A298) );
 a18597a <=( (not A267)  and  a18596a );
 a18598a <=( a18597a  and  a18592a );
 a18601a <=( A167  and  A168 );
 a18605a <=( (not A233)  and  A200 );
 a18606a <=( A199  and  a18605a );
 a18607a <=( a18606a  and  a18601a );
 a18611a <=( (not A265)  and  (not A236) );
 a18612a <=( (not A235)  and  a18611a );
 a18616a <=( (not A300)  and  A298 );
 a18617a <=( (not A266)  and  a18616a );
 a18618a <=( a18617a  and  a18612a );
 a18621a <=( A167  and  A168 );
 a18625a <=( (not A233)  and  A200 );
 a18626a <=( A199  and  a18625a );
 a18627a <=( a18626a  and  a18621a );
 a18631a <=( (not A265)  and  (not A236) );
 a18632a <=( (not A235)  and  a18631a );
 a18636a <=( A299  and  A298 );
 a18637a <=( (not A266)  and  a18636a );
 a18638a <=( a18637a  and  a18632a );
 a18641a <=( A167  and  A168 );
 a18645a <=( (not A233)  and  A200 );
 a18646a <=( A199  and  a18645a );
 a18647a <=( a18646a  and  a18641a );
 a18651a <=( (not A265)  and  (not A236) );
 a18652a <=( (not A235)  and  a18651a );
 a18656a <=( (not A299)  and  (not A298) );
 a18657a <=( (not A266)  and  a18656a );
 a18658a <=( a18657a  and  a18652a );
 a18661a <=( A167  and  A168 );
 a18665a <=( (not A233)  and  A200 );
 a18666a <=( A199  and  a18665a );
 a18667a <=( a18666a  and  a18661a );
 a18671a <=( A266  and  A265 );
 a18672a <=( (not A234)  and  a18671a );
 a18676a <=( (not A302)  and  (not A301) );
 a18677a <=( A298  and  a18676a );
 a18678a <=( a18677a  and  a18672a );
 a18681a <=( A167  and  A168 );
 a18685a <=( (not A233)  and  A200 );
 a18686a <=( A199  and  a18685a );
 a18687a <=( a18686a  and  a18681a );
 a18691a <=( (not A268)  and  (not A266) );
 a18692a <=( (not A234)  and  a18691a );
 a18696a <=( (not A300)  and  A298 );
 a18697a <=( (not A269)  and  a18696a );
 a18698a <=( a18697a  and  a18692a );
 a18701a <=( A167  and  A168 );
 a18705a <=( (not A233)  and  A200 );
 a18706a <=( A199  and  a18705a );
 a18707a <=( a18706a  and  a18701a );
 a18711a <=( (not A268)  and  (not A266) );
 a18712a <=( (not A234)  and  a18711a );
 a18716a <=( A299  and  A298 );
 a18717a <=( (not A269)  and  a18716a );
 a18718a <=( a18717a  and  a18712a );
 a18721a <=( A167  and  A168 );
 a18725a <=( (not A233)  and  A200 );
 a18726a <=( A199  and  a18725a );
 a18727a <=( a18726a  and  a18721a );
 a18731a <=( (not A268)  and  (not A266) );
 a18732a <=( (not A234)  and  a18731a );
 a18736a <=( (not A299)  and  (not A298) );
 a18737a <=( (not A269)  and  a18736a );
 a18738a <=( a18737a  and  a18732a );
 a18741a <=( A167  and  A168 );
 a18745a <=( (not A233)  and  A200 );
 a18746a <=( A199  and  a18745a );
 a18747a <=( a18746a  and  a18741a );
 a18751a <=( (not A267)  and  (not A266) );
 a18752a <=( (not A234)  and  a18751a );
 a18756a <=( (not A302)  and  (not A301) );
 a18757a <=( A298  and  a18756a );
 a18758a <=( a18757a  and  a18752a );
 a18761a <=( A167  and  A168 );
 a18765a <=( (not A233)  and  A200 );
 a18766a <=( A199  and  a18765a );
 a18767a <=( a18766a  and  a18761a );
 a18771a <=( (not A266)  and  (not A265) );
 a18772a <=( (not A234)  and  a18771a );
 a18776a <=( (not A302)  and  (not A301) );
 a18777a <=( A298  and  a18776a );
 a18778a <=( a18777a  and  a18772a );
 a18781a <=( A167  and  A168 );
 a18785a <=( (not A232)  and  A200 );
 a18786a <=( A199  and  a18785a );
 a18787a <=( a18786a  and  a18781a );
 a18791a <=( A266  and  A265 );
 a18792a <=( (not A233)  and  a18791a );
 a18796a <=( (not A302)  and  (not A301) );
 a18797a <=( A298  and  a18796a );
 a18798a <=( a18797a  and  a18792a );
 a18801a <=( A167  and  A168 );
 a18805a <=( (not A232)  and  A200 );
 a18806a <=( A199  and  a18805a );
 a18807a <=( a18806a  and  a18801a );
 a18811a <=( (not A268)  and  (not A266) );
 a18812a <=( (not A233)  and  a18811a );
 a18816a <=( (not A300)  and  A298 );
 a18817a <=( (not A269)  and  a18816a );
 a18818a <=( a18817a  and  a18812a );
 a18821a <=( A167  and  A168 );
 a18825a <=( (not A232)  and  A200 );
 a18826a <=( A199  and  a18825a );
 a18827a <=( a18826a  and  a18821a );
 a18831a <=( (not A268)  and  (not A266) );
 a18832a <=( (not A233)  and  a18831a );
 a18836a <=( A299  and  A298 );
 a18837a <=( (not A269)  and  a18836a );
 a18838a <=( a18837a  and  a18832a );
 a18841a <=( A167  and  A168 );
 a18845a <=( (not A232)  and  A200 );
 a18846a <=( A199  and  a18845a );
 a18847a <=( a18846a  and  a18841a );
 a18851a <=( (not A268)  and  (not A266) );
 a18852a <=( (not A233)  and  a18851a );
 a18856a <=( (not A299)  and  (not A298) );
 a18857a <=( (not A269)  and  a18856a );
 a18858a <=( a18857a  and  a18852a );
 a18861a <=( A167  and  A168 );
 a18865a <=( (not A232)  and  A200 );
 a18866a <=( A199  and  a18865a );
 a18867a <=( a18866a  and  a18861a );
 a18871a <=( (not A267)  and  (not A266) );
 a18872a <=( (not A233)  and  a18871a );
 a18876a <=( (not A302)  and  (not A301) );
 a18877a <=( A298  and  a18876a );
 a18878a <=( a18877a  and  a18872a );
 a18881a <=( A167  and  A168 );
 a18885a <=( (not A232)  and  A200 );
 a18886a <=( A199  and  a18885a );
 a18887a <=( a18886a  and  a18881a );
 a18891a <=( (not A266)  and  (not A265) );
 a18892a <=( (not A233)  and  a18891a );
 a18896a <=( (not A302)  and  (not A301) );
 a18897a <=( A298  and  a18896a );
 a18898a <=( a18897a  and  a18892a );
 a18901a <=( A167  and  A168 );
 a18905a <=( (not A203)  and  (not A202) );
 a18906a <=( (not A200)  and  a18905a );
 a18907a <=( a18906a  and  a18901a );
 a18911a <=( A265  and  A233 );
 a18912a <=( A232  and  a18911a );
 a18916a <=( (not A300)  and  (not A299) );
 a18917a <=( (not A267)  and  a18916a );
 a18918a <=( a18917a  and  a18912a );
 a18921a <=( A167  and  A168 );
 a18925a <=( (not A203)  and  (not A202) );
 a18926a <=( (not A200)  and  a18925a );
 a18927a <=( a18926a  and  a18921a );
 a18931a <=( A265  and  A233 );
 a18932a <=( A232  and  a18931a );
 a18936a <=( A299  and  A298 );
 a18937a <=( (not A267)  and  a18936a );
 a18938a <=( a18937a  and  a18932a );
 a18941a <=( A167  and  A168 );
 a18945a <=( (not A203)  and  (not A202) );
 a18946a <=( (not A200)  and  a18945a );
 a18947a <=( a18946a  and  a18941a );
 a18951a <=( A265  and  A233 );
 a18952a <=( A232  and  a18951a );
 a18956a <=( (not A299)  and  (not A298) );
 a18957a <=( (not A267)  and  a18956a );
 a18958a <=( a18957a  and  a18952a );
 a18961a <=( A167  and  A168 );
 a18965a <=( (not A203)  and  (not A202) );
 a18966a <=( (not A200)  and  a18965a );
 a18967a <=( a18966a  and  a18961a );
 a18971a <=( A265  and  A233 );
 a18972a <=( A232  and  a18971a );
 a18976a <=( (not A300)  and  (not A299) );
 a18977a <=( A266  and  a18976a );
 a18978a <=( a18977a  and  a18972a );
 a18981a <=( A167  and  A168 );
 a18985a <=( (not A203)  and  (not A202) );
 a18986a <=( (not A200)  and  a18985a );
 a18987a <=( a18986a  and  a18981a );
 a18991a <=( A265  and  A233 );
 a18992a <=( A232  and  a18991a );
 a18996a <=( A299  and  A298 );
 a18997a <=( A266  and  a18996a );
 a18998a <=( a18997a  and  a18992a );
 a19001a <=( A167  and  A168 );
 a19005a <=( (not A203)  and  (not A202) );
 a19006a <=( (not A200)  and  a19005a );
 a19007a <=( a19006a  and  a19001a );
 a19011a <=( A265  and  A233 );
 a19012a <=( A232  and  a19011a );
 a19016a <=( (not A299)  and  (not A298) );
 a19017a <=( A266  and  a19016a );
 a19018a <=( a19017a  and  a19012a );
 a19021a <=( A167  and  A168 );
 a19025a <=( (not A203)  and  (not A202) );
 a19026a <=( (not A200)  and  a19025a );
 a19027a <=( a19026a  and  a19021a );
 a19031a <=( (not A265)  and  A233 );
 a19032a <=( A232  and  a19031a );
 a19036a <=( (not A300)  and  (not A299) );
 a19037a <=( (not A266)  and  a19036a );
 a19038a <=( a19037a  and  a19032a );
 a19041a <=( A167  and  A168 );
 a19045a <=( (not A203)  and  (not A202) );
 a19046a <=( (not A200)  and  a19045a );
 a19047a <=( a19046a  and  a19041a );
 a19051a <=( (not A265)  and  A233 );
 a19052a <=( A232  and  a19051a );
 a19056a <=( A299  and  A298 );
 a19057a <=( (not A266)  and  a19056a );
 a19058a <=( a19057a  and  a19052a );
 a19061a <=( A167  and  A168 );
 a19065a <=( (not A203)  and  (not A202) );
 a19066a <=( (not A200)  and  a19065a );
 a19067a <=( a19066a  and  a19061a );
 a19071a <=( (not A265)  and  A233 );
 a19072a <=( A232  and  a19071a );
 a19076a <=( (not A299)  and  (not A298) );
 a19077a <=( (not A266)  and  a19076a );
 a19078a <=( a19077a  and  a19072a );
 a19081a <=( A167  and  A168 );
 a19085a <=( (not A203)  and  (not A202) );
 a19086a <=( (not A200)  and  a19085a );
 a19087a <=( a19086a  and  a19081a );
 a19091a <=( A298  and  A233 );
 a19092a <=( (not A232)  and  a19091a );
 a19096a <=( A301  and  A300 );
 a19097a <=( (not A299)  and  a19096a );
 a19098a <=( a19097a  and  a19092a );
 a19101a <=( A167  and  A168 );
 a19105a <=( (not A203)  and  (not A202) );
 a19106a <=( (not A200)  and  a19105a );
 a19107a <=( a19106a  and  a19101a );
 a19111a <=( A298  and  A233 );
 a19112a <=( (not A232)  and  a19111a );
 a19116a <=( A302  and  A300 );
 a19117a <=( (not A299)  and  a19116a );
 a19118a <=( a19117a  and  a19112a );
 a19121a <=( A167  and  A168 );
 a19125a <=( (not A203)  and  (not A202) );
 a19126a <=( (not A200)  and  a19125a );
 a19127a <=( a19126a  and  a19121a );
 a19131a <=( A265  and  A233 );
 a19132a <=( (not A232)  and  a19131a );
 a19136a <=( A268  and  A267 );
 a19137a <=( (not A266)  and  a19136a );
 a19138a <=( a19137a  and  a19132a );
 a19141a <=( A167  and  A168 );
 a19145a <=( (not A203)  and  (not A202) );
 a19146a <=( (not A200)  and  a19145a );
 a19147a <=( a19146a  and  a19141a );
 a19151a <=( A265  and  A233 );
 a19152a <=( (not A232)  and  a19151a );
 a19156a <=( A269  and  A267 );
 a19157a <=( (not A266)  and  a19156a );
 a19158a <=( a19157a  and  a19152a );
 a19161a <=( A167  and  A168 );
 a19165a <=( (not A203)  and  (not A202) );
 a19166a <=( (not A200)  and  a19165a );
 a19167a <=( a19166a  and  a19161a );
 a19171a <=( A265  and  (not A234) );
 a19172a <=( (not A233)  and  a19171a );
 a19176a <=( (not A300)  and  A298 );
 a19177a <=( A266  and  a19176a );
 a19178a <=( a19177a  and  a19172a );
 a19181a <=( A167  and  A168 );
 a19185a <=( (not A203)  and  (not A202) );
 a19186a <=( (not A200)  and  a19185a );
 a19187a <=( a19186a  and  a19181a );
 a19191a <=( A265  and  (not A234) );
 a19192a <=( (not A233)  and  a19191a );
 a19196a <=( A299  and  A298 );
 a19197a <=( A266  and  a19196a );
 a19198a <=( a19197a  and  a19192a );
 a19201a <=( A167  and  A168 );
 a19205a <=( (not A203)  and  (not A202) );
 a19206a <=( (not A200)  and  a19205a );
 a19207a <=( a19206a  and  a19201a );
 a19211a <=( A265  and  (not A234) );
 a19212a <=( (not A233)  and  a19211a );
 a19216a <=( (not A299)  and  (not A298) );
 a19217a <=( A266  and  a19216a );
 a19218a <=( a19217a  and  a19212a );
 a19221a <=( A167  and  A168 );
 a19225a <=( (not A203)  and  (not A202) );
 a19226a <=( (not A200)  and  a19225a );
 a19227a <=( a19226a  and  a19221a );
 a19231a <=( (not A266)  and  (not A234) );
 a19232a <=( (not A233)  and  a19231a );
 a19236a <=( (not A300)  and  A298 );
 a19237a <=( (not A267)  and  a19236a );
 a19238a <=( a19237a  and  a19232a );
 a19241a <=( A167  and  A168 );
 a19245a <=( (not A203)  and  (not A202) );
 a19246a <=( (not A200)  and  a19245a );
 a19247a <=( a19246a  and  a19241a );
 a19251a <=( (not A266)  and  (not A234) );
 a19252a <=( (not A233)  and  a19251a );
 a19256a <=( A299  and  A298 );
 a19257a <=( (not A267)  and  a19256a );
 a19258a <=( a19257a  and  a19252a );
 a19261a <=( A167  and  A168 );
 a19265a <=( (not A203)  and  (not A202) );
 a19266a <=( (not A200)  and  a19265a );
 a19267a <=( a19266a  and  a19261a );
 a19271a <=( (not A266)  and  (not A234) );
 a19272a <=( (not A233)  and  a19271a );
 a19276a <=( (not A299)  and  (not A298) );
 a19277a <=( (not A267)  and  a19276a );
 a19278a <=( a19277a  and  a19272a );
 a19281a <=( A167  and  A168 );
 a19285a <=( (not A203)  and  (not A202) );
 a19286a <=( (not A200)  and  a19285a );
 a19287a <=( a19286a  and  a19281a );
 a19291a <=( (not A265)  and  (not A234) );
 a19292a <=( (not A233)  and  a19291a );
 a19296a <=( (not A300)  and  A298 );
 a19297a <=( (not A266)  and  a19296a );
 a19298a <=( a19297a  and  a19292a );
 a19301a <=( A167  and  A168 );
 a19305a <=( (not A203)  and  (not A202) );
 a19306a <=( (not A200)  and  a19305a );
 a19307a <=( a19306a  and  a19301a );
 a19311a <=( (not A265)  and  (not A234) );
 a19312a <=( (not A233)  and  a19311a );
 a19316a <=( A299  and  A298 );
 a19317a <=( (not A266)  and  a19316a );
 a19318a <=( a19317a  and  a19312a );
 a19321a <=( A167  and  A168 );
 a19325a <=( (not A203)  and  (not A202) );
 a19326a <=( (not A200)  and  a19325a );
 a19327a <=( a19326a  and  a19321a );
 a19331a <=( (not A265)  and  (not A234) );
 a19332a <=( (not A233)  and  a19331a );
 a19336a <=( (not A299)  and  (not A298) );
 a19337a <=( (not A266)  and  a19336a );
 a19338a <=( a19337a  and  a19332a );
 a19341a <=( A167  and  A168 );
 a19345a <=( (not A203)  and  (not A202) );
 a19346a <=( (not A200)  and  a19345a );
 a19347a <=( a19346a  and  a19341a );
 a19351a <=( A234  and  (not A233) );
 a19352a <=( A232  and  a19351a );
 a19356a <=( A299  and  (not A298) );
 a19357a <=( A235  and  a19356a );
 a19358a <=( a19357a  and  a19352a );
 a19361a <=( A167  and  A168 );
 a19365a <=( (not A203)  and  (not A202) );
 a19366a <=( (not A200)  and  a19365a );
 a19367a <=( a19366a  and  a19361a );
 a19371a <=( A234  and  (not A233) );
 a19372a <=( A232  and  a19371a );
 a19376a <=( A266  and  (not A265) );
 a19377a <=( A235  and  a19376a );
 a19378a <=( a19377a  and  a19372a );
 a19381a <=( A167  and  A168 );
 a19385a <=( (not A203)  and  (not A202) );
 a19386a <=( (not A200)  and  a19385a );
 a19387a <=( a19386a  and  a19381a );
 a19391a <=( A234  and  (not A233) );
 a19392a <=( A232  and  a19391a );
 a19396a <=( A299  and  (not A298) );
 a19397a <=( A236  and  a19396a );
 a19398a <=( a19397a  and  a19392a );
 a19401a <=( A167  and  A168 );
 a19405a <=( (not A203)  and  (not A202) );
 a19406a <=( (not A200)  and  a19405a );
 a19407a <=( a19406a  and  a19401a );
 a19411a <=( A234  and  (not A233) );
 a19412a <=( A232  and  a19411a );
 a19416a <=( A266  and  (not A265) );
 a19417a <=( A236  and  a19416a );
 a19418a <=( a19417a  and  a19412a );
 a19421a <=( A167  and  A168 );
 a19425a <=( (not A203)  and  (not A202) );
 a19426a <=( (not A200)  and  a19425a );
 a19427a <=( a19426a  and  a19421a );
 a19431a <=( A265  and  (not A233) );
 a19432a <=( (not A232)  and  a19431a );
 a19436a <=( (not A300)  and  A298 );
 a19437a <=( A266  and  a19436a );
 a19438a <=( a19437a  and  a19432a );
 a19441a <=( A167  and  A168 );
 a19445a <=( (not A203)  and  (not A202) );
 a19446a <=( (not A200)  and  a19445a );
 a19447a <=( a19446a  and  a19441a );
 a19451a <=( A265  and  (not A233) );
 a19452a <=( (not A232)  and  a19451a );
 a19456a <=( A299  and  A298 );
 a19457a <=( A266  and  a19456a );
 a19458a <=( a19457a  and  a19452a );
 a19461a <=( A167  and  A168 );
 a19465a <=( (not A203)  and  (not A202) );
 a19466a <=( (not A200)  and  a19465a );
 a19467a <=( a19466a  and  a19461a );
 a19471a <=( A265  and  (not A233) );
 a19472a <=( (not A232)  and  a19471a );
 a19476a <=( (not A299)  and  (not A298) );
 a19477a <=( A266  and  a19476a );
 a19478a <=( a19477a  and  a19472a );
 a19481a <=( A167  and  A168 );
 a19485a <=( (not A203)  and  (not A202) );
 a19486a <=( (not A200)  and  a19485a );
 a19487a <=( a19486a  and  a19481a );
 a19491a <=( (not A266)  and  (not A233) );
 a19492a <=( (not A232)  and  a19491a );
 a19496a <=( (not A300)  and  A298 );
 a19497a <=( (not A267)  and  a19496a );
 a19498a <=( a19497a  and  a19492a );
 a19501a <=( A167  and  A168 );
 a19505a <=( (not A203)  and  (not A202) );
 a19506a <=( (not A200)  and  a19505a );
 a19507a <=( a19506a  and  a19501a );
 a19511a <=( (not A266)  and  (not A233) );
 a19512a <=( (not A232)  and  a19511a );
 a19516a <=( A299  and  A298 );
 a19517a <=( (not A267)  and  a19516a );
 a19518a <=( a19517a  and  a19512a );
 a19521a <=( A167  and  A168 );
 a19525a <=( (not A203)  and  (not A202) );
 a19526a <=( (not A200)  and  a19525a );
 a19527a <=( a19526a  and  a19521a );
 a19531a <=( (not A266)  and  (not A233) );
 a19532a <=( (not A232)  and  a19531a );
 a19536a <=( (not A299)  and  (not A298) );
 a19537a <=( (not A267)  and  a19536a );
 a19538a <=( a19537a  and  a19532a );
 a19541a <=( A167  and  A168 );
 a19545a <=( (not A203)  and  (not A202) );
 a19546a <=( (not A200)  and  a19545a );
 a19547a <=( a19546a  and  a19541a );
 a19551a <=( (not A265)  and  (not A233) );
 a19552a <=( (not A232)  and  a19551a );
 a19556a <=( (not A300)  and  A298 );
 a19557a <=( (not A266)  and  a19556a );
 a19558a <=( a19557a  and  a19552a );
 a19561a <=( A167  and  A168 );
 a19565a <=( (not A203)  and  (not A202) );
 a19566a <=( (not A200)  and  a19565a );
 a19567a <=( a19566a  and  a19561a );
 a19571a <=( (not A265)  and  (not A233) );
 a19572a <=( (not A232)  and  a19571a );
 a19576a <=( A299  and  A298 );
 a19577a <=( (not A266)  and  a19576a );
 a19578a <=( a19577a  and  a19572a );
 a19581a <=( A167  and  A168 );
 a19585a <=( (not A203)  and  (not A202) );
 a19586a <=( (not A200)  and  a19585a );
 a19587a <=( a19586a  and  a19581a );
 a19591a <=( (not A265)  and  (not A233) );
 a19592a <=( (not A232)  and  a19591a );
 a19596a <=( (not A299)  and  (not A298) );
 a19597a <=( (not A266)  and  a19596a );
 a19598a <=( a19597a  and  a19592a );
 a19601a <=( A167  and  A168 );
 a19605a <=( A232  and  (not A201) );
 a19606a <=( (not A200)  and  a19605a );
 a19607a <=( a19606a  and  a19601a );
 a19611a <=( (not A268)  and  A265 );
 a19612a <=( A233  and  a19611a );
 a19616a <=( (not A300)  and  (not A299) );
 a19617a <=( (not A269)  and  a19616a );
 a19618a <=( a19617a  and  a19612a );
 a19621a <=( A167  and  A168 );
 a19625a <=( A232  and  (not A201) );
 a19626a <=( (not A200)  and  a19625a );
 a19627a <=( a19626a  and  a19621a );
 a19631a <=( (not A268)  and  A265 );
 a19632a <=( A233  and  a19631a );
 a19636a <=( A299  and  A298 );
 a19637a <=( (not A269)  and  a19636a );
 a19638a <=( a19637a  and  a19632a );
 a19641a <=( A167  and  A168 );
 a19645a <=( A232  and  (not A201) );
 a19646a <=( (not A200)  and  a19645a );
 a19647a <=( a19646a  and  a19641a );
 a19651a <=( (not A268)  and  A265 );
 a19652a <=( A233  and  a19651a );
 a19656a <=( (not A299)  and  (not A298) );
 a19657a <=( (not A269)  and  a19656a );
 a19658a <=( a19657a  and  a19652a );
 a19661a <=( A167  and  A168 );
 a19665a <=( A232  and  (not A201) );
 a19666a <=( (not A200)  and  a19665a );
 a19667a <=( a19666a  and  a19661a );
 a19671a <=( (not A267)  and  A265 );
 a19672a <=( A233  and  a19671a );
 a19676a <=( (not A302)  and  (not A301) );
 a19677a <=( (not A299)  and  a19676a );
 a19678a <=( a19677a  and  a19672a );
 a19681a <=( A167  and  A168 );
 a19685a <=( A232  and  (not A201) );
 a19686a <=( (not A200)  and  a19685a );
 a19687a <=( a19686a  and  a19681a );
 a19691a <=( A266  and  A265 );
 a19692a <=( A233  and  a19691a );
 a19696a <=( (not A302)  and  (not A301) );
 a19697a <=( (not A299)  and  a19696a );
 a19698a <=( a19697a  and  a19692a );
 a19701a <=( A167  and  A168 );
 a19705a <=( A232  and  (not A201) );
 a19706a <=( (not A200)  and  a19705a );
 a19707a <=( a19706a  and  a19701a );
 a19711a <=( (not A266)  and  (not A265) );
 a19712a <=( A233  and  a19711a );
 a19716a <=( (not A302)  and  (not A301) );
 a19717a <=( (not A299)  and  a19716a );
 a19718a <=( a19717a  and  a19712a );
 a19721a <=( A167  and  A168 );
 a19725a <=( (not A233)  and  (not A201) );
 a19726a <=( (not A200)  and  a19725a );
 a19727a <=( a19726a  and  a19721a );
 a19731a <=( A265  and  (not A236) );
 a19732a <=( (not A235)  and  a19731a );
 a19736a <=( (not A300)  and  A298 );
 a19737a <=( A266  and  a19736a );
 a19738a <=( a19737a  and  a19732a );
 a19741a <=( A167  and  A168 );
 a19745a <=( (not A233)  and  (not A201) );
 a19746a <=( (not A200)  and  a19745a );
 a19747a <=( a19746a  and  a19741a );
 a19751a <=( A265  and  (not A236) );
 a19752a <=( (not A235)  and  a19751a );
 a19756a <=( A299  and  A298 );
 a19757a <=( A266  and  a19756a );
 a19758a <=( a19757a  and  a19752a );
 a19761a <=( A167  and  A168 );
 a19765a <=( (not A233)  and  (not A201) );
 a19766a <=( (not A200)  and  a19765a );
 a19767a <=( a19766a  and  a19761a );
 a19771a <=( A265  and  (not A236) );
 a19772a <=( (not A235)  and  a19771a );
 a19776a <=( (not A299)  and  (not A298) );
 a19777a <=( A266  and  a19776a );
 a19778a <=( a19777a  and  a19772a );
 a19781a <=( A167  and  A168 );
 a19785a <=( (not A233)  and  (not A201) );
 a19786a <=( (not A200)  and  a19785a );
 a19787a <=( a19786a  and  a19781a );
 a19791a <=( (not A266)  and  (not A236) );
 a19792a <=( (not A235)  and  a19791a );
 a19796a <=( (not A300)  and  A298 );
 a19797a <=( (not A267)  and  a19796a );
 a19798a <=( a19797a  and  a19792a );
 a19801a <=( A167  and  A168 );
 a19805a <=( (not A233)  and  (not A201) );
 a19806a <=( (not A200)  and  a19805a );
 a19807a <=( a19806a  and  a19801a );
 a19811a <=( (not A266)  and  (not A236) );
 a19812a <=( (not A235)  and  a19811a );
 a19816a <=( A299  and  A298 );
 a19817a <=( (not A267)  and  a19816a );
 a19818a <=( a19817a  and  a19812a );
 a19821a <=( A167  and  A168 );
 a19825a <=( (not A233)  and  (not A201) );
 a19826a <=( (not A200)  and  a19825a );
 a19827a <=( a19826a  and  a19821a );
 a19831a <=( (not A266)  and  (not A236) );
 a19832a <=( (not A235)  and  a19831a );
 a19836a <=( (not A299)  and  (not A298) );
 a19837a <=( (not A267)  and  a19836a );
 a19838a <=( a19837a  and  a19832a );
 a19841a <=( A167  and  A168 );
 a19845a <=( (not A233)  and  (not A201) );
 a19846a <=( (not A200)  and  a19845a );
 a19847a <=( a19846a  and  a19841a );
 a19851a <=( (not A265)  and  (not A236) );
 a19852a <=( (not A235)  and  a19851a );
 a19856a <=( (not A300)  and  A298 );
 a19857a <=( (not A266)  and  a19856a );
 a19858a <=( a19857a  and  a19852a );
 a19861a <=( A167  and  A168 );
 a19865a <=( (not A233)  and  (not A201) );
 a19866a <=( (not A200)  and  a19865a );
 a19867a <=( a19866a  and  a19861a );
 a19871a <=( (not A265)  and  (not A236) );
 a19872a <=( (not A235)  and  a19871a );
 a19876a <=( A299  and  A298 );
 a19877a <=( (not A266)  and  a19876a );
 a19878a <=( a19877a  and  a19872a );
 a19881a <=( A167  and  A168 );
 a19885a <=( (not A233)  and  (not A201) );
 a19886a <=( (not A200)  and  a19885a );
 a19887a <=( a19886a  and  a19881a );
 a19891a <=( (not A265)  and  (not A236) );
 a19892a <=( (not A235)  and  a19891a );
 a19896a <=( (not A299)  and  (not A298) );
 a19897a <=( (not A266)  and  a19896a );
 a19898a <=( a19897a  and  a19892a );
 a19901a <=( A167  and  A168 );
 a19905a <=( (not A233)  and  (not A201) );
 a19906a <=( (not A200)  and  a19905a );
 a19907a <=( a19906a  and  a19901a );
 a19911a <=( A266  and  A265 );
 a19912a <=( (not A234)  and  a19911a );
 a19916a <=( (not A302)  and  (not A301) );
 a19917a <=( A298  and  a19916a );
 a19918a <=( a19917a  and  a19912a );
 a19921a <=( A167  and  A168 );
 a19925a <=( (not A233)  and  (not A201) );
 a19926a <=( (not A200)  and  a19925a );
 a19927a <=( a19926a  and  a19921a );
 a19931a <=( (not A268)  and  (not A266) );
 a19932a <=( (not A234)  and  a19931a );
 a19936a <=( (not A300)  and  A298 );
 a19937a <=( (not A269)  and  a19936a );
 a19938a <=( a19937a  and  a19932a );
 a19941a <=( A167  and  A168 );
 a19945a <=( (not A233)  and  (not A201) );
 a19946a <=( (not A200)  and  a19945a );
 a19947a <=( a19946a  and  a19941a );
 a19951a <=( (not A268)  and  (not A266) );
 a19952a <=( (not A234)  and  a19951a );
 a19956a <=( A299  and  A298 );
 a19957a <=( (not A269)  and  a19956a );
 a19958a <=( a19957a  and  a19952a );
 a19961a <=( A167  and  A168 );
 a19965a <=( (not A233)  and  (not A201) );
 a19966a <=( (not A200)  and  a19965a );
 a19967a <=( a19966a  and  a19961a );
 a19971a <=( (not A268)  and  (not A266) );
 a19972a <=( (not A234)  and  a19971a );
 a19976a <=( (not A299)  and  (not A298) );
 a19977a <=( (not A269)  and  a19976a );
 a19978a <=( a19977a  and  a19972a );
 a19981a <=( A167  and  A168 );
 a19985a <=( (not A233)  and  (not A201) );
 a19986a <=( (not A200)  and  a19985a );
 a19987a <=( a19986a  and  a19981a );
 a19991a <=( (not A267)  and  (not A266) );
 a19992a <=( (not A234)  and  a19991a );
 a19996a <=( (not A302)  and  (not A301) );
 a19997a <=( A298  and  a19996a );
 a19998a <=( a19997a  and  a19992a );
 a20001a <=( A167  and  A168 );
 a20005a <=( (not A233)  and  (not A201) );
 a20006a <=( (not A200)  and  a20005a );
 a20007a <=( a20006a  and  a20001a );
 a20011a <=( (not A266)  and  (not A265) );
 a20012a <=( (not A234)  and  a20011a );
 a20016a <=( (not A302)  and  (not A301) );
 a20017a <=( A298  and  a20016a );
 a20018a <=( a20017a  and  a20012a );
 a20021a <=( A167  and  A168 );
 a20025a <=( (not A232)  and  (not A201) );
 a20026a <=( (not A200)  and  a20025a );
 a20027a <=( a20026a  and  a20021a );
 a20031a <=( A266  and  A265 );
 a20032a <=( (not A233)  and  a20031a );
 a20036a <=( (not A302)  and  (not A301) );
 a20037a <=( A298  and  a20036a );
 a20038a <=( a20037a  and  a20032a );
 a20041a <=( A167  and  A168 );
 a20045a <=( (not A232)  and  (not A201) );
 a20046a <=( (not A200)  and  a20045a );
 a20047a <=( a20046a  and  a20041a );
 a20051a <=( (not A268)  and  (not A266) );
 a20052a <=( (not A233)  and  a20051a );
 a20056a <=( (not A300)  and  A298 );
 a20057a <=( (not A269)  and  a20056a );
 a20058a <=( a20057a  and  a20052a );
 a20061a <=( A167  and  A168 );
 a20065a <=( (not A232)  and  (not A201) );
 a20066a <=( (not A200)  and  a20065a );
 a20067a <=( a20066a  and  a20061a );
 a20071a <=( (not A268)  and  (not A266) );
 a20072a <=( (not A233)  and  a20071a );
 a20076a <=( A299  and  A298 );
 a20077a <=( (not A269)  and  a20076a );
 a20078a <=( a20077a  and  a20072a );
 a20081a <=( A167  and  A168 );
 a20085a <=( (not A232)  and  (not A201) );
 a20086a <=( (not A200)  and  a20085a );
 a20087a <=( a20086a  and  a20081a );
 a20091a <=( (not A268)  and  (not A266) );
 a20092a <=( (not A233)  and  a20091a );
 a20096a <=( (not A299)  and  (not A298) );
 a20097a <=( (not A269)  and  a20096a );
 a20098a <=( a20097a  and  a20092a );
 a20101a <=( A167  and  A168 );
 a20105a <=( (not A232)  and  (not A201) );
 a20106a <=( (not A200)  and  a20105a );
 a20107a <=( a20106a  and  a20101a );
 a20111a <=( (not A267)  and  (not A266) );
 a20112a <=( (not A233)  and  a20111a );
 a20116a <=( (not A302)  and  (not A301) );
 a20117a <=( A298  and  a20116a );
 a20118a <=( a20117a  and  a20112a );
 a20121a <=( A167  and  A168 );
 a20125a <=( (not A232)  and  (not A201) );
 a20126a <=( (not A200)  and  a20125a );
 a20127a <=( a20126a  and  a20121a );
 a20131a <=( (not A266)  and  (not A265) );
 a20132a <=( (not A233)  and  a20131a );
 a20136a <=( (not A302)  and  (not A301) );
 a20137a <=( A298  and  a20136a );
 a20138a <=( a20137a  and  a20132a );
 a20141a <=( A167  and  A168 );
 a20145a <=( A232  and  (not A200) );
 a20146a <=( (not A199)  and  a20145a );
 a20147a <=( a20146a  and  a20141a );
 a20151a <=( (not A268)  and  A265 );
 a20152a <=( A233  and  a20151a );
 a20156a <=( (not A300)  and  (not A299) );
 a20157a <=( (not A269)  and  a20156a );
 a20158a <=( a20157a  and  a20152a );
 a20161a <=( A167  and  A168 );
 a20165a <=( A232  and  (not A200) );
 a20166a <=( (not A199)  and  a20165a );
 a20167a <=( a20166a  and  a20161a );
 a20171a <=( (not A268)  and  A265 );
 a20172a <=( A233  and  a20171a );
 a20176a <=( A299  and  A298 );
 a20177a <=( (not A269)  and  a20176a );
 a20178a <=( a20177a  and  a20172a );
 a20181a <=( A167  and  A168 );
 a20185a <=( A232  and  (not A200) );
 a20186a <=( (not A199)  and  a20185a );
 a20187a <=( a20186a  and  a20181a );
 a20191a <=( (not A268)  and  A265 );
 a20192a <=( A233  and  a20191a );
 a20196a <=( (not A299)  and  (not A298) );
 a20197a <=( (not A269)  and  a20196a );
 a20198a <=( a20197a  and  a20192a );
 a20201a <=( A167  and  A168 );
 a20205a <=( A232  and  (not A200) );
 a20206a <=( (not A199)  and  a20205a );
 a20207a <=( a20206a  and  a20201a );
 a20211a <=( (not A267)  and  A265 );
 a20212a <=( A233  and  a20211a );
 a20216a <=( (not A302)  and  (not A301) );
 a20217a <=( (not A299)  and  a20216a );
 a20218a <=( a20217a  and  a20212a );
 a20221a <=( A167  and  A168 );
 a20225a <=( A232  and  (not A200) );
 a20226a <=( (not A199)  and  a20225a );
 a20227a <=( a20226a  and  a20221a );
 a20231a <=( A266  and  A265 );
 a20232a <=( A233  and  a20231a );
 a20236a <=( (not A302)  and  (not A301) );
 a20237a <=( (not A299)  and  a20236a );
 a20238a <=( a20237a  and  a20232a );
 a20241a <=( A167  and  A168 );
 a20245a <=( A232  and  (not A200) );
 a20246a <=( (not A199)  and  a20245a );
 a20247a <=( a20246a  and  a20241a );
 a20251a <=( (not A266)  and  (not A265) );
 a20252a <=( A233  and  a20251a );
 a20256a <=( (not A302)  and  (not A301) );
 a20257a <=( (not A299)  and  a20256a );
 a20258a <=( a20257a  and  a20252a );
 a20261a <=( A167  and  A168 );
 a20265a <=( (not A233)  and  (not A200) );
 a20266a <=( (not A199)  and  a20265a );
 a20267a <=( a20266a  and  a20261a );
 a20271a <=( A265  and  (not A236) );
 a20272a <=( (not A235)  and  a20271a );
 a20276a <=( (not A300)  and  A298 );
 a20277a <=( A266  and  a20276a );
 a20278a <=( a20277a  and  a20272a );
 a20281a <=( A167  and  A168 );
 a20285a <=( (not A233)  and  (not A200) );
 a20286a <=( (not A199)  and  a20285a );
 a20287a <=( a20286a  and  a20281a );
 a20291a <=( A265  and  (not A236) );
 a20292a <=( (not A235)  and  a20291a );
 a20296a <=( A299  and  A298 );
 a20297a <=( A266  and  a20296a );
 a20298a <=( a20297a  and  a20292a );
 a20301a <=( A167  and  A168 );
 a20305a <=( (not A233)  and  (not A200) );
 a20306a <=( (not A199)  and  a20305a );
 a20307a <=( a20306a  and  a20301a );
 a20311a <=( A265  and  (not A236) );
 a20312a <=( (not A235)  and  a20311a );
 a20316a <=( (not A299)  and  (not A298) );
 a20317a <=( A266  and  a20316a );
 a20318a <=( a20317a  and  a20312a );
 a20321a <=( A167  and  A168 );
 a20325a <=( (not A233)  and  (not A200) );
 a20326a <=( (not A199)  and  a20325a );
 a20327a <=( a20326a  and  a20321a );
 a20331a <=( (not A266)  and  (not A236) );
 a20332a <=( (not A235)  and  a20331a );
 a20336a <=( (not A300)  and  A298 );
 a20337a <=( (not A267)  and  a20336a );
 a20338a <=( a20337a  and  a20332a );
 a20341a <=( A167  and  A168 );
 a20345a <=( (not A233)  and  (not A200) );
 a20346a <=( (not A199)  and  a20345a );
 a20347a <=( a20346a  and  a20341a );
 a20351a <=( (not A266)  and  (not A236) );
 a20352a <=( (not A235)  and  a20351a );
 a20356a <=( A299  and  A298 );
 a20357a <=( (not A267)  and  a20356a );
 a20358a <=( a20357a  and  a20352a );
 a20361a <=( A167  and  A168 );
 a20365a <=( (not A233)  and  (not A200) );
 a20366a <=( (not A199)  and  a20365a );
 a20367a <=( a20366a  and  a20361a );
 a20371a <=( (not A266)  and  (not A236) );
 a20372a <=( (not A235)  and  a20371a );
 a20376a <=( (not A299)  and  (not A298) );
 a20377a <=( (not A267)  and  a20376a );
 a20378a <=( a20377a  and  a20372a );
 a20381a <=( A167  and  A168 );
 a20385a <=( (not A233)  and  (not A200) );
 a20386a <=( (not A199)  and  a20385a );
 a20387a <=( a20386a  and  a20381a );
 a20391a <=( (not A265)  and  (not A236) );
 a20392a <=( (not A235)  and  a20391a );
 a20396a <=( (not A300)  and  A298 );
 a20397a <=( (not A266)  and  a20396a );
 a20398a <=( a20397a  and  a20392a );
 a20401a <=( A167  and  A168 );
 a20405a <=( (not A233)  and  (not A200) );
 a20406a <=( (not A199)  and  a20405a );
 a20407a <=( a20406a  and  a20401a );
 a20411a <=( (not A265)  and  (not A236) );
 a20412a <=( (not A235)  and  a20411a );
 a20416a <=( A299  and  A298 );
 a20417a <=( (not A266)  and  a20416a );
 a20418a <=( a20417a  and  a20412a );
 a20421a <=( A167  and  A168 );
 a20425a <=( (not A233)  and  (not A200) );
 a20426a <=( (not A199)  and  a20425a );
 a20427a <=( a20426a  and  a20421a );
 a20431a <=( (not A265)  and  (not A236) );
 a20432a <=( (not A235)  and  a20431a );
 a20436a <=( (not A299)  and  (not A298) );
 a20437a <=( (not A266)  and  a20436a );
 a20438a <=( a20437a  and  a20432a );
 a20441a <=( A167  and  A168 );
 a20445a <=( (not A233)  and  (not A200) );
 a20446a <=( (not A199)  and  a20445a );
 a20447a <=( a20446a  and  a20441a );
 a20451a <=( A266  and  A265 );
 a20452a <=( (not A234)  and  a20451a );
 a20456a <=( (not A302)  and  (not A301) );
 a20457a <=( A298  and  a20456a );
 a20458a <=( a20457a  and  a20452a );
 a20461a <=( A167  and  A168 );
 a20465a <=( (not A233)  and  (not A200) );
 a20466a <=( (not A199)  and  a20465a );
 a20467a <=( a20466a  and  a20461a );
 a20471a <=( (not A268)  and  (not A266) );
 a20472a <=( (not A234)  and  a20471a );
 a20476a <=( (not A300)  and  A298 );
 a20477a <=( (not A269)  and  a20476a );
 a20478a <=( a20477a  and  a20472a );
 a20481a <=( A167  and  A168 );
 a20485a <=( (not A233)  and  (not A200) );
 a20486a <=( (not A199)  and  a20485a );
 a20487a <=( a20486a  and  a20481a );
 a20491a <=( (not A268)  and  (not A266) );
 a20492a <=( (not A234)  and  a20491a );
 a20496a <=( A299  and  A298 );
 a20497a <=( (not A269)  and  a20496a );
 a20498a <=( a20497a  and  a20492a );
 a20501a <=( A167  and  A168 );
 a20505a <=( (not A233)  and  (not A200) );
 a20506a <=( (not A199)  and  a20505a );
 a20507a <=( a20506a  and  a20501a );
 a20511a <=( (not A268)  and  (not A266) );
 a20512a <=( (not A234)  and  a20511a );
 a20516a <=( (not A299)  and  (not A298) );
 a20517a <=( (not A269)  and  a20516a );
 a20518a <=( a20517a  and  a20512a );
 a20521a <=( A167  and  A168 );
 a20525a <=( (not A233)  and  (not A200) );
 a20526a <=( (not A199)  and  a20525a );
 a20527a <=( a20526a  and  a20521a );
 a20531a <=( (not A267)  and  (not A266) );
 a20532a <=( (not A234)  and  a20531a );
 a20536a <=( (not A302)  and  (not A301) );
 a20537a <=( A298  and  a20536a );
 a20538a <=( a20537a  and  a20532a );
 a20541a <=( A167  and  A168 );
 a20545a <=( (not A233)  and  (not A200) );
 a20546a <=( (not A199)  and  a20545a );
 a20547a <=( a20546a  and  a20541a );
 a20551a <=( (not A266)  and  (not A265) );
 a20552a <=( (not A234)  and  a20551a );
 a20556a <=( (not A302)  and  (not A301) );
 a20557a <=( A298  and  a20556a );
 a20558a <=( a20557a  and  a20552a );
 a20561a <=( A167  and  A168 );
 a20565a <=( (not A232)  and  (not A200) );
 a20566a <=( (not A199)  and  a20565a );
 a20567a <=( a20566a  and  a20561a );
 a20571a <=( A266  and  A265 );
 a20572a <=( (not A233)  and  a20571a );
 a20576a <=( (not A302)  and  (not A301) );
 a20577a <=( A298  and  a20576a );
 a20578a <=( a20577a  and  a20572a );
 a20581a <=( A167  and  A168 );
 a20585a <=( (not A232)  and  (not A200) );
 a20586a <=( (not A199)  and  a20585a );
 a20587a <=( a20586a  and  a20581a );
 a20591a <=( (not A268)  and  (not A266) );
 a20592a <=( (not A233)  and  a20591a );
 a20596a <=( (not A300)  and  A298 );
 a20597a <=( (not A269)  and  a20596a );
 a20598a <=( a20597a  and  a20592a );
 a20601a <=( A167  and  A168 );
 a20605a <=( (not A232)  and  (not A200) );
 a20606a <=( (not A199)  and  a20605a );
 a20607a <=( a20606a  and  a20601a );
 a20611a <=( (not A268)  and  (not A266) );
 a20612a <=( (not A233)  and  a20611a );
 a20616a <=( A299  and  A298 );
 a20617a <=( (not A269)  and  a20616a );
 a20618a <=( a20617a  and  a20612a );
 a20621a <=( A167  and  A168 );
 a20625a <=( (not A232)  and  (not A200) );
 a20626a <=( (not A199)  and  a20625a );
 a20627a <=( a20626a  and  a20621a );
 a20631a <=( (not A268)  and  (not A266) );
 a20632a <=( (not A233)  and  a20631a );
 a20636a <=( (not A299)  and  (not A298) );
 a20637a <=( (not A269)  and  a20636a );
 a20638a <=( a20637a  and  a20632a );
 a20641a <=( A167  and  A168 );
 a20645a <=( (not A232)  and  (not A200) );
 a20646a <=( (not A199)  and  a20645a );
 a20647a <=( a20646a  and  a20641a );
 a20651a <=( (not A267)  and  (not A266) );
 a20652a <=( (not A233)  and  a20651a );
 a20656a <=( (not A302)  and  (not A301) );
 a20657a <=( A298  and  a20656a );
 a20658a <=( a20657a  and  a20652a );
 a20661a <=( A167  and  A168 );
 a20665a <=( (not A232)  and  (not A200) );
 a20666a <=( (not A199)  and  a20665a );
 a20667a <=( a20666a  and  a20661a );
 a20671a <=( (not A266)  and  (not A265) );
 a20672a <=( (not A233)  and  a20671a );
 a20676a <=( (not A302)  and  (not A301) );
 a20677a <=( A298  and  a20676a );
 a20678a <=( a20677a  and  a20672a );
 a20681a <=( (not A167)  and  A170 );
 a20685a <=( A200  and  (not A199) );
 a20686a <=( (not A166)  and  a20685a );
 a20687a <=( a20686a  and  a20681a );
 a20691a <=( A265  and  A233 );
 a20692a <=( A232  and  a20691a );
 a20696a <=( (not A300)  and  (not A299) );
 a20697a <=( (not A267)  and  a20696a );
 a20698a <=( a20697a  and  a20692a );
 a20701a <=( (not A167)  and  A170 );
 a20705a <=( A200  and  (not A199) );
 a20706a <=( (not A166)  and  a20705a );
 a20707a <=( a20706a  and  a20701a );
 a20711a <=( A265  and  A233 );
 a20712a <=( A232  and  a20711a );
 a20716a <=( A299  and  A298 );
 a20717a <=( (not A267)  and  a20716a );
 a20718a <=( a20717a  and  a20712a );
 a20721a <=( (not A167)  and  A170 );
 a20725a <=( A200  and  (not A199) );
 a20726a <=( (not A166)  and  a20725a );
 a20727a <=( a20726a  and  a20721a );
 a20731a <=( A265  and  A233 );
 a20732a <=( A232  and  a20731a );
 a20736a <=( (not A299)  and  (not A298) );
 a20737a <=( (not A267)  and  a20736a );
 a20738a <=( a20737a  and  a20732a );
 a20741a <=( (not A167)  and  A170 );
 a20745a <=( A200  and  (not A199) );
 a20746a <=( (not A166)  and  a20745a );
 a20747a <=( a20746a  and  a20741a );
 a20751a <=( A265  and  A233 );
 a20752a <=( A232  and  a20751a );
 a20756a <=( (not A300)  and  (not A299) );
 a20757a <=( A266  and  a20756a );
 a20758a <=( a20757a  and  a20752a );
 a20761a <=( (not A167)  and  A170 );
 a20765a <=( A200  and  (not A199) );
 a20766a <=( (not A166)  and  a20765a );
 a20767a <=( a20766a  and  a20761a );
 a20771a <=( A265  and  A233 );
 a20772a <=( A232  and  a20771a );
 a20776a <=( A299  and  A298 );
 a20777a <=( A266  and  a20776a );
 a20778a <=( a20777a  and  a20772a );
 a20781a <=( (not A167)  and  A170 );
 a20785a <=( A200  and  (not A199) );
 a20786a <=( (not A166)  and  a20785a );
 a20787a <=( a20786a  and  a20781a );
 a20791a <=( A265  and  A233 );
 a20792a <=( A232  and  a20791a );
 a20796a <=( (not A299)  and  (not A298) );
 a20797a <=( A266  and  a20796a );
 a20798a <=( a20797a  and  a20792a );
 a20801a <=( (not A167)  and  A170 );
 a20805a <=( A200  and  (not A199) );
 a20806a <=( (not A166)  and  a20805a );
 a20807a <=( a20806a  and  a20801a );
 a20811a <=( (not A265)  and  A233 );
 a20812a <=( A232  and  a20811a );
 a20816a <=( (not A300)  and  (not A299) );
 a20817a <=( (not A266)  and  a20816a );
 a20818a <=( a20817a  and  a20812a );
 a20821a <=( (not A167)  and  A170 );
 a20825a <=( A200  and  (not A199) );
 a20826a <=( (not A166)  and  a20825a );
 a20827a <=( a20826a  and  a20821a );
 a20831a <=( (not A265)  and  A233 );
 a20832a <=( A232  and  a20831a );
 a20836a <=( A299  and  A298 );
 a20837a <=( (not A266)  and  a20836a );
 a20838a <=( a20837a  and  a20832a );
 a20841a <=( (not A167)  and  A170 );
 a20845a <=( A200  and  (not A199) );
 a20846a <=( (not A166)  and  a20845a );
 a20847a <=( a20846a  and  a20841a );
 a20851a <=( (not A265)  and  A233 );
 a20852a <=( A232  and  a20851a );
 a20856a <=( (not A299)  and  (not A298) );
 a20857a <=( (not A266)  and  a20856a );
 a20858a <=( a20857a  and  a20852a );
 a20861a <=( (not A167)  and  A170 );
 a20865a <=( A200  and  (not A199) );
 a20866a <=( (not A166)  and  a20865a );
 a20867a <=( a20866a  and  a20861a );
 a20871a <=( A298  and  A233 );
 a20872a <=( (not A232)  and  a20871a );
 a20876a <=( A301  and  A300 );
 a20877a <=( (not A299)  and  a20876a );
 a20878a <=( a20877a  and  a20872a );
 a20881a <=( (not A167)  and  A170 );
 a20885a <=( A200  and  (not A199) );
 a20886a <=( (not A166)  and  a20885a );
 a20887a <=( a20886a  and  a20881a );
 a20891a <=( A298  and  A233 );
 a20892a <=( (not A232)  and  a20891a );
 a20896a <=( A302  and  A300 );
 a20897a <=( (not A299)  and  a20896a );
 a20898a <=( a20897a  and  a20892a );
 a20901a <=( (not A167)  and  A170 );
 a20905a <=( A200  and  (not A199) );
 a20906a <=( (not A166)  and  a20905a );
 a20907a <=( a20906a  and  a20901a );
 a20911a <=( A265  and  A233 );
 a20912a <=( (not A232)  and  a20911a );
 a20916a <=( A268  and  A267 );
 a20917a <=( (not A266)  and  a20916a );
 a20918a <=( a20917a  and  a20912a );
 a20921a <=( (not A167)  and  A170 );
 a20925a <=( A200  and  (not A199) );
 a20926a <=( (not A166)  and  a20925a );
 a20927a <=( a20926a  and  a20921a );
 a20931a <=( A265  and  A233 );
 a20932a <=( (not A232)  and  a20931a );
 a20936a <=( A269  and  A267 );
 a20937a <=( (not A266)  and  a20936a );
 a20938a <=( a20937a  and  a20932a );
 a20941a <=( (not A167)  and  A170 );
 a20945a <=( A200  and  (not A199) );
 a20946a <=( (not A166)  and  a20945a );
 a20947a <=( a20946a  and  a20941a );
 a20951a <=( A265  and  (not A234) );
 a20952a <=( (not A233)  and  a20951a );
 a20956a <=( (not A300)  and  A298 );
 a20957a <=( A266  and  a20956a );
 a20958a <=( a20957a  and  a20952a );
 a20961a <=( (not A167)  and  A170 );
 a20965a <=( A200  and  (not A199) );
 a20966a <=( (not A166)  and  a20965a );
 a20967a <=( a20966a  and  a20961a );
 a20971a <=( A265  and  (not A234) );
 a20972a <=( (not A233)  and  a20971a );
 a20976a <=( A299  and  A298 );
 a20977a <=( A266  and  a20976a );
 a20978a <=( a20977a  and  a20972a );
 a20981a <=( (not A167)  and  A170 );
 a20985a <=( A200  and  (not A199) );
 a20986a <=( (not A166)  and  a20985a );
 a20987a <=( a20986a  and  a20981a );
 a20991a <=( A265  and  (not A234) );
 a20992a <=( (not A233)  and  a20991a );
 a20996a <=( (not A299)  and  (not A298) );
 a20997a <=( A266  and  a20996a );
 a20998a <=( a20997a  and  a20992a );
 a21001a <=( (not A167)  and  A170 );
 a21005a <=( A200  and  (not A199) );
 a21006a <=( (not A166)  and  a21005a );
 a21007a <=( a21006a  and  a21001a );
 a21011a <=( (not A266)  and  (not A234) );
 a21012a <=( (not A233)  and  a21011a );
 a21016a <=( (not A300)  and  A298 );
 a21017a <=( (not A267)  and  a21016a );
 a21018a <=( a21017a  and  a21012a );
 a21021a <=( (not A167)  and  A170 );
 a21025a <=( A200  and  (not A199) );
 a21026a <=( (not A166)  and  a21025a );
 a21027a <=( a21026a  and  a21021a );
 a21031a <=( (not A266)  and  (not A234) );
 a21032a <=( (not A233)  and  a21031a );
 a21036a <=( A299  and  A298 );
 a21037a <=( (not A267)  and  a21036a );
 a21038a <=( a21037a  and  a21032a );
 a21041a <=( (not A167)  and  A170 );
 a21045a <=( A200  and  (not A199) );
 a21046a <=( (not A166)  and  a21045a );
 a21047a <=( a21046a  and  a21041a );
 a21051a <=( (not A266)  and  (not A234) );
 a21052a <=( (not A233)  and  a21051a );
 a21056a <=( (not A299)  and  (not A298) );
 a21057a <=( (not A267)  and  a21056a );
 a21058a <=( a21057a  and  a21052a );
 a21061a <=( (not A167)  and  A170 );
 a21065a <=( A200  and  (not A199) );
 a21066a <=( (not A166)  and  a21065a );
 a21067a <=( a21066a  and  a21061a );
 a21071a <=( (not A265)  and  (not A234) );
 a21072a <=( (not A233)  and  a21071a );
 a21076a <=( (not A300)  and  A298 );
 a21077a <=( (not A266)  and  a21076a );
 a21078a <=( a21077a  and  a21072a );
 a21081a <=( (not A167)  and  A170 );
 a21085a <=( A200  and  (not A199) );
 a21086a <=( (not A166)  and  a21085a );
 a21087a <=( a21086a  and  a21081a );
 a21091a <=( (not A265)  and  (not A234) );
 a21092a <=( (not A233)  and  a21091a );
 a21096a <=( A299  and  A298 );
 a21097a <=( (not A266)  and  a21096a );
 a21098a <=( a21097a  and  a21092a );
 a21101a <=( (not A167)  and  A170 );
 a21105a <=( A200  and  (not A199) );
 a21106a <=( (not A166)  and  a21105a );
 a21107a <=( a21106a  and  a21101a );
 a21111a <=( (not A265)  and  (not A234) );
 a21112a <=( (not A233)  and  a21111a );
 a21116a <=( (not A299)  and  (not A298) );
 a21117a <=( (not A266)  and  a21116a );
 a21118a <=( a21117a  and  a21112a );
 a21121a <=( (not A167)  and  A170 );
 a21125a <=( A200  and  (not A199) );
 a21126a <=( (not A166)  and  a21125a );
 a21127a <=( a21126a  and  a21121a );
 a21131a <=( A234  and  (not A233) );
 a21132a <=( A232  and  a21131a );
 a21136a <=( A299  and  (not A298) );
 a21137a <=( A235  and  a21136a );
 a21138a <=( a21137a  and  a21132a );
 a21141a <=( (not A167)  and  A170 );
 a21145a <=( A200  and  (not A199) );
 a21146a <=( (not A166)  and  a21145a );
 a21147a <=( a21146a  and  a21141a );
 a21151a <=( A234  and  (not A233) );
 a21152a <=( A232  and  a21151a );
 a21156a <=( A266  and  (not A265) );
 a21157a <=( A235  and  a21156a );
 a21158a <=( a21157a  and  a21152a );
 a21161a <=( (not A167)  and  A170 );
 a21165a <=( A200  and  (not A199) );
 a21166a <=( (not A166)  and  a21165a );
 a21167a <=( a21166a  and  a21161a );
 a21171a <=( A234  and  (not A233) );
 a21172a <=( A232  and  a21171a );
 a21176a <=( A299  and  (not A298) );
 a21177a <=( A236  and  a21176a );
 a21178a <=( a21177a  and  a21172a );
 a21181a <=( (not A167)  and  A170 );
 a21185a <=( A200  and  (not A199) );
 a21186a <=( (not A166)  and  a21185a );
 a21187a <=( a21186a  and  a21181a );
 a21191a <=( A234  and  (not A233) );
 a21192a <=( A232  and  a21191a );
 a21196a <=( A266  and  (not A265) );
 a21197a <=( A236  and  a21196a );
 a21198a <=( a21197a  and  a21192a );
 a21201a <=( (not A167)  and  A170 );
 a21205a <=( A200  and  (not A199) );
 a21206a <=( (not A166)  and  a21205a );
 a21207a <=( a21206a  and  a21201a );
 a21211a <=( A265  and  (not A233) );
 a21212a <=( (not A232)  and  a21211a );
 a21216a <=( (not A300)  and  A298 );
 a21217a <=( A266  and  a21216a );
 a21218a <=( a21217a  and  a21212a );
 a21221a <=( (not A167)  and  A170 );
 a21225a <=( A200  and  (not A199) );
 a21226a <=( (not A166)  and  a21225a );
 a21227a <=( a21226a  and  a21221a );
 a21231a <=( A265  and  (not A233) );
 a21232a <=( (not A232)  and  a21231a );
 a21236a <=( A299  and  A298 );
 a21237a <=( A266  and  a21236a );
 a21238a <=( a21237a  and  a21232a );
 a21241a <=( (not A167)  and  A170 );
 a21245a <=( A200  and  (not A199) );
 a21246a <=( (not A166)  and  a21245a );
 a21247a <=( a21246a  and  a21241a );
 a21251a <=( A265  and  (not A233) );
 a21252a <=( (not A232)  and  a21251a );
 a21256a <=( (not A299)  and  (not A298) );
 a21257a <=( A266  and  a21256a );
 a21258a <=( a21257a  and  a21252a );
 a21261a <=( (not A167)  and  A170 );
 a21265a <=( A200  and  (not A199) );
 a21266a <=( (not A166)  and  a21265a );
 a21267a <=( a21266a  and  a21261a );
 a21271a <=( (not A266)  and  (not A233) );
 a21272a <=( (not A232)  and  a21271a );
 a21276a <=( (not A300)  and  A298 );
 a21277a <=( (not A267)  and  a21276a );
 a21278a <=( a21277a  and  a21272a );
 a21281a <=( (not A167)  and  A170 );
 a21285a <=( A200  and  (not A199) );
 a21286a <=( (not A166)  and  a21285a );
 a21287a <=( a21286a  and  a21281a );
 a21291a <=( (not A266)  and  (not A233) );
 a21292a <=( (not A232)  and  a21291a );
 a21296a <=( A299  and  A298 );
 a21297a <=( (not A267)  and  a21296a );
 a21298a <=( a21297a  and  a21292a );
 a21301a <=( (not A167)  and  A170 );
 a21305a <=( A200  and  (not A199) );
 a21306a <=( (not A166)  and  a21305a );
 a21307a <=( a21306a  and  a21301a );
 a21311a <=( (not A266)  and  (not A233) );
 a21312a <=( (not A232)  and  a21311a );
 a21316a <=( (not A299)  and  (not A298) );
 a21317a <=( (not A267)  and  a21316a );
 a21318a <=( a21317a  and  a21312a );
 a21321a <=( (not A167)  and  A170 );
 a21325a <=( A200  and  (not A199) );
 a21326a <=( (not A166)  and  a21325a );
 a21327a <=( a21326a  and  a21321a );
 a21331a <=( (not A265)  and  (not A233) );
 a21332a <=( (not A232)  and  a21331a );
 a21336a <=( (not A300)  and  A298 );
 a21337a <=( (not A266)  and  a21336a );
 a21338a <=( a21337a  and  a21332a );
 a21341a <=( (not A167)  and  A170 );
 a21345a <=( A200  and  (not A199) );
 a21346a <=( (not A166)  and  a21345a );
 a21347a <=( a21346a  and  a21341a );
 a21351a <=( (not A265)  and  (not A233) );
 a21352a <=( (not A232)  and  a21351a );
 a21356a <=( A299  and  A298 );
 a21357a <=( (not A266)  and  a21356a );
 a21358a <=( a21357a  and  a21352a );
 a21361a <=( (not A167)  and  A170 );
 a21365a <=( A200  and  (not A199) );
 a21366a <=( (not A166)  and  a21365a );
 a21367a <=( a21366a  and  a21361a );
 a21371a <=( (not A265)  and  (not A233) );
 a21372a <=( (not A232)  and  a21371a );
 a21376a <=( (not A299)  and  (not A298) );
 a21377a <=( (not A266)  and  a21376a );
 a21378a <=( a21377a  and  a21372a );
 a21381a <=( (not A167)  and  A170 );
 a21385a <=( (not A200)  and  A199 );
 a21386a <=( (not A166)  and  a21385a );
 a21387a <=( a21386a  and  a21381a );
 a21391a <=( (not A232)  and  A202 );
 a21392a <=( A201  and  a21391a );
 a21396a <=( A299  and  (not A298) );
 a21397a <=( A233  and  a21396a );
 a21398a <=( a21397a  and  a21392a );
 a21401a <=( (not A167)  and  A170 );
 a21405a <=( (not A200)  and  A199 );
 a21406a <=( (not A166)  and  a21405a );
 a21407a <=( a21406a  and  a21401a );
 a21411a <=( (not A232)  and  A202 );
 a21412a <=( A201  and  a21411a );
 a21416a <=( A266  and  (not A265) );
 a21417a <=( A233  and  a21416a );
 a21418a <=( a21417a  and  a21412a );
 a21421a <=( (not A167)  and  A170 );
 a21425a <=( (not A200)  and  A199 );
 a21426a <=( (not A166)  and  a21425a );
 a21427a <=( a21426a  and  a21421a );
 a21431a <=( (not A232)  and  A203 );
 a21432a <=( A201  and  a21431a );
 a21436a <=( A299  and  (not A298) );
 a21437a <=( A233  and  a21436a );
 a21438a <=( a21437a  and  a21432a );
 a21441a <=( (not A167)  and  A170 );
 a21445a <=( (not A200)  and  A199 );
 a21446a <=( (not A166)  and  a21445a );
 a21447a <=( a21446a  and  a21441a );
 a21451a <=( (not A232)  and  A203 );
 a21452a <=( A201  and  a21451a );
 a21456a <=( A266  and  (not A265) );
 a21457a <=( A233  and  a21456a );
 a21458a <=( a21457a  and  a21452a );
 a21461a <=( A169  and  (not A170) );
 a21465a <=( (not A200)  and  A166 );
 a21466a <=( A167  and  a21465a );
 a21467a <=( a21466a  and  a21461a );
 a21471a <=( (not A232)  and  (not A203) );
 a21472a <=( (not A202)  and  a21471a );
 a21476a <=( A299  and  (not A298) );
 a21477a <=( A233  and  a21476a );
 a21478a <=( a21477a  and  a21472a );
 a21481a <=( A169  and  (not A170) );
 a21485a <=( (not A200)  and  A166 );
 a21486a <=( A167  and  a21485a );
 a21487a <=( a21486a  and  a21481a );
 a21491a <=( (not A232)  and  (not A203) );
 a21492a <=( (not A202)  and  a21491a );
 a21496a <=( A266  and  (not A265) );
 a21497a <=( A233  and  a21496a );
 a21498a <=( a21497a  and  a21492a );
 a21501a <=( A169  and  (not A170) );
 a21505a <=( (not A200)  and  (not A166) );
 a21506a <=( (not A167)  and  a21505a );
 a21507a <=( a21506a  and  a21501a );
 a21511a <=( (not A232)  and  (not A203) );
 a21512a <=( (not A202)  and  a21511a );
 a21516a <=( A299  and  (not A298) );
 a21517a <=( A233  and  a21516a );
 a21518a <=( a21517a  and  a21512a );
 a21521a <=( A169  and  (not A170) );
 a21525a <=( (not A200)  and  (not A166) );
 a21526a <=( (not A167)  and  a21525a );
 a21527a <=( a21526a  and  a21521a );
 a21531a <=( (not A232)  and  (not A203) );
 a21532a <=( (not A202)  and  a21531a );
 a21536a <=( A266  and  (not A265) );
 a21537a <=( A233  and  a21536a );
 a21538a <=( a21537a  and  a21532a );
 a21541a <=( (not A167)  and  (not A169) );
 a21545a <=( A200  and  (not A199) );
 a21546a <=( (not A166)  and  a21545a );
 a21547a <=( a21546a  and  a21541a );
 a21551a <=( A265  and  A233 );
 a21552a <=( A232  and  a21551a );
 a21556a <=( (not A300)  and  (not A299) );
 a21557a <=( (not A267)  and  a21556a );
 a21558a <=( a21557a  and  a21552a );
 a21561a <=( (not A167)  and  (not A169) );
 a21565a <=( A200  and  (not A199) );
 a21566a <=( (not A166)  and  a21565a );
 a21567a <=( a21566a  and  a21561a );
 a21571a <=( A265  and  A233 );
 a21572a <=( A232  and  a21571a );
 a21576a <=( A299  and  A298 );
 a21577a <=( (not A267)  and  a21576a );
 a21578a <=( a21577a  and  a21572a );
 a21581a <=( (not A167)  and  (not A169) );
 a21585a <=( A200  and  (not A199) );
 a21586a <=( (not A166)  and  a21585a );
 a21587a <=( a21586a  and  a21581a );
 a21591a <=( A265  and  A233 );
 a21592a <=( A232  and  a21591a );
 a21596a <=( (not A299)  and  (not A298) );
 a21597a <=( (not A267)  and  a21596a );
 a21598a <=( a21597a  and  a21592a );
 a21601a <=( (not A167)  and  (not A169) );
 a21605a <=( A200  and  (not A199) );
 a21606a <=( (not A166)  and  a21605a );
 a21607a <=( a21606a  and  a21601a );
 a21611a <=( A265  and  A233 );
 a21612a <=( A232  and  a21611a );
 a21616a <=( (not A300)  and  (not A299) );
 a21617a <=( A266  and  a21616a );
 a21618a <=( a21617a  and  a21612a );
 a21621a <=( (not A167)  and  (not A169) );
 a21625a <=( A200  and  (not A199) );
 a21626a <=( (not A166)  and  a21625a );
 a21627a <=( a21626a  and  a21621a );
 a21631a <=( A265  and  A233 );
 a21632a <=( A232  and  a21631a );
 a21636a <=( A299  and  A298 );
 a21637a <=( A266  and  a21636a );
 a21638a <=( a21637a  and  a21632a );
 a21641a <=( (not A167)  and  (not A169) );
 a21645a <=( A200  and  (not A199) );
 a21646a <=( (not A166)  and  a21645a );
 a21647a <=( a21646a  and  a21641a );
 a21651a <=( A265  and  A233 );
 a21652a <=( A232  and  a21651a );
 a21656a <=( (not A299)  and  (not A298) );
 a21657a <=( A266  and  a21656a );
 a21658a <=( a21657a  and  a21652a );
 a21661a <=( (not A167)  and  (not A169) );
 a21665a <=( A200  and  (not A199) );
 a21666a <=( (not A166)  and  a21665a );
 a21667a <=( a21666a  and  a21661a );
 a21671a <=( (not A265)  and  A233 );
 a21672a <=( A232  and  a21671a );
 a21676a <=( (not A300)  and  (not A299) );
 a21677a <=( (not A266)  and  a21676a );
 a21678a <=( a21677a  and  a21672a );
 a21681a <=( (not A167)  and  (not A169) );
 a21685a <=( A200  and  (not A199) );
 a21686a <=( (not A166)  and  a21685a );
 a21687a <=( a21686a  and  a21681a );
 a21691a <=( (not A265)  and  A233 );
 a21692a <=( A232  and  a21691a );
 a21696a <=( A299  and  A298 );
 a21697a <=( (not A266)  and  a21696a );
 a21698a <=( a21697a  and  a21692a );
 a21701a <=( (not A167)  and  (not A169) );
 a21705a <=( A200  and  (not A199) );
 a21706a <=( (not A166)  and  a21705a );
 a21707a <=( a21706a  and  a21701a );
 a21711a <=( (not A265)  and  A233 );
 a21712a <=( A232  and  a21711a );
 a21716a <=( (not A299)  and  (not A298) );
 a21717a <=( (not A266)  and  a21716a );
 a21718a <=( a21717a  and  a21712a );
 a21721a <=( (not A167)  and  (not A169) );
 a21725a <=( A200  and  (not A199) );
 a21726a <=( (not A166)  and  a21725a );
 a21727a <=( a21726a  and  a21721a );
 a21731a <=( A298  and  A233 );
 a21732a <=( (not A232)  and  a21731a );
 a21736a <=( A301  and  A300 );
 a21737a <=( (not A299)  and  a21736a );
 a21738a <=( a21737a  and  a21732a );
 a21741a <=( (not A167)  and  (not A169) );
 a21745a <=( A200  and  (not A199) );
 a21746a <=( (not A166)  and  a21745a );
 a21747a <=( a21746a  and  a21741a );
 a21751a <=( A298  and  A233 );
 a21752a <=( (not A232)  and  a21751a );
 a21756a <=( A302  and  A300 );
 a21757a <=( (not A299)  and  a21756a );
 a21758a <=( a21757a  and  a21752a );
 a21761a <=( (not A167)  and  (not A169) );
 a21765a <=( A200  and  (not A199) );
 a21766a <=( (not A166)  and  a21765a );
 a21767a <=( a21766a  and  a21761a );
 a21771a <=( A265  and  A233 );
 a21772a <=( (not A232)  and  a21771a );
 a21776a <=( A268  and  A267 );
 a21777a <=( (not A266)  and  a21776a );
 a21778a <=( a21777a  and  a21772a );
 a21781a <=( (not A167)  and  (not A169) );
 a21785a <=( A200  and  (not A199) );
 a21786a <=( (not A166)  and  a21785a );
 a21787a <=( a21786a  and  a21781a );
 a21791a <=( A265  and  A233 );
 a21792a <=( (not A232)  and  a21791a );
 a21796a <=( A269  and  A267 );
 a21797a <=( (not A266)  and  a21796a );
 a21798a <=( a21797a  and  a21792a );
 a21801a <=( (not A167)  and  (not A169) );
 a21805a <=( A200  and  (not A199) );
 a21806a <=( (not A166)  and  a21805a );
 a21807a <=( a21806a  and  a21801a );
 a21811a <=( A265  and  (not A234) );
 a21812a <=( (not A233)  and  a21811a );
 a21816a <=( (not A300)  and  A298 );
 a21817a <=( A266  and  a21816a );
 a21818a <=( a21817a  and  a21812a );
 a21821a <=( (not A167)  and  (not A169) );
 a21825a <=( A200  and  (not A199) );
 a21826a <=( (not A166)  and  a21825a );
 a21827a <=( a21826a  and  a21821a );
 a21831a <=( A265  and  (not A234) );
 a21832a <=( (not A233)  and  a21831a );
 a21836a <=( A299  and  A298 );
 a21837a <=( A266  and  a21836a );
 a21838a <=( a21837a  and  a21832a );
 a21841a <=( (not A167)  and  (not A169) );
 a21845a <=( A200  and  (not A199) );
 a21846a <=( (not A166)  and  a21845a );
 a21847a <=( a21846a  and  a21841a );
 a21851a <=( A265  and  (not A234) );
 a21852a <=( (not A233)  and  a21851a );
 a21856a <=( (not A299)  and  (not A298) );
 a21857a <=( A266  and  a21856a );
 a21858a <=( a21857a  and  a21852a );
 a21861a <=( (not A167)  and  (not A169) );
 a21865a <=( A200  and  (not A199) );
 a21866a <=( (not A166)  and  a21865a );
 a21867a <=( a21866a  and  a21861a );
 a21871a <=( (not A266)  and  (not A234) );
 a21872a <=( (not A233)  and  a21871a );
 a21876a <=( (not A300)  and  A298 );
 a21877a <=( (not A267)  and  a21876a );
 a21878a <=( a21877a  and  a21872a );
 a21881a <=( (not A167)  and  (not A169) );
 a21885a <=( A200  and  (not A199) );
 a21886a <=( (not A166)  and  a21885a );
 a21887a <=( a21886a  and  a21881a );
 a21891a <=( (not A266)  and  (not A234) );
 a21892a <=( (not A233)  and  a21891a );
 a21896a <=( A299  and  A298 );
 a21897a <=( (not A267)  and  a21896a );
 a21898a <=( a21897a  and  a21892a );
 a21901a <=( (not A167)  and  (not A169) );
 a21905a <=( A200  and  (not A199) );
 a21906a <=( (not A166)  and  a21905a );
 a21907a <=( a21906a  and  a21901a );
 a21911a <=( (not A266)  and  (not A234) );
 a21912a <=( (not A233)  and  a21911a );
 a21916a <=( (not A299)  and  (not A298) );
 a21917a <=( (not A267)  and  a21916a );
 a21918a <=( a21917a  and  a21912a );
 a21921a <=( (not A167)  and  (not A169) );
 a21925a <=( A200  and  (not A199) );
 a21926a <=( (not A166)  and  a21925a );
 a21927a <=( a21926a  and  a21921a );
 a21931a <=( (not A265)  and  (not A234) );
 a21932a <=( (not A233)  and  a21931a );
 a21936a <=( (not A300)  and  A298 );
 a21937a <=( (not A266)  and  a21936a );
 a21938a <=( a21937a  and  a21932a );
 a21941a <=( (not A167)  and  (not A169) );
 a21945a <=( A200  and  (not A199) );
 a21946a <=( (not A166)  and  a21945a );
 a21947a <=( a21946a  and  a21941a );
 a21951a <=( (not A265)  and  (not A234) );
 a21952a <=( (not A233)  and  a21951a );
 a21956a <=( A299  and  A298 );
 a21957a <=( (not A266)  and  a21956a );
 a21958a <=( a21957a  and  a21952a );
 a21961a <=( (not A167)  and  (not A169) );
 a21965a <=( A200  and  (not A199) );
 a21966a <=( (not A166)  and  a21965a );
 a21967a <=( a21966a  and  a21961a );
 a21971a <=( (not A265)  and  (not A234) );
 a21972a <=( (not A233)  and  a21971a );
 a21976a <=( (not A299)  and  (not A298) );
 a21977a <=( (not A266)  and  a21976a );
 a21978a <=( a21977a  and  a21972a );
 a21981a <=( (not A167)  and  (not A169) );
 a21985a <=( A200  and  (not A199) );
 a21986a <=( (not A166)  and  a21985a );
 a21987a <=( a21986a  and  a21981a );
 a21991a <=( A234  and  (not A233) );
 a21992a <=( A232  and  a21991a );
 a21996a <=( A299  and  (not A298) );
 a21997a <=( A235  and  a21996a );
 a21998a <=( a21997a  and  a21992a );
 a22001a <=( (not A167)  and  (not A169) );
 a22005a <=( A200  and  (not A199) );
 a22006a <=( (not A166)  and  a22005a );
 a22007a <=( a22006a  and  a22001a );
 a22011a <=( A234  and  (not A233) );
 a22012a <=( A232  and  a22011a );
 a22016a <=( A266  and  (not A265) );
 a22017a <=( A235  and  a22016a );
 a22018a <=( a22017a  and  a22012a );
 a22021a <=( (not A167)  and  (not A169) );
 a22025a <=( A200  and  (not A199) );
 a22026a <=( (not A166)  and  a22025a );
 a22027a <=( a22026a  and  a22021a );
 a22031a <=( A234  and  (not A233) );
 a22032a <=( A232  and  a22031a );
 a22036a <=( A299  and  (not A298) );
 a22037a <=( A236  and  a22036a );
 a22038a <=( a22037a  and  a22032a );
 a22041a <=( (not A167)  and  (not A169) );
 a22045a <=( A200  and  (not A199) );
 a22046a <=( (not A166)  and  a22045a );
 a22047a <=( a22046a  and  a22041a );
 a22051a <=( A234  and  (not A233) );
 a22052a <=( A232  and  a22051a );
 a22056a <=( A266  and  (not A265) );
 a22057a <=( A236  and  a22056a );
 a22058a <=( a22057a  and  a22052a );
 a22061a <=( (not A167)  and  (not A169) );
 a22065a <=( A200  and  (not A199) );
 a22066a <=( (not A166)  and  a22065a );
 a22067a <=( a22066a  and  a22061a );
 a22071a <=( A265  and  (not A233) );
 a22072a <=( (not A232)  and  a22071a );
 a22076a <=( (not A300)  and  A298 );
 a22077a <=( A266  and  a22076a );
 a22078a <=( a22077a  and  a22072a );
 a22081a <=( (not A167)  and  (not A169) );
 a22085a <=( A200  and  (not A199) );
 a22086a <=( (not A166)  and  a22085a );
 a22087a <=( a22086a  and  a22081a );
 a22091a <=( A265  and  (not A233) );
 a22092a <=( (not A232)  and  a22091a );
 a22096a <=( A299  and  A298 );
 a22097a <=( A266  and  a22096a );
 a22098a <=( a22097a  and  a22092a );
 a22101a <=( (not A167)  and  (not A169) );
 a22105a <=( A200  and  (not A199) );
 a22106a <=( (not A166)  and  a22105a );
 a22107a <=( a22106a  and  a22101a );
 a22111a <=( A265  and  (not A233) );
 a22112a <=( (not A232)  and  a22111a );
 a22116a <=( (not A299)  and  (not A298) );
 a22117a <=( A266  and  a22116a );
 a22118a <=( a22117a  and  a22112a );
 a22121a <=( (not A167)  and  (not A169) );
 a22125a <=( A200  and  (not A199) );
 a22126a <=( (not A166)  and  a22125a );
 a22127a <=( a22126a  and  a22121a );
 a22131a <=( (not A266)  and  (not A233) );
 a22132a <=( (not A232)  and  a22131a );
 a22136a <=( (not A300)  and  A298 );
 a22137a <=( (not A267)  and  a22136a );
 a22138a <=( a22137a  and  a22132a );
 a22141a <=( (not A167)  and  (not A169) );
 a22145a <=( A200  and  (not A199) );
 a22146a <=( (not A166)  and  a22145a );
 a22147a <=( a22146a  and  a22141a );
 a22151a <=( (not A266)  and  (not A233) );
 a22152a <=( (not A232)  and  a22151a );
 a22156a <=( A299  and  A298 );
 a22157a <=( (not A267)  and  a22156a );
 a22158a <=( a22157a  and  a22152a );
 a22161a <=( (not A167)  and  (not A169) );
 a22165a <=( A200  and  (not A199) );
 a22166a <=( (not A166)  and  a22165a );
 a22167a <=( a22166a  and  a22161a );
 a22171a <=( (not A266)  and  (not A233) );
 a22172a <=( (not A232)  and  a22171a );
 a22176a <=( (not A299)  and  (not A298) );
 a22177a <=( (not A267)  and  a22176a );
 a22178a <=( a22177a  and  a22172a );
 a22181a <=( (not A167)  and  (not A169) );
 a22185a <=( A200  and  (not A199) );
 a22186a <=( (not A166)  and  a22185a );
 a22187a <=( a22186a  and  a22181a );
 a22191a <=( (not A265)  and  (not A233) );
 a22192a <=( (not A232)  and  a22191a );
 a22196a <=( (not A300)  and  A298 );
 a22197a <=( (not A266)  and  a22196a );
 a22198a <=( a22197a  and  a22192a );
 a22201a <=( (not A167)  and  (not A169) );
 a22205a <=( A200  and  (not A199) );
 a22206a <=( (not A166)  and  a22205a );
 a22207a <=( a22206a  and  a22201a );
 a22211a <=( (not A265)  and  (not A233) );
 a22212a <=( (not A232)  and  a22211a );
 a22216a <=( A299  and  A298 );
 a22217a <=( (not A266)  and  a22216a );
 a22218a <=( a22217a  and  a22212a );
 a22221a <=( (not A167)  and  (not A169) );
 a22225a <=( A200  and  (not A199) );
 a22226a <=( (not A166)  and  a22225a );
 a22227a <=( a22226a  and  a22221a );
 a22231a <=( (not A265)  and  (not A233) );
 a22232a <=( (not A232)  and  a22231a );
 a22236a <=( (not A299)  and  (not A298) );
 a22237a <=( (not A266)  and  a22236a );
 a22238a <=( a22237a  and  a22232a );
 a22241a <=( (not A167)  and  (not A169) );
 a22245a <=( (not A200)  and  A199 );
 a22246a <=( (not A166)  and  a22245a );
 a22247a <=( a22246a  and  a22241a );
 a22251a <=( (not A232)  and  A202 );
 a22252a <=( A201  and  a22251a );
 a22256a <=( A299  and  (not A298) );
 a22257a <=( A233  and  a22256a );
 a22258a <=( a22257a  and  a22252a );
 a22261a <=( (not A167)  and  (not A169) );
 a22265a <=( (not A200)  and  A199 );
 a22266a <=( (not A166)  and  a22265a );
 a22267a <=( a22266a  and  a22261a );
 a22271a <=( (not A232)  and  A202 );
 a22272a <=( A201  and  a22271a );
 a22276a <=( A266  and  (not A265) );
 a22277a <=( A233  and  a22276a );
 a22278a <=( a22277a  and  a22272a );
 a22281a <=( (not A167)  and  (not A169) );
 a22285a <=( (not A200)  and  A199 );
 a22286a <=( (not A166)  and  a22285a );
 a22287a <=( a22286a  and  a22281a );
 a22291a <=( (not A232)  and  A203 );
 a22292a <=( A201  and  a22291a );
 a22296a <=( A299  and  (not A298) );
 a22297a <=( A233  and  a22296a );
 a22298a <=( a22297a  and  a22292a );
 a22301a <=( (not A167)  and  (not A169) );
 a22305a <=( (not A200)  and  A199 );
 a22306a <=( (not A166)  and  a22305a );
 a22307a <=( a22306a  and  a22301a );
 a22311a <=( (not A232)  and  A203 );
 a22312a <=( A201  and  a22311a );
 a22316a <=( A266  and  (not A265) );
 a22317a <=( A233  and  a22316a );
 a22318a <=( a22317a  and  a22312a );
 a22321a <=( (not A169)  and  A170 );
 a22325a <=( (not A200)  and  (not A166) );
 a22326a <=( A167  and  a22325a );
 a22327a <=( a22326a  and  a22321a );
 a22331a <=( (not A232)  and  (not A203) );
 a22332a <=( (not A202)  and  a22331a );
 a22336a <=( A299  and  (not A298) );
 a22337a <=( A233  and  a22336a );
 a22338a <=( a22337a  and  a22332a );
 a22341a <=( (not A169)  and  A170 );
 a22345a <=( (not A200)  and  (not A166) );
 a22346a <=( A167  and  a22345a );
 a22347a <=( a22346a  and  a22341a );
 a22351a <=( (not A232)  and  (not A203) );
 a22352a <=( (not A202)  and  a22351a );
 a22356a <=( A266  and  (not A265) );
 a22357a <=( A233  and  a22356a );
 a22358a <=( a22357a  and  a22352a );
 a22361a <=( (not A169)  and  A170 );
 a22365a <=( (not A200)  and  A166 );
 a22366a <=( (not A167)  and  a22365a );
 a22367a <=( a22366a  and  a22361a );
 a22371a <=( (not A232)  and  (not A203) );
 a22372a <=( (not A202)  and  a22371a );
 a22376a <=( A299  and  (not A298) );
 a22377a <=( A233  and  a22376a );
 a22378a <=( a22377a  and  a22372a );
 a22381a <=( (not A169)  and  A170 );
 a22385a <=( (not A200)  and  A166 );
 a22386a <=( (not A167)  and  a22385a );
 a22387a <=( a22386a  and  a22381a );
 a22391a <=( (not A232)  and  (not A203) );
 a22392a <=( (not A202)  and  a22391a );
 a22396a <=( A266  and  (not A265) );
 a22397a <=( A233  and  a22396a );
 a22398a <=( a22397a  and  a22392a );
 a22401a <=( (not A169)  and  (not A170) );
 a22405a <=( (not A200)  and  A199 );
 a22406a <=( (not A168)  and  a22405a );
 a22407a <=( a22406a  and  a22401a );
 a22411a <=( (not A232)  and  A202 );
 a22412a <=( A201  and  a22411a );
 a22416a <=( A299  and  (not A298) );
 a22417a <=( A233  and  a22416a );
 a22418a <=( a22417a  and  a22412a );
 a22421a <=( (not A169)  and  (not A170) );
 a22425a <=( (not A200)  and  A199 );
 a22426a <=( (not A168)  and  a22425a );
 a22427a <=( a22426a  and  a22421a );
 a22431a <=( (not A232)  and  A202 );
 a22432a <=( A201  and  a22431a );
 a22436a <=( A266  and  (not A265) );
 a22437a <=( A233  and  a22436a );
 a22438a <=( a22437a  and  a22432a );
 a22441a <=( (not A169)  and  (not A170) );
 a22445a <=( (not A200)  and  A199 );
 a22446a <=( (not A168)  and  a22445a );
 a22447a <=( a22446a  and  a22441a );
 a22451a <=( (not A232)  and  A203 );
 a22452a <=( A201  and  a22451a );
 a22456a <=( A299  and  (not A298) );
 a22457a <=( A233  and  a22456a );
 a22458a <=( a22457a  and  a22452a );
 a22461a <=( (not A169)  and  (not A170) );
 a22465a <=( (not A200)  and  A199 );
 a22466a <=( (not A168)  and  a22465a );
 a22467a <=( a22466a  and  a22461a );
 a22471a <=( (not A232)  and  A203 );
 a22472a <=( A201  and  a22471a );
 a22476a <=( A266  and  (not A265) );
 a22477a <=( A233  and  a22476a );
 a22478a <=( a22477a  and  a22472a );
 a22482a <=( A199  and  A166 );
 a22483a <=( A168  and  a22482a );
 a22487a <=( A233  and  A232 );
 a22488a <=( A200  and  a22487a );
 a22489a <=( a22488a  and  a22483a );
 a22493a <=( (not A269)  and  (not A268) );
 a22494a <=( A265  and  a22493a );
 a22498a <=( (not A302)  and  (not A301) );
 a22499a <=( (not A299)  and  a22498a );
 a22500a <=( a22499a  and  a22494a );
 a22504a <=( A199  and  A166 );
 a22505a <=( A168  and  a22504a );
 a22509a <=( (not A235)  and  (not A233) );
 a22510a <=( A200  and  a22509a );
 a22511a <=( a22510a  and  a22505a );
 a22515a <=( A266  and  A265 );
 a22516a <=( (not A236)  and  a22515a );
 a22520a <=( (not A302)  and  (not A301) );
 a22521a <=( A298  and  a22520a );
 a22522a <=( a22521a  and  a22516a );
 a22526a <=( A199  and  A166 );
 a22527a <=( A168  and  a22526a );
 a22531a <=( (not A235)  and  (not A233) );
 a22532a <=( A200  and  a22531a );
 a22533a <=( a22532a  and  a22527a );
 a22537a <=( (not A268)  and  (not A266) );
 a22538a <=( (not A236)  and  a22537a );
 a22542a <=( (not A300)  and  A298 );
 a22543a <=( (not A269)  and  a22542a );
 a22544a <=( a22543a  and  a22538a );
 a22548a <=( A199  and  A166 );
 a22549a <=( A168  and  a22548a );
 a22553a <=( (not A235)  and  (not A233) );
 a22554a <=( A200  and  a22553a );
 a22555a <=( a22554a  and  a22549a );
 a22559a <=( (not A268)  and  (not A266) );
 a22560a <=( (not A236)  and  a22559a );
 a22564a <=( A299  and  A298 );
 a22565a <=( (not A269)  and  a22564a );
 a22566a <=( a22565a  and  a22560a );
 a22570a <=( A199  and  A166 );
 a22571a <=( A168  and  a22570a );
 a22575a <=( (not A235)  and  (not A233) );
 a22576a <=( A200  and  a22575a );
 a22577a <=( a22576a  and  a22571a );
 a22581a <=( (not A268)  and  (not A266) );
 a22582a <=( (not A236)  and  a22581a );
 a22586a <=( (not A299)  and  (not A298) );
 a22587a <=( (not A269)  and  a22586a );
 a22588a <=( a22587a  and  a22582a );
 a22592a <=( A199  and  A166 );
 a22593a <=( A168  and  a22592a );
 a22597a <=( (not A235)  and  (not A233) );
 a22598a <=( A200  and  a22597a );
 a22599a <=( a22598a  and  a22593a );
 a22603a <=( (not A267)  and  (not A266) );
 a22604a <=( (not A236)  and  a22603a );
 a22608a <=( (not A302)  and  (not A301) );
 a22609a <=( A298  and  a22608a );
 a22610a <=( a22609a  and  a22604a );
 a22614a <=( A199  and  A166 );
 a22615a <=( A168  and  a22614a );
 a22619a <=( (not A235)  and  (not A233) );
 a22620a <=( A200  and  a22619a );
 a22621a <=( a22620a  and  a22615a );
 a22625a <=( (not A266)  and  (not A265) );
 a22626a <=( (not A236)  and  a22625a );
 a22630a <=( (not A302)  and  (not A301) );
 a22631a <=( A298  and  a22630a );
 a22632a <=( a22631a  and  a22626a );
 a22636a <=( A199  and  A166 );
 a22637a <=( A168  and  a22636a );
 a22641a <=( (not A234)  and  (not A233) );
 a22642a <=( A200  and  a22641a );
 a22643a <=( a22642a  and  a22637a );
 a22647a <=( (not A269)  and  (not A268) );
 a22648a <=( (not A266)  and  a22647a );
 a22652a <=( (not A302)  and  (not A301) );
 a22653a <=( A298  and  a22652a );
 a22654a <=( a22653a  and  a22648a );
 a22658a <=( A199  and  A166 );
 a22659a <=( A168  and  a22658a );
 a22663a <=( (not A233)  and  A232 );
 a22664a <=( A200  and  a22663a );
 a22665a <=( a22664a  and  a22659a );
 a22669a <=( A298  and  A235 );
 a22670a <=( A234  and  a22669a );
 a22674a <=( A301  and  A300 );
 a22675a <=( (not A299)  and  a22674a );
 a22676a <=( a22675a  and  a22670a );
 a22680a <=( A199  and  A166 );
 a22681a <=( A168  and  a22680a );
 a22685a <=( (not A233)  and  A232 );
 a22686a <=( A200  and  a22685a );
 a22687a <=( a22686a  and  a22681a );
 a22691a <=( A298  and  A235 );
 a22692a <=( A234  and  a22691a );
 a22696a <=( A302  and  A300 );
 a22697a <=( (not A299)  and  a22696a );
 a22698a <=( a22697a  and  a22692a );
 a22702a <=( A199  and  A166 );
 a22703a <=( A168  and  a22702a );
 a22707a <=( (not A233)  and  A232 );
 a22708a <=( A200  and  a22707a );
 a22709a <=( a22708a  and  a22703a );
 a22713a <=( A265  and  A235 );
 a22714a <=( A234  and  a22713a );
 a22718a <=( A268  and  A267 );
 a22719a <=( (not A266)  and  a22718a );
 a22720a <=( a22719a  and  a22714a );
 a22724a <=( A199  and  A166 );
 a22725a <=( A168  and  a22724a );
 a22729a <=( (not A233)  and  A232 );
 a22730a <=( A200  and  a22729a );
 a22731a <=( a22730a  and  a22725a );
 a22735a <=( A265  and  A235 );
 a22736a <=( A234  and  a22735a );
 a22740a <=( A269  and  A267 );
 a22741a <=( (not A266)  and  a22740a );
 a22742a <=( a22741a  and  a22736a );
 a22746a <=( A199  and  A166 );
 a22747a <=( A168  and  a22746a );
 a22751a <=( (not A233)  and  A232 );
 a22752a <=( A200  and  a22751a );
 a22753a <=( a22752a  and  a22747a );
 a22757a <=( A298  and  A236 );
 a22758a <=( A234  and  a22757a );
 a22762a <=( A301  and  A300 );
 a22763a <=( (not A299)  and  a22762a );
 a22764a <=( a22763a  and  a22758a );
 a22768a <=( A199  and  A166 );
 a22769a <=( A168  and  a22768a );
 a22773a <=( (not A233)  and  A232 );
 a22774a <=( A200  and  a22773a );
 a22775a <=( a22774a  and  a22769a );
 a22779a <=( A298  and  A236 );
 a22780a <=( A234  and  a22779a );
 a22784a <=( A302  and  A300 );
 a22785a <=( (not A299)  and  a22784a );
 a22786a <=( a22785a  and  a22780a );
 a22790a <=( A199  and  A166 );
 a22791a <=( A168  and  a22790a );
 a22795a <=( (not A233)  and  A232 );
 a22796a <=( A200  and  a22795a );
 a22797a <=( a22796a  and  a22791a );
 a22801a <=( A265  and  A236 );
 a22802a <=( A234  and  a22801a );
 a22806a <=( A268  and  A267 );
 a22807a <=( (not A266)  and  a22806a );
 a22808a <=( a22807a  and  a22802a );
 a22812a <=( A199  and  A166 );
 a22813a <=( A168  and  a22812a );
 a22817a <=( (not A233)  and  A232 );
 a22818a <=( A200  and  a22817a );
 a22819a <=( a22818a  and  a22813a );
 a22823a <=( A265  and  A236 );
 a22824a <=( A234  and  a22823a );
 a22828a <=( A269  and  A267 );
 a22829a <=( (not A266)  and  a22828a );
 a22830a <=( a22829a  and  a22824a );
 a22834a <=( A199  and  A166 );
 a22835a <=( A168  and  a22834a );
 a22839a <=( (not A233)  and  (not A232) );
 a22840a <=( A200  and  a22839a );
 a22841a <=( a22840a  and  a22835a );
 a22845a <=( (not A269)  and  (not A268) );
 a22846a <=( (not A266)  and  a22845a );
 a22850a <=( (not A302)  and  (not A301) );
 a22851a <=( A298  and  a22850a );
 a22852a <=( a22851a  and  a22846a );
 a22856a <=( (not A200)  and  A166 );
 a22857a <=( A168  and  a22856a );
 a22861a <=( A232  and  (not A203) );
 a22862a <=( (not A202)  and  a22861a );
 a22863a <=( a22862a  and  a22857a );
 a22867a <=( (not A268)  and  A265 );
 a22868a <=( A233  and  a22867a );
 a22872a <=( (not A300)  and  (not A299) );
 a22873a <=( (not A269)  and  a22872a );
 a22874a <=( a22873a  and  a22868a );
 a22878a <=( (not A200)  and  A166 );
 a22879a <=( A168  and  a22878a );
 a22883a <=( A232  and  (not A203) );
 a22884a <=( (not A202)  and  a22883a );
 a22885a <=( a22884a  and  a22879a );
 a22889a <=( (not A268)  and  A265 );
 a22890a <=( A233  and  a22889a );
 a22894a <=( A299  and  A298 );
 a22895a <=( (not A269)  and  a22894a );
 a22896a <=( a22895a  and  a22890a );
 a22900a <=( (not A200)  and  A166 );
 a22901a <=( A168  and  a22900a );
 a22905a <=( A232  and  (not A203) );
 a22906a <=( (not A202)  and  a22905a );
 a22907a <=( a22906a  and  a22901a );
 a22911a <=( (not A268)  and  A265 );
 a22912a <=( A233  and  a22911a );
 a22916a <=( (not A299)  and  (not A298) );
 a22917a <=( (not A269)  and  a22916a );
 a22918a <=( a22917a  and  a22912a );
 a22922a <=( (not A200)  and  A166 );
 a22923a <=( A168  and  a22922a );
 a22927a <=( A232  and  (not A203) );
 a22928a <=( (not A202)  and  a22927a );
 a22929a <=( a22928a  and  a22923a );
 a22933a <=( (not A267)  and  A265 );
 a22934a <=( A233  and  a22933a );
 a22938a <=( (not A302)  and  (not A301) );
 a22939a <=( (not A299)  and  a22938a );
 a22940a <=( a22939a  and  a22934a );
 a22944a <=( (not A200)  and  A166 );
 a22945a <=( A168  and  a22944a );
 a22949a <=( A232  and  (not A203) );
 a22950a <=( (not A202)  and  a22949a );
 a22951a <=( a22950a  and  a22945a );
 a22955a <=( A266  and  A265 );
 a22956a <=( A233  and  a22955a );
 a22960a <=( (not A302)  and  (not A301) );
 a22961a <=( (not A299)  and  a22960a );
 a22962a <=( a22961a  and  a22956a );
 a22966a <=( (not A200)  and  A166 );
 a22967a <=( A168  and  a22966a );
 a22971a <=( A232  and  (not A203) );
 a22972a <=( (not A202)  and  a22971a );
 a22973a <=( a22972a  and  a22967a );
 a22977a <=( (not A266)  and  (not A265) );
 a22978a <=( A233  and  a22977a );
 a22982a <=( (not A302)  and  (not A301) );
 a22983a <=( (not A299)  and  a22982a );
 a22984a <=( a22983a  and  a22978a );
 a22988a <=( (not A200)  and  A166 );
 a22989a <=( A168  and  a22988a );
 a22993a <=( (not A233)  and  (not A203) );
 a22994a <=( (not A202)  and  a22993a );
 a22995a <=( a22994a  and  a22989a );
 a22999a <=( A265  and  (not A236) );
 a23000a <=( (not A235)  and  a22999a );
 a23004a <=( (not A300)  and  A298 );
 a23005a <=( A266  and  a23004a );
 a23006a <=( a23005a  and  a23000a );
 a23010a <=( (not A200)  and  A166 );
 a23011a <=( A168  and  a23010a );
 a23015a <=( (not A233)  and  (not A203) );
 a23016a <=( (not A202)  and  a23015a );
 a23017a <=( a23016a  and  a23011a );
 a23021a <=( A265  and  (not A236) );
 a23022a <=( (not A235)  and  a23021a );
 a23026a <=( A299  and  A298 );
 a23027a <=( A266  and  a23026a );
 a23028a <=( a23027a  and  a23022a );
 a23032a <=( (not A200)  and  A166 );
 a23033a <=( A168  and  a23032a );
 a23037a <=( (not A233)  and  (not A203) );
 a23038a <=( (not A202)  and  a23037a );
 a23039a <=( a23038a  and  a23033a );
 a23043a <=( A265  and  (not A236) );
 a23044a <=( (not A235)  and  a23043a );
 a23048a <=( (not A299)  and  (not A298) );
 a23049a <=( A266  and  a23048a );
 a23050a <=( a23049a  and  a23044a );
 a23054a <=( (not A200)  and  A166 );
 a23055a <=( A168  and  a23054a );
 a23059a <=( (not A233)  and  (not A203) );
 a23060a <=( (not A202)  and  a23059a );
 a23061a <=( a23060a  and  a23055a );
 a23065a <=( (not A266)  and  (not A236) );
 a23066a <=( (not A235)  and  a23065a );
 a23070a <=( (not A300)  and  A298 );
 a23071a <=( (not A267)  and  a23070a );
 a23072a <=( a23071a  and  a23066a );
 a23076a <=( (not A200)  and  A166 );
 a23077a <=( A168  and  a23076a );
 a23081a <=( (not A233)  and  (not A203) );
 a23082a <=( (not A202)  and  a23081a );
 a23083a <=( a23082a  and  a23077a );
 a23087a <=( (not A266)  and  (not A236) );
 a23088a <=( (not A235)  and  a23087a );
 a23092a <=( A299  and  A298 );
 a23093a <=( (not A267)  and  a23092a );
 a23094a <=( a23093a  and  a23088a );
 a23098a <=( (not A200)  and  A166 );
 a23099a <=( A168  and  a23098a );
 a23103a <=( (not A233)  and  (not A203) );
 a23104a <=( (not A202)  and  a23103a );
 a23105a <=( a23104a  and  a23099a );
 a23109a <=( (not A266)  and  (not A236) );
 a23110a <=( (not A235)  and  a23109a );
 a23114a <=( (not A299)  and  (not A298) );
 a23115a <=( (not A267)  and  a23114a );
 a23116a <=( a23115a  and  a23110a );
 a23120a <=( (not A200)  and  A166 );
 a23121a <=( A168  and  a23120a );
 a23125a <=( (not A233)  and  (not A203) );
 a23126a <=( (not A202)  and  a23125a );
 a23127a <=( a23126a  and  a23121a );
 a23131a <=( (not A265)  and  (not A236) );
 a23132a <=( (not A235)  and  a23131a );
 a23136a <=( (not A300)  and  A298 );
 a23137a <=( (not A266)  and  a23136a );
 a23138a <=( a23137a  and  a23132a );
 a23142a <=( (not A200)  and  A166 );
 a23143a <=( A168  and  a23142a );
 a23147a <=( (not A233)  and  (not A203) );
 a23148a <=( (not A202)  and  a23147a );
 a23149a <=( a23148a  and  a23143a );
 a23153a <=( (not A265)  and  (not A236) );
 a23154a <=( (not A235)  and  a23153a );
 a23158a <=( A299  and  A298 );
 a23159a <=( (not A266)  and  a23158a );
 a23160a <=( a23159a  and  a23154a );
 a23164a <=( (not A200)  and  A166 );
 a23165a <=( A168  and  a23164a );
 a23169a <=( (not A233)  and  (not A203) );
 a23170a <=( (not A202)  and  a23169a );
 a23171a <=( a23170a  and  a23165a );
 a23175a <=( (not A265)  and  (not A236) );
 a23176a <=( (not A235)  and  a23175a );
 a23180a <=( (not A299)  and  (not A298) );
 a23181a <=( (not A266)  and  a23180a );
 a23182a <=( a23181a  and  a23176a );
 a23186a <=( (not A200)  and  A166 );
 a23187a <=( A168  and  a23186a );
 a23191a <=( (not A233)  and  (not A203) );
 a23192a <=( (not A202)  and  a23191a );
 a23193a <=( a23192a  and  a23187a );
 a23197a <=( A266  and  A265 );
 a23198a <=( (not A234)  and  a23197a );
 a23202a <=( (not A302)  and  (not A301) );
 a23203a <=( A298  and  a23202a );
 a23204a <=( a23203a  and  a23198a );
 a23208a <=( (not A200)  and  A166 );
 a23209a <=( A168  and  a23208a );
 a23213a <=( (not A233)  and  (not A203) );
 a23214a <=( (not A202)  and  a23213a );
 a23215a <=( a23214a  and  a23209a );
 a23219a <=( (not A268)  and  (not A266) );
 a23220a <=( (not A234)  and  a23219a );
 a23224a <=( (not A300)  and  A298 );
 a23225a <=( (not A269)  and  a23224a );
 a23226a <=( a23225a  and  a23220a );
 a23230a <=( (not A200)  and  A166 );
 a23231a <=( A168  and  a23230a );
 a23235a <=( (not A233)  and  (not A203) );
 a23236a <=( (not A202)  and  a23235a );
 a23237a <=( a23236a  and  a23231a );
 a23241a <=( (not A268)  and  (not A266) );
 a23242a <=( (not A234)  and  a23241a );
 a23246a <=( A299  and  A298 );
 a23247a <=( (not A269)  and  a23246a );
 a23248a <=( a23247a  and  a23242a );
 a23252a <=( (not A200)  and  A166 );
 a23253a <=( A168  and  a23252a );
 a23257a <=( (not A233)  and  (not A203) );
 a23258a <=( (not A202)  and  a23257a );
 a23259a <=( a23258a  and  a23253a );
 a23263a <=( (not A268)  and  (not A266) );
 a23264a <=( (not A234)  and  a23263a );
 a23268a <=( (not A299)  and  (not A298) );
 a23269a <=( (not A269)  and  a23268a );
 a23270a <=( a23269a  and  a23264a );
 a23274a <=( (not A200)  and  A166 );
 a23275a <=( A168  and  a23274a );
 a23279a <=( (not A233)  and  (not A203) );
 a23280a <=( (not A202)  and  a23279a );
 a23281a <=( a23280a  and  a23275a );
 a23285a <=( (not A267)  and  (not A266) );
 a23286a <=( (not A234)  and  a23285a );
 a23290a <=( (not A302)  and  (not A301) );
 a23291a <=( A298  and  a23290a );
 a23292a <=( a23291a  and  a23286a );
 a23296a <=( (not A200)  and  A166 );
 a23297a <=( A168  and  a23296a );
 a23301a <=( (not A233)  and  (not A203) );
 a23302a <=( (not A202)  and  a23301a );
 a23303a <=( a23302a  and  a23297a );
 a23307a <=( (not A266)  and  (not A265) );
 a23308a <=( (not A234)  and  a23307a );
 a23312a <=( (not A302)  and  (not A301) );
 a23313a <=( A298  and  a23312a );
 a23314a <=( a23313a  and  a23308a );
 a23318a <=( (not A200)  and  A166 );
 a23319a <=( A168  and  a23318a );
 a23323a <=( (not A232)  and  (not A203) );
 a23324a <=( (not A202)  and  a23323a );
 a23325a <=( a23324a  and  a23319a );
 a23329a <=( A266  and  A265 );
 a23330a <=( (not A233)  and  a23329a );
 a23334a <=( (not A302)  and  (not A301) );
 a23335a <=( A298  and  a23334a );
 a23336a <=( a23335a  and  a23330a );
 a23340a <=( (not A200)  and  A166 );
 a23341a <=( A168  and  a23340a );
 a23345a <=( (not A232)  and  (not A203) );
 a23346a <=( (not A202)  and  a23345a );
 a23347a <=( a23346a  and  a23341a );
 a23351a <=( (not A268)  and  (not A266) );
 a23352a <=( (not A233)  and  a23351a );
 a23356a <=( (not A300)  and  A298 );
 a23357a <=( (not A269)  and  a23356a );
 a23358a <=( a23357a  and  a23352a );
 a23362a <=( (not A200)  and  A166 );
 a23363a <=( A168  and  a23362a );
 a23367a <=( (not A232)  and  (not A203) );
 a23368a <=( (not A202)  and  a23367a );
 a23369a <=( a23368a  and  a23363a );
 a23373a <=( (not A268)  and  (not A266) );
 a23374a <=( (not A233)  and  a23373a );
 a23378a <=( A299  and  A298 );
 a23379a <=( (not A269)  and  a23378a );
 a23380a <=( a23379a  and  a23374a );
 a23384a <=( (not A200)  and  A166 );
 a23385a <=( A168  and  a23384a );
 a23389a <=( (not A232)  and  (not A203) );
 a23390a <=( (not A202)  and  a23389a );
 a23391a <=( a23390a  and  a23385a );
 a23395a <=( (not A268)  and  (not A266) );
 a23396a <=( (not A233)  and  a23395a );
 a23400a <=( (not A299)  and  (not A298) );
 a23401a <=( (not A269)  and  a23400a );
 a23402a <=( a23401a  and  a23396a );
 a23406a <=( (not A200)  and  A166 );
 a23407a <=( A168  and  a23406a );
 a23411a <=( (not A232)  and  (not A203) );
 a23412a <=( (not A202)  and  a23411a );
 a23413a <=( a23412a  and  a23407a );
 a23417a <=( (not A267)  and  (not A266) );
 a23418a <=( (not A233)  and  a23417a );
 a23422a <=( (not A302)  and  (not A301) );
 a23423a <=( A298  and  a23422a );
 a23424a <=( a23423a  and  a23418a );
 a23428a <=( (not A200)  and  A166 );
 a23429a <=( A168  and  a23428a );
 a23433a <=( (not A232)  and  (not A203) );
 a23434a <=( (not A202)  and  a23433a );
 a23435a <=( a23434a  and  a23429a );
 a23439a <=( (not A266)  and  (not A265) );
 a23440a <=( (not A233)  and  a23439a );
 a23444a <=( (not A302)  and  (not A301) );
 a23445a <=( A298  and  a23444a );
 a23446a <=( a23445a  and  a23440a );
 a23450a <=( (not A200)  and  A166 );
 a23451a <=( A168  and  a23450a );
 a23455a <=( A233  and  A232 );
 a23456a <=( (not A201)  and  a23455a );
 a23457a <=( a23456a  and  a23451a );
 a23461a <=( (not A269)  and  (not A268) );
 a23462a <=( A265  and  a23461a );
 a23466a <=( (not A302)  and  (not A301) );
 a23467a <=( (not A299)  and  a23466a );
 a23468a <=( a23467a  and  a23462a );
 a23472a <=( (not A200)  and  A166 );
 a23473a <=( A168  and  a23472a );
 a23477a <=( (not A235)  and  (not A233) );
 a23478a <=( (not A201)  and  a23477a );
 a23479a <=( a23478a  and  a23473a );
 a23483a <=( A266  and  A265 );
 a23484a <=( (not A236)  and  a23483a );
 a23488a <=( (not A302)  and  (not A301) );
 a23489a <=( A298  and  a23488a );
 a23490a <=( a23489a  and  a23484a );
 a23494a <=( (not A200)  and  A166 );
 a23495a <=( A168  and  a23494a );
 a23499a <=( (not A235)  and  (not A233) );
 a23500a <=( (not A201)  and  a23499a );
 a23501a <=( a23500a  and  a23495a );
 a23505a <=( (not A268)  and  (not A266) );
 a23506a <=( (not A236)  and  a23505a );
 a23510a <=( (not A300)  and  A298 );
 a23511a <=( (not A269)  and  a23510a );
 a23512a <=( a23511a  and  a23506a );
 a23516a <=( (not A200)  and  A166 );
 a23517a <=( A168  and  a23516a );
 a23521a <=( (not A235)  and  (not A233) );
 a23522a <=( (not A201)  and  a23521a );
 a23523a <=( a23522a  and  a23517a );
 a23527a <=( (not A268)  and  (not A266) );
 a23528a <=( (not A236)  and  a23527a );
 a23532a <=( A299  and  A298 );
 a23533a <=( (not A269)  and  a23532a );
 a23534a <=( a23533a  and  a23528a );
 a23538a <=( (not A200)  and  A166 );
 a23539a <=( A168  and  a23538a );
 a23543a <=( (not A235)  and  (not A233) );
 a23544a <=( (not A201)  and  a23543a );
 a23545a <=( a23544a  and  a23539a );
 a23549a <=( (not A268)  and  (not A266) );
 a23550a <=( (not A236)  and  a23549a );
 a23554a <=( (not A299)  and  (not A298) );
 a23555a <=( (not A269)  and  a23554a );
 a23556a <=( a23555a  and  a23550a );
 a23560a <=( (not A200)  and  A166 );
 a23561a <=( A168  and  a23560a );
 a23565a <=( (not A235)  and  (not A233) );
 a23566a <=( (not A201)  and  a23565a );
 a23567a <=( a23566a  and  a23561a );
 a23571a <=( (not A267)  and  (not A266) );
 a23572a <=( (not A236)  and  a23571a );
 a23576a <=( (not A302)  and  (not A301) );
 a23577a <=( A298  and  a23576a );
 a23578a <=( a23577a  and  a23572a );
 a23582a <=( (not A200)  and  A166 );
 a23583a <=( A168  and  a23582a );
 a23587a <=( (not A235)  and  (not A233) );
 a23588a <=( (not A201)  and  a23587a );
 a23589a <=( a23588a  and  a23583a );
 a23593a <=( (not A266)  and  (not A265) );
 a23594a <=( (not A236)  and  a23593a );
 a23598a <=( (not A302)  and  (not A301) );
 a23599a <=( A298  and  a23598a );
 a23600a <=( a23599a  and  a23594a );
 a23604a <=( (not A200)  and  A166 );
 a23605a <=( A168  and  a23604a );
 a23609a <=( (not A234)  and  (not A233) );
 a23610a <=( (not A201)  and  a23609a );
 a23611a <=( a23610a  and  a23605a );
 a23615a <=( (not A269)  and  (not A268) );
 a23616a <=( (not A266)  and  a23615a );
 a23620a <=( (not A302)  and  (not A301) );
 a23621a <=( A298  and  a23620a );
 a23622a <=( a23621a  and  a23616a );
 a23626a <=( (not A200)  and  A166 );
 a23627a <=( A168  and  a23626a );
 a23631a <=( (not A233)  and  A232 );
 a23632a <=( (not A201)  and  a23631a );
 a23633a <=( a23632a  and  a23627a );
 a23637a <=( A298  and  A235 );
 a23638a <=( A234  and  a23637a );
 a23642a <=( A301  and  A300 );
 a23643a <=( (not A299)  and  a23642a );
 a23644a <=( a23643a  and  a23638a );
 a23648a <=( (not A200)  and  A166 );
 a23649a <=( A168  and  a23648a );
 a23653a <=( (not A233)  and  A232 );
 a23654a <=( (not A201)  and  a23653a );
 a23655a <=( a23654a  and  a23649a );
 a23659a <=( A298  and  A235 );
 a23660a <=( A234  and  a23659a );
 a23664a <=( A302  and  A300 );
 a23665a <=( (not A299)  and  a23664a );
 a23666a <=( a23665a  and  a23660a );
 a23670a <=( (not A200)  and  A166 );
 a23671a <=( A168  and  a23670a );
 a23675a <=( (not A233)  and  A232 );
 a23676a <=( (not A201)  and  a23675a );
 a23677a <=( a23676a  and  a23671a );
 a23681a <=( A265  and  A235 );
 a23682a <=( A234  and  a23681a );
 a23686a <=( A268  and  A267 );
 a23687a <=( (not A266)  and  a23686a );
 a23688a <=( a23687a  and  a23682a );
 a23692a <=( (not A200)  and  A166 );
 a23693a <=( A168  and  a23692a );
 a23697a <=( (not A233)  and  A232 );
 a23698a <=( (not A201)  and  a23697a );
 a23699a <=( a23698a  and  a23693a );
 a23703a <=( A265  and  A235 );
 a23704a <=( A234  and  a23703a );
 a23708a <=( A269  and  A267 );
 a23709a <=( (not A266)  and  a23708a );
 a23710a <=( a23709a  and  a23704a );
 a23714a <=( (not A200)  and  A166 );
 a23715a <=( A168  and  a23714a );
 a23719a <=( (not A233)  and  A232 );
 a23720a <=( (not A201)  and  a23719a );
 a23721a <=( a23720a  and  a23715a );
 a23725a <=( A298  and  A236 );
 a23726a <=( A234  and  a23725a );
 a23730a <=( A301  and  A300 );
 a23731a <=( (not A299)  and  a23730a );
 a23732a <=( a23731a  and  a23726a );
 a23736a <=( (not A200)  and  A166 );
 a23737a <=( A168  and  a23736a );
 a23741a <=( (not A233)  and  A232 );
 a23742a <=( (not A201)  and  a23741a );
 a23743a <=( a23742a  and  a23737a );
 a23747a <=( A298  and  A236 );
 a23748a <=( A234  and  a23747a );
 a23752a <=( A302  and  A300 );
 a23753a <=( (not A299)  and  a23752a );
 a23754a <=( a23753a  and  a23748a );
 a23758a <=( (not A200)  and  A166 );
 a23759a <=( A168  and  a23758a );
 a23763a <=( (not A233)  and  A232 );
 a23764a <=( (not A201)  and  a23763a );
 a23765a <=( a23764a  and  a23759a );
 a23769a <=( A265  and  A236 );
 a23770a <=( A234  and  a23769a );
 a23774a <=( A268  and  A267 );
 a23775a <=( (not A266)  and  a23774a );
 a23776a <=( a23775a  and  a23770a );
 a23780a <=( (not A200)  and  A166 );
 a23781a <=( A168  and  a23780a );
 a23785a <=( (not A233)  and  A232 );
 a23786a <=( (not A201)  and  a23785a );
 a23787a <=( a23786a  and  a23781a );
 a23791a <=( A265  and  A236 );
 a23792a <=( A234  and  a23791a );
 a23796a <=( A269  and  A267 );
 a23797a <=( (not A266)  and  a23796a );
 a23798a <=( a23797a  and  a23792a );
 a23802a <=( (not A200)  and  A166 );
 a23803a <=( A168  and  a23802a );
 a23807a <=( (not A233)  and  (not A232) );
 a23808a <=( (not A201)  and  a23807a );
 a23809a <=( a23808a  and  a23803a );
 a23813a <=( (not A269)  and  (not A268) );
 a23814a <=( (not A266)  and  a23813a );
 a23818a <=( (not A302)  and  (not A301) );
 a23819a <=( A298  and  a23818a );
 a23820a <=( a23819a  and  a23814a );
 a23824a <=( (not A199)  and  A166 );
 a23825a <=( A168  and  a23824a );
 a23829a <=( A233  and  A232 );
 a23830a <=( (not A200)  and  a23829a );
 a23831a <=( a23830a  and  a23825a );
 a23835a <=( (not A269)  and  (not A268) );
 a23836a <=( A265  and  a23835a );
 a23840a <=( (not A302)  and  (not A301) );
 a23841a <=( (not A299)  and  a23840a );
 a23842a <=( a23841a  and  a23836a );
 a23846a <=( (not A199)  and  A166 );
 a23847a <=( A168  and  a23846a );
 a23851a <=( (not A235)  and  (not A233) );
 a23852a <=( (not A200)  and  a23851a );
 a23853a <=( a23852a  and  a23847a );
 a23857a <=( A266  and  A265 );
 a23858a <=( (not A236)  and  a23857a );
 a23862a <=( (not A302)  and  (not A301) );
 a23863a <=( A298  and  a23862a );
 a23864a <=( a23863a  and  a23858a );
 a23868a <=( (not A199)  and  A166 );
 a23869a <=( A168  and  a23868a );
 a23873a <=( (not A235)  and  (not A233) );
 a23874a <=( (not A200)  and  a23873a );
 a23875a <=( a23874a  and  a23869a );
 a23879a <=( (not A268)  and  (not A266) );
 a23880a <=( (not A236)  and  a23879a );
 a23884a <=( (not A300)  and  A298 );
 a23885a <=( (not A269)  and  a23884a );
 a23886a <=( a23885a  and  a23880a );
 a23890a <=( (not A199)  and  A166 );
 a23891a <=( A168  and  a23890a );
 a23895a <=( (not A235)  and  (not A233) );
 a23896a <=( (not A200)  and  a23895a );
 a23897a <=( a23896a  and  a23891a );
 a23901a <=( (not A268)  and  (not A266) );
 a23902a <=( (not A236)  and  a23901a );
 a23906a <=( A299  and  A298 );
 a23907a <=( (not A269)  and  a23906a );
 a23908a <=( a23907a  and  a23902a );
 a23912a <=( (not A199)  and  A166 );
 a23913a <=( A168  and  a23912a );
 a23917a <=( (not A235)  and  (not A233) );
 a23918a <=( (not A200)  and  a23917a );
 a23919a <=( a23918a  and  a23913a );
 a23923a <=( (not A268)  and  (not A266) );
 a23924a <=( (not A236)  and  a23923a );
 a23928a <=( (not A299)  and  (not A298) );
 a23929a <=( (not A269)  and  a23928a );
 a23930a <=( a23929a  and  a23924a );
 a23934a <=( (not A199)  and  A166 );
 a23935a <=( A168  and  a23934a );
 a23939a <=( (not A235)  and  (not A233) );
 a23940a <=( (not A200)  and  a23939a );
 a23941a <=( a23940a  and  a23935a );
 a23945a <=( (not A267)  and  (not A266) );
 a23946a <=( (not A236)  and  a23945a );
 a23950a <=( (not A302)  and  (not A301) );
 a23951a <=( A298  and  a23950a );
 a23952a <=( a23951a  and  a23946a );
 a23956a <=( (not A199)  and  A166 );
 a23957a <=( A168  and  a23956a );
 a23961a <=( (not A235)  and  (not A233) );
 a23962a <=( (not A200)  and  a23961a );
 a23963a <=( a23962a  and  a23957a );
 a23967a <=( (not A266)  and  (not A265) );
 a23968a <=( (not A236)  and  a23967a );
 a23972a <=( (not A302)  and  (not A301) );
 a23973a <=( A298  and  a23972a );
 a23974a <=( a23973a  and  a23968a );
 a23978a <=( (not A199)  and  A166 );
 a23979a <=( A168  and  a23978a );
 a23983a <=( (not A234)  and  (not A233) );
 a23984a <=( (not A200)  and  a23983a );
 a23985a <=( a23984a  and  a23979a );
 a23989a <=( (not A269)  and  (not A268) );
 a23990a <=( (not A266)  and  a23989a );
 a23994a <=( (not A302)  and  (not A301) );
 a23995a <=( A298  and  a23994a );
 a23996a <=( a23995a  and  a23990a );
 a24000a <=( (not A199)  and  A166 );
 a24001a <=( A168  and  a24000a );
 a24005a <=( (not A233)  and  A232 );
 a24006a <=( (not A200)  and  a24005a );
 a24007a <=( a24006a  and  a24001a );
 a24011a <=( A298  and  A235 );
 a24012a <=( A234  and  a24011a );
 a24016a <=( A301  and  A300 );
 a24017a <=( (not A299)  and  a24016a );
 a24018a <=( a24017a  and  a24012a );
 a24022a <=( (not A199)  and  A166 );
 a24023a <=( A168  and  a24022a );
 a24027a <=( (not A233)  and  A232 );
 a24028a <=( (not A200)  and  a24027a );
 a24029a <=( a24028a  and  a24023a );
 a24033a <=( A298  and  A235 );
 a24034a <=( A234  and  a24033a );
 a24038a <=( A302  and  A300 );
 a24039a <=( (not A299)  and  a24038a );
 a24040a <=( a24039a  and  a24034a );
 a24044a <=( (not A199)  and  A166 );
 a24045a <=( A168  and  a24044a );
 a24049a <=( (not A233)  and  A232 );
 a24050a <=( (not A200)  and  a24049a );
 a24051a <=( a24050a  and  a24045a );
 a24055a <=( A265  and  A235 );
 a24056a <=( A234  and  a24055a );
 a24060a <=( A268  and  A267 );
 a24061a <=( (not A266)  and  a24060a );
 a24062a <=( a24061a  and  a24056a );
 a24066a <=( (not A199)  and  A166 );
 a24067a <=( A168  and  a24066a );
 a24071a <=( (not A233)  and  A232 );
 a24072a <=( (not A200)  and  a24071a );
 a24073a <=( a24072a  and  a24067a );
 a24077a <=( A265  and  A235 );
 a24078a <=( A234  and  a24077a );
 a24082a <=( A269  and  A267 );
 a24083a <=( (not A266)  and  a24082a );
 a24084a <=( a24083a  and  a24078a );
 a24088a <=( (not A199)  and  A166 );
 a24089a <=( A168  and  a24088a );
 a24093a <=( (not A233)  and  A232 );
 a24094a <=( (not A200)  and  a24093a );
 a24095a <=( a24094a  and  a24089a );
 a24099a <=( A298  and  A236 );
 a24100a <=( A234  and  a24099a );
 a24104a <=( A301  and  A300 );
 a24105a <=( (not A299)  and  a24104a );
 a24106a <=( a24105a  and  a24100a );
 a24110a <=( (not A199)  and  A166 );
 a24111a <=( A168  and  a24110a );
 a24115a <=( (not A233)  and  A232 );
 a24116a <=( (not A200)  and  a24115a );
 a24117a <=( a24116a  and  a24111a );
 a24121a <=( A298  and  A236 );
 a24122a <=( A234  and  a24121a );
 a24126a <=( A302  and  A300 );
 a24127a <=( (not A299)  and  a24126a );
 a24128a <=( a24127a  and  a24122a );
 a24132a <=( (not A199)  and  A166 );
 a24133a <=( A168  and  a24132a );
 a24137a <=( (not A233)  and  A232 );
 a24138a <=( (not A200)  and  a24137a );
 a24139a <=( a24138a  and  a24133a );
 a24143a <=( A265  and  A236 );
 a24144a <=( A234  and  a24143a );
 a24148a <=( A268  and  A267 );
 a24149a <=( (not A266)  and  a24148a );
 a24150a <=( a24149a  and  a24144a );
 a24154a <=( (not A199)  and  A166 );
 a24155a <=( A168  and  a24154a );
 a24159a <=( (not A233)  and  A232 );
 a24160a <=( (not A200)  and  a24159a );
 a24161a <=( a24160a  and  a24155a );
 a24165a <=( A265  and  A236 );
 a24166a <=( A234  and  a24165a );
 a24170a <=( A269  and  A267 );
 a24171a <=( (not A266)  and  a24170a );
 a24172a <=( a24171a  and  a24166a );
 a24176a <=( (not A199)  and  A166 );
 a24177a <=( A168  and  a24176a );
 a24181a <=( (not A233)  and  (not A232) );
 a24182a <=( (not A200)  and  a24181a );
 a24183a <=( a24182a  and  a24177a );
 a24187a <=( (not A269)  and  (not A268) );
 a24188a <=( (not A266)  and  a24187a );
 a24192a <=( (not A302)  and  (not A301) );
 a24193a <=( A298  and  a24192a );
 a24194a <=( a24193a  and  a24188a );
 a24198a <=( A199  and  A167 );
 a24199a <=( A168  and  a24198a );
 a24203a <=( A233  and  A232 );
 a24204a <=( A200  and  a24203a );
 a24205a <=( a24204a  and  a24199a );
 a24209a <=( (not A269)  and  (not A268) );
 a24210a <=( A265  and  a24209a );
 a24214a <=( (not A302)  and  (not A301) );
 a24215a <=( (not A299)  and  a24214a );
 a24216a <=( a24215a  and  a24210a );
 a24220a <=( A199  and  A167 );
 a24221a <=( A168  and  a24220a );
 a24225a <=( (not A235)  and  (not A233) );
 a24226a <=( A200  and  a24225a );
 a24227a <=( a24226a  and  a24221a );
 a24231a <=( A266  and  A265 );
 a24232a <=( (not A236)  and  a24231a );
 a24236a <=( (not A302)  and  (not A301) );
 a24237a <=( A298  and  a24236a );
 a24238a <=( a24237a  and  a24232a );
 a24242a <=( A199  and  A167 );
 a24243a <=( A168  and  a24242a );
 a24247a <=( (not A235)  and  (not A233) );
 a24248a <=( A200  and  a24247a );
 a24249a <=( a24248a  and  a24243a );
 a24253a <=( (not A268)  and  (not A266) );
 a24254a <=( (not A236)  and  a24253a );
 a24258a <=( (not A300)  and  A298 );
 a24259a <=( (not A269)  and  a24258a );
 a24260a <=( a24259a  and  a24254a );
 a24264a <=( A199  and  A167 );
 a24265a <=( A168  and  a24264a );
 a24269a <=( (not A235)  and  (not A233) );
 a24270a <=( A200  and  a24269a );
 a24271a <=( a24270a  and  a24265a );
 a24275a <=( (not A268)  and  (not A266) );
 a24276a <=( (not A236)  and  a24275a );
 a24280a <=( A299  and  A298 );
 a24281a <=( (not A269)  and  a24280a );
 a24282a <=( a24281a  and  a24276a );
 a24286a <=( A199  and  A167 );
 a24287a <=( A168  and  a24286a );
 a24291a <=( (not A235)  and  (not A233) );
 a24292a <=( A200  and  a24291a );
 a24293a <=( a24292a  and  a24287a );
 a24297a <=( (not A268)  and  (not A266) );
 a24298a <=( (not A236)  and  a24297a );
 a24302a <=( (not A299)  and  (not A298) );
 a24303a <=( (not A269)  and  a24302a );
 a24304a <=( a24303a  and  a24298a );
 a24308a <=( A199  and  A167 );
 a24309a <=( A168  and  a24308a );
 a24313a <=( (not A235)  and  (not A233) );
 a24314a <=( A200  and  a24313a );
 a24315a <=( a24314a  and  a24309a );
 a24319a <=( (not A267)  and  (not A266) );
 a24320a <=( (not A236)  and  a24319a );
 a24324a <=( (not A302)  and  (not A301) );
 a24325a <=( A298  and  a24324a );
 a24326a <=( a24325a  and  a24320a );
 a24330a <=( A199  and  A167 );
 a24331a <=( A168  and  a24330a );
 a24335a <=( (not A235)  and  (not A233) );
 a24336a <=( A200  and  a24335a );
 a24337a <=( a24336a  and  a24331a );
 a24341a <=( (not A266)  and  (not A265) );
 a24342a <=( (not A236)  and  a24341a );
 a24346a <=( (not A302)  and  (not A301) );
 a24347a <=( A298  and  a24346a );
 a24348a <=( a24347a  and  a24342a );
 a24352a <=( A199  and  A167 );
 a24353a <=( A168  and  a24352a );
 a24357a <=( (not A234)  and  (not A233) );
 a24358a <=( A200  and  a24357a );
 a24359a <=( a24358a  and  a24353a );
 a24363a <=( (not A269)  and  (not A268) );
 a24364a <=( (not A266)  and  a24363a );
 a24368a <=( (not A302)  and  (not A301) );
 a24369a <=( A298  and  a24368a );
 a24370a <=( a24369a  and  a24364a );
 a24374a <=( A199  and  A167 );
 a24375a <=( A168  and  a24374a );
 a24379a <=( (not A233)  and  A232 );
 a24380a <=( A200  and  a24379a );
 a24381a <=( a24380a  and  a24375a );
 a24385a <=( A298  and  A235 );
 a24386a <=( A234  and  a24385a );
 a24390a <=( A301  and  A300 );
 a24391a <=( (not A299)  and  a24390a );
 a24392a <=( a24391a  and  a24386a );
 a24396a <=( A199  and  A167 );
 a24397a <=( A168  and  a24396a );
 a24401a <=( (not A233)  and  A232 );
 a24402a <=( A200  and  a24401a );
 a24403a <=( a24402a  and  a24397a );
 a24407a <=( A298  and  A235 );
 a24408a <=( A234  and  a24407a );
 a24412a <=( A302  and  A300 );
 a24413a <=( (not A299)  and  a24412a );
 a24414a <=( a24413a  and  a24408a );
 a24418a <=( A199  and  A167 );
 a24419a <=( A168  and  a24418a );
 a24423a <=( (not A233)  and  A232 );
 a24424a <=( A200  and  a24423a );
 a24425a <=( a24424a  and  a24419a );
 a24429a <=( A265  and  A235 );
 a24430a <=( A234  and  a24429a );
 a24434a <=( A268  and  A267 );
 a24435a <=( (not A266)  and  a24434a );
 a24436a <=( a24435a  and  a24430a );
 a24440a <=( A199  and  A167 );
 a24441a <=( A168  and  a24440a );
 a24445a <=( (not A233)  and  A232 );
 a24446a <=( A200  and  a24445a );
 a24447a <=( a24446a  and  a24441a );
 a24451a <=( A265  and  A235 );
 a24452a <=( A234  and  a24451a );
 a24456a <=( A269  and  A267 );
 a24457a <=( (not A266)  and  a24456a );
 a24458a <=( a24457a  and  a24452a );
 a24462a <=( A199  and  A167 );
 a24463a <=( A168  and  a24462a );
 a24467a <=( (not A233)  and  A232 );
 a24468a <=( A200  and  a24467a );
 a24469a <=( a24468a  and  a24463a );
 a24473a <=( A298  and  A236 );
 a24474a <=( A234  and  a24473a );
 a24478a <=( A301  and  A300 );
 a24479a <=( (not A299)  and  a24478a );
 a24480a <=( a24479a  and  a24474a );
 a24484a <=( A199  and  A167 );
 a24485a <=( A168  and  a24484a );
 a24489a <=( (not A233)  and  A232 );
 a24490a <=( A200  and  a24489a );
 a24491a <=( a24490a  and  a24485a );
 a24495a <=( A298  and  A236 );
 a24496a <=( A234  and  a24495a );
 a24500a <=( A302  and  A300 );
 a24501a <=( (not A299)  and  a24500a );
 a24502a <=( a24501a  and  a24496a );
 a24506a <=( A199  and  A167 );
 a24507a <=( A168  and  a24506a );
 a24511a <=( (not A233)  and  A232 );
 a24512a <=( A200  and  a24511a );
 a24513a <=( a24512a  and  a24507a );
 a24517a <=( A265  and  A236 );
 a24518a <=( A234  and  a24517a );
 a24522a <=( A268  and  A267 );
 a24523a <=( (not A266)  and  a24522a );
 a24524a <=( a24523a  and  a24518a );
 a24528a <=( A199  and  A167 );
 a24529a <=( A168  and  a24528a );
 a24533a <=( (not A233)  and  A232 );
 a24534a <=( A200  and  a24533a );
 a24535a <=( a24534a  and  a24529a );
 a24539a <=( A265  and  A236 );
 a24540a <=( A234  and  a24539a );
 a24544a <=( A269  and  A267 );
 a24545a <=( (not A266)  and  a24544a );
 a24546a <=( a24545a  and  a24540a );
 a24550a <=( A199  and  A167 );
 a24551a <=( A168  and  a24550a );
 a24555a <=( (not A233)  and  (not A232) );
 a24556a <=( A200  and  a24555a );
 a24557a <=( a24556a  and  a24551a );
 a24561a <=( (not A269)  and  (not A268) );
 a24562a <=( (not A266)  and  a24561a );
 a24566a <=( (not A302)  and  (not A301) );
 a24567a <=( A298  and  a24566a );
 a24568a <=( a24567a  and  a24562a );
 a24572a <=( (not A200)  and  A167 );
 a24573a <=( A168  and  a24572a );
 a24577a <=( A232  and  (not A203) );
 a24578a <=( (not A202)  and  a24577a );
 a24579a <=( a24578a  and  a24573a );
 a24583a <=( (not A268)  and  A265 );
 a24584a <=( A233  and  a24583a );
 a24588a <=( (not A300)  and  (not A299) );
 a24589a <=( (not A269)  and  a24588a );
 a24590a <=( a24589a  and  a24584a );
 a24594a <=( (not A200)  and  A167 );
 a24595a <=( A168  and  a24594a );
 a24599a <=( A232  and  (not A203) );
 a24600a <=( (not A202)  and  a24599a );
 a24601a <=( a24600a  and  a24595a );
 a24605a <=( (not A268)  and  A265 );
 a24606a <=( A233  and  a24605a );
 a24610a <=( A299  and  A298 );
 a24611a <=( (not A269)  and  a24610a );
 a24612a <=( a24611a  and  a24606a );
 a24616a <=( (not A200)  and  A167 );
 a24617a <=( A168  and  a24616a );
 a24621a <=( A232  and  (not A203) );
 a24622a <=( (not A202)  and  a24621a );
 a24623a <=( a24622a  and  a24617a );
 a24627a <=( (not A268)  and  A265 );
 a24628a <=( A233  and  a24627a );
 a24632a <=( (not A299)  and  (not A298) );
 a24633a <=( (not A269)  and  a24632a );
 a24634a <=( a24633a  and  a24628a );
 a24638a <=( (not A200)  and  A167 );
 a24639a <=( A168  and  a24638a );
 a24643a <=( A232  and  (not A203) );
 a24644a <=( (not A202)  and  a24643a );
 a24645a <=( a24644a  and  a24639a );
 a24649a <=( (not A267)  and  A265 );
 a24650a <=( A233  and  a24649a );
 a24654a <=( (not A302)  and  (not A301) );
 a24655a <=( (not A299)  and  a24654a );
 a24656a <=( a24655a  and  a24650a );
 a24660a <=( (not A200)  and  A167 );
 a24661a <=( A168  and  a24660a );
 a24665a <=( A232  and  (not A203) );
 a24666a <=( (not A202)  and  a24665a );
 a24667a <=( a24666a  and  a24661a );
 a24671a <=( A266  and  A265 );
 a24672a <=( A233  and  a24671a );
 a24676a <=( (not A302)  and  (not A301) );
 a24677a <=( (not A299)  and  a24676a );
 a24678a <=( a24677a  and  a24672a );
 a24682a <=( (not A200)  and  A167 );
 a24683a <=( A168  and  a24682a );
 a24687a <=( A232  and  (not A203) );
 a24688a <=( (not A202)  and  a24687a );
 a24689a <=( a24688a  and  a24683a );
 a24693a <=( (not A266)  and  (not A265) );
 a24694a <=( A233  and  a24693a );
 a24698a <=( (not A302)  and  (not A301) );
 a24699a <=( (not A299)  and  a24698a );
 a24700a <=( a24699a  and  a24694a );
 a24704a <=( (not A200)  and  A167 );
 a24705a <=( A168  and  a24704a );
 a24709a <=( (not A233)  and  (not A203) );
 a24710a <=( (not A202)  and  a24709a );
 a24711a <=( a24710a  and  a24705a );
 a24715a <=( A265  and  (not A236) );
 a24716a <=( (not A235)  and  a24715a );
 a24720a <=( (not A300)  and  A298 );
 a24721a <=( A266  and  a24720a );
 a24722a <=( a24721a  and  a24716a );
 a24726a <=( (not A200)  and  A167 );
 a24727a <=( A168  and  a24726a );
 a24731a <=( (not A233)  and  (not A203) );
 a24732a <=( (not A202)  and  a24731a );
 a24733a <=( a24732a  and  a24727a );
 a24737a <=( A265  and  (not A236) );
 a24738a <=( (not A235)  and  a24737a );
 a24742a <=( A299  and  A298 );
 a24743a <=( A266  and  a24742a );
 a24744a <=( a24743a  and  a24738a );
 a24748a <=( (not A200)  and  A167 );
 a24749a <=( A168  and  a24748a );
 a24753a <=( (not A233)  and  (not A203) );
 a24754a <=( (not A202)  and  a24753a );
 a24755a <=( a24754a  and  a24749a );
 a24759a <=( A265  and  (not A236) );
 a24760a <=( (not A235)  and  a24759a );
 a24764a <=( (not A299)  and  (not A298) );
 a24765a <=( A266  and  a24764a );
 a24766a <=( a24765a  and  a24760a );
 a24770a <=( (not A200)  and  A167 );
 a24771a <=( A168  and  a24770a );
 a24775a <=( (not A233)  and  (not A203) );
 a24776a <=( (not A202)  and  a24775a );
 a24777a <=( a24776a  and  a24771a );
 a24781a <=( (not A266)  and  (not A236) );
 a24782a <=( (not A235)  and  a24781a );
 a24786a <=( (not A300)  and  A298 );
 a24787a <=( (not A267)  and  a24786a );
 a24788a <=( a24787a  and  a24782a );
 a24792a <=( (not A200)  and  A167 );
 a24793a <=( A168  and  a24792a );
 a24797a <=( (not A233)  and  (not A203) );
 a24798a <=( (not A202)  and  a24797a );
 a24799a <=( a24798a  and  a24793a );
 a24803a <=( (not A266)  and  (not A236) );
 a24804a <=( (not A235)  and  a24803a );
 a24808a <=( A299  and  A298 );
 a24809a <=( (not A267)  and  a24808a );
 a24810a <=( a24809a  and  a24804a );
 a24814a <=( (not A200)  and  A167 );
 a24815a <=( A168  and  a24814a );
 a24819a <=( (not A233)  and  (not A203) );
 a24820a <=( (not A202)  and  a24819a );
 a24821a <=( a24820a  and  a24815a );
 a24825a <=( (not A266)  and  (not A236) );
 a24826a <=( (not A235)  and  a24825a );
 a24830a <=( (not A299)  and  (not A298) );
 a24831a <=( (not A267)  and  a24830a );
 a24832a <=( a24831a  and  a24826a );
 a24836a <=( (not A200)  and  A167 );
 a24837a <=( A168  and  a24836a );
 a24841a <=( (not A233)  and  (not A203) );
 a24842a <=( (not A202)  and  a24841a );
 a24843a <=( a24842a  and  a24837a );
 a24847a <=( (not A265)  and  (not A236) );
 a24848a <=( (not A235)  and  a24847a );
 a24852a <=( (not A300)  and  A298 );
 a24853a <=( (not A266)  and  a24852a );
 a24854a <=( a24853a  and  a24848a );
 a24858a <=( (not A200)  and  A167 );
 a24859a <=( A168  and  a24858a );
 a24863a <=( (not A233)  and  (not A203) );
 a24864a <=( (not A202)  and  a24863a );
 a24865a <=( a24864a  and  a24859a );
 a24869a <=( (not A265)  and  (not A236) );
 a24870a <=( (not A235)  and  a24869a );
 a24874a <=( A299  and  A298 );
 a24875a <=( (not A266)  and  a24874a );
 a24876a <=( a24875a  and  a24870a );
 a24880a <=( (not A200)  and  A167 );
 a24881a <=( A168  and  a24880a );
 a24885a <=( (not A233)  and  (not A203) );
 a24886a <=( (not A202)  and  a24885a );
 a24887a <=( a24886a  and  a24881a );
 a24891a <=( (not A265)  and  (not A236) );
 a24892a <=( (not A235)  and  a24891a );
 a24896a <=( (not A299)  and  (not A298) );
 a24897a <=( (not A266)  and  a24896a );
 a24898a <=( a24897a  and  a24892a );
 a24902a <=( (not A200)  and  A167 );
 a24903a <=( A168  and  a24902a );
 a24907a <=( (not A233)  and  (not A203) );
 a24908a <=( (not A202)  and  a24907a );
 a24909a <=( a24908a  and  a24903a );
 a24913a <=( A266  and  A265 );
 a24914a <=( (not A234)  and  a24913a );
 a24918a <=( (not A302)  and  (not A301) );
 a24919a <=( A298  and  a24918a );
 a24920a <=( a24919a  and  a24914a );
 a24924a <=( (not A200)  and  A167 );
 a24925a <=( A168  and  a24924a );
 a24929a <=( (not A233)  and  (not A203) );
 a24930a <=( (not A202)  and  a24929a );
 a24931a <=( a24930a  and  a24925a );
 a24935a <=( (not A268)  and  (not A266) );
 a24936a <=( (not A234)  and  a24935a );
 a24940a <=( (not A300)  and  A298 );
 a24941a <=( (not A269)  and  a24940a );
 a24942a <=( a24941a  and  a24936a );
 a24946a <=( (not A200)  and  A167 );
 a24947a <=( A168  and  a24946a );
 a24951a <=( (not A233)  and  (not A203) );
 a24952a <=( (not A202)  and  a24951a );
 a24953a <=( a24952a  and  a24947a );
 a24957a <=( (not A268)  and  (not A266) );
 a24958a <=( (not A234)  and  a24957a );
 a24962a <=( A299  and  A298 );
 a24963a <=( (not A269)  and  a24962a );
 a24964a <=( a24963a  and  a24958a );
 a24968a <=( (not A200)  and  A167 );
 a24969a <=( A168  and  a24968a );
 a24973a <=( (not A233)  and  (not A203) );
 a24974a <=( (not A202)  and  a24973a );
 a24975a <=( a24974a  and  a24969a );
 a24979a <=( (not A268)  and  (not A266) );
 a24980a <=( (not A234)  and  a24979a );
 a24984a <=( (not A299)  and  (not A298) );
 a24985a <=( (not A269)  and  a24984a );
 a24986a <=( a24985a  and  a24980a );
 a24990a <=( (not A200)  and  A167 );
 a24991a <=( A168  and  a24990a );
 a24995a <=( (not A233)  and  (not A203) );
 a24996a <=( (not A202)  and  a24995a );
 a24997a <=( a24996a  and  a24991a );
 a25001a <=( (not A267)  and  (not A266) );
 a25002a <=( (not A234)  and  a25001a );
 a25006a <=( (not A302)  and  (not A301) );
 a25007a <=( A298  and  a25006a );
 a25008a <=( a25007a  and  a25002a );
 a25012a <=( (not A200)  and  A167 );
 a25013a <=( A168  and  a25012a );
 a25017a <=( (not A233)  and  (not A203) );
 a25018a <=( (not A202)  and  a25017a );
 a25019a <=( a25018a  and  a25013a );
 a25023a <=( (not A266)  and  (not A265) );
 a25024a <=( (not A234)  and  a25023a );
 a25028a <=( (not A302)  and  (not A301) );
 a25029a <=( A298  and  a25028a );
 a25030a <=( a25029a  and  a25024a );
 a25034a <=( (not A200)  and  A167 );
 a25035a <=( A168  and  a25034a );
 a25039a <=( (not A232)  and  (not A203) );
 a25040a <=( (not A202)  and  a25039a );
 a25041a <=( a25040a  and  a25035a );
 a25045a <=( A266  and  A265 );
 a25046a <=( (not A233)  and  a25045a );
 a25050a <=( (not A302)  and  (not A301) );
 a25051a <=( A298  and  a25050a );
 a25052a <=( a25051a  and  a25046a );
 a25056a <=( (not A200)  and  A167 );
 a25057a <=( A168  and  a25056a );
 a25061a <=( (not A232)  and  (not A203) );
 a25062a <=( (not A202)  and  a25061a );
 a25063a <=( a25062a  and  a25057a );
 a25067a <=( (not A268)  and  (not A266) );
 a25068a <=( (not A233)  and  a25067a );
 a25072a <=( (not A300)  and  A298 );
 a25073a <=( (not A269)  and  a25072a );
 a25074a <=( a25073a  and  a25068a );
 a25078a <=( (not A200)  and  A167 );
 a25079a <=( A168  and  a25078a );
 a25083a <=( (not A232)  and  (not A203) );
 a25084a <=( (not A202)  and  a25083a );
 a25085a <=( a25084a  and  a25079a );
 a25089a <=( (not A268)  and  (not A266) );
 a25090a <=( (not A233)  and  a25089a );
 a25094a <=( A299  and  A298 );
 a25095a <=( (not A269)  and  a25094a );
 a25096a <=( a25095a  and  a25090a );
 a25100a <=( (not A200)  and  A167 );
 a25101a <=( A168  and  a25100a );
 a25105a <=( (not A232)  and  (not A203) );
 a25106a <=( (not A202)  and  a25105a );
 a25107a <=( a25106a  and  a25101a );
 a25111a <=( (not A268)  and  (not A266) );
 a25112a <=( (not A233)  and  a25111a );
 a25116a <=( (not A299)  and  (not A298) );
 a25117a <=( (not A269)  and  a25116a );
 a25118a <=( a25117a  and  a25112a );
 a25122a <=( (not A200)  and  A167 );
 a25123a <=( A168  and  a25122a );
 a25127a <=( (not A232)  and  (not A203) );
 a25128a <=( (not A202)  and  a25127a );
 a25129a <=( a25128a  and  a25123a );
 a25133a <=( (not A267)  and  (not A266) );
 a25134a <=( (not A233)  and  a25133a );
 a25138a <=( (not A302)  and  (not A301) );
 a25139a <=( A298  and  a25138a );
 a25140a <=( a25139a  and  a25134a );
 a25144a <=( (not A200)  and  A167 );
 a25145a <=( A168  and  a25144a );
 a25149a <=( (not A232)  and  (not A203) );
 a25150a <=( (not A202)  and  a25149a );
 a25151a <=( a25150a  and  a25145a );
 a25155a <=( (not A266)  and  (not A265) );
 a25156a <=( (not A233)  and  a25155a );
 a25160a <=( (not A302)  and  (not A301) );
 a25161a <=( A298  and  a25160a );
 a25162a <=( a25161a  and  a25156a );
 a25166a <=( (not A200)  and  A167 );
 a25167a <=( A168  and  a25166a );
 a25171a <=( A233  and  A232 );
 a25172a <=( (not A201)  and  a25171a );
 a25173a <=( a25172a  and  a25167a );
 a25177a <=( (not A269)  and  (not A268) );
 a25178a <=( A265  and  a25177a );
 a25182a <=( (not A302)  and  (not A301) );
 a25183a <=( (not A299)  and  a25182a );
 a25184a <=( a25183a  and  a25178a );
 a25188a <=( (not A200)  and  A167 );
 a25189a <=( A168  and  a25188a );
 a25193a <=( (not A235)  and  (not A233) );
 a25194a <=( (not A201)  and  a25193a );
 a25195a <=( a25194a  and  a25189a );
 a25199a <=( A266  and  A265 );
 a25200a <=( (not A236)  and  a25199a );
 a25204a <=( (not A302)  and  (not A301) );
 a25205a <=( A298  and  a25204a );
 a25206a <=( a25205a  and  a25200a );
 a25210a <=( (not A200)  and  A167 );
 a25211a <=( A168  and  a25210a );
 a25215a <=( (not A235)  and  (not A233) );
 a25216a <=( (not A201)  and  a25215a );
 a25217a <=( a25216a  and  a25211a );
 a25221a <=( (not A268)  and  (not A266) );
 a25222a <=( (not A236)  and  a25221a );
 a25226a <=( (not A300)  and  A298 );
 a25227a <=( (not A269)  and  a25226a );
 a25228a <=( a25227a  and  a25222a );
 a25232a <=( (not A200)  and  A167 );
 a25233a <=( A168  and  a25232a );
 a25237a <=( (not A235)  and  (not A233) );
 a25238a <=( (not A201)  and  a25237a );
 a25239a <=( a25238a  and  a25233a );
 a25243a <=( (not A268)  and  (not A266) );
 a25244a <=( (not A236)  and  a25243a );
 a25248a <=( A299  and  A298 );
 a25249a <=( (not A269)  and  a25248a );
 a25250a <=( a25249a  and  a25244a );
 a25254a <=( (not A200)  and  A167 );
 a25255a <=( A168  and  a25254a );
 a25259a <=( (not A235)  and  (not A233) );
 a25260a <=( (not A201)  and  a25259a );
 a25261a <=( a25260a  and  a25255a );
 a25265a <=( (not A268)  and  (not A266) );
 a25266a <=( (not A236)  and  a25265a );
 a25270a <=( (not A299)  and  (not A298) );
 a25271a <=( (not A269)  and  a25270a );
 a25272a <=( a25271a  and  a25266a );
 a25276a <=( (not A200)  and  A167 );
 a25277a <=( A168  and  a25276a );
 a25281a <=( (not A235)  and  (not A233) );
 a25282a <=( (not A201)  and  a25281a );
 a25283a <=( a25282a  and  a25277a );
 a25287a <=( (not A267)  and  (not A266) );
 a25288a <=( (not A236)  and  a25287a );
 a25292a <=( (not A302)  and  (not A301) );
 a25293a <=( A298  and  a25292a );
 a25294a <=( a25293a  and  a25288a );
 a25298a <=( (not A200)  and  A167 );
 a25299a <=( A168  and  a25298a );
 a25303a <=( (not A235)  and  (not A233) );
 a25304a <=( (not A201)  and  a25303a );
 a25305a <=( a25304a  and  a25299a );
 a25309a <=( (not A266)  and  (not A265) );
 a25310a <=( (not A236)  and  a25309a );
 a25314a <=( (not A302)  and  (not A301) );
 a25315a <=( A298  and  a25314a );
 a25316a <=( a25315a  and  a25310a );
 a25320a <=( (not A200)  and  A167 );
 a25321a <=( A168  and  a25320a );
 a25325a <=( (not A234)  and  (not A233) );
 a25326a <=( (not A201)  and  a25325a );
 a25327a <=( a25326a  and  a25321a );
 a25331a <=( (not A269)  and  (not A268) );
 a25332a <=( (not A266)  and  a25331a );
 a25336a <=( (not A302)  and  (not A301) );
 a25337a <=( A298  and  a25336a );
 a25338a <=( a25337a  and  a25332a );
 a25342a <=( (not A200)  and  A167 );
 a25343a <=( A168  and  a25342a );
 a25347a <=( (not A233)  and  A232 );
 a25348a <=( (not A201)  and  a25347a );
 a25349a <=( a25348a  and  a25343a );
 a25353a <=( A298  and  A235 );
 a25354a <=( A234  and  a25353a );
 a25358a <=( A301  and  A300 );
 a25359a <=( (not A299)  and  a25358a );
 a25360a <=( a25359a  and  a25354a );
 a25364a <=( (not A200)  and  A167 );
 a25365a <=( A168  and  a25364a );
 a25369a <=( (not A233)  and  A232 );
 a25370a <=( (not A201)  and  a25369a );
 a25371a <=( a25370a  and  a25365a );
 a25375a <=( A298  and  A235 );
 a25376a <=( A234  and  a25375a );
 a25380a <=( A302  and  A300 );
 a25381a <=( (not A299)  and  a25380a );
 a25382a <=( a25381a  and  a25376a );
 a25386a <=( (not A200)  and  A167 );
 a25387a <=( A168  and  a25386a );
 a25391a <=( (not A233)  and  A232 );
 a25392a <=( (not A201)  and  a25391a );
 a25393a <=( a25392a  and  a25387a );
 a25397a <=( A265  and  A235 );
 a25398a <=( A234  and  a25397a );
 a25402a <=( A268  and  A267 );
 a25403a <=( (not A266)  and  a25402a );
 a25404a <=( a25403a  and  a25398a );
 a25408a <=( (not A200)  and  A167 );
 a25409a <=( A168  and  a25408a );
 a25413a <=( (not A233)  and  A232 );
 a25414a <=( (not A201)  and  a25413a );
 a25415a <=( a25414a  and  a25409a );
 a25419a <=( A265  and  A235 );
 a25420a <=( A234  and  a25419a );
 a25424a <=( A269  and  A267 );
 a25425a <=( (not A266)  and  a25424a );
 a25426a <=( a25425a  and  a25420a );
 a25430a <=( (not A200)  and  A167 );
 a25431a <=( A168  and  a25430a );
 a25435a <=( (not A233)  and  A232 );
 a25436a <=( (not A201)  and  a25435a );
 a25437a <=( a25436a  and  a25431a );
 a25441a <=( A298  and  A236 );
 a25442a <=( A234  and  a25441a );
 a25446a <=( A301  and  A300 );
 a25447a <=( (not A299)  and  a25446a );
 a25448a <=( a25447a  and  a25442a );
 a25452a <=( (not A200)  and  A167 );
 a25453a <=( A168  and  a25452a );
 a25457a <=( (not A233)  and  A232 );
 a25458a <=( (not A201)  and  a25457a );
 a25459a <=( a25458a  and  a25453a );
 a25463a <=( A298  and  A236 );
 a25464a <=( A234  and  a25463a );
 a25468a <=( A302  and  A300 );
 a25469a <=( (not A299)  and  a25468a );
 a25470a <=( a25469a  and  a25464a );
 a25474a <=( (not A200)  and  A167 );
 a25475a <=( A168  and  a25474a );
 a25479a <=( (not A233)  and  A232 );
 a25480a <=( (not A201)  and  a25479a );
 a25481a <=( a25480a  and  a25475a );
 a25485a <=( A265  and  A236 );
 a25486a <=( A234  and  a25485a );
 a25490a <=( A268  and  A267 );
 a25491a <=( (not A266)  and  a25490a );
 a25492a <=( a25491a  and  a25486a );
 a25496a <=( (not A200)  and  A167 );
 a25497a <=( A168  and  a25496a );
 a25501a <=( (not A233)  and  A232 );
 a25502a <=( (not A201)  and  a25501a );
 a25503a <=( a25502a  and  a25497a );
 a25507a <=( A265  and  A236 );
 a25508a <=( A234  and  a25507a );
 a25512a <=( A269  and  A267 );
 a25513a <=( (not A266)  and  a25512a );
 a25514a <=( a25513a  and  a25508a );
 a25518a <=( (not A200)  and  A167 );
 a25519a <=( A168  and  a25518a );
 a25523a <=( (not A233)  and  (not A232) );
 a25524a <=( (not A201)  and  a25523a );
 a25525a <=( a25524a  and  a25519a );
 a25529a <=( (not A269)  and  (not A268) );
 a25530a <=( (not A266)  and  a25529a );
 a25534a <=( (not A302)  and  (not A301) );
 a25535a <=( A298  and  a25534a );
 a25536a <=( a25535a  and  a25530a );
 a25540a <=( (not A199)  and  A167 );
 a25541a <=( A168  and  a25540a );
 a25545a <=( A233  and  A232 );
 a25546a <=( (not A200)  and  a25545a );
 a25547a <=( a25546a  and  a25541a );
 a25551a <=( (not A269)  and  (not A268) );
 a25552a <=( A265  and  a25551a );
 a25556a <=( (not A302)  and  (not A301) );
 a25557a <=( (not A299)  and  a25556a );
 a25558a <=( a25557a  and  a25552a );
 a25562a <=( (not A199)  and  A167 );
 a25563a <=( A168  and  a25562a );
 a25567a <=( (not A235)  and  (not A233) );
 a25568a <=( (not A200)  and  a25567a );
 a25569a <=( a25568a  and  a25563a );
 a25573a <=( A266  and  A265 );
 a25574a <=( (not A236)  and  a25573a );
 a25578a <=( (not A302)  and  (not A301) );
 a25579a <=( A298  and  a25578a );
 a25580a <=( a25579a  and  a25574a );
 a25584a <=( (not A199)  and  A167 );
 a25585a <=( A168  and  a25584a );
 a25589a <=( (not A235)  and  (not A233) );
 a25590a <=( (not A200)  and  a25589a );
 a25591a <=( a25590a  and  a25585a );
 a25595a <=( (not A268)  and  (not A266) );
 a25596a <=( (not A236)  and  a25595a );
 a25600a <=( (not A300)  and  A298 );
 a25601a <=( (not A269)  and  a25600a );
 a25602a <=( a25601a  and  a25596a );
 a25606a <=( (not A199)  and  A167 );
 a25607a <=( A168  and  a25606a );
 a25611a <=( (not A235)  and  (not A233) );
 a25612a <=( (not A200)  and  a25611a );
 a25613a <=( a25612a  and  a25607a );
 a25617a <=( (not A268)  and  (not A266) );
 a25618a <=( (not A236)  and  a25617a );
 a25622a <=( A299  and  A298 );
 a25623a <=( (not A269)  and  a25622a );
 a25624a <=( a25623a  and  a25618a );
 a25628a <=( (not A199)  and  A167 );
 a25629a <=( A168  and  a25628a );
 a25633a <=( (not A235)  and  (not A233) );
 a25634a <=( (not A200)  and  a25633a );
 a25635a <=( a25634a  and  a25629a );
 a25639a <=( (not A268)  and  (not A266) );
 a25640a <=( (not A236)  and  a25639a );
 a25644a <=( (not A299)  and  (not A298) );
 a25645a <=( (not A269)  and  a25644a );
 a25646a <=( a25645a  and  a25640a );
 a25650a <=( (not A199)  and  A167 );
 a25651a <=( A168  and  a25650a );
 a25655a <=( (not A235)  and  (not A233) );
 a25656a <=( (not A200)  and  a25655a );
 a25657a <=( a25656a  and  a25651a );
 a25661a <=( (not A267)  and  (not A266) );
 a25662a <=( (not A236)  and  a25661a );
 a25666a <=( (not A302)  and  (not A301) );
 a25667a <=( A298  and  a25666a );
 a25668a <=( a25667a  and  a25662a );
 a25672a <=( (not A199)  and  A167 );
 a25673a <=( A168  and  a25672a );
 a25677a <=( (not A235)  and  (not A233) );
 a25678a <=( (not A200)  and  a25677a );
 a25679a <=( a25678a  and  a25673a );
 a25683a <=( (not A266)  and  (not A265) );
 a25684a <=( (not A236)  and  a25683a );
 a25688a <=( (not A302)  and  (not A301) );
 a25689a <=( A298  and  a25688a );
 a25690a <=( a25689a  and  a25684a );
 a25694a <=( (not A199)  and  A167 );
 a25695a <=( A168  and  a25694a );
 a25699a <=( (not A234)  and  (not A233) );
 a25700a <=( (not A200)  and  a25699a );
 a25701a <=( a25700a  and  a25695a );
 a25705a <=( (not A269)  and  (not A268) );
 a25706a <=( (not A266)  and  a25705a );
 a25710a <=( (not A302)  and  (not A301) );
 a25711a <=( A298  and  a25710a );
 a25712a <=( a25711a  and  a25706a );
 a25716a <=( (not A199)  and  A167 );
 a25717a <=( A168  and  a25716a );
 a25721a <=( (not A233)  and  A232 );
 a25722a <=( (not A200)  and  a25721a );
 a25723a <=( a25722a  and  a25717a );
 a25727a <=( A298  and  A235 );
 a25728a <=( A234  and  a25727a );
 a25732a <=( A301  and  A300 );
 a25733a <=( (not A299)  and  a25732a );
 a25734a <=( a25733a  and  a25728a );
 a25738a <=( (not A199)  and  A167 );
 a25739a <=( A168  and  a25738a );
 a25743a <=( (not A233)  and  A232 );
 a25744a <=( (not A200)  and  a25743a );
 a25745a <=( a25744a  and  a25739a );
 a25749a <=( A298  and  A235 );
 a25750a <=( A234  and  a25749a );
 a25754a <=( A302  and  A300 );
 a25755a <=( (not A299)  and  a25754a );
 a25756a <=( a25755a  and  a25750a );
 a25760a <=( (not A199)  and  A167 );
 a25761a <=( A168  and  a25760a );
 a25765a <=( (not A233)  and  A232 );
 a25766a <=( (not A200)  and  a25765a );
 a25767a <=( a25766a  and  a25761a );
 a25771a <=( A265  and  A235 );
 a25772a <=( A234  and  a25771a );
 a25776a <=( A268  and  A267 );
 a25777a <=( (not A266)  and  a25776a );
 a25778a <=( a25777a  and  a25772a );
 a25782a <=( (not A199)  and  A167 );
 a25783a <=( A168  and  a25782a );
 a25787a <=( (not A233)  and  A232 );
 a25788a <=( (not A200)  and  a25787a );
 a25789a <=( a25788a  and  a25783a );
 a25793a <=( A265  and  A235 );
 a25794a <=( A234  and  a25793a );
 a25798a <=( A269  and  A267 );
 a25799a <=( (not A266)  and  a25798a );
 a25800a <=( a25799a  and  a25794a );
 a25804a <=( (not A199)  and  A167 );
 a25805a <=( A168  and  a25804a );
 a25809a <=( (not A233)  and  A232 );
 a25810a <=( (not A200)  and  a25809a );
 a25811a <=( a25810a  and  a25805a );
 a25815a <=( A298  and  A236 );
 a25816a <=( A234  and  a25815a );
 a25820a <=( A301  and  A300 );
 a25821a <=( (not A299)  and  a25820a );
 a25822a <=( a25821a  and  a25816a );
 a25826a <=( (not A199)  and  A167 );
 a25827a <=( A168  and  a25826a );
 a25831a <=( (not A233)  and  A232 );
 a25832a <=( (not A200)  and  a25831a );
 a25833a <=( a25832a  and  a25827a );
 a25837a <=( A298  and  A236 );
 a25838a <=( A234  and  a25837a );
 a25842a <=( A302  and  A300 );
 a25843a <=( (not A299)  and  a25842a );
 a25844a <=( a25843a  and  a25838a );
 a25848a <=( (not A199)  and  A167 );
 a25849a <=( A168  and  a25848a );
 a25853a <=( (not A233)  and  A232 );
 a25854a <=( (not A200)  and  a25853a );
 a25855a <=( a25854a  and  a25849a );
 a25859a <=( A265  and  A236 );
 a25860a <=( A234  and  a25859a );
 a25864a <=( A268  and  A267 );
 a25865a <=( (not A266)  and  a25864a );
 a25866a <=( a25865a  and  a25860a );
 a25870a <=( (not A199)  and  A167 );
 a25871a <=( A168  and  a25870a );
 a25875a <=( (not A233)  and  A232 );
 a25876a <=( (not A200)  and  a25875a );
 a25877a <=( a25876a  and  a25871a );
 a25881a <=( A265  and  A236 );
 a25882a <=( A234  and  a25881a );
 a25886a <=( A269  and  A267 );
 a25887a <=( (not A266)  and  a25886a );
 a25888a <=( a25887a  and  a25882a );
 a25892a <=( (not A199)  and  A167 );
 a25893a <=( A168  and  a25892a );
 a25897a <=( (not A233)  and  (not A232) );
 a25898a <=( (not A200)  and  a25897a );
 a25899a <=( a25898a  and  a25893a );
 a25903a <=( (not A269)  and  (not A268) );
 a25904a <=( (not A266)  and  a25903a );
 a25908a <=( (not A302)  and  (not A301) );
 a25909a <=( A298  and  a25908a );
 a25910a <=( a25909a  and  a25904a );
 a25914a <=( (not A166)  and  (not A167) );
 a25915a <=( A170  and  a25914a );
 a25919a <=( A232  and  A200 );
 a25920a <=( (not A199)  and  a25919a );
 a25921a <=( a25920a  and  a25915a );
 a25925a <=( (not A268)  and  A265 );
 a25926a <=( A233  and  a25925a );
 a25930a <=( (not A300)  and  (not A299) );
 a25931a <=( (not A269)  and  a25930a );
 a25932a <=( a25931a  and  a25926a );
 a25936a <=( (not A166)  and  (not A167) );
 a25937a <=( A170  and  a25936a );
 a25941a <=( A232  and  A200 );
 a25942a <=( (not A199)  and  a25941a );
 a25943a <=( a25942a  and  a25937a );
 a25947a <=( (not A268)  and  A265 );
 a25948a <=( A233  and  a25947a );
 a25952a <=( A299  and  A298 );
 a25953a <=( (not A269)  and  a25952a );
 a25954a <=( a25953a  and  a25948a );
 a25958a <=( (not A166)  and  (not A167) );
 a25959a <=( A170  and  a25958a );
 a25963a <=( A232  and  A200 );
 a25964a <=( (not A199)  and  a25963a );
 a25965a <=( a25964a  and  a25959a );
 a25969a <=( (not A268)  and  A265 );
 a25970a <=( A233  and  a25969a );
 a25974a <=( (not A299)  and  (not A298) );
 a25975a <=( (not A269)  and  a25974a );
 a25976a <=( a25975a  and  a25970a );
 a25980a <=( (not A166)  and  (not A167) );
 a25981a <=( A170  and  a25980a );
 a25985a <=( A232  and  A200 );
 a25986a <=( (not A199)  and  a25985a );
 a25987a <=( a25986a  and  a25981a );
 a25991a <=( (not A267)  and  A265 );
 a25992a <=( A233  and  a25991a );
 a25996a <=( (not A302)  and  (not A301) );
 a25997a <=( (not A299)  and  a25996a );
 a25998a <=( a25997a  and  a25992a );
 a26002a <=( (not A166)  and  (not A167) );
 a26003a <=( A170  and  a26002a );
 a26007a <=( A232  and  A200 );
 a26008a <=( (not A199)  and  a26007a );
 a26009a <=( a26008a  and  a26003a );
 a26013a <=( A266  and  A265 );
 a26014a <=( A233  and  a26013a );
 a26018a <=( (not A302)  and  (not A301) );
 a26019a <=( (not A299)  and  a26018a );
 a26020a <=( a26019a  and  a26014a );
 a26024a <=( (not A166)  and  (not A167) );
 a26025a <=( A170  and  a26024a );
 a26029a <=( A232  and  A200 );
 a26030a <=( (not A199)  and  a26029a );
 a26031a <=( a26030a  and  a26025a );
 a26035a <=( (not A266)  and  (not A265) );
 a26036a <=( A233  and  a26035a );
 a26040a <=( (not A302)  and  (not A301) );
 a26041a <=( (not A299)  and  a26040a );
 a26042a <=( a26041a  and  a26036a );
 a26046a <=( (not A166)  and  (not A167) );
 a26047a <=( A170  and  a26046a );
 a26051a <=( (not A233)  and  A200 );
 a26052a <=( (not A199)  and  a26051a );
 a26053a <=( a26052a  and  a26047a );
 a26057a <=( A265  and  (not A236) );
 a26058a <=( (not A235)  and  a26057a );
 a26062a <=( (not A300)  and  A298 );
 a26063a <=( A266  and  a26062a );
 a26064a <=( a26063a  and  a26058a );
 a26068a <=( (not A166)  and  (not A167) );
 a26069a <=( A170  and  a26068a );
 a26073a <=( (not A233)  and  A200 );
 a26074a <=( (not A199)  and  a26073a );
 a26075a <=( a26074a  and  a26069a );
 a26079a <=( A265  and  (not A236) );
 a26080a <=( (not A235)  and  a26079a );
 a26084a <=( A299  and  A298 );
 a26085a <=( A266  and  a26084a );
 a26086a <=( a26085a  and  a26080a );
 a26090a <=( (not A166)  and  (not A167) );
 a26091a <=( A170  and  a26090a );
 a26095a <=( (not A233)  and  A200 );
 a26096a <=( (not A199)  and  a26095a );
 a26097a <=( a26096a  and  a26091a );
 a26101a <=( A265  and  (not A236) );
 a26102a <=( (not A235)  and  a26101a );
 a26106a <=( (not A299)  and  (not A298) );
 a26107a <=( A266  and  a26106a );
 a26108a <=( a26107a  and  a26102a );
 a26112a <=( (not A166)  and  (not A167) );
 a26113a <=( A170  and  a26112a );
 a26117a <=( (not A233)  and  A200 );
 a26118a <=( (not A199)  and  a26117a );
 a26119a <=( a26118a  and  a26113a );
 a26123a <=( (not A266)  and  (not A236) );
 a26124a <=( (not A235)  and  a26123a );
 a26128a <=( (not A300)  and  A298 );
 a26129a <=( (not A267)  and  a26128a );
 a26130a <=( a26129a  and  a26124a );
 a26134a <=( (not A166)  and  (not A167) );
 a26135a <=( A170  and  a26134a );
 a26139a <=( (not A233)  and  A200 );
 a26140a <=( (not A199)  and  a26139a );
 a26141a <=( a26140a  and  a26135a );
 a26145a <=( (not A266)  and  (not A236) );
 a26146a <=( (not A235)  and  a26145a );
 a26150a <=( A299  and  A298 );
 a26151a <=( (not A267)  and  a26150a );
 a26152a <=( a26151a  and  a26146a );
 a26156a <=( (not A166)  and  (not A167) );
 a26157a <=( A170  and  a26156a );
 a26161a <=( (not A233)  and  A200 );
 a26162a <=( (not A199)  and  a26161a );
 a26163a <=( a26162a  and  a26157a );
 a26167a <=( (not A266)  and  (not A236) );
 a26168a <=( (not A235)  and  a26167a );
 a26172a <=( (not A299)  and  (not A298) );
 a26173a <=( (not A267)  and  a26172a );
 a26174a <=( a26173a  and  a26168a );
 a26178a <=( (not A166)  and  (not A167) );
 a26179a <=( A170  and  a26178a );
 a26183a <=( (not A233)  and  A200 );
 a26184a <=( (not A199)  and  a26183a );
 a26185a <=( a26184a  and  a26179a );
 a26189a <=( (not A265)  and  (not A236) );
 a26190a <=( (not A235)  and  a26189a );
 a26194a <=( (not A300)  and  A298 );
 a26195a <=( (not A266)  and  a26194a );
 a26196a <=( a26195a  and  a26190a );
 a26200a <=( (not A166)  and  (not A167) );
 a26201a <=( A170  and  a26200a );
 a26205a <=( (not A233)  and  A200 );
 a26206a <=( (not A199)  and  a26205a );
 a26207a <=( a26206a  and  a26201a );
 a26211a <=( (not A265)  and  (not A236) );
 a26212a <=( (not A235)  and  a26211a );
 a26216a <=( A299  and  A298 );
 a26217a <=( (not A266)  and  a26216a );
 a26218a <=( a26217a  and  a26212a );
 a26222a <=( (not A166)  and  (not A167) );
 a26223a <=( A170  and  a26222a );
 a26227a <=( (not A233)  and  A200 );
 a26228a <=( (not A199)  and  a26227a );
 a26229a <=( a26228a  and  a26223a );
 a26233a <=( (not A265)  and  (not A236) );
 a26234a <=( (not A235)  and  a26233a );
 a26238a <=( (not A299)  and  (not A298) );
 a26239a <=( (not A266)  and  a26238a );
 a26240a <=( a26239a  and  a26234a );
 a26244a <=( (not A166)  and  (not A167) );
 a26245a <=( A170  and  a26244a );
 a26249a <=( (not A233)  and  A200 );
 a26250a <=( (not A199)  and  a26249a );
 a26251a <=( a26250a  and  a26245a );
 a26255a <=( A266  and  A265 );
 a26256a <=( (not A234)  and  a26255a );
 a26260a <=( (not A302)  and  (not A301) );
 a26261a <=( A298  and  a26260a );
 a26262a <=( a26261a  and  a26256a );
 a26266a <=( (not A166)  and  (not A167) );
 a26267a <=( A170  and  a26266a );
 a26271a <=( (not A233)  and  A200 );
 a26272a <=( (not A199)  and  a26271a );
 a26273a <=( a26272a  and  a26267a );
 a26277a <=( (not A268)  and  (not A266) );
 a26278a <=( (not A234)  and  a26277a );
 a26282a <=( (not A300)  and  A298 );
 a26283a <=( (not A269)  and  a26282a );
 a26284a <=( a26283a  and  a26278a );
 a26288a <=( (not A166)  and  (not A167) );
 a26289a <=( A170  and  a26288a );
 a26293a <=( (not A233)  and  A200 );
 a26294a <=( (not A199)  and  a26293a );
 a26295a <=( a26294a  and  a26289a );
 a26299a <=( (not A268)  and  (not A266) );
 a26300a <=( (not A234)  and  a26299a );
 a26304a <=( A299  and  A298 );
 a26305a <=( (not A269)  and  a26304a );
 a26306a <=( a26305a  and  a26300a );
 a26310a <=( (not A166)  and  (not A167) );
 a26311a <=( A170  and  a26310a );
 a26315a <=( (not A233)  and  A200 );
 a26316a <=( (not A199)  and  a26315a );
 a26317a <=( a26316a  and  a26311a );
 a26321a <=( (not A268)  and  (not A266) );
 a26322a <=( (not A234)  and  a26321a );
 a26326a <=( (not A299)  and  (not A298) );
 a26327a <=( (not A269)  and  a26326a );
 a26328a <=( a26327a  and  a26322a );
 a26332a <=( (not A166)  and  (not A167) );
 a26333a <=( A170  and  a26332a );
 a26337a <=( (not A233)  and  A200 );
 a26338a <=( (not A199)  and  a26337a );
 a26339a <=( a26338a  and  a26333a );
 a26343a <=( (not A267)  and  (not A266) );
 a26344a <=( (not A234)  and  a26343a );
 a26348a <=( (not A302)  and  (not A301) );
 a26349a <=( A298  and  a26348a );
 a26350a <=( a26349a  and  a26344a );
 a26354a <=( (not A166)  and  (not A167) );
 a26355a <=( A170  and  a26354a );
 a26359a <=( (not A233)  and  A200 );
 a26360a <=( (not A199)  and  a26359a );
 a26361a <=( a26360a  and  a26355a );
 a26365a <=( (not A266)  and  (not A265) );
 a26366a <=( (not A234)  and  a26365a );
 a26370a <=( (not A302)  and  (not A301) );
 a26371a <=( A298  and  a26370a );
 a26372a <=( a26371a  and  a26366a );
 a26376a <=( (not A166)  and  (not A167) );
 a26377a <=( A170  and  a26376a );
 a26381a <=( (not A232)  and  A200 );
 a26382a <=( (not A199)  and  a26381a );
 a26383a <=( a26382a  and  a26377a );
 a26387a <=( A266  and  A265 );
 a26388a <=( (not A233)  and  a26387a );
 a26392a <=( (not A302)  and  (not A301) );
 a26393a <=( A298  and  a26392a );
 a26394a <=( a26393a  and  a26388a );
 a26398a <=( (not A166)  and  (not A167) );
 a26399a <=( A170  and  a26398a );
 a26403a <=( (not A232)  and  A200 );
 a26404a <=( (not A199)  and  a26403a );
 a26405a <=( a26404a  and  a26399a );
 a26409a <=( (not A268)  and  (not A266) );
 a26410a <=( (not A233)  and  a26409a );
 a26414a <=( (not A300)  and  A298 );
 a26415a <=( (not A269)  and  a26414a );
 a26416a <=( a26415a  and  a26410a );
 a26420a <=( (not A166)  and  (not A167) );
 a26421a <=( A170  and  a26420a );
 a26425a <=( (not A232)  and  A200 );
 a26426a <=( (not A199)  and  a26425a );
 a26427a <=( a26426a  and  a26421a );
 a26431a <=( (not A268)  and  (not A266) );
 a26432a <=( (not A233)  and  a26431a );
 a26436a <=( A299  and  A298 );
 a26437a <=( (not A269)  and  a26436a );
 a26438a <=( a26437a  and  a26432a );
 a26442a <=( (not A166)  and  (not A167) );
 a26443a <=( A170  and  a26442a );
 a26447a <=( (not A232)  and  A200 );
 a26448a <=( (not A199)  and  a26447a );
 a26449a <=( a26448a  and  a26443a );
 a26453a <=( (not A268)  and  (not A266) );
 a26454a <=( (not A233)  and  a26453a );
 a26458a <=( (not A299)  and  (not A298) );
 a26459a <=( (not A269)  and  a26458a );
 a26460a <=( a26459a  and  a26454a );
 a26464a <=( (not A166)  and  (not A167) );
 a26465a <=( A170  and  a26464a );
 a26469a <=( (not A232)  and  A200 );
 a26470a <=( (not A199)  and  a26469a );
 a26471a <=( a26470a  and  a26465a );
 a26475a <=( (not A267)  and  (not A266) );
 a26476a <=( (not A233)  and  a26475a );
 a26480a <=( (not A302)  and  (not A301) );
 a26481a <=( A298  and  a26480a );
 a26482a <=( a26481a  and  a26476a );
 a26486a <=( (not A166)  and  (not A167) );
 a26487a <=( A170  and  a26486a );
 a26491a <=( (not A232)  and  A200 );
 a26492a <=( (not A199)  and  a26491a );
 a26493a <=( a26492a  and  a26487a );
 a26497a <=( (not A266)  and  (not A265) );
 a26498a <=( (not A233)  and  a26497a );
 a26502a <=( (not A302)  and  (not A301) );
 a26503a <=( A298  and  a26502a );
 a26504a <=( a26503a  and  a26498a );
 a26508a <=( A167  and  (not A168) );
 a26509a <=( A170  and  a26508a );
 a26513a <=( A200  and  (not A199) );
 a26514a <=( A166  and  a26513a );
 a26515a <=( a26514a  and  a26509a );
 a26519a <=( A265  and  A233 );
 a26520a <=( A232  and  a26519a );
 a26524a <=( (not A300)  and  (not A299) );
 a26525a <=( (not A267)  and  a26524a );
 a26526a <=( a26525a  and  a26520a );
 a26530a <=( A167  and  (not A168) );
 a26531a <=( A170  and  a26530a );
 a26535a <=( A200  and  (not A199) );
 a26536a <=( A166  and  a26535a );
 a26537a <=( a26536a  and  a26531a );
 a26541a <=( A265  and  A233 );
 a26542a <=( A232  and  a26541a );
 a26546a <=( A299  and  A298 );
 a26547a <=( (not A267)  and  a26546a );
 a26548a <=( a26547a  and  a26542a );
 a26552a <=( A167  and  (not A168) );
 a26553a <=( A170  and  a26552a );
 a26557a <=( A200  and  (not A199) );
 a26558a <=( A166  and  a26557a );
 a26559a <=( a26558a  and  a26553a );
 a26563a <=( A265  and  A233 );
 a26564a <=( A232  and  a26563a );
 a26568a <=( (not A299)  and  (not A298) );
 a26569a <=( (not A267)  and  a26568a );
 a26570a <=( a26569a  and  a26564a );
 a26574a <=( A167  and  (not A168) );
 a26575a <=( A170  and  a26574a );
 a26579a <=( A200  and  (not A199) );
 a26580a <=( A166  and  a26579a );
 a26581a <=( a26580a  and  a26575a );
 a26585a <=( A265  and  A233 );
 a26586a <=( A232  and  a26585a );
 a26590a <=( (not A300)  and  (not A299) );
 a26591a <=( A266  and  a26590a );
 a26592a <=( a26591a  and  a26586a );
 a26596a <=( A167  and  (not A168) );
 a26597a <=( A170  and  a26596a );
 a26601a <=( A200  and  (not A199) );
 a26602a <=( A166  and  a26601a );
 a26603a <=( a26602a  and  a26597a );
 a26607a <=( A265  and  A233 );
 a26608a <=( A232  and  a26607a );
 a26612a <=( A299  and  A298 );
 a26613a <=( A266  and  a26612a );
 a26614a <=( a26613a  and  a26608a );
 a26618a <=( A167  and  (not A168) );
 a26619a <=( A170  and  a26618a );
 a26623a <=( A200  and  (not A199) );
 a26624a <=( A166  and  a26623a );
 a26625a <=( a26624a  and  a26619a );
 a26629a <=( A265  and  A233 );
 a26630a <=( A232  and  a26629a );
 a26634a <=( (not A299)  and  (not A298) );
 a26635a <=( A266  and  a26634a );
 a26636a <=( a26635a  and  a26630a );
 a26640a <=( A167  and  (not A168) );
 a26641a <=( A170  and  a26640a );
 a26645a <=( A200  and  (not A199) );
 a26646a <=( A166  and  a26645a );
 a26647a <=( a26646a  and  a26641a );
 a26651a <=( (not A265)  and  A233 );
 a26652a <=( A232  and  a26651a );
 a26656a <=( (not A300)  and  (not A299) );
 a26657a <=( (not A266)  and  a26656a );
 a26658a <=( a26657a  and  a26652a );
 a26662a <=( A167  and  (not A168) );
 a26663a <=( A170  and  a26662a );
 a26667a <=( A200  and  (not A199) );
 a26668a <=( A166  and  a26667a );
 a26669a <=( a26668a  and  a26663a );
 a26673a <=( (not A265)  and  A233 );
 a26674a <=( A232  and  a26673a );
 a26678a <=( A299  and  A298 );
 a26679a <=( (not A266)  and  a26678a );
 a26680a <=( a26679a  and  a26674a );
 a26684a <=( A167  and  (not A168) );
 a26685a <=( A170  and  a26684a );
 a26689a <=( A200  and  (not A199) );
 a26690a <=( A166  and  a26689a );
 a26691a <=( a26690a  and  a26685a );
 a26695a <=( (not A265)  and  A233 );
 a26696a <=( A232  and  a26695a );
 a26700a <=( (not A299)  and  (not A298) );
 a26701a <=( (not A266)  and  a26700a );
 a26702a <=( a26701a  and  a26696a );
 a26706a <=( A167  and  (not A168) );
 a26707a <=( A170  and  a26706a );
 a26711a <=( A200  and  (not A199) );
 a26712a <=( A166  and  a26711a );
 a26713a <=( a26712a  and  a26707a );
 a26717a <=( A298  and  A233 );
 a26718a <=( (not A232)  and  a26717a );
 a26722a <=( A301  and  A300 );
 a26723a <=( (not A299)  and  a26722a );
 a26724a <=( a26723a  and  a26718a );
 a26728a <=( A167  and  (not A168) );
 a26729a <=( A170  and  a26728a );
 a26733a <=( A200  and  (not A199) );
 a26734a <=( A166  and  a26733a );
 a26735a <=( a26734a  and  a26729a );
 a26739a <=( A298  and  A233 );
 a26740a <=( (not A232)  and  a26739a );
 a26744a <=( A302  and  A300 );
 a26745a <=( (not A299)  and  a26744a );
 a26746a <=( a26745a  and  a26740a );
 a26750a <=( A167  and  (not A168) );
 a26751a <=( A170  and  a26750a );
 a26755a <=( A200  and  (not A199) );
 a26756a <=( A166  and  a26755a );
 a26757a <=( a26756a  and  a26751a );
 a26761a <=( A265  and  A233 );
 a26762a <=( (not A232)  and  a26761a );
 a26766a <=( A268  and  A267 );
 a26767a <=( (not A266)  and  a26766a );
 a26768a <=( a26767a  and  a26762a );
 a26772a <=( A167  and  (not A168) );
 a26773a <=( A170  and  a26772a );
 a26777a <=( A200  and  (not A199) );
 a26778a <=( A166  and  a26777a );
 a26779a <=( a26778a  and  a26773a );
 a26783a <=( A265  and  A233 );
 a26784a <=( (not A232)  and  a26783a );
 a26788a <=( A269  and  A267 );
 a26789a <=( (not A266)  and  a26788a );
 a26790a <=( a26789a  and  a26784a );
 a26794a <=( A167  and  (not A168) );
 a26795a <=( A170  and  a26794a );
 a26799a <=( A200  and  (not A199) );
 a26800a <=( A166  and  a26799a );
 a26801a <=( a26800a  and  a26795a );
 a26805a <=( A265  and  (not A234) );
 a26806a <=( (not A233)  and  a26805a );
 a26810a <=( (not A300)  and  A298 );
 a26811a <=( A266  and  a26810a );
 a26812a <=( a26811a  and  a26806a );
 a26816a <=( A167  and  (not A168) );
 a26817a <=( A170  and  a26816a );
 a26821a <=( A200  and  (not A199) );
 a26822a <=( A166  and  a26821a );
 a26823a <=( a26822a  and  a26817a );
 a26827a <=( A265  and  (not A234) );
 a26828a <=( (not A233)  and  a26827a );
 a26832a <=( A299  and  A298 );
 a26833a <=( A266  and  a26832a );
 a26834a <=( a26833a  and  a26828a );
 a26838a <=( A167  and  (not A168) );
 a26839a <=( A170  and  a26838a );
 a26843a <=( A200  and  (not A199) );
 a26844a <=( A166  and  a26843a );
 a26845a <=( a26844a  and  a26839a );
 a26849a <=( A265  and  (not A234) );
 a26850a <=( (not A233)  and  a26849a );
 a26854a <=( (not A299)  and  (not A298) );
 a26855a <=( A266  and  a26854a );
 a26856a <=( a26855a  and  a26850a );
 a26860a <=( A167  and  (not A168) );
 a26861a <=( A170  and  a26860a );
 a26865a <=( A200  and  (not A199) );
 a26866a <=( A166  and  a26865a );
 a26867a <=( a26866a  and  a26861a );
 a26871a <=( (not A266)  and  (not A234) );
 a26872a <=( (not A233)  and  a26871a );
 a26876a <=( (not A300)  and  A298 );
 a26877a <=( (not A267)  and  a26876a );
 a26878a <=( a26877a  and  a26872a );
 a26882a <=( A167  and  (not A168) );
 a26883a <=( A170  and  a26882a );
 a26887a <=( A200  and  (not A199) );
 a26888a <=( A166  and  a26887a );
 a26889a <=( a26888a  and  a26883a );
 a26893a <=( (not A266)  and  (not A234) );
 a26894a <=( (not A233)  and  a26893a );
 a26898a <=( A299  and  A298 );
 a26899a <=( (not A267)  and  a26898a );
 a26900a <=( a26899a  and  a26894a );
 a26904a <=( A167  and  (not A168) );
 a26905a <=( A170  and  a26904a );
 a26909a <=( A200  and  (not A199) );
 a26910a <=( A166  and  a26909a );
 a26911a <=( a26910a  and  a26905a );
 a26915a <=( (not A266)  and  (not A234) );
 a26916a <=( (not A233)  and  a26915a );
 a26920a <=( (not A299)  and  (not A298) );
 a26921a <=( (not A267)  and  a26920a );
 a26922a <=( a26921a  and  a26916a );
 a26926a <=( A167  and  (not A168) );
 a26927a <=( A170  and  a26926a );
 a26931a <=( A200  and  (not A199) );
 a26932a <=( A166  and  a26931a );
 a26933a <=( a26932a  and  a26927a );
 a26937a <=( (not A265)  and  (not A234) );
 a26938a <=( (not A233)  and  a26937a );
 a26942a <=( (not A300)  and  A298 );
 a26943a <=( (not A266)  and  a26942a );
 a26944a <=( a26943a  and  a26938a );
 a26948a <=( A167  and  (not A168) );
 a26949a <=( A170  and  a26948a );
 a26953a <=( A200  and  (not A199) );
 a26954a <=( A166  and  a26953a );
 a26955a <=( a26954a  and  a26949a );
 a26959a <=( (not A265)  and  (not A234) );
 a26960a <=( (not A233)  and  a26959a );
 a26964a <=( A299  and  A298 );
 a26965a <=( (not A266)  and  a26964a );
 a26966a <=( a26965a  and  a26960a );
 a26970a <=( A167  and  (not A168) );
 a26971a <=( A170  and  a26970a );
 a26975a <=( A200  and  (not A199) );
 a26976a <=( A166  and  a26975a );
 a26977a <=( a26976a  and  a26971a );
 a26981a <=( (not A265)  and  (not A234) );
 a26982a <=( (not A233)  and  a26981a );
 a26986a <=( (not A299)  and  (not A298) );
 a26987a <=( (not A266)  and  a26986a );
 a26988a <=( a26987a  and  a26982a );
 a26992a <=( A167  and  (not A168) );
 a26993a <=( A170  and  a26992a );
 a26997a <=( A200  and  (not A199) );
 a26998a <=( A166  and  a26997a );
 a26999a <=( a26998a  and  a26993a );
 a27003a <=( A234  and  (not A233) );
 a27004a <=( A232  and  a27003a );
 a27008a <=( A299  and  (not A298) );
 a27009a <=( A235  and  a27008a );
 a27010a <=( a27009a  and  a27004a );
 a27014a <=( A167  and  (not A168) );
 a27015a <=( A170  and  a27014a );
 a27019a <=( A200  and  (not A199) );
 a27020a <=( A166  and  a27019a );
 a27021a <=( a27020a  and  a27015a );
 a27025a <=( A234  and  (not A233) );
 a27026a <=( A232  and  a27025a );
 a27030a <=( A266  and  (not A265) );
 a27031a <=( A235  and  a27030a );
 a27032a <=( a27031a  and  a27026a );
 a27036a <=( A167  and  (not A168) );
 a27037a <=( A170  and  a27036a );
 a27041a <=( A200  and  (not A199) );
 a27042a <=( A166  and  a27041a );
 a27043a <=( a27042a  and  a27037a );
 a27047a <=( A234  and  (not A233) );
 a27048a <=( A232  and  a27047a );
 a27052a <=( A299  and  (not A298) );
 a27053a <=( A236  and  a27052a );
 a27054a <=( a27053a  and  a27048a );
 a27058a <=( A167  and  (not A168) );
 a27059a <=( A170  and  a27058a );
 a27063a <=( A200  and  (not A199) );
 a27064a <=( A166  and  a27063a );
 a27065a <=( a27064a  and  a27059a );
 a27069a <=( A234  and  (not A233) );
 a27070a <=( A232  and  a27069a );
 a27074a <=( A266  and  (not A265) );
 a27075a <=( A236  and  a27074a );
 a27076a <=( a27075a  and  a27070a );
 a27080a <=( A167  and  (not A168) );
 a27081a <=( A170  and  a27080a );
 a27085a <=( A200  and  (not A199) );
 a27086a <=( A166  and  a27085a );
 a27087a <=( a27086a  and  a27081a );
 a27091a <=( A265  and  (not A233) );
 a27092a <=( (not A232)  and  a27091a );
 a27096a <=( (not A300)  and  A298 );
 a27097a <=( A266  and  a27096a );
 a27098a <=( a27097a  and  a27092a );
 a27102a <=( A167  and  (not A168) );
 a27103a <=( A170  and  a27102a );
 a27107a <=( A200  and  (not A199) );
 a27108a <=( A166  and  a27107a );
 a27109a <=( a27108a  and  a27103a );
 a27113a <=( A265  and  (not A233) );
 a27114a <=( (not A232)  and  a27113a );
 a27118a <=( A299  and  A298 );
 a27119a <=( A266  and  a27118a );
 a27120a <=( a27119a  and  a27114a );
 a27124a <=( A167  and  (not A168) );
 a27125a <=( A170  and  a27124a );
 a27129a <=( A200  and  (not A199) );
 a27130a <=( A166  and  a27129a );
 a27131a <=( a27130a  and  a27125a );
 a27135a <=( A265  and  (not A233) );
 a27136a <=( (not A232)  and  a27135a );
 a27140a <=( (not A299)  and  (not A298) );
 a27141a <=( A266  and  a27140a );
 a27142a <=( a27141a  and  a27136a );
 a27146a <=( A167  and  (not A168) );
 a27147a <=( A170  and  a27146a );
 a27151a <=( A200  and  (not A199) );
 a27152a <=( A166  and  a27151a );
 a27153a <=( a27152a  and  a27147a );
 a27157a <=( (not A266)  and  (not A233) );
 a27158a <=( (not A232)  and  a27157a );
 a27162a <=( (not A300)  and  A298 );
 a27163a <=( (not A267)  and  a27162a );
 a27164a <=( a27163a  and  a27158a );
 a27168a <=( A167  and  (not A168) );
 a27169a <=( A170  and  a27168a );
 a27173a <=( A200  and  (not A199) );
 a27174a <=( A166  and  a27173a );
 a27175a <=( a27174a  and  a27169a );
 a27179a <=( (not A266)  and  (not A233) );
 a27180a <=( (not A232)  and  a27179a );
 a27184a <=( A299  and  A298 );
 a27185a <=( (not A267)  and  a27184a );
 a27186a <=( a27185a  and  a27180a );
 a27190a <=( A167  and  (not A168) );
 a27191a <=( A170  and  a27190a );
 a27195a <=( A200  and  (not A199) );
 a27196a <=( A166  and  a27195a );
 a27197a <=( a27196a  and  a27191a );
 a27201a <=( (not A266)  and  (not A233) );
 a27202a <=( (not A232)  and  a27201a );
 a27206a <=( (not A299)  and  (not A298) );
 a27207a <=( (not A267)  and  a27206a );
 a27208a <=( a27207a  and  a27202a );
 a27212a <=( A167  and  (not A168) );
 a27213a <=( A170  and  a27212a );
 a27217a <=( A200  and  (not A199) );
 a27218a <=( A166  and  a27217a );
 a27219a <=( a27218a  and  a27213a );
 a27223a <=( (not A265)  and  (not A233) );
 a27224a <=( (not A232)  and  a27223a );
 a27228a <=( (not A300)  and  A298 );
 a27229a <=( (not A266)  and  a27228a );
 a27230a <=( a27229a  and  a27224a );
 a27234a <=( A167  and  (not A168) );
 a27235a <=( A170  and  a27234a );
 a27239a <=( A200  and  (not A199) );
 a27240a <=( A166  and  a27239a );
 a27241a <=( a27240a  and  a27235a );
 a27245a <=( (not A265)  and  (not A233) );
 a27246a <=( (not A232)  and  a27245a );
 a27250a <=( A299  and  A298 );
 a27251a <=( (not A266)  and  a27250a );
 a27252a <=( a27251a  and  a27246a );
 a27256a <=( A167  and  (not A168) );
 a27257a <=( A170  and  a27256a );
 a27261a <=( A200  and  (not A199) );
 a27262a <=( A166  and  a27261a );
 a27263a <=( a27262a  and  a27257a );
 a27267a <=( (not A265)  and  (not A233) );
 a27268a <=( (not A232)  and  a27267a );
 a27272a <=( (not A299)  and  (not A298) );
 a27273a <=( (not A266)  and  a27272a );
 a27274a <=( a27273a  and  a27268a );
 a27278a <=( A167  and  (not A168) );
 a27279a <=( (not A170)  and  a27278a );
 a27283a <=( A200  and  (not A199) );
 a27284a <=( (not A166)  and  a27283a );
 a27285a <=( a27284a  and  a27279a );
 a27289a <=( A265  and  A233 );
 a27290a <=( A232  and  a27289a );
 a27294a <=( (not A300)  and  (not A299) );
 a27295a <=( (not A267)  and  a27294a );
 a27296a <=( a27295a  and  a27290a );
 a27300a <=( A167  and  (not A168) );
 a27301a <=( (not A170)  and  a27300a );
 a27305a <=( A200  and  (not A199) );
 a27306a <=( (not A166)  and  a27305a );
 a27307a <=( a27306a  and  a27301a );
 a27311a <=( A265  and  A233 );
 a27312a <=( A232  and  a27311a );
 a27316a <=( A299  and  A298 );
 a27317a <=( (not A267)  and  a27316a );
 a27318a <=( a27317a  and  a27312a );
 a27322a <=( A167  and  (not A168) );
 a27323a <=( (not A170)  and  a27322a );
 a27327a <=( A200  and  (not A199) );
 a27328a <=( (not A166)  and  a27327a );
 a27329a <=( a27328a  and  a27323a );
 a27333a <=( A265  and  A233 );
 a27334a <=( A232  and  a27333a );
 a27338a <=( (not A299)  and  (not A298) );
 a27339a <=( (not A267)  and  a27338a );
 a27340a <=( a27339a  and  a27334a );
 a27344a <=( A167  and  (not A168) );
 a27345a <=( (not A170)  and  a27344a );
 a27349a <=( A200  and  (not A199) );
 a27350a <=( (not A166)  and  a27349a );
 a27351a <=( a27350a  and  a27345a );
 a27355a <=( A265  and  A233 );
 a27356a <=( A232  and  a27355a );
 a27360a <=( (not A300)  and  (not A299) );
 a27361a <=( A266  and  a27360a );
 a27362a <=( a27361a  and  a27356a );
 a27366a <=( A167  and  (not A168) );
 a27367a <=( (not A170)  and  a27366a );
 a27371a <=( A200  and  (not A199) );
 a27372a <=( (not A166)  and  a27371a );
 a27373a <=( a27372a  and  a27367a );
 a27377a <=( A265  and  A233 );
 a27378a <=( A232  and  a27377a );
 a27382a <=( A299  and  A298 );
 a27383a <=( A266  and  a27382a );
 a27384a <=( a27383a  and  a27378a );
 a27388a <=( A167  and  (not A168) );
 a27389a <=( (not A170)  and  a27388a );
 a27393a <=( A200  and  (not A199) );
 a27394a <=( (not A166)  and  a27393a );
 a27395a <=( a27394a  and  a27389a );
 a27399a <=( A265  and  A233 );
 a27400a <=( A232  and  a27399a );
 a27404a <=( (not A299)  and  (not A298) );
 a27405a <=( A266  and  a27404a );
 a27406a <=( a27405a  and  a27400a );
 a27410a <=( A167  and  (not A168) );
 a27411a <=( (not A170)  and  a27410a );
 a27415a <=( A200  and  (not A199) );
 a27416a <=( (not A166)  and  a27415a );
 a27417a <=( a27416a  and  a27411a );
 a27421a <=( (not A265)  and  A233 );
 a27422a <=( A232  and  a27421a );
 a27426a <=( (not A300)  and  (not A299) );
 a27427a <=( (not A266)  and  a27426a );
 a27428a <=( a27427a  and  a27422a );
 a27432a <=( A167  and  (not A168) );
 a27433a <=( (not A170)  and  a27432a );
 a27437a <=( A200  and  (not A199) );
 a27438a <=( (not A166)  and  a27437a );
 a27439a <=( a27438a  and  a27433a );
 a27443a <=( (not A265)  and  A233 );
 a27444a <=( A232  and  a27443a );
 a27448a <=( A299  and  A298 );
 a27449a <=( (not A266)  and  a27448a );
 a27450a <=( a27449a  and  a27444a );
 a27454a <=( A167  and  (not A168) );
 a27455a <=( (not A170)  and  a27454a );
 a27459a <=( A200  and  (not A199) );
 a27460a <=( (not A166)  and  a27459a );
 a27461a <=( a27460a  and  a27455a );
 a27465a <=( (not A265)  and  A233 );
 a27466a <=( A232  and  a27465a );
 a27470a <=( (not A299)  and  (not A298) );
 a27471a <=( (not A266)  and  a27470a );
 a27472a <=( a27471a  and  a27466a );
 a27476a <=( A167  and  (not A168) );
 a27477a <=( (not A170)  and  a27476a );
 a27481a <=( A200  and  (not A199) );
 a27482a <=( (not A166)  and  a27481a );
 a27483a <=( a27482a  and  a27477a );
 a27487a <=( A298  and  A233 );
 a27488a <=( (not A232)  and  a27487a );
 a27492a <=( A301  and  A300 );
 a27493a <=( (not A299)  and  a27492a );
 a27494a <=( a27493a  and  a27488a );
 a27498a <=( A167  and  (not A168) );
 a27499a <=( (not A170)  and  a27498a );
 a27503a <=( A200  and  (not A199) );
 a27504a <=( (not A166)  and  a27503a );
 a27505a <=( a27504a  and  a27499a );
 a27509a <=( A298  and  A233 );
 a27510a <=( (not A232)  and  a27509a );
 a27514a <=( A302  and  A300 );
 a27515a <=( (not A299)  and  a27514a );
 a27516a <=( a27515a  and  a27510a );
 a27520a <=( A167  and  (not A168) );
 a27521a <=( (not A170)  and  a27520a );
 a27525a <=( A200  and  (not A199) );
 a27526a <=( (not A166)  and  a27525a );
 a27527a <=( a27526a  and  a27521a );
 a27531a <=( A265  and  A233 );
 a27532a <=( (not A232)  and  a27531a );
 a27536a <=( A268  and  A267 );
 a27537a <=( (not A266)  and  a27536a );
 a27538a <=( a27537a  and  a27532a );
 a27542a <=( A167  and  (not A168) );
 a27543a <=( (not A170)  and  a27542a );
 a27547a <=( A200  and  (not A199) );
 a27548a <=( (not A166)  and  a27547a );
 a27549a <=( a27548a  and  a27543a );
 a27553a <=( A265  and  A233 );
 a27554a <=( (not A232)  and  a27553a );
 a27558a <=( A269  and  A267 );
 a27559a <=( (not A266)  and  a27558a );
 a27560a <=( a27559a  and  a27554a );
 a27564a <=( A167  and  (not A168) );
 a27565a <=( (not A170)  and  a27564a );
 a27569a <=( A200  and  (not A199) );
 a27570a <=( (not A166)  and  a27569a );
 a27571a <=( a27570a  and  a27565a );
 a27575a <=( A265  and  (not A234) );
 a27576a <=( (not A233)  and  a27575a );
 a27580a <=( (not A300)  and  A298 );
 a27581a <=( A266  and  a27580a );
 a27582a <=( a27581a  and  a27576a );
 a27586a <=( A167  and  (not A168) );
 a27587a <=( (not A170)  and  a27586a );
 a27591a <=( A200  and  (not A199) );
 a27592a <=( (not A166)  and  a27591a );
 a27593a <=( a27592a  and  a27587a );
 a27597a <=( A265  and  (not A234) );
 a27598a <=( (not A233)  and  a27597a );
 a27602a <=( A299  and  A298 );
 a27603a <=( A266  and  a27602a );
 a27604a <=( a27603a  and  a27598a );
 a27608a <=( A167  and  (not A168) );
 a27609a <=( (not A170)  and  a27608a );
 a27613a <=( A200  and  (not A199) );
 a27614a <=( (not A166)  and  a27613a );
 a27615a <=( a27614a  and  a27609a );
 a27619a <=( A265  and  (not A234) );
 a27620a <=( (not A233)  and  a27619a );
 a27624a <=( (not A299)  and  (not A298) );
 a27625a <=( A266  and  a27624a );
 a27626a <=( a27625a  and  a27620a );
 a27630a <=( A167  and  (not A168) );
 a27631a <=( (not A170)  and  a27630a );
 a27635a <=( A200  and  (not A199) );
 a27636a <=( (not A166)  and  a27635a );
 a27637a <=( a27636a  and  a27631a );
 a27641a <=( (not A266)  and  (not A234) );
 a27642a <=( (not A233)  and  a27641a );
 a27646a <=( (not A300)  and  A298 );
 a27647a <=( (not A267)  and  a27646a );
 a27648a <=( a27647a  and  a27642a );
 a27652a <=( A167  and  (not A168) );
 a27653a <=( (not A170)  and  a27652a );
 a27657a <=( A200  and  (not A199) );
 a27658a <=( (not A166)  and  a27657a );
 a27659a <=( a27658a  and  a27653a );
 a27663a <=( (not A266)  and  (not A234) );
 a27664a <=( (not A233)  and  a27663a );
 a27668a <=( A299  and  A298 );
 a27669a <=( (not A267)  and  a27668a );
 a27670a <=( a27669a  and  a27664a );
 a27674a <=( A167  and  (not A168) );
 a27675a <=( (not A170)  and  a27674a );
 a27679a <=( A200  and  (not A199) );
 a27680a <=( (not A166)  and  a27679a );
 a27681a <=( a27680a  and  a27675a );
 a27685a <=( (not A266)  and  (not A234) );
 a27686a <=( (not A233)  and  a27685a );
 a27690a <=( (not A299)  and  (not A298) );
 a27691a <=( (not A267)  and  a27690a );
 a27692a <=( a27691a  and  a27686a );
 a27696a <=( A167  and  (not A168) );
 a27697a <=( (not A170)  and  a27696a );
 a27701a <=( A200  and  (not A199) );
 a27702a <=( (not A166)  and  a27701a );
 a27703a <=( a27702a  and  a27697a );
 a27707a <=( (not A265)  and  (not A234) );
 a27708a <=( (not A233)  and  a27707a );
 a27712a <=( (not A300)  and  A298 );
 a27713a <=( (not A266)  and  a27712a );
 a27714a <=( a27713a  and  a27708a );
 a27718a <=( A167  and  (not A168) );
 a27719a <=( (not A170)  and  a27718a );
 a27723a <=( A200  and  (not A199) );
 a27724a <=( (not A166)  and  a27723a );
 a27725a <=( a27724a  and  a27719a );
 a27729a <=( (not A265)  and  (not A234) );
 a27730a <=( (not A233)  and  a27729a );
 a27734a <=( A299  and  A298 );
 a27735a <=( (not A266)  and  a27734a );
 a27736a <=( a27735a  and  a27730a );
 a27740a <=( A167  and  (not A168) );
 a27741a <=( (not A170)  and  a27740a );
 a27745a <=( A200  and  (not A199) );
 a27746a <=( (not A166)  and  a27745a );
 a27747a <=( a27746a  and  a27741a );
 a27751a <=( (not A265)  and  (not A234) );
 a27752a <=( (not A233)  and  a27751a );
 a27756a <=( (not A299)  and  (not A298) );
 a27757a <=( (not A266)  and  a27756a );
 a27758a <=( a27757a  and  a27752a );
 a27762a <=( A167  and  (not A168) );
 a27763a <=( (not A170)  and  a27762a );
 a27767a <=( A200  and  (not A199) );
 a27768a <=( (not A166)  and  a27767a );
 a27769a <=( a27768a  and  a27763a );
 a27773a <=( A234  and  (not A233) );
 a27774a <=( A232  and  a27773a );
 a27778a <=( A299  and  (not A298) );
 a27779a <=( A235  and  a27778a );
 a27780a <=( a27779a  and  a27774a );
 a27784a <=( A167  and  (not A168) );
 a27785a <=( (not A170)  and  a27784a );
 a27789a <=( A200  and  (not A199) );
 a27790a <=( (not A166)  and  a27789a );
 a27791a <=( a27790a  and  a27785a );
 a27795a <=( A234  and  (not A233) );
 a27796a <=( A232  and  a27795a );
 a27800a <=( A266  and  (not A265) );
 a27801a <=( A235  and  a27800a );
 a27802a <=( a27801a  and  a27796a );
 a27806a <=( A167  and  (not A168) );
 a27807a <=( (not A170)  and  a27806a );
 a27811a <=( A200  and  (not A199) );
 a27812a <=( (not A166)  and  a27811a );
 a27813a <=( a27812a  and  a27807a );
 a27817a <=( A234  and  (not A233) );
 a27818a <=( A232  and  a27817a );
 a27822a <=( A299  and  (not A298) );
 a27823a <=( A236  and  a27822a );
 a27824a <=( a27823a  and  a27818a );
 a27828a <=( A167  and  (not A168) );
 a27829a <=( (not A170)  and  a27828a );
 a27833a <=( A200  and  (not A199) );
 a27834a <=( (not A166)  and  a27833a );
 a27835a <=( a27834a  and  a27829a );
 a27839a <=( A234  and  (not A233) );
 a27840a <=( A232  and  a27839a );
 a27844a <=( A266  and  (not A265) );
 a27845a <=( A236  and  a27844a );
 a27846a <=( a27845a  and  a27840a );
 a27850a <=( A167  and  (not A168) );
 a27851a <=( (not A170)  and  a27850a );
 a27855a <=( A200  and  (not A199) );
 a27856a <=( (not A166)  and  a27855a );
 a27857a <=( a27856a  and  a27851a );
 a27861a <=( A265  and  (not A233) );
 a27862a <=( (not A232)  and  a27861a );
 a27866a <=( (not A300)  and  A298 );
 a27867a <=( A266  and  a27866a );
 a27868a <=( a27867a  and  a27862a );
 a27872a <=( A167  and  (not A168) );
 a27873a <=( (not A170)  and  a27872a );
 a27877a <=( A200  and  (not A199) );
 a27878a <=( (not A166)  and  a27877a );
 a27879a <=( a27878a  and  a27873a );
 a27883a <=( A265  and  (not A233) );
 a27884a <=( (not A232)  and  a27883a );
 a27888a <=( A299  and  A298 );
 a27889a <=( A266  and  a27888a );
 a27890a <=( a27889a  and  a27884a );
 a27894a <=( A167  and  (not A168) );
 a27895a <=( (not A170)  and  a27894a );
 a27899a <=( A200  and  (not A199) );
 a27900a <=( (not A166)  and  a27899a );
 a27901a <=( a27900a  and  a27895a );
 a27905a <=( A265  and  (not A233) );
 a27906a <=( (not A232)  and  a27905a );
 a27910a <=( (not A299)  and  (not A298) );
 a27911a <=( A266  and  a27910a );
 a27912a <=( a27911a  and  a27906a );
 a27916a <=( A167  and  (not A168) );
 a27917a <=( (not A170)  and  a27916a );
 a27921a <=( A200  and  (not A199) );
 a27922a <=( (not A166)  and  a27921a );
 a27923a <=( a27922a  and  a27917a );
 a27927a <=( (not A266)  and  (not A233) );
 a27928a <=( (not A232)  and  a27927a );
 a27932a <=( (not A300)  and  A298 );
 a27933a <=( (not A267)  and  a27932a );
 a27934a <=( a27933a  and  a27928a );
 a27938a <=( A167  and  (not A168) );
 a27939a <=( (not A170)  and  a27938a );
 a27943a <=( A200  and  (not A199) );
 a27944a <=( (not A166)  and  a27943a );
 a27945a <=( a27944a  and  a27939a );
 a27949a <=( (not A266)  and  (not A233) );
 a27950a <=( (not A232)  and  a27949a );
 a27954a <=( A299  and  A298 );
 a27955a <=( (not A267)  and  a27954a );
 a27956a <=( a27955a  and  a27950a );
 a27960a <=( A167  and  (not A168) );
 a27961a <=( (not A170)  and  a27960a );
 a27965a <=( A200  and  (not A199) );
 a27966a <=( (not A166)  and  a27965a );
 a27967a <=( a27966a  and  a27961a );
 a27971a <=( (not A266)  and  (not A233) );
 a27972a <=( (not A232)  and  a27971a );
 a27976a <=( (not A299)  and  (not A298) );
 a27977a <=( (not A267)  and  a27976a );
 a27978a <=( a27977a  and  a27972a );
 a27982a <=( A167  and  (not A168) );
 a27983a <=( (not A170)  and  a27982a );
 a27987a <=( A200  and  (not A199) );
 a27988a <=( (not A166)  and  a27987a );
 a27989a <=( a27988a  and  a27983a );
 a27993a <=( (not A265)  and  (not A233) );
 a27994a <=( (not A232)  and  a27993a );
 a27998a <=( (not A300)  and  A298 );
 a27999a <=( (not A266)  and  a27998a );
 a28000a <=( a27999a  and  a27994a );
 a28004a <=( A167  and  (not A168) );
 a28005a <=( (not A170)  and  a28004a );
 a28009a <=( A200  and  (not A199) );
 a28010a <=( (not A166)  and  a28009a );
 a28011a <=( a28010a  and  a28005a );
 a28015a <=( (not A265)  and  (not A233) );
 a28016a <=( (not A232)  and  a28015a );
 a28020a <=( A299  and  A298 );
 a28021a <=( (not A266)  and  a28020a );
 a28022a <=( a28021a  and  a28016a );
 a28026a <=( A167  and  (not A168) );
 a28027a <=( (not A170)  and  a28026a );
 a28031a <=( A200  and  (not A199) );
 a28032a <=( (not A166)  and  a28031a );
 a28033a <=( a28032a  and  a28027a );
 a28037a <=( (not A265)  and  (not A233) );
 a28038a <=( (not A232)  and  a28037a );
 a28042a <=( (not A299)  and  (not A298) );
 a28043a <=( (not A266)  and  a28042a );
 a28044a <=( a28043a  and  a28038a );
 a28048a <=( (not A167)  and  (not A168) );
 a28049a <=( (not A170)  and  a28048a );
 a28053a <=( A200  and  (not A199) );
 a28054a <=( A166  and  a28053a );
 a28055a <=( a28054a  and  a28049a );
 a28059a <=( A265  and  A233 );
 a28060a <=( A232  and  a28059a );
 a28064a <=( (not A300)  and  (not A299) );
 a28065a <=( (not A267)  and  a28064a );
 a28066a <=( a28065a  and  a28060a );
 a28070a <=( (not A167)  and  (not A168) );
 a28071a <=( (not A170)  and  a28070a );
 a28075a <=( A200  and  (not A199) );
 a28076a <=( A166  and  a28075a );
 a28077a <=( a28076a  and  a28071a );
 a28081a <=( A265  and  A233 );
 a28082a <=( A232  and  a28081a );
 a28086a <=( A299  and  A298 );
 a28087a <=( (not A267)  and  a28086a );
 a28088a <=( a28087a  and  a28082a );
 a28092a <=( (not A167)  and  (not A168) );
 a28093a <=( (not A170)  and  a28092a );
 a28097a <=( A200  and  (not A199) );
 a28098a <=( A166  and  a28097a );
 a28099a <=( a28098a  and  a28093a );
 a28103a <=( A265  and  A233 );
 a28104a <=( A232  and  a28103a );
 a28108a <=( (not A299)  and  (not A298) );
 a28109a <=( (not A267)  and  a28108a );
 a28110a <=( a28109a  and  a28104a );
 a28114a <=( (not A167)  and  (not A168) );
 a28115a <=( (not A170)  and  a28114a );
 a28119a <=( A200  and  (not A199) );
 a28120a <=( A166  and  a28119a );
 a28121a <=( a28120a  and  a28115a );
 a28125a <=( A265  and  A233 );
 a28126a <=( A232  and  a28125a );
 a28130a <=( (not A300)  and  (not A299) );
 a28131a <=( A266  and  a28130a );
 a28132a <=( a28131a  and  a28126a );
 a28136a <=( (not A167)  and  (not A168) );
 a28137a <=( (not A170)  and  a28136a );
 a28141a <=( A200  and  (not A199) );
 a28142a <=( A166  and  a28141a );
 a28143a <=( a28142a  and  a28137a );
 a28147a <=( A265  and  A233 );
 a28148a <=( A232  and  a28147a );
 a28152a <=( A299  and  A298 );
 a28153a <=( A266  and  a28152a );
 a28154a <=( a28153a  and  a28148a );
 a28158a <=( (not A167)  and  (not A168) );
 a28159a <=( (not A170)  and  a28158a );
 a28163a <=( A200  and  (not A199) );
 a28164a <=( A166  and  a28163a );
 a28165a <=( a28164a  and  a28159a );
 a28169a <=( A265  and  A233 );
 a28170a <=( A232  and  a28169a );
 a28174a <=( (not A299)  and  (not A298) );
 a28175a <=( A266  and  a28174a );
 a28176a <=( a28175a  and  a28170a );
 a28180a <=( (not A167)  and  (not A168) );
 a28181a <=( (not A170)  and  a28180a );
 a28185a <=( A200  and  (not A199) );
 a28186a <=( A166  and  a28185a );
 a28187a <=( a28186a  and  a28181a );
 a28191a <=( (not A265)  and  A233 );
 a28192a <=( A232  and  a28191a );
 a28196a <=( (not A300)  and  (not A299) );
 a28197a <=( (not A266)  and  a28196a );
 a28198a <=( a28197a  and  a28192a );
 a28202a <=( (not A167)  and  (not A168) );
 a28203a <=( (not A170)  and  a28202a );
 a28207a <=( A200  and  (not A199) );
 a28208a <=( A166  and  a28207a );
 a28209a <=( a28208a  and  a28203a );
 a28213a <=( (not A265)  and  A233 );
 a28214a <=( A232  and  a28213a );
 a28218a <=( A299  and  A298 );
 a28219a <=( (not A266)  and  a28218a );
 a28220a <=( a28219a  and  a28214a );
 a28224a <=( (not A167)  and  (not A168) );
 a28225a <=( (not A170)  and  a28224a );
 a28229a <=( A200  and  (not A199) );
 a28230a <=( A166  and  a28229a );
 a28231a <=( a28230a  and  a28225a );
 a28235a <=( (not A265)  and  A233 );
 a28236a <=( A232  and  a28235a );
 a28240a <=( (not A299)  and  (not A298) );
 a28241a <=( (not A266)  and  a28240a );
 a28242a <=( a28241a  and  a28236a );
 a28246a <=( (not A167)  and  (not A168) );
 a28247a <=( (not A170)  and  a28246a );
 a28251a <=( A200  and  (not A199) );
 a28252a <=( A166  and  a28251a );
 a28253a <=( a28252a  and  a28247a );
 a28257a <=( A298  and  A233 );
 a28258a <=( (not A232)  and  a28257a );
 a28262a <=( A301  and  A300 );
 a28263a <=( (not A299)  and  a28262a );
 a28264a <=( a28263a  and  a28258a );
 a28268a <=( (not A167)  and  (not A168) );
 a28269a <=( (not A170)  and  a28268a );
 a28273a <=( A200  and  (not A199) );
 a28274a <=( A166  and  a28273a );
 a28275a <=( a28274a  and  a28269a );
 a28279a <=( A298  and  A233 );
 a28280a <=( (not A232)  and  a28279a );
 a28284a <=( A302  and  A300 );
 a28285a <=( (not A299)  and  a28284a );
 a28286a <=( a28285a  and  a28280a );
 a28290a <=( (not A167)  and  (not A168) );
 a28291a <=( (not A170)  and  a28290a );
 a28295a <=( A200  and  (not A199) );
 a28296a <=( A166  and  a28295a );
 a28297a <=( a28296a  and  a28291a );
 a28301a <=( A265  and  A233 );
 a28302a <=( (not A232)  and  a28301a );
 a28306a <=( A268  and  A267 );
 a28307a <=( (not A266)  and  a28306a );
 a28308a <=( a28307a  and  a28302a );
 a28312a <=( (not A167)  and  (not A168) );
 a28313a <=( (not A170)  and  a28312a );
 a28317a <=( A200  and  (not A199) );
 a28318a <=( A166  and  a28317a );
 a28319a <=( a28318a  and  a28313a );
 a28323a <=( A265  and  A233 );
 a28324a <=( (not A232)  and  a28323a );
 a28328a <=( A269  and  A267 );
 a28329a <=( (not A266)  and  a28328a );
 a28330a <=( a28329a  and  a28324a );
 a28334a <=( (not A167)  and  (not A168) );
 a28335a <=( (not A170)  and  a28334a );
 a28339a <=( A200  and  (not A199) );
 a28340a <=( A166  and  a28339a );
 a28341a <=( a28340a  and  a28335a );
 a28345a <=( A265  and  (not A234) );
 a28346a <=( (not A233)  and  a28345a );
 a28350a <=( (not A300)  and  A298 );
 a28351a <=( A266  and  a28350a );
 a28352a <=( a28351a  and  a28346a );
 a28356a <=( (not A167)  and  (not A168) );
 a28357a <=( (not A170)  and  a28356a );
 a28361a <=( A200  and  (not A199) );
 a28362a <=( A166  and  a28361a );
 a28363a <=( a28362a  and  a28357a );
 a28367a <=( A265  and  (not A234) );
 a28368a <=( (not A233)  and  a28367a );
 a28372a <=( A299  and  A298 );
 a28373a <=( A266  and  a28372a );
 a28374a <=( a28373a  and  a28368a );
 a28378a <=( (not A167)  and  (not A168) );
 a28379a <=( (not A170)  and  a28378a );
 a28383a <=( A200  and  (not A199) );
 a28384a <=( A166  and  a28383a );
 a28385a <=( a28384a  and  a28379a );
 a28389a <=( A265  and  (not A234) );
 a28390a <=( (not A233)  and  a28389a );
 a28394a <=( (not A299)  and  (not A298) );
 a28395a <=( A266  and  a28394a );
 a28396a <=( a28395a  and  a28390a );
 a28400a <=( (not A167)  and  (not A168) );
 a28401a <=( (not A170)  and  a28400a );
 a28405a <=( A200  and  (not A199) );
 a28406a <=( A166  and  a28405a );
 a28407a <=( a28406a  and  a28401a );
 a28411a <=( (not A266)  and  (not A234) );
 a28412a <=( (not A233)  and  a28411a );
 a28416a <=( (not A300)  and  A298 );
 a28417a <=( (not A267)  and  a28416a );
 a28418a <=( a28417a  and  a28412a );
 a28422a <=( (not A167)  and  (not A168) );
 a28423a <=( (not A170)  and  a28422a );
 a28427a <=( A200  and  (not A199) );
 a28428a <=( A166  and  a28427a );
 a28429a <=( a28428a  and  a28423a );
 a28433a <=( (not A266)  and  (not A234) );
 a28434a <=( (not A233)  and  a28433a );
 a28438a <=( A299  and  A298 );
 a28439a <=( (not A267)  and  a28438a );
 a28440a <=( a28439a  and  a28434a );
 a28444a <=( (not A167)  and  (not A168) );
 a28445a <=( (not A170)  and  a28444a );
 a28449a <=( A200  and  (not A199) );
 a28450a <=( A166  and  a28449a );
 a28451a <=( a28450a  and  a28445a );
 a28455a <=( (not A266)  and  (not A234) );
 a28456a <=( (not A233)  and  a28455a );
 a28460a <=( (not A299)  and  (not A298) );
 a28461a <=( (not A267)  and  a28460a );
 a28462a <=( a28461a  and  a28456a );
 a28466a <=( (not A167)  and  (not A168) );
 a28467a <=( (not A170)  and  a28466a );
 a28471a <=( A200  and  (not A199) );
 a28472a <=( A166  and  a28471a );
 a28473a <=( a28472a  and  a28467a );
 a28477a <=( (not A265)  and  (not A234) );
 a28478a <=( (not A233)  and  a28477a );
 a28482a <=( (not A300)  and  A298 );
 a28483a <=( (not A266)  and  a28482a );
 a28484a <=( a28483a  and  a28478a );
 a28488a <=( (not A167)  and  (not A168) );
 a28489a <=( (not A170)  and  a28488a );
 a28493a <=( A200  and  (not A199) );
 a28494a <=( A166  and  a28493a );
 a28495a <=( a28494a  and  a28489a );
 a28499a <=( (not A265)  and  (not A234) );
 a28500a <=( (not A233)  and  a28499a );
 a28504a <=( A299  and  A298 );
 a28505a <=( (not A266)  and  a28504a );
 a28506a <=( a28505a  and  a28500a );
 a28510a <=( (not A167)  and  (not A168) );
 a28511a <=( (not A170)  and  a28510a );
 a28515a <=( A200  and  (not A199) );
 a28516a <=( A166  and  a28515a );
 a28517a <=( a28516a  and  a28511a );
 a28521a <=( (not A265)  and  (not A234) );
 a28522a <=( (not A233)  and  a28521a );
 a28526a <=( (not A299)  and  (not A298) );
 a28527a <=( (not A266)  and  a28526a );
 a28528a <=( a28527a  and  a28522a );
 a28532a <=( (not A167)  and  (not A168) );
 a28533a <=( (not A170)  and  a28532a );
 a28537a <=( A200  and  (not A199) );
 a28538a <=( A166  and  a28537a );
 a28539a <=( a28538a  and  a28533a );
 a28543a <=( A234  and  (not A233) );
 a28544a <=( A232  and  a28543a );
 a28548a <=( A299  and  (not A298) );
 a28549a <=( A235  and  a28548a );
 a28550a <=( a28549a  and  a28544a );
 a28554a <=( (not A167)  and  (not A168) );
 a28555a <=( (not A170)  and  a28554a );
 a28559a <=( A200  and  (not A199) );
 a28560a <=( A166  and  a28559a );
 a28561a <=( a28560a  and  a28555a );
 a28565a <=( A234  and  (not A233) );
 a28566a <=( A232  and  a28565a );
 a28570a <=( A266  and  (not A265) );
 a28571a <=( A235  and  a28570a );
 a28572a <=( a28571a  and  a28566a );
 a28576a <=( (not A167)  and  (not A168) );
 a28577a <=( (not A170)  and  a28576a );
 a28581a <=( A200  and  (not A199) );
 a28582a <=( A166  and  a28581a );
 a28583a <=( a28582a  and  a28577a );
 a28587a <=( A234  and  (not A233) );
 a28588a <=( A232  and  a28587a );
 a28592a <=( A299  and  (not A298) );
 a28593a <=( A236  and  a28592a );
 a28594a <=( a28593a  and  a28588a );
 a28598a <=( (not A167)  and  (not A168) );
 a28599a <=( (not A170)  and  a28598a );
 a28603a <=( A200  and  (not A199) );
 a28604a <=( A166  and  a28603a );
 a28605a <=( a28604a  and  a28599a );
 a28609a <=( A234  and  (not A233) );
 a28610a <=( A232  and  a28609a );
 a28614a <=( A266  and  (not A265) );
 a28615a <=( A236  and  a28614a );
 a28616a <=( a28615a  and  a28610a );
 a28620a <=( (not A167)  and  (not A168) );
 a28621a <=( (not A170)  and  a28620a );
 a28625a <=( A200  and  (not A199) );
 a28626a <=( A166  and  a28625a );
 a28627a <=( a28626a  and  a28621a );
 a28631a <=( A265  and  (not A233) );
 a28632a <=( (not A232)  and  a28631a );
 a28636a <=( (not A300)  and  A298 );
 a28637a <=( A266  and  a28636a );
 a28638a <=( a28637a  and  a28632a );
 a28642a <=( (not A167)  and  (not A168) );
 a28643a <=( (not A170)  and  a28642a );
 a28647a <=( A200  and  (not A199) );
 a28648a <=( A166  and  a28647a );
 a28649a <=( a28648a  and  a28643a );
 a28653a <=( A265  and  (not A233) );
 a28654a <=( (not A232)  and  a28653a );
 a28658a <=( A299  and  A298 );
 a28659a <=( A266  and  a28658a );
 a28660a <=( a28659a  and  a28654a );
 a28664a <=( (not A167)  and  (not A168) );
 a28665a <=( (not A170)  and  a28664a );
 a28669a <=( A200  and  (not A199) );
 a28670a <=( A166  and  a28669a );
 a28671a <=( a28670a  and  a28665a );
 a28675a <=( A265  and  (not A233) );
 a28676a <=( (not A232)  and  a28675a );
 a28680a <=( (not A299)  and  (not A298) );
 a28681a <=( A266  and  a28680a );
 a28682a <=( a28681a  and  a28676a );
 a28686a <=( (not A167)  and  (not A168) );
 a28687a <=( (not A170)  and  a28686a );
 a28691a <=( A200  and  (not A199) );
 a28692a <=( A166  and  a28691a );
 a28693a <=( a28692a  and  a28687a );
 a28697a <=( (not A266)  and  (not A233) );
 a28698a <=( (not A232)  and  a28697a );
 a28702a <=( (not A300)  and  A298 );
 a28703a <=( (not A267)  and  a28702a );
 a28704a <=( a28703a  and  a28698a );
 a28708a <=( (not A167)  and  (not A168) );
 a28709a <=( (not A170)  and  a28708a );
 a28713a <=( A200  and  (not A199) );
 a28714a <=( A166  and  a28713a );
 a28715a <=( a28714a  and  a28709a );
 a28719a <=( (not A266)  and  (not A233) );
 a28720a <=( (not A232)  and  a28719a );
 a28724a <=( A299  and  A298 );
 a28725a <=( (not A267)  and  a28724a );
 a28726a <=( a28725a  and  a28720a );
 a28730a <=( (not A167)  and  (not A168) );
 a28731a <=( (not A170)  and  a28730a );
 a28735a <=( A200  and  (not A199) );
 a28736a <=( A166  and  a28735a );
 a28737a <=( a28736a  and  a28731a );
 a28741a <=( (not A266)  and  (not A233) );
 a28742a <=( (not A232)  and  a28741a );
 a28746a <=( (not A299)  and  (not A298) );
 a28747a <=( (not A267)  and  a28746a );
 a28748a <=( a28747a  and  a28742a );
 a28752a <=( (not A167)  and  (not A168) );
 a28753a <=( (not A170)  and  a28752a );
 a28757a <=( A200  and  (not A199) );
 a28758a <=( A166  and  a28757a );
 a28759a <=( a28758a  and  a28753a );
 a28763a <=( (not A265)  and  (not A233) );
 a28764a <=( (not A232)  and  a28763a );
 a28768a <=( (not A300)  and  A298 );
 a28769a <=( (not A266)  and  a28768a );
 a28770a <=( a28769a  and  a28764a );
 a28774a <=( (not A167)  and  (not A168) );
 a28775a <=( (not A170)  and  a28774a );
 a28779a <=( A200  and  (not A199) );
 a28780a <=( A166  and  a28779a );
 a28781a <=( a28780a  and  a28775a );
 a28785a <=( (not A265)  and  (not A233) );
 a28786a <=( (not A232)  and  a28785a );
 a28790a <=( A299  and  A298 );
 a28791a <=( (not A266)  and  a28790a );
 a28792a <=( a28791a  and  a28786a );
 a28796a <=( (not A167)  and  (not A168) );
 a28797a <=( (not A170)  and  a28796a );
 a28801a <=( A200  and  (not A199) );
 a28802a <=( A166  and  a28801a );
 a28803a <=( a28802a  and  a28797a );
 a28807a <=( (not A265)  and  (not A233) );
 a28808a <=( (not A232)  and  a28807a );
 a28812a <=( (not A299)  and  (not A298) );
 a28813a <=( (not A266)  and  a28812a );
 a28814a <=( a28813a  and  a28808a );
 a28818a <=( A167  and  (not A168) );
 a28819a <=( A169  and  a28818a );
 a28823a <=( A200  and  (not A199) );
 a28824a <=( (not A166)  and  a28823a );
 a28825a <=( a28824a  and  a28819a );
 a28829a <=( A265  and  A233 );
 a28830a <=( A232  and  a28829a );
 a28834a <=( (not A300)  and  (not A299) );
 a28835a <=( (not A267)  and  a28834a );
 a28836a <=( a28835a  and  a28830a );
 a28840a <=( A167  and  (not A168) );
 a28841a <=( A169  and  a28840a );
 a28845a <=( A200  and  (not A199) );
 a28846a <=( (not A166)  and  a28845a );
 a28847a <=( a28846a  and  a28841a );
 a28851a <=( A265  and  A233 );
 a28852a <=( A232  and  a28851a );
 a28856a <=( A299  and  A298 );
 a28857a <=( (not A267)  and  a28856a );
 a28858a <=( a28857a  and  a28852a );
 a28862a <=( A167  and  (not A168) );
 a28863a <=( A169  and  a28862a );
 a28867a <=( A200  and  (not A199) );
 a28868a <=( (not A166)  and  a28867a );
 a28869a <=( a28868a  and  a28863a );
 a28873a <=( A265  and  A233 );
 a28874a <=( A232  and  a28873a );
 a28878a <=( (not A299)  and  (not A298) );
 a28879a <=( (not A267)  and  a28878a );
 a28880a <=( a28879a  and  a28874a );
 a28884a <=( A167  and  (not A168) );
 a28885a <=( A169  and  a28884a );
 a28889a <=( A200  and  (not A199) );
 a28890a <=( (not A166)  and  a28889a );
 a28891a <=( a28890a  and  a28885a );
 a28895a <=( A265  and  A233 );
 a28896a <=( A232  and  a28895a );
 a28900a <=( (not A300)  and  (not A299) );
 a28901a <=( A266  and  a28900a );
 a28902a <=( a28901a  and  a28896a );
 a28906a <=( A167  and  (not A168) );
 a28907a <=( A169  and  a28906a );
 a28911a <=( A200  and  (not A199) );
 a28912a <=( (not A166)  and  a28911a );
 a28913a <=( a28912a  and  a28907a );
 a28917a <=( A265  and  A233 );
 a28918a <=( A232  and  a28917a );
 a28922a <=( A299  and  A298 );
 a28923a <=( A266  and  a28922a );
 a28924a <=( a28923a  and  a28918a );
 a28928a <=( A167  and  (not A168) );
 a28929a <=( A169  and  a28928a );
 a28933a <=( A200  and  (not A199) );
 a28934a <=( (not A166)  and  a28933a );
 a28935a <=( a28934a  and  a28929a );
 a28939a <=( A265  and  A233 );
 a28940a <=( A232  and  a28939a );
 a28944a <=( (not A299)  and  (not A298) );
 a28945a <=( A266  and  a28944a );
 a28946a <=( a28945a  and  a28940a );
 a28950a <=( A167  and  (not A168) );
 a28951a <=( A169  and  a28950a );
 a28955a <=( A200  and  (not A199) );
 a28956a <=( (not A166)  and  a28955a );
 a28957a <=( a28956a  and  a28951a );
 a28961a <=( (not A265)  and  A233 );
 a28962a <=( A232  and  a28961a );
 a28966a <=( (not A300)  and  (not A299) );
 a28967a <=( (not A266)  and  a28966a );
 a28968a <=( a28967a  and  a28962a );
 a28972a <=( A167  and  (not A168) );
 a28973a <=( A169  and  a28972a );
 a28977a <=( A200  and  (not A199) );
 a28978a <=( (not A166)  and  a28977a );
 a28979a <=( a28978a  and  a28973a );
 a28983a <=( (not A265)  and  A233 );
 a28984a <=( A232  and  a28983a );
 a28988a <=( A299  and  A298 );
 a28989a <=( (not A266)  and  a28988a );
 a28990a <=( a28989a  and  a28984a );
 a28994a <=( A167  and  (not A168) );
 a28995a <=( A169  and  a28994a );
 a28999a <=( A200  and  (not A199) );
 a29000a <=( (not A166)  and  a28999a );
 a29001a <=( a29000a  and  a28995a );
 a29005a <=( (not A265)  and  A233 );
 a29006a <=( A232  and  a29005a );
 a29010a <=( (not A299)  and  (not A298) );
 a29011a <=( (not A266)  and  a29010a );
 a29012a <=( a29011a  and  a29006a );
 a29016a <=( A167  and  (not A168) );
 a29017a <=( A169  and  a29016a );
 a29021a <=( A200  and  (not A199) );
 a29022a <=( (not A166)  and  a29021a );
 a29023a <=( a29022a  and  a29017a );
 a29027a <=( A298  and  A233 );
 a29028a <=( (not A232)  and  a29027a );
 a29032a <=( A301  and  A300 );
 a29033a <=( (not A299)  and  a29032a );
 a29034a <=( a29033a  and  a29028a );
 a29038a <=( A167  and  (not A168) );
 a29039a <=( A169  and  a29038a );
 a29043a <=( A200  and  (not A199) );
 a29044a <=( (not A166)  and  a29043a );
 a29045a <=( a29044a  and  a29039a );
 a29049a <=( A298  and  A233 );
 a29050a <=( (not A232)  and  a29049a );
 a29054a <=( A302  and  A300 );
 a29055a <=( (not A299)  and  a29054a );
 a29056a <=( a29055a  and  a29050a );
 a29060a <=( A167  and  (not A168) );
 a29061a <=( A169  and  a29060a );
 a29065a <=( A200  and  (not A199) );
 a29066a <=( (not A166)  and  a29065a );
 a29067a <=( a29066a  and  a29061a );
 a29071a <=( A265  and  A233 );
 a29072a <=( (not A232)  and  a29071a );
 a29076a <=( A268  and  A267 );
 a29077a <=( (not A266)  and  a29076a );
 a29078a <=( a29077a  and  a29072a );
 a29082a <=( A167  and  (not A168) );
 a29083a <=( A169  and  a29082a );
 a29087a <=( A200  and  (not A199) );
 a29088a <=( (not A166)  and  a29087a );
 a29089a <=( a29088a  and  a29083a );
 a29093a <=( A265  and  A233 );
 a29094a <=( (not A232)  and  a29093a );
 a29098a <=( A269  and  A267 );
 a29099a <=( (not A266)  and  a29098a );
 a29100a <=( a29099a  and  a29094a );
 a29104a <=( A167  and  (not A168) );
 a29105a <=( A169  and  a29104a );
 a29109a <=( A200  and  (not A199) );
 a29110a <=( (not A166)  and  a29109a );
 a29111a <=( a29110a  and  a29105a );
 a29115a <=( A265  and  (not A234) );
 a29116a <=( (not A233)  and  a29115a );
 a29120a <=( (not A300)  and  A298 );
 a29121a <=( A266  and  a29120a );
 a29122a <=( a29121a  and  a29116a );
 a29126a <=( A167  and  (not A168) );
 a29127a <=( A169  and  a29126a );
 a29131a <=( A200  and  (not A199) );
 a29132a <=( (not A166)  and  a29131a );
 a29133a <=( a29132a  and  a29127a );
 a29137a <=( A265  and  (not A234) );
 a29138a <=( (not A233)  and  a29137a );
 a29142a <=( A299  and  A298 );
 a29143a <=( A266  and  a29142a );
 a29144a <=( a29143a  and  a29138a );
 a29148a <=( A167  and  (not A168) );
 a29149a <=( A169  and  a29148a );
 a29153a <=( A200  and  (not A199) );
 a29154a <=( (not A166)  and  a29153a );
 a29155a <=( a29154a  and  a29149a );
 a29159a <=( A265  and  (not A234) );
 a29160a <=( (not A233)  and  a29159a );
 a29164a <=( (not A299)  and  (not A298) );
 a29165a <=( A266  and  a29164a );
 a29166a <=( a29165a  and  a29160a );
 a29170a <=( A167  and  (not A168) );
 a29171a <=( A169  and  a29170a );
 a29175a <=( A200  and  (not A199) );
 a29176a <=( (not A166)  and  a29175a );
 a29177a <=( a29176a  and  a29171a );
 a29181a <=( (not A266)  and  (not A234) );
 a29182a <=( (not A233)  and  a29181a );
 a29186a <=( (not A300)  and  A298 );
 a29187a <=( (not A267)  and  a29186a );
 a29188a <=( a29187a  and  a29182a );
 a29192a <=( A167  and  (not A168) );
 a29193a <=( A169  and  a29192a );
 a29197a <=( A200  and  (not A199) );
 a29198a <=( (not A166)  and  a29197a );
 a29199a <=( a29198a  and  a29193a );
 a29203a <=( (not A266)  and  (not A234) );
 a29204a <=( (not A233)  and  a29203a );
 a29208a <=( A299  and  A298 );
 a29209a <=( (not A267)  and  a29208a );
 a29210a <=( a29209a  and  a29204a );
 a29214a <=( A167  and  (not A168) );
 a29215a <=( A169  and  a29214a );
 a29219a <=( A200  and  (not A199) );
 a29220a <=( (not A166)  and  a29219a );
 a29221a <=( a29220a  and  a29215a );
 a29225a <=( (not A266)  and  (not A234) );
 a29226a <=( (not A233)  and  a29225a );
 a29230a <=( (not A299)  and  (not A298) );
 a29231a <=( (not A267)  and  a29230a );
 a29232a <=( a29231a  and  a29226a );
 a29236a <=( A167  and  (not A168) );
 a29237a <=( A169  and  a29236a );
 a29241a <=( A200  and  (not A199) );
 a29242a <=( (not A166)  and  a29241a );
 a29243a <=( a29242a  and  a29237a );
 a29247a <=( (not A265)  and  (not A234) );
 a29248a <=( (not A233)  and  a29247a );
 a29252a <=( (not A300)  and  A298 );
 a29253a <=( (not A266)  and  a29252a );
 a29254a <=( a29253a  and  a29248a );
 a29258a <=( A167  and  (not A168) );
 a29259a <=( A169  and  a29258a );
 a29263a <=( A200  and  (not A199) );
 a29264a <=( (not A166)  and  a29263a );
 a29265a <=( a29264a  and  a29259a );
 a29269a <=( (not A265)  and  (not A234) );
 a29270a <=( (not A233)  and  a29269a );
 a29274a <=( A299  and  A298 );
 a29275a <=( (not A266)  and  a29274a );
 a29276a <=( a29275a  and  a29270a );
 a29280a <=( A167  and  (not A168) );
 a29281a <=( A169  and  a29280a );
 a29285a <=( A200  and  (not A199) );
 a29286a <=( (not A166)  and  a29285a );
 a29287a <=( a29286a  and  a29281a );
 a29291a <=( (not A265)  and  (not A234) );
 a29292a <=( (not A233)  and  a29291a );
 a29296a <=( (not A299)  and  (not A298) );
 a29297a <=( (not A266)  and  a29296a );
 a29298a <=( a29297a  and  a29292a );
 a29302a <=( A167  and  (not A168) );
 a29303a <=( A169  and  a29302a );
 a29307a <=( A200  and  (not A199) );
 a29308a <=( (not A166)  and  a29307a );
 a29309a <=( a29308a  and  a29303a );
 a29313a <=( A234  and  (not A233) );
 a29314a <=( A232  and  a29313a );
 a29318a <=( A299  and  (not A298) );
 a29319a <=( A235  and  a29318a );
 a29320a <=( a29319a  and  a29314a );
 a29324a <=( A167  and  (not A168) );
 a29325a <=( A169  and  a29324a );
 a29329a <=( A200  and  (not A199) );
 a29330a <=( (not A166)  and  a29329a );
 a29331a <=( a29330a  and  a29325a );
 a29335a <=( A234  and  (not A233) );
 a29336a <=( A232  and  a29335a );
 a29340a <=( A266  and  (not A265) );
 a29341a <=( A235  and  a29340a );
 a29342a <=( a29341a  and  a29336a );
 a29346a <=( A167  and  (not A168) );
 a29347a <=( A169  and  a29346a );
 a29351a <=( A200  and  (not A199) );
 a29352a <=( (not A166)  and  a29351a );
 a29353a <=( a29352a  and  a29347a );
 a29357a <=( A234  and  (not A233) );
 a29358a <=( A232  and  a29357a );
 a29362a <=( A299  and  (not A298) );
 a29363a <=( A236  and  a29362a );
 a29364a <=( a29363a  and  a29358a );
 a29368a <=( A167  and  (not A168) );
 a29369a <=( A169  and  a29368a );
 a29373a <=( A200  and  (not A199) );
 a29374a <=( (not A166)  and  a29373a );
 a29375a <=( a29374a  and  a29369a );
 a29379a <=( A234  and  (not A233) );
 a29380a <=( A232  and  a29379a );
 a29384a <=( A266  and  (not A265) );
 a29385a <=( A236  and  a29384a );
 a29386a <=( a29385a  and  a29380a );
 a29390a <=( A167  and  (not A168) );
 a29391a <=( A169  and  a29390a );
 a29395a <=( A200  and  (not A199) );
 a29396a <=( (not A166)  and  a29395a );
 a29397a <=( a29396a  and  a29391a );
 a29401a <=( A265  and  (not A233) );
 a29402a <=( (not A232)  and  a29401a );
 a29406a <=( (not A300)  and  A298 );
 a29407a <=( A266  and  a29406a );
 a29408a <=( a29407a  and  a29402a );
 a29412a <=( A167  and  (not A168) );
 a29413a <=( A169  and  a29412a );
 a29417a <=( A200  and  (not A199) );
 a29418a <=( (not A166)  and  a29417a );
 a29419a <=( a29418a  and  a29413a );
 a29423a <=( A265  and  (not A233) );
 a29424a <=( (not A232)  and  a29423a );
 a29428a <=( A299  and  A298 );
 a29429a <=( A266  and  a29428a );
 a29430a <=( a29429a  and  a29424a );
 a29434a <=( A167  and  (not A168) );
 a29435a <=( A169  and  a29434a );
 a29439a <=( A200  and  (not A199) );
 a29440a <=( (not A166)  and  a29439a );
 a29441a <=( a29440a  and  a29435a );
 a29445a <=( A265  and  (not A233) );
 a29446a <=( (not A232)  and  a29445a );
 a29450a <=( (not A299)  and  (not A298) );
 a29451a <=( A266  and  a29450a );
 a29452a <=( a29451a  and  a29446a );
 a29456a <=( A167  and  (not A168) );
 a29457a <=( A169  and  a29456a );
 a29461a <=( A200  and  (not A199) );
 a29462a <=( (not A166)  and  a29461a );
 a29463a <=( a29462a  and  a29457a );
 a29467a <=( (not A266)  and  (not A233) );
 a29468a <=( (not A232)  and  a29467a );
 a29472a <=( (not A300)  and  A298 );
 a29473a <=( (not A267)  and  a29472a );
 a29474a <=( a29473a  and  a29468a );
 a29478a <=( A167  and  (not A168) );
 a29479a <=( A169  and  a29478a );
 a29483a <=( A200  and  (not A199) );
 a29484a <=( (not A166)  and  a29483a );
 a29485a <=( a29484a  and  a29479a );
 a29489a <=( (not A266)  and  (not A233) );
 a29490a <=( (not A232)  and  a29489a );
 a29494a <=( A299  and  A298 );
 a29495a <=( (not A267)  and  a29494a );
 a29496a <=( a29495a  and  a29490a );
 a29500a <=( A167  and  (not A168) );
 a29501a <=( A169  and  a29500a );
 a29505a <=( A200  and  (not A199) );
 a29506a <=( (not A166)  and  a29505a );
 a29507a <=( a29506a  and  a29501a );
 a29511a <=( (not A266)  and  (not A233) );
 a29512a <=( (not A232)  and  a29511a );
 a29516a <=( (not A299)  and  (not A298) );
 a29517a <=( (not A267)  and  a29516a );
 a29518a <=( a29517a  and  a29512a );
 a29522a <=( A167  and  (not A168) );
 a29523a <=( A169  and  a29522a );
 a29527a <=( A200  and  (not A199) );
 a29528a <=( (not A166)  and  a29527a );
 a29529a <=( a29528a  and  a29523a );
 a29533a <=( (not A265)  and  (not A233) );
 a29534a <=( (not A232)  and  a29533a );
 a29538a <=( (not A300)  and  A298 );
 a29539a <=( (not A266)  and  a29538a );
 a29540a <=( a29539a  and  a29534a );
 a29544a <=( A167  and  (not A168) );
 a29545a <=( A169  and  a29544a );
 a29549a <=( A200  and  (not A199) );
 a29550a <=( (not A166)  and  a29549a );
 a29551a <=( a29550a  and  a29545a );
 a29555a <=( (not A265)  and  (not A233) );
 a29556a <=( (not A232)  and  a29555a );
 a29560a <=( A299  and  A298 );
 a29561a <=( (not A266)  and  a29560a );
 a29562a <=( a29561a  and  a29556a );
 a29566a <=( A167  and  (not A168) );
 a29567a <=( A169  and  a29566a );
 a29571a <=( A200  and  (not A199) );
 a29572a <=( (not A166)  and  a29571a );
 a29573a <=( a29572a  and  a29567a );
 a29577a <=( (not A265)  and  (not A233) );
 a29578a <=( (not A232)  and  a29577a );
 a29582a <=( (not A299)  and  (not A298) );
 a29583a <=( (not A266)  and  a29582a );
 a29584a <=( a29583a  and  a29578a );
 a29588a <=( A167  and  (not A168) );
 a29589a <=( A169  and  a29588a );
 a29593a <=( (not A200)  and  A199 );
 a29594a <=( (not A166)  and  a29593a );
 a29595a <=( a29594a  and  a29589a );
 a29599a <=( (not A232)  and  A202 );
 a29600a <=( A201  and  a29599a );
 a29604a <=( A299  and  (not A298) );
 a29605a <=( A233  and  a29604a );
 a29606a <=( a29605a  and  a29600a );
 a29610a <=( A167  and  (not A168) );
 a29611a <=( A169  and  a29610a );
 a29615a <=( (not A200)  and  A199 );
 a29616a <=( (not A166)  and  a29615a );
 a29617a <=( a29616a  and  a29611a );
 a29621a <=( (not A232)  and  A202 );
 a29622a <=( A201  and  a29621a );
 a29626a <=( A266  and  (not A265) );
 a29627a <=( A233  and  a29626a );
 a29628a <=( a29627a  and  a29622a );
 a29632a <=( A167  and  (not A168) );
 a29633a <=( A169  and  a29632a );
 a29637a <=( (not A200)  and  A199 );
 a29638a <=( (not A166)  and  a29637a );
 a29639a <=( a29638a  and  a29633a );
 a29643a <=( (not A232)  and  A203 );
 a29644a <=( A201  and  a29643a );
 a29648a <=( A299  and  (not A298) );
 a29649a <=( A233  and  a29648a );
 a29650a <=( a29649a  and  a29644a );
 a29654a <=( A167  and  (not A168) );
 a29655a <=( A169  and  a29654a );
 a29659a <=( (not A200)  and  A199 );
 a29660a <=( (not A166)  and  a29659a );
 a29661a <=( a29660a  and  a29655a );
 a29665a <=( (not A232)  and  A203 );
 a29666a <=( A201  and  a29665a );
 a29670a <=( A266  and  (not A265) );
 a29671a <=( A233  and  a29670a );
 a29672a <=( a29671a  and  a29666a );
 a29676a <=( (not A167)  and  (not A168) );
 a29677a <=( A169  and  a29676a );
 a29681a <=( A200  and  (not A199) );
 a29682a <=( A166  and  a29681a );
 a29683a <=( a29682a  and  a29677a );
 a29687a <=( A265  and  A233 );
 a29688a <=( A232  and  a29687a );
 a29692a <=( (not A300)  and  (not A299) );
 a29693a <=( (not A267)  and  a29692a );
 a29694a <=( a29693a  and  a29688a );
 a29698a <=( (not A167)  and  (not A168) );
 a29699a <=( A169  and  a29698a );
 a29703a <=( A200  and  (not A199) );
 a29704a <=( A166  and  a29703a );
 a29705a <=( a29704a  and  a29699a );
 a29709a <=( A265  and  A233 );
 a29710a <=( A232  and  a29709a );
 a29714a <=( A299  and  A298 );
 a29715a <=( (not A267)  and  a29714a );
 a29716a <=( a29715a  and  a29710a );
 a29720a <=( (not A167)  and  (not A168) );
 a29721a <=( A169  and  a29720a );
 a29725a <=( A200  and  (not A199) );
 a29726a <=( A166  and  a29725a );
 a29727a <=( a29726a  and  a29721a );
 a29731a <=( A265  and  A233 );
 a29732a <=( A232  and  a29731a );
 a29736a <=( (not A299)  and  (not A298) );
 a29737a <=( (not A267)  and  a29736a );
 a29738a <=( a29737a  and  a29732a );
 a29742a <=( (not A167)  and  (not A168) );
 a29743a <=( A169  and  a29742a );
 a29747a <=( A200  and  (not A199) );
 a29748a <=( A166  and  a29747a );
 a29749a <=( a29748a  and  a29743a );
 a29753a <=( A265  and  A233 );
 a29754a <=( A232  and  a29753a );
 a29758a <=( (not A300)  and  (not A299) );
 a29759a <=( A266  and  a29758a );
 a29760a <=( a29759a  and  a29754a );
 a29764a <=( (not A167)  and  (not A168) );
 a29765a <=( A169  and  a29764a );
 a29769a <=( A200  and  (not A199) );
 a29770a <=( A166  and  a29769a );
 a29771a <=( a29770a  and  a29765a );
 a29775a <=( A265  and  A233 );
 a29776a <=( A232  and  a29775a );
 a29780a <=( A299  and  A298 );
 a29781a <=( A266  and  a29780a );
 a29782a <=( a29781a  and  a29776a );
 a29786a <=( (not A167)  and  (not A168) );
 a29787a <=( A169  and  a29786a );
 a29791a <=( A200  and  (not A199) );
 a29792a <=( A166  and  a29791a );
 a29793a <=( a29792a  and  a29787a );
 a29797a <=( A265  and  A233 );
 a29798a <=( A232  and  a29797a );
 a29802a <=( (not A299)  and  (not A298) );
 a29803a <=( A266  and  a29802a );
 a29804a <=( a29803a  and  a29798a );
 a29808a <=( (not A167)  and  (not A168) );
 a29809a <=( A169  and  a29808a );
 a29813a <=( A200  and  (not A199) );
 a29814a <=( A166  and  a29813a );
 a29815a <=( a29814a  and  a29809a );
 a29819a <=( (not A265)  and  A233 );
 a29820a <=( A232  and  a29819a );
 a29824a <=( (not A300)  and  (not A299) );
 a29825a <=( (not A266)  and  a29824a );
 a29826a <=( a29825a  and  a29820a );
 a29830a <=( (not A167)  and  (not A168) );
 a29831a <=( A169  and  a29830a );
 a29835a <=( A200  and  (not A199) );
 a29836a <=( A166  and  a29835a );
 a29837a <=( a29836a  and  a29831a );
 a29841a <=( (not A265)  and  A233 );
 a29842a <=( A232  and  a29841a );
 a29846a <=( A299  and  A298 );
 a29847a <=( (not A266)  and  a29846a );
 a29848a <=( a29847a  and  a29842a );
 a29852a <=( (not A167)  and  (not A168) );
 a29853a <=( A169  and  a29852a );
 a29857a <=( A200  and  (not A199) );
 a29858a <=( A166  and  a29857a );
 a29859a <=( a29858a  and  a29853a );
 a29863a <=( (not A265)  and  A233 );
 a29864a <=( A232  and  a29863a );
 a29868a <=( (not A299)  and  (not A298) );
 a29869a <=( (not A266)  and  a29868a );
 a29870a <=( a29869a  and  a29864a );
 a29874a <=( (not A167)  and  (not A168) );
 a29875a <=( A169  and  a29874a );
 a29879a <=( A200  and  (not A199) );
 a29880a <=( A166  and  a29879a );
 a29881a <=( a29880a  and  a29875a );
 a29885a <=( A298  and  A233 );
 a29886a <=( (not A232)  and  a29885a );
 a29890a <=( A301  and  A300 );
 a29891a <=( (not A299)  and  a29890a );
 a29892a <=( a29891a  and  a29886a );
 a29896a <=( (not A167)  and  (not A168) );
 a29897a <=( A169  and  a29896a );
 a29901a <=( A200  and  (not A199) );
 a29902a <=( A166  and  a29901a );
 a29903a <=( a29902a  and  a29897a );
 a29907a <=( A298  and  A233 );
 a29908a <=( (not A232)  and  a29907a );
 a29912a <=( A302  and  A300 );
 a29913a <=( (not A299)  and  a29912a );
 a29914a <=( a29913a  and  a29908a );
 a29918a <=( (not A167)  and  (not A168) );
 a29919a <=( A169  and  a29918a );
 a29923a <=( A200  and  (not A199) );
 a29924a <=( A166  and  a29923a );
 a29925a <=( a29924a  and  a29919a );
 a29929a <=( A265  and  A233 );
 a29930a <=( (not A232)  and  a29929a );
 a29934a <=( A268  and  A267 );
 a29935a <=( (not A266)  and  a29934a );
 a29936a <=( a29935a  and  a29930a );
 a29940a <=( (not A167)  and  (not A168) );
 a29941a <=( A169  and  a29940a );
 a29945a <=( A200  and  (not A199) );
 a29946a <=( A166  and  a29945a );
 a29947a <=( a29946a  and  a29941a );
 a29951a <=( A265  and  A233 );
 a29952a <=( (not A232)  and  a29951a );
 a29956a <=( A269  and  A267 );
 a29957a <=( (not A266)  and  a29956a );
 a29958a <=( a29957a  and  a29952a );
 a29962a <=( (not A167)  and  (not A168) );
 a29963a <=( A169  and  a29962a );
 a29967a <=( A200  and  (not A199) );
 a29968a <=( A166  and  a29967a );
 a29969a <=( a29968a  and  a29963a );
 a29973a <=( A265  and  (not A234) );
 a29974a <=( (not A233)  and  a29973a );
 a29978a <=( (not A300)  and  A298 );
 a29979a <=( A266  and  a29978a );
 a29980a <=( a29979a  and  a29974a );
 a29984a <=( (not A167)  and  (not A168) );
 a29985a <=( A169  and  a29984a );
 a29989a <=( A200  and  (not A199) );
 a29990a <=( A166  and  a29989a );
 a29991a <=( a29990a  and  a29985a );
 a29995a <=( A265  and  (not A234) );
 a29996a <=( (not A233)  and  a29995a );
 a30000a <=( A299  and  A298 );
 a30001a <=( A266  and  a30000a );
 a30002a <=( a30001a  and  a29996a );
 a30006a <=( (not A167)  and  (not A168) );
 a30007a <=( A169  and  a30006a );
 a30011a <=( A200  and  (not A199) );
 a30012a <=( A166  and  a30011a );
 a30013a <=( a30012a  and  a30007a );
 a30017a <=( A265  and  (not A234) );
 a30018a <=( (not A233)  and  a30017a );
 a30022a <=( (not A299)  and  (not A298) );
 a30023a <=( A266  and  a30022a );
 a30024a <=( a30023a  and  a30018a );
 a30028a <=( (not A167)  and  (not A168) );
 a30029a <=( A169  and  a30028a );
 a30033a <=( A200  and  (not A199) );
 a30034a <=( A166  and  a30033a );
 a30035a <=( a30034a  and  a30029a );
 a30039a <=( (not A266)  and  (not A234) );
 a30040a <=( (not A233)  and  a30039a );
 a30044a <=( (not A300)  and  A298 );
 a30045a <=( (not A267)  and  a30044a );
 a30046a <=( a30045a  and  a30040a );
 a30050a <=( (not A167)  and  (not A168) );
 a30051a <=( A169  and  a30050a );
 a30055a <=( A200  and  (not A199) );
 a30056a <=( A166  and  a30055a );
 a30057a <=( a30056a  and  a30051a );
 a30061a <=( (not A266)  and  (not A234) );
 a30062a <=( (not A233)  and  a30061a );
 a30066a <=( A299  and  A298 );
 a30067a <=( (not A267)  and  a30066a );
 a30068a <=( a30067a  and  a30062a );
 a30072a <=( (not A167)  and  (not A168) );
 a30073a <=( A169  and  a30072a );
 a30077a <=( A200  and  (not A199) );
 a30078a <=( A166  and  a30077a );
 a30079a <=( a30078a  and  a30073a );
 a30083a <=( (not A266)  and  (not A234) );
 a30084a <=( (not A233)  and  a30083a );
 a30088a <=( (not A299)  and  (not A298) );
 a30089a <=( (not A267)  and  a30088a );
 a30090a <=( a30089a  and  a30084a );
 a30094a <=( (not A167)  and  (not A168) );
 a30095a <=( A169  and  a30094a );
 a30099a <=( A200  and  (not A199) );
 a30100a <=( A166  and  a30099a );
 a30101a <=( a30100a  and  a30095a );
 a30105a <=( (not A265)  and  (not A234) );
 a30106a <=( (not A233)  and  a30105a );
 a30110a <=( (not A300)  and  A298 );
 a30111a <=( (not A266)  and  a30110a );
 a30112a <=( a30111a  and  a30106a );
 a30116a <=( (not A167)  and  (not A168) );
 a30117a <=( A169  and  a30116a );
 a30121a <=( A200  and  (not A199) );
 a30122a <=( A166  and  a30121a );
 a30123a <=( a30122a  and  a30117a );
 a30127a <=( (not A265)  and  (not A234) );
 a30128a <=( (not A233)  and  a30127a );
 a30132a <=( A299  and  A298 );
 a30133a <=( (not A266)  and  a30132a );
 a30134a <=( a30133a  and  a30128a );
 a30138a <=( (not A167)  and  (not A168) );
 a30139a <=( A169  and  a30138a );
 a30143a <=( A200  and  (not A199) );
 a30144a <=( A166  and  a30143a );
 a30145a <=( a30144a  and  a30139a );
 a30149a <=( (not A265)  and  (not A234) );
 a30150a <=( (not A233)  and  a30149a );
 a30154a <=( (not A299)  and  (not A298) );
 a30155a <=( (not A266)  and  a30154a );
 a30156a <=( a30155a  and  a30150a );
 a30160a <=( (not A167)  and  (not A168) );
 a30161a <=( A169  and  a30160a );
 a30165a <=( A200  and  (not A199) );
 a30166a <=( A166  and  a30165a );
 a30167a <=( a30166a  and  a30161a );
 a30171a <=( A234  and  (not A233) );
 a30172a <=( A232  and  a30171a );
 a30176a <=( A299  and  (not A298) );
 a30177a <=( A235  and  a30176a );
 a30178a <=( a30177a  and  a30172a );
 a30182a <=( (not A167)  and  (not A168) );
 a30183a <=( A169  and  a30182a );
 a30187a <=( A200  and  (not A199) );
 a30188a <=( A166  and  a30187a );
 a30189a <=( a30188a  and  a30183a );
 a30193a <=( A234  and  (not A233) );
 a30194a <=( A232  and  a30193a );
 a30198a <=( A266  and  (not A265) );
 a30199a <=( A235  and  a30198a );
 a30200a <=( a30199a  and  a30194a );
 a30204a <=( (not A167)  and  (not A168) );
 a30205a <=( A169  and  a30204a );
 a30209a <=( A200  and  (not A199) );
 a30210a <=( A166  and  a30209a );
 a30211a <=( a30210a  and  a30205a );
 a30215a <=( A234  and  (not A233) );
 a30216a <=( A232  and  a30215a );
 a30220a <=( A299  and  (not A298) );
 a30221a <=( A236  and  a30220a );
 a30222a <=( a30221a  and  a30216a );
 a30226a <=( (not A167)  and  (not A168) );
 a30227a <=( A169  and  a30226a );
 a30231a <=( A200  and  (not A199) );
 a30232a <=( A166  and  a30231a );
 a30233a <=( a30232a  and  a30227a );
 a30237a <=( A234  and  (not A233) );
 a30238a <=( A232  and  a30237a );
 a30242a <=( A266  and  (not A265) );
 a30243a <=( A236  and  a30242a );
 a30244a <=( a30243a  and  a30238a );
 a30248a <=( (not A167)  and  (not A168) );
 a30249a <=( A169  and  a30248a );
 a30253a <=( A200  and  (not A199) );
 a30254a <=( A166  and  a30253a );
 a30255a <=( a30254a  and  a30249a );
 a30259a <=( A265  and  (not A233) );
 a30260a <=( (not A232)  and  a30259a );
 a30264a <=( (not A300)  and  A298 );
 a30265a <=( A266  and  a30264a );
 a30266a <=( a30265a  and  a30260a );
 a30270a <=( (not A167)  and  (not A168) );
 a30271a <=( A169  and  a30270a );
 a30275a <=( A200  and  (not A199) );
 a30276a <=( A166  and  a30275a );
 a30277a <=( a30276a  and  a30271a );
 a30281a <=( A265  and  (not A233) );
 a30282a <=( (not A232)  and  a30281a );
 a30286a <=( A299  and  A298 );
 a30287a <=( A266  and  a30286a );
 a30288a <=( a30287a  and  a30282a );
 a30292a <=( (not A167)  and  (not A168) );
 a30293a <=( A169  and  a30292a );
 a30297a <=( A200  and  (not A199) );
 a30298a <=( A166  and  a30297a );
 a30299a <=( a30298a  and  a30293a );
 a30303a <=( A265  and  (not A233) );
 a30304a <=( (not A232)  and  a30303a );
 a30308a <=( (not A299)  and  (not A298) );
 a30309a <=( A266  and  a30308a );
 a30310a <=( a30309a  and  a30304a );
 a30314a <=( (not A167)  and  (not A168) );
 a30315a <=( A169  and  a30314a );
 a30319a <=( A200  and  (not A199) );
 a30320a <=( A166  and  a30319a );
 a30321a <=( a30320a  and  a30315a );
 a30325a <=( (not A266)  and  (not A233) );
 a30326a <=( (not A232)  and  a30325a );
 a30330a <=( (not A300)  and  A298 );
 a30331a <=( (not A267)  and  a30330a );
 a30332a <=( a30331a  and  a30326a );
 a30336a <=( (not A167)  and  (not A168) );
 a30337a <=( A169  and  a30336a );
 a30341a <=( A200  and  (not A199) );
 a30342a <=( A166  and  a30341a );
 a30343a <=( a30342a  and  a30337a );
 a30347a <=( (not A266)  and  (not A233) );
 a30348a <=( (not A232)  and  a30347a );
 a30352a <=( A299  and  A298 );
 a30353a <=( (not A267)  and  a30352a );
 a30354a <=( a30353a  and  a30348a );
 a30358a <=( (not A167)  and  (not A168) );
 a30359a <=( A169  and  a30358a );
 a30363a <=( A200  and  (not A199) );
 a30364a <=( A166  and  a30363a );
 a30365a <=( a30364a  and  a30359a );
 a30369a <=( (not A266)  and  (not A233) );
 a30370a <=( (not A232)  and  a30369a );
 a30374a <=( (not A299)  and  (not A298) );
 a30375a <=( (not A267)  and  a30374a );
 a30376a <=( a30375a  and  a30370a );
 a30380a <=( (not A167)  and  (not A168) );
 a30381a <=( A169  and  a30380a );
 a30385a <=( A200  and  (not A199) );
 a30386a <=( A166  and  a30385a );
 a30387a <=( a30386a  and  a30381a );
 a30391a <=( (not A265)  and  (not A233) );
 a30392a <=( (not A232)  and  a30391a );
 a30396a <=( (not A300)  and  A298 );
 a30397a <=( (not A266)  and  a30396a );
 a30398a <=( a30397a  and  a30392a );
 a30402a <=( (not A167)  and  (not A168) );
 a30403a <=( A169  and  a30402a );
 a30407a <=( A200  and  (not A199) );
 a30408a <=( A166  and  a30407a );
 a30409a <=( a30408a  and  a30403a );
 a30413a <=( (not A265)  and  (not A233) );
 a30414a <=( (not A232)  and  a30413a );
 a30418a <=( A299  and  A298 );
 a30419a <=( (not A266)  and  a30418a );
 a30420a <=( a30419a  and  a30414a );
 a30424a <=( (not A167)  and  (not A168) );
 a30425a <=( A169  and  a30424a );
 a30429a <=( A200  and  (not A199) );
 a30430a <=( A166  and  a30429a );
 a30431a <=( a30430a  and  a30425a );
 a30435a <=( (not A265)  and  (not A233) );
 a30436a <=( (not A232)  and  a30435a );
 a30440a <=( (not A299)  and  (not A298) );
 a30441a <=( (not A266)  and  a30440a );
 a30442a <=( a30441a  and  a30436a );
 a30446a <=( (not A167)  and  (not A168) );
 a30447a <=( A169  and  a30446a );
 a30451a <=( (not A200)  and  A199 );
 a30452a <=( A166  and  a30451a );
 a30453a <=( a30452a  and  a30447a );
 a30457a <=( (not A232)  and  A202 );
 a30458a <=( A201  and  a30457a );
 a30462a <=( A299  and  (not A298) );
 a30463a <=( A233  and  a30462a );
 a30464a <=( a30463a  and  a30458a );
 a30468a <=( (not A167)  and  (not A168) );
 a30469a <=( A169  and  a30468a );
 a30473a <=( (not A200)  and  A199 );
 a30474a <=( A166  and  a30473a );
 a30475a <=( a30474a  and  a30469a );
 a30479a <=( (not A232)  and  A202 );
 a30480a <=( A201  and  a30479a );
 a30484a <=( A266  and  (not A265) );
 a30485a <=( A233  and  a30484a );
 a30486a <=( a30485a  and  a30480a );
 a30490a <=( (not A167)  and  (not A168) );
 a30491a <=( A169  and  a30490a );
 a30495a <=( (not A200)  and  A199 );
 a30496a <=( A166  and  a30495a );
 a30497a <=( a30496a  and  a30491a );
 a30501a <=( (not A232)  and  A203 );
 a30502a <=( A201  and  a30501a );
 a30506a <=( A299  and  (not A298) );
 a30507a <=( A233  and  a30506a );
 a30508a <=( a30507a  and  a30502a );
 a30512a <=( (not A167)  and  (not A168) );
 a30513a <=( A169  and  a30512a );
 a30517a <=( (not A200)  and  A199 );
 a30518a <=( A166  and  a30517a );
 a30519a <=( a30518a  and  a30513a );
 a30523a <=( (not A232)  and  A203 );
 a30524a <=( A201  and  a30523a );
 a30528a <=( A266  and  (not A265) );
 a30529a <=( A233  and  a30528a );
 a30530a <=( a30529a  and  a30524a );
 a30534a <=( (not A168)  and  A169 );
 a30535a <=( A170  and  a30534a );
 a30539a <=( (not A200)  and  A199 );
 a30540a <=( A166  and  a30539a );
 a30541a <=( a30540a  and  a30535a );
 a30545a <=( (not A232)  and  A202 );
 a30546a <=( A201  and  a30545a );
 a30550a <=( A299  and  (not A298) );
 a30551a <=( A233  and  a30550a );
 a30552a <=( a30551a  and  a30546a );
 a30556a <=( (not A168)  and  A169 );
 a30557a <=( A170  and  a30556a );
 a30561a <=( (not A200)  and  A199 );
 a30562a <=( A166  and  a30561a );
 a30563a <=( a30562a  and  a30557a );
 a30567a <=( (not A232)  and  A202 );
 a30568a <=( A201  and  a30567a );
 a30572a <=( A266  and  (not A265) );
 a30573a <=( A233  and  a30572a );
 a30574a <=( a30573a  and  a30568a );
 a30578a <=( (not A168)  and  A169 );
 a30579a <=( A170  and  a30578a );
 a30583a <=( (not A200)  and  A199 );
 a30584a <=( A166  and  a30583a );
 a30585a <=( a30584a  and  a30579a );
 a30589a <=( (not A232)  and  A203 );
 a30590a <=( A201  and  a30589a );
 a30594a <=( A299  and  (not A298) );
 a30595a <=( A233  and  a30594a );
 a30596a <=( a30595a  and  a30590a );
 a30600a <=( (not A168)  and  A169 );
 a30601a <=( A170  and  a30600a );
 a30605a <=( (not A200)  and  A199 );
 a30606a <=( A166  and  a30605a );
 a30607a <=( a30606a  and  a30601a );
 a30611a <=( (not A232)  and  A203 );
 a30612a <=( A201  and  a30611a );
 a30616a <=( A266  and  (not A265) );
 a30617a <=( A233  and  a30616a );
 a30618a <=( a30617a  and  a30612a );
 a30622a <=( A167  and  A169 );
 a30623a <=( (not A170)  and  a30622a );
 a30627a <=( A200  and  A199 );
 a30628a <=( A166  and  a30627a );
 a30629a <=( a30628a  and  a30623a );
 a30633a <=( A265  and  A233 );
 a30634a <=( A232  and  a30633a );
 a30638a <=( (not A300)  and  (not A299) );
 a30639a <=( (not A267)  and  a30638a );
 a30640a <=( a30639a  and  a30634a );
 a30644a <=( A167  and  A169 );
 a30645a <=( (not A170)  and  a30644a );
 a30649a <=( A200  and  A199 );
 a30650a <=( A166  and  a30649a );
 a30651a <=( a30650a  and  a30645a );
 a30655a <=( A265  and  A233 );
 a30656a <=( A232  and  a30655a );
 a30660a <=( A299  and  A298 );
 a30661a <=( (not A267)  and  a30660a );
 a30662a <=( a30661a  and  a30656a );
 a30666a <=( A167  and  A169 );
 a30667a <=( (not A170)  and  a30666a );
 a30671a <=( A200  and  A199 );
 a30672a <=( A166  and  a30671a );
 a30673a <=( a30672a  and  a30667a );
 a30677a <=( A265  and  A233 );
 a30678a <=( A232  and  a30677a );
 a30682a <=( (not A299)  and  (not A298) );
 a30683a <=( (not A267)  and  a30682a );
 a30684a <=( a30683a  and  a30678a );
 a30688a <=( A167  and  A169 );
 a30689a <=( (not A170)  and  a30688a );
 a30693a <=( A200  and  A199 );
 a30694a <=( A166  and  a30693a );
 a30695a <=( a30694a  and  a30689a );
 a30699a <=( A265  and  A233 );
 a30700a <=( A232  and  a30699a );
 a30704a <=( (not A300)  and  (not A299) );
 a30705a <=( A266  and  a30704a );
 a30706a <=( a30705a  and  a30700a );
 a30710a <=( A167  and  A169 );
 a30711a <=( (not A170)  and  a30710a );
 a30715a <=( A200  and  A199 );
 a30716a <=( A166  and  a30715a );
 a30717a <=( a30716a  and  a30711a );
 a30721a <=( A265  and  A233 );
 a30722a <=( A232  and  a30721a );
 a30726a <=( A299  and  A298 );
 a30727a <=( A266  and  a30726a );
 a30728a <=( a30727a  and  a30722a );
 a30732a <=( A167  and  A169 );
 a30733a <=( (not A170)  and  a30732a );
 a30737a <=( A200  and  A199 );
 a30738a <=( A166  and  a30737a );
 a30739a <=( a30738a  and  a30733a );
 a30743a <=( A265  and  A233 );
 a30744a <=( A232  and  a30743a );
 a30748a <=( (not A299)  and  (not A298) );
 a30749a <=( A266  and  a30748a );
 a30750a <=( a30749a  and  a30744a );
 a30754a <=( A167  and  A169 );
 a30755a <=( (not A170)  and  a30754a );
 a30759a <=( A200  and  A199 );
 a30760a <=( A166  and  a30759a );
 a30761a <=( a30760a  and  a30755a );
 a30765a <=( (not A265)  and  A233 );
 a30766a <=( A232  and  a30765a );
 a30770a <=( (not A300)  and  (not A299) );
 a30771a <=( (not A266)  and  a30770a );
 a30772a <=( a30771a  and  a30766a );
 a30776a <=( A167  and  A169 );
 a30777a <=( (not A170)  and  a30776a );
 a30781a <=( A200  and  A199 );
 a30782a <=( A166  and  a30781a );
 a30783a <=( a30782a  and  a30777a );
 a30787a <=( (not A265)  and  A233 );
 a30788a <=( A232  and  a30787a );
 a30792a <=( A299  and  A298 );
 a30793a <=( (not A266)  and  a30792a );
 a30794a <=( a30793a  and  a30788a );
 a30798a <=( A167  and  A169 );
 a30799a <=( (not A170)  and  a30798a );
 a30803a <=( A200  and  A199 );
 a30804a <=( A166  and  a30803a );
 a30805a <=( a30804a  and  a30799a );
 a30809a <=( (not A265)  and  A233 );
 a30810a <=( A232  and  a30809a );
 a30814a <=( (not A299)  and  (not A298) );
 a30815a <=( (not A266)  and  a30814a );
 a30816a <=( a30815a  and  a30810a );
 a30820a <=( A167  and  A169 );
 a30821a <=( (not A170)  and  a30820a );
 a30825a <=( A200  and  A199 );
 a30826a <=( A166  and  a30825a );
 a30827a <=( a30826a  and  a30821a );
 a30831a <=( A298  and  A233 );
 a30832a <=( (not A232)  and  a30831a );
 a30836a <=( A301  and  A300 );
 a30837a <=( (not A299)  and  a30836a );
 a30838a <=( a30837a  and  a30832a );
 a30842a <=( A167  and  A169 );
 a30843a <=( (not A170)  and  a30842a );
 a30847a <=( A200  and  A199 );
 a30848a <=( A166  and  a30847a );
 a30849a <=( a30848a  and  a30843a );
 a30853a <=( A298  and  A233 );
 a30854a <=( (not A232)  and  a30853a );
 a30858a <=( A302  and  A300 );
 a30859a <=( (not A299)  and  a30858a );
 a30860a <=( a30859a  and  a30854a );
 a30864a <=( A167  and  A169 );
 a30865a <=( (not A170)  and  a30864a );
 a30869a <=( A200  and  A199 );
 a30870a <=( A166  and  a30869a );
 a30871a <=( a30870a  and  a30865a );
 a30875a <=( A265  and  A233 );
 a30876a <=( (not A232)  and  a30875a );
 a30880a <=( A268  and  A267 );
 a30881a <=( (not A266)  and  a30880a );
 a30882a <=( a30881a  and  a30876a );
 a30886a <=( A167  and  A169 );
 a30887a <=( (not A170)  and  a30886a );
 a30891a <=( A200  and  A199 );
 a30892a <=( A166  and  a30891a );
 a30893a <=( a30892a  and  a30887a );
 a30897a <=( A265  and  A233 );
 a30898a <=( (not A232)  and  a30897a );
 a30902a <=( A269  and  A267 );
 a30903a <=( (not A266)  and  a30902a );
 a30904a <=( a30903a  and  a30898a );
 a30908a <=( A167  and  A169 );
 a30909a <=( (not A170)  and  a30908a );
 a30913a <=( A200  and  A199 );
 a30914a <=( A166  and  a30913a );
 a30915a <=( a30914a  and  a30909a );
 a30919a <=( A265  and  (not A234) );
 a30920a <=( (not A233)  and  a30919a );
 a30924a <=( (not A300)  and  A298 );
 a30925a <=( A266  and  a30924a );
 a30926a <=( a30925a  and  a30920a );
 a30930a <=( A167  and  A169 );
 a30931a <=( (not A170)  and  a30930a );
 a30935a <=( A200  and  A199 );
 a30936a <=( A166  and  a30935a );
 a30937a <=( a30936a  and  a30931a );
 a30941a <=( A265  and  (not A234) );
 a30942a <=( (not A233)  and  a30941a );
 a30946a <=( A299  and  A298 );
 a30947a <=( A266  and  a30946a );
 a30948a <=( a30947a  and  a30942a );
 a30952a <=( A167  and  A169 );
 a30953a <=( (not A170)  and  a30952a );
 a30957a <=( A200  and  A199 );
 a30958a <=( A166  and  a30957a );
 a30959a <=( a30958a  and  a30953a );
 a30963a <=( A265  and  (not A234) );
 a30964a <=( (not A233)  and  a30963a );
 a30968a <=( (not A299)  and  (not A298) );
 a30969a <=( A266  and  a30968a );
 a30970a <=( a30969a  and  a30964a );
 a30974a <=( A167  and  A169 );
 a30975a <=( (not A170)  and  a30974a );
 a30979a <=( A200  and  A199 );
 a30980a <=( A166  and  a30979a );
 a30981a <=( a30980a  and  a30975a );
 a30985a <=( (not A266)  and  (not A234) );
 a30986a <=( (not A233)  and  a30985a );
 a30990a <=( (not A300)  and  A298 );
 a30991a <=( (not A267)  and  a30990a );
 a30992a <=( a30991a  and  a30986a );
 a30996a <=( A167  and  A169 );
 a30997a <=( (not A170)  and  a30996a );
 a31001a <=( A200  and  A199 );
 a31002a <=( A166  and  a31001a );
 a31003a <=( a31002a  and  a30997a );
 a31007a <=( (not A266)  and  (not A234) );
 a31008a <=( (not A233)  and  a31007a );
 a31012a <=( A299  and  A298 );
 a31013a <=( (not A267)  and  a31012a );
 a31014a <=( a31013a  and  a31008a );
 a31018a <=( A167  and  A169 );
 a31019a <=( (not A170)  and  a31018a );
 a31023a <=( A200  and  A199 );
 a31024a <=( A166  and  a31023a );
 a31025a <=( a31024a  and  a31019a );
 a31029a <=( (not A266)  and  (not A234) );
 a31030a <=( (not A233)  and  a31029a );
 a31034a <=( (not A299)  and  (not A298) );
 a31035a <=( (not A267)  and  a31034a );
 a31036a <=( a31035a  and  a31030a );
 a31040a <=( A167  and  A169 );
 a31041a <=( (not A170)  and  a31040a );
 a31045a <=( A200  and  A199 );
 a31046a <=( A166  and  a31045a );
 a31047a <=( a31046a  and  a31041a );
 a31051a <=( (not A265)  and  (not A234) );
 a31052a <=( (not A233)  and  a31051a );
 a31056a <=( (not A300)  and  A298 );
 a31057a <=( (not A266)  and  a31056a );
 a31058a <=( a31057a  and  a31052a );
 a31062a <=( A167  and  A169 );
 a31063a <=( (not A170)  and  a31062a );
 a31067a <=( A200  and  A199 );
 a31068a <=( A166  and  a31067a );
 a31069a <=( a31068a  and  a31063a );
 a31073a <=( (not A265)  and  (not A234) );
 a31074a <=( (not A233)  and  a31073a );
 a31078a <=( A299  and  A298 );
 a31079a <=( (not A266)  and  a31078a );
 a31080a <=( a31079a  and  a31074a );
 a31084a <=( A167  and  A169 );
 a31085a <=( (not A170)  and  a31084a );
 a31089a <=( A200  and  A199 );
 a31090a <=( A166  and  a31089a );
 a31091a <=( a31090a  and  a31085a );
 a31095a <=( (not A265)  and  (not A234) );
 a31096a <=( (not A233)  and  a31095a );
 a31100a <=( (not A299)  and  (not A298) );
 a31101a <=( (not A266)  and  a31100a );
 a31102a <=( a31101a  and  a31096a );
 a31106a <=( A167  and  A169 );
 a31107a <=( (not A170)  and  a31106a );
 a31111a <=( A200  and  A199 );
 a31112a <=( A166  and  a31111a );
 a31113a <=( a31112a  and  a31107a );
 a31117a <=( A234  and  (not A233) );
 a31118a <=( A232  and  a31117a );
 a31122a <=( A299  and  (not A298) );
 a31123a <=( A235  and  a31122a );
 a31124a <=( a31123a  and  a31118a );
 a31128a <=( A167  and  A169 );
 a31129a <=( (not A170)  and  a31128a );
 a31133a <=( A200  and  A199 );
 a31134a <=( A166  and  a31133a );
 a31135a <=( a31134a  and  a31129a );
 a31139a <=( A234  and  (not A233) );
 a31140a <=( A232  and  a31139a );
 a31144a <=( A266  and  (not A265) );
 a31145a <=( A235  and  a31144a );
 a31146a <=( a31145a  and  a31140a );
 a31150a <=( A167  and  A169 );
 a31151a <=( (not A170)  and  a31150a );
 a31155a <=( A200  and  A199 );
 a31156a <=( A166  and  a31155a );
 a31157a <=( a31156a  and  a31151a );
 a31161a <=( A234  and  (not A233) );
 a31162a <=( A232  and  a31161a );
 a31166a <=( A299  and  (not A298) );
 a31167a <=( A236  and  a31166a );
 a31168a <=( a31167a  and  a31162a );
 a31172a <=( A167  and  A169 );
 a31173a <=( (not A170)  and  a31172a );
 a31177a <=( A200  and  A199 );
 a31178a <=( A166  and  a31177a );
 a31179a <=( a31178a  and  a31173a );
 a31183a <=( A234  and  (not A233) );
 a31184a <=( A232  and  a31183a );
 a31188a <=( A266  and  (not A265) );
 a31189a <=( A236  and  a31188a );
 a31190a <=( a31189a  and  a31184a );
 a31194a <=( A167  and  A169 );
 a31195a <=( (not A170)  and  a31194a );
 a31199a <=( A200  and  A199 );
 a31200a <=( A166  and  a31199a );
 a31201a <=( a31200a  and  a31195a );
 a31205a <=( A265  and  (not A233) );
 a31206a <=( (not A232)  and  a31205a );
 a31210a <=( (not A300)  and  A298 );
 a31211a <=( A266  and  a31210a );
 a31212a <=( a31211a  and  a31206a );
 a31216a <=( A167  and  A169 );
 a31217a <=( (not A170)  and  a31216a );
 a31221a <=( A200  and  A199 );
 a31222a <=( A166  and  a31221a );
 a31223a <=( a31222a  and  a31217a );
 a31227a <=( A265  and  (not A233) );
 a31228a <=( (not A232)  and  a31227a );
 a31232a <=( A299  and  A298 );
 a31233a <=( A266  and  a31232a );
 a31234a <=( a31233a  and  a31228a );
 a31238a <=( A167  and  A169 );
 a31239a <=( (not A170)  and  a31238a );
 a31243a <=( A200  and  A199 );
 a31244a <=( A166  and  a31243a );
 a31245a <=( a31244a  and  a31239a );
 a31249a <=( A265  and  (not A233) );
 a31250a <=( (not A232)  and  a31249a );
 a31254a <=( (not A299)  and  (not A298) );
 a31255a <=( A266  and  a31254a );
 a31256a <=( a31255a  and  a31250a );
 a31260a <=( A167  and  A169 );
 a31261a <=( (not A170)  and  a31260a );
 a31265a <=( A200  and  A199 );
 a31266a <=( A166  and  a31265a );
 a31267a <=( a31266a  and  a31261a );
 a31271a <=( (not A266)  and  (not A233) );
 a31272a <=( (not A232)  and  a31271a );
 a31276a <=( (not A300)  and  A298 );
 a31277a <=( (not A267)  and  a31276a );
 a31278a <=( a31277a  and  a31272a );
 a31282a <=( A167  and  A169 );
 a31283a <=( (not A170)  and  a31282a );
 a31287a <=( A200  and  A199 );
 a31288a <=( A166  and  a31287a );
 a31289a <=( a31288a  and  a31283a );
 a31293a <=( (not A266)  and  (not A233) );
 a31294a <=( (not A232)  and  a31293a );
 a31298a <=( A299  and  A298 );
 a31299a <=( (not A267)  and  a31298a );
 a31300a <=( a31299a  and  a31294a );
 a31304a <=( A167  and  A169 );
 a31305a <=( (not A170)  and  a31304a );
 a31309a <=( A200  and  A199 );
 a31310a <=( A166  and  a31309a );
 a31311a <=( a31310a  and  a31305a );
 a31315a <=( (not A266)  and  (not A233) );
 a31316a <=( (not A232)  and  a31315a );
 a31320a <=( (not A299)  and  (not A298) );
 a31321a <=( (not A267)  and  a31320a );
 a31322a <=( a31321a  and  a31316a );
 a31326a <=( A167  and  A169 );
 a31327a <=( (not A170)  and  a31326a );
 a31331a <=( A200  and  A199 );
 a31332a <=( A166  and  a31331a );
 a31333a <=( a31332a  and  a31327a );
 a31337a <=( (not A265)  and  (not A233) );
 a31338a <=( (not A232)  and  a31337a );
 a31342a <=( (not A300)  and  A298 );
 a31343a <=( (not A266)  and  a31342a );
 a31344a <=( a31343a  and  a31338a );
 a31348a <=( A167  and  A169 );
 a31349a <=( (not A170)  and  a31348a );
 a31353a <=( A200  and  A199 );
 a31354a <=( A166  and  a31353a );
 a31355a <=( a31354a  and  a31349a );
 a31359a <=( (not A265)  and  (not A233) );
 a31360a <=( (not A232)  and  a31359a );
 a31364a <=( A299  and  A298 );
 a31365a <=( (not A266)  and  a31364a );
 a31366a <=( a31365a  and  a31360a );
 a31370a <=( A167  and  A169 );
 a31371a <=( (not A170)  and  a31370a );
 a31375a <=( A200  and  A199 );
 a31376a <=( A166  and  a31375a );
 a31377a <=( a31376a  and  a31371a );
 a31381a <=( (not A265)  and  (not A233) );
 a31382a <=( (not A232)  and  a31381a );
 a31386a <=( (not A299)  and  (not A298) );
 a31387a <=( (not A266)  and  a31386a );
 a31388a <=( a31387a  and  a31382a );
 a31392a <=( A167  and  A169 );
 a31393a <=( (not A170)  and  a31392a );
 a31397a <=( (not A201)  and  (not A200) );
 a31398a <=( A166  and  a31397a );
 a31399a <=( a31398a  and  a31393a );
 a31403a <=( A265  and  A233 );
 a31404a <=( A232  and  a31403a );
 a31408a <=( (not A300)  and  (not A299) );
 a31409a <=( (not A267)  and  a31408a );
 a31410a <=( a31409a  and  a31404a );
 a31414a <=( A167  and  A169 );
 a31415a <=( (not A170)  and  a31414a );
 a31419a <=( (not A201)  and  (not A200) );
 a31420a <=( A166  and  a31419a );
 a31421a <=( a31420a  and  a31415a );
 a31425a <=( A265  and  A233 );
 a31426a <=( A232  and  a31425a );
 a31430a <=( A299  and  A298 );
 a31431a <=( (not A267)  and  a31430a );
 a31432a <=( a31431a  and  a31426a );
 a31436a <=( A167  and  A169 );
 a31437a <=( (not A170)  and  a31436a );
 a31441a <=( (not A201)  and  (not A200) );
 a31442a <=( A166  and  a31441a );
 a31443a <=( a31442a  and  a31437a );
 a31447a <=( A265  and  A233 );
 a31448a <=( A232  and  a31447a );
 a31452a <=( (not A299)  and  (not A298) );
 a31453a <=( (not A267)  and  a31452a );
 a31454a <=( a31453a  and  a31448a );
 a31458a <=( A167  and  A169 );
 a31459a <=( (not A170)  and  a31458a );
 a31463a <=( (not A201)  and  (not A200) );
 a31464a <=( A166  and  a31463a );
 a31465a <=( a31464a  and  a31459a );
 a31469a <=( A265  and  A233 );
 a31470a <=( A232  and  a31469a );
 a31474a <=( (not A300)  and  (not A299) );
 a31475a <=( A266  and  a31474a );
 a31476a <=( a31475a  and  a31470a );
 a31480a <=( A167  and  A169 );
 a31481a <=( (not A170)  and  a31480a );
 a31485a <=( (not A201)  and  (not A200) );
 a31486a <=( A166  and  a31485a );
 a31487a <=( a31486a  and  a31481a );
 a31491a <=( A265  and  A233 );
 a31492a <=( A232  and  a31491a );
 a31496a <=( A299  and  A298 );
 a31497a <=( A266  and  a31496a );
 a31498a <=( a31497a  and  a31492a );
 a31502a <=( A167  and  A169 );
 a31503a <=( (not A170)  and  a31502a );
 a31507a <=( (not A201)  and  (not A200) );
 a31508a <=( A166  and  a31507a );
 a31509a <=( a31508a  and  a31503a );
 a31513a <=( A265  and  A233 );
 a31514a <=( A232  and  a31513a );
 a31518a <=( (not A299)  and  (not A298) );
 a31519a <=( A266  and  a31518a );
 a31520a <=( a31519a  and  a31514a );
 a31524a <=( A167  and  A169 );
 a31525a <=( (not A170)  and  a31524a );
 a31529a <=( (not A201)  and  (not A200) );
 a31530a <=( A166  and  a31529a );
 a31531a <=( a31530a  and  a31525a );
 a31535a <=( (not A265)  and  A233 );
 a31536a <=( A232  and  a31535a );
 a31540a <=( (not A300)  and  (not A299) );
 a31541a <=( (not A266)  and  a31540a );
 a31542a <=( a31541a  and  a31536a );
 a31546a <=( A167  and  A169 );
 a31547a <=( (not A170)  and  a31546a );
 a31551a <=( (not A201)  and  (not A200) );
 a31552a <=( A166  and  a31551a );
 a31553a <=( a31552a  and  a31547a );
 a31557a <=( (not A265)  and  A233 );
 a31558a <=( A232  and  a31557a );
 a31562a <=( A299  and  A298 );
 a31563a <=( (not A266)  and  a31562a );
 a31564a <=( a31563a  and  a31558a );
 a31568a <=( A167  and  A169 );
 a31569a <=( (not A170)  and  a31568a );
 a31573a <=( (not A201)  and  (not A200) );
 a31574a <=( A166  and  a31573a );
 a31575a <=( a31574a  and  a31569a );
 a31579a <=( (not A265)  and  A233 );
 a31580a <=( A232  and  a31579a );
 a31584a <=( (not A299)  and  (not A298) );
 a31585a <=( (not A266)  and  a31584a );
 a31586a <=( a31585a  and  a31580a );
 a31590a <=( A167  and  A169 );
 a31591a <=( (not A170)  and  a31590a );
 a31595a <=( (not A201)  and  (not A200) );
 a31596a <=( A166  and  a31595a );
 a31597a <=( a31596a  and  a31591a );
 a31601a <=( A298  and  A233 );
 a31602a <=( (not A232)  and  a31601a );
 a31606a <=( A301  and  A300 );
 a31607a <=( (not A299)  and  a31606a );
 a31608a <=( a31607a  and  a31602a );
 a31612a <=( A167  and  A169 );
 a31613a <=( (not A170)  and  a31612a );
 a31617a <=( (not A201)  and  (not A200) );
 a31618a <=( A166  and  a31617a );
 a31619a <=( a31618a  and  a31613a );
 a31623a <=( A298  and  A233 );
 a31624a <=( (not A232)  and  a31623a );
 a31628a <=( A302  and  A300 );
 a31629a <=( (not A299)  and  a31628a );
 a31630a <=( a31629a  and  a31624a );
 a31634a <=( A167  and  A169 );
 a31635a <=( (not A170)  and  a31634a );
 a31639a <=( (not A201)  and  (not A200) );
 a31640a <=( A166  and  a31639a );
 a31641a <=( a31640a  and  a31635a );
 a31645a <=( A265  and  A233 );
 a31646a <=( (not A232)  and  a31645a );
 a31650a <=( A268  and  A267 );
 a31651a <=( (not A266)  and  a31650a );
 a31652a <=( a31651a  and  a31646a );
 a31656a <=( A167  and  A169 );
 a31657a <=( (not A170)  and  a31656a );
 a31661a <=( (not A201)  and  (not A200) );
 a31662a <=( A166  and  a31661a );
 a31663a <=( a31662a  and  a31657a );
 a31667a <=( A265  and  A233 );
 a31668a <=( (not A232)  and  a31667a );
 a31672a <=( A269  and  A267 );
 a31673a <=( (not A266)  and  a31672a );
 a31674a <=( a31673a  and  a31668a );
 a31678a <=( A167  and  A169 );
 a31679a <=( (not A170)  and  a31678a );
 a31683a <=( (not A201)  and  (not A200) );
 a31684a <=( A166  and  a31683a );
 a31685a <=( a31684a  and  a31679a );
 a31689a <=( A265  and  (not A234) );
 a31690a <=( (not A233)  and  a31689a );
 a31694a <=( (not A300)  and  A298 );
 a31695a <=( A266  and  a31694a );
 a31696a <=( a31695a  and  a31690a );
 a31700a <=( A167  and  A169 );
 a31701a <=( (not A170)  and  a31700a );
 a31705a <=( (not A201)  and  (not A200) );
 a31706a <=( A166  and  a31705a );
 a31707a <=( a31706a  and  a31701a );
 a31711a <=( A265  and  (not A234) );
 a31712a <=( (not A233)  and  a31711a );
 a31716a <=( A299  and  A298 );
 a31717a <=( A266  and  a31716a );
 a31718a <=( a31717a  and  a31712a );
 a31722a <=( A167  and  A169 );
 a31723a <=( (not A170)  and  a31722a );
 a31727a <=( (not A201)  and  (not A200) );
 a31728a <=( A166  and  a31727a );
 a31729a <=( a31728a  and  a31723a );
 a31733a <=( A265  and  (not A234) );
 a31734a <=( (not A233)  and  a31733a );
 a31738a <=( (not A299)  and  (not A298) );
 a31739a <=( A266  and  a31738a );
 a31740a <=( a31739a  and  a31734a );
 a31744a <=( A167  and  A169 );
 a31745a <=( (not A170)  and  a31744a );
 a31749a <=( (not A201)  and  (not A200) );
 a31750a <=( A166  and  a31749a );
 a31751a <=( a31750a  and  a31745a );
 a31755a <=( (not A266)  and  (not A234) );
 a31756a <=( (not A233)  and  a31755a );
 a31760a <=( (not A300)  and  A298 );
 a31761a <=( (not A267)  and  a31760a );
 a31762a <=( a31761a  and  a31756a );
 a31766a <=( A167  and  A169 );
 a31767a <=( (not A170)  and  a31766a );
 a31771a <=( (not A201)  and  (not A200) );
 a31772a <=( A166  and  a31771a );
 a31773a <=( a31772a  and  a31767a );
 a31777a <=( (not A266)  and  (not A234) );
 a31778a <=( (not A233)  and  a31777a );
 a31782a <=( A299  and  A298 );
 a31783a <=( (not A267)  and  a31782a );
 a31784a <=( a31783a  and  a31778a );
 a31788a <=( A167  and  A169 );
 a31789a <=( (not A170)  and  a31788a );
 a31793a <=( (not A201)  and  (not A200) );
 a31794a <=( A166  and  a31793a );
 a31795a <=( a31794a  and  a31789a );
 a31799a <=( (not A266)  and  (not A234) );
 a31800a <=( (not A233)  and  a31799a );
 a31804a <=( (not A299)  and  (not A298) );
 a31805a <=( (not A267)  and  a31804a );
 a31806a <=( a31805a  and  a31800a );
 a31810a <=( A167  and  A169 );
 a31811a <=( (not A170)  and  a31810a );
 a31815a <=( (not A201)  and  (not A200) );
 a31816a <=( A166  and  a31815a );
 a31817a <=( a31816a  and  a31811a );
 a31821a <=( (not A265)  and  (not A234) );
 a31822a <=( (not A233)  and  a31821a );
 a31826a <=( (not A300)  and  A298 );
 a31827a <=( (not A266)  and  a31826a );
 a31828a <=( a31827a  and  a31822a );
 a31832a <=( A167  and  A169 );
 a31833a <=( (not A170)  and  a31832a );
 a31837a <=( (not A201)  and  (not A200) );
 a31838a <=( A166  and  a31837a );
 a31839a <=( a31838a  and  a31833a );
 a31843a <=( (not A265)  and  (not A234) );
 a31844a <=( (not A233)  and  a31843a );
 a31848a <=( A299  and  A298 );
 a31849a <=( (not A266)  and  a31848a );
 a31850a <=( a31849a  and  a31844a );
 a31854a <=( A167  and  A169 );
 a31855a <=( (not A170)  and  a31854a );
 a31859a <=( (not A201)  and  (not A200) );
 a31860a <=( A166  and  a31859a );
 a31861a <=( a31860a  and  a31855a );
 a31865a <=( (not A265)  and  (not A234) );
 a31866a <=( (not A233)  and  a31865a );
 a31870a <=( (not A299)  and  (not A298) );
 a31871a <=( (not A266)  and  a31870a );
 a31872a <=( a31871a  and  a31866a );
 a31876a <=( A167  and  A169 );
 a31877a <=( (not A170)  and  a31876a );
 a31881a <=( (not A201)  and  (not A200) );
 a31882a <=( A166  and  a31881a );
 a31883a <=( a31882a  and  a31877a );
 a31887a <=( A234  and  (not A233) );
 a31888a <=( A232  and  a31887a );
 a31892a <=( A299  and  (not A298) );
 a31893a <=( A235  and  a31892a );
 a31894a <=( a31893a  and  a31888a );
 a31898a <=( A167  and  A169 );
 a31899a <=( (not A170)  and  a31898a );
 a31903a <=( (not A201)  and  (not A200) );
 a31904a <=( A166  and  a31903a );
 a31905a <=( a31904a  and  a31899a );
 a31909a <=( A234  and  (not A233) );
 a31910a <=( A232  and  a31909a );
 a31914a <=( A266  and  (not A265) );
 a31915a <=( A235  and  a31914a );
 a31916a <=( a31915a  and  a31910a );
 a31920a <=( A167  and  A169 );
 a31921a <=( (not A170)  and  a31920a );
 a31925a <=( (not A201)  and  (not A200) );
 a31926a <=( A166  and  a31925a );
 a31927a <=( a31926a  and  a31921a );
 a31931a <=( A234  and  (not A233) );
 a31932a <=( A232  and  a31931a );
 a31936a <=( A299  and  (not A298) );
 a31937a <=( A236  and  a31936a );
 a31938a <=( a31937a  and  a31932a );
 a31942a <=( A167  and  A169 );
 a31943a <=( (not A170)  and  a31942a );
 a31947a <=( (not A201)  and  (not A200) );
 a31948a <=( A166  and  a31947a );
 a31949a <=( a31948a  and  a31943a );
 a31953a <=( A234  and  (not A233) );
 a31954a <=( A232  and  a31953a );
 a31958a <=( A266  and  (not A265) );
 a31959a <=( A236  and  a31958a );
 a31960a <=( a31959a  and  a31954a );
 a31964a <=( A167  and  A169 );
 a31965a <=( (not A170)  and  a31964a );
 a31969a <=( (not A201)  and  (not A200) );
 a31970a <=( A166  and  a31969a );
 a31971a <=( a31970a  and  a31965a );
 a31975a <=( A265  and  (not A233) );
 a31976a <=( (not A232)  and  a31975a );
 a31980a <=( (not A300)  and  A298 );
 a31981a <=( A266  and  a31980a );
 a31982a <=( a31981a  and  a31976a );
 a31986a <=( A167  and  A169 );
 a31987a <=( (not A170)  and  a31986a );
 a31991a <=( (not A201)  and  (not A200) );
 a31992a <=( A166  and  a31991a );
 a31993a <=( a31992a  and  a31987a );
 a31997a <=( A265  and  (not A233) );
 a31998a <=( (not A232)  and  a31997a );
 a32002a <=( A299  and  A298 );
 a32003a <=( A266  and  a32002a );
 a32004a <=( a32003a  and  a31998a );
 a32008a <=( A167  and  A169 );
 a32009a <=( (not A170)  and  a32008a );
 a32013a <=( (not A201)  and  (not A200) );
 a32014a <=( A166  and  a32013a );
 a32015a <=( a32014a  and  a32009a );
 a32019a <=( A265  and  (not A233) );
 a32020a <=( (not A232)  and  a32019a );
 a32024a <=( (not A299)  and  (not A298) );
 a32025a <=( A266  and  a32024a );
 a32026a <=( a32025a  and  a32020a );
 a32030a <=( A167  and  A169 );
 a32031a <=( (not A170)  and  a32030a );
 a32035a <=( (not A201)  and  (not A200) );
 a32036a <=( A166  and  a32035a );
 a32037a <=( a32036a  and  a32031a );
 a32041a <=( (not A266)  and  (not A233) );
 a32042a <=( (not A232)  and  a32041a );
 a32046a <=( (not A300)  and  A298 );
 a32047a <=( (not A267)  and  a32046a );
 a32048a <=( a32047a  and  a32042a );
 a32052a <=( A167  and  A169 );
 a32053a <=( (not A170)  and  a32052a );
 a32057a <=( (not A201)  and  (not A200) );
 a32058a <=( A166  and  a32057a );
 a32059a <=( a32058a  and  a32053a );
 a32063a <=( (not A266)  and  (not A233) );
 a32064a <=( (not A232)  and  a32063a );
 a32068a <=( A299  and  A298 );
 a32069a <=( (not A267)  and  a32068a );
 a32070a <=( a32069a  and  a32064a );
 a32074a <=( A167  and  A169 );
 a32075a <=( (not A170)  and  a32074a );
 a32079a <=( (not A201)  and  (not A200) );
 a32080a <=( A166  and  a32079a );
 a32081a <=( a32080a  and  a32075a );
 a32085a <=( (not A266)  and  (not A233) );
 a32086a <=( (not A232)  and  a32085a );
 a32090a <=( (not A299)  and  (not A298) );
 a32091a <=( (not A267)  and  a32090a );
 a32092a <=( a32091a  and  a32086a );
 a32096a <=( A167  and  A169 );
 a32097a <=( (not A170)  and  a32096a );
 a32101a <=( (not A201)  and  (not A200) );
 a32102a <=( A166  and  a32101a );
 a32103a <=( a32102a  and  a32097a );
 a32107a <=( (not A265)  and  (not A233) );
 a32108a <=( (not A232)  and  a32107a );
 a32112a <=( (not A300)  and  A298 );
 a32113a <=( (not A266)  and  a32112a );
 a32114a <=( a32113a  and  a32108a );
 a32118a <=( A167  and  A169 );
 a32119a <=( (not A170)  and  a32118a );
 a32123a <=( (not A201)  and  (not A200) );
 a32124a <=( A166  and  a32123a );
 a32125a <=( a32124a  and  a32119a );
 a32129a <=( (not A265)  and  (not A233) );
 a32130a <=( (not A232)  and  a32129a );
 a32134a <=( A299  and  A298 );
 a32135a <=( (not A266)  and  a32134a );
 a32136a <=( a32135a  and  a32130a );
 a32140a <=( A167  and  A169 );
 a32141a <=( (not A170)  and  a32140a );
 a32145a <=( (not A201)  and  (not A200) );
 a32146a <=( A166  and  a32145a );
 a32147a <=( a32146a  and  a32141a );
 a32151a <=( (not A265)  and  (not A233) );
 a32152a <=( (not A232)  and  a32151a );
 a32156a <=( (not A299)  and  (not A298) );
 a32157a <=( (not A266)  and  a32156a );
 a32158a <=( a32157a  and  a32152a );
 a32162a <=( A167  and  A169 );
 a32163a <=( (not A170)  and  a32162a );
 a32167a <=( (not A200)  and  (not A199) );
 a32168a <=( A166  and  a32167a );
 a32169a <=( a32168a  and  a32163a );
 a32173a <=( A265  and  A233 );
 a32174a <=( A232  and  a32173a );
 a32178a <=( (not A300)  and  (not A299) );
 a32179a <=( (not A267)  and  a32178a );
 a32180a <=( a32179a  and  a32174a );
 a32184a <=( A167  and  A169 );
 a32185a <=( (not A170)  and  a32184a );
 a32189a <=( (not A200)  and  (not A199) );
 a32190a <=( A166  and  a32189a );
 a32191a <=( a32190a  and  a32185a );
 a32195a <=( A265  and  A233 );
 a32196a <=( A232  and  a32195a );
 a32200a <=( A299  and  A298 );
 a32201a <=( (not A267)  and  a32200a );
 a32202a <=( a32201a  and  a32196a );
 a32206a <=( A167  and  A169 );
 a32207a <=( (not A170)  and  a32206a );
 a32211a <=( (not A200)  and  (not A199) );
 a32212a <=( A166  and  a32211a );
 a32213a <=( a32212a  and  a32207a );
 a32217a <=( A265  and  A233 );
 a32218a <=( A232  and  a32217a );
 a32222a <=( (not A299)  and  (not A298) );
 a32223a <=( (not A267)  and  a32222a );
 a32224a <=( a32223a  and  a32218a );
 a32228a <=( A167  and  A169 );
 a32229a <=( (not A170)  and  a32228a );
 a32233a <=( (not A200)  and  (not A199) );
 a32234a <=( A166  and  a32233a );
 a32235a <=( a32234a  and  a32229a );
 a32239a <=( A265  and  A233 );
 a32240a <=( A232  and  a32239a );
 a32244a <=( (not A300)  and  (not A299) );
 a32245a <=( A266  and  a32244a );
 a32246a <=( a32245a  and  a32240a );
 a32250a <=( A167  and  A169 );
 a32251a <=( (not A170)  and  a32250a );
 a32255a <=( (not A200)  and  (not A199) );
 a32256a <=( A166  and  a32255a );
 a32257a <=( a32256a  and  a32251a );
 a32261a <=( A265  and  A233 );
 a32262a <=( A232  and  a32261a );
 a32266a <=( A299  and  A298 );
 a32267a <=( A266  and  a32266a );
 a32268a <=( a32267a  and  a32262a );
 a32272a <=( A167  and  A169 );
 a32273a <=( (not A170)  and  a32272a );
 a32277a <=( (not A200)  and  (not A199) );
 a32278a <=( A166  and  a32277a );
 a32279a <=( a32278a  and  a32273a );
 a32283a <=( A265  and  A233 );
 a32284a <=( A232  and  a32283a );
 a32288a <=( (not A299)  and  (not A298) );
 a32289a <=( A266  and  a32288a );
 a32290a <=( a32289a  and  a32284a );
 a32294a <=( A167  and  A169 );
 a32295a <=( (not A170)  and  a32294a );
 a32299a <=( (not A200)  and  (not A199) );
 a32300a <=( A166  and  a32299a );
 a32301a <=( a32300a  and  a32295a );
 a32305a <=( (not A265)  and  A233 );
 a32306a <=( A232  and  a32305a );
 a32310a <=( (not A300)  and  (not A299) );
 a32311a <=( (not A266)  and  a32310a );
 a32312a <=( a32311a  and  a32306a );
 a32316a <=( A167  and  A169 );
 a32317a <=( (not A170)  and  a32316a );
 a32321a <=( (not A200)  and  (not A199) );
 a32322a <=( A166  and  a32321a );
 a32323a <=( a32322a  and  a32317a );
 a32327a <=( (not A265)  and  A233 );
 a32328a <=( A232  and  a32327a );
 a32332a <=( A299  and  A298 );
 a32333a <=( (not A266)  and  a32332a );
 a32334a <=( a32333a  and  a32328a );
 a32338a <=( A167  and  A169 );
 a32339a <=( (not A170)  and  a32338a );
 a32343a <=( (not A200)  and  (not A199) );
 a32344a <=( A166  and  a32343a );
 a32345a <=( a32344a  and  a32339a );
 a32349a <=( (not A265)  and  A233 );
 a32350a <=( A232  and  a32349a );
 a32354a <=( (not A299)  and  (not A298) );
 a32355a <=( (not A266)  and  a32354a );
 a32356a <=( a32355a  and  a32350a );
 a32360a <=( A167  and  A169 );
 a32361a <=( (not A170)  and  a32360a );
 a32365a <=( (not A200)  and  (not A199) );
 a32366a <=( A166  and  a32365a );
 a32367a <=( a32366a  and  a32361a );
 a32371a <=( A298  and  A233 );
 a32372a <=( (not A232)  and  a32371a );
 a32376a <=( A301  and  A300 );
 a32377a <=( (not A299)  and  a32376a );
 a32378a <=( a32377a  and  a32372a );
 a32382a <=( A167  and  A169 );
 a32383a <=( (not A170)  and  a32382a );
 a32387a <=( (not A200)  and  (not A199) );
 a32388a <=( A166  and  a32387a );
 a32389a <=( a32388a  and  a32383a );
 a32393a <=( A298  and  A233 );
 a32394a <=( (not A232)  and  a32393a );
 a32398a <=( A302  and  A300 );
 a32399a <=( (not A299)  and  a32398a );
 a32400a <=( a32399a  and  a32394a );
 a32404a <=( A167  and  A169 );
 a32405a <=( (not A170)  and  a32404a );
 a32409a <=( (not A200)  and  (not A199) );
 a32410a <=( A166  and  a32409a );
 a32411a <=( a32410a  and  a32405a );
 a32415a <=( A265  and  A233 );
 a32416a <=( (not A232)  and  a32415a );
 a32420a <=( A268  and  A267 );
 a32421a <=( (not A266)  and  a32420a );
 a32422a <=( a32421a  and  a32416a );
 a32426a <=( A167  and  A169 );
 a32427a <=( (not A170)  and  a32426a );
 a32431a <=( (not A200)  and  (not A199) );
 a32432a <=( A166  and  a32431a );
 a32433a <=( a32432a  and  a32427a );
 a32437a <=( A265  and  A233 );
 a32438a <=( (not A232)  and  a32437a );
 a32442a <=( A269  and  A267 );
 a32443a <=( (not A266)  and  a32442a );
 a32444a <=( a32443a  and  a32438a );
 a32448a <=( A167  and  A169 );
 a32449a <=( (not A170)  and  a32448a );
 a32453a <=( (not A200)  and  (not A199) );
 a32454a <=( A166  and  a32453a );
 a32455a <=( a32454a  and  a32449a );
 a32459a <=( A265  and  (not A234) );
 a32460a <=( (not A233)  and  a32459a );
 a32464a <=( (not A300)  and  A298 );
 a32465a <=( A266  and  a32464a );
 a32466a <=( a32465a  and  a32460a );
 a32470a <=( A167  and  A169 );
 a32471a <=( (not A170)  and  a32470a );
 a32475a <=( (not A200)  and  (not A199) );
 a32476a <=( A166  and  a32475a );
 a32477a <=( a32476a  and  a32471a );
 a32481a <=( A265  and  (not A234) );
 a32482a <=( (not A233)  and  a32481a );
 a32486a <=( A299  and  A298 );
 a32487a <=( A266  and  a32486a );
 a32488a <=( a32487a  and  a32482a );
 a32492a <=( A167  and  A169 );
 a32493a <=( (not A170)  and  a32492a );
 a32497a <=( (not A200)  and  (not A199) );
 a32498a <=( A166  and  a32497a );
 a32499a <=( a32498a  and  a32493a );
 a32503a <=( A265  and  (not A234) );
 a32504a <=( (not A233)  and  a32503a );
 a32508a <=( (not A299)  and  (not A298) );
 a32509a <=( A266  and  a32508a );
 a32510a <=( a32509a  and  a32504a );
 a32514a <=( A167  and  A169 );
 a32515a <=( (not A170)  and  a32514a );
 a32519a <=( (not A200)  and  (not A199) );
 a32520a <=( A166  and  a32519a );
 a32521a <=( a32520a  and  a32515a );
 a32525a <=( (not A266)  and  (not A234) );
 a32526a <=( (not A233)  and  a32525a );
 a32530a <=( (not A300)  and  A298 );
 a32531a <=( (not A267)  and  a32530a );
 a32532a <=( a32531a  and  a32526a );
 a32536a <=( A167  and  A169 );
 a32537a <=( (not A170)  and  a32536a );
 a32541a <=( (not A200)  and  (not A199) );
 a32542a <=( A166  and  a32541a );
 a32543a <=( a32542a  and  a32537a );
 a32547a <=( (not A266)  and  (not A234) );
 a32548a <=( (not A233)  and  a32547a );
 a32552a <=( A299  and  A298 );
 a32553a <=( (not A267)  and  a32552a );
 a32554a <=( a32553a  and  a32548a );
 a32558a <=( A167  and  A169 );
 a32559a <=( (not A170)  and  a32558a );
 a32563a <=( (not A200)  and  (not A199) );
 a32564a <=( A166  and  a32563a );
 a32565a <=( a32564a  and  a32559a );
 a32569a <=( (not A266)  and  (not A234) );
 a32570a <=( (not A233)  and  a32569a );
 a32574a <=( (not A299)  and  (not A298) );
 a32575a <=( (not A267)  and  a32574a );
 a32576a <=( a32575a  and  a32570a );
 a32580a <=( A167  and  A169 );
 a32581a <=( (not A170)  and  a32580a );
 a32585a <=( (not A200)  and  (not A199) );
 a32586a <=( A166  and  a32585a );
 a32587a <=( a32586a  and  a32581a );
 a32591a <=( (not A265)  and  (not A234) );
 a32592a <=( (not A233)  and  a32591a );
 a32596a <=( (not A300)  and  A298 );
 a32597a <=( (not A266)  and  a32596a );
 a32598a <=( a32597a  and  a32592a );
 a32602a <=( A167  and  A169 );
 a32603a <=( (not A170)  and  a32602a );
 a32607a <=( (not A200)  and  (not A199) );
 a32608a <=( A166  and  a32607a );
 a32609a <=( a32608a  and  a32603a );
 a32613a <=( (not A265)  and  (not A234) );
 a32614a <=( (not A233)  and  a32613a );
 a32618a <=( A299  and  A298 );
 a32619a <=( (not A266)  and  a32618a );
 a32620a <=( a32619a  and  a32614a );
 a32624a <=( A167  and  A169 );
 a32625a <=( (not A170)  and  a32624a );
 a32629a <=( (not A200)  and  (not A199) );
 a32630a <=( A166  and  a32629a );
 a32631a <=( a32630a  and  a32625a );
 a32635a <=( (not A265)  and  (not A234) );
 a32636a <=( (not A233)  and  a32635a );
 a32640a <=( (not A299)  and  (not A298) );
 a32641a <=( (not A266)  and  a32640a );
 a32642a <=( a32641a  and  a32636a );
 a32646a <=( A167  and  A169 );
 a32647a <=( (not A170)  and  a32646a );
 a32651a <=( (not A200)  and  (not A199) );
 a32652a <=( A166  and  a32651a );
 a32653a <=( a32652a  and  a32647a );
 a32657a <=( A234  and  (not A233) );
 a32658a <=( A232  and  a32657a );
 a32662a <=( A299  and  (not A298) );
 a32663a <=( A235  and  a32662a );
 a32664a <=( a32663a  and  a32658a );
 a32668a <=( A167  and  A169 );
 a32669a <=( (not A170)  and  a32668a );
 a32673a <=( (not A200)  and  (not A199) );
 a32674a <=( A166  and  a32673a );
 a32675a <=( a32674a  and  a32669a );
 a32679a <=( A234  and  (not A233) );
 a32680a <=( A232  and  a32679a );
 a32684a <=( A266  and  (not A265) );
 a32685a <=( A235  and  a32684a );
 a32686a <=( a32685a  and  a32680a );
 a32690a <=( A167  and  A169 );
 a32691a <=( (not A170)  and  a32690a );
 a32695a <=( (not A200)  and  (not A199) );
 a32696a <=( A166  and  a32695a );
 a32697a <=( a32696a  and  a32691a );
 a32701a <=( A234  and  (not A233) );
 a32702a <=( A232  and  a32701a );
 a32706a <=( A299  and  (not A298) );
 a32707a <=( A236  and  a32706a );
 a32708a <=( a32707a  and  a32702a );
 a32712a <=( A167  and  A169 );
 a32713a <=( (not A170)  and  a32712a );
 a32717a <=( (not A200)  and  (not A199) );
 a32718a <=( A166  and  a32717a );
 a32719a <=( a32718a  and  a32713a );
 a32723a <=( A234  and  (not A233) );
 a32724a <=( A232  and  a32723a );
 a32728a <=( A266  and  (not A265) );
 a32729a <=( A236  and  a32728a );
 a32730a <=( a32729a  and  a32724a );
 a32734a <=( A167  and  A169 );
 a32735a <=( (not A170)  and  a32734a );
 a32739a <=( (not A200)  and  (not A199) );
 a32740a <=( A166  and  a32739a );
 a32741a <=( a32740a  and  a32735a );
 a32745a <=( A265  and  (not A233) );
 a32746a <=( (not A232)  and  a32745a );
 a32750a <=( (not A300)  and  A298 );
 a32751a <=( A266  and  a32750a );
 a32752a <=( a32751a  and  a32746a );
 a32756a <=( A167  and  A169 );
 a32757a <=( (not A170)  and  a32756a );
 a32761a <=( (not A200)  and  (not A199) );
 a32762a <=( A166  and  a32761a );
 a32763a <=( a32762a  and  a32757a );
 a32767a <=( A265  and  (not A233) );
 a32768a <=( (not A232)  and  a32767a );
 a32772a <=( A299  and  A298 );
 a32773a <=( A266  and  a32772a );
 a32774a <=( a32773a  and  a32768a );
 a32778a <=( A167  and  A169 );
 a32779a <=( (not A170)  and  a32778a );
 a32783a <=( (not A200)  and  (not A199) );
 a32784a <=( A166  and  a32783a );
 a32785a <=( a32784a  and  a32779a );
 a32789a <=( A265  and  (not A233) );
 a32790a <=( (not A232)  and  a32789a );
 a32794a <=( (not A299)  and  (not A298) );
 a32795a <=( A266  and  a32794a );
 a32796a <=( a32795a  and  a32790a );
 a32800a <=( A167  and  A169 );
 a32801a <=( (not A170)  and  a32800a );
 a32805a <=( (not A200)  and  (not A199) );
 a32806a <=( A166  and  a32805a );
 a32807a <=( a32806a  and  a32801a );
 a32811a <=( (not A266)  and  (not A233) );
 a32812a <=( (not A232)  and  a32811a );
 a32816a <=( (not A300)  and  A298 );
 a32817a <=( (not A267)  and  a32816a );
 a32818a <=( a32817a  and  a32812a );
 a32822a <=( A167  and  A169 );
 a32823a <=( (not A170)  and  a32822a );
 a32827a <=( (not A200)  and  (not A199) );
 a32828a <=( A166  and  a32827a );
 a32829a <=( a32828a  and  a32823a );
 a32833a <=( (not A266)  and  (not A233) );
 a32834a <=( (not A232)  and  a32833a );
 a32838a <=( A299  and  A298 );
 a32839a <=( (not A267)  and  a32838a );
 a32840a <=( a32839a  and  a32834a );
 a32844a <=( A167  and  A169 );
 a32845a <=( (not A170)  and  a32844a );
 a32849a <=( (not A200)  and  (not A199) );
 a32850a <=( A166  and  a32849a );
 a32851a <=( a32850a  and  a32845a );
 a32855a <=( (not A266)  and  (not A233) );
 a32856a <=( (not A232)  and  a32855a );
 a32860a <=( (not A299)  and  (not A298) );
 a32861a <=( (not A267)  and  a32860a );
 a32862a <=( a32861a  and  a32856a );
 a32866a <=( A167  and  A169 );
 a32867a <=( (not A170)  and  a32866a );
 a32871a <=( (not A200)  and  (not A199) );
 a32872a <=( A166  and  a32871a );
 a32873a <=( a32872a  and  a32867a );
 a32877a <=( (not A265)  and  (not A233) );
 a32878a <=( (not A232)  and  a32877a );
 a32882a <=( (not A300)  and  A298 );
 a32883a <=( (not A266)  and  a32882a );
 a32884a <=( a32883a  and  a32878a );
 a32888a <=( A167  and  A169 );
 a32889a <=( (not A170)  and  a32888a );
 a32893a <=( (not A200)  and  (not A199) );
 a32894a <=( A166  and  a32893a );
 a32895a <=( a32894a  and  a32889a );
 a32899a <=( (not A265)  and  (not A233) );
 a32900a <=( (not A232)  and  a32899a );
 a32904a <=( A299  and  A298 );
 a32905a <=( (not A266)  and  a32904a );
 a32906a <=( a32905a  and  a32900a );
 a32910a <=( A167  and  A169 );
 a32911a <=( (not A170)  and  a32910a );
 a32915a <=( (not A200)  and  (not A199) );
 a32916a <=( A166  and  a32915a );
 a32917a <=( a32916a  and  a32911a );
 a32921a <=( (not A265)  and  (not A233) );
 a32922a <=( (not A232)  and  a32921a );
 a32926a <=( (not A299)  and  (not A298) );
 a32927a <=( (not A266)  and  a32926a );
 a32928a <=( a32927a  and  a32922a );
 a32932a <=( (not A167)  and  A169 );
 a32933a <=( (not A170)  and  a32932a );
 a32937a <=( A200  and  A199 );
 a32938a <=( (not A166)  and  a32937a );
 a32939a <=( a32938a  and  a32933a );
 a32943a <=( A265  and  A233 );
 a32944a <=( A232  and  a32943a );
 a32948a <=( (not A300)  and  (not A299) );
 a32949a <=( (not A267)  and  a32948a );
 a32950a <=( a32949a  and  a32944a );
 a32954a <=( (not A167)  and  A169 );
 a32955a <=( (not A170)  and  a32954a );
 a32959a <=( A200  and  A199 );
 a32960a <=( (not A166)  and  a32959a );
 a32961a <=( a32960a  and  a32955a );
 a32965a <=( A265  and  A233 );
 a32966a <=( A232  and  a32965a );
 a32970a <=( A299  and  A298 );
 a32971a <=( (not A267)  and  a32970a );
 a32972a <=( a32971a  and  a32966a );
 a32976a <=( (not A167)  and  A169 );
 a32977a <=( (not A170)  and  a32976a );
 a32981a <=( A200  and  A199 );
 a32982a <=( (not A166)  and  a32981a );
 a32983a <=( a32982a  and  a32977a );
 a32987a <=( A265  and  A233 );
 a32988a <=( A232  and  a32987a );
 a32992a <=( (not A299)  and  (not A298) );
 a32993a <=( (not A267)  and  a32992a );
 a32994a <=( a32993a  and  a32988a );
 a32998a <=( (not A167)  and  A169 );
 a32999a <=( (not A170)  and  a32998a );
 a33003a <=( A200  and  A199 );
 a33004a <=( (not A166)  and  a33003a );
 a33005a <=( a33004a  and  a32999a );
 a33009a <=( A265  and  A233 );
 a33010a <=( A232  and  a33009a );
 a33014a <=( (not A300)  and  (not A299) );
 a33015a <=( A266  and  a33014a );
 a33016a <=( a33015a  and  a33010a );
 a33020a <=( (not A167)  and  A169 );
 a33021a <=( (not A170)  and  a33020a );
 a33025a <=( A200  and  A199 );
 a33026a <=( (not A166)  and  a33025a );
 a33027a <=( a33026a  and  a33021a );
 a33031a <=( A265  and  A233 );
 a33032a <=( A232  and  a33031a );
 a33036a <=( A299  and  A298 );
 a33037a <=( A266  and  a33036a );
 a33038a <=( a33037a  and  a33032a );
 a33042a <=( (not A167)  and  A169 );
 a33043a <=( (not A170)  and  a33042a );
 a33047a <=( A200  and  A199 );
 a33048a <=( (not A166)  and  a33047a );
 a33049a <=( a33048a  and  a33043a );
 a33053a <=( A265  and  A233 );
 a33054a <=( A232  and  a33053a );
 a33058a <=( (not A299)  and  (not A298) );
 a33059a <=( A266  and  a33058a );
 a33060a <=( a33059a  and  a33054a );
 a33064a <=( (not A167)  and  A169 );
 a33065a <=( (not A170)  and  a33064a );
 a33069a <=( A200  and  A199 );
 a33070a <=( (not A166)  and  a33069a );
 a33071a <=( a33070a  and  a33065a );
 a33075a <=( (not A265)  and  A233 );
 a33076a <=( A232  and  a33075a );
 a33080a <=( (not A300)  and  (not A299) );
 a33081a <=( (not A266)  and  a33080a );
 a33082a <=( a33081a  and  a33076a );
 a33086a <=( (not A167)  and  A169 );
 a33087a <=( (not A170)  and  a33086a );
 a33091a <=( A200  and  A199 );
 a33092a <=( (not A166)  and  a33091a );
 a33093a <=( a33092a  and  a33087a );
 a33097a <=( (not A265)  and  A233 );
 a33098a <=( A232  and  a33097a );
 a33102a <=( A299  and  A298 );
 a33103a <=( (not A266)  and  a33102a );
 a33104a <=( a33103a  and  a33098a );
 a33108a <=( (not A167)  and  A169 );
 a33109a <=( (not A170)  and  a33108a );
 a33113a <=( A200  and  A199 );
 a33114a <=( (not A166)  and  a33113a );
 a33115a <=( a33114a  and  a33109a );
 a33119a <=( (not A265)  and  A233 );
 a33120a <=( A232  and  a33119a );
 a33124a <=( (not A299)  and  (not A298) );
 a33125a <=( (not A266)  and  a33124a );
 a33126a <=( a33125a  and  a33120a );
 a33130a <=( (not A167)  and  A169 );
 a33131a <=( (not A170)  and  a33130a );
 a33135a <=( A200  and  A199 );
 a33136a <=( (not A166)  and  a33135a );
 a33137a <=( a33136a  and  a33131a );
 a33141a <=( A298  and  A233 );
 a33142a <=( (not A232)  and  a33141a );
 a33146a <=( A301  and  A300 );
 a33147a <=( (not A299)  and  a33146a );
 a33148a <=( a33147a  and  a33142a );
 a33152a <=( (not A167)  and  A169 );
 a33153a <=( (not A170)  and  a33152a );
 a33157a <=( A200  and  A199 );
 a33158a <=( (not A166)  and  a33157a );
 a33159a <=( a33158a  and  a33153a );
 a33163a <=( A298  and  A233 );
 a33164a <=( (not A232)  and  a33163a );
 a33168a <=( A302  and  A300 );
 a33169a <=( (not A299)  and  a33168a );
 a33170a <=( a33169a  and  a33164a );
 a33174a <=( (not A167)  and  A169 );
 a33175a <=( (not A170)  and  a33174a );
 a33179a <=( A200  and  A199 );
 a33180a <=( (not A166)  and  a33179a );
 a33181a <=( a33180a  and  a33175a );
 a33185a <=( A265  and  A233 );
 a33186a <=( (not A232)  and  a33185a );
 a33190a <=( A268  and  A267 );
 a33191a <=( (not A266)  and  a33190a );
 a33192a <=( a33191a  and  a33186a );
 a33196a <=( (not A167)  and  A169 );
 a33197a <=( (not A170)  and  a33196a );
 a33201a <=( A200  and  A199 );
 a33202a <=( (not A166)  and  a33201a );
 a33203a <=( a33202a  and  a33197a );
 a33207a <=( A265  and  A233 );
 a33208a <=( (not A232)  and  a33207a );
 a33212a <=( A269  and  A267 );
 a33213a <=( (not A266)  and  a33212a );
 a33214a <=( a33213a  and  a33208a );
 a33218a <=( (not A167)  and  A169 );
 a33219a <=( (not A170)  and  a33218a );
 a33223a <=( A200  and  A199 );
 a33224a <=( (not A166)  and  a33223a );
 a33225a <=( a33224a  and  a33219a );
 a33229a <=( A265  and  (not A234) );
 a33230a <=( (not A233)  and  a33229a );
 a33234a <=( (not A300)  and  A298 );
 a33235a <=( A266  and  a33234a );
 a33236a <=( a33235a  and  a33230a );
 a33240a <=( (not A167)  and  A169 );
 a33241a <=( (not A170)  and  a33240a );
 a33245a <=( A200  and  A199 );
 a33246a <=( (not A166)  and  a33245a );
 a33247a <=( a33246a  and  a33241a );
 a33251a <=( A265  and  (not A234) );
 a33252a <=( (not A233)  and  a33251a );
 a33256a <=( A299  and  A298 );
 a33257a <=( A266  and  a33256a );
 a33258a <=( a33257a  and  a33252a );
 a33262a <=( (not A167)  and  A169 );
 a33263a <=( (not A170)  and  a33262a );
 a33267a <=( A200  and  A199 );
 a33268a <=( (not A166)  and  a33267a );
 a33269a <=( a33268a  and  a33263a );
 a33273a <=( A265  and  (not A234) );
 a33274a <=( (not A233)  and  a33273a );
 a33278a <=( (not A299)  and  (not A298) );
 a33279a <=( A266  and  a33278a );
 a33280a <=( a33279a  and  a33274a );
 a33284a <=( (not A167)  and  A169 );
 a33285a <=( (not A170)  and  a33284a );
 a33289a <=( A200  and  A199 );
 a33290a <=( (not A166)  and  a33289a );
 a33291a <=( a33290a  and  a33285a );
 a33295a <=( (not A266)  and  (not A234) );
 a33296a <=( (not A233)  and  a33295a );
 a33300a <=( (not A300)  and  A298 );
 a33301a <=( (not A267)  and  a33300a );
 a33302a <=( a33301a  and  a33296a );
 a33306a <=( (not A167)  and  A169 );
 a33307a <=( (not A170)  and  a33306a );
 a33311a <=( A200  and  A199 );
 a33312a <=( (not A166)  and  a33311a );
 a33313a <=( a33312a  and  a33307a );
 a33317a <=( (not A266)  and  (not A234) );
 a33318a <=( (not A233)  and  a33317a );
 a33322a <=( A299  and  A298 );
 a33323a <=( (not A267)  and  a33322a );
 a33324a <=( a33323a  and  a33318a );
 a33328a <=( (not A167)  and  A169 );
 a33329a <=( (not A170)  and  a33328a );
 a33333a <=( A200  and  A199 );
 a33334a <=( (not A166)  and  a33333a );
 a33335a <=( a33334a  and  a33329a );
 a33339a <=( (not A266)  and  (not A234) );
 a33340a <=( (not A233)  and  a33339a );
 a33344a <=( (not A299)  and  (not A298) );
 a33345a <=( (not A267)  and  a33344a );
 a33346a <=( a33345a  and  a33340a );
 a33350a <=( (not A167)  and  A169 );
 a33351a <=( (not A170)  and  a33350a );
 a33355a <=( A200  and  A199 );
 a33356a <=( (not A166)  and  a33355a );
 a33357a <=( a33356a  and  a33351a );
 a33361a <=( (not A265)  and  (not A234) );
 a33362a <=( (not A233)  and  a33361a );
 a33366a <=( (not A300)  and  A298 );
 a33367a <=( (not A266)  and  a33366a );
 a33368a <=( a33367a  and  a33362a );
 a33372a <=( (not A167)  and  A169 );
 a33373a <=( (not A170)  and  a33372a );
 a33377a <=( A200  and  A199 );
 a33378a <=( (not A166)  and  a33377a );
 a33379a <=( a33378a  and  a33373a );
 a33383a <=( (not A265)  and  (not A234) );
 a33384a <=( (not A233)  and  a33383a );
 a33388a <=( A299  and  A298 );
 a33389a <=( (not A266)  and  a33388a );
 a33390a <=( a33389a  and  a33384a );
 a33394a <=( (not A167)  and  A169 );
 a33395a <=( (not A170)  and  a33394a );
 a33399a <=( A200  and  A199 );
 a33400a <=( (not A166)  and  a33399a );
 a33401a <=( a33400a  and  a33395a );
 a33405a <=( (not A265)  and  (not A234) );
 a33406a <=( (not A233)  and  a33405a );
 a33410a <=( (not A299)  and  (not A298) );
 a33411a <=( (not A266)  and  a33410a );
 a33412a <=( a33411a  and  a33406a );
 a33416a <=( (not A167)  and  A169 );
 a33417a <=( (not A170)  and  a33416a );
 a33421a <=( A200  and  A199 );
 a33422a <=( (not A166)  and  a33421a );
 a33423a <=( a33422a  and  a33417a );
 a33427a <=( A234  and  (not A233) );
 a33428a <=( A232  and  a33427a );
 a33432a <=( A299  and  (not A298) );
 a33433a <=( A235  and  a33432a );
 a33434a <=( a33433a  and  a33428a );
 a33438a <=( (not A167)  and  A169 );
 a33439a <=( (not A170)  and  a33438a );
 a33443a <=( A200  and  A199 );
 a33444a <=( (not A166)  and  a33443a );
 a33445a <=( a33444a  and  a33439a );
 a33449a <=( A234  and  (not A233) );
 a33450a <=( A232  and  a33449a );
 a33454a <=( A266  and  (not A265) );
 a33455a <=( A235  and  a33454a );
 a33456a <=( a33455a  and  a33450a );
 a33460a <=( (not A167)  and  A169 );
 a33461a <=( (not A170)  and  a33460a );
 a33465a <=( A200  and  A199 );
 a33466a <=( (not A166)  and  a33465a );
 a33467a <=( a33466a  and  a33461a );
 a33471a <=( A234  and  (not A233) );
 a33472a <=( A232  and  a33471a );
 a33476a <=( A299  and  (not A298) );
 a33477a <=( A236  and  a33476a );
 a33478a <=( a33477a  and  a33472a );
 a33482a <=( (not A167)  and  A169 );
 a33483a <=( (not A170)  and  a33482a );
 a33487a <=( A200  and  A199 );
 a33488a <=( (not A166)  and  a33487a );
 a33489a <=( a33488a  and  a33483a );
 a33493a <=( A234  and  (not A233) );
 a33494a <=( A232  and  a33493a );
 a33498a <=( A266  and  (not A265) );
 a33499a <=( A236  and  a33498a );
 a33500a <=( a33499a  and  a33494a );
 a33504a <=( (not A167)  and  A169 );
 a33505a <=( (not A170)  and  a33504a );
 a33509a <=( A200  and  A199 );
 a33510a <=( (not A166)  and  a33509a );
 a33511a <=( a33510a  and  a33505a );
 a33515a <=( A265  and  (not A233) );
 a33516a <=( (not A232)  and  a33515a );
 a33520a <=( (not A300)  and  A298 );
 a33521a <=( A266  and  a33520a );
 a33522a <=( a33521a  and  a33516a );
 a33526a <=( (not A167)  and  A169 );
 a33527a <=( (not A170)  and  a33526a );
 a33531a <=( A200  and  A199 );
 a33532a <=( (not A166)  and  a33531a );
 a33533a <=( a33532a  and  a33527a );
 a33537a <=( A265  and  (not A233) );
 a33538a <=( (not A232)  and  a33537a );
 a33542a <=( A299  and  A298 );
 a33543a <=( A266  and  a33542a );
 a33544a <=( a33543a  and  a33538a );
 a33548a <=( (not A167)  and  A169 );
 a33549a <=( (not A170)  and  a33548a );
 a33553a <=( A200  and  A199 );
 a33554a <=( (not A166)  and  a33553a );
 a33555a <=( a33554a  and  a33549a );
 a33559a <=( A265  and  (not A233) );
 a33560a <=( (not A232)  and  a33559a );
 a33564a <=( (not A299)  and  (not A298) );
 a33565a <=( A266  and  a33564a );
 a33566a <=( a33565a  and  a33560a );
 a33570a <=( (not A167)  and  A169 );
 a33571a <=( (not A170)  and  a33570a );
 a33575a <=( A200  and  A199 );
 a33576a <=( (not A166)  and  a33575a );
 a33577a <=( a33576a  and  a33571a );
 a33581a <=( (not A266)  and  (not A233) );
 a33582a <=( (not A232)  and  a33581a );
 a33586a <=( (not A300)  and  A298 );
 a33587a <=( (not A267)  and  a33586a );
 a33588a <=( a33587a  and  a33582a );
 a33592a <=( (not A167)  and  A169 );
 a33593a <=( (not A170)  and  a33592a );
 a33597a <=( A200  and  A199 );
 a33598a <=( (not A166)  and  a33597a );
 a33599a <=( a33598a  and  a33593a );
 a33603a <=( (not A266)  and  (not A233) );
 a33604a <=( (not A232)  and  a33603a );
 a33608a <=( A299  and  A298 );
 a33609a <=( (not A267)  and  a33608a );
 a33610a <=( a33609a  and  a33604a );
 a33614a <=( (not A167)  and  A169 );
 a33615a <=( (not A170)  and  a33614a );
 a33619a <=( A200  and  A199 );
 a33620a <=( (not A166)  and  a33619a );
 a33621a <=( a33620a  and  a33615a );
 a33625a <=( (not A266)  and  (not A233) );
 a33626a <=( (not A232)  and  a33625a );
 a33630a <=( (not A299)  and  (not A298) );
 a33631a <=( (not A267)  and  a33630a );
 a33632a <=( a33631a  and  a33626a );
 a33636a <=( (not A167)  and  A169 );
 a33637a <=( (not A170)  and  a33636a );
 a33641a <=( A200  and  A199 );
 a33642a <=( (not A166)  and  a33641a );
 a33643a <=( a33642a  and  a33637a );
 a33647a <=( (not A265)  and  (not A233) );
 a33648a <=( (not A232)  and  a33647a );
 a33652a <=( (not A300)  and  A298 );
 a33653a <=( (not A266)  and  a33652a );
 a33654a <=( a33653a  and  a33648a );
 a33658a <=( (not A167)  and  A169 );
 a33659a <=( (not A170)  and  a33658a );
 a33663a <=( A200  and  A199 );
 a33664a <=( (not A166)  and  a33663a );
 a33665a <=( a33664a  and  a33659a );
 a33669a <=( (not A265)  and  (not A233) );
 a33670a <=( (not A232)  and  a33669a );
 a33674a <=( A299  and  A298 );
 a33675a <=( (not A266)  and  a33674a );
 a33676a <=( a33675a  and  a33670a );
 a33680a <=( (not A167)  and  A169 );
 a33681a <=( (not A170)  and  a33680a );
 a33685a <=( A200  and  A199 );
 a33686a <=( (not A166)  and  a33685a );
 a33687a <=( a33686a  and  a33681a );
 a33691a <=( (not A265)  and  (not A233) );
 a33692a <=( (not A232)  and  a33691a );
 a33696a <=( (not A299)  and  (not A298) );
 a33697a <=( (not A266)  and  a33696a );
 a33698a <=( a33697a  and  a33692a );
 a33702a <=( (not A167)  and  A169 );
 a33703a <=( (not A170)  and  a33702a );
 a33707a <=( (not A201)  and  (not A200) );
 a33708a <=( (not A166)  and  a33707a );
 a33709a <=( a33708a  and  a33703a );
 a33713a <=( A265  and  A233 );
 a33714a <=( A232  and  a33713a );
 a33718a <=( (not A300)  and  (not A299) );
 a33719a <=( (not A267)  and  a33718a );
 a33720a <=( a33719a  and  a33714a );
 a33724a <=( (not A167)  and  A169 );
 a33725a <=( (not A170)  and  a33724a );
 a33729a <=( (not A201)  and  (not A200) );
 a33730a <=( (not A166)  and  a33729a );
 a33731a <=( a33730a  and  a33725a );
 a33735a <=( A265  and  A233 );
 a33736a <=( A232  and  a33735a );
 a33740a <=( A299  and  A298 );
 a33741a <=( (not A267)  and  a33740a );
 a33742a <=( a33741a  and  a33736a );
 a33746a <=( (not A167)  and  A169 );
 a33747a <=( (not A170)  and  a33746a );
 a33751a <=( (not A201)  and  (not A200) );
 a33752a <=( (not A166)  and  a33751a );
 a33753a <=( a33752a  and  a33747a );
 a33757a <=( A265  and  A233 );
 a33758a <=( A232  and  a33757a );
 a33762a <=( (not A299)  and  (not A298) );
 a33763a <=( (not A267)  and  a33762a );
 a33764a <=( a33763a  and  a33758a );
 a33768a <=( (not A167)  and  A169 );
 a33769a <=( (not A170)  and  a33768a );
 a33773a <=( (not A201)  and  (not A200) );
 a33774a <=( (not A166)  and  a33773a );
 a33775a <=( a33774a  and  a33769a );
 a33779a <=( A265  and  A233 );
 a33780a <=( A232  and  a33779a );
 a33784a <=( (not A300)  and  (not A299) );
 a33785a <=( A266  and  a33784a );
 a33786a <=( a33785a  and  a33780a );
 a33790a <=( (not A167)  and  A169 );
 a33791a <=( (not A170)  and  a33790a );
 a33795a <=( (not A201)  and  (not A200) );
 a33796a <=( (not A166)  and  a33795a );
 a33797a <=( a33796a  and  a33791a );
 a33801a <=( A265  and  A233 );
 a33802a <=( A232  and  a33801a );
 a33806a <=( A299  and  A298 );
 a33807a <=( A266  and  a33806a );
 a33808a <=( a33807a  and  a33802a );
 a33812a <=( (not A167)  and  A169 );
 a33813a <=( (not A170)  and  a33812a );
 a33817a <=( (not A201)  and  (not A200) );
 a33818a <=( (not A166)  and  a33817a );
 a33819a <=( a33818a  and  a33813a );
 a33823a <=( A265  and  A233 );
 a33824a <=( A232  and  a33823a );
 a33828a <=( (not A299)  and  (not A298) );
 a33829a <=( A266  and  a33828a );
 a33830a <=( a33829a  and  a33824a );
 a33834a <=( (not A167)  and  A169 );
 a33835a <=( (not A170)  and  a33834a );
 a33839a <=( (not A201)  and  (not A200) );
 a33840a <=( (not A166)  and  a33839a );
 a33841a <=( a33840a  and  a33835a );
 a33845a <=( (not A265)  and  A233 );
 a33846a <=( A232  and  a33845a );
 a33850a <=( (not A300)  and  (not A299) );
 a33851a <=( (not A266)  and  a33850a );
 a33852a <=( a33851a  and  a33846a );
 a33856a <=( (not A167)  and  A169 );
 a33857a <=( (not A170)  and  a33856a );
 a33861a <=( (not A201)  and  (not A200) );
 a33862a <=( (not A166)  and  a33861a );
 a33863a <=( a33862a  and  a33857a );
 a33867a <=( (not A265)  and  A233 );
 a33868a <=( A232  and  a33867a );
 a33872a <=( A299  and  A298 );
 a33873a <=( (not A266)  and  a33872a );
 a33874a <=( a33873a  and  a33868a );
 a33878a <=( (not A167)  and  A169 );
 a33879a <=( (not A170)  and  a33878a );
 a33883a <=( (not A201)  and  (not A200) );
 a33884a <=( (not A166)  and  a33883a );
 a33885a <=( a33884a  and  a33879a );
 a33889a <=( (not A265)  and  A233 );
 a33890a <=( A232  and  a33889a );
 a33894a <=( (not A299)  and  (not A298) );
 a33895a <=( (not A266)  and  a33894a );
 a33896a <=( a33895a  and  a33890a );
 a33900a <=( (not A167)  and  A169 );
 a33901a <=( (not A170)  and  a33900a );
 a33905a <=( (not A201)  and  (not A200) );
 a33906a <=( (not A166)  and  a33905a );
 a33907a <=( a33906a  and  a33901a );
 a33911a <=( A298  and  A233 );
 a33912a <=( (not A232)  and  a33911a );
 a33916a <=( A301  and  A300 );
 a33917a <=( (not A299)  and  a33916a );
 a33918a <=( a33917a  and  a33912a );
 a33922a <=( (not A167)  and  A169 );
 a33923a <=( (not A170)  and  a33922a );
 a33927a <=( (not A201)  and  (not A200) );
 a33928a <=( (not A166)  and  a33927a );
 a33929a <=( a33928a  and  a33923a );
 a33933a <=( A298  and  A233 );
 a33934a <=( (not A232)  and  a33933a );
 a33938a <=( A302  and  A300 );
 a33939a <=( (not A299)  and  a33938a );
 a33940a <=( a33939a  and  a33934a );
 a33944a <=( (not A167)  and  A169 );
 a33945a <=( (not A170)  and  a33944a );
 a33949a <=( (not A201)  and  (not A200) );
 a33950a <=( (not A166)  and  a33949a );
 a33951a <=( a33950a  and  a33945a );
 a33955a <=( A265  and  A233 );
 a33956a <=( (not A232)  and  a33955a );
 a33960a <=( A268  and  A267 );
 a33961a <=( (not A266)  and  a33960a );
 a33962a <=( a33961a  and  a33956a );
 a33966a <=( (not A167)  and  A169 );
 a33967a <=( (not A170)  and  a33966a );
 a33971a <=( (not A201)  and  (not A200) );
 a33972a <=( (not A166)  and  a33971a );
 a33973a <=( a33972a  and  a33967a );
 a33977a <=( A265  and  A233 );
 a33978a <=( (not A232)  and  a33977a );
 a33982a <=( A269  and  A267 );
 a33983a <=( (not A266)  and  a33982a );
 a33984a <=( a33983a  and  a33978a );
 a33988a <=( (not A167)  and  A169 );
 a33989a <=( (not A170)  and  a33988a );
 a33993a <=( (not A201)  and  (not A200) );
 a33994a <=( (not A166)  and  a33993a );
 a33995a <=( a33994a  and  a33989a );
 a33999a <=( A265  and  (not A234) );
 a34000a <=( (not A233)  and  a33999a );
 a34004a <=( (not A300)  and  A298 );
 a34005a <=( A266  and  a34004a );
 a34006a <=( a34005a  and  a34000a );
 a34010a <=( (not A167)  and  A169 );
 a34011a <=( (not A170)  and  a34010a );
 a34015a <=( (not A201)  and  (not A200) );
 a34016a <=( (not A166)  and  a34015a );
 a34017a <=( a34016a  and  a34011a );
 a34021a <=( A265  and  (not A234) );
 a34022a <=( (not A233)  and  a34021a );
 a34026a <=( A299  and  A298 );
 a34027a <=( A266  and  a34026a );
 a34028a <=( a34027a  and  a34022a );
 a34032a <=( (not A167)  and  A169 );
 a34033a <=( (not A170)  and  a34032a );
 a34037a <=( (not A201)  and  (not A200) );
 a34038a <=( (not A166)  and  a34037a );
 a34039a <=( a34038a  and  a34033a );
 a34043a <=( A265  and  (not A234) );
 a34044a <=( (not A233)  and  a34043a );
 a34048a <=( (not A299)  and  (not A298) );
 a34049a <=( A266  and  a34048a );
 a34050a <=( a34049a  and  a34044a );
 a34054a <=( (not A167)  and  A169 );
 a34055a <=( (not A170)  and  a34054a );
 a34059a <=( (not A201)  and  (not A200) );
 a34060a <=( (not A166)  and  a34059a );
 a34061a <=( a34060a  and  a34055a );
 a34065a <=( (not A266)  and  (not A234) );
 a34066a <=( (not A233)  and  a34065a );
 a34070a <=( (not A300)  and  A298 );
 a34071a <=( (not A267)  and  a34070a );
 a34072a <=( a34071a  and  a34066a );
 a34076a <=( (not A167)  and  A169 );
 a34077a <=( (not A170)  and  a34076a );
 a34081a <=( (not A201)  and  (not A200) );
 a34082a <=( (not A166)  and  a34081a );
 a34083a <=( a34082a  and  a34077a );
 a34087a <=( (not A266)  and  (not A234) );
 a34088a <=( (not A233)  and  a34087a );
 a34092a <=( A299  and  A298 );
 a34093a <=( (not A267)  and  a34092a );
 a34094a <=( a34093a  and  a34088a );
 a34098a <=( (not A167)  and  A169 );
 a34099a <=( (not A170)  and  a34098a );
 a34103a <=( (not A201)  and  (not A200) );
 a34104a <=( (not A166)  and  a34103a );
 a34105a <=( a34104a  and  a34099a );
 a34109a <=( (not A266)  and  (not A234) );
 a34110a <=( (not A233)  and  a34109a );
 a34114a <=( (not A299)  and  (not A298) );
 a34115a <=( (not A267)  and  a34114a );
 a34116a <=( a34115a  and  a34110a );
 a34120a <=( (not A167)  and  A169 );
 a34121a <=( (not A170)  and  a34120a );
 a34125a <=( (not A201)  and  (not A200) );
 a34126a <=( (not A166)  and  a34125a );
 a34127a <=( a34126a  and  a34121a );
 a34131a <=( (not A265)  and  (not A234) );
 a34132a <=( (not A233)  and  a34131a );
 a34136a <=( (not A300)  and  A298 );
 a34137a <=( (not A266)  and  a34136a );
 a34138a <=( a34137a  and  a34132a );
 a34142a <=( (not A167)  and  A169 );
 a34143a <=( (not A170)  and  a34142a );
 a34147a <=( (not A201)  and  (not A200) );
 a34148a <=( (not A166)  and  a34147a );
 a34149a <=( a34148a  and  a34143a );
 a34153a <=( (not A265)  and  (not A234) );
 a34154a <=( (not A233)  and  a34153a );
 a34158a <=( A299  and  A298 );
 a34159a <=( (not A266)  and  a34158a );
 a34160a <=( a34159a  and  a34154a );
 a34164a <=( (not A167)  and  A169 );
 a34165a <=( (not A170)  and  a34164a );
 a34169a <=( (not A201)  and  (not A200) );
 a34170a <=( (not A166)  and  a34169a );
 a34171a <=( a34170a  and  a34165a );
 a34175a <=( (not A265)  and  (not A234) );
 a34176a <=( (not A233)  and  a34175a );
 a34180a <=( (not A299)  and  (not A298) );
 a34181a <=( (not A266)  and  a34180a );
 a34182a <=( a34181a  and  a34176a );
 a34186a <=( (not A167)  and  A169 );
 a34187a <=( (not A170)  and  a34186a );
 a34191a <=( (not A201)  and  (not A200) );
 a34192a <=( (not A166)  and  a34191a );
 a34193a <=( a34192a  and  a34187a );
 a34197a <=( A234  and  (not A233) );
 a34198a <=( A232  and  a34197a );
 a34202a <=( A299  and  (not A298) );
 a34203a <=( A235  and  a34202a );
 a34204a <=( a34203a  and  a34198a );
 a34208a <=( (not A167)  and  A169 );
 a34209a <=( (not A170)  and  a34208a );
 a34213a <=( (not A201)  and  (not A200) );
 a34214a <=( (not A166)  and  a34213a );
 a34215a <=( a34214a  and  a34209a );
 a34219a <=( A234  and  (not A233) );
 a34220a <=( A232  and  a34219a );
 a34224a <=( A266  and  (not A265) );
 a34225a <=( A235  and  a34224a );
 a34226a <=( a34225a  and  a34220a );
 a34230a <=( (not A167)  and  A169 );
 a34231a <=( (not A170)  and  a34230a );
 a34235a <=( (not A201)  and  (not A200) );
 a34236a <=( (not A166)  and  a34235a );
 a34237a <=( a34236a  and  a34231a );
 a34241a <=( A234  and  (not A233) );
 a34242a <=( A232  and  a34241a );
 a34246a <=( A299  and  (not A298) );
 a34247a <=( A236  and  a34246a );
 a34248a <=( a34247a  and  a34242a );
 a34252a <=( (not A167)  and  A169 );
 a34253a <=( (not A170)  and  a34252a );
 a34257a <=( (not A201)  and  (not A200) );
 a34258a <=( (not A166)  and  a34257a );
 a34259a <=( a34258a  and  a34253a );
 a34263a <=( A234  and  (not A233) );
 a34264a <=( A232  and  a34263a );
 a34268a <=( A266  and  (not A265) );
 a34269a <=( A236  and  a34268a );
 a34270a <=( a34269a  and  a34264a );
 a34274a <=( (not A167)  and  A169 );
 a34275a <=( (not A170)  and  a34274a );
 a34279a <=( (not A201)  and  (not A200) );
 a34280a <=( (not A166)  and  a34279a );
 a34281a <=( a34280a  and  a34275a );
 a34285a <=( A265  and  (not A233) );
 a34286a <=( (not A232)  and  a34285a );
 a34290a <=( (not A300)  and  A298 );
 a34291a <=( A266  and  a34290a );
 a34292a <=( a34291a  and  a34286a );
 a34296a <=( (not A167)  and  A169 );
 a34297a <=( (not A170)  and  a34296a );
 a34301a <=( (not A201)  and  (not A200) );
 a34302a <=( (not A166)  and  a34301a );
 a34303a <=( a34302a  and  a34297a );
 a34307a <=( A265  and  (not A233) );
 a34308a <=( (not A232)  and  a34307a );
 a34312a <=( A299  and  A298 );
 a34313a <=( A266  and  a34312a );
 a34314a <=( a34313a  and  a34308a );
 a34318a <=( (not A167)  and  A169 );
 a34319a <=( (not A170)  and  a34318a );
 a34323a <=( (not A201)  and  (not A200) );
 a34324a <=( (not A166)  and  a34323a );
 a34325a <=( a34324a  and  a34319a );
 a34329a <=( A265  and  (not A233) );
 a34330a <=( (not A232)  and  a34329a );
 a34334a <=( (not A299)  and  (not A298) );
 a34335a <=( A266  and  a34334a );
 a34336a <=( a34335a  and  a34330a );
 a34340a <=( (not A167)  and  A169 );
 a34341a <=( (not A170)  and  a34340a );
 a34345a <=( (not A201)  and  (not A200) );
 a34346a <=( (not A166)  and  a34345a );
 a34347a <=( a34346a  and  a34341a );
 a34351a <=( (not A266)  and  (not A233) );
 a34352a <=( (not A232)  and  a34351a );
 a34356a <=( (not A300)  and  A298 );
 a34357a <=( (not A267)  and  a34356a );
 a34358a <=( a34357a  and  a34352a );
 a34362a <=( (not A167)  and  A169 );
 a34363a <=( (not A170)  and  a34362a );
 a34367a <=( (not A201)  and  (not A200) );
 a34368a <=( (not A166)  and  a34367a );
 a34369a <=( a34368a  and  a34363a );
 a34373a <=( (not A266)  and  (not A233) );
 a34374a <=( (not A232)  and  a34373a );
 a34378a <=( A299  and  A298 );
 a34379a <=( (not A267)  and  a34378a );
 a34380a <=( a34379a  and  a34374a );
 a34384a <=( (not A167)  and  A169 );
 a34385a <=( (not A170)  and  a34384a );
 a34389a <=( (not A201)  and  (not A200) );
 a34390a <=( (not A166)  and  a34389a );
 a34391a <=( a34390a  and  a34385a );
 a34395a <=( (not A266)  and  (not A233) );
 a34396a <=( (not A232)  and  a34395a );
 a34400a <=( (not A299)  and  (not A298) );
 a34401a <=( (not A267)  and  a34400a );
 a34402a <=( a34401a  and  a34396a );
 a34406a <=( (not A167)  and  A169 );
 a34407a <=( (not A170)  and  a34406a );
 a34411a <=( (not A201)  and  (not A200) );
 a34412a <=( (not A166)  and  a34411a );
 a34413a <=( a34412a  and  a34407a );
 a34417a <=( (not A265)  and  (not A233) );
 a34418a <=( (not A232)  and  a34417a );
 a34422a <=( (not A300)  and  A298 );
 a34423a <=( (not A266)  and  a34422a );
 a34424a <=( a34423a  and  a34418a );
 a34428a <=( (not A167)  and  A169 );
 a34429a <=( (not A170)  and  a34428a );
 a34433a <=( (not A201)  and  (not A200) );
 a34434a <=( (not A166)  and  a34433a );
 a34435a <=( a34434a  and  a34429a );
 a34439a <=( (not A265)  and  (not A233) );
 a34440a <=( (not A232)  and  a34439a );
 a34444a <=( A299  and  A298 );
 a34445a <=( (not A266)  and  a34444a );
 a34446a <=( a34445a  and  a34440a );
 a34450a <=( (not A167)  and  A169 );
 a34451a <=( (not A170)  and  a34450a );
 a34455a <=( (not A201)  and  (not A200) );
 a34456a <=( (not A166)  and  a34455a );
 a34457a <=( a34456a  and  a34451a );
 a34461a <=( (not A265)  and  (not A233) );
 a34462a <=( (not A232)  and  a34461a );
 a34466a <=( (not A299)  and  (not A298) );
 a34467a <=( (not A266)  and  a34466a );
 a34468a <=( a34467a  and  a34462a );
 a34472a <=( (not A167)  and  A169 );
 a34473a <=( (not A170)  and  a34472a );
 a34477a <=( (not A200)  and  (not A199) );
 a34478a <=( (not A166)  and  a34477a );
 a34479a <=( a34478a  and  a34473a );
 a34483a <=( A265  and  A233 );
 a34484a <=( A232  and  a34483a );
 a34488a <=( (not A300)  and  (not A299) );
 a34489a <=( (not A267)  and  a34488a );
 a34490a <=( a34489a  and  a34484a );
 a34494a <=( (not A167)  and  A169 );
 a34495a <=( (not A170)  and  a34494a );
 a34499a <=( (not A200)  and  (not A199) );
 a34500a <=( (not A166)  and  a34499a );
 a34501a <=( a34500a  and  a34495a );
 a34505a <=( A265  and  A233 );
 a34506a <=( A232  and  a34505a );
 a34510a <=( A299  and  A298 );
 a34511a <=( (not A267)  and  a34510a );
 a34512a <=( a34511a  and  a34506a );
 a34516a <=( (not A167)  and  A169 );
 a34517a <=( (not A170)  and  a34516a );
 a34521a <=( (not A200)  and  (not A199) );
 a34522a <=( (not A166)  and  a34521a );
 a34523a <=( a34522a  and  a34517a );
 a34527a <=( A265  and  A233 );
 a34528a <=( A232  and  a34527a );
 a34532a <=( (not A299)  and  (not A298) );
 a34533a <=( (not A267)  and  a34532a );
 a34534a <=( a34533a  and  a34528a );
 a34538a <=( (not A167)  and  A169 );
 a34539a <=( (not A170)  and  a34538a );
 a34543a <=( (not A200)  and  (not A199) );
 a34544a <=( (not A166)  and  a34543a );
 a34545a <=( a34544a  and  a34539a );
 a34549a <=( A265  and  A233 );
 a34550a <=( A232  and  a34549a );
 a34554a <=( (not A300)  and  (not A299) );
 a34555a <=( A266  and  a34554a );
 a34556a <=( a34555a  and  a34550a );
 a34560a <=( (not A167)  and  A169 );
 a34561a <=( (not A170)  and  a34560a );
 a34565a <=( (not A200)  and  (not A199) );
 a34566a <=( (not A166)  and  a34565a );
 a34567a <=( a34566a  and  a34561a );
 a34571a <=( A265  and  A233 );
 a34572a <=( A232  and  a34571a );
 a34576a <=( A299  and  A298 );
 a34577a <=( A266  and  a34576a );
 a34578a <=( a34577a  and  a34572a );
 a34582a <=( (not A167)  and  A169 );
 a34583a <=( (not A170)  and  a34582a );
 a34587a <=( (not A200)  and  (not A199) );
 a34588a <=( (not A166)  and  a34587a );
 a34589a <=( a34588a  and  a34583a );
 a34593a <=( A265  and  A233 );
 a34594a <=( A232  and  a34593a );
 a34598a <=( (not A299)  and  (not A298) );
 a34599a <=( A266  and  a34598a );
 a34600a <=( a34599a  and  a34594a );
 a34604a <=( (not A167)  and  A169 );
 a34605a <=( (not A170)  and  a34604a );
 a34609a <=( (not A200)  and  (not A199) );
 a34610a <=( (not A166)  and  a34609a );
 a34611a <=( a34610a  and  a34605a );
 a34615a <=( (not A265)  and  A233 );
 a34616a <=( A232  and  a34615a );
 a34620a <=( (not A300)  and  (not A299) );
 a34621a <=( (not A266)  and  a34620a );
 a34622a <=( a34621a  and  a34616a );
 a34626a <=( (not A167)  and  A169 );
 a34627a <=( (not A170)  and  a34626a );
 a34631a <=( (not A200)  and  (not A199) );
 a34632a <=( (not A166)  and  a34631a );
 a34633a <=( a34632a  and  a34627a );
 a34637a <=( (not A265)  and  A233 );
 a34638a <=( A232  and  a34637a );
 a34642a <=( A299  and  A298 );
 a34643a <=( (not A266)  and  a34642a );
 a34644a <=( a34643a  and  a34638a );
 a34648a <=( (not A167)  and  A169 );
 a34649a <=( (not A170)  and  a34648a );
 a34653a <=( (not A200)  and  (not A199) );
 a34654a <=( (not A166)  and  a34653a );
 a34655a <=( a34654a  and  a34649a );
 a34659a <=( (not A265)  and  A233 );
 a34660a <=( A232  and  a34659a );
 a34664a <=( (not A299)  and  (not A298) );
 a34665a <=( (not A266)  and  a34664a );
 a34666a <=( a34665a  and  a34660a );
 a34670a <=( (not A167)  and  A169 );
 a34671a <=( (not A170)  and  a34670a );
 a34675a <=( (not A200)  and  (not A199) );
 a34676a <=( (not A166)  and  a34675a );
 a34677a <=( a34676a  and  a34671a );
 a34681a <=( A298  and  A233 );
 a34682a <=( (not A232)  and  a34681a );
 a34686a <=( A301  and  A300 );
 a34687a <=( (not A299)  and  a34686a );
 a34688a <=( a34687a  and  a34682a );
 a34692a <=( (not A167)  and  A169 );
 a34693a <=( (not A170)  and  a34692a );
 a34697a <=( (not A200)  and  (not A199) );
 a34698a <=( (not A166)  and  a34697a );
 a34699a <=( a34698a  and  a34693a );
 a34703a <=( A298  and  A233 );
 a34704a <=( (not A232)  and  a34703a );
 a34708a <=( A302  and  A300 );
 a34709a <=( (not A299)  and  a34708a );
 a34710a <=( a34709a  and  a34704a );
 a34714a <=( (not A167)  and  A169 );
 a34715a <=( (not A170)  and  a34714a );
 a34719a <=( (not A200)  and  (not A199) );
 a34720a <=( (not A166)  and  a34719a );
 a34721a <=( a34720a  and  a34715a );
 a34725a <=( A265  and  A233 );
 a34726a <=( (not A232)  and  a34725a );
 a34730a <=( A268  and  A267 );
 a34731a <=( (not A266)  and  a34730a );
 a34732a <=( a34731a  and  a34726a );
 a34736a <=( (not A167)  and  A169 );
 a34737a <=( (not A170)  and  a34736a );
 a34741a <=( (not A200)  and  (not A199) );
 a34742a <=( (not A166)  and  a34741a );
 a34743a <=( a34742a  and  a34737a );
 a34747a <=( A265  and  A233 );
 a34748a <=( (not A232)  and  a34747a );
 a34752a <=( A269  and  A267 );
 a34753a <=( (not A266)  and  a34752a );
 a34754a <=( a34753a  and  a34748a );
 a34758a <=( (not A167)  and  A169 );
 a34759a <=( (not A170)  and  a34758a );
 a34763a <=( (not A200)  and  (not A199) );
 a34764a <=( (not A166)  and  a34763a );
 a34765a <=( a34764a  and  a34759a );
 a34769a <=( A265  and  (not A234) );
 a34770a <=( (not A233)  and  a34769a );
 a34774a <=( (not A300)  and  A298 );
 a34775a <=( A266  and  a34774a );
 a34776a <=( a34775a  and  a34770a );
 a34780a <=( (not A167)  and  A169 );
 a34781a <=( (not A170)  and  a34780a );
 a34785a <=( (not A200)  and  (not A199) );
 a34786a <=( (not A166)  and  a34785a );
 a34787a <=( a34786a  and  a34781a );
 a34791a <=( A265  and  (not A234) );
 a34792a <=( (not A233)  and  a34791a );
 a34796a <=( A299  and  A298 );
 a34797a <=( A266  and  a34796a );
 a34798a <=( a34797a  and  a34792a );
 a34802a <=( (not A167)  and  A169 );
 a34803a <=( (not A170)  and  a34802a );
 a34807a <=( (not A200)  and  (not A199) );
 a34808a <=( (not A166)  and  a34807a );
 a34809a <=( a34808a  and  a34803a );
 a34813a <=( A265  and  (not A234) );
 a34814a <=( (not A233)  and  a34813a );
 a34818a <=( (not A299)  and  (not A298) );
 a34819a <=( A266  and  a34818a );
 a34820a <=( a34819a  and  a34814a );
 a34824a <=( (not A167)  and  A169 );
 a34825a <=( (not A170)  and  a34824a );
 a34829a <=( (not A200)  and  (not A199) );
 a34830a <=( (not A166)  and  a34829a );
 a34831a <=( a34830a  and  a34825a );
 a34835a <=( (not A266)  and  (not A234) );
 a34836a <=( (not A233)  and  a34835a );
 a34840a <=( (not A300)  and  A298 );
 a34841a <=( (not A267)  and  a34840a );
 a34842a <=( a34841a  and  a34836a );
 a34846a <=( (not A167)  and  A169 );
 a34847a <=( (not A170)  and  a34846a );
 a34851a <=( (not A200)  and  (not A199) );
 a34852a <=( (not A166)  and  a34851a );
 a34853a <=( a34852a  and  a34847a );
 a34857a <=( (not A266)  and  (not A234) );
 a34858a <=( (not A233)  and  a34857a );
 a34862a <=( A299  and  A298 );
 a34863a <=( (not A267)  and  a34862a );
 a34864a <=( a34863a  and  a34858a );
 a34868a <=( (not A167)  and  A169 );
 a34869a <=( (not A170)  and  a34868a );
 a34873a <=( (not A200)  and  (not A199) );
 a34874a <=( (not A166)  and  a34873a );
 a34875a <=( a34874a  and  a34869a );
 a34879a <=( (not A266)  and  (not A234) );
 a34880a <=( (not A233)  and  a34879a );
 a34884a <=( (not A299)  and  (not A298) );
 a34885a <=( (not A267)  and  a34884a );
 a34886a <=( a34885a  and  a34880a );
 a34890a <=( (not A167)  and  A169 );
 a34891a <=( (not A170)  and  a34890a );
 a34895a <=( (not A200)  and  (not A199) );
 a34896a <=( (not A166)  and  a34895a );
 a34897a <=( a34896a  and  a34891a );
 a34901a <=( (not A265)  and  (not A234) );
 a34902a <=( (not A233)  and  a34901a );
 a34906a <=( (not A300)  and  A298 );
 a34907a <=( (not A266)  and  a34906a );
 a34908a <=( a34907a  and  a34902a );
 a34912a <=( (not A167)  and  A169 );
 a34913a <=( (not A170)  and  a34912a );
 a34917a <=( (not A200)  and  (not A199) );
 a34918a <=( (not A166)  and  a34917a );
 a34919a <=( a34918a  and  a34913a );
 a34923a <=( (not A265)  and  (not A234) );
 a34924a <=( (not A233)  and  a34923a );
 a34928a <=( A299  and  A298 );
 a34929a <=( (not A266)  and  a34928a );
 a34930a <=( a34929a  and  a34924a );
 a34934a <=( (not A167)  and  A169 );
 a34935a <=( (not A170)  and  a34934a );
 a34939a <=( (not A200)  and  (not A199) );
 a34940a <=( (not A166)  and  a34939a );
 a34941a <=( a34940a  and  a34935a );
 a34945a <=( (not A265)  and  (not A234) );
 a34946a <=( (not A233)  and  a34945a );
 a34950a <=( (not A299)  and  (not A298) );
 a34951a <=( (not A266)  and  a34950a );
 a34952a <=( a34951a  and  a34946a );
 a34956a <=( (not A167)  and  A169 );
 a34957a <=( (not A170)  and  a34956a );
 a34961a <=( (not A200)  and  (not A199) );
 a34962a <=( (not A166)  and  a34961a );
 a34963a <=( a34962a  and  a34957a );
 a34967a <=( A234  and  (not A233) );
 a34968a <=( A232  and  a34967a );
 a34972a <=( A299  and  (not A298) );
 a34973a <=( A235  and  a34972a );
 a34974a <=( a34973a  and  a34968a );
 a34978a <=( (not A167)  and  A169 );
 a34979a <=( (not A170)  and  a34978a );
 a34983a <=( (not A200)  and  (not A199) );
 a34984a <=( (not A166)  and  a34983a );
 a34985a <=( a34984a  and  a34979a );
 a34989a <=( A234  and  (not A233) );
 a34990a <=( A232  and  a34989a );
 a34994a <=( A266  and  (not A265) );
 a34995a <=( A235  and  a34994a );
 a34996a <=( a34995a  and  a34990a );
 a35000a <=( (not A167)  and  A169 );
 a35001a <=( (not A170)  and  a35000a );
 a35005a <=( (not A200)  and  (not A199) );
 a35006a <=( (not A166)  and  a35005a );
 a35007a <=( a35006a  and  a35001a );
 a35011a <=( A234  and  (not A233) );
 a35012a <=( A232  and  a35011a );
 a35016a <=( A299  and  (not A298) );
 a35017a <=( A236  and  a35016a );
 a35018a <=( a35017a  and  a35012a );
 a35022a <=( (not A167)  and  A169 );
 a35023a <=( (not A170)  and  a35022a );
 a35027a <=( (not A200)  and  (not A199) );
 a35028a <=( (not A166)  and  a35027a );
 a35029a <=( a35028a  and  a35023a );
 a35033a <=( A234  and  (not A233) );
 a35034a <=( A232  and  a35033a );
 a35038a <=( A266  and  (not A265) );
 a35039a <=( A236  and  a35038a );
 a35040a <=( a35039a  and  a35034a );
 a35044a <=( (not A167)  and  A169 );
 a35045a <=( (not A170)  and  a35044a );
 a35049a <=( (not A200)  and  (not A199) );
 a35050a <=( (not A166)  and  a35049a );
 a35051a <=( a35050a  and  a35045a );
 a35055a <=( A265  and  (not A233) );
 a35056a <=( (not A232)  and  a35055a );
 a35060a <=( (not A300)  and  A298 );
 a35061a <=( A266  and  a35060a );
 a35062a <=( a35061a  and  a35056a );
 a35066a <=( (not A167)  and  A169 );
 a35067a <=( (not A170)  and  a35066a );
 a35071a <=( (not A200)  and  (not A199) );
 a35072a <=( (not A166)  and  a35071a );
 a35073a <=( a35072a  and  a35067a );
 a35077a <=( A265  and  (not A233) );
 a35078a <=( (not A232)  and  a35077a );
 a35082a <=( A299  and  A298 );
 a35083a <=( A266  and  a35082a );
 a35084a <=( a35083a  and  a35078a );
 a35088a <=( (not A167)  and  A169 );
 a35089a <=( (not A170)  and  a35088a );
 a35093a <=( (not A200)  and  (not A199) );
 a35094a <=( (not A166)  and  a35093a );
 a35095a <=( a35094a  and  a35089a );
 a35099a <=( A265  and  (not A233) );
 a35100a <=( (not A232)  and  a35099a );
 a35104a <=( (not A299)  and  (not A298) );
 a35105a <=( A266  and  a35104a );
 a35106a <=( a35105a  and  a35100a );
 a35110a <=( (not A167)  and  A169 );
 a35111a <=( (not A170)  and  a35110a );
 a35115a <=( (not A200)  and  (not A199) );
 a35116a <=( (not A166)  and  a35115a );
 a35117a <=( a35116a  and  a35111a );
 a35121a <=( (not A266)  and  (not A233) );
 a35122a <=( (not A232)  and  a35121a );
 a35126a <=( (not A300)  and  A298 );
 a35127a <=( (not A267)  and  a35126a );
 a35128a <=( a35127a  and  a35122a );
 a35132a <=( (not A167)  and  A169 );
 a35133a <=( (not A170)  and  a35132a );
 a35137a <=( (not A200)  and  (not A199) );
 a35138a <=( (not A166)  and  a35137a );
 a35139a <=( a35138a  and  a35133a );
 a35143a <=( (not A266)  and  (not A233) );
 a35144a <=( (not A232)  and  a35143a );
 a35148a <=( A299  and  A298 );
 a35149a <=( (not A267)  and  a35148a );
 a35150a <=( a35149a  and  a35144a );
 a35154a <=( (not A167)  and  A169 );
 a35155a <=( (not A170)  and  a35154a );
 a35159a <=( (not A200)  and  (not A199) );
 a35160a <=( (not A166)  and  a35159a );
 a35161a <=( a35160a  and  a35155a );
 a35165a <=( (not A266)  and  (not A233) );
 a35166a <=( (not A232)  and  a35165a );
 a35170a <=( (not A299)  and  (not A298) );
 a35171a <=( (not A267)  and  a35170a );
 a35172a <=( a35171a  and  a35166a );
 a35176a <=( (not A167)  and  A169 );
 a35177a <=( (not A170)  and  a35176a );
 a35181a <=( (not A200)  and  (not A199) );
 a35182a <=( (not A166)  and  a35181a );
 a35183a <=( a35182a  and  a35177a );
 a35187a <=( (not A265)  and  (not A233) );
 a35188a <=( (not A232)  and  a35187a );
 a35192a <=( (not A300)  and  A298 );
 a35193a <=( (not A266)  and  a35192a );
 a35194a <=( a35193a  and  a35188a );
 a35198a <=( (not A167)  and  A169 );
 a35199a <=( (not A170)  and  a35198a );
 a35203a <=( (not A200)  and  (not A199) );
 a35204a <=( (not A166)  and  a35203a );
 a35205a <=( a35204a  and  a35199a );
 a35209a <=( (not A265)  and  (not A233) );
 a35210a <=( (not A232)  and  a35209a );
 a35214a <=( A299  and  A298 );
 a35215a <=( (not A266)  and  a35214a );
 a35216a <=( a35215a  and  a35210a );
 a35220a <=( (not A167)  and  A169 );
 a35221a <=( (not A170)  and  a35220a );
 a35225a <=( (not A200)  and  (not A199) );
 a35226a <=( (not A166)  and  a35225a );
 a35227a <=( a35226a  and  a35221a );
 a35231a <=( (not A265)  and  (not A233) );
 a35232a <=( (not A232)  and  a35231a );
 a35236a <=( (not A299)  and  (not A298) );
 a35237a <=( (not A266)  and  a35236a );
 a35238a <=( a35237a  and  a35232a );
 a35242a <=( (not A166)  and  (not A167) );
 a35243a <=( (not A169)  and  a35242a );
 a35247a <=( A232  and  A200 );
 a35248a <=( (not A199)  and  a35247a );
 a35249a <=( a35248a  and  a35243a );
 a35253a <=( (not A268)  and  A265 );
 a35254a <=( A233  and  a35253a );
 a35258a <=( (not A300)  and  (not A299) );
 a35259a <=( (not A269)  and  a35258a );
 a35260a <=( a35259a  and  a35254a );
 a35264a <=( (not A166)  and  (not A167) );
 a35265a <=( (not A169)  and  a35264a );
 a35269a <=( A232  and  A200 );
 a35270a <=( (not A199)  and  a35269a );
 a35271a <=( a35270a  and  a35265a );
 a35275a <=( (not A268)  and  A265 );
 a35276a <=( A233  and  a35275a );
 a35280a <=( A299  and  A298 );
 a35281a <=( (not A269)  and  a35280a );
 a35282a <=( a35281a  and  a35276a );
 a35286a <=( (not A166)  and  (not A167) );
 a35287a <=( (not A169)  and  a35286a );
 a35291a <=( A232  and  A200 );
 a35292a <=( (not A199)  and  a35291a );
 a35293a <=( a35292a  and  a35287a );
 a35297a <=( (not A268)  and  A265 );
 a35298a <=( A233  and  a35297a );
 a35302a <=( (not A299)  and  (not A298) );
 a35303a <=( (not A269)  and  a35302a );
 a35304a <=( a35303a  and  a35298a );
 a35308a <=( (not A166)  and  (not A167) );
 a35309a <=( (not A169)  and  a35308a );
 a35313a <=( A232  and  A200 );
 a35314a <=( (not A199)  and  a35313a );
 a35315a <=( a35314a  and  a35309a );
 a35319a <=( (not A267)  and  A265 );
 a35320a <=( A233  and  a35319a );
 a35324a <=( (not A302)  and  (not A301) );
 a35325a <=( (not A299)  and  a35324a );
 a35326a <=( a35325a  and  a35320a );
 a35330a <=( (not A166)  and  (not A167) );
 a35331a <=( (not A169)  and  a35330a );
 a35335a <=( A232  and  A200 );
 a35336a <=( (not A199)  and  a35335a );
 a35337a <=( a35336a  and  a35331a );
 a35341a <=( A266  and  A265 );
 a35342a <=( A233  and  a35341a );
 a35346a <=( (not A302)  and  (not A301) );
 a35347a <=( (not A299)  and  a35346a );
 a35348a <=( a35347a  and  a35342a );
 a35352a <=( (not A166)  and  (not A167) );
 a35353a <=( (not A169)  and  a35352a );
 a35357a <=( A232  and  A200 );
 a35358a <=( (not A199)  and  a35357a );
 a35359a <=( a35358a  and  a35353a );
 a35363a <=( (not A266)  and  (not A265) );
 a35364a <=( A233  and  a35363a );
 a35368a <=( (not A302)  and  (not A301) );
 a35369a <=( (not A299)  and  a35368a );
 a35370a <=( a35369a  and  a35364a );
 a35374a <=( (not A166)  and  (not A167) );
 a35375a <=( (not A169)  and  a35374a );
 a35379a <=( (not A233)  and  A200 );
 a35380a <=( (not A199)  and  a35379a );
 a35381a <=( a35380a  and  a35375a );
 a35385a <=( A265  and  (not A236) );
 a35386a <=( (not A235)  and  a35385a );
 a35390a <=( (not A300)  and  A298 );
 a35391a <=( A266  and  a35390a );
 a35392a <=( a35391a  and  a35386a );
 a35396a <=( (not A166)  and  (not A167) );
 a35397a <=( (not A169)  and  a35396a );
 a35401a <=( (not A233)  and  A200 );
 a35402a <=( (not A199)  and  a35401a );
 a35403a <=( a35402a  and  a35397a );
 a35407a <=( A265  and  (not A236) );
 a35408a <=( (not A235)  and  a35407a );
 a35412a <=( A299  and  A298 );
 a35413a <=( A266  and  a35412a );
 a35414a <=( a35413a  and  a35408a );
 a35418a <=( (not A166)  and  (not A167) );
 a35419a <=( (not A169)  and  a35418a );
 a35423a <=( (not A233)  and  A200 );
 a35424a <=( (not A199)  and  a35423a );
 a35425a <=( a35424a  and  a35419a );
 a35429a <=( A265  and  (not A236) );
 a35430a <=( (not A235)  and  a35429a );
 a35434a <=( (not A299)  and  (not A298) );
 a35435a <=( A266  and  a35434a );
 a35436a <=( a35435a  and  a35430a );
 a35440a <=( (not A166)  and  (not A167) );
 a35441a <=( (not A169)  and  a35440a );
 a35445a <=( (not A233)  and  A200 );
 a35446a <=( (not A199)  and  a35445a );
 a35447a <=( a35446a  and  a35441a );
 a35451a <=( (not A266)  and  (not A236) );
 a35452a <=( (not A235)  and  a35451a );
 a35456a <=( (not A300)  and  A298 );
 a35457a <=( (not A267)  and  a35456a );
 a35458a <=( a35457a  and  a35452a );
 a35462a <=( (not A166)  and  (not A167) );
 a35463a <=( (not A169)  and  a35462a );
 a35467a <=( (not A233)  and  A200 );
 a35468a <=( (not A199)  and  a35467a );
 a35469a <=( a35468a  and  a35463a );
 a35473a <=( (not A266)  and  (not A236) );
 a35474a <=( (not A235)  and  a35473a );
 a35478a <=( A299  and  A298 );
 a35479a <=( (not A267)  and  a35478a );
 a35480a <=( a35479a  and  a35474a );
 a35484a <=( (not A166)  and  (not A167) );
 a35485a <=( (not A169)  and  a35484a );
 a35489a <=( (not A233)  and  A200 );
 a35490a <=( (not A199)  and  a35489a );
 a35491a <=( a35490a  and  a35485a );
 a35495a <=( (not A266)  and  (not A236) );
 a35496a <=( (not A235)  and  a35495a );
 a35500a <=( (not A299)  and  (not A298) );
 a35501a <=( (not A267)  and  a35500a );
 a35502a <=( a35501a  and  a35496a );
 a35506a <=( (not A166)  and  (not A167) );
 a35507a <=( (not A169)  and  a35506a );
 a35511a <=( (not A233)  and  A200 );
 a35512a <=( (not A199)  and  a35511a );
 a35513a <=( a35512a  and  a35507a );
 a35517a <=( (not A265)  and  (not A236) );
 a35518a <=( (not A235)  and  a35517a );
 a35522a <=( (not A300)  and  A298 );
 a35523a <=( (not A266)  and  a35522a );
 a35524a <=( a35523a  and  a35518a );
 a35528a <=( (not A166)  and  (not A167) );
 a35529a <=( (not A169)  and  a35528a );
 a35533a <=( (not A233)  and  A200 );
 a35534a <=( (not A199)  and  a35533a );
 a35535a <=( a35534a  and  a35529a );
 a35539a <=( (not A265)  and  (not A236) );
 a35540a <=( (not A235)  and  a35539a );
 a35544a <=( A299  and  A298 );
 a35545a <=( (not A266)  and  a35544a );
 a35546a <=( a35545a  and  a35540a );
 a35550a <=( (not A166)  and  (not A167) );
 a35551a <=( (not A169)  and  a35550a );
 a35555a <=( (not A233)  and  A200 );
 a35556a <=( (not A199)  and  a35555a );
 a35557a <=( a35556a  and  a35551a );
 a35561a <=( (not A265)  and  (not A236) );
 a35562a <=( (not A235)  and  a35561a );
 a35566a <=( (not A299)  and  (not A298) );
 a35567a <=( (not A266)  and  a35566a );
 a35568a <=( a35567a  and  a35562a );
 a35572a <=( (not A166)  and  (not A167) );
 a35573a <=( (not A169)  and  a35572a );
 a35577a <=( (not A233)  and  A200 );
 a35578a <=( (not A199)  and  a35577a );
 a35579a <=( a35578a  and  a35573a );
 a35583a <=( A266  and  A265 );
 a35584a <=( (not A234)  and  a35583a );
 a35588a <=( (not A302)  and  (not A301) );
 a35589a <=( A298  and  a35588a );
 a35590a <=( a35589a  and  a35584a );
 a35594a <=( (not A166)  and  (not A167) );
 a35595a <=( (not A169)  and  a35594a );
 a35599a <=( (not A233)  and  A200 );
 a35600a <=( (not A199)  and  a35599a );
 a35601a <=( a35600a  and  a35595a );
 a35605a <=( (not A268)  and  (not A266) );
 a35606a <=( (not A234)  and  a35605a );
 a35610a <=( (not A300)  and  A298 );
 a35611a <=( (not A269)  and  a35610a );
 a35612a <=( a35611a  and  a35606a );
 a35616a <=( (not A166)  and  (not A167) );
 a35617a <=( (not A169)  and  a35616a );
 a35621a <=( (not A233)  and  A200 );
 a35622a <=( (not A199)  and  a35621a );
 a35623a <=( a35622a  and  a35617a );
 a35627a <=( (not A268)  and  (not A266) );
 a35628a <=( (not A234)  and  a35627a );
 a35632a <=( A299  and  A298 );
 a35633a <=( (not A269)  and  a35632a );
 a35634a <=( a35633a  and  a35628a );
 a35638a <=( (not A166)  and  (not A167) );
 a35639a <=( (not A169)  and  a35638a );
 a35643a <=( (not A233)  and  A200 );
 a35644a <=( (not A199)  and  a35643a );
 a35645a <=( a35644a  and  a35639a );
 a35649a <=( (not A268)  and  (not A266) );
 a35650a <=( (not A234)  and  a35649a );
 a35654a <=( (not A299)  and  (not A298) );
 a35655a <=( (not A269)  and  a35654a );
 a35656a <=( a35655a  and  a35650a );
 a35660a <=( (not A166)  and  (not A167) );
 a35661a <=( (not A169)  and  a35660a );
 a35665a <=( (not A233)  and  A200 );
 a35666a <=( (not A199)  and  a35665a );
 a35667a <=( a35666a  and  a35661a );
 a35671a <=( (not A267)  and  (not A266) );
 a35672a <=( (not A234)  and  a35671a );
 a35676a <=( (not A302)  and  (not A301) );
 a35677a <=( A298  and  a35676a );
 a35678a <=( a35677a  and  a35672a );
 a35682a <=( (not A166)  and  (not A167) );
 a35683a <=( (not A169)  and  a35682a );
 a35687a <=( (not A233)  and  A200 );
 a35688a <=( (not A199)  and  a35687a );
 a35689a <=( a35688a  and  a35683a );
 a35693a <=( (not A266)  and  (not A265) );
 a35694a <=( (not A234)  and  a35693a );
 a35698a <=( (not A302)  and  (not A301) );
 a35699a <=( A298  and  a35698a );
 a35700a <=( a35699a  and  a35694a );
 a35704a <=( (not A166)  and  (not A167) );
 a35705a <=( (not A169)  and  a35704a );
 a35709a <=( (not A232)  and  A200 );
 a35710a <=( (not A199)  and  a35709a );
 a35711a <=( a35710a  and  a35705a );
 a35715a <=( A266  and  A265 );
 a35716a <=( (not A233)  and  a35715a );
 a35720a <=( (not A302)  and  (not A301) );
 a35721a <=( A298  and  a35720a );
 a35722a <=( a35721a  and  a35716a );
 a35726a <=( (not A166)  and  (not A167) );
 a35727a <=( (not A169)  and  a35726a );
 a35731a <=( (not A232)  and  A200 );
 a35732a <=( (not A199)  and  a35731a );
 a35733a <=( a35732a  and  a35727a );
 a35737a <=( (not A268)  and  (not A266) );
 a35738a <=( (not A233)  and  a35737a );
 a35742a <=( (not A300)  and  A298 );
 a35743a <=( (not A269)  and  a35742a );
 a35744a <=( a35743a  and  a35738a );
 a35748a <=( (not A166)  and  (not A167) );
 a35749a <=( (not A169)  and  a35748a );
 a35753a <=( (not A232)  and  A200 );
 a35754a <=( (not A199)  and  a35753a );
 a35755a <=( a35754a  and  a35749a );
 a35759a <=( (not A268)  and  (not A266) );
 a35760a <=( (not A233)  and  a35759a );
 a35764a <=( A299  and  A298 );
 a35765a <=( (not A269)  and  a35764a );
 a35766a <=( a35765a  and  a35760a );
 a35770a <=( (not A166)  and  (not A167) );
 a35771a <=( (not A169)  and  a35770a );
 a35775a <=( (not A232)  and  A200 );
 a35776a <=( (not A199)  and  a35775a );
 a35777a <=( a35776a  and  a35771a );
 a35781a <=( (not A268)  and  (not A266) );
 a35782a <=( (not A233)  and  a35781a );
 a35786a <=( (not A299)  and  (not A298) );
 a35787a <=( (not A269)  and  a35786a );
 a35788a <=( a35787a  and  a35782a );
 a35792a <=( (not A166)  and  (not A167) );
 a35793a <=( (not A169)  and  a35792a );
 a35797a <=( (not A232)  and  A200 );
 a35798a <=( (not A199)  and  a35797a );
 a35799a <=( a35798a  and  a35793a );
 a35803a <=( (not A267)  and  (not A266) );
 a35804a <=( (not A233)  and  a35803a );
 a35808a <=( (not A302)  and  (not A301) );
 a35809a <=( A298  and  a35808a );
 a35810a <=( a35809a  and  a35804a );
 a35814a <=( (not A166)  and  (not A167) );
 a35815a <=( (not A169)  and  a35814a );
 a35819a <=( (not A232)  and  A200 );
 a35820a <=( (not A199)  and  a35819a );
 a35821a <=( a35820a  and  a35815a );
 a35825a <=( (not A266)  and  (not A265) );
 a35826a <=( (not A233)  and  a35825a );
 a35830a <=( (not A302)  and  (not A301) );
 a35831a <=( A298  and  a35830a );
 a35832a <=( a35831a  and  a35826a );
 a35836a <=( A167  and  (not A168) );
 a35837a <=( (not A169)  and  a35836a );
 a35841a <=( A200  and  (not A199) );
 a35842a <=( A166  and  a35841a );
 a35843a <=( a35842a  and  a35837a );
 a35847a <=( A265  and  A233 );
 a35848a <=( A232  and  a35847a );
 a35852a <=( (not A300)  and  (not A299) );
 a35853a <=( (not A267)  and  a35852a );
 a35854a <=( a35853a  and  a35848a );
 a35858a <=( A167  and  (not A168) );
 a35859a <=( (not A169)  and  a35858a );
 a35863a <=( A200  and  (not A199) );
 a35864a <=( A166  and  a35863a );
 a35865a <=( a35864a  and  a35859a );
 a35869a <=( A265  and  A233 );
 a35870a <=( A232  and  a35869a );
 a35874a <=( A299  and  A298 );
 a35875a <=( (not A267)  and  a35874a );
 a35876a <=( a35875a  and  a35870a );
 a35880a <=( A167  and  (not A168) );
 a35881a <=( (not A169)  and  a35880a );
 a35885a <=( A200  and  (not A199) );
 a35886a <=( A166  and  a35885a );
 a35887a <=( a35886a  and  a35881a );
 a35891a <=( A265  and  A233 );
 a35892a <=( A232  and  a35891a );
 a35896a <=( (not A299)  and  (not A298) );
 a35897a <=( (not A267)  and  a35896a );
 a35898a <=( a35897a  and  a35892a );
 a35902a <=( A167  and  (not A168) );
 a35903a <=( (not A169)  and  a35902a );
 a35907a <=( A200  and  (not A199) );
 a35908a <=( A166  and  a35907a );
 a35909a <=( a35908a  and  a35903a );
 a35913a <=( A265  and  A233 );
 a35914a <=( A232  and  a35913a );
 a35918a <=( (not A300)  and  (not A299) );
 a35919a <=( A266  and  a35918a );
 a35920a <=( a35919a  and  a35914a );
 a35924a <=( A167  and  (not A168) );
 a35925a <=( (not A169)  and  a35924a );
 a35929a <=( A200  and  (not A199) );
 a35930a <=( A166  and  a35929a );
 a35931a <=( a35930a  and  a35925a );
 a35935a <=( A265  and  A233 );
 a35936a <=( A232  and  a35935a );
 a35940a <=( A299  and  A298 );
 a35941a <=( A266  and  a35940a );
 a35942a <=( a35941a  and  a35936a );
 a35946a <=( A167  and  (not A168) );
 a35947a <=( (not A169)  and  a35946a );
 a35951a <=( A200  and  (not A199) );
 a35952a <=( A166  and  a35951a );
 a35953a <=( a35952a  and  a35947a );
 a35957a <=( A265  and  A233 );
 a35958a <=( A232  and  a35957a );
 a35962a <=( (not A299)  and  (not A298) );
 a35963a <=( A266  and  a35962a );
 a35964a <=( a35963a  and  a35958a );
 a35968a <=( A167  and  (not A168) );
 a35969a <=( (not A169)  and  a35968a );
 a35973a <=( A200  and  (not A199) );
 a35974a <=( A166  and  a35973a );
 a35975a <=( a35974a  and  a35969a );
 a35979a <=( (not A265)  and  A233 );
 a35980a <=( A232  and  a35979a );
 a35984a <=( (not A300)  and  (not A299) );
 a35985a <=( (not A266)  and  a35984a );
 a35986a <=( a35985a  and  a35980a );
 a35990a <=( A167  and  (not A168) );
 a35991a <=( (not A169)  and  a35990a );
 a35995a <=( A200  and  (not A199) );
 a35996a <=( A166  and  a35995a );
 a35997a <=( a35996a  and  a35991a );
 a36001a <=( (not A265)  and  A233 );
 a36002a <=( A232  and  a36001a );
 a36006a <=( A299  and  A298 );
 a36007a <=( (not A266)  and  a36006a );
 a36008a <=( a36007a  and  a36002a );
 a36012a <=( A167  and  (not A168) );
 a36013a <=( (not A169)  and  a36012a );
 a36017a <=( A200  and  (not A199) );
 a36018a <=( A166  and  a36017a );
 a36019a <=( a36018a  and  a36013a );
 a36023a <=( (not A265)  and  A233 );
 a36024a <=( A232  and  a36023a );
 a36028a <=( (not A299)  and  (not A298) );
 a36029a <=( (not A266)  and  a36028a );
 a36030a <=( a36029a  and  a36024a );
 a36034a <=( A167  and  (not A168) );
 a36035a <=( (not A169)  and  a36034a );
 a36039a <=( A200  and  (not A199) );
 a36040a <=( A166  and  a36039a );
 a36041a <=( a36040a  and  a36035a );
 a36045a <=( A298  and  A233 );
 a36046a <=( (not A232)  and  a36045a );
 a36050a <=( A301  and  A300 );
 a36051a <=( (not A299)  and  a36050a );
 a36052a <=( a36051a  and  a36046a );
 a36056a <=( A167  and  (not A168) );
 a36057a <=( (not A169)  and  a36056a );
 a36061a <=( A200  and  (not A199) );
 a36062a <=( A166  and  a36061a );
 a36063a <=( a36062a  and  a36057a );
 a36067a <=( A298  and  A233 );
 a36068a <=( (not A232)  and  a36067a );
 a36072a <=( A302  and  A300 );
 a36073a <=( (not A299)  and  a36072a );
 a36074a <=( a36073a  and  a36068a );
 a36078a <=( A167  and  (not A168) );
 a36079a <=( (not A169)  and  a36078a );
 a36083a <=( A200  and  (not A199) );
 a36084a <=( A166  and  a36083a );
 a36085a <=( a36084a  and  a36079a );
 a36089a <=( A265  and  A233 );
 a36090a <=( (not A232)  and  a36089a );
 a36094a <=( A268  and  A267 );
 a36095a <=( (not A266)  and  a36094a );
 a36096a <=( a36095a  and  a36090a );
 a36100a <=( A167  and  (not A168) );
 a36101a <=( (not A169)  and  a36100a );
 a36105a <=( A200  and  (not A199) );
 a36106a <=( A166  and  a36105a );
 a36107a <=( a36106a  and  a36101a );
 a36111a <=( A265  and  A233 );
 a36112a <=( (not A232)  and  a36111a );
 a36116a <=( A269  and  A267 );
 a36117a <=( (not A266)  and  a36116a );
 a36118a <=( a36117a  and  a36112a );
 a36122a <=( A167  and  (not A168) );
 a36123a <=( (not A169)  and  a36122a );
 a36127a <=( A200  and  (not A199) );
 a36128a <=( A166  and  a36127a );
 a36129a <=( a36128a  and  a36123a );
 a36133a <=( A265  and  (not A234) );
 a36134a <=( (not A233)  and  a36133a );
 a36138a <=( (not A300)  and  A298 );
 a36139a <=( A266  and  a36138a );
 a36140a <=( a36139a  and  a36134a );
 a36144a <=( A167  and  (not A168) );
 a36145a <=( (not A169)  and  a36144a );
 a36149a <=( A200  and  (not A199) );
 a36150a <=( A166  and  a36149a );
 a36151a <=( a36150a  and  a36145a );
 a36155a <=( A265  and  (not A234) );
 a36156a <=( (not A233)  and  a36155a );
 a36160a <=( A299  and  A298 );
 a36161a <=( A266  and  a36160a );
 a36162a <=( a36161a  and  a36156a );
 a36166a <=( A167  and  (not A168) );
 a36167a <=( (not A169)  and  a36166a );
 a36171a <=( A200  and  (not A199) );
 a36172a <=( A166  and  a36171a );
 a36173a <=( a36172a  and  a36167a );
 a36177a <=( A265  and  (not A234) );
 a36178a <=( (not A233)  and  a36177a );
 a36182a <=( (not A299)  and  (not A298) );
 a36183a <=( A266  and  a36182a );
 a36184a <=( a36183a  and  a36178a );
 a36188a <=( A167  and  (not A168) );
 a36189a <=( (not A169)  and  a36188a );
 a36193a <=( A200  and  (not A199) );
 a36194a <=( A166  and  a36193a );
 a36195a <=( a36194a  and  a36189a );
 a36199a <=( (not A266)  and  (not A234) );
 a36200a <=( (not A233)  and  a36199a );
 a36204a <=( (not A300)  and  A298 );
 a36205a <=( (not A267)  and  a36204a );
 a36206a <=( a36205a  and  a36200a );
 a36210a <=( A167  and  (not A168) );
 a36211a <=( (not A169)  and  a36210a );
 a36215a <=( A200  and  (not A199) );
 a36216a <=( A166  and  a36215a );
 a36217a <=( a36216a  and  a36211a );
 a36221a <=( (not A266)  and  (not A234) );
 a36222a <=( (not A233)  and  a36221a );
 a36226a <=( A299  and  A298 );
 a36227a <=( (not A267)  and  a36226a );
 a36228a <=( a36227a  and  a36222a );
 a36232a <=( A167  and  (not A168) );
 a36233a <=( (not A169)  and  a36232a );
 a36237a <=( A200  and  (not A199) );
 a36238a <=( A166  and  a36237a );
 a36239a <=( a36238a  and  a36233a );
 a36243a <=( (not A266)  and  (not A234) );
 a36244a <=( (not A233)  and  a36243a );
 a36248a <=( (not A299)  and  (not A298) );
 a36249a <=( (not A267)  and  a36248a );
 a36250a <=( a36249a  and  a36244a );
 a36254a <=( A167  and  (not A168) );
 a36255a <=( (not A169)  and  a36254a );
 a36259a <=( A200  and  (not A199) );
 a36260a <=( A166  and  a36259a );
 a36261a <=( a36260a  and  a36255a );
 a36265a <=( (not A265)  and  (not A234) );
 a36266a <=( (not A233)  and  a36265a );
 a36270a <=( (not A300)  and  A298 );
 a36271a <=( (not A266)  and  a36270a );
 a36272a <=( a36271a  and  a36266a );
 a36276a <=( A167  and  (not A168) );
 a36277a <=( (not A169)  and  a36276a );
 a36281a <=( A200  and  (not A199) );
 a36282a <=( A166  and  a36281a );
 a36283a <=( a36282a  and  a36277a );
 a36287a <=( (not A265)  and  (not A234) );
 a36288a <=( (not A233)  and  a36287a );
 a36292a <=( A299  and  A298 );
 a36293a <=( (not A266)  and  a36292a );
 a36294a <=( a36293a  and  a36288a );
 a36298a <=( A167  and  (not A168) );
 a36299a <=( (not A169)  and  a36298a );
 a36303a <=( A200  and  (not A199) );
 a36304a <=( A166  and  a36303a );
 a36305a <=( a36304a  and  a36299a );
 a36309a <=( (not A265)  and  (not A234) );
 a36310a <=( (not A233)  and  a36309a );
 a36314a <=( (not A299)  and  (not A298) );
 a36315a <=( (not A266)  and  a36314a );
 a36316a <=( a36315a  and  a36310a );
 a36320a <=( A167  and  (not A168) );
 a36321a <=( (not A169)  and  a36320a );
 a36325a <=( A200  and  (not A199) );
 a36326a <=( A166  and  a36325a );
 a36327a <=( a36326a  and  a36321a );
 a36331a <=( A234  and  (not A233) );
 a36332a <=( A232  and  a36331a );
 a36336a <=( A299  and  (not A298) );
 a36337a <=( A235  and  a36336a );
 a36338a <=( a36337a  and  a36332a );
 a36342a <=( A167  and  (not A168) );
 a36343a <=( (not A169)  and  a36342a );
 a36347a <=( A200  and  (not A199) );
 a36348a <=( A166  and  a36347a );
 a36349a <=( a36348a  and  a36343a );
 a36353a <=( A234  and  (not A233) );
 a36354a <=( A232  and  a36353a );
 a36358a <=( A266  and  (not A265) );
 a36359a <=( A235  and  a36358a );
 a36360a <=( a36359a  and  a36354a );
 a36364a <=( A167  and  (not A168) );
 a36365a <=( (not A169)  and  a36364a );
 a36369a <=( A200  and  (not A199) );
 a36370a <=( A166  and  a36369a );
 a36371a <=( a36370a  and  a36365a );
 a36375a <=( A234  and  (not A233) );
 a36376a <=( A232  and  a36375a );
 a36380a <=( A299  and  (not A298) );
 a36381a <=( A236  and  a36380a );
 a36382a <=( a36381a  and  a36376a );
 a36386a <=( A167  and  (not A168) );
 a36387a <=( (not A169)  and  a36386a );
 a36391a <=( A200  and  (not A199) );
 a36392a <=( A166  and  a36391a );
 a36393a <=( a36392a  and  a36387a );
 a36397a <=( A234  and  (not A233) );
 a36398a <=( A232  and  a36397a );
 a36402a <=( A266  and  (not A265) );
 a36403a <=( A236  and  a36402a );
 a36404a <=( a36403a  and  a36398a );
 a36408a <=( A167  and  (not A168) );
 a36409a <=( (not A169)  and  a36408a );
 a36413a <=( A200  and  (not A199) );
 a36414a <=( A166  and  a36413a );
 a36415a <=( a36414a  and  a36409a );
 a36419a <=( A265  and  (not A233) );
 a36420a <=( (not A232)  and  a36419a );
 a36424a <=( (not A300)  and  A298 );
 a36425a <=( A266  and  a36424a );
 a36426a <=( a36425a  and  a36420a );
 a36430a <=( A167  and  (not A168) );
 a36431a <=( (not A169)  and  a36430a );
 a36435a <=( A200  and  (not A199) );
 a36436a <=( A166  and  a36435a );
 a36437a <=( a36436a  and  a36431a );
 a36441a <=( A265  and  (not A233) );
 a36442a <=( (not A232)  and  a36441a );
 a36446a <=( A299  and  A298 );
 a36447a <=( A266  and  a36446a );
 a36448a <=( a36447a  and  a36442a );
 a36452a <=( A167  and  (not A168) );
 a36453a <=( (not A169)  and  a36452a );
 a36457a <=( A200  and  (not A199) );
 a36458a <=( A166  and  a36457a );
 a36459a <=( a36458a  and  a36453a );
 a36463a <=( A265  and  (not A233) );
 a36464a <=( (not A232)  and  a36463a );
 a36468a <=( (not A299)  and  (not A298) );
 a36469a <=( A266  and  a36468a );
 a36470a <=( a36469a  and  a36464a );
 a36474a <=( A167  and  (not A168) );
 a36475a <=( (not A169)  and  a36474a );
 a36479a <=( A200  and  (not A199) );
 a36480a <=( A166  and  a36479a );
 a36481a <=( a36480a  and  a36475a );
 a36485a <=( (not A266)  and  (not A233) );
 a36486a <=( (not A232)  and  a36485a );
 a36490a <=( (not A300)  and  A298 );
 a36491a <=( (not A267)  and  a36490a );
 a36492a <=( a36491a  and  a36486a );
 a36496a <=( A167  and  (not A168) );
 a36497a <=( (not A169)  and  a36496a );
 a36501a <=( A200  and  (not A199) );
 a36502a <=( A166  and  a36501a );
 a36503a <=( a36502a  and  a36497a );
 a36507a <=( (not A266)  and  (not A233) );
 a36508a <=( (not A232)  and  a36507a );
 a36512a <=( A299  and  A298 );
 a36513a <=( (not A267)  and  a36512a );
 a36514a <=( a36513a  and  a36508a );
 a36518a <=( A167  and  (not A168) );
 a36519a <=( (not A169)  and  a36518a );
 a36523a <=( A200  and  (not A199) );
 a36524a <=( A166  and  a36523a );
 a36525a <=( a36524a  and  a36519a );
 a36529a <=( (not A266)  and  (not A233) );
 a36530a <=( (not A232)  and  a36529a );
 a36534a <=( (not A299)  and  (not A298) );
 a36535a <=( (not A267)  and  a36534a );
 a36536a <=( a36535a  and  a36530a );
 a36540a <=( A167  and  (not A168) );
 a36541a <=( (not A169)  and  a36540a );
 a36545a <=( A200  and  (not A199) );
 a36546a <=( A166  and  a36545a );
 a36547a <=( a36546a  and  a36541a );
 a36551a <=( (not A265)  and  (not A233) );
 a36552a <=( (not A232)  and  a36551a );
 a36556a <=( (not A300)  and  A298 );
 a36557a <=( (not A266)  and  a36556a );
 a36558a <=( a36557a  and  a36552a );
 a36562a <=( A167  and  (not A168) );
 a36563a <=( (not A169)  and  a36562a );
 a36567a <=( A200  and  (not A199) );
 a36568a <=( A166  and  a36567a );
 a36569a <=( a36568a  and  a36563a );
 a36573a <=( (not A265)  and  (not A233) );
 a36574a <=( (not A232)  and  a36573a );
 a36578a <=( A299  and  A298 );
 a36579a <=( (not A266)  and  a36578a );
 a36580a <=( a36579a  and  a36574a );
 a36584a <=( A167  and  (not A168) );
 a36585a <=( (not A169)  and  a36584a );
 a36589a <=( A200  and  (not A199) );
 a36590a <=( A166  and  a36589a );
 a36591a <=( a36590a  and  a36585a );
 a36595a <=( (not A265)  and  (not A233) );
 a36596a <=( (not A232)  and  a36595a );
 a36600a <=( (not A299)  and  (not A298) );
 a36601a <=( (not A266)  and  a36600a );
 a36602a <=( a36601a  and  a36596a );
 a36606a <=( A167  and  (not A168) );
 a36607a <=( (not A169)  and  a36606a );
 a36611a <=( (not A200)  and  A199 );
 a36612a <=( A166  and  a36611a );
 a36613a <=( a36612a  and  a36607a );
 a36617a <=( (not A232)  and  A202 );
 a36618a <=( A201  and  a36617a );
 a36622a <=( A299  and  (not A298) );
 a36623a <=( A233  and  a36622a );
 a36624a <=( a36623a  and  a36618a );
 a36628a <=( A167  and  (not A168) );
 a36629a <=( (not A169)  and  a36628a );
 a36633a <=( (not A200)  and  A199 );
 a36634a <=( A166  and  a36633a );
 a36635a <=( a36634a  and  a36629a );
 a36639a <=( (not A232)  and  A202 );
 a36640a <=( A201  and  a36639a );
 a36644a <=( A266  and  (not A265) );
 a36645a <=( A233  and  a36644a );
 a36646a <=( a36645a  and  a36640a );
 a36650a <=( A167  and  (not A168) );
 a36651a <=( (not A169)  and  a36650a );
 a36655a <=( (not A200)  and  A199 );
 a36656a <=( A166  and  a36655a );
 a36657a <=( a36656a  and  a36651a );
 a36661a <=( (not A232)  and  A203 );
 a36662a <=( A201  and  a36661a );
 a36666a <=( A299  and  (not A298) );
 a36667a <=( A233  and  a36666a );
 a36668a <=( a36667a  and  a36662a );
 a36672a <=( A167  and  (not A168) );
 a36673a <=( (not A169)  and  a36672a );
 a36677a <=( (not A200)  and  A199 );
 a36678a <=( A166  and  a36677a );
 a36679a <=( a36678a  and  a36673a );
 a36683a <=( (not A232)  and  A203 );
 a36684a <=( A201  and  a36683a );
 a36688a <=( A266  and  (not A265) );
 a36689a <=( A233  and  a36688a );
 a36690a <=( a36689a  and  a36684a );
 a36694a <=( A167  and  (not A169) );
 a36695a <=( A170  and  a36694a );
 a36699a <=( A200  and  A199 );
 a36700a <=( (not A166)  and  a36699a );
 a36701a <=( a36700a  and  a36695a );
 a36705a <=( A265  and  A233 );
 a36706a <=( A232  and  a36705a );
 a36710a <=( (not A300)  and  (not A299) );
 a36711a <=( (not A267)  and  a36710a );
 a36712a <=( a36711a  and  a36706a );
 a36716a <=( A167  and  (not A169) );
 a36717a <=( A170  and  a36716a );
 a36721a <=( A200  and  A199 );
 a36722a <=( (not A166)  and  a36721a );
 a36723a <=( a36722a  and  a36717a );
 a36727a <=( A265  and  A233 );
 a36728a <=( A232  and  a36727a );
 a36732a <=( A299  and  A298 );
 a36733a <=( (not A267)  and  a36732a );
 a36734a <=( a36733a  and  a36728a );
 a36738a <=( A167  and  (not A169) );
 a36739a <=( A170  and  a36738a );
 a36743a <=( A200  and  A199 );
 a36744a <=( (not A166)  and  a36743a );
 a36745a <=( a36744a  and  a36739a );
 a36749a <=( A265  and  A233 );
 a36750a <=( A232  and  a36749a );
 a36754a <=( (not A299)  and  (not A298) );
 a36755a <=( (not A267)  and  a36754a );
 a36756a <=( a36755a  and  a36750a );
 a36760a <=( A167  and  (not A169) );
 a36761a <=( A170  and  a36760a );
 a36765a <=( A200  and  A199 );
 a36766a <=( (not A166)  and  a36765a );
 a36767a <=( a36766a  and  a36761a );
 a36771a <=( A265  and  A233 );
 a36772a <=( A232  and  a36771a );
 a36776a <=( (not A300)  and  (not A299) );
 a36777a <=( A266  and  a36776a );
 a36778a <=( a36777a  and  a36772a );
 a36782a <=( A167  and  (not A169) );
 a36783a <=( A170  and  a36782a );
 a36787a <=( A200  and  A199 );
 a36788a <=( (not A166)  and  a36787a );
 a36789a <=( a36788a  and  a36783a );
 a36793a <=( A265  and  A233 );
 a36794a <=( A232  and  a36793a );
 a36798a <=( A299  and  A298 );
 a36799a <=( A266  and  a36798a );
 a36800a <=( a36799a  and  a36794a );
 a36804a <=( A167  and  (not A169) );
 a36805a <=( A170  and  a36804a );
 a36809a <=( A200  and  A199 );
 a36810a <=( (not A166)  and  a36809a );
 a36811a <=( a36810a  and  a36805a );
 a36815a <=( A265  and  A233 );
 a36816a <=( A232  and  a36815a );
 a36820a <=( (not A299)  and  (not A298) );
 a36821a <=( A266  and  a36820a );
 a36822a <=( a36821a  and  a36816a );
 a36826a <=( A167  and  (not A169) );
 a36827a <=( A170  and  a36826a );
 a36831a <=( A200  and  A199 );
 a36832a <=( (not A166)  and  a36831a );
 a36833a <=( a36832a  and  a36827a );
 a36837a <=( (not A265)  and  A233 );
 a36838a <=( A232  and  a36837a );
 a36842a <=( (not A300)  and  (not A299) );
 a36843a <=( (not A266)  and  a36842a );
 a36844a <=( a36843a  and  a36838a );
 a36848a <=( A167  and  (not A169) );
 a36849a <=( A170  and  a36848a );
 a36853a <=( A200  and  A199 );
 a36854a <=( (not A166)  and  a36853a );
 a36855a <=( a36854a  and  a36849a );
 a36859a <=( (not A265)  and  A233 );
 a36860a <=( A232  and  a36859a );
 a36864a <=( A299  and  A298 );
 a36865a <=( (not A266)  and  a36864a );
 a36866a <=( a36865a  and  a36860a );
 a36870a <=( A167  and  (not A169) );
 a36871a <=( A170  and  a36870a );
 a36875a <=( A200  and  A199 );
 a36876a <=( (not A166)  and  a36875a );
 a36877a <=( a36876a  and  a36871a );
 a36881a <=( (not A265)  and  A233 );
 a36882a <=( A232  and  a36881a );
 a36886a <=( (not A299)  and  (not A298) );
 a36887a <=( (not A266)  and  a36886a );
 a36888a <=( a36887a  and  a36882a );
 a36892a <=( A167  and  (not A169) );
 a36893a <=( A170  and  a36892a );
 a36897a <=( A200  and  A199 );
 a36898a <=( (not A166)  and  a36897a );
 a36899a <=( a36898a  and  a36893a );
 a36903a <=( A298  and  A233 );
 a36904a <=( (not A232)  and  a36903a );
 a36908a <=( A301  and  A300 );
 a36909a <=( (not A299)  and  a36908a );
 a36910a <=( a36909a  and  a36904a );
 a36914a <=( A167  and  (not A169) );
 a36915a <=( A170  and  a36914a );
 a36919a <=( A200  and  A199 );
 a36920a <=( (not A166)  and  a36919a );
 a36921a <=( a36920a  and  a36915a );
 a36925a <=( A298  and  A233 );
 a36926a <=( (not A232)  and  a36925a );
 a36930a <=( A302  and  A300 );
 a36931a <=( (not A299)  and  a36930a );
 a36932a <=( a36931a  and  a36926a );
 a36936a <=( A167  and  (not A169) );
 a36937a <=( A170  and  a36936a );
 a36941a <=( A200  and  A199 );
 a36942a <=( (not A166)  and  a36941a );
 a36943a <=( a36942a  and  a36937a );
 a36947a <=( A265  and  A233 );
 a36948a <=( (not A232)  and  a36947a );
 a36952a <=( A268  and  A267 );
 a36953a <=( (not A266)  and  a36952a );
 a36954a <=( a36953a  and  a36948a );
 a36958a <=( A167  and  (not A169) );
 a36959a <=( A170  and  a36958a );
 a36963a <=( A200  and  A199 );
 a36964a <=( (not A166)  and  a36963a );
 a36965a <=( a36964a  and  a36959a );
 a36969a <=( A265  and  A233 );
 a36970a <=( (not A232)  and  a36969a );
 a36974a <=( A269  and  A267 );
 a36975a <=( (not A266)  and  a36974a );
 a36976a <=( a36975a  and  a36970a );
 a36980a <=( A167  and  (not A169) );
 a36981a <=( A170  and  a36980a );
 a36985a <=( A200  and  A199 );
 a36986a <=( (not A166)  and  a36985a );
 a36987a <=( a36986a  and  a36981a );
 a36991a <=( A265  and  (not A234) );
 a36992a <=( (not A233)  and  a36991a );
 a36996a <=( (not A300)  and  A298 );
 a36997a <=( A266  and  a36996a );
 a36998a <=( a36997a  and  a36992a );
 a37002a <=( A167  and  (not A169) );
 a37003a <=( A170  and  a37002a );
 a37007a <=( A200  and  A199 );
 a37008a <=( (not A166)  and  a37007a );
 a37009a <=( a37008a  and  a37003a );
 a37013a <=( A265  and  (not A234) );
 a37014a <=( (not A233)  and  a37013a );
 a37018a <=( A299  and  A298 );
 a37019a <=( A266  and  a37018a );
 a37020a <=( a37019a  and  a37014a );
 a37024a <=( A167  and  (not A169) );
 a37025a <=( A170  and  a37024a );
 a37029a <=( A200  and  A199 );
 a37030a <=( (not A166)  and  a37029a );
 a37031a <=( a37030a  and  a37025a );
 a37035a <=( A265  and  (not A234) );
 a37036a <=( (not A233)  and  a37035a );
 a37040a <=( (not A299)  and  (not A298) );
 a37041a <=( A266  and  a37040a );
 a37042a <=( a37041a  and  a37036a );
 a37046a <=( A167  and  (not A169) );
 a37047a <=( A170  and  a37046a );
 a37051a <=( A200  and  A199 );
 a37052a <=( (not A166)  and  a37051a );
 a37053a <=( a37052a  and  a37047a );
 a37057a <=( (not A266)  and  (not A234) );
 a37058a <=( (not A233)  and  a37057a );
 a37062a <=( (not A300)  and  A298 );
 a37063a <=( (not A267)  and  a37062a );
 a37064a <=( a37063a  and  a37058a );
 a37068a <=( A167  and  (not A169) );
 a37069a <=( A170  and  a37068a );
 a37073a <=( A200  and  A199 );
 a37074a <=( (not A166)  and  a37073a );
 a37075a <=( a37074a  and  a37069a );
 a37079a <=( (not A266)  and  (not A234) );
 a37080a <=( (not A233)  and  a37079a );
 a37084a <=( A299  and  A298 );
 a37085a <=( (not A267)  and  a37084a );
 a37086a <=( a37085a  and  a37080a );
 a37090a <=( A167  and  (not A169) );
 a37091a <=( A170  and  a37090a );
 a37095a <=( A200  and  A199 );
 a37096a <=( (not A166)  and  a37095a );
 a37097a <=( a37096a  and  a37091a );
 a37101a <=( (not A266)  and  (not A234) );
 a37102a <=( (not A233)  and  a37101a );
 a37106a <=( (not A299)  and  (not A298) );
 a37107a <=( (not A267)  and  a37106a );
 a37108a <=( a37107a  and  a37102a );
 a37112a <=( A167  and  (not A169) );
 a37113a <=( A170  and  a37112a );
 a37117a <=( A200  and  A199 );
 a37118a <=( (not A166)  and  a37117a );
 a37119a <=( a37118a  and  a37113a );
 a37123a <=( (not A265)  and  (not A234) );
 a37124a <=( (not A233)  and  a37123a );
 a37128a <=( (not A300)  and  A298 );
 a37129a <=( (not A266)  and  a37128a );
 a37130a <=( a37129a  and  a37124a );
 a37134a <=( A167  and  (not A169) );
 a37135a <=( A170  and  a37134a );
 a37139a <=( A200  and  A199 );
 a37140a <=( (not A166)  and  a37139a );
 a37141a <=( a37140a  and  a37135a );
 a37145a <=( (not A265)  and  (not A234) );
 a37146a <=( (not A233)  and  a37145a );
 a37150a <=( A299  and  A298 );
 a37151a <=( (not A266)  and  a37150a );
 a37152a <=( a37151a  and  a37146a );
 a37156a <=( A167  and  (not A169) );
 a37157a <=( A170  and  a37156a );
 a37161a <=( A200  and  A199 );
 a37162a <=( (not A166)  and  a37161a );
 a37163a <=( a37162a  and  a37157a );
 a37167a <=( (not A265)  and  (not A234) );
 a37168a <=( (not A233)  and  a37167a );
 a37172a <=( (not A299)  and  (not A298) );
 a37173a <=( (not A266)  and  a37172a );
 a37174a <=( a37173a  and  a37168a );
 a37178a <=( A167  and  (not A169) );
 a37179a <=( A170  and  a37178a );
 a37183a <=( A200  and  A199 );
 a37184a <=( (not A166)  and  a37183a );
 a37185a <=( a37184a  and  a37179a );
 a37189a <=( A234  and  (not A233) );
 a37190a <=( A232  and  a37189a );
 a37194a <=( A299  and  (not A298) );
 a37195a <=( A235  and  a37194a );
 a37196a <=( a37195a  and  a37190a );
 a37200a <=( A167  and  (not A169) );
 a37201a <=( A170  and  a37200a );
 a37205a <=( A200  and  A199 );
 a37206a <=( (not A166)  and  a37205a );
 a37207a <=( a37206a  and  a37201a );
 a37211a <=( A234  and  (not A233) );
 a37212a <=( A232  and  a37211a );
 a37216a <=( A266  and  (not A265) );
 a37217a <=( A235  and  a37216a );
 a37218a <=( a37217a  and  a37212a );
 a37222a <=( A167  and  (not A169) );
 a37223a <=( A170  and  a37222a );
 a37227a <=( A200  and  A199 );
 a37228a <=( (not A166)  and  a37227a );
 a37229a <=( a37228a  and  a37223a );
 a37233a <=( A234  and  (not A233) );
 a37234a <=( A232  and  a37233a );
 a37238a <=( A299  and  (not A298) );
 a37239a <=( A236  and  a37238a );
 a37240a <=( a37239a  and  a37234a );
 a37244a <=( A167  and  (not A169) );
 a37245a <=( A170  and  a37244a );
 a37249a <=( A200  and  A199 );
 a37250a <=( (not A166)  and  a37249a );
 a37251a <=( a37250a  and  a37245a );
 a37255a <=( A234  and  (not A233) );
 a37256a <=( A232  and  a37255a );
 a37260a <=( A266  and  (not A265) );
 a37261a <=( A236  and  a37260a );
 a37262a <=( a37261a  and  a37256a );
 a37266a <=( A167  and  (not A169) );
 a37267a <=( A170  and  a37266a );
 a37271a <=( A200  and  A199 );
 a37272a <=( (not A166)  and  a37271a );
 a37273a <=( a37272a  and  a37267a );
 a37277a <=( A265  and  (not A233) );
 a37278a <=( (not A232)  and  a37277a );
 a37282a <=( (not A300)  and  A298 );
 a37283a <=( A266  and  a37282a );
 a37284a <=( a37283a  and  a37278a );
 a37288a <=( A167  and  (not A169) );
 a37289a <=( A170  and  a37288a );
 a37293a <=( A200  and  A199 );
 a37294a <=( (not A166)  and  a37293a );
 a37295a <=( a37294a  and  a37289a );
 a37299a <=( A265  and  (not A233) );
 a37300a <=( (not A232)  and  a37299a );
 a37304a <=( A299  and  A298 );
 a37305a <=( A266  and  a37304a );
 a37306a <=( a37305a  and  a37300a );
 a37310a <=( A167  and  (not A169) );
 a37311a <=( A170  and  a37310a );
 a37315a <=( A200  and  A199 );
 a37316a <=( (not A166)  and  a37315a );
 a37317a <=( a37316a  and  a37311a );
 a37321a <=( A265  and  (not A233) );
 a37322a <=( (not A232)  and  a37321a );
 a37326a <=( (not A299)  and  (not A298) );
 a37327a <=( A266  and  a37326a );
 a37328a <=( a37327a  and  a37322a );
 a37332a <=( A167  and  (not A169) );
 a37333a <=( A170  and  a37332a );
 a37337a <=( A200  and  A199 );
 a37338a <=( (not A166)  and  a37337a );
 a37339a <=( a37338a  and  a37333a );
 a37343a <=( (not A266)  and  (not A233) );
 a37344a <=( (not A232)  and  a37343a );
 a37348a <=( (not A300)  and  A298 );
 a37349a <=( (not A267)  and  a37348a );
 a37350a <=( a37349a  and  a37344a );
 a37354a <=( A167  and  (not A169) );
 a37355a <=( A170  and  a37354a );
 a37359a <=( A200  and  A199 );
 a37360a <=( (not A166)  and  a37359a );
 a37361a <=( a37360a  and  a37355a );
 a37365a <=( (not A266)  and  (not A233) );
 a37366a <=( (not A232)  and  a37365a );
 a37370a <=( A299  and  A298 );
 a37371a <=( (not A267)  and  a37370a );
 a37372a <=( a37371a  and  a37366a );
 a37376a <=( A167  and  (not A169) );
 a37377a <=( A170  and  a37376a );
 a37381a <=( A200  and  A199 );
 a37382a <=( (not A166)  and  a37381a );
 a37383a <=( a37382a  and  a37377a );
 a37387a <=( (not A266)  and  (not A233) );
 a37388a <=( (not A232)  and  a37387a );
 a37392a <=( (not A299)  and  (not A298) );
 a37393a <=( (not A267)  and  a37392a );
 a37394a <=( a37393a  and  a37388a );
 a37398a <=( A167  and  (not A169) );
 a37399a <=( A170  and  a37398a );
 a37403a <=( A200  and  A199 );
 a37404a <=( (not A166)  and  a37403a );
 a37405a <=( a37404a  and  a37399a );
 a37409a <=( (not A265)  and  (not A233) );
 a37410a <=( (not A232)  and  a37409a );
 a37414a <=( (not A300)  and  A298 );
 a37415a <=( (not A266)  and  a37414a );
 a37416a <=( a37415a  and  a37410a );
 a37420a <=( A167  and  (not A169) );
 a37421a <=( A170  and  a37420a );
 a37425a <=( A200  and  A199 );
 a37426a <=( (not A166)  and  a37425a );
 a37427a <=( a37426a  and  a37421a );
 a37431a <=( (not A265)  and  (not A233) );
 a37432a <=( (not A232)  and  a37431a );
 a37436a <=( A299  and  A298 );
 a37437a <=( (not A266)  and  a37436a );
 a37438a <=( a37437a  and  a37432a );
 a37442a <=( A167  and  (not A169) );
 a37443a <=( A170  and  a37442a );
 a37447a <=( A200  and  A199 );
 a37448a <=( (not A166)  and  a37447a );
 a37449a <=( a37448a  and  a37443a );
 a37453a <=( (not A265)  and  (not A233) );
 a37454a <=( (not A232)  and  a37453a );
 a37458a <=( (not A299)  and  (not A298) );
 a37459a <=( (not A266)  and  a37458a );
 a37460a <=( a37459a  and  a37454a );
 a37464a <=( A167  and  (not A169) );
 a37465a <=( A170  and  a37464a );
 a37469a <=( (not A201)  and  (not A200) );
 a37470a <=( (not A166)  and  a37469a );
 a37471a <=( a37470a  and  a37465a );
 a37475a <=( A265  and  A233 );
 a37476a <=( A232  and  a37475a );
 a37480a <=( (not A300)  and  (not A299) );
 a37481a <=( (not A267)  and  a37480a );
 a37482a <=( a37481a  and  a37476a );
 a37486a <=( A167  and  (not A169) );
 a37487a <=( A170  and  a37486a );
 a37491a <=( (not A201)  and  (not A200) );
 a37492a <=( (not A166)  and  a37491a );
 a37493a <=( a37492a  and  a37487a );
 a37497a <=( A265  and  A233 );
 a37498a <=( A232  and  a37497a );
 a37502a <=( A299  and  A298 );
 a37503a <=( (not A267)  and  a37502a );
 a37504a <=( a37503a  and  a37498a );
 a37508a <=( A167  and  (not A169) );
 a37509a <=( A170  and  a37508a );
 a37513a <=( (not A201)  and  (not A200) );
 a37514a <=( (not A166)  and  a37513a );
 a37515a <=( a37514a  and  a37509a );
 a37519a <=( A265  and  A233 );
 a37520a <=( A232  and  a37519a );
 a37524a <=( (not A299)  and  (not A298) );
 a37525a <=( (not A267)  and  a37524a );
 a37526a <=( a37525a  and  a37520a );
 a37530a <=( A167  and  (not A169) );
 a37531a <=( A170  and  a37530a );
 a37535a <=( (not A201)  and  (not A200) );
 a37536a <=( (not A166)  and  a37535a );
 a37537a <=( a37536a  and  a37531a );
 a37541a <=( A265  and  A233 );
 a37542a <=( A232  and  a37541a );
 a37546a <=( (not A300)  and  (not A299) );
 a37547a <=( A266  and  a37546a );
 a37548a <=( a37547a  and  a37542a );
 a37552a <=( A167  and  (not A169) );
 a37553a <=( A170  and  a37552a );
 a37557a <=( (not A201)  and  (not A200) );
 a37558a <=( (not A166)  and  a37557a );
 a37559a <=( a37558a  and  a37553a );
 a37563a <=( A265  and  A233 );
 a37564a <=( A232  and  a37563a );
 a37568a <=( A299  and  A298 );
 a37569a <=( A266  and  a37568a );
 a37570a <=( a37569a  and  a37564a );
 a37574a <=( A167  and  (not A169) );
 a37575a <=( A170  and  a37574a );
 a37579a <=( (not A201)  and  (not A200) );
 a37580a <=( (not A166)  and  a37579a );
 a37581a <=( a37580a  and  a37575a );
 a37585a <=( A265  and  A233 );
 a37586a <=( A232  and  a37585a );
 a37590a <=( (not A299)  and  (not A298) );
 a37591a <=( A266  and  a37590a );
 a37592a <=( a37591a  and  a37586a );
 a37596a <=( A167  and  (not A169) );
 a37597a <=( A170  and  a37596a );
 a37601a <=( (not A201)  and  (not A200) );
 a37602a <=( (not A166)  and  a37601a );
 a37603a <=( a37602a  and  a37597a );
 a37607a <=( (not A265)  and  A233 );
 a37608a <=( A232  and  a37607a );
 a37612a <=( (not A300)  and  (not A299) );
 a37613a <=( (not A266)  and  a37612a );
 a37614a <=( a37613a  and  a37608a );
 a37618a <=( A167  and  (not A169) );
 a37619a <=( A170  and  a37618a );
 a37623a <=( (not A201)  and  (not A200) );
 a37624a <=( (not A166)  and  a37623a );
 a37625a <=( a37624a  and  a37619a );
 a37629a <=( (not A265)  and  A233 );
 a37630a <=( A232  and  a37629a );
 a37634a <=( A299  and  A298 );
 a37635a <=( (not A266)  and  a37634a );
 a37636a <=( a37635a  and  a37630a );
 a37640a <=( A167  and  (not A169) );
 a37641a <=( A170  and  a37640a );
 a37645a <=( (not A201)  and  (not A200) );
 a37646a <=( (not A166)  and  a37645a );
 a37647a <=( a37646a  and  a37641a );
 a37651a <=( (not A265)  and  A233 );
 a37652a <=( A232  and  a37651a );
 a37656a <=( (not A299)  and  (not A298) );
 a37657a <=( (not A266)  and  a37656a );
 a37658a <=( a37657a  and  a37652a );
 a37662a <=( A167  and  (not A169) );
 a37663a <=( A170  and  a37662a );
 a37667a <=( (not A201)  and  (not A200) );
 a37668a <=( (not A166)  and  a37667a );
 a37669a <=( a37668a  and  a37663a );
 a37673a <=( A298  and  A233 );
 a37674a <=( (not A232)  and  a37673a );
 a37678a <=( A301  and  A300 );
 a37679a <=( (not A299)  and  a37678a );
 a37680a <=( a37679a  and  a37674a );
 a37684a <=( A167  and  (not A169) );
 a37685a <=( A170  and  a37684a );
 a37689a <=( (not A201)  and  (not A200) );
 a37690a <=( (not A166)  and  a37689a );
 a37691a <=( a37690a  and  a37685a );
 a37695a <=( A298  and  A233 );
 a37696a <=( (not A232)  and  a37695a );
 a37700a <=( A302  and  A300 );
 a37701a <=( (not A299)  and  a37700a );
 a37702a <=( a37701a  and  a37696a );
 a37706a <=( A167  and  (not A169) );
 a37707a <=( A170  and  a37706a );
 a37711a <=( (not A201)  and  (not A200) );
 a37712a <=( (not A166)  and  a37711a );
 a37713a <=( a37712a  and  a37707a );
 a37717a <=( A265  and  A233 );
 a37718a <=( (not A232)  and  a37717a );
 a37722a <=( A268  and  A267 );
 a37723a <=( (not A266)  and  a37722a );
 a37724a <=( a37723a  and  a37718a );
 a37728a <=( A167  and  (not A169) );
 a37729a <=( A170  and  a37728a );
 a37733a <=( (not A201)  and  (not A200) );
 a37734a <=( (not A166)  and  a37733a );
 a37735a <=( a37734a  and  a37729a );
 a37739a <=( A265  and  A233 );
 a37740a <=( (not A232)  and  a37739a );
 a37744a <=( A269  and  A267 );
 a37745a <=( (not A266)  and  a37744a );
 a37746a <=( a37745a  and  a37740a );
 a37750a <=( A167  and  (not A169) );
 a37751a <=( A170  and  a37750a );
 a37755a <=( (not A201)  and  (not A200) );
 a37756a <=( (not A166)  and  a37755a );
 a37757a <=( a37756a  and  a37751a );
 a37761a <=( A265  and  (not A234) );
 a37762a <=( (not A233)  and  a37761a );
 a37766a <=( (not A300)  and  A298 );
 a37767a <=( A266  and  a37766a );
 a37768a <=( a37767a  and  a37762a );
 a37772a <=( A167  and  (not A169) );
 a37773a <=( A170  and  a37772a );
 a37777a <=( (not A201)  and  (not A200) );
 a37778a <=( (not A166)  and  a37777a );
 a37779a <=( a37778a  and  a37773a );
 a37783a <=( A265  and  (not A234) );
 a37784a <=( (not A233)  and  a37783a );
 a37788a <=( A299  and  A298 );
 a37789a <=( A266  and  a37788a );
 a37790a <=( a37789a  and  a37784a );
 a37794a <=( A167  and  (not A169) );
 a37795a <=( A170  and  a37794a );
 a37799a <=( (not A201)  and  (not A200) );
 a37800a <=( (not A166)  and  a37799a );
 a37801a <=( a37800a  and  a37795a );
 a37805a <=( A265  and  (not A234) );
 a37806a <=( (not A233)  and  a37805a );
 a37810a <=( (not A299)  and  (not A298) );
 a37811a <=( A266  and  a37810a );
 a37812a <=( a37811a  and  a37806a );
 a37816a <=( A167  and  (not A169) );
 a37817a <=( A170  and  a37816a );
 a37821a <=( (not A201)  and  (not A200) );
 a37822a <=( (not A166)  and  a37821a );
 a37823a <=( a37822a  and  a37817a );
 a37827a <=( (not A266)  and  (not A234) );
 a37828a <=( (not A233)  and  a37827a );
 a37832a <=( (not A300)  and  A298 );
 a37833a <=( (not A267)  and  a37832a );
 a37834a <=( a37833a  and  a37828a );
 a37838a <=( A167  and  (not A169) );
 a37839a <=( A170  and  a37838a );
 a37843a <=( (not A201)  and  (not A200) );
 a37844a <=( (not A166)  and  a37843a );
 a37845a <=( a37844a  and  a37839a );
 a37849a <=( (not A266)  and  (not A234) );
 a37850a <=( (not A233)  and  a37849a );
 a37854a <=( A299  and  A298 );
 a37855a <=( (not A267)  and  a37854a );
 a37856a <=( a37855a  and  a37850a );
 a37860a <=( A167  and  (not A169) );
 a37861a <=( A170  and  a37860a );
 a37865a <=( (not A201)  and  (not A200) );
 a37866a <=( (not A166)  and  a37865a );
 a37867a <=( a37866a  and  a37861a );
 a37871a <=( (not A266)  and  (not A234) );
 a37872a <=( (not A233)  and  a37871a );
 a37876a <=( (not A299)  and  (not A298) );
 a37877a <=( (not A267)  and  a37876a );
 a37878a <=( a37877a  and  a37872a );
 a37882a <=( A167  and  (not A169) );
 a37883a <=( A170  and  a37882a );
 a37887a <=( (not A201)  and  (not A200) );
 a37888a <=( (not A166)  and  a37887a );
 a37889a <=( a37888a  and  a37883a );
 a37893a <=( (not A265)  and  (not A234) );
 a37894a <=( (not A233)  and  a37893a );
 a37898a <=( (not A300)  and  A298 );
 a37899a <=( (not A266)  and  a37898a );
 a37900a <=( a37899a  and  a37894a );
 a37904a <=( A167  and  (not A169) );
 a37905a <=( A170  and  a37904a );
 a37909a <=( (not A201)  and  (not A200) );
 a37910a <=( (not A166)  and  a37909a );
 a37911a <=( a37910a  and  a37905a );
 a37915a <=( (not A265)  and  (not A234) );
 a37916a <=( (not A233)  and  a37915a );
 a37920a <=( A299  and  A298 );
 a37921a <=( (not A266)  and  a37920a );
 a37922a <=( a37921a  and  a37916a );
 a37926a <=( A167  and  (not A169) );
 a37927a <=( A170  and  a37926a );
 a37931a <=( (not A201)  and  (not A200) );
 a37932a <=( (not A166)  and  a37931a );
 a37933a <=( a37932a  and  a37927a );
 a37937a <=( (not A265)  and  (not A234) );
 a37938a <=( (not A233)  and  a37937a );
 a37942a <=( (not A299)  and  (not A298) );
 a37943a <=( (not A266)  and  a37942a );
 a37944a <=( a37943a  and  a37938a );
 a37948a <=( A167  and  (not A169) );
 a37949a <=( A170  and  a37948a );
 a37953a <=( (not A201)  and  (not A200) );
 a37954a <=( (not A166)  and  a37953a );
 a37955a <=( a37954a  and  a37949a );
 a37959a <=( A234  and  (not A233) );
 a37960a <=( A232  and  a37959a );
 a37964a <=( A299  and  (not A298) );
 a37965a <=( A235  and  a37964a );
 a37966a <=( a37965a  and  a37960a );
 a37970a <=( A167  and  (not A169) );
 a37971a <=( A170  and  a37970a );
 a37975a <=( (not A201)  and  (not A200) );
 a37976a <=( (not A166)  and  a37975a );
 a37977a <=( a37976a  and  a37971a );
 a37981a <=( A234  and  (not A233) );
 a37982a <=( A232  and  a37981a );
 a37986a <=( A266  and  (not A265) );
 a37987a <=( A235  and  a37986a );
 a37988a <=( a37987a  and  a37982a );
 a37992a <=( A167  and  (not A169) );
 a37993a <=( A170  and  a37992a );
 a37997a <=( (not A201)  and  (not A200) );
 a37998a <=( (not A166)  and  a37997a );
 a37999a <=( a37998a  and  a37993a );
 a38003a <=( A234  and  (not A233) );
 a38004a <=( A232  and  a38003a );
 a38008a <=( A299  and  (not A298) );
 a38009a <=( A236  and  a38008a );
 a38010a <=( a38009a  and  a38004a );
 a38014a <=( A167  and  (not A169) );
 a38015a <=( A170  and  a38014a );
 a38019a <=( (not A201)  and  (not A200) );
 a38020a <=( (not A166)  and  a38019a );
 a38021a <=( a38020a  and  a38015a );
 a38025a <=( A234  and  (not A233) );
 a38026a <=( A232  and  a38025a );
 a38030a <=( A266  and  (not A265) );
 a38031a <=( A236  and  a38030a );
 a38032a <=( a38031a  and  a38026a );
 a38036a <=( A167  and  (not A169) );
 a38037a <=( A170  and  a38036a );
 a38041a <=( (not A201)  and  (not A200) );
 a38042a <=( (not A166)  and  a38041a );
 a38043a <=( a38042a  and  a38037a );
 a38047a <=( A265  and  (not A233) );
 a38048a <=( (not A232)  and  a38047a );
 a38052a <=( (not A300)  and  A298 );
 a38053a <=( A266  and  a38052a );
 a38054a <=( a38053a  and  a38048a );
 a38058a <=( A167  and  (not A169) );
 a38059a <=( A170  and  a38058a );
 a38063a <=( (not A201)  and  (not A200) );
 a38064a <=( (not A166)  and  a38063a );
 a38065a <=( a38064a  and  a38059a );
 a38069a <=( A265  and  (not A233) );
 a38070a <=( (not A232)  and  a38069a );
 a38074a <=( A299  and  A298 );
 a38075a <=( A266  and  a38074a );
 a38076a <=( a38075a  and  a38070a );
 a38080a <=( A167  and  (not A169) );
 a38081a <=( A170  and  a38080a );
 a38085a <=( (not A201)  and  (not A200) );
 a38086a <=( (not A166)  and  a38085a );
 a38087a <=( a38086a  and  a38081a );
 a38091a <=( A265  and  (not A233) );
 a38092a <=( (not A232)  and  a38091a );
 a38096a <=( (not A299)  and  (not A298) );
 a38097a <=( A266  and  a38096a );
 a38098a <=( a38097a  and  a38092a );
 a38102a <=( A167  and  (not A169) );
 a38103a <=( A170  and  a38102a );
 a38107a <=( (not A201)  and  (not A200) );
 a38108a <=( (not A166)  and  a38107a );
 a38109a <=( a38108a  and  a38103a );
 a38113a <=( (not A266)  and  (not A233) );
 a38114a <=( (not A232)  and  a38113a );
 a38118a <=( (not A300)  and  A298 );
 a38119a <=( (not A267)  and  a38118a );
 a38120a <=( a38119a  and  a38114a );
 a38124a <=( A167  and  (not A169) );
 a38125a <=( A170  and  a38124a );
 a38129a <=( (not A201)  and  (not A200) );
 a38130a <=( (not A166)  and  a38129a );
 a38131a <=( a38130a  and  a38125a );
 a38135a <=( (not A266)  and  (not A233) );
 a38136a <=( (not A232)  and  a38135a );
 a38140a <=( A299  and  A298 );
 a38141a <=( (not A267)  and  a38140a );
 a38142a <=( a38141a  and  a38136a );
 a38146a <=( A167  and  (not A169) );
 a38147a <=( A170  and  a38146a );
 a38151a <=( (not A201)  and  (not A200) );
 a38152a <=( (not A166)  and  a38151a );
 a38153a <=( a38152a  and  a38147a );
 a38157a <=( (not A266)  and  (not A233) );
 a38158a <=( (not A232)  and  a38157a );
 a38162a <=( (not A299)  and  (not A298) );
 a38163a <=( (not A267)  and  a38162a );
 a38164a <=( a38163a  and  a38158a );
 a38168a <=( A167  and  (not A169) );
 a38169a <=( A170  and  a38168a );
 a38173a <=( (not A201)  and  (not A200) );
 a38174a <=( (not A166)  and  a38173a );
 a38175a <=( a38174a  and  a38169a );
 a38179a <=( (not A265)  and  (not A233) );
 a38180a <=( (not A232)  and  a38179a );
 a38184a <=( (not A300)  and  A298 );
 a38185a <=( (not A266)  and  a38184a );
 a38186a <=( a38185a  and  a38180a );
 a38190a <=( A167  and  (not A169) );
 a38191a <=( A170  and  a38190a );
 a38195a <=( (not A201)  and  (not A200) );
 a38196a <=( (not A166)  and  a38195a );
 a38197a <=( a38196a  and  a38191a );
 a38201a <=( (not A265)  and  (not A233) );
 a38202a <=( (not A232)  and  a38201a );
 a38206a <=( A299  and  A298 );
 a38207a <=( (not A266)  and  a38206a );
 a38208a <=( a38207a  and  a38202a );
 a38212a <=( A167  and  (not A169) );
 a38213a <=( A170  and  a38212a );
 a38217a <=( (not A201)  and  (not A200) );
 a38218a <=( (not A166)  and  a38217a );
 a38219a <=( a38218a  and  a38213a );
 a38223a <=( (not A265)  and  (not A233) );
 a38224a <=( (not A232)  and  a38223a );
 a38228a <=( (not A299)  and  (not A298) );
 a38229a <=( (not A266)  and  a38228a );
 a38230a <=( a38229a  and  a38224a );
 a38234a <=( A167  and  (not A169) );
 a38235a <=( A170  and  a38234a );
 a38239a <=( (not A200)  and  (not A199) );
 a38240a <=( (not A166)  and  a38239a );
 a38241a <=( a38240a  and  a38235a );
 a38245a <=( A265  and  A233 );
 a38246a <=( A232  and  a38245a );
 a38250a <=( (not A300)  and  (not A299) );
 a38251a <=( (not A267)  and  a38250a );
 a38252a <=( a38251a  and  a38246a );
 a38256a <=( A167  and  (not A169) );
 a38257a <=( A170  and  a38256a );
 a38261a <=( (not A200)  and  (not A199) );
 a38262a <=( (not A166)  and  a38261a );
 a38263a <=( a38262a  and  a38257a );
 a38267a <=( A265  and  A233 );
 a38268a <=( A232  and  a38267a );
 a38272a <=( A299  and  A298 );
 a38273a <=( (not A267)  and  a38272a );
 a38274a <=( a38273a  and  a38268a );
 a38278a <=( A167  and  (not A169) );
 a38279a <=( A170  and  a38278a );
 a38283a <=( (not A200)  and  (not A199) );
 a38284a <=( (not A166)  and  a38283a );
 a38285a <=( a38284a  and  a38279a );
 a38289a <=( A265  and  A233 );
 a38290a <=( A232  and  a38289a );
 a38294a <=( (not A299)  and  (not A298) );
 a38295a <=( (not A267)  and  a38294a );
 a38296a <=( a38295a  and  a38290a );
 a38300a <=( A167  and  (not A169) );
 a38301a <=( A170  and  a38300a );
 a38305a <=( (not A200)  and  (not A199) );
 a38306a <=( (not A166)  and  a38305a );
 a38307a <=( a38306a  and  a38301a );
 a38311a <=( A265  and  A233 );
 a38312a <=( A232  and  a38311a );
 a38316a <=( (not A300)  and  (not A299) );
 a38317a <=( A266  and  a38316a );
 a38318a <=( a38317a  and  a38312a );
 a38322a <=( A167  and  (not A169) );
 a38323a <=( A170  and  a38322a );
 a38327a <=( (not A200)  and  (not A199) );
 a38328a <=( (not A166)  and  a38327a );
 a38329a <=( a38328a  and  a38323a );
 a38333a <=( A265  and  A233 );
 a38334a <=( A232  and  a38333a );
 a38338a <=( A299  and  A298 );
 a38339a <=( A266  and  a38338a );
 a38340a <=( a38339a  and  a38334a );
 a38344a <=( A167  and  (not A169) );
 a38345a <=( A170  and  a38344a );
 a38349a <=( (not A200)  and  (not A199) );
 a38350a <=( (not A166)  and  a38349a );
 a38351a <=( a38350a  and  a38345a );
 a38355a <=( A265  and  A233 );
 a38356a <=( A232  and  a38355a );
 a38360a <=( (not A299)  and  (not A298) );
 a38361a <=( A266  and  a38360a );
 a38362a <=( a38361a  and  a38356a );
 a38366a <=( A167  and  (not A169) );
 a38367a <=( A170  and  a38366a );
 a38371a <=( (not A200)  and  (not A199) );
 a38372a <=( (not A166)  and  a38371a );
 a38373a <=( a38372a  and  a38367a );
 a38377a <=( (not A265)  and  A233 );
 a38378a <=( A232  and  a38377a );
 a38382a <=( (not A300)  and  (not A299) );
 a38383a <=( (not A266)  and  a38382a );
 a38384a <=( a38383a  and  a38378a );
 a38388a <=( A167  and  (not A169) );
 a38389a <=( A170  and  a38388a );
 a38393a <=( (not A200)  and  (not A199) );
 a38394a <=( (not A166)  and  a38393a );
 a38395a <=( a38394a  and  a38389a );
 a38399a <=( (not A265)  and  A233 );
 a38400a <=( A232  and  a38399a );
 a38404a <=( A299  and  A298 );
 a38405a <=( (not A266)  and  a38404a );
 a38406a <=( a38405a  and  a38400a );
 a38410a <=( A167  and  (not A169) );
 a38411a <=( A170  and  a38410a );
 a38415a <=( (not A200)  and  (not A199) );
 a38416a <=( (not A166)  and  a38415a );
 a38417a <=( a38416a  and  a38411a );
 a38421a <=( (not A265)  and  A233 );
 a38422a <=( A232  and  a38421a );
 a38426a <=( (not A299)  and  (not A298) );
 a38427a <=( (not A266)  and  a38426a );
 a38428a <=( a38427a  and  a38422a );
 a38432a <=( A167  and  (not A169) );
 a38433a <=( A170  and  a38432a );
 a38437a <=( (not A200)  and  (not A199) );
 a38438a <=( (not A166)  and  a38437a );
 a38439a <=( a38438a  and  a38433a );
 a38443a <=( A298  and  A233 );
 a38444a <=( (not A232)  and  a38443a );
 a38448a <=( A301  and  A300 );
 a38449a <=( (not A299)  and  a38448a );
 a38450a <=( a38449a  and  a38444a );
 a38454a <=( A167  and  (not A169) );
 a38455a <=( A170  and  a38454a );
 a38459a <=( (not A200)  and  (not A199) );
 a38460a <=( (not A166)  and  a38459a );
 a38461a <=( a38460a  and  a38455a );
 a38465a <=( A298  and  A233 );
 a38466a <=( (not A232)  and  a38465a );
 a38470a <=( A302  and  A300 );
 a38471a <=( (not A299)  and  a38470a );
 a38472a <=( a38471a  and  a38466a );
 a38476a <=( A167  and  (not A169) );
 a38477a <=( A170  and  a38476a );
 a38481a <=( (not A200)  and  (not A199) );
 a38482a <=( (not A166)  and  a38481a );
 a38483a <=( a38482a  and  a38477a );
 a38487a <=( A265  and  A233 );
 a38488a <=( (not A232)  and  a38487a );
 a38492a <=( A268  and  A267 );
 a38493a <=( (not A266)  and  a38492a );
 a38494a <=( a38493a  and  a38488a );
 a38498a <=( A167  and  (not A169) );
 a38499a <=( A170  and  a38498a );
 a38503a <=( (not A200)  and  (not A199) );
 a38504a <=( (not A166)  and  a38503a );
 a38505a <=( a38504a  and  a38499a );
 a38509a <=( A265  and  A233 );
 a38510a <=( (not A232)  and  a38509a );
 a38514a <=( A269  and  A267 );
 a38515a <=( (not A266)  and  a38514a );
 a38516a <=( a38515a  and  a38510a );
 a38520a <=( A167  and  (not A169) );
 a38521a <=( A170  and  a38520a );
 a38525a <=( (not A200)  and  (not A199) );
 a38526a <=( (not A166)  and  a38525a );
 a38527a <=( a38526a  and  a38521a );
 a38531a <=( A265  and  (not A234) );
 a38532a <=( (not A233)  and  a38531a );
 a38536a <=( (not A300)  and  A298 );
 a38537a <=( A266  and  a38536a );
 a38538a <=( a38537a  and  a38532a );
 a38542a <=( A167  and  (not A169) );
 a38543a <=( A170  and  a38542a );
 a38547a <=( (not A200)  and  (not A199) );
 a38548a <=( (not A166)  and  a38547a );
 a38549a <=( a38548a  and  a38543a );
 a38553a <=( A265  and  (not A234) );
 a38554a <=( (not A233)  and  a38553a );
 a38558a <=( A299  and  A298 );
 a38559a <=( A266  and  a38558a );
 a38560a <=( a38559a  and  a38554a );
 a38564a <=( A167  and  (not A169) );
 a38565a <=( A170  and  a38564a );
 a38569a <=( (not A200)  and  (not A199) );
 a38570a <=( (not A166)  and  a38569a );
 a38571a <=( a38570a  and  a38565a );
 a38575a <=( A265  and  (not A234) );
 a38576a <=( (not A233)  and  a38575a );
 a38580a <=( (not A299)  and  (not A298) );
 a38581a <=( A266  and  a38580a );
 a38582a <=( a38581a  and  a38576a );
 a38586a <=( A167  and  (not A169) );
 a38587a <=( A170  and  a38586a );
 a38591a <=( (not A200)  and  (not A199) );
 a38592a <=( (not A166)  and  a38591a );
 a38593a <=( a38592a  and  a38587a );
 a38597a <=( (not A266)  and  (not A234) );
 a38598a <=( (not A233)  and  a38597a );
 a38602a <=( (not A300)  and  A298 );
 a38603a <=( (not A267)  and  a38602a );
 a38604a <=( a38603a  and  a38598a );
 a38608a <=( A167  and  (not A169) );
 a38609a <=( A170  and  a38608a );
 a38613a <=( (not A200)  and  (not A199) );
 a38614a <=( (not A166)  and  a38613a );
 a38615a <=( a38614a  and  a38609a );
 a38619a <=( (not A266)  and  (not A234) );
 a38620a <=( (not A233)  and  a38619a );
 a38624a <=( A299  and  A298 );
 a38625a <=( (not A267)  and  a38624a );
 a38626a <=( a38625a  and  a38620a );
 a38630a <=( A167  and  (not A169) );
 a38631a <=( A170  and  a38630a );
 a38635a <=( (not A200)  and  (not A199) );
 a38636a <=( (not A166)  and  a38635a );
 a38637a <=( a38636a  and  a38631a );
 a38641a <=( (not A266)  and  (not A234) );
 a38642a <=( (not A233)  and  a38641a );
 a38646a <=( (not A299)  and  (not A298) );
 a38647a <=( (not A267)  and  a38646a );
 a38648a <=( a38647a  and  a38642a );
 a38652a <=( A167  and  (not A169) );
 a38653a <=( A170  and  a38652a );
 a38657a <=( (not A200)  and  (not A199) );
 a38658a <=( (not A166)  and  a38657a );
 a38659a <=( a38658a  and  a38653a );
 a38663a <=( (not A265)  and  (not A234) );
 a38664a <=( (not A233)  and  a38663a );
 a38668a <=( (not A300)  and  A298 );
 a38669a <=( (not A266)  and  a38668a );
 a38670a <=( a38669a  and  a38664a );
 a38674a <=( A167  and  (not A169) );
 a38675a <=( A170  and  a38674a );
 a38679a <=( (not A200)  and  (not A199) );
 a38680a <=( (not A166)  and  a38679a );
 a38681a <=( a38680a  and  a38675a );
 a38685a <=( (not A265)  and  (not A234) );
 a38686a <=( (not A233)  and  a38685a );
 a38690a <=( A299  and  A298 );
 a38691a <=( (not A266)  and  a38690a );
 a38692a <=( a38691a  and  a38686a );
 a38696a <=( A167  and  (not A169) );
 a38697a <=( A170  and  a38696a );
 a38701a <=( (not A200)  and  (not A199) );
 a38702a <=( (not A166)  and  a38701a );
 a38703a <=( a38702a  and  a38697a );
 a38707a <=( (not A265)  and  (not A234) );
 a38708a <=( (not A233)  and  a38707a );
 a38712a <=( (not A299)  and  (not A298) );
 a38713a <=( (not A266)  and  a38712a );
 a38714a <=( a38713a  and  a38708a );
 a38718a <=( A167  and  (not A169) );
 a38719a <=( A170  and  a38718a );
 a38723a <=( (not A200)  and  (not A199) );
 a38724a <=( (not A166)  and  a38723a );
 a38725a <=( a38724a  and  a38719a );
 a38729a <=( A234  and  (not A233) );
 a38730a <=( A232  and  a38729a );
 a38734a <=( A299  and  (not A298) );
 a38735a <=( A235  and  a38734a );
 a38736a <=( a38735a  and  a38730a );
 a38740a <=( A167  and  (not A169) );
 a38741a <=( A170  and  a38740a );
 a38745a <=( (not A200)  and  (not A199) );
 a38746a <=( (not A166)  and  a38745a );
 a38747a <=( a38746a  and  a38741a );
 a38751a <=( A234  and  (not A233) );
 a38752a <=( A232  and  a38751a );
 a38756a <=( A266  and  (not A265) );
 a38757a <=( A235  and  a38756a );
 a38758a <=( a38757a  and  a38752a );
 a38762a <=( A167  and  (not A169) );
 a38763a <=( A170  and  a38762a );
 a38767a <=( (not A200)  and  (not A199) );
 a38768a <=( (not A166)  and  a38767a );
 a38769a <=( a38768a  and  a38763a );
 a38773a <=( A234  and  (not A233) );
 a38774a <=( A232  and  a38773a );
 a38778a <=( A299  and  (not A298) );
 a38779a <=( A236  and  a38778a );
 a38780a <=( a38779a  and  a38774a );
 a38784a <=( A167  and  (not A169) );
 a38785a <=( A170  and  a38784a );
 a38789a <=( (not A200)  and  (not A199) );
 a38790a <=( (not A166)  and  a38789a );
 a38791a <=( a38790a  and  a38785a );
 a38795a <=( A234  and  (not A233) );
 a38796a <=( A232  and  a38795a );
 a38800a <=( A266  and  (not A265) );
 a38801a <=( A236  and  a38800a );
 a38802a <=( a38801a  and  a38796a );
 a38806a <=( A167  and  (not A169) );
 a38807a <=( A170  and  a38806a );
 a38811a <=( (not A200)  and  (not A199) );
 a38812a <=( (not A166)  and  a38811a );
 a38813a <=( a38812a  and  a38807a );
 a38817a <=( A265  and  (not A233) );
 a38818a <=( (not A232)  and  a38817a );
 a38822a <=( (not A300)  and  A298 );
 a38823a <=( A266  and  a38822a );
 a38824a <=( a38823a  and  a38818a );
 a38828a <=( A167  and  (not A169) );
 a38829a <=( A170  and  a38828a );
 a38833a <=( (not A200)  and  (not A199) );
 a38834a <=( (not A166)  and  a38833a );
 a38835a <=( a38834a  and  a38829a );
 a38839a <=( A265  and  (not A233) );
 a38840a <=( (not A232)  and  a38839a );
 a38844a <=( A299  and  A298 );
 a38845a <=( A266  and  a38844a );
 a38846a <=( a38845a  and  a38840a );
 a38850a <=( A167  and  (not A169) );
 a38851a <=( A170  and  a38850a );
 a38855a <=( (not A200)  and  (not A199) );
 a38856a <=( (not A166)  and  a38855a );
 a38857a <=( a38856a  and  a38851a );
 a38861a <=( A265  and  (not A233) );
 a38862a <=( (not A232)  and  a38861a );
 a38866a <=( (not A299)  and  (not A298) );
 a38867a <=( A266  and  a38866a );
 a38868a <=( a38867a  and  a38862a );
 a38872a <=( A167  and  (not A169) );
 a38873a <=( A170  and  a38872a );
 a38877a <=( (not A200)  and  (not A199) );
 a38878a <=( (not A166)  and  a38877a );
 a38879a <=( a38878a  and  a38873a );
 a38883a <=( (not A266)  and  (not A233) );
 a38884a <=( (not A232)  and  a38883a );
 a38888a <=( (not A300)  and  A298 );
 a38889a <=( (not A267)  and  a38888a );
 a38890a <=( a38889a  and  a38884a );
 a38894a <=( A167  and  (not A169) );
 a38895a <=( A170  and  a38894a );
 a38899a <=( (not A200)  and  (not A199) );
 a38900a <=( (not A166)  and  a38899a );
 a38901a <=( a38900a  and  a38895a );
 a38905a <=( (not A266)  and  (not A233) );
 a38906a <=( (not A232)  and  a38905a );
 a38910a <=( A299  and  A298 );
 a38911a <=( (not A267)  and  a38910a );
 a38912a <=( a38911a  and  a38906a );
 a38916a <=( A167  and  (not A169) );
 a38917a <=( A170  and  a38916a );
 a38921a <=( (not A200)  and  (not A199) );
 a38922a <=( (not A166)  and  a38921a );
 a38923a <=( a38922a  and  a38917a );
 a38927a <=( (not A266)  and  (not A233) );
 a38928a <=( (not A232)  and  a38927a );
 a38932a <=( (not A299)  and  (not A298) );
 a38933a <=( (not A267)  and  a38932a );
 a38934a <=( a38933a  and  a38928a );
 a38938a <=( A167  and  (not A169) );
 a38939a <=( A170  and  a38938a );
 a38943a <=( (not A200)  and  (not A199) );
 a38944a <=( (not A166)  and  a38943a );
 a38945a <=( a38944a  and  a38939a );
 a38949a <=( (not A265)  and  (not A233) );
 a38950a <=( (not A232)  and  a38949a );
 a38954a <=( (not A300)  and  A298 );
 a38955a <=( (not A266)  and  a38954a );
 a38956a <=( a38955a  and  a38950a );
 a38960a <=( A167  and  (not A169) );
 a38961a <=( A170  and  a38960a );
 a38965a <=( (not A200)  and  (not A199) );
 a38966a <=( (not A166)  and  a38965a );
 a38967a <=( a38966a  and  a38961a );
 a38971a <=( (not A265)  and  (not A233) );
 a38972a <=( (not A232)  and  a38971a );
 a38976a <=( A299  and  A298 );
 a38977a <=( (not A266)  and  a38976a );
 a38978a <=( a38977a  and  a38972a );
 a38982a <=( A167  and  (not A169) );
 a38983a <=( A170  and  a38982a );
 a38987a <=( (not A200)  and  (not A199) );
 a38988a <=( (not A166)  and  a38987a );
 a38989a <=( a38988a  and  a38983a );
 a38993a <=( (not A265)  and  (not A233) );
 a38994a <=( (not A232)  and  a38993a );
 a38998a <=( (not A299)  and  (not A298) );
 a38999a <=( (not A266)  and  a38998a );
 a39000a <=( a38999a  and  a38994a );
 a39004a <=( (not A167)  and  (not A169) );
 a39005a <=( A170  and  a39004a );
 a39009a <=( A200  and  A199 );
 a39010a <=( A166  and  a39009a );
 a39011a <=( a39010a  and  a39005a );
 a39015a <=( A265  and  A233 );
 a39016a <=( A232  and  a39015a );
 a39020a <=( (not A300)  and  (not A299) );
 a39021a <=( (not A267)  and  a39020a );
 a39022a <=( a39021a  and  a39016a );
 a39026a <=( (not A167)  and  (not A169) );
 a39027a <=( A170  and  a39026a );
 a39031a <=( A200  and  A199 );
 a39032a <=( A166  and  a39031a );
 a39033a <=( a39032a  and  a39027a );
 a39037a <=( A265  and  A233 );
 a39038a <=( A232  and  a39037a );
 a39042a <=( A299  and  A298 );
 a39043a <=( (not A267)  and  a39042a );
 a39044a <=( a39043a  and  a39038a );
 a39048a <=( (not A167)  and  (not A169) );
 a39049a <=( A170  and  a39048a );
 a39053a <=( A200  and  A199 );
 a39054a <=( A166  and  a39053a );
 a39055a <=( a39054a  and  a39049a );
 a39059a <=( A265  and  A233 );
 a39060a <=( A232  and  a39059a );
 a39064a <=( (not A299)  and  (not A298) );
 a39065a <=( (not A267)  and  a39064a );
 a39066a <=( a39065a  and  a39060a );
 a39070a <=( (not A167)  and  (not A169) );
 a39071a <=( A170  and  a39070a );
 a39075a <=( A200  and  A199 );
 a39076a <=( A166  and  a39075a );
 a39077a <=( a39076a  and  a39071a );
 a39081a <=( A265  and  A233 );
 a39082a <=( A232  and  a39081a );
 a39086a <=( (not A300)  and  (not A299) );
 a39087a <=( A266  and  a39086a );
 a39088a <=( a39087a  and  a39082a );
 a39092a <=( (not A167)  and  (not A169) );
 a39093a <=( A170  and  a39092a );
 a39097a <=( A200  and  A199 );
 a39098a <=( A166  and  a39097a );
 a39099a <=( a39098a  and  a39093a );
 a39103a <=( A265  and  A233 );
 a39104a <=( A232  and  a39103a );
 a39108a <=( A299  and  A298 );
 a39109a <=( A266  and  a39108a );
 a39110a <=( a39109a  and  a39104a );
 a39114a <=( (not A167)  and  (not A169) );
 a39115a <=( A170  and  a39114a );
 a39119a <=( A200  and  A199 );
 a39120a <=( A166  and  a39119a );
 a39121a <=( a39120a  and  a39115a );
 a39125a <=( A265  and  A233 );
 a39126a <=( A232  and  a39125a );
 a39130a <=( (not A299)  and  (not A298) );
 a39131a <=( A266  and  a39130a );
 a39132a <=( a39131a  and  a39126a );
 a39136a <=( (not A167)  and  (not A169) );
 a39137a <=( A170  and  a39136a );
 a39141a <=( A200  and  A199 );
 a39142a <=( A166  and  a39141a );
 a39143a <=( a39142a  and  a39137a );
 a39147a <=( (not A265)  and  A233 );
 a39148a <=( A232  and  a39147a );
 a39152a <=( (not A300)  and  (not A299) );
 a39153a <=( (not A266)  and  a39152a );
 a39154a <=( a39153a  and  a39148a );
 a39158a <=( (not A167)  and  (not A169) );
 a39159a <=( A170  and  a39158a );
 a39163a <=( A200  and  A199 );
 a39164a <=( A166  and  a39163a );
 a39165a <=( a39164a  and  a39159a );
 a39169a <=( (not A265)  and  A233 );
 a39170a <=( A232  and  a39169a );
 a39174a <=( A299  and  A298 );
 a39175a <=( (not A266)  and  a39174a );
 a39176a <=( a39175a  and  a39170a );
 a39180a <=( (not A167)  and  (not A169) );
 a39181a <=( A170  and  a39180a );
 a39185a <=( A200  and  A199 );
 a39186a <=( A166  and  a39185a );
 a39187a <=( a39186a  and  a39181a );
 a39191a <=( (not A265)  and  A233 );
 a39192a <=( A232  and  a39191a );
 a39196a <=( (not A299)  and  (not A298) );
 a39197a <=( (not A266)  and  a39196a );
 a39198a <=( a39197a  and  a39192a );
 a39202a <=( (not A167)  and  (not A169) );
 a39203a <=( A170  and  a39202a );
 a39207a <=( A200  and  A199 );
 a39208a <=( A166  and  a39207a );
 a39209a <=( a39208a  and  a39203a );
 a39213a <=( A298  and  A233 );
 a39214a <=( (not A232)  and  a39213a );
 a39218a <=( A301  and  A300 );
 a39219a <=( (not A299)  and  a39218a );
 a39220a <=( a39219a  and  a39214a );
 a39224a <=( (not A167)  and  (not A169) );
 a39225a <=( A170  and  a39224a );
 a39229a <=( A200  and  A199 );
 a39230a <=( A166  and  a39229a );
 a39231a <=( a39230a  and  a39225a );
 a39235a <=( A298  and  A233 );
 a39236a <=( (not A232)  and  a39235a );
 a39240a <=( A302  and  A300 );
 a39241a <=( (not A299)  and  a39240a );
 a39242a <=( a39241a  and  a39236a );
 a39246a <=( (not A167)  and  (not A169) );
 a39247a <=( A170  and  a39246a );
 a39251a <=( A200  and  A199 );
 a39252a <=( A166  and  a39251a );
 a39253a <=( a39252a  and  a39247a );
 a39257a <=( A265  and  A233 );
 a39258a <=( (not A232)  and  a39257a );
 a39262a <=( A268  and  A267 );
 a39263a <=( (not A266)  and  a39262a );
 a39264a <=( a39263a  and  a39258a );
 a39268a <=( (not A167)  and  (not A169) );
 a39269a <=( A170  and  a39268a );
 a39273a <=( A200  and  A199 );
 a39274a <=( A166  and  a39273a );
 a39275a <=( a39274a  and  a39269a );
 a39279a <=( A265  and  A233 );
 a39280a <=( (not A232)  and  a39279a );
 a39284a <=( A269  and  A267 );
 a39285a <=( (not A266)  and  a39284a );
 a39286a <=( a39285a  and  a39280a );
 a39290a <=( (not A167)  and  (not A169) );
 a39291a <=( A170  and  a39290a );
 a39295a <=( A200  and  A199 );
 a39296a <=( A166  and  a39295a );
 a39297a <=( a39296a  and  a39291a );
 a39301a <=( A265  and  (not A234) );
 a39302a <=( (not A233)  and  a39301a );
 a39306a <=( (not A300)  and  A298 );
 a39307a <=( A266  and  a39306a );
 a39308a <=( a39307a  and  a39302a );
 a39312a <=( (not A167)  and  (not A169) );
 a39313a <=( A170  and  a39312a );
 a39317a <=( A200  and  A199 );
 a39318a <=( A166  and  a39317a );
 a39319a <=( a39318a  and  a39313a );
 a39323a <=( A265  and  (not A234) );
 a39324a <=( (not A233)  and  a39323a );
 a39328a <=( A299  and  A298 );
 a39329a <=( A266  and  a39328a );
 a39330a <=( a39329a  and  a39324a );
 a39334a <=( (not A167)  and  (not A169) );
 a39335a <=( A170  and  a39334a );
 a39339a <=( A200  and  A199 );
 a39340a <=( A166  and  a39339a );
 a39341a <=( a39340a  and  a39335a );
 a39345a <=( A265  and  (not A234) );
 a39346a <=( (not A233)  and  a39345a );
 a39350a <=( (not A299)  and  (not A298) );
 a39351a <=( A266  and  a39350a );
 a39352a <=( a39351a  and  a39346a );
 a39356a <=( (not A167)  and  (not A169) );
 a39357a <=( A170  and  a39356a );
 a39361a <=( A200  and  A199 );
 a39362a <=( A166  and  a39361a );
 a39363a <=( a39362a  and  a39357a );
 a39367a <=( (not A266)  and  (not A234) );
 a39368a <=( (not A233)  and  a39367a );
 a39372a <=( (not A300)  and  A298 );
 a39373a <=( (not A267)  and  a39372a );
 a39374a <=( a39373a  and  a39368a );
 a39378a <=( (not A167)  and  (not A169) );
 a39379a <=( A170  and  a39378a );
 a39383a <=( A200  and  A199 );
 a39384a <=( A166  and  a39383a );
 a39385a <=( a39384a  and  a39379a );
 a39389a <=( (not A266)  and  (not A234) );
 a39390a <=( (not A233)  and  a39389a );
 a39394a <=( A299  and  A298 );
 a39395a <=( (not A267)  and  a39394a );
 a39396a <=( a39395a  and  a39390a );
 a39400a <=( (not A167)  and  (not A169) );
 a39401a <=( A170  and  a39400a );
 a39405a <=( A200  and  A199 );
 a39406a <=( A166  and  a39405a );
 a39407a <=( a39406a  and  a39401a );
 a39411a <=( (not A266)  and  (not A234) );
 a39412a <=( (not A233)  and  a39411a );
 a39416a <=( (not A299)  and  (not A298) );
 a39417a <=( (not A267)  and  a39416a );
 a39418a <=( a39417a  and  a39412a );
 a39422a <=( (not A167)  and  (not A169) );
 a39423a <=( A170  and  a39422a );
 a39427a <=( A200  and  A199 );
 a39428a <=( A166  and  a39427a );
 a39429a <=( a39428a  and  a39423a );
 a39433a <=( (not A265)  and  (not A234) );
 a39434a <=( (not A233)  and  a39433a );
 a39438a <=( (not A300)  and  A298 );
 a39439a <=( (not A266)  and  a39438a );
 a39440a <=( a39439a  and  a39434a );
 a39444a <=( (not A167)  and  (not A169) );
 a39445a <=( A170  and  a39444a );
 a39449a <=( A200  and  A199 );
 a39450a <=( A166  and  a39449a );
 a39451a <=( a39450a  and  a39445a );
 a39455a <=( (not A265)  and  (not A234) );
 a39456a <=( (not A233)  and  a39455a );
 a39460a <=( A299  and  A298 );
 a39461a <=( (not A266)  and  a39460a );
 a39462a <=( a39461a  and  a39456a );
 a39466a <=( (not A167)  and  (not A169) );
 a39467a <=( A170  and  a39466a );
 a39471a <=( A200  and  A199 );
 a39472a <=( A166  and  a39471a );
 a39473a <=( a39472a  and  a39467a );
 a39477a <=( (not A265)  and  (not A234) );
 a39478a <=( (not A233)  and  a39477a );
 a39482a <=( (not A299)  and  (not A298) );
 a39483a <=( (not A266)  and  a39482a );
 a39484a <=( a39483a  and  a39478a );
 a39488a <=( (not A167)  and  (not A169) );
 a39489a <=( A170  and  a39488a );
 a39493a <=( A200  and  A199 );
 a39494a <=( A166  and  a39493a );
 a39495a <=( a39494a  and  a39489a );
 a39499a <=( A234  and  (not A233) );
 a39500a <=( A232  and  a39499a );
 a39504a <=( A299  and  (not A298) );
 a39505a <=( A235  and  a39504a );
 a39506a <=( a39505a  and  a39500a );
 a39510a <=( (not A167)  and  (not A169) );
 a39511a <=( A170  and  a39510a );
 a39515a <=( A200  and  A199 );
 a39516a <=( A166  and  a39515a );
 a39517a <=( a39516a  and  a39511a );
 a39521a <=( A234  and  (not A233) );
 a39522a <=( A232  and  a39521a );
 a39526a <=( A266  and  (not A265) );
 a39527a <=( A235  and  a39526a );
 a39528a <=( a39527a  and  a39522a );
 a39532a <=( (not A167)  and  (not A169) );
 a39533a <=( A170  and  a39532a );
 a39537a <=( A200  and  A199 );
 a39538a <=( A166  and  a39537a );
 a39539a <=( a39538a  and  a39533a );
 a39543a <=( A234  and  (not A233) );
 a39544a <=( A232  and  a39543a );
 a39548a <=( A299  and  (not A298) );
 a39549a <=( A236  and  a39548a );
 a39550a <=( a39549a  and  a39544a );
 a39554a <=( (not A167)  and  (not A169) );
 a39555a <=( A170  and  a39554a );
 a39559a <=( A200  and  A199 );
 a39560a <=( A166  and  a39559a );
 a39561a <=( a39560a  and  a39555a );
 a39565a <=( A234  and  (not A233) );
 a39566a <=( A232  and  a39565a );
 a39570a <=( A266  and  (not A265) );
 a39571a <=( A236  and  a39570a );
 a39572a <=( a39571a  and  a39566a );
 a39576a <=( (not A167)  and  (not A169) );
 a39577a <=( A170  and  a39576a );
 a39581a <=( A200  and  A199 );
 a39582a <=( A166  and  a39581a );
 a39583a <=( a39582a  and  a39577a );
 a39587a <=( A265  and  (not A233) );
 a39588a <=( (not A232)  and  a39587a );
 a39592a <=( (not A300)  and  A298 );
 a39593a <=( A266  and  a39592a );
 a39594a <=( a39593a  and  a39588a );
 a39598a <=( (not A167)  and  (not A169) );
 a39599a <=( A170  and  a39598a );
 a39603a <=( A200  and  A199 );
 a39604a <=( A166  and  a39603a );
 a39605a <=( a39604a  and  a39599a );
 a39609a <=( A265  and  (not A233) );
 a39610a <=( (not A232)  and  a39609a );
 a39614a <=( A299  and  A298 );
 a39615a <=( A266  and  a39614a );
 a39616a <=( a39615a  and  a39610a );
 a39620a <=( (not A167)  and  (not A169) );
 a39621a <=( A170  and  a39620a );
 a39625a <=( A200  and  A199 );
 a39626a <=( A166  and  a39625a );
 a39627a <=( a39626a  and  a39621a );
 a39631a <=( A265  and  (not A233) );
 a39632a <=( (not A232)  and  a39631a );
 a39636a <=( (not A299)  and  (not A298) );
 a39637a <=( A266  and  a39636a );
 a39638a <=( a39637a  and  a39632a );
 a39642a <=( (not A167)  and  (not A169) );
 a39643a <=( A170  and  a39642a );
 a39647a <=( A200  and  A199 );
 a39648a <=( A166  and  a39647a );
 a39649a <=( a39648a  and  a39643a );
 a39653a <=( (not A266)  and  (not A233) );
 a39654a <=( (not A232)  and  a39653a );
 a39658a <=( (not A300)  and  A298 );
 a39659a <=( (not A267)  and  a39658a );
 a39660a <=( a39659a  and  a39654a );
 a39664a <=( (not A167)  and  (not A169) );
 a39665a <=( A170  and  a39664a );
 a39669a <=( A200  and  A199 );
 a39670a <=( A166  and  a39669a );
 a39671a <=( a39670a  and  a39665a );
 a39675a <=( (not A266)  and  (not A233) );
 a39676a <=( (not A232)  and  a39675a );
 a39680a <=( A299  and  A298 );
 a39681a <=( (not A267)  and  a39680a );
 a39682a <=( a39681a  and  a39676a );
 a39686a <=( (not A167)  and  (not A169) );
 a39687a <=( A170  and  a39686a );
 a39691a <=( A200  and  A199 );
 a39692a <=( A166  and  a39691a );
 a39693a <=( a39692a  and  a39687a );
 a39697a <=( (not A266)  and  (not A233) );
 a39698a <=( (not A232)  and  a39697a );
 a39702a <=( (not A299)  and  (not A298) );
 a39703a <=( (not A267)  and  a39702a );
 a39704a <=( a39703a  and  a39698a );
 a39708a <=( (not A167)  and  (not A169) );
 a39709a <=( A170  and  a39708a );
 a39713a <=( A200  and  A199 );
 a39714a <=( A166  and  a39713a );
 a39715a <=( a39714a  and  a39709a );
 a39719a <=( (not A265)  and  (not A233) );
 a39720a <=( (not A232)  and  a39719a );
 a39724a <=( (not A300)  and  A298 );
 a39725a <=( (not A266)  and  a39724a );
 a39726a <=( a39725a  and  a39720a );
 a39730a <=( (not A167)  and  (not A169) );
 a39731a <=( A170  and  a39730a );
 a39735a <=( A200  and  A199 );
 a39736a <=( A166  and  a39735a );
 a39737a <=( a39736a  and  a39731a );
 a39741a <=( (not A265)  and  (not A233) );
 a39742a <=( (not A232)  and  a39741a );
 a39746a <=( A299  and  A298 );
 a39747a <=( (not A266)  and  a39746a );
 a39748a <=( a39747a  and  a39742a );
 a39752a <=( (not A167)  and  (not A169) );
 a39753a <=( A170  and  a39752a );
 a39757a <=( A200  and  A199 );
 a39758a <=( A166  and  a39757a );
 a39759a <=( a39758a  and  a39753a );
 a39763a <=( (not A265)  and  (not A233) );
 a39764a <=( (not A232)  and  a39763a );
 a39768a <=( (not A299)  and  (not A298) );
 a39769a <=( (not A266)  and  a39768a );
 a39770a <=( a39769a  and  a39764a );
 a39774a <=( (not A167)  and  (not A169) );
 a39775a <=( A170  and  a39774a );
 a39779a <=( (not A201)  and  (not A200) );
 a39780a <=( A166  and  a39779a );
 a39781a <=( a39780a  and  a39775a );
 a39785a <=( A265  and  A233 );
 a39786a <=( A232  and  a39785a );
 a39790a <=( (not A300)  and  (not A299) );
 a39791a <=( (not A267)  and  a39790a );
 a39792a <=( a39791a  and  a39786a );
 a39796a <=( (not A167)  and  (not A169) );
 a39797a <=( A170  and  a39796a );
 a39801a <=( (not A201)  and  (not A200) );
 a39802a <=( A166  and  a39801a );
 a39803a <=( a39802a  and  a39797a );
 a39807a <=( A265  and  A233 );
 a39808a <=( A232  and  a39807a );
 a39812a <=( A299  and  A298 );
 a39813a <=( (not A267)  and  a39812a );
 a39814a <=( a39813a  and  a39808a );
 a39818a <=( (not A167)  and  (not A169) );
 a39819a <=( A170  and  a39818a );
 a39823a <=( (not A201)  and  (not A200) );
 a39824a <=( A166  and  a39823a );
 a39825a <=( a39824a  and  a39819a );
 a39829a <=( A265  and  A233 );
 a39830a <=( A232  and  a39829a );
 a39834a <=( (not A299)  and  (not A298) );
 a39835a <=( (not A267)  and  a39834a );
 a39836a <=( a39835a  and  a39830a );
 a39840a <=( (not A167)  and  (not A169) );
 a39841a <=( A170  and  a39840a );
 a39845a <=( (not A201)  and  (not A200) );
 a39846a <=( A166  and  a39845a );
 a39847a <=( a39846a  and  a39841a );
 a39851a <=( A265  and  A233 );
 a39852a <=( A232  and  a39851a );
 a39856a <=( (not A300)  and  (not A299) );
 a39857a <=( A266  and  a39856a );
 a39858a <=( a39857a  and  a39852a );
 a39862a <=( (not A167)  and  (not A169) );
 a39863a <=( A170  and  a39862a );
 a39867a <=( (not A201)  and  (not A200) );
 a39868a <=( A166  and  a39867a );
 a39869a <=( a39868a  and  a39863a );
 a39873a <=( A265  and  A233 );
 a39874a <=( A232  and  a39873a );
 a39878a <=( A299  and  A298 );
 a39879a <=( A266  and  a39878a );
 a39880a <=( a39879a  and  a39874a );
 a39884a <=( (not A167)  and  (not A169) );
 a39885a <=( A170  and  a39884a );
 a39889a <=( (not A201)  and  (not A200) );
 a39890a <=( A166  and  a39889a );
 a39891a <=( a39890a  and  a39885a );
 a39895a <=( A265  and  A233 );
 a39896a <=( A232  and  a39895a );
 a39900a <=( (not A299)  and  (not A298) );
 a39901a <=( A266  and  a39900a );
 a39902a <=( a39901a  and  a39896a );
 a39906a <=( (not A167)  and  (not A169) );
 a39907a <=( A170  and  a39906a );
 a39911a <=( (not A201)  and  (not A200) );
 a39912a <=( A166  and  a39911a );
 a39913a <=( a39912a  and  a39907a );
 a39917a <=( (not A265)  and  A233 );
 a39918a <=( A232  and  a39917a );
 a39922a <=( (not A300)  and  (not A299) );
 a39923a <=( (not A266)  and  a39922a );
 a39924a <=( a39923a  and  a39918a );
 a39928a <=( (not A167)  and  (not A169) );
 a39929a <=( A170  and  a39928a );
 a39933a <=( (not A201)  and  (not A200) );
 a39934a <=( A166  and  a39933a );
 a39935a <=( a39934a  and  a39929a );
 a39939a <=( (not A265)  and  A233 );
 a39940a <=( A232  and  a39939a );
 a39944a <=( A299  and  A298 );
 a39945a <=( (not A266)  and  a39944a );
 a39946a <=( a39945a  and  a39940a );
 a39950a <=( (not A167)  and  (not A169) );
 a39951a <=( A170  and  a39950a );
 a39955a <=( (not A201)  and  (not A200) );
 a39956a <=( A166  and  a39955a );
 a39957a <=( a39956a  and  a39951a );
 a39961a <=( (not A265)  and  A233 );
 a39962a <=( A232  and  a39961a );
 a39966a <=( (not A299)  and  (not A298) );
 a39967a <=( (not A266)  and  a39966a );
 a39968a <=( a39967a  and  a39962a );
 a39972a <=( (not A167)  and  (not A169) );
 a39973a <=( A170  and  a39972a );
 a39977a <=( (not A201)  and  (not A200) );
 a39978a <=( A166  and  a39977a );
 a39979a <=( a39978a  and  a39973a );
 a39983a <=( A298  and  A233 );
 a39984a <=( (not A232)  and  a39983a );
 a39988a <=( A301  and  A300 );
 a39989a <=( (not A299)  and  a39988a );
 a39990a <=( a39989a  and  a39984a );
 a39994a <=( (not A167)  and  (not A169) );
 a39995a <=( A170  and  a39994a );
 a39999a <=( (not A201)  and  (not A200) );
 a40000a <=( A166  and  a39999a );
 a40001a <=( a40000a  and  a39995a );
 a40005a <=( A298  and  A233 );
 a40006a <=( (not A232)  and  a40005a );
 a40010a <=( A302  and  A300 );
 a40011a <=( (not A299)  and  a40010a );
 a40012a <=( a40011a  and  a40006a );
 a40016a <=( (not A167)  and  (not A169) );
 a40017a <=( A170  and  a40016a );
 a40021a <=( (not A201)  and  (not A200) );
 a40022a <=( A166  and  a40021a );
 a40023a <=( a40022a  and  a40017a );
 a40027a <=( A265  and  A233 );
 a40028a <=( (not A232)  and  a40027a );
 a40032a <=( A268  and  A267 );
 a40033a <=( (not A266)  and  a40032a );
 a40034a <=( a40033a  and  a40028a );
 a40038a <=( (not A167)  and  (not A169) );
 a40039a <=( A170  and  a40038a );
 a40043a <=( (not A201)  and  (not A200) );
 a40044a <=( A166  and  a40043a );
 a40045a <=( a40044a  and  a40039a );
 a40049a <=( A265  and  A233 );
 a40050a <=( (not A232)  and  a40049a );
 a40054a <=( A269  and  A267 );
 a40055a <=( (not A266)  and  a40054a );
 a40056a <=( a40055a  and  a40050a );
 a40060a <=( (not A167)  and  (not A169) );
 a40061a <=( A170  and  a40060a );
 a40065a <=( (not A201)  and  (not A200) );
 a40066a <=( A166  and  a40065a );
 a40067a <=( a40066a  and  a40061a );
 a40071a <=( A265  and  (not A234) );
 a40072a <=( (not A233)  and  a40071a );
 a40076a <=( (not A300)  and  A298 );
 a40077a <=( A266  and  a40076a );
 a40078a <=( a40077a  and  a40072a );
 a40082a <=( (not A167)  and  (not A169) );
 a40083a <=( A170  and  a40082a );
 a40087a <=( (not A201)  and  (not A200) );
 a40088a <=( A166  and  a40087a );
 a40089a <=( a40088a  and  a40083a );
 a40093a <=( A265  and  (not A234) );
 a40094a <=( (not A233)  and  a40093a );
 a40098a <=( A299  and  A298 );
 a40099a <=( A266  and  a40098a );
 a40100a <=( a40099a  and  a40094a );
 a40104a <=( (not A167)  and  (not A169) );
 a40105a <=( A170  and  a40104a );
 a40109a <=( (not A201)  and  (not A200) );
 a40110a <=( A166  and  a40109a );
 a40111a <=( a40110a  and  a40105a );
 a40115a <=( A265  and  (not A234) );
 a40116a <=( (not A233)  and  a40115a );
 a40120a <=( (not A299)  and  (not A298) );
 a40121a <=( A266  and  a40120a );
 a40122a <=( a40121a  and  a40116a );
 a40126a <=( (not A167)  and  (not A169) );
 a40127a <=( A170  and  a40126a );
 a40131a <=( (not A201)  and  (not A200) );
 a40132a <=( A166  and  a40131a );
 a40133a <=( a40132a  and  a40127a );
 a40137a <=( (not A266)  and  (not A234) );
 a40138a <=( (not A233)  and  a40137a );
 a40142a <=( (not A300)  and  A298 );
 a40143a <=( (not A267)  and  a40142a );
 a40144a <=( a40143a  and  a40138a );
 a40148a <=( (not A167)  and  (not A169) );
 a40149a <=( A170  and  a40148a );
 a40153a <=( (not A201)  and  (not A200) );
 a40154a <=( A166  and  a40153a );
 a40155a <=( a40154a  and  a40149a );
 a40159a <=( (not A266)  and  (not A234) );
 a40160a <=( (not A233)  and  a40159a );
 a40164a <=( A299  and  A298 );
 a40165a <=( (not A267)  and  a40164a );
 a40166a <=( a40165a  and  a40160a );
 a40170a <=( (not A167)  and  (not A169) );
 a40171a <=( A170  and  a40170a );
 a40175a <=( (not A201)  and  (not A200) );
 a40176a <=( A166  and  a40175a );
 a40177a <=( a40176a  and  a40171a );
 a40181a <=( (not A266)  and  (not A234) );
 a40182a <=( (not A233)  and  a40181a );
 a40186a <=( (not A299)  and  (not A298) );
 a40187a <=( (not A267)  and  a40186a );
 a40188a <=( a40187a  and  a40182a );
 a40192a <=( (not A167)  and  (not A169) );
 a40193a <=( A170  and  a40192a );
 a40197a <=( (not A201)  and  (not A200) );
 a40198a <=( A166  and  a40197a );
 a40199a <=( a40198a  and  a40193a );
 a40203a <=( (not A265)  and  (not A234) );
 a40204a <=( (not A233)  and  a40203a );
 a40208a <=( (not A300)  and  A298 );
 a40209a <=( (not A266)  and  a40208a );
 a40210a <=( a40209a  and  a40204a );
 a40214a <=( (not A167)  and  (not A169) );
 a40215a <=( A170  and  a40214a );
 a40219a <=( (not A201)  and  (not A200) );
 a40220a <=( A166  and  a40219a );
 a40221a <=( a40220a  and  a40215a );
 a40225a <=( (not A265)  and  (not A234) );
 a40226a <=( (not A233)  and  a40225a );
 a40230a <=( A299  and  A298 );
 a40231a <=( (not A266)  and  a40230a );
 a40232a <=( a40231a  and  a40226a );
 a40236a <=( (not A167)  and  (not A169) );
 a40237a <=( A170  and  a40236a );
 a40241a <=( (not A201)  and  (not A200) );
 a40242a <=( A166  and  a40241a );
 a40243a <=( a40242a  and  a40237a );
 a40247a <=( (not A265)  and  (not A234) );
 a40248a <=( (not A233)  and  a40247a );
 a40252a <=( (not A299)  and  (not A298) );
 a40253a <=( (not A266)  and  a40252a );
 a40254a <=( a40253a  and  a40248a );
 a40258a <=( (not A167)  and  (not A169) );
 a40259a <=( A170  and  a40258a );
 a40263a <=( (not A201)  and  (not A200) );
 a40264a <=( A166  and  a40263a );
 a40265a <=( a40264a  and  a40259a );
 a40269a <=( A234  and  (not A233) );
 a40270a <=( A232  and  a40269a );
 a40274a <=( A299  and  (not A298) );
 a40275a <=( A235  and  a40274a );
 a40276a <=( a40275a  and  a40270a );
 a40280a <=( (not A167)  and  (not A169) );
 a40281a <=( A170  and  a40280a );
 a40285a <=( (not A201)  and  (not A200) );
 a40286a <=( A166  and  a40285a );
 a40287a <=( a40286a  and  a40281a );
 a40291a <=( A234  and  (not A233) );
 a40292a <=( A232  and  a40291a );
 a40296a <=( A266  and  (not A265) );
 a40297a <=( A235  and  a40296a );
 a40298a <=( a40297a  and  a40292a );
 a40302a <=( (not A167)  and  (not A169) );
 a40303a <=( A170  and  a40302a );
 a40307a <=( (not A201)  and  (not A200) );
 a40308a <=( A166  and  a40307a );
 a40309a <=( a40308a  and  a40303a );
 a40313a <=( A234  and  (not A233) );
 a40314a <=( A232  and  a40313a );
 a40318a <=( A299  and  (not A298) );
 a40319a <=( A236  and  a40318a );
 a40320a <=( a40319a  and  a40314a );
 a40324a <=( (not A167)  and  (not A169) );
 a40325a <=( A170  and  a40324a );
 a40329a <=( (not A201)  and  (not A200) );
 a40330a <=( A166  and  a40329a );
 a40331a <=( a40330a  and  a40325a );
 a40335a <=( A234  and  (not A233) );
 a40336a <=( A232  and  a40335a );
 a40340a <=( A266  and  (not A265) );
 a40341a <=( A236  and  a40340a );
 a40342a <=( a40341a  and  a40336a );
 a40346a <=( (not A167)  and  (not A169) );
 a40347a <=( A170  and  a40346a );
 a40351a <=( (not A201)  and  (not A200) );
 a40352a <=( A166  and  a40351a );
 a40353a <=( a40352a  and  a40347a );
 a40357a <=( A265  and  (not A233) );
 a40358a <=( (not A232)  and  a40357a );
 a40362a <=( (not A300)  and  A298 );
 a40363a <=( A266  and  a40362a );
 a40364a <=( a40363a  and  a40358a );
 a40368a <=( (not A167)  and  (not A169) );
 a40369a <=( A170  and  a40368a );
 a40373a <=( (not A201)  and  (not A200) );
 a40374a <=( A166  and  a40373a );
 a40375a <=( a40374a  and  a40369a );
 a40379a <=( A265  and  (not A233) );
 a40380a <=( (not A232)  and  a40379a );
 a40384a <=( A299  and  A298 );
 a40385a <=( A266  and  a40384a );
 a40386a <=( a40385a  and  a40380a );
 a40390a <=( (not A167)  and  (not A169) );
 a40391a <=( A170  and  a40390a );
 a40395a <=( (not A201)  and  (not A200) );
 a40396a <=( A166  and  a40395a );
 a40397a <=( a40396a  and  a40391a );
 a40401a <=( A265  and  (not A233) );
 a40402a <=( (not A232)  and  a40401a );
 a40406a <=( (not A299)  and  (not A298) );
 a40407a <=( A266  and  a40406a );
 a40408a <=( a40407a  and  a40402a );
 a40412a <=( (not A167)  and  (not A169) );
 a40413a <=( A170  and  a40412a );
 a40417a <=( (not A201)  and  (not A200) );
 a40418a <=( A166  and  a40417a );
 a40419a <=( a40418a  and  a40413a );
 a40423a <=( (not A266)  and  (not A233) );
 a40424a <=( (not A232)  and  a40423a );
 a40428a <=( (not A300)  and  A298 );
 a40429a <=( (not A267)  and  a40428a );
 a40430a <=( a40429a  and  a40424a );
 a40434a <=( (not A167)  and  (not A169) );
 a40435a <=( A170  and  a40434a );
 a40439a <=( (not A201)  and  (not A200) );
 a40440a <=( A166  and  a40439a );
 a40441a <=( a40440a  and  a40435a );
 a40445a <=( (not A266)  and  (not A233) );
 a40446a <=( (not A232)  and  a40445a );
 a40450a <=( A299  and  A298 );
 a40451a <=( (not A267)  and  a40450a );
 a40452a <=( a40451a  and  a40446a );
 a40456a <=( (not A167)  and  (not A169) );
 a40457a <=( A170  and  a40456a );
 a40461a <=( (not A201)  and  (not A200) );
 a40462a <=( A166  and  a40461a );
 a40463a <=( a40462a  and  a40457a );
 a40467a <=( (not A266)  and  (not A233) );
 a40468a <=( (not A232)  and  a40467a );
 a40472a <=( (not A299)  and  (not A298) );
 a40473a <=( (not A267)  and  a40472a );
 a40474a <=( a40473a  and  a40468a );
 a40478a <=( (not A167)  and  (not A169) );
 a40479a <=( A170  and  a40478a );
 a40483a <=( (not A201)  and  (not A200) );
 a40484a <=( A166  and  a40483a );
 a40485a <=( a40484a  and  a40479a );
 a40489a <=( (not A265)  and  (not A233) );
 a40490a <=( (not A232)  and  a40489a );
 a40494a <=( (not A300)  and  A298 );
 a40495a <=( (not A266)  and  a40494a );
 a40496a <=( a40495a  and  a40490a );
 a40500a <=( (not A167)  and  (not A169) );
 a40501a <=( A170  and  a40500a );
 a40505a <=( (not A201)  and  (not A200) );
 a40506a <=( A166  and  a40505a );
 a40507a <=( a40506a  and  a40501a );
 a40511a <=( (not A265)  and  (not A233) );
 a40512a <=( (not A232)  and  a40511a );
 a40516a <=( A299  and  A298 );
 a40517a <=( (not A266)  and  a40516a );
 a40518a <=( a40517a  and  a40512a );
 a40522a <=( (not A167)  and  (not A169) );
 a40523a <=( A170  and  a40522a );
 a40527a <=( (not A201)  and  (not A200) );
 a40528a <=( A166  and  a40527a );
 a40529a <=( a40528a  and  a40523a );
 a40533a <=( (not A265)  and  (not A233) );
 a40534a <=( (not A232)  and  a40533a );
 a40538a <=( (not A299)  and  (not A298) );
 a40539a <=( (not A266)  and  a40538a );
 a40540a <=( a40539a  and  a40534a );
 a40544a <=( (not A167)  and  (not A169) );
 a40545a <=( A170  and  a40544a );
 a40549a <=( (not A200)  and  (not A199) );
 a40550a <=( A166  and  a40549a );
 a40551a <=( a40550a  and  a40545a );
 a40555a <=( A265  and  A233 );
 a40556a <=( A232  and  a40555a );
 a40560a <=( (not A300)  and  (not A299) );
 a40561a <=( (not A267)  and  a40560a );
 a40562a <=( a40561a  and  a40556a );
 a40566a <=( (not A167)  and  (not A169) );
 a40567a <=( A170  and  a40566a );
 a40571a <=( (not A200)  and  (not A199) );
 a40572a <=( A166  and  a40571a );
 a40573a <=( a40572a  and  a40567a );
 a40577a <=( A265  and  A233 );
 a40578a <=( A232  and  a40577a );
 a40582a <=( A299  and  A298 );
 a40583a <=( (not A267)  and  a40582a );
 a40584a <=( a40583a  and  a40578a );
 a40588a <=( (not A167)  and  (not A169) );
 a40589a <=( A170  and  a40588a );
 a40593a <=( (not A200)  and  (not A199) );
 a40594a <=( A166  and  a40593a );
 a40595a <=( a40594a  and  a40589a );
 a40599a <=( A265  and  A233 );
 a40600a <=( A232  and  a40599a );
 a40604a <=( (not A299)  and  (not A298) );
 a40605a <=( (not A267)  and  a40604a );
 a40606a <=( a40605a  and  a40600a );
 a40610a <=( (not A167)  and  (not A169) );
 a40611a <=( A170  and  a40610a );
 a40615a <=( (not A200)  and  (not A199) );
 a40616a <=( A166  and  a40615a );
 a40617a <=( a40616a  and  a40611a );
 a40621a <=( A265  and  A233 );
 a40622a <=( A232  and  a40621a );
 a40626a <=( (not A300)  and  (not A299) );
 a40627a <=( A266  and  a40626a );
 a40628a <=( a40627a  and  a40622a );
 a40632a <=( (not A167)  and  (not A169) );
 a40633a <=( A170  and  a40632a );
 a40637a <=( (not A200)  and  (not A199) );
 a40638a <=( A166  and  a40637a );
 a40639a <=( a40638a  and  a40633a );
 a40643a <=( A265  and  A233 );
 a40644a <=( A232  and  a40643a );
 a40648a <=( A299  and  A298 );
 a40649a <=( A266  and  a40648a );
 a40650a <=( a40649a  and  a40644a );
 a40654a <=( (not A167)  and  (not A169) );
 a40655a <=( A170  and  a40654a );
 a40659a <=( (not A200)  and  (not A199) );
 a40660a <=( A166  and  a40659a );
 a40661a <=( a40660a  and  a40655a );
 a40665a <=( A265  and  A233 );
 a40666a <=( A232  and  a40665a );
 a40670a <=( (not A299)  and  (not A298) );
 a40671a <=( A266  and  a40670a );
 a40672a <=( a40671a  and  a40666a );
 a40676a <=( (not A167)  and  (not A169) );
 a40677a <=( A170  and  a40676a );
 a40681a <=( (not A200)  and  (not A199) );
 a40682a <=( A166  and  a40681a );
 a40683a <=( a40682a  and  a40677a );
 a40687a <=( (not A265)  and  A233 );
 a40688a <=( A232  and  a40687a );
 a40692a <=( (not A300)  and  (not A299) );
 a40693a <=( (not A266)  and  a40692a );
 a40694a <=( a40693a  and  a40688a );
 a40698a <=( (not A167)  and  (not A169) );
 a40699a <=( A170  and  a40698a );
 a40703a <=( (not A200)  and  (not A199) );
 a40704a <=( A166  and  a40703a );
 a40705a <=( a40704a  and  a40699a );
 a40709a <=( (not A265)  and  A233 );
 a40710a <=( A232  and  a40709a );
 a40714a <=( A299  and  A298 );
 a40715a <=( (not A266)  and  a40714a );
 a40716a <=( a40715a  and  a40710a );
 a40720a <=( (not A167)  and  (not A169) );
 a40721a <=( A170  and  a40720a );
 a40725a <=( (not A200)  and  (not A199) );
 a40726a <=( A166  and  a40725a );
 a40727a <=( a40726a  and  a40721a );
 a40731a <=( (not A265)  and  A233 );
 a40732a <=( A232  and  a40731a );
 a40736a <=( (not A299)  and  (not A298) );
 a40737a <=( (not A266)  and  a40736a );
 a40738a <=( a40737a  and  a40732a );
 a40742a <=( (not A167)  and  (not A169) );
 a40743a <=( A170  and  a40742a );
 a40747a <=( (not A200)  and  (not A199) );
 a40748a <=( A166  and  a40747a );
 a40749a <=( a40748a  and  a40743a );
 a40753a <=( A298  and  A233 );
 a40754a <=( (not A232)  and  a40753a );
 a40758a <=( A301  and  A300 );
 a40759a <=( (not A299)  and  a40758a );
 a40760a <=( a40759a  and  a40754a );
 a40764a <=( (not A167)  and  (not A169) );
 a40765a <=( A170  and  a40764a );
 a40769a <=( (not A200)  and  (not A199) );
 a40770a <=( A166  and  a40769a );
 a40771a <=( a40770a  and  a40765a );
 a40775a <=( A298  and  A233 );
 a40776a <=( (not A232)  and  a40775a );
 a40780a <=( A302  and  A300 );
 a40781a <=( (not A299)  and  a40780a );
 a40782a <=( a40781a  and  a40776a );
 a40786a <=( (not A167)  and  (not A169) );
 a40787a <=( A170  and  a40786a );
 a40791a <=( (not A200)  and  (not A199) );
 a40792a <=( A166  and  a40791a );
 a40793a <=( a40792a  and  a40787a );
 a40797a <=( A265  and  A233 );
 a40798a <=( (not A232)  and  a40797a );
 a40802a <=( A268  and  A267 );
 a40803a <=( (not A266)  and  a40802a );
 a40804a <=( a40803a  and  a40798a );
 a40808a <=( (not A167)  and  (not A169) );
 a40809a <=( A170  and  a40808a );
 a40813a <=( (not A200)  and  (not A199) );
 a40814a <=( A166  and  a40813a );
 a40815a <=( a40814a  and  a40809a );
 a40819a <=( A265  and  A233 );
 a40820a <=( (not A232)  and  a40819a );
 a40824a <=( A269  and  A267 );
 a40825a <=( (not A266)  and  a40824a );
 a40826a <=( a40825a  and  a40820a );
 a40830a <=( (not A167)  and  (not A169) );
 a40831a <=( A170  and  a40830a );
 a40835a <=( (not A200)  and  (not A199) );
 a40836a <=( A166  and  a40835a );
 a40837a <=( a40836a  and  a40831a );
 a40841a <=( A265  and  (not A234) );
 a40842a <=( (not A233)  and  a40841a );
 a40846a <=( (not A300)  and  A298 );
 a40847a <=( A266  and  a40846a );
 a40848a <=( a40847a  and  a40842a );
 a40852a <=( (not A167)  and  (not A169) );
 a40853a <=( A170  and  a40852a );
 a40857a <=( (not A200)  and  (not A199) );
 a40858a <=( A166  and  a40857a );
 a40859a <=( a40858a  and  a40853a );
 a40863a <=( A265  and  (not A234) );
 a40864a <=( (not A233)  and  a40863a );
 a40868a <=( A299  and  A298 );
 a40869a <=( A266  and  a40868a );
 a40870a <=( a40869a  and  a40864a );
 a40874a <=( (not A167)  and  (not A169) );
 a40875a <=( A170  and  a40874a );
 a40879a <=( (not A200)  and  (not A199) );
 a40880a <=( A166  and  a40879a );
 a40881a <=( a40880a  and  a40875a );
 a40885a <=( A265  and  (not A234) );
 a40886a <=( (not A233)  and  a40885a );
 a40890a <=( (not A299)  and  (not A298) );
 a40891a <=( A266  and  a40890a );
 a40892a <=( a40891a  and  a40886a );
 a40896a <=( (not A167)  and  (not A169) );
 a40897a <=( A170  and  a40896a );
 a40901a <=( (not A200)  and  (not A199) );
 a40902a <=( A166  and  a40901a );
 a40903a <=( a40902a  and  a40897a );
 a40907a <=( (not A266)  and  (not A234) );
 a40908a <=( (not A233)  and  a40907a );
 a40912a <=( (not A300)  and  A298 );
 a40913a <=( (not A267)  and  a40912a );
 a40914a <=( a40913a  and  a40908a );
 a40918a <=( (not A167)  and  (not A169) );
 a40919a <=( A170  and  a40918a );
 a40923a <=( (not A200)  and  (not A199) );
 a40924a <=( A166  and  a40923a );
 a40925a <=( a40924a  and  a40919a );
 a40929a <=( (not A266)  and  (not A234) );
 a40930a <=( (not A233)  and  a40929a );
 a40934a <=( A299  and  A298 );
 a40935a <=( (not A267)  and  a40934a );
 a40936a <=( a40935a  and  a40930a );
 a40940a <=( (not A167)  and  (not A169) );
 a40941a <=( A170  and  a40940a );
 a40945a <=( (not A200)  and  (not A199) );
 a40946a <=( A166  and  a40945a );
 a40947a <=( a40946a  and  a40941a );
 a40951a <=( (not A266)  and  (not A234) );
 a40952a <=( (not A233)  and  a40951a );
 a40956a <=( (not A299)  and  (not A298) );
 a40957a <=( (not A267)  and  a40956a );
 a40958a <=( a40957a  and  a40952a );
 a40962a <=( (not A167)  and  (not A169) );
 a40963a <=( A170  and  a40962a );
 a40967a <=( (not A200)  and  (not A199) );
 a40968a <=( A166  and  a40967a );
 a40969a <=( a40968a  and  a40963a );
 a40973a <=( (not A265)  and  (not A234) );
 a40974a <=( (not A233)  and  a40973a );
 a40978a <=( (not A300)  and  A298 );
 a40979a <=( (not A266)  and  a40978a );
 a40980a <=( a40979a  and  a40974a );
 a40984a <=( (not A167)  and  (not A169) );
 a40985a <=( A170  and  a40984a );
 a40989a <=( (not A200)  and  (not A199) );
 a40990a <=( A166  and  a40989a );
 a40991a <=( a40990a  and  a40985a );
 a40995a <=( (not A265)  and  (not A234) );
 a40996a <=( (not A233)  and  a40995a );
 a41000a <=( A299  and  A298 );
 a41001a <=( (not A266)  and  a41000a );
 a41002a <=( a41001a  and  a40996a );
 a41006a <=( (not A167)  and  (not A169) );
 a41007a <=( A170  and  a41006a );
 a41011a <=( (not A200)  and  (not A199) );
 a41012a <=( A166  and  a41011a );
 a41013a <=( a41012a  and  a41007a );
 a41017a <=( (not A265)  and  (not A234) );
 a41018a <=( (not A233)  and  a41017a );
 a41022a <=( (not A299)  and  (not A298) );
 a41023a <=( (not A266)  and  a41022a );
 a41024a <=( a41023a  and  a41018a );
 a41028a <=( (not A167)  and  (not A169) );
 a41029a <=( A170  and  a41028a );
 a41033a <=( (not A200)  and  (not A199) );
 a41034a <=( A166  and  a41033a );
 a41035a <=( a41034a  and  a41029a );
 a41039a <=( A234  and  (not A233) );
 a41040a <=( A232  and  a41039a );
 a41044a <=( A299  and  (not A298) );
 a41045a <=( A235  and  a41044a );
 a41046a <=( a41045a  and  a41040a );
 a41050a <=( (not A167)  and  (not A169) );
 a41051a <=( A170  and  a41050a );
 a41055a <=( (not A200)  and  (not A199) );
 a41056a <=( A166  and  a41055a );
 a41057a <=( a41056a  and  a41051a );
 a41061a <=( A234  and  (not A233) );
 a41062a <=( A232  and  a41061a );
 a41066a <=( A266  and  (not A265) );
 a41067a <=( A235  and  a41066a );
 a41068a <=( a41067a  and  a41062a );
 a41072a <=( (not A167)  and  (not A169) );
 a41073a <=( A170  and  a41072a );
 a41077a <=( (not A200)  and  (not A199) );
 a41078a <=( A166  and  a41077a );
 a41079a <=( a41078a  and  a41073a );
 a41083a <=( A234  and  (not A233) );
 a41084a <=( A232  and  a41083a );
 a41088a <=( A299  and  (not A298) );
 a41089a <=( A236  and  a41088a );
 a41090a <=( a41089a  and  a41084a );
 a41094a <=( (not A167)  and  (not A169) );
 a41095a <=( A170  and  a41094a );
 a41099a <=( (not A200)  and  (not A199) );
 a41100a <=( A166  and  a41099a );
 a41101a <=( a41100a  and  a41095a );
 a41105a <=( A234  and  (not A233) );
 a41106a <=( A232  and  a41105a );
 a41110a <=( A266  and  (not A265) );
 a41111a <=( A236  and  a41110a );
 a41112a <=( a41111a  and  a41106a );
 a41116a <=( (not A167)  and  (not A169) );
 a41117a <=( A170  and  a41116a );
 a41121a <=( (not A200)  and  (not A199) );
 a41122a <=( A166  and  a41121a );
 a41123a <=( a41122a  and  a41117a );
 a41127a <=( A265  and  (not A233) );
 a41128a <=( (not A232)  and  a41127a );
 a41132a <=( (not A300)  and  A298 );
 a41133a <=( A266  and  a41132a );
 a41134a <=( a41133a  and  a41128a );
 a41138a <=( (not A167)  and  (not A169) );
 a41139a <=( A170  and  a41138a );
 a41143a <=( (not A200)  and  (not A199) );
 a41144a <=( A166  and  a41143a );
 a41145a <=( a41144a  and  a41139a );
 a41149a <=( A265  and  (not A233) );
 a41150a <=( (not A232)  and  a41149a );
 a41154a <=( A299  and  A298 );
 a41155a <=( A266  and  a41154a );
 a41156a <=( a41155a  and  a41150a );
 a41160a <=( (not A167)  and  (not A169) );
 a41161a <=( A170  and  a41160a );
 a41165a <=( (not A200)  and  (not A199) );
 a41166a <=( A166  and  a41165a );
 a41167a <=( a41166a  and  a41161a );
 a41171a <=( A265  and  (not A233) );
 a41172a <=( (not A232)  and  a41171a );
 a41176a <=( (not A299)  and  (not A298) );
 a41177a <=( A266  and  a41176a );
 a41178a <=( a41177a  and  a41172a );
 a41182a <=( (not A167)  and  (not A169) );
 a41183a <=( A170  and  a41182a );
 a41187a <=( (not A200)  and  (not A199) );
 a41188a <=( A166  and  a41187a );
 a41189a <=( a41188a  and  a41183a );
 a41193a <=( (not A266)  and  (not A233) );
 a41194a <=( (not A232)  and  a41193a );
 a41198a <=( (not A300)  and  A298 );
 a41199a <=( (not A267)  and  a41198a );
 a41200a <=( a41199a  and  a41194a );
 a41204a <=( (not A167)  and  (not A169) );
 a41205a <=( A170  and  a41204a );
 a41209a <=( (not A200)  and  (not A199) );
 a41210a <=( A166  and  a41209a );
 a41211a <=( a41210a  and  a41205a );
 a41215a <=( (not A266)  and  (not A233) );
 a41216a <=( (not A232)  and  a41215a );
 a41220a <=( A299  and  A298 );
 a41221a <=( (not A267)  and  a41220a );
 a41222a <=( a41221a  and  a41216a );
 a41226a <=( (not A167)  and  (not A169) );
 a41227a <=( A170  and  a41226a );
 a41231a <=( (not A200)  and  (not A199) );
 a41232a <=( A166  and  a41231a );
 a41233a <=( a41232a  and  a41227a );
 a41237a <=( (not A266)  and  (not A233) );
 a41238a <=( (not A232)  and  a41237a );
 a41242a <=( (not A299)  and  (not A298) );
 a41243a <=( (not A267)  and  a41242a );
 a41244a <=( a41243a  and  a41238a );
 a41248a <=( (not A167)  and  (not A169) );
 a41249a <=( A170  and  a41248a );
 a41253a <=( (not A200)  and  (not A199) );
 a41254a <=( A166  and  a41253a );
 a41255a <=( a41254a  and  a41249a );
 a41259a <=( (not A265)  and  (not A233) );
 a41260a <=( (not A232)  and  a41259a );
 a41264a <=( (not A300)  and  A298 );
 a41265a <=( (not A266)  and  a41264a );
 a41266a <=( a41265a  and  a41260a );
 a41270a <=( (not A167)  and  (not A169) );
 a41271a <=( A170  and  a41270a );
 a41275a <=( (not A200)  and  (not A199) );
 a41276a <=( A166  and  a41275a );
 a41277a <=( a41276a  and  a41271a );
 a41281a <=( (not A265)  and  (not A233) );
 a41282a <=( (not A232)  and  a41281a );
 a41286a <=( A299  and  A298 );
 a41287a <=( (not A266)  and  a41286a );
 a41288a <=( a41287a  and  a41282a );
 a41292a <=( (not A167)  and  (not A169) );
 a41293a <=( A170  and  a41292a );
 a41297a <=( (not A200)  and  (not A199) );
 a41298a <=( A166  and  a41297a );
 a41299a <=( a41298a  and  a41293a );
 a41303a <=( (not A265)  and  (not A233) );
 a41304a <=( (not A232)  and  a41303a );
 a41308a <=( (not A299)  and  (not A298) );
 a41309a <=( (not A266)  and  a41308a );
 a41310a <=( a41309a  and  a41304a );
 a41314a <=( A199  and  A166 );
 a41315a <=( A168  and  a41314a );
 a41319a <=( (not A235)  and  (not A233) );
 a41320a <=( A200  and  a41319a );
 a41321a <=( a41320a  and  a41315a );
 a41325a <=( (not A268)  and  (not A266) );
 a41326a <=( (not A236)  and  a41325a );
 a41329a <=( A298  and  (not A269) );
 a41332a <=( (not A302)  and  (not A301) );
 a41333a <=( a41332a  and  a41329a );
 a41334a <=( a41333a  and  a41326a );
 a41338a <=( (not A200)  and  A166 );
 a41339a <=( A168  and  a41338a );
 a41343a <=( A232  and  (not A203) );
 a41344a <=( (not A202)  and  a41343a );
 a41345a <=( a41344a  and  a41339a );
 a41349a <=( (not A268)  and  A265 );
 a41350a <=( A233  and  a41349a );
 a41353a <=( (not A299)  and  (not A269) );
 a41356a <=( (not A302)  and  (not A301) );
 a41357a <=( a41356a  and  a41353a );
 a41358a <=( a41357a  and  a41350a );
 a41362a <=( (not A200)  and  A166 );
 a41363a <=( A168  and  a41362a );
 a41367a <=( (not A233)  and  (not A203) );
 a41368a <=( (not A202)  and  a41367a );
 a41369a <=( a41368a  and  a41363a );
 a41373a <=( A265  and  (not A236) );
 a41374a <=( (not A235)  and  a41373a );
 a41377a <=( A298  and  A266 );
 a41380a <=( (not A302)  and  (not A301) );
 a41381a <=( a41380a  and  a41377a );
 a41382a <=( a41381a  and  a41374a );
 a41386a <=( (not A200)  and  A166 );
 a41387a <=( A168  and  a41386a );
 a41391a <=( (not A233)  and  (not A203) );
 a41392a <=( (not A202)  and  a41391a );
 a41393a <=( a41392a  and  a41387a );
 a41397a <=( (not A266)  and  (not A236) );
 a41398a <=( (not A235)  and  a41397a );
 a41401a <=( (not A269)  and  (not A268) );
 a41404a <=( (not A300)  and  A298 );
 a41405a <=( a41404a  and  a41401a );
 a41406a <=( a41405a  and  a41398a );
 a41410a <=( (not A200)  and  A166 );
 a41411a <=( A168  and  a41410a );
 a41415a <=( (not A233)  and  (not A203) );
 a41416a <=( (not A202)  and  a41415a );
 a41417a <=( a41416a  and  a41411a );
 a41421a <=( (not A266)  and  (not A236) );
 a41422a <=( (not A235)  and  a41421a );
 a41425a <=( (not A269)  and  (not A268) );
 a41428a <=( A299  and  A298 );
 a41429a <=( a41428a  and  a41425a );
 a41430a <=( a41429a  and  a41422a );
 a41434a <=( (not A200)  and  A166 );
 a41435a <=( A168  and  a41434a );
 a41439a <=( (not A233)  and  (not A203) );
 a41440a <=( (not A202)  and  a41439a );
 a41441a <=( a41440a  and  a41435a );
 a41445a <=( (not A266)  and  (not A236) );
 a41446a <=( (not A235)  and  a41445a );
 a41449a <=( (not A269)  and  (not A268) );
 a41452a <=( (not A299)  and  (not A298) );
 a41453a <=( a41452a  and  a41449a );
 a41454a <=( a41453a  and  a41446a );
 a41458a <=( (not A200)  and  A166 );
 a41459a <=( A168  and  a41458a );
 a41463a <=( (not A233)  and  (not A203) );
 a41464a <=( (not A202)  and  a41463a );
 a41465a <=( a41464a  and  a41459a );
 a41469a <=( (not A266)  and  (not A236) );
 a41470a <=( (not A235)  and  a41469a );
 a41473a <=( A298  and  (not A267) );
 a41476a <=( (not A302)  and  (not A301) );
 a41477a <=( a41476a  and  a41473a );
 a41478a <=( a41477a  and  a41470a );
 a41482a <=( (not A200)  and  A166 );
 a41483a <=( A168  and  a41482a );
 a41487a <=( (not A233)  and  (not A203) );
 a41488a <=( (not A202)  and  a41487a );
 a41489a <=( a41488a  and  a41483a );
 a41493a <=( (not A265)  and  (not A236) );
 a41494a <=( (not A235)  and  a41493a );
 a41497a <=( A298  and  (not A266) );
 a41500a <=( (not A302)  and  (not A301) );
 a41501a <=( a41500a  and  a41497a );
 a41502a <=( a41501a  and  a41494a );
 a41506a <=( (not A200)  and  A166 );
 a41507a <=( A168  and  a41506a );
 a41511a <=( (not A233)  and  (not A203) );
 a41512a <=( (not A202)  and  a41511a );
 a41513a <=( a41512a  and  a41507a );
 a41517a <=( (not A268)  and  (not A266) );
 a41518a <=( (not A234)  and  a41517a );
 a41521a <=( A298  and  (not A269) );
 a41524a <=( (not A302)  and  (not A301) );
 a41525a <=( a41524a  and  a41521a );
 a41526a <=( a41525a  and  a41518a );
 a41530a <=( (not A200)  and  A166 );
 a41531a <=( A168  and  a41530a );
 a41535a <=( A232  and  (not A203) );
 a41536a <=( (not A202)  and  a41535a );
 a41537a <=( a41536a  and  a41531a );
 a41541a <=( A235  and  A234 );
 a41542a <=( (not A233)  and  a41541a );
 a41545a <=( (not A299)  and  A298 );
 a41548a <=( A301  and  A300 );
 a41549a <=( a41548a  and  a41545a );
 a41550a <=( a41549a  and  a41542a );
 a41554a <=( (not A200)  and  A166 );
 a41555a <=( A168  and  a41554a );
 a41559a <=( A232  and  (not A203) );
 a41560a <=( (not A202)  and  a41559a );
 a41561a <=( a41560a  and  a41555a );
 a41565a <=( A235  and  A234 );
 a41566a <=( (not A233)  and  a41565a );
 a41569a <=( (not A299)  and  A298 );
 a41572a <=( A302  and  A300 );
 a41573a <=( a41572a  and  a41569a );
 a41574a <=( a41573a  and  a41566a );
 a41578a <=( (not A200)  and  A166 );
 a41579a <=( A168  and  a41578a );
 a41583a <=( A232  and  (not A203) );
 a41584a <=( (not A202)  and  a41583a );
 a41585a <=( a41584a  and  a41579a );
 a41589a <=( A235  and  A234 );
 a41590a <=( (not A233)  and  a41589a );
 a41593a <=( (not A266)  and  A265 );
 a41596a <=( A268  and  A267 );
 a41597a <=( a41596a  and  a41593a );
 a41598a <=( a41597a  and  a41590a );
 a41602a <=( (not A200)  and  A166 );
 a41603a <=( A168  and  a41602a );
 a41607a <=( A232  and  (not A203) );
 a41608a <=( (not A202)  and  a41607a );
 a41609a <=( a41608a  and  a41603a );
 a41613a <=( A235  and  A234 );
 a41614a <=( (not A233)  and  a41613a );
 a41617a <=( (not A266)  and  A265 );
 a41620a <=( A269  and  A267 );
 a41621a <=( a41620a  and  a41617a );
 a41622a <=( a41621a  and  a41614a );
 a41626a <=( (not A200)  and  A166 );
 a41627a <=( A168  and  a41626a );
 a41631a <=( A232  and  (not A203) );
 a41632a <=( (not A202)  and  a41631a );
 a41633a <=( a41632a  and  a41627a );
 a41637a <=( A236  and  A234 );
 a41638a <=( (not A233)  and  a41637a );
 a41641a <=( (not A299)  and  A298 );
 a41644a <=( A301  and  A300 );
 a41645a <=( a41644a  and  a41641a );
 a41646a <=( a41645a  and  a41638a );
 a41650a <=( (not A200)  and  A166 );
 a41651a <=( A168  and  a41650a );
 a41655a <=( A232  and  (not A203) );
 a41656a <=( (not A202)  and  a41655a );
 a41657a <=( a41656a  and  a41651a );
 a41661a <=( A236  and  A234 );
 a41662a <=( (not A233)  and  a41661a );
 a41665a <=( (not A299)  and  A298 );
 a41668a <=( A302  and  A300 );
 a41669a <=( a41668a  and  a41665a );
 a41670a <=( a41669a  and  a41662a );
 a41674a <=( (not A200)  and  A166 );
 a41675a <=( A168  and  a41674a );
 a41679a <=( A232  and  (not A203) );
 a41680a <=( (not A202)  and  a41679a );
 a41681a <=( a41680a  and  a41675a );
 a41685a <=( A236  and  A234 );
 a41686a <=( (not A233)  and  a41685a );
 a41689a <=( (not A266)  and  A265 );
 a41692a <=( A268  and  A267 );
 a41693a <=( a41692a  and  a41689a );
 a41694a <=( a41693a  and  a41686a );
 a41698a <=( (not A200)  and  A166 );
 a41699a <=( A168  and  a41698a );
 a41703a <=( A232  and  (not A203) );
 a41704a <=( (not A202)  and  a41703a );
 a41705a <=( a41704a  and  a41699a );
 a41709a <=( A236  and  A234 );
 a41710a <=( (not A233)  and  a41709a );
 a41713a <=( (not A266)  and  A265 );
 a41716a <=( A269  and  A267 );
 a41717a <=( a41716a  and  a41713a );
 a41718a <=( a41717a  and  a41710a );
 a41722a <=( (not A200)  and  A166 );
 a41723a <=( A168  and  a41722a );
 a41727a <=( (not A232)  and  (not A203) );
 a41728a <=( (not A202)  and  a41727a );
 a41729a <=( a41728a  and  a41723a );
 a41733a <=( (not A268)  and  (not A266) );
 a41734a <=( (not A233)  and  a41733a );
 a41737a <=( A298  and  (not A269) );
 a41740a <=( (not A302)  and  (not A301) );
 a41741a <=( a41740a  and  a41737a );
 a41742a <=( a41741a  and  a41734a );
 a41746a <=( (not A200)  and  A166 );
 a41747a <=( A168  and  a41746a );
 a41751a <=( (not A235)  and  (not A233) );
 a41752a <=( (not A201)  and  a41751a );
 a41753a <=( a41752a  and  a41747a );
 a41757a <=( (not A268)  and  (not A266) );
 a41758a <=( (not A236)  and  a41757a );
 a41761a <=( A298  and  (not A269) );
 a41764a <=( (not A302)  and  (not A301) );
 a41765a <=( a41764a  and  a41761a );
 a41766a <=( a41765a  and  a41758a );
 a41770a <=( (not A199)  and  A166 );
 a41771a <=( A168  and  a41770a );
 a41775a <=( (not A235)  and  (not A233) );
 a41776a <=( (not A200)  and  a41775a );
 a41777a <=( a41776a  and  a41771a );
 a41781a <=( (not A268)  and  (not A266) );
 a41782a <=( (not A236)  and  a41781a );
 a41785a <=( A298  and  (not A269) );
 a41788a <=( (not A302)  and  (not A301) );
 a41789a <=( a41788a  and  a41785a );
 a41790a <=( a41789a  and  a41782a );
 a41794a <=( A199  and  A167 );
 a41795a <=( A168  and  a41794a );
 a41799a <=( (not A235)  and  (not A233) );
 a41800a <=( A200  and  a41799a );
 a41801a <=( a41800a  and  a41795a );
 a41805a <=( (not A268)  and  (not A266) );
 a41806a <=( (not A236)  and  a41805a );
 a41809a <=( A298  and  (not A269) );
 a41812a <=( (not A302)  and  (not A301) );
 a41813a <=( a41812a  and  a41809a );
 a41814a <=( a41813a  and  a41806a );
 a41818a <=( (not A200)  and  A167 );
 a41819a <=( A168  and  a41818a );
 a41823a <=( A232  and  (not A203) );
 a41824a <=( (not A202)  and  a41823a );
 a41825a <=( a41824a  and  a41819a );
 a41829a <=( (not A268)  and  A265 );
 a41830a <=( A233  and  a41829a );
 a41833a <=( (not A299)  and  (not A269) );
 a41836a <=( (not A302)  and  (not A301) );
 a41837a <=( a41836a  and  a41833a );
 a41838a <=( a41837a  and  a41830a );
 a41842a <=( (not A200)  and  A167 );
 a41843a <=( A168  and  a41842a );
 a41847a <=( (not A233)  and  (not A203) );
 a41848a <=( (not A202)  and  a41847a );
 a41849a <=( a41848a  and  a41843a );
 a41853a <=( A265  and  (not A236) );
 a41854a <=( (not A235)  and  a41853a );
 a41857a <=( A298  and  A266 );
 a41860a <=( (not A302)  and  (not A301) );
 a41861a <=( a41860a  and  a41857a );
 a41862a <=( a41861a  and  a41854a );
 a41866a <=( (not A200)  and  A167 );
 a41867a <=( A168  and  a41866a );
 a41871a <=( (not A233)  and  (not A203) );
 a41872a <=( (not A202)  and  a41871a );
 a41873a <=( a41872a  and  a41867a );
 a41877a <=( (not A266)  and  (not A236) );
 a41878a <=( (not A235)  and  a41877a );
 a41881a <=( (not A269)  and  (not A268) );
 a41884a <=( (not A300)  and  A298 );
 a41885a <=( a41884a  and  a41881a );
 a41886a <=( a41885a  and  a41878a );
 a41890a <=( (not A200)  and  A167 );
 a41891a <=( A168  and  a41890a );
 a41895a <=( (not A233)  and  (not A203) );
 a41896a <=( (not A202)  and  a41895a );
 a41897a <=( a41896a  and  a41891a );
 a41901a <=( (not A266)  and  (not A236) );
 a41902a <=( (not A235)  and  a41901a );
 a41905a <=( (not A269)  and  (not A268) );
 a41908a <=( A299  and  A298 );
 a41909a <=( a41908a  and  a41905a );
 a41910a <=( a41909a  and  a41902a );
 a41914a <=( (not A200)  and  A167 );
 a41915a <=( A168  and  a41914a );
 a41919a <=( (not A233)  and  (not A203) );
 a41920a <=( (not A202)  and  a41919a );
 a41921a <=( a41920a  and  a41915a );
 a41925a <=( (not A266)  and  (not A236) );
 a41926a <=( (not A235)  and  a41925a );
 a41929a <=( (not A269)  and  (not A268) );
 a41932a <=( (not A299)  and  (not A298) );
 a41933a <=( a41932a  and  a41929a );
 a41934a <=( a41933a  and  a41926a );
 a41938a <=( (not A200)  and  A167 );
 a41939a <=( A168  and  a41938a );
 a41943a <=( (not A233)  and  (not A203) );
 a41944a <=( (not A202)  and  a41943a );
 a41945a <=( a41944a  and  a41939a );
 a41949a <=( (not A266)  and  (not A236) );
 a41950a <=( (not A235)  and  a41949a );
 a41953a <=( A298  and  (not A267) );
 a41956a <=( (not A302)  and  (not A301) );
 a41957a <=( a41956a  and  a41953a );
 a41958a <=( a41957a  and  a41950a );
 a41962a <=( (not A200)  and  A167 );
 a41963a <=( A168  and  a41962a );
 a41967a <=( (not A233)  and  (not A203) );
 a41968a <=( (not A202)  and  a41967a );
 a41969a <=( a41968a  and  a41963a );
 a41973a <=( (not A265)  and  (not A236) );
 a41974a <=( (not A235)  and  a41973a );
 a41977a <=( A298  and  (not A266) );
 a41980a <=( (not A302)  and  (not A301) );
 a41981a <=( a41980a  and  a41977a );
 a41982a <=( a41981a  and  a41974a );
 a41986a <=( (not A200)  and  A167 );
 a41987a <=( A168  and  a41986a );
 a41991a <=( (not A233)  and  (not A203) );
 a41992a <=( (not A202)  and  a41991a );
 a41993a <=( a41992a  and  a41987a );
 a41997a <=( (not A268)  and  (not A266) );
 a41998a <=( (not A234)  and  a41997a );
 a42001a <=( A298  and  (not A269) );
 a42004a <=( (not A302)  and  (not A301) );
 a42005a <=( a42004a  and  a42001a );
 a42006a <=( a42005a  and  a41998a );
 a42010a <=( (not A200)  and  A167 );
 a42011a <=( A168  and  a42010a );
 a42015a <=( A232  and  (not A203) );
 a42016a <=( (not A202)  and  a42015a );
 a42017a <=( a42016a  and  a42011a );
 a42021a <=( A235  and  A234 );
 a42022a <=( (not A233)  and  a42021a );
 a42025a <=( (not A299)  and  A298 );
 a42028a <=( A301  and  A300 );
 a42029a <=( a42028a  and  a42025a );
 a42030a <=( a42029a  and  a42022a );
 a42034a <=( (not A200)  and  A167 );
 a42035a <=( A168  and  a42034a );
 a42039a <=( A232  and  (not A203) );
 a42040a <=( (not A202)  and  a42039a );
 a42041a <=( a42040a  and  a42035a );
 a42045a <=( A235  and  A234 );
 a42046a <=( (not A233)  and  a42045a );
 a42049a <=( (not A299)  and  A298 );
 a42052a <=( A302  and  A300 );
 a42053a <=( a42052a  and  a42049a );
 a42054a <=( a42053a  and  a42046a );
 a42058a <=( (not A200)  and  A167 );
 a42059a <=( A168  and  a42058a );
 a42063a <=( A232  and  (not A203) );
 a42064a <=( (not A202)  and  a42063a );
 a42065a <=( a42064a  and  a42059a );
 a42069a <=( A235  and  A234 );
 a42070a <=( (not A233)  and  a42069a );
 a42073a <=( (not A266)  and  A265 );
 a42076a <=( A268  and  A267 );
 a42077a <=( a42076a  and  a42073a );
 a42078a <=( a42077a  and  a42070a );
 a42082a <=( (not A200)  and  A167 );
 a42083a <=( A168  and  a42082a );
 a42087a <=( A232  and  (not A203) );
 a42088a <=( (not A202)  and  a42087a );
 a42089a <=( a42088a  and  a42083a );
 a42093a <=( A235  and  A234 );
 a42094a <=( (not A233)  and  a42093a );
 a42097a <=( (not A266)  and  A265 );
 a42100a <=( A269  and  A267 );
 a42101a <=( a42100a  and  a42097a );
 a42102a <=( a42101a  and  a42094a );
 a42106a <=( (not A200)  and  A167 );
 a42107a <=( A168  and  a42106a );
 a42111a <=( A232  and  (not A203) );
 a42112a <=( (not A202)  and  a42111a );
 a42113a <=( a42112a  and  a42107a );
 a42117a <=( A236  and  A234 );
 a42118a <=( (not A233)  and  a42117a );
 a42121a <=( (not A299)  and  A298 );
 a42124a <=( A301  and  A300 );
 a42125a <=( a42124a  and  a42121a );
 a42126a <=( a42125a  and  a42118a );
 a42130a <=( (not A200)  and  A167 );
 a42131a <=( A168  and  a42130a );
 a42135a <=( A232  and  (not A203) );
 a42136a <=( (not A202)  and  a42135a );
 a42137a <=( a42136a  and  a42131a );
 a42141a <=( A236  and  A234 );
 a42142a <=( (not A233)  and  a42141a );
 a42145a <=( (not A299)  and  A298 );
 a42148a <=( A302  and  A300 );
 a42149a <=( a42148a  and  a42145a );
 a42150a <=( a42149a  and  a42142a );
 a42154a <=( (not A200)  and  A167 );
 a42155a <=( A168  and  a42154a );
 a42159a <=( A232  and  (not A203) );
 a42160a <=( (not A202)  and  a42159a );
 a42161a <=( a42160a  and  a42155a );
 a42165a <=( A236  and  A234 );
 a42166a <=( (not A233)  and  a42165a );
 a42169a <=( (not A266)  and  A265 );
 a42172a <=( A268  and  A267 );
 a42173a <=( a42172a  and  a42169a );
 a42174a <=( a42173a  and  a42166a );
 a42178a <=( (not A200)  and  A167 );
 a42179a <=( A168  and  a42178a );
 a42183a <=( A232  and  (not A203) );
 a42184a <=( (not A202)  and  a42183a );
 a42185a <=( a42184a  and  a42179a );
 a42189a <=( A236  and  A234 );
 a42190a <=( (not A233)  and  a42189a );
 a42193a <=( (not A266)  and  A265 );
 a42196a <=( A269  and  A267 );
 a42197a <=( a42196a  and  a42193a );
 a42198a <=( a42197a  and  a42190a );
 a42202a <=( (not A200)  and  A167 );
 a42203a <=( A168  and  a42202a );
 a42207a <=( (not A232)  and  (not A203) );
 a42208a <=( (not A202)  and  a42207a );
 a42209a <=( a42208a  and  a42203a );
 a42213a <=( (not A268)  and  (not A266) );
 a42214a <=( (not A233)  and  a42213a );
 a42217a <=( A298  and  (not A269) );
 a42220a <=( (not A302)  and  (not A301) );
 a42221a <=( a42220a  and  a42217a );
 a42222a <=( a42221a  and  a42214a );
 a42226a <=( (not A200)  and  A167 );
 a42227a <=( A168  and  a42226a );
 a42231a <=( (not A235)  and  (not A233) );
 a42232a <=( (not A201)  and  a42231a );
 a42233a <=( a42232a  and  a42227a );
 a42237a <=( (not A268)  and  (not A266) );
 a42238a <=( (not A236)  and  a42237a );
 a42241a <=( A298  and  (not A269) );
 a42244a <=( (not A302)  and  (not A301) );
 a42245a <=( a42244a  and  a42241a );
 a42246a <=( a42245a  and  a42238a );
 a42250a <=( (not A199)  and  A167 );
 a42251a <=( A168  and  a42250a );
 a42255a <=( (not A235)  and  (not A233) );
 a42256a <=( (not A200)  and  a42255a );
 a42257a <=( a42256a  and  a42251a );
 a42261a <=( (not A268)  and  (not A266) );
 a42262a <=( (not A236)  and  a42261a );
 a42265a <=( A298  and  (not A269) );
 a42268a <=( (not A302)  and  (not A301) );
 a42269a <=( a42268a  and  a42265a );
 a42270a <=( a42269a  and  a42262a );
 a42274a <=( (not A166)  and  (not A167) );
 a42275a <=( A170  and  a42274a );
 a42279a <=( A232  and  A200 );
 a42280a <=( (not A199)  and  a42279a );
 a42281a <=( a42280a  and  a42275a );
 a42285a <=( (not A268)  and  A265 );
 a42286a <=( A233  and  a42285a );
 a42289a <=( (not A299)  and  (not A269) );
 a42292a <=( (not A302)  and  (not A301) );
 a42293a <=( a42292a  and  a42289a );
 a42294a <=( a42293a  and  a42286a );
 a42298a <=( (not A166)  and  (not A167) );
 a42299a <=( A170  and  a42298a );
 a42303a <=( (not A233)  and  A200 );
 a42304a <=( (not A199)  and  a42303a );
 a42305a <=( a42304a  and  a42299a );
 a42309a <=( A265  and  (not A236) );
 a42310a <=( (not A235)  and  a42309a );
 a42313a <=( A298  and  A266 );
 a42316a <=( (not A302)  and  (not A301) );
 a42317a <=( a42316a  and  a42313a );
 a42318a <=( a42317a  and  a42310a );
 a42322a <=( (not A166)  and  (not A167) );
 a42323a <=( A170  and  a42322a );
 a42327a <=( (not A233)  and  A200 );
 a42328a <=( (not A199)  and  a42327a );
 a42329a <=( a42328a  and  a42323a );
 a42333a <=( (not A266)  and  (not A236) );
 a42334a <=( (not A235)  and  a42333a );
 a42337a <=( (not A269)  and  (not A268) );
 a42340a <=( (not A300)  and  A298 );
 a42341a <=( a42340a  and  a42337a );
 a42342a <=( a42341a  and  a42334a );
 a42346a <=( (not A166)  and  (not A167) );
 a42347a <=( A170  and  a42346a );
 a42351a <=( (not A233)  and  A200 );
 a42352a <=( (not A199)  and  a42351a );
 a42353a <=( a42352a  and  a42347a );
 a42357a <=( (not A266)  and  (not A236) );
 a42358a <=( (not A235)  and  a42357a );
 a42361a <=( (not A269)  and  (not A268) );
 a42364a <=( A299  and  A298 );
 a42365a <=( a42364a  and  a42361a );
 a42366a <=( a42365a  and  a42358a );
 a42370a <=( (not A166)  and  (not A167) );
 a42371a <=( A170  and  a42370a );
 a42375a <=( (not A233)  and  A200 );
 a42376a <=( (not A199)  and  a42375a );
 a42377a <=( a42376a  and  a42371a );
 a42381a <=( (not A266)  and  (not A236) );
 a42382a <=( (not A235)  and  a42381a );
 a42385a <=( (not A269)  and  (not A268) );
 a42388a <=( (not A299)  and  (not A298) );
 a42389a <=( a42388a  and  a42385a );
 a42390a <=( a42389a  and  a42382a );
 a42394a <=( (not A166)  and  (not A167) );
 a42395a <=( A170  and  a42394a );
 a42399a <=( (not A233)  and  A200 );
 a42400a <=( (not A199)  and  a42399a );
 a42401a <=( a42400a  and  a42395a );
 a42405a <=( (not A266)  and  (not A236) );
 a42406a <=( (not A235)  and  a42405a );
 a42409a <=( A298  and  (not A267) );
 a42412a <=( (not A302)  and  (not A301) );
 a42413a <=( a42412a  and  a42409a );
 a42414a <=( a42413a  and  a42406a );
 a42418a <=( (not A166)  and  (not A167) );
 a42419a <=( A170  and  a42418a );
 a42423a <=( (not A233)  and  A200 );
 a42424a <=( (not A199)  and  a42423a );
 a42425a <=( a42424a  and  a42419a );
 a42429a <=( (not A265)  and  (not A236) );
 a42430a <=( (not A235)  and  a42429a );
 a42433a <=( A298  and  (not A266) );
 a42436a <=( (not A302)  and  (not A301) );
 a42437a <=( a42436a  and  a42433a );
 a42438a <=( a42437a  and  a42430a );
 a42442a <=( (not A166)  and  (not A167) );
 a42443a <=( A170  and  a42442a );
 a42447a <=( (not A233)  and  A200 );
 a42448a <=( (not A199)  and  a42447a );
 a42449a <=( a42448a  and  a42443a );
 a42453a <=( (not A268)  and  (not A266) );
 a42454a <=( (not A234)  and  a42453a );
 a42457a <=( A298  and  (not A269) );
 a42460a <=( (not A302)  and  (not A301) );
 a42461a <=( a42460a  and  a42457a );
 a42462a <=( a42461a  and  a42454a );
 a42466a <=( (not A166)  and  (not A167) );
 a42467a <=( A170  and  a42466a );
 a42471a <=( A232  and  A200 );
 a42472a <=( (not A199)  and  a42471a );
 a42473a <=( a42472a  and  a42467a );
 a42477a <=( A235  and  A234 );
 a42478a <=( (not A233)  and  a42477a );
 a42481a <=( (not A299)  and  A298 );
 a42484a <=( A301  and  A300 );
 a42485a <=( a42484a  and  a42481a );
 a42486a <=( a42485a  and  a42478a );
 a42490a <=( (not A166)  and  (not A167) );
 a42491a <=( A170  and  a42490a );
 a42495a <=( A232  and  A200 );
 a42496a <=( (not A199)  and  a42495a );
 a42497a <=( a42496a  and  a42491a );
 a42501a <=( A235  and  A234 );
 a42502a <=( (not A233)  and  a42501a );
 a42505a <=( (not A299)  and  A298 );
 a42508a <=( A302  and  A300 );
 a42509a <=( a42508a  and  a42505a );
 a42510a <=( a42509a  and  a42502a );
 a42514a <=( (not A166)  and  (not A167) );
 a42515a <=( A170  and  a42514a );
 a42519a <=( A232  and  A200 );
 a42520a <=( (not A199)  and  a42519a );
 a42521a <=( a42520a  and  a42515a );
 a42525a <=( A235  and  A234 );
 a42526a <=( (not A233)  and  a42525a );
 a42529a <=( (not A266)  and  A265 );
 a42532a <=( A268  and  A267 );
 a42533a <=( a42532a  and  a42529a );
 a42534a <=( a42533a  and  a42526a );
 a42538a <=( (not A166)  and  (not A167) );
 a42539a <=( A170  and  a42538a );
 a42543a <=( A232  and  A200 );
 a42544a <=( (not A199)  and  a42543a );
 a42545a <=( a42544a  and  a42539a );
 a42549a <=( A235  and  A234 );
 a42550a <=( (not A233)  and  a42549a );
 a42553a <=( (not A266)  and  A265 );
 a42556a <=( A269  and  A267 );
 a42557a <=( a42556a  and  a42553a );
 a42558a <=( a42557a  and  a42550a );
 a42562a <=( (not A166)  and  (not A167) );
 a42563a <=( A170  and  a42562a );
 a42567a <=( A232  and  A200 );
 a42568a <=( (not A199)  and  a42567a );
 a42569a <=( a42568a  and  a42563a );
 a42573a <=( A236  and  A234 );
 a42574a <=( (not A233)  and  a42573a );
 a42577a <=( (not A299)  and  A298 );
 a42580a <=( A301  and  A300 );
 a42581a <=( a42580a  and  a42577a );
 a42582a <=( a42581a  and  a42574a );
 a42586a <=( (not A166)  and  (not A167) );
 a42587a <=( A170  and  a42586a );
 a42591a <=( A232  and  A200 );
 a42592a <=( (not A199)  and  a42591a );
 a42593a <=( a42592a  and  a42587a );
 a42597a <=( A236  and  A234 );
 a42598a <=( (not A233)  and  a42597a );
 a42601a <=( (not A299)  and  A298 );
 a42604a <=( A302  and  A300 );
 a42605a <=( a42604a  and  a42601a );
 a42606a <=( a42605a  and  a42598a );
 a42610a <=( (not A166)  and  (not A167) );
 a42611a <=( A170  and  a42610a );
 a42615a <=( A232  and  A200 );
 a42616a <=( (not A199)  and  a42615a );
 a42617a <=( a42616a  and  a42611a );
 a42621a <=( A236  and  A234 );
 a42622a <=( (not A233)  and  a42621a );
 a42625a <=( (not A266)  and  A265 );
 a42628a <=( A268  and  A267 );
 a42629a <=( a42628a  and  a42625a );
 a42630a <=( a42629a  and  a42622a );
 a42634a <=( (not A166)  and  (not A167) );
 a42635a <=( A170  and  a42634a );
 a42639a <=( A232  and  A200 );
 a42640a <=( (not A199)  and  a42639a );
 a42641a <=( a42640a  and  a42635a );
 a42645a <=( A236  and  A234 );
 a42646a <=( (not A233)  and  a42645a );
 a42649a <=( (not A266)  and  A265 );
 a42652a <=( A269  and  A267 );
 a42653a <=( a42652a  and  a42649a );
 a42654a <=( a42653a  and  a42646a );
 a42658a <=( (not A166)  and  (not A167) );
 a42659a <=( A170  and  a42658a );
 a42663a <=( (not A232)  and  A200 );
 a42664a <=( (not A199)  and  a42663a );
 a42665a <=( a42664a  and  a42659a );
 a42669a <=( (not A268)  and  (not A266) );
 a42670a <=( (not A233)  and  a42669a );
 a42673a <=( A298  and  (not A269) );
 a42676a <=( (not A302)  and  (not A301) );
 a42677a <=( a42676a  and  a42673a );
 a42678a <=( a42677a  and  a42670a );
 a42682a <=( (not A166)  and  (not A167) );
 a42683a <=( A170  and  a42682a );
 a42687a <=( A201  and  (not A200) );
 a42688a <=( A199  and  a42687a );
 a42689a <=( a42688a  and  a42683a );
 a42693a <=( A233  and  A232 );
 a42694a <=( A202  and  a42693a );
 a42697a <=( (not A267)  and  A265 );
 a42700a <=( (not A300)  and  (not A299) );
 a42701a <=( a42700a  and  a42697a );
 a42702a <=( a42701a  and  a42694a );
 a42706a <=( (not A166)  and  (not A167) );
 a42707a <=( A170  and  a42706a );
 a42711a <=( A201  and  (not A200) );
 a42712a <=( A199  and  a42711a );
 a42713a <=( a42712a  and  a42707a );
 a42717a <=( A233  and  A232 );
 a42718a <=( A202  and  a42717a );
 a42721a <=( (not A267)  and  A265 );
 a42724a <=( A299  and  A298 );
 a42725a <=( a42724a  and  a42721a );
 a42726a <=( a42725a  and  a42718a );
 a42730a <=( (not A166)  and  (not A167) );
 a42731a <=( A170  and  a42730a );
 a42735a <=( A201  and  (not A200) );
 a42736a <=( A199  and  a42735a );
 a42737a <=( a42736a  and  a42731a );
 a42741a <=( A233  and  A232 );
 a42742a <=( A202  and  a42741a );
 a42745a <=( (not A267)  and  A265 );
 a42748a <=( (not A299)  and  (not A298) );
 a42749a <=( a42748a  and  a42745a );
 a42750a <=( a42749a  and  a42742a );
 a42754a <=( (not A166)  and  (not A167) );
 a42755a <=( A170  and  a42754a );
 a42759a <=( A201  and  (not A200) );
 a42760a <=( A199  and  a42759a );
 a42761a <=( a42760a  and  a42755a );
 a42765a <=( A233  and  A232 );
 a42766a <=( A202  and  a42765a );
 a42769a <=( A266  and  A265 );
 a42772a <=( (not A300)  and  (not A299) );
 a42773a <=( a42772a  and  a42769a );
 a42774a <=( a42773a  and  a42766a );
 a42778a <=( (not A166)  and  (not A167) );
 a42779a <=( A170  and  a42778a );
 a42783a <=( A201  and  (not A200) );
 a42784a <=( A199  and  a42783a );
 a42785a <=( a42784a  and  a42779a );
 a42789a <=( A233  and  A232 );
 a42790a <=( A202  and  a42789a );
 a42793a <=( A266  and  A265 );
 a42796a <=( A299  and  A298 );
 a42797a <=( a42796a  and  a42793a );
 a42798a <=( a42797a  and  a42790a );
 a42802a <=( (not A166)  and  (not A167) );
 a42803a <=( A170  and  a42802a );
 a42807a <=( A201  and  (not A200) );
 a42808a <=( A199  and  a42807a );
 a42809a <=( a42808a  and  a42803a );
 a42813a <=( A233  and  A232 );
 a42814a <=( A202  and  a42813a );
 a42817a <=( A266  and  A265 );
 a42820a <=( (not A299)  and  (not A298) );
 a42821a <=( a42820a  and  a42817a );
 a42822a <=( a42821a  and  a42814a );
 a42826a <=( (not A166)  and  (not A167) );
 a42827a <=( A170  and  a42826a );
 a42831a <=( A201  and  (not A200) );
 a42832a <=( A199  and  a42831a );
 a42833a <=( a42832a  and  a42827a );
 a42837a <=( A233  and  A232 );
 a42838a <=( A202  and  a42837a );
 a42841a <=( (not A266)  and  (not A265) );
 a42844a <=( (not A300)  and  (not A299) );
 a42845a <=( a42844a  and  a42841a );
 a42846a <=( a42845a  and  a42838a );
 a42850a <=( (not A166)  and  (not A167) );
 a42851a <=( A170  and  a42850a );
 a42855a <=( A201  and  (not A200) );
 a42856a <=( A199  and  a42855a );
 a42857a <=( a42856a  and  a42851a );
 a42861a <=( A233  and  A232 );
 a42862a <=( A202  and  a42861a );
 a42865a <=( (not A266)  and  (not A265) );
 a42868a <=( A299  and  A298 );
 a42869a <=( a42868a  and  a42865a );
 a42870a <=( a42869a  and  a42862a );
 a42874a <=( (not A166)  and  (not A167) );
 a42875a <=( A170  and  a42874a );
 a42879a <=( A201  and  (not A200) );
 a42880a <=( A199  and  a42879a );
 a42881a <=( a42880a  and  a42875a );
 a42885a <=( A233  and  A232 );
 a42886a <=( A202  and  a42885a );
 a42889a <=( (not A266)  and  (not A265) );
 a42892a <=( (not A299)  and  (not A298) );
 a42893a <=( a42892a  and  a42889a );
 a42894a <=( a42893a  and  a42886a );
 a42898a <=( (not A166)  and  (not A167) );
 a42899a <=( A170  and  a42898a );
 a42903a <=( A201  and  (not A200) );
 a42904a <=( A199  and  a42903a );
 a42905a <=( a42904a  and  a42899a );
 a42909a <=( A233  and  (not A232) );
 a42910a <=( A202  and  a42909a );
 a42913a <=( (not A299)  and  A298 );
 a42916a <=( A301  and  A300 );
 a42917a <=( a42916a  and  a42913a );
 a42918a <=( a42917a  and  a42910a );
 a42922a <=( (not A166)  and  (not A167) );
 a42923a <=( A170  and  a42922a );
 a42927a <=( A201  and  (not A200) );
 a42928a <=( A199  and  a42927a );
 a42929a <=( a42928a  and  a42923a );
 a42933a <=( A233  and  (not A232) );
 a42934a <=( A202  and  a42933a );
 a42937a <=( (not A299)  and  A298 );
 a42940a <=( A302  and  A300 );
 a42941a <=( a42940a  and  a42937a );
 a42942a <=( a42941a  and  a42934a );
 a42946a <=( (not A166)  and  (not A167) );
 a42947a <=( A170  and  a42946a );
 a42951a <=( A201  and  (not A200) );
 a42952a <=( A199  and  a42951a );
 a42953a <=( a42952a  and  a42947a );
 a42957a <=( A233  and  (not A232) );
 a42958a <=( A202  and  a42957a );
 a42961a <=( (not A266)  and  A265 );
 a42964a <=( A268  and  A267 );
 a42965a <=( a42964a  and  a42961a );
 a42966a <=( a42965a  and  a42958a );
 a42970a <=( (not A166)  and  (not A167) );
 a42971a <=( A170  and  a42970a );
 a42975a <=( A201  and  (not A200) );
 a42976a <=( A199  and  a42975a );
 a42977a <=( a42976a  and  a42971a );
 a42981a <=( A233  and  (not A232) );
 a42982a <=( A202  and  a42981a );
 a42985a <=( (not A266)  and  A265 );
 a42988a <=( A269  and  A267 );
 a42989a <=( a42988a  and  a42985a );
 a42990a <=( a42989a  and  a42982a );
 a42994a <=( (not A166)  and  (not A167) );
 a42995a <=( A170  and  a42994a );
 a42999a <=( A201  and  (not A200) );
 a43000a <=( A199  and  a42999a );
 a43001a <=( a43000a  and  a42995a );
 a43005a <=( (not A234)  and  (not A233) );
 a43006a <=( A202  and  a43005a );
 a43009a <=( A266  and  A265 );
 a43012a <=( (not A300)  and  A298 );
 a43013a <=( a43012a  and  a43009a );
 a43014a <=( a43013a  and  a43006a );
 a43018a <=( (not A166)  and  (not A167) );
 a43019a <=( A170  and  a43018a );
 a43023a <=( A201  and  (not A200) );
 a43024a <=( A199  and  a43023a );
 a43025a <=( a43024a  and  a43019a );
 a43029a <=( (not A234)  and  (not A233) );
 a43030a <=( A202  and  a43029a );
 a43033a <=( A266  and  A265 );
 a43036a <=( A299  and  A298 );
 a43037a <=( a43036a  and  a43033a );
 a43038a <=( a43037a  and  a43030a );
 a43042a <=( (not A166)  and  (not A167) );
 a43043a <=( A170  and  a43042a );
 a43047a <=( A201  and  (not A200) );
 a43048a <=( A199  and  a43047a );
 a43049a <=( a43048a  and  a43043a );
 a43053a <=( (not A234)  and  (not A233) );
 a43054a <=( A202  and  a43053a );
 a43057a <=( A266  and  A265 );
 a43060a <=( (not A299)  and  (not A298) );
 a43061a <=( a43060a  and  a43057a );
 a43062a <=( a43061a  and  a43054a );
 a43066a <=( (not A166)  and  (not A167) );
 a43067a <=( A170  and  a43066a );
 a43071a <=( A201  and  (not A200) );
 a43072a <=( A199  and  a43071a );
 a43073a <=( a43072a  and  a43067a );
 a43077a <=( (not A234)  and  (not A233) );
 a43078a <=( A202  and  a43077a );
 a43081a <=( (not A267)  and  (not A266) );
 a43084a <=( (not A300)  and  A298 );
 a43085a <=( a43084a  and  a43081a );
 a43086a <=( a43085a  and  a43078a );
 a43090a <=( (not A166)  and  (not A167) );
 a43091a <=( A170  and  a43090a );
 a43095a <=( A201  and  (not A200) );
 a43096a <=( A199  and  a43095a );
 a43097a <=( a43096a  and  a43091a );
 a43101a <=( (not A234)  and  (not A233) );
 a43102a <=( A202  and  a43101a );
 a43105a <=( (not A267)  and  (not A266) );
 a43108a <=( A299  and  A298 );
 a43109a <=( a43108a  and  a43105a );
 a43110a <=( a43109a  and  a43102a );
 a43114a <=( (not A166)  and  (not A167) );
 a43115a <=( A170  and  a43114a );
 a43119a <=( A201  and  (not A200) );
 a43120a <=( A199  and  a43119a );
 a43121a <=( a43120a  and  a43115a );
 a43125a <=( (not A234)  and  (not A233) );
 a43126a <=( A202  and  a43125a );
 a43129a <=( (not A267)  and  (not A266) );
 a43132a <=( (not A299)  and  (not A298) );
 a43133a <=( a43132a  and  a43129a );
 a43134a <=( a43133a  and  a43126a );
 a43138a <=( (not A166)  and  (not A167) );
 a43139a <=( A170  and  a43138a );
 a43143a <=( A201  and  (not A200) );
 a43144a <=( A199  and  a43143a );
 a43145a <=( a43144a  and  a43139a );
 a43149a <=( (not A234)  and  (not A233) );
 a43150a <=( A202  and  a43149a );
 a43153a <=( (not A266)  and  (not A265) );
 a43156a <=( (not A300)  and  A298 );
 a43157a <=( a43156a  and  a43153a );
 a43158a <=( a43157a  and  a43150a );
 a43162a <=( (not A166)  and  (not A167) );
 a43163a <=( A170  and  a43162a );
 a43167a <=( A201  and  (not A200) );
 a43168a <=( A199  and  a43167a );
 a43169a <=( a43168a  and  a43163a );
 a43173a <=( (not A234)  and  (not A233) );
 a43174a <=( A202  and  a43173a );
 a43177a <=( (not A266)  and  (not A265) );
 a43180a <=( A299  and  A298 );
 a43181a <=( a43180a  and  a43177a );
 a43182a <=( a43181a  and  a43174a );
 a43186a <=( (not A166)  and  (not A167) );
 a43187a <=( A170  and  a43186a );
 a43191a <=( A201  and  (not A200) );
 a43192a <=( A199  and  a43191a );
 a43193a <=( a43192a  and  a43187a );
 a43197a <=( (not A234)  and  (not A233) );
 a43198a <=( A202  and  a43197a );
 a43201a <=( (not A266)  and  (not A265) );
 a43204a <=( (not A299)  and  (not A298) );
 a43205a <=( a43204a  and  a43201a );
 a43206a <=( a43205a  and  a43198a );
 a43210a <=( (not A166)  and  (not A167) );
 a43211a <=( A170  and  a43210a );
 a43215a <=( A201  and  (not A200) );
 a43216a <=( A199  and  a43215a );
 a43217a <=( a43216a  and  a43211a );
 a43221a <=( (not A233)  and  A232 );
 a43222a <=( A202  and  a43221a );
 a43225a <=( A235  and  A234 );
 a43228a <=( A299  and  (not A298) );
 a43229a <=( a43228a  and  a43225a );
 a43230a <=( a43229a  and  a43222a );
 a43234a <=( (not A166)  and  (not A167) );
 a43235a <=( A170  and  a43234a );
 a43239a <=( A201  and  (not A200) );
 a43240a <=( A199  and  a43239a );
 a43241a <=( a43240a  and  a43235a );
 a43245a <=( (not A233)  and  A232 );
 a43246a <=( A202  and  a43245a );
 a43249a <=( A235  and  A234 );
 a43252a <=( A266  and  (not A265) );
 a43253a <=( a43252a  and  a43249a );
 a43254a <=( a43253a  and  a43246a );
 a43258a <=( (not A166)  and  (not A167) );
 a43259a <=( A170  and  a43258a );
 a43263a <=( A201  and  (not A200) );
 a43264a <=( A199  and  a43263a );
 a43265a <=( a43264a  and  a43259a );
 a43269a <=( (not A233)  and  A232 );
 a43270a <=( A202  and  a43269a );
 a43273a <=( A236  and  A234 );
 a43276a <=( A299  and  (not A298) );
 a43277a <=( a43276a  and  a43273a );
 a43278a <=( a43277a  and  a43270a );
 a43282a <=( (not A166)  and  (not A167) );
 a43283a <=( A170  and  a43282a );
 a43287a <=( A201  and  (not A200) );
 a43288a <=( A199  and  a43287a );
 a43289a <=( a43288a  and  a43283a );
 a43293a <=( (not A233)  and  A232 );
 a43294a <=( A202  and  a43293a );
 a43297a <=( A236  and  A234 );
 a43300a <=( A266  and  (not A265) );
 a43301a <=( a43300a  and  a43297a );
 a43302a <=( a43301a  and  a43294a );
 a43306a <=( (not A166)  and  (not A167) );
 a43307a <=( A170  and  a43306a );
 a43311a <=( A201  and  (not A200) );
 a43312a <=( A199  and  a43311a );
 a43313a <=( a43312a  and  a43307a );
 a43317a <=( (not A233)  and  (not A232) );
 a43318a <=( A202  and  a43317a );
 a43321a <=( A266  and  A265 );
 a43324a <=( (not A300)  and  A298 );
 a43325a <=( a43324a  and  a43321a );
 a43326a <=( a43325a  and  a43318a );
 a43330a <=( (not A166)  and  (not A167) );
 a43331a <=( A170  and  a43330a );
 a43335a <=( A201  and  (not A200) );
 a43336a <=( A199  and  a43335a );
 a43337a <=( a43336a  and  a43331a );
 a43341a <=( (not A233)  and  (not A232) );
 a43342a <=( A202  and  a43341a );
 a43345a <=( A266  and  A265 );
 a43348a <=( A299  and  A298 );
 a43349a <=( a43348a  and  a43345a );
 a43350a <=( a43349a  and  a43342a );
 a43354a <=( (not A166)  and  (not A167) );
 a43355a <=( A170  and  a43354a );
 a43359a <=( A201  and  (not A200) );
 a43360a <=( A199  and  a43359a );
 a43361a <=( a43360a  and  a43355a );
 a43365a <=( (not A233)  and  (not A232) );
 a43366a <=( A202  and  a43365a );
 a43369a <=( A266  and  A265 );
 a43372a <=( (not A299)  and  (not A298) );
 a43373a <=( a43372a  and  a43369a );
 a43374a <=( a43373a  and  a43366a );
 a43378a <=( (not A166)  and  (not A167) );
 a43379a <=( A170  and  a43378a );
 a43383a <=( A201  and  (not A200) );
 a43384a <=( A199  and  a43383a );
 a43385a <=( a43384a  and  a43379a );
 a43389a <=( (not A233)  and  (not A232) );
 a43390a <=( A202  and  a43389a );
 a43393a <=( (not A267)  and  (not A266) );
 a43396a <=( (not A300)  and  A298 );
 a43397a <=( a43396a  and  a43393a );
 a43398a <=( a43397a  and  a43390a );
 a43402a <=( (not A166)  and  (not A167) );
 a43403a <=( A170  and  a43402a );
 a43407a <=( A201  and  (not A200) );
 a43408a <=( A199  and  a43407a );
 a43409a <=( a43408a  and  a43403a );
 a43413a <=( (not A233)  and  (not A232) );
 a43414a <=( A202  and  a43413a );
 a43417a <=( (not A267)  and  (not A266) );
 a43420a <=( A299  and  A298 );
 a43421a <=( a43420a  and  a43417a );
 a43422a <=( a43421a  and  a43414a );
 a43426a <=( (not A166)  and  (not A167) );
 a43427a <=( A170  and  a43426a );
 a43431a <=( A201  and  (not A200) );
 a43432a <=( A199  and  a43431a );
 a43433a <=( a43432a  and  a43427a );
 a43437a <=( (not A233)  and  (not A232) );
 a43438a <=( A202  and  a43437a );
 a43441a <=( (not A267)  and  (not A266) );
 a43444a <=( (not A299)  and  (not A298) );
 a43445a <=( a43444a  and  a43441a );
 a43446a <=( a43445a  and  a43438a );
 a43450a <=( (not A166)  and  (not A167) );
 a43451a <=( A170  and  a43450a );
 a43455a <=( A201  and  (not A200) );
 a43456a <=( A199  and  a43455a );
 a43457a <=( a43456a  and  a43451a );
 a43461a <=( (not A233)  and  (not A232) );
 a43462a <=( A202  and  a43461a );
 a43465a <=( (not A266)  and  (not A265) );
 a43468a <=( (not A300)  and  A298 );
 a43469a <=( a43468a  and  a43465a );
 a43470a <=( a43469a  and  a43462a );
 a43474a <=( (not A166)  and  (not A167) );
 a43475a <=( A170  and  a43474a );
 a43479a <=( A201  and  (not A200) );
 a43480a <=( A199  and  a43479a );
 a43481a <=( a43480a  and  a43475a );
 a43485a <=( (not A233)  and  (not A232) );
 a43486a <=( A202  and  a43485a );
 a43489a <=( (not A266)  and  (not A265) );
 a43492a <=( A299  and  A298 );
 a43493a <=( a43492a  and  a43489a );
 a43494a <=( a43493a  and  a43486a );
 a43498a <=( (not A166)  and  (not A167) );
 a43499a <=( A170  and  a43498a );
 a43503a <=( A201  and  (not A200) );
 a43504a <=( A199  and  a43503a );
 a43505a <=( a43504a  and  a43499a );
 a43509a <=( (not A233)  and  (not A232) );
 a43510a <=( A202  and  a43509a );
 a43513a <=( (not A266)  and  (not A265) );
 a43516a <=( (not A299)  and  (not A298) );
 a43517a <=( a43516a  and  a43513a );
 a43518a <=( a43517a  and  a43510a );
 a43522a <=( (not A166)  and  (not A167) );
 a43523a <=( A170  and  a43522a );
 a43527a <=( A201  and  (not A200) );
 a43528a <=( A199  and  a43527a );
 a43529a <=( a43528a  and  a43523a );
 a43533a <=( A233  and  A232 );
 a43534a <=( A203  and  a43533a );
 a43537a <=( (not A267)  and  A265 );
 a43540a <=( (not A300)  and  (not A299) );
 a43541a <=( a43540a  and  a43537a );
 a43542a <=( a43541a  and  a43534a );
 a43546a <=( (not A166)  and  (not A167) );
 a43547a <=( A170  and  a43546a );
 a43551a <=( A201  and  (not A200) );
 a43552a <=( A199  and  a43551a );
 a43553a <=( a43552a  and  a43547a );
 a43557a <=( A233  and  A232 );
 a43558a <=( A203  and  a43557a );
 a43561a <=( (not A267)  and  A265 );
 a43564a <=( A299  and  A298 );
 a43565a <=( a43564a  and  a43561a );
 a43566a <=( a43565a  and  a43558a );
 a43570a <=( (not A166)  and  (not A167) );
 a43571a <=( A170  and  a43570a );
 a43575a <=( A201  and  (not A200) );
 a43576a <=( A199  and  a43575a );
 a43577a <=( a43576a  and  a43571a );
 a43581a <=( A233  and  A232 );
 a43582a <=( A203  and  a43581a );
 a43585a <=( (not A267)  and  A265 );
 a43588a <=( (not A299)  and  (not A298) );
 a43589a <=( a43588a  and  a43585a );
 a43590a <=( a43589a  and  a43582a );
 a43594a <=( (not A166)  and  (not A167) );
 a43595a <=( A170  and  a43594a );
 a43599a <=( A201  and  (not A200) );
 a43600a <=( A199  and  a43599a );
 a43601a <=( a43600a  and  a43595a );
 a43605a <=( A233  and  A232 );
 a43606a <=( A203  and  a43605a );
 a43609a <=( A266  and  A265 );
 a43612a <=( (not A300)  and  (not A299) );
 a43613a <=( a43612a  and  a43609a );
 a43614a <=( a43613a  and  a43606a );
 a43618a <=( (not A166)  and  (not A167) );
 a43619a <=( A170  and  a43618a );
 a43623a <=( A201  and  (not A200) );
 a43624a <=( A199  and  a43623a );
 a43625a <=( a43624a  and  a43619a );
 a43629a <=( A233  and  A232 );
 a43630a <=( A203  and  a43629a );
 a43633a <=( A266  and  A265 );
 a43636a <=( A299  and  A298 );
 a43637a <=( a43636a  and  a43633a );
 a43638a <=( a43637a  and  a43630a );
 a43642a <=( (not A166)  and  (not A167) );
 a43643a <=( A170  and  a43642a );
 a43647a <=( A201  and  (not A200) );
 a43648a <=( A199  and  a43647a );
 a43649a <=( a43648a  and  a43643a );
 a43653a <=( A233  and  A232 );
 a43654a <=( A203  and  a43653a );
 a43657a <=( A266  and  A265 );
 a43660a <=( (not A299)  and  (not A298) );
 a43661a <=( a43660a  and  a43657a );
 a43662a <=( a43661a  and  a43654a );
 a43666a <=( (not A166)  and  (not A167) );
 a43667a <=( A170  and  a43666a );
 a43671a <=( A201  and  (not A200) );
 a43672a <=( A199  and  a43671a );
 a43673a <=( a43672a  and  a43667a );
 a43677a <=( A233  and  A232 );
 a43678a <=( A203  and  a43677a );
 a43681a <=( (not A266)  and  (not A265) );
 a43684a <=( (not A300)  and  (not A299) );
 a43685a <=( a43684a  and  a43681a );
 a43686a <=( a43685a  and  a43678a );
 a43690a <=( (not A166)  and  (not A167) );
 a43691a <=( A170  and  a43690a );
 a43695a <=( A201  and  (not A200) );
 a43696a <=( A199  and  a43695a );
 a43697a <=( a43696a  and  a43691a );
 a43701a <=( A233  and  A232 );
 a43702a <=( A203  and  a43701a );
 a43705a <=( (not A266)  and  (not A265) );
 a43708a <=( A299  and  A298 );
 a43709a <=( a43708a  and  a43705a );
 a43710a <=( a43709a  and  a43702a );
 a43714a <=( (not A166)  and  (not A167) );
 a43715a <=( A170  and  a43714a );
 a43719a <=( A201  and  (not A200) );
 a43720a <=( A199  and  a43719a );
 a43721a <=( a43720a  and  a43715a );
 a43725a <=( A233  and  A232 );
 a43726a <=( A203  and  a43725a );
 a43729a <=( (not A266)  and  (not A265) );
 a43732a <=( (not A299)  and  (not A298) );
 a43733a <=( a43732a  and  a43729a );
 a43734a <=( a43733a  and  a43726a );
 a43738a <=( (not A166)  and  (not A167) );
 a43739a <=( A170  and  a43738a );
 a43743a <=( A201  and  (not A200) );
 a43744a <=( A199  and  a43743a );
 a43745a <=( a43744a  and  a43739a );
 a43749a <=( A233  and  (not A232) );
 a43750a <=( A203  and  a43749a );
 a43753a <=( (not A299)  and  A298 );
 a43756a <=( A301  and  A300 );
 a43757a <=( a43756a  and  a43753a );
 a43758a <=( a43757a  and  a43750a );
 a43762a <=( (not A166)  and  (not A167) );
 a43763a <=( A170  and  a43762a );
 a43767a <=( A201  and  (not A200) );
 a43768a <=( A199  and  a43767a );
 a43769a <=( a43768a  and  a43763a );
 a43773a <=( A233  and  (not A232) );
 a43774a <=( A203  and  a43773a );
 a43777a <=( (not A299)  and  A298 );
 a43780a <=( A302  and  A300 );
 a43781a <=( a43780a  and  a43777a );
 a43782a <=( a43781a  and  a43774a );
 a43786a <=( (not A166)  and  (not A167) );
 a43787a <=( A170  and  a43786a );
 a43791a <=( A201  and  (not A200) );
 a43792a <=( A199  and  a43791a );
 a43793a <=( a43792a  and  a43787a );
 a43797a <=( A233  and  (not A232) );
 a43798a <=( A203  and  a43797a );
 a43801a <=( (not A266)  and  A265 );
 a43804a <=( A268  and  A267 );
 a43805a <=( a43804a  and  a43801a );
 a43806a <=( a43805a  and  a43798a );
 a43810a <=( (not A166)  and  (not A167) );
 a43811a <=( A170  and  a43810a );
 a43815a <=( A201  and  (not A200) );
 a43816a <=( A199  and  a43815a );
 a43817a <=( a43816a  and  a43811a );
 a43821a <=( A233  and  (not A232) );
 a43822a <=( A203  and  a43821a );
 a43825a <=( (not A266)  and  A265 );
 a43828a <=( A269  and  A267 );
 a43829a <=( a43828a  and  a43825a );
 a43830a <=( a43829a  and  a43822a );
 a43834a <=( (not A166)  and  (not A167) );
 a43835a <=( A170  and  a43834a );
 a43839a <=( A201  and  (not A200) );
 a43840a <=( A199  and  a43839a );
 a43841a <=( a43840a  and  a43835a );
 a43845a <=( (not A234)  and  (not A233) );
 a43846a <=( A203  and  a43845a );
 a43849a <=( A266  and  A265 );
 a43852a <=( (not A300)  and  A298 );
 a43853a <=( a43852a  and  a43849a );
 a43854a <=( a43853a  and  a43846a );
 a43858a <=( (not A166)  and  (not A167) );
 a43859a <=( A170  and  a43858a );
 a43863a <=( A201  and  (not A200) );
 a43864a <=( A199  and  a43863a );
 a43865a <=( a43864a  and  a43859a );
 a43869a <=( (not A234)  and  (not A233) );
 a43870a <=( A203  and  a43869a );
 a43873a <=( A266  and  A265 );
 a43876a <=( A299  and  A298 );
 a43877a <=( a43876a  and  a43873a );
 a43878a <=( a43877a  and  a43870a );
 a43882a <=( (not A166)  and  (not A167) );
 a43883a <=( A170  and  a43882a );
 a43887a <=( A201  and  (not A200) );
 a43888a <=( A199  and  a43887a );
 a43889a <=( a43888a  and  a43883a );
 a43893a <=( (not A234)  and  (not A233) );
 a43894a <=( A203  and  a43893a );
 a43897a <=( A266  and  A265 );
 a43900a <=( (not A299)  and  (not A298) );
 a43901a <=( a43900a  and  a43897a );
 a43902a <=( a43901a  and  a43894a );
 a43906a <=( (not A166)  and  (not A167) );
 a43907a <=( A170  and  a43906a );
 a43911a <=( A201  and  (not A200) );
 a43912a <=( A199  and  a43911a );
 a43913a <=( a43912a  and  a43907a );
 a43917a <=( (not A234)  and  (not A233) );
 a43918a <=( A203  and  a43917a );
 a43921a <=( (not A267)  and  (not A266) );
 a43924a <=( (not A300)  and  A298 );
 a43925a <=( a43924a  and  a43921a );
 a43926a <=( a43925a  and  a43918a );
 a43930a <=( (not A166)  and  (not A167) );
 a43931a <=( A170  and  a43930a );
 a43935a <=( A201  and  (not A200) );
 a43936a <=( A199  and  a43935a );
 a43937a <=( a43936a  and  a43931a );
 a43941a <=( (not A234)  and  (not A233) );
 a43942a <=( A203  and  a43941a );
 a43945a <=( (not A267)  and  (not A266) );
 a43948a <=( A299  and  A298 );
 a43949a <=( a43948a  and  a43945a );
 a43950a <=( a43949a  and  a43942a );
 a43954a <=( (not A166)  and  (not A167) );
 a43955a <=( A170  and  a43954a );
 a43959a <=( A201  and  (not A200) );
 a43960a <=( A199  and  a43959a );
 a43961a <=( a43960a  and  a43955a );
 a43965a <=( (not A234)  and  (not A233) );
 a43966a <=( A203  and  a43965a );
 a43969a <=( (not A267)  and  (not A266) );
 a43972a <=( (not A299)  and  (not A298) );
 a43973a <=( a43972a  and  a43969a );
 a43974a <=( a43973a  and  a43966a );
 a43978a <=( (not A166)  and  (not A167) );
 a43979a <=( A170  and  a43978a );
 a43983a <=( A201  and  (not A200) );
 a43984a <=( A199  and  a43983a );
 a43985a <=( a43984a  and  a43979a );
 a43989a <=( (not A234)  and  (not A233) );
 a43990a <=( A203  and  a43989a );
 a43993a <=( (not A266)  and  (not A265) );
 a43996a <=( (not A300)  and  A298 );
 a43997a <=( a43996a  and  a43993a );
 a43998a <=( a43997a  and  a43990a );
 a44002a <=( (not A166)  and  (not A167) );
 a44003a <=( A170  and  a44002a );
 a44007a <=( A201  and  (not A200) );
 a44008a <=( A199  and  a44007a );
 a44009a <=( a44008a  and  a44003a );
 a44013a <=( (not A234)  and  (not A233) );
 a44014a <=( A203  and  a44013a );
 a44017a <=( (not A266)  and  (not A265) );
 a44020a <=( A299  and  A298 );
 a44021a <=( a44020a  and  a44017a );
 a44022a <=( a44021a  and  a44014a );
 a44026a <=( (not A166)  and  (not A167) );
 a44027a <=( A170  and  a44026a );
 a44031a <=( A201  and  (not A200) );
 a44032a <=( A199  and  a44031a );
 a44033a <=( a44032a  and  a44027a );
 a44037a <=( (not A234)  and  (not A233) );
 a44038a <=( A203  and  a44037a );
 a44041a <=( (not A266)  and  (not A265) );
 a44044a <=( (not A299)  and  (not A298) );
 a44045a <=( a44044a  and  a44041a );
 a44046a <=( a44045a  and  a44038a );
 a44050a <=( (not A166)  and  (not A167) );
 a44051a <=( A170  and  a44050a );
 a44055a <=( A201  and  (not A200) );
 a44056a <=( A199  and  a44055a );
 a44057a <=( a44056a  and  a44051a );
 a44061a <=( (not A233)  and  A232 );
 a44062a <=( A203  and  a44061a );
 a44065a <=( A235  and  A234 );
 a44068a <=( A299  and  (not A298) );
 a44069a <=( a44068a  and  a44065a );
 a44070a <=( a44069a  and  a44062a );
 a44074a <=( (not A166)  and  (not A167) );
 a44075a <=( A170  and  a44074a );
 a44079a <=( A201  and  (not A200) );
 a44080a <=( A199  and  a44079a );
 a44081a <=( a44080a  and  a44075a );
 a44085a <=( (not A233)  and  A232 );
 a44086a <=( A203  and  a44085a );
 a44089a <=( A235  and  A234 );
 a44092a <=( A266  and  (not A265) );
 a44093a <=( a44092a  and  a44089a );
 a44094a <=( a44093a  and  a44086a );
 a44098a <=( (not A166)  and  (not A167) );
 a44099a <=( A170  and  a44098a );
 a44103a <=( A201  and  (not A200) );
 a44104a <=( A199  and  a44103a );
 a44105a <=( a44104a  and  a44099a );
 a44109a <=( (not A233)  and  A232 );
 a44110a <=( A203  and  a44109a );
 a44113a <=( A236  and  A234 );
 a44116a <=( A299  and  (not A298) );
 a44117a <=( a44116a  and  a44113a );
 a44118a <=( a44117a  and  a44110a );
 a44122a <=( (not A166)  and  (not A167) );
 a44123a <=( A170  and  a44122a );
 a44127a <=( A201  and  (not A200) );
 a44128a <=( A199  and  a44127a );
 a44129a <=( a44128a  and  a44123a );
 a44133a <=( (not A233)  and  A232 );
 a44134a <=( A203  and  a44133a );
 a44137a <=( A236  and  A234 );
 a44140a <=( A266  and  (not A265) );
 a44141a <=( a44140a  and  a44137a );
 a44142a <=( a44141a  and  a44134a );
 a44146a <=( (not A166)  and  (not A167) );
 a44147a <=( A170  and  a44146a );
 a44151a <=( A201  and  (not A200) );
 a44152a <=( A199  and  a44151a );
 a44153a <=( a44152a  and  a44147a );
 a44157a <=( (not A233)  and  (not A232) );
 a44158a <=( A203  and  a44157a );
 a44161a <=( A266  and  A265 );
 a44164a <=( (not A300)  and  A298 );
 a44165a <=( a44164a  and  a44161a );
 a44166a <=( a44165a  and  a44158a );
 a44170a <=( (not A166)  and  (not A167) );
 a44171a <=( A170  and  a44170a );
 a44175a <=( A201  and  (not A200) );
 a44176a <=( A199  and  a44175a );
 a44177a <=( a44176a  and  a44171a );
 a44181a <=( (not A233)  and  (not A232) );
 a44182a <=( A203  and  a44181a );
 a44185a <=( A266  and  A265 );
 a44188a <=( A299  and  A298 );
 a44189a <=( a44188a  and  a44185a );
 a44190a <=( a44189a  and  a44182a );
 a44194a <=( (not A166)  and  (not A167) );
 a44195a <=( A170  and  a44194a );
 a44199a <=( A201  and  (not A200) );
 a44200a <=( A199  and  a44199a );
 a44201a <=( a44200a  and  a44195a );
 a44205a <=( (not A233)  and  (not A232) );
 a44206a <=( A203  and  a44205a );
 a44209a <=( A266  and  A265 );
 a44212a <=( (not A299)  and  (not A298) );
 a44213a <=( a44212a  and  a44209a );
 a44214a <=( a44213a  and  a44206a );
 a44218a <=( (not A166)  and  (not A167) );
 a44219a <=( A170  and  a44218a );
 a44223a <=( A201  and  (not A200) );
 a44224a <=( A199  and  a44223a );
 a44225a <=( a44224a  and  a44219a );
 a44229a <=( (not A233)  and  (not A232) );
 a44230a <=( A203  and  a44229a );
 a44233a <=( (not A267)  and  (not A266) );
 a44236a <=( (not A300)  and  A298 );
 a44237a <=( a44236a  and  a44233a );
 a44238a <=( a44237a  and  a44230a );
 a44242a <=( (not A166)  and  (not A167) );
 a44243a <=( A170  and  a44242a );
 a44247a <=( A201  and  (not A200) );
 a44248a <=( A199  and  a44247a );
 a44249a <=( a44248a  and  a44243a );
 a44253a <=( (not A233)  and  (not A232) );
 a44254a <=( A203  and  a44253a );
 a44257a <=( (not A267)  and  (not A266) );
 a44260a <=( A299  and  A298 );
 a44261a <=( a44260a  and  a44257a );
 a44262a <=( a44261a  and  a44254a );
 a44266a <=( (not A166)  and  (not A167) );
 a44267a <=( A170  and  a44266a );
 a44271a <=( A201  and  (not A200) );
 a44272a <=( A199  and  a44271a );
 a44273a <=( a44272a  and  a44267a );
 a44277a <=( (not A233)  and  (not A232) );
 a44278a <=( A203  and  a44277a );
 a44281a <=( (not A267)  and  (not A266) );
 a44284a <=( (not A299)  and  (not A298) );
 a44285a <=( a44284a  and  a44281a );
 a44286a <=( a44285a  and  a44278a );
 a44290a <=( (not A166)  and  (not A167) );
 a44291a <=( A170  and  a44290a );
 a44295a <=( A201  and  (not A200) );
 a44296a <=( A199  and  a44295a );
 a44297a <=( a44296a  and  a44291a );
 a44301a <=( (not A233)  and  (not A232) );
 a44302a <=( A203  and  a44301a );
 a44305a <=( (not A266)  and  (not A265) );
 a44308a <=( (not A300)  and  A298 );
 a44309a <=( a44308a  and  a44305a );
 a44310a <=( a44309a  and  a44302a );
 a44314a <=( (not A166)  and  (not A167) );
 a44315a <=( A170  and  a44314a );
 a44319a <=( A201  and  (not A200) );
 a44320a <=( A199  and  a44319a );
 a44321a <=( a44320a  and  a44315a );
 a44325a <=( (not A233)  and  (not A232) );
 a44326a <=( A203  and  a44325a );
 a44329a <=( (not A266)  and  (not A265) );
 a44332a <=( A299  and  A298 );
 a44333a <=( a44332a  and  a44329a );
 a44334a <=( a44333a  and  a44326a );
 a44338a <=( (not A166)  and  (not A167) );
 a44339a <=( A170  and  a44338a );
 a44343a <=( A201  and  (not A200) );
 a44344a <=( A199  and  a44343a );
 a44345a <=( a44344a  and  a44339a );
 a44349a <=( (not A233)  and  (not A232) );
 a44350a <=( A203  and  a44349a );
 a44353a <=( (not A266)  and  (not A265) );
 a44356a <=( (not A299)  and  (not A298) );
 a44357a <=( a44356a  and  a44353a );
 a44358a <=( a44357a  and  a44350a );
 a44362a <=( A167  and  (not A168) );
 a44363a <=( A170  and  a44362a );
 a44367a <=( A200  and  (not A199) );
 a44368a <=( A166  and  a44367a );
 a44369a <=( a44368a  and  a44363a );
 a44373a <=( A265  and  A233 );
 a44374a <=( A232  and  a44373a );
 a44377a <=( (not A269)  and  (not A268) );
 a44380a <=( (not A300)  and  (not A299) );
 a44381a <=( a44380a  and  a44377a );
 a44382a <=( a44381a  and  a44374a );
 a44386a <=( A167  and  (not A168) );
 a44387a <=( A170  and  a44386a );
 a44391a <=( A200  and  (not A199) );
 a44392a <=( A166  and  a44391a );
 a44393a <=( a44392a  and  a44387a );
 a44397a <=( A265  and  A233 );
 a44398a <=( A232  and  a44397a );
 a44401a <=( (not A269)  and  (not A268) );
 a44404a <=( A299  and  A298 );
 a44405a <=( a44404a  and  a44401a );
 a44406a <=( a44405a  and  a44398a );
 a44410a <=( A167  and  (not A168) );
 a44411a <=( A170  and  a44410a );
 a44415a <=( A200  and  (not A199) );
 a44416a <=( A166  and  a44415a );
 a44417a <=( a44416a  and  a44411a );
 a44421a <=( A265  and  A233 );
 a44422a <=( A232  and  a44421a );
 a44425a <=( (not A269)  and  (not A268) );
 a44428a <=( (not A299)  and  (not A298) );
 a44429a <=( a44428a  and  a44425a );
 a44430a <=( a44429a  and  a44422a );
 a44434a <=( A167  and  (not A168) );
 a44435a <=( A170  and  a44434a );
 a44439a <=( A200  and  (not A199) );
 a44440a <=( A166  and  a44439a );
 a44441a <=( a44440a  and  a44435a );
 a44445a <=( A265  and  A233 );
 a44446a <=( A232  and  a44445a );
 a44449a <=( (not A299)  and  (not A267) );
 a44452a <=( (not A302)  and  (not A301) );
 a44453a <=( a44452a  and  a44449a );
 a44454a <=( a44453a  and  a44446a );
 a44458a <=( A167  and  (not A168) );
 a44459a <=( A170  and  a44458a );
 a44463a <=( A200  and  (not A199) );
 a44464a <=( A166  and  a44463a );
 a44465a <=( a44464a  and  a44459a );
 a44469a <=( A265  and  A233 );
 a44470a <=( A232  and  a44469a );
 a44473a <=( (not A299)  and  A266 );
 a44476a <=( (not A302)  and  (not A301) );
 a44477a <=( a44476a  and  a44473a );
 a44478a <=( a44477a  and  a44470a );
 a44482a <=( A167  and  (not A168) );
 a44483a <=( A170  and  a44482a );
 a44487a <=( A200  and  (not A199) );
 a44488a <=( A166  and  a44487a );
 a44489a <=( a44488a  and  a44483a );
 a44493a <=( (not A265)  and  A233 );
 a44494a <=( A232  and  a44493a );
 a44497a <=( (not A299)  and  (not A266) );
 a44500a <=( (not A302)  and  (not A301) );
 a44501a <=( a44500a  and  a44497a );
 a44502a <=( a44501a  and  a44494a );
 a44506a <=( A167  and  (not A168) );
 a44507a <=( A170  and  a44506a );
 a44511a <=( A200  and  (not A199) );
 a44512a <=( A166  and  a44511a );
 a44513a <=( a44512a  and  a44507a );
 a44517a <=( (not A236)  and  (not A235) );
 a44518a <=( (not A233)  and  a44517a );
 a44521a <=( A266  and  A265 );
 a44524a <=( (not A300)  and  A298 );
 a44525a <=( a44524a  and  a44521a );
 a44526a <=( a44525a  and  a44518a );
 a44530a <=( A167  and  (not A168) );
 a44531a <=( A170  and  a44530a );
 a44535a <=( A200  and  (not A199) );
 a44536a <=( A166  and  a44535a );
 a44537a <=( a44536a  and  a44531a );
 a44541a <=( (not A236)  and  (not A235) );
 a44542a <=( (not A233)  and  a44541a );
 a44545a <=( A266  and  A265 );
 a44548a <=( A299  and  A298 );
 a44549a <=( a44548a  and  a44545a );
 a44550a <=( a44549a  and  a44542a );
 a44554a <=( A167  and  (not A168) );
 a44555a <=( A170  and  a44554a );
 a44559a <=( A200  and  (not A199) );
 a44560a <=( A166  and  a44559a );
 a44561a <=( a44560a  and  a44555a );
 a44565a <=( (not A236)  and  (not A235) );
 a44566a <=( (not A233)  and  a44565a );
 a44569a <=( A266  and  A265 );
 a44572a <=( (not A299)  and  (not A298) );
 a44573a <=( a44572a  and  a44569a );
 a44574a <=( a44573a  and  a44566a );
 a44578a <=( A167  and  (not A168) );
 a44579a <=( A170  and  a44578a );
 a44583a <=( A200  and  (not A199) );
 a44584a <=( A166  and  a44583a );
 a44585a <=( a44584a  and  a44579a );
 a44589a <=( (not A236)  and  (not A235) );
 a44590a <=( (not A233)  and  a44589a );
 a44593a <=( (not A267)  and  (not A266) );
 a44596a <=( (not A300)  and  A298 );
 a44597a <=( a44596a  and  a44593a );
 a44598a <=( a44597a  and  a44590a );
 a44602a <=( A167  and  (not A168) );
 a44603a <=( A170  and  a44602a );
 a44607a <=( A200  and  (not A199) );
 a44608a <=( A166  and  a44607a );
 a44609a <=( a44608a  and  a44603a );
 a44613a <=( (not A236)  and  (not A235) );
 a44614a <=( (not A233)  and  a44613a );
 a44617a <=( (not A267)  and  (not A266) );
 a44620a <=( A299  and  A298 );
 a44621a <=( a44620a  and  a44617a );
 a44622a <=( a44621a  and  a44614a );
 a44626a <=( A167  and  (not A168) );
 a44627a <=( A170  and  a44626a );
 a44631a <=( A200  and  (not A199) );
 a44632a <=( A166  and  a44631a );
 a44633a <=( a44632a  and  a44627a );
 a44637a <=( (not A236)  and  (not A235) );
 a44638a <=( (not A233)  and  a44637a );
 a44641a <=( (not A267)  and  (not A266) );
 a44644a <=( (not A299)  and  (not A298) );
 a44645a <=( a44644a  and  a44641a );
 a44646a <=( a44645a  and  a44638a );
 a44650a <=( A167  and  (not A168) );
 a44651a <=( A170  and  a44650a );
 a44655a <=( A200  and  (not A199) );
 a44656a <=( A166  and  a44655a );
 a44657a <=( a44656a  and  a44651a );
 a44661a <=( (not A236)  and  (not A235) );
 a44662a <=( (not A233)  and  a44661a );
 a44665a <=( (not A266)  and  (not A265) );
 a44668a <=( (not A300)  and  A298 );
 a44669a <=( a44668a  and  a44665a );
 a44670a <=( a44669a  and  a44662a );
 a44674a <=( A167  and  (not A168) );
 a44675a <=( A170  and  a44674a );
 a44679a <=( A200  and  (not A199) );
 a44680a <=( A166  and  a44679a );
 a44681a <=( a44680a  and  a44675a );
 a44685a <=( (not A236)  and  (not A235) );
 a44686a <=( (not A233)  and  a44685a );
 a44689a <=( (not A266)  and  (not A265) );
 a44692a <=( A299  and  A298 );
 a44693a <=( a44692a  and  a44689a );
 a44694a <=( a44693a  and  a44686a );
 a44698a <=( A167  and  (not A168) );
 a44699a <=( A170  and  a44698a );
 a44703a <=( A200  and  (not A199) );
 a44704a <=( A166  and  a44703a );
 a44705a <=( a44704a  and  a44699a );
 a44709a <=( (not A236)  and  (not A235) );
 a44710a <=( (not A233)  and  a44709a );
 a44713a <=( (not A266)  and  (not A265) );
 a44716a <=( (not A299)  and  (not A298) );
 a44717a <=( a44716a  and  a44713a );
 a44718a <=( a44717a  and  a44710a );
 a44722a <=( A167  and  (not A168) );
 a44723a <=( A170  and  a44722a );
 a44727a <=( A200  and  (not A199) );
 a44728a <=( A166  and  a44727a );
 a44729a <=( a44728a  and  a44723a );
 a44733a <=( A265  and  (not A234) );
 a44734a <=( (not A233)  and  a44733a );
 a44737a <=( A298  and  A266 );
 a44740a <=( (not A302)  and  (not A301) );
 a44741a <=( a44740a  and  a44737a );
 a44742a <=( a44741a  and  a44734a );
 a44746a <=( A167  and  (not A168) );
 a44747a <=( A170  and  a44746a );
 a44751a <=( A200  and  (not A199) );
 a44752a <=( A166  and  a44751a );
 a44753a <=( a44752a  and  a44747a );
 a44757a <=( (not A266)  and  (not A234) );
 a44758a <=( (not A233)  and  a44757a );
 a44761a <=( (not A269)  and  (not A268) );
 a44764a <=( (not A300)  and  A298 );
 a44765a <=( a44764a  and  a44761a );
 a44766a <=( a44765a  and  a44758a );
 a44770a <=( A167  and  (not A168) );
 a44771a <=( A170  and  a44770a );
 a44775a <=( A200  and  (not A199) );
 a44776a <=( A166  and  a44775a );
 a44777a <=( a44776a  and  a44771a );
 a44781a <=( (not A266)  and  (not A234) );
 a44782a <=( (not A233)  and  a44781a );
 a44785a <=( (not A269)  and  (not A268) );
 a44788a <=( A299  and  A298 );
 a44789a <=( a44788a  and  a44785a );
 a44790a <=( a44789a  and  a44782a );
 a44794a <=( A167  and  (not A168) );
 a44795a <=( A170  and  a44794a );
 a44799a <=( A200  and  (not A199) );
 a44800a <=( A166  and  a44799a );
 a44801a <=( a44800a  and  a44795a );
 a44805a <=( (not A266)  and  (not A234) );
 a44806a <=( (not A233)  and  a44805a );
 a44809a <=( (not A269)  and  (not A268) );
 a44812a <=( (not A299)  and  (not A298) );
 a44813a <=( a44812a  and  a44809a );
 a44814a <=( a44813a  and  a44806a );
 a44818a <=( A167  and  (not A168) );
 a44819a <=( A170  and  a44818a );
 a44823a <=( A200  and  (not A199) );
 a44824a <=( A166  and  a44823a );
 a44825a <=( a44824a  and  a44819a );
 a44829a <=( (not A266)  and  (not A234) );
 a44830a <=( (not A233)  and  a44829a );
 a44833a <=( A298  and  (not A267) );
 a44836a <=( (not A302)  and  (not A301) );
 a44837a <=( a44836a  and  a44833a );
 a44838a <=( a44837a  and  a44830a );
 a44842a <=( A167  and  (not A168) );
 a44843a <=( A170  and  a44842a );
 a44847a <=( A200  and  (not A199) );
 a44848a <=( A166  and  a44847a );
 a44849a <=( a44848a  and  a44843a );
 a44853a <=( (not A265)  and  (not A234) );
 a44854a <=( (not A233)  and  a44853a );
 a44857a <=( A298  and  (not A266) );
 a44860a <=( (not A302)  and  (not A301) );
 a44861a <=( a44860a  and  a44857a );
 a44862a <=( a44861a  and  a44854a );
 a44866a <=( A167  and  (not A168) );
 a44867a <=( A170  and  a44866a );
 a44871a <=( A200  and  (not A199) );
 a44872a <=( A166  and  a44871a );
 a44873a <=( a44872a  and  a44867a );
 a44877a <=( A265  and  (not A233) );
 a44878a <=( (not A232)  and  a44877a );
 a44881a <=( A298  and  A266 );
 a44884a <=( (not A302)  and  (not A301) );
 a44885a <=( a44884a  and  a44881a );
 a44886a <=( a44885a  and  a44878a );
 a44890a <=( A167  and  (not A168) );
 a44891a <=( A170  and  a44890a );
 a44895a <=( A200  and  (not A199) );
 a44896a <=( A166  and  a44895a );
 a44897a <=( a44896a  and  a44891a );
 a44901a <=( (not A266)  and  (not A233) );
 a44902a <=( (not A232)  and  a44901a );
 a44905a <=( (not A269)  and  (not A268) );
 a44908a <=( (not A300)  and  A298 );
 a44909a <=( a44908a  and  a44905a );
 a44910a <=( a44909a  and  a44902a );
 a44914a <=( A167  and  (not A168) );
 a44915a <=( A170  and  a44914a );
 a44919a <=( A200  and  (not A199) );
 a44920a <=( A166  and  a44919a );
 a44921a <=( a44920a  and  a44915a );
 a44925a <=( (not A266)  and  (not A233) );
 a44926a <=( (not A232)  and  a44925a );
 a44929a <=( (not A269)  and  (not A268) );
 a44932a <=( A299  and  A298 );
 a44933a <=( a44932a  and  a44929a );
 a44934a <=( a44933a  and  a44926a );
 a44938a <=( A167  and  (not A168) );
 a44939a <=( A170  and  a44938a );
 a44943a <=( A200  and  (not A199) );
 a44944a <=( A166  and  a44943a );
 a44945a <=( a44944a  and  a44939a );
 a44949a <=( (not A266)  and  (not A233) );
 a44950a <=( (not A232)  and  a44949a );
 a44953a <=( (not A269)  and  (not A268) );
 a44956a <=( (not A299)  and  (not A298) );
 a44957a <=( a44956a  and  a44953a );
 a44958a <=( a44957a  and  a44950a );
 a44962a <=( A167  and  (not A168) );
 a44963a <=( A170  and  a44962a );
 a44967a <=( A200  and  (not A199) );
 a44968a <=( A166  and  a44967a );
 a44969a <=( a44968a  and  a44963a );
 a44973a <=( (not A266)  and  (not A233) );
 a44974a <=( (not A232)  and  a44973a );
 a44977a <=( A298  and  (not A267) );
 a44980a <=( (not A302)  and  (not A301) );
 a44981a <=( a44980a  and  a44977a );
 a44982a <=( a44981a  and  a44974a );
 a44986a <=( A167  and  (not A168) );
 a44987a <=( A170  and  a44986a );
 a44991a <=( A200  and  (not A199) );
 a44992a <=( A166  and  a44991a );
 a44993a <=( a44992a  and  a44987a );
 a44997a <=( (not A265)  and  (not A233) );
 a44998a <=( (not A232)  and  a44997a );
 a45001a <=( A298  and  (not A266) );
 a45004a <=( (not A302)  and  (not A301) );
 a45005a <=( a45004a  and  a45001a );
 a45006a <=( a45005a  and  a44998a );
 a45010a <=( A167  and  (not A168) );
 a45011a <=( (not A170)  and  a45010a );
 a45015a <=( A200  and  (not A199) );
 a45016a <=( (not A166)  and  a45015a );
 a45017a <=( a45016a  and  a45011a );
 a45021a <=( A265  and  A233 );
 a45022a <=( A232  and  a45021a );
 a45025a <=( (not A269)  and  (not A268) );
 a45028a <=( (not A300)  and  (not A299) );
 a45029a <=( a45028a  and  a45025a );
 a45030a <=( a45029a  and  a45022a );
 a45034a <=( A167  and  (not A168) );
 a45035a <=( (not A170)  and  a45034a );
 a45039a <=( A200  and  (not A199) );
 a45040a <=( (not A166)  and  a45039a );
 a45041a <=( a45040a  and  a45035a );
 a45045a <=( A265  and  A233 );
 a45046a <=( A232  and  a45045a );
 a45049a <=( (not A269)  and  (not A268) );
 a45052a <=( A299  and  A298 );
 a45053a <=( a45052a  and  a45049a );
 a45054a <=( a45053a  and  a45046a );
 a45058a <=( A167  and  (not A168) );
 a45059a <=( (not A170)  and  a45058a );
 a45063a <=( A200  and  (not A199) );
 a45064a <=( (not A166)  and  a45063a );
 a45065a <=( a45064a  and  a45059a );
 a45069a <=( A265  and  A233 );
 a45070a <=( A232  and  a45069a );
 a45073a <=( (not A269)  and  (not A268) );
 a45076a <=( (not A299)  and  (not A298) );
 a45077a <=( a45076a  and  a45073a );
 a45078a <=( a45077a  and  a45070a );
 a45082a <=( A167  and  (not A168) );
 a45083a <=( (not A170)  and  a45082a );
 a45087a <=( A200  and  (not A199) );
 a45088a <=( (not A166)  and  a45087a );
 a45089a <=( a45088a  and  a45083a );
 a45093a <=( A265  and  A233 );
 a45094a <=( A232  and  a45093a );
 a45097a <=( (not A299)  and  (not A267) );
 a45100a <=( (not A302)  and  (not A301) );
 a45101a <=( a45100a  and  a45097a );
 a45102a <=( a45101a  and  a45094a );
 a45106a <=( A167  and  (not A168) );
 a45107a <=( (not A170)  and  a45106a );
 a45111a <=( A200  and  (not A199) );
 a45112a <=( (not A166)  and  a45111a );
 a45113a <=( a45112a  and  a45107a );
 a45117a <=( A265  and  A233 );
 a45118a <=( A232  and  a45117a );
 a45121a <=( (not A299)  and  A266 );
 a45124a <=( (not A302)  and  (not A301) );
 a45125a <=( a45124a  and  a45121a );
 a45126a <=( a45125a  and  a45118a );
 a45130a <=( A167  and  (not A168) );
 a45131a <=( (not A170)  and  a45130a );
 a45135a <=( A200  and  (not A199) );
 a45136a <=( (not A166)  and  a45135a );
 a45137a <=( a45136a  and  a45131a );
 a45141a <=( (not A265)  and  A233 );
 a45142a <=( A232  and  a45141a );
 a45145a <=( (not A299)  and  (not A266) );
 a45148a <=( (not A302)  and  (not A301) );
 a45149a <=( a45148a  and  a45145a );
 a45150a <=( a45149a  and  a45142a );
 a45154a <=( A167  and  (not A168) );
 a45155a <=( (not A170)  and  a45154a );
 a45159a <=( A200  and  (not A199) );
 a45160a <=( (not A166)  and  a45159a );
 a45161a <=( a45160a  and  a45155a );
 a45165a <=( (not A236)  and  (not A235) );
 a45166a <=( (not A233)  and  a45165a );
 a45169a <=( A266  and  A265 );
 a45172a <=( (not A300)  and  A298 );
 a45173a <=( a45172a  and  a45169a );
 a45174a <=( a45173a  and  a45166a );
 a45178a <=( A167  and  (not A168) );
 a45179a <=( (not A170)  and  a45178a );
 a45183a <=( A200  and  (not A199) );
 a45184a <=( (not A166)  and  a45183a );
 a45185a <=( a45184a  and  a45179a );
 a45189a <=( (not A236)  and  (not A235) );
 a45190a <=( (not A233)  and  a45189a );
 a45193a <=( A266  and  A265 );
 a45196a <=( A299  and  A298 );
 a45197a <=( a45196a  and  a45193a );
 a45198a <=( a45197a  and  a45190a );
 a45202a <=( A167  and  (not A168) );
 a45203a <=( (not A170)  and  a45202a );
 a45207a <=( A200  and  (not A199) );
 a45208a <=( (not A166)  and  a45207a );
 a45209a <=( a45208a  and  a45203a );
 a45213a <=( (not A236)  and  (not A235) );
 a45214a <=( (not A233)  and  a45213a );
 a45217a <=( A266  and  A265 );
 a45220a <=( (not A299)  and  (not A298) );
 a45221a <=( a45220a  and  a45217a );
 a45222a <=( a45221a  and  a45214a );
 a45226a <=( A167  and  (not A168) );
 a45227a <=( (not A170)  and  a45226a );
 a45231a <=( A200  and  (not A199) );
 a45232a <=( (not A166)  and  a45231a );
 a45233a <=( a45232a  and  a45227a );
 a45237a <=( (not A236)  and  (not A235) );
 a45238a <=( (not A233)  and  a45237a );
 a45241a <=( (not A267)  and  (not A266) );
 a45244a <=( (not A300)  and  A298 );
 a45245a <=( a45244a  and  a45241a );
 a45246a <=( a45245a  and  a45238a );
 a45250a <=( A167  and  (not A168) );
 a45251a <=( (not A170)  and  a45250a );
 a45255a <=( A200  and  (not A199) );
 a45256a <=( (not A166)  and  a45255a );
 a45257a <=( a45256a  and  a45251a );
 a45261a <=( (not A236)  and  (not A235) );
 a45262a <=( (not A233)  and  a45261a );
 a45265a <=( (not A267)  and  (not A266) );
 a45268a <=( A299  and  A298 );
 a45269a <=( a45268a  and  a45265a );
 a45270a <=( a45269a  and  a45262a );
 a45274a <=( A167  and  (not A168) );
 a45275a <=( (not A170)  and  a45274a );
 a45279a <=( A200  and  (not A199) );
 a45280a <=( (not A166)  and  a45279a );
 a45281a <=( a45280a  and  a45275a );
 a45285a <=( (not A236)  and  (not A235) );
 a45286a <=( (not A233)  and  a45285a );
 a45289a <=( (not A267)  and  (not A266) );
 a45292a <=( (not A299)  and  (not A298) );
 a45293a <=( a45292a  and  a45289a );
 a45294a <=( a45293a  and  a45286a );
 a45298a <=( A167  and  (not A168) );
 a45299a <=( (not A170)  and  a45298a );
 a45303a <=( A200  and  (not A199) );
 a45304a <=( (not A166)  and  a45303a );
 a45305a <=( a45304a  and  a45299a );
 a45309a <=( (not A236)  and  (not A235) );
 a45310a <=( (not A233)  and  a45309a );
 a45313a <=( (not A266)  and  (not A265) );
 a45316a <=( (not A300)  and  A298 );
 a45317a <=( a45316a  and  a45313a );
 a45318a <=( a45317a  and  a45310a );
 a45322a <=( A167  and  (not A168) );
 a45323a <=( (not A170)  and  a45322a );
 a45327a <=( A200  and  (not A199) );
 a45328a <=( (not A166)  and  a45327a );
 a45329a <=( a45328a  and  a45323a );
 a45333a <=( (not A236)  and  (not A235) );
 a45334a <=( (not A233)  and  a45333a );
 a45337a <=( (not A266)  and  (not A265) );
 a45340a <=( A299  and  A298 );
 a45341a <=( a45340a  and  a45337a );
 a45342a <=( a45341a  and  a45334a );
 a45346a <=( A167  and  (not A168) );
 a45347a <=( (not A170)  and  a45346a );
 a45351a <=( A200  and  (not A199) );
 a45352a <=( (not A166)  and  a45351a );
 a45353a <=( a45352a  and  a45347a );
 a45357a <=( (not A236)  and  (not A235) );
 a45358a <=( (not A233)  and  a45357a );
 a45361a <=( (not A266)  and  (not A265) );
 a45364a <=( (not A299)  and  (not A298) );
 a45365a <=( a45364a  and  a45361a );
 a45366a <=( a45365a  and  a45358a );
 a45370a <=( A167  and  (not A168) );
 a45371a <=( (not A170)  and  a45370a );
 a45375a <=( A200  and  (not A199) );
 a45376a <=( (not A166)  and  a45375a );
 a45377a <=( a45376a  and  a45371a );
 a45381a <=( A265  and  (not A234) );
 a45382a <=( (not A233)  and  a45381a );
 a45385a <=( A298  and  A266 );
 a45388a <=( (not A302)  and  (not A301) );
 a45389a <=( a45388a  and  a45385a );
 a45390a <=( a45389a  and  a45382a );
 a45394a <=( A167  and  (not A168) );
 a45395a <=( (not A170)  and  a45394a );
 a45399a <=( A200  and  (not A199) );
 a45400a <=( (not A166)  and  a45399a );
 a45401a <=( a45400a  and  a45395a );
 a45405a <=( (not A266)  and  (not A234) );
 a45406a <=( (not A233)  and  a45405a );
 a45409a <=( (not A269)  and  (not A268) );
 a45412a <=( (not A300)  and  A298 );
 a45413a <=( a45412a  and  a45409a );
 a45414a <=( a45413a  and  a45406a );
 a45418a <=( A167  and  (not A168) );
 a45419a <=( (not A170)  and  a45418a );
 a45423a <=( A200  and  (not A199) );
 a45424a <=( (not A166)  and  a45423a );
 a45425a <=( a45424a  and  a45419a );
 a45429a <=( (not A266)  and  (not A234) );
 a45430a <=( (not A233)  and  a45429a );
 a45433a <=( (not A269)  and  (not A268) );
 a45436a <=( A299  and  A298 );
 a45437a <=( a45436a  and  a45433a );
 a45438a <=( a45437a  and  a45430a );
 a45442a <=( A167  and  (not A168) );
 a45443a <=( (not A170)  and  a45442a );
 a45447a <=( A200  and  (not A199) );
 a45448a <=( (not A166)  and  a45447a );
 a45449a <=( a45448a  and  a45443a );
 a45453a <=( (not A266)  and  (not A234) );
 a45454a <=( (not A233)  and  a45453a );
 a45457a <=( (not A269)  and  (not A268) );
 a45460a <=( (not A299)  and  (not A298) );
 a45461a <=( a45460a  and  a45457a );
 a45462a <=( a45461a  and  a45454a );
 a45466a <=( A167  and  (not A168) );
 a45467a <=( (not A170)  and  a45466a );
 a45471a <=( A200  and  (not A199) );
 a45472a <=( (not A166)  and  a45471a );
 a45473a <=( a45472a  and  a45467a );
 a45477a <=( (not A266)  and  (not A234) );
 a45478a <=( (not A233)  and  a45477a );
 a45481a <=( A298  and  (not A267) );
 a45484a <=( (not A302)  and  (not A301) );
 a45485a <=( a45484a  and  a45481a );
 a45486a <=( a45485a  and  a45478a );
 a45490a <=( A167  and  (not A168) );
 a45491a <=( (not A170)  and  a45490a );
 a45495a <=( A200  and  (not A199) );
 a45496a <=( (not A166)  and  a45495a );
 a45497a <=( a45496a  and  a45491a );
 a45501a <=( (not A265)  and  (not A234) );
 a45502a <=( (not A233)  and  a45501a );
 a45505a <=( A298  and  (not A266) );
 a45508a <=( (not A302)  and  (not A301) );
 a45509a <=( a45508a  and  a45505a );
 a45510a <=( a45509a  and  a45502a );
 a45514a <=( A167  and  (not A168) );
 a45515a <=( (not A170)  and  a45514a );
 a45519a <=( A200  and  (not A199) );
 a45520a <=( (not A166)  and  a45519a );
 a45521a <=( a45520a  and  a45515a );
 a45525a <=( A265  and  (not A233) );
 a45526a <=( (not A232)  and  a45525a );
 a45529a <=( A298  and  A266 );
 a45532a <=( (not A302)  and  (not A301) );
 a45533a <=( a45532a  and  a45529a );
 a45534a <=( a45533a  and  a45526a );
 a45538a <=( A167  and  (not A168) );
 a45539a <=( (not A170)  and  a45538a );
 a45543a <=( A200  and  (not A199) );
 a45544a <=( (not A166)  and  a45543a );
 a45545a <=( a45544a  and  a45539a );
 a45549a <=( (not A266)  and  (not A233) );
 a45550a <=( (not A232)  and  a45549a );
 a45553a <=( (not A269)  and  (not A268) );
 a45556a <=( (not A300)  and  A298 );
 a45557a <=( a45556a  and  a45553a );
 a45558a <=( a45557a  and  a45550a );
 a45562a <=( A167  and  (not A168) );
 a45563a <=( (not A170)  and  a45562a );
 a45567a <=( A200  and  (not A199) );
 a45568a <=( (not A166)  and  a45567a );
 a45569a <=( a45568a  and  a45563a );
 a45573a <=( (not A266)  and  (not A233) );
 a45574a <=( (not A232)  and  a45573a );
 a45577a <=( (not A269)  and  (not A268) );
 a45580a <=( A299  and  A298 );
 a45581a <=( a45580a  and  a45577a );
 a45582a <=( a45581a  and  a45574a );
 a45586a <=( A167  and  (not A168) );
 a45587a <=( (not A170)  and  a45586a );
 a45591a <=( A200  and  (not A199) );
 a45592a <=( (not A166)  and  a45591a );
 a45593a <=( a45592a  and  a45587a );
 a45597a <=( (not A266)  and  (not A233) );
 a45598a <=( (not A232)  and  a45597a );
 a45601a <=( (not A269)  and  (not A268) );
 a45604a <=( (not A299)  and  (not A298) );
 a45605a <=( a45604a  and  a45601a );
 a45606a <=( a45605a  and  a45598a );
 a45610a <=( A167  and  (not A168) );
 a45611a <=( (not A170)  and  a45610a );
 a45615a <=( A200  and  (not A199) );
 a45616a <=( (not A166)  and  a45615a );
 a45617a <=( a45616a  and  a45611a );
 a45621a <=( (not A266)  and  (not A233) );
 a45622a <=( (not A232)  and  a45621a );
 a45625a <=( A298  and  (not A267) );
 a45628a <=( (not A302)  and  (not A301) );
 a45629a <=( a45628a  and  a45625a );
 a45630a <=( a45629a  and  a45622a );
 a45634a <=( A167  and  (not A168) );
 a45635a <=( (not A170)  and  a45634a );
 a45639a <=( A200  and  (not A199) );
 a45640a <=( (not A166)  and  a45639a );
 a45641a <=( a45640a  and  a45635a );
 a45645a <=( (not A265)  and  (not A233) );
 a45646a <=( (not A232)  and  a45645a );
 a45649a <=( A298  and  (not A266) );
 a45652a <=( (not A302)  and  (not A301) );
 a45653a <=( a45652a  and  a45649a );
 a45654a <=( a45653a  and  a45646a );
 a45658a <=( (not A167)  and  (not A168) );
 a45659a <=( (not A170)  and  a45658a );
 a45663a <=( A200  and  (not A199) );
 a45664a <=( A166  and  a45663a );
 a45665a <=( a45664a  and  a45659a );
 a45669a <=( A265  and  A233 );
 a45670a <=( A232  and  a45669a );
 a45673a <=( (not A269)  and  (not A268) );
 a45676a <=( (not A300)  and  (not A299) );
 a45677a <=( a45676a  and  a45673a );
 a45678a <=( a45677a  and  a45670a );
 a45682a <=( (not A167)  and  (not A168) );
 a45683a <=( (not A170)  and  a45682a );
 a45687a <=( A200  and  (not A199) );
 a45688a <=( A166  and  a45687a );
 a45689a <=( a45688a  and  a45683a );
 a45693a <=( A265  and  A233 );
 a45694a <=( A232  and  a45693a );
 a45697a <=( (not A269)  and  (not A268) );
 a45700a <=( A299  and  A298 );
 a45701a <=( a45700a  and  a45697a );
 a45702a <=( a45701a  and  a45694a );
 a45706a <=( (not A167)  and  (not A168) );
 a45707a <=( (not A170)  and  a45706a );
 a45711a <=( A200  and  (not A199) );
 a45712a <=( A166  and  a45711a );
 a45713a <=( a45712a  and  a45707a );
 a45717a <=( A265  and  A233 );
 a45718a <=( A232  and  a45717a );
 a45721a <=( (not A269)  and  (not A268) );
 a45724a <=( (not A299)  and  (not A298) );
 a45725a <=( a45724a  and  a45721a );
 a45726a <=( a45725a  and  a45718a );
 a45730a <=( (not A167)  and  (not A168) );
 a45731a <=( (not A170)  and  a45730a );
 a45735a <=( A200  and  (not A199) );
 a45736a <=( A166  and  a45735a );
 a45737a <=( a45736a  and  a45731a );
 a45741a <=( A265  and  A233 );
 a45742a <=( A232  and  a45741a );
 a45745a <=( (not A299)  and  (not A267) );
 a45748a <=( (not A302)  and  (not A301) );
 a45749a <=( a45748a  and  a45745a );
 a45750a <=( a45749a  and  a45742a );
 a45754a <=( (not A167)  and  (not A168) );
 a45755a <=( (not A170)  and  a45754a );
 a45759a <=( A200  and  (not A199) );
 a45760a <=( A166  and  a45759a );
 a45761a <=( a45760a  and  a45755a );
 a45765a <=( A265  and  A233 );
 a45766a <=( A232  and  a45765a );
 a45769a <=( (not A299)  and  A266 );
 a45772a <=( (not A302)  and  (not A301) );
 a45773a <=( a45772a  and  a45769a );
 a45774a <=( a45773a  and  a45766a );
 a45778a <=( (not A167)  and  (not A168) );
 a45779a <=( (not A170)  and  a45778a );
 a45783a <=( A200  and  (not A199) );
 a45784a <=( A166  and  a45783a );
 a45785a <=( a45784a  and  a45779a );
 a45789a <=( (not A265)  and  A233 );
 a45790a <=( A232  and  a45789a );
 a45793a <=( (not A299)  and  (not A266) );
 a45796a <=( (not A302)  and  (not A301) );
 a45797a <=( a45796a  and  a45793a );
 a45798a <=( a45797a  and  a45790a );
 a45802a <=( (not A167)  and  (not A168) );
 a45803a <=( (not A170)  and  a45802a );
 a45807a <=( A200  and  (not A199) );
 a45808a <=( A166  and  a45807a );
 a45809a <=( a45808a  and  a45803a );
 a45813a <=( (not A236)  and  (not A235) );
 a45814a <=( (not A233)  and  a45813a );
 a45817a <=( A266  and  A265 );
 a45820a <=( (not A300)  and  A298 );
 a45821a <=( a45820a  and  a45817a );
 a45822a <=( a45821a  and  a45814a );
 a45826a <=( (not A167)  and  (not A168) );
 a45827a <=( (not A170)  and  a45826a );
 a45831a <=( A200  and  (not A199) );
 a45832a <=( A166  and  a45831a );
 a45833a <=( a45832a  and  a45827a );
 a45837a <=( (not A236)  and  (not A235) );
 a45838a <=( (not A233)  and  a45837a );
 a45841a <=( A266  and  A265 );
 a45844a <=( A299  and  A298 );
 a45845a <=( a45844a  and  a45841a );
 a45846a <=( a45845a  and  a45838a );
 a45850a <=( (not A167)  and  (not A168) );
 a45851a <=( (not A170)  and  a45850a );
 a45855a <=( A200  and  (not A199) );
 a45856a <=( A166  and  a45855a );
 a45857a <=( a45856a  and  a45851a );
 a45861a <=( (not A236)  and  (not A235) );
 a45862a <=( (not A233)  and  a45861a );
 a45865a <=( A266  and  A265 );
 a45868a <=( (not A299)  and  (not A298) );
 a45869a <=( a45868a  and  a45865a );
 a45870a <=( a45869a  and  a45862a );
 a45874a <=( (not A167)  and  (not A168) );
 a45875a <=( (not A170)  and  a45874a );
 a45879a <=( A200  and  (not A199) );
 a45880a <=( A166  and  a45879a );
 a45881a <=( a45880a  and  a45875a );
 a45885a <=( (not A236)  and  (not A235) );
 a45886a <=( (not A233)  and  a45885a );
 a45889a <=( (not A267)  and  (not A266) );
 a45892a <=( (not A300)  and  A298 );
 a45893a <=( a45892a  and  a45889a );
 a45894a <=( a45893a  and  a45886a );
 a45898a <=( (not A167)  and  (not A168) );
 a45899a <=( (not A170)  and  a45898a );
 a45903a <=( A200  and  (not A199) );
 a45904a <=( A166  and  a45903a );
 a45905a <=( a45904a  and  a45899a );
 a45909a <=( (not A236)  and  (not A235) );
 a45910a <=( (not A233)  and  a45909a );
 a45913a <=( (not A267)  and  (not A266) );
 a45916a <=( A299  and  A298 );
 a45917a <=( a45916a  and  a45913a );
 a45918a <=( a45917a  and  a45910a );
 a45922a <=( (not A167)  and  (not A168) );
 a45923a <=( (not A170)  and  a45922a );
 a45927a <=( A200  and  (not A199) );
 a45928a <=( A166  and  a45927a );
 a45929a <=( a45928a  and  a45923a );
 a45933a <=( (not A236)  and  (not A235) );
 a45934a <=( (not A233)  and  a45933a );
 a45937a <=( (not A267)  and  (not A266) );
 a45940a <=( (not A299)  and  (not A298) );
 a45941a <=( a45940a  and  a45937a );
 a45942a <=( a45941a  and  a45934a );
 a45946a <=( (not A167)  and  (not A168) );
 a45947a <=( (not A170)  and  a45946a );
 a45951a <=( A200  and  (not A199) );
 a45952a <=( A166  and  a45951a );
 a45953a <=( a45952a  and  a45947a );
 a45957a <=( (not A236)  and  (not A235) );
 a45958a <=( (not A233)  and  a45957a );
 a45961a <=( (not A266)  and  (not A265) );
 a45964a <=( (not A300)  and  A298 );
 a45965a <=( a45964a  and  a45961a );
 a45966a <=( a45965a  and  a45958a );
 a45970a <=( (not A167)  and  (not A168) );
 a45971a <=( (not A170)  and  a45970a );
 a45975a <=( A200  and  (not A199) );
 a45976a <=( A166  and  a45975a );
 a45977a <=( a45976a  and  a45971a );
 a45981a <=( (not A236)  and  (not A235) );
 a45982a <=( (not A233)  and  a45981a );
 a45985a <=( (not A266)  and  (not A265) );
 a45988a <=( A299  and  A298 );
 a45989a <=( a45988a  and  a45985a );
 a45990a <=( a45989a  and  a45982a );
 a45994a <=( (not A167)  and  (not A168) );
 a45995a <=( (not A170)  and  a45994a );
 a45999a <=( A200  and  (not A199) );
 a46000a <=( A166  and  a45999a );
 a46001a <=( a46000a  and  a45995a );
 a46005a <=( (not A236)  and  (not A235) );
 a46006a <=( (not A233)  and  a46005a );
 a46009a <=( (not A266)  and  (not A265) );
 a46012a <=( (not A299)  and  (not A298) );
 a46013a <=( a46012a  and  a46009a );
 a46014a <=( a46013a  and  a46006a );
 a46018a <=( (not A167)  and  (not A168) );
 a46019a <=( (not A170)  and  a46018a );
 a46023a <=( A200  and  (not A199) );
 a46024a <=( A166  and  a46023a );
 a46025a <=( a46024a  and  a46019a );
 a46029a <=( A265  and  (not A234) );
 a46030a <=( (not A233)  and  a46029a );
 a46033a <=( A298  and  A266 );
 a46036a <=( (not A302)  and  (not A301) );
 a46037a <=( a46036a  and  a46033a );
 a46038a <=( a46037a  and  a46030a );
 a46042a <=( (not A167)  and  (not A168) );
 a46043a <=( (not A170)  and  a46042a );
 a46047a <=( A200  and  (not A199) );
 a46048a <=( A166  and  a46047a );
 a46049a <=( a46048a  and  a46043a );
 a46053a <=( (not A266)  and  (not A234) );
 a46054a <=( (not A233)  and  a46053a );
 a46057a <=( (not A269)  and  (not A268) );
 a46060a <=( (not A300)  and  A298 );
 a46061a <=( a46060a  and  a46057a );
 a46062a <=( a46061a  and  a46054a );
 a46066a <=( (not A167)  and  (not A168) );
 a46067a <=( (not A170)  and  a46066a );
 a46071a <=( A200  and  (not A199) );
 a46072a <=( A166  and  a46071a );
 a46073a <=( a46072a  and  a46067a );
 a46077a <=( (not A266)  and  (not A234) );
 a46078a <=( (not A233)  and  a46077a );
 a46081a <=( (not A269)  and  (not A268) );
 a46084a <=( A299  and  A298 );
 a46085a <=( a46084a  and  a46081a );
 a46086a <=( a46085a  and  a46078a );
 a46090a <=( (not A167)  and  (not A168) );
 a46091a <=( (not A170)  and  a46090a );
 a46095a <=( A200  and  (not A199) );
 a46096a <=( A166  and  a46095a );
 a46097a <=( a46096a  and  a46091a );
 a46101a <=( (not A266)  and  (not A234) );
 a46102a <=( (not A233)  and  a46101a );
 a46105a <=( (not A269)  and  (not A268) );
 a46108a <=( (not A299)  and  (not A298) );
 a46109a <=( a46108a  and  a46105a );
 a46110a <=( a46109a  and  a46102a );
 a46114a <=( (not A167)  and  (not A168) );
 a46115a <=( (not A170)  and  a46114a );
 a46119a <=( A200  and  (not A199) );
 a46120a <=( A166  and  a46119a );
 a46121a <=( a46120a  and  a46115a );
 a46125a <=( (not A266)  and  (not A234) );
 a46126a <=( (not A233)  and  a46125a );
 a46129a <=( A298  and  (not A267) );
 a46132a <=( (not A302)  and  (not A301) );
 a46133a <=( a46132a  and  a46129a );
 a46134a <=( a46133a  and  a46126a );
 a46138a <=( (not A167)  and  (not A168) );
 a46139a <=( (not A170)  and  a46138a );
 a46143a <=( A200  and  (not A199) );
 a46144a <=( A166  and  a46143a );
 a46145a <=( a46144a  and  a46139a );
 a46149a <=( (not A265)  and  (not A234) );
 a46150a <=( (not A233)  and  a46149a );
 a46153a <=( A298  and  (not A266) );
 a46156a <=( (not A302)  and  (not A301) );
 a46157a <=( a46156a  and  a46153a );
 a46158a <=( a46157a  and  a46150a );
 a46162a <=( (not A167)  and  (not A168) );
 a46163a <=( (not A170)  and  a46162a );
 a46167a <=( A200  and  (not A199) );
 a46168a <=( A166  and  a46167a );
 a46169a <=( a46168a  and  a46163a );
 a46173a <=( A265  and  (not A233) );
 a46174a <=( (not A232)  and  a46173a );
 a46177a <=( A298  and  A266 );
 a46180a <=( (not A302)  and  (not A301) );
 a46181a <=( a46180a  and  a46177a );
 a46182a <=( a46181a  and  a46174a );
 a46186a <=( (not A167)  and  (not A168) );
 a46187a <=( (not A170)  and  a46186a );
 a46191a <=( A200  and  (not A199) );
 a46192a <=( A166  and  a46191a );
 a46193a <=( a46192a  and  a46187a );
 a46197a <=( (not A266)  and  (not A233) );
 a46198a <=( (not A232)  and  a46197a );
 a46201a <=( (not A269)  and  (not A268) );
 a46204a <=( (not A300)  and  A298 );
 a46205a <=( a46204a  and  a46201a );
 a46206a <=( a46205a  and  a46198a );
 a46210a <=( (not A167)  and  (not A168) );
 a46211a <=( (not A170)  and  a46210a );
 a46215a <=( A200  and  (not A199) );
 a46216a <=( A166  and  a46215a );
 a46217a <=( a46216a  and  a46211a );
 a46221a <=( (not A266)  and  (not A233) );
 a46222a <=( (not A232)  and  a46221a );
 a46225a <=( (not A269)  and  (not A268) );
 a46228a <=( A299  and  A298 );
 a46229a <=( a46228a  and  a46225a );
 a46230a <=( a46229a  and  a46222a );
 a46234a <=( (not A167)  and  (not A168) );
 a46235a <=( (not A170)  and  a46234a );
 a46239a <=( A200  and  (not A199) );
 a46240a <=( A166  and  a46239a );
 a46241a <=( a46240a  and  a46235a );
 a46245a <=( (not A266)  and  (not A233) );
 a46246a <=( (not A232)  and  a46245a );
 a46249a <=( (not A269)  and  (not A268) );
 a46252a <=( (not A299)  and  (not A298) );
 a46253a <=( a46252a  and  a46249a );
 a46254a <=( a46253a  and  a46246a );
 a46258a <=( (not A167)  and  (not A168) );
 a46259a <=( (not A170)  and  a46258a );
 a46263a <=( A200  and  (not A199) );
 a46264a <=( A166  and  a46263a );
 a46265a <=( a46264a  and  a46259a );
 a46269a <=( (not A266)  and  (not A233) );
 a46270a <=( (not A232)  and  a46269a );
 a46273a <=( A298  and  (not A267) );
 a46276a <=( (not A302)  and  (not A301) );
 a46277a <=( a46276a  and  a46273a );
 a46278a <=( a46277a  and  a46270a );
 a46282a <=( (not A167)  and  (not A168) );
 a46283a <=( (not A170)  and  a46282a );
 a46287a <=( A200  and  (not A199) );
 a46288a <=( A166  and  a46287a );
 a46289a <=( a46288a  and  a46283a );
 a46293a <=( (not A265)  and  (not A233) );
 a46294a <=( (not A232)  and  a46293a );
 a46297a <=( A298  and  (not A266) );
 a46300a <=( (not A302)  and  (not A301) );
 a46301a <=( a46300a  and  a46297a );
 a46302a <=( a46301a  and  a46294a );
 a46306a <=( A167  and  (not A168) );
 a46307a <=( A169  and  a46306a );
 a46311a <=( A200  and  (not A199) );
 a46312a <=( (not A166)  and  a46311a );
 a46313a <=( a46312a  and  a46307a );
 a46317a <=( A265  and  A233 );
 a46318a <=( A232  and  a46317a );
 a46321a <=( (not A269)  and  (not A268) );
 a46324a <=( (not A300)  and  (not A299) );
 a46325a <=( a46324a  and  a46321a );
 a46326a <=( a46325a  and  a46318a );
 a46330a <=( A167  and  (not A168) );
 a46331a <=( A169  and  a46330a );
 a46335a <=( A200  and  (not A199) );
 a46336a <=( (not A166)  and  a46335a );
 a46337a <=( a46336a  and  a46331a );
 a46341a <=( A265  and  A233 );
 a46342a <=( A232  and  a46341a );
 a46345a <=( (not A269)  and  (not A268) );
 a46348a <=( A299  and  A298 );
 a46349a <=( a46348a  and  a46345a );
 a46350a <=( a46349a  and  a46342a );
 a46354a <=( A167  and  (not A168) );
 a46355a <=( A169  and  a46354a );
 a46359a <=( A200  and  (not A199) );
 a46360a <=( (not A166)  and  a46359a );
 a46361a <=( a46360a  and  a46355a );
 a46365a <=( A265  and  A233 );
 a46366a <=( A232  and  a46365a );
 a46369a <=( (not A269)  and  (not A268) );
 a46372a <=( (not A299)  and  (not A298) );
 a46373a <=( a46372a  and  a46369a );
 a46374a <=( a46373a  and  a46366a );
 a46378a <=( A167  and  (not A168) );
 a46379a <=( A169  and  a46378a );
 a46383a <=( A200  and  (not A199) );
 a46384a <=( (not A166)  and  a46383a );
 a46385a <=( a46384a  and  a46379a );
 a46389a <=( A265  and  A233 );
 a46390a <=( A232  and  a46389a );
 a46393a <=( (not A299)  and  (not A267) );
 a46396a <=( (not A302)  and  (not A301) );
 a46397a <=( a46396a  and  a46393a );
 a46398a <=( a46397a  and  a46390a );
 a46402a <=( A167  and  (not A168) );
 a46403a <=( A169  and  a46402a );
 a46407a <=( A200  and  (not A199) );
 a46408a <=( (not A166)  and  a46407a );
 a46409a <=( a46408a  and  a46403a );
 a46413a <=( A265  and  A233 );
 a46414a <=( A232  and  a46413a );
 a46417a <=( (not A299)  and  A266 );
 a46420a <=( (not A302)  and  (not A301) );
 a46421a <=( a46420a  and  a46417a );
 a46422a <=( a46421a  and  a46414a );
 a46426a <=( A167  and  (not A168) );
 a46427a <=( A169  and  a46426a );
 a46431a <=( A200  and  (not A199) );
 a46432a <=( (not A166)  and  a46431a );
 a46433a <=( a46432a  and  a46427a );
 a46437a <=( (not A265)  and  A233 );
 a46438a <=( A232  and  a46437a );
 a46441a <=( (not A299)  and  (not A266) );
 a46444a <=( (not A302)  and  (not A301) );
 a46445a <=( a46444a  and  a46441a );
 a46446a <=( a46445a  and  a46438a );
 a46450a <=( A167  and  (not A168) );
 a46451a <=( A169  and  a46450a );
 a46455a <=( A200  and  (not A199) );
 a46456a <=( (not A166)  and  a46455a );
 a46457a <=( a46456a  and  a46451a );
 a46461a <=( (not A236)  and  (not A235) );
 a46462a <=( (not A233)  and  a46461a );
 a46465a <=( A266  and  A265 );
 a46468a <=( (not A300)  and  A298 );
 a46469a <=( a46468a  and  a46465a );
 a46470a <=( a46469a  and  a46462a );
 a46474a <=( A167  and  (not A168) );
 a46475a <=( A169  and  a46474a );
 a46479a <=( A200  and  (not A199) );
 a46480a <=( (not A166)  and  a46479a );
 a46481a <=( a46480a  and  a46475a );
 a46485a <=( (not A236)  and  (not A235) );
 a46486a <=( (not A233)  and  a46485a );
 a46489a <=( A266  and  A265 );
 a46492a <=( A299  and  A298 );
 a46493a <=( a46492a  and  a46489a );
 a46494a <=( a46493a  and  a46486a );
 a46498a <=( A167  and  (not A168) );
 a46499a <=( A169  and  a46498a );
 a46503a <=( A200  and  (not A199) );
 a46504a <=( (not A166)  and  a46503a );
 a46505a <=( a46504a  and  a46499a );
 a46509a <=( (not A236)  and  (not A235) );
 a46510a <=( (not A233)  and  a46509a );
 a46513a <=( A266  and  A265 );
 a46516a <=( (not A299)  and  (not A298) );
 a46517a <=( a46516a  and  a46513a );
 a46518a <=( a46517a  and  a46510a );
 a46522a <=( A167  and  (not A168) );
 a46523a <=( A169  and  a46522a );
 a46527a <=( A200  and  (not A199) );
 a46528a <=( (not A166)  and  a46527a );
 a46529a <=( a46528a  and  a46523a );
 a46533a <=( (not A236)  and  (not A235) );
 a46534a <=( (not A233)  and  a46533a );
 a46537a <=( (not A267)  and  (not A266) );
 a46540a <=( (not A300)  and  A298 );
 a46541a <=( a46540a  and  a46537a );
 a46542a <=( a46541a  and  a46534a );
 a46546a <=( A167  and  (not A168) );
 a46547a <=( A169  and  a46546a );
 a46551a <=( A200  and  (not A199) );
 a46552a <=( (not A166)  and  a46551a );
 a46553a <=( a46552a  and  a46547a );
 a46557a <=( (not A236)  and  (not A235) );
 a46558a <=( (not A233)  and  a46557a );
 a46561a <=( (not A267)  and  (not A266) );
 a46564a <=( A299  and  A298 );
 a46565a <=( a46564a  and  a46561a );
 a46566a <=( a46565a  and  a46558a );
 a46570a <=( A167  and  (not A168) );
 a46571a <=( A169  and  a46570a );
 a46575a <=( A200  and  (not A199) );
 a46576a <=( (not A166)  and  a46575a );
 a46577a <=( a46576a  and  a46571a );
 a46581a <=( (not A236)  and  (not A235) );
 a46582a <=( (not A233)  and  a46581a );
 a46585a <=( (not A267)  and  (not A266) );
 a46588a <=( (not A299)  and  (not A298) );
 a46589a <=( a46588a  and  a46585a );
 a46590a <=( a46589a  and  a46582a );
 a46594a <=( A167  and  (not A168) );
 a46595a <=( A169  and  a46594a );
 a46599a <=( A200  and  (not A199) );
 a46600a <=( (not A166)  and  a46599a );
 a46601a <=( a46600a  and  a46595a );
 a46605a <=( (not A236)  and  (not A235) );
 a46606a <=( (not A233)  and  a46605a );
 a46609a <=( (not A266)  and  (not A265) );
 a46612a <=( (not A300)  and  A298 );
 a46613a <=( a46612a  and  a46609a );
 a46614a <=( a46613a  and  a46606a );
 a46618a <=( A167  and  (not A168) );
 a46619a <=( A169  and  a46618a );
 a46623a <=( A200  and  (not A199) );
 a46624a <=( (not A166)  and  a46623a );
 a46625a <=( a46624a  and  a46619a );
 a46629a <=( (not A236)  and  (not A235) );
 a46630a <=( (not A233)  and  a46629a );
 a46633a <=( (not A266)  and  (not A265) );
 a46636a <=( A299  and  A298 );
 a46637a <=( a46636a  and  a46633a );
 a46638a <=( a46637a  and  a46630a );
 a46642a <=( A167  and  (not A168) );
 a46643a <=( A169  and  a46642a );
 a46647a <=( A200  and  (not A199) );
 a46648a <=( (not A166)  and  a46647a );
 a46649a <=( a46648a  and  a46643a );
 a46653a <=( (not A236)  and  (not A235) );
 a46654a <=( (not A233)  and  a46653a );
 a46657a <=( (not A266)  and  (not A265) );
 a46660a <=( (not A299)  and  (not A298) );
 a46661a <=( a46660a  and  a46657a );
 a46662a <=( a46661a  and  a46654a );
 a46666a <=( A167  and  (not A168) );
 a46667a <=( A169  and  a46666a );
 a46671a <=( A200  and  (not A199) );
 a46672a <=( (not A166)  and  a46671a );
 a46673a <=( a46672a  and  a46667a );
 a46677a <=( A265  and  (not A234) );
 a46678a <=( (not A233)  and  a46677a );
 a46681a <=( A298  and  A266 );
 a46684a <=( (not A302)  and  (not A301) );
 a46685a <=( a46684a  and  a46681a );
 a46686a <=( a46685a  and  a46678a );
 a46690a <=( A167  and  (not A168) );
 a46691a <=( A169  and  a46690a );
 a46695a <=( A200  and  (not A199) );
 a46696a <=( (not A166)  and  a46695a );
 a46697a <=( a46696a  and  a46691a );
 a46701a <=( (not A266)  and  (not A234) );
 a46702a <=( (not A233)  and  a46701a );
 a46705a <=( (not A269)  and  (not A268) );
 a46708a <=( (not A300)  and  A298 );
 a46709a <=( a46708a  and  a46705a );
 a46710a <=( a46709a  and  a46702a );
 a46714a <=( A167  and  (not A168) );
 a46715a <=( A169  and  a46714a );
 a46719a <=( A200  and  (not A199) );
 a46720a <=( (not A166)  and  a46719a );
 a46721a <=( a46720a  and  a46715a );
 a46725a <=( (not A266)  and  (not A234) );
 a46726a <=( (not A233)  and  a46725a );
 a46729a <=( (not A269)  and  (not A268) );
 a46732a <=( A299  and  A298 );
 a46733a <=( a46732a  and  a46729a );
 a46734a <=( a46733a  and  a46726a );
 a46738a <=( A167  and  (not A168) );
 a46739a <=( A169  and  a46738a );
 a46743a <=( A200  and  (not A199) );
 a46744a <=( (not A166)  and  a46743a );
 a46745a <=( a46744a  and  a46739a );
 a46749a <=( (not A266)  and  (not A234) );
 a46750a <=( (not A233)  and  a46749a );
 a46753a <=( (not A269)  and  (not A268) );
 a46756a <=( (not A299)  and  (not A298) );
 a46757a <=( a46756a  and  a46753a );
 a46758a <=( a46757a  and  a46750a );
 a46762a <=( A167  and  (not A168) );
 a46763a <=( A169  and  a46762a );
 a46767a <=( A200  and  (not A199) );
 a46768a <=( (not A166)  and  a46767a );
 a46769a <=( a46768a  and  a46763a );
 a46773a <=( (not A266)  and  (not A234) );
 a46774a <=( (not A233)  and  a46773a );
 a46777a <=( A298  and  (not A267) );
 a46780a <=( (not A302)  and  (not A301) );
 a46781a <=( a46780a  and  a46777a );
 a46782a <=( a46781a  and  a46774a );
 a46786a <=( A167  and  (not A168) );
 a46787a <=( A169  and  a46786a );
 a46791a <=( A200  and  (not A199) );
 a46792a <=( (not A166)  and  a46791a );
 a46793a <=( a46792a  and  a46787a );
 a46797a <=( (not A265)  and  (not A234) );
 a46798a <=( (not A233)  and  a46797a );
 a46801a <=( A298  and  (not A266) );
 a46804a <=( (not A302)  and  (not A301) );
 a46805a <=( a46804a  and  a46801a );
 a46806a <=( a46805a  and  a46798a );
 a46810a <=( A167  and  (not A168) );
 a46811a <=( A169  and  a46810a );
 a46815a <=( A200  and  (not A199) );
 a46816a <=( (not A166)  and  a46815a );
 a46817a <=( a46816a  and  a46811a );
 a46821a <=( A265  and  (not A233) );
 a46822a <=( (not A232)  and  a46821a );
 a46825a <=( A298  and  A266 );
 a46828a <=( (not A302)  and  (not A301) );
 a46829a <=( a46828a  and  a46825a );
 a46830a <=( a46829a  and  a46822a );
 a46834a <=( A167  and  (not A168) );
 a46835a <=( A169  and  a46834a );
 a46839a <=( A200  and  (not A199) );
 a46840a <=( (not A166)  and  a46839a );
 a46841a <=( a46840a  and  a46835a );
 a46845a <=( (not A266)  and  (not A233) );
 a46846a <=( (not A232)  and  a46845a );
 a46849a <=( (not A269)  and  (not A268) );
 a46852a <=( (not A300)  and  A298 );
 a46853a <=( a46852a  and  a46849a );
 a46854a <=( a46853a  and  a46846a );
 a46858a <=( A167  and  (not A168) );
 a46859a <=( A169  and  a46858a );
 a46863a <=( A200  and  (not A199) );
 a46864a <=( (not A166)  and  a46863a );
 a46865a <=( a46864a  and  a46859a );
 a46869a <=( (not A266)  and  (not A233) );
 a46870a <=( (not A232)  and  a46869a );
 a46873a <=( (not A269)  and  (not A268) );
 a46876a <=( A299  and  A298 );
 a46877a <=( a46876a  and  a46873a );
 a46878a <=( a46877a  and  a46870a );
 a46882a <=( A167  and  (not A168) );
 a46883a <=( A169  and  a46882a );
 a46887a <=( A200  and  (not A199) );
 a46888a <=( (not A166)  and  a46887a );
 a46889a <=( a46888a  and  a46883a );
 a46893a <=( (not A266)  and  (not A233) );
 a46894a <=( (not A232)  and  a46893a );
 a46897a <=( (not A269)  and  (not A268) );
 a46900a <=( (not A299)  and  (not A298) );
 a46901a <=( a46900a  and  a46897a );
 a46902a <=( a46901a  and  a46894a );
 a46906a <=( A167  and  (not A168) );
 a46907a <=( A169  and  a46906a );
 a46911a <=( A200  and  (not A199) );
 a46912a <=( (not A166)  and  a46911a );
 a46913a <=( a46912a  and  a46907a );
 a46917a <=( (not A266)  and  (not A233) );
 a46918a <=( (not A232)  and  a46917a );
 a46921a <=( A298  and  (not A267) );
 a46924a <=( (not A302)  and  (not A301) );
 a46925a <=( a46924a  and  a46921a );
 a46926a <=( a46925a  and  a46918a );
 a46930a <=( A167  and  (not A168) );
 a46931a <=( A169  and  a46930a );
 a46935a <=( A200  and  (not A199) );
 a46936a <=( (not A166)  and  a46935a );
 a46937a <=( a46936a  and  a46931a );
 a46941a <=( (not A265)  and  (not A233) );
 a46942a <=( (not A232)  and  a46941a );
 a46945a <=( A298  and  (not A266) );
 a46948a <=( (not A302)  and  (not A301) );
 a46949a <=( a46948a  and  a46945a );
 a46950a <=( a46949a  and  a46942a );
 a46954a <=( (not A167)  and  (not A168) );
 a46955a <=( A169  and  a46954a );
 a46959a <=( A200  and  (not A199) );
 a46960a <=( A166  and  a46959a );
 a46961a <=( a46960a  and  a46955a );
 a46965a <=( A265  and  A233 );
 a46966a <=( A232  and  a46965a );
 a46969a <=( (not A269)  and  (not A268) );
 a46972a <=( (not A300)  and  (not A299) );
 a46973a <=( a46972a  and  a46969a );
 a46974a <=( a46973a  and  a46966a );
 a46978a <=( (not A167)  and  (not A168) );
 a46979a <=( A169  and  a46978a );
 a46983a <=( A200  and  (not A199) );
 a46984a <=( A166  and  a46983a );
 a46985a <=( a46984a  and  a46979a );
 a46989a <=( A265  and  A233 );
 a46990a <=( A232  and  a46989a );
 a46993a <=( (not A269)  and  (not A268) );
 a46996a <=( A299  and  A298 );
 a46997a <=( a46996a  and  a46993a );
 a46998a <=( a46997a  and  a46990a );
 a47002a <=( (not A167)  and  (not A168) );
 a47003a <=( A169  and  a47002a );
 a47007a <=( A200  and  (not A199) );
 a47008a <=( A166  and  a47007a );
 a47009a <=( a47008a  and  a47003a );
 a47013a <=( A265  and  A233 );
 a47014a <=( A232  and  a47013a );
 a47017a <=( (not A269)  and  (not A268) );
 a47020a <=( (not A299)  and  (not A298) );
 a47021a <=( a47020a  and  a47017a );
 a47022a <=( a47021a  and  a47014a );
 a47026a <=( (not A167)  and  (not A168) );
 a47027a <=( A169  and  a47026a );
 a47031a <=( A200  and  (not A199) );
 a47032a <=( A166  and  a47031a );
 a47033a <=( a47032a  and  a47027a );
 a47037a <=( A265  and  A233 );
 a47038a <=( A232  and  a47037a );
 a47041a <=( (not A299)  and  (not A267) );
 a47044a <=( (not A302)  and  (not A301) );
 a47045a <=( a47044a  and  a47041a );
 a47046a <=( a47045a  and  a47038a );
 a47050a <=( (not A167)  and  (not A168) );
 a47051a <=( A169  and  a47050a );
 a47055a <=( A200  and  (not A199) );
 a47056a <=( A166  and  a47055a );
 a47057a <=( a47056a  and  a47051a );
 a47061a <=( A265  and  A233 );
 a47062a <=( A232  and  a47061a );
 a47065a <=( (not A299)  and  A266 );
 a47068a <=( (not A302)  and  (not A301) );
 a47069a <=( a47068a  and  a47065a );
 a47070a <=( a47069a  and  a47062a );
 a47074a <=( (not A167)  and  (not A168) );
 a47075a <=( A169  and  a47074a );
 a47079a <=( A200  and  (not A199) );
 a47080a <=( A166  and  a47079a );
 a47081a <=( a47080a  and  a47075a );
 a47085a <=( (not A265)  and  A233 );
 a47086a <=( A232  and  a47085a );
 a47089a <=( (not A299)  and  (not A266) );
 a47092a <=( (not A302)  and  (not A301) );
 a47093a <=( a47092a  and  a47089a );
 a47094a <=( a47093a  and  a47086a );
 a47098a <=( (not A167)  and  (not A168) );
 a47099a <=( A169  and  a47098a );
 a47103a <=( A200  and  (not A199) );
 a47104a <=( A166  and  a47103a );
 a47105a <=( a47104a  and  a47099a );
 a47109a <=( (not A236)  and  (not A235) );
 a47110a <=( (not A233)  and  a47109a );
 a47113a <=( A266  and  A265 );
 a47116a <=( (not A300)  and  A298 );
 a47117a <=( a47116a  and  a47113a );
 a47118a <=( a47117a  and  a47110a );
 a47122a <=( (not A167)  and  (not A168) );
 a47123a <=( A169  and  a47122a );
 a47127a <=( A200  and  (not A199) );
 a47128a <=( A166  and  a47127a );
 a47129a <=( a47128a  and  a47123a );
 a47133a <=( (not A236)  and  (not A235) );
 a47134a <=( (not A233)  and  a47133a );
 a47137a <=( A266  and  A265 );
 a47140a <=( A299  and  A298 );
 a47141a <=( a47140a  and  a47137a );
 a47142a <=( a47141a  and  a47134a );
 a47146a <=( (not A167)  and  (not A168) );
 a47147a <=( A169  and  a47146a );
 a47151a <=( A200  and  (not A199) );
 a47152a <=( A166  and  a47151a );
 a47153a <=( a47152a  and  a47147a );
 a47157a <=( (not A236)  and  (not A235) );
 a47158a <=( (not A233)  and  a47157a );
 a47161a <=( A266  and  A265 );
 a47164a <=( (not A299)  and  (not A298) );
 a47165a <=( a47164a  and  a47161a );
 a47166a <=( a47165a  and  a47158a );
 a47170a <=( (not A167)  and  (not A168) );
 a47171a <=( A169  and  a47170a );
 a47175a <=( A200  and  (not A199) );
 a47176a <=( A166  and  a47175a );
 a47177a <=( a47176a  and  a47171a );
 a47181a <=( (not A236)  and  (not A235) );
 a47182a <=( (not A233)  and  a47181a );
 a47185a <=( (not A267)  and  (not A266) );
 a47188a <=( (not A300)  and  A298 );
 a47189a <=( a47188a  and  a47185a );
 a47190a <=( a47189a  and  a47182a );
 a47194a <=( (not A167)  and  (not A168) );
 a47195a <=( A169  and  a47194a );
 a47199a <=( A200  and  (not A199) );
 a47200a <=( A166  and  a47199a );
 a47201a <=( a47200a  and  a47195a );
 a47205a <=( (not A236)  and  (not A235) );
 a47206a <=( (not A233)  and  a47205a );
 a47209a <=( (not A267)  and  (not A266) );
 a47212a <=( A299  and  A298 );
 a47213a <=( a47212a  and  a47209a );
 a47214a <=( a47213a  and  a47206a );
 a47218a <=( (not A167)  and  (not A168) );
 a47219a <=( A169  and  a47218a );
 a47223a <=( A200  and  (not A199) );
 a47224a <=( A166  and  a47223a );
 a47225a <=( a47224a  and  a47219a );
 a47229a <=( (not A236)  and  (not A235) );
 a47230a <=( (not A233)  and  a47229a );
 a47233a <=( (not A267)  and  (not A266) );
 a47236a <=( (not A299)  and  (not A298) );
 a47237a <=( a47236a  and  a47233a );
 a47238a <=( a47237a  and  a47230a );
 a47242a <=( (not A167)  and  (not A168) );
 a47243a <=( A169  and  a47242a );
 a47247a <=( A200  and  (not A199) );
 a47248a <=( A166  and  a47247a );
 a47249a <=( a47248a  and  a47243a );
 a47253a <=( (not A236)  and  (not A235) );
 a47254a <=( (not A233)  and  a47253a );
 a47257a <=( (not A266)  and  (not A265) );
 a47260a <=( (not A300)  and  A298 );
 a47261a <=( a47260a  and  a47257a );
 a47262a <=( a47261a  and  a47254a );
 a47266a <=( (not A167)  and  (not A168) );
 a47267a <=( A169  and  a47266a );
 a47271a <=( A200  and  (not A199) );
 a47272a <=( A166  and  a47271a );
 a47273a <=( a47272a  and  a47267a );
 a47277a <=( (not A236)  and  (not A235) );
 a47278a <=( (not A233)  and  a47277a );
 a47281a <=( (not A266)  and  (not A265) );
 a47284a <=( A299  and  A298 );
 a47285a <=( a47284a  and  a47281a );
 a47286a <=( a47285a  and  a47278a );
 a47290a <=( (not A167)  and  (not A168) );
 a47291a <=( A169  and  a47290a );
 a47295a <=( A200  and  (not A199) );
 a47296a <=( A166  and  a47295a );
 a47297a <=( a47296a  and  a47291a );
 a47301a <=( (not A236)  and  (not A235) );
 a47302a <=( (not A233)  and  a47301a );
 a47305a <=( (not A266)  and  (not A265) );
 a47308a <=( (not A299)  and  (not A298) );
 a47309a <=( a47308a  and  a47305a );
 a47310a <=( a47309a  and  a47302a );
 a47314a <=( (not A167)  and  (not A168) );
 a47315a <=( A169  and  a47314a );
 a47319a <=( A200  and  (not A199) );
 a47320a <=( A166  and  a47319a );
 a47321a <=( a47320a  and  a47315a );
 a47325a <=( A265  and  (not A234) );
 a47326a <=( (not A233)  and  a47325a );
 a47329a <=( A298  and  A266 );
 a47332a <=( (not A302)  and  (not A301) );
 a47333a <=( a47332a  and  a47329a );
 a47334a <=( a47333a  and  a47326a );
 a47338a <=( (not A167)  and  (not A168) );
 a47339a <=( A169  and  a47338a );
 a47343a <=( A200  and  (not A199) );
 a47344a <=( A166  and  a47343a );
 a47345a <=( a47344a  and  a47339a );
 a47349a <=( (not A266)  and  (not A234) );
 a47350a <=( (not A233)  and  a47349a );
 a47353a <=( (not A269)  and  (not A268) );
 a47356a <=( (not A300)  and  A298 );
 a47357a <=( a47356a  and  a47353a );
 a47358a <=( a47357a  and  a47350a );
 a47362a <=( (not A167)  and  (not A168) );
 a47363a <=( A169  and  a47362a );
 a47367a <=( A200  and  (not A199) );
 a47368a <=( A166  and  a47367a );
 a47369a <=( a47368a  and  a47363a );
 a47373a <=( (not A266)  and  (not A234) );
 a47374a <=( (not A233)  and  a47373a );
 a47377a <=( (not A269)  and  (not A268) );
 a47380a <=( A299  and  A298 );
 a47381a <=( a47380a  and  a47377a );
 a47382a <=( a47381a  and  a47374a );
 a47386a <=( (not A167)  and  (not A168) );
 a47387a <=( A169  and  a47386a );
 a47391a <=( A200  and  (not A199) );
 a47392a <=( A166  and  a47391a );
 a47393a <=( a47392a  and  a47387a );
 a47397a <=( (not A266)  and  (not A234) );
 a47398a <=( (not A233)  and  a47397a );
 a47401a <=( (not A269)  and  (not A268) );
 a47404a <=( (not A299)  and  (not A298) );
 a47405a <=( a47404a  and  a47401a );
 a47406a <=( a47405a  and  a47398a );
 a47410a <=( (not A167)  and  (not A168) );
 a47411a <=( A169  and  a47410a );
 a47415a <=( A200  and  (not A199) );
 a47416a <=( A166  and  a47415a );
 a47417a <=( a47416a  and  a47411a );
 a47421a <=( (not A266)  and  (not A234) );
 a47422a <=( (not A233)  and  a47421a );
 a47425a <=( A298  and  (not A267) );
 a47428a <=( (not A302)  and  (not A301) );
 a47429a <=( a47428a  and  a47425a );
 a47430a <=( a47429a  and  a47422a );
 a47434a <=( (not A167)  and  (not A168) );
 a47435a <=( A169  and  a47434a );
 a47439a <=( A200  and  (not A199) );
 a47440a <=( A166  and  a47439a );
 a47441a <=( a47440a  and  a47435a );
 a47445a <=( (not A265)  and  (not A234) );
 a47446a <=( (not A233)  and  a47445a );
 a47449a <=( A298  and  (not A266) );
 a47452a <=( (not A302)  and  (not A301) );
 a47453a <=( a47452a  and  a47449a );
 a47454a <=( a47453a  and  a47446a );
 a47458a <=( (not A167)  and  (not A168) );
 a47459a <=( A169  and  a47458a );
 a47463a <=( A200  and  (not A199) );
 a47464a <=( A166  and  a47463a );
 a47465a <=( a47464a  and  a47459a );
 a47469a <=( A265  and  (not A233) );
 a47470a <=( (not A232)  and  a47469a );
 a47473a <=( A298  and  A266 );
 a47476a <=( (not A302)  and  (not A301) );
 a47477a <=( a47476a  and  a47473a );
 a47478a <=( a47477a  and  a47470a );
 a47482a <=( (not A167)  and  (not A168) );
 a47483a <=( A169  and  a47482a );
 a47487a <=( A200  and  (not A199) );
 a47488a <=( A166  and  a47487a );
 a47489a <=( a47488a  and  a47483a );
 a47493a <=( (not A266)  and  (not A233) );
 a47494a <=( (not A232)  and  a47493a );
 a47497a <=( (not A269)  and  (not A268) );
 a47500a <=( (not A300)  and  A298 );
 a47501a <=( a47500a  and  a47497a );
 a47502a <=( a47501a  and  a47494a );
 a47506a <=( (not A167)  and  (not A168) );
 a47507a <=( A169  and  a47506a );
 a47511a <=( A200  and  (not A199) );
 a47512a <=( A166  and  a47511a );
 a47513a <=( a47512a  and  a47507a );
 a47517a <=( (not A266)  and  (not A233) );
 a47518a <=( (not A232)  and  a47517a );
 a47521a <=( (not A269)  and  (not A268) );
 a47524a <=( A299  and  A298 );
 a47525a <=( a47524a  and  a47521a );
 a47526a <=( a47525a  and  a47518a );
 a47530a <=( (not A167)  and  (not A168) );
 a47531a <=( A169  and  a47530a );
 a47535a <=( A200  and  (not A199) );
 a47536a <=( A166  and  a47535a );
 a47537a <=( a47536a  and  a47531a );
 a47541a <=( (not A266)  and  (not A233) );
 a47542a <=( (not A232)  and  a47541a );
 a47545a <=( (not A269)  and  (not A268) );
 a47548a <=( (not A299)  and  (not A298) );
 a47549a <=( a47548a  and  a47545a );
 a47550a <=( a47549a  and  a47542a );
 a47554a <=( (not A167)  and  (not A168) );
 a47555a <=( A169  and  a47554a );
 a47559a <=( A200  and  (not A199) );
 a47560a <=( A166  and  a47559a );
 a47561a <=( a47560a  and  a47555a );
 a47565a <=( (not A266)  and  (not A233) );
 a47566a <=( (not A232)  and  a47565a );
 a47569a <=( A298  and  (not A267) );
 a47572a <=( (not A302)  and  (not A301) );
 a47573a <=( a47572a  and  a47569a );
 a47574a <=( a47573a  and  a47566a );
 a47578a <=( (not A167)  and  (not A168) );
 a47579a <=( A169  and  a47578a );
 a47583a <=( A200  and  (not A199) );
 a47584a <=( A166  and  a47583a );
 a47585a <=( a47584a  and  a47579a );
 a47589a <=( (not A265)  and  (not A233) );
 a47590a <=( (not A232)  and  a47589a );
 a47593a <=( A298  and  (not A266) );
 a47596a <=( (not A302)  and  (not A301) );
 a47597a <=( a47596a  and  a47593a );
 a47598a <=( a47597a  and  a47590a );
 a47602a <=( (not A168)  and  A169 );
 a47603a <=( A170  and  a47602a );
 a47607a <=( A201  and  (not A200) );
 a47608a <=( A199  and  a47607a );
 a47609a <=( a47608a  and  a47603a );
 a47613a <=( A233  and  A232 );
 a47614a <=( A202  and  a47613a );
 a47617a <=( (not A267)  and  A265 );
 a47620a <=( (not A300)  and  (not A299) );
 a47621a <=( a47620a  and  a47617a );
 a47622a <=( a47621a  and  a47614a );
 a47626a <=( (not A168)  and  A169 );
 a47627a <=( A170  and  a47626a );
 a47631a <=( A201  and  (not A200) );
 a47632a <=( A199  and  a47631a );
 a47633a <=( a47632a  and  a47627a );
 a47637a <=( A233  and  A232 );
 a47638a <=( A202  and  a47637a );
 a47641a <=( (not A267)  and  A265 );
 a47644a <=( A299  and  A298 );
 a47645a <=( a47644a  and  a47641a );
 a47646a <=( a47645a  and  a47638a );
 a47650a <=( (not A168)  and  A169 );
 a47651a <=( A170  and  a47650a );
 a47655a <=( A201  and  (not A200) );
 a47656a <=( A199  and  a47655a );
 a47657a <=( a47656a  and  a47651a );
 a47661a <=( A233  and  A232 );
 a47662a <=( A202  and  a47661a );
 a47665a <=( (not A267)  and  A265 );
 a47668a <=( (not A299)  and  (not A298) );
 a47669a <=( a47668a  and  a47665a );
 a47670a <=( a47669a  and  a47662a );
 a47674a <=( (not A168)  and  A169 );
 a47675a <=( A170  and  a47674a );
 a47679a <=( A201  and  (not A200) );
 a47680a <=( A199  and  a47679a );
 a47681a <=( a47680a  and  a47675a );
 a47685a <=( A233  and  A232 );
 a47686a <=( A202  and  a47685a );
 a47689a <=( A266  and  A265 );
 a47692a <=( (not A300)  and  (not A299) );
 a47693a <=( a47692a  and  a47689a );
 a47694a <=( a47693a  and  a47686a );
 a47698a <=( (not A168)  and  A169 );
 a47699a <=( A170  and  a47698a );
 a47703a <=( A201  and  (not A200) );
 a47704a <=( A199  and  a47703a );
 a47705a <=( a47704a  and  a47699a );
 a47709a <=( A233  and  A232 );
 a47710a <=( A202  and  a47709a );
 a47713a <=( A266  and  A265 );
 a47716a <=( A299  and  A298 );
 a47717a <=( a47716a  and  a47713a );
 a47718a <=( a47717a  and  a47710a );
 a47722a <=( (not A168)  and  A169 );
 a47723a <=( A170  and  a47722a );
 a47727a <=( A201  and  (not A200) );
 a47728a <=( A199  and  a47727a );
 a47729a <=( a47728a  and  a47723a );
 a47733a <=( A233  and  A232 );
 a47734a <=( A202  and  a47733a );
 a47737a <=( A266  and  A265 );
 a47740a <=( (not A299)  and  (not A298) );
 a47741a <=( a47740a  and  a47737a );
 a47742a <=( a47741a  and  a47734a );
 a47746a <=( (not A168)  and  A169 );
 a47747a <=( A170  and  a47746a );
 a47751a <=( A201  and  (not A200) );
 a47752a <=( A199  and  a47751a );
 a47753a <=( a47752a  and  a47747a );
 a47757a <=( A233  and  A232 );
 a47758a <=( A202  and  a47757a );
 a47761a <=( (not A266)  and  (not A265) );
 a47764a <=( (not A300)  and  (not A299) );
 a47765a <=( a47764a  and  a47761a );
 a47766a <=( a47765a  and  a47758a );
 a47770a <=( (not A168)  and  A169 );
 a47771a <=( A170  and  a47770a );
 a47775a <=( A201  and  (not A200) );
 a47776a <=( A199  and  a47775a );
 a47777a <=( a47776a  and  a47771a );
 a47781a <=( A233  and  A232 );
 a47782a <=( A202  and  a47781a );
 a47785a <=( (not A266)  and  (not A265) );
 a47788a <=( A299  and  A298 );
 a47789a <=( a47788a  and  a47785a );
 a47790a <=( a47789a  and  a47782a );
 a47794a <=( (not A168)  and  A169 );
 a47795a <=( A170  and  a47794a );
 a47799a <=( A201  and  (not A200) );
 a47800a <=( A199  and  a47799a );
 a47801a <=( a47800a  and  a47795a );
 a47805a <=( A233  and  A232 );
 a47806a <=( A202  and  a47805a );
 a47809a <=( (not A266)  and  (not A265) );
 a47812a <=( (not A299)  and  (not A298) );
 a47813a <=( a47812a  and  a47809a );
 a47814a <=( a47813a  and  a47806a );
 a47818a <=( (not A168)  and  A169 );
 a47819a <=( A170  and  a47818a );
 a47823a <=( A201  and  (not A200) );
 a47824a <=( A199  and  a47823a );
 a47825a <=( a47824a  and  a47819a );
 a47829a <=( (not A234)  and  (not A233) );
 a47830a <=( A202  and  a47829a );
 a47833a <=( A266  and  A265 );
 a47836a <=( (not A300)  and  A298 );
 a47837a <=( a47836a  and  a47833a );
 a47838a <=( a47837a  and  a47830a );
 a47842a <=( (not A168)  and  A169 );
 a47843a <=( A170  and  a47842a );
 a47847a <=( A201  and  (not A200) );
 a47848a <=( A199  and  a47847a );
 a47849a <=( a47848a  and  a47843a );
 a47853a <=( (not A234)  and  (not A233) );
 a47854a <=( A202  and  a47853a );
 a47857a <=( A266  and  A265 );
 a47860a <=( A299  and  A298 );
 a47861a <=( a47860a  and  a47857a );
 a47862a <=( a47861a  and  a47854a );
 a47866a <=( (not A168)  and  A169 );
 a47867a <=( A170  and  a47866a );
 a47871a <=( A201  and  (not A200) );
 a47872a <=( A199  and  a47871a );
 a47873a <=( a47872a  and  a47867a );
 a47877a <=( (not A234)  and  (not A233) );
 a47878a <=( A202  and  a47877a );
 a47881a <=( A266  and  A265 );
 a47884a <=( (not A299)  and  (not A298) );
 a47885a <=( a47884a  and  a47881a );
 a47886a <=( a47885a  and  a47878a );
 a47890a <=( (not A168)  and  A169 );
 a47891a <=( A170  and  a47890a );
 a47895a <=( A201  and  (not A200) );
 a47896a <=( A199  and  a47895a );
 a47897a <=( a47896a  and  a47891a );
 a47901a <=( (not A234)  and  (not A233) );
 a47902a <=( A202  and  a47901a );
 a47905a <=( (not A267)  and  (not A266) );
 a47908a <=( (not A300)  and  A298 );
 a47909a <=( a47908a  and  a47905a );
 a47910a <=( a47909a  and  a47902a );
 a47914a <=( (not A168)  and  A169 );
 a47915a <=( A170  and  a47914a );
 a47919a <=( A201  and  (not A200) );
 a47920a <=( A199  and  a47919a );
 a47921a <=( a47920a  and  a47915a );
 a47925a <=( (not A234)  and  (not A233) );
 a47926a <=( A202  and  a47925a );
 a47929a <=( (not A267)  and  (not A266) );
 a47932a <=( A299  and  A298 );
 a47933a <=( a47932a  and  a47929a );
 a47934a <=( a47933a  and  a47926a );
 a47938a <=( (not A168)  and  A169 );
 a47939a <=( A170  and  a47938a );
 a47943a <=( A201  and  (not A200) );
 a47944a <=( A199  and  a47943a );
 a47945a <=( a47944a  and  a47939a );
 a47949a <=( (not A234)  and  (not A233) );
 a47950a <=( A202  and  a47949a );
 a47953a <=( (not A267)  and  (not A266) );
 a47956a <=( (not A299)  and  (not A298) );
 a47957a <=( a47956a  and  a47953a );
 a47958a <=( a47957a  and  a47950a );
 a47962a <=( (not A168)  and  A169 );
 a47963a <=( A170  and  a47962a );
 a47967a <=( A201  and  (not A200) );
 a47968a <=( A199  and  a47967a );
 a47969a <=( a47968a  and  a47963a );
 a47973a <=( (not A234)  and  (not A233) );
 a47974a <=( A202  and  a47973a );
 a47977a <=( (not A266)  and  (not A265) );
 a47980a <=( (not A300)  and  A298 );
 a47981a <=( a47980a  and  a47977a );
 a47982a <=( a47981a  and  a47974a );
 a47986a <=( (not A168)  and  A169 );
 a47987a <=( A170  and  a47986a );
 a47991a <=( A201  and  (not A200) );
 a47992a <=( A199  and  a47991a );
 a47993a <=( a47992a  and  a47987a );
 a47997a <=( (not A234)  and  (not A233) );
 a47998a <=( A202  and  a47997a );
 a48001a <=( (not A266)  and  (not A265) );
 a48004a <=( A299  and  A298 );
 a48005a <=( a48004a  and  a48001a );
 a48006a <=( a48005a  and  a47998a );
 a48010a <=( (not A168)  and  A169 );
 a48011a <=( A170  and  a48010a );
 a48015a <=( A201  and  (not A200) );
 a48016a <=( A199  and  a48015a );
 a48017a <=( a48016a  and  a48011a );
 a48021a <=( (not A234)  and  (not A233) );
 a48022a <=( A202  and  a48021a );
 a48025a <=( (not A266)  and  (not A265) );
 a48028a <=( (not A299)  and  (not A298) );
 a48029a <=( a48028a  and  a48025a );
 a48030a <=( a48029a  and  a48022a );
 a48034a <=( (not A168)  and  A169 );
 a48035a <=( A170  and  a48034a );
 a48039a <=( A201  and  (not A200) );
 a48040a <=( A199  and  a48039a );
 a48041a <=( a48040a  and  a48035a );
 a48045a <=( (not A233)  and  A232 );
 a48046a <=( A202  and  a48045a );
 a48049a <=( A235  and  A234 );
 a48052a <=( A299  and  (not A298) );
 a48053a <=( a48052a  and  a48049a );
 a48054a <=( a48053a  and  a48046a );
 a48058a <=( (not A168)  and  A169 );
 a48059a <=( A170  and  a48058a );
 a48063a <=( A201  and  (not A200) );
 a48064a <=( A199  and  a48063a );
 a48065a <=( a48064a  and  a48059a );
 a48069a <=( (not A233)  and  A232 );
 a48070a <=( A202  and  a48069a );
 a48073a <=( A235  and  A234 );
 a48076a <=( A266  and  (not A265) );
 a48077a <=( a48076a  and  a48073a );
 a48078a <=( a48077a  and  a48070a );
 a48082a <=( (not A168)  and  A169 );
 a48083a <=( A170  and  a48082a );
 a48087a <=( A201  and  (not A200) );
 a48088a <=( A199  and  a48087a );
 a48089a <=( a48088a  and  a48083a );
 a48093a <=( (not A233)  and  A232 );
 a48094a <=( A202  and  a48093a );
 a48097a <=( A236  and  A234 );
 a48100a <=( A299  and  (not A298) );
 a48101a <=( a48100a  and  a48097a );
 a48102a <=( a48101a  and  a48094a );
 a48106a <=( (not A168)  and  A169 );
 a48107a <=( A170  and  a48106a );
 a48111a <=( A201  and  (not A200) );
 a48112a <=( A199  and  a48111a );
 a48113a <=( a48112a  and  a48107a );
 a48117a <=( (not A233)  and  A232 );
 a48118a <=( A202  and  a48117a );
 a48121a <=( A236  and  A234 );
 a48124a <=( A266  and  (not A265) );
 a48125a <=( a48124a  and  a48121a );
 a48126a <=( a48125a  and  a48118a );
 a48130a <=( (not A168)  and  A169 );
 a48131a <=( A170  and  a48130a );
 a48135a <=( A201  and  (not A200) );
 a48136a <=( A199  and  a48135a );
 a48137a <=( a48136a  and  a48131a );
 a48141a <=( (not A233)  and  (not A232) );
 a48142a <=( A202  and  a48141a );
 a48145a <=( A266  and  A265 );
 a48148a <=( (not A300)  and  A298 );
 a48149a <=( a48148a  and  a48145a );
 a48150a <=( a48149a  and  a48142a );
 a48154a <=( (not A168)  and  A169 );
 a48155a <=( A170  and  a48154a );
 a48159a <=( A201  and  (not A200) );
 a48160a <=( A199  and  a48159a );
 a48161a <=( a48160a  and  a48155a );
 a48165a <=( (not A233)  and  (not A232) );
 a48166a <=( A202  and  a48165a );
 a48169a <=( A266  and  A265 );
 a48172a <=( A299  and  A298 );
 a48173a <=( a48172a  and  a48169a );
 a48174a <=( a48173a  and  a48166a );
 a48178a <=( (not A168)  and  A169 );
 a48179a <=( A170  and  a48178a );
 a48183a <=( A201  and  (not A200) );
 a48184a <=( A199  and  a48183a );
 a48185a <=( a48184a  and  a48179a );
 a48189a <=( (not A233)  and  (not A232) );
 a48190a <=( A202  and  a48189a );
 a48193a <=( A266  and  A265 );
 a48196a <=( (not A299)  and  (not A298) );
 a48197a <=( a48196a  and  a48193a );
 a48198a <=( a48197a  and  a48190a );
 a48202a <=( (not A168)  and  A169 );
 a48203a <=( A170  and  a48202a );
 a48207a <=( A201  and  (not A200) );
 a48208a <=( A199  and  a48207a );
 a48209a <=( a48208a  and  a48203a );
 a48213a <=( (not A233)  and  (not A232) );
 a48214a <=( A202  and  a48213a );
 a48217a <=( (not A267)  and  (not A266) );
 a48220a <=( (not A300)  and  A298 );
 a48221a <=( a48220a  and  a48217a );
 a48222a <=( a48221a  and  a48214a );
 a48226a <=( (not A168)  and  A169 );
 a48227a <=( A170  and  a48226a );
 a48231a <=( A201  and  (not A200) );
 a48232a <=( A199  and  a48231a );
 a48233a <=( a48232a  and  a48227a );
 a48237a <=( (not A233)  and  (not A232) );
 a48238a <=( A202  and  a48237a );
 a48241a <=( (not A267)  and  (not A266) );
 a48244a <=( A299  and  A298 );
 a48245a <=( a48244a  and  a48241a );
 a48246a <=( a48245a  and  a48238a );
 a48250a <=( (not A168)  and  A169 );
 a48251a <=( A170  and  a48250a );
 a48255a <=( A201  and  (not A200) );
 a48256a <=( A199  and  a48255a );
 a48257a <=( a48256a  and  a48251a );
 a48261a <=( (not A233)  and  (not A232) );
 a48262a <=( A202  and  a48261a );
 a48265a <=( (not A267)  and  (not A266) );
 a48268a <=( (not A299)  and  (not A298) );
 a48269a <=( a48268a  and  a48265a );
 a48270a <=( a48269a  and  a48262a );
 a48274a <=( (not A168)  and  A169 );
 a48275a <=( A170  and  a48274a );
 a48279a <=( A201  and  (not A200) );
 a48280a <=( A199  and  a48279a );
 a48281a <=( a48280a  and  a48275a );
 a48285a <=( (not A233)  and  (not A232) );
 a48286a <=( A202  and  a48285a );
 a48289a <=( (not A266)  and  (not A265) );
 a48292a <=( (not A300)  and  A298 );
 a48293a <=( a48292a  and  a48289a );
 a48294a <=( a48293a  and  a48286a );
 a48298a <=( (not A168)  and  A169 );
 a48299a <=( A170  and  a48298a );
 a48303a <=( A201  and  (not A200) );
 a48304a <=( A199  and  a48303a );
 a48305a <=( a48304a  and  a48299a );
 a48309a <=( (not A233)  and  (not A232) );
 a48310a <=( A202  and  a48309a );
 a48313a <=( (not A266)  and  (not A265) );
 a48316a <=( A299  and  A298 );
 a48317a <=( a48316a  and  a48313a );
 a48318a <=( a48317a  and  a48310a );
 a48322a <=( (not A168)  and  A169 );
 a48323a <=( A170  and  a48322a );
 a48327a <=( A201  and  (not A200) );
 a48328a <=( A199  and  a48327a );
 a48329a <=( a48328a  and  a48323a );
 a48333a <=( (not A233)  and  (not A232) );
 a48334a <=( A202  and  a48333a );
 a48337a <=( (not A266)  and  (not A265) );
 a48340a <=( (not A299)  and  (not A298) );
 a48341a <=( a48340a  and  a48337a );
 a48342a <=( a48341a  and  a48334a );
 a48346a <=( (not A168)  and  A169 );
 a48347a <=( A170  and  a48346a );
 a48351a <=( A201  and  (not A200) );
 a48352a <=( A199  and  a48351a );
 a48353a <=( a48352a  and  a48347a );
 a48357a <=( A233  and  A232 );
 a48358a <=( A203  and  a48357a );
 a48361a <=( (not A267)  and  A265 );
 a48364a <=( (not A300)  and  (not A299) );
 a48365a <=( a48364a  and  a48361a );
 a48366a <=( a48365a  and  a48358a );
 a48370a <=( (not A168)  and  A169 );
 a48371a <=( A170  and  a48370a );
 a48375a <=( A201  and  (not A200) );
 a48376a <=( A199  and  a48375a );
 a48377a <=( a48376a  and  a48371a );
 a48381a <=( A233  and  A232 );
 a48382a <=( A203  and  a48381a );
 a48385a <=( (not A267)  and  A265 );
 a48388a <=( A299  and  A298 );
 a48389a <=( a48388a  and  a48385a );
 a48390a <=( a48389a  and  a48382a );
 a48394a <=( (not A168)  and  A169 );
 a48395a <=( A170  and  a48394a );
 a48399a <=( A201  and  (not A200) );
 a48400a <=( A199  and  a48399a );
 a48401a <=( a48400a  and  a48395a );
 a48405a <=( A233  and  A232 );
 a48406a <=( A203  and  a48405a );
 a48409a <=( (not A267)  and  A265 );
 a48412a <=( (not A299)  and  (not A298) );
 a48413a <=( a48412a  and  a48409a );
 a48414a <=( a48413a  and  a48406a );
 a48418a <=( (not A168)  and  A169 );
 a48419a <=( A170  and  a48418a );
 a48423a <=( A201  and  (not A200) );
 a48424a <=( A199  and  a48423a );
 a48425a <=( a48424a  and  a48419a );
 a48429a <=( A233  and  A232 );
 a48430a <=( A203  and  a48429a );
 a48433a <=( A266  and  A265 );
 a48436a <=( (not A300)  and  (not A299) );
 a48437a <=( a48436a  and  a48433a );
 a48438a <=( a48437a  and  a48430a );
 a48442a <=( (not A168)  and  A169 );
 a48443a <=( A170  and  a48442a );
 a48447a <=( A201  and  (not A200) );
 a48448a <=( A199  and  a48447a );
 a48449a <=( a48448a  and  a48443a );
 a48453a <=( A233  and  A232 );
 a48454a <=( A203  and  a48453a );
 a48457a <=( A266  and  A265 );
 a48460a <=( A299  and  A298 );
 a48461a <=( a48460a  and  a48457a );
 a48462a <=( a48461a  and  a48454a );
 a48466a <=( (not A168)  and  A169 );
 a48467a <=( A170  and  a48466a );
 a48471a <=( A201  and  (not A200) );
 a48472a <=( A199  and  a48471a );
 a48473a <=( a48472a  and  a48467a );
 a48477a <=( A233  and  A232 );
 a48478a <=( A203  and  a48477a );
 a48481a <=( A266  and  A265 );
 a48484a <=( (not A299)  and  (not A298) );
 a48485a <=( a48484a  and  a48481a );
 a48486a <=( a48485a  and  a48478a );
 a48490a <=( (not A168)  and  A169 );
 a48491a <=( A170  and  a48490a );
 a48495a <=( A201  and  (not A200) );
 a48496a <=( A199  and  a48495a );
 a48497a <=( a48496a  and  a48491a );
 a48501a <=( A233  and  A232 );
 a48502a <=( A203  and  a48501a );
 a48505a <=( (not A266)  and  (not A265) );
 a48508a <=( (not A300)  and  (not A299) );
 a48509a <=( a48508a  and  a48505a );
 a48510a <=( a48509a  and  a48502a );
 a48514a <=( (not A168)  and  A169 );
 a48515a <=( A170  and  a48514a );
 a48519a <=( A201  and  (not A200) );
 a48520a <=( A199  and  a48519a );
 a48521a <=( a48520a  and  a48515a );
 a48525a <=( A233  and  A232 );
 a48526a <=( A203  and  a48525a );
 a48529a <=( (not A266)  and  (not A265) );
 a48532a <=( A299  and  A298 );
 a48533a <=( a48532a  and  a48529a );
 a48534a <=( a48533a  and  a48526a );
 a48538a <=( (not A168)  and  A169 );
 a48539a <=( A170  and  a48538a );
 a48543a <=( A201  and  (not A200) );
 a48544a <=( A199  and  a48543a );
 a48545a <=( a48544a  and  a48539a );
 a48549a <=( A233  and  A232 );
 a48550a <=( A203  and  a48549a );
 a48553a <=( (not A266)  and  (not A265) );
 a48556a <=( (not A299)  and  (not A298) );
 a48557a <=( a48556a  and  a48553a );
 a48558a <=( a48557a  and  a48550a );
 a48562a <=( (not A168)  and  A169 );
 a48563a <=( A170  and  a48562a );
 a48567a <=( A201  and  (not A200) );
 a48568a <=( A199  and  a48567a );
 a48569a <=( a48568a  and  a48563a );
 a48573a <=( (not A234)  and  (not A233) );
 a48574a <=( A203  and  a48573a );
 a48577a <=( A266  and  A265 );
 a48580a <=( (not A300)  and  A298 );
 a48581a <=( a48580a  and  a48577a );
 a48582a <=( a48581a  and  a48574a );
 a48586a <=( (not A168)  and  A169 );
 a48587a <=( A170  and  a48586a );
 a48591a <=( A201  and  (not A200) );
 a48592a <=( A199  and  a48591a );
 a48593a <=( a48592a  and  a48587a );
 a48597a <=( (not A234)  and  (not A233) );
 a48598a <=( A203  and  a48597a );
 a48601a <=( A266  and  A265 );
 a48604a <=( A299  and  A298 );
 a48605a <=( a48604a  and  a48601a );
 a48606a <=( a48605a  and  a48598a );
 a48610a <=( (not A168)  and  A169 );
 a48611a <=( A170  and  a48610a );
 a48615a <=( A201  and  (not A200) );
 a48616a <=( A199  and  a48615a );
 a48617a <=( a48616a  and  a48611a );
 a48621a <=( (not A234)  and  (not A233) );
 a48622a <=( A203  and  a48621a );
 a48625a <=( A266  and  A265 );
 a48628a <=( (not A299)  and  (not A298) );
 a48629a <=( a48628a  and  a48625a );
 a48630a <=( a48629a  and  a48622a );
 a48634a <=( (not A168)  and  A169 );
 a48635a <=( A170  and  a48634a );
 a48639a <=( A201  and  (not A200) );
 a48640a <=( A199  and  a48639a );
 a48641a <=( a48640a  and  a48635a );
 a48645a <=( (not A234)  and  (not A233) );
 a48646a <=( A203  and  a48645a );
 a48649a <=( (not A267)  and  (not A266) );
 a48652a <=( (not A300)  and  A298 );
 a48653a <=( a48652a  and  a48649a );
 a48654a <=( a48653a  and  a48646a );
 a48658a <=( (not A168)  and  A169 );
 a48659a <=( A170  and  a48658a );
 a48663a <=( A201  and  (not A200) );
 a48664a <=( A199  and  a48663a );
 a48665a <=( a48664a  and  a48659a );
 a48669a <=( (not A234)  and  (not A233) );
 a48670a <=( A203  and  a48669a );
 a48673a <=( (not A267)  and  (not A266) );
 a48676a <=( A299  and  A298 );
 a48677a <=( a48676a  and  a48673a );
 a48678a <=( a48677a  and  a48670a );
 a48682a <=( (not A168)  and  A169 );
 a48683a <=( A170  and  a48682a );
 a48687a <=( A201  and  (not A200) );
 a48688a <=( A199  and  a48687a );
 a48689a <=( a48688a  and  a48683a );
 a48693a <=( (not A234)  and  (not A233) );
 a48694a <=( A203  and  a48693a );
 a48697a <=( (not A267)  and  (not A266) );
 a48700a <=( (not A299)  and  (not A298) );
 a48701a <=( a48700a  and  a48697a );
 a48702a <=( a48701a  and  a48694a );
 a48706a <=( (not A168)  and  A169 );
 a48707a <=( A170  and  a48706a );
 a48711a <=( A201  and  (not A200) );
 a48712a <=( A199  and  a48711a );
 a48713a <=( a48712a  and  a48707a );
 a48717a <=( (not A234)  and  (not A233) );
 a48718a <=( A203  and  a48717a );
 a48721a <=( (not A266)  and  (not A265) );
 a48724a <=( (not A300)  and  A298 );
 a48725a <=( a48724a  and  a48721a );
 a48726a <=( a48725a  and  a48718a );
 a48730a <=( (not A168)  and  A169 );
 a48731a <=( A170  and  a48730a );
 a48735a <=( A201  and  (not A200) );
 a48736a <=( A199  and  a48735a );
 a48737a <=( a48736a  and  a48731a );
 a48741a <=( (not A234)  and  (not A233) );
 a48742a <=( A203  and  a48741a );
 a48745a <=( (not A266)  and  (not A265) );
 a48748a <=( A299  and  A298 );
 a48749a <=( a48748a  and  a48745a );
 a48750a <=( a48749a  and  a48742a );
 a48754a <=( (not A168)  and  A169 );
 a48755a <=( A170  and  a48754a );
 a48759a <=( A201  and  (not A200) );
 a48760a <=( A199  and  a48759a );
 a48761a <=( a48760a  and  a48755a );
 a48765a <=( (not A234)  and  (not A233) );
 a48766a <=( A203  and  a48765a );
 a48769a <=( (not A266)  and  (not A265) );
 a48772a <=( (not A299)  and  (not A298) );
 a48773a <=( a48772a  and  a48769a );
 a48774a <=( a48773a  and  a48766a );
 a48778a <=( (not A168)  and  A169 );
 a48779a <=( A170  and  a48778a );
 a48783a <=( A201  and  (not A200) );
 a48784a <=( A199  and  a48783a );
 a48785a <=( a48784a  and  a48779a );
 a48789a <=( (not A233)  and  A232 );
 a48790a <=( A203  and  a48789a );
 a48793a <=( A235  and  A234 );
 a48796a <=( A299  and  (not A298) );
 a48797a <=( a48796a  and  a48793a );
 a48798a <=( a48797a  and  a48790a );
 a48802a <=( (not A168)  and  A169 );
 a48803a <=( A170  and  a48802a );
 a48807a <=( A201  and  (not A200) );
 a48808a <=( A199  and  a48807a );
 a48809a <=( a48808a  and  a48803a );
 a48813a <=( (not A233)  and  A232 );
 a48814a <=( A203  and  a48813a );
 a48817a <=( A235  and  A234 );
 a48820a <=( A266  and  (not A265) );
 a48821a <=( a48820a  and  a48817a );
 a48822a <=( a48821a  and  a48814a );
 a48826a <=( (not A168)  and  A169 );
 a48827a <=( A170  and  a48826a );
 a48831a <=( A201  and  (not A200) );
 a48832a <=( A199  and  a48831a );
 a48833a <=( a48832a  and  a48827a );
 a48837a <=( (not A233)  and  A232 );
 a48838a <=( A203  and  a48837a );
 a48841a <=( A236  and  A234 );
 a48844a <=( A299  and  (not A298) );
 a48845a <=( a48844a  and  a48841a );
 a48846a <=( a48845a  and  a48838a );
 a48850a <=( (not A168)  and  A169 );
 a48851a <=( A170  and  a48850a );
 a48855a <=( A201  and  (not A200) );
 a48856a <=( A199  and  a48855a );
 a48857a <=( a48856a  and  a48851a );
 a48861a <=( (not A233)  and  A232 );
 a48862a <=( A203  and  a48861a );
 a48865a <=( A236  and  A234 );
 a48868a <=( A266  and  (not A265) );
 a48869a <=( a48868a  and  a48865a );
 a48870a <=( a48869a  and  a48862a );
 a48874a <=( (not A168)  and  A169 );
 a48875a <=( A170  and  a48874a );
 a48879a <=( A201  and  (not A200) );
 a48880a <=( A199  and  a48879a );
 a48881a <=( a48880a  and  a48875a );
 a48885a <=( (not A233)  and  (not A232) );
 a48886a <=( A203  and  a48885a );
 a48889a <=( A266  and  A265 );
 a48892a <=( (not A300)  and  A298 );
 a48893a <=( a48892a  and  a48889a );
 a48894a <=( a48893a  and  a48886a );
 a48898a <=( (not A168)  and  A169 );
 a48899a <=( A170  and  a48898a );
 a48903a <=( A201  and  (not A200) );
 a48904a <=( A199  and  a48903a );
 a48905a <=( a48904a  and  a48899a );
 a48909a <=( (not A233)  and  (not A232) );
 a48910a <=( A203  and  a48909a );
 a48913a <=( A266  and  A265 );
 a48916a <=( A299  and  A298 );
 a48917a <=( a48916a  and  a48913a );
 a48918a <=( a48917a  and  a48910a );
 a48922a <=( (not A168)  and  A169 );
 a48923a <=( A170  and  a48922a );
 a48927a <=( A201  and  (not A200) );
 a48928a <=( A199  and  a48927a );
 a48929a <=( a48928a  and  a48923a );
 a48933a <=( (not A233)  and  (not A232) );
 a48934a <=( A203  and  a48933a );
 a48937a <=( A266  and  A265 );
 a48940a <=( (not A299)  and  (not A298) );
 a48941a <=( a48940a  and  a48937a );
 a48942a <=( a48941a  and  a48934a );
 a48946a <=( (not A168)  and  A169 );
 a48947a <=( A170  and  a48946a );
 a48951a <=( A201  and  (not A200) );
 a48952a <=( A199  and  a48951a );
 a48953a <=( a48952a  and  a48947a );
 a48957a <=( (not A233)  and  (not A232) );
 a48958a <=( A203  and  a48957a );
 a48961a <=( (not A267)  and  (not A266) );
 a48964a <=( (not A300)  and  A298 );
 a48965a <=( a48964a  and  a48961a );
 a48966a <=( a48965a  and  a48958a );
 a48970a <=( (not A168)  and  A169 );
 a48971a <=( A170  and  a48970a );
 a48975a <=( A201  and  (not A200) );
 a48976a <=( A199  and  a48975a );
 a48977a <=( a48976a  and  a48971a );
 a48981a <=( (not A233)  and  (not A232) );
 a48982a <=( A203  and  a48981a );
 a48985a <=( (not A267)  and  (not A266) );
 a48988a <=( A299  and  A298 );
 a48989a <=( a48988a  and  a48985a );
 a48990a <=( a48989a  and  a48982a );
 a48994a <=( (not A168)  and  A169 );
 a48995a <=( A170  and  a48994a );
 a48999a <=( A201  and  (not A200) );
 a49000a <=( A199  and  a48999a );
 a49001a <=( a49000a  and  a48995a );
 a49005a <=( (not A233)  and  (not A232) );
 a49006a <=( A203  and  a49005a );
 a49009a <=( (not A267)  and  (not A266) );
 a49012a <=( (not A299)  and  (not A298) );
 a49013a <=( a49012a  and  a49009a );
 a49014a <=( a49013a  and  a49006a );
 a49018a <=( (not A168)  and  A169 );
 a49019a <=( A170  and  a49018a );
 a49023a <=( A201  and  (not A200) );
 a49024a <=( A199  and  a49023a );
 a49025a <=( a49024a  and  a49019a );
 a49029a <=( (not A233)  and  (not A232) );
 a49030a <=( A203  and  a49029a );
 a49033a <=( (not A266)  and  (not A265) );
 a49036a <=( (not A300)  and  A298 );
 a49037a <=( a49036a  and  a49033a );
 a49038a <=( a49037a  and  a49030a );
 a49042a <=( (not A168)  and  A169 );
 a49043a <=( A170  and  a49042a );
 a49047a <=( A201  and  (not A200) );
 a49048a <=( A199  and  a49047a );
 a49049a <=( a49048a  and  a49043a );
 a49053a <=( (not A233)  and  (not A232) );
 a49054a <=( A203  and  a49053a );
 a49057a <=( (not A266)  and  (not A265) );
 a49060a <=( A299  and  A298 );
 a49061a <=( a49060a  and  a49057a );
 a49062a <=( a49061a  and  a49054a );
 a49066a <=( (not A168)  and  A169 );
 a49067a <=( A170  and  a49066a );
 a49071a <=( A201  and  (not A200) );
 a49072a <=( A199  and  a49071a );
 a49073a <=( a49072a  and  a49067a );
 a49077a <=( (not A233)  and  (not A232) );
 a49078a <=( A203  and  a49077a );
 a49081a <=( (not A266)  and  (not A265) );
 a49084a <=( (not A299)  and  (not A298) );
 a49085a <=( a49084a  and  a49081a );
 a49086a <=( a49085a  and  a49078a );
 a49090a <=( A167  and  A169 );
 a49091a <=( (not A170)  and  a49090a );
 a49095a <=( A200  and  A199 );
 a49096a <=( A166  and  a49095a );
 a49097a <=( a49096a  and  a49091a );
 a49101a <=( A265  and  A233 );
 a49102a <=( A232  and  a49101a );
 a49105a <=( (not A269)  and  (not A268) );
 a49108a <=( (not A300)  and  (not A299) );
 a49109a <=( a49108a  and  a49105a );
 a49110a <=( a49109a  and  a49102a );
 a49114a <=( A167  and  A169 );
 a49115a <=( (not A170)  and  a49114a );
 a49119a <=( A200  and  A199 );
 a49120a <=( A166  and  a49119a );
 a49121a <=( a49120a  and  a49115a );
 a49125a <=( A265  and  A233 );
 a49126a <=( A232  and  a49125a );
 a49129a <=( (not A269)  and  (not A268) );
 a49132a <=( A299  and  A298 );
 a49133a <=( a49132a  and  a49129a );
 a49134a <=( a49133a  and  a49126a );
 a49138a <=( A167  and  A169 );
 a49139a <=( (not A170)  and  a49138a );
 a49143a <=( A200  and  A199 );
 a49144a <=( A166  and  a49143a );
 a49145a <=( a49144a  and  a49139a );
 a49149a <=( A265  and  A233 );
 a49150a <=( A232  and  a49149a );
 a49153a <=( (not A269)  and  (not A268) );
 a49156a <=( (not A299)  and  (not A298) );
 a49157a <=( a49156a  and  a49153a );
 a49158a <=( a49157a  and  a49150a );
 a49162a <=( A167  and  A169 );
 a49163a <=( (not A170)  and  a49162a );
 a49167a <=( A200  and  A199 );
 a49168a <=( A166  and  a49167a );
 a49169a <=( a49168a  and  a49163a );
 a49173a <=( A265  and  A233 );
 a49174a <=( A232  and  a49173a );
 a49177a <=( (not A299)  and  (not A267) );
 a49180a <=( (not A302)  and  (not A301) );
 a49181a <=( a49180a  and  a49177a );
 a49182a <=( a49181a  and  a49174a );
 a49186a <=( A167  and  A169 );
 a49187a <=( (not A170)  and  a49186a );
 a49191a <=( A200  and  A199 );
 a49192a <=( A166  and  a49191a );
 a49193a <=( a49192a  and  a49187a );
 a49197a <=( A265  and  A233 );
 a49198a <=( A232  and  a49197a );
 a49201a <=( (not A299)  and  A266 );
 a49204a <=( (not A302)  and  (not A301) );
 a49205a <=( a49204a  and  a49201a );
 a49206a <=( a49205a  and  a49198a );
 a49210a <=( A167  and  A169 );
 a49211a <=( (not A170)  and  a49210a );
 a49215a <=( A200  and  A199 );
 a49216a <=( A166  and  a49215a );
 a49217a <=( a49216a  and  a49211a );
 a49221a <=( (not A265)  and  A233 );
 a49222a <=( A232  and  a49221a );
 a49225a <=( (not A299)  and  (not A266) );
 a49228a <=( (not A302)  and  (not A301) );
 a49229a <=( a49228a  and  a49225a );
 a49230a <=( a49229a  and  a49222a );
 a49234a <=( A167  and  A169 );
 a49235a <=( (not A170)  and  a49234a );
 a49239a <=( A200  and  A199 );
 a49240a <=( A166  and  a49239a );
 a49241a <=( a49240a  and  a49235a );
 a49245a <=( (not A236)  and  (not A235) );
 a49246a <=( (not A233)  and  a49245a );
 a49249a <=( A266  and  A265 );
 a49252a <=( (not A300)  and  A298 );
 a49253a <=( a49252a  and  a49249a );
 a49254a <=( a49253a  and  a49246a );
 a49258a <=( A167  and  A169 );
 a49259a <=( (not A170)  and  a49258a );
 a49263a <=( A200  and  A199 );
 a49264a <=( A166  and  a49263a );
 a49265a <=( a49264a  and  a49259a );
 a49269a <=( (not A236)  and  (not A235) );
 a49270a <=( (not A233)  and  a49269a );
 a49273a <=( A266  and  A265 );
 a49276a <=( A299  and  A298 );
 a49277a <=( a49276a  and  a49273a );
 a49278a <=( a49277a  and  a49270a );
 a49282a <=( A167  and  A169 );
 a49283a <=( (not A170)  and  a49282a );
 a49287a <=( A200  and  A199 );
 a49288a <=( A166  and  a49287a );
 a49289a <=( a49288a  and  a49283a );
 a49293a <=( (not A236)  and  (not A235) );
 a49294a <=( (not A233)  and  a49293a );
 a49297a <=( A266  and  A265 );
 a49300a <=( (not A299)  and  (not A298) );
 a49301a <=( a49300a  and  a49297a );
 a49302a <=( a49301a  and  a49294a );
 a49306a <=( A167  and  A169 );
 a49307a <=( (not A170)  and  a49306a );
 a49311a <=( A200  and  A199 );
 a49312a <=( A166  and  a49311a );
 a49313a <=( a49312a  and  a49307a );
 a49317a <=( (not A236)  and  (not A235) );
 a49318a <=( (not A233)  and  a49317a );
 a49321a <=( (not A267)  and  (not A266) );
 a49324a <=( (not A300)  and  A298 );
 a49325a <=( a49324a  and  a49321a );
 a49326a <=( a49325a  and  a49318a );
 a49330a <=( A167  and  A169 );
 a49331a <=( (not A170)  and  a49330a );
 a49335a <=( A200  and  A199 );
 a49336a <=( A166  and  a49335a );
 a49337a <=( a49336a  and  a49331a );
 a49341a <=( (not A236)  and  (not A235) );
 a49342a <=( (not A233)  and  a49341a );
 a49345a <=( (not A267)  and  (not A266) );
 a49348a <=( A299  and  A298 );
 a49349a <=( a49348a  and  a49345a );
 a49350a <=( a49349a  and  a49342a );
 a49354a <=( A167  and  A169 );
 a49355a <=( (not A170)  and  a49354a );
 a49359a <=( A200  and  A199 );
 a49360a <=( A166  and  a49359a );
 a49361a <=( a49360a  and  a49355a );
 a49365a <=( (not A236)  and  (not A235) );
 a49366a <=( (not A233)  and  a49365a );
 a49369a <=( (not A267)  and  (not A266) );
 a49372a <=( (not A299)  and  (not A298) );
 a49373a <=( a49372a  and  a49369a );
 a49374a <=( a49373a  and  a49366a );
 a49378a <=( A167  and  A169 );
 a49379a <=( (not A170)  and  a49378a );
 a49383a <=( A200  and  A199 );
 a49384a <=( A166  and  a49383a );
 a49385a <=( a49384a  and  a49379a );
 a49389a <=( (not A236)  and  (not A235) );
 a49390a <=( (not A233)  and  a49389a );
 a49393a <=( (not A266)  and  (not A265) );
 a49396a <=( (not A300)  and  A298 );
 a49397a <=( a49396a  and  a49393a );
 a49398a <=( a49397a  and  a49390a );
 a49402a <=( A167  and  A169 );
 a49403a <=( (not A170)  and  a49402a );
 a49407a <=( A200  and  A199 );
 a49408a <=( A166  and  a49407a );
 a49409a <=( a49408a  and  a49403a );
 a49413a <=( (not A236)  and  (not A235) );
 a49414a <=( (not A233)  and  a49413a );
 a49417a <=( (not A266)  and  (not A265) );
 a49420a <=( A299  and  A298 );
 a49421a <=( a49420a  and  a49417a );
 a49422a <=( a49421a  and  a49414a );
 a49426a <=( A167  and  A169 );
 a49427a <=( (not A170)  and  a49426a );
 a49431a <=( A200  and  A199 );
 a49432a <=( A166  and  a49431a );
 a49433a <=( a49432a  and  a49427a );
 a49437a <=( (not A236)  and  (not A235) );
 a49438a <=( (not A233)  and  a49437a );
 a49441a <=( (not A266)  and  (not A265) );
 a49444a <=( (not A299)  and  (not A298) );
 a49445a <=( a49444a  and  a49441a );
 a49446a <=( a49445a  and  a49438a );
 a49450a <=( A167  and  A169 );
 a49451a <=( (not A170)  and  a49450a );
 a49455a <=( A200  and  A199 );
 a49456a <=( A166  and  a49455a );
 a49457a <=( a49456a  and  a49451a );
 a49461a <=( A265  and  (not A234) );
 a49462a <=( (not A233)  and  a49461a );
 a49465a <=( A298  and  A266 );
 a49468a <=( (not A302)  and  (not A301) );
 a49469a <=( a49468a  and  a49465a );
 a49470a <=( a49469a  and  a49462a );
 a49474a <=( A167  and  A169 );
 a49475a <=( (not A170)  and  a49474a );
 a49479a <=( A200  and  A199 );
 a49480a <=( A166  and  a49479a );
 a49481a <=( a49480a  and  a49475a );
 a49485a <=( (not A266)  and  (not A234) );
 a49486a <=( (not A233)  and  a49485a );
 a49489a <=( (not A269)  and  (not A268) );
 a49492a <=( (not A300)  and  A298 );
 a49493a <=( a49492a  and  a49489a );
 a49494a <=( a49493a  and  a49486a );
 a49498a <=( A167  and  A169 );
 a49499a <=( (not A170)  and  a49498a );
 a49503a <=( A200  and  A199 );
 a49504a <=( A166  and  a49503a );
 a49505a <=( a49504a  and  a49499a );
 a49509a <=( (not A266)  and  (not A234) );
 a49510a <=( (not A233)  and  a49509a );
 a49513a <=( (not A269)  and  (not A268) );
 a49516a <=( A299  and  A298 );
 a49517a <=( a49516a  and  a49513a );
 a49518a <=( a49517a  and  a49510a );
 a49522a <=( A167  and  A169 );
 a49523a <=( (not A170)  and  a49522a );
 a49527a <=( A200  and  A199 );
 a49528a <=( A166  and  a49527a );
 a49529a <=( a49528a  and  a49523a );
 a49533a <=( (not A266)  and  (not A234) );
 a49534a <=( (not A233)  and  a49533a );
 a49537a <=( (not A269)  and  (not A268) );
 a49540a <=( (not A299)  and  (not A298) );
 a49541a <=( a49540a  and  a49537a );
 a49542a <=( a49541a  and  a49534a );
 a49546a <=( A167  and  A169 );
 a49547a <=( (not A170)  and  a49546a );
 a49551a <=( A200  and  A199 );
 a49552a <=( A166  and  a49551a );
 a49553a <=( a49552a  and  a49547a );
 a49557a <=( (not A266)  and  (not A234) );
 a49558a <=( (not A233)  and  a49557a );
 a49561a <=( A298  and  (not A267) );
 a49564a <=( (not A302)  and  (not A301) );
 a49565a <=( a49564a  and  a49561a );
 a49566a <=( a49565a  and  a49558a );
 a49570a <=( A167  and  A169 );
 a49571a <=( (not A170)  and  a49570a );
 a49575a <=( A200  and  A199 );
 a49576a <=( A166  and  a49575a );
 a49577a <=( a49576a  and  a49571a );
 a49581a <=( (not A265)  and  (not A234) );
 a49582a <=( (not A233)  and  a49581a );
 a49585a <=( A298  and  (not A266) );
 a49588a <=( (not A302)  and  (not A301) );
 a49589a <=( a49588a  and  a49585a );
 a49590a <=( a49589a  and  a49582a );
 a49594a <=( A167  and  A169 );
 a49595a <=( (not A170)  and  a49594a );
 a49599a <=( A200  and  A199 );
 a49600a <=( A166  and  a49599a );
 a49601a <=( a49600a  and  a49595a );
 a49605a <=( A265  and  (not A233) );
 a49606a <=( (not A232)  and  a49605a );
 a49609a <=( A298  and  A266 );
 a49612a <=( (not A302)  and  (not A301) );
 a49613a <=( a49612a  and  a49609a );
 a49614a <=( a49613a  and  a49606a );
 a49618a <=( A167  and  A169 );
 a49619a <=( (not A170)  and  a49618a );
 a49623a <=( A200  and  A199 );
 a49624a <=( A166  and  a49623a );
 a49625a <=( a49624a  and  a49619a );
 a49629a <=( (not A266)  and  (not A233) );
 a49630a <=( (not A232)  and  a49629a );
 a49633a <=( (not A269)  and  (not A268) );
 a49636a <=( (not A300)  and  A298 );
 a49637a <=( a49636a  and  a49633a );
 a49638a <=( a49637a  and  a49630a );
 a49642a <=( A167  and  A169 );
 a49643a <=( (not A170)  and  a49642a );
 a49647a <=( A200  and  A199 );
 a49648a <=( A166  and  a49647a );
 a49649a <=( a49648a  and  a49643a );
 a49653a <=( (not A266)  and  (not A233) );
 a49654a <=( (not A232)  and  a49653a );
 a49657a <=( (not A269)  and  (not A268) );
 a49660a <=( A299  and  A298 );
 a49661a <=( a49660a  and  a49657a );
 a49662a <=( a49661a  and  a49654a );
 a49666a <=( A167  and  A169 );
 a49667a <=( (not A170)  and  a49666a );
 a49671a <=( A200  and  A199 );
 a49672a <=( A166  and  a49671a );
 a49673a <=( a49672a  and  a49667a );
 a49677a <=( (not A266)  and  (not A233) );
 a49678a <=( (not A232)  and  a49677a );
 a49681a <=( (not A269)  and  (not A268) );
 a49684a <=( (not A299)  and  (not A298) );
 a49685a <=( a49684a  and  a49681a );
 a49686a <=( a49685a  and  a49678a );
 a49690a <=( A167  and  A169 );
 a49691a <=( (not A170)  and  a49690a );
 a49695a <=( A200  and  A199 );
 a49696a <=( A166  and  a49695a );
 a49697a <=( a49696a  and  a49691a );
 a49701a <=( (not A266)  and  (not A233) );
 a49702a <=( (not A232)  and  a49701a );
 a49705a <=( A298  and  (not A267) );
 a49708a <=( (not A302)  and  (not A301) );
 a49709a <=( a49708a  and  a49705a );
 a49710a <=( a49709a  and  a49702a );
 a49714a <=( A167  and  A169 );
 a49715a <=( (not A170)  and  a49714a );
 a49719a <=( A200  and  A199 );
 a49720a <=( A166  and  a49719a );
 a49721a <=( a49720a  and  a49715a );
 a49725a <=( (not A265)  and  (not A233) );
 a49726a <=( (not A232)  and  a49725a );
 a49729a <=( A298  and  (not A266) );
 a49732a <=( (not A302)  and  (not A301) );
 a49733a <=( a49732a  and  a49729a );
 a49734a <=( a49733a  and  a49726a );
 a49738a <=( A167  and  A169 );
 a49739a <=( (not A170)  and  a49738a );
 a49743a <=( (not A202)  and  (not A200) );
 a49744a <=( A166  and  a49743a );
 a49745a <=( a49744a  and  a49739a );
 a49749a <=( A233  and  A232 );
 a49750a <=( (not A203)  and  a49749a );
 a49753a <=( (not A267)  and  A265 );
 a49756a <=( (not A300)  and  (not A299) );
 a49757a <=( a49756a  and  a49753a );
 a49758a <=( a49757a  and  a49750a );
 a49762a <=( A167  and  A169 );
 a49763a <=( (not A170)  and  a49762a );
 a49767a <=( (not A202)  and  (not A200) );
 a49768a <=( A166  and  a49767a );
 a49769a <=( a49768a  and  a49763a );
 a49773a <=( A233  and  A232 );
 a49774a <=( (not A203)  and  a49773a );
 a49777a <=( (not A267)  and  A265 );
 a49780a <=( A299  and  A298 );
 a49781a <=( a49780a  and  a49777a );
 a49782a <=( a49781a  and  a49774a );
 a49786a <=( A167  and  A169 );
 a49787a <=( (not A170)  and  a49786a );
 a49791a <=( (not A202)  and  (not A200) );
 a49792a <=( A166  and  a49791a );
 a49793a <=( a49792a  and  a49787a );
 a49797a <=( A233  and  A232 );
 a49798a <=( (not A203)  and  a49797a );
 a49801a <=( (not A267)  and  A265 );
 a49804a <=( (not A299)  and  (not A298) );
 a49805a <=( a49804a  and  a49801a );
 a49806a <=( a49805a  and  a49798a );
 a49810a <=( A167  and  A169 );
 a49811a <=( (not A170)  and  a49810a );
 a49815a <=( (not A202)  and  (not A200) );
 a49816a <=( A166  and  a49815a );
 a49817a <=( a49816a  and  a49811a );
 a49821a <=( A233  and  A232 );
 a49822a <=( (not A203)  and  a49821a );
 a49825a <=( A266  and  A265 );
 a49828a <=( (not A300)  and  (not A299) );
 a49829a <=( a49828a  and  a49825a );
 a49830a <=( a49829a  and  a49822a );
 a49834a <=( A167  and  A169 );
 a49835a <=( (not A170)  and  a49834a );
 a49839a <=( (not A202)  and  (not A200) );
 a49840a <=( A166  and  a49839a );
 a49841a <=( a49840a  and  a49835a );
 a49845a <=( A233  and  A232 );
 a49846a <=( (not A203)  and  a49845a );
 a49849a <=( A266  and  A265 );
 a49852a <=( A299  and  A298 );
 a49853a <=( a49852a  and  a49849a );
 a49854a <=( a49853a  and  a49846a );
 a49858a <=( A167  and  A169 );
 a49859a <=( (not A170)  and  a49858a );
 a49863a <=( (not A202)  and  (not A200) );
 a49864a <=( A166  and  a49863a );
 a49865a <=( a49864a  and  a49859a );
 a49869a <=( A233  and  A232 );
 a49870a <=( (not A203)  and  a49869a );
 a49873a <=( A266  and  A265 );
 a49876a <=( (not A299)  and  (not A298) );
 a49877a <=( a49876a  and  a49873a );
 a49878a <=( a49877a  and  a49870a );
 a49882a <=( A167  and  A169 );
 a49883a <=( (not A170)  and  a49882a );
 a49887a <=( (not A202)  and  (not A200) );
 a49888a <=( A166  and  a49887a );
 a49889a <=( a49888a  and  a49883a );
 a49893a <=( A233  and  A232 );
 a49894a <=( (not A203)  and  a49893a );
 a49897a <=( (not A266)  and  (not A265) );
 a49900a <=( (not A300)  and  (not A299) );
 a49901a <=( a49900a  and  a49897a );
 a49902a <=( a49901a  and  a49894a );
 a49906a <=( A167  and  A169 );
 a49907a <=( (not A170)  and  a49906a );
 a49911a <=( (not A202)  and  (not A200) );
 a49912a <=( A166  and  a49911a );
 a49913a <=( a49912a  and  a49907a );
 a49917a <=( A233  and  A232 );
 a49918a <=( (not A203)  and  a49917a );
 a49921a <=( (not A266)  and  (not A265) );
 a49924a <=( A299  and  A298 );
 a49925a <=( a49924a  and  a49921a );
 a49926a <=( a49925a  and  a49918a );
 a49930a <=( A167  and  A169 );
 a49931a <=( (not A170)  and  a49930a );
 a49935a <=( (not A202)  and  (not A200) );
 a49936a <=( A166  and  a49935a );
 a49937a <=( a49936a  and  a49931a );
 a49941a <=( A233  and  A232 );
 a49942a <=( (not A203)  and  a49941a );
 a49945a <=( (not A266)  and  (not A265) );
 a49948a <=( (not A299)  and  (not A298) );
 a49949a <=( a49948a  and  a49945a );
 a49950a <=( a49949a  and  a49942a );
 a49954a <=( A167  and  A169 );
 a49955a <=( (not A170)  and  a49954a );
 a49959a <=( (not A202)  and  (not A200) );
 a49960a <=( A166  and  a49959a );
 a49961a <=( a49960a  and  a49955a );
 a49965a <=( A233  and  (not A232) );
 a49966a <=( (not A203)  and  a49965a );
 a49969a <=( (not A299)  and  A298 );
 a49972a <=( A301  and  A300 );
 a49973a <=( a49972a  and  a49969a );
 a49974a <=( a49973a  and  a49966a );
 a49978a <=( A167  and  A169 );
 a49979a <=( (not A170)  and  a49978a );
 a49983a <=( (not A202)  and  (not A200) );
 a49984a <=( A166  and  a49983a );
 a49985a <=( a49984a  and  a49979a );
 a49989a <=( A233  and  (not A232) );
 a49990a <=( (not A203)  and  a49989a );
 a49993a <=( (not A299)  and  A298 );
 a49996a <=( A302  and  A300 );
 a49997a <=( a49996a  and  a49993a );
 a49998a <=( a49997a  and  a49990a );
 a50002a <=( A167  and  A169 );
 a50003a <=( (not A170)  and  a50002a );
 a50007a <=( (not A202)  and  (not A200) );
 a50008a <=( A166  and  a50007a );
 a50009a <=( a50008a  and  a50003a );
 a50013a <=( A233  and  (not A232) );
 a50014a <=( (not A203)  and  a50013a );
 a50017a <=( (not A266)  and  A265 );
 a50020a <=( A268  and  A267 );
 a50021a <=( a50020a  and  a50017a );
 a50022a <=( a50021a  and  a50014a );
 a50026a <=( A167  and  A169 );
 a50027a <=( (not A170)  and  a50026a );
 a50031a <=( (not A202)  and  (not A200) );
 a50032a <=( A166  and  a50031a );
 a50033a <=( a50032a  and  a50027a );
 a50037a <=( A233  and  (not A232) );
 a50038a <=( (not A203)  and  a50037a );
 a50041a <=( (not A266)  and  A265 );
 a50044a <=( A269  and  A267 );
 a50045a <=( a50044a  and  a50041a );
 a50046a <=( a50045a  and  a50038a );
 a50050a <=( A167  and  A169 );
 a50051a <=( (not A170)  and  a50050a );
 a50055a <=( (not A202)  and  (not A200) );
 a50056a <=( A166  and  a50055a );
 a50057a <=( a50056a  and  a50051a );
 a50061a <=( (not A234)  and  (not A233) );
 a50062a <=( (not A203)  and  a50061a );
 a50065a <=( A266  and  A265 );
 a50068a <=( (not A300)  and  A298 );
 a50069a <=( a50068a  and  a50065a );
 a50070a <=( a50069a  and  a50062a );
 a50074a <=( A167  and  A169 );
 a50075a <=( (not A170)  and  a50074a );
 a50079a <=( (not A202)  and  (not A200) );
 a50080a <=( A166  and  a50079a );
 a50081a <=( a50080a  and  a50075a );
 a50085a <=( (not A234)  and  (not A233) );
 a50086a <=( (not A203)  and  a50085a );
 a50089a <=( A266  and  A265 );
 a50092a <=( A299  and  A298 );
 a50093a <=( a50092a  and  a50089a );
 a50094a <=( a50093a  and  a50086a );
 a50098a <=( A167  and  A169 );
 a50099a <=( (not A170)  and  a50098a );
 a50103a <=( (not A202)  and  (not A200) );
 a50104a <=( A166  and  a50103a );
 a50105a <=( a50104a  and  a50099a );
 a50109a <=( (not A234)  and  (not A233) );
 a50110a <=( (not A203)  and  a50109a );
 a50113a <=( A266  and  A265 );
 a50116a <=( (not A299)  and  (not A298) );
 a50117a <=( a50116a  and  a50113a );
 a50118a <=( a50117a  and  a50110a );
 a50122a <=( A167  and  A169 );
 a50123a <=( (not A170)  and  a50122a );
 a50127a <=( (not A202)  and  (not A200) );
 a50128a <=( A166  and  a50127a );
 a50129a <=( a50128a  and  a50123a );
 a50133a <=( (not A234)  and  (not A233) );
 a50134a <=( (not A203)  and  a50133a );
 a50137a <=( (not A267)  and  (not A266) );
 a50140a <=( (not A300)  and  A298 );
 a50141a <=( a50140a  and  a50137a );
 a50142a <=( a50141a  and  a50134a );
 a50146a <=( A167  and  A169 );
 a50147a <=( (not A170)  and  a50146a );
 a50151a <=( (not A202)  and  (not A200) );
 a50152a <=( A166  and  a50151a );
 a50153a <=( a50152a  and  a50147a );
 a50157a <=( (not A234)  and  (not A233) );
 a50158a <=( (not A203)  and  a50157a );
 a50161a <=( (not A267)  and  (not A266) );
 a50164a <=( A299  and  A298 );
 a50165a <=( a50164a  and  a50161a );
 a50166a <=( a50165a  and  a50158a );
 a50170a <=( A167  and  A169 );
 a50171a <=( (not A170)  and  a50170a );
 a50175a <=( (not A202)  and  (not A200) );
 a50176a <=( A166  and  a50175a );
 a50177a <=( a50176a  and  a50171a );
 a50181a <=( (not A234)  and  (not A233) );
 a50182a <=( (not A203)  and  a50181a );
 a50185a <=( (not A267)  and  (not A266) );
 a50188a <=( (not A299)  and  (not A298) );
 a50189a <=( a50188a  and  a50185a );
 a50190a <=( a50189a  and  a50182a );
 a50194a <=( A167  and  A169 );
 a50195a <=( (not A170)  and  a50194a );
 a50199a <=( (not A202)  and  (not A200) );
 a50200a <=( A166  and  a50199a );
 a50201a <=( a50200a  and  a50195a );
 a50205a <=( (not A234)  and  (not A233) );
 a50206a <=( (not A203)  and  a50205a );
 a50209a <=( (not A266)  and  (not A265) );
 a50212a <=( (not A300)  and  A298 );
 a50213a <=( a50212a  and  a50209a );
 a50214a <=( a50213a  and  a50206a );
 a50218a <=( A167  and  A169 );
 a50219a <=( (not A170)  and  a50218a );
 a50223a <=( (not A202)  and  (not A200) );
 a50224a <=( A166  and  a50223a );
 a50225a <=( a50224a  and  a50219a );
 a50229a <=( (not A234)  and  (not A233) );
 a50230a <=( (not A203)  and  a50229a );
 a50233a <=( (not A266)  and  (not A265) );
 a50236a <=( A299  and  A298 );
 a50237a <=( a50236a  and  a50233a );
 a50238a <=( a50237a  and  a50230a );
 a50242a <=( A167  and  A169 );
 a50243a <=( (not A170)  and  a50242a );
 a50247a <=( (not A202)  and  (not A200) );
 a50248a <=( A166  and  a50247a );
 a50249a <=( a50248a  and  a50243a );
 a50253a <=( (not A234)  and  (not A233) );
 a50254a <=( (not A203)  and  a50253a );
 a50257a <=( (not A266)  and  (not A265) );
 a50260a <=( (not A299)  and  (not A298) );
 a50261a <=( a50260a  and  a50257a );
 a50262a <=( a50261a  and  a50254a );
 a50266a <=( A167  and  A169 );
 a50267a <=( (not A170)  and  a50266a );
 a50271a <=( (not A202)  and  (not A200) );
 a50272a <=( A166  and  a50271a );
 a50273a <=( a50272a  and  a50267a );
 a50277a <=( (not A233)  and  A232 );
 a50278a <=( (not A203)  and  a50277a );
 a50281a <=( A235  and  A234 );
 a50284a <=( A299  and  (not A298) );
 a50285a <=( a50284a  and  a50281a );
 a50286a <=( a50285a  and  a50278a );
 a50290a <=( A167  and  A169 );
 a50291a <=( (not A170)  and  a50290a );
 a50295a <=( (not A202)  and  (not A200) );
 a50296a <=( A166  and  a50295a );
 a50297a <=( a50296a  and  a50291a );
 a50301a <=( (not A233)  and  A232 );
 a50302a <=( (not A203)  and  a50301a );
 a50305a <=( A235  and  A234 );
 a50308a <=( A266  and  (not A265) );
 a50309a <=( a50308a  and  a50305a );
 a50310a <=( a50309a  and  a50302a );
 a50314a <=( A167  and  A169 );
 a50315a <=( (not A170)  and  a50314a );
 a50319a <=( (not A202)  and  (not A200) );
 a50320a <=( A166  and  a50319a );
 a50321a <=( a50320a  and  a50315a );
 a50325a <=( (not A233)  and  A232 );
 a50326a <=( (not A203)  and  a50325a );
 a50329a <=( A236  and  A234 );
 a50332a <=( A299  and  (not A298) );
 a50333a <=( a50332a  and  a50329a );
 a50334a <=( a50333a  and  a50326a );
 a50338a <=( A167  and  A169 );
 a50339a <=( (not A170)  and  a50338a );
 a50343a <=( (not A202)  and  (not A200) );
 a50344a <=( A166  and  a50343a );
 a50345a <=( a50344a  and  a50339a );
 a50349a <=( (not A233)  and  A232 );
 a50350a <=( (not A203)  and  a50349a );
 a50353a <=( A236  and  A234 );
 a50356a <=( A266  and  (not A265) );
 a50357a <=( a50356a  and  a50353a );
 a50358a <=( a50357a  and  a50350a );
 a50362a <=( A167  and  A169 );
 a50363a <=( (not A170)  and  a50362a );
 a50367a <=( (not A202)  and  (not A200) );
 a50368a <=( A166  and  a50367a );
 a50369a <=( a50368a  and  a50363a );
 a50373a <=( (not A233)  and  (not A232) );
 a50374a <=( (not A203)  and  a50373a );
 a50377a <=( A266  and  A265 );
 a50380a <=( (not A300)  and  A298 );
 a50381a <=( a50380a  and  a50377a );
 a50382a <=( a50381a  and  a50374a );
 a50386a <=( A167  and  A169 );
 a50387a <=( (not A170)  and  a50386a );
 a50391a <=( (not A202)  and  (not A200) );
 a50392a <=( A166  and  a50391a );
 a50393a <=( a50392a  and  a50387a );
 a50397a <=( (not A233)  and  (not A232) );
 a50398a <=( (not A203)  and  a50397a );
 a50401a <=( A266  and  A265 );
 a50404a <=( A299  and  A298 );
 a50405a <=( a50404a  and  a50401a );
 a50406a <=( a50405a  and  a50398a );
 a50410a <=( A167  and  A169 );
 a50411a <=( (not A170)  and  a50410a );
 a50415a <=( (not A202)  and  (not A200) );
 a50416a <=( A166  and  a50415a );
 a50417a <=( a50416a  and  a50411a );
 a50421a <=( (not A233)  and  (not A232) );
 a50422a <=( (not A203)  and  a50421a );
 a50425a <=( A266  and  A265 );
 a50428a <=( (not A299)  and  (not A298) );
 a50429a <=( a50428a  and  a50425a );
 a50430a <=( a50429a  and  a50422a );
 a50434a <=( A167  and  A169 );
 a50435a <=( (not A170)  and  a50434a );
 a50439a <=( (not A202)  and  (not A200) );
 a50440a <=( A166  and  a50439a );
 a50441a <=( a50440a  and  a50435a );
 a50445a <=( (not A233)  and  (not A232) );
 a50446a <=( (not A203)  and  a50445a );
 a50449a <=( (not A267)  and  (not A266) );
 a50452a <=( (not A300)  and  A298 );
 a50453a <=( a50452a  and  a50449a );
 a50454a <=( a50453a  and  a50446a );
 a50458a <=( A167  and  A169 );
 a50459a <=( (not A170)  and  a50458a );
 a50463a <=( (not A202)  and  (not A200) );
 a50464a <=( A166  and  a50463a );
 a50465a <=( a50464a  and  a50459a );
 a50469a <=( (not A233)  and  (not A232) );
 a50470a <=( (not A203)  and  a50469a );
 a50473a <=( (not A267)  and  (not A266) );
 a50476a <=( A299  and  A298 );
 a50477a <=( a50476a  and  a50473a );
 a50478a <=( a50477a  and  a50470a );
 a50482a <=( A167  and  A169 );
 a50483a <=( (not A170)  and  a50482a );
 a50487a <=( (not A202)  and  (not A200) );
 a50488a <=( A166  and  a50487a );
 a50489a <=( a50488a  and  a50483a );
 a50493a <=( (not A233)  and  (not A232) );
 a50494a <=( (not A203)  and  a50493a );
 a50497a <=( (not A267)  and  (not A266) );
 a50500a <=( (not A299)  and  (not A298) );
 a50501a <=( a50500a  and  a50497a );
 a50502a <=( a50501a  and  a50494a );
 a50506a <=( A167  and  A169 );
 a50507a <=( (not A170)  and  a50506a );
 a50511a <=( (not A202)  and  (not A200) );
 a50512a <=( A166  and  a50511a );
 a50513a <=( a50512a  and  a50507a );
 a50517a <=( (not A233)  and  (not A232) );
 a50518a <=( (not A203)  and  a50517a );
 a50521a <=( (not A266)  and  (not A265) );
 a50524a <=( (not A300)  and  A298 );
 a50525a <=( a50524a  and  a50521a );
 a50526a <=( a50525a  and  a50518a );
 a50530a <=( A167  and  A169 );
 a50531a <=( (not A170)  and  a50530a );
 a50535a <=( (not A202)  and  (not A200) );
 a50536a <=( A166  and  a50535a );
 a50537a <=( a50536a  and  a50531a );
 a50541a <=( (not A233)  and  (not A232) );
 a50542a <=( (not A203)  and  a50541a );
 a50545a <=( (not A266)  and  (not A265) );
 a50548a <=( A299  and  A298 );
 a50549a <=( a50548a  and  a50545a );
 a50550a <=( a50549a  and  a50542a );
 a50554a <=( A167  and  A169 );
 a50555a <=( (not A170)  and  a50554a );
 a50559a <=( (not A202)  and  (not A200) );
 a50560a <=( A166  and  a50559a );
 a50561a <=( a50560a  and  a50555a );
 a50565a <=( (not A233)  and  (not A232) );
 a50566a <=( (not A203)  and  a50565a );
 a50569a <=( (not A266)  and  (not A265) );
 a50572a <=( (not A299)  and  (not A298) );
 a50573a <=( a50572a  and  a50569a );
 a50574a <=( a50573a  and  a50566a );
 a50578a <=( A167  and  A169 );
 a50579a <=( (not A170)  and  a50578a );
 a50583a <=( (not A201)  and  (not A200) );
 a50584a <=( A166  and  a50583a );
 a50585a <=( a50584a  and  a50579a );
 a50589a <=( A265  and  A233 );
 a50590a <=( A232  and  a50589a );
 a50593a <=( (not A269)  and  (not A268) );
 a50596a <=( (not A300)  and  (not A299) );
 a50597a <=( a50596a  and  a50593a );
 a50598a <=( a50597a  and  a50590a );
 a50602a <=( A167  and  A169 );
 a50603a <=( (not A170)  and  a50602a );
 a50607a <=( (not A201)  and  (not A200) );
 a50608a <=( A166  and  a50607a );
 a50609a <=( a50608a  and  a50603a );
 a50613a <=( A265  and  A233 );
 a50614a <=( A232  and  a50613a );
 a50617a <=( (not A269)  and  (not A268) );
 a50620a <=( A299  and  A298 );
 a50621a <=( a50620a  and  a50617a );
 a50622a <=( a50621a  and  a50614a );
 a50626a <=( A167  and  A169 );
 a50627a <=( (not A170)  and  a50626a );
 a50631a <=( (not A201)  and  (not A200) );
 a50632a <=( A166  and  a50631a );
 a50633a <=( a50632a  and  a50627a );
 a50637a <=( A265  and  A233 );
 a50638a <=( A232  and  a50637a );
 a50641a <=( (not A269)  and  (not A268) );
 a50644a <=( (not A299)  and  (not A298) );
 a50645a <=( a50644a  and  a50641a );
 a50646a <=( a50645a  and  a50638a );
 a50650a <=( A167  and  A169 );
 a50651a <=( (not A170)  and  a50650a );
 a50655a <=( (not A201)  and  (not A200) );
 a50656a <=( A166  and  a50655a );
 a50657a <=( a50656a  and  a50651a );
 a50661a <=( A265  and  A233 );
 a50662a <=( A232  and  a50661a );
 a50665a <=( (not A299)  and  (not A267) );
 a50668a <=( (not A302)  and  (not A301) );
 a50669a <=( a50668a  and  a50665a );
 a50670a <=( a50669a  and  a50662a );
 a50674a <=( A167  and  A169 );
 a50675a <=( (not A170)  and  a50674a );
 a50679a <=( (not A201)  and  (not A200) );
 a50680a <=( A166  and  a50679a );
 a50681a <=( a50680a  and  a50675a );
 a50685a <=( A265  and  A233 );
 a50686a <=( A232  and  a50685a );
 a50689a <=( (not A299)  and  A266 );
 a50692a <=( (not A302)  and  (not A301) );
 a50693a <=( a50692a  and  a50689a );
 a50694a <=( a50693a  and  a50686a );
 a50698a <=( A167  and  A169 );
 a50699a <=( (not A170)  and  a50698a );
 a50703a <=( (not A201)  and  (not A200) );
 a50704a <=( A166  and  a50703a );
 a50705a <=( a50704a  and  a50699a );
 a50709a <=( (not A265)  and  A233 );
 a50710a <=( A232  and  a50709a );
 a50713a <=( (not A299)  and  (not A266) );
 a50716a <=( (not A302)  and  (not A301) );
 a50717a <=( a50716a  and  a50713a );
 a50718a <=( a50717a  and  a50710a );
 a50722a <=( A167  and  A169 );
 a50723a <=( (not A170)  and  a50722a );
 a50727a <=( (not A201)  and  (not A200) );
 a50728a <=( A166  and  a50727a );
 a50729a <=( a50728a  and  a50723a );
 a50733a <=( (not A236)  and  (not A235) );
 a50734a <=( (not A233)  and  a50733a );
 a50737a <=( A266  and  A265 );
 a50740a <=( (not A300)  and  A298 );
 a50741a <=( a50740a  and  a50737a );
 a50742a <=( a50741a  and  a50734a );
 a50746a <=( A167  and  A169 );
 a50747a <=( (not A170)  and  a50746a );
 a50751a <=( (not A201)  and  (not A200) );
 a50752a <=( A166  and  a50751a );
 a50753a <=( a50752a  and  a50747a );
 a50757a <=( (not A236)  and  (not A235) );
 a50758a <=( (not A233)  and  a50757a );
 a50761a <=( A266  and  A265 );
 a50764a <=( A299  and  A298 );
 a50765a <=( a50764a  and  a50761a );
 a50766a <=( a50765a  and  a50758a );
 a50770a <=( A167  and  A169 );
 a50771a <=( (not A170)  and  a50770a );
 a50775a <=( (not A201)  and  (not A200) );
 a50776a <=( A166  and  a50775a );
 a50777a <=( a50776a  and  a50771a );
 a50781a <=( (not A236)  and  (not A235) );
 a50782a <=( (not A233)  and  a50781a );
 a50785a <=( A266  and  A265 );
 a50788a <=( (not A299)  and  (not A298) );
 a50789a <=( a50788a  and  a50785a );
 a50790a <=( a50789a  and  a50782a );
 a50794a <=( A167  and  A169 );
 a50795a <=( (not A170)  and  a50794a );
 a50799a <=( (not A201)  and  (not A200) );
 a50800a <=( A166  and  a50799a );
 a50801a <=( a50800a  and  a50795a );
 a50805a <=( (not A236)  and  (not A235) );
 a50806a <=( (not A233)  and  a50805a );
 a50809a <=( (not A267)  and  (not A266) );
 a50812a <=( (not A300)  and  A298 );
 a50813a <=( a50812a  and  a50809a );
 a50814a <=( a50813a  and  a50806a );
 a50818a <=( A167  and  A169 );
 a50819a <=( (not A170)  and  a50818a );
 a50823a <=( (not A201)  and  (not A200) );
 a50824a <=( A166  and  a50823a );
 a50825a <=( a50824a  and  a50819a );
 a50829a <=( (not A236)  and  (not A235) );
 a50830a <=( (not A233)  and  a50829a );
 a50833a <=( (not A267)  and  (not A266) );
 a50836a <=( A299  and  A298 );
 a50837a <=( a50836a  and  a50833a );
 a50838a <=( a50837a  and  a50830a );
 a50842a <=( A167  and  A169 );
 a50843a <=( (not A170)  and  a50842a );
 a50847a <=( (not A201)  and  (not A200) );
 a50848a <=( A166  and  a50847a );
 a50849a <=( a50848a  and  a50843a );
 a50853a <=( (not A236)  and  (not A235) );
 a50854a <=( (not A233)  and  a50853a );
 a50857a <=( (not A267)  and  (not A266) );
 a50860a <=( (not A299)  and  (not A298) );
 a50861a <=( a50860a  and  a50857a );
 a50862a <=( a50861a  and  a50854a );
 a50866a <=( A167  and  A169 );
 a50867a <=( (not A170)  and  a50866a );
 a50871a <=( (not A201)  and  (not A200) );
 a50872a <=( A166  and  a50871a );
 a50873a <=( a50872a  and  a50867a );
 a50877a <=( (not A236)  and  (not A235) );
 a50878a <=( (not A233)  and  a50877a );
 a50881a <=( (not A266)  and  (not A265) );
 a50884a <=( (not A300)  and  A298 );
 a50885a <=( a50884a  and  a50881a );
 a50886a <=( a50885a  and  a50878a );
 a50890a <=( A167  and  A169 );
 a50891a <=( (not A170)  and  a50890a );
 a50895a <=( (not A201)  and  (not A200) );
 a50896a <=( A166  and  a50895a );
 a50897a <=( a50896a  and  a50891a );
 a50901a <=( (not A236)  and  (not A235) );
 a50902a <=( (not A233)  and  a50901a );
 a50905a <=( (not A266)  and  (not A265) );
 a50908a <=( A299  and  A298 );
 a50909a <=( a50908a  and  a50905a );
 a50910a <=( a50909a  and  a50902a );
 a50914a <=( A167  and  A169 );
 a50915a <=( (not A170)  and  a50914a );
 a50919a <=( (not A201)  and  (not A200) );
 a50920a <=( A166  and  a50919a );
 a50921a <=( a50920a  and  a50915a );
 a50925a <=( (not A236)  and  (not A235) );
 a50926a <=( (not A233)  and  a50925a );
 a50929a <=( (not A266)  and  (not A265) );
 a50932a <=( (not A299)  and  (not A298) );
 a50933a <=( a50932a  and  a50929a );
 a50934a <=( a50933a  and  a50926a );
 a50938a <=( A167  and  A169 );
 a50939a <=( (not A170)  and  a50938a );
 a50943a <=( (not A201)  and  (not A200) );
 a50944a <=( A166  and  a50943a );
 a50945a <=( a50944a  and  a50939a );
 a50949a <=( A265  and  (not A234) );
 a50950a <=( (not A233)  and  a50949a );
 a50953a <=( A298  and  A266 );
 a50956a <=( (not A302)  and  (not A301) );
 a50957a <=( a50956a  and  a50953a );
 a50958a <=( a50957a  and  a50950a );
 a50962a <=( A167  and  A169 );
 a50963a <=( (not A170)  and  a50962a );
 a50967a <=( (not A201)  and  (not A200) );
 a50968a <=( A166  and  a50967a );
 a50969a <=( a50968a  and  a50963a );
 a50973a <=( (not A266)  and  (not A234) );
 a50974a <=( (not A233)  and  a50973a );
 a50977a <=( (not A269)  and  (not A268) );
 a50980a <=( (not A300)  and  A298 );
 a50981a <=( a50980a  and  a50977a );
 a50982a <=( a50981a  and  a50974a );
 a50986a <=( A167  and  A169 );
 a50987a <=( (not A170)  and  a50986a );
 a50991a <=( (not A201)  and  (not A200) );
 a50992a <=( A166  and  a50991a );
 a50993a <=( a50992a  and  a50987a );
 a50997a <=( (not A266)  and  (not A234) );
 a50998a <=( (not A233)  and  a50997a );
 a51001a <=( (not A269)  and  (not A268) );
 a51004a <=( A299  and  A298 );
 a51005a <=( a51004a  and  a51001a );
 a51006a <=( a51005a  and  a50998a );
 a51010a <=( A167  and  A169 );
 a51011a <=( (not A170)  and  a51010a );
 a51015a <=( (not A201)  and  (not A200) );
 a51016a <=( A166  and  a51015a );
 a51017a <=( a51016a  and  a51011a );
 a51021a <=( (not A266)  and  (not A234) );
 a51022a <=( (not A233)  and  a51021a );
 a51025a <=( (not A269)  and  (not A268) );
 a51028a <=( (not A299)  and  (not A298) );
 a51029a <=( a51028a  and  a51025a );
 a51030a <=( a51029a  and  a51022a );
 a51034a <=( A167  and  A169 );
 a51035a <=( (not A170)  and  a51034a );
 a51039a <=( (not A201)  and  (not A200) );
 a51040a <=( A166  and  a51039a );
 a51041a <=( a51040a  and  a51035a );
 a51045a <=( (not A266)  and  (not A234) );
 a51046a <=( (not A233)  and  a51045a );
 a51049a <=( A298  and  (not A267) );
 a51052a <=( (not A302)  and  (not A301) );
 a51053a <=( a51052a  and  a51049a );
 a51054a <=( a51053a  and  a51046a );
 a51058a <=( A167  and  A169 );
 a51059a <=( (not A170)  and  a51058a );
 a51063a <=( (not A201)  and  (not A200) );
 a51064a <=( A166  and  a51063a );
 a51065a <=( a51064a  and  a51059a );
 a51069a <=( (not A265)  and  (not A234) );
 a51070a <=( (not A233)  and  a51069a );
 a51073a <=( A298  and  (not A266) );
 a51076a <=( (not A302)  and  (not A301) );
 a51077a <=( a51076a  and  a51073a );
 a51078a <=( a51077a  and  a51070a );
 a51082a <=( A167  and  A169 );
 a51083a <=( (not A170)  and  a51082a );
 a51087a <=( (not A201)  and  (not A200) );
 a51088a <=( A166  and  a51087a );
 a51089a <=( a51088a  and  a51083a );
 a51093a <=( A265  and  (not A233) );
 a51094a <=( (not A232)  and  a51093a );
 a51097a <=( A298  and  A266 );
 a51100a <=( (not A302)  and  (not A301) );
 a51101a <=( a51100a  and  a51097a );
 a51102a <=( a51101a  and  a51094a );
 a51106a <=( A167  and  A169 );
 a51107a <=( (not A170)  and  a51106a );
 a51111a <=( (not A201)  and  (not A200) );
 a51112a <=( A166  and  a51111a );
 a51113a <=( a51112a  and  a51107a );
 a51117a <=( (not A266)  and  (not A233) );
 a51118a <=( (not A232)  and  a51117a );
 a51121a <=( (not A269)  and  (not A268) );
 a51124a <=( (not A300)  and  A298 );
 a51125a <=( a51124a  and  a51121a );
 a51126a <=( a51125a  and  a51118a );
 a51130a <=( A167  and  A169 );
 a51131a <=( (not A170)  and  a51130a );
 a51135a <=( (not A201)  and  (not A200) );
 a51136a <=( A166  and  a51135a );
 a51137a <=( a51136a  and  a51131a );
 a51141a <=( (not A266)  and  (not A233) );
 a51142a <=( (not A232)  and  a51141a );
 a51145a <=( (not A269)  and  (not A268) );
 a51148a <=( A299  and  A298 );
 a51149a <=( a51148a  and  a51145a );
 a51150a <=( a51149a  and  a51142a );
 a51154a <=( A167  and  A169 );
 a51155a <=( (not A170)  and  a51154a );
 a51159a <=( (not A201)  and  (not A200) );
 a51160a <=( A166  and  a51159a );
 a51161a <=( a51160a  and  a51155a );
 a51165a <=( (not A266)  and  (not A233) );
 a51166a <=( (not A232)  and  a51165a );
 a51169a <=( (not A269)  and  (not A268) );
 a51172a <=( (not A299)  and  (not A298) );
 a51173a <=( a51172a  and  a51169a );
 a51174a <=( a51173a  and  a51166a );
 a51178a <=( A167  and  A169 );
 a51179a <=( (not A170)  and  a51178a );
 a51183a <=( (not A201)  and  (not A200) );
 a51184a <=( A166  and  a51183a );
 a51185a <=( a51184a  and  a51179a );
 a51189a <=( (not A266)  and  (not A233) );
 a51190a <=( (not A232)  and  a51189a );
 a51193a <=( A298  and  (not A267) );
 a51196a <=( (not A302)  and  (not A301) );
 a51197a <=( a51196a  and  a51193a );
 a51198a <=( a51197a  and  a51190a );
 a51202a <=( A167  and  A169 );
 a51203a <=( (not A170)  and  a51202a );
 a51207a <=( (not A201)  and  (not A200) );
 a51208a <=( A166  and  a51207a );
 a51209a <=( a51208a  and  a51203a );
 a51213a <=( (not A265)  and  (not A233) );
 a51214a <=( (not A232)  and  a51213a );
 a51217a <=( A298  and  (not A266) );
 a51220a <=( (not A302)  and  (not A301) );
 a51221a <=( a51220a  and  a51217a );
 a51222a <=( a51221a  and  a51214a );
 a51226a <=( A167  and  A169 );
 a51227a <=( (not A170)  and  a51226a );
 a51231a <=( (not A200)  and  (not A199) );
 a51232a <=( A166  and  a51231a );
 a51233a <=( a51232a  and  a51227a );
 a51237a <=( A265  and  A233 );
 a51238a <=( A232  and  a51237a );
 a51241a <=( (not A269)  and  (not A268) );
 a51244a <=( (not A300)  and  (not A299) );
 a51245a <=( a51244a  and  a51241a );
 a51246a <=( a51245a  and  a51238a );
 a51250a <=( A167  and  A169 );
 a51251a <=( (not A170)  and  a51250a );
 a51255a <=( (not A200)  and  (not A199) );
 a51256a <=( A166  and  a51255a );
 a51257a <=( a51256a  and  a51251a );
 a51261a <=( A265  and  A233 );
 a51262a <=( A232  and  a51261a );
 a51265a <=( (not A269)  and  (not A268) );
 a51268a <=( A299  and  A298 );
 a51269a <=( a51268a  and  a51265a );
 a51270a <=( a51269a  and  a51262a );
 a51274a <=( A167  and  A169 );
 a51275a <=( (not A170)  and  a51274a );
 a51279a <=( (not A200)  and  (not A199) );
 a51280a <=( A166  and  a51279a );
 a51281a <=( a51280a  and  a51275a );
 a51285a <=( A265  and  A233 );
 a51286a <=( A232  and  a51285a );
 a51289a <=( (not A269)  and  (not A268) );
 a51292a <=( (not A299)  and  (not A298) );
 a51293a <=( a51292a  and  a51289a );
 a51294a <=( a51293a  and  a51286a );
 a51298a <=( A167  and  A169 );
 a51299a <=( (not A170)  and  a51298a );
 a51303a <=( (not A200)  and  (not A199) );
 a51304a <=( A166  and  a51303a );
 a51305a <=( a51304a  and  a51299a );
 a51309a <=( A265  and  A233 );
 a51310a <=( A232  and  a51309a );
 a51313a <=( (not A299)  and  (not A267) );
 a51316a <=( (not A302)  and  (not A301) );
 a51317a <=( a51316a  and  a51313a );
 a51318a <=( a51317a  and  a51310a );
 a51322a <=( A167  and  A169 );
 a51323a <=( (not A170)  and  a51322a );
 a51327a <=( (not A200)  and  (not A199) );
 a51328a <=( A166  and  a51327a );
 a51329a <=( a51328a  and  a51323a );
 a51333a <=( A265  and  A233 );
 a51334a <=( A232  and  a51333a );
 a51337a <=( (not A299)  and  A266 );
 a51340a <=( (not A302)  and  (not A301) );
 a51341a <=( a51340a  and  a51337a );
 a51342a <=( a51341a  and  a51334a );
 a51346a <=( A167  and  A169 );
 a51347a <=( (not A170)  and  a51346a );
 a51351a <=( (not A200)  and  (not A199) );
 a51352a <=( A166  and  a51351a );
 a51353a <=( a51352a  and  a51347a );
 a51357a <=( (not A265)  and  A233 );
 a51358a <=( A232  and  a51357a );
 a51361a <=( (not A299)  and  (not A266) );
 a51364a <=( (not A302)  and  (not A301) );
 a51365a <=( a51364a  and  a51361a );
 a51366a <=( a51365a  and  a51358a );
 a51370a <=( A167  and  A169 );
 a51371a <=( (not A170)  and  a51370a );
 a51375a <=( (not A200)  and  (not A199) );
 a51376a <=( A166  and  a51375a );
 a51377a <=( a51376a  and  a51371a );
 a51381a <=( (not A236)  and  (not A235) );
 a51382a <=( (not A233)  and  a51381a );
 a51385a <=( A266  and  A265 );
 a51388a <=( (not A300)  and  A298 );
 a51389a <=( a51388a  and  a51385a );
 a51390a <=( a51389a  and  a51382a );
 a51394a <=( A167  and  A169 );
 a51395a <=( (not A170)  and  a51394a );
 a51399a <=( (not A200)  and  (not A199) );
 a51400a <=( A166  and  a51399a );
 a51401a <=( a51400a  and  a51395a );
 a51405a <=( (not A236)  and  (not A235) );
 a51406a <=( (not A233)  and  a51405a );
 a51409a <=( A266  and  A265 );
 a51412a <=( A299  and  A298 );
 a51413a <=( a51412a  and  a51409a );
 a51414a <=( a51413a  and  a51406a );
 a51418a <=( A167  and  A169 );
 a51419a <=( (not A170)  and  a51418a );
 a51423a <=( (not A200)  and  (not A199) );
 a51424a <=( A166  and  a51423a );
 a51425a <=( a51424a  and  a51419a );
 a51429a <=( (not A236)  and  (not A235) );
 a51430a <=( (not A233)  and  a51429a );
 a51433a <=( A266  and  A265 );
 a51436a <=( (not A299)  and  (not A298) );
 a51437a <=( a51436a  and  a51433a );
 a51438a <=( a51437a  and  a51430a );
 a51442a <=( A167  and  A169 );
 a51443a <=( (not A170)  and  a51442a );
 a51447a <=( (not A200)  and  (not A199) );
 a51448a <=( A166  and  a51447a );
 a51449a <=( a51448a  and  a51443a );
 a51453a <=( (not A236)  and  (not A235) );
 a51454a <=( (not A233)  and  a51453a );
 a51457a <=( (not A267)  and  (not A266) );
 a51460a <=( (not A300)  and  A298 );
 a51461a <=( a51460a  and  a51457a );
 a51462a <=( a51461a  and  a51454a );
 a51466a <=( A167  and  A169 );
 a51467a <=( (not A170)  and  a51466a );
 a51471a <=( (not A200)  and  (not A199) );
 a51472a <=( A166  and  a51471a );
 a51473a <=( a51472a  and  a51467a );
 a51477a <=( (not A236)  and  (not A235) );
 a51478a <=( (not A233)  and  a51477a );
 a51481a <=( (not A267)  and  (not A266) );
 a51484a <=( A299  and  A298 );
 a51485a <=( a51484a  and  a51481a );
 a51486a <=( a51485a  and  a51478a );
 a51490a <=( A167  and  A169 );
 a51491a <=( (not A170)  and  a51490a );
 a51495a <=( (not A200)  and  (not A199) );
 a51496a <=( A166  and  a51495a );
 a51497a <=( a51496a  and  a51491a );
 a51501a <=( (not A236)  and  (not A235) );
 a51502a <=( (not A233)  and  a51501a );
 a51505a <=( (not A267)  and  (not A266) );
 a51508a <=( (not A299)  and  (not A298) );
 a51509a <=( a51508a  and  a51505a );
 a51510a <=( a51509a  and  a51502a );
 a51514a <=( A167  and  A169 );
 a51515a <=( (not A170)  and  a51514a );
 a51519a <=( (not A200)  and  (not A199) );
 a51520a <=( A166  and  a51519a );
 a51521a <=( a51520a  and  a51515a );
 a51525a <=( (not A236)  and  (not A235) );
 a51526a <=( (not A233)  and  a51525a );
 a51529a <=( (not A266)  and  (not A265) );
 a51532a <=( (not A300)  and  A298 );
 a51533a <=( a51532a  and  a51529a );
 a51534a <=( a51533a  and  a51526a );
 a51538a <=( A167  and  A169 );
 a51539a <=( (not A170)  and  a51538a );
 a51543a <=( (not A200)  and  (not A199) );
 a51544a <=( A166  and  a51543a );
 a51545a <=( a51544a  and  a51539a );
 a51549a <=( (not A236)  and  (not A235) );
 a51550a <=( (not A233)  and  a51549a );
 a51553a <=( (not A266)  and  (not A265) );
 a51556a <=( A299  and  A298 );
 a51557a <=( a51556a  and  a51553a );
 a51558a <=( a51557a  and  a51550a );
 a51562a <=( A167  and  A169 );
 a51563a <=( (not A170)  and  a51562a );
 a51567a <=( (not A200)  and  (not A199) );
 a51568a <=( A166  and  a51567a );
 a51569a <=( a51568a  and  a51563a );
 a51573a <=( (not A236)  and  (not A235) );
 a51574a <=( (not A233)  and  a51573a );
 a51577a <=( (not A266)  and  (not A265) );
 a51580a <=( (not A299)  and  (not A298) );
 a51581a <=( a51580a  and  a51577a );
 a51582a <=( a51581a  and  a51574a );
 a51586a <=( A167  and  A169 );
 a51587a <=( (not A170)  and  a51586a );
 a51591a <=( (not A200)  and  (not A199) );
 a51592a <=( A166  and  a51591a );
 a51593a <=( a51592a  and  a51587a );
 a51597a <=( A265  and  (not A234) );
 a51598a <=( (not A233)  and  a51597a );
 a51601a <=( A298  and  A266 );
 a51604a <=( (not A302)  and  (not A301) );
 a51605a <=( a51604a  and  a51601a );
 a51606a <=( a51605a  and  a51598a );
 a51610a <=( A167  and  A169 );
 a51611a <=( (not A170)  and  a51610a );
 a51615a <=( (not A200)  and  (not A199) );
 a51616a <=( A166  and  a51615a );
 a51617a <=( a51616a  and  a51611a );
 a51621a <=( (not A266)  and  (not A234) );
 a51622a <=( (not A233)  and  a51621a );
 a51625a <=( (not A269)  and  (not A268) );
 a51628a <=( (not A300)  and  A298 );
 a51629a <=( a51628a  and  a51625a );
 a51630a <=( a51629a  and  a51622a );
 a51634a <=( A167  and  A169 );
 a51635a <=( (not A170)  and  a51634a );
 a51639a <=( (not A200)  and  (not A199) );
 a51640a <=( A166  and  a51639a );
 a51641a <=( a51640a  and  a51635a );
 a51645a <=( (not A266)  and  (not A234) );
 a51646a <=( (not A233)  and  a51645a );
 a51649a <=( (not A269)  and  (not A268) );
 a51652a <=( A299  and  A298 );
 a51653a <=( a51652a  and  a51649a );
 a51654a <=( a51653a  and  a51646a );
 a51658a <=( A167  and  A169 );
 a51659a <=( (not A170)  and  a51658a );
 a51663a <=( (not A200)  and  (not A199) );
 a51664a <=( A166  and  a51663a );
 a51665a <=( a51664a  and  a51659a );
 a51669a <=( (not A266)  and  (not A234) );
 a51670a <=( (not A233)  and  a51669a );
 a51673a <=( (not A269)  and  (not A268) );
 a51676a <=( (not A299)  and  (not A298) );
 a51677a <=( a51676a  and  a51673a );
 a51678a <=( a51677a  and  a51670a );
 a51682a <=( A167  and  A169 );
 a51683a <=( (not A170)  and  a51682a );
 a51687a <=( (not A200)  and  (not A199) );
 a51688a <=( A166  and  a51687a );
 a51689a <=( a51688a  and  a51683a );
 a51693a <=( (not A266)  and  (not A234) );
 a51694a <=( (not A233)  and  a51693a );
 a51697a <=( A298  and  (not A267) );
 a51700a <=( (not A302)  and  (not A301) );
 a51701a <=( a51700a  and  a51697a );
 a51702a <=( a51701a  and  a51694a );
 a51706a <=( A167  and  A169 );
 a51707a <=( (not A170)  and  a51706a );
 a51711a <=( (not A200)  and  (not A199) );
 a51712a <=( A166  and  a51711a );
 a51713a <=( a51712a  and  a51707a );
 a51717a <=( (not A265)  and  (not A234) );
 a51718a <=( (not A233)  and  a51717a );
 a51721a <=( A298  and  (not A266) );
 a51724a <=( (not A302)  and  (not A301) );
 a51725a <=( a51724a  and  a51721a );
 a51726a <=( a51725a  and  a51718a );
 a51730a <=( A167  and  A169 );
 a51731a <=( (not A170)  and  a51730a );
 a51735a <=( (not A200)  and  (not A199) );
 a51736a <=( A166  and  a51735a );
 a51737a <=( a51736a  and  a51731a );
 a51741a <=( A265  and  (not A233) );
 a51742a <=( (not A232)  and  a51741a );
 a51745a <=( A298  and  A266 );
 a51748a <=( (not A302)  and  (not A301) );
 a51749a <=( a51748a  and  a51745a );
 a51750a <=( a51749a  and  a51742a );
 a51754a <=( A167  and  A169 );
 a51755a <=( (not A170)  and  a51754a );
 a51759a <=( (not A200)  and  (not A199) );
 a51760a <=( A166  and  a51759a );
 a51761a <=( a51760a  and  a51755a );
 a51765a <=( (not A266)  and  (not A233) );
 a51766a <=( (not A232)  and  a51765a );
 a51769a <=( (not A269)  and  (not A268) );
 a51772a <=( (not A300)  and  A298 );
 a51773a <=( a51772a  and  a51769a );
 a51774a <=( a51773a  and  a51766a );
 a51778a <=( A167  and  A169 );
 a51779a <=( (not A170)  and  a51778a );
 a51783a <=( (not A200)  and  (not A199) );
 a51784a <=( A166  and  a51783a );
 a51785a <=( a51784a  and  a51779a );
 a51789a <=( (not A266)  and  (not A233) );
 a51790a <=( (not A232)  and  a51789a );
 a51793a <=( (not A269)  and  (not A268) );
 a51796a <=( A299  and  A298 );
 a51797a <=( a51796a  and  a51793a );
 a51798a <=( a51797a  and  a51790a );
 a51802a <=( A167  and  A169 );
 a51803a <=( (not A170)  and  a51802a );
 a51807a <=( (not A200)  and  (not A199) );
 a51808a <=( A166  and  a51807a );
 a51809a <=( a51808a  and  a51803a );
 a51813a <=( (not A266)  and  (not A233) );
 a51814a <=( (not A232)  and  a51813a );
 a51817a <=( (not A269)  and  (not A268) );
 a51820a <=( (not A299)  and  (not A298) );
 a51821a <=( a51820a  and  a51817a );
 a51822a <=( a51821a  and  a51814a );
 a51826a <=( A167  and  A169 );
 a51827a <=( (not A170)  and  a51826a );
 a51831a <=( (not A200)  and  (not A199) );
 a51832a <=( A166  and  a51831a );
 a51833a <=( a51832a  and  a51827a );
 a51837a <=( (not A266)  and  (not A233) );
 a51838a <=( (not A232)  and  a51837a );
 a51841a <=( A298  and  (not A267) );
 a51844a <=( (not A302)  and  (not A301) );
 a51845a <=( a51844a  and  a51841a );
 a51846a <=( a51845a  and  a51838a );
 a51850a <=( A167  and  A169 );
 a51851a <=( (not A170)  and  a51850a );
 a51855a <=( (not A200)  and  (not A199) );
 a51856a <=( A166  and  a51855a );
 a51857a <=( a51856a  and  a51851a );
 a51861a <=( (not A265)  and  (not A233) );
 a51862a <=( (not A232)  and  a51861a );
 a51865a <=( A298  and  (not A266) );
 a51868a <=( (not A302)  and  (not A301) );
 a51869a <=( a51868a  and  a51865a );
 a51870a <=( a51869a  and  a51862a );
 a51874a <=( (not A167)  and  A169 );
 a51875a <=( (not A170)  and  a51874a );
 a51879a <=( A200  and  A199 );
 a51880a <=( (not A166)  and  a51879a );
 a51881a <=( a51880a  and  a51875a );
 a51885a <=( A265  and  A233 );
 a51886a <=( A232  and  a51885a );
 a51889a <=( (not A269)  and  (not A268) );
 a51892a <=( (not A300)  and  (not A299) );
 a51893a <=( a51892a  and  a51889a );
 a51894a <=( a51893a  and  a51886a );
 a51898a <=( (not A167)  and  A169 );
 a51899a <=( (not A170)  and  a51898a );
 a51903a <=( A200  and  A199 );
 a51904a <=( (not A166)  and  a51903a );
 a51905a <=( a51904a  and  a51899a );
 a51909a <=( A265  and  A233 );
 a51910a <=( A232  and  a51909a );
 a51913a <=( (not A269)  and  (not A268) );
 a51916a <=( A299  and  A298 );
 a51917a <=( a51916a  and  a51913a );
 a51918a <=( a51917a  and  a51910a );
 a51922a <=( (not A167)  and  A169 );
 a51923a <=( (not A170)  and  a51922a );
 a51927a <=( A200  and  A199 );
 a51928a <=( (not A166)  and  a51927a );
 a51929a <=( a51928a  and  a51923a );
 a51933a <=( A265  and  A233 );
 a51934a <=( A232  and  a51933a );
 a51937a <=( (not A269)  and  (not A268) );
 a51940a <=( (not A299)  and  (not A298) );
 a51941a <=( a51940a  and  a51937a );
 a51942a <=( a51941a  and  a51934a );
 a51946a <=( (not A167)  and  A169 );
 a51947a <=( (not A170)  and  a51946a );
 a51951a <=( A200  and  A199 );
 a51952a <=( (not A166)  and  a51951a );
 a51953a <=( a51952a  and  a51947a );
 a51957a <=( A265  and  A233 );
 a51958a <=( A232  and  a51957a );
 a51961a <=( (not A299)  and  (not A267) );
 a51964a <=( (not A302)  and  (not A301) );
 a51965a <=( a51964a  and  a51961a );
 a51966a <=( a51965a  and  a51958a );
 a51970a <=( (not A167)  and  A169 );
 a51971a <=( (not A170)  and  a51970a );
 a51975a <=( A200  and  A199 );
 a51976a <=( (not A166)  and  a51975a );
 a51977a <=( a51976a  and  a51971a );
 a51981a <=( A265  and  A233 );
 a51982a <=( A232  and  a51981a );
 a51985a <=( (not A299)  and  A266 );
 a51988a <=( (not A302)  and  (not A301) );
 a51989a <=( a51988a  and  a51985a );
 a51990a <=( a51989a  and  a51982a );
 a51994a <=( (not A167)  and  A169 );
 a51995a <=( (not A170)  and  a51994a );
 a51999a <=( A200  and  A199 );
 a52000a <=( (not A166)  and  a51999a );
 a52001a <=( a52000a  and  a51995a );
 a52005a <=( (not A265)  and  A233 );
 a52006a <=( A232  and  a52005a );
 a52009a <=( (not A299)  and  (not A266) );
 a52012a <=( (not A302)  and  (not A301) );
 a52013a <=( a52012a  and  a52009a );
 a52014a <=( a52013a  and  a52006a );
 a52018a <=( (not A167)  and  A169 );
 a52019a <=( (not A170)  and  a52018a );
 a52023a <=( A200  and  A199 );
 a52024a <=( (not A166)  and  a52023a );
 a52025a <=( a52024a  and  a52019a );
 a52029a <=( (not A236)  and  (not A235) );
 a52030a <=( (not A233)  and  a52029a );
 a52033a <=( A266  and  A265 );
 a52036a <=( (not A300)  and  A298 );
 a52037a <=( a52036a  and  a52033a );
 a52038a <=( a52037a  and  a52030a );
 a52042a <=( (not A167)  and  A169 );
 a52043a <=( (not A170)  and  a52042a );
 a52047a <=( A200  and  A199 );
 a52048a <=( (not A166)  and  a52047a );
 a52049a <=( a52048a  and  a52043a );
 a52053a <=( (not A236)  and  (not A235) );
 a52054a <=( (not A233)  and  a52053a );
 a52057a <=( A266  and  A265 );
 a52060a <=( A299  and  A298 );
 a52061a <=( a52060a  and  a52057a );
 a52062a <=( a52061a  and  a52054a );
 a52066a <=( (not A167)  and  A169 );
 a52067a <=( (not A170)  and  a52066a );
 a52071a <=( A200  and  A199 );
 a52072a <=( (not A166)  and  a52071a );
 a52073a <=( a52072a  and  a52067a );
 a52077a <=( (not A236)  and  (not A235) );
 a52078a <=( (not A233)  and  a52077a );
 a52081a <=( A266  and  A265 );
 a52084a <=( (not A299)  and  (not A298) );
 a52085a <=( a52084a  and  a52081a );
 a52086a <=( a52085a  and  a52078a );
 a52090a <=( (not A167)  and  A169 );
 a52091a <=( (not A170)  and  a52090a );
 a52095a <=( A200  and  A199 );
 a52096a <=( (not A166)  and  a52095a );
 a52097a <=( a52096a  and  a52091a );
 a52101a <=( (not A236)  and  (not A235) );
 a52102a <=( (not A233)  and  a52101a );
 a52105a <=( (not A267)  and  (not A266) );
 a52108a <=( (not A300)  and  A298 );
 a52109a <=( a52108a  and  a52105a );
 a52110a <=( a52109a  and  a52102a );
 a52114a <=( (not A167)  and  A169 );
 a52115a <=( (not A170)  and  a52114a );
 a52119a <=( A200  and  A199 );
 a52120a <=( (not A166)  and  a52119a );
 a52121a <=( a52120a  and  a52115a );
 a52125a <=( (not A236)  and  (not A235) );
 a52126a <=( (not A233)  and  a52125a );
 a52129a <=( (not A267)  and  (not A266) );
 a52132a <=( A299  and  A298 );
 a52133a <=( a52132a  and  a52129a );
 a52134a <=( a52133a  and  a52126a );
 a52138a <=( (not A167)  and  A169 );
 a52139a <=( (not A170)  and  a52138a );
 a52143a <=( A200  and  A199 );
 a52144a <=( (not A166)  and  a52143a );
 a52145a <=( a52144a  and  a52139a );
 a52149a <=( (not A236)  and  (not A235) );
 a52150a <=( (not A233)  and  a52149a );
 a52153a <=( (not A267)  and  (not A266) );
 a52156a <=( (not A299)  and  (not A298) );
 a52157a <=( a52156a  and  a52153a );
 a52158a <=( a52157a  and  a52150a );
 a52162a <=( (not A167)  and  A169 );
 a52163a <=( (not A170)  and  a52162a );
 a52167a <=( A200  and  A199 );
 a52168a <=( (not A166)  and  a52167a );
 a52169a <=( a52168a  and  a52163a );
 a52173a <=( (not A236)  and  (not A235) );
 a52174a <=( (not A233)  and  a52173a );
 a52177a <=( (not A266)  and  (not A265) );
 a52180a <=( (not A300)  and  A298 );
 a52181a <=( a52180a  and  a52177a );
 a52182a <=( a52181a  and  a52174a );
 a52186a <=( (not A167)  and  A169 );
 a52187a <=( (not A170)  and  a52186a );
 a52191a <=( A200  and  A199 );
 a52192a <=( (not A166)  and  a52191a );
 a52193a <=( a52192a  and  a52187a );
 a52197a <=( (not A236)  and  (not A235) );
 a52198a <=( (not A233)  and  a52197a );
 a52201a <=( (not A266)  and  (not A265) );
 a52204a <=( A299  and  A298 );
 a52205a <=( a52204a  and  a52201a );
 a52206a <=( a52205a  and  a52198a );
 a52210a <=( (not A167)  and  A169 );
 a52211a <=( (not A170)  and  a52210a );
 a52215a <=( A200  and  A199 );
 a52216a <=( (not A166)  and  a52215a );
 a52217a <=( a52216a  and  a52211a );
 a52221a <=( (not A236)  and  (not A235) );
 a52222a <=( (not A233)  and  a52221a );
 a52225a <=( (not A266)  and  (not A265) );
 a52228a <=( (not A299)  and  (not A298) );
 a52229a <=( a52228a  and  a52225a );
 a52230a <=( a52229a  and  a52222a );
 a52234a <=( (not A167)  and  A169 );
 a52235a <=( (not A170)  and  a52234a );
 a52239a <=( A200  and  A199 );
 a52240a <=( (not A166)  and  a52239a );
 a52241a <=( a52240a  and  a52235a );
 a52245a <=( A265  and  (not A234) );
 a52246a <=( (not A233)  and  a52245a );
 a52249a <=( A298  and  A266 );
 a52252a <=( (not A302)  and  (not A301) );
 a52253a <=( a52252a  and  a52249a );
 a52254a <=( a52253a  and  a52246a );
 a52258a <=( (not A167)  and  A169 );
 a52259a <=( (not A170)  and  a52258a );
 a52263a <=( A200  and  A199 );
 a52264a <=( (not A166)  and  a52263a );
 a52265a <=( a52264a  and  a52259a );
 a52269a <=( (not A266)  and  (not A234) );
 a52270a <=( (not A233)  and  a52269a );
 a52273a <=( (not A269)  and  (not A268) );
 a52276a <=( (not A300)  and  A298 );
 a52277a <=( a52276a  and  a52273a );
 a52278a <=( a52277a  and  a52270a );
 a52282a <=( (not A167)  and  A169 );
 a52283a <=( (not A170)  and  a52282a );
 a52287a <=( A200  and  A199 );
 a52288a <=( (not A166)  and  a52287a );
 a52289a <=( a52288a  and  a52283a );
 a52293a <=( (not A266)  and  (not A234) );
 a52294a <=( (not A233)  and  a52293a );
 a52297a <=( (not A269)  and  (not A268) );
 a52300a <=( A299  and  A298 );
 a52301a <=( a52300a  and  a52297a );
 a52302a <=( a52301a  and  a52294a );
 a52306a <=( (not A167)  and  A169 );
 a52307a <=( (not A170)  and  a52306a );
 a52311a <=( A200  and  A199 );
 a52312a <=( (not A166)  and  a52311a );
 a52313a <=( a52312a  and  a52307a );
 a52317a <=( (not A266)  and  (not A234) );
 a52318a <=( (not A233)  and  a52317a );
 a52321a <=( (not A269)  and  (not A268) );
 a52324a <=( (not A299)  and  (not A298) );
 a52325a <=( a52324a  and  a52321a );
 a52326a <=( a52325a  and  a52318a );
 a52330a <=( (not A167)  and  A169 );
 a52331a <=( (not A170)  and  a52330a );
 a52335a <=( A200  and  A199 );
 a52336a <=( (not A166)  and  a52335a );
 a52337a <=( a52336a  and  a52331a );
 a52341a <=( (not A266)  and  (not A234) );
 a52342a <=( (not A233)  and  a52341a );
 a52345a <=( A298  and  (not A267) );
 a52348a <=( (not A302)  and  (not A301) );
 a52349a <=( a52348a  and  a52345a );
 a52350a <=( a52349a  and  a52342a );
 a52354a <=( (not A167)  and  A169 );
 a52355a <=( (not A170)  and  a52354a );
 a52359a <=( A200  and  A199 );
 a52360a <=( (not A166)  and  a52359a );
 a52361a <=( a52360a  and  a52355a );
 a52365a <=( (not A265)  and  (not A234) );
 a52366a <=( (not A233)  and  a52365a );
 a52369a <=( A298  and  (not A266) );
 a52372a <=( (not A302)  and  (not A301) );
 a52373a <=( a52372a  and  a52369a );
 a52374a <=( a52373a  and  a52366a );
 a52378a <=( (not A167)  and  A169 );
 a52379a <=( (not A170)  and  a52378a );
 a52383a <=( A200  and  A199 );
 a52384a <=( (not A166)  and  a52383a );
 a52385a <=( a52384a  and  a52379a );
 a52389a <=( A265  and  (not A233) );
 a52390a <=( (not A232)  and  a52389a );
 a52393a <=( A298  and  A266 );
 a52396a <=( (not A302)  and  (not A301) );
 a52397a <=( a52396a  and  a52393a );
 a52398a <=( a52397a  and  a52390a );
 a52402a <=( (not A167)  and  A169 );
 a52403a <=( (not A170)  and  a52402a );
 a52407a <=( A200  and  A199 );
 a52408a <=( (not A166)  and  a52407a );
 a52409a <=( a52408a  and  a52403a );
 a52413a <=( (not A266)  and  (not A233) );
 a52414a <=( (not A232)  and  a52413a );
 a52417a <=( (not A269)  and  (not A268) );
 a52420a <=( (not A300)  and  A298 );
 a52421a <=( a52420a  and  a52417a );
 a52422a <=( a52421a  and  a52414a );
 a52426a <=( (not A167)  and  A169 );
 a52427a <=( (not A170)  and  a52426a );
 a52431a <=( A200  and  A199 );
 a52432a <=( (not A166)  and  a52431a );
 a52433a <=( a52432a  and  a52427a );
 a52437a <=( (not A266)  and  (not A233) );
 a52438a <=( (not A232)  and  a52437a );
 a52441a <=( (not A269)  and  (not A268) );
 a52444a <=( A299  and  A298 );
 a52445a <=( a52444a  and  a52441a );
 a52446a <=( a52445a  and  a52438a );
 a52450a <=( (not A167)  and  A169 );
 a52451a <=( (not A170)  and  a52450a );
 a52455a <=( A200  and  A199 );
 a52456a <=( (not A166)  and  a52455a );
 a52457a <=( a52456a  and  a52451a );
 a52461a <=( (not A266)  and  (not A233) );
 a52462a <=( (not A232)  and  a52461a );
 a52465a <=( (not A269)  and  (not A268) );
 a52468a <=( (not A299)  and  (not A298) );
 a52469a <=( a52468a  and  a52465a );
 a52470a <=( a52469a  and  a52462a );
 a52474a <=( (not A167)  and  A169 );
 a52475a <=( (not A170)  and  a52474a );
 a52479a <=( A200  and  A199 );
 a52480a <=( (not A166)  and  a52479a );
 a52481a <=( a52480a  and  a52475a );
 a52485a <=( (not A266)  and  (not A233) );
 a52486a <=( (not A232)  and  a52485a );
 a52489a <=( A298  and  (not A267) );
 a52492a <=( (not A302)  and  (not A301) );
 a52493a <=( a52492a  and  a52489a );
 a52494a <=( a52493a  and  a52486a );
 a52498a <=( (not A167)  and  A169 );
 a52499a <=( (not A170)  and  a52498a );
 a52503a <=( A200  and  A199 );
 a52504a <=( (not A166)  and  a52503a );
 a52505a <=( a52504a  and  a52499a );
 a52509a <=( (not A265)  and  (not A233) );
 a52510a <=( (not A232)  and  a52509a );
 a52513a <=( A298  and  (not A266) );
 a52516a <=( (not A302)  and  (not A301) );
 a52517a <=( a52516a  and  a52513a );
 a52518a <=( a52517a  and  a52510a );
 a52522a <=( (not A167)  and  A169 );
 a52523a <=( (not A170)  and  a52522a );
 a52527a <=( (not A202)  and  (not A200) );
 a52528a <=( (not A166)  and  a52527a );
 a52529a <=( a52528a  and  a52523a );
 a52533a <=( A233  and  A232 );
 a52534a <=( (not A203)  and  a52533a );
 a52537a <=( (not A267)  and  A265 );
 a52540a <=( (not A300)  and  (not A299) );
 a52541a <=( a52540a  and  a52537a );
 a52542a <=( a52541a  and  a52534a );
 a52546a <=( (not A167)  and  A169 );
 a52547a <=( (not A170)  and  a52546a );
 a52551a <=( (not A202)  and  (not A200) );
 a52552a <=( (not A166)  and  a52551a );
 a52553a <=( a52552a  and  a52547a );
 a52557a <=( A233  and  A232 );
 a52558a <=( (not A203)  and  a52557a );
 a52561a <=( (not A267)  and  A265 );
 a52564a <=( A299  and  A298 );
 a52565a <=( a52564a  and  a52561a );
 a52566a <=( a52565a  and  a52558a );
 a52570a <=( (not A167)  and  A169 );
 a52571a <=( (not A170)  and  a52570a );
 a52575a <=( (not A202)  and  (not A200) );
 a52576a <=( (not A166)  and  a52575a );
 a52577a <=( a52576a  and  a52571a );
 a52581a <=( A233  and  A232 );
 a52582a <=( (not A203)  and  a52581a );
 a52585a <=( (not A267)  and  A265 );
 a52588a <=( (not A299)  and  (not A298) );
 a52589a <=( a52588a  and  a52585a );
 a52590a <=( a52589a  and  a52582a );
 a52594a <=( (not A167)  and  A169 );
 a52595a <=( (not A170)  and  a52594a );
 a52599a <=( (not A202)  and  (not A200) );
 a52600a <=( (not A166)  and  a52599a );
 a52601a <=( a52600a  and  a52595a );
 a52605a <=( A233  and  A232 );
 a52606a <=( (not A203)  and  a52605a );
 a52609a <=( A266  and  A265 );
 a52612a <=( (not A300)  and  (not A299) );
 a52613a <=( a52612a  and  a52609a );
 a52614a <=( a52613a  and  a52606a );
 a52618a <=( (not A167)  and  A169 );
 a52619a <=( (not A170)  and  a52618a );
 a52623a <=( (not A202)  and  (not A200) );
 a52624a <=( (not A166)  and  a52623a );
 a52625a <=( a52624a  and  a52619a );
 a52629a <=( A233  and  A232 );
 a52630a <=( (not A203)  and  a52629a );
 a52633a <=( A266  and  A265 );
 a52636a <=( A299  and  A298 );
 a52637a <=( a52636a  and  a52633a );
 a52638a <=( a52637a  and  a52630a );
 a52642a <=( (not A167)  and  A169 );
 a52643a <=( (not A170)  and  a52642a );
 a52647a <=( (not A202)  and  (not A200) );
 a52648a <=( (not A166)  and  a52647a );
 a52649a <=( a52648a  and  a52643a );
 a52653a <=( A233  and  A232 );
 a52654a <=( (not A203)  and  a52653a );
 a52657a <=( A266  and  A265 );
 a52660a <=( (not A299)  and  (not A298) );
 a52661a <=( a52660a  and  a52657a );
 a52662a <=( a52661a  and  a52654a );
 a52666a <=( (not A167)  and  A169 );
 a52667a <=( (not A170)  and  a52666a );
 a52671a <=( (not A202)  and  (not A200) );
 a52672a <=( (not A166)  and  a52671a );
 a52673a <=( a52672a  and  a52667a );
 a52677a <=( A233  and  A232 );
 a52678a <=( (not A203)  and  a52677a );
 a52681a <=( (not A266)  and  (not A265) );
 a52684a <=( (not A300)  and  (not A299) );
 a52685a <=( a52684a  and  a52681a );
 a52686a <=( a52685a  and  a52678a );
 a52690a <=( (not A167)  and  A169 );
 a52691a <=( (not A170)  and  a52690a );
 a52695a <=( (not A202)  and  (not A200) );
 a52696a <=( (not A166)  and  a52695a );
 a52697a <=( a52696a  and  a52691a );
 a52701a <=( A233  and  A232 );
 a52702a <=( (not A203)  and  a52701a );
 a52705a <=( (not A266)  and  (not A265) );
 a52708a <=( A299  and  A298 );
 a52709a <=( a52708a  and  a52705a );
 a52710a <=( a52709a  and  a52702a );
 a52714a <=( (not A167)  and  A169 );
 a52715a <=( (not A170)  and  a52714a );
 a52719a <=( (not A202)  and  (not A200) );
 a52720a <=( (not A166)  and  a52719a );
 a52721a <=( a52720a  and  a52715a );
 a52725a <=( A233  and  A232 );
 a52726a <=( (not A203)  and  a52725a );
 a52729a <=( (not A266)  and  (not A265) );
 a52732a <=( (not A299)  and  (not A298) );
 a52733a <=( a52732a  and  a52729a );
 a52734a <=( a52733a  and  a52726a );
 a52738a <=( (not A167)  and  A169 );
 a52739a <=( (not A170)  and  a52738a );
 a52743a <=( (not A202)  and  (not A200) );
 a52744a <=( (not A166)  and  a52743a );
 a52745a <=( a52744a  and  a52739a );
 a52749a <=( A233  and  (not A232) );
 a52750a <=( (not A203)  and  a52749a );
 a52753a <=( (not A299)  and  A298 );
 a52756a <=( A301  and  A300 );
 a52757a <=( a52756a  and  a52753a );
 a52758a <=( a52757a  and  a52750a );
 a52762a <=( (not A167)  and  A169 );
 a52763a <=( (not A170)  and  a52762a );
 a52767a <=( (not A202)  and  (not A200) );
 a52768a <=( (not A166)  and  a52767a );
 a52769a <=( a52768a  and  a52763a );
 a52773a <=( A233  and  (not A232) );
 a52774a <=( (not A203)  and  a52773a );
 a52777a <=( (not A299)  and  A298 );
 a52780a <=( A302  and  A300 );
 a52781a <=( a52780a  and  a52777a );
 a52782a <=( a52781a  and  a52774a );
 a52786a <=( (not A167)  and  A169 );
 a52787a <=( (not A170)  and  a52786a );
 a52791a <=( (not A202)  and  (not A200) );
 a52792a <=( (not A166)  and  a52791a );
 a52793a <=( a52792a  and  a52787a );
 a52797a <=( A233  and  (not A232) );
 a52798a <=( (not A203)  and  a52797a );
 a52801a <=( (not A266)  and  A265 );
 a52804a <=( A268  and  A267 );
 a52805a <=( a52804a  and  a52801a );
 a52806a <=( a52805a  and  a52798a );
 a52810a <=( (not A167)  and  A169 );
 a52811a <=( (not A170)  and  a52810a );
 a52815a <=( (not A202)  and  (not A200) );
 a52816a <=( (not A166)  and  a52815a );
 a52817a <=( a52816a  and  a52811a );
 a52821a <=( A233  and  (not A232) );
 a52822a <=( (not A203)  and  a52821a );
 a52825a <=( (not A266)  and  A265 );
 a52828a <=( A269  and  A267 );
 a52829a <=( a52828a  and  a52825a );
 a52830a <=( a52829a  and  a52822a );
 a52834a <=( (not A167)  and  A169 );
 a52835a <=( (not A170)  and  a52834a );
 a52839a <=( (not A202)  and  (not A200) );
 a52840a <=( (not A166)  and  a52839a );
 a52841a <=( a52840a  and  a52835a );
 a52845a <=( (not A234)  and  (not A233) );
 a52846a <=( (not A203)  and  a52845a );
 a52849a <=( A266  and  A265 );
 a52852a <=( (not A300)  and  A298 );
 a52853a <=( a52852a  and  a52849a );
 a52854a <=( a52853a  and  a52846a );
 a52858a <=( (not A167)  and  A169 );
 a52859a <=( (not A170)  and  a52858a );
 a52863a <=( (not A202)  and  (not A200) );
 a52864a <=( (not A166)  and  a52863a );
 a52865a <=( a52864a  and  a52859a );
 a52869a <=( (not A234)  and  (not A233) );
 a52870a <=( (not A203)  and  a52869a );
 a52873a <=( A266  and  A265 );
 a52876a <=( A299  and  A298 );
 a52877a <=( a52876a  and  a52873a );
 a52878a <=( a52877a  and  a52870a );
 a52882a <=( (not A167)  and  A169 );
 a52883a <=( (not A170)  and  a52882a );
 a52887a <=( (not A202)  and  (not A200) );
 a52888a <=( (not A166)  and  a52887a );
 a52889a <=( a52888a  and  a52883a );
 a52893a <=( (not A234)  and  (not A233) );
 a52894a <=( (not A203)  and  a52893a );
 a52897a <=( A266  and  A265 );
 a52900a <=( (not A299)  and  (not A298) );
 a52901a <=( a52900a  and  a52897a );
 a52902a <=( a52901a  and  a52894a );
 a52906a <=( (not A167)  and  A169 );
 a52907a <=( (not A170)  and  a52906a );
 a52911a <=( (not A202)  and  (not A200) );
 a52912a <=( (not A166)  and  a52911a );
 a52913a <=( a52912a  and  a52907a );
 a52917a <=( (not A234)  and  (not A233) );
 a52918a <=( (not A203)  and  a52917a );
 a52921a <=( (not A267)  and  (not A266) );
 a52924a <=( (not A300)  and  A298 );
 a52925a <=( a52924a  and  a52921a );
 a52926a <=( a52925a  and  a52918a );
 a52930a <=( (not A167)  and  A169 );
 a52931a <=( (not A170)  and  a52930a );
 a52935a <=( (not A202)  and  (not A200) );
 a52936a <=( (not A166)  and  a52935a );
 a52937a <=( a52936a  and  a52931a );
 a52941a <=( (not A234)  and  (not A233) );
 a52942a <=( (not A203)  and  a52941a );
 a52945a <=( (not A267)  and  (not A266) );
 a52948a <=( A299  and  A298 );
 a52949a <=( a52948a  and  a52945a );
 a52950a <=( a52949a  and  a52942a );
 a52954a <=( (not A167)  and  A169 );
 a52955a <=( (not A170)  and  a52954a );
 a52959a <=( (not A202)  and  (not A200) );
 a52960a <=( (not A166)  and  a52959a );
 a52961a <=( a52960a  and  a52955a );
 a52965a <=( (not A234)  and  (not A233) );
 a52966a <=( (not A203)  and  a52965a );
 a52969a <=( (not A267)  and  (not A266) );
 a52972a <=( (not A299)  and  (not A298) );
 a52973a <=( a52972a  and  a52969a );
 a52974a <=( a52973a  and  a52966a );
 a52978a <=( (not A167)  and  A169 );
 a52979a <=( (not A170)  and  a52978a );
 a52983a <=( (not A202)  and  (not A200) );
 a52984a <=( (not A166)  and  a52983a );
 a52985a <=( a52984a  and  a52979a );
 a52989a <=( (not A234)  and  (not A233) );
 a52990a <=( (not A203)  and  a52989a );
 a52993a <=( (not A266)  and  (not A265) );
 a52996a <=( (not A300)  and  A298 );
 a52997a <=( a52996a  and  a52993a );
 a52998a <=( a52997a  and  a52990a );
 a53002a <=( (not A167)  and  A169 );
 a53003a <=( (not A170)  and  a53002a );
 a53007a <=( (not A202)  and  (not A200) );
 a53008a <=( (not A166)  and  a53007a );
 a53009a <=( a53008a  and  a53003a );
 a53013a <=( (not A234)  and  (not A233) );
 a53014a <=( (not A203)  and  a53013a );
 a53017a <=( (not A266)  and  (not A265) );
 a53020a <=( A299  and  A298 );
 a53021a <=( a53020a  and  a53017a );
 a53022a <=( a53021a  and  a53014a );
 a53026a <=( (not A167)  and  A169 );
 a53027a <=( (not A170)  and  a53026a );
 a53031a <=( (not A202)  and  (not A200) );
 a53032a <=( (not A166)  and  a53031a );
 a53033a <=( a53032a  and  a53027a );
 a53037a <=( (not A234)  and  (not A233) );
 a53038a <=( (not A203)  and  a53037a );
 a53041a <=( (not A266)  and  (not A265) );
 a53044a <=( (not A299)  and  (not A298) );
 a53045a <=( a53044a  and  a53041a );
 a53046a <=( a53045a  and  a53038a );
 a53050a <=( (not A167)  and  A169 );
 a53051a <=( (not A170)  and  a53050a );
 a53055a <=( (not A202)  and  (not A200) );
 a53056a <=( (not A166)  and  a53055a );
 a53057a <=( a53056a  and  a53051a );
 a53061a <=( (not A233)  and  A232 );
 a53062a <=( (not A203)  and  a53061a );
 a53065a <=( A235  and  A234 );
 a53068a <=( A299  and  (not A298) );
 a53069a <=( a53068a  and  a53065a );
 a53070a <=( a53069a  and  a53062a );
 a53074a <=( (not A167)  and  A169 );
 a53075a <=( (not A170)  and  a53074a );
 a53079a <=( (not A202)  and  (not A200) );
 a53080a <=( (not A166)  and  a53079a );
 a53081a <=( a53080a  and  a53075a );
 a53085a <=( (not A233)  and  A232 );
 a53086a <=( (not A203)  and  a53085a );
 a53089a <=( A235  and  A234 );
 a53092a <=( A266  and  (not A265) );
 a53093a <=( a53092a  and  a53089a );
 a53094a <=( a53093a  and  a53086a );
 a53098a <=( (not A167)  and  A169 );
 a53099a <=( (not A170)  and  a53098a );
 a53103a <=( (not A202)  and  (not A200) );
 a53104a <=( (not A166)  and  a53103a );
 a53105a <=( a53104a  and  a53099a );
 a53109a <=( (not A233)  and  A232 );
 a53110a <=( (not A203)  and  a53109a );
 a53113a <=( A236  and  A234 );
 a53116a <=( A299  and  (not A298) );
 a53117a <=( a53116a  and  a53113a );
 a53118a <=( a53117a  and  a53110a );
 a53122a <=( (not A167)  and  A169 );
 a53123a <=( (not A170)  and  a53122a );
 a53127a <=( (not A202)  and  (not A200) );
 a53128a <=( (not A166)  and  a53127a );
 a53129a <=( a53128a  and  a53123a );
 a53133a <=( (not A233)  and  A232 );
 a53134a <=( (not A203)  and  a53133a );
 a53137a <=( A236  and  A234 );
 a53140a <=( A266  and  (not A265) );
 a53141a <=( a53140a  and  a53137a );
 a53142a <=( a53141a  and  a53134a );
 a53146a <=( (not A167)  and  A169 );
 a53147a <=( (not A170)  and  a53146a );
 a53151a <=( (not A202)  and  (not A200) );
 a53152a <=( (not A166)  and  a53151a );
 a53153a <=( a53152a  and  a53147a );
 a53157a <=( (not A233)  and  (not A232) );
 a53158a <=( (not A203)  and  a53157a );
 a53161a <=( A266  and  A265 );
 a53164a <=( (not A300)  and  A298 );
 a53165a <=( a53164a  and  a53161a );
 a53166a <=( a53165a  and  a53158a );
 a53170a <=( (not A167)  and  A169 );
 a53171a <=( (not A170)  and  a53170a );
 a53175a <=( (not A202)  and  (not A200) );
 a53176a <=( (not A166)  and  a53175a );
 a53177a <=( a53176a  and  a53171a );
 a53181a <=( (not A233)  and  (not A232) );
 a53182a <=( (not A203)  and  a53181a );
 a53185a <=( A266  and  A265 );
 a53188a <=( A299  and  A298 );
 a53189a <=( a53188a  and  a53185a );
 a53190a <=( a53189a  and  a53182a );
 a53194a <=( (not A167)  and  A169 );
 a53195a <=( (not A170)  and  a53194a );
 a53199a <=( (not A202)  and  (not A200) );
 a53200a <=( (not A166)  and  a53199a );
 a53201a <=( a53200a  and  a53195a );
 a53205a <=( (not A233)  and  (not A232) );
 a53206a <=( (not A203)  and  a53205a );
 a53209a <=( A266  and  A265 );
 a53212a <=( (not A299)  and  (not A298) );
 a53213a <=( a53212a  and  a53209a );
 a53214a <=( a53213a  and  a53206a );
 a53218a <=( (not A167)  and  A169 );
 a53219a <=( (not A170)  and  a53218a );
 a53223a <=( (not A202)  and  (not A200) );
 a53224a <=( (not A166)  and  a53223a );
 a53225a <=( a53224a  and  a53219a );
 a53229a <=( (not A233)  and  (not A232) );
 a53230a <=( (not A203)  and  a53229a );
 a53233a <=( (not A267)  and  (not A266) );
 a53236a <=( (not A300)  and  A298 );
 a53237a <=( a53236a  and  a53233a );
 a53238a <=( a53237a  and  a53230a );
 a53242a <=( (not A167)  and  A169 );
 a53243a <=( (not A170)  and  a53242a );
 a53247a <=( (not A202)  and  (not A200) );
 a53248a <=( (not A166)  and  a53247a );
 a53249a <=( a53248a  and  a53243a );
 a53253a <=( (not A233)  and  (not A232) );
 a53254a <=( (not A203)  and  a53253a );
 a53257a <=( (not A267)  and  (not A266) );
 a53260a <=( A299  and  A298 );
 a53261a <=( a53260a  and  a53257a );
 a53262a <=( a53261a  and  a53254a );
 a53266a <=( (not A167)  and  A169 );
 a53267a <=( (not A170)  and  a53266a );
 a53271a <=( (not A202)  and  (not A200) );
 a53272a <=( (not A166)  and  a53271a );
 a53273a <=( a53272a  and  a53267a );
 a53277a <=( (not A233)  and  (not A232) );
 a53278a <=( (not A203)  and  a53277a );
 a53281a <=( (not A267)  and  (not A266) );
 a53284a <=( (not A299)  and  (not A298) );
 a53285a <=( a53284a  and  a53281a );
 a53286a <=( a53285a  and  a53278a );
 a53290a <=( (not A167)  and  A169 );
 a53291a <=( (not A170)  and  a53290a );
 a53295a <=( (not A202)  and  (not A200) );
 a53296a <=( (not A166)  and  a53295a );
 a53297a <=( a53296a  and  a53291a );
 a53301a <=( (not A233)  and  (not A232) );
 a53302a <=( (not A203)  and  a53301a );
 a53305a <=( (not A266)  and  (not A265) );
 a53308a <=( (not A300)  and  A298 );
 a53309a <=( a53308a  and  a53305a );
 a53310a <=( a53309a  and  a53302a );
 a53314a <=( (not A167)  and  A169 );
 a53315a <=( (not A170)  and  a53314a );
 a53319a <=( (not A202)  and  (not A200) );
 a53320a <=( (not A166)  and  a53319a );
 a53321a <=( a53320a  and  a53315a );
 a53325a <=( (not A233)  and  (not A232) );
 a53326a <=( (not A203)  and  a53325a );
 a53329a <=( (not A266)  and  (not A265) );
 a53332a <=( A299  and  A298 );
 a53333a <=( a53332a  and  a53329a );
 a53334a <=( a53333a  and  a53326a );
 a53338a <=( (not A167)  and  A169 );
 a53339a <=( (not A170)  and  a53338a );
 a53343a <=( (not A202)  and  (not A200) );
 a53344a <=( (not A166)  and  a53343a );
 a53345a <=( a53344a  and  a53339a );
 a53349a <=( (not A233)  and  (not A232) );
 a53350a <=( (not A203)  and  a53349a );
 a53353a <=( (not A266)  and  (not A265) );
 a53356a <=( (not A299)  and  (not A298) );
 a53357a <=( a53356a  and  a53353a );
 a53358a <=( a53357a  and  a53350a );
 a53362a <=( (not A167)  and  A169 );
 a53363a <=( (not A170)  and  a53362a );
 a53367a <=( (not A201)  and  (not A200) );
 a53368a <=( (not A166)  and  a53367a );
 a53369a <=( a53368a  and  a53363a );
 a53373a <=( A265  and  A233 );
 a53374a <=( A232  and  a53373a );
 a53377a <=( (not A269)  and  (not A268) );
 a53380a <=( (not A300)  and  (not A299) );
 a53381a <=( a53380a  and  a53377a );
 a53382a <=( a53381a  and  a53374a );
 a53386a <=( (not A167)  and  A169 );
 a53387a <=( (not A170)  and  a53386a );
 a53391a <=( (not A201)  and  (not A200) );
 a53392a <=( (not A166)  and  a53391a );
 a53393a <=( a53392a  and  a53387a );
 a53397a <=( A265  and  A233 );
 a53398a <=( A232  and  a53397a );
 a53401a <=( (not A269)  and  (not A268) );
 a53404a <=( A299  and  A298 );
 a53405a <=( a53404a  and  a53401a );
 a53406a <=( a53405a  and  a53398a );
 a53410a <=( (not A167)  and  A169 );
 a53411a <=( (not A170)  and  a53410a );
 a53415a <=( (not A201)  and  (not A200) );
 a53416a <=( (not A166)  and  a53415a );
 a53417a <=( a53416a  and  a53411a );
 a53421a <=( A265  and  A233 );
 a53422a <=( A232  and  a53421a );
 a53425a <=( (not A269)  and  (not A268) );
 a53428a <=( (not A299)  and  (not A298) );
 a53429a <=( a53428a  and  a53425a );
 a53430a <=( a53429a  and  a53422a );
 a53434a <=( (not A167)  and  A169 );
 a53435a <=( (not A170)  and  a53434a );
 a53439a <=( (not A201)  and  (not A200) );
 a53440a <=( (not A166)  and  a53439a );
 a53441a <=( a53440a  and  a53435a );
 a53445a <=( A265  and  A233 );
 a53446a <=( A232  and  a53445a );
 a53449a <=( (not A299)  and  (not A267) );
 a53452a <=( (not A302)  and  (not A301) );
 a53453a <=( a53452a  and  a53449a );
 a53454a <=( a53453a  and  a53446a );
 a53458a <=( (not A167)  and  A169 );
 a53459a <=( (not A170)  and  a53458a );
 a53463a <=( (not A201)  and  (not A200) );
 a53464a <=( (not A166)  and  a53463a );
 a53465a <=( a53464a  and  a53459a );
 a53469a <=( A265  and  A233 );
 a53470a <=( A232  and  a53469a );
 a53473a <=( (not A299)  and  A266 );
 a53476a <=( (not A302)  and  (not A301) );
 a53477a <=( a53476a  and  a53473a );
 a53478a <=( a53477a  and  a53470a );
 a53482a <=( (not A167)  and  A169 );
 a53483a <=( (not A170)  and  a53482a );
 a53487a <=( (not A201)  and  (not A200) );
 a53488a <=( (not A166)  and  a53487a );
 a53489a <=( a53488a  and  a53483a );
 a53493a <=( (not A265)  and  A233 );
 a53494a <=( A232  and  a53493a );
 a53497a <=( (not A299)  and  (not A266) );
 a53500a <=( (not A302)  and  (not A301) );
 a53501a <=( a53500a  and  a53497a );
 a53502a <=( a53501a  and  a53494a );
 a53506a <=( (not A167)  and  A169 );
 a53507a <=( (not A170)  and  a53506a );
 a53511a <=( (not A201)  and  (not A200) );
 a53512a <=( (not A166)  and  a53511a );
 a53513a <=( a53512a  and  a53507a );
 a53517a <=( (not A236)  and  (not A235) );
 a53518a <=( (not A233)  and  a53517a );
 a53521a <=( A266  and  A265 );
 a53524a <=( (not A300)  and  A298 );
 a53525a <=( a53524a  and  a53521a );
 a53526a <=( a53525a  and  a53518a );
 a53530a <=( (not A167)  and  A169 );
 a53531a <=( (not A170)  and  a53530a );
 a53535a <=( (not A201)  and  (not A200) );
 a53536a <=( (not A166)  and  a53535a );
 a53537a <=( a53536a  and  a53531a );
 a53541a <=( (not A236)  and  (not A235) );
 a53542a <=( (not A233)  and  a53541a );
 a53545a <=( A266  and  A265 );
 a53548a <=( A299  and  A298 );
 a53549a <=( a53548a  and  a53545a );
 a53550a <=( a53549a  and  a53542a );
 a53554a <=( (not A167)  and  A169 );
 a53555a <=( (not A170)  and  a53554a );
 a53559a <=( (not A201)  and  (not A200) );
 a53560a <=( (not A166)  and  a53559a );
 a53561a <=( a53560a  and  a53555a );
 a53565a <=( (not A236)  and  (not A235) );
 a53566a <=( (not A233)  and  a53565a );
 a53569a <=( A266  and  A265 );
 a53572a <=( (not A299)  and  (not A298) );
 a53573a <=( a53572a  and  a53569a );
 a53574a <=( a53573a  and  a53566a );
 a53578a <=( (not A167)  and  A169 );
 a53579a <=( (not A170)  and  a53578a );
 a53583a <=( (not A201)  and  (not A200) );
 a53584a <=( (not A166)  and  a53583a );
 a53585a <=( a53584a  and  a53579a );
 a53589a <=( (not A236)  and  (not A235) );
 a53590a <=( (not A233)  and  a53589a );
 a53593a <=( (not A267)  and  (not A266) );
 a53596a <=( (not A300)  and  A298 );
 a53597a <=( a53596a  and  a53593a );
 a53598a <=( a53597a  and  a53590a );
 a53602a <=( (not A167)  and  A169 );
 a53603a <=( (not A170)  and  a53602a );
 a53607a <=( (not A201)  and  (not A200) );
 a53608a <=( (not A166)  and  a53607a );
 a53609a <=( a53608a  and  a53603a );
 a53613a <=( (not A236)  and  (not A235) );
 a53614a <=( (not A233)  and  a53613a );
 a53617a <=( (not A267)  and  (not A266) );
 a53620a <=( A299  and  A298 );
 a53621a <=( a53620a  and  a53617a );
 a53622a <=( a53621a  and  a53614a );
 a53626a <=( (not A167)  and  A169 );
 a53627a <=( (not A170)  and  a53626a );
 a53631a <=( (not A201)  and  (not A200) );
 a53632a <=( (not A166)  and  a53631a );
 a53633a <=( a53632a  and  a53627a );
 a53637a <=( (not A236)  and  (not A235) );
 a53638a <=( (not A233)  and  a53637a );
 a53641a <=( (not A267)  and  (not A266) );
 a53644a <=( (not A299)  and  (not A298) );
 a53645a <=( a53644a  and  a53641a );
 a53646a <=( a53645a  and  a53638a );
 a53650a <=( (not A167)  and  A169 );
 a53651a <=( (not A170)  and  a53650a );
 a53655a <=( (not A201)  and  (not A200) );
 a53656a <=( (not A166)  and  a53655a );
 a53657a <=( a53656a  and  a53651a );
 a53661a <=( (not A236)  and  (not A235) );
 a53662a <=( (not A233)  and  a53661a );
 a53665a <=( (not A266)  and  (not A265) );
 a53668a <=( (not A300)  and  A298 );
 a53669a <=( a53668a  and  a53665a );
 a53670a <=( a53669a  and  a53662a );
 a53674a <=( (not A167)  and  A169 );
 a53675a <=( (not A170)  and  a53674a );
 a53679a <=( (not A201)  and  (not A200) );
 a53680a <=( (not A166)  and  a53679a );
 a53681a <=( a53680a  and  a53675a );
 a53685a <=( (not A236)  and  (not A235) );
 a53686a <=( (not A233)  and  a53685a );
 a53689a <=( (not A266)  and  (not A265) );
 a53692a <=( A299  and  A298 );
 a53693a <=( a53692a  and  a53689a );
 a53694a <=( a53693a  and  a53686a );
 a53698a <=( (not A167)  and  A169 );
 a53699a <=( (not A170)  and  a53698a );
 a53703a <=( (not A201)  and  (not A200) );
 a53704a <=( (not A166)  and  a53703a );
 a53705a <=( a53704a  and  a53699a );
 a53709a <=( (not A236)  and  (not A235) );
 a53710a <=( (not A233)  and  a53709a );
 a53713a <=( (not A266)  and  (not A265) );
 a53716a <=( (not A299)  and  (not A298) );
 a53717a <=( a53716a  and  a53713a );
 a53718a <=( a53717a  and  a53710a );
 a53722a <=( (not A167)  and  A169 );
 a53723a <=( (not A170)  and  a53722a );
 a53727a <=( (not A201)  and  (not A200) );
 a53728a <=( (not A166)  and  a53727a );
 a53729a <=( a53728a  and  a53723a );
 a53733a <=( A265  and  (not A234) );
 a53734a <=( (not A233)  and  a53733a );
 a53737a <=( A298  and  A266 );
 a53740a <=( (not A302)  and  (not A301) );
 a53741a <=( a53740a  and  a53737a );
 a53742a <=( a53741a  and  a53734a );
 a53746a <=( (not A167)  and  A169 );
 a53747a <=( (not A170)  and  a53746a );
 a53751a <=( (not A201)  and  (not A200) );
 a53752a <=( (not A166)  and  a53751a );
 a53753a <=( a53752a  and  a53747a );
 a53757a <=( (not A266)  and  (not A234) );
 a53758a <=( (not A233)  and  a53757a );
 a53761a <=( (not A269)  and  (not A268) );
 a53764a <=( (not A300)  and  A298 );
 a53765a <=( a53764a  and  a53761a );
 a53766a <=( a53765a  and  a53758a );
 a53770a <=( (not A167)  and  A169 );
 a53771a <=( (not A170)  and  a53770a );
 a53775a <=( (not A201)  and  (not A200) );
 a53776a <=( (not A166)  and  a53775a );
 a53777a <=( a53776a  and  a53771a );
 a53781a <=( (not A266)  and  (not A234) );
 a53782a <=( (not A233)  and  a53781a );
 a53785a <=( (not A269)  and  (not A268) );
 a53788a <=( A299  and  A298 );
 a53789a <=( a53788a  and  a53785a );
 a53790a <=( a53789a  and  a53782a );
 a53794a <=( (not A167)  and  A169 );
 a53795a <=( (not A170)  and  a53794a );
 a53799a <=( (not A201)  and  (not A200) );
 a53800a <=( (not A166)  and  a53799a );
 a53801a <=( a53800a  and  a53795a );
 a53805a <=( (not A266)  and  (not A234) );
 a53806a <=( (not A233)  and  a53805a );
 a53809a <=( (not A269)  and  (not A268) );
 a53812a <=( (not A299)  and  (not A298) );
 a53813a <=( a53812a  and  a53809a );
 a53814a <=( a53813a  and  a53806a );
 a53818a <=( (not A167)  and  A169 );
 a53819a <=( (not A170)  and  a53818a );
 a53823a <=( (not A201)  and  (not A200) );
 a53824a <=( (not A166)  and  a53823a );
 a53825a <=( a53824a  and  a53819a );
 a53829a <=( (not A266)  and  (not A234) );
 a53830a <=( (not A233)  and  a53829a );
 a53833a <=( A298  and  (not A267) );
 a53836a <=( (not A302)  and  (not A301) );
 a53837a <=( a53836a  and  a53833a );
 a53838a <=( a53837a  and  a53830a );
 a53842a <=( (not A167)  and  A169 );
 a53843a <=( (not A170)  and  a53842a );
 a53847a <=( (not A201)  and  (not A200) );
 a53848a <=( (not A166)  and  a53847a );
 a53849a <=( a53848a  and  a53843a );
 a53853a <=( (not A265)  and  (not A234) );
 a53854a <=( (not A233)  and  a53853a );
 a53857a <=( A298  and  (not A266) );
 a53860a <=( (not A302)  and  (not A301) );
 a53861a <=( a53860a  and  a53857a );
 a53862a <=( a53861a  and  a53854a );
 a53866a <=( (not A167)  and  A169 );
 a53867a <=( (not A170)  and  a53866a );
 a53871a <=( (not A201)  and  (not A200) );
 a53872a <=( (not A166)  and  a53871a );
 a53873a <=( a53872a  and  a53867a );
 a53877a <=( A265  and  (not A233) );
 a53878a <=( (not A232)  and  a53877a );
 a53881a <=( A298  and  A266 );
 a53884a <=( (not A302)  and  (not A301) );
 a53885a <=( a53884a  and  a53881a );
 a53886a <=( a53885a  and  a53878a );
 a53890a <=( (not A167)  and  A169 );
 a53891a <=( (not A170)  and  a53890a );
 a53895a <=( (not A201)  and  (not A200) );
 a53896a <=( (not A166)  and  a53895a );
 a53897a <=( a53896a  and  a53891a );
 a53901a <=( (not A266)  and  (not A233) );
 a53902a <=( (not A232)  and  a53901a );
 a53905a <=( (not A269)  and  (not A268) );
 a53908a <=( (not A300)  and  A298 );
 a53909a <=( a53908a  and  a53905a );
 a53910a <=( a53909a  and  a53902a );
 a53914a <=( (not A167)  and  A169 );
 a53915a <=( (not A170)  and  a53914a );
 a53919a <=( (not A201)  and  (not A200) );
 a53920a <=( (not A166)  and  a53919a );
 a53921a <=( a53920a  and  a53915a );
 a53925a <=( (not A266)  and  (not A233) );
 a53926a <=( (not A232)  and  a53925a );
 a53929a <=( (not A269)  and  (not A268) );
 a53932a <=( A299  and  A298 );
 a53933a <=( a53932a  and  a53929a );
 a53934a <=( a53933a  and  a53926a );
 a53938a <=( (not A167)  and  A169 );
 a53939a <=( (not A170)  and  a53938a );
 a53943a <=( (not A201)  and  (not A200) );
 a53944a <=( (not A166)  and  a53943a );
 a53945a <=( a53944a  and  a53939a );
 a53949a <=( (not A266)  and  (not A233) );
 a53950a <=( (not A232)  and  a53949a );
 a53953a <=( (not A269)  and  (not A268) );
 a53956a <=( (not A299)  and  (not A298) );
 a53957a <=( a53956a  and  a53953a );
 a53958a <=( a53957a  and  a53950a );
 a53962a <=( (not A167)  and  A169 );
 a53963a <=( (not A170)  and  a53962a );
 a53967a <=( (not A201)  and  (not A200) );
 a53968a <=( (not A166)  and  a53967a );
 a53969a <=( a53968a  and  a53963a );
 a53973a <=( (not A266)  and  (not A233) );
 a53974a <=( (not A232)  and  a53973a );
 a53977a <=( A298  and  (not A267) );
 a53980a <=( (not A302)  and  (not A301) );
 a53981a <=( a53980a  and  a53977a );
 a53982a <=( a53981a  and  a53974a );
 a53986a <=( (not A167)  and  A169 );
 a53987a <=( (not A170)  and  a53986a );
 a53991a <=( (not A201)  and  (not A200) );
 a53992a <=( (not A166)  and  a53991a );
 a53993a <=( a53992a  and  a53987a );
 a53997a <=( (not A265)  and  (not A233) );
 a53998a <=( (not A232)  and  a53997a );
 a54001a <=( A298  and  (not A266) );
 a54004a <=( (not A302)  and  (not A301) );
 a54005a <=( a54004a  and  a54001a );
 a54006a <=( a54005a  and  a53998a );
 a54010a <=( (not A167)  and  A169 );
 a54011a <=( (not A170)  and  a54010a );
 a54015a <=( (not A200)  and  (not A199) );
 a54016a <=( (not A166)  and  a54015a );
 a54017a <=( a54016a  and  a54011a );
 a54021a <=( A265  and  A233 );
 a54022a <=( A232  and  a54021a );
 a54025a <=( (not A269)  and  (not A268) );
 a54028a <=( (not A300)  and  (not A299) );
 a54029a <=( a54028a  and  a54025a );
 a54030a <=( a54029a  and  a54022a );
 a54034a <=( (not A167)  and  A169 );
 a54035a <=( (not A170)  and  a54034a );
 a54039a <=( (not A200)  and  (not A199) );
 a54040a <=( (not A166)  and  a54039a );
 a54041a <=( a54040a  and  a54035a );
 a54045a <=( A265  and  A233 );
 a54046a <=( A232  and  a54045a );
 a54049a <=( (not A269)  and  (not A268) );
 a54052a <=( A299  and  A298 );
 a54053a <=( a54052a  and  a54049a );
 a54054a <=( a54053a  and  a54046a );
 a54058a <=( (not A167)  and  A169 );
 a54059a <=( (not A170)  and  a54058a );
 a54063a <=( (not A200)  and  (not A199) );
 a54064a <=( (not A166)  and  a54063a );
 a54065a <=( a54064a  and  a54059a );
 a54069a <=( A265  and  A233 );
 a54070a <=( A232  and  a54069a );
 a54073a <=( (not A269)  and  (not A268) );
 a54076a <=( (not A299)  and  (not A298) );
 a54077a <=( a54076a  and  a54073a );
 a54078a <=( a54077a  and  a54070a );
 a54082a <=( (not A167)  and  A169 );
 a54083a <=( (not A170)  and  a54082a );
 a54087a <=( (not A200)  and  (not A199) );
 a54088a <=( (not A166)  and  a54087a );
 a54089a <=( a54088a  and  a54083a );
 a54093a <=( A265  and  A233 );
 a54094a <=( A232  and  a54093a );
 a54097a <=( (not A299)  and  (not A267) );
 a54100a <=( (not A302)  and  (not A301) );
 a54101a <=( a54100a  and  a54097a );
 a54102a <=( a54101a  and  a54094a );
 a54106a <=( (not A167)  and  A169 );
 a54107a <=( (not A170)  and  a54106a );
 a54111a <=( (not A200)  and  (not A199) );
 a54112a <=( (not A166)  and  a54111a );
 a54113a <=( a54112a  and  a54107a );
 a54117a <=( A265  and  A233 );
 a54118a <=( A232  and  a54117a );
 a54121a <=( (not A299)  and  A266 );
 a54124a <=( (not A302)  and  (not A301) );
 a54125a <=( a54124a  and  a54121a );
 a54126a <=( a54125a  and  a54118a );
 a54130a <=( (not A167)  and  A169 );
 a54131a <=( (not A170)  and  a54130a );
 a54135a <=( (not A200)  and  (not A199) );
 a54136a <=( (not A166)  and  a54135a );
 a54137a <=( a54136a  and  a54131a );
 a54141a <=( (not A265)  and  A233 );
 a54142a <=( A232  and  a54141a );
 a54145a <=( (not A299)  and  (not A266) );
 a54148a <=( (not A302)  and  (not A301) );
 a54149a <=( a54148a  and  a54145a );
 a54150a <=( a54149a  and  a54142a );
 a54154a <=( (not A167)  and  A169 );
 a54155a <=( (not A170)  and  a54154a );
 a54159a <=( (not A200)  and  (not A199) );
 a54160a <=( (not A166)  and  a54159a );
 a54161a <=( a54160a  and  a54155a );
 a54165a <=( (not A236)  and  (not A235) );
 a54166a <=( (not A233)  and  a54165a );
 a54169a <=( A266  and  A265 );
 a54172a <=( (not A300)  and  A298 );
 a54173a <=( a54172a  and  a54169a );
 a54174a <=( a54173a  and  a54166a );
 a54178a <=( (not A167)  and  A169 );
 a54179a <=( (not A170)  and  a54178a );
 a54183a <=( (not A200)  and  (not A199) );
 a54184a <=( (not A166)  and  a54183a );
 a54185a <=( a54184a  and  a54179a );
 a54189a <=( (not A236)  and  (not A235) );
 a54190a <=( (not A233)  and  a54189a );
 a54193a <=( A266  and  A265 );
 a54196a <=( A299  and  A298 );
 a54197a <=( a54196a  and  a54193a );
 a54198a <=( a54197a  and  a54190a );
 a54202a <=( (not A167)  and  A169 );
 a54203a <=( (not A170)  and  a54202a );
 a54207a <=( (not A200)  and  (not A199) );
 a54208a <=( (not A166)  and  a54207a );
 a54209a <=( a54208a  and  a54203a );
 a54213a <=( (not A236)  and  (not A235) );
 a54214a <=( (not A233)  and  a54213a );
 a54217a <=( A266  and  A265 );
 a54220a <=( (not A299)  and  (not A298) );
 a54221a <=( a54220a  and  a54217a );
 a54222a <=( a54221a  and  a54214a );
 a54226a <=( (not A167)  and  A169 );
 a54227a <=( (not A170)  and  a54226a );
 a54231a <=( (not A200)  and  (not A199) );
 a54232a <=( (not A166)  and  a54231a );
 a54233a <=( a54232a  and  a54227a );
 a54237a <=( (not A236)  and  (not A235) );
 a54238a <=( (not A233)  and  a54237a );
 a54241a <=( (not A267)  and  (not A266) );
 a54244a <=( (not A300)  and  A298 );
 a54245a <=( a54244a  and  a54241a );
 a54246a <=( a54245a  and  a54238a );
 a54250a <=( (not A167)  and  A169 );
 a54251a <=( (not A170)  and  a54250a );
 a54255a <=( (not A200)  and  (not A199) );
 a54256a <=( (not A166)  and  a54255a );
 a54257a <=( a54256a  and  a54251a );
 a54261a <=( (not A236)  and  (not A235) );
 a54262a <=( (not A233)  and  a54261a );
 a54265a <=( (not A267)  and  (not A266) );
 a54268a <=( A299  and  A298 );
 a54269a <=( a54268a  and  a54265a );
 a54270a <=( a54269a  and  a54262a );
 a54274a <=( (not A167)  and  A169 );
 a54275a <=( (not A170)  and  a54274a );
 a54279a <=( (not A200)  and  (not A199) );
 a54280a <=( (not A166)  and  a54279a );
 a54281a <=( a54280a  and  a54275a );
 a54285a <=( (not A236)  and  (not A235) );
 a54286a <=( (not A233)  and  a54285a );
 a54289a <=( (not A267)  and  (not A266) );
 a54292a <=( (not A299)  and  (not A298) );
 a54293a <=( a54292a  and  a54289a );
 a54294a <=( a54293a  and  a54286a );
 a54298a <=( (not A167)  and  A169 );
 a54299a <=( (not A170)  and  a54298a );
 a54303a <=( (not A200)  and  (not A199) );
 a54304a <=( (not A166)  and  a54303a );
 a54305a <=( a54304a  and  a54299a );
 a54309a <=( (not A236)  and  (not A235) );
 a54310a <=( (not A233)  and  a54309a );
 a54313a <=( (not A266)  and  (not A265) );
 a54316a <=( (not A300)  and  A298 );
 a54317a <=( a54316a  and  a54313a );
 a54318a <=( a54317a  and  a54310a );
 a54322a <=( (not A167)  and  A169 );
 a54323a <=( (not A170)  and  a54322a );
 a54327a <=( (not A200)  and  (not A199) );
 a54328a <=( (not A166)  and  a54327a );
 a54329a <=( a54328a  and  a54323a );
 a54333a <=( (not A236)  and  (not A235) );
 a54334a <=( (not A233)  and  a54333a );
 a54337a <=( (not A266)  and  (not A265) );
 a54340a <=( A299  and  A298 );
 a54341a <=( a54340a  and  a54337a );
 a54342a <=( a54341a  and  a54334a );
 a54346a <=( (not A167)  and  A169 );
 a54347a <=( (not A170)  and  a54346a );
 a54351a <=( (not A200)  and  (not A199) );
 a54352a <=( (not A166)  and  a54351a );
 a54353a <=( a54352a  and  a54347a );
 a54357a <=( (not A236)  and  (not A235) );
 a54358a <=( (not A233)  and  a54357a );
 a54361a <=( (not A266)  and  (not A265) );
 a54364a <=( (not A299)  and  (not A298) );
 a54365a <=( a54364a  and  a54361a );
 a54366a <=( a54365a  and  a54358a );
 a54370a <=( (not A167)  and  A169 );
 a54371a <=( (not A170)  and  a54370a );
 a54375a <=( (not A200)  and  (not A199) );
 a54376a <=( (not A166)  and  a54375a );
 a54377a <=( a54376a  and  a54371a );
 a54381a <=( A265  and  (not A234) );
 a54382a <=( (not A233)  and  a54381a );
 a54385a <=( A298  and  A266 );
 a54388a <=( (not A302)  and  (not A301) );
 a54389a <=( a54388a  and  a54385a );
 a54390a <=( a54389a  and  a54382a );
 a54394a <=( (not A167)  and  A169 );
 a54395a <=( (not A170)  and  a54394a );
 a54399a <=( (not A200)  and  (not A199) );
 a54400a <=( (not A166)  and  a54399a );
 a54401a <=( a54400a  and  a54395a );
 a54405a <=( (not A266)  and  (not A234) );
 a54406a <=( (not A233)  and  a54405a );
 a54409a <=( (not A269)  and  (not A268) );
 a54412a <=( (not A300)  and  A298 );
 a54413a <=( a54412a  and  a54409a );
 a54414a <=( a54413a  and  a54406a );
 a54418a <=( (not A167)  and  A169 );
 a54419a <=( (not A170)  and  a54418a );
 a54423a <=( (not A200)  and  (not A199) );
 a54424a <=( (not A166)  and  a54423a );
 a54425a <=( a54424a  and  a54419a );
 a54429a <=( (not A266)  and  (not A234) );
 a54430a <=( (not A233)  and  a54429a );
 a54433a <=( (not A269)  and  (not A268) );
 a54436a <=( A299  and  A298 );
 a54437a <=( a54436a  and  a54433a );
 a54438a <=( a54437a  and  a54430a );
 a54442a <=( (not A167)  and  A169 );
 a54443a <=( (not A170)  and  a54442a );
 a54447a <=( (not A200)  and  (not A199) );
 a54448a <=( (not A166)  and  a54447a );
 a54449a <=( a54448a  and  a54443a );
 a54453a <=( (not A266)  and  (not A234) );
 a54454a <=( (not A233)  and  a54453a );
 a54457a <=( (not A269)  and  (not A268) );
 a54460a <=( (not A299)  and  (not A298) );
 a54461a <=( a54460a  and  a54457a );
 a54462a <=( a54461a  and  a54454a );
 a54466a <=( (not A167)  and  A169 );
 a54467a <=( (not A170)  and  a54466a );
 a54471a <=( (not A200)  and  (not A199) );
 a54472a <=( (not A166)  and  a54471a );
 a54473a <=( a54472a  and  a54467a );
 a54477a <=( (not A266)  and  (not A234) );
 a54478a <=( (not A233)  and  a54477a );
 a54481a <=( A298  and  (not A267) );
 a54484a <=( (not A302)  and  (not A301) );
 a54485a <=( a54484a  and  a54481a );
 a54486a <=( a54485a  and  a54478a );
 a54490a <=( (not A167)  and  A169 );
 a54491a <=( (not A170)  and  a54490a );
 a54495a <=( (not A200)  and  (not A199) );
 a54496a <=( (not A166)  and  a54495a );
 a54497a <=( a54496a  and  a54491a );
 a54501a <=( (not A265)  and  (not A234) );
 a54502a <=( (not A233)  and  a54501a );
 a54505a <=( A298  and  (not A266) );
 a54508a <=( (not A302)  and  (not A301) );
 a54509a <=( a54508a  and  a54505a );
 a54510a <=( a54509a  and  a54502a );
 a54514a <=( (not A167)  and  A169 );
 a54515a <=( (not A170)  and  a54514a );
 a54519a <=( (not A200)  and  (not A199) );
 a54520a <=( (not A166)  and  a54519a );
 a54521a <=( a54520a  and  a54515a );
 a54525a <=( A265  and  (not A233) );
 a54526a <=( (not A232)  and  a54525a );
 a54529a <=( A298  and  A266 );
 a54532a <=( (not A302)  and  (not A301) );
 a54533a <=( a54532a  and  a54529a );
 a54534a <=( a54533a  and  a54526a );
 a54538a <=( (not A167)  and  A169 );
 a54539a <=( (not A170)  and  a54538a );
 a54543a <=( (not A200)  and  (not A199) );
 a54544a <=( (not A166)  and  a54543a );
 a54545a <=( a54544a  and  a54539a );
 a54549a <=( (not A266)  and  (not A233) );
 a54550a <=( (not A232)  and  a54549a );
 a54553a <=( (not A269)  and  (not A268) );
 a54556a <=( (not A300)  and  A298 );
 a54557a <=( a54556a  and  a54553a );
 a54558a <=( a54557a  and  a54550a );
 a54562a <=( (not A167)  and  A169 );
 a54563a <=( (not A170)  and  a54562a );
 a54567a <=( (not A200)  and  (not A199) );
 a54568a <=( (not A166)  and  a54567a );
 a54569a <=( a54568a  and  a54563a );
 a54573a <=( (not A266)  and  (not A233) );
 a54574a <=( (not A232)  and  a54573a );
 a54577a <=( (not A269)  and  (not A268) );
 a54580a <=( A299  and  A298 );
 a54581a <=( a54580a  and  a54577a );
 a54582a <=( a54581a  and  a54574a );
 a54586a <=( (not A167)  and  A169 );
 a54587a <=( (not A170)  and  a54586a );
 a54591a <=( (not A200)  and  (not A199) );
 a54592a <=( (not A166)  and  a54591a );
 a54593a <=( a54592a  and  a54587a );
 a54597a <=( (not A266)  and  (not A233) );
 a54598a <=( (not A232)  and  a54597a );
 a54601a <=( (not A269)  and  (not A268) );
 a54604a <=( (not A299)  and  (not A298) );
 a54605a <=( a54604a  and  a54601a );
 a54606a <=( a54605a  and  a54598a );
 a54610a <=( (not A167)  and  A169 );
 a54611a <=( (not A170)  and  a54610a );
 a54615a <=( (not A200)  and  (not A199) );
 a54616a <=( (not A166)  and  a54615a );
 a54617a <=( a54616a  and  a54611a );
 a54621a <=( (not A266)  and  (not A233) );
 a54622a <=( (not A232)  and  a54621a );
 a54625a <=( A298  and  (not A267) );
 a54628a <=( (not A302)  and  (not A301) );
 a54629a <=( a54628a  and  a54625a );
 a54630a <=( a54629a  and  a54622a );
 a54634a <=( (not A167)  and  A169 );
 a54635a <=( (not A170)  and  a54634a );
 a54639a <=( (not A200)  and  (not A199) );
 a54640a <=( (not A166)  and  a54639a );
 a54641a <=( a54640a  and  a54635a );
 a54645a <=( (not A265)  and  (not A233) );
 a54646a <=( (not A232)  and  a54645a );
 a54649a <=( A298  and  (not A266) );
 a54652a <=( (not A302)  and  (not A301) );
 a54653a <=( a54652a  and  a54649a );
 a54654a <=( a54653a  and  a54646a );
 a54658a <=( (not A166)  and  (not A167) );
 a54659a <=( (not A169)  and  a54658a );
 a54663a <=( A232  and  A200 );
 a54664a <=( (not A199)  and  a54663a );
 a54665a <=( a54664a  and  a54659a );
 a54669a <=( (not A268)  and  A265 );
 a54670a <=( A233  and  a54669a );
 a54673a <=( (not A299)  and  (not A269) );
 a54676a <=( (not A302)  and  (not A301) );
 a54677a <=( a54676a  and  a54673a );
 a54678a <=( a54677a  and  a54670a );
 a54682a <=( (not A166)  and  (not A167) );
 a54683a <=( (not A169)  and  a54682a );
 a54687a <=( (not A233)  and  A200 );
 a54688a <=( (not A199)  and  a54687a );
 a54689a <=( a54688a  and  a54683a );
 a54693a <=( A265  and  (not A236) );
 a54694a <=( (not A235)  and  a54693a );
 a54697a <=( A298  and  A266 );
 a54700a <=( (not A302)  and  (not A301) );
 a54701a <=( a54700a  and  a54697a );
 a54702a <=( a54701a  and  a54694a );
 a54706a <=( (not A166)  and  (not A167) );
 a54707a <=( (not A169)  and  a54706a );
 a54711a <=( (not A233)  and  A200 );
 a54712a <=( (not A199)  and  a54711a );
 a54713a <=( a54712a  and  a54707a );
 a54717a <=( (not A266)  and  (not A236) );
 a54718a <=( (not A235)  and  a54717a );
 a54721a <=( (not A269)  and  (not A268) );
 a54724a <=( (not A300)  and  A298 );
 a54725a <=( a54724a  and  a54721a );
 a54726a <=( a54725a  and  a54718a );
 a54730a <=( (not A166)  and  (not A167) );
 a54731a <=( (not A169)  and  a54730a );
 a54735a <=( (not A233)  and  A200 );
 a54736a <=( (not A199)  and  a54735a );
 a54737a <=( a54736a  and  a54731a );
 a54741a <=( (not A266)  and  (not A236) );
 a54742a <=( (not A235)  and  a54741a );
 a54745a <=( (not A269)  and  (not A268) );
 a54748a <=( A299  and  A298 );
 a54749a <=( a54748a  and  a54745a );
 a54750a <=( a54749a  and  a54742a );
 a54754a <=( (not A166)  and  (not A167) );
 a54755a <=( (not A169)  and  a54754a );
 a54759a <=( (not A233)  and  A200 );
 a54760a <=( (not A199)  and  a54759a );
 a54761a <=( a54760a  and  a54755a );
 a54765a <=( (not A266)  and  (not A236) );
 a54766a <=( (not A235)  and  a54765a );
 a54769a <=( (not A269)  and  (not A268) );
 a54772a <=( (not A299)  and  (not A298) );
 a54773a <=( a54772a  and  a54769a );
 a54774a <=( a54773a  and  a54766a );
 a54778a <=( (not A166)  and  (not A167) );
 a54779a <=( (not A169)  and  a54778a );
 a54783a <=( (not A233)  and  A200 );
 a54784a <=( (not A199)  and  a54783a );
 a54785a <=( a54784a  and  a54779a );
 a54789a <=( (not A266)  and  (not A236) );
 a54790a <=( (not A235)  and  a54789a );
 a54793a <=( A298  and  (not A267) );
 a54796a <=( (not A302)  and  (not A301) );
 a54797a <=( a54796a  and  a54793a );
 a54798a <=( a54797a  and  a54790a );
 a54802a <=( (not A166)  and  (not A167) );
 a54803a <=( (not A169)  and  a54802a );
 a54807a <=( (not A233)  and  A200 );
 a54808a <=( (not A199)  and  a54807a );
 a54809a <=( a54808a  and  a54803a );
 a54813a <=( (not A265)  and  (not A236) );
 a54814a <=( (not A235)  and  a54813a );
 a54817a <=( A298  and  (not A266) );
 a54820a <=( (not A302)  and  (not A301) );
 a54821a <=( a54820a  and  a54817a );
 a54822a <=( a54821a  and  a54814a );
 a54826a <=( (not A166)  and  (not A167) );
 a54827a <=( (not A169)  and  a54826a );
 a54831a <=( (not A233)  and  A200 );
 a54832a <=( (not A199)  and  a54831a );
 a54833a <=( a54832a  and  a54827a );
 a54837a <=( (not A268)  and  (not A266) );
 a54838a <=( (not A234)  and  a54837a );
 a54841a <=( A298  and  (not A269) );
 a54844a <=( (not A302)  and  (not A301) );
 a54845a <=( a54844a  and  a54841a );
 a54846a <=( a54845a  and  a54838a );
 a54850a <=( (not A166)  and  (not A167) );
 a54851a <=( (not A169)  and  a54850a );
 a54855a <=( A232  and  A200 );
 a54856a <=( (not A199)  and  a54855a );
 a54857a <=( a54856a  and  a54851a );
 a54861a <=( A235  and  A234 );
 a54862a <=( (not A233)  and  a54861a );
 a54865a <=( (not A299)  and  A298 );
 a54868a <=( A301  and  A300 );
 a54869a <=( a54868a  and  a54865a );
 a54870a <=( a54869a  and  a54862a );
 a54874a <=( (not A166)  and  (not A167) );
 a54875a <=( (not A169)  and  a54874a );
 a54879a <=( A232  and  A200 );
 a54880a <=( (not A199)  and  a54879a );
 a54881a <=( a54880a  and  a54875a );
 a54885a <=( A235  and  A234 );
 a54886a <=( (not A233)  and  a54885a );
 a54889a <=( (not A299)  and  A298 );
 a54892a <=( A302  and  A300 );
 a54893a <=( a54892a  and  a54889a );
 a54894a <=( a54893a  and  a54886a );
 a54898a <=( (not A166)  and  (not A167) );
 a54899a <=( (not A169)  and  a54898a );
 a54903a <=( A232  and  A200 );
 a54904a <=( (not A199)  and  a54903a );
 a54905a <=( a54904a  and  a54899a );
 a54909a <=( A235  and  A234 );
 a54910a <=( (not A233)  and  a54909a );
 a54913a <=( (not A266)  and  A265 );
 a54916a <=( A268  and  A267 );
 a54917a <=( a54916a  and  a54913a );
 a54918a <=( a54917a  and  a54910a );
 a54922a <=( (not A166)  and  (not A167) );
 a54923a <=( (not A169)  and  a54922a );
 a54927a <=( A232  and  A200 );
 a54928a <=( (not A199)  and  a54927a );
 a54929a <=( a54928a  and  a54923a );
 a54933a <=( A235  and  A234 );
 a54934a <=( (not A233)  and  a54933a );
 a54937a <=( (not A266)  and  A265 );
 a54940a <=( A269  and  A267 );
 a54941a <=( a54940a  and  a54937a );
 a54942a <=( a54941a  and  a54934a );
 a54946a <=( (not A166)  and  (not A167) );
 a54947a <=( (not A169)  and  a54946a );
 a54951a <=( A232  and  A200 );
 a54952a <=( (not A199)  and  a54951a );
 a54953a <=( a54952a  and  a54947a );
 a54957a <=( A236  and  A234 );
 a54958a <=( (not A233)  and  a54957a );
 a54961a <=( (not A299)  and  A298 );
 a54964a <=( A301  and  A300 );
 a54965a <=( a54964a  and  a54961a );
 a54966a <=( a54965a  and  a54958a );
 a54970a <=( (not A166)  and  (not A167) );
 a54971a <=( (not A169)  and  a54970a );
 a54975a <=( A232  and  A200 );
 a54976a <=( (not A199)  and  a54975a );
 a54977a <=( a54976a  and  a54971a );
 a54981a <=( A236  and  A234 );
 a54982a <=( (not A233)  and  a54981a );
 a54985a <=( (not A299)  and  A298 );
 a54988a <=( A302  and  A300 );
 a54989a <=( a54988a  and  a54985a );
 a54990a <=( a54989a  and  a54982a );
 a54994a <=( (not A166)  and  (not A167) );
 a54995a <=( (not A169)  and  a54994a );
 a54999a <=( A232  and  A200 );
 a55000a <=( (not A199)  and  a54999a );
 a55001a <=( a55000a  and  a54995a );
 a55005a <=( A236  and  A234 );
 a55006a <=( (not A233)  and  a55005a );
 a55009a <=( (not A266)  and  A265 );
 a55012a <=( A268  and  A267 );
 a55013a <=( a55012a  and  a55009a );
 a55014a <=( a55013a  and  a55006a );
 a55018a <=( (not A166)  and  (not A167) );
 a55019a <=( (not A169)  and  a55018a );
 a55023a <=( A232  and  A200 );
 a55024a <=( (not A199)  and  a55023a );
 a55025a <=( a55024a  and  a55019a );
 a55029a <=( A236  and  A234 );
 a55030a <=( (not A233)  and  a55029a );
 a55033a <=( (not A266)  and  A265 );
 a55036a <=( A269  and  A267 );
 a55037a <=( a55036a  and  a55033a );
 a55038a <=( a55037a  and  a55030a );
 a55042a <=( (not A166)  and  (not A167) );
 a55043a <=( (not A169)  and  a55042a );
 a55047a <=( (not A232)  and  A200 );
 a55048a <=( (not A199)  and  a55047a );
 a55049a <=( a55048a  and  a55043a );
 a55053a <=( (not A268)  and  (not A266) );
 a55054a <=( (not A233)  and  a55053a );
 a55057a <=( A298  and  (not A269) );
 a55060a <=( (not A302)  and  (not A301) );
 a55061a <=( a55060a  and  a55057a );
 a55062a <=( a55061a  and  a55054a );
 a55066a <=( (not A166)  and  (not A167) );
 a55067a <=( (not A169)  and  a55066a );
 a55071a <=( A201  and  (not A200) );
 a55072a <=( A199  and  a55071a );
 a55073a <=( a55072a  and  a55067a );
 a55077a <=( A233  and  A232 );
 a55078a <=( A202  and  a55077a );
 a55081a <=( (not A267)  and  A265 );
 a55084a <=( (not A300)  and  (not A299) );
 a55085a <=( a55084a  and  a55081a );
 a55086a <=( a55085a  and  a55078a );
 a55090a <=( (not A166)  and  (not A167) );
 a55091a <=( (not A169)  and  a55090a );
 a55095a <=( A201  and  (not A200) );
 a55096a <=( A199  and  a55095a );
 a55097a <=( a55096a  and  a55091a );
 a55101a <=( A233  and  A232 );
 a55102a <=( A202  and  a55101a );
 a55105a <=( (not A267)  and  A265 );
 a55108a <=( A299  and  A298 );
 a55109a <=( a55108a  and  a55105a );
 a55110a <=( a55109a  and  a55102a );
 a55114a <=( (not A166)  and  (not A167) );
 a55115a <=( (not A169)  and  a55114a );
 a55119a <=( A201  and  (not A200) );
 a55120a <=( A199  and  a55119a );
 a55121a <=( a55120a  and  a55115a );
 a55125a <=( A233  and  A232 );
 a55126a <=( A202  and  a55125a );
 a55129a <=( (not A267)  and  A265 );
 a55132a <=( (not A299)  and  (not A298) );
 a55133a <=( a55132a  and  a55129a );
 a55134a <=( a55133a  and  a55126a );
 a55138a <=( (not A166)  and  (not A167) );
 a55139a <=( (not A169)  and  a55138a );
 a55143a <=( A201  and  (not A200) );
 a55144a <=( A199  and  a55143a );
 a55145a <=( a55144a  and  a55139a );
 a55149a <=( A233  and  A232 );
 a55150a <=( A202  and  a55149a );
 a55153a <=( A266  and  A265 );
 a55156a <=( (not A300)  and  (not A299) );
 a55157a <=( a55156a  and  a55153a );
 a55158a <=( a55157a  and  a55150a );
 a55162a <=( (not A166)  and  (not A167) );
 a55163a <=( (not A169)  and  a55162a );
 a55167a <=( A201  and  (not A200) );
 a55168a <=( A199  and  a55167a );
 a55169a <=( a55168a  and  a55163a );
 a55173a <=( A233  and  A232 );
 a55174a <=( A202  and  a55173a );
 a55177a <=( A266  and  A265 );
 a55180a <=( A299  and  A298 );
 a55181a <=( a55180a  and  a55177a );
 a55182a <=( a55181a  and  a55174a );
 a55186a <=( (not A166)  and  (not A167) );
 a55187a <=( (not A169)  and  a55186a );
 a55191a <=( A201  and  (not A200) );
 a55192a <=( A199  and  a55191a );
 a55193a <=( a55192a  and  a55187a );
 a55197a <=( A233  and  A232 );
 a55198a <=( A202  and  a55197a );
 a55201a <=( A266  and  A265 );
 a55204a <=( (not A299)  and  (not A298) );
 a55205a <=( a55204a  and  a55201a );
 a55206a <=( a55205a  and  a55198a );
 a55210a <=( (not A166)  and  (not A167) );
 a55211a <=( (not A169)  and  a55210a );
 a55215a <=( A201  and  (not A200) );
 a55216a <=( A199  and  a55215a );
 a55217a <=( a55216a  and  a55211a );
 a55221a <=( A233  and  A232 );
 a55222a <=( A202  and  a55221a );
 a55225a <=( (not A266)  and  (not A265) );
 a55228a <=( (not A300)  and  (not A299) );
 a55229a <=( a55228a  and  a55225a );
 a55230a <=( a55229a  and  a55222a );
 a55234a <=( (not A166)  and  (not A167) );
 a55235a <=( (not A169)  and  a55234a );
 a55239a <=( A201  and  (not A200) );
 a55240a <=( A199  and  a55239a );
 a55241a <=( a55240a  and  a55235a );
 a55245a <=( A233  and  A232 );
 a55246a <=( A202  and  a55245a );
 a55249a <=( (not A266)  and  (not A265) );
 a55252a <=( A299  and  A298 );
 a55253a <=( a55252a  and  a55249a );
 a55254a <=( a55253a  and  a55246a );
 a55258a <=( (not A166)  and  (not A167) );
 a55259a <=( (not A169)  and  a55258a );
 a55263a <=( A201  and  (not A200) );
 a55264a <=( A199  and  a55263a );
 a55265a <=( a55264a  and  a55259a );
 a55269a <=( A233  and  A232 );
 a55270a <=( A202  and  a55269a );
 a55273a <=( (not A266)  and  (not A265) );
 a55276a <=( (not A299)  and  (not A298) );
 a55277a <=( a55276a  and  a55273a );
 a55278a <=( a55277a  and  a55270a );
 a55282a <=( (not A166)  and  (not A167) );
 a55283a <=( (not A169)  and  a55282a );
 a55287a <=( A201  and  (not A200) );
 a55288a <=( A199  and  a55287a );
 a55289a <=( a55288a  and  a55283a );
 a55293a <=( A233  and  (not A232) );
 a55294a <=( A202  and  a55293a );
 a55297a <=( (not A299)  and  A298 );
 a55300a <=( A301  and  A300 );
 a55301a <=( a55300a  and  a55297a );
 a55302a <=( a55301a  and  a55294a );
 a55306a <=( (not A166)  and  (not A167) );
 a55307a <=( (not A169)  and  a55306a );
 a55311a <=( A201  and  (not A200) );
 a55312a <=( A199  and  a55311a );
 a55313a <=( a55312a  and  a55307a );
 a55317a <=( A233  and  (not A232) );
 a55318a <=( A202  and  a55317a );
 a55321a <=( (not A299)  and  A298 );
 a55324a <=( A302  and  A300 );
 a55325a <=( a55324a  and  a55321a );
 a55326a <=( a55325a  and  a55318a );
 a55330a <=( (not A166)  and  (not A167) );
 a55331a <=( (not A169)  and  a55330a );
 a55335a <=( A201  and  (not A200) );
 a55336a <=( A199  and  a55335a );
 a55337a <=( a55336a  and  a55331a );
 a55341a <=( A233  and  (not A232) );
 a55342a <=( A202  and  a55341a );
 a55345a <=( (not A266)  and  A265 );
 a55348a <=( A268  and  A267 );
 a55349a <=( a55348a  and  a55345a );
 a55350a <=( a55349a  and  a55342a );
 a55354a <=( (not A166)  and  (not A167) );
 a55355a <=( (not A169)  and  a55354a );
 a55359a <=( A201  and  (not A200) );
 a55360a <=( A199  and  a55359a );
 a55361a <=( a55360a  and  a55355a );
 a55365a <=( A233  and  (not A232) );
 a55366a <=( A202  and  a55365a );
 a55369a <=( (not A266)  and  A265 );
 a55372a <=( A269  and  A267 );
 a55373a <=( a55372a  and  a55369a );
 a55374a <=( a55373a  and  a55366a );
 a55378a <=( (not A166)  and  (not A167) );
 a55379a <=( (not A169)  and  a55378a );
 a55383a <=( A201  and  (not A200) );
 a55384a <=( A199  and  a55383a );
 a55385a <=( a55384a  and  a55379a );
 a55389a <=( (not A234)  and  (not A233) );
 a55390a <=( A202  and  a55389a );
 a55393a <=( A266  and  A265 );
 a55396a <=( (not A300)  and  A298 );
 a55397a <=( a55396a  and  a55393a );
 a55398a <=( a55397a  and  a55390a );
 a55402a <=( (not A166)  and  (not A167) );
 a55403a <=( (not A169)  and  a55402a );
 a55407a <=( A201  and  (not A200) );
 a55408a <=( A199  and  a55407a );
 a55409a <=( a55408a  and  a55403a );
 a55413a <=( (not A234)  and  (not A233) );
 a55414a <=( A202  and  a55413a );
 a55417a <=( A266  and  A265 );
 a55420a <=( A299  and  A298 );
 a55421a <=( a55420a  and  a55417a );
 a55422a <=( a55421a  and  a55414a );
 a55426a <=( (not A166)  and  (not A167) );
 a55427a <=( (not A169)  and  a55426a );
 a55431a <=( A201  and  (not A200) );
 a55432a <=( A199  and  a55431a );
 a55433a <=( a55432a  and  a55427a );
 a55437a <=( (not A234)  and  (not A233) );
 a55438a <=( A202  and  a55437a );
 a55441a <=( A266  and  A265 );
 a55444a <=( (not A299)  and  (not A298) );
 a55445a <=( a55444a  and  a55441a );
 a55446a <=( a55445a  and  a55438a );
 a55450a <=( (not A166)  and  (not A167) );
 a55451a <=( (not A169)  and  a55450a );
 a55455a <=( A201  and  (not A200) );
 a55456a <=( A199  and  a55455a );
 a55457a <=( a55456a  and  a55451a );
 a55461a <=( (not A234)  and  (not A233) );
 a55462a <=( A202  and  a55461a );
 a55465a <=( (not A267)  and  (not A266) );
 a55468a <=( (not A300)  and  A298 );
 a55469a <=( a55468a  and  a55465a );
 a55470a <=( a55469a  and  a55462a );
 a55474a <=( (not A166)  and  (not A167) );
 a55475a <=( (not A169)  and  a55474a );
 a55479a <=( A201  and  (not A200) );
 a55480a <=( A199  and  a55479a );
 a55481a <=( a55480a  and  a55475a );
 a55485a <=( (not A234)  and  (not A233) );
 a55486a <=( A202  and  a55485a );
 a55489a <=( (not A267)  and  (not A266) );
 a55492a <=( A299  and  A298 );
 a55493a <=( a55492a  and  a55489a );
 a55494a <=( a55493a  and  a55486a );
 a55498a <=( (not A166)  and  (not A167) );
 a55499a <=( (not A169)  and  a55498a );
 a55503a <=( A201  and  (not A200) );
 a55504a <=( A199  and  a55503a );
 a55505a <=( a55504a  and  a55499a );
 a55509a <=( (not A234)  and  (not A233) );
 a55510a <=( A202  and  a55509a );
 a55513a <=( (not A267)  and  (not A266) );
 a55516a <=( (not A299)  and  (not A298) );
 a55517a <=( a55516a  and  a55513a );
 a55518a <=( a55517a  and  a55510a );
 a55522a <=( (not A166)  and  (not A167) );
 a55523a <=( (not A169)  and  a55522a );
 a55527a <=( A201  and  (not A200) );
 a55528a <=( A199  and  a55527a );
 a55529a <=( a55528a  and  a55523a );
 a55533a <=( (not A234)  and  (not A233) );
 a55534a <=( A202  and  a55533a );
 a55537a <=( (not A266)  and  (not A265) );
 a55540a <=( (not A300)  and  A298 );
 a55541a <=( a55540a  and  a55537a );
 a55542a <=( a55541a  and  a55534a );
 a55546a <=( (not A166)  and  (not A167) );
 a55547a <=( (not A169)  and  a55546a );
 a55551a <=( A201  and  (not A200) );
 a55552a <=( A199  and  a55551a );
 a55553a <=( a55552a  and  a55547a );
 a55557a <=( (not A234)  and  (not A233) );
 a55558a <=( A202  and  a55557a );
 a55561a <=( (not A266)  and  (not A265) );
 a55564a <=( A299  and  A298 );
 a55565a <=( a55564a  and  a55561a );
 a55566a <=( a55565a  and  a55558a );
 a55570a <=( (not A166)  and  (not A167) );
 a55571a <=( (not A169)  and  a55570a );
 a55575a <=( A201  and  (not A200) );
 a55576a <=( A199  and  a55575a );
 a55577a <=( a55576a  and  a55571a );
 a55581a <=( (not A234)  and  (not A233) );
 a55582a <=( A202  and  a55581a );
 a55585a <=( (not A266)  and  (not A265) );
 a55588a <=( (not A299)  and  (not A298) );
 a55589a <=( a55588a  and  a55585a );
 a55590a <=( a55589a  and  a55582a );
 a55594a <=( (not A166)  and  (not A167) );
 a55595a <=( (not A169)  and  a55594a );
 a55599a <=( A201  and  (not A200) );
 a55600a <=( A199  and  a55599a );
 a55601a <=( a55600a  and  a55595a );
 a55605a <=( (not A233)  and  A232 );
 a55606a <=( A202  and  a55605a );
 a55609a <=( A235  and  A234 );
 a55612a <=( A299  and  (not A298) );
 a55613a <=( a55612a  and  a55609a );
 a55614a <=( a55613a  and  a55606a );
 a55618a <=( (not A166)  and  (not A167) );
 a55619a <=( (not A169)  and  a55618a );
 a55623a <=( A201  and  (not A200) );
 a55624a <=( A199  and  a55623a );
 a55625a <=( a55624a  and  a55619a );
 a55629a <=( (not A233)  and  A232 );
 a55630a <=( A202  and  a55629a );
 a55633a <=( A235  and  A234 );
 a55636a <=( A266  and  (not A265) );
 a55637a <=( a55636a  and  a55633a );
 a55638a <=( a55637a  and  a55630a );
 a55642a <=( (not A166)  and  (not A167) );
 a55643a <=( (not A169)  and  a55642a );
 a55647a <=( A201  and  (not A200) );
 a55648a <=( A199  and  a55647a );
 a55649a <=( a55648a  and  a55643a );
 a55653a <=( (not A233)  and  A232 );
 a55654a <=( A202  and  a55653a );
 a55657a <=( A236  and  A234 );
 a55660a <=( A299  and  (not A298) );
 a55661a <=( a55660a  and  a55657a );
 a55662a <=( a55661a  and  a55654a );
 a55666a <=( (not A166)  and  (not A167) );
 a55667a <=( (not A169)  and  a55666a );
 a55671a <=( A201  and  (not A200) );
 a55672a <=( A199  and  a55671a );
 a55673a <=( a55672a  and  a55667a );
 a55677a <=( (not A233)  and  A232 );
 a55678a <=( A202  and  a55677a );
 a55681a <=( A236  and  A234 );
 a55684a <=( A266  and  (not A265) );
 a55685a <=( a55684a  and  a55681a );
 a55686a <=( a55685a  and  a55678a );
 a55690a <=( (not A166)  and  (not A167) );
 a55691a <=( (not A169)  and  a55690a );
 a55695a <=( A201  and  (not A200) );
 a55696a <=( A199  and  a55695a );
 a55697a <=( a55696a  and  a55691a );
 a55701a <=( (not A233)  and  (not A232) );
 a55702a <=( A202  and  a55701a );
 a55705a <=( A266  and  A265 );
 a55708a <=( (not A300)  and  A298 );
 a55709a <=( a55708a  and  a55705a );
 a55710a <=( a55709a  and  a55702a );
 a55714a <=( (not A166)  and  (not A167) );
 a55715a <=( (not A169)  and  a55714a );
 a55719a <=( A201  and  (not A200) );
 a55720a <=( A199  and  a55719a );
 a55721a <=( a55720a  and  a55715a );
 a55725a <=( (not A233)  and  (not A232) );
 a55726a <=( A202  and  a55725a );
 a55729a <=( A266  and  A265 );
 a55732a <=( A299  and  A298 );
 a55733a <=( a55732a  and  a55729a );
 a55734a <=( a55733a  and  a55726a );
 a55738a <=( (not A166)  and  (not A167) );
 a55739a <=( (not A169)  and  a55738a );
 a55743a <=( A201  and  (not A200) );
 a55744a <=( A199  and  a55743a );
 a55745a <=( a55744a  and  a55739a );
 a55749a <=( (not A233)  and  (not A232) );
 a55750a <=( A202  and  a55749a );
 a55753a <=( A266  and  A265 );
 a55756a <=( (not A299)  and  (not A298) );
 a55757a <=( a55756a  and  a55753a );
 a55758a <=( a55757a  and  a55750a );
 a55762a <=( (not A166)  and  (not A167) );
 a55763a <=( (not A169)  and  a55762a );
 a55767a <=( A201  and  (not A200) );
 a55768a <=( A199  and  a55767a );
 a55769a <=( a55768a  and  a55763a );
 a55773a <=( (not A233)  and  (not A232) );
 a55774a <=( A202  and  a55773a );
 a55777a <=( (not A267)  and  (not A266) );
 a55780a <=( (not A300)  and  A298 );
 a55781a <=( a55780a  and  a55777a );
 a55782a <=( a55781a  and  a55774a );
 a55786a <=( (not A166)  and  (not A167) );
 a55787a <=( (not A169)  and  a55786a );
 a55791a <=( A201  and  (not A200) );
 a55792a <=( A199  and  a55791a );
 a55793a <=( a55792a  and  a55787a );
 a55797a <=( (not A233)  and  (not A232) );
 a55798a <=( A202  and  a55797a );
 a55801a <=( (not A267)  and  (not A266) );
 a55804a <=( A299  and  A298 );
 a55805a <=( a55804a  and  a55801a );
 a55806a <=( a55805a  and  a55798a );
 a55810a <=( (not A166)  and  (not A167) );
 a55811a <=( (not A169)  and  a55810a );
 a55815a <=( A201  and  (not A200) );
 a55816a <=( A199  and  a55815a );
 a55817a <=( a55816a  and  a55811a );
 a55821a <=( (not A233)  and  (not A232) );
 a55822a <=( A202  and  a55821a );
 a55825a <=( (not A267)  and  (not A266) );
 a55828a <=( (not A299)  and  (not A298) );
 a55829a <=( a55828a  and  a55825a );
 a55830a <=( a55829a  and  a55822a );
 a55834a <=( (not A166)  and  (not A167) );
 a55835a <=( (not A169)  and  a55834a );
 a55839a <=( A201  and  (not A200) );
 a55840a <=( A199  and  a55839a );
 a55841a <=( a55840a  and  a55835a );
 a55845a <=( (not A233)  and  (not A232) );
 a55846a <=( A202  and  a55845a );
 a55849a <=( (not A266)  and  (not A265) );
 a55852a <=( (not A300)  and  A298 );
 a55853a <=( a55852a  and  a55849a );
 a55854a <=( a55853a  and  a55846a );
 a55858a <=( (not A166)  and  (not A167) );
 a55859a <=( (not A169)  and  a55858a );
 a55863a <=( A201  and  (not A200) );
 a55864a <=( A199  and  a55863a );
 a55865a <=( a55864a  and  a55859a );
 a55869a <=( (not A233)  and  (not A232) );
 a55870a <=( A202  and  a55869a );
 a55873a <=( (not A266)  and  (not A265) );
 a55876a <=( A299  and  A298 );
 a55877a <=( a55876a  and  a55873a );
 a55878a <=( a55877a  and  a55870a );
 a55882a <=( (not A166)  and  (not A167) );
 a55883a <=( (not A169)  and  a55882a );
 a55887a <=( A201  and  (not A200) );
 a55888a <=( A199  and  a55887a );
 a55889a <=( a55888a  and  a55883a );
 a55893a <=( (not A233)  and  (not A232) );
 a55894a <=( A202  and  a55893a );
 a55897a <=( (not A266)  and  (not A265) );
 a55900a <=( (not A299)  and  (not A298) );
 a55901a <=( a55900a  and  a55897a );
 a55902a <=( a55901a  and  a55894a );
 a55906a <=( (not A166)  and  (not A167) );
 a55907a <=( (not A169)  and  a55906a );
 a55911a <=( A201  and  (not A200) );
 a55912a <=( A199  and  a55911a );
 a55913a <=( a55912a  and  a55907a );
 a55917a <=( A233  and  A232 );
 a55918a <=( A203  and  a55917a );
 a55921a <=( (not A267)  and  A265 );
 a55924a <=( (not A300)  and  (not A299) );
 a55925a <=( a55924a  and  a55921a );
 a55926a <=( a55925a  and  a55918a );
 a55930a <=( (not A166)  and  (not A167) );
 a55931a <=( (not A169)  and  a55930a );
 a55935a <=( A201  and  (not A200) );
 a55936a <=( A199  and  a55935a );
 a55937a <=( a55936a  and  a55931a );
 a55941a <=( A233  and  A232 );
 a55942a <=( A203  and  a55941a );
 a55945a <=( (not A267)  and  A265 );
 a55948a <=( A299  and  A298 );
 a55949a <=( a55948a  and  a55945a );
 a55950a <=( a55949a  and  a55942a );
 a55954a <=( (not A166)  and  (not A167) );
 a55955a <=( (not A169)  and  a55954a );
 a55959a <=( A201  and  (not A200) );
 a55960a <=( A199  and  a55959a );
 a55961a <=( a55960a  and  a55955a );
 a55965a <=( A233  and  A232 );
 a55966a <=( A203  and  a55965a );
 a55969a <=( (not A267)  and  A265 );
 a55972a <=( (not A299)  and  (not A298) );
 a55973a <=( a55972a  and  a55969a );
 a55974a <=( a55973a  and  a55966a );
 a55978a <=( (not A166)  and  (not A167) );
 a55979a <=( (not A169)  and  a55978a );
 a55983a <=( A201  and  (not A200) );
 a55984a <=( A199  and  a55983a );
 a55985a <=( a55984a  and  a55979a );
 a55989a <=( A233  and  A232 );
 a55990a <=( A203  and  a55989a );
 a55993a <=( A266  and  A265 );
 a55996a <=( (not A300)  and  (not A299) );
 a55997a <=( a55996a  and  a55993a );
 a55998a <=( a55997a  and  a55990a );
 a56002a <=( (not A166)  and  (not A167) );
 a56003a <=( (not A169)  and  a56002a );
 a56007a <=( A201  and  (not A200) );
 a56008a <=( A199  and  a56007a );
 a56009a <=( a56008a  and  a56003a );
 a56013a <=( A233  and  A232 );
 a56014a <=( A203  and  a56013a );
 a56017a <=( A266  and  A265 );
 a56020a <=( A299  and  A298 );
 a56021a <=( a56020a  and  a56017a );
 a56022a <=( a56021a  and  a56014a );
 a56026a <=( (not A166)  and  (not A167) );
 a56027a <=( (not A169)  and  a56026a );
 a56031a <=( A201  and  (not A200) );
 a56032a <=( A199  and  a56031a );
 a56033a <=( a56032a  and  a56027a );
 a56037a <=( A233  and  A232 );
 a56038a <=( A203  and  a56037a );
 a56041a <=( A266  and  A265 );
 a56044a <=( (not A299)  and  (not A298) );
 a56045a <=( a56044a  and  a56041a );
 a56046a <=( a56045a  and  a56038a );
 a56050a <=( (not A166)  and  (not A167) );
 a56051a <=( (not A169)  and  a56050a );
 a56055a <=( A201  and  (not A200) );
 a56056a <=( A199  and  a56055a );
 a56057a <=( a56056a  and  a56051a );
 a56061a <=( A233  and  A232 );
 a56062a <=( A203  and  a56061a );
 a56065a <=( (not A266)  and  (not A265) );
 a56068a <=( (not A300)  and  (not A299) );
 a56069a <=( a56068a  and  a56065a );
 a56070a <=( a56069a  and  a56062a );
 a56074a <=( (not A166)  and  (not A167) );
 a56075a <=( (not A169)  and  a56074a );
 a56079a <=( A201  and  (not A200) );
 a56080a <=( A199  and  a56079a );
 a56081a <=( a56080a  and  a56075a );
 a56085a <=( A233  and  A232 );
 a56086a <=( A203  and  a56085a );
 a56089a <=( (not A266)  and  (not A265) );
 a56092a <=( A299  and  A298 );
 a56093a <=( a56092a  and  a56089a );
 a56094a <=( a56093a  and  a56086a );
 a56098a <=( (not A166)  and  (not A167) );
 a56099a <=( (not A169)  and  a56098a );
 a56103a <=( A201  and  (not A200) );
 a56104a <=( A199  and  a56103a );
 a56105a <=( a56104a  and  a56099a );
 a56109a <=( A233  and  A232 );
 a56110a <=( A203  and  a56109a );
 a56113a <=( (not A266)  and  (not A265) );
 a56116a <=( (not A299)  and  (not A298) );
 a56117a <=( a56116a  and  a56113a );
 a56118a <=( a56117a  and  a56110a );
 a56122a <=( (not A166)  and  (not A167) );
 a56123a <=( (not A169)  and  a56122a );
 a56127a <=( A201  and  (not A200) );
 a56128a <=( A199  and  a56127a );
 a56129a <=( a56128a  and  a56123a );
 a56133a <=( A233  and  (not A232) );
 a56134a <=( A203  and  a56133a );
 a56137a <=( (not A299)  and  A298 );
 a56140a <=( A301  and  A300 );
 a56141a <=( a56140a  and  a56137a );
 a56142a <=( a56141a  and  a56134a );
 a56146a <=( (not A166)  and  (not A167) );
 a56147a <=( (not A169)  and  a56146a );
 a56151a <=( A201  and  (not A200) );
 a56152a <=( A199  and  a56151a );
 a56153a <=( a56152a  and  a56147a );
 a56157a <=( A233  and  (not A232) );
 a56158a <=( A203  and  a56157a );
 a56161a <=( (not A299)  and  A298 );
 a56164a <=( A302  and  A300 );
 a56165a <=( a56164a  and  a56161a );
 a56166a <=( a56165a  and  a56158a );
 a56170a <=( (not A166)  and  (not A167) );
 a56171a <=( (not A169)  and  a56170a );
 a56175a <=( A201  and  (not A200) );
 a56176a <=( A199  and  a56175a );
 a56177a <=( a56176a  and  a56171a );
 a56181a <=( A233  and  (not A232) );
 a56182a <=( A203  and  a56181a );
 a56185a <=( (not A266)  and  A265 );
 a56188a <=( A268  and  A267 );
 a56189a <=( a56188a  and  a56185a );
 a56190a <=( a56189a  and  a56182a );
 a56194a <=( (not A166)  and  (not A167) );
 a56195a <=( (not A169)  and  a56194a );
 a56199a <=( A201  and  (not A200) );
 a56200a <=( A199  and  a56199a );
 a56201a <=( a56200a  and  a56195a );
 a56205a <=( A233  and  (not A232) );
 a56206a <=( A203  and  a56205a );
 a56209a <=( (not A266)  and  A265 );
 a56212a <=( A269  and  A267 );
 a56213a <=( a56212a  and  a56209a );
 a56214a <=( a56213a  and  a56206a );
 a56218a <=( (not A166)  and  (not A167) );
 a56219a <=( (not A169)  and  a56218a );
 a56223a <=( A201  and  (not A200) );
 a56224a <=( A199  and  a56223a );
 a56225a <=( a56224a  and  a56219a );
 a56229a <=( (not A234)  and  (not A233) );
 a56230a <=( A203  and  a56229a );
 a56233a <=( A266  and  A265 );
 a56236a <=( (not A300)  and  A298 );
 a56237a <=( a56236a  and  a56233a );
 a56238a <=( a56237a  and  a56230a );
 a56242a <=( (not A166)  and  (not A167) );
 a56243a <=( (not A169)  and  a56242a );
 a56247a <=( A201  and  (not A200) );
 a56248a <=( A199  and  a56247a );
 a56249a <=( a56248a  and  a56243a );
 a56253a <=( (not A234)  and  (not A233) );
 a56254a <=( A203  and  a56253a );
 a56257a <=( A266  and  A265 );
 a56260a <=( A299  and  A298 );
 a56261a <=( a56260a  and  a56257a );
 a56262a <=( a56261a  and  a56254a );
 a56266a <=( (not A166)  and  (not A167) );
 a56267a <=( (not A169)  and  a56266a );
 a56271a <=( A201  and  (not A200) );
 a56272a <=( A199  and  a56271a );
 a56273a <=( a56272a  and  a56267a );
 a56277a <=( (not A234)  and  (not A233) );
 a56278a <=( A203  and  a56277a );
 a56281a <=( A266  and  A265 );
 a56284a <=( (not A299)  and  (not A298) );
 a56285a <=( a56284a  and  a56281a );
 a56286a <=( a56285a  and  a56278a );
 a56290a <=( (not A166)  and  (not A167) );
 a56291a <=( (not A169)  and  a56290a );
 a56295a <=( A201  and  (not A200) );
 a56296a <=( A199  and  a56295a );
 a56297a <=( a56296a  and  a56291a );
 a56301a <=( (not A234)  and  (not A233) );
 a56302a <=( A203  and  a56301a );
 a56305a <=( (not A267)  and  (not A266) );
 a56308a <=( (not A300)  and  A298 );
 a56309a <=( a56308a  and  a56305a );
 a56310a <=( a56309a  and  a56302a );
 a56314a <=( (not A166)  and  (not A167) );
 a56315a <=( (not A169)  and  a56314a );
 a56319a <=( A201  and  (not A200) );
 a56320a <=( A199  and  a56319a );
 a56321a <=( a56320a  and  a56315a );
 a56325a <=( (not A234)  and  (not A233) );
 a56326a <=( A203  and  a56325a );
 a56329a <=( (not A267)  and  (not A266) );
 a56332a <=( A299  and  A298 );
 a56333a <=( a56332a  and  a56329a );
 a56334a <=( a56333a  and  a56326a );
 a56338a <=( (not A166)  and  (not A167) );
 a56339a <=( (not A169)  and  a56338a );
 a56343a <=( A201  and  (not A200) );
 a56344a <=( A199  and  a56343a );
 a56345a <=( a56344a  and  a56339a );
 a56349a <=( (not A234)  and  (not A233) );
 a56350a <=( A203  and  a56349a );
 a56353a <=( (not A267)  and  (not A266) );
 a56356a <=( (not A299)  and  (not A298) );
 a56357a <=( a56356a  and  a56353a );
 a56358a <=( a56357a  and  a56350a );
 a56362a <=( (not A166)  and  (not A167) );
 a56363a <=( (not A169)  and  a56362a );
 a56367a <=( A201  and  (not A200) );
 a56368a <=( A199  and  a56367a );
 a56369a <=( a56368a  and  a56363a );
 a56373a <=( (not A234)  and  (not A233) );
 a56374a <=( A203  and  a56373a );
 a56377a <=( (not A266)  and  (not A265) );
 a56380a <=( (not A300)  and  A298 );
 a56381a <=( a56380a  and  a56377a );
 a56382a <=( a56381a  and  a56374a );
 a56386a <=( (not A166)  and  (not A167) );
 a56387a <=( (not A169)  and  a56386a );
 a56391a <=( A201  and  (not A200) );
 a56392a <=( A199  and  a56391a );
 a56393a <=( a56392a  and  a56387a );
 a56397a <=( (not A234)  and  (not A233) );
 a56398a <=( A203  and  a56397a );
 a56401a <=( (not A266)  and  (not A265) );
 a56404a <=( A299  and  A298 );
 a56405a <=( a56404a  and  a56401a );
 a56406a <=( a56405a  and  a56398a );
 a56410a <=( (not A166)  and  (not A167) );
 a56411a <=( (not A169)  and  a56410a );
 a56415a <=( A201  and  (not A200) );
 a56416a <=( A199  and  a56415a );
 a56417a <=( a56416a  and  a56411a );
 a56421a <=( (not A234)  and  (not A233) );
 a56422a <=( A203  and  a56421a );
 a56425a <=( (not A266)  and  (not A265) );
 a56428a <=( (not A299)  and  (not A298) );
 a56429a <=( a56428a  and  a56425a );
 a56430a <=( a56429a  and  a56422a );
 a56434a <=( (not A166)  and  (not A167) );
 a56435a <=( (not A169)  and  a56434a );
 a56439a <=( A201  and  (not A200) );
 a56440a <=( A199  and  a56439a );
 a56441a <=( a56440a  and  a56435a );
 a56445a <=( (not A233)  and  A232 );
 a56446a <=( A203  and  a56445a );
 a56449a <=( A235  and  A234 );
 a56452a <=( A299  and  (not A298) );
 a56453a <=( a56452a  and  a56449a );
 a56454a <=( a56453a  and  a56446a );
 a56458a <=( (not A166)  and  (not A167) );
 a56459a <=( (not A169)  and  a56458a );
 a56463a <=( A201  and  (not A200) );
 a56464a <=( A199  and  a56463a );
 a56465a <=( a56464a  and  a56459a );
 a56469a <=( (not A233)  and  A232 );
 a56470a <=( A203  and  a56469a );
 a56473a <=( A235  and  A234 );
 a56476a <=( A266  and  (not A265) );
 a56477a <=( a56476a  and  a56473a );
 a56478a <=( a56477a  and  a56470a );
 a56482a <=( (not A166)  and  (not A167) );
 a56483a <=( (not A169)  and  a56482a );
 a56487a <=( A201  and  (not A200) );
 a56488a <=( A199  and  a56487a );
 a56489a <=( a56488a  and  a56483a );
 a56493a <=( (not A233)  and  A232 );
 a56494a <=( A203  and  a56493a );
 a56497a <=( A236  and  A234 );
 a56500a <=( A299  and  (not A298) );
 a56501a <=( a56500a  and  a56497a );
 a56502a <=( a56501a  and  a56494a );
 a56506a <=( (not A166)  and  (not A167) );
 a56507a <=( (not A169)  and  a56506a );
 a56511a <=( A201  and  (not A200) );
 a56512a <=( A199  and  a56511a );
 a56513a <=( a56512a  and  a56507a );
 a56517a <=( (not A233)  and  A232 );
 a56518a <=( A203  and  a56517a );
 a56521a <=( A236  and  A234 );
 a56524a <=( A266  and  (not A265) );
 a56525a <=( a56524a  and  a56521a );
 a56526a <=( a56525a  and  a56518a );
 a56530a <=( (not A166)  and  (not A167) );
 a56531a <=( (not A169)  and  a56530a );
 a56535a <=( A201  and  (not A200) );
 a56536a <=( A199  and  a56535a );
 a56537a <=( a56536a  and  a56531a );
 a56541a <=( (not A233)  and  (not A232) );
 a56542a <=( A203  and  a56541a );
 a56545a <=( A266  and  A265 );
 a56548a <=( (not A300)  and  A298 );
 a56549a <=( a56548a  and  a56545a );
 a56550a <=( a56549a  and  a56542a );
 a56554a <=( (not A166)  and  (not A167) );
 a56555a <=( (not A169)  and  a56554a );
 a56559a <=( A201  and  (not A200) );
 a56560a <=( A199  and  a56559a );
 a56561a <=( a56560a  and  a56555a );
 a56565a <=( (not A233)  and  (not A232) );
 a56566a <=( A203  and  a56565a );
 a56569a <=( A266  and  A265 );
 a56572a <=( A299  and  A298 );
 a56573a <=( a56572a  and  a56569a );
 a56574a <=( a56573a  and  a56566a );
 a56578a <=( (not A166)  and  (not A167) );
 a56579a <=( (not A169)  and  a56578a );
 a56583a <=( A201  and  (not A200) );
 a56584a <=( A199  and  a56583a );
 a56585a <=( a56584a  and  a56579a );
 a56589a <=( (not A233)  and  (not A232) );
 a56590a <=( A203  and  a56589a );
 a56593a <=( A266  and  A265 );
 a56596a <=( (not A299)  and  (not A298) );
 a56597a <=( a56596a  and  a56593a );
 a56598a <=( a56597a  and  a56590a );
 a56602a <=( (not A166)  and  (not A167) );
 a56603a <=( (not A169)  and  a56602a );
 a56607a <=( A201  and  (not A200) );
 a56608a <=( A199  and  a56607a );
 a56609a <=( a56608a  and  a56603a );
 a56613a <=( (not A233)  and  (not A232) );
 a56614a <=( A203  and  a56613a );
 a56617a <=( (not A267)  and  (not A266) );
 a56620a <=( (not A300)  and  A298 );
 a56621a <=( a56620a  and  a56617a );
 a56622a <=( a56621a  and  a56614a );
 a56626a <=( (not A166)  and  (not A167) );
 a56627a <=( (not A169)  and  a56626a );
 a56631a <=( A201  and  (not A200) );
 a56632a <=( A199  and  a56631a );
 a56633a <=( a56632a  and  a56627a );
 a56637a <=( (not A233)  and  (not A232) );
 a56638a <=( A203  and  a56637a );
 a56641a <=( (not A267)  and  (not A266) );
 a56644a <=( A299  and  A298 );
 a56645a <=( a56644a  and  a56641a );
 a56646a <=( a56645a  and  a56638a );
 a56650a <=( (not A166)  and  (not A167) );
 a56651a <=( (not A169)  and  a56650a );
 a56655a <=( A201  and  (not A200) );
 a56656a <=( A199  and  a56655a );
 a56657a <=( a56656a  and  a56651a );
 a56661a <=( (not A233)  and  (not A232) );
 a56662a <=( A203  and  a56661a );
 a56665a <=( (not A267)  and  (not A266) );
 a56668a <=( (not A299)  and  (not A298) );
 a56669a <=( a56668a  and  a56665a );
 a56670a <=( a56669a  and  a56662a );
 a56674a <=( (not A166)  and  (not A167) );
 a56675a <=( (not A169)  and  a56674a );
 a56679a <=( A201  and  (not A200) );
 a56680a <=( A199  and  a56679a );
 a56681a <=( a56680a  and  a56675a );
 a56685a <=( (not A233)  and  (not A232) );
 a56686a <=( A203  and  a56685a );
 a56689a <=( (not A266)  and  (not A265) );
 a56692a <=( (not A300)  and  A298 );
 a56693a <=( a56692a  and  a56689a );
 a56694a <=( a56693a  and  a56686a );
 a56698a <=( (not A166)  and  (not A167) );
 a56699a <=( (not A169)  and  a56698a );
 a56703a <=( A201  and  (not A200) );
 a56704a <=( A199  and  a56703a );
 a56705a <=( a56704a  and  a56699a );
 a56709a <=( (not A233)  and  (not A232) );
 a56710a <=( A203  and  a56709a );
 a56713a <=( (not A266)  and  (not A265) );
 a56716a <=( A299  and  A298 );
 a56717a <=( a56716a  and  a56713a );
 a56718a <=( a56717a  and  a56710a );
 a56722a <=( (not A166)  and  (not A167) );
 a56723a <=( (not A169)  and  a56722a );
 a56727a <=( A201  and  (not A200) );
 a56728a <=( A199  and  a56727a );
 a56729a <=( a56728a  and  a56723a );
 a56733a <=( (not A233)  and  (not A232) );
 a56734a <=( A203  and  a56733a );
 a56737a <=( (not A266)  and  (not A265) );
 a56740a <=( (not A299)  and  (not A298) );
 a56741a <=( a56740a  and  a56737a );
 a56742a <=( a56741a  and  a56734a );
 a56746a <=( A167  and  (not A168) );
 a56747a <=( (not A169)  and  a56746a );
 a56751a <=( A200  and  (not A199) );
 a56752a <=( A166  and  a56751a );
 a56753a <=( a56752a  and  a56747a );
 a56757a <=( A265  and  A233 );
 a56758a <=( A232  and  a56757a );
 a56761a <=( (not A269)  and  (not A268) );
 a56764a <=( (not A300)  and  (not A299) );
 a56765a <=( a56764a  and  a56761a );
 a56766a <=( a56765a  and  a56758a );
 a56770a <=( A167  and  (not A168) );
 a56771a <=( (not A169)  and  a56770a );
 a56775a <=( A200  and  (not A199) );
 a56776a <=( A166  and  a56775a );
 a56777a <=( a56776a  and  a56771a );
 a56781a <=( A265  and  A233 );
 a56782a <=( A232  and  a56781a );
 a56785a <=( (not A269)  and  (not A268) );
 a56788a <=( A299  and  A298 );
 a56789a <=( a56788a  and  a56785a );
 a56790a <=( a56789a  and  a56782a );
 a56794a <=( A167  and  (not A168) );
 a56795a <=( (not A169)  and  a56794a );
 a56799a <=( A200  and  (not A199) );
 a56800a <=( A166  and  a56799a );
 a56801a <=( a56800a  and  a56795a );
 a56805a <=( A265  and  A233 );
 a56806a <=( A232  and  a56805a );
 a56809a <=( (not A269)  and  (not A268) );
 a56812a <=( (not A299)  and  (not A298) );
 a56813a <=( a56812a  and  a56809a );
 a56814a <=( a56813a  and  a56806a );
 a56818a <=( A167  and  (not A168) );
 a56819a <=( (not A169)  and  a56818a );
 a56823a <=( A200  and  (not A199) );
 a56824a <=( A166  and  a56823a );
 a56825a <=( a56824a  and  a56819a );
 a56829a <=( A265  and  A233 );
 a56830a <=( A232  and  a56829a );
 a56833a <=( (not A299)  and  (not A267) );
 a56836a <=( (not A302)  and  (not A301) );
 a56837a <=( a56836a  and  a56833a );
 a56838a <=( a56837a  and  a56830a );
 a56842a <=( A167  and  (not A168) );
 a56843a <=( (not A169)  and  a56842a );
 a56847a <=( A200  and  (not A199) );
 a56848a <=( A166  and  a56847a );
 a56849a <=( a56848a  and  a56843a );
 a56853a <=( A265  and  A233 );
 a56854a <=( A232  and  a56853a );
 a56857a <=( (not A299)  and  A266 );
 a56860a <=( (not A302)  and  (not A301) );
 a56861a <=( a56860a  and  a56857a );
 a56862a <=( a56861a  and  a56854a );
 a56866a <=( A167  and  (not A168) );
 a56867a <=( (not A169)  and  a56866a );
 a56871a <=( A200  and  (not A199) );
 a56872a <=( A166  and  a56871a );
 a56873a <=( a56872a  and  a56867a );
 a56877a <=( (not A265)  and  A233 );
 a56878a <=( A232  and  a56877a );
 a56881a <=( (not A299)  and  (not A266) );
 a56884a <=( (not A302)  and  (not A301) );
 a56885a <=( a56884a  and  a56881a );
 a56886a <=( a56885a  and  a56878a );
 a56890a <=( A167  and  (not A168) );
 a56891a <=( (not A169)  and  a56890a );
 a56895a <=( A200  and  (not A199) );
 a56896a <=( A166  and  a56895a );
 a56897a <=( a56896a  and  a56891a );
 a56901a <=( (not A236)  and  (not A235) );
 a56902a <=( (not A233)  and  a56901a );
 a56905a <=( A266  and  A265 );
 a56908a <=( (not A300)  and  A298 );
 a56909a <=( a56908a  and  a56905a );
 a56910a <=( a56909a  and  a56902a );
 a56914a <=( A167  and  (not A168) );
 a56915a <=( (not A169)  and  a56914a );
 a56919a <=( A200  and  (not A199) );
 a56920a <=( A166  and  a56919a );
 a56921a <=( a56920a  and  a56915a );
 a56925a <=( (not A236)  and  (not A235) );
 a56926a <=( (not A233)  and  a56925a );
 a56929a <=( A266  and  A265 );
 a56932a <=( A299  and  A298 );
 a56933a <=( a56932a  and  a56929a );
 a56934a <=( a56933a  and  a56926a );
 a56938a <=( A167  and  (not A168) );
 a56939a <=( (not A169)  and  a56938a );
 a56943a <=( A200  and  (not A199) );
 a56944a <=( A166  and  a56943a );
 a56945a <=( a56944a  and  a56939a );
 a56949a <=( (not A236)  and  (not A235) );
 a56950a <=( (not A233)  and  a56949a );
 a56953a <=( A266  and  A265 );
 a56956a <=( (not A299)  and  (not A298) );
 a56957a <=( a56956a  and  a56953a );
 a56958a <=( a56957a  and  a56950a );
 a56962a <=( A167  and  (not A168) );
 a56963a <=( (not A169)  and  a56962a );
 a56967a <=( A200  and  (not A199) );
 a56968a <=( A166  and  a56967a );
 a56969a <=( a56968a  and  a56963a );
 a56973a <=( (not A236)  and  (not A235) );
 a56974a <=( (not A233)  and  a56973a );
 a56977a <=( (not A267)  and  (not A266) );
 a56980a <=( (not A300)  and  A298 );
 a56981a <=( a56980a  and  a56977a );
 a56982a <=( a56981a  and  a56974a );
 a56986a <=( A167  and  (not A168) );
 a56987a <=( (not A169)  and  a56986a );
 a56991a <=( A200  and  (not A199) );
 a56992a <=( A166  and  a56991a );
 a56993a <=( a56992a  and  a56987a );
 a56997a <=( (not A236)  and  (not A235) );
 a56998a <=( (not A233)  and  a56997a );
 a57001a <=( (not A267)  and  (not A266) );
 a57004a <=( A299  and  A298 );
 a57005a <=( a57004a  and  a57001a );
 a57006a <=( a57005a  and  a56998a );
 a57010a <=( A167  and  (not A168) );
 a57011a <=( (not A169)  and  a57010a );
 a57015a <=( A200  and  (not A199) );
 a57016a <=( A166  and  a57015a );
 a57017a <=( a57016a  and  a57011a );
 a57021a <=( (not A236)  and  (not A235) );
 a57022a <=( (not A233)  and  a57021a );
 a57025a <=( (not A267)  and  (not A266) );
 a57028a <=( (not A299)  and  (not A298) );
 a57029a <=( a57028a  and  a57025a );
 a57030a <=( a57029a  and  a57022a );
 a57034a <=( A167  and  (not A168) );
 a57035a <=( (not A169)  and  a57034a );
 a57039a <=( A200  and  (not A199) );
 a57040a <=( A166  and  a57039a );
 a57041a <=( a57040a  and  a57035a );
 a57045a <=( (not A236)  and  (not A235) );
 a57046a <=( (not A233)  and  a57045a );
 a57049a <=( (not A266)  and  (not A265) );
 a57052a <=( (not A300)  and  A298 );
 a57053a <=( a57052a  and  a57049a );
 a57054a <=( a57053a  and  a57046a );
 a57058a <=( A167  and  (not A168) );
 a57059a <=( (not A169)  and  a57058a );
 a57063a <=( A200  and  (not A199) );
 a57064a <=( A166  and  a57063a );
 a57065a <=( a57064a  and  a57059a );
 a57069a <=( (not A236)  and  (not A235) );
 a57070a <=( (not A233)  and  a57069a );
 a57073a <=( (not A266)  and  (not A265) );
 a57076a <=( A299  and  A298 );
 a57077a <=( a57076a  and  a57073a );
 a57078a <=( a57077a  and  a57070a );
 a57082a <=( A167  and  (not A168) );
 a57083a <=( (not A169)  and  a57082a );
 a57087a <=( A200  and  (not A199) );
 a57088a <=( A166  and  a57087a );
 a57089a <=( a57088a  and  a57083a );
 a57093a <=( (not A236)  and  (not A235) );
 a57094a <=( (not A233)  and  a57093a );
 a57097a <=( (not A266)  and  (not A265) );
 a57100a <=( (not A299)  and  (not A298) );
 a57101a <=( a57100a  and  a57097a );
 a57102a <=( a57101a  and  a57094a );
 a57106a <=( A167  and  (not A168) );
 a57107a <=( (not A169)  and  a57106a );
 a57111a <=( A200  and  (not A199) );
 a57112a <=( A166  and  a57111a );
 a57113a <=( a57112a  and  a57107a );
 a57117a <=( A265  and  (not A234) );
 a57118a <=( (not A233)  and  a57117a );
 a57121a <=( A298  and  A266 );
 a57124a <=( (not A302)  and  (not A301) );
 a57125a <=( a57124a  and  a57121a );
 a57126a <=( a57125a  and  a57118a );
 a57130a <=( A167  and  (not A168) );
 a57131a <=( (not A169)  and  a57130a );
 a57135a <=( A200  and  (not A199) );
 a57136a <=( A166  and  a57135a );
 a57137a <=( a57136a  and  a57131a );
 a57141a <=( (not A266)  and  (not A234) );
 a57142a <=( (not A233)  and  a57141a );
 a57145a <=( (not A269)  and  (not A268) );
 a57148a <=( (not A300)  and  A298 );
 a57149a <=( a57148a  and  a57145a );
 a57150a <=( a57149a  and  a57142a );
 a57154a <=( A167  and  (not A168) );
 a57155a <=( (not A169)  and  a57154a );
 a57159a <=( A200  and  (not A199) );
 a57160a <=( A166  and  a57159a );
 a57161a <=( a57160a  and  a57155a );
 a57165a <=( (not A266)  and  (not A234) );
 a57166a <=( (not A233)  and  a57165a );
 a57169a <=( (not A269)  and  (not A268) );
 a57172a <=( A299  and  A298 );
 a57173a <=( a57172a  and  a57169a );
 a57174a <=( a57173a  and  a57166a );
 a57178a <=( A167  and  (not A168) );
 a57179a <=( (not A169)  and  a57178a );
 a57183a <=( A200  and  (not A199) );
 a57184a <=( A166  and  a57183a );
 a57185a <=( a57184a  and  a57179a );
 a57189a <=( (not A266)  and  (not A234) );
 a57190a <=( (not A233)  and  a57189a );
 a57193a <=( (not A269)  and  (not A268) );
 a57196a <=( (not A299)  and  (not A298) );
 a57197a <=( a57196a  and  a57193a );
 a57198a <=( a57197a  and  a57190a );
 a57202a <=( A167  and  (not A168) );
 a57203a <=( (not A169)  and  a57202a );
 a57207a <=( A200  and  (not A199) );
 a57208a <=( A166  and  a57207a );
 a57209a <=( a57208a  and  a57203a );
 a57213a <=( (not A266)  and  (not A234) );
 a57214a <=( (not A233)  and  a57213a );
 a57217a <=( A298  and  (not A267) );
 a57220a <=( (not A302)  and  (not A301) );
 a57221a <=( a57220a  and  a57217a );
 a57222a <=( a57221a  and  a57214a );
 a57226a <=( A167  and  (not A168) );
 a57227a <=( (not A169)  and  a57226a );
 a57231a <=( A200  and  (not A199) );
 a57232a <=( A166  and  a57231a );
 a57233a <=( a57232a  and  a57227a );
 a57237a <=( (not A265)  and  (not A234) );
 a57238a <=( (not A233)  and  a57237a );
 a57241a <=( A298  and  (not A266) );
 a57244a <=( (not A302)  and  (not A301) );
 a57245a <=( a57244a  and  a57241a );
 a57246a <=( a57245a  and  a57238a );
 a57250a <=( A167  and  (not A168) );
 a57251a <=( (not A169)  and  a57250a );
 a57255a <=( A200  and  (not A199) );
 a57256a <=( A166  and  a57255a );
 a57257a <=( a57256a  and  a57251a );
 a57261a <=( A265  and  (not A233) );
 a57262a <=( (not A232)  and  a57261a );
 a57265a <=( A298  and  A266 );
 a57268a <=( (not A302)  and  (not A301) );
 a57269a <=( a57268a  and  a57265a );
 a57270a <=( a57269a  and  a57262a );
 a57274a <=( A167  and  (not A168) );
 a57275a <=( (not A169)  and  a57274a );
 a57279a <=( A200  and  (not A199) );
 a57280a <=( A166  and  a57279a );
 a57281a <=( a57280a  and  a57275a );
 a57285a <=( (not A266)  and  (not A233) );
 a57286a <=( (not A232)  and  a57285a );
 a57289a <=( (not A269)  and  (not A268) );
 a57292a <=( (not A300)  and  A298 );
 a57293a <=( a57292a  and  a57289a );
 a57294a <=( a57293a  and  a57286a );
 a57298a <=( A167  and  (not A168) );
 a57299a <=( (not A169)  and  a57298a );
 a57303a <=( A200  and  (not A199) );
 a57304a <=( A166  and  a57303a );
 a57305a <=( a57304a  and  a57299a );
 a57309a <=( (not A266)  and  (not A233) );
 a57310a <=( (not A232)  and  a57309a );
 a57313a <=( (not A269)  and  (not A268) );
 a57316a <=( A299  and  A298 );
 a57317a <=( a57316a  and  a57313a );
 a57318a <=( a57317a  and  a57310a );
 a57322a <=( A167  and  (not A168) );
 a57323a <=( (not A169)  and  a57322a );
 a57327a <=( A200  and  (not A199) );
 a57328a <=( A166  and  a57327a );
 a57329a <=( a57328a  and  a57323a );
 a57333a <=( (not A266)  and  (not A233) );
 a57334a <=( (not A232)  and  a57333a );
 a57337a <=( (not A269)  and  (not A268) );
 a57340a <=( (not A299)  and  (not A298) );
 a57341a <=( a57340a  and  a57337a );
 a57342a <=( a57341a  and  a57334a );
 a57346a <=( A167  and  (not A168) );
 a57347a <=( (not A169)  and  a57346a );
 a57351a <=( A200  and  (not A199) );
 a57352a <=( A166  and  a57351a );
 a57353a <=( a57352a  and  a57347a );
 a57357a <=( (not A266)  and  (not A233) );
 a57358a <=( (not A232)  and  a57357a );
 a57361a <=( A298  and  (not A267) );
 a57364a <=( (not A302)  and  (not A301) );
 a57365a <=( a57364a  and  a57361a );
 a57366a <=( a57365a  and  a57358a );
 a57370a <=( A167  and  (not A168) );
 a57371a <=( (not A169)  and  a57370a );
 a57375a <=( A200  and  (not A199) );
 a57376a <=( A166  and  a57375a );
 a57377a <=( a57376a  and  a57371a );
 a57381a <=( (not A265)  and  (not A233) );
 a57382a <=( (not A232)  and  a57381a );
 a57385a <=( A298  and  (not A266) );
 a57388a <=( (not A302)  and  (not A301) );
 a57389a <=( a57388a  and  a57385a );
 a57390a <=( a57389a  and  a57382a );
 a57394a <=( A167  and  (not A169) );
 a57395a <=( A170  and  a57394a );
 a57399a <=( A200  and  A199 );
 a57400a <=( (not A166)  and  a57399a );
 a57401a <=( a57400a  and  a57395a );
 a57405a <=( A265  and  A233 );
 a57406a <=( A232  and  a57405a );
 a57409a <=( (not A269)  and  (not A268) );
 a57412a <=( (not A300)  and  (not A299) );
 a57413a <=( a57412a  and  a57409a );
 a57414a <=( a57413a  and  a57406a );
 a57418a <=( A167  and  (not A169) );
 a57419a <=( A170  and  a57418a );
 a57423a <=( A200  and  A199 );
 a57424a <=( (not A166)  and  a57423a );
 a57425a <=( a57424a  and  a57419a );
 a57429a <=( A265  and  A233 );
 a57430a <=( A232  and  a57429a );
 a57433a <=( (not A269)  and  (not A268) );
 a57436a <=( A299  and  A298 );
 a57437a <=( a57436a  and  a57433a );
 a57438a <=( a57437a  and  a57430a );
 a57442a <=( A167  and  (not A169) );
 a57443a <=( A170  and  a57442a );
 a57447a <=( A200  and  A199 );
 a57448a <=( (not A166)  and  a57447a );
 a57449a <=( a57448a  and  a57443a );
 a57453a <=( A265  and  A233 );
 a57454a <=( A232  and  a57453a );
 a57457a <=( (not A269)  and  (not A268) );
 a57460a <=( (not A299)  and  (not A298) );
 a57461a <=( a57460a  and  a57457a );
 a57462a <=( a57461a  and  a57454a );
 a57466a <=( A167  and  (not A169) );
 a57467a <=( A170  and  a57466a );
 a57471a <=( A200  and  A199 );
 a57472a <=( (not A166)  and  a57471a );
 a57473a <=( a57472a  and  a57467a );
 a57477a <=( A265  and  A233 );
 a57478a <=( A232  and  a57477a );
 a57481a <=( (not A299)  and  (not A267) );
 a57484a <=( (not A302)  and  (not A301) );
 a57485a <=( a57484a  and  a57481a );
 a57486a <=( a57485a  and  a57478a );
 a57490a <=( A167  and  (not A169) );
 a57491a <=( A170  and  a57490a );
 a57495a <=( A200  and  A199 );
 a57496a <=( (not A166)  and  a57495a );
 a57497a <=( a57496a  and  a57491a );
 a57501a <=( A265  and  A233 );
 a57502a <=( A232  and  a57501a );
 a57505a <=( (not A299)  and  A266 );
 a57508a <=( (not A302)  and  (not A301) );
 a57509a <=( a57508a  and  a57505a );
 a57510a <=( a57509a  and  a57502a );
 a57514a <=( A167  and  (not A169) );
 a57515a <=( A170  and  a57514a );
 a57519a <=( A200  and  A199 );
 a57520a <=( (not A166)  and  a57519a );
 a57521a <=( a57520a  and  a57515a );
 a57525a <=( (not A265)  and  A233 );
 a57526a <=( A232  and  a57525a );
 a57529a <=( (not A299)  and  (not A266) );
 a57532a <=( (not A302)  and  (not A301) );
 a57533a <=( a57532a  and  a57529a );
 a57534a <=( a57533a  and  a57526a );
 a57538a <=( A167  and  (not A169) );
 a57539a <=( A170  and  a57538a );
 a57543a <=( A200  and  A199 );
 a57544a <=( (not A166)  and  a57543a );
 a57545a <=( a57544a  and  a57539a );
 a57549a <=( (not A236)  and  (not A235) );
 a57550a <=( (not A233)  and  a57549a );
 a57553a <=( A266  and  A265 );
 a57556a <=( (not A300)  and  A298 );
 a57557a <=( a57556a  and  a57553a );
 a57558a <=( a57557a  and  a57550a );
 a57562a <=( A167  and  (not A169) );
 a57563a <=( A170  and  a57562a );
 a57567a <=( A200  and  A199 );
 a57568a <=( (not A166)  and  a57567a );
 a57569a <=( a57568a  and  a57563a );
 a57573a <=( (not A236)  and  (not A235) );
 a57574a <=( (not A233)  and  a57573a );
 a57577a <=( A266  and  A265 );
 a57580a <=( A299  and  A298 );
 a57581a <=( a57580a  and  a57577a );
 a57582a <=( a57581a  and  a57574a );
 a57586a <=( A167  and  (not A169) );
 a57587a <=( A170  and  a57586a );
 a57591a <=( A200  and  A199 );
 a57592a <=( (not A166)  and  a57591a );
 a57593a <=( a57592a  and  a57587a );
 a57597a <=( (not A236)  and  (not A235) );
 a57598a <=( (not A233)  and  a57597a );
 a57601a <=( A266  and  A265 );
 a57604a <=( (not A299)  and  (not A298) );
 a57605a <=( a57604a  and  a57601a );
 a57606a <=( a57605a  and  a57598a );
 a57610a <=( A167  and  (not A169) );
 a57611a <=( A170  and  a57610a );
 a57615a <=( A200  and  A199 );
 a57616a <=( (not A166)  and  a57615a );
 a57617a <=( a57616a  and  a57611a );
 a57621a <=( (not A236)  and  (not A235) );
 a57622a <=( (not A233)  and  a57621a );
 a57625a <=( (not A267)  and  (not A266) );
 a57628a <=( (not A300)  and  A298 );
 a57629a <=( a57628a  and  a57625a );
 a57630a <=( a57629a  and  a57622a );
 a57634a <=( A167  and  (not A169) );
 a57635a <=( A170  and  a57634a );
 a57639a <=( A200  and  A199 );
 a57640a <=( (not A166)  and  a57639a );
 a57641a <=( a57640a  and  a57635a );
 a57645a <=( (not A236)  and  (not A235) );
 a57646a <=( (not A233)  and  a57645a );
 a57649a <=( (not A267)  and  (not A266) );
 a57652a <=( A299  and  A298 );
 a57653a <=( a57652a  and  a57649a );
 a57654a <=( a57653a  and  a57646a );
 a57658a <=( A167  and  (not A169) );
 a57659a <=( A170  and  a57658a );
 a57663a <=( A200  and  A199 );
 a57664a <=( (not A166)  and  a57663a );
 a57665a <=( a57664a  and  a57659a );
 a57669a <=( (not A236)  and  (not A235) );
 a57670a <=( (not A233)  and  a57669a );
 a57673a <=( (not A267)  and  (not A266) );
 a57676a <=( (not A299)  and  (not A298) );
 a57677a <=( a57676a  and  a57673a );
 a57678a <=( a57677a  and  a57670a );
 a57682a <=( A167  and  (not A169) );
 a57683a <=( A170  and  a57682a );
 a57687a <=( A200  and  A199 );
 a57688a <=( (not A166)  and  a57687a );
 a57689a <=( a57688a  and  a57683a );
 a57693a <=( (not A236)  and  (not A235) );
 a57694a <=( (not A233)  and  a57693a );
 a57697a <=( (not A266)  and  (not A265) );
 a57700a <=( (not A300)  and  A298 );
 a57701a <=( a57700a  and  a57697a );
 a57702a <=( a57701a  and  a57694a );
 a57706a <=( A167  and  (not A169) );
 a57707a <=( A170  and  a57706a );
 a57711a <=( A200  and  A199 );
 a57712a <=( (not A166)  and  a57711a );
 a57713a <=( a57712a  and  a57707a );
 a57717a <=( (not A236)  and  (not A235) );
 a57718a <=( (not A233)  and  a57717a );
 a57721a <=( (not A266)  and  (not A265) );
 a57724a <=( A299  and  A298 );
 a57725a <=( a57724a  and  a57721a );
 a57726a <=( a57725a  and  a57718a );
 a57730a <=( A167  and  (not A169) );
 a57731a <=( A170  and  a57730a );
 a57735a <=( A200  and  A199 );
 a57736a <=( (not A166)  and  a57735a );
 a57737a <=( a57736a  and  a57731a );
 a57741a <=( (not A236)  and  (not A235) );
 a57742a <=( (not A233)  and  a57741a );
 a57745a <=( (not A266)  and  (not A265) );
 a57748a <=( (not A299)  and  (not A298) );
 a57749a <=( a57748a  and  a57745a );
 a57750a <=( a57749a  and  a57742a );
 a57754a <=( A167  and  (not A169) );
 a57755a <=( A170  and  a57754a );
 a57759a <=( A200  and  A199 );
 a57760a <=( (not A166)  and  a57759a );
 a57761a <=( a57760a  and  a57755a );
 a57765a <=( A265  and  (not A234) );
 a57766a <=( (not A233)  and  a57765a );
 a57769a <=( A298  and  A266 );
 a57772a <=( (not A302)  and  (not A301) );
 a57773a <=( a57772a  and  a57769a );
 a57774a <=( a57773a  and  a57766a );
 a57778a <=( A167  and  (not A169) );
 a57779a <=( A170  and  a57778a );
 a57783a <=( A200  and  A199 );
 a57784a <=( (not A166)  and  a57783a );
 a57785a <=( a57784a  and  a57779a );
 a57789a <=( (not A266)  and  (not A234) );
 a57790a <=( (not A233)  and  a57789a );
 a57793a <=( (not A269)  and  (not A268) );
 a57796a <=( (not A300)  and  A298 );
 a57797a <=( a57796a  and  a57793a );
 a57798a <=( a57797a  and  a57790a );
 a57802a <=( A167  and  (not A169) );
 a57803a <=( A170  and  a57802a );
 a57807a <=( A200  and  A199 );
 a57808a <=( (not A166)  and  a57807a );
 a57809a <=( a57808a  and  a57803a );
 a57813a <=( (not A266)  and  (not A234) );
 a57814a <=( (not A233)  and  a57813a );
 a57817a <=( (not A269)  and  (not A268) );
 a57820a <=( A299  and  A298 );
 a57821a <=( a57820a  and  a57817a );
 a57822a <=( a57821a  and  a57814a );
 a57826a <=( A167  and  (not A169) );
 a57827a <=( A170  and  a57826a );
 a57831a <=( A200  and  A199 );
 a57832a <=( (not A166)  and  a57831a );
 a57833a <=( a57832a  and  a57827a );
 a57837a <=( (not A266)  and  (not A234) );
 a57838a <=( (not A233)  and  a57837a );
 a57841a <=( (not A269)  and  (not A268) );
 a57844a <=( (not A299)  and  (not A298) );
 a57845a <=( a57844a  and  a57841a );
 a57846a <=( a57845a  and  a57838a );
 a57850a <=( A167  and  (not A169) );
 a57851a <=( A170  and  a57850a );
 a57855a <=( A200  and  A199 );
 a57856a <=( (not A166)  and  a57855a );
 a57857a <=( a57856a  and  a57851a );
 a57861a <=( (not A266)  and  (not A234) );
 a57862a <=( (not A233)  and  a57861a );
 a57865a <=( A298  and  (not A267) );
 a57868a <=( (not A302)  and  (not A301) );
 a57869a <=( a57868a  and  a57865a );
 a57870a <=( a57869a  and  a57862a );
 a57874a <=( A167  and  (not A169) );
 a57875a <=( A170  and  a57874a );
 a57879a <=( A200  and  A199 );
 a57880a <=( (not A166)  and  a57879a );
 a57881a <=( a57880a  and  a57875a );
 a57885a <=( (not A265)  and  (not A234) );
 a57886a <=( (not A233)  and  a57885a );
 a57889a <=( A298  and  (not A266) );
 a57892a <=( (not A302)  and  (not A301) );
 a57893a <=( a57892a  and  a57889a );
 a57894a <=( a57893a  and  a57886a );
 a57898a <=( A167  and  (not A169) );
 a57899a <=( A170  and  a57898a );
 a57903a <=( A200  and  A199 );
 a57904a <=( (not A166)  and  a57903a );
 a57905a <=( a57904a  and  a57899a );
 a57909a <=( A265  and  (not A233) );
 a57910a <=( (not A232)  and  a57909a );
 a57913a <=( A298  and  A266 );
 a57916a <=( (not A302)  and  (not A301) );
 a57917a <=( a57916a  and  a57913a );
 a57918a <=( a57917a  and  a57910a );
 a57922a <=( A167  and  (not A169) );
 a57923a <=( A170  and  a57922a );
 a57927a <=( A200  and  A199 );
 a57928a <=( (not A166)  and  a57927a );
 a57929a <=( a57928a  and  a57923a );
 a57933a <=( (not A266)  and  (not A233) );
 a57934a <=( (not A232)  and  a57933a );
 a57937a <=( (not A269)  and  (not A268) );
 a57940a <=( (not A300)  and  A298 );
 a57941a <=( a57940a  and  a57937a );
 a57942a <=( a57941a  and  a57934a );
 a57946a <=( A167  and  (not A169) );
 a57947a <=( A170  and  a57946a );
 a57951a <=( A200  and  A199 );
 a57952a <=( (not A166)  and  a57951a );
 a57953a <=( a57952a  and  a57947a );
 a57957a <=( (not A266)  and  (not A233) );
 a57958a <=( (not A232)  and  a57957a );
 a57961a <=( (not A269)  and  (not A268) );
 a57964a <=( A299  and  A298 );
 a57965a <=( a57964a  and  a57961a );
 a57966a <=( a57965a  and  a57958a );
 a57970a <=( A167  and  (not A169) );
 a57971a <=( A170  and  a57970a );
 a57975a <=( A200  and  A199 );
 a57976a <=( (not A166)  and  a57975a );
 a57977a <=( a57976a  and  a57971a );
 a57981a <=( (not A266)  and  (not A233) );
 a57982a <=( (not A232)  and  a57981a );
 a57985a <=( (not A269)  and  (not A268) );
 a57988a <=( (not A299)  and  (not A298) );
 a57989a <=( a57988a  and  a57985a );
 a57990a <=( a57989a  and  a57982a );
 a57994a <=( A167  and  (not A169) );
 a57995a <=( A170  and  a57994a );
 a57999a <=( A200  and  A199 );
 a58000a <=( (not A166)  and  a57999a );
 a58001a <=( a58000a  and  a57995a );
 a58005a <=( (not A266)  and  (not A233) );
 a58006a <=( (not A232)  and  a58005a );
 a58009a <=( A298  and  (not A267) );
 a58012a <=( (not A302)  and  (not A301) );
 a58013a <=( a58012a  and  a58009a );
 a58014a <=( a58013a  and  a58006a );
 a58018a <=( A167  and  (not A169) );
 a58019a <=( A170  and  a58018a );
 a58023a <=( A200  and  A199 );
 a58024a <=( (not A166)  and  a58023a );
 a58025a <=( a58024a  and  a58019a );
 a58029a <=( (not A265)  and  (not A233) );
 a58030a <=( (not A232)  and  a58029a );
 a58033a <=( A298  and  (not A266) );
 a58036a <=( (not A302)  and  (not A301) );
 a58037a <=( a58036a  and  a58033a );
 a58038a <=( a58037a  and  a58030a );
 a58042a <=( A167  and  (not A169) );
 a58043a <=( A170  and  a58042a );
 a58047a <=( (not A202)  and  (not A200) );
 a58048a <=( (not A166)  and  a58047a );
 a58049a <=( a58048a  and  a58043a );
 a58053a <=( A233  and  A232 );
 a58054a <=( (not A203)  and  a58053a );
 a58057a <=( (not A267)  and  A265 );
 a58060a <=( (not A300)  and  (not A299) );
 a58061a <=( a58060a  and  a58057a );
 a58062a <=( a58061a  and  a58054a );
 a58066a <=( A167  and  (not A169) );
 a58067a <=( A170  and  a58066a );
 a58071a <=( (not A202)  and  (not A200) );
 a58072a <=( (not A166)  and  a58071a );
 a58073a <=( a58072a  and  a58067a );
 a58077a <=( A233  and  A232 );
 a58078a <=( (not A203)  and  a58077a );
 a58081a <=( (not A267)  and  A265 );
 a58084a <=( A299  and  A298 );
 a58085a <=( a58084a  and  a58081a );
 a58086a <=( a58085a  and  a58078a );
 a58090a <=( A167  and  (not A169) );
 a58091a <=( A170  and  a58090a );
 a58095a <=( (not A202)  and  (not A200) );
 a58096a <=( (not A166)  and  a58095a );
 a58097a <=( a58096a  and  a58091a );
 a58101a <=( A233  and  A232 );
 a58102a <=( (not A203)  and  a58101a );
 a58105a <=( (not A267)  and  A265 );
 a58108a <=( (not A299)  and  (not A298) );
 a58109a <=( a58108a  and  a58105a );
 a58110a <=( a58109a  and  a58102a );
 a58114a <=( A167  and  (not A169) );
 a58115a <=( A170  and  a58114a );
 a58119a <=( (not A202)  and  (not A200) );
 a58120a <=( (not A166)  and  a58119a );
 a58121a <=( a58120a  and  a58115a );
 a58125a <=( A233  and  A232 );
 a58126a <=( (not A203)  and  a58125a );
 a58129a <=( A266  and  A265 );
 a58132a <=( (not A300)  and  (not A299) );
 a58133a <=( a58132a  and  a58129a );
 a58134a <=( a58133a  and  a58126a );
 a58138a <=( A167  and  (not A169) );
 a58139a <=( A170  and  a58138a );
 a58143a <=( (not A202)  and  (not A200) );
 a58144a <=( (not A166)  and  a58143a );
 a58145a <=( a58144a  and  a58139a );
 a58149a <=( A233  and  A232 );
 a58150a <=( (not A203)  and  a58149a );
 a58153a <=( A266  and  A265 );
 a58156a <=( A299  and  A298 );
 a58157a <=( a58156a  and  a58153a );
 a58158a <=( a58157a  and  a58150a );
 a58162a <=( A167  and  (not A169) );
 a58163a <=( A170  and  a58162a );
 a58167a <=( (not A202)  and  (not A200) );
 a58168a <=( (not A166)  and  a58167a );
 a58169a <=( a58168a  and  a58163a );
 a58173a <=( A233  and  A232 );
 a58174a <=( (not A203)  and  a58173a );
 a58177a <=( A266  and  A265 );
 a58180a <=( (not A299)  and  (not A298) );
 a58181a <=( a58180a  and  a58177a );
 a58182a <=( a58181a  and  a58174a );
 a58186a <=( A167  and  (not A169) );
 a58187a <=( A170  and  a58186a );
 a58191a <=( (not A202)  and  (not A200) );
 a58192a <=( (not A166)  and  a58191a );
 a58193a <=( a58192a  and  a58187a );
 a58197a <=( A233  and  A232 );
 a58198a <=( (not A203)  and  a58197a );
 a58201a <=( (not A266)  and  (not A265) );
 a58204a <=( (not A300)  and  (not A299) );
 a58205a <=( a58204a  and  a58201a );
 a58206a <=( a58205a  and  a58198a );
 a58210a <=( A167  and  (not A169) );
 a58211a <=( A170  and  a58210a );
 a58215a <=( (not A202)  and  (not A200) );
 a58216a <=( (not A166)  and  a58215a );
 a58217a <=( a58216a  and  a58211a );
 a58221a <=( A233  and  A232 );
 a58222a <=( (not A203)  and  a58221a );
 a58225a <=( (not A266)  and  (not A265) );
 a58228a <=( A299  and  A298 );
 a58229a <=( a58228a  and  a58225a );
 a58230a <=( a58229a  and  a58222a );
 a58234a <=( A167  and  (not A169) );
 a58235a <=( A170  and  a58234a );
 a58239a <=( (not A202)  and  (not A200) );
 a58240a <=( (not A166)  and  a58239a );
 a58241a <=( a58240a  and  a58235a );
 a58245a <=( A233  and  A232 );
 a58246a <=( (not A203)  and  a58245a );
 a58249a <=( (not A266)  and  (not A265) );
 a58252a <=( (not A299)  and  (not A298) );
 a58253a <=( a58252a  and  a58249a );
 a58254a <=( a58253a  and  a58246a );
 a58258a <=( A167  and  (not A169) );
 a58259a <=( A170  and  a58258a );
 a58263a <=( (not A202)  and  (not A200) );
 a58264a <=( (not A166)  and  a58263a );
 a58265a <=( a58264a  and  a58259a );
 a58269a <=( A233  and  (not A232) );
 a58270a <=( (not A203)  and  a58269a );
 a58273a <=( (not A299)  and  A298 );
 a58276a <=( A301  and  A300 );
 a58277a <=( a58276a  and  a58273a );
 a58278a <=( a58277a  and  a58270a );
 a58282a <=( A167  and  (not A169) );
 a58283a <=( A170  and  a58282a );
 a58287a <=( (not A202)  and  (not A200) );
 a58288a <=( (not A166)  and  a58287a );
 a58289a <=( a58288a  and  a58283a );
 a58293a <=( A233  and  (not A232) );
 a58294a <=( (not A203)  and  a58293a );
 a58297a <=( (not A299)  and  A298 );
 a58300a <=( A302  and  A300 );
 a58301a <=( a58300a  and  a58297a );
 a58302a <=( a58301a  and  a58294a );
 a58306a <=( A167  and  (not A169) );
 a58307a <=( A170  and  a58306a );
 a58311a <=( (not A202)  and  (not A200) );
 a58312a <=( (not A166)  and  a58311a );
 a58313a <=( a58312a  and  a58307a );
 a58317a <=( A233  and  (not A232) );
 a58318a <=( (not A203)  and  a58317a );
 a58321a <=( (not A266)  and  A265 );
 a58324a <=( A268  and  A267 );
 a58325a <=( a58324a  and  a58321a );
 a58326a <=( a58325a  and  a58318a );
 a58330a <=( A167  and  (not A169) );
 a58331a <=( A170  and  a58330a );
 a58335a <=( (not A202)  and  (not A200) );
 a58336a <=( (not A166)  and  a58335a );
 a58337a <=( a58336a  and  a58331a );
 a58341a <=( A233  and  (not A232) );
 a58342a <=( (not A203)  and  a58341a );
 a58345a <=( (not A266)  and  A265 );
 a58348a <=( A269  and  A267 );
 a58349a <=( a58348a  and  a58345a );
 a58350a <=( a58349a  and  a58342a );
 a58354a <=( A167  and  (not A169) );
 a58355a <=( A170  and  a58354a );
 a58359a <=( (not A202)  and  (not A200) );
 a58360a <=( (not A166)  and  a58359a );
 a58361a <=( a58360a  and  a58355a );
 a58365a <=( (not A234)  and  (not A233) );
 a58366a <=( (not A203)  and  a58365a );
 a58369a <=( A266  and  A265 );
 a58372a <=( (not A300)  and  A298 );
 a58373a <=( a58372a  and  a58369a );
 a58374a <=( a58373a  and  a58366a );
 a58378a <=( A167  and  (not A169) );
 a58379a <=( A170  and  a58378a );
 a58383a <=( (not A202)  and  (not A200) );
 a58384a <=( (not A166)  and  a58383a );
 a58385a <=( a58384a  and  a58379a );
 a58389a <=( (not A234)  and  (not A233) );
 a58390a <=( (not A203)  and  a58389a );
 a58393a <=( A266  and  A265 );
 a58396a <=( A299  and  A298 );
 a58397a <=( a58396a  and  a58393a );
 a58398a <=( a58397a  and  a58390a );
 a58402a <=( A167  and  (not A169) );
 a58403a <=( A170  and  a58402a );
 a58407a <=( (not A202)  and  (not A200) );
 a58408a <=( (not A166)  and  a58407a );
 a58409a <=( a58408a  and  a58403a );
 a58413a <=( (not A234)  and  (not A233) );
 a58414a <=( (not A203)  and  a58413a );
 a58417a <=( A266  and  A265 );
 a58420a <=( (not A299)  and  (not A298) );
 a58421a <=( a58420a  and  a58417a );
 a58422a <=( a58421a  and  a58414a );
 a58426a <=( A167  and  (not A169) );
 a58427a <=( A170  and  a58426a );
 a58431a <=( (not A202)  and  (not A200) );
 a58432a <=( (not A166)  and  a58431a );
 a58433a <=( a58432a  and  a58427a );
 a58437a <=( (not A234)  and  (not A233) );
 a58438a <=( (not A203)  and  a58437a );
 a58441a <=( (not A267)  and  (not A266) );
 a58444a <=( (not A300)  and  A298 );
 a58445a <=( a58444a  and  a58441a );
 a58446a <=( a58445a  and  a58438a );
 a58450a <=( A167  and  (not A169) );
 a58451a <=( A170  and  a58450a );
 a58455a <=( (not A202)  and  (not A200) );
 a58456a <=( (not A166)  and  a58455a );
 a58457a <=( a58456a  and  a58451a );
 a58461a <=( (not A234)  and  (not A233) );
 a58462a <=( (not A203)  and  a58461a );
 a58465a <=( (not A267)  and  (not A266) );
 a58468a <=( A299  and  A298 );
 a58469a <=( a58468a  and  a58465a );
 a58470a <=( a58469a  and  a58462a );
 a58474a <=( A167  and  (not A169) );
 a58475a <=( A170  and  a58474a );
 a58479a <=( (not A202)  and  (not A200) );
 a58480a <=( (not A166)  and  a58479a );
 a58481a <=( a58480a  and  a58475a );
 a58485a <=( (not A234)  and  (not A233) );
 a58486a <=( (not A203)  and  a58485a );
 a58489a <=( (not A267)  and  (not A266) );
 a58492a <=( (not A299)  and  (not A298) );
 a58493a <=( a58492a  and  a58489a );
 a58494a <=( a58493a  and  a58486a );
 a58498a <=( A167  and  (not A169) );
 a58499a <=( A170  and  a58498a );
 a58503a <=( (not A202)  and  (not A200) );
 a58504a <=( (not A166)  and  a58503a );
 a58505a <=( a58504a  and  a58499a );
 a58509a <=( (not A234)  and  (not A233) );
 a58510a <=( (not A203)  and  a58509a );
 a58513a <=( (not A266)  and  (not A265) );
 a58516a <=( (not A300)  and  A298 );
 a58517a <=( a58516a  and  a58513a );
 a58518a <=( a58517a  and  a58510a );
 a58522a <=( A167  and  (not A169) );
 a58523a <=( A170  and  a58522a );
 a58527a <=( (not A202)  and  (not A200) );
 a58528a <=( (not A166)  and  a58527a );
 a58529a <=( a58528a  and  a58523a );
 a58533a <=( (not A234)  and  (not A233) );
 a58534a <=( (not A203)  and  a58533a );
 a58537a <=( (not A266)  and  (not A265) );
 a58540a <=( A299  and  A298 );
 a58541a <=( a58540a  and  a58537a );
 a58542a <=( a58541a  and  a58534a );
 a58546a <=( A167  and  (not A169) );
 a58547a <=( A170  and  a58546a );
 a58551a <=( (not A202)  and  (not A200) );
 a58552a <=( (not A166)  and  a58551a );
 a58553a <=( a58552a  and  a58547a );
 a58557a <=( (not A234)  and  (not A233) );
 a58558a <=( (not A203)  and  a58557a );
 a58561a <=( (not A266)  and  (not A265) );
 a58564a <=( (not A299)  and  (not A298) );
 a58565a <=( a58564a  and  a58561a );
 a58566a <=( a58565a  and  a58558a );
 a58570a <=( A167  and  (not A169) );
 a58571a <=( A170  and  a58570a );
 a58575a <=( (not A202)  and  (not A200) );
 a58576a <=( (not A166)  and  a58575a );
 a58577a <=( a58576a  and  a58571a );
 a58581a <=( (not A233)  and  A232 );
 a58582a <=( (not A203)  and  a58581a );
 a58585a <=( A235  and  A234 );
 a58588a <=( A299  and  (not A298) );
 a58589a <=( a58588a  and  a58585a );
 a58590a <=( a58589a  and  a58582a );
 a58594a <=( A167  and  (not A169) );
 a58595a <=( A170  and  a58594a );
 a58599a <=( (not A202)  and  (not A200) );
 a58600a <=( (not A166)  and  a58599a );
 a58601a <=( a58600a  and  a58595a );
 a58605a <=( (not A233)  and  A232 );
 a58606a <=( (not A203)  and  a58605a );
 a58609a <=( A235  and  A234 );
 a58612a <=( A266  and  (not A265) );
 a58613a <=( a58612a  and  a58609a );
 a58614a <=( a58613a  and  a58606a );
 a58618a <=( A167  and  (not A169) );
 a58619a <=( A170  and  a58618a );
 a58623a <=( (not A202)  and  (not A200) );
 a58624a <=( (not A166)  and  a58623a );
 a58625a <=( a58624a  and  a58619a );
 a58629a <=( (not A233)  and  A232 );
 a58630a <=( (not A203)  and  a58629a );
 a58633a <=( A236  and  A234 );
 a58636a <=( A299  and  (not A298) );
 a58637a <=( a58636a  and  a58633a );
 a58638a <=( a58637a  and  a58630a );
 a58642a <=( A167  and  (not A169) );
 a58643a <=( A170  and  a58642a );
 a58647a <=( (not A202)  and  (not A200) );
 a58648a <=( (not A166)  and  a58647a );
 a58649a <=( a58648a  and  a58643a );
 a58653a <=( (not A233)  and  A232 );
 a58654a <=( (not A203)  and  a58653a );
 a58657a <=( A236  and  A234 );
 a58660a <=( A266  and  (not A265) );
 a58661a <=( a58660a  and  a58657a );
 a58662a <=( a58661a  and  a58654a );
 a58666a <=( A167  and  (not A169) );
 a58667a <=( A170  and  a58666a );
 a58671a <=( (not A202)  and  (not A200) );
 a58672a <=( (not A166)  and  a58671a );
 a58673a <=( a58672a  and  a58667a );
 a58677a <=( (not A233)  and  (not A232) );
 a58678a <=( (not A203)  and  a58677a );
 a58681a <=( A266  and  A265 );
 a58684a <=( (not A300)  and  A298 );
 a58685a <=( a58684a  and  a58681a );
 a58686a <=( a58685a  and  a58678a );
 a58690a <=( A167  and  (not A169) );
 a58691a <=( A170  and  a58690a );
 a58695a <=( (not A202)  and  (not A200) );
 a58696a <=( (not A166)  and  a58695a );
 a58697a <=( a58696a  and  a58691a );
 a58701a <=( (not A233)  and  (not A232) );
 a58702a <=( (not A203)  and  a58701a );
 a58705a <=( A266  and  A265 );
 a58708a <=( A299  and  A298 );
 a58709a <=( a58708a  and  a58705a );
 a58710a <=( a58709a  and  a58702a );
 a58714a <=( A167  and  (not A169) );
 a58715a <=( A170  and  a58714a );
 a58719a <=( (not A202)  and  (not A200) );
 a58720a <=( (not A166)  and  a58719a );
 a58721a <=( a58720a  and  a58715a );
 a58725a <=( (not A233)  and  (not A232) );
 a58726a <=( (not A203)  and  a58725a );
 a58729a <=( A266  and  A265 );
 a58732a <=( (not A299)  and  (not A298) );
 a58733a <=( a58732a  and  a58729a );
 a58734a <=( a58733a  and  a58726a );
 a58738a <=( A167  and  (not A169) );
 a58739a <=( A170  and  a58738a );
 a58743a <=( (not A202)  and  (not A200) );
 a58744a <=( (not A166)  and  a58743a );
 a58745a <=( a58744a  and  a58739a );
 a58749a <=( (not A233)  and  (not A232) );
 a58750a <=( (not A203)  and  a58749a );
 a58753a <=( (not A267)  and  (not A266) );
 a58756a <=( (not A300)  and  A298 );
 a58757a <=( a58756a  and  a58753a );
 a58758a <=( a58757a  and  a58750a );
 a58762a <=( A167  and  (not A169) );
 a58763a <=( A170  and  a58762a );
 a58767a <=( (not A202)  and  (not A200) );
 a58768a <=( (not A166)  and  a58767a );
 a58769a <=( a58768a  and  a58763a );
 a58773a <=( (not A233)  and  (not A232) );
 a58774a <=( (not A203)  and  a58773a );
 a58777a <=( (not A267)  and  (not A266) );
 a58780a <=( A299  and  A298 );
 a58781a <=( a58780a  and  a58777a );
 a58782a <=( a58781a  and  a58774a );
 a58786a <=( A167  and  (not A169) );
 a58787a <=( A170  and  a58786a );
 a58791a <=( (not A202)  and  (not A200) );
 a58792a <=( (not A166)  and  a58791a );
 a58793a <=( a58792a  and  a58787a );
 a58797a <=( (not A233)  and  (not A232) );
 a58798a <=( (not A203)  and  a58797a );
 a58801a <=( (not A267)  and  (not A266) );
 a58804a <=( (not A299)  and  (not A298) );
 a58805a <=( a58804a  and  a58801a );
 a58806a <=( a58805a  and  a58798a );
 a58810a <=( A167  and  (not A169) );
 a58811a <=( A170  and  a58810a );
 a58815a <=( (not A202)  and  (not A200) );
 a58816a <=( (not A166)  and  a58815a );
 a58817a <=( a58816a  and  a58811a );
 a58821a <=( (not A233)  and  (not A232) );
 a58822a <=( (not A203)  and  a58821a );
 a58825a <=( (not A266)  and  (not A265) );
 a58828a <=( (not A300)  and  A298 );
 a58829a <=( a58828a  and  a58825a );
 a58830a <=( a58829a  and  a58822a );
 a58834a <=( A167  and  (not A169) );
 a58835a <=( A170  and  a58834a );
 a58839a <=( (not A202)  and  (not A200) );
 a58840a <=( (not A166)  and  a58839a );
 a58841a <=( a58840a  and  a58835a );
 a58845a <=( (not A233)  and  (not A232) );
 a58846a <=( (not A203)  and  a58845a );
 a58849a <=( (not A266)  and  (not A265) );
 a58852a <=( A299  and  A298 );
 a58853a <=( a58852a  and  a58849a );
 a58854a <=( a58853a  and  a58846a );
 a58858a <=( A167  and  (not A169) );
 a58859a <=( A170  and  a58858a );
 a58863a <=( (not A202)  and  (not A200) );
 a58864a <=( (not A166)  and  a58863a );
 a58865a <=( a58864a  and  a58859a );
 a58869a <=( (not A233)  and  (not A232) );
 a58870a <=( (not A203)  and  a58869a );
 a58873a <=( (not A266)  and  (not A265) );
 a58876a <=( (not A299)  and  (not A298) );
 a58877a <=( a58876a  and  a58873a );
 a58878a <=( a58877a  and  a58870a );
 a58882a <=( A167  and  (not A169) );
 a58883a <=( A170  and  a58882a );
 a58887a <=( (not A201)  and  (not A200) );
 a58888a <=( (not A166)  and  a58887a );
 a58889a <=( a58888a  and  a58883a );
 a58893a <=( A265  and  A233 );
 a58894a <=( A232  and  a58893a );
 a58897a <=( (not A269)  and  (not A268) );
 a58900a <=( (not A300)  and  (not A299) );
 a58901a <=( a58900a  and  a58897a );
 a58902a <=( a58901a  and  a58894a );
 a58906a <=( A167  and  (not A169) );
 a58907a <=( A170  and  a58906a );
 a58911a <=( (not A201)  and  (not A200) );
 a58912a <=( (not A166)  and  a58911a );
 a58913a <=( a58912a  and  a58907a );
 a58917a <=( A265  and  A233 );
 a58918a <=( A232  and  a58917a );
 a58921a <=( (not A269)  and  (not A268) );
 a58924a <=( A299  and  A298 );
 a58925a <=( a58924a  and  a58921a );
 a58926a <=( a58925a  and  a58918a );
 a58930a <=( A167  and  (not A169) );
 a58931a <=( A170  and  a58930a );
 a58935a <=( (not A201)  and  (not A200) );
 a58936a <=( (not A166)  and  a58935a );
 a58937a <=( a58936a  and  a58931a );
 a58941a <=( A265  and  A233 );
 a58942a <=( A232  and  a58941a );
 a58945a <=( (not A269)  and  (not A268) );
 a58948a <=( (not A299)  and  (not A298) );
 a58949a <=( a58948a  and  a58945a );
 a58950a <=( a58949a  and  a58942a );
 a58954a <=( A167  and  (not A169) );
 a58955a <=( A170  and  a58954a );
 a58959a <=( (not A201)  and  (not A200) );
 a58960a <=( (not A166)  and  a58959a );
 a58961a <=( a58960a  and  a58955a );
 a58965a <=( A265  and  A233 );
 a58966a <=( A232  and  a58965a );
 a58969a <=( (not A299)  and  (not A267) );
 a58972a <=( (not A302)  and  (not A301) );
 a58973a <=( a58972a  and  a58969a );
 a58974a <=( a58973a  and  a58966a );
 a58978a <=( A167  and  (not A169) );
 a58979a <=( A170  and  a58978a );
 a58983a <=( (not A201)  and  (not A200) );
 a58984a <=( (not A166)  and  a58983a );
 a58985a <=( a58984a  and  a58979a );
 a58989a <=( A265  and  A233 );
 a58990a <=( A232  and  a58989a );
 a58993a <=( (not A299)  and  A266 );
 a58996a <=( (not A302)  and  (not A301) );
 a58997a <=( a58996a  and  a58993a );
 a58998a <=( a58997a  and  a58990a );
 a59002a <=( A167  and  (not A169) );
 a59003a <=( A170  and  a59002a );
 a59007a <=( (not A201)  and  (not A200) );
 a59008a <=( (not A166)  and  a59007a );
 a59009a <=( a59008a  and  a59003a );
 a59013a <=( (not A265)  and  A233 );
 a59014a <=( A232  and  a59013a );
 a59017a <=( (not A299)  and  (not A266) );
 a59020a <=( (not A302)  and  (not A301) );
 a59021a <=( a59020a  and  a59017a );
 a59022a <=( a59021a  and  a59014a );
 a59026a <=( A167  and  (not A169) );
 a59027a <=( A170  and  a59026a );
 a59031a <=( (not A201)  and  (not A200) );
 a59032a <=( (not A166)  and  a59031a );
 a59033a <=( a59032a  and  a59027a );
 a59037a <=( (not A236)  and  (not A235) );
 a59038a <=( (not A233)  and  a59037a );
 a59041a <=( A266  and  A265 );
 a59044a <=( (not A300)  and  A298 );
 a59045a <=( a59044a  and  a59041a );
 a59046a <=( a59045a  and  a59038a );
 a59050a <=( A167  and  (not A169) );
 a59051a <=( A170  and  a59050a );
 a59055a <=( (not A201)  and  (not A200) );
 a59056a <=( (not A166)  and  a59055a );
 a59057a <=( a59056a  and  a59051a );
 a59061a <=( (not A236)  and  (not A235) );
 a59062a <=( (not A233)  and  a59061a );
 a59065a <=( A266  and  A265 );
 a59068a <=( A299  and  A298 );
 a59069a <=( a59068a  and  a59065a );
 a59070a <=( a59069a  and  a59062a );
 a59074a <=( A167  and  (not A169) );
 a59075a <=( A170  and  a59074a );
 a59079a <=( (not A201)  and  (not A200) );
 a59080a <=( (not A166)  and  a59079a );
 a59081a <=( a59080a  and  a59075a );
 a59085a <=( (not A236)  and  (not A235) );
 a59086a <=( (not A233)  and  a59085a );
 a59089a <=( A266  and  A265 );
 a59092a <=( (not A299)  and  (not A298) );
 a59093a <=( a59092a  and  a59089a );
 a59094a <=( a59093a  and  a59086a );
 a59098a <=( A167  and  (not A169) );
 a59099a <=( A170  and  a59098a );
 a59103a <=( (not A201)  and  (not A200) );
 a59104a <=( (not A166)  and  a59103a );
 a59105a <=( a59104a  and  a59099a );
 a59109a <=( (not A236)  and  (not A235) );
 a59110a <=( (not A233)  and  a59109a );
 a59113a <=( (not A267)  and  (not A266) );
 a59116a <=( (not A300)  and  A298 );
 a59117a <=( a59116a  and  a59113a );
 a59118a <=( a59117a  and  a59110a );
 a59122a <=( A167  and  (not A169) );
 a59123a <=( A170  and  a59122a );
 a59127a <=( (not A201)  and  (not A200) );
 a59128a <=( (not A166)  and  a59127a );
 a59129a <=( a59128a  and  a59123a );
 a59133a <=( (not A236)  and  (not A235) );
 a59134a <=( (not A233)  and  a59133a );
 a59137a <=( (not A267)  and  (not A266) );
 a59140a <=( A299  and  A298 );
 a59141a <=( a59140a  and  a59137a );
 a59142a <=( a59141a  and  a59134a );
 a59146a <=( A167  and  (not A169) );
 a59147a <=( A170  and  a59146a );
 a59151a <=( (not A201)  and  (not A200) );
 a59152a <=( (not A166)  and  a59151a );
 a59153a <=( a59152a  and  a59147a );
 a59157a <=( (not A236)  and  (not A235) );
 a59158a <=( (not A233)  and  a59157a );
 a59161a <=( (not A267)  and  (not A266) );
 a59164a <=( (not A299)  and  (not A298) );
 a59165a <=( a59164a  and  a59161a );
 a59166a <=( a59165a  and  a59158a );
 a59170a <=( A167  and  (not A169) );
 a59171a <=( A170  and  a59170a );
 a59175a <=( (not A201)  and  (not A200) );
 a59176a <=( (not A166)  and  a59175a );
 a59177a <=( a59176a  and  a59171a );
 a59181a <=( (not A236)  and  (not A235) );
 a59182a <=( (not A233)  and  a59181a );
 a59185a <=( (not A266)  and  (not A265) );
 a59188a <=( (not A300)  and  A298 );
 a59189a <=( a59188a  and  a59185a );
 a59190a <=( a59189a  and  a59182a );
 a59194a <=( A167  and  (not A169) );
 a59195a <=( A170  and  a59194a );
 a59199a <=( (not A201)  and  (not A200) );
 a59200a <=( (not A166)  and  a59199a );
 a59201a <=( a59200a  and  a59195a );
 a59205a <=( (not A236)  and  (not A235) );
 a59206a <=( (not A233)  and  a59205a );
 a59209a <=( (not A266)  and  (not A265) );
 a59212a <=( A299  and  A298 );
 a59213a <=( a59212a  and  a59209a );
 a59214a <=( a59213a  and  a59206a );
 a59218a <=( A167  and  (not A169) );
 a59219a <=( A170  and  a59218a );
 a59223a <=( (not A201)  and  (not A200) );
 a59224a <=( (not A166)  and  a59223a );
 a59225a <=( a59224a  and  a59219a );
 a59229a <=( (not A236)  and  (not A235) );
 a59230a <=( (not A233)  and  a59229a );
 a59233a <=( (not A266)  and  (not A265) );
 a59236a <=( (not A299)  and  (not A298) );
 a59237a <=( a59236a  and  a59233a );
 a59238a <=( a59237a  and  a59230a );
 a59242a <=( A167  and  (not A169) );
 a59243a <=( A170  and  a59242a );
 a59247a <=( (not A201)  and  (not A200) );
 a59248a <=( (not A166)  and  a59247a );
 a59249a <=( a59248a  and  a59243a );
 a59253a <=( A265  and  (not A234) );
 a59254a <=( (not A233)  and  a59253a );
 a59257a <=( A298  and  A266 );
 a59260a <=( (not A302)  and  (not A301) );
 a59261a <=( a59260a  and  a59257a );
 a59262a <=( a59261a  and  a59254a );
 a59266a <=( A167  and  (not A169) );
 a59267a <=( A170  and  a59266a );
 a59271a <=( (not A201)  and  (not A200) );
 a59272a <=( (not A166)  and  a59271a );
 a59273a <=( a59272a  and  a59267a );
 a59277a <=( (not A266)  and  (not A234) );
 a59278a <=( (not A233)  and  a59277a );
 a59281a <=( (not A269)  and  (not A268) );
 a59284a <=( (not A300)  and  A298 );
 a59285a <=( a59284a  and  a59281a );
 a59286a <=( a59285a  and  a59278a );
 a59290a <=( A167  and  (not A169) );
 a59291a <=( A170  and  a59290a );
 a59295a <=( (not A201)  and  (not A200) );
 a59296a <=( (not A166)  and  a59295a );
 a59297a <=( a59296a  and  a59291a );
 a59301a <=( (not A266)  and  (not A234) );
 a59302a <=( (not A233)  and  a59301a );
 a59305a <=( (not A269)  and  (not A268) );
 a59308a <=( A299  and  A298 );
 a59309a <=( a59308a  and  a59305a );
 a59310a <=( a59309a  and  a59302a );
 a59314a <=( A167  and  (not A169) );
 a59315a <=( A170  and  a59314a );
 a59319a <=( (not A201)  and  (not A200) );
 a59320a <=( (not A166)  and  a59319a );
 a59321a <=( a59320a  and  a59315a );
 a59325a <=( (not A266)  and  (not A234) );
 a59326a <=( (not A233)  and  a59325a );
 a59329a <=( (not A269)  and  (not A268) );
 a59332a <=( (not A299)  and  (not A298) );
 a59333a <=( a59332a  and  a59329a );
 a59334a <=( a59333a  and  a59326a );
 a59338a <=( A167  and  (not A169) );
 a59339a <=( A170  and  a59338a );
 a59343a <=( (not A201)  and  (not A200) );
 a59344a <=( (not A166)  and  a59343a );
 a59345a <=( a59344a  and  a59339a );
 a59349a <=( (not A266)  and  (not A234) );
 a59350a <=( (not A233)  and  a59349a );
 a59353a <=( A298  and  (not A267) );
 a59356a <=( (not A302)  and  (not A301) );
 a59357a <=( a59356a  and  a59353a );
 a59358a <=( a59357a  and  a59350a );
 a59362a <=( A167  and  (not A169) );
 a59363a <=( A170  and  a59362a );
 a59367a <=( (not A201)  and  (not A200) );
 a59368a <=( (not A166)  and  a59367a );
 a59369a <=( a59368a  and  a59363a );
 a59373a <=( (not A265)  and  (not A234) );
 a59374a <=( (not A233)  and  a59373a );
 a59377a <=( A298  and  (not A266) );
 a59380a <=( (not A302)  and  (not A301) );
 a59381a <=( a59380a  and  a59377a );
 a59382a <=( a59381a  and  a59374a );
 a59386a <=( A167  and  (not A169) );
 a59387a <=( A170  and  a59386a );
 a59391a <=( (not A201)  and  (not A200) );
 a59392a <=( (not A166)  and  a59391a );
 a59393a <=( a59392a  and  a59387a );
 a59397a <=( A265  and  (not A233) );
 a59398a <=( (not A232)  and  a59397a );
 a59401a <=( A298  and  A266 );
 a59404a <=( (not A302)  and  (not A301) );
 a59405a <=( a59404a  and  a59401a );
 a59406a <=( a59405a  and  a59398a );
 a59410a <=( A167  and  (not A169) );
 a59411a <=( A170  and  a59410a );
 a59415a <=( (not A201)  and  (not A200) );
 a59416a <=( (not A166)  and  a59415a );
 a59417a <=( a59416a  and  a59411a );
 a59421a <=( (not A266)  and  (not A233) );
 a59422a <=( (not A232)  and  a59421a );
 a59425a <=( (not A269)  and  (not A268) );
 a59428a <=( (not A300)  and  A298 );
 a59429a <=( a59428a  and  a59425a );
 a59430a <=( a59429a  and  a59422a );
 a59434a <=( A167  and  (not A169) );
 a59435a <=( A170  and  a59434a );
 a59439a <=( (not A201)  and  (not A200) );
 a59440a <=( (not A166)  and  a59439a );
 a59441a <=( a59440a  and  a59435a );
 a59445a <=( (not A266)  and  (not A233) );
 a59446a <=( (not A232)  and  a59445a );
 a59449a <=( (not A269)  and  (not A268) );
 a59452a <=( A299  and  A298 );
 a59453a <=( a59452a  and  a59449a );
 a59454a <=( a59453a  and  a59446a );
 a59458a <=( A167  and  (not A169) );
 a59459a <=( A170  and  a59458a );
 a59463a <=( (not A201)  and  (not A200) );
 a59464a <=( (not A166)  and  a59463a );
 a59465a <=( a59464a  and  a59459a );
 a59469a <=( (not A266)  and  (not A233) );
 a59470a <=( (not A232)  and  a59469a );
 a59473a <=( (not A269)  and  (not A268) );
 a59476a <=( (not A299)  and  (not A298) );
 a59477a <=( a59476a  and  a59473a );
 a59478a <=( a59477a  and  a59470a );
 a59482a <=( A167  and  (not A169) );
 a59483a <=( A170  and  a59482a );
 a59487a <=( (not A201)  and  (not A200) );
 a59488a <=( (not A166)  and  a59487a );
 a59489a <=( a59488a  and  a59483a );
 a59493a <=( (not A266)  and  (not A233) );
 a59494a <=( (not A232)  and  a59493a );
 a59497a <=( A298  and  (not A267) );
 a59500a <=( (not A302)  and  (not A301) );
 a59501a <=( a59500a  and  a59497a );
 a59502a <=( a59501a  and  a59494a );
 a59506a <=( A167  and  (not A169) );
 a59507a <=( A170  and  a59506a );
 a59511a <=( (not A201)  and  (not A200) );
 a59512a <=( (not A166)  and  a59511a );
 a59513a <=( a59512a  and  a59507a );
 a59517a <=( (not A265)  and  (not A233) );
 a59518a <=( (not A232)  and  a59517a );
 a59521a <=( A298  and  (not A266) );
 a59524a <=( (not A302)  and  (not A301) );
 a59525a <=( a59524a  and  a59521a );
 a59526a <=( a59525a  and  a59518a );
 a59530a <=( A167  and  (not A169) );
 a59531a <=( A170  and  a59530a );
 a59535a <=( (not A200)  and  (not A199) );
 a59536a <=( (not A166)  and  a59535a );
 a59537a <=( a59536a  and  a59531a );
 a59541a <=( A265  and  A233 );
 a59542a <=( A232  and  a59541a );
 a59545a <=( (not A269)  and  (not A268) );
 a59548a <=( (not A300)  and  (not A299) );
 a59549a <=( a59548a  and  a59545a );
 a59550a <=( a59549a  and  a59542a );
 a59554a <=( A167  and  (not A169) );
 a59555a <=( A170  and  a59554a );
 a59559a <=( (not A200)  and  (not A199) );
 a59560a <=( (not A166)  and  a59559a );
 a59561a <=( a59560a  and  a59555a );
 a59565a <=( A265  and  A233 );
 a59566a <=( A232  and  a59565a );
 a59569a <=( (not A269)  and  (not A268) );
 a59572a <=( A299  and  A298 );
 a59573a <=( a59572a  and  a59569a );
 a59574a <=( a59573a  and  a59566a );
 a59578a <=( A167  and  (not A169) );
 a59579a <=( A170  and  a59578a );
 a59583a <=( (not A200)  and  (not A199) );
 a59584a <=( (not A166)  and  a59583a );
 a59585a <=( a59584a  and  a59579a );
 a59589a <=( A265  and  A233 );
 a59590a <=( A232  and  a59589a );
 a59593a <=( (not A269)  and  (not A268) );
 a59596a <=( (not A299)  and  (not A298) );
 a59597a <=( a59596a  and  a59593a );
 a59598a <=( a59597a  and  a59590a );
 a59602a <=( A167  and  (not A169) );
 a59603a <=( A170  and  a59602a );
 a59607a <=( (not A200)  and  (not A199) );
 a59608a <=( (not A166)  and  a59607a );
 a59609a <=( a59608a  and  a59603a );
 a59613a <=( A265  and  A233 );
 a59614a <=( A232  and  a59613a );
 a59617a <=( (not A299)  and  (not A267) );
 a59620a <=( (not A302)  and  (not A301) );
 a59621a <=( a59620a  and  a59617a );
 a59622a <=( a59621a  and  a59614a );
 a59626a <=( A167  and  (not A169) );
 a59627a <=( A170  and  a59626a );
 a59631a <=( (not A200)  and  (not A199) );
 a59632a <=( (not A166)  and  a59631a );
 a59633a <=( a59632a  and  a59627a );
 a59637a <=( A265  and  A233 );
 a59638a <=( A232  and  a59637a );
 a59641a <=( (not A299)  and  A266 );
 a59644a <=( (not A302)  and  (not A301) );
 a59645a <=( a59644a  and  a59641a );
 a59646a <=( a59645a  and  a59638a );
 a59650a <=( A167  and  (not A169) );
 a59651a <=( A170  and  a59650a );
 a59655a <=( (not A200)  and  (not A199) );
 a59656a <=( (not A166)  and  a59655a );
 a59657a <=( a59656a  and  a59651a );
 a59661a <=( (not A265)  and  A233 );
 a59662a <=( A232  and  a59661a );
 a59665a <=( (not A299)  and  (not A266) );
 a59668a <=( (not A302)  and  (not A301) );
 a59669a <=( a59668a  and  a59665a );
 a59670a <=( a59669a  and  a59662a );
 a59674a <=( A167  and  (not A169) );
 a59675a <=( A170  and  a59674a );
 a59679a <=( (not A200)  and  (not A199) );
 a59680a <=( (not A166)  and  a59679a );
 a59681a <=( a59680a  and  a59675a );
 a59685a <=( (not A236)  and  (not A235) );
 a59686a <=( (not A233)  and  a59685a );
 a59689a <=( A266  and  A265 );
 a59692a <=( (not A300)  and  A298 );
 a59693a <=( a59692a  and  a59689a );
 a59694a <=( a59693a  and  a59686a );
 a59698a <=( A167  and  (not A169) );
 a59699a <=( A170  and  a59698a );
 a59703a <=( (not A200)  and  (not A199) );
 a59704a <=( (not A166)  and  a59703a );
 a59705a <=( a59704a  and  a59699a );
 a59709a <=( (not A236)  and  (not A235) );
 a59710a <=( (not A233)  and  a59709a );
 a59713a <=( A266  and  A265 );
 a59716a <=( A299  and  A298 );
 a59717a <=( a59716a  and  a59713a );
 a59718a <=( a59717a  and  a59710a );
 a59722a <=( A167  and  (not A169) );
 a59723a <=( A170  and  a59722a );
 a59727a <=( (not A200)  and  (not A199) );
 a59728a <=( (not A166)  and  a59727a );
 a59729a <=( a59728a  and  a59723a );
 a59733a <=( (not A236)  and  (not A235) );
 a59734a <=( (not A233)  and  a59733a );
 a59737a <=( A266  and  A265 );
 a59740a <=( (not A299)  and  (not A298) );
 a59741a <=( a59740a  and  a59737a );
 a59742a <=( a59741a  and  a59734a );
 a59746a <=( A167  and  (not A169) );
 a59747a <=( A170  and  a59746a );
 a59751a <=( (not A200)  and  (not A199) );
 a59752a <=( (not A166)  and  a59751a );
 a59753a <=( a59752a  and  a59747a );
 a59757a <=( (not A236)  and  (not A235) );
 a59758a <=( (not A233)  and  a59757a );
 a59761a <=( (not A267)  and  (not A266) );
 a59764a <=( (not A300)  and  A298 );
 a59765a <=( a59764a  and  a59761a );
 a59766a <=( a59765a  and  a59758a );
 a59770a <=( A167  and  (not A169) );
 a59771a <=( A170  and  a59770a );
 a59775a <=( (not A200)  and  (not A199) );
 a59776a <=( (not A166)  and  a59775a );
 a59777a <=( a59776a  and  a59771a );
 a59781a <=( (not A236)  and  (not A235) );
 a59782a <=( (not A233)  and  a59781a );
 a59785a <=( (not A267)  and  (not A266) );
 a59788a <=( A299  and  A298 );
 a59789a <=( a59788a  and  a59785a );
 a59790a <=( a59789a  and  a59782a );
 a59794a <=( A167  and  (not A169) );
 a59795a <=( A170  and  a59794a );
 a59799a <=( (not A200)  and  (not A199) );
 a59800a <=( (not A166)  and  a59799a );
 a59801a <=( a59800a  and  a59795a );
 a59805a <=( (not A236)  and  (not A235) );
 a59806a <=( (not A233)  and  a59805a );
 a59809a <=( (not A267)  and  (not A266) );
 a59812a <=( (not A299)  and  (not A298) );
 a59813a <=( a59812a  and  a59809a );
 a59814a <=( a59813a  and  a59806a );
 a59818a <=( A167  and  (not A169) );
 a59819a <=( A170  and  a59818a );
 a59823a <=( (not A200)  and  (not A199) );
 a59824a <=( (not A166)  and  a59823a );
 a59825a <=( a59824a  and  a59819a );
 a59829a <=( (not A236)  and  (not A235) );
 a59830a <=( (not A233)  and  a59829a );
 a59833a <=( (not A266)  and  (not A265) );
 a59836a <=( (not A300)  and  A298 );
 a59837a <=( a59836a  and  a59833a );
 a59838a <=( a59837a  and  a59830a );
 a59842a <=( A167  and  (not A169) );
 a59843a <=( A170  and  a59842a );
 a59847a <=( (not A200)  and  (not A199) );
 a59848a <=( (not A166)  and  a59847a );
 a59849a <=( a59848a  and  a59843a );
 a59853a <=( (not A236)  and  (not A235) );
 a59854a <=( (not A233)  and  a59853a );
 a59857a <=( (not A266)  and  (not A265) );
 a59860a <=( A299  and  A298 );
 a59861a <=( a59860a  and  a59857a );
 a59862a <=( a59861a  and  a59854a );
 a59866a <=( A167  and  (not A169) );
 a59867a <=( A170  and  a59866a );
 a59871a <=( (not A200)  and  (not A199) );
 a59872a <=( (not A166)  and  a59871a );
 a59873a <=( a59872a  and  a59867a );
 a59877a <=( (not A236)  and  (not A235) );
 a59878a <=( (not A233)  and  a59877a );
 a59881a <=( (not A266)  and  (not A265) );
 a59884a <=( (not A299)  and  (not A298) );
 a59885a <=( a59884a  and  a59881a );
 a59886a <=( a59885a  and  a59878a );
 a59890a <=( A167  and  (not A169) );
 a59891a <=( A170  and  a59890a );
 a59895a <=( (not A200)  and  (not A199) );
 a59896a <=( (not A166)  and  a59895a );
 a59897a <=( a59896a  and  a59891a );
 a59901a <=( A265  and  (not A234) );
 a59902a <=( (not A233)  and  a59901a );
 a59905a <=( A298  and  A266 );
 a59908a <=( (not A302)  and  (not A301) );
 a59909a <=( a59908a  and  a59905a );
 a59910a <=( a59909a  and  a59902a );
 a59914a <=( A167  and  (not A169) );
 a59915a <=( A170  and  a59914a );
 a59919a <=( (not A200)  and  (not A199) );
 a59920a <=( (not A166)  and  a59919a );
 a59921a <=( a59920a  and  a59915a );
 a59925a <=( (not A266)  and  (not A234) );
 a59926a <=( (not A233)  and  a59925a );
 a59929a <=( (not A269)  and  (not A268) );
 a59932a <=( (not A300)  and  A298 );
 a59933a <=( a59932a  and  a59929a );
 a59934a <=( a59933a  and  a59926a );
 a59938a <=( A167  and  (not A169) );
 a59939a <=( A170  and  a59938a );
 a59943a <=( (not A200)  and  (not A199) );
 a59944a <=( (not A166)  and  a59943a );
 a59945a <=( a59944a  and  a59939a );
 a59949a <=( (not A266)  and  (not A234) );
 a59950a <=( (not A233)  and  a59949a );
 a59953a <=( (not A269)  and  (not A268) );
 a59956a <=( A299  and  A298 );
 a59957a <=( a59956a  and  a59953a );
 a59958a <=( a59957a  and  a59950a );
 a59962a <=( A167  and  (not A169) );
 a59963a <=( A170  and  a59962a );
 a59967a <=( (not A200)  and  (not A199) );
 a59968a <=( (not A166)  and  a59967a );
 a59969a <=( a59968a  and  a59963a );
 a59973a <=( (not A266)  and  (not A234) );
 a59974a <=( (not A233)  and  a59973a );
 a59977a <=( (not A269)  and  (not A268) );
 a59980a <=( (not A299)  and  (not A298) );
 a59981a <=( a59980a  and  a59977a );
 a59982a <=( a59981a  and  a59974a );
 a59986a <=( A167  and  (not A169) );
 a59987a <=( A170  and  a59986a );
 a59991a <=( (not A200)  and  (not A199) );
 a59992a <=( (not A166)  and  a59991a );
 a59993a <=( a59992a  and  a59987a );
 a59997a <=( (not A266)  and  (not A234) );
 a59998a <=( (not A233)  and  a59997a );
 a60001a <=( A298  and  (not A267) );
 a60004a <=( (not A302)  and  (not A301) );
 a60005a <=( a60004a  and  a60001a );
 a60006a <=( a60005a  and  a59998a );
 a60010a <=( A167  and  (not A169) );
 a60011a <=( A170  and  a60010a );
 a60015a <=( (not A200)  and  (not A199) );
 a60016a <=( (not A166)  and  a60015a );
 a60017a <=( a60016a  and  a60011a );
 a60021a <=( (not A265)  and  (not A234) );
 a60022a <=( (not A233)  and  a60021a );
 a60025a <=( A298  and  (not A266) );
 a60028a <=( (not A302)  and  (not A301) );
 a60029a <=( a60028a  and  a60025a );
 a60030a <=( a60029a  and  a60022a );
 a60034a <=( A167  and  (not A169) );
 a60035a <=( A170  and  a60034a );
 a60039a <=( (not A200)  and  (not A199) );
 a60040a <=( (not A166)  and  a60039a );
 a60041a <=( a60040a  and  a60035a );
 a60045a <=( A265  and  (not A233) );
 a60046a <=( (not A232)  and  a60045a );
 a60049a <=( A298  and  A266 );
 a60052a <=( (not A302)  and  (not A301) );
 a60053a <=( a60052a  and  a60049a );
 a60054a <=( a60053a  and  a60046a );
 a60058a <=( A167  and  (not A169) );
 a60059a <=( A170  and  a60058a );
 a60063a <=( (not A200)  and  (not A199) );
 a60064a <=( (not A166)  and  a60063a );
 a60065a <=( a60064a  and  a60059a );
 a60069a <=( (not A266)  and  (not A233) );
 a60070a <=( (not A232)  and  a60069a );
 a60073a <=( (not A269)  and  (not A268) );
 a60076a <=( (not A300)  and  A298 );
 a60077a <=( a60076a  and  a60073a );
 a60078a <=( a60077a  and  a60070a );
 a60082a <=( A167  and  (not A169) );
 a60083a <=( A170  and  a60082a );
 a60087a <=( (not A200)  and  (not A199) );
 a60088a <=( (not A166)  and  a60087a );
 a60089a <=( a60088a  and  a60083a );
 a60093a <=( (not A266)  and  (not A233) );
 a60094a <=( (not A232)  and  a60093a );
 a60097a <=( (not A269)  and  (not A268) );
 a60100a <=( A299  and  A298 );
 a60101a <=( a60100a  and  a60097a );
 a60102a <=( a60101a  and  a60094a );
 a60106a <=( A167  and  (not A169) );
 a60107a <=( A170  and  a60106a );
 a60111a <=( (not A200)  and  (not A199) );
 a60112a <=( (not A166)  and  a60111a );
 a60113a <=( a60112a  and  a60107a );
 a60117a <=( (not A266)  and  (not A233) );
 a60118a <=( (not A232)  and  a60117a );
 a60121a <=( (not A269)  and  (not A268) );
 a60124a <=( (not A299)  and  (not A298) );
 a60125a <=( a60124a  and  a60121a );
 a60126a <=( a60125a  and  a60118a );
 a60130a <=( A167  and  (not A169) );
 a60131a <=( A170  and  a60130a );
 a60135a <=( (not A200)  and  (not A199) );
 a60136a <=( (not A166)  and  a60135a );
 a60137a <=( a60136a  and  a60131a );
 a60141a <=( (not A266)  and  (not A233) );
 a60142a <=( (not A232)  and  a60141a );
 a60145a <=( A298  and  (not A267) );
 a60148a <=( (not A302)  and  (not A301) );
 a60149a <=( a60148a  and  a60145a );
 a60150a <=( a60149a  and  a60142a );
 a60154a <=( A167  and  (not A169) );
 a60155a <=( A170  and  a60154a );
 a60159a <=( (not A200)  and  (not A199) );
 a60160a <=( (not A166)  and  a60159a );
 a60161a <=( a60160a  and  a60155a );
 a60165a <=( (not A265)  and  (not A233) );
 a60166a <=( (not A232)  and  a60165a );
 a60169a <=( A298  and  (not A266) );
 a60172a <=( (not A302)  and  (not A301) );
 a60173a <=( a60172a  and  a60169a );
 a60174a <=( a60173a  and  a60166a );
 a60178a <=( (not A167)  and  (not A169) );
 a60179a <=( A170  and  a60178a );
 a60183a <=( A200  and  A199 );
 a60184a <=( A166  and  a60183a );
 a60185a <=( a60184a  and  a60179a );
 a60189a <=( A265  and  A233 );
 a60190a <=( A232  and  a60189a );
 a60193a <=( (not A269)  and  (not A268) );
 a60196a <=( (not A300)  and  (not A299) );
 a60197a <=( a60196a  and  a60193a );
 a60198a <=( a60197a  and  a60190a );
 a60202a <=( (not A167)  and  (not A169) );
 a60203a <=( A170  and  a60202a );
 a60207a <=( A200  and  A199 );
 a60208a <=( A166  and  a60207a );
 a60209a <=( a60208a  and  a60203a );
 a60213a <=( A265  and  A233 );
 a60214a <=( A232  and  a60213a );
 a60217a <=( (not A269)  and  (not A268) );
 a60220a <=( A299  and  A298 );
 a60221a <=( a60220a  and  a60217a );
 a60222a <=( a60221a  and  a60214a );
 a60226a <=( (not A167)  and  (not A169) );
 a60227a <=( A170  and  a60226a );
 a60231a <=( A200  and  A199 );
 a60232a <=( A166  and  a60231a );
 a60233a <=( a60232a  and  a60227a );
 a60237a <=( A265  and  A233 );
 a60238a <=( A232  and  a60237a );
 a60241a <=( (not A269)  and  (not A268) );
 a60244a <=( (not A299)  and  (not A298) );
 a60245a <=( a60244a  and  a60241a );
 a60246a <=( a60245a  and  a60238a );
 a60250a <=( (not A167)  and  (not A169) );
 a60251a <=( A170  and  a60250a );
 a60255a <=( A200  and  A199 );
 a60256a <=( A166  and  a60255a );
 a60257a <=( a60256a  and  a60251a );
 a60261a <=( A265  and  A233 );
 a60262a <=( A232  and  a60261a );
 a60265a <=( (not A299)  and  (not A267) );
 a60268a <=( (not A302)  and  (not A301) );
 a60269a <=( a60268a  and  a60265a );
 a60270a <=( a60269a  and  a60262a );
 a60274a <=( (not A167)  and  (not A169) );
 a60275a <=( A170  and  a60274a );
 a60279a <=( A200  and  A199 );
 a60280a <=( A166  and  a60279a );
 a60281a <=( a60280a  and  a60275a );
 a60285a <=( A265  and  A233 );
 a60286a <=( A232  and  a60285a );
 a60289a <=( (not A299)  and  A266 );
 a60292a <=( (not A302)  and  (not A301) );
 a60293a <=( a60292a  and  a60289a );
 a60294a <=( a60293a  and  a60286a );
 a60298a <=( (not A167)  and  (not A169) );
 a60299a <=( A170  and  a60298a );
 a60303a <=( A200  and  A199 );
 a60304a <=( A166  and  a60303a );
 a60305a <=( a60304a  and  a60299a );
 a60309a <=( (not A265)  and  A233 );
 a60310a <=( A232  and  a60309a );
 a60313a <=( (not A299)  and  (not A266) );
 a60316a <=( (not A302)  and  (not A301) );
 a60317a <=( a60316a  and  a60313a );
 a60318a <=( a60317a  and  a60310a );
 a60322a <=( (not A167)  and  (not A169) );
 a60323a <=( A170  and  a60322a );
 a60327a <=( A200  and  A199 );
 a60328a <=( A166  and  a60327a );
 a60329a <=( a60328a  and  a60323a );
 a60333a <=( (not A236)  and  (not A235) );
 a60334a <=( (not A233)  and  a60333a );
 a60337a <=( A266  and  A265 );
 a60340a <=( (not A300)  and  A298 );
 a60341a <=( a60340a  and  a60337a );
 a60342a <=( a60341a  and  a60334a );
 a60346a <=( (not A167)  and  (not A169) );
 a60347a <=( A170  and  a60346a );
 a60351a <=( A200  and  A199 );
 a60352a <=( A166  and  a60351a );
 a60353a <=( a60352a  and  a60347a );
 a60357a <=( (not A236)  and  (not A235) );
 a60358a <=( (not A233)  and  a60357a );
 a60361a <=( A266  and  A265 );
 a60364a <=( A299  and  A298 );
 a60365a <=( a60364a  and  a60361a );
 a60366a <=( a60365a  and  a60358a );
 a60370a <=( (not A167)  and  (not A169) );
 a60371a <=( A170  and  a60370a );
 a60375a <=( A200  and  A199 );
 a60376a <=( A166  and  a60375a );
 a60377a <=( a60376a  and  a60371a );
 a60381a <=( (not A236)  and  (not A235) );
 a60382a <=( (not A233)  and  a60381a );
 a60385a <=( A266  and  A265 );
 a60388a <=( (not A299)  and  (not A298) );
 a60389a <=( a60388a  and  a60385a );
 a60390a <=( a60389a  and  a60382a );
 a60394a <=( (not A167)  and  (not A169) );
 a60395a <=( A170  and  a60394a );
 a60399a <=( A200  and  A199 );
 a60400a <=( A166  and  a60399a );
 a60401a <=( a60400a  and  a60395a );
 a60405a <=( (not A236)  and  (not A235) );
 a60406a <=( (not A233)  and  a60405a );
 a60409a <=( (not A267)  and  (not A266) );
 a60412a <=( (not A300)  and  A298 );
 a60413a <=( a60412a  and  a60409a );
 a60414a <=( a60413a  and  a60406a );
 a60418a <=( (not A167)  and  (not A169) );
 a60419a <=( A170  and  a60418a );
 a60423a <=( A200  and  A199 );
 a60424a <=( A166  and  a60423a );
 a60425a <=( a60424a  and  a60419a );
 a60429a <=( (not A236)  and  (not A235) );
 a60430a <=( (not A233)  and  a60429a );
 a60433a <=( (not A267)  and  (not A266) );
 a60436a <=( A299  and  A298 );
 a60437a <=( a60436a  and  a60433a );
 a60438a <=( a60437a  and  a60430a );
 a60442a <=( (not A167)  and  (not A169) );
 a60443a <=( A170  and  a60442a );
 a60447a <=( A200  and  A199 );
 a60448a <=( A166  and  a60447a );
 a60449a <=( a60448a  and  a60443a );
 a60453a <=( (not A236)  and  (not A235) );
 a60454a <=( (not A233)  and  a60453a );
 a60457a <=( (not A267)  and  (not A266) );
 a60460a <=( (not A299)  and  (not A298) );
 a60461a <=( a60460a  and  a60457a );
 a60462a <=( a60461a  and  a60454a );
 a60466a <=( (not A167)  and  (not A169) );
 a60467a <=( A170  and  a60466a );
 a60471a <=( A200  and  A199 );
 a60472a <=( A166  and  a60471a );
 a60473a <=( a60472a  and  a60467a );
 a60477a <=( (not A236)  and  (not A235) );
 a60478a <=( (not A233)  and  a60477a );
 a60481a <=( (not A266)  and  (not A265) );
 a60484a <=( (not A300)  and  A298 );
 a60485a <=( a60484a  and  a60481a );
 a60486a <=( a60485a  and  a60478a );
 a60490a <=( (not A167)  and  (not A169) );
 a60491a <=( A170  and  a60490a );
 a60495a <=( A200  and  A199 );
 a60496a <=( A166  and  a60495a );
 a60497a <=( a60496a  and  a60491a );
 a60501a <=( (not A236)  and  (not A235) );
 a60502a <=( (not A233)  and  a60501a );
 a60505a <=( (not A266)  and  (not A265) );
 a60508a <=( A299  and  A298 );
 a60509a <=( a60508a  and  a60505a );
 a60510a <=( a60509a  and  a60502a );
 a60514a <=( (not A167)  and  (not A169) );
 a60515a <=( A170  and  a60514a );
 a60519a <=( A200  and  A199 );
 a60520a <=( A166  and  a60519a );
 a60521a <=( a60520a  and  a60515a );
 a60525a <=( (not A236)  and  (not A235) );
 a60526a <=( (not A233)  and  a60525a );
 a60529a <=( (not A266)  and  (not A265) );
 a60532a <=( (not A299)  and  (not A298) );
 a60533a <=( a60532a  and  a60529a );
 a60534a <=( a60533a  and  a60526a );
 a60538a <=( (not A167)  and  (not A169) );
 a60539a <=( A170  and  a60538a );
 a60543a <=( A200  and  A199 );
 a60544a <=( A166  and  a60543a );
 a60545a <=( a60544a  and  a60539a );
 a60549a <=( A265  and  (not A234) );
 a60550a <=( (not A233)  and  a60549a );
 a60553a <=( A298  and  A266 );
 a60556a <=( (not A302)  and  (not A301) );
 a60557a <=( a60556a  and  a60553a );
 a60558a <=( a60557a  and  a60550a );
 a60562a <=( (not A167)  and  (not A169) );
 a60563a <=( A170  and  a60562a );
 a60567a <=( A200  and  A199 );
 a60568a <=( A166  and  a60567a );
 a60569a <=( a60568a  and  a60563a );
 a60573a <=( (not A266)  and  (not A234) );
 a60574a <=( (not A233)  and  a60573a );
 a60577a <=( (not A269)  and  (not A268) );
 a60580a <=( (not A300)  and  A298 );
 a60581a <=( a60580a  and  a60577a );
 a60582a <=( a60581a  and  a60574a );
 a60586a <=( (not A167)  and  (not A169) );
 a60587a <=( A170  and  a60586a );
 a60591a <=( A200  and  A199 );
 a60592a <=( A166  and  a60591a );
 a60593a <=( a60592a  and  a60587a );
 a60597a <=( (not A266)  and  (not A234) );
 a60598a <=( (not A233)  and  a60597a );
 a60601a <=( (not A269)  and  (not A268) );
 a60604a <=( A299  and  A298 );
 a60605a <=( a60604a  and  a60601a );
 a60606a <=( a60605a  and  a60598a );
 a60610a <=( (not A167)  and  (not A169) );
 a60611a <=( A170  and  a60610a );
 a60615a <=( A200  and  A199 );
 a60616a <=( A166  and  a60615a );
 a60617a <=( a60616a  and  a60611a );
 a60621a <=( (not A266)  and  (not A234) );
 a60622a <=( (not A233)  and  a60621a );
 a60625a <=( (not A269)  and  (not A268) );
 a60628a <=( (not A299)  and  (not A298) );
 a60629a <=( a60628a  and  a60625a );
 a60630a <=( a60629a  and  a60622a );
 a60634a <=( (not A167)  and  (not A169) );
 a60635a <=( A170  and  a60634a );
 a60639a <=( A200  and  A199 );
 a60640a <=( A166  and  a60639a );
 a60641a <=( a60640a  and  a60635a );
 a60645a <=( (not A266)  and  (not A234) );
 a60646a <=( (not A233)  and  a60645a );
 a60649a <=( A298  and  (not A267) );
 a60652a <=( (not A302)  and  (not A301) );
 a60653a <=( a60652a  and  a60649a );
 a60654a <=( a60653a  and  a60646a );
 a60658a <=( (not A167)  and  (not A169) );
 a60659a <=( A170  and  a60658a );
 a60663a <=( A200  and  A199 );
 a60664a <=( A166  and  a60663a );
 a60665a <=( a60664a  and  a60659a );
 a60669a <=( (not A265)  and  (not A234) );
 a60670a <=( (not A233)  and  a60669a );
 a60673a <=( A298  and  (not A266) );
 a60676a <=( (not A302)  and  (not A301) );
 a60677a <=( a60676a  and  a60673a );
 a60678a <=( a60677a  and  a60670a );
 a60682a <=( (not A167)  and  (not A169) );
 a60683a <=( A170  and  a60682a );
 a60687a <=( A200  and  A199 );
 a60688a <=( A166  and  a60687a );
 a60689a <=( a60688a  and  a60683a );
 a60693a <=( A265  and  (not A233) );
 a60694a <=( (not A232)  and  a60693a );
 a60697a <=( A298  and  A266 );
 a60700a <=( (not A302)  and  (not A301) );
 a60701a <=( a60700a  and  a60697a );
 a60702a <=( a60701a  and  a60694a );
 a60706a <=( (not A167)  and  (not A169) );
 a60707a <=( A170  and  a60706a );
 a60711a <=( A200  and  A199 );
 a60712a <=( A166  and  a60711a );
 a60713a <=( a60712a  and  a60707a );
 a60717a <=( (not A266)  and  (not A233) );
 a60718a <=( (not A232)  and  a60717a );
 a60721a <=( (not A269)  and  (not A268) );
 a60724a <=( (not A300)  and  A298 );
 a60725a <=( a60724a  and  a60721a );
 a60726a <=( a60725a  and  a60718a );
 a60730a <=( (not A167)  and  (not A169) );
 a60731a <=( A170  and  a60730a );
 a60735a <=( A200  and  A199 );
 a60736a <=( A166  and  a60735a );
 a60737a <=( a60736a  and  a60731a );
 a60741a <=( (not A266)  and  (not A233) );
 a60742a <=( (not A232)  and  a60741a );
 a60745a <=( (not A269)  and  (not A268) );
 a60748a <=( A299  and  A298 );
 a60749a <=( a60748a  and  a60745a );
 a60750a <=( a60749a  and  a60742a );
 a60754a <=( (not A167)  and  (not A169) );
 a60755a <=( A170  and  a60754a );
 a60759a <=( A200  and  A199 );
 a60760a <=( A166  and  a60759a );
 a60761a <=( a60760a  and  a60755a );
 a60765a <=( (not A266)  and  (not A233) );
 a60766a <=( (not A232)  and  a60765a );
 a60769a <=( (not A269)  and  (not A268) );
 a60772a <=( (not A299)  and  (not A298) );
 a60773a <=( a60772a  and  a60769a );
 a60774a <=( a60773a  and  a60766a );
 a60778a <=( (not A167)  and  (not A169) );
 a60779a <=( A170  and  a60778a );
 a60783a <=( A200  and  A199 );
 a60784a <=( A166  and  a60783a );
 a60785a <=( a60784a  and  a60779a );
 a60789a <=( (not A266)  and  (not A233) );
 a60790a <=( (not A232)  and  a60789a );
 a60793a <=( A298  and  (not A267) );
 a60796a <=( (not A302)  and  (not A301) );
 a60797a <=( a60796a  and  a60793a );
 a60798a <=( a60797a  and  a60790a );
 a60802a <=( (not A167)  and  (not A169) );
 a60803a <=( A170  and  a60802a );
 a60807a <=( A200  and  A199 );
 a60808a <=( A166  and  a60807a );
 a60809a <=( a60808a  and  a60803a );
 a60813a <=( (not A265)  and  (not A233) );
 a60814a <=( (not A232)  and  a60813a );
 a60817a <=( A298  and  (not A266) );
 a60820a <=( (not A302)  and  (not A301) );
 a60821a <=( a60820a  and  a60817a );
 a60822a <=( a60821a  and  a60814a );
 a60826a <=( (not A167)  and  (not A169) );
 a60827a <=( A170  and  a60826a );
 a60831a <=( (not A202)  and  (not A200) );
 a60832a <=( A166  and  a60831a );
 a60833a <=( a60832a  and  a60827a );
 a60837a <=( A233  and  A232 );
 a60838a <=( (not A203)  and  a60837a );
 a60841a <=( (not A267)  and  A265 );
 a60844a <=( (not A300)  and  (not A299) );
 a60845a <=( a60844a  and  a60841a );
 a60846a <=( a60845a  and  a60838a );
 a60850a <=( (not A167)  and  (not A169) );
 a60851a <=( A170  and  a60850a );
 a60855a <=( (not A202)  and  (not A200) );
 a60856a <=( A166  and  a60855a );
 a60857a <=( a60856a  and  a60851a );
 a60861a <=( A233  and  A232 );
 a60862a <=( (not A203)  and  a60861a );
 a60865a <=( (not A267)  and  A265 );
 a60868a <=( A299  and  A298 );
 a60869a <=( a60868a  and  a60865a );
 a60870a <=( a60869a  and  a60862a );
 a60874a <=( (not A167)  and  (not A169) );
 a60875a <=( A170  and  a60874a );
 a60879a <=( (not A202)  and  (not A200) );
 a60880a <=( A166  and  a60879a );
 a60881a <=( a60880a  and  a60875a );
 a60885a <=( A233  and  A232 );
 a60886a <=( (not A203)  and  a60885a );
 a60889a <=( (not A267)  and  A265 );
 a60892a <=( (not A299)  and  (not A298) );
 a60893a <=( a60892a  and  a60889a );
 a60894a <=( a60893a  and  a60886a );
 a60898a <=( (not A167)  and  (not A169) );
 a60899a <=( A170  and  a60898a );
 a60903a <=( (not A202)  and  (not A200) );
 a60904a <=( A166  and  a60903a );
 a60905a <=( a60904a  and  a60899a );
 a60909a <=( A233  and  A232 );
 a60910a <=( (not A203)  and  a60909a );
 a60913a <=( A266  and  A265 );
 a60916a <=( (not A300)  and  (not A299) );
 a60917a <=( a60916a  and  a60913a );
 a60918a <=( a60917a  and  a60910a );
 a60922a <=( (not A167)  and  (not A169) );
 a60923a <=( A170  and  a60922a );
 a60927a <=( (not A202)  and  (not A200) );
 a60928a <=( A166  and  a60927a );
 a60929a <=( a60928a  and  a60923a );
 a60933a <=( A233  and  A232 );
 a60934a <=( (not A203)  and  a60933a );
 a60937a <=( A266  and  A265 );
 a60940a <=( A299  and  A298 );
 a60941a <=( a60940a  and  a60937a );
 a60942a <=( a60941a  and  a60934a );
 a60946a <=( (not A167)  and  (not A169) );
 a60947a <=( A170  and  a60946a );
 a60951a <=( (not A202)  and  (not A200) );
 a60952a <=( A166  and  a60951a );
 a60953a <=( a60952a  and  a60947a );
 a60957a <=( A233  and  A232 );
 a60958a <=( (not A203)  and  a60957a );
 a60961a <=( A266  and  A265 );
 a60964a <=( (not A299)  and  (not A298) );
 a60965a <=( a60964a  and  a60961a );
 a60966a <=( a60965a  and  a60958a );
 a60970a <=( (not A167)  and  (not A169) );
 a60971a <=( A170  and  a60970a );
 a60975a <=( (not A202)  and  (not A200) );
 a60976a <=( A166  and  a60975a );
 a60977a <=( a60976a  and  a60971a );
 a60981a <=( A233  and  A232 );
 a60982a <=( (not A203)  and  a60981a );
 a60985a <=( (not A266)  and  (not A265) );
 a60988a <=( (not A300)  and  (not A299) );
 a60989a <=( a60988a  and  a60985a );
 a60990a <=( a60989a  and  a60982a );
 a60994a <=( (not A167)  and  (not A169) );
 a60995a <=( A170  and  a60994a );
 a60999a <=( (not A202)  and  (not A200) );
 a61000a <=( A166  and  a60999a );
 a61001a <=( a61000a  and  a60995a );
 a61005a <=( A233  and  A232 );
 a61006a <=( (not A203)  and  a61005a );
 a61009a <=( (not A266)  and  (not A265) );
 a61012a <=( A299  and  A298 );
 a61013a <=( a61012a  and  a61009a );
 a61014a <=( a61013a  and  a61006a );
 a61018a <=( (not A167)  and  (not A169) );
 a61019a <=( A170  and  a61018a );
 a61023a <=( (not A202)  and  (not A200) );
 a61024a <=( A166  and  a61023a );
 a61025a <=( a61024a  and  a61019a );
 a61029a <=( A233  and  A232 );
 a61030a <=( (not A203)  and  a61029a );
 a61033a <=( (not A266)  and  (not A265) );
 a61036a <=( (not A299)  and  (not A298) );
 a61037a <=( a61036a  and  a61033a );
 a61038a <=( a61037a  and  a61030a );
 a61042a <=( (not A167)  and  (not A169) );
 a61043a <=( A170  and  a61042a );
 a61047a <=( (not A202)  and  (not A200) );
 a61048a <=( A166  and  a61047a );
 a61049a <=( a61048a  and  a61043a );
 a61053a <=( A233  and  (not A232) );
 a61054a <=( (not A203)  and  a61053a );
 a61057a <=( (not A299)  and  A298 );
 a61060a <=( A301  and  A300 );
 a61061a <=( a61060a  and  a61057a );
 a61062a <=( a61061a  and  a61054a );
 a61066a <=( (not A167)  and  (not A169) );
 a61067a <=( A170  and  a61066a );
 a61071a <=( (not A202)  and  (not A200) );
 a61072a <=( A166  and  a61071a );
 a61073a <=( a61072a  and  a61067a );
 a61077a <=( A233  and  (not A232) );
 a61078a <=( (not A203)  and  a61077a );
 a61081a <=( (not A299)  and  A298 );
 a61084a <=( A302  and  A300 );
 a61085a <=( a61084a  and  a61081a );
 a61086a <=( a61085a  and  a61078a );
 a61090a <=( (not A167)  and  (not A169) );
 a61091a <=( A170  and  a61090a );
 a61095a <=( (not A202)  and  (not A200) );
 a61096a <=( A166  and  a61095a );
 a61097a <=( a61096a  and  a61091a );
 a61101a <=( A233  and  (not A232) );
 a61102a <=( (not A203)  and  a61101a );
 a61105a <=( (not A266)  and  A265 );
 a61108a <=( A268  and  A267 );
 a61109a <=( a61108a  and  a61105a );
 a61110a <=( a61109a  and  a61102a );
 a61114a <=( (not A167)  and  (not A169) );
 a61115a <=( A170  and  a61114a );
 a61119a <=( (not A202)  and  (not A200) );
 a61120a <=( A166  and  a61119a );
 a61121a <=( a61120a  and  a61115a );
 a61125a <=( A233  and  (not A232) );
 a61126a <=( (not A203)  and  a61125a );
 a61129a <=( (not A266)  and  A265 );
 a61132a <=( A269  and  A267 );
 a61133a <=( a61132a  and  a61129a );
 a61134a <=( a61133a  and  a61126a );
 a61138a <=( (not A167)  and  (not A169) );
 a61139a <=( A170  and  a61138a );
 a61143a <=( (not A202)  and  (not A200) );
 a61144a <=( A166  and  a61143a );
 a61145a <=( a61144a  and  a61139a );
 a61149a <=( (not A234)  and  (not A233) );
 a61150a <=( (not A203)  and  a61149a );
 a61153a <=( A266  and  A265 );
 a61156a <=( (not A300)  and  A298 );
 a61157a <=( a61156a  and  a61153a );
 a61158a <=( a61157a  and  a61150a );
 a61162a <=( (not A167)  and  (not A169) );
 a61163a <=( A170  and  a61162a );
 a61167a <=( (not A202)  and  (not A200) );
 a61168a <=( A166  and  a61167a );
 a61169a <=( a61168a  and  a61163a );
 a61173a <=( (not A234)  and  (not A233) );
 a61174a <=( (not A203)  and  a61173a );
 a61177a <=( A266  and  A265 );
 a61180a <=( A299  and  A298 );
 a61181a <=( a61180a  and  a61177a );
 a61182a <=( a61181a  and  a61174a );
 a61186a <=( (not A167)  and  (not A169) );
 a61187a <=( A170  and  a61186a );
 a61191a <=( (not A202)  and  (not A200) );
 a61192a <=( A166  and  a61191a );
 a61193a <=( a61192a  and  a61187a );
 a61197a <=( (not A234)  and  (not A233) );
 a61198a <=( (not A203)  and  a61197a );
 a61201a <=( A266  and  A265 );
 a61204a <=( (not A299)  and  (not A298) );
 a61205a <=( a61204a  and  a61201a );
 a61206a <=( a61205a  and  a61198a );
 a61210a <=( (not A167)  and  (not A169) );
 a61211a <=( A170  and  a61210a );
 a61215a <=( (not A202)  and  (not A200) );
 a61216a <=( A166  and  a61215a );
 a61217a <=( a61216a  and  a61211a );
 a61221a <=( (not A234)  and  (not A233) );
 a61222a <=( (not A203)  and  a61221a );
 a61225a <=( (not A267)  and  (not A266) );
 a61228a <=( (not A300)  and  A298 );
 a61229a <=( a61228a  and  a61225a );
 a61230a <=( a61229a  and  a61222a );
 a61234a <=( (not A167)  and  (not A169) );
 a61235a <=( A170  and  a61234a );
 a61239a <=( (not A202)  and  (not A200) );
 a61240a <=( A166  and  a61239a );
 a61241a <=( a61240a  and  a61235a );
 a61245a <=( (not A234)  and  (not A233) );
 a61246a <=( (not A203)  and  a61245a );
 a61249a <=( (not A267)  and  (not A266) );
 a61252a <=( A299  and  A298 );
 a61253a <=( a61252a  and  a61249a );
 a61254a <=( a61253a  and  a61246a );
 a61258a <=( (not A167)  and  (not A169) );
 a61259a <=( A170  and  a61258a );
 a61263a <=( (not A202)  and  (not A200) );
 a61264a <=( A166  and  a61263a );
 a61265a <=( a61264a  and  a61259a );
 a61269a <=( (not A234)  and  (not A233) );
 a61270a <=( (not A203)  and  a61269a );
 a61273a <=( (not A267)  and  (not A266) );
 a61276a <=( (not A299)  and  (not A298) );
 a61277a <=( a61276a  and  a61273a );
 a61278a <=( a61277a  and  a61270a );
 a61282a <=( (not A167)  and  (not A169) );
 a61283a <=( A170  and  a61282a );
 a61287a <=( (not A202)  and  (not A200) );
 a61288a <=( A166  and  a61287a );
 a61289a <=( a61288a  and  a61283a );
 a61293a <=( (not A234)  and  (not A233) );
 a61294a <=( (not A203)  and  a61293a );
 a61297a <=( (not A266)  and  (not A265) );
 a61300a <=( (not A300)  and  A298 );
 a61301a <=( a61300a  and  a61297a );
 a61302a <=( a61301a  and  a61294a );
 a61306a <=( (not A167)  and  (not A169) );
 a61307a <=( A170  and  a61306a );
 a61311a <=( (not A202)  and  (not A200) );
 a61312a <=( A166  and  a61311a );
 a61313a <=( a61312a  and  a61307a );
 a61317a <=( (not A234)  and  (not A233) );
 a61318a <=( (not A203)  and  a61317a );
 a61321a <=( (not A266)  and  (not A265) );
 a61324a <=( A299  and  A298 );
 a61325a <=( a61324a  and  a61321a );
 a61326a <=( a61325a  and  a61318a );
 a61330a <=( (not A167)  and  (not A169) );
 a61331a <=( A170  and  a61330a );
 a61335a <=( (not A202)  and  (not A200) );
 a61336a <=( A166  and  a61335a );
 a61337a <=( a61336a  and  a61331a );
 a61341a <=( (not A234)  and  (not A233) );
 a61342a <=( (not A203)  and  a61341a );
 a61345a <=( (not A266)  and  (not A265) );
 a61348a <=( (not A299)  and  (not A298) );
 a61349a <=( a61348a  and  a61345a );
 a61350a <=( a61349a  and  a61342a );
 a61354a <=( (not A167)  and  (not A169) );
 a61355a <=( A170  and  a61354a );
 a61359a <=( (not A202)  and  (not A200) );
 a61360a <=( A166  and  a61359a );
 a61361a <=( a61360a  and  a61355a );
 a61365a <=( (not A233)  and  A232 );
 a61366a <=( (not A203)  and  a61365a );
 a61369a <=( A235  and  A234 );
 a61372a <=( A299  and  (not A298) );
 a61373a <=( a61372a  and  a61369a );
 a61374a <=( a61373a  and  a61366a );
 a61378a <=( (not A167)  and  (not A169) );
 a61379a <=( A170  and  a61378a );
 a61383a <=( (not A202)  and  (not A200) );
 a61384a <=( A166  and  a61383a );
 a61385a <=( a61384a  and  a61379a );
 a61389a <=( (not A233)  and  A232 );
 a61390a <=( (not A203)  and  a61389a );
 a61393a <=( A235  and  A234 );
 a61396a <=( A266  and  (not A265) );
 a61397a <=( a61396a  and  a61393a );
 a61398a <=( a61397a  and  a61390a );
 a61402a <=( (not A167)  and  (not A169) );
 a61403a <=( A170  and  a61402a );
 a61407a <=( (not A202)  and  (not A200) );
 a61408a <=( A166  and  a61407a );
 a61409a <=( a61408a  and  a61403a );
 a61413a <=( (not A233)  and  A232 );
 a61414a <=( (not A203)  and  a61413a );
 a61417a <=( A236  and  A234 );
 a61420a <=( A299  and  (not A298) );
 a61421a <=( a61420a  and  a61417a );
 a61422a <=( a61421a  and  a61414a );
 a61426a <=( (not A167)  and  (not A169) );
 a61427a <=( A170  and  a61426a );
 a61431a <=( (not A202)  and  (not A200) );
 a61432a <=( A166  and  a61431a );
 a61433a <=( a61432a  and  a61427a );
 a61437a <=( (not A233)  and  A232 );
 a61438a <=( (not A203)  and  a61437a );
 a61441a <=( A236  and  A234 );
 a61444a <=( A266  and  (not A265) );
 a61445a <=( a61444a  and  a61441a );
 a61446a <=( a61445a  and  a61438a );
 a61450a <=( (not A167)  and  (not A169) );
 a61451a <=( A170  and  a61450a );
 a61455a <=( (not A202)  and  (not A200) );
 a61456a <=( A166  and  a61455a );
 a61457a <=( a61456a  and  a61451a );
 a61461a <=( (not A233)  and  (not A232) );
 a61462a <=( (not A203)  and  a61461a );
 a61465a <=( A266  and  A265 );
 a61468a <=( (not A300)  and  A298 );
 a61469a <=( a61468a  and  a61465a );
 a61470a <=( a61469a  and  a61462a );
 a61474a <=( (not A167)  and  (not A169) );
 a61475a <=( A170  and  a61474a );
 a61479a <=( (not A202)  and  (not A200) );
 a61480a <=( A166  and  a61479a );
 a61481a <=( a61480a  and  a61475a );
 a61485a <=( (not A233)  and  (not A232) );
 a61486a <=( (not A203)  and  a61485a );
 a61489a <=( A266  and  A265 );
 a61492a <=( A299  and  A298 );
 a61493a <=( a61492a  and  a61489a );
 a61494a <=( a61493a  and  a61486a );
 a61498a <=( (not A167)  and  (not A169) );
 a61499a <=( A170  and  a61498a );
 a61503a <=( (not A202)  and  (not A200) );
 a61504a <=( A166  and  a61503a );
 a61505a <=( a61504a  and  a61499a );
 a61509a <=( (not A233)  and  (not A232) );
 a61510a <=( (not A203)  and  a61509a );
 a61513a <=( A266  and  A265 );
 a61516a <=( (not A299)  and  (not A298) );
 a61517a <=( a61516a  and  a61513a );
 a61518a <=( a61517a  and  a61510a );
 a61522a <=( (not A167)  and  (not A169) );
 a61523a <=( A170  and  a61522a );
 a61527a <=( (not A202)  and  (not A200) );
 a61528a <=( A166  and  a61527a );
 a61529a <=( a61528a  and  a61523a );
 a61533a <=( (not A233)  and  (not A232) );
 a61534a <=( (not A203)  and  a61533a );
 a61537a <=( (not A267)  and  (not A266) );
 a61540a <=( (not A300)  and  A298 );
 a61541a <=( a61540a  and  a61537a );
 a61542a <=( a61541a  and  a61534a );
 a61546a <=( (not A167)  and  (not A169) );
 a61547a <=( A170  and  a61546a );
 a61551a <=( (not A202)  and  (not A200) );
 a61552a <=( A166  and  a61551a );
 a61553a <=( a61552a  and  a61547a );
 a61557a <=( (not A233)  and  (not A232) );
 a61558a <=( (not A203)  and  a61557a );
 a61561a <=( (not A267)  and  (not A266) );
 a61564a <=( A299  and  A298 );
 a61565a <=( a61564a  and  a61561a );
 a61566a <=( a61565a  and  a61558a );
 a61570a <=( (not A167)  and  (not A169) );
 a61571a <=( A170  and  a61570a );
 a61575a <=( (not A202)  and  (not A200) );
 a61576a <=( A166  and  a61575a );
 a61577a <=( a61576a  and  a61571a );
 a61581a <=( (not A233)  and  (not A232) );
 a61582a <=( (not A203)  and  a61581a );
 a61585a <=( (not A267)  and  (not A266) );
 a61588a <=( (not A299)  and  (not A298) );
 a61589a <=( a61588a  and  a61585a );
 a61590a <=( a61589a  and  a61582a );
 a61594a <=( (not A167)  and  (not A169) );
 a61595a <=( A170  and  a61594a );
 a61599a <=( (not A202)  and  (not A200) );
 a61600a <=( A166  and  a61599a );
 a61601a <=( a61600a  and  a61595a );
 a61605a <=( (not A233)  and  (not A232) );
 a61606a <=( (not A203)  and  a61605a );
 a61609a <=( (not A266)  and  (not A265) );
 a61612a <=( (not A300)  and  A298 );
 a61613a <=( a61612a  and  a61609a );
 a61614a <=( a61613a  and  a61606a );
 a61618a <=( (not A167)  and  (not A169) );
 a61619a <=( A170  and  a61618a );
 a61623a <=( (not A202)  and  (not A200) );
 a61624a <=( A166  and  a61623a );
 a61625a <=( a61624a  and  a61619a );
 a61629a <=( (not A233)  and  (not A232) );
 a61630a <=( (not A203)  and  a61629a );
 a61633a <=( (not A266)  and  (not A265) );
 a61636a <=( A299  and  A298 );
 a61637a <=( a61636a  and  a61633a );
 a61638a <=( a61637a  and  a61630a );
 a61642a <=( (not A167)  and  (not A169) );
 a61643a <=( A170  and  a61642a );
 a61647a <=( (not A202)  and  (not A200) );
 a61648a <=( A166  and  a61647a );
 a61649a <=( a61648a  and  a61643a );
 a61653a <=( (not A233)  and  (not A232) );
 a61654a <=( (not A203)  and  a61653a );
 a61657a <=( (not A266)  and  (not A265) );
 a61660a <=( (not A299)  and  (not A298) );
 a61661a <=( a61660a  and  a61657a );
 a61662a <=( a61661a  and  a61654a );
 a61666a <=( (not A167)  and  (not A169) );
 a61667a <=( A170  and  a61666a );
 a61671a <=( (not A201)  and  (not A200) );
 a61672a <=( A166  and  a61671a );
 a61673a <=( a61672a  and  a61667a );
 a61677a <=( A265  and  A233 );
 a61678a <=( A232  and  a61677a );
 a61681a <=( (not A269)  and  (not A268) );
 a61684a <=( (not A300)  and  (not A299) );
 a61685a <=( a61684a  and  a61681a );
 a61686a <=( a61685a  and  a61678a );
 a61690a <=( (not A167)  and  (not A169) );
 a61691a <=( A170  and  a61690a );
 a61695a <=( (not A201)  and  (not A200) );
 a61696a <=( A166  and  a61695a );
 a61697a <=( a61696a  and  a61691a );
 a61701a <=( A265  and  A233 );
 a61702a <=( A232  and  a61701a );
 a61705a <=( (not A269)  and  (not A268) );
 a61708a <=( A299  and  A298 );
 a61709a <=( a61708a  and  a61705a );
 a61710a <=( a61709a  and  a61702a );
 a61714a <=( (not A167)  and  (not A169) );
 a61715a <=( A170  and  a61714a );
 a61719a <=( (not A201)  and  (not A200) );
 a61720a <=( A166  and  a61719a );
 a61721a <=( a61720a  and  a61715a );
 a61725a <=( A265  and  A233 );
 a61726a <=( A232  and  a61725a );
 a61729a <=( (not A269)  and  (not A268) );
 a61732a <=( (not A299)  and  (not A298) );
 a61733a <=( a61732a  and  a61729a );
 a61734a <=( a61733a  and  a61726a );
 a61738a <=( (not A167)  and  (not A169) );
 a61739a <=( A170  and  a61738a );
 a61743a <=( (not A201)  and  (not A200) );
 a61744a <=( A166  and  a61743a );
 a61745a <=( a61744a  and  a61739a );
 a61749a <=( A265  and  A233 );
 a61750a <=( A232  and  a61749a );
 a61753a <=( (not A299)  and  (not A267) );
 a61756a <=( (not A302)  and  (not A301) );
 a61757a <=( a61756a  and  a61753a );
 a61758a <=( a61757a  and  a61750a );
 a61762a <=( (not A167)  and  (not A169) );
 a61763a <=( A170  and  a61762a );
 a61767a <=( (not A201)  and  (not A200) );
 a61768a <=( A166  and  a61767a );
 a61769a <=( a61768a  and  a61763a );
 a61773a <=( A265  and  A233 );
 a61774a <=( A232  and  a61773a );
 a61777a <=( (not A299)  and  A266 );
 a61780a <=( (not A302)  and  (not A301) );
 a61781a <=( a61780a  and  a61777a );
 a61782a <=( a61781a  and  a61774a );
 a61786a <=( (not A167)  and  (not A169) );
 a61787a <=( A170  and  a61786a );
 a61791a <=( (not A201)  and  (not A200) );
 a61792a <=( A166  and  a61791a );
 a61793a <=( a61792a  and  a61787a );
 a61797a <=( (not A265)  and  A233 );
 a61798a <=( A232  and  a61797a );
 a61801a <=( (not A299)  and  (not A266) );
 a61804a <=( (not A302)  and  (not A301) );
 a61805a <=( a61804a  and  a61801a );
 a61806a <=( a61805a  and  a61798a );
 a61810a <=( (not A167)  and  (not A169) );
 a61811a <=( A170  and  a61810a );
 a61815a <=( (not A201)  and  (not A200) );
 a61816a <=( A166  and  a61815a );
 a61817a <=( a61816a  and  a61811a );
 a61821a <=( (not A236)  and  (not A235) );
 a61822a <=( (not A233)  and  a61821a );
 a61825a <=( A266  and  A265 );
 a61828a <=( (not A300)  and  A298 );
 a61829a <=( a61828a  and  a61825a );
 a61830a <=( a61829a  and  a61822a );
 a61834a <=( (not A167)  and  (not A169) );
 a61835a <=( A170  and  a61834a );
 a61839a <=( (not A201)  and  (not A200) );
 a61840a <=( A166  and  a61839a );
 a61841a <=( a61840a  and  a61835a );
 a61845a <=( (not A236)  and  (not A235) );
 a61846a <=( (not A233)  and  a61845a );
 a61849a <=( A266  and  A265 );
 a61852a <=( A299  and  A298 );
 a61853a <=( a61852a  and  a61849a );
 a61854a <=( a61853a  and  a61846a );
 a61858a <=( (not A167)  and  (not A169) );
 a61859a <=( A170  and  a61858a );
 a61863a <=( (not A201)  and  (not A200) );
 a61864a <=( A166  and  a61863a );
 a61865a <=( a61864a  and  a61859a );
 a61869a <=( (not A236)  and  (not A235) );
 a61870a <=( (not A233)  and  a61869a );
 a61873a <=( A266  and  A265 );
 a61876a <=( (not A299)  and  (not A298) );
 a61877a <=( a61876a  and  a61873a );
 a61878a <=( a61877a  and  a61870a );
 a61882a <=( (not A167)  and  (not A169) );
 a61883a <=( A170  and  a61882a );
 a61887a <=( (not A201)  and  (not A200) );
 a61888a <=( A166  and  a61887a );
 a61889a <=( a61888a  and  a61883a );
 a61893a <=( (not A236)  and  (not A235) );
 a61894a <=( (not A233)  and  a61893a );
 a61897a <=( (not A267)  and  (not A266) );
 a61900a <=( (not A300)  and  A298 );
 a61901a <=( a61900a  and  a61897a );
 a61902a <=( a61901a  and  a61894a );
 a61906a <=( (not A167)  and  (not A169) );
 a61907a <=( A170  and  a61906a );
 a61911a <=( (not A201)  and  (not A200) );
 a61912a <=( A166  and  a61911a );
 a61913a <=( a61912a  and  a61907a );
 a61917a <=( (not A236)  and  (not A235) );
 a61918a <=( (not A233)  and  a61917a );
 a61921a <=( (not A267)  and  (not A266) );
 a61924a <=( A299  and  A298 );
 a61925a <=( a61924a  and  a61921a );
 a61926a <=( a61925a  and  a61918a );
 a61930a <=( (not A167)  and  (not A169) );
 a61931a <=( A170  and  a61930a );
 a61935a <=( (not A201)  and  (not A200) );
 a61936a <=( A166  and  a61935a );
 a61937a <=( a61936a  and  a61931a );
 a61941a <=( (not A236)  and  (not A235) );
 a61942a <=( (not A233)  and  a61941a );
 a61945a <=( (not A267)  and  (not A266) );
 a61948a <=( (not A299)  and  (not A298) );
 a61949a <=( a61948a  and  a61945a );
 a61950a <=( a61949a  and  a61942a );
 a61954a <=( (not A167)  and  (not A169) );
 a61955a <=( A170  and  a61954a );
 a61959a <=( (not A201)  and  (not A200) );
 a61960a <=( A166  and  a61959a );
 a61961a <=( a61960a  and  a61955a );
 a61965a <=( (not A236)  and  (not A235) );
 a61966a <=( (not A233)  and  a61965a );
 a61969a <=( (not A266)  and  (not A265) );
 a61972a <=( (not A300)  and  A298 );
 a61973a <=( a61972a  and  a61969a );
 a61974a <=( a61973a  and  a61966a );
 a61978a <=( (not A167)  and  (not A169) );
 a61979a <=( A170  and  a61978a );
 a61983a <=( (not A201)  and  (not A200) );
 a61984a <=( A166  and  a61983a );
 a61985a <=( a61984a  and  a61979a );
 a61989a <=( (not A236)  and  (not A235) );
 a61990a <=( (not A233)  and  a61989a );
 a61993a <=( (not A266)  and  (not A265) );
 a61996a <=( A299  and  A298 );
 a61997a <=( a61996a  and  a61993a );
 a61998a <=( a61997a  and  a61990a );
 a62002a <=( (not A167)  and  (not A169) );
 a62003a <=( A170  and  a62002a );
 a62007a <=( (not A201)  and  (not A200) );
 a62008a <=( A166  and  a62007a );
 a62009a <=( a62008a  and  a62003a );
 a62013a <=( (not A236)  and  (not A235) );
 a62014a <=( (not A233)  and  a62013a );
 a62017a <=( (not A266)  and  (not A265) );
 a62020a <=( (not A299)  and  (not A298) );
 a62021a <=( a62020a  and  a62017a );
 a62022a <=( a62021a  and  a62014a );
 a62026a <=( (not A167)  and  (not A169) );
 a62027a <=( A170  and  a62026a );
 a62031a <=( (not A201)  and  (not A200) );
 a62032a <=( A166  and  a62031a );
 a62033a <=( a62032a  and  a62027a );
 a62037a <=( A265  and  (not A234) );
 a62038a <=( (not A233)  and  a62037a );
 a62041a <=( A298  and  A266 );
 a62044a <=( (not A302)  and  (not A301) );
 a62045a <=( a62044a  and  a62041a );
 a62046a <=( a62045a  and  a62038a );
 a62050a <=( (not A167)  and  (not A169) );
 a62051a <=( A170  and  a62050a );
 a62055a <=( (not A201)  and  (not A200) );
 a62056a <=( A166  and  a62055a );
 a62057a <=( a62056a  and  a62051a );
 a62061a <=( (not A266)  and  (not A234) );
 a62062a <=( (not A233)  and  a62061a );
 a62065a <=( (not A269)  and  (not A268) );
 a62068a <=( (not A300)  and  A298 );
 a62069a <=( a62068a  and  a62065a );
 a62070a <=( a62069a  and  a62062a );
 a62074a <=( (not A167)  and  (not A169) );
 a62075a <=( A170  and  a62074a );
 a62079a <=( (not A201)  and  (not A200) );
 a62080a <=( A166  and  a62079a );
 a62081a <=( a62080a  and  a62075a );
 a62085a <=( (not A266)  and  (not A234) );
 a62086a <=( (not A233)  and  a62085a );
 a62089a <=( (not A269)  and  (not A268) );
 a62092a <=( A299  and  A298 );
 a62093a <=( a62092a  and  a62089a );
 a62094a <=( a62093a  and  a62086a );
 a62098a <=( (not A167)  and  (not A169) );
 a62099a <=( A170  and  a62098a );
 a62103a <=( (not A201)  and  (not A200) );
 a62104a <=( A166  and  a62103a );
 a62105a <=( a62104a  and  a62099a );
 a62109a <=( (not A266)  and  (not A234) );
 a62110a <=( (not A233)  and  a62109a );
 a62113a <=( (not A269)  and  (not A268) );
 a62116a <=( (not A299)  and  (not A298) );
 a62117a <=( a62116a  and  a62113a );
 a62118a <=( a62117a  and  a62110a );
 a62122a <=( (not A167)  and  (not A169) );
 a62123a <=( A170  and  a62122a );
 a62127a <=( (not A201)  and  (not A200) );
 a62128a <=( A166  and  a62127a );
 a62129a <=( a62128a  and  a62123a );
 a62133a <=( (not A266)  and  (not A234) );
 a62134a <=( (not A233)  and  a62133a );
 a62137a <=( A298  and  (not A267) );
 a62140a <=( (not A302)  and  (not A301) );
 a62141a <=( a62140a  and  a62137a );
 a62142a <=( a62141a  and  a62134a );
 a62146a <=( (not A167)  and  (not A169) );
 a62147a <=( A170  and  a62146a );
 a62151a <=( (not A201)  and  (not A200) );
 a62152a <=( A166  and  a62151a );
 a62153a <=( a62152a  and  a62147a );
 a62157a <=( (not A265)  and  (not A234) );
 a62158a <=( (not A233)  and  a62157a );
 a62161a <=( A298  and  (not A266) );
 a62164a <=( (not A302)  and  (not A301) );
 a62165a <=( a62164a  and  a62161a );
 a62166a <=( a62165a  and  a62158a );
 a62170a <=( (not A167)  and  (not A169) );
 a62171a <=( A170  and  a62170a );
 a62175a <=( (not A201)  and  (not A200) );
 a62176a <=( A166  and  a62175a );
 a62177a <=( a62176a  and  a62171a );
 a62181a <=( A265  and  (not A233) );
 a62182a <=( (not A232)  and  a62181a );
 a62185a <=( A298  and  A266 );
 a62188a <=( (not A302)  and  (not A301) );
 a62189a <=( a62188a  and  a62185a );
 a62190a <=( a62189a  and  a62182a );
 a62194a <=( (not A167)  and  (not A169) );
 a62195a <=( A170  and  a62194a );
 a62199a <=( (not A201)  and  (not A200) );
 a62200a <=( A166  and  a62199a );
 a62201a <=( a62200a  and  a62195a );
 a62205a <=( (not A266)  and  (not A233) );
 a62206a <=( (not A232)  and  a62205a );
 a62209a <=( (not A269)  and  (not A268) );
 a62212a <=( (not A300)  and  A298 );
 a62213a <=( a62212a  and  a62209a );
 a62214a <=( a62213a  and  a62206a );
 a62218a <=( (not A167)  and  (not A169) );
 a62219a <=( A170  and  a62218a );
 a62223a <=( (not A201)  and  (not A200) );
 a62224a <=( A166  and  a62223a );
 a62225a <=( a62224a  and  a62219a );
 a62229a <=( (not A266)  and  (not A233) );
 a62230a <=( (not A232)  and  a62229a );
 a62233a <=( (not A269)  and  (not A268) );
 a62236a <=( A299  and  A298 );
 a62237a <=( a62236a  and  a62233a );
 a62238a <=( a62237a  and  a62230a );
 a62242a <=( (not A167)  and  (not A169) );
 a62243a <=( A170  and  a62242a );
 a62247a <=( (not A201)  and  (not A200) );
 a62248a <=( A166  and  a62247a );
 a62249a <=( a62248a  and  a62243a );
 a62253a <=( (not A266)  and  (not A233) );
 a62254a <=( (not A232)  and  a62253a );
 a62257a <=( (not A269)  and  (not A268) );
 a62260a <=( (not A299)  and  (not A298) );
 a62261a <=( a62260a  and  a62257a );
 a62262a <=( a62261a  and  a62254a );
 a62266a <=( (not A167)  and  (not A169) );
 a62267a <=( A170  and  a62266a );
 a62271a <=( (not A201)  and  (not A200) );
 a62272a <=( A166  and  a62271a );
 a62273a <=( a62272a  and  a62267a );
 a62277a <=( (not A266)  and  (not A233) );
 a62278a <=( (not A232)  and  a62277a );
 a62281a <=( A298  and  (not A267) );
 a62284a <=( (not A302)  and  (not A301) );
 a62285a <=( a62284a  and  a62281a );
 a62286a <=( a62285a  and  a62278a );
 a62290a <=( (not A167)  and  (not A169) );
 a62291a <=( A170  and  a62290a );
 a62295a <=( (not A201)  and  (not A200) );
 a62296a <=( A166  and  a62295a );
 a62297a <=( a62296a  and  a62291a );
 a62301a <=( (not A265)  and  (not A233) );
 a62302a <=( (not A232)  and  a62301a );
 a62305a <=( A298  and  (not A266) );
 a62308a <=( (not A302)  and  (not A301) );
 a62309a <=( a62308a  and  a62305a );
 a62310a <=( a62309a  and  a62302a );
 a62314a <=( (not A167)  and  (not A169) );
 a62315a <=( A170  and  a62314a );
 a62319a <=( (not A200)  and  (not A199) );
 a62320a <=( A166  and  a62319a );
 a62321a <=( a62320a  and  a62315a );
 a62325a <=( A265  and  A233 );
 a62326a <=( A232  and  a62325a );
 a62329a <=( (not A269)  and  (not A268) );
 a62332a <=( (not A300)  and  (not A299) );
 a62333a <=( a62332a  and  a62329a );
 a62334a <=( a62333a  and  a62326a );
 a62338a <=( (not A167)  and  (not A169) );
 a62339a <=( A170  and  a62338a );
 a62343a <=( (not A200)  and  (not A199) );
 a62344a <=( A166  and  a62343a );
 a62345a <=( a62344a  and  a62339a );
 a62349a <=( A265  and  A233 );
 a62350a <=( A232  and  a62349a );
 a62353a <=( (not A269)  and  (not A268) );
 a62356a <=( A299  and  A298 );
 a62357a <=( a62356a  and  a62353a );
 a62358a <=( a62357a  and  a62350a );
 a62362a <=( (not A167)  and  (not A169) );
 a62363a <=( A170  and  a62362a );
 a62367a <=( (not A200)  and  (not A199) );
 a62368a <=( A166  and  a62367a );
 a62369a <=( a62368a  and  a62363a );
 a62373a <=( A265  and  A233 );
 a62374a <=( A232  and  a62373a );
 a62377a <=( (not A269)  and  (not A268) );
 a62380a <=( (not A299)  and  (not A298) );
 a62381a <=( a62380a  and  a62377a );
 a62382a <=( a62381a  and  a62374a );
 a62386a <=( (not A167)  and  (not A169) );
 a62387a <=( A170  and  a62386a );
 a62391a <=( (not A200)  and  (not A199) );
 a62392a <=( A166  and  a62391a );
 a62393a <=( a62392a  and  a62387a );
 a62397a <=( A265  and  A233 );
 a62398a <=( A232  and  a62397a );
 a62401a <=( (not A299)  and  (not A267) );
 a62404a <=( (not A302)  and  (not A301) );
 a62405a <=( a62404a  and  a62401a );
 a62406a <=( a62405a  and  a62398a );
 a62410a <=( (not A167)  and  (not A169) );
 a62411a <=( A170  and  a62410a );
 a62415a <=( (not A200)  and  (not A199) );
 a62416a <=( A166  and  a62415a );
 a62417a <=( a62416a  and  a62411a );
 a62421a <=( A265  and  A233 );
 a62422a <=( A232  and  a62421a );
 a62425a <=( (not A299)  and  A266 );
 a62428a <=( (not A302)  and  (not A301) );
 a62429a <=( a62428a  and  a62425a );
 a62430a <=( a62429a  and  a62422a );
 a62434a <=( (not A167)  and  (not A169) );
 a62435a <=( A170  and  a62434a );
 a62439a <=( (not A200)  and  (not A199) );
 a62440a <=( A166  and  a62439a );
 a62441a <=( a62440a  and  a62435a );
 a62445a <=( (not A265)  and  A233 );
 a62446a <=( A232  and  a62445a );
 a62449a <=( (not A299)  and  (not A266) );
 a62452a <=( (not A302)  and  (not A301) );
 a62453a <=( a62452a  and  a62449a );
 a62454a <=( a62453a  and  a62446a );
 a62458a <=( (not A167)  and  (not A169) );
 a62459a <=( A170  and  a62458a );
 a62463a <=( (not A200)  and  (not A199) );
 a62464a <=( A166  and  a62463a );
 a62465a <=( a62464a  and  a62459a );
 a62469a <=( (not A236)  and  (not A235) );
 a62470a <=( (not A233)  and  a62469a );
 a62473a <=( A266  and  A265 );
 a62476a <=( (not A300)  and  A298 );
 a62477a <=( a62476a  and  a62473a );
 a62478a <=( a62477a  and  a62470a );
 a62482a <=( (not A167)  and  (not A169) );
 a62483a <=( A170  and  a62482a );
 a62487a <=( (not A200)  and  (not A199) );
 a62488a <=( A166  and  a62487a );
 a62489a <=( a62488a  and  a62483a );
 a62493a <=( (not A236)  and  (not A235) );
 a62494a <=( (not A233)  and  a62493a );
 a62497a <=( A266  and  A265 );
 a62500a <=( A299  and  A298 );
 a62501a <=( a62500a  and  a62497a );
 a62502a <=( a62501a  and  a62494a );
 a62506a <=( (not A167)  and  (not A169) );
 a62507a <=( A170  and  a62506a );
 a62511a <=( (not A200)  and  (not A199) );
 a62512a <=( A166  and  a62511a );
 a62513a <=( a62512a  and  a62507a );
 a62517a <=( (not A236)  and  (not A235) );
 a62518a <=( (not A233)  and  a62517a );
 a62521a <=( A266  and  A265 );
 a62524a <=( (not A299)  and  (not A298) );
 a62525a <=( a62524a  and  a62521a );
 a62526a <=( a62525a  and  a62518a );
 a62530a <=( (not A167)  and  (not A169) );
 a62531a <=( A170  and  a62530a );
 a62535a <=( (not A200)  and  (not A199) );
 a62536a <=( A166  and  a62535a );
 a62537a <=( a62536a  and  a62531a );
 a62541a <=( (not A236)  and  (not A235) );
 a62542a <=( (not A233)  and  a62541a );
 a62545a <=( (not A267)  and  (not A266) );
 a62548a <=( (not A300)  and  A298 );
 a62549a <=( a62548a  and  a62545a );
 a62550a <=( a62549a  and  a62542a );
 a62554a <=( (not A167)  and  (not A169) );
 a62555a <=( A170  and  a62554a );
 a62559a <=( (not A200)  and  (not A199) );
 a62560a <=( A166  and  a62559a );
 a62561a <=( a62560a  and  a62555a );
 a62565a <=( (not A236)  and  (not A235) );
 a62566a <=( (not A233)  and  a62565a );
 a62569a <=( (not A267)  and  (not A266) );
 a62572a <=( A299  and  A298 );
 a62573a <=( a62572a  and  a62569a );
 a62574a <=( a62573a  and  a62566a );
 a62578a <=( (not A167)  and  (not A169) );
 a62579a <=( A170  and  a62578a );
 a62583a <=( (not A200)  and  (not A199) );
 a62584a <=( A166  and  a62583a );
 a62585a <=( a62584a  and  a62579a );
 a62589a <=( (not A236)  and  (not A235) );
 a62590a <=( (not A233)  and  a62589a );
 a62593a <=( (not A267)  and  (not A266) );
 a62596a <=( (not A299)  and  (not A298) );
 a62597a <=( a62596a  and  a62593a );
 a62598a <=( a62597a  and  a62590a );
 a62602a <=( (not A167)  and  (not A169) );
 a62603a <=( A170  and  a62602a );
 a62607a <=( (not A200)  and  (not A199) );
 a62608a <=( A166  and  a62607a );
 a62609a <=( a62608a  and  a62603a );
 a62613a <=( (not A236)  and  (not A235) );
 a62614a <=( (not A233)  and  a62613a );
 a62617a <=( (not A266)  and  (not A265) );
 a62620a <=( (not A300)  and  A298 );
 a62621a <=( a62620a  and  a62617a );
 a62622a <=( a62621a  and  a62614a );
 a62626a <=( (not A167)  and  (not A169) );
 a62627a <=( A170  and  a62626a );
 a62631a <=( (not A200)  and  (not A199) );
 a62632a <=( A166  and  a62631a );
 a62633a <=( a62632a  and  a62627a );
 a62637a <=( (not A236)  and  (not A235) );
 a62638a <=( (not A233)  and  a62637a );
 a62641a <=( (not A266)  and  (not A265) );
 a62644a <=( A299  and  A298 );
 a62645a <=( a62644a  and  a62641a );
 a62646a <=( a62645a  and  a62638a );
 a62650a <=( (not A167)  and  (not A169) );
 a62651a <=( A170  and  a62650a );
 a62655a <=( (not A200)  and  (not A199) );
 a62656a <=( A166  and  a62655a );
 a62657a <=( a62656a  and  a62651a );
 a62661a <=( (not A236)  and  (not A235) );
 a62662a <=( (not A233)  and  a62661a );
 a62665a <=( (not A266)  and  (not A265) );
 a62668a <=( (not A299)  and  (not A298) );
 a62669a <=( a62668a  and  a62665a );
 a62670a <=( a62669a  and  a62662a );
 a62674a <=( (not A167)  and  (not A169) );
 a62675a <=( A170  and  a62674a );
 a62679a <=( (not A200)  and  (not A199) );
 a62680a <=( A166  and  a62679a );
 a62681a <=( a62680a  and  a62675a );
 a62685a <=( A265  and  (not A234) );
 a62686a <=( (not A233)  and  a62685a );
 a62689a <=( A298  and  A266 );
 a62692a <=( (not A302)  and  (not A301) );
 a62693a <=( a62692a  and  a62689a );
 a62694a <=( a62693a  and  a62686a );
 a62698a <=( (not A167)  and  (not A169) );
 a62699a <=( A170  and  a62698a );
 a62703a <=( (not A200)  and  (not A199) );
 a62704a <=( A166  and  a62703a );
 a62705a <=( a62704a  and  a62699a );
 a62709a <=( (not A266)  and  (not A234) );
 a62710a <=( (not A233)  and  a62709a );
 a62713a <=( (not A269)  and  (not A268) );
 a62716a <=( (not A300)  and  A298 );
 a62717a <=( a62716a  and  a62713a );
 a62718a <=( a62717a  and  a62710a );
 a62722a <=( (not A167)  and  (not A169) );
 a62723a <=( A170  and  a62722a );
 a62727a <=( (not A200)  and  (not A199) );
 a62728a <=( A166  and  a62727a );
 a62729a <=( a62728a  and  a62723a );
 a62733a <=( (not A266)  and  (not A234) );
 a62734a <=( (not A233)  and  a62733a );
 a62737a <=( (not A269)  and  (not A268) );
 a62740a <=( A299  and  A298 );
 a62741a <=( a62740a  and  a62737a );
 a62742a <=( a62741a  and  a62734a );
 a62746a <=( (not A167)  and  (not A169) );
 a62747a <=( A170  and  a62746a );
 a62751a <=( (not A200)  and  (not A199) );
 a62752a <=( A166  and  a62751a );
 a62753a <=( a62752a  and  a62747a );
 a62757a <=( (not A266)  and  (not A234) );
 a62758a <=( (not A233)  and  a62757a );
 a62761a <=( (not A269)  and  (not A268) );
 a62764a <=( (not A299)  and  (not A298) );
 a62765a <=( a62764a  and  a62761a );
 a62766a <=( a62765a  and  a62758a );
 a62770a <=( (not A167)  and  (not A169) );
 a62771a <=( A170  and  a62770a );
 a62775a <=( (not A200)  and  (not A199) );
 a62776a <=( A166  and  a62775a );
 a62777a <=( a62776a  and  a62771a );
 a62781a <=( (not A266)  and  (not A234) );
 a62782a <=( (not A233)  and  a62781a );
 a62785a <=( A298  and  (not A267) );
 a62788a <=( (not A302)  and  (not A301) );
 a62789a <=( a62788a  and  a62785a );
 a62790a <=( a62789a  and  a62782a );
 a62794a <=( (not A167)  and  (not A169) );
 a62795a <=( A170  and  a62794a );
 a62799a <=( (not A200)  and  (not A199) );
 a62800a <=( A166  and  a62799a );
 a62801a <=( a62800a  and  a62795a );
 a62805a <=( (not A265)  and  (not A234) );
 a62806a <=( (not A233)  and  a62805a );
 a62809a <=( A298  and  (not A266) );
 a62812a <=( (not A302)  and  (not A301) );
 a62813a <=( a62812a  and  a62809a );
 a62814a <=( a62813a  and  a62806a );
 a62818a <=( (not A167)  and  (not A169) );
 a62819a <=( A170  and  a62818a );
 a62823a <=( (not A200)  and  (not A199) );
 a62824a <=( A166  and  a62823a );
 a62825a <=( a62824a  and  a62819a );
 a62829a <=( A265  and  (not A233) );
 a62830a <=( (not A232)  and  a62829a );
 a62833a <=( A298  and  A266 );
 a62836a <=( (not A302)  and  (not A301) );
 a62837a <=( a62836a  and  a62833a );
 a62838a <=( a62837a  and  a62830a );
 a62842a <=( (not A167)  and  (not A169) );
 a62843a <=( A170  and  a62842a );
 a62847a <=( (not A200)  and  (not A199) );
 a62848a <=( A166  and  a62847a );
 a62849a <=( a62848a  and  a62843a );
 a62853a <=( (not A266)  and  (not A233) );
 a62854a <=( (not A232)  and  a62853a );
 a62857a <=( (not A269)  and  (not A268) );
 a62860a <=( (not A300)  and  A298 );
 a62861a <=( a62860a  and  a62857a );
 a62862a <=( a62861a  and  a62854a );
 a62866a <=( (not A167)  and  (not A169) );
 a62867a <=( A170  and  a62866a );
 a62871a <=( (not A200)  and  (not A199) );
 a62872a <=( A166  and  a62871a );
 a62873a <=( a62872a  and  a62867a );
 a62877a <=( (not A266)  and  (not A233) );
 a62878a <=( (not A232)  and  a62877a );
 a62881a <=( (not A269)  and  (not A268) );
 a62884a <=( A299  and  A298 );
 a62885a <=( a62884a  and  a62881a );
 a62886a <=( a62885a  and  a62878a );
 a62890a <=( (not A167)  and  (not A169) );
 a62891a <=( A170  and  a62890a );
 a62895a <=( (not A200)  and  (not A199) );
 a62896a <=( A166  and  a62895a );
 a62897a <=( a62896a  and  a62891a );
 a62901a <=( (not A266)  and  (not A233) );
 a62902a <=( (not A232)  and  a62901a );
 a62905a <=( (not A269)  and  (not A268) );
 a62908a <=( (not A299)  and  (not A298) );
 a62909a <=( a62908a  and  a62905a );
 a62910a <=( a62909a  and  a62902a );
 a62914a <=( (not A167)  and  (not A169) );
 a62915a <=( A170  and  a62914a );
 a62919a <=( (not A200)  and  (not A199) );
 a62920a <=( A166  and  a62919a );
 a62921a <=( a62920a  and  a62915a );
 a62925a <=( (not A266)  and  (not A233) );
 a62926a <=( (not A232)  and  a62925a );
 a62929a <=( A298  and  (not A267) );
 a62932a <=( (not A302)  and  (not A301) );
 a62933a <=( a62932a  and  a62929a );
 a62934a <=( a62933a  and  a62926a );
 a62938a <=( (not A167)  and  (not A169) );
 a62939a <=( A170  and  a62938a );
 a62943a <=( (not A200)  and  (not A199) );
 a62944a <=( A166  and  a62943a );
 a62945a <=( a62944a  and  a62939a );
 a62949a <=( (not A265)  and  (not A233) );
 a62950a <=( (not A232)  and  a62949a );
 a62953a <=( A298  and  (not A266) );
 a62956a <=( (not A302)  and  (not A301) );
 a62957a <=( a62956a  and  a62953a );
 a62958a <=( a62957a  and  a62950a );
 a62962a <=( (not A168)  and  (not A169) );
 a62963a <=( (not A170)  and  a62962a );
 a62967a <=( A201  and  (not A200) );
 a62968a <=( A199  and  a62967a );
 a62969a <=( a62968a  and  a62963a );
 a62973a <=( A233  and  A232 );
 a62974a <=( A202  and  a62973a );
 a62977a <=( (not A267)  and  A265 );
 a62980a <=( (not A300)  and  (not A299) );
 a62981a <=( a62980a  and  a62977a );
 a62982a <=( a62981a  and  a62974a );
 a62986a <=( (not A168)  and  (not A169) );
 a62987a <=( (not A170)  and  a62986a );
 a62991a <=( A201  and  (not A200) );
 a62992a <=( A199  and  a62991a );
 a62993a <=( a62992a  and  a62987a );
 a62997a <=( A233  and  A232 );
 a62998a <=( A202  and  a62997a );
 a63001a <=( (not A267)  and  A265 );
 a63004a <=( A299  and  A298 );
 a63005a <=( a63004a  and  a63001a );
 a63006a <=( a63005a  and  a62998a );
 a63010a <=( (not A168)  and  (not A169) );
 a63011a <=( (not A170)  and  a63010a );
 a63015a <=( A201  and  (not A200) );
 a63016a <=( A199  and  a63015a );
 a63017a <=( a63016a  and  a63011a );
 a63021a <=( A233  and  A232 );
 a63022a <=( A202  and  a63021a );
 a63025a <=( (not A267)  and  A265 );
 a63028a <=( (not A299)  and  (not A298) );
 a63029a <=( a63028a  and  a63025a );
 a63030a <=( a63029a  and  a63022a );
 a63034a <=( (not A168)  and  (not A169) );
 a63035a <=( (not A170)  and  a63034a );
 a63039a <=( A201  and  (not A200) );
 a63040a <=( A199  and  a63039a );
 a63041a <=( a63040a  and  a63035a );
 a63045a <=( A233  and  A232 );
 a63046a <=( A202  and  a63045a );
 a63049a <=( A266  and  A265 );
 a63052a <=( (not A300)  and  (not A299) );
 a63053a <=( a63052a  and  a63049a );
 a63054a <=( a63053a  and  a63046a );
 a63058a <=( (not A168)  and  (not A169) );
 a63059a <=( (not A170)  and  a63058a );
 a63063a <=( A201  and  (not A200) );
 a63064a <=( A199  and  a63063a );
 a63065a <=( a63064a  and  a63059a );
 a63069a <=( A233  and  A232 );
 a63070a <=( A202  and  a63069a );
 a63073a <=( A266  and  A265 );
 a63076a <=( A299  and  A298 );
 a63077a <=( a63076a  and  a63073a );
 a63078a <=( a63077a  and  a63070a );
 a63082a <=( (not A168)  and  (not A169) );
 a63083a <=( (not A170)  and  a63082a );
 a63087a <=( A201  and  (not A200) );
 a63088a <=( A199  and  a63087a );
 a63089a <=( a63088a  and  a63083a );
 a63093a <=( A233  and  A232 );
 a63094a <=( A202  and  a63093a );
 a63097a <=( A266  and  A265 );
 a63100a <=( (not A299)  and  (not A298) );
 a63101a <=( a63100a  and  a63097a );
 a63102a <=( a63101a  and  a63094a );
 a63106a <=( (not A168)  and  (not A169) );
 a63107a <=( (not A170)  and  a63106a );
 a63111a <=( A201  and  (not A200) );
 a63112a <=( A199  and  a63111a );
 a63113a <=( a63112a  and  a63107a );
 a63117a <=( A233  and  A232 );
 a63118a <=( A202  and  a63117a );
 a63121a <=( (not A266)  and  (not A265) );
 a63124a <=( (not A300)  and  (not A299) );
 a63125a <=( a63124a  and  a63121a );
 a63126a <=( a63125a  and  a63118a );
 a63130a <=( (not A168)  and  (not A169) );
 a63131a <=( (not A170)  and  a63130a );
 a63135a <=( A201  and  (not A200) );
 a63136a <=( A199  and  a63135a );
 a63137a <=( a63136a  and  a63131a );
 a63141a <=( A233  and  A232 );
 a63142a <=( A202  and  a63141a );
 a63145a <=( (not A266)  and  (not A265) );
 a63148a <=( A299  and  A298 );
 a63149a <=( a63148a  and  a63145a );
 a63150a <=( a63149a  and  a63142a );
 a63154a <=( (not A168)  and  (not A169) );
 a63155a <=( (not A170)  and  a63154a );
 a63159a <=( A201  and  (not A200) );
 a63160a <=( A199  and  a63159a );
 a63161a <=( a63160a  and  a63155a );
 a63165a <=( A233  and  A232 );
 a63166a <=( A202  and  a63165a );
 a63169a <=( (not A266)  and  (not A265) );
 a63172a <=( (not A299)  and  (not A298) );
 a63173a <=( a63172a  and  a63169a );
 a63174a <=( a63173a  and  a63166a );
 a63178a <=( (not A168)  and  (not A169) );
 a63179a <=( (not A170)  and  a63178a );
 a63183a <=( A201  and  (not A200) );
 a63184a <=( A199  and  a63183a );
 a63185a <=( a63184a  and  a63179a );
 a63189a <=( A233  and  (not A232) );
 a63190a <=( A202  and  a63189a );
 a63193a <=( (not A299)  and  A298 );
 a63196a <=( A301  and  A300 );
 a63197a <=( a63196a  and  a63193a );
 a63198a <=( a63197a  and  a63190a );
 a63202a <=( (not A168)  and  (not A169) );
 a63203a <=( (not A170)  and  a63202a );
 a63207a <=( A201  and  (not A200) );
 a63208a <=( A199  and  a63207a );
 a63209a <=( a63208a  and  a63203a );
 a63213a <=( A233  and  (not A232) );
 a63214a <=( A202  and  a63213a );
 a63217a <=( (not A299)  and  A298 );
 a63220a <=( A302  and  A300 );
 a63221a <=( a63220a  and  a63217a );
 a63222a <=( a63221a  and  a63214a );
 a63226a <=( (not A168)  and  (not A169) );
 a63227a <=( (not A170)  and  a63226a );
 a63231a <=( A201  and  (not A200) );
 a63232a <=( A199  and  a63231a );
 a63233a <=( a63232a  and  a63227a );
 a63237a <=( A233  and  (not A232) );
 a63238a <=( A202  and  a63237a );
 a63241a <=( (not A266)  and  A265 );
 a63244a <=( A268  and  A267 );
 a63245a <=( a63244a  and  a63241a );
 a63246a <=( a63245a  and  a63238a );
 a63250a <=( (not A168)  and  (not A169) );
 a63251a <=( (not A170)  and  a63250a );
 a63255a <=( A201  and  (not A200) );
 a63256a <=( A199  and  a63255a );
 a63257a <=( a63256a  and  a63251a );
 a63261a <=( A233  and  (not A232) );
 a63262a <=( A202  and  a63261a );
 a63265a <=( (not A266)  and  A265 );
 a63268a <=( A269  and  A267 );
 a63269a <=( a63268a  and  a63265a );
 a63270a <=( a63269a  and  a63262a );
 a63274a <=( (not A168)  and  (not A169) );
 a63275a <=( (not A170)  and  a63274a );
 a63279a <=( A201  and  (not A200) );
 a63280a <=( A199  and  a63279a );
 a63281a <=( a63280a  and  a63275a );
 a63285a <=( (not A234)  and  (not A233) );
 a63286a <=( A202  and  a63285a );
 a63289a <=( A266  and  A265 );
 a63292a <=( (not A300)  and  A298 );
 a63293a <=( a63292a  and  a63289a );
 a63294a <=( a63293a  and  a63286a );
 a63298a <=( (not A168)  and  (not A169) );
 a63299a <=( (not A170)  and  a63298a );
 a63303a <=( A201  and  (not A200) );
 a63304a <=( A199  and  a63303a );
 a63305a <=( a63304a  and  a63299a );
 a63309a <=( (not A234)  and  (not A233) );
 a63310a <=( A202  and  a63309a );
 a63313a <=( A266  and  A265 );
 a63316a <=( A299  and  A298 );
 a63317a <=( a63316a  and  a63313a );
 a63318a <=( a63317a  and  a63310a );
 a63322a <=( (not A168)  and  (not A169) );
 a63323a <=( (not A170)  and  a63322a );
 a63327a <=( A201  and  (not A200) );
 a63328a <=( A199  and  a63327a );
 a63329a <=( a63328a  and  a63323a );
 a63333a <=( (not A234)  and  (not A233) );
 a63334a <=( A202  and  a63333a );
 a63337a <=( A266  and  A265 );
 a63340a <=( (not A299)  and  (not A298) );
 a63341a <=( a63340a  and  a63337a );
 a63342a <=( a63341a  and  a63334a );
 a63346a <=( (not A168)  and  (not A169) );
 a63347a <=( (not A170)  and  a63346a );
 a63351a <=( A201  and  (not A200) );
 a63352a <=( A199  and  a63351a );
 a63353a <=( a63352a  and  a63347a );
 a63357a <=( (not A234)  and  (not A233) );
 a63358a <=( A202  and  a63357a );
 a63361a <=( (not A267)  and  (not A266) );
 a63364a <=( (not A300)  and  A298 );
 a63365a <=( a63364a  and  a63361a );
 a63366a <=( a63365a  and  a63358a );
 a63370a <=( (not A168)  and  (not A169) );
 a63371a <=( (not A170)  and  a63370a );
 a63375a <=( A201  and  (not A200) );
 a63376a <=( A199  and  a63375a );
 a63377a <=( a63376a  and  a63371a );
 a63381a <=( (not A234)  and  (not A233) );
 a63382a <=( A202  and  a63381a );
 a63385a <=( (not A267)  and  (not A266) );
 a63388a <=( A299  and  A298 );
 a63389a <=( a63388a  and  a63385a );
 a63390a <=( a63389a  and  a63382a );
 a63394a <=( (not A168)  and  (not A169) );
 a63395a <=( (not A170)  and  a63394a );
 a63399a <=( A201  and  (not A200) );
 a63400a <=( A199  and  a63399a );
 a63401a <=( a63400a  and  a63395a );
 a63405a <=( (not A234)  and  (not A233) );
 a63406a <=( A202  and  a63405a );
 a63409a <=( (not A267)  and  (not A266) );
 a63412a <=( (not A299)  and  (not A298) );
 a63413a <=( a63412a  and  a63409a );
 a63414a <=( a63413a  and  a63406a );
 a63418a <=( (not A168)  and  (not A169) );
 a63419a <=( (not A170)  and  a63418a );
 a63423a <=( A201  and  (not A200) );
 a63424a <=( A199  and  a63423a );
 a63425a <=( a63424a  and  a63419a );
 a63429a <=( (not A234)  and  (not A233) );
 a63430a <=( A202  and  a63429a );
 a63433a <=( (not A266)  and  (not A265) );
 a63436a <=( (not A300)  and  A298 );
 a63437a <=( a63436a  and  a63433a );
 a63438a <=( a63437a  and  a63430a );
 a63442a <=( (not A168)  and  (not A169) );
 a63443a <=( (not A170)  and  a63442a );
 a63447a <=( A201  and  (not A200) );
 a63448a <=( A199  and  a63447a );
 a63449a <=( a63448a  and  a63443a );
 a63453a <=( (not A234)  and  (not A233) );
 a63454a <=( A202  and  a63453a );
 a63457a <=( (not A266)  and  (not A265) );
 a63460a <=( A299  and  A298 );
 a63461a <=( a63460a  and  a63457a );
 a63462a <=( a63461a  and  a63454a );
 a63466a <=( (not A168)  and  (not A169) );
 a63467a <=( (not A170)  and  a63466a );
 a63471a <=( A201  and  (not A200) );
 a63472a <=( A199  and  a63471a );
 a63473a <=( a63472a  and  a63467a );
 a63477a <=( (not A234)  and  (not A233) );
 a63478a <=( A202  and  a63477a );
 a63481a <=( (not A266)  and  (not A265) );
 a63484a <=( (not A299)  and  (not A298) );
 a63485a <=( a63484a  and  a63481a );
 a63486a <=( a63485a  and  a63478a );
 a63490a <=( (not A168)  and  (not A169) );
 a63491a <=( (not A170)  and  a63490a );
 a63495a <=( A201  and  (not A200) );
 a63496a <=( A199  and  a63495a );
 a63497a <=( a63496a  and  a63491a );
 a63501a <=( (not A233)  and  A232 );
 a63502a <=( A202  and  a63501a );
 a63505a <=( A235  and  A234 );
 a63508a <=( A299  and  (not A298) );
 a63509a <=( a63508a  and  a63505a );
 a63510a <=( a63509a  and  a63502a );
 a63514a <=( (not A168)  and  (not A169) );
 a63515a <=( (not A170)  and  a63514a );
 a63519a <=( A201  and  (not A200) );
 a63520a <=( A199  and  a63519a );
 a63521a <=( a63520a  and  a63515a );
 a63525a <=( (not A233)  and  A232 );
 a63526a <=( A202  and  a63525a );
 a63529a <=( A235  and  A234 );
 a63532a <=( A266  and  (not A265) );
 a63533a <=( a63532a  and  a63529a );
 a63534a <=( a63533a  and  a63526a );
 a63538a <=( (not A168)  and  (not A169) );
 a63539a <=( (not A170)  and  a63538a );
 a63543a <=( A201  and  (not A200) );
 a63544a <=( A199  and  a63543a );
 a63545a <=( a63544a  and  a63539a );
 a63549a <=( (not A233)  and  A232 );
 a63550a <=( A202  and  a63549a );
 a63553a <=( A236  and  A234 );
 a63556a <=( A299  and  (not A298) );
 a63557a <=( a63556a  and  a63553a );
 a63558a <=( a63557a  and  a63550a );
 a63562a <=( (not A168)  and  (not A169) );
 a63563a <=( (not A170)  and  a63562a );
 a63567a <=( A201  and  (not A200) );
 a63568a <=( A199  and  a63567a );
 a63569a <=( a63568a  and  a63563a );
 a63573a <=( (not A233)  and  A232 );
 a63574a <=( A202  and  a63573a );
 a63577a <=( A236  and  A234 );
 a63580a <=( A266  and  (not A265) );
 a63581a <=( a63580a  and  a63577a );
 a63582a <=( a63581a  and  a63574a );
 a63586a <=( (not A168)  and  (not A169) );
 a63587a <=( (not A170)  and  a63586a );
 a63591a <=( A201  and  (not A200) );
 a63592a <=( A199  and  a63591a );
 a63593a <=( a63592a  and  a63587a );
 a63597a <=( (not A233)  and  (not A232) );
 a63598a <=( A202  and  a63597a );
 a63601a <=( A266  and  A265 );
 a63604a <=( (not A300)  and  A298 );
 a63605a <=( a63604a  and  a63601a );
 a63606a <=( a63605a  and  a63598a );
 a63610a <=( (not A168)  and  (not A169) );
 a63611a <=( (not A170)  and  a63610a );
 a63615a <=( A201  and  (not A200) );
 a63616a <=( A199  and  a63615a );
 a63617a <=( a63616a  and  a63611a );
 a63621a <=( (not A233)  and  (not A232) );
 a63622a <=( A202  and  a63621a );
 a63625a <=( A266  and  A265 );
 a63628a <=( A299  and  A298 );
 a63629a <=( a63628a  and  a63625a );
 a63630a <=( a63629a  and  a63622a );
 a63634a <=( (not A168)  and  (not A169) );
 a63635a <=( (not A170)  and  a63634a );
 a63639a <=( A201  and  (not A200) );
 a63640a <=( A199  and  a63639a );
 a63641a <=( a63640a  and  a63635a );
 a63645a <=( (not A233)  and  (not A232) );
 a63646a <=( A202  and  a63645a );
 a63649a <=( A266  and  A265 );
 a63652a <=( (not A299)  and  (not A298) );
 a63653a <=( a63652a  and  a63649a );
 a63654a <=( a63653a  and  a63646a );
 a63658a <=( (not A168)  and  (not A169) );
 a63659a <=( (not A170)  and  a63658a );
 a63663a <=( A201  and  (not A200) );
 a63664a <=( A199  and  a63663a );
 a63665a <=( a63664a  and  a63659a );
 a63669a <=( (not A233)  and  (not A232) );
 a63670a <=( A202  and  a63669a );
 a63673a <=( (not A267)  and  (not A266) );
 a63676a <=( (not A300)  and  A298 );
 a63677a <=( a63676a  and  a63673a );
 a63678a <=( a63677a  and  a63670a );
 a63682a <=( (not A168)  and  (not A169) );
 a63683a <=( (not A170)  and  a63682a );
 a63687a <=( A201  and  (not A200) );
 a63688a <=( A199  and  a63687a );
 a63689a <=( a63688a  and  a63683a );
 a63693a <=( (not A233)  and  (not A232) );
 a63694a <=( A202  and  a63693a );
 a63697a <=( (not A267)  and  (not A266) );
 a63700a <=( A299  and  A298 );
 a63701a <=( a63700a  and  a63697a );
 a63702a <=( a63701a  and  a63694a );
 a63706a <=( (not A168)  and  (not A169) );
 a63707a <=( (not A170)  and  a63706a );
 a63711a <=( A201  and  (not A200) );
 a63712a <=( A199  and  a63711a );
 a63713a <=( a63712a  and  a63707a );
 a63717a <=( (not A233)  and  (not A232) );
 a63718a <=( A202  and  a63717a );
 a63721a <=( (not A267)  and  (not A266) );
 a63724a <=( (not A299)  and  (not A298) );
 a63725a <=( a63724a  and  a63721a );
 a63726a <=( a63725a  and  a63718a );
 a63730a <=( (not A168)  and  (not A169) );
 a63731a <=( (not A170)  and  a63730a );
 a63735a <=( A201  and  (not A200) );
 a63736a <=( A199  and  a63735a );
 a63737a <=( a63736a  and  a63731a );
 a63741a <=( (not A233)  and  (not A232) );
 a63742a <=( A202  and  a63741a );
 a63745a <=( (not A266)  and  (not A265) );
 a63748a <=( (not A300)  and  A298 );
 a63749a <=( a63748a  and  a63745a );
 a63750a <=( a63749a  and  a63742a );
 a63754a <=( (not A168)  and  (not A169) );
 a63755a <=( (not A170)  and  a63754a );
 a63759a <=( A201  and  (not A200) );
 a63760a <=( A199  and  a63759a );
 a63761a <=( a63760a  and  a63755a );
 a63765a <=( (not A233)  and  (not A232) );
 a63766a <=( A202  and  a63765a );
 a63769a <=( (not A266)  and  (not A265) );
 a63772a <=( A299  and  A298 );
 a63773a <=( a63772a  and  a63769a );
 a63774a <=( a63773a  and  a63766a );
 a63778a <=( (not A168)  and  (not A169) );
 a63779a <=( (not A170)  and  a63778a );
 a63783a <=( A201  and  (not A200) );
 a63784a <=( A199  and  a63783a );
 a63785a <=( a63784a  and  a63779a );
 a63789a <=( (not A233)  and  (not A232) );
 a63790a <=( A202  and  a63789a );
 a63793a <=( (not A266)  and  (not A265) );
 a63796a <=( (not A299)  and  (not A298) );
 a63797a <=( a63796a  and  a63793a );
 a63798a <=( a63797a  and  a63790a );
 a63802a <=( (not A168)  and  (not A169) );
 a63803a <=( (not A170)  and  a63802a );
 a63807a <=( A201  and  (not A200) );
 a63808a <=( A199  and  a63807a );
 a63809a <=( a63808a  and  a63803a );
 a63813a <=( A233  and  A232 );
 a63814a <=( A203  and  a63813a );
 a63817a <=( (not A267)  and  A265 );
 a63820a <=( (not A300)  and  (not A299) );
 a63821a <=( a63820a  and  a63817a );
 a63822a <=( a63821a  and  a63814a );
 a63826a <=( (not A168)  and  (not A169) );
 a63827a <=( (not A170)  and  a63826a );
 a63831a <=( A201  and  (not A200) );
 a63832a <=( A199  and  a63831a );
 a63833a <=( a63832a  and  a63827a );
 a63837a <=( A233  and  A232 );
 a63838a <=( A203  and  a63837a );
 a63841a <=( (not A267)  and  A265 );
 a63844a <=( A299  and  A298 );
 a63845a <=( a63844a  and  a63841a );
 a63846a <=( a63845a  and  a63838a );
 a63850a <=( (not A168)  and  (not A169) );
 a63851a <=( (not A170)  and  a63850a );
 a63855a <=( A201  and  (not A200) );
 a63856a <=( A199  and  a63855a );
 a63857a <=( a63856a  and  a63851a );
 a63861a <=( A233  and  A232 );
 a63862a <=( A203  and  a63861a );
 a63865a <=( (not A267)  and  A265 );
 a63868a <=( (not A299)  and  (not A298) );
 a63869a <=( a63868a  and  a63865a );
 a63870a <=( a63869a  and  a63862a );
 a63874a <=( (not A168)  and  (not A169) );
 a63875a <=( (not A170)  and  a63874a );
 a63879a <=( A201  and  (not A200) );
 a63880a <=( A199  and  a63879a );
 a63881a <=( a63880a  and  a63875a );
 a63885a <=( A233  and  A232 );
 a63886a <=( A203  and  a63885a );
 a63889a <=( A266  and  A265 );
 a63892a <=( (not A300)  and  (not A299) );
 a63893a <=( a63892a  and  a63889a );
 a63894a <=( a63893a  and  a63886a );
 a63898a <=( (not A168)  and  (not A169) );
 a63899a <=( (not A170)  and  a63898a );
 a63903a <=( A201  and  (not A200) );
 a63904a <=( A199  and  a63903a );
 a63905a <=( a63904a  and  a63899a );
 a63909a <=( A233  and  A232 );
 a63910a <=( A203  and  a63909a );
 a63913a <=( A266  and  A265 );
 a63916a <=( A299  and  A298 );
 a63917a <=( a63916a  and  a63913a );
 a63918a <=( a63917a  and  a63910a );
 a63922a <=( (not A168)  and  (not A169) );
 a63923a <=( (not A170)  and  a63922a );
 a63927a <=( A201  and  (not A200) );
 a63928a <=( A199  and  a63927a );
 a63929a <=( a63928a  and  a63923a );
 a63933a <=( A233  and  A232 );
 a63934a <=( A203  and  a63933a );
 a63937a <=( A266  and  A265 );
 a63940a <=( (not A299)  and  (not A298) );
 a63941a <=( a63940a  and  a63937a );
 a63942a <=( a63941a  and  a63934a );
 a63946a <=( (not A168)  and  (not A169) );
 a63947a <=( (not A170)  and  a63946a );
 a63951a <=( A201  and  (not A200) );
 a63952a <=( A199  and  a63951a );
 a63953a <=( a63952a  and  a63947a );
 a63957a <=( A233  and  A232 );
 a63958a <=( A203  and  a63957a );
 a63961a <=( (not A266)  and  (not A265) );
 a63964a <=( (not A300)  and  (not A299) );
 a63965a <=( a63964a  and  a63961a );
 a63966a <=( a63965a  and  a63958a );
 a63970a <=( (not A168)  and  (not A169) );
 a63971a <=( (not A170)  and  a63970a );
 a63975a <=( A201  and  (not A200) );
 a63976a <=( A199  and  a63975a );
 a63977a <=( a63976a  and  a63971a );
 a63981a <=( A233  and  A232 );
 a63982a <=( A203  and  a63981a );
 a63985a <=( (not A266)  and  (not A265) );
 a63988a <=( A299  and  A298 );
 a63989a <=( a63988a  and  a63985a );
 a63990a <=( a63989a  and  a63982a );
 a63994a <=( (not A168)  and  (not A169) );
 a63995a <=( (not A170)  and  a63994a );
 a63999a <=( A201  and  (not A200) );
 a64000a <=( A199  and  a63999a );
 a64001a <=( a64000a  and  a63995a );
 a64005a <=( A233  and  A232 );
 a64006a <=( A203  and  a64005a );
 a64009a <=( (not A266)  and  (not A265) );
 a64012a <=( (not A299)  and  (not A298) );
 a64013a <=( a64012a  and  a64009a );
 a64014a <=( a64013a  and  a64006a );
 a64018a <=( (not A168)  and  (not A169) );
 a64019a <=( (not A170)  and  a64018a );
 a64023a <=( A201  and  (not A200) );
 a64024a <=( A199  and  a64023a );
 a64025a <=( a64024a  and  a64019a );
 a64029a <=( A233  and  (not A232) );
 a64030a <=( A203  and  a64029a );
 a64033a <=( (not A299)  and  A298 );
 a64036a <=( A301  and  A300 );
 a64037a <=( a64036a  and  a64033a );
 a64038a <=( a64037a  and  a64030a );
 a64042a <=( (not A168)  and  (not A169) );
 a64043a <=( (not A170)  and  a64042a );
 a64047a <=( A201  and  (not A200) );
 a64048a <=( A199  and  a64047a );
 a64049a <=( a64048a  and  a64043a );
 a64053a <=( A233  and  (not A232) );
 a64054a <=( A203  and  a64053a );
 a64057a <=( (not A299)  and  A298 );
 a64060a <=( A302  and  A300 );
 a64061a <=( a64060a  and  a64057a );
 a64062a <=( a64061a  and  a64054a );
 a64066a <=( (not A168)  and  (not A169) );
 a64067a <=( (not A170)  and  a64066a );
 a64071a <=( A201  and  (not A200) );
 a64072a <=( A199  and  a64071a );
 a64073a <=( a64072a  and  a64067a );
 a64077a <=( A233  and  (not A232) );
 a64078a <=( A203  and  a64077a );
 a64081a <=( (not A266)  and  A265 );
 a64084a <=( A268  and  A267 );
 a64085a <=( a64084a  and  a64081a );
 a64086a <=( a64085a  and  a64078a );
 a64090a <=( (not A168)  and  (not A169) );
 a64091a <=( (not A170)  and  a64090a );
 a64095a <=( A201  and  (not A200) );
 a64096a <=( A199  and  a64095a );
 a64097a <=( a64096a  and  a64091a );
 a64101a <=( A233  and  (not A232) );
 a64102a <=( A203  and  a64101a );
 a64105a <=( (not A266)  and  A265 );
 a64108a <=( A269  and  A267 );
 a64109a <=( a64108a  and  a64105a );
 a64110a <=( a64109a  and  a64102a );
 a64114a <=( (not A168)  and  (not A169) );
 a64115a <=( (not A170)  and  a64114a );
 a64119a <=( A201  and  (not A200) );
 a64120a <=( A199  and  a64119a );
 a64121a <=( a64120a  and  a64115a );
 a64125a <=( (not A234)  and  (not A233) );
 a64126a <=( A203  and  a64125a );
 a64129a <=( A266  and  A265 );
 a64132a <=( (not A300)  and  A298 );
 a64133a <=( a64132a  and  a64129a );
 a64134a <=( a64133a  and  a64126a );
 a64138a <=( (not A168)  and  (not A169) );
 a64139a <=( (not A170)  and  a64138a );
 a64143a <=( A201  and  (not A200) );
 a64144a <=( A199  and  a64143a );
 a64145a <=( a64144a  and  a64139a );
 a64149a <=( (not A234)  and  (not A233) );
 a64150a <=( A203  and  a64149a );
 a64153a <=( A266  and  A265 );
 a64156a <=( A299  and  A298 );
 a64157a <=( a64156a  and  a64153a );
 a64158a <=( a64157a  and  a64150a );
 a64162a <=( (not A168)  and  (not A169) );
 a64163a <=( (not A170)  and  a64162a );
 a64167a <=( A201  and  (not A200) );
 a64168a <=( A199  and  a64167a );
 a64169a <=( a64168a  and  a64163a );
 a64173a <=( (not A234)  and  (not A233) );
 a64174a <=( A203  and  a64173a );
 a64177a <=( A266  and  A265 );
 a64180a <=( (not A299)  and  (not A298) );
 a64181a <=( a64180a  and  a64177a );
 a64182a <=( a64181a  and  a64174a );
 a64186a <=( (not A168)  and  (not A169) );
 a64187a <=( (not A170)  and  a64186a );
 a64191a <=( A201  and  (not A200) );
 a64192a <=( A199  and  a64191a );
 a64193a <=( a64192a  and  a64187a );
 a64197a <=( (not A234)  and  (not A233) );
 a64198a <=( A203  and  a64197a );
 a64201a <=( (not A267)  and  (not A266) );
 a64204a <=( (not A300)  and  A298 );
 a64205a <=( a64204a  and  a64201a );
 a64206a <=( a64205a  and  a64198a );
 a64210a <=( (not A168)  and  (not A169) );
 a64211a <=( (not A170)  and  a64210a );
 a64215a <=( A201  and  (not A200) );
 a64216a <=( A199  and  a64215a );
 a64217a <=( a64216a  and  a64211a );
 a64221a <=( (not A234)  and  (not A233) );
 a64222a <=( A203  and  a64221a );
 a64225a <=( (not A267)  and  (not A266) );
 a64228a <=( A299  and  A298 );
 a64229a <=( a64228a  and  a64225a );
 a64230a <=( a64229a  and  a64222a );
 a64234a <=( (not A168)  and  (not A169) );
 a64235a <=( (not A170)  and  a64234a );
 a64239a <=( A201  and  (not A200) );
 a64240a <=( A199  and  a64239a );
 a64241a <=( a64240a  and  a64235a );
 a64245a <=( (not A234)  and  (not A233) );
 a64246a <=( A203  and  a64245a );
 a64249a <=( (not A267)  and  (not A266) );
 a64252a <=( (not A299)  and  (not A298) );
 a64253a <=( a64252a  and  a64249a );
 a64254a <=( a64253a  and  a64246a );
 a64258a <=( (not A168)  and  (not A169) );
 a64259a <=( (not A170)  and  a64258a );
 a64263a <=( A201  and  (not A200) );
 a64264a <=( A199  and  a64263a );
 a64265a <=( a64264a  and  a64259a );
 a64269a <=( (not A234)  and  (not A233) );
 a64270a <=( A203  and  a64269a );
 a64273a <=( (not A266)  and  (not A265) );
 a64276a <=( (not A300)  and  A298 );
 a64277a <=( a64276a  and  a64273a );
 a64278a <=( a64277a  and  a64270a );
 a64282a <=( (not A168)  and  (not A169) );
 a64283a <=( (not A170)  and  a64282a );
 a64287a <=( A201  and  (not A200) );
 a64288a <=( A199  and  a64287a );
 a64289a <=( a64288a  and  a64283a );
 a64293a <=( (not A234)  and  (not A233) );
 a64294a <=( A203  and  a64293a );
 a64297a <=( (not A266)  and  (not A265) );
 a64300a <=( A299  and  A298 );
 a64301a <=( a64300a  and  a64297a );
 a64302a <=( a64301a  and  a64294a );
 a64306a <=( (not A168)  and  (not A169) );
 a64307a <=( (not A170)  and  a64306a );
 a64311a <=( A201  and  (not A200) );
 a64312a <=( A199  and  a64311a );
 a64313a <=( a64312a  and  a64307a );
 a64317a <=( (not A234)  and  (not A233) );
 a64318a <=( A203  and  a64317a );
 a64321a <=( (not A266)  and  (not A265) );
 a64324a <=( (not A299)  and  (not A298) );
 a64325a <=( a64324a  and  a64321a );
 a64326a <=( a64325a  and  a64318a );
 a64330a <=( (not A168)  and  (not A169) );
 a64331a <=( (not A170)  and  a64330a );
 a64335a <=( A201  and  (not A200) );
 a64336a <=( A199  and  a64335a );
 a64337a <=( a64336a  and  a64331a );
 a64341a <=( (not A233)  and  A232 );
 a64342a <=( A203  and  a64341a );
 a64345a <=( A235  and  A234 );
 a64348a <=( A299  and  (not A298) );
 a64349a <=( a64348a  and  a64345a );
 a64350a <=( a64349a  and  a64342a );
 a64354a <=( (not A168)  and  (not A169) );
 a64355a <=( (not A170)  and  a64354a );
 a64359a <=( A201  and  (not A200) );
 a64360a <=( A199  and  a64359a );
 a64361a <=( a64360a  and  a64355a );
 a64365a <=( (not A233)  and  A232 );
 a64366a <=( A203  and  a64365a );
 a64369a <=( A235  and  A234 );
 a64372a <=( A266  and  (not A265) );
 a64373a <=( a64372a  and  a64369a );
 a64374a <=( a64373a  and  a64366a );
 a64378a <=( (not A168)  and  (not A169) );
 a64379a <=( (not A170)  and  a64378a );
 a64383a <=( A201  and  (not A200) );
 a64384a <=( A199  and  a64383a );
 a64385a <=( a64384a  and  a64379a );
 a64389a <=( (not A233)  and  A232 );
 a64390a <=( A203  and  a64389a );
 a64393a <=( A236  and  A234 );
 a64396a <=( A299  and  (not A298) );
 a64397a <=( a64396a  and  a64393a );
 a64398a <=( a64397a  and  a64390a );
 a64402a <=( (not A168)  and  (not A169) );
 a64403a <=( (not A170)  and  a64402a );
 a64407a <=( A201  and  (not A200) );
 a64408a <=( A199  and  a64407a );
 a64409a <=( a64408a  and  a64403a );
 a64413a <=( (not A233)  and  A232 );
 a64414a <=( A203  and  a64413a );
 a64417a <=( A236  and  A234 );
 a64420a <=( A266  and  (not A265) );
 a64421a <=( a64420a  and  a64417a );
 a64422a <=( a64421a  and  a64414a );
 a64426a <=( (not A168)  and  (not A169) );
 a64427a <=( (not A170)  and  a64426a );
 a64431a <=( A201  and  (not A200) );
 a64432a <=( A199  and  a64431a );
 a64433a <=( a64432a  and  a64427a );
 a64437a <=( (not A233)  and  (not A232) );
 a64438a <=( A203  and  a64437a );
 a64441a <=( A266  and  A265 );
 a64444a <=( (not A300)  and  A298 );
 a64445a <=( a64444a  and  a64441a );
 a64446a <=( a64445a  and  a64438a );
 a64450a <=( (not A168)  and  (not A169) );
 a64451a <=( (not A170)  and  a64450a );
 a64455a <=( A201  and  (not A200) );
 a64456a <=( A199  and  a64455a );
 a64457a <=( a64456a  and  a64451a );
 a64461a <=( (not A233)  and  (not A232) );
 a64462a <=( A203  and  a64461a );
 a64465a <=( A266  and  A265 );
 a64468a <=( A299  and  A298 );
 a64469a <=( a64468a  and  a64465a );
 a64470a <=( a64469a  and  a64462a );
 a64474a <=( (not A168)  and  (not A169) );
 a64475a <=( (not A170)  and  a64474a );
 a64479a <=( A201  and  (not A200) );
 a64480a <=( A199  and  a64479a );
 a64481a <=( a64480a  and  a64475a );
 a64485a <=( (not A233)  and  (not A232) );
 a64486a <=( A203  and  a64485a );
 a64489a <=( A266  and  A265 );
 a64492a <=( (not A299)  and  (not A298) );
 a64493a <=( a64492a  and  a64489a );
 a64494a <=( a64493a  and  a64486a );
 a64498a <=( (not A168)  and  (not A169) );
 a64499a <=( (not A170)  and  a64498a );
 a64503a <=( A201  and  (not A200) );
 a64504a <=( A199  and  a64503a );
 a64505a <=( a64504a  and  a64499a );
 a64509a <=( (not A233)  and  (not A232) );
 a64510a <=( A203  and  a64509a );
 a64513a <=( (not A267)  and  (not A266) );
 a64516a <=( (not A300)  and  A298 );
 a64517a <=( a64516a  and  a64513a );
 a64518a <=( a64517a  and  a64510a );
 a64522a <=( (not A168)  and  (not A169) );
 a64523a <=( (not A170)  and  a64522a );
 a64527a <=( A201  and  (not A200) );
 a64528a <=( A199  and  a64527a );
 a64529a <=( a64528a  and  a64523a );
 a64533a <=( (not A233)  and  (not A232) );
 a64534a <=( A203  and  a64533a );
 a64537a <=( (not A267)  and  (not A266) );
 a64540a <=( A299  and  A298 );
 a64541a <=( a64540a  and  a64537a );
 a64542a <=( a64541a  and  a64534a );
 a64546a <=( (not A168)  and  (not A169) );
 a64547a <=( (not A170)  and  a64546a );
 a64551a <=( A201  and  (not A200) );
 a64552a <=( A199  and  a64551a );
 a64553a <=( a64552a  and  a64547a );
 a64557a <=( (not A233)  and  (not A232) );
 a64558a <=( A203  and  a64557a );
 a64561a <=( (not A267)  and  (not A266) );
 a64564a <=( (not A299)  and  (not A298) );
 a64565a <=( a64564a  and  a64561a );
 a64566a <=( a64565a  and  a64558a );
 a64570a <=( (not A168)  and  (not A169) );
 a64571a <=( (not A170)  and  a64570a );
 a64575a <=( A201  and  (not A200) );
 a64576a <=( A199  and  a64575a );
 a64577a <=( a64576a  and  a64571a );
 a64581a <=( (not A233)  and  (not A232) );
 a64582a <=( A203  and  a64581a );
 a64585a <=( (not A266)  and  (not A265) );
 a64588a <=( (not A300)  and  A298 );
 a64589a <=( a64588a  and  a64585a );
 a64590a <=( a64589a  and  a64582a );
 a64594a <=( (not A168)  and  (not A169) );
 a64595a <=( (not A170)  and  a64594a );
 a64599a <=( A201  and  (not A200) );
 a64600a <=( A199  and  a64599a );
 a64601a <=( a64600a  and  a64595a );
 a64605a <=( (not A233)  and  (not A232) );
 a64606a <=( A203  and  a64605a );
 a64609a <=( (not A266)  and  (not A265) );
 a64612a <=( A299  and  A298 );
 a64613a <=( a64612a  and  a64609a );
 a64614a <=( a64613a  and  a64606a );
 a64618a <=( (not A168)  and  (not A169) );
 a64619a <=( (not A170)  and  a64618a );
 a64623a <=( A201  and  (not A200) );
 a64624a <=( A199  and  a64623a );
 a64625a <=( a64624a  and  a64619a );
 a64629a <=( (not A233)  and  (not A232) );
 a64630a <=( A203  and  a64629a );
 a64633a <=( (not A266)  and  (not A265) );
 a64636a <=( (not A299)  and  (not A298) );
 a64637a <=( a64636a  and  a64633a );
 a64638a <=( a64637a  and  a64630a );
 a64642a <=( (not A200)  and  A166 );
 a64643a <=( A168  and  a64642a );
 a64646a <=( (not A203)  and  (not A202) );
 a64649a <=( (not A235)  and  (not A233) );
 a64650a <=( a64649a  and  a64646a );
 a64651a <=( a64650a  and  a64643a );
 a64655a <=( (not A268)  and  (not A266) );
 a64656a <=( (not A236)  and  a64655a );
 a64659a <=( A298  and  (not A269) );
 a64662a <=( (not A302)  and  (not A301) );
 a64663a <=( a64662a  and  a64659a );
 a64664a <=( a64663a  and  a64656a );
 a64668a <=( (not A200)  and  A167 );
 a64669a <=( A168  and  a64668a );
 a64672a <=( (not A203)  and  (not A202) );
 a64675a <=( (not A235)  and  (not A233) );
 a64676a <=( a64675a  and  a64672a );
 a64677a <=( a64676a  and  a64669a );
 a64681a <=( (not A268)  and  (not A266) );
 a64682a <=( (not A236)  and  a64681a );
 a64685a <=( A298  and  (not A269) );
 a64688a <=( (not A302)  and  (not A301) );
 a64689a <=( a64688a  and  a64685a );
 a64690a <=( a64689a  and  a64682a );
 a64694a <=( (not A166)  and  (not A167) );
 a64695a <=( A170  and  a64694a );
 a64698a <=( A200  and  (not A199) );
 a64701a <=( (not A235)  and  (not A233) );
 a64702a <=( a64701a  and  a64698a );
 a64703a <=( a64702a  and  a64695a );
 a64707a <=( (not A268)  and  (not A266) );
 a64708a <=( (not A236)  and  a64707a );
 a64711a <=( A298  and  (not A269) );
 a64714a <=( (not A302)  and  (not A301) );
 a64715a <=( a64714a  and  a64711a );
 a64716a <=( a64715a  and  a64708a );
 a64720a <=( (not A166)  and  (not A167) );
 a64721a <=( A170  and  a64720a );
 a64724a <=( (not A200)  and  A199 );
 a64727a <=( A202  and  A201 );
 a64728a <=( a64727a  and  a64724a );
 a64729a <=( a64728a  and  a64721a );
 a64733a <=( A265  and  A233 );
 a64734a <=( A232  and  a64733a );
 a64737a <=( (not A269)  and  (not A268) );
 a64740a <=( (not A300)  and  (not A299) );
 a64741a <=( a64740a  and  a64737a );
 a64742a <=( a64741a  and  a64734a );
 a64746a <=( (not A166)  and  (not A167) );
 a64747a <=( A170  and  a64746a );
 a64750a <=( (not A200)  and  A199 );
 a64753a <=( A202  and  A201 );
 a64754a <=( a64753a  and  a64750a );
 a64755a <=( a64754a  and  a64747a );
 a64759a <=( A265  and  A233 );
 a64760a <=( A232  and  a64759a );
 a64763a <=( (not A269)  and  (not A268) );
 a64766a <=( A299  and  A298 );
 a64767a <=( a64766a  and  a64763a );
 a64768a <=( a64767a  and  a64760a );
 a64772a <=( (not A166)  and  (not A167) );
 a64773a <=( A170  and  a64772a );
 a64776a <=( (not A200)  and  A199 );
 a64779a <=( A202  and  A201 );
 a64780a <=( a64779a  and  a64776a );
 a64781a <=( a64780a  and  a64773a );
 a64785a <=( A265  and  A233 );
 a64786a <=( A232  and  a64785a );
 a64789a <=( (not A269)  and  (not A268) );
 a64792a <=( (not A299)  and  (not A298) );
 a64793a <=( a64792a  and  a64789a );
 a64794a <=( a64793a  and  a64786a );
 a64798a <=( (not A166)  and  (not A167) );
 a64799a <=( A170  and  a64798a );
 a64802a <=( (not A200)  and  A199 );
 a64805a <=( A202  and  A201 );
 a64806a <=( a64805a  and  a64802a );
 a64807a <=( a64806a  and  a64799a );
 a64811a <=( A265  and  A233 );
 a64812a <=( A232  and  a64811a );
 a64815a <=( (not A299)  and  (not A267) );
 a64818a <=( (not A302)  and  (not A301) );
 a64819a <=( a64818a  and  a64815a );
 a64820a <=( a64819a  and  a64812a );
 a64824a <=( (not A166)  and  (not A167) );
 a64825a <=( A170  and  a64824a );
 a64828a <=( (not A200)  and  A199 );
 a64831a <=( A202  and  A201 );
 a64832a <=( a64831a  and  a64828a );
 a64833a <=( a64832a  and  a64825a );
 a64837a <=( A265  and  A233 );
 a64838a <=( A232  and  a64837a );
 a64841a <=( (not A299)  and  A266 );
 a64844a <=( (not A302)  and  (not A301) );
 a64845a <=( a64844a  and  a64841a );
 a64846a <=( a64845a  and  a64838a );
 a64850a <=( (not A166)  and  (not A167) );
 a64851a <=( A170  and  a64850a );
 a64854a <=( (not A200)  and  A199 );
 a64857a <=( A202  and  A201 );
 a64858a <=( a64857a  and  a64854a );
 a64859a <=( a64858a  and  a64851a );
 a64863a <=( (not A265)  and  A233 );
 a64864a <=( A232  and  a64863a );
 a64867a <=( (not A299)  and  (not A266) );
 a64870a <=( (not A302)  and  (not A301) );
 a64871a <=( a64870a  and  a64867a );
 a64872a <=( a64871a  and  a64864a );
 a64876a <=( (not A166)  and  (not A167) );
 a64877a <=( A170  and  a64876a );
 a64880a <=( (not A200)  and  A199 );
 a64883a <=( A202  and  A201 );
 a64884a <=( a64883a  and  a64880a );
 a64885a <=( a64884a  and  a64877a );
 a64889a <=( (not A236)  and  (not A235) );
 a64890a <=( (not A233)  and  a64889a );
 a64893a <=( A266  and  A265 );
 a64896a <=( (not A300)  and  A298 );
 a64897a <=( a64896a  and  a64893a );
 a64898a <=( a64897a  and  a64890a );
 a64902a <=( (not A166)  and  (not A167) );
 a64903a <=( A170  and  a64902a );
 a64906a <=( (not A200)  and  A199 );
 a64909a <=( A202  and  A201 );
 a64910a <=( a64909a  and  a64906a );
 a64911a <=( a64910a  and  a64903a );
 a64915a <=( (not A236)  and  (not A235) );
 a64916a <=( (not A233)  and  a64915a );
 a64919a <=( A266  and  A265 );
 a64922a <=( A299  and  A298 );
 a64923a <=( a64922a  and  a64919a );
 a64924a <=( a64923a  and  a64916a );
 a64928a <=( (not A166)  and  (not A167) );
 a64929a <=( A170  and  a64928a );
 a64932a <=( (not A200)  and  A199 );
 a64935a <=( A202  and  A201 );
 a64936a <=( a64935a  and  a64932a );
 a64937a <=( a64936a  and  a64929a );
 a64941a <=( (not A236)  and  (not A235) );
 a64942a <=( (not A233)  and  a64941a );
 a64945a <=( A266  and  A265 );
 a64948a <=( (not A299)  and  (not A298) );
 a64949a <=( a64948a  and  a64945a );
 a64950a <=( a64949a  and  a64942a );
 a64954a <=( (not A166)  and  (not A167) );
 a64955a <=( A170  and  a64954a );
 a64958a <=( (not A200)  and  A199 );
 a64961a <=( A202  and  A201 );
 a64962a <=( a64961a  and  a64958a );
 a64963a <=( a64962a  and  a64955a );
 a64967a <=( (not A236)  and  (not A235) );
 a64968a <=( (not A233)  and  a64967a );
 a64971a <=( (not A267)  and  (not A266) );
 a64974a <=( (not A300)  and  A298 );
 a64975a <=( a64974a  and  a64971a );
 a64976a <=( a64975a  and  a64968a );
 a64980a <=( (not A166)  and  (not A167) );
 a64981a <=( A170  and  a64980a );
 a64984a <=( (not A200)  and  A199 );
 a64987a <=( A202  and  A201 );
 a64988a <=( a64987a  and  a64984a );
 a64989a <=( a64988a  and  a64981a );
 a64993a <=( (not A236)  and  (not A235) );
 a64994a <=( (not A233)  and  a64993a );
 a64997a <=( (not A267)  and  (not A266) );
 a65000a <=( A299  and  A298 );
 a65001a <=( a65000a  and  a64997a );
 a65002a <=( a65001a  and  a64994a );
 a65006a <=( (not A166)  and  (not A167) );
 a65007a <=( A170  and  a65006a );
 a65010a <=( (not A200)  and  A199 );
 a65013a <=( A202  and  A201 );
 a65014a <=( a65013a  and  a65010a );
 a65015a <=( a65014a  and  a65007a );
 a65019a <=( (not A236)  and  (not A235) );
 a65020a <=( (not A233)  and  a65019a );
 a65023a <=( (not A267)  and  (not A266) );
 a65026a <=( (not A299)  and  (not A298) );
 a65027a <=( a65026a  and  a65023a );
 a65028a <=( a65027a  and  a65020a );
 a65032a <=( (not A166)  and  (not A167) );
 a65033a <=( A170  and  a65032a );
 a65036a <=( (not A200)  and  A199 );
 a65039a <=( A202  and  A201 );
 a65040a <=( a65039a  and  a65036a );
 a65041a <=( a65040a  and  a65033a );
 a65045a <=( (not A236)  and  (not A235) );
 a65046a <=( (not A233)  and  a65045a );
 a65049a <=( (not A266)  and  (not A265) );
 a65052a <=( (not A300)  and  A298 );
 a65053a <=( a65052a  and  a65049a );
 a65054a <=( a65053a  and  a65046a );
 a65058a <=( (not A166)  and  (not A167) );
 a65059a <=( A170  and  a65058a );
 a65062a <=( (not A200)  and  A199 );
 a65065a <=( A202  and  A201 );
 a65066a <=( a65065a  and  a65062a );
 a65067a <=( a65066a  and  a65059a );
 a65071a <=( (not A236)  and  (not A235) );
 a65072a <=( (not A233)  and  a65071a );
 a65075a <=( (not A266)  and  (not A265) );
 a65078a <=( A299  and  A298 );
 a65079a <=( a65078a  and  a65075a );
 a65080a <=( a65079a  and  a65072a );
 a65084a <=( (not A166)  and  (not A167) );
 a65085a <=( A170  and  a65084a );
 a65088a <=( (not A200)  and  A199 );
 a65091a <=( A202  and  A201 );
 a65092a <=( a65091a  and  a65088a );
 a65093a <=( a65092a  and  a65085a );
 a65097a <=( (not A236)  and  (not A235) );
 a65098a <=( (not A233)  and  a65097a );
 a65101a <=( (not A266)  and  (not A265) );
 a65104a <=( (not A299)  and  (not A298) );
 a65105a <=( a65104a  and  a65101a );
 a65106a <=( a65105a  and  a65098a );
 a65110a <=( (not A166)  and  (not A167) );
 a65111a <=( A170  and  a65110a );
 a65114a <=( (not A200)  and  A199 );
 a65117a <=( A202  and  A201 );
 a65118a <=( a65117a  and  a65114a );
 a65119a <=( a65118a  and  a65111a );
 a65123a <=( A265  and  (not A234) );
 a65124a <=( (not A233)  and  a65123a );
 a65127a <=( A298  and  A266 );
 a65130a <=( (not A302)  and  (not A301) );
 a65131a <=( a65130a  and  a65127a );
 a65132a <=( a65131a  and  a65124a );
 a65136a <=( (not A166)  and  (not A167) );
 a65137a <=( A170  and  a65136a );
 a65140a <=( (not A200)  and  A199 );
 a65143a <=( A202  and  A201 );
 a65144a <=( a65143a  and  a65140a );
 a65145a <=( a65144a  and  a65137a );
 a65149a <=( (not A266)  and  (not A234) );
 a65150a <=( (not A233)  and  a65149a );
 a65153a <=( (not A269)  and  (not A268) );
 a65156a <=( (not A300)  and  A298 );
 a65157a <=( a65156a  and  a65153a );
 a65158a <=( a65157a  and  a65150a );
 a65162a <=( (not A166)  and  (not A167) );
 a65163a <=( A170  and  a65162a );
 a65166a <=( (not A200)  and  A199 );
 a65169a <=( A202  and  A201 );
 a65170a <=( a65169a  and  a65166a );
 a65171a <=( a65170a  and  a65163a );
 a65175a <=( (not A266)  and  (not A234) );
 a65176a <=( (not A233)  and  a65175a );
 a65179a <=( (not A269)  and  (not A268) );
 a65182a <=( A299  and  A298 );
 a65183a <=( a65182a  and  a65179a );
 a65184a <=( a65183a  and  a65176a );
 a65188a <=( (not A166)  and  (not A167) );
 a65189a <=( A170  and  a65188a );
 a65192a <=( (not A200)  and  A199 );
 a65195a <=( A202  and  A201 );
 a65196a <=( a65195a  and  a65192a );
 a65197a <=( a65196a  and  a65189a );
 a65201a <=( (not A266)  and  (not A234) );
 a65202a <=( (not A233)  and  a65201a );
 a65205a <=( (not A269)  and  (not A268) );
 a65208a <=( (not A299)  and  (not A298) );
 a65209a <=( a65208a  and  a65205a );
 a65210a <=( a65209a  and  a65202a );
 a65214a <=( (not A166)  and  (not A167) );
 a65215a <=( A170  and  a65214a );
 a65218a <=( (not A200)  and  A199 );
 a65221a <=( A202  and  A201 );
 a65222a <=( a65221a  and  a65218a );
 a65223a <=( a65222a  and  a65215a );
 a65227a <=( (not A266)  and  (not A234) );
 a65228a <=( (not A233)  and  a65227a );
 a65231a <=( A298  and  (not A267) );
 a65234a <=( (not A302)  and  (not A301) );
 a65235a <=( a65234a  and  a65231a );
 a65236a <=( a65235a  and  a65228a );
 a65240a <=( (not A166)  and  (not A167) );
 a65241a <=( A170  and  a65240a );
 a65244a <=( (not A200)  and  A199 );
 a65247a <=( A202  and  A201 );
 a65248a <=( a65247a  and  a65244a );
 a65249a <=( a65248a  and  a65241a );
 a65253a <=( (not A265)  and  (not A234) );
 a65254a <=( (not A233)  and  a65253a );
 a65257a <=( A298  and  (not A266) );
 a65260a <=( (not A302)  and  (not A301) );
 a65261a <=( a65260a  and  a65257a );
 a65262a <=( a65261a  and  a65254a );
 a65266a <=( (not A166)  and  (not A167) );
 a65267a <=( A170  and  a65266a );
 a65270a <=( (not A200)  and  A199 );
 a65273a <=( A202  and  A201 );
 a65274a <=( a65273a  and  a65270a );
 a65275a <=( a65274a  and  a65267a );
 a65279a <=( A265  and  (not A233) );
 a65280a <=( (not A232)  and  a65279a );
 a65283a <=( A298  and  A266 );
 a65286a <=( (not A302)  and  (not A301) );
 a65287a <=( a65286a  and  a65283a );
 a65288a <=( a65287a  and  a65280a );
 a65292a <=( (not A166)  and  (not A167) );
 a65293a <=( A170  and  a65292a );
 a65296a <=( (not A200)  and  A199 );
 a65299a <=( A202  and  A201 );
 a65300a <=( a65299a  and  a65296a );
 a65301a <=( a65300a  and  a65293a );
 a65305a <=( (not A266)  and  (not A233) );
 a65306a <=( (not A232)  and  a65305a );
 a65309a <=( (not A269)  and  (not A268) );
 a65312a <=( (not A300)  and  A298 );
 a65313a <=( a65312a  and  a65309a );
 a65314a <=( a65313a  and  a65306a );
 a65318a <=( (not A166)  and  (not A167) );
 a65319a <=( A170  and  a65318a );
 a65322a <=( (not A200)  and  A199 );
 a65325a <=( A202  and  A201 );
 a65326a <=( a65325a  and  a65322a );
 a65327a <=( a65326a  and  a65319a );
 a65331a <=( (not A266)  and  (not A233) );
 a65332a <=( (not A232)  and  a65331a );
 a65335a <=( (not A269)  and  (not A268) );
 a65338a <=( A299  and  A298 );
 a65339a <=( a65338a  and  a65335a );
 a65340a <=( a65339a  and  a65332a );
 a65344a <=( (not A166)  and  (not A167) );
 a65345a <=( A170  and  a65344a );
 a65348a <=( (not A200)  and  A199 );
 a65351a <=( A202  and  A201 );
 a65352a <=( a65351a  and  a65348a );
 a65353a <=( a65352a  and  a65345a );
 a65357a <=( (not A266)  and  (not A233) );
 a65358a <=( (not A232)  and  a65357a );
 a65361a <=( (not A269)  and  (not A268) );
 a65364a <=( (not A299)  and  (not A298) );
 a65365a <=( a65364a  and  a65361a );
 a65366a <=( a65365a  and  a65358a );
 a65370a <=( (not A166)  and  (not A167) );
 a65371a <=( A170  and  a65370a );
 a65374a <=( (not A200)  and  A199 );
 a65377a <=( A202  and  A201 );
 a65378a <=( a65377a  and  a65374a );
 a65379a <=( a65378a  and  a65371a );
 a65383a <=( (not A266)  and  (not A233) );
 a65384a <=( (not A232)  and  a65383a );
 a65387a <=( A298  and  (not A267) );
 a65390a <=( (not A302)  and  (not A301) );
 a65391a <=( a65390a  and  a65387a );
 a65392a <=( a65391a  and  a65384a );
 a65396a <=( (not A166)  and  (not A167) );
 a65397a <=( A170  and  a65396a );
 a65400a <=( (not A200)  and  A199 );
 a65403a <=( A202  and  A201 );
 a65404a <=( a65403a  and  a65400a );
 a65405a <=( a65404a  and  a65397a );
 a65409a <=( (not A265)  and  (not A233) );
 a65410a <=( (not A232)  and  a65409a );
 a65413a <=( A298  and  (not A266) );
 a65416a <=( (not A302)  and  (not A301) );
 a65417a <=( a65416a  and  a65413a );
 a65418a <=( a65417a  and  a65410a );
 a65422a <=( (not A166)  and  (not A167) );
 a65423a <=( A170  and  a65422a );
 a65426a <=( (not A200)  and  A199 );
 a65429a <=( A203  and  A201 );
 a65430a <=( a65429a  and  a65426a );
 a65431a <=( a65430a  and  a65423a );
 a65435a <=( A265  and  A233 );
 a65436a <=( A232  and  a65435a );
 a65439a <=( (not A269)  and  (not A268) );
 a65442a <=( (not A300)  and  (not A299) );
 a65443a <=( a65442a  and  a65439a );
 a65444a <=( a65443a  and  a65436a );
 a65448a <=( (not A166)  and  (not A167) );
 a65449a <=( A170  and  a65448a );
 a65452a <=( (not A200)  and  A199 );
 a65455a <=( A203  and  A201 );
 a65456a <=( a65455a  and  a65452a );
 a65457a <=( a65456a  and  a65449a );
 a65461a <=( A265  and  A233 );
 a65462a <=( A232  and  a65461a );
 a65465a <=( (not A269)  and  (not A268) );
 a65468a <=( A299  and  A298 );
 a65469a <=( a65468a  and  a65465a );
 a65470a <=( a65469a  and  a65462a );
 a65474a <=( (not A166)  and  (not A167) );
 a65475a <=( A170  and  a65474a );
 a65478a <=( (not A200)  and  A199 );
 a65481a <=( A203  and  A201 );
 a65482a <=( a65481a  and  a65478a );
 a65483a <=( a65482a  and  a65475a );
 a65487a <=( A265  and  A233 );
 a65488a <=( A232  and  a65487a );
 a65491a <=( (not A269)  and  (not A268) );
 a65494a <=( (not A299)  and  (not A298) );
 a65495a <=( a65494a  and  a65491a );
 a65496a <=( a65495a  and  a65488a );
 a65500a <=( (not A166)  and  (not A167) );
 a65501a <=( A170  and  a65500a );
 a65504a <=( (not A200)  and  A199 );
 a65507a <=( A203  and  A201 );
 a65508a <=( a65507a  and  a65504a );
 a65509a <=( a65508a  and  a65501a );
 a65513a <=( A265  and  A233 );
 a65514a <=( A232  and  a65513a );
 a65517a <=( (not A299)  and  (not A267) );
 a65520a <=( (not A302)  and  (not A301) );
 a65521a <=( a65520a  and  a65517a );
 a65522a <=( a65521a  and  a65514a );
 a65526a <=( (not A166)  and  (not A167) );
 a65527a <=( A170  and  a65526a );
 a65530a <=( (not A200)  and  A199 );
 a65533a <=( A203  and  A201 );
 a65534a <=( a65533a  and  a65530a );
 a65535a <=( a65534a  and  a65527a );
 a65539a <=( A265  and  A233 );
 a65540a <=( A232  and  a65539a );
 a65543a <=( (not A299)  and  A266 );
 a65546a <=( (not A302)  and  (not A301) );
 a65547a <=( a65546a  and  a65543a );
 a65548a <=( a65547a  and  a65540a );
 a65552a <=( (not A166)  and  (not A167) );
 a65553a <=( A170  and  a65552a );
 a65556a <=( (not A200)  and  A199 );
 a65559a <=( A203  and  A201 );
 a65560a <=( a65559a  and  a65556a );
 a65561a <=( a65560a  and  a65553a );
 a65565a <=( (not A265)  and  A233 );
 a65566a <=( A232  and  a65565a );
 a65569a <=( (not A299)  and  (not A266) );
 a65572a <=( (not A302)  and  (not A301) );
 a65573a <=( a65572a  and  a65569a );
 a65574a <=( a65573a  and  a65566a );
 a65578a <=( (not A166)  and  (not A167) );
 a65579a <=( A170  and  a65578a );
 a65582a <=( (not A200)  and  A199 );
 a65585a <=( A203  and  A201 );
 a65586a <=( a65585a  and  a65582a );
 a65587a <=( a65586a  and  a65579a );
 a65591a <=( (not A236)  and  (not A235) );
 a65592a <=( (not A233)  and  a65591a );
 a65595a <=( A266  and  A265 );
 a65598a <=( (not A300)  and  A298 );
 a65599a <=( a65598a  and  a65595a );
 a65600a <=( a65599a  and  a65592a );
 a65604a <=( (not A166)  and  (not A167) );
 a65605a <=( A170  and  a65604a );
 a65608a <=( (not A200)  and  A199 );
 a65611a <=( A203  and  A201 );
 a65612a <=( a65611a  and  a65608a );
 a65613a <=( a65612a  and  a65605a );
 a65617a <=( (not A236)  and  (not A235) );
 a65618a <=( (not A233)  and  a65617a );
 a65621a <=( A266  and  A265 );
 a65624a <=( A299  and  A298 );
 a65625a <=( a65624a  and  a65621a );
 a65626a <=( a65625a  and  a65618a );
 a65630a <=( (not A166)  and  (not A167) );
 a65631a <=( A170  and  a65630a );
 a65634a <=( (not A200)  and  A199 );
 a65637a <=( A203  and  A201 );
 a65638a <=( a65637a  and  a65634a );
 a65639a <=( a65638a  and  a65631a );
 a65643a <=( (not A236)  and  (not A235) );
 a65644a <=( (not A233)  and  a65643a );
 a65647a <=( A266  and  A265 );
 a65650a <=( (not A299)  and  (not A298) );
 a65651a <=( a65650a  and  a65647a );
 a65652a <=( a65651a  and  a65644a );
 a65656a <=( (not A166)  and  (not A167) );
 a65657a <=( A170  and  a65656a );
 a65660a <=( (not A200)  and  A199 );
 a65663a <=( A203  and  A201 );
 a65664a <=( a65663a  and  a65660a );
 a65665a <=( a65664a  and  a65657a );
 a65669a <=( (not A236)  and  (not A235) );
 a65670a <=( (not A233)  and  a65669a );
 a65673a <=( (not A267)  and  (not A266) );
 a65676a <=( (not A300)  and  A298 );
 a65677a <=( a65676a  and  a65673a );
 a65678a <=( a65677a  and  a65670a );
 a65682a <=( (not A166)  and  (not A167) );
 a65683a <=( A170  and  a65682a );
 a65686a <=( (not A200)  and  A199 );
 a65689a <=( A203  and  A201 );
 a65690a <=( a65689a  and  a65686a );
 a65691a <=( a65690a  and  a65683a );
 a65695a <=( (not A236)  and  (not A235) );
 a65696a <=( (not A233)  and  a65695a );
 a65699a <=( (not A267)  and  (not A266) );
 a65702a <=( A299  and  A298 );
 a65703a <=( a65702a  and  a65699a );
 a65704a <=( a65703a  and  a65696a );
 a65708a <=( (not A166)  and  (not A167) );
 a65709a <=( A170  and  a65708a );
 a65712a <=( (not A200)  and  A199 );
 a65715a <=( A203  and  A201 );
 a65716a <=( a65715a  and  a65712a );
 a65717a <=( a65716a  and  a65709a );
 a65721a <=( (not A236)  and  (not A235) );
 a65722a <=( (not A233)  and  a65721a );
 a65725a <=( (not A267)  and  (not A266) );
 a65728a <=( (not A299)  and  (not A298) );
 a65729a <=( a65728a  and  a65725a );
 a65730a <=( a65729a  and  a65722a );
 a65734a <=( (not A166)  and  (not A167) );
 a65735a <=( A170  and  a65734a );
 a65738a <=( (not A200)  and  A199 );
 a65741a <=( A203  and  A201 );
 a65742a <=( a65741a  and  a65738a );
 a65743a <=( a65742a  and  a65735a );
 a65747a <=( (not A236)  and  (not A235) );
 a65748a <=( (not A233)  and  a65747a );
 a65751a <=( (not A266)  and  (not A265) );
 a65754a <=( (not A300)  and  A298 );
 a65755a <=( a65754a  and  a65751a );
 a65756a <=( a65755a  and  a65748a );
 a65760a <=( (not A166)  and  (not A167) );
 a65761a <=( A170  and  a65760a );
 a65764a <=( (not A200)  and  A199 );
 a65767a <=( A203  and  A201 );
 a65768a <=( a65767a  and  a65764a );
 a65769a <=( a65768a  and  a65761a );
 a65773a <=( (not A236)  and  (not A235) );
 a65774a <=( (not A233)  and  a65773a );
 a65777a <=( (not A266)  and  (not A265) );
 a65780a <=( A299  and  A298 );
 a65781a <=( a65780a  and  a65777a );
 a65782a <=( a65781a  and  a65774a );
 a65786a <=( (not A166)  and  (not A167) );
 a65787a <=( A170  and  a65786a );
 a65790a <=( (not A200)  and  A199 );
 a65793a <=( A203  and  A201 );
 a65794a <=( a65793a  and  a65790a );
 a65795a <=( a65794a  and  a65787a );
 a65799a <=( (not A236)  and  (not A235) );
 a65800a <=( (not A233)  and  a65799a );
 a65803a <=( (not A266)  and  (not A265) );
 a65806a <=( (not A299)  and  (not A298) );
 a65807a <=( a65806a  and  a65803a );
 a65808a <=( a65807a  and  a65800a );
 a65812a <=( (not A166)  and  (not A167) );
 a65813a <=( A170  and  a65812a );
 a65816a <=( (not A200)  and  A199 );
 a65819a <=( A203  and  A201 );
 a65820a <=( a65819a  and  a65816a );
 a65821a <=( a65820a  and  a65813a );
 a65825a <=( A265  and  (not A234) );
 a65826a <=( (not A233)  and  a65825a );
 a65829a <=( A298  and  A266 );
 a65832a <=( (not A302)  and  (not A301) );
 a65833a <=( a65832a  and  a65829a );
 a65834a <=( a65833a  and  a65826a );
 a65838a <=( (not A166)  and  (not A167) );
 a65839a <=( A170  and  a65838a );
 a65842a <=( (not A200)  and  A199 );
 a65845a <=( A203  and  A201 );
 a65846a <=( a65845a  and  a65842a );
 a65847a <=( a65846a  and  a65839a );
 a65851a <=( (not A266)  and  (not A234) );
 a65852a <=( (not A233)  and  a65851a );
 a65855a <=( (not A269)  and  (not A268) );
 a65858a <=( (not A300)  and  A298 );
 a65859a <=( a65858a  and  a65855a );
 a65860a <=( a65859a  and  a65852a );
 a65864a <=( (not A166)  and  (not A167) );
 a65865a <=( A170  and  a65864a );
 a65868a <=( (not A200)  and  A199 );
 a65871a <=( A203  and  A201 );
 a65872a <=( a65871a  and  a65868a );
 a65873a <=( a65872a  and  a65865a );
 a65877a <=( (not A266)  and  (not A234) );
 a65878a <=( (not A233)  and  a65877a );
 a65881a <=( (not A269)  and  (not A268) );
 a65884a <=( A299  and  A298 );
 a65885a <=( a65884a  and  a65881a );
 a65886a <=( a65885a  and  a65878a );
 a65890a <=( (not A166)  and  (not A167) );
 a65891a <=( A170  and  a65890a );
 a65894a <=( (not A200)  and  A199 );
 a65897a <=( A203  and  A201 );
 a65898a <=( a65897a  and  a65894a );
 a65899a <=( a65898a  and  a65891a );
 a65903a <=( (not A266)  and  (not A234) );
 a65904a <=( (not A233)  and  a65903a );
 a65907a <=( (not A269)  and  (not A268) );
 a65910a <=( (not A299)  and  (not A298) );
 a65911a <=( a65910a  and  a65907a );
 a65912a <=( a65911a  and  a65904a );
 a65916a <=( (not A166)  and  (not A167) );
 a65917a <=( A170  and  a65916a );
 a65920a <=( (not A200)  and  A199 );
 a65923a <=( A203  and  A201 );
 a65924a <=( a65923a  and  a65920a );
 a65925a <=( a65924a  and  a65917a );
 a65929a <=( (not A266)  and  (not A234) );
 a65930a <=( (not A233)  and  a65929a );
 a65933a <=( A298  and  (not A267) );
 a65936a <=( (not A302)  and  (not A301) );
 a65937a <=( a65936a  and  a65933a );
 a65938a <=( a65937a  and  a65930a );
 a65942a <=( (not A166)  and  (not A167) );
 a65943a <=( A170  and  a65942a );
 a65946a <=( (not A200)  and  A199 );
 a65949a <=( A203  and  A201 );
 a65950a <=( a65949a  and  a65946a );
 a65951a <=( a65950a  and  a65943a );
 a65955a <=( (not A265)  and  (not A234) );
 a65956a <=( (not A233)  and  a65955a );
 a65959a <=( A298  and  (not A266) );
 a65962a <=( (not A302)  and  (not A301) );
 a65963a <=( a65962a  and  a65959a );
 a65964a <=( a65963a  and  a65956a );
 a65968a <=( (not A166)  and  (not A167) );
 a65969a <=( A170  and  a65968a );
 a65972a <=( (not A200)  and  A199 );
 a65975a <=( A203  and  A201 );
 a65976a <=( a65975a  and  a65972a );
 a65977a <=( a65976a  and  a65969a );
 a65981a <=( A265  and  (not A233) );
 a65982a <=( (not A232)  and  a65981a );
 a65985a <=( A298  and  A266 );
 a65988a <=( (not A302)  and  (not A301) );
 a65989a <=( a65988a  and  a65985a );
 a65990a <=( a65989a  and  a65982a );
 a65994a <=( (not A166)  and  (not A167) );
 a65995a <=( A170  and  a65994a );
 a65998a <=( (not A200)  and  A199 );
 a66001a <=( A203  and  A201 );
 a66002a <=( a66001a  and  a65998a );
 a66003a <=( a66002a  and  a65995a );
 a66007a <=( (not A266)  and  (not A233) );
 a66008a <=( (not A232)  and  a66007a );
 a66011a <=( (not A269)  and  (not A268) );
 a66014a <=( (not A300)  and  A298 );
 a66015a <=( a66014a  and  a66011a );
 a66016a <=( a66015a  and  a66008a );
 a66020a <=( (not A166)  and  (not A167) );
 a66021a <=( A170  and  a66020a );
 a66024a <=( (not A200)  and  A199 );
 a66027a <=( A203  and  A201 );
 a66028a <=( a66027a  and  a66024a );
 a66029a <=( a66028a  and  a66021a );
 a66033a <=( (not A266)  and  (not A233) );
 a66034a <=( (not A232)  and  a66033a );
 a66037a <=( (not A269)  and  (not A268) );
 a66040a <=( A299  and  A298 );
 a66041a <=( a66040a  and  a66037a );
 a66042a <=( a66041a  and  a66034a );
 a66046a <=( (not A166)  and  (not A167) );
 a66047a <=( A170  and  a66046a );
 a66050a <=( (not A200)  and  A199 );
 a66053a <=( A203  and  A201 );
 a66054a <=( a66053a  and  a66050a );
 a66055a <=( a66054a  and  a66047a );
 a66059a <=( (not A266)  and  (not A233) );
 a66060a <=( (not A232)  and  a66059a );
 a66063a <=( (not A269)  and  (not A268) );
 a66066a <=( (not A299)  and  (not A298) );
 a66067a <=( a66066a  and  a66063a );
 a66068a <=( a66067a  and  a66060a );
 a66072a <=( (not A166)  and  (not A167) );
 a66073a <=( A170  and  a66072a );
 a66076a <=( (not A200)  and  A199 );
 a66079a <=( A203  and  A201 );
 a66080a <=( a66079a  and  a66076a );
 a66081a <=( a66080a  and  a66073a );
 a66085a <=( (not A266)  and  (not A233) );
 a66086a <=( (not A232)  and  a66085a );
 a66089a <=( A298  and  (not A267) );
 a66092a <=( (not A302)  and  (not A301) );
 a66093a <=( a66092a  and  a66089a );
 a66094a <=( a66093a  and  a66086a );
 a66098a <=( (not A166)  and  (not A167) );
 a66099a <=( A170  and  a66098a );
 a66102a <=( (not A200)  and  A199 );
 a66105a <=( A203  and  A201 );
 a66106a <=( a66105a  and  a66102a );
 a66107a <=( a66106a  and  a66099a );
 a66111a <=( (not A265)  and  (not A233) );
 a66112a <=( (not A232)  and  a66111a );
 a66115a <=( A298  and  (not A266) );
 a66118a <=( (not A302)  and  (not A301) );
 a66119a <=( a66118a  and  a66115a );
 a66120a <=( a66119a  and  a66112a );
 a66124a <=( A167  and  (not A168) );
 a66125a <=( A170  and  a66124a );
 a66128a <=( (not A199)  and  A166 );
 a66131a <=( A232  and  A200 );
 a66132a <=( a66131a  and  a66128a );
 a66133a <=( a66132a  and  a66125a );
 a66137a <=( (not A268)  and  A265 );
 a66138a <=( A233  and  a66137a );
 a66141a <=( (not A299)  and  (not A269) );
 a66144a <=( (not A302)  and  (not A301) );
 a66145a <=( a66144a  and  a66141a );
 a66146a <=( a66145a  and  a66138a );
 a66150a <=( A167  and  (not A168) );
 a66151a <=( A170  and  a66150a );
 a66154a <=( (not A199)  and  A166 );
 a66157a <=( (not A233)  and  A200 );
 a66158a <=( a66157a  and  a66154a );
 a66159a <=( a66158a  and  a66151a );
 a66163a <=( A265  and  (not A236) );
 a66164a <=( (not A235)  and  a66163a );
 a66167a <=( A298  and  A266 );
 a66170a <=( (not A302)  and  (not A301) );
 a66171a <=( a66170a  and  a66167a );
 a66172a <=( a66171a  and  a66164a );
 a66176a <=( A167  and  (not A168) );
 a66177a <=( A170  and  a66176a );
 a66180a <=( (not A199)  and  A166 );
 a66183a <=( (not A233)  and  A200 );
 a66184a <=( a66183a  and  a66180a );
 a66185a <=( a66184a  and  a66177a );
 a66189a <=( (not A266)  and  (not A236) );
 a66190a <=( (not A235)  and  a66189a );
 a66193a <=( (not A269)  and  (not A268) );
 a66196a <=( (not A300)  and  A298 );
 a66197a <=( a66196a  and  a66193a );
 a66198a <=( a66197a  and  a66190a );
 a66202a <=( A167  and  (not A168) );
 a66203a <=( A170  and  a66202a );
 a66206a <=( (not A199)  and  A166 );
 a66209a <=( (not A233)  and  A200 );
 a66210a <=( a66209a  and  a66206a );
 a66211a <=( a66210a  and  a66203a );
 a66215a <=( (not A266)  and  (not A236) );
 a66216a <=( (not A235)  and  a66215a );
 a66219a <=( (not A269)  and  (not A268) );
 a66222a <=( A299  and  A298 );
 a66223a <=( a66222a  and  a66219a );
 a66224a <=( a66223a  and  a66216a );
 a66228a <=( A167  and  (not A168) );
 a66229a <=( A170  and  a66228a );
 a66232a <=( (not A199)  and  A166 );
 a66235a <=( (not A233)  and  A200 );
 a66236a <=( a66235a  and  a66232a );
 a66237a <=( a66236a  and  a66229a );
 a66241a <=( (not A266)  and  (not A236) );
 a66242a <=( (not A235)  and  a66241a );
 a66245a <=( (not A269)  and  (not A268) );
 a66248a <=( (not A299)  and  (not A298) );
 a66249a <=( a66248a  and  a66245a );
 a66250a <=( a66249a  and  a66242a );
 a66254a <=( A167  and  (not A168) );
 a66255a <=( A170  and  a66254a );
 a66258a <=( (not A199)  and  A166 );
 a66261a <=( (not A233)  and  A200 );
 a66262a <=( a66261a  and  a66258a );
 a66263a <=( a66262a  and  a66255a );
 a66267a <=( (not A266)  and  (not A236) );
 a66268a <=( (not A235)  and  a66267a );
 a66271a <=( A298  and  (not A267) );
 a66274a <=( (not A302)  and  (not A301) );
 a66275a <=( a66274a  and  a66271a );
 a66276a <=( a66275a  and  a66268a );
 a66280a <=( A167  and  (not A168) );
 a66281a <=( A170  and  a66280a );
 a66284a <=( (not A199)  and  A166 );
 a66287a <=( (not A233)  and  A200 );
 a66288a <=( a66287a  and  a66284a );
 a66289a <=( a66288a  and  a66281a );
 a66293a <=( (not A265)  and  (not A236) );
 a66294a <=( (not A235)  and  a66293a );
 a66297a <=( A298  and  (not A266) );
 a66300a <=( (not A302)  and  (not A301) );
 a66301a <=( a66300a  and  a66297a );
 a66302a <=( a66301a  and  a66294a );
 a66306a <=( A167  and  (not A168) );
 a66307a <=( A170  and  a66306a );
 a66310a <=( (not A199)  and  A166 );
 a66313a <=( (not A233)  and  A200 );
 a66314a <=( a66313a  and  a66310a );
 a66315a <=( a66314a  and  a66307a );
 a66319a <=( (not A268)  and  (not A266) );
 a66320a <=( (not A234)  and  a66319a );
 a66323a <=( A298  and  (not A269) );
 a66326a <=( (not A302)  and  (not A301) );
 a66327a <=( a66326a  and  a66323a );
 a66328a <=( a66327a  and  a66320a );
 a66332a <=( A167  and  (not A168) );
 a66333a <=( A170  and  a66332a );
 a66336a <=( (not A199)  and  A166 );
 a66339a <=( A232  and  A200 );
 a66340a <=( a66339a  and  a66336a );
 a66341a <=( a66340a  and  a66333a );
 a66345a <=( A235  and  A234 );
 a66346a <=( (not A233)  and  a66345a );
 a66349a <=( (not A299)  and  A298 );
 a66352a <=( A301  and  A300 );
 a66353a <=( a66352a  and  a66349a );
 a66354a <=( a66353a  and  a66346a );
 a66358a <=( A167  and  (not A168) );
 a66359a <=( A170  and  a66358a );
 a66362a <=( (not A199)  and  A166 );
 a66365a <=( A232  and  A200 );
 a66366a <=( a66365a  and  a66362a );
 a66367a <=( a66366a  and  a66359a );
 a66371a <=( A235  and  A234 );
 a66372a <=( (not A233)  and  a66371a );
 a66375a <=( (not A299)  and  A298 );
 a66378a <=( A302  and  A300 );
 a66379a <=( a66378a  and  a66375a );
 a66380a <=( a66379a  and  a66372a );
 a66384a <=( A167  and  (not A168) );
 a66385a <=( A170  and  a66384a );
 a66388a <=( (not A199)  and  A166 );
 a66391a <=( A232  and  A200 );
 a66392a <=( a66391a  and  a66388a );
 a66393a <=( a66392a  and  a66385a );
 a66397a <=( A235  and  A234 );
 a66398a <=( (not A233)  and  a66397a );
 a66401a <=( (not A266)  and  A265 );
 a66404a <=( A268  and  A267 );
 a66405a <=( a66404a  and  a66401a );
 a66406a <=( a66405a  and  a66398a );
 a66410a <=( A167  and  (not A168) );
 a66411a <=( A170  and  a66410a );
 a66414a <=( (not A199)  and  A166 );
 a66417a <=( A232  and  A200 );
 a66418a <=( a66417a  and  a66414a );
 a66419a <=( a66418a  and  a66411a );
 a66423a <=( A235  and  A234 );
 a66424a <=( (not A233)  and  a66423a );
 a66427a <=( (not A266)  and  A265 );
 a66430a <=( A269  and  A267 );
 a66431a <=( a66430a  and  a66427a );
 a66432a <=( a66431a  and  a66424a );
 a66436a <=( A167  and  (not A168) );
 a66437a <=( A170  and  a66436a );
 a66440a <=( (not A199)  and  A166 );
 a66443a <=( A232  and  A200 );
 a66444a <=( a66443a  and  a66440a );
 a66445a <=( a66444a  and  a66437a );
 a66449a <=( A236  and  A234 );
 a66450a <=( (not A233)  and  a66449a );
 a66453a <=( (not A299)  and  A298 );
 a66456a <=( A301  and  A300 );
 a66457a <=( a66456a  and  a66453a );
 a66458a <=( a66457a  and  a66450a );
 a66462a <=( A167  and  (not A168) );
 a66463a <=( A170  and  a66462a );
 a66466a <=( (not A199)  and  A166 );
 a66469a <=( A232  and  A200 );
 a66470a <=( a66469a  and  a66466a );
 a66471a <=( a66470a  and  a66463a );
 a66475a <=( A236  and  A234 );
 a66476a <=( (not A233)  and  a66475a );
 a66479a <=( (not A299)  and  A298 );
 a66482a <=( A302  and  A300 );
 a66483a <=( a66482a  and  a66479a );
 a66484a <=( a66483a  and  a66476a );
 a66488a <=( A167  and  (not A168) );
 a66489a <=( A170  and  a66488a );
 a66492a <=( (not A199)  and  A166 );
 a66495a <=( A232  and  A200 );
 a66496a <=( a66495a  and  a66492a );
 a66497a <=( a66496a  and  a66489a );
 a66501a <=( A236  and  A234 );
 a66502a <=( (not A233)  and  a66501a );
 a66505a <=( (not A266)  and  A265 );
 a66508a <=( A268  and  A267 );
 a66509a <=( a66508a  and  a66505a );
 a66510a <=( a66509a  and  a66502a );
 a66514a <=( A167  and  (not A168) );
 a66515a <=( A170  and  a66514a );
 a66518a <=( (not A199)  and  A166 );
 a66521a <=( A232  and  A200 );
 a66522a <=( a66521a  and  a66518a );
 a66523a <=( a66522a  and  a66515a );
 a66527a <=( A236  and  A234 );
 a66528a <=( (not A233)  and  a66527a );
 a66531a <=( (not A266)  and  A265 );
 a66534a <=( A269  and  A267 );
 a66535a <=( a66534a  and  a66531a );
 a66536a <=( a66535a  and  a66528a );
 a66540a <=( A167  and  (not A168) );
 a66541a <=( A170  and  a66540a );
 a66544a <=( (not A199)  and  A166 );
 a66547a <=( (not A232)  and  A200 );
 a66548a <=( a66547a  and  a66544a );
 a66549a <=( a66548a  and  a66541a );
 a66553a <=( (not A268)  and  (not A266) );
 a66554a <=( (not A233)  and  a66553a );
 a66557a <=( A298  and  (not A269) );
 a66560a <=( (not A302)  and  (not A301) );
 a66561a <=( a66560a  and  a66557a );
 a66562a <=( a66561a  and  a66554a );
 a66566a <=( A167  and  (not A168) );
 a66567a <=( (not A170)  and  a66566a );
 a66570a <=( (not A199)  and  (not A166) );
 a66573a <=( A232  and  A200 );
 a66574a <=( a66573a  and  a66570a );
 a66575a <=( a66574a  and  a66567a );
 a66579a <=( (not A268)  and  A265 );
 a66580a <=( A233  and  a66579a );
 a66583a <=( (not A299)  and  (not A269) );
 a66586a <=( (not A302)  and  (not A301) );
 a66587a <=( a66586a  and  a66583a );
 a66588a <=( a66587a  and  a66580a );
 a66592a <=( A167  and  (not A168) );
 a66593a <=( (not A170)  and  a66592a );
 a66596a <=( (not A199)  and  (not A166) );
 a66599a <=( (not A233)  and  A200 );
 a66600a <=( a66599a  and  a66596a );
 a66601a <=( a66600a  and  a66593a );
 a66605a <=( A265  and  (not A236) );
 a66606a <=( (not A235)  and  a66605a );
 a66609a <=( A298  and  A266 );
 a66612a <=( (not A302)  and  (not A301) );
 a66613a <=( a66612a  and  a66609a );
 a66614a <=( a66613a  and  a66606a );
 a66618a <=( A167  and  (not A168) );
 a66619a <=( (not A170)  and  a66618a );
 a66622a <=( (not A199)  and  (not A166) );
 a66625a <=( (not A233)  and  A200 );
 a66626a <=( a66625a  and  a66622a );
 a66627a <=( a66626a  and  a66619a );
 a66631a <=( (not A266)  and  (not A236) );
 a66632a <=( (not A235)  and  a66631a );
 a66635a <=( (not A269)  and  (not A268) );
 a66638a <=( (not A300)  and  A298 );
 a66639a <=( a66638a  and  a66635a );
 a66640a <=( a66639a  and  a66632a );
 a66644a <=( A167  and  (not A168) );
 a66645a <=( (not A170)  and  a66644a );
 a66648a <=( (not A199)  and  (not A166) );
 a66651a <=( (not A233)  and  A200 );
 a66652a <=( a66651a  and  a66648a );
 a66653a <=( a66652a  and  a66645a );
 a66657a <=( (not A266)  and  (not A236) );
 a66658a <=( (not A235)  and  a66657a );
 a66661a <=( (not A269)  and  (not A268) );
 a66664a <=( A299  and  A298 );
 a66665a <=( a66664a  and  a66661a );
 a66666a <=( a66665a  and  a66658a );
 a66670a <=( A167  and  (not A168) );
 a66671a <=( (not A170)  and  a66670a );
 a66674a <=( (not A199)  and  (not A166) );
 a66677a <=( (not A233)  and  A200 );
 a66678a <=( a66677a  and  a66674a );
 a66679a <=( a66678a  and  a66671a );
 a66683a <=( (not A266)  and  (not A236) );
 a66684a <=( (not A235)  and  a66683a );
 a66687a <=( (not A269)  and  (not A268) );
 a66690a <=( (not A299)  and  (not A298) );
 a66691a <=( a66690a  and  a66687a );
 a66692a <=( a66691a  and  a66684a );
 a66696a <=( A167  and  (not A168) );
 a66697a <=( (not A170)  and  a66696a );
 a66700a <=( (not A199)  and  (not A166) );
 a66703a <=( (not A233)  and  A200 );
 a66704a <=( a66703a  and  a66700a );
 a66705a <=( a66704a  and  a66697a );
 a66709a <=( (not A266)  and  (not A236) );
 a66710a <=( (not A235)  and  a66709a );
 a66713a <=( A298  and  (not A267) );
 a66716a <=( (not A302)  and  (not A301) );
 a66717a <=( a66716a  and  a66713a );
 a66718a <=( a66717a  and  a66710a );
 a66722a <=( A167  and  (not A168) );
 a66723a <=( (not A170)  and  a66722a );
 a66726a <=( (not A199)  and  (not A166) );
 a66729a <=( (not A233)  and  A200 );
 a66730a <=( a66729a  and  a66726a );
 a66731a <=( a66730a  and  a66723a );
 a66735a <=( (not A265)  and  (not A236) );
 a66736a <=( (not A235)  and  a66735a );
 a66739a <=( A298  and  (not A266) );
 a66742a <=( (not A302)  and  (not A301) );
 a66743a <=( a66742a  and  a66739a );
 a66744a <=( a66743a  and  a66736a );
 a66748a <=( A167  and  (not A168) );
 a66749a <=( (not A170)  and  a66748a );
 a66752a <=( (not A199)  and  (not A166) );
 a66755a <=( (not A233)  and  A200 );
 a66756a <=( a66755a  and  a66752a );
 a66757a <=( a66756a  and  a66749a );
 a66761a <=( (not A268)  and  (not A266) );
 a66762a <=( (not A234)  and  a66761a );
 a66765a <=( A298  and  (not A269) );
 a66768a <=( (not A302)  and  (not A301) );
 a66769a <=( a66768a  and  a66765a );
 a66770a <=( a66769a  and  a66762a );
 a66774a <=( A167  and  (not A168) );
 a66775a <=( (not A170)  and  a66774a );
 a66778a <=( (not A199)  and  (not A166) );
 a66781a <=( A232  and  A200 );
 a66782a <=( a66781a  and  a66778a );
 a66783a <=( a66782a  and  a66775a );
 a66787a <=( A235  and  A234 );
 a66788a <=( (not A233)  and  a66787a );
 a66791a <=( (not A299)  and  A298 );
 a66794a <=( A301  and  A300 );
 a66795a <=( a66794a  and  a66791a );
 a66796a <=( a66795a  and  a66788a );
 a66800a <=( A167  and  (not A168) );
 a66801a <=( (not A170)  and  a66800a );
 a66804a <=( (not A199)  and  (not A166) );
 a66807a <=( A232  and  A200 );
 a66808a <=( a66807a  and  a66804a );
 a66809a <=( a66808a  and  a66801a );
 a66813a <=( A235  and  A234 );
 a66814a <=( (not A233)  and  a66813a );
 a66817a <=( (not A299)  and  A298 );
 a66820a <=( A302  and  A300 );
 a66821a <=( a66820a  and  a66817a );
 a66822a <=( a66821a  and  a66814a );
 a66826a <=( A167  and  (not A168) );
 a66827a <=( (not A170)  and  a66826a );
 a66830a <=( (not A199)  and  (not A166) );
 a66833a <=( A232  and  A200 );
 a66834a <=( a66833a  and  a66830a );
 a66835a <=( a66834a  and  a66827a );
 a66839a <=( A235  and  A234 );
 a66840a <=( (not A233)  and  a66839a );
 a66843a <=( (not A266)  and  A265 );
 a66846a <=( A268  and  A267 );
 a66847a <=( a66846a  and  a66843a );
 a66848a <=( a66847a  and  a66840a );
 a66852a <=( A167  and  (not A168) );
 a66853a <=( (not A170)  and  a66852a );
 a66856a <=( (not A199)  and  (not A166) );
 a66859a <=( A232  and  A200 );
 a66860a <=( a66859a  and  a66856a );
 a66861a <=( a66860a  and  a66853a );
 a66865a <=( A235  and  A234 );
 a66866a <=( (not A233)  and  a66865a );
 a66869a <=( (not A266)  and  A265 );
 a66872a <=( A269  and  A267 );
 a66873a <=( a66872a  and  a66869a );
 a66874a <=( a66873a  and  a66866a );
 a66878a <=( A167  and  (not A168) );
 a66879a <=( (not A170)  and  a66878a );
 a66882a <=( (not A199)  and  (not A166) );
 a66885a <=( A232  and  A200 );
 a66886a <=( a66885a  and  a66882a );
 a66887a <=( a66886a  and  a66879a );
 a66891a <=( A236  and  A234 );
 a66892a <=( (not A233)  and  a66891a );
 a66895a <=( (not A299)  and  A298 );
 a66898a <=( A301  and  A300 );
 a66899a <=( a66898a  and  a66895a );
 a66900a <=( a66899a  and  a66892a );
 a66904a <=( A167  and  (not A168) );
 a66905a <=( (not A170)  and  a66904a );
 a66908a <=( (not A199)  and  (not A166) );
 a66911a <=( A232  and  A200 );
 a66912a <=( a66911a  and  a66908a );
 a66913a <=( a66912a  and  a66905a );
 a66917a <=( A236  and  A234 );
 a66918a <=( (not A233)  and  a66917a );
 a66921a <=( (not A299)  and  A298 );
 a66924a <=( A302  and  A300 );
 a66925a <=( a66924a  and  a66921a );
 a66926a <=( a66925a  and  a66918a );
 a66930a <=( A167  and  (not A168) );
 a66931a <=( (not A170)  and  a66930a );
 a66934a <=( (not A199)  and  (not A166) );
 a66937a <=( A232  and  A200 );
 a66938a <=( a66937a  and  a66934a );
 a66939a <=( a66938a  and  a66931a );
 a66943a <=( A236  and  A234 );
 a66944a <=( (not A233)  and  a66943a );
 a66947a <=( (not A266)  and  A265 );
 a66950a <=( A268  and  A267 );
 a66951a <=( a66950a  and  a66947a );
 a66952a <=( a66951a  and  a66944a );
 a66956a <=( A167  and  (not A168) );
 a66957a <=( (not A170)  and  a66956a );
 a66960a <=( (not A199)  and  (not A166) );
 a66963a <=( A232  and  A200 );
 a66964a <=( a66963a  and  a66960a );
 a66965a <=( a66964a  and  a66957a );
 a66969a <=( A236  and  A234 );
 a66970a <=( (not A233)  and  a66969a );
 a66973a <=( (not A266)  and  A265 );
 a66976a <=( A269  and  A267 );
 a66977a <=( a66976a  and  a66973a );
 a66978a <=( a66977a  and  a66970a );
 a66982a <=( A167  and  (not A168) );
 a66983a <=( (not A170)  and  a66982a );
 a66986a <=( (not A199)  and  (not A166) );
 a66989a <=( (not A232)  and  A200 );
 a66990a <=( a66989a  and  a66986a );
 a66991a <=( a66990a  and  a66983a );
 a66995a <=( (not A268)  and  (not A266) );
 a66996a <=( (not A233)  and  a66995a );
 a66999a <=( A298  and  (not A269) );
 a67002a <=( (not A302)  and  (not A301) );
 a67003a <=( a67002a  and  a66999a );
 a67004a <=( a67003a  and  a66996a );
 a67008a <=( (not A167)  and  (not A168) );
 a67009a <=( (not A170)  and  a67008a );
 a67012a <=( (not A199)  and  A166 );
 a67015a <=( A232  and  A200 );
 a67016a <=( a67015a  and  a67012a );
 a67017a <=( a67016a  and  a67009a );
 a67021a <=( (not A268)  and  A265 );
 a67022a <=( A233  and  a67021a );
 a67025a <=( (not A299)  and  (not A269) );
 a67028a <=( (not A302)  and  (not A301) );
 a67029a <=( a67028a  and  a67025a );
 a67030a <=( a67029a  and  a67022a );
 a67034a <=( (not A167)  and  (not A168) );
 a67035a <=( (not A170)  and  a67034a );
 a67038a <=( (not A199)  and  A166 );
 a67041a <=( (not A233)  and  A200 );
 a67042a <=( a67041a  and  a67038a );
 a67043a <=( a67042a  and  a67035a );
 a67047a <=( A265  and  (not A236) );
 a67048a <=( (not A235)  and  a67047a );
 a67051a <=( A298  and  A266 );
 a67054a <=( (not A302)  and  (not A301) );
 a67055a <=( a67054a  and  a67051a );
 a67056a <=( a67055a  and  a67048a );
 a67060a <=( (not A167)  and  (not A168) );
 a67061a <=( (not A170)  and  a67060a );
 a67064a <=( (not A199)  and  A166 );
 a67067a <=( (not A233)  and  A200 );
 a67068a <=( a67067a  and  a67064a );
 a67069a <=( a67068a  and  a67061a );
 a67073a <=( (not A266)  and  (not A236) );
 a67074a <=( (not A235)  and  a67073a );
 a67077a <=( (not A269)  and  (not A268) );
 a67080a <=( (not A300)  and  A298 );
 a67081a <=( a67080a  and  a67077a );
 a67082a <=( a67081a  and  a67074a );
 a67086a <=( (not A167)  and  (not A168) );
 a67087a <=( (not A170)  and  a67086a );
 a67090a <=( (not A199)  and  A166 );
 a67093a <=( (not A233)  and  A200 );
 a67094a <=( a67093a  and  a67090a );
 a67095a <=( a67094a  and  a67087a );
 a67099a <=( (not A266)  and  (not A236) );
 a67100a <=( (not A235)  and  a67099a );
 a67103a <=( (not A269)  and  (not A268) );
 a67106a <=( A299  and  A298 );
 a67107a <=( a67106a  and  a67103a );
 a67108a <=( a67107a  and  a67100a );
 a67112a <=( (not A167)  and  (not A168) );
 a67113a <=( (not A170)  and  a67112a );
 a67116a <=( (not A199)  and  A166 );
 a67119a <=( (not A233)  and  A200 );
 a67120a <=( a67119a  and  a67116a );
 a67121a <=( a67120a  and  a67113a );
 a67125a <=( (not A266)  and  (not A236) );
 a67126a <=( (not A235)  and  a67125a );
 a67129a <=( (not A269)  and  (not A268) );
 a67132a <=( (not A299)  and  (not A298) );
 a67133a <=( a67132a  and  a67129a );
 a67134a <=( a67133a  and  a67126a );
 a67138a <=( (not A167)  and  (not A168) );
 a67139a <=( (not A170)  and  a67138a );
 a67142a <=( (not A199)  and  A166 );
 a67145a <=( (not A233)  and  A200 );
 a67146a <=( a67145a  and  a67142a );
 a67147a <=( a67146a  and  a67139a );
 a67151a <=( (not A266)  and  (not A236) );
 a67152a <=( (not A235)  and  a67151a );
 a67155a <=( A298  and  (not A267) );
 a67158a <=( (not A302)  and  (not A301) );
 a67159a <=( a67158a  and  a67155a );
 a67160a <=( a67159a  and  a67152a );
 a67164a <=( (not A167)  and  (not A168) );
 a67165a <=( (not A170)  and  a67164a );
 a67168a <=( (not A199)  and  A166 );
 a67171a <=( (not A233)  and  A200 );
 a67172a <=( a67171a  and  a67168a );
 a67173a <=( a67172a  and  a67165a );
 a67177a <=( (not A265)  and  (not A236) );
 a67178a <=( (not A235)  and  a67177a );
 a67181a <=( A298  and  (not A266) );
 a67184a <=( (not A302)  and  (not A301) );
 a67185a <=( a67184a  and  a67181a );
 a67186a <=( a67185a  and  a67178a );
 a67190a <=( (not A167)  and  (not A168) );
 a67191a <=( (not A170)  and  a67190a );
 a67194a <=( (not A199)  and  A166 );
 a67197a <=( (not A233)  and  A200 );
 a67198a <=( a67197a  and  a67194a );
 a67199a <=( a67198a  and  a67191a );
 a67203a <=( (not A268)  and  (not A266) );
 a67204a <=( (not A234)  and  a67203a );
 a67207a <=( A298  and  (not A269) );
 a67210a <=( (not A302)  and  (not A301) );
 a67211a <=( a67210a  and  a67207a );
 a67212a <=( a67211a  and  a67204a );
 a67216a <=( (not A167)  and  (not A168) );
 a67217a <=( (not A170)  and  a67216a );
 a67220a <=( (not A199)  and  A166 );
 a67223a <=( A232  and  A200 );
 a67224a <=( a67223a  and  a67220a );
 a67225a <=( a67224a  and  a67217a );
 a67229a <=( A235  and  A234 );
 a67230a <=( (not A233)  and  a67229a );
 a67233a <=( (not A299)  and  A298 );
 a67236a <=( A301  and  A300 );
 a67237a <=( a67236a  and  a67233a );
 a67238a <=( a67237a  and  a67230a );
 a67242a <=( (not A167)  and  (not A168) );
 a67243a <=( (not A170)  and  a67242a );
 a67246a <=( (not A199)  and  A166 );
 a67249a <=( A232  and  A200 );
 a67250a <=( a67249a  and  a67246a );
 a67251a <=( a67250a  and  a67243a );
 a67255a <=( A235  and  A234 );
 a67256a <=( (not A233)  and  a67255a );
 a67259a <=( (not A299)  and  A298 );
 a67262a <=( A302  and  A300 );
 a67263a <=( a67262a  and  a67259a );
 a67264a <=( a67263a  and  a67256a );
 a67268a <=( (not A167)  and  (not A168) );
 a67269a <=( (not A170)  and  a67268a );
 a67272a <=( (not A199)  and  A166 );
 a67275a <=( A232  and  A200 );
 a67276a <=( a67275a  and  a67272a );
 a67277a <=( a67276a  and  a67269a );
 a67281a <=( A235  and  A234 );
 a67282a <=( (not A233)  and  a67281a );
 a67285a <=( (not A266)  and  A265 );
 a67288a <=( A268  and  A267 );
 a67289a <=( a67288a  and  a67285a );
 a67290a <=( a67289a  and  a67282a );
 a67294a <=( (not A167)  and  (not A168) );
 a67295a <=( (not A170)  and  a67294a );
 a67298a <=( (not A199)  and  A166 );
 a67301a <=( A232  and  A200 );
 a67302a <=( a67301a  and  a67298a );
 a67303a <=( a67302a  and  a67295a );
 a67307a <=( A235  and  A234 );
 a67308a <=( (not A233)  and  a67307a );
 a67311a <=( (not A266)  and  A265 );
 a67314a <=( A269  and  A267 );
 a67315a <=( a67314a  and  a67311a );
 a67316a <=( a67315a  and  a67308a );
 a67320a <=( (not A167)  and  (not A168) );
 a67321a <=( (not A170)  and  a67320a );
 a67324a <=( (not A199)  and  A166 );
 a67327a <=( A232  and  A200 );
 a67328a <=( a67327a  and  a67324a );
 a67329a <=( a67328a  and  a67321a );
 a67333a <=( A236  and  A234 );
 a67334a <=( (not A233)  and  a67333a );
 a67337a <=( (not A299)  and  A298 );
 a67340a <=( A301  and  A300 );
 a67341a <=( a67340a  and  a67337a );
 a67342a <=( a67341a  and  a67334a );
 a67346a <=( (not A167)  and  (not A168) );
 a67347a <=( (not A170)  and  a67346a );
 a67350a <=( (not A199)  and  A166 );
 a67353a <=( A232  and  A200 );
 a67354a <=( a67353a  and  a67350a );
 a67355a <=( a67354a  and  a67347a );
 a67359a <=( A236  and  A234 );
 a67360a <=( (not A233)  and  a67359a );
 a67363a <=( (not A299)  and  A298 );
 a67366a <=( A302  and  A300 );
 a67367a <=( a67366a  and  a67363a );
 a67368a <=( a67367a  and  a67360a );
 a67372a <=( (not A167)  and  (not A168) );
 a67373a <=( (not A170)  and  a67372a );
 a67376a <=( (not A199)  and  A166 );
 a67379a <=( A232  and  A200 );
 a67380a <=( a67379a  and  a67376a );
 a67381a <=( a67380a  and  a67373a );
 a67385a <=( A236  and  A234 );
 a67386a <=( (not A233)  and  a67385a );
 a67389a <=( (not A266)  and  A265 );
 a67392a <=( A268  and  A267 );
 a67393a <=( a67392a  and  a67389a );
 a67394a <=( a67393a  and  a67386a );
 a67398a <=( (not A167)  and  (not A168) );
 a67399a <=( (not A170)  and  a67398a );
 a67402a <=( (not A199)  and  A166 );
 a67405a <=( A232  and  A200 );
 a67406a <=( a67405a  and  a67402a );
 a67407a <=( a67406a  and  a67399a );
 a67411a <=( A236  and  A234 );
 a67412a <=( (not A233)  and  a67411a );
 a67415a <=( (not A266)  and  A265 );
 a67418a <=( A269  and  A267 );
 a67419a <=( a67418a  and  a67415a );
 a67420a <=( a67419a  and  a67412a );
 a67424a <=( (not A167)  and  (not A168) );
 a67425a <=( (not A170)  and  a67424a );
 a67428a <=( (not A199)  and  A166 );
 a67431a <=( (not A232)  and  A200 );
 a67432a <=( a67431a  and  a67428a );
 a67433a <=( a67432a  and  a67425a );
 a67437a <=( (not A268)  and  (not A266) );
 a67438a <=( (not A233)  and  a67437a );
 a67441a <=( A298  and  (not A269) );
 a67444a <=( (not A302)  and  (not A301) );
 a67445a <=( a67444a  and  a67441a );
 a67446a <=( a67445a  and  a67438a );
 a67450a <=( A167  and  (not A168) );
 a67451a <=( A169  and  a67450a );
 a67454a <=( (not A199)  and  (not A166) );
 a67457a <=( A232  and  A200 );
 a67458a <=( a67457a  and  a67454a );
 a67459a <=( a67458a  and  a67451a );
 a67463a <=( (not A268)  and  A265 );
 a67464a <=( A233  and  a67463a );
 a67467a <=( (not A299)  and  (not A269) );
 a67470a <=( (not A302)  and  (not A301) );
 a67471a <=( a67470a  and  a67467a );
 a67472a <=( a67471a  and  a67464a );
 a67476a <=( A167  and  (not A168) );
 a67477a <=( A169  and  a67476a );
 a67480a <=( (not A199)  and  (not A166) );
 a67483a <=( (not A233)  and  A200 );
 a67484a <=( a67483a  and  a67480a );
 a67485a <=( a67484a  and  a67477a );
 a67489a <=( A265  and  (not A236) );
 a67490a <=( (not A235)  and  a67489a );
 a67493a <=( A298  and  A266 );
 a67496a <=( (not A302)  and  (not A301) );
 a67497a <=( a67496a  and  a67493a );
 a67498a <=( a67497a  and  a67490a );
 a67502a <=( A167  and  (not A168) );
 a67503a <=( A169  and  a67502a );
 a67506a <=( (not A199)  and  (not A166) );
 a67509a <=( (not A233)  and  A200 );
 a67510a <=( a67509a  and  a67506a );
 a67511a <=( a67510a  and  a67503a );
 a67515a <=( (not A266)  and  (not A236) );
 a67516a <=( (not A235)  and  a67515a );
 a67519a <=( (not A269)  and  (not A268) );
 a67522a <=( (not A300)  and  A298 );
 a67523a <=( a67522a  and  a67519a );
 a67524a <=( a67523a  and  a67516a );
 a67528a <=( A167  and  (not A168) );
 a67529a <=( A169  and  a67528a );
 a67532a <=( (not A199)  and  (not A166) );
 a67535a <=( (not A233)  and  A200 );
 a67536a <=( a67535a  and  a67532a );
 a67537a <=( a67536a  and  a67529a );
 a67541a <=( (not A266)  and  (not A236) );
 a67542a <=( (not A235)  and  a67541a );
 a67545a <=( (not A269)  and  (not A268) );
 a67548a <=( A299  and  A298 );
 a67549a <=( a67548a  and  a67545a );
 a67550a <=( a67549a  and  a67542a );
 a67554a <=( A167  and  (not A168) );
 a67555a <=( A169  and  a67554a );
 a67558a <=( (not A199)  and  (not A166) );
 a67561a <=( (not A233)  and  A200 );
 a67562a <=( a67561a  and  a67558a );
 a67563a <=( a67562a  and  a67555a );
 a67567a <=( (not A266)  and  (not A236) );
 a67568a <=( (not A235)  and  a67567a );
 a67571a <=( (not A269)  and  (not A268) );
 a67574a <=( (not A299)  and  (not A298) );
 a67575a <=( a67574a  and  a67571a );
 a67576a <=( a67575a  and  a67568a );
 a67580a <=( A167  and  (not A168) );
 a67581a <=( A169  and  a67580a );
 a67584a <=( (not A199)  and  (not A166) );
 a67587a <=( (not A233)  and  A200 );
 a67588a <=( a67587a  and  a67584a );
 a67589a <=( a67588a  and  a67581a );
 a67593a <=( (not A266)  and  (not A236) );
 a67594a <=( (not A235)  and  a67593a );
 a67597a <=( A298  and  (not A267) );
 a67600a <=( (not A302)  and  (not A301) );
 a67601a <=( a67600a  and  a67597a );
 a67602a <=( a67601a  and  a67594a );
 a67606a <=( A167  and  (not A168) );
 a67607a <=( A169  and  a67606a );
 a67610a <=( (not A199)  and  (not A166) );
 a67613a <=( (not A233)  and  A200 );
 a67614a <=( a67613a  and  a67610a );
 a67615a <=( a67614a  and  a67607a );
 a67619a <=( (not A265)  and  (not A236) );
 a67620a <=( (not A235)  and  a67619a );
 a67623a <=( A298  and  (not A266) );
 a67626a <=( (not A302)  and  (not A301) );
 a67627a <=( a67626a  and  a67623a );
 a67628a <=( a67627a  and  a67620a );
 a67632a <=( A167  and  (not A168) );
 a67633a <=( A169  and  a67632a );
 a67636a <=( (not A199)  and  (not A166) );
 a67639a <=( (not A233)  and  A200 );
 a67640a <=( a67639a  and  a67636a );
 a67641a <=( a67640a  and  a67633a );
 a67645a <=( (not A268)  and  (not A266) );
 a67646a <=( (not A234)  and  a67645a );
 a67649a <=( A298  and  (not A269) );
 a67652a <=( (not A302)  and  (not A301) );
 a67653a <=( a67652a  and  a67649a );
 a67654a <=( a67653a  and  a67646a );
 a67658a <=( A167  and  (not A168) );
 a67659a <=( A169  and  a67658a );
 a67662a <=( (not A199)  and  (not A166) );
 a67665a <=( A232  and  A200 );
 a67666a <=( a67665a  and  a67662a );
 a67667a <=( a67666a  and  a67659a );
 a67671a <=( A235  and  A234 );
 a67672a <=( (not A233)  and  a67671a );
 a67675a <=( (not A299)  and  A298 );
 a67678a <=( A301  and  A300 );
 a67679a <=( a67678a  and  a67675a );
 a67680a <=( a67679a  and  a67672a );
 a67684a <=( A167  and  (not A168) );
 a67685a <=( A169  and  a67684a );
 a67688a <=( (not A199)  and  (not A166) );
 a67691a <=( A232  and  A200 );
 a67692a <=( a67691a  and  a67688a );
 a67693a <=( a67692a  and  a67685a );
 a67697a <=( A235  and  A234 );
 a67698a <=( (not A233)  and  a67697a );
 a67701a <=( (not A299)  and  A298 );
 a67704a <=( A302  and  A300 );
 a67705a <=( a67704a  and  a67701a );
 a67706a <=( a67705a  and  a67698a );
 a67710a <=( A167  and  (not A168) );
 a67711a <=( A169  and  a67710a );
 a67714a <=( (not A199)  and  (not A166) );
 a67717a <=( A232  and  A200 );
 a67718a <=( a67717a  and  a67714a );
 a67719a <=( a67718a  and  a67711a );
 a67723a <=( A235  and  A234 );
 a67724a <=( (not A233)  and  a67723a );
 a67727a <=( (not A266)  and  A265 );
 a67730a <=( A268  and  A267 );
 a67731a <=( a67730a  and  a67727a );
 a67732a <=( a67731a  and  a67724a );
 a67736a <=( A167  and  (not A168) );
 a67737a <=( A169  and  a67736a );
 a67740a <=( (not A199)  and  (not A166) );
 a67743a <=( A232  and  A200 );
 a67744a <=( a67743a  and  a67740a );
 a67745a <=( a67744a  and  a67737a );
 a67749a <=( A235  and  A234 );
 a67750a <=( (not A233)  and  a67749a );
 a67753a <=( (not A266)  and  A265 );
 a67756a <=( A269  and  A267 );
 a67757a <=( a67756a  and  a67753a );
 a67758a <=( a67757a  and  a67750a );
 a67762a <=( A167  and  (not A168) );
 a67763a <=( A169  and  a67762a );
 a67766a <=( (not A199)  and  (not A166) );
 a67769a <=( A232  and  A200 );
 a67770a <=( a67769a  and  a67766a );
 a67771a <=( a67770a  and  a67763a );
 a67775a <=( A236  and  A234 );
 a67776a <=( (not A233)  and  a67775a );
 a67779a <=( (not A299)  and  A298 );
 a67782a <=( A301  and  A300 );
 a67783a <=( a67782a  and  a67779a );
 a67784a <=( a67783a  and  a67776a );
 a67788a <=( A167  and  (not A168) );
 a67789a <=( A169  and  a67788a );
 a67792a <=( (not A199)  and  (not A166) );
 a67795a <=( A232  and  A200 );
 a67796a <=( a67795a  and  a67792a );
 a67797a <=( a67796a  and  a67789a );
 a67801a <=( A236  and  A234 );
 a67802a <=( (not A233)  and  a67801a );
 a67805a <=( (not A299)  and  A298 );
 a67808a <=( A302  and  A300 );
 a67809a <=( a67808a  and  a67805a );
 a67810a <=( a67809a  and  a67802a );
 a67814a <=( A167  and  (not A168) );
 a67815a <=( A169  and  a67814a );
 a67818a <=( (not A199)  and  (not A166) );
 a67821a <=( A232  and  A200 );
 a67822a <=( a67821a  and  a67818a );
 a67823a <=( a67822a  and  a67815a );
 a67827a <=( A236  and  A234 );
 a67828a <=( (not A233)  and  a67827a );
 a67831a <=( (not A266)  and  A265 );
 a67834a <=( A268  and  A267 );
 a67835a <=( a67834a  and  a67831a );
 a67836a <=( a67835a  and  a67828a );
 a67840a <=( A167  and  (not A168) );
 a67841a <=( A169  and  a67840a );
 a67844a <=( (not A199)  and  (not A166) );
 a67847a <=( A232  and  A200 );
 a67848a <=( a67847a  and  a67844a );
 a67849a <=( a67848a  and  a67841a );
 a67853a <=( A236  and  A234 );
 a67854a <=( (not A233)  and  a67853a );
 a67857a <=( (not A266)  and  A265 );
 a67860a <=( A269  and  A267 );
 a67861a <=( a67860a  and  a67857a );
 a67862a <=( a67861a  and  a67854a );
 a67866a <=( A167  and  (not A168) );
 a67867a <=( A169  and  a67866a );
 a67870a <=( (not A199)  and  (not A166) );
 a67873a <=( (not A232)  and  A200 );
 a67874a <=( a67873a  and  a67870a );
 a67875a <=( a67874a  and  a67867a );
 a67879a <=( (not A268)  and  (not A266) );
 a67880a <=( (not A233)  and  a67879a );
 a67883a <=( A298  and  (not A269) );
 a67886a <=( (not A302)  and  (not A301) );
 a67887a <=( a67886a  and  a67883a );
 a67888a <=( a67887a  and  a67880a );
 a67892a <=( A167  and  (not A168) );
 a67893a <=( A169  and  a67892a );
 a67896a <=( A199  and  (not A166) );
 a67899a <=( A201  and  (not A200) );
 a67900a <=( a67899a  and  a67896a );
 a67901a <=( a67900a  and  a67893a );
 a67905a <=( A233  and  A232 );
 a67906a <=( A202  and  a67905a );
 a67909a <=( (not A267)  and  A265 );
 a67912a <=( (not A300)  and  (not A299) );
 a67913a <=( a67912a  and  a67909a );
 a67914a <=( a67913a  and  a67906a );
 a67918a <=( A167  and  (not A168) );
 a67919a <=( A169  and  a67918a );
 a67922a <=( A199  and  (not A166) );
 a67925a <=( A201  and  (not A200) );
 a67926a <=( a67925a  and  a67922a );
 a67927a <=( a67926a  and  a67919a );
 a67931a <=( A233  and  A232 );
 a67932a <=( A202  and  a67931a );
 a67935a <=( (not A267)  and  A265 );
 a67938a <=( A299  and  A298 );
 a67939a <=( a67938a  and  a67935a );
 a67940a <=( a67939a  and  a67932a );
 a67944a <=( A167  and  (not A168) );
 a67945a <=( A169  and  a67944a );
 a67948a <=( A199  and  (not A166) );
 a67951a <=( A201  and  (not A200) );
 a67952a <=( a67951a  and  a67948a );
 a67953a <=( a67952a  and  a67945a );
 a67957a <=( A233  and  A232 );
 a67958a <=( A202  and  a67957a );
 a67961a <=( (not A267)  and  A265 );
 a67964a <=( (not A299)  and  (not A298) );
 a67965a <=( a67964a  and  a67961a );
 a67966a <=( a67965a  and  a67958a );
 a67970a <=( A167  and  (not A168) );
 a67971a <=( A169  and  a67970a );
 a67974a <=( A199  and  (not A166) );
 a67977a <=( A201  and  (not A200) );
 a67978a <=( a67977a  and  a67974a );
 a67979a <=( a67978a  and  a67971a );
 a67983a <=( A233  and  A232 );
 a67984a <=( A202  and  a67983a );
 a67987a <=( A266  and  A265 );
 a67990a <=( (not A300)  and  (not A299) );
 a67991a <=( a67990a  and  a67987a );
 a67992a <=( a67991a  and  a67984a );
 a67996a <=( A167  and  (not A168) );
 a67997a <=( A169  and  a67996a );
 a68000a <=( A199  and  (not A166) );
 a68003a <=( A201  and  (not A200) );
 a68004a <=( a68003a  and  a68000a );
 a68005a <=( a68004a  and  a67997a );
 a68009a <=( A233  and  A232 );
 a68010a <=( A202  and  a68009a );
 a68013a <=( A266  and  A265 );
 a68016a <=( A299  and  A298 );
 a68017a <=( a68016a  and  a68013a );
 a68018a <=( a68017a  and  a68010a );
 a68022a <=( A167  and  (not A168) );
 a68023a <=( A169  and  a68022a );
 a68026a <=( A199  and  (not A166) );
 a68029a <=( A201  and  (not A200) );
 a68030a <=( a68029a  and  a68026a );
 a68031a <=( a68030a  and  a68023a );
 a68035a <=( A233  and  A232 );
 a68036a <=( A202  and  a68035a );
 a68039a <=( A266  and  A265 );
 a68042a <=( (not A299)  and  (not A298) );
 a68043a <=( a68042a  and  a68039a );
 a68044a <=( a68043a  and  a68036a );
 a68048a <=( A167  and  (not A168) );
 a68049a <=( A169  and  a68048a );
 a68052a <=( A199  and  (not A166) );
 a68055a <=( A201  and  (not A200) );
 a68056a <=( a68055a  and  a68052a );
 a68057a <=( a68056a  and  a68049a );
 a68061a <=( A233  and  A232 );
 a68062a <=( A202  and  a68061a );
 a68065a <=( (not A266)  and  (not A265) );
 a68068a <=( (not A300)  and  (not A299) );
 a68069a <=( a68068a  and  a68065a );
 a68070a <=( a68069a  and  a68062a );
 a68074a <=( A167  and  (not A168) );
 a68075a <=( A169  and  a68074a );
 a68078a <=( A199  and  (not A166) );
 a68081a <=( A201  and  (not A200) );
 a68082a <=( a68081a  and  a68078a );
 a68083a <=( a68082a  and  a68075a );
 a68087a <=( A233  and  A232 );
 a68088a <=( A202  and  a68087a );
 a68091a <=( (not A266)  and  (not A265) );
 a68094a <=( A299  and  A298 );
 a68095a <=( a68094a  and  a68091a );
 a68096a <=( a68095a  and  a68088a );
 a68100a <=( A167  and  (not A168) );
 a68101a <=( A169  and  a68100a );
 a68104a <=( A199  and  (not A166) );
 a68107a <=( A201  and  (not A200) );
 a68108a <=( a68107a  and  a68104a );
 a68109a <=( a68108a  and  a68101a );
 a68113a <=( A233  and  A232 );
 a68114a <=( A202  and  a68113a );
 a68117a <=( (not A266)  and  (not A265) );
 a68120a <=( (not A299)  and  (not A298) );
 a68121a <=( a68120a  and  a68117a );
 a68122a <=( a68121a  and  a68114a );
 a68126a <=( A167  and  (not A168) );
 a68127a <=( A169  and  a68126a );
 a68130a <=( A199  and  (not A166) );
 a68133a <=( A201  and  (not A200) );
 a68134a <=( a68133a  and  a68130a );
 a68135a <=( a68134a  and  a68127a );
 a68139a <=( A233  and  (not A232) );
 a68140a <=( A202  and  a68139a );
 a68143a <=( (not A299)  and  A298 );
 a68146a <=( A301  and  A300 );
 a68147a <=( a68146a  and  a68143a );
 a68148a <=( a68147a  and  a68140a );
 a68152a <=( A167  and  (not A168) );
 a68153a <=( A169  and  a68152a );
 a68156a <=( A199  and  (not A166) );
 a68159a <=( A201  and  (not A200) );
 a68160a <=( a68159a  and  a68156a );
 a68161a <=( a68160a  and  a68153a );
 a68165a <=( A233  and  (not A232) );
 a68166a <=( A202  and  a68165a );
 a68169a <=( (not A299)  and  A298 );
 a68172a <=( A302  and  A300 );
 a68173a <=( a68172a  and  a68169a );
 a68174a <=( a68173a  and  a68166a );
 a68178a <=( A167  and  (not A168) );
 a68179a <=( A169  and  a68178a );
 a68182a <=( A199  and  (not A166) );
 a68185a <=( A201  and  (not A200) );
 a68186a <=( a68185a  and  a68182a );
 a68187a <=( a68186a  and  a68179a );
 a68191a <=( A233  and  (not A232) );
 a68192a <=( A202  and  a68191a );
 a68195a <=( (not A266)  and  A265 );
 a68198a <=( A268  and  A267 );
 a68199a <=( a68198a  and  a68195a );
 a68200a <=( a68199a  and  a68192a );
 a68204a <=( A167  and  (not A168) );
 a68205a <=( A169  and  a68204a );
 a68208a <=( A199  and  (not A166) );
 a68211a <=( A201  and  (not A200) );
 a68212a <=( a68211a  and  a68208a );
 a68213a <=( a68212a  and  a68205a );
 a68217a <=( A233  and  (not A232) );
 a68218a <=( A202  and  a68217a );
 a68221a <=( (not A266)  and  A265 );
 a68224a <=( A269  and  A267 );
 a68225a <=( a68224a  and  a68221a );
 a68226a <=( a68225a  and  a68218a );
 a68230a <=( A167  and  (not A168) );
 a68231a <=( A169  and  a68230a );
 a68234a <=( A199  and  (not A166) );
 a68237a <=( A201  and  (not A200) );
 a68238a <=( a68237a  and  a68234a );
 a68239a <=( a68238a  and  a68231a );
 a68243a <=( (not A234)  and  (not A233) );
 a68244a <=( A202  and  a68243a );
 a68247a <=( A266  and  A265 );
 a68250a <=( (not A300)  and  A298 );
 a68251a <=( a68250a  and  a68247a );
 a68252a <=( a68251a  and  a68244a );
 a68256a <=( A167  and  (not A168) );
 a68257a <=( A169  and  a68256a );
 a68260a <=( A199  and  (not A166) );
 a68263a <=( A201  and  (not A200) );
 a68264a <=( a68263a  and  a68260a );
 a68265a <=( a68264a  and  a68257a );
 a68269a <=( (not A234)  and  (not A233) );
 a68270a <=( A202  and  a68269a );
 a68273a <=( A266  and  A265 );
 a68276a <=( A299  and  A298 );
 a68277a <=( a68276a  and  a68273a );
 a68278a <=( a68277a  and  a68270a );
 a68282a <=( A167  and  (not A168) );
 a68283a <=( A169  and  a68282a );
 a68286a <=( A199  and  (not A166) );
 a68289a <=( A201  and  (not A200) );
 a68290a <=( a68289a  and  a68286a );
 a68291a <=( a68290a  and  a68283a );
 a68295a <=( (not A234)  and  (not A233) );
 a68296a <=( A202  and  a68295a );
 a68299a <=( A266  and  A265 );
 a68302a <=( (not A299)  and  (not A298) );
 a68303a <=( a68302a  and  a68299a );
 a68304a <=( a68303a  and  a68296a );
 a68308a <=( A167  and  (not A168) );
 a68309a <=( A169  and  a68308a );
 a68312a <=( A199  and  (not A166) );
 a68315a <=( A201  and  (not A200) );
 a68316a <=( a68315a  and  a68312a );
 a68317a <=( a68316a  and  a68309a );
 a68321a <=( (not A234)  and  (not A233) );
 a68322a <=( A202  and  a68321a );
 a68325a <=( (not A267)  and  (not A266) );
 a68328a <=( (not A300)  and  A298 );
 a68329a <=( a68328a  and  a68325a );
 a68330a <=( a68329a  and  a68322a );
 a68334a <=( A167  and  (not A168) );
 a68335a <=( A169  and  a68334a );
 a68338a <=( A199  and  (not A166) );
 a68341a <=( A201  and  (not A200) );
 a68342a <=( a68341a  and  a68338a );
 a68343a <=( a68342a  and  a68335a );
 a68347a <=( (not A234)  and  (not A233) );
 a68348a <=( A202  and  a68347a );
 a68351a <=( (not A267)  and  (not A266) );
 a68354a <=( A299  and  A298 );
 a68355a <=( a68354a  and  a68351a );
 a68356a <=( a68355a  and  a68348a );
 a68360a <=( A167  and  (not A168) );
 a68361a <=( A169  and  a68360a );
 a68364a <=( A199  and  (not A166) );
 a68367a <=( A201  and  (not A200) );
 a68368a <=( a68367a  and  a68364a );
 a68369a <=( a68368a  and  a68361a );
 a68373a <=( (not A234)  and  (not A233) );
 a68374a <=( A202  and  a68373a );
 a68377a <=( (not A267)  and  (not A266) );
 a68380a <=( (not A299)  and  (not A298) );
 a68381a <=( a68380a  and  a68377a );
 a68382a <=( a68381a  and  a68374a );
 a68386a <=( A167  and  (not A168) );
 a68387a <=( A169  and  a68386a );
 a68390a <=( A199  and  (not A166) );
 a68393a <=( A201  and  (not A200) );
 a68394a <=( a68393a  and  a68390a );
 a68395a <=( a68394a  and  a68387a );
 a68399a <=( (not A234)  and  (not A233) );
 a68400a <=( A202  and  a68399a );
 a68403a <=( (not A266)  and  (not A265) );
 a68406a <=( (not A300)  and  A298 );
 a68407a <=( a68406a  and  a68403a );
 a68408a <=( a68407a  and  a68400a );
 a68412a <=( A167  and  (not A168) );
 a68413a <=( A169  and  a68412a );
 a68416a <=( A199  and  (not A166) );
 a68419a <=( A201  and  (not A200) );
 a68420a <=( a68419a  and  a68416a );
 a68421a <=( a68420a  and  a68413a );
 a68425a <=( (not A234)  and  (not A233) );
 a68426a <=( A202  and  a68425a );
 a68429a <=( (not A266)  and  (not A265) );
 a68432a <=( A299  and  A298 );
 a68433a <=( a68432a  and  a68429a );
 a68434a <=( a68433a  and  a68426a );
 a68438a <=( A167  and  (not A168) );
 a68439a <=( A169  and  a68438a );
 a68442a <=( A199  and  (not A166) );
 a68445a <=( A201  and  (not A200) );
 a68446a <=( a68445a  and  a68442a );
 a68447a <=( a68446a  and  a68439a );
 a68451a <=( (not A234)  and  (not A233) );
 a68452a <=( A202  and  a68451a );
 a68455a <=( (not A266)  and  (not A265) );
 a68458a <=( (not A299)  and  (not A298) );
 a68459a <=( a68458a  and  a68455a );
 a68460a <=( a68459a  and  a68452a );
 a68464a <=( A167  and  (not A168) );
 a68465a <=( A169  and  a68464a );
 a68468a <=( A199  and  (not A166) );
 a68471a <=( A201  and  (not A200) );
 a68472a <=( a68471a  and  a68468a );
 a68473a <=( a68472a  and  a68465a );
 a68477a <=( (not A233)  and  A232 );
 a68478a <=( A202  and  a68477a );
 a68481a <=( A235  and  A234 );
 a68484a <=( A299  and  (not A298) );
 a68485a <=( a68484a  and  a68481a );
 a68486a <=( a68485a  and  a68478a );
 a68490a <=( A167  and  (not A168) );
 a68491a <=( A169  and  a68490a );
 a68494a <=( A199  and  (not A166) );
 a68497a <=( A201  and  (not A200) );
 a68498a <=( a68497a  and  a68494a );
 a68499a <=( a68498a  and  a68491a );
 a68503a <=( (not A233)  and  A232 );
 a68504a <=( A202  and  a68503a );
 a68507a <=( A235  and  A234 );
 a68510a <=( A266  and  (not A265) );
 a68511a <=( a68510a  and  a68507a );
 a68512a <=( a68511a  and  a68504a );
 a68516a <=( A167  and  (not A168) );
 a68517a <=( A169  and  a68516a );
 a68520a <=( A199  and  (not A166) );
 a68523a <=( A201  and  (not A200) );
 a68524a <=( a68523a  and  a68520a );
 a68525a <=( a68524a  and  a68517a );
 a68529a <=( (not A233)  and  A232 );
 a68530a <=( A202  and  a68529a );
 a68533a <=( A236  and  A234 );
 a68536a <=( A299  and  (not A298) );
 a68537a <=( a68536a  and  a68533a );
 a68538a <=( a68537a  and  a68530a );
 a68542a <=( A167  and  (not A168) );
 a68543a <=( A169  and  a68542a );
 a68546a <=( A199  and  (not A166) );
 a68549a <=( A201  and  (not A200) );
 a68550a <=( a68549a  and  a68546a );
 a68551a <=( a68550a  and  a68543a );
 a68555a <=( (not A233)  and  A232 );
 a68556a <=( A202  and  a68555a );
 a68559a <=( A236  and  A234 );
 a68562a <=( A266  and  (not A265) );
 a68563a <=( a68562a  and  a68559a );
 a68564a <=( a68563a  and  a68556a );
 a68568a <=( A167  and  (not A168) );
 a68569a <=( A169  and  a68568a );
 a68572a <=( A199  and  (not A166) );
 a68575a <=( A201  and  (not A200) );
 a68576a <=( a68575a  and  a68572a );
 a68577a <=( a68576a  and  a68569a );
 a68581a <=( (not A233)  and  (not A232) );
 a68582a <=( A202  and  a68581a );
 a68585a <=( A266  and  A265 );
 a68588a <=( (not A300)  and  A298 );
 a68589a <=( a68588a  and  a68585a );
 a68590a <=( a68589a  and  a68582a );
 a68594a <=( A167  and  (not A168) );
 a68595a <=( A169  and  a68594a );
 a68598a <=( A199  and  (not A166) );
 a68601a <=( A201  and  (not A200) );
 a68602a <=( a68601a  and  a68598a );
 a68603a <=( a68602a  and  a68595a );
 a68607a <=( (not A233)  and  (not A232) );
 a68608a <=( A202  and  a68607a );
 a68611a <=( A266  and  A265 );
 a68614a <=( A299  and  A298 );
 a68615a <=( a68614a  and  a68611a );
 a68616a <=( a68615a  and  a68608a );
 a68620a <=( A167  and  (not A168) );
 a68621a <=( A169  and  a68620a );
 a68624a <=( A199  and  (not A166) );
 a68627a <=( A201  and  (not A200) );
 a68628a <=( a68627a  and  a68624a );
 a68629a <=( a68628a  and  a68621a );
 a68633a <=( (not A233)  and  (not A232) );
 a68634a <=( A202  and  a68633a );
 a68637a <=( A266  and  A265 );
 a68640a <=( (not A299)  and  (not A298) );
 a68641a <=( a68640a  and  a68637a );
 a68642a <=( a68641a  and  a68634a );
 a68646a <=( A167  and  (not A168) );
 a68647a <=( A169  and  a68646a );
 a68650a <=( A199  and  (not A166) );
 a68653a <=( A201  and  (not A200) );
 a68654a <=( a68653a  and  a68650a );
 a68655a <=( a68654a  and  a68647a );
 a68659a <=( (not A233)  and  (not A232) );
 a68660a <=( A202  and  a68659a );
 a68663a <=( (not A267)  and  (not A266) );
 a68666a <=( (not A300)  and  A298 );
 a68667a <=( a68666a  and  a68663a );
 a68668a <=( a68667a  and  a68660a );
 a68672a <=( A167  and  (not A168) );
 a68673a <=( A169  and  a68672a );
 a68676a <=( A199  and  (not A166) );
 a68679a <=( A201  and  (not A200) );
 a68680a <=( a68679a  and  a68676a );
 a68681a <=( a68680a  and  a68673a );
 a68685a <=( (not A233)  and  (not A232) );
 a68686a <=( A202  and  a68685a );
 a68689a <=( (not A267)  and  (not A266) );
 a68692a <=( A299  and  A298 );
 a68693a <=( a68692a  and  a68689a );
 a68694a <=( a68693a  and  a68686a );
 a68698a <=( A167  and  (not A168) );
 a68699a <=( A169  and  a68698a );
 a68702a <=( A199  and  (not A166) );
 a68705a <=( A201  and  (not A200) );
 a68706a <=( a68705a  and  a68702a );
 a68707a <=( a68706a  and  a68699a );
 a68711a <=( (not A233)  and  (not A232) );
 a68712a <=( A202  and  a68711a );
 a68715a <=( (not A267)  and  (not A266) );
 a68718a <=( (not A299)  and  (not A298) );
 a68719a <=( a68718a  and  a68715a );
 a68720a <=( a68719a  and  a68712a );
 a68724a <=( A167  and  (not A168) );
 a68725a <=( A169  and  a68724a );
 a68728a <=( A199  and  (not A166) );
 a68731a <=( A201  and  (not A200) );
 a68732a <=( a68731a  and  a68728a );
 a68733a <=( a68732a  and  a68725a );
 a68737a <=( (not A233)  and  (not A232) );
 a68738a <=( A202  and  a68737a );
 a68741a <=( (not A266)  and  (not A265) );
 a68744a <=( (not A300)  and  A298 );
 a68745a <=( a68744a  and  a68741a );
 a68746a <=( a68745a  and  a68738a );
 a68750a <=( A167  and  (not A168) );
 a68751a <=( A169  and  a68750a );
 a68754a <=( A199  and  (not A166) );
 a68757a <=( A201  and  (not A200) );
 a68758a <=( a68757a  and  a68754a );
 a68759a <=( a68758a  and  a68751a );
 a68763a <=( (not A233)  and  (not A232) );
 a68764a <=( A202  and  a68763a );
 a68767a <=( (not A266)  and  (not A265) );
 a68770a <=( A299  and  A298 );
 a68771a <=( a68770a  and  a68767a );
 a68772a <=( a68771a  and  a68764a );
 a68776a <=( A167  and  (not A168) );
 a68777a <=( A169  and  a68776a );
 a68780a <=( A199  and  (not A166) );
 a68783a <=( A201  and  (not A200) );
 a68784a <=( a68783a  and  a68780a );
 a68785a <=( a68784a  and  a68777a );
 a68789a <=( (not A233)  and  (not A232) );
 a68790a <=( A202  and  a68789a );
 a68793a <=( (not A266)  and  (not A265) );
 a68796a <=( (not A299)  and  (not A298) );
 a68797a <=( a68796a  and  a68793a );
 a68798a <=( a68797a  and  a68790a );
 a68802a <=( A167  and  (not A168) );
 a68803a <=( A169  and  a68802a );
 a68806a <=( A199  and  (not A166) );
 a68809a <=( A201  and  (not A200) );
 a68810a <=( a68809a  and  a68806a );
 a68811a <=( a68810a  and  a68803a );
 a68815a <=( A233  and  A232 );
 a68816a <=( A203  and  a68815a );
 a68819a <=( (not A267)  and  A265 );
 a68822a <=( (not A300)  and  (not A299) );
 a68823a <=( a68822a  and  a68819a );
 a68824a <=( a68823a  and  a68816a );
 a68828a <=( A167  and  (not A168) );
 a68829a <=( A169  and  a68828a );
 a68832a <=( A199  and  (not A166) );
 a68835a <=( A201  and  (not A200) );
 a68836a <=( a68835a  and  a68832a );
 a68837a <=( a68836a  and  a68829a );
 a68841a <=( A233  and  A232 );
 a68842a <=( A203  and  a68841a );
 a68845a <=( (not A267)  and  A265 );
 a68848a <=( A299  and  A298 );
 a68849a <=( a68848a  and  a68845a );
 a68850a <=( a68849a  and  a68842a );
 a68854a <=( A167  and  (not A168) );
 a68855a <=( A169  and  a68854a );
 a68858a <=( A199  and  (not A166) );
 a68861a <=( A201  and  (not A200) );
 a68862a <=( a68861a  and  a68858a );
 a68863a <=( a68862a  and  a68855a );
 a68867a <=( A233  and  A232 );
 a68868a <=( A203  and  a68867a );
 a68871a <=( (not A267)  and  A265 );
 a68874a <=( (not A299)  and  (not A298) );
 a68875a <=( a68874a  and  a68871a );
 a68876a <=( a68875a  and  a68868a );
 a68880a <=( A167  and  (not A168) );
 a68881a <=( A169  and  a68880a );
 a68884a <=( A199  and  (not A166) );
 a68887a <=( A201  and  (not A200) );
 a68888a <=( a68887a  and  a68884a );
 a68889a <=( a68888a  and  a68881a );
 a68893a <=( A233  and  A232 );
 a68894a <=( A203  and  a68893a );
 a68897a <=( A266  and  A265 );
 a68900a <=( (not A300)  and  (not A299) );
 a68901a <=( a68900a  and  a68897a );
 a68902a <=( a68901a  and  a68894a );
 a68906a <=( A167  and  (not A168) );
 a68907a <=( A169  and  a68906a );
 a68910a <=( A199  and  (not A166) );
 a68913a <=( A201  and  (not A200) );
 a68914a <=( a68913a  and  a68910a );
 a68915a <=( a68914a  and  a68907a );
 a68919a <=( A233  and  A232 );
 a68920a <=( A203  and  a68919a );
 a68923a <=( A266  and  A265 );
 a68926a <=( A299  and  A298 );
 a68927a <=( a68926a  and  a68923a );
 a68928a <=( a68927a  and  a68920a );
 a68932a <=( A167  and  (not A168) );
 a68933a <=( A169  and  a68932a );
 a68936a <=( A199  and  (not A166) );
 a68939a <=( A201  and  (not A200) );
 a68940a <=( a68939a  and  a68936a );
 a68941a <=( a68940a  and  a68933a );
 a68945a <=( A233  and  A232 );
 a68946a <=( A203  and  a68945a );
 a68949a <=( A266  and  A265 );
 a68952a <=( (not A299)  and  (not A298) );
 a68953a <=( a68952a  and  a68949a );
 a68954a <=( a68953a  and  a68946a );
 a68958a <=( A167  and  (not A168) );
 a68959a <=( A169  and  a68958a );
 a68962a <=( A199  and  (not A166) );
 a68965a <=( A201  and  (not A200) );
 a68966a <=( a68965a  and  a68962a );
 a68967a <=( a68966a  and  a68959a );
 a68971a <=( A233  and  A232 );
 a68972a <=( A203  and  a68971a );
 a68975a <=( (not A266)  and  (not A265) );
 a68978a <=( (not A300)  and  (not A299) );
 a68979a <=( a68978a  and  a68975a );
 a68980a <=( a68979a  and  a68972a );
 a68984a <=( A167  and  (not A168) );
 a68985a <=( A169  and  a68984a );
 a68988a <=( A199  and  (not A166) );
 a68991a <=( A201  and  (not A200) );
 a68992a <=( a68991a  and  a68988a );
 a68993a <=( a68992a  and  a68985a );
 a68997a <=( A233  and  A232 );
 a68998a <=( A203  and  a68997a );
 a69001a <=( (not A266)  and  (not A265) );
 a69004a <=( A299  and  A298 );
 a69005a <=( a69004a  and  a69001a );
 a69006a <=( a69005a  and  a68998a );
 a69010a <=( A167  and  (not A168) );
 a69011a <=( A169  and  a69010a );
 a69014a <=( A199  and  (not A166) );
 a69017a <=( A201  and  (not A200) );
 a69018a <=( a69017a  and  a69014a );
 a69019a <=( a69018a  and  a69011a );
 a69023a <=( A233  and  A232 );
 a69024a <=( A203  and  a69023a );
 a69027a <=( (not A266)  and  (not A265) );
 a69030a <=( (not A299)  and  (not A298) );
 a69031a <=( a69030a  and  a69027a );
 a69032a <=( a69031a  and  a69024a );
 a69036a <=( A167  and  (not A168) );
 a69037a <=( A169  and  a69036a );
 a69040a <=( A199  and  (not A166) );
 a69043a <=( A201  and  (not A200) );
 a69044a <=( a69043a  and  a69040a );
 a69045a <=( a69044a  and  a69037a );
 a69049a <=( A233  and  (not A232) );
 a69050a <=( A203  and  a69049a );
 a69053a <=( (not A299)  and  A298 );
 a69056a <=( A301  and  A300 );
 a69057a <=( a69056a  and  a69053a );
 a69058a <=( a69057a  and  a69050a );
 a69062a <=( A167  and  (not A168) );
 a69063a <=( A169  and  a69062a );
 a69066a <=( A199  and  (not A166) );
 a69069a <=( A201  and  (not A200) );
 a69070a <=( a69069a  and  a69066a );
 a69071a <=( a69070a  and  a69063a );
 a69075a <=( A233  and  (not A232) );
 a69076a <=( A203  and  a69075a );
 a69079a <=( (not A299)  and  A298 );
 a69082a <=( A302  and  A300 );
 a69083a <=( a69082a  and  a69079a );
 a69084a <=( a69083a  and  a69076a );
 a69088a <=( A167  and  (not A168) );
 a69089a <=( A169  and  a69088a );
 a69092a <=( A199  and  (not A166) );
 a69095a <=( A201  and  (not A200) );
 a69096a <=( a69095a  and  a69092a );
 a69097a <=( a69096a  and  a69089a );
 a69101a <=( A233  and  (not A232) );
 a69102a <=( A203  and  a69101a );
 a69105a <=( (not A266)  and  A265 );
 a69108a <=( A268  and  A267 );
 a69109a <=( a69108a  and  a69105a );
 a69110a <=( a69109a  and  a69102a );
 a69114a <=( A167  and  (not A168) );
 a69115a <=( A169  and  a69114a );
 a69118a <=( A199  and  (not A166) );
 a69121a <=( A201  and  (not A200) );
 a69122a <=( a69121a  and  a69118a );
 a69123a <=( a69122a  and  a69115a );
 a69127a <=( A233  and  (not A232) );
 a69128a <=( A203  and  a69127a );
 a69131a <=( (not A266)  and  A265 );
 a69134a <=( A269  and  A267 );
 a69135a <=( a69134a  and  a69131a );
 a69136a <=( a69135a  and  a69128a );
 a69140a <=( A167  and  (not A168) );
 a69141a <=( A169  and  a69140a );
 a69144a <=( A199  and  (not A166) );
 a69147a <=( A201  and  (not A200) );
 a69148a <=( a69147a  and  a69144a );
 a69149a <=( a69148a  and  a69141a );
 a69153a <=( (not A234)  and  (not A233) );
 a69154a <=( A203  and  a69153a );
 a69157a <=( A266  and  A265 );
 a69160a <=( (not A300)  and  A298 );
 a69161a <=( a69160a  and  a69157a );
 a69162a <=( a69161a  and  a69154a );
 a69166a <=( A167  and  (not A168) );
 a69167a <=( A169  and  a69166a );
 a69170a <=( A199  and  (not A166) );
 a69173a <=( A201  and  (not A200) );
 a69174a <=( a69173a  and  a69170a );
 a69175a <=( a69174a  and  a69167a );
 a69179a <=( (not A234)  and  (not A233) );
 a69180a <=( A203  and  a69179a );
 a69183a <=( A266  and  A265 );
 a69186a <=( A299  and  A298 );
 a69187a <=( a69186a  and  a69183a );
 a69188a <=( a69187a  and  a69180a );
 a69192a <=( A167  and  (not A168) );
 a69193a <=( A169  and  a69192a );
 a69196a <=( A199  and  (not A166) );
 a69199a <=( A201  and  (not A200) );
 a69200a <=( a69199a  and  a69196a );
 a69201a <=( a69200a  and  a69193a );
 a69205a <=( (not A234)  and  (not A233) );
 a69206a <=( A203  and  a69205a );
 a69209a <=( A266  and  A265 );
 a69212a <=( (not A299)  and  (not A298) );
 a69213a <=( a69212a  and  a69209a );
 a69214a <=( a69213a  and  a69206a );
 a69218a <=( A167  and  (not A168) );
 a69219a <=( A169  and  a69218a );
 a69222a <=( A199  and  (not A166) );
 a69225a <=( A201  and  (not A200) );
 a69226a <=( a69225a  and  a69222a );
 a69227a <=( a69226a  and  a69219a );
 a69231a <=( (not A234)  and  (not A233) );
 a69232a <=( A203  and  a69231a );
 a69235a <=( (not A267)  and  (not A266) );
 a69238a <=( (not A300)  and  A298 );
 a69239a <=( a69238a  and  a69235a );
 a69240a <=( a69239a  and  a69232a );
 a69244a <=( A167  and  (not A168) );
 a69245a <=( A169  and  a69244a );
 a69248a <=( A199  and  (not A166) );
 a69251a <=( A201  and  (not A200) );
 a69252a <=( a69251a  and  a69248a );
 a69253a <=( a69252a  and  a69245a );
 a69257a <=( (not A234)  and  (not A233) );
 a69258a <=( A203  and  a69257a );
 a69261a <=( (not A267)  and  (not A266) );
 a69264a <=( A299  and  A298 );
 a69265a <=( a69264a  and  a69261a );
 a69266a <=( a69265a  and  a69258a );
 a69270a <=( A167  and  (not A168) );
 a69271a <=( A169  and  a69270a );
 a69274a <=( A199  and  (not A166) );
 a69277a <=( A201  and  (not A200) );
 a69278a <=( a69277a  and  a69274a );
 a69279a <=( a69278a  and  a69271a );
 a69283a <=( (not A234)  and  (not A233) );
 a69284a <=( A203  and  a69283a );
 a69287a <=( (not A267)  and  (not A266) );
 a69290a <=( (not A299)  and  (not A298) );
 a69291a <=( a69290a  and  a69287a );
 a69292a <=( a69291a  and  a69284a );
 a69296a <=( A167  and  (not A168) );
 a69297a <=( A169  and  a69296a );
 a69300a <=( A199  and  (not A166) );
 a69303a <=( A201  and  (not A200) );
 a69304a <=( a69303a  and  a69300a );
 a69305a <=( a69304a  and  a69297a );
 a69309a <=( (not A234)  and  (not A233) );
 a69310a <=( A203  and  a69309a );
 a69313a <=( (not A266)  and  (not A265) );
 a69316a <=( (not A300)  and  A298 );
 a69317a <=( a69316a  and  a69313a );
 a69318a <=( a69317a  and  a69310a );
 a69322a <=( A167  and  (not A168) );
 a69323a <=( A169  and  a69322a );
 a69326a <=( A199  and  (not A166) );
 a69329a <=( A201  and  (not A200) );
 a69330a <=( a69329a  and  a69326a );
 a69331a <=( a69330a  and  a69323a );
 a69335a <=( (not A234)  and  (not A233) );
 a69336a <=( A203  and  a69335a );
 a69339a <=( (not A266)  and  (not A265) );
 a69342a <=( A299  and  A298 );
 a69343a <=( a69342a  and  a69339a );
 a69344a <=( a69343a  and  a69336a );
 a69348a <=( A167  and  (not A168) );
 a69349a <=( A169  and  a69348a );
 a69352a <=( A199  and  (not A166) );
 a69355a <=( A201  and  (not A200) );
 a69356a <=( a69355a  and  a69352a );
 a69357a <=( a69356a  and  a69349a );
 a69361a <=( (not A234)  and  (not A233) );
 a69362a <=( A203  and  a69361a );
 a69365a <=( (not A266)  and  (not A265) );
 a69368a <=( (not A299)  and  (not A298) );
 a69369a <=( a69368a  and  a69365a );
 a69370a <=( a69369a  and  a69362a );
 a69374a <=( A167  and  (not A168) );
 a69375a <=( A169  and  a69374a );
 a69378a <=( A199  and  (not A166) );
 a69381a <=( A201  and  (not A200) );
 a69382a <=( a69381a  and  a69378a );
 a69383a <=( a69382a  and  a69375a );
 a69387a <=( (not A233)  and  A232 );
 a69388a <=( A203  and  a69387a );
 a69391a <=( A235  and  A234 );
 a69394a <=( A299  and  (not A298) );
 a69395a <=( a69394a  and  a69391a );
 a69396a <=( a69395a  and  a69388a );
 a69400a <=( A167  and  (not A168) );
 a69401a <=( A169  and  a69400a );
 a69404a <=( A199  and  (not A166) );
 a69407a <=( A201  and  (not A200) );
 a69408a <=( a69407a  and  a69404a );
 a69409a <=( a69408a  and  a69401a );
 a69413a <=( (not A233)  and  A232 );
 a69414a <=( A203  and  a69413a );
 a69417a <=( A235  and  A234 );
 a69420a <=( A266  and  (not A265) );
 a69421a <=( a69420a  and  a69417a );
 a69422a <=( a69421a  and  a69414a );
 a69426a <=( A167  and  (not A168) );
 a69427a <=( A169  and  a69426a );
 a69430a <=( A199  and  (not A166) );
 a69433a <=( A201  and  (not A200) );
 a69434a <=( a69433a  and  a69430a );
 a69435a <=( a69434a  and  a69427a );
 a69439a <=( (not A233)  and  A232 );
 a69440a <=( A203  and  a69439a );
 a69443a <=( A236  and  A234 );
 a69446a <=( A299  and  (not A298) );
 a69447a <=( a69446a  and  a69443a );
 a69448a <=( a69447a  and  a69440a );
 a69452a <=( A167  and  (not A168) );
 a69453a <=( A169  and  a69452a );
 a69456a <=( A199  and  (not A166) );
 a69459a <=( A201  and  (not A200) );
 a69460a <=( a69459a  and  a69456a );
 a69461a <=( a69460a  and  a69453a );
 a69465a <=( (not A233)  and  A232 );
 a69466a <=( A203  and  a69465a );
 a69469a <=( A236  and  A234 );
 a69472a <=( A266  and  (not A265) );
 a69473a <=( a69472a  and  a69469a );
 a69474a <=( a69473a  and  a69466a );
 a69478a <=( A167  and  (not A168) );
 a69479a <=( A169  and  a69478a );
 a69482a <=( A199  and  (not A166) );
 a69485a <=( A201  and  (not A200) );
 a69486a <=( a69485a  and  a69482a );
 a69487a <=( a69486a  and  a69479a );
 a69491a <=( (not A233)  and  (not A232) );
 a69492a <=( A203  and  a69491a );
 a69495a <=( A266  and  A265 );
 a69498a <=( (not A300)  and  A298 );
 a69499a <=( a69498a  and  a69495a );
 a69500a <=( a69499a  and  a69492a );
 a69504a <=( A167  and  (not A168) );
 a69505a <=( A169  and  a69504a );
 a69508a <=( A199  and  (not A166) );
 a69511a <=( A201  and  (not A200) );
 a69512a <=( a69511a  and  a69508a );
 a69513a <=( a69512a  and  a69505a );
 a69517a <=( (not A233)  and  (not A232) );
 a69518a <=( A203  and  a69517a );
 a69521a <=( A266  and  A265 );
 a69524a <=( A299  and  A298 );
 a69525a <=( a69524a  and  a69521a );
 a69526a <=( a69525a  and  a69518a );
 a69530a <=( A167  and  (not A168) );
 a69531a <=( A169  and  a69530a );
 a69534a <=( A199  and  (not A166) );
 a69537a <=( A201  and  (not A200) );
 a69538a <=( a69537a  and  a69534a );
 a69539a <=( a69538a  and  a69531a );
 a69543a <=( (not A233)  and  (not A232) );
 a69544a <=( A203  and  a69543a );
 a69547a <=( A266  and  A265 );
 a69550a <=( (not A299)  and  (not A298) );
 a69551a <=( a69550a  and  a69547a );
 a69552a <=( a69551a  and  a69544a );
 a69556a <=( A167  and  (not A168) );
 a69557a <=( A169  and  a69556a );
 a69560a <=( A199  and  (not A166) );
 a69563a <=( A201  and  (not A200) );
 a69564a <=( a69563a  and  a69560a );
 a69565a <=( a69564a  and  a69557a );
 a69569a <=( (not A233)  and  (not A232) );
 a69570a <=( A203  and  a69569a );
 a69573a <=( (not A267)  and  (not A266) );
 a69576a <=( (not A300)  and  A298 );
 a69577a <=( a69576a  and  a69573a );
 a69578a <=( a69577a  and  a69570a );
 a69582a <=( A167  and  (not A168) );
 a69583a <=( A169  and  a69582a );
 a69586a <=( A199  and  (not A166) );
 a69589a <=( A201  and  (not A200) );
 a69590a <=( a69589a  and  a69586a );
 a69591a <=( a69590a  and  a69583a );
 a69595a <=( (not A233)  and  (not A232) );
 a69596a <=( A203  and  a69595a );
 a69599a <=( (not A267)  and  (not A266) );
 a69602a <=( A299  and  A298 );
 a69603a <=( a69602a  and  a69599a );
 a69604a <=( a69603a  and  a69596a );
 a69608a <=( A167  and  (not A168) );
 a69609a <=( A169  and  a69608a );
 a69612a <=( A199  and  (not A166) );
 a69615a <=( A201  and  (not A200) );
 a69616a <=( a69615a  and  a69612a );
 a69617a <=( a69616a  and  a69609a );
 a69621a <=( (not A233)  and  (not A232) );
 a69622a <=( A203  and  a69621a );
 a69625a <=( (not A267)  and  (not A266) );
 a69628a <=( (not A299)  and  (not A298) );
 a69629a <=( a69628a  and  a69625a );
 a69630a <=( a69629a  and  a69622a );
 a69634a <=( A167  and  (not A168) );
 a69635a <=( A169  and  a69634a );
 a69638a <=( A199  and  (not A166) );
 a69641a <=( A201  and  (not A200) );
 a69642a <=( a69641a  and  a69638a );
 a69643a <=( a69642a  and  a69635a );
 a69647a <=( (not A233)  and  (not A232) );
 a69648a <=( A203  and  a69647a );
 a69651a <=( (not A266)  and  (not A265) );
 a69654a <=( (not A300)  and  A298 );
 a69655a <=( a69654a  and  a69651a );
 a69656a <=( a69655a  and  a69648a );
 a69660a <=( A167  and  (not A168) );
 a69661a <=( A169  and  a69660a );
 a69664a <=( A199  and  (not A166) );
 a69667a <=( A201  and  (not A200) );
 a69668a <=( a69667a  and  a69664a );
 a69669a <=( a69668a  and  a69661a );
 a69673a <=( (not A233)  and  (not A232) );
 a69674a <=( A203  and  a69673a );
 a69677a <=( (not A266)  and  (not A265) );
 a69680a <=( A299  and  A298 );
 a69681a <=( a69680a  and  a69677a );
 a69682a <=( a69681a  and  a69674a );
 a69686a <=( A167  and  (not A168) );
 a69687a <=( A169  and  a69686a );
 a69690a <=( A199  and  (not A166) );
 a69693a <=( A201  and  (not A200) );
 a69694a <=( a69693a  and  a69690a );
 a69695a <=( a69694a  and  a69687a );
 a69699a <=( (not A233)  and  (not A232) );
 a69700a <=( A203  and  a69699a );
 a69703a <=( (not A266)  and  (not A265) );
 a69706a <=( (not A299)  and  (not A298) );
 a69707a <=( a69706a  and  a69703a );
 a69708a <=( a69707a  and  a69700a );
 a69712a <=( (not A167)  and  (not A168) );
 a69713a <=( A169  and  a69712a );
 a69716a <=( (not A199)  and  A166 );
 a69719a <=( A232  and  A200 );
 a69720a <=( a69719a  and  a69716a );
 a69721a <=( a69720a  and  a69713a );
 a69725a <=( (not A268)  and  A265 );
 a69726a <=( A233  and  a69725a );
 a69729a <=( (not A299)  and  (not A269) );
 a69732a <=( (not A302)  and  (not A301) );
 a69733a <=( a69732a  and  a69729a );
 a69734a <=( a69733a  and  a69726a );
 a69738a <=( (not A167)  and  (not A168) );
 a69739a <=( A169  and  a69738a );
 a69742a <=( (not A199)  and  A166 );
 a69745a <=( (not A233)  and  A200 );
 a69746a <=( a69745a  and  a69742a );
 a69747a <=( a69746a  and  a69739a );
 a69751a <=( A265  and  (not A236) );
 a69752a <=( (not A235)  and  a69751a );
 a69755a <=( A298  and  A266 );
 a69758a <=( (not A302)  and  (not A301) );
 a69759a <=( a69758a  and  a69755a );
 a69760a <=( a69759a  and  a69752a );
 a69764a <=( (not A167)  and  (not A168) );
 a69765a <=( A169  and  a69764a );
 a69768a <=( (not A199)  and  A166 );
 a69771a <=( (not A233)  and  A200 );
 a69772a <=( a69771a  and  a69768a );
 a69773a <=( a69772a  and  a69765a );
 a69777a <=( (not A266)  and  (not A236) );
 a69778a <=( (not A235)  and  a69777a );
 a69781a <=( (not A269)  and  (not A268) );
 a69784a <=( (not A300)  and  A298 );
 a69785a <=( a69784a  and  a69781a );
 a69786a <=( a69785a  and  a69778a );
 a69790a <=( (not A167)  and  (not A168) );
 a69791a <=( A169  and  a69790a );
 a69794a <=( (not A199)  and  A166 );
 a69797a <=( (not A233)  and  A200 );
 a69798a <=( a69797a  and  a69794a );
 a69799a <=( a69798a  and  a69791a );
 a69803a <=( (not A266)  and  (not A236) );
 a69804a <=( (not A235)  and  a69803a );
 a69807a <=( (not A269)  and  (not A268) );
 a69810a <=( A299  and  A298 );
 a69811a <=( a69810a  and  a69807a );
 a69812a <=( a69811a  and  a69804a );
 a69816a <=( (not A167)  and  (not A168) );
 a69817a <=( A169  and  a69816a );
 a69820a <=( (not A199)  and  A166 );
 a69823a <=( (not A233)  and  A200 );
 a69824a <=( a69823a  and  a69820a );
 a69825a <=( a69824a  and  a69817a );
 a69829a <=( (not A266)  and  (not A236) );
 a69830a <=( (not A235)  and  a69829a );
 a69833a <=( (not A269)  and  (not A268) );
 a69836a <=( (not A299)  and  (not A298) );
 a69837a <=( a69836a  and  a69833a );
 a69838a <=( a69837a  and  a69830a );
 a69842a <=( (not A167)  and  (not A168) );
 a69843a <=( A169  and  a69842a );
 a69846a <=( (not A199)  and  A166 );
 a69849a <=( (not A233)  and  A200 );
 a69850a <=( a69849a  and  a69846a );
 a69851a <=( a69850a  and  a69843a );
 a69855a <=( (not A266)  and  (not A236) );
 a69856a <=( (not A235)  and  a69855a );
 a69859a <=( A298  and  (not A267) );
 a69862a <=( (not A302)  and  (not A301) );
 a69863a <=( a69862a  and  a69859a );
 a69864a <=( a69863a  and  a69856a );
 a69868a <=( (not A167)  and  (not A168) );
 a69869a <=( A169  and  a69868a );
 a69872a <=( (not A199)  and  A166 );
 a69875a <=( (not A233)  and  A200 );
 a69876a <=( a69875a  and  a69872a );
 a69877a <=( a69876a  and  a69869a );
 a69881a <=( (not A265)  and  (not A236) );
 a69882a <=( (not A235)  and  a69881a );
 a69885a <=( A298  and  (not A266) );
 a69888a <=( (not A302)  and  (not A301) );
 a69889a <=( a69888a  and  a69885a );
 a69890a <=( a69889a  and  a69882a );
 a69894a <=( (not A167)  and  (not A168) );
 a69895a <=( A169  and  a69894a );
 a69898a <=( (not A199)  and  A166 );
 a69901a <=( (not A233)  and  A200 );
 a69902a <=( a69901a  and  a69898a );
 a69903a <=( a69902a  and  a69895a );
 a69907a <=( (not A268)  and  (not A266) );
 a69908a <=( (not A234)  and  a69907a );
 a69911a <=( A298  and  (not A269) );
 a69914a <=( (not A302)  and  (not A301) );
 a69915a <=( a69914a  and  a69911a );
 a69916a <=( a69915a  and  a69908a );
 a69920a <=( (not A167)  and  (not A168) );
 a69921a <=( A169  and  a69920a );
 a69924a <=( (not A199)  and  A166 );
 a69927a <=( A232  and  A200 );
 a69928a <=( a69927a  and  a69924a );
 a69929a <=( a69928a  and  a69921a );
 a69933a <=( A235  and  A234 );
 a69934a <=( (not A233)  and  a69933a );
 a69937a <=( (not A299)  and  A298 );
 a69940a <=( A301  and  A300 );
 a69941a <=( a69940a  and  a69937a );
 a69942a <=( a69941a  and  a69934a );
 a69946a <=( (not A167)  and  (not A168) );
 a69947a <=( A169  and  a69946a );
 a69950a <=( (not A199)  and  A166 );
 a69953a <=( A232  and  A200 );
 a69954a <=( a69953a  and  a69950a );
 a69955a <=( a69954a  and  a69947a );
 a69959a <=( A235  and  A234 );
 a69960a <=( (not A233)  and  a69959a );
 a69963a <=( (not A299)  and  A298 );
 a69966a <=( A302  and  A300 );
 a69967a <=( a69966a  and  a69963a );
 a69968a <=( a69967a  and  a69960a );
 a69972a <=( (not A167)  and  (not A168) );
 a69973a <=( A169  and  a69972a );
 a69976a <=( (not A199)  and  A166 );
 a69979a <=( A232  and  A200 );
 a69980a <=( a69979a  and  a69976a );
 a69981a <=( a69980a  and  a69973a );
 a69985a <=( A235  and  A234 );
 a69986a <=( (not A233)  and  a69985a );
 a69989a <=( (not A266)  and  A265 );
 a69992a <=( A268  and  A267 );
 a69993a <=( a69992a  and  a69989a );
 a69994a <=( a69993a  and  a69986a );
 a69998a <=( (not A167)  and  (not A168) );
 a69999a <=( A169  and  a69998a );
 a70002a <=( (not A199)  and  A166 );
 a70005a <=( A232  and  A200 );
 a70006a <=( a70005a  and  a70002a );
 a70007a <=( a70006a  and  a69999a );
 a70011a <=( A235  and  A234 );
 a70012a <=( (not A233)  and  a70011a );
 a70015a <=( (not A266)  and  A265 );
 a70018a <=( A269  and  A267 );
 a70019a <=( a70018a  and  a70015a );
 a70020a <=( a70019a  and  a70012a );
 a70024a <=( (not A167)  and  (not A168) );
 a70025a <=( A169  and  a70024a );
 a70028a <=( (not A199)  and  A166 );
 a70031a <=( A232  and  A200 );
 a70032a <=( a70031a  and  a70028a );
 a70033a <=( a70032a  and  a70025a );
 a70037a <=( A236  and  A234 );
 a70038a <=( (not A233)  and  a70037a );
 a70041a <=( (not A299)  and  A298 );
 a70044a <=( A301  and  A300 );
 a70045a <=( a70044a  and  a70041a );
 a70046a <=( a70045a  and  a70038a );
 a70050a <=( (not A167)  and  (not A168) );
 a70051a <=( A169  and  a70050a );
 a70054a <=( (not A199)  and  A166 );
 a70057a <=( A232  and  A200 );
 a70058a <=( a70057a  and  a70054a );
 a70059a <=( a70058a  and  a70051a );
 a70063a <=( A236  and  A234 );
 a70064a <=( (not A233)  and  a70063a );
 a70067a <=( (not A299)  and  A298 );
 a70070a <=( A302  and  A300 );
 a70071a <=( a70070a  and  a70067a );
 a70072a <=( a70071a  and  a70064a );
 a70076a <=( (not A167)  and  (not A168) );
 a70077a <=( A169  and  a70076a );
 a70080a <=( (not A199)  and  A166 );
 a70083a <=( A232  and  A200 );
 a70084a <=( a70083a  and  a70080a );
 a70085a <=( a70084a  and  a70077a );
 a70089a <=( A236  and  A234 );
 a70090a <=( (not A233)  and  a70089a );
 a70093a <=( (not A266)  and  A265 );
 a70096a <=( A268  and  A267 );
 a70097a <=( a70096a  and  a70093a );
 a70098a <=( a70097a  and  a70090a );
 a70102a <=( (not A167)  and  (not A168) );
 a70103a <=( A169  and  a70102a );
 a70106a <=( (not A199)  and  A166 );
 a70109a <=( A232  and  A200 );
 a70110a <=( a70109a  and  a70106a );
 a70111a <=( a70110a  and  a70103a );
 a70115a <=( A236  and  A234 );
 a70116a <=( (not A233)  and  a70115a );
 a70119a <=( (not A266)  and  A265 );
 a70122a <=( A269  and  A267 );
 a70123a <=( a70122a  and  a70119a );
 a70124a <=( a70123a  and  a70116a );
 a70128a <=( (not A167)  and  (not A168) );
 a70129a <=( A169  and  a70128a );
 a70132a <=( (not A199)  and  A166 );
 a70135a <=( (not A232)  and  A200 );
 a70136a <=( a70135a  and  a70132a );
 a70137a <=( a70136a  and  a70129a );
 a70141a <=( (not A268)  and  (not A266) );
 a70142a <=( (not A233)  and  a70141a );
 a70145a <=( A298  and  (not A269) );
 a70148a <=( (not A302)  and  (not A301) );
 a70149a <=( a70148a  and  a70145a );
 a70150a <=( a70149a  and  a70142a );
 a70154a <=( (not A167)  and  (not A168) );
 a70155a <=( A169  and  a70154a );
 a70158a <=( A199  and  A166 );
 a70161a <=( A201  and  (not A200) );
 a70162a <=( a70161a  and  a70158a );
 a70163a <=( a70162a  and  a70155a );
 a70167a <=( A233  and  A232 );
 a70168a <=( A202  and  a70167a );
 a70171a <=( (not A267)  and  A265 );
 a70174a <=( (not A300)  and  (not A299) );
 a70175a <=( a70174a  and  a70171a );
 a70176a <=( a70175a  and  a70168a );
 a70180a <=( (not A167)  and  (not A168) );
 a70181a <=( A169  and  a70180a );
 a70184a <=( A199  and  A166 );
 a70187a <=( A201  and  (not A200) );
 a70188a <=( a70187a  and  a70184a );
 a70189a <=( a70188a  and  a70181a );
 a70193a <=( A233  and  A232 );
 a70194a <=( A202  and  a70193a );
 a70197a <=( (not A267)  and  A265 );
 a70200a <=( A299  and  A298 );
 a70201a <=( a70200a  and  a70197a );
 a70202a <=( a70201a  and  a70194a );
 a70206a <=( (not A167)  and  (not A168) );
 a70207a <=( A169  and  a70206a );
 a70210a <=( A199  and  A166 );
 a70213a <=( A201  and  (not A200) );
 a70214a <=( a70213a  and  a70210a );
 a70215a <=( a70214a  and  a70207a );
 a70219a <=( A233  and  A232 );
 a70220a <=( A202  and  a70219a );
 a70223a <=( (not A267)  and  A265 );
 a70226a <=( (not A299)  and  (not A298) );
 a70227a <=( a70226a  and  a70223a );
 a70228a <=( a70227a  and  a70220a );
 a70232a <=( (not A167)  and  (not A168) );
 a70233a <=( A169  and  a70232a );
 a70236a <=( A199  and  A166 );
 a70239a <=( A201  and  (not A200) );
 a70240a <=( a70239a  and  a70236a );
 a70241a <=( a70240a  and  a70233a );
 a70245a <=( A233  and  A232 );
 a70246a <=( A202  and  a70245a );
 a70249a <=( A266  and  A265 );
 a70252a <=( (not A300)  and  (not A299) );
 a70253a <=( a70252a  and  a70249a );
 a70254a <=( a70253a  and  a70246a );
 a70258a <=( (not A167)  and  (not A168) );
 a70259a <=( A169  and  a70258a );
 a70262a <=( A199  and  A166 );
 a70265a <=( A201  and  (not A200) );
 a70266a <=( a70265a  and  a70262a );
 a70267a <=( a70266a  and  a70259a );
 a70271a <=( A233  and  A232 );
 a70272a <=( A202  and  a70271a );
 a70275a <=( A266  and  A265 );
 a70278a <=( A299  and  A298 );
 a70279a <=( a70278a  and  a70275a );
 a70280a <=( a70279a  and  a70272a );
 a70284a <=( (not A167)  and  (not A168) );
 a70285a <=( A169  and  a70284a );
 a70288a <=( A199  and  A166 );
 a70291a <=( A201  and  (not A200) );
 a70292a <=( a70291a  and  a70288a );
 a70293a <=( a70292a  and  a70285a );
 a70297a <=( A233  and  A232 );
 a70298a <=( A202  and  a70297a );
 a70301a <=( A266  and  A265 );
 a70304a <=( (not A299)  and  (not A298) );
 a70305a <=( a70304a  and  a70301a );
 a70306a <=( a70305a  and  a70298a );
 a70310a <=( (not A167)  and  (not A168) );
 a70311a <=( A169  and  a70310a );
 a70314a <=( A199  and  A166 );
 a70317a <=( A201  and  (not A200) );
 a70318a <=( a70317a  and  a70314a );
 a70319a <=( a70318a  and  a70311a );
 a70323a <=( A233  and  A232 );
 a70324a <=( A202  and  a70323a );
 a70327a <=( (not A266)  and  (not A265) );
 a70330a <=( (not A300)  and  (not A299) );
 a70331a <=( a70330a  and  a70327a );
 a70332a <=( a70331a  and  a70324a );
 a70336a <=( (not A167)  and  (not A168) );
 a70337a <=( A169  and  a70336a );
 a70340a <=( A199  and  A166 );
 a70343a <=( A201  and  (not A200) );
 a70344a <=( a70343a  and  a70340a );
 a70345a <=( a70344a  and  a70337a );
 a70349a <=( A233  and  A232 );
 a70350a <=( A202  and  a70349a );
 a70353a <=( (not A266)  and  (not A265) );
 a70356a <=( A299  and  A298 );
 a70357a <=( a70356a  and  a70353a );
 a70358a <=( a70357a  and  a70350a );
 a70362a <=( (not A167)  and  (not A168) );
 a70363a <=( A169  and  a70362a );
 a70366a <=( A199  and  A166 );
 a70369a <=( A201  and  (not A200) );
 a70370a <=( a70369a  and  a70366a );
 a70371a <=( a70370a  and  a70363a );
 a70375a <=( A233  and  A232 );
 a70376a <=( A202  and  a70375a );
 a70379a <=( (not A266)  and  (not A265) );
 a70382a <=( (not A299)  and  (not A298) );
 a70383a <=( a70382a  and  a70379a );
 a70384a <=( a70383a  and  a70376a );
 a70388a <=( (not A167)  and  (not A168) );
 a70389a <=( A169  and  a70388a );
 a70392a <=( A199  and  A166 );
 a70395a <=( A201  and  (not A200) );
 a70396a <=( a70395a  and  a70392a );
 a70397a <=( a70396a  and  a70389a );
 a70401a <=( A233  and  (not A232) );
 a70402a <=( A202  and  a70401a );
 a70405a <=( (not A299)  and  A298 );
 a70408a <=( A301  and  A300 );
 a70409a <=( a70408a  and  a70405a );
 a70410a <=( a70409a  and  a70402a );
 a70414a <=( (not A167)  and  (not A168) );
 a70415a <=( A169  and  a70414a );
 a70418a <=( A199  and  A166 );
 a70421a <=( A201  and  (not A200) );
 a70422a <=( a70421a  and  a70418a );
 a70423a <=( a70422a  and  a70415a );
 a70427a <=( A233  and  (not A232) );
 a70428a <=( A202  and  a70427a );
 a70431a <=( (not A299)  and  A298 );
 a70434a <=( A302  and  A300 );
 a70435a <=( a70434a  and  a70431a );
 a70436a <=( a70435a  and  a70428a );
 a70440a <=( (not A167)  and  (not A168) );
 a70441a <=( A169  and  a70440a );
 a70444a <=( A199  and  A166 );
 a70447a <=( A201  and  (not A200) );
 a70448a <=( a70447a  and  a70444a );
 a70449a <=( a70448a  and  a70441a );
 a70453a <=( A233  and  (not A232) );
 a70454a <=( A202  and  a70453a );
 a70457a <=( (not A266)  and  A265 );
 a70460a <=( A268  and  A267 );
 a70461a <=( a70460a  and  a70457a );
 a70462a <=( a70461a  and  a70454a );
 a70466a <=( (not A167)  and  (not A168) );
 a70467a <=( A169  and  a70466a );
 a70470a <=( A199  and  A166 );
 a70473a <=( A201  and  (not A200) );
 a70474a <=( a70473a  and  a70470a );
 a70475a <=( a70474a  and  a70467a );
 a70479a <=( A233  and  (not A232) );
 a70480a <=( A202  and  a70479a );
 a70483a <=( (not A266)  and  A265 );
 a70486a <=( A269  and  A267 );
 a70487a <=( a70486a  and  a70483a );
 a70488a <=( a70487a  and  a70480a );
 a70492a <=( (not A167)  and  (not A168) );
 a70493a <=( A169  and  a70492a );
 a70496a <=( A199  and  A166 );
 a70499a <=( A201  and  (not A200) );
 a70500a <=( a70499a  and  a70496a );
 a70501a <=( a70500a  and  a70493a );
 a70505a <=( (not A234)  and  (not A233) );
 a70506a <=( A202  and  a70505a );
 a70509a <=( A266  and  A265 );
 a70512a <=( (not A300)  and  A298 );
 a70513a <=( a70512a  and  a70509a );
 a70514a <=( a70513a  and  a70506a );
 a70518a <=( (not A167)  and  (not A168) );
 a70519a <=( A169  and  a70518a );
 a70522a <=( A199  and  A166 );
 a70525a <=( A201  and  (not A200) );
 a70526a <=( a70525a  and  a70522a );
 a70527a <=( a70526a  and  a70519a );
 a70531a <=( (not A234)  and  (not A233) );
 a70532a <=( A202  and  a70531a );
 a70535a <=( A266  and  A265 );
 a70538a <=( A299  and  A298 );
 a70539a <=( a70538a  and  a70535a );
 a70540a <=( a70539a  and  a70532a );
 a70544a <=( (not A167)  and  (not A168) );
 a70545a <=( A169  and  a70544a );
 a70548a <=( A199  and  A166 );
 a70551a <=( A201  and  (not A200) );
 a70552a <=( a70551a  and  a70548a );
 a70553a <=( a70552a  and  a70545a );
 a70557a <=( (not A234)  and  (not A233) );
 a70558a <=( A202  and  a70557a );
 a70561a <=( A266  and  A265 );
 a70564a <=( (not A299)  and  (not A298) );
 a70565a <=( a70564a  and  a70561a );
 a70566a <=( a70565a  and  a70558a );
 a70570a <=( (not A167)  and  (not A168) );
 a70571a <=( A169  and  a70570a );
 a70574a <=( A199  and  A166 );
 a70577a <=( A201  and  (not A200) );
 a70578a <=( a70577a  and  a70574a );
 a70579a <=( a70578a  and  a70571a );
 a70583a <=( (not A234)  and  (not A233) );
 a70584a <=( A202  and  a70583a );
 a70587a <=( (not A267)  and  (not A266) );
 a70590a <=( (not A300)  and  A298 );
 a70591a <=( a70590a  and  a70587a );
 a70592a <=( a70591a  and  a70584a );
 a70596a <=( (not A167)  and  (not A168) );
 a70597a <=( A169  and  a70596a );
 a70600a <=( A199  and  A166 );
 a70603a <=( A201  and  (not A200) );
 a70604a <=( a70603a  and  a70600a );
 a70605a <=( a70604a  and  a70597a );
 a70609a <=( (not A234)  and  (not A233) );
 a70610a <=( A202  and  a70609a );
 a70613a <=( (not A267)  and  (not A266) );
 a70616a <=( A299  and  A298 );
 a70617a <=( a70616a  and  a70613a );
 a70618a <=( a70617a  and  a70610a );
 a70622a <=( (not A167)  and  (not A168) );
 a70623a <=( A169  and  a70622a );
 a70626a <=( A199  and  A166 );
 a70629a <=( A201  and  (not A200) );
 a70630a <=( a70629a  and  a70626a );
 a70631a <=( a70630a  and  a70623a );
 a70635a <=( (not A234)  and  (not A233) );
 a70636a <=( A202  and  a70635a );
 a70639a <=( (not A267)  and  (not A266) );
 a70642a <=( (not A299)  and  (not A298) );
 a70643a <=( a70642a  and  a70639a );
 a70644a <=( a70643a  and  a70636a );
 a70648a <=( (not A167)  and  (not A168) );
 a70649a <=( A169  and  a70648a );
 a70652a <=( A199  and  A166 );
 a70655a <=( A201  and  (not A200) );
 a70656a <=( a70655a  and  a70652a );
 a70657a <=( a70656a  and  a70649a );
 a70661a <=( (not A234)  and  (not A233) );
 a70662a <=( A202  and  a70661a );
 a70665a <=( (not A266)  and  (not A265) );
 a70668a <=( (not A300)  and  A298 );
 a70669a <=( a70668a  and  a70665a );
 a70670a <=( a70669a  and  a70662a );
 a70674a <=( (not A167)  and  (not A168) );
 a70675a <=( A169  and  a70674a );
 a70678a <=( A199  and  A166 );
 a70681a <=( A201  and  (not A200) );
 a70682a <=( a70681a  and  a70678a );
 a70683a <=( a70682a  and  a70675a );
 a70687a <=( (not A234)  and  (not A233) );
 a70688a <=( A202  and  a70687a );
 a70691a <=( (not A266)  and  (not A265) );
 a70694a <=( A299  and  A298 );
 a70695a <=( a70694a  and  a70691a );
 a70696a <=( a70695a  and  a70688a );
 a70700a <=( (not A167)  and  (not A168) );
 a70701a <=( A169  and  a70700a );
 a70704a <=( A199  and  A166 );
 a70707a <=( A201  and  (not A200) );
 a70708a <=( a70707a  and  a70704a );
 a70709a <=( a70708a  and  a70701a );
 a70713a <=( (not A234)  and  (not A233) );
 a70714a <=( A202  and  a70713a );
 a70717a <=( (not A266)  and  (not A265) );
 a70720a <=( (not A299)  and  (not A298) );
 a70721a <=( a70720a  and  a70717a );
 a70722a <=( a70721a  and  a70714a );
 a70726a <=( (not A167)  and  (not A168) );
 a70727a <=( A169  and  a70726a );
 a70730a <=( A199  and  A166 );
 a70733a <=( A201  and  (not A200) );
 a70734a <=( a70733a  and  a70730a );
 a70735a <=( a70734a  and  a70727a );
 a70739a <=( (not A233)  and  A232 );
 a70740a <=( A202  and  a70739a );
 a70743a <=( A235  and  A234 );
 a70746a <=( A299  and  (not A298) );
 a70747a <=( a70746a  and  a70743a );
 a70748a <=( a70747a  and  a70740a );
 a70752a <=( (not A167)  and  (not A168) );
 a70753a <=( A169  and  a70752a );
 a70756a <=( A199  and  A166 );
 a70759a <=( A201  and  (not A200) );
 a70760a <=( a70759a  and  a70756a );
 a70761a <=( a70760a  and  a70753a );
 a70765a <=( (not A233)  and  A232 );
 a70766a <=( A202  and  a70765a );
 a70769a <=( A235  and  A234 );
 a70772a <=( A266  and  (not A265) );
 a70773a <=( a70772a  and  a70769a );
 a70774a <=( a70773a  and  a70766a );
 a70778a <=( (not A167)  and  (not A168) );
 a70779a <=( A169  and  a70778a );
 a70782a <=( A199  and  A166 );
 a70785a <=( A201  and  (not A200) );
 a70786a <=( a70785a  and  a70782a );
 a70787a <=( a70786a  and  a70779a );
 a70791a <=( (not A233)  and  A232 );
 a70792a <=( A202  and  a70791a );
 a70795a <=( A236  and  A234 );
 a70798a <=( A299  and  (not A298) );
 a70799a <=( a70798a  and  a70795a );
 a70800a <=( a70799a  and  a70792a );
 a70804a <=( (not A167)  and  (not A168) );
 a70805a <=( A169  and  a70804a );
 a70808a <=( A199  and  A166 );
 a70811a <=( A201  and  (not A200) );
 a70812a <=( a70811a  and  a70808a );
 a70813a <=( a70812a  and  a70805a );
 a70817a <=( (not A233)  and  A232 );
 a70818a <=( A202  and  a70817a );
 a70821a <=( A236  and  A234 );
 a70824a <=( A266  and  (not A265) );
 a70825a <=( a70824a  and  a70821a );
 a70826a <=( a70825a  and  a70818a );
 a70830a <=( (not A167)  and  (not A168) );
 a70831a <=( A169  and  a70830a );
 a70834a <=( A199  and  A166 );
 a70837a <=( A201  and  (not A200) );
 a70838a <=( a70837a  and  a70834a );
 a70839a <=( a70838a  and  a70831a );
 a70843a <=( (not A233)  and  (not A232) );
 a70844a <=( A202  and  a70843a );
 a70847a <=( A266  and  A265 );
 a70850a <=( (not A300)  and  A298 );
 a70851a <=( a70850a  and  a70847a );
 a70852a <=( a70851a  and  a70844a );
 a70856a <=( (not A167)  and  (not A168) );
 a70857a <=( A169  and  a70856a );
 a70860a <=( A199  and  A166 );
 a70863a <=( A201  and  (not A200) );
 a70864a <=( a70863a  and  a70860a );
 a70865a <=( a70864a  and  a70857a );
 a70869a <=( (not A233)  and  (not A232) );
 a70870a <=( A202  and  a70869a );
 a70873a <=( A266  and  A265 );
 a70876a <=( A299  and  A298 );
 a70877a <=( a70876a  and  a70873a );
 a70878a <=( a70877a  and  a70870a );
 a70882a <=( (not A167)  and  (not A168) );
 a70883a <=( A169  and  a70882a );
 a70886a <=( A199  and  A166 );
 a70889a <=( A201  and  (not A200) );
 a70890a <=( a70889a  and  a70886a );
 a70891a <=( a70890a  and  a70883a );
 a70895a <=( (not A233)  and  (not A232) );
 a70896a <=( A202  and  a70895a );
 a70899a <=( A266  and  A265 );
 a70902a <=( (not A299)  and  (not A298) );
 a70903a <=( a70902a  and  a70899a );
 a70904a <=( a70903a  and  a70896a );
 a70908a <=( (not A167)  and  (not A168) );
 a70909a <=( A169  and  a70908a );
 a70912a <=( A199  and  A166 );
 a70915a <=( A201  and  (not A200) );
 a70916a <=( a70915a  and  a70912a );
 a70917a <=( a70916a  and  a70909a );
 a70921a <=( (not A233)  and  (not A232) );
 a70922a <=( A202  and  a70921a );
 a70925a <=( (not A267)  and  (not A266) );
 a70928a <=( (not A300)  and  A298 );
 a70929a <=( a70928a  and  a70925a );
 a70930a <=( a70929a  and  a70922a );
 a70934a <=( (not A167)  and  (not A168) );
 a70935a <=( A169  and  a70934a );
 a70938a <=( A199  and  A166 );
 a70941a <=( A201  and  (not A200) );
 a70942a <=( a70941a  and  a70938a );
 a70943a <=( a70942a  and  a70935a );
 a70947a <=( (not A233)  and  (not A232) );
 a70948a <=( A202  and  a70947a );
 a70951a <=( (not A267)  and  (not A266) );
 a70954a <=( A299  and  A298 );
 a70955a <=( a70954a  and  a70951a );
 a70956a <=( a70955a  and  a70948a );
 a70960a <=( (not A167)  and  (not A168) );
 a70961a <=( A169  and  a70960a );
 a70964a <=( A199  and  A166 );
 a70967a <=( A201  and  (not A200) );
 a70968a <=( a70967a  and  a70964a );
 a70969a <=( a70968a  and  a70961a );
 a70973a <=( (not A233)  and  (not A232) );
 a70974a <=( A202  and  a70973a );
 a70977a <=( (not A267)  and  (not A266) );
 a70980a <=( (not A299)  and  (not A298) );
 a70981a <=( a70980a  and  a70977a );
 a70982a <=( a70981a  and  a70974a );
 a70986a <=( (not A167)  and  (not A168) );
 a70987a <=( A169  and  a70986a );
 a70990a <=( A199  and  A166 );
 a70993a <=( A201  and  (not A200) );
 a70994a <=( a70993a  and  a70990a );
 a70995a <=( a70994a  and  a70987a );
 a70999a <=( (not A233)  and  (not A232) );
 a71000a <=( A202  and  a70999a );
 a71003a <=( (not A266)  and  (not A265) );
 a71006a <=( (not A300)  and  A298 );
 a71007a <=( a71006a  and  a71003a );
 a71008a <=( a71007a  and  a71000a );
 a71012a <=( (not A167)  and  (not A168) );
 a71013a <=( A169  and  a71012a );
 a71016a <=( A199  and  A166 );
 a71019a <=( A201  and  (not A200) );
 a71020a <=( a71019a  and  a71016a );
 a71021a <=( a71020a  and  a71013a );
 a71025a <=( (not A233)  and  (not A232) );
 a71026a <=( A202  and  a71025a );
 a71029a <=( (not A266)  and  (not A265) );
 a71032a <=( A299  and  A298 );
 a71033a <=( a71032a  and  a71029a );
 a71034a <=( a71033a  and  a71026a );
 a71038a <=( (not A167)  and  (not A168) );
 a71039a <=( A169  and  a71038a );
 a71042a <=( A199  and  A166 );
 a71045a <=( A201  and  (not A200) );
 a71046a <=( a71045a  and  a71042a );
 a71047a <=( a71046a  and  a71039a );
 a71051a <=( (not A233)  and  (not A232) );
 a71052a <=( A202  and  a71051a );
 a71055a <=( (not A266)  and  (not A265) );
 a71058a <=( (not A299)  and  (not A298) );
 a71059a <=( a71058a  and  a71055a );
 a71060a <=( a71059a  and  a71052a );
 a71064a <=( (not A167)  and  (not A168) );
 a71065a <=( A169  and  a71064a );
 a71068a <=( A199  and  A166 );
 a71071a <=( A201  and  (not A200) );
 a71072a <=( a71071a  and  a71068a );
 a71073a <=( a71072a  and  a71065a );
 a71077a <=( A233  and  A232 );
 a71078a <=( A203  and  a71077a );
 a71081a <=( (not A267)  and  A265 );
 a71084a <=( (not A300)  and  (not A299) );
 a71085a <=( a71084a  and  a71081a );
 a71086a <=( a71085a  and  a71078a );
 a71090a <=( (not A167)  and  (not A168) );
 a71091a <=( A169  and  a71090a );
 a71094a <=( A199  and  A166 );
 a71097a <=( A201  and  (not A200) );
 a71098a <=( a71097a  and  a71094a );
 a71099a <=( a71098a  and  a71091a );
 a71103a <=( A233  and  A232 );
 a71104a <=( A203  and  a71103a );
 a71107a <=( (not A267)  and  A265 );
 a71110a <=( A299  and  A298 );
 a71111a <=( a71110a  and  a71107a );
 a71112a <=( a71111a  and  a71104a );
 a71116a <=( (not A167)  and  (not A168) );
 a71117a <=( A169  and  a71116a );
 a71120a <=( A199  and  A166 );
 a71123a <=( A201  and  (not A200) );
 a71124a <=( a71123a  and  a71120a );
 a71125a <=( a71124a  and  a71117a );
 a71129a <=( A233  and  A232 );
 a71130a <=( A203  and  a71129a );
 a71133a <=( (not A267)  and  A265 );
 a71136a <=( (not A299)  and  (not A298) );
 a71137a <=( a71136a  and  a71133a );
 a71138a <=( a71137a  and  a71130a );
 a71142a <=( (not A167)  and  (not A168) );
 a71143a <=( A169  and  a71142a );
 a71146a <=( A199  and  A166 );
 a71149a <=( A201  and  (not A200) );
 a71150a <=( a71149a  and  a71146a );
 a71151a <=( a71150a  and  a71143a );
 a71155a <=( A233  and  A232 );
 a71156a <=( A203  and  a71155a );
 a71159a <=( A266  and  A265 );
 a71162a <=( (not A300)  and  (not A299) );
 a71163a <=( a71162a  and  a71159a );
 a71164a <=( a71163a  and  a71156a );
 a71168a <=( (not A167)  and  (not A168) );
 a71169a <=( A169  and  a71168a );
 a71172a <=( A199  and  A166 );
 a71175a <=( A201  and  (not A200) );
 a71176a <=( a71175a  and  a71172a );
 a71177a <=( a71176a  and  a71169a );
 a71181a <=( A233  and  A232 );
 a71182a <=( A203  and  a71181a );
 a71185a <=( A266  and  A265 );
 a71188a <=( A299  and  A298 );
 a71189a <=( a71188a  and  a71185a );
 a71190a <=( a71189a  and  a71182a );
 a71194a <=( (not A167)  and  (not A168) );
 a71195a <=( A169  and  a71194a );
 a71198a <=( A199  and  A166 );
 a71201a <=( A201  and  (not A200) );
 a71202a <=( a71201a  and  a71198a );
 a71203a <=( a71202a  and  a71195a );
 a71207a <=( A233  and  A232 );
 a71208a <=( A203  and  a71207a );
 a71211a <=( A266  and  A265 );
 a71214a <=( (not A299)  and  (not A298) );
 a71215a <=( a71214a  and  a71211a );
 a71216a <=( a71215a  and  a71208a );
 a71220a <=( (not A167)  and  (not A168) );
 a71221a <=( A169  and  a71220a );
 a71224a <=( A199  and  A166 );
 a71227a <=( A201  and  (not A200) );
 a71228a <=( a71227a  and  a71224a );
 a71229a <=( a71228a  and  a71221a );
 a71233a <=( A233  and  A232 );
 a71234a <=( A203  and  a71233a );
 a71237a <=( (not A266)  and  (not A265) );
 a71240a <=( (not A300)  and  (not A299) );
 a71241a <=( a71240a  and  a71237a );
 a71242a <=( a71241a  and  a71234a );
 a71246a <=( (not A167)  and  (not A168) );
 a71247a <=( A169  and  a71246a );
 a71250a <=( A199  and  A166 );
 a71253a <=( A201  and  (not A200) );
 a71254a <=( a71253a  and  a71250a );
 a71255a <=( a71254a  and  a71247a );
 a71259a <=( A233  and  A232 );
 a71260a <=( A203  and  a71259a );
 a71263a <=( (not A266)  and  (not A265) );
 a71266a <=( A299  and  A298 );
 a71267a <=( a71266a  and  a71263a );
 a71268a <=( a71267a  and  a71260a );
 a71272a <=( (not A167)  and  (not A168) );
 a71273a <=( A169  and  a71272a );
 a71276a <=( A199  and  A166 );
 a71279a <=( A201  and  (not A200) );
 a71280a <=( a71279a  and  a71276a );
 a71281a <=( a71280a  and  a71273a );
 a71285a <=( A233  and  A232 );
 a71286a <=( A203  and  a71285a );
 a71289a <=( (not A266)  and  (not A265) );
 a71292a <=( (not A299)  and  (not A298) );
 a71293a <=( a71292a  and  a71289a );
 a71294a <=( a71293a  and  a71286a );
 a71298a <=( (not A167)  and  (not A168) );
 a71299a <=( A169  and  a71298a );
 a71302a <=( A199  and  A166 );
 a71305a <=( A201  and  (not A200) );
 a71306a <=( a71305a  and  a71302a );
 a71307a <=( a71306a  and  a71299a );
 a71311a <=( A233  and  (not A232) );
 a71312a <=( A203  and  a71311a );
 a71315a <=( (not A299)  and  A298 );
 a71318a <=( A301  and  A300 );
 a71319a <=( a71318a  and  a71315a );
 a71320a <=( a71319a  and  a71312a );
 a71324a <=( (not A167)  and  (not A168) );
 a71325a <=( A169  and  a71324a );
 a71328a <=( A199  and  A166 );
 a71331a <=( A201  and  (not A200) );
 a71332a <=( a71331a  and  a71328a );
 a71333a <=( a71332a  and  a71325a );
 a71337a <=( A233  and  (not A232) );
 a71338a <=( A203  and  a71337a );
 a71341a <=( (not A299)  and  A298 );
 a71344a <=( A302  and  A300 );
 a71345a <=( a71344a  and  a71341a );
 a71346a <=( a71345a  and  a71338a );
 a71350a <=( (not A167)  and  (not A168) );
 a71351a <=( A169  and  a71350a );
 a71354a <=( A199  and  A166 );
 a71357a <=( A201  and  (not A200) );
 a71358a <=( a71357a  and  a71354a );
 a71359a <=( a71358a  and  a71351a );
 a71363a <=( A233  and  (not A232) );
 a71364a <=( A203  and  a71363a );
 a71367a <=( (not A266)  and  A265 );
 a71370a <=( A268  and  A267 );
 a71371a <=( a71370a  and  a71367a );
 a71372a <=( a71371a  and  a71364a );
 a71376a <=( (not A167)  and  (not A168) );
 a71377a <=( A169  and  a71376a );
 a71380a <=( A199  and  A166 );
 a71383a <=( A201  and  (not A200) );
 a71384a <=( a71383a  and  a71380a );
 a71385a <=( a71384a  and  a71377a );
 a71389a <=( A233  and  (not A232) );
 a71390a <=( A203  and  a71389a );
 a71393a <=( (not A266)  and  A265 );
 a71396a <=( A269  and  A267 );
 a71397a <=( a71396a  and  a71393a );
 a71398a <=( a71397a  and  a71390a );
 a71402a <=( (not A167)  and  (not A168) );
 a71403a <=( A169  and  a71402a );
 a71406a <=( A199  and  A166 );
 a71409a <=( A201  and  (not A200) );
 a71410a <=( a71409a  and  a71406a );
 a71411a <=( a71410a  and  a71403a );
 a71415a <=( (not A234)  and  (not A233) );
 a71416a <=( A203  and  a71415a );
 a71419a <=( A266  and  A265 );
 a71422a <=( (not A300)  and  A298 );
 a71423a <=( a71422a  and  a71419a );
 a71424a <=( a71423a  and  a71416a );
 a71428a <=( (not A167)  and  (not A168) );
 a71429a <=( A169  and  a71428a );
 a71432a <=( A199  and  A166 );
 a71435a <=( A201  and  (not A200) );
 a71436a <=( a71435a  and  a71432a );
 a71437a <=( a71436a  and  a71429a );
 a71441a <=( (not A234)  and  (not A233) );
 a71442a <=( A203  and  a71441a );
 a71445a <=( A266  and  A265 );
 a71448a <=( A299  and  A298 );
 a71449a <=( a71448a  and  a71445a );
 a71450a <=( a71449a  and  a71442a );
 a71454a <=( (not A167)  and  (not A168) );
 a71455a <=( A169  and  a71454a );
 a71458a <=( A199  and  A166 );
 a71461a <=( A201  and  (not A200) );
 a71462a <=( a71461a  and  a71458a );
 a71463a <=( a71462a  and  a71455a );
 a71467a <=( (not A234)  and  (not A233) );
 a71468a <=( A203  and  a71467a );
 a71471a <=( A266  and  A265 );
 a71474a <=( (not A299)  and  (not A298) );
 a71475a <=( a71474a  and  a71471a );
 a71476a <=( a71475a  and  a71468a );
 a71480a <=( (not A167)  and  (not A168) );
 a71481a <=( A169  and  a71480a );
 a71484a <=( A199  and  A166 );
 a71487a <=( A201  and  (not A200) );
 a71488a <=( a71487a  and  a71484a );
 a71489a <=( a71488a  and  a71481a );
 a71493a <=( (not A234)  and  (not A233) );
 a71494a <=( A203  and  a71493a );
 a71497a <=( (not A267)  and  (not A266) );
 a71500a <=( (not A300)  and  A298 );
 a71501a <=( a71500a  and  a71497a );
 a71502a <=( a71501a  and  a71494a );
 a71506a <=( (not A167)  and  (not A168) );
 a71507a <=( A169  and  a71506a );
 a71510a <=( A199  and  A166 );
 a71513a <=( A201  and  (not A200) );
 a71514a <=( a71513a  and  a71510a );
 a71515a <=( a71514a  and  a71507a );
 a71519a <=( (not A234)  and  (not A233) );
 a71520a <=( A203  and  a71519a );
 a71523a <=( (not A267)  and  (not A266) );
 a71526a <=( A299  and  A298 );
 a71527a <=( a71526a  and  a71523a );
 a71528a <=( a71527a  and  a71520a );
 a71532a <=( (not A167)  and  (not A168) );
 a71533a <=( A169  and  a71532a );
 a71536a <=( A199  and  A166 );
 a71539a <=( A201  and  (not A200) );
 a71540a <=( a71539a  and  a71536a );
 a71541a <=( a71540a  and  a71533a );
 a71545a <=( (not A234)  and  (not A233) );
 a71546a <=( A203  and  a71545a );
 a71549a <=( (not A267)  and  (not A266) );
 a71552a <=( (not A299)  and  (not A298) );
 a71553a <=( a71552a  and  a71549a );
 a71554a <=( a71553a  and  a71546a );
 a71558a <=( (not A167)  and  (not A168) );
 a71559a <=( A169  and  a71558a );
 a71562a <=( A199  and  A166 );
 a71565a <=( A201  and  (not A200) );
 a71566a <=( a71565a  and  a71562a );
 a71567a <=( a71566a  and  a71559a );
 a71571a <=( (not A234)  and  (not A233) );
 a71572a <=( A203  and  a71571a );
 a71575a <=( (not A266)  and  (not A265) );
 a71578a <=( (not A300)  and  A298 );
 a71579a <=( a71578a  and  a71575a );
 a71580a <=( a71579a  and  a71572a );
 a71584a <=( (not A167)  and  (not A168) );
 a71585a <=( A169  and  a71584a );
 a71588a <=( A199  and  A166 );
 a71591a <=( A201  and  (not A200) );
 a71592a <=( a71591a  and  a71588a );
 a71593a <=( a71592a  and  a71585a );
 a71597a <=( (not A234)  and  (not A233) );
 a71598a <=( A203  and  a71597a );
 a71601a <=( (not A266)  and  (not A265) );
 a71604a <=( A299  and  A298 );
 a71605a <=( a71604a  and  a71601a );
 a71606a <=( a71605a  and  a71598a );
 a71610a <=( (not A167)  and  (not A168) );
 a71611a <=( A169  and  a71610a );
 a71614a <=( A199  and  A166 );
 a71617a <=( A201  and  (not A200) );
 a71618a <=( a71617a  and  a71614a );
 a71619a <=( a71618a  and  a71611a );
 a71623a <=( (not A234)  and  (not A233) );
 a71624a <=( A203  and  a71623a );
 a71627a <=( (not A266)  and  (not A265) );
 a71630a <=( (not A299)  and  (not A298) );
 a71631a <=( a71630a  and  a71627a );
 a71632a <=( a71631a  and  a71624a );
 a71636a <=( (not A167)  and  (not A168) );
 a71637a <=( A169  and  a71636a );
 a71640a <=( A199  and  A166 );
 a71643a <=( A201  and  (not A200) );
 a71644a <=( a71643a  and  a71640a );
 a71645a <=( a71644a  and  a71637a );
 a71649a <=( (not A233)  and  A232 );
 a71650a <=( A203  and  a71649a );
 a71653a <=( A235  and  A234 );
 a71656a <=( A299  and  (not A298) );
 a71657a <=( a71656a  and  a71653a );
 a71658a <=( a71657a  and  a71650a );
 a71662a <=( (not A167)  and  (not A168) );
 a71663a <=( A169  and  a71662a );
 a71666a <=( A199  and  A166 );
 a71669a <=( A201  and  (not A200) );
 a71670a <=( a71669a  and  a71666a );
 a71671a <=( a71670a  and  a71663a );
 a71675a <=( (not A233)  and  A232 );
 a71676a <=( A203  and  a71675a );
 a71679a <=( A235  and  A234 );
 a71682a <=( A266  and  (not A265) );
 a71683a <=( a71682a  and  a71679a );
 a71684a <=( a71683a  and  a71676a );
 a71688a <=( (not A167)  and  (not A168) );
 a71689a <=( A169  and  a71688a );
 a71692a <=( A199  and  A166 );
 a71695a <=( A201  and  (not A200) );
 a71696a <=( a71695a  and  a71692a );
 a71697a <=( a71696a  and  a71689a );
 a71701a <=( (not A233)  and  A232 );
 a71702a <=( A203  and  a71701a );
 a71705a <=( A236  and  A234 );
 a71708a <=( A299  and  (not A298) );
 a71709a <=( a71708a  and  a71705a );
 a71710a <=( a71709a  and  a71702a );
 a71714a <=( (not A167)  and  (not A168) );
 a71715a <=( A169  and  a71714a );
 a71718a <=( A199  and  A166 );
 a71721a <=( A201  and  (not A200) );
 a71722a <=( a71721a  and  a71718a );
 a71723a <=( a71722a  and  a71715a );
 a71727a <=( (not A233)  and  A232 );
 a71728a <=( A203  and  a71727a );
 a71731a <=( A236  and  A234 );
 a71734a <=( A266  and  (not A265) );
 a71735a <=( a71734a  and  a71731a );
 a71736a <=( a71735a  and  a71728a );
 a71740a <=( (not A167)  and  (not A168) );
 a71741a <=( A169  and  a71740a );
 a71744a <=( A199  and  A166 );
 a71747a <=( A201  and  (not A200) );
 a71748a <=( a71747a  and  a71744a );
 a71749a <=( a71748a  and  a71741a );
 a71753a <=( (not A233)  and  (not A232) );
 a71754a <=( A203  and  a71753a );
 a71757a <=( A266  and  A265 );
 a71760a <=( (not A300)  and  A298 );
 a71761a <=( a71760a  and  a71757a );
 a71762a <=( a71761a  and  a71754a );
 a71766a <=( (not A167)  and  (not A168) );
 a71767a <=( A169  and  a71766a );
 a71770a <=( A199  and  A166 );
 a71773a <=( A201  and  (not A200) );
 a71774a <=( a71773a  and  a71770a );
 a71775a <=( a71774a  and  a71767a );
 a71779a <=( (not A233)  and  (not A232) );
 a71780a <=( A203  and  a71779a );
 a71783a <=( A266  and  A265 );
 a71786a <=( A299  and  A298 );
 a71787a <=( a71786a  and  a71783a );
 a71788a <=( a71787a  and  a71780a );
 a71792a <=( (not A167)  and  (not A168) );
 a71793a <=( A169  and  a71792a );
 a71796a <=( A199  and  A166 );
 a71799a <=( A201  and  (not A200) );
 a71800a <=( a71799a  and  a71796a );
 a71801a <=( a71800a  and  a71793a );
 a71805a <=( (not A233)  and  (not A232) );
 a71806a <=( A203  and  a71805a );
 a71809a <=( A266  and  A265 );
 a71812a <=( (not A299)  and  (not A298) );
 a71813a <=( a71812a  and  a71809a );
 a71814a <=( a71813a  and  a71806a );
 a71818a <=( (not A167)  and  (not A168) );
 a71819a <=( A169  and  a71818a );
 a71822a <=( A199  and  A166 );
 a71825a <=( A201  and  (not A200) );
 a71826a <=( a71825a  and  a71822a );
 a71827a <=( a71826a  and  a71819a );
 a71831a <=( (not A233)  and  (not A232) );
 a71832a <=( A203  and  a71831a );
 a71835a <=( (not A267)  and  (not A266) );
 a71838a <=( (not A300)  and  A298 );
 a71839a <=( a71838a  and  a71835a );
 a71840a <=( a71839a  and  a71832a );
 a71844a <=( (not A167)  and  (not A168) );
 a71845a <=( A169  and  a71844a );
 a71848a <=( A199  and  A166 );
 a71851a <=( A201  and  (not A200) );
 a71852a <=( a71851a  and  a71848a );
 a71853a <=( a71852a  and  a71845a );
 a71857a <=( (not A233)  and  (not A232) );
 a71858a <=( A203  and  a71857a );
 a71861a <=( (not A267)  and  (not A266) );
 a71864a <=( A299  and  A298 );
 a71865a <=( a71864a  and  a71861a );
 a71866a <=( a71865a  and  a71858a );
 a71870a <=( (not A167)  and  (not A168) );
 a71871a <=( A169  and  a71870a );
 a71874a <=( A199  and  A166 );
 a71877a <=( A201  and  (not A200) );
 a71878a <=( a71877a  and  a71874a );
 a71879a <=( a71878a  and  a71871a );
 a71883a <=( (not A233)  and  (not A232) );
 a71884a <=( A203  and  a71883a );
 a71887a <=( (not A267)  and  (not A266) );
 a71890a <=( (not A299)  and  (not A298) );
 a71891a <=( a71890a  and  a71887a );
 a71892a <=( a71891a  and  a71884a );
 a71896a <=( (not A167)  and  (not A168) );
 a71897a <=( A169  and  a71896a );
 a71900a <=( A199  and  A166 );
 a71903a <=( A201  and  (not A200) );
 a71904a <=( a71903a  and  a71900a );
 a71905a <=( a71904a  and  a71897a );
 a71909a <=( (not A233)  and  (not A232) );
 a71910a <=( A203  and  a71909a );
 a71913a <=( (not A266)  and  (not A265) );
 a71916a <=( (not A300)  and  A298 );
 a71917a <=( a71916a  and  a71913a );
 a71918a <=( a71917a  and  a71910a );
 a71922a <=( (not A167)  and  (not A168) );
 a71923a <=( A169  and  a71922a );
 a71926a <=( A199  and  A166 );
 a71929a <=( A201  and  (not A200) );
 a71930a <=( a71929a  and  a71926a );
 a71931a <=( a71930a  and  a71923a );
 a71935a <=( (not A233)  and  (not A232) );
 a71936a <=( A203  and  a71935a );
 a71939a <=( (not A266)  and  (not A265) );
 a71942a <=( A299  and  A298 );
 a71943a <=( a71942a  and  a71939a );
 a71944a <=( a71943a  and  a71936a );
 a71948a <=( (not A167)  and  (not A168) );
 a71949a <=( A169  and  a71948a );
 a71952a <=( A199  and  A166 );
 a71955a <=( A201  and  (not A200) );
 a71956a <=( a71955a  and  a71952a );
 a71957a <=( a71956a  and  a71949a );
 a71961a <=( (not A233)  and  (not A232) );
 a71962a <=( A203  and  a71961a );
 a71965a <=( (not A266)  and  (not A265) );
 a71968a <=( (not A299)  and  (not A298) );
 a71969a <=( a71968a  and  a71965a );
 a71970a <=( a71969a  and  a71962a );
 a71974a <=( (not A168)  and  A169 );
 a71975a <=( A170  and  a71974a );
 a71978a <=( (not A200)  and  A199 );
 a71981a <=( A202  and  A201 );
 a71982a <=( a71981a  and  a71978a );
 a71983a <=( a71982a  and  a71975a );
 a71987a <=( A265  and  A233 );
 a71988a <=( A232  and  a71987a );
 a71991a <=( (not A269)  and  (not A268) );
 a71994a <=( (not A300)  and  (not A299) );
 a71995a <=( a71994a  and  a71991a );
 a71996a <=( a71995a  and  a71988a );
 a72000a <=( (not A168)  and  A169 );
 a72001a <=( A170  and  a72000a );
 a72004a <=( (not A200)  and  A199 );
 a72007a <=( A202  and  A201 );
 a72008a <=( a72007a  and  a72004a );
 a72009a <=( a72008a  and  a72001a );
 a72013a <=( A265  and  A233 );
 a72014a <=( A232  and  a72013a );
 a72017a <=( (not A269)  and  (not A268) );
 a72020a <=( A299  and  A298 );
 a72021a <=( a72020a  and  a72017a );
 a72022a <=( a72021a  and  a72014a );
 a72026a <=( (not A168)  and  A169 );
 a72027a <=( A170  and  a72026a );
 a72030a <=( (not A200)  and  A199 );
 a72033a <=( A202  and  A201 );
 a72034a <=( a72033a  and  a72030a );
 a72035a <=( a72034a  and  a72027a );
 a72039a <=( A265  and  A233 );
 a72040a <=( A232  and  a72039a );
 a72043a <=( (not A269)  and  (not A268) );
 a72046a <=( (not A299)  and  (not A298) );
 a72047a <=( a72046a  and  a72043a );
 a72048a <=( a72047a  and  a72040a );
 a72052a <=( (not A168)  and  A169 );
 a72053a <=( A170  and  a72052a );
 a72056a <=( (not A200)  and  A199 );
 a72059a <=( A202  and  A201 );
 a72060a <=( a72059a  and  a72056a );
 a72061a <=( a72060a  and  a72053a );
 a72065a <=( A265  and  A233 );
 a72066a <=( A232  and  a72065a );
 a72069a <=( (not A299)  and  (not A267) );
 a72072a <=( (not A302)  and  (not A301) );
 a72073a <=( a72072a  and  a72069a );
 a72074a <=( a72073a  and  a72066a );
 a72078a <=( (not A168)  and  A169 );
 a72079a <=( A170  and  a72078a );
 a72082a <=( (not A200)  and  A199 );
 a72085a <=( A202  and  A201 );
 a72086a <=( a72085a  and  a72082a );
 a72087a <=( a72086a  and  a72079a );
 a72091a <=( A265  and  A233 );
 a72092a <=( A232  and  a72091a );
 a72095a <=( (not A299)  and  A266 );
 a72098a <=( (not A302)  and  (not A301) );
 a72099a <=( a72098a  and  a72095a );
 a72100a <=( a72099a  and  a72092a );
 a72104a <=( (not A168)  and  A169 );
 a72105a <=( A170  and  a72104a );
 a72108a <=( (not A200)  and  A199 );
 a72111a <=( A202  and  A201 );
 a72112a <=( a72111a  and  a72108a );
 a72113a <=( a72112a  and  a72105a );
 a72117a <=( (not A265)  and  A233 );
 a72118a <=( A232  and  a72117a );
 a72121a <=( (not A299)  and  (not A266) );
 a72124a <=( (not A302)  and  (not A301) );
 a72125a <=( a72124a  and  a72121a );
 a72126a <=( a72125a  and  a72118a );
 a72130a <=( (not A168)  and  A169 );
 a72131a <=( A170  and  a72130a );
 a72134a <=( (not A200)  and  A199 );
 a72137a <=( A202  and  A201 );
 a72138a <=( a72137a  and  a72134a );
 a72139a <=( a72138a  and  a72131a );
 a72143a <=( (not A236)  and  (not A235) );
 a72144a <=( (not A233)  and  a72143a );
 a72147a <=( A266  and  A265 );
 a72150a <=( (not A300)  and  A298 );
 a72151a <=( a72150a  and  a72147a );
 a72152a <=( a72151a  and  a72144a );
 a72156a <=( (not A168)  and  A169 );
 a72157a <=( A170  and  a72156a );
 a72160a <=( (not A200)  and  A199 );
 a72163a <=( A202  and  A201 );
 a72164a <=( a72163a  and  a72160a );
 a72165a <=( a72164a  and  a72157a );
 a72169a <=( (not A236)  and  (not A235) );
 a72170a <=( (not A233)  and  a72169a );
 a72173a <=( A266  and  A265 );
 a72176a <=( A299  and  A298 );
 a72177a <=( a72176a  and  a72173a );
 a72178a <=( a72177a  and  a72170a );
 a72182a <=( (not A168)  and  A169 );
 a72183a <=( A170  and  a72182a );
 a72186a <=( (not A200)  and  A199 );
 a72189a <=( A202  and  A201 );
 a72190a <=( a72189a  and  a72186a );
 a72191a <=( a72190a  and  a72183a );
 a72195a <=( (not A236)  and  (not A235) );
 a72196a <=( (not A233)  and  a72195a );
 a72199a <=( A266  and  A265 );
 a72202a <=( (not A299)  and  (not A298) );
 a72203a <=( a72202a  and  a72199a );
 a72204a <=( a72203a  and  a72196a );
 a72208a <=( (not A168)  and  A169 );
 a72209a <=( A170  and  a72208a );
 a72212a <=( (not A200)  and  A199 );
 a72215a <=( A202  and  A201 );
 a72216a <=( a72215a  and  a72212a );
 a72217a <=( a72216a  and  a72209a );
 a72221a <=( (not A236)  and  (not A235) );
 a72222a <=( (not A233)  and  a72221a );
 a72225a <=( (not A267)  and  (not A266) );
 a72228a <=( (not A300)  and  A298 );
 a72229a <=( a72228a  and  a72225a );
 a72230a <=( a72229a  and  a72222a );
 a72234a <=( (not A168)  and  A169 );
 a72235a <=( A170  and  a72234a );
 a72238a <=( (not A200)  and  A199 );
 a72241a <=( A202  and  A201 );
 a72242a <=( a72241a  and  a72238a );
 a72243a <=( a72242a  and  a72235a );
 a72247a <=( (not A236)  and  (not A235) );
 a72248a <=( (not A233)  and  a72247a );
 a72251a <=( (not A267)  and  (not A266) );
 a72254a <=( A299  and  A298 );
 a72255a <=( a72254a  and  a72251a );
 a72256a <=( a72255a  and  a72248a );
 a72260a <=( (not A168)  and  A169 );
 a72261a <=( A170  and  a72260a );
 a72264a <=( (not A200)  and  A199 );
 a72267a <=( A202  and  A201 );
 a72268a <=( a72267a  and  a72264a );
 a72269a <=( a72268a  and  a72261a );
 a72273a <=( (not A236)  and  (not A235) );
 a72274a <=( (not A233)  and  a72273a );
 a72277a <=( (not A267)  and  (not A266) );
 a72280a <=( (not A299)  and  (not A298) );
 a72281a <=( a72280a  and  a72277a );
 a72282a <=( a72281a  and  a72274a );
 a72286a <=( (not A168)  and  A169 );
 a72287a <=( A170  and  a72286a );
 a72290a <=( (not A200)  and  A199 );
 a72293a <=( A202  and  A201 );
 a72294a <=( a72293a  and  a72290a );
 a72295a <=( a72294a  and  a72287a );
 a72299a <=( (not A236)  and  (not A235) );
 a72300a <=( (not A233)  and  a72299a );
 a72303a <=( (not A266)  and  (not A265) );
 a72306a <=( (not A300)  and  A298 );
 a72307a <=( a72306a  and  a72303a );
 a72308a <=( a72307a  and  a72300a );
 a72312a <=( (not A168)  and  A169 );
 a72313a <=( A170  and  a72312a );
 a72316a <=( (not A200)  and  A199 );
 a72319a <=( A202  and  A201 );
 a72320a <=( a72319a  and  a72316a );
 a72321a <=( a72320a  and  a72313a );
 a72325a <=( (not A236)  and  (not A235) );
 a72326a <=( (not A233)  and  a72325a );
 a72329a <=( (not A266)  and  (not A265) );
 a72332a <=( A299  and  A298 );
 a72333a <=( a72332a  and  a72329a );
 a72334a <=( a72333a  and  a72326a );
 a72338a <=( (not A168)  and  A169 );
 a72339a <=( A170  and  a72338a );
 a72342a <=( (not A200)  and  A199 );
 a72345a <=( A202  and  A201 );
 a72346a <=( a72345a  and  a72342a );
 a72347a <=( a72346a  and  a72339a );
 a72351a <=( (not A236)  and  (not A235) );
 a72352a <=( (not A233)  and  a72351a );
 a72355a <=( (not A266)  and  (not A265) );
 a72358a <=( (not A299)  and  (not A298) );
 a72359a <=( a72358a  and  a72355a );
 a72360a <=( a72359a  and  a72352a );
 a72364a <=( (not A168)  and  A169 );
 a72365a <=( A170  and  a72364a );
 a72368a <=( (not A200)  and  A199 );
 a72371a <=( A202  and  A201 );
 a72372a <=( a72371a  and  a72368a );
 a72373a <=( a72372a  and  a72365a );
 a72377a <=( A265  and  (not A234) );
 a72378a <=( (not A233)  and  a72377a );
 a72381a <=( A298  and  A266 );
 a72384a <=( (not A302)  and  (not A301) );
 a72385a <=( a72384a  and  a72381a );
 a72386a <=( a72385a  and  a72378a );
 a72390a <=( (not A168)  and  A169 );
 a72391a <=( A170  and  a72390a );
 a72394a <=( (not A200)  and  A199 );
 a72397a <=( A202  and  A201 );
 a72398a <=( a72397a  and  a72394a );
 a72399a <=( a72398a  and  a72391a );
 a72403a <=( (not A266)  and  (not A234) );
 a72404a <=( (not A233)  and  a72403a );
 a72407a <=( (not A269)  and  (not A268) );
 a72410a <=( (not A300)  and  A298 );
 a72411a <=( a72410a  and  a72407a );
 a72412a <=( a72411a  and  a72404a );
 a72416a <=( (not A168)  and  A169 );
 a72417a <=( A170  and  a72416a );
 a72420a <=( (not A200)  and  A199 );
 a72423a <=( A202  and  A201 );
 a72424a <=( a72423a  and  a72420a );
 a72425a <=( a72424a  and  a72417a );
 a72429a <=( (not A266)  and  (not A234) );
 a72430a <=( (not A233)  and  a72429a );
 a72433a <=( (not A269)  and  (not A268) );
 a72436a <=( A299  and  A298 );
 a72437a <=( a72436a  and  a72433a );
 a72438a <=( a72437a  and  a72430a );
 a72442a <=( (not A168)  and  A169 );
 a72443a <=( A170  and  a72442a );
 a72446a <=( (not A200)  and  A199 );
 a72449a <=( A202  and  A201 );
 a72450a <=( a72449a  and  a72446a );
 a72451a <=( a72450a  and  a72443a );
 a72455a <=( (not A266)  and  (not A234) );
 a72456a <=( (not A233)  and  a72455a );
 a72459a <=( (not A269)  and  (not A268) );
 a72462a <=( (not A299)  and  (not A298) );
 a72463a <=( a72462a  and  a72459a );
 a72464a <=( a72463a  and  a72456a );
 a72468a <=( (not A168)  and  A169 );
 a72469a <=( A170  and  a72468a );
 a72472a <=( (not A200)  and  A199 );
 a72475a <=( A202  and  A201 );
 a72476a <=( a72475a  and  a72472a );
 a72477a <=( a72476a  and  a72469a );
 a72481a <=( (not A266)  and  (not A234) );
 a72482a <=( (not A233)  and  a72481a );
 a72485a <=( A298  and  (not A267) );
 a72488a <=( (not A302)  and  (not A301) );
 a72489a <=( a72488a  and  a72485a );
 a72490a <=( a72489a  and  a72482a );
 a72494a <=( (not A168)  and  A169 );
 a72495a <=( A170  and  a72494a );
 a72498a <=( (not A200)  and  A199 );
 a72501a <=( A202  and  A201 );
 a72502a <=( a72501a  and  a72498a );
 a72503a <=( a72502a  and  a72495a );
 a72507a <=( (not A265)  and  (not A234) );
 a72508a <=( (not A233)  and  a72507a );
 a72511a <=( A298  and  (not A266) );
 a72514a <=( (not A302)  and  (not A301) );
 a72515a <=( a72514a  and  a72511a );
 a72516a <=( a72515a  and  a72508a );
 a72520a <=( (not A168)  and  A169 );
 a72521a <=( A170  and  a72520a );
 a72524a <=( (not A200)  and  A199 );
 a72527a <=( A202  and  A201 );
 a72528a <=( a72527a  and  a72524a );
 a72529a <=( a72528a  and  a72521a );
 a72533a <=( A265  and  (not A233) );
 a72534a <=( (not A232)  and  a72533a );
 a72537a <=( A298  and  A266 );
 a72540a <=( (not A302)  and  (not A301) );
 a72541a <=( a72540a  and  a72537a );
 a72542a <=( a72541a  and  a72534a );
 a72546a <=( (not A168)  and  A169 );
 a72547a <=( A170  and  a72546a );
 a72550a <=( (not A200)  and  A199 );
 a72553a <=( A202  and  A201 );
 a72554a <=( a72553a  and  a72550a );
 a72555a <=( a72554a  and  a72547a );
 a72559a <=( (not A266)  and  (not A233) );
 a72560a <=( (not A232)  and  a72559a );
 a72563a <=( (not A269)  and  (not A268) );
 a72566a <=( (not A300)  and  A298 );
 a72567a <=( a72566a  and  a72563a );
 a72568a <=( a72567a  and  a72560a );
 a72572a <=( (not A168)  and  A169 );
 a72573a <=( A170  and  a72572a );
 a72576a <=( (not A200)  and  A199 );
 a72579a <=( A202  and  A201 );
 a72580a <=( a72579a  and  a72576a );
 a72581a <=( a72580a  and  a72573a );
 a72585a <=( (not A266)  and  (not A233) );
 a72586a <=( (not A232)  and  a72585a );
 a72589a <=( (not A269)  and  (not A268) );
 a72592a <=( A299  and  A298 );
 a72593a <=( a72592a  and  a72589a );
 a72594a <=( a72593a  and  a72586a );
 a72598a <=( (not A168)  and  A169 );
 a72599a <=( A170  and  a72598a );
 a72602a <=( (not A200)  and  A199 );
 a72605a <=( A202  and  A201 );
 a72606a <=( a72605a  and  a72602a );
 a72607a <=( a72606a  and  a72599a );
 a72611a <=( (not A266)  and  (not A233) );
 a72612a <=( (not A232)  and  a72611a );
 a72615a <=( (not A269)  and  (not A268) );
 a72618a <=( (not A299)  and  (not A298) );
 a72619a <=( a72618a  and  a72615a );
 a72620a <=( a72619a  and  a72612a );
 a72624a <=( (not A168)  and  A169 );
 a72625a <=( A170  and  a72624a );
 a72628a <=( (not A200)  and  A199 );
 a72631a <=( A202  and  A201 );
 a72632a <=( a72631a  and  a72628a );
 a72633a <=( a72632a  and  a72625a );
 a72637a <=( (not A266)  and  (not A233) );
 a72638a <=( (not A232)  and  a72637a );
 a72641a <=( A298  and  (not A267) );
 a72644a <=( (not A302)  and  (not A301) );
 a72645a <=( a72644a  and  a72641a );
 a72646a <=( a72645a  and  a72638a );
 a72650a <=( (not A168)  and  A169 );
 a72651a <=( A170  and  a72650a );
 a72654a <=( (not A200)  and  A199 );
 a72657a <=( A202  and  A201 );
 a72658a <=( a72657a  and  a72654a );
 a72659a <=( a72658a  and  a72651a );
 a72663a <=( (not A265)  and  (not A233) );
 a72664a <=( (not A232)  and  a72663a );
 a72667a <=( A298  and  (not A266) );
 a72670a <=( (not A302)  and  (not A301) );
 a72671a <=( a72670a  and  a72667a );
 a72672a <=( a72671a  and  a72664a );
 a72676a <=( (not A168)  and  A169 );
 a72677a <=( A170  and  a72676a );
 a72680a <=( (not A200)  and  A199 );
 a72683a <=( A203  and  A201 );
 a72684a <=( a72683a  and  a72680a );
 a72685a <=( a72684a  and  a72677a );
 a72689a <=( A265  and  A233 );
 a72690a <=( A232  and  a72689a );
 a72693a <=( (not A269)  and  (not A268) );
 a72696a <=( (not A300)  and  (not A299) );
 a72697a <=( a72696a  and  a72693a );
 a72698a <=( a72697a  and  a72690a );
 a72702a <=( (not A168)  and  A169 );
 a72703a <=( A170  and  a72702a );
 a72706a <=( (not A200)  and  A199 );
 a72709a <=( A203  and  A201 );
 a72710a <=( a72709a  and  a72706a );
 a72711a <=( a72710a  and  a72703a );
 a72715a <=( A265  and  A233 );
 a72716a <=( A232  and  a72715a );
 a72719a <=( (not A269)  and  (not A268) );
 a72722a <=( A299  and  A298 );
 a72723a <=( a72722a  and  a72719a );
 a72724a <=( a72723a  and  a72716a );
 a72728a <=( (not A168)  and  A169 );
 a72729a <=( A170  and  a72728a );
 a72732a <=( (not A200)  and  A199 );
 a72735a <=( A203  and  A201 );
 a72736a <=( a72735a  and  a72732a );
 a72737a <=( a72736a  and  a72729a );
 a72741a <=( A265  and  A233 );
 a72742a <=( A232  and  a72741a );
 a72745a <=( (not A269)  and  (not A268) );
 a72748a <=( (not A299)  and  (not A298) );
 a72749a <=( a72748a  and  a72745a );
 a72750a <=( a72749a  and  a72742a );
 a72754a <=( (not A168)  and  A169 );
 a72755a <=( A170  and  a72754a );
 a72758a <=( (not A200)  and  A199 );
 a72761a <=( A203  and  A201 );
 a72762a <=( a72761a  and  a72758a );
 a72763a <=( a72762a  and  a72755a );
 a72767a <=( A265  and  A233 );
 a72768a <=( A232  and  a72767a );
 a72771a <=( (not A299)  and  (not A267) );
 a72774a <=( (not A302)  and  (not A301) );
 a72775a <=( a72774a  and  a72771a );
 a72776a <=( a72775a  and  a72768a );
 a72780a <=( (not A168)  and  A169 );
 a72781a <=( A170  and  a72780a );
 a72784a <=( (not A200)  and  A199 );
 a72787a <=( A203  and  A201 );
 a72788a <=( a72787a  and  a72784a );
 a72789a <=( a72788a  and  a72781a );
 a72793a <=( A265  and  A233 );
 a72794a <=( A232  and  a72793a );
 a72797a <=( (not A299)  and  A266 );
 a72800a <=( (not A302)  and  (not A301) );
 a72801a <=( a72800a  and  a72797a );
 a72802a <=( a72801a  and  a72794a );
 a72806a <=( (not A168)  and  A169 );
 a72807a <=( A170  and  a72806a );
 a72810a <=( (not A200)  and  A199 );
 a72813a <=( A203  and  A201 );
 a72814a <=( a72813a  and  a72810a );
 a72815a <=( a72814a  and  a72807a );
 a72819a <=( (not A265)  and  A233 );
 a72820a <=( A232  and  a72819a );
 a72823a <=( (not A299)  and  (not A266) );
 a72826a <=( (not A302)  and  (not A301) );
 a72827a <=( a72826a  and  a72823a );
 a72828a <=( a72827a  and  a72820a );
 a72832a <=( (not A168)  and  A169 );
 a72833a <=( A170  and  a72832a );
 a72836a <=( (not A200)  and  A199 );
 a72839a <=( A203  and  A201 );
 a72840a <=( a72839a  and  a72836a );
 a72841a <=( a72840a  and  a72833a );
 a72845a <=( (not A236)  and  (not A235) );
 a72846a <=( (not A233)  and  a72845a );
 a72849a <=( A266  and  A265 );
 a72852a <=( (not A300)  and  A298 );
 a72853a <=( a72852a  and  a72849a );
 a72854a <=( a72853a  and  a72846a );
 a72858a <=( (not A168)  and  A169 );
 a72859a <=( A170  and  a72858a );
 a72862a <=( (not A200)  and  A199 );
 a72865a <=( A203  and  A201 );
 a72866a <=( a72865a  and  a72862a );
 a72867a <=( a72866a  and  a72859a );
 a72871a <=( (not A236)  and  (not A235) );
 a72872a <=( (not A233)  and  a72871a );
 a72875a <=( A266  and  A265 );
 a72878a <=( A299  and  A298 );
 a72879a <=( a72878a  and  a72875a );
 a72880a <=( a72879a  and  a72872a );
 a72884a <=( (not A168)  and  A169 );
 a72885a <=( A170  and  a72884a );
 a72888a <=( (not A200)  and  A199 );
 a72891a <=( A203  and  A201 );
 a72892a <=( a72891a  and  a72888a );
 a72893a <=( a72892a  and  a72885a );
 a72897a <=( (not A236)  and  (not A235) );
 a72898a <=( (not A233)  and  a72897a );
 a72901a <=( A266  and  A265 );
 a72904a <=( (not A299)  and  (not A298) );
 a72905a <=( a72904a  and  a72901a );
 a72906a <=( a72905a  and  a72898a );
 a72910a <=( (not A168)  and  A169 );
 a72911a <=( A170  and  a72910a );
 a72914a <=( (not A200)  and  A199 );
 a72917a <=( A203  and  A201 );
 a72918a <=( a72917a  and  a72914a );
 a72919a <=( a72918a  and  a72911a );
 a72923a <=( (not A236)  and  (not A235) );
 a72924a <=( (not A233)  and  a72923a );
 a72927a <=( (not A267)  and  (not A266) );
 a72930a <=( (not A300)  and  A298 );
 a72931a <=( a72930a  and  a72927a );
 a72932a <=( a72931a  and  a72924a );
 a72936a <=( (not A168)  and  A169 );
 a72937a <=( A170  and  a72936a );
 a72940a <=( (not A200)  and  A199 );
 a72943a <=( A203  and  A201 );
 a72944a <=( a72943a  and  a72940a );
 a72945a <=( a72944a  and  a72937a );
 a72949a <=( (not A236)  and  (not A235) );
 a72950a <=( (not A233)  and  a72949a );
 a72953a <=( (not A267)  and  (not A266) );
 a72956a <=( A299  and  A298 );
 a72957a <=( a72956a  and  a72953a );
 a72958a <=( a72957a  and  a72950a );
 a72962a <=( (not A168)  and  A169 );
 a72963a <=( A170  and  a72962a );
 a72966a <=( (not A200)  and  A199 );
 a72969a <=( A203  and  A201 );
 a72970a <=( a72969a  and  a72966a );
 a72971a <=( a72970a  and  a72963a );
 a72975a <=( (not A236)  and  (not A235) );
 a72976a <=( (not A233)  and  a72975a );
 a72979a <=( (not A267)  and  (not A266) );
 a72982a <=( (not A299)  and  (not A298) );
 a72983a <=( a72982a  and  a72979a );
 a72984a <=( a72983a  and  a72976a );
 a72988a <=( (not A168)  and  A169 );
 a72989a <=( A170  and  a72988a );
 a72992a <=( (not A200)  and  A199 );
 a72995a <=( A203  and  A201 );
 a72996a <=( a72995a  and  a72992a );
 a72997a <=( a72996a  and  a72989a );
 a73001a <=( (not A236)  and  (not A235) );
 a73002a <=( (not A233)  and  a73001a );
 a73005a <=( (not A266)  and  (not A265) );
 a73008a <=( (not A300)  and  A298 );
 a73009a <=( a73008a  and  a73005a );
 a73010a <=( a73009a  and  a73002a );
 a73014a <=( (not A168)  and  A169 );
 a73015a <=( A170  and  a73014a );
 a73018a <=( (not A200)  and  A199 );
 a73021a <=( A203  and  A201 );
 a73022a <=( a73021a  and  a73018a );
 a73023a <=( a73022a  and  a73015a );
 a73027a <=( (not A236)  and  (not A235) );
 a73028a <=( (not A233)  and  a73027a );
 a73031a <=( (not A266)  and  (not A265) );
 a73034a <=( A299  and  A298 );
 a73035a <=( a73034a  and  a73031a );
 a73036a <=( a73035a  and  a73028a );
 a73040a <=( (not A168)  and  A169 );
 a73041a <=( A170  and  a73040a );
 a73044a <=( (not A200)  and  A199 );
 a73047a <=( A203  and  A201 );
 a73048a <=( a73047a  and  a73044a );
 a73049a <=( a73048a  and  a73041a );
 a73053a <=( (not A236)  and  (not A235) );
 a73054a <=( (not A233)  and  a73053a );
 a73057a <=( (not A266)  and  (not A265) );
 a73060a <=( (not A299)  and  (not A298) );
 a73061a <=( a73060a  and  a73057a );
 a73062a <=( a73061a  and  a73054a );
 a73066a <=( (not A168)  and  A169 );
 a73067a <=( A170  and  a73066a );
 a73070a <=( (not A200)  and  A199 );
 a73073a <=( A203  and  A201 );
 a73074a <=( a73073a  and  a73070a );
 a73075a <=( a73074a  and  a73067a );
 a73079a <=( A265  and  (not A234) );
 a73080a <=( (not A233)  and  a73079a );
 a73083a <=( A298  and  A266 );
 a73086a <=( (not A302)  and  (not A301) );
 a73087a <=( a73086a  and  a73083a );
 a73088a <=( a73087a  and  a73080a );
 a73092a <=( (not A168)  and  A169 );
 a73093a <=( A170  and  a73092a );
 a73096a <=( (not A200)  and  A199 );
 a73099a <=( A203  and  A201 );
 a73100a <=( a73099a  and  a73096a );
 a73101a <=( a73100a  and  a73093a );
 a73105a <=( (not A266)  and  (not A234) );
 a73106a <=( (not A233)  and  a73105a );
 a73109a <=( (not A269)  and  (not A268) );
 a73112a <=( (not A300)  and  A298 );
 a73113a <=( a73112a  and  a73109a );
 a73114a <=( a73113a  and  a73106a );
 a73118a <=( (not A168)  and  A169 );
 a73119a <=( A170  and  a73118a );
 a73122a <=( (not A200)  and  A199 );
 a73125a <=( A203  and  A201 );
 a73126a <=( a73125a  and  a73122a );
 a73127a <=( a73126a  and  a73119a );
 a73131a <=( (not A266)  and  (not A234) );
 a73132a <=( (not A233)  and  a73131a );
 a73135a <=( (not A269)  and  (not A268) );
 a73138a <=( A299  and  A298 );
 a73139a <=( a73138a  and  a73135a );
 a73140a <=( a73139a  and  a73132a );
 a73144a <=( (not A168)  and  A169 );
 a73145a <=( A170  and  a73144a );
 a73148a <=( (not A200)  and  A199 );
 a73151a <=( A203  and  A201 );
 a73152a <=( a73151a  and  a73148a );
 a73153a <=( a73152a  and  a73145a );
 a73157a <=( (not A266)  and  (not A234) );
 a73158a <=( (not A233)  and  a73157a );
 a73161a <=( (not A269)  and  (not A268) );
 a73164a <=( (not A299)  and  (not A298) );
 a73165a <=( a73164a  and  a73161a );
 a73166a <=( a73165a  and  a73158a );
 a73170a <=( (not A168)  and  A169 );
 a73171a <=( A170  and  a73170a );
 a73174a <=( (not A200)  and  A199 );
 a73177a <=( A203  and  A201 );
 a73178a <=( a73177a  and  a73174a );
 a73179a <=( a73178a  and  a73171a );
 a73183a <=( (not A266)  and  (not A234) );
 a73184a <=( (not A233)  and  a73183a );
 a73187a <=( A298  and  (not A267) );
 a73190a <=( (not A302)  and  (not A301) );
 a73191a <=( a73190a  and  a73187a );
 a73192a <=( a73191a  and  a73184a );
 a73196a <=( (not A168)  and  A169 );
 a73197a <=( A170  and  a73196a );
 a73200a <=( (not A200)  and  A199 );
 a73203a <=( A203  and  A201 );
 a73204a <=( a73203a  and  a73200a );
 a73205a <=( a73204a  and  a73197a );
 a73209a <=( (not A265)  and  (not A234) );
 a73210a <=( (not A233)  and  a73209a );
 a73213a <=( A298  and  (not A266) );
 a73216a <=( (not A302)  and  (not A301) );
 a73217a <=( a73216a  and  a73213a );
 a73218a <=( a73217a  and  a73210a );
 a73222a <=( (not A168)  and  A169 );
 a73223a <=( A170  and  a73222a );
 a73226a <=( (not A200)  and  A199 );
 a73229a <=( A203  and  A201 );
 a73230a <=( a73229a  and  a73226a );
 a73231a <=( a73230a  and  a73223a );
 a73235a <=( A265  and  (not A233) );
 a73236a <=( (not A232)  and  a73235a );
 a73239a <=( A298  and  A266 );
 a73242a <=( (not A302)  and  (not A301) );
 a73243a <=( a73242a  and  a73239a );
 a73244a <=( a73243a  and  a73236a );
 a73248a <=( (not A168)  and  A169 );
 a73249a <=( A170  and  a73248a );
 a73252a <=( (not A200)  and  A199 );
 a73255a <=( A203  and  A201 );
 a73256a <=( a73255a  and  a73252a );
 a73257a <=( a73256a  and  a73249a );
 a73261a <=( (not A266)  and  (not A233) );
 a73262a <=( (not A232)  and  a73261a );
 a73265a <=( (not A269)  and  (not A268) );
 a73268a <=( (not A300)  and  A298 );
 a73269a <=( a73268a  and  a73265a );
 a73270a <=( a73269a  and  a73262a );
 a73274a <=( (not A168)  and  A169 );
 a73275a <=( A170  and  a73274a );
 a73278a <=( (not A200)  and  A199 );
 a73281a <=( A203  and  A201 );
 a73282a <=( a73281a  and  a73278a );
 a73283a <=( a73282a  and  a73275a );
 a73287a <=( (not A266)  and  (not A233) );
 a73288a <=( (not A232)  and  a73287a );
 a73291a <=( (not A269)  and  (not A268) );
 a73294a <=( A299  and  A298 );
 a73295a <=( a73294a  and  a73291a );
 a73296a <=( a73295a  and  a73288a );
 a73300a <=( (not A168)  and  A169 );
 a73301a <=( A170  and  a73300a );
 a73304a <=( (not A200)  and  A199 );
 a73307a <=( A203  and  A201 );
 a73308a <=( a73307a  and  a73304a );
 a73309a <=( a73308a  and  a73301a );
 a73313a <=( (not A266)  and  (not A233) );
 a73314a <=( (not A232)  and  a73313a );
 a73317a <=( (not A269)  and  (not A268) );
 a73320a <=( (not A299)  and  (not A298) );
 a73321a <=( a73320a  and  a73317a );
 a73322a <=( a73321a  and  a73314a );
 a73326a <=( (not A168)  and  A169 );
 a73327a <=( A170  and  a73326a );
 a73330a <=( (not A200)  and  A199 );
 a73333a <=( A203  and  A201 );
 a73334a <=( a73333a  and  a73330a );
 a73335a <=( a73334a  and  a73327a );
 a73339a <=( (not A266)  and  (not A233) );
 a73340a <=( (not A232)  and  a73339a );
 a73343a <=( A298  and  (not A267) );
 a73346a <=( (not A302)  and  (not A301) );
 a73347a <=( a73346a  and  a73343a );
 a73348a <=( a73347a  and  a73340a );
 a73352a <=( (not A168)  and  A169 );
 a73353a <=( A170  and  a73352a );
 a73356a <=( (not A200)  and  A199 );
 a73359a <=( A203  and  A201 );
 a73360a <=( a73359a  and  a73356a );
 a73361a <=( a73360a  and  a73353a );
 a73365a <=( (not A265)  and  (not A233) );
 a73366a <=( (not A232)  and  a73365a );
 a73369a <=( A298  and  (not A266) );
 a73372a <=( (not A302)  and  (not A301) );
 a73373a <=( a73372a  and  a73369a );
 a73374a <=( a73373a  and  a73366a );
 a73378a <=( (not A168)  and  A169 );
 a73379a <=( A170  and  a73378a );
 a73382a <=( A199  and  A166 );
 a73385a <=( A201  and  (not A200) );
 a73386a <=( a73385a  and  a73382a );
 a73387a <=( a73386a  and  a73379a );
 a73391a <=( A233  and  (not A232) );
 a73392a <=( A202  and  a73391a );
 a73395a <=( (not A299)  and  A298 );
 a73398a <=( A301  and  A300 );
 a73399a <=( a73398a  and  a73395a );
 a73400a <=( a73399a  and  a73392a );
 a73404a <=( (not A168)  and  A169 );
 a73405a <=( A170  and  a73404a );
 a73408a <=( A199  and  A166 );
 a73411a <=( A201  and  (not A200) );
 a73412a <=( a73411a  and  a73408a );
 a73413a <=( a73412a  and  a73405a );
 a73417a <=( A233  and  (not A232) );
 a73418a <=( A202  and  a73417a );
 a73421a <=( (not A299)  and  A298 );
 a73424a <=( A302  and  A300 );
 a73425a <=( a73424a  and  a73421a );
 a73426a <=( a73425a  and  a73418a );
 a73430a <=( (not A168)  and  A169 );
 a73431a <=( A170  and  a73430a );
 a73434a <=( A199  and  A166 );
 a73437a <=( A201  and  (not A200) );
 a73438a <=( a73437a  and  a73434a );
 a73439a <=( a73438a  and  a73431a );
 a73443a <=( A233  and  (not A232) );
 a73444a <=( A202  and  a73443a );
 a73447a <=( (not A266)  and  A265 );
 a73450a <=( A268  and  A267 );
 a73451a <=( a73450a  and  a73447a );
 a73452a <=( a73451a  and  a73444a );
 a73456a <=( (not A168)  and  A169 );
 a73457a <=( A170  and  a73456a );
 a73460a <=( A199  and  A166 );
 a73463a <=( A201  and  (not A200) );
 a73464a <=( a73463a  and  a73460a );
 a73465a <=( a73464a  and  a73457a );
 a73469a <=( A233  and  (not A232) );
 a73470a <=( A202  and  a73469a );
 a73473a <=( (not A266)  and  A265 );
 a73476a <=( A269  and  A267 );
 a73477a <=( a73476a  and  a73473a );
 a73478a <=( a73477a  and  a73470a );
 a73482a <=( (not A168)  and  A169 );
 a73483a <=( A170  and  a73482a );
 a73486a <=( A199  and  A166 );
 a73489a <=( A201  and  (not A200) );
 a73490a <=( a73489a  and  a73486a );
 a73491a <=( a73490a  and  a73483a );
 a73495a <=( A233  and  (not A232) );
 a73496a <=( A203  and  a73495a );
 a73499a <=( (not A299)  and  A298 );
 a73502a <=( A301  and  A300 );
 a73503a <=( a73502a  and  a73499a );
 a73504a <=( a73503a  and  a73496a );
 a73508a <=( (not A168)  and  A169 );
 a73509a <=( A170  and  a73508a );
 a73512a <=( A199  and  A166 );
 a73515a <=( A201  and  (not A200) );
 a73516a <=( a73515a  and  a73512a );
 a73517a <=( a73516a  and  a73509a );
 a73521a <=( A233  and  (not A232) );
 a73522a <=( A203  and  a73521a );
 a73525a <=( (not A299)  and  A298 );
 a73528a <=( A302  and  A300 );
 a73529a <=( a73528a  and  a73525a );
 a73530a <=( a73529a  and  a73522a );
 a73534a <=( (not A168)  and  A169 );
 a73535a <=( A170  and  a73534a );
 a73538a <=( A199  and  A166 );
 a73541a <=( A201  and  (not A200) );
 a73542a <=( a73541a  and  a73538a );
 a73543a <=( a73542a  and  a73535a );
 a73547a <=( A233  and  (not A232) );
 a73548a <=( A203  and  a73547a );
 a73551a <=( (not A266)  and  A265 );
 a73554a <=( A268  and  A267 );
 a73555a <=( a73554a  and  a73551a );
 a73556a <=( a73555a  and  a73548a );
 a73560a <=( (not A168)  and  A169 );
 a73561a <=( A170  and  a73560a );
 a73564a <=( A199  and  A166 );
 a73567a <=( A201  and  (not A200) );
 a73568a <=( a73567a  and  a73564a );
 a73569a <=( a73568a  and  a73561a );
 a73573a <=( A233  and  (not A232) );
 a73574a <=( A203  and  a73573a );
 a73577a <=( (not A266)  and  A265 );
 a73580a <=( A269  and  A267 );
 a73581a <=( a73580a  and  a73577a );
 a73582a <=( a73581a  and  a73574a );
 a73586a <=( A167  and  A169 );
 a73587a <=( (not A170)  and  a73586a );
 a73590a <=( A199  and  A166 );
 a73593a <=( A232  and  A200 );
 a73594a <=( a73593a  and  a73590a );
 a73595a <=( a73594a  and  a73587a );
 a73599a <=( (not A268)  and  A265 );
 a73600a <=( A233  and  a73599a );
 a73603a <=( (not A299)  and  (not A269) );
 a73606a <=( (not A302)  and  (not A301) );
 a73607a <=( a73606a  and  a73603a );
 a73608a <=( a73607a  and  a73600a );
 a73612a <=( A167  and  A169 );
 a73613a <=( (not A170)  and  a73612a );
 a73616a <=( A199  and  A166 );
 a73619a <=( (not A233)  and  A200 );
 a73620a <=( a73619a  and  a73616a );
 a73621a <=( a73620a  and  a73613a );
 a73625a <=( A265  and  (not A236) );
 a73626a <=( (not A235)  and  a73625a );
 a73629a <=( A298  and  A266 );
 a73632a <=( (not A302)  and  (not A301) );
 a73633a <=( a73632a  and  a73629a );
 a73634a <=( a73633a  and  a73626a );
 a73638a <=( A167  and  A169 );
 a73639a <=( (not A170)  and  a73638a );
 a73642a <=( A199  and  A166 );
 a73645a <=( (not A233)  and  A200 );
 a73646a <=( a73645a  and  a73642a );
 a73647a <=( a73646a  and  a73639a );
 a73651a <=( (not A266)  and  (not A236) );
 a73652a <=( (not A235)  and  a73651a );
 a73655a <=( (not A269)  and  (not A268) );
 a73658a <=( (not A300)  and  A298 );
 a73659a <=( a73658a  and  a73655a );
 a73660a <=( a73659a  and  a73652a );
 a73664a <=( A167  and  A169 );
 a73665a <=( (not A170)  and  a73664a );
 a73668a <=( A199  and  A166 );
 a73671a <=( (not A233)  and  A200 );
 a73672a <=( a73671a  and  a73668a );
 a73673a <=( a73672a  and  a73665a );
 a73677a <=( (not A266)  and  (not A236) );
 a73678a <=( (not A235)  and  a73677a );
 a73681a <=( (not A269)  and  (not A268) );
 a73684a <=( A299  and  A298 );
 a73685a <=( a73684a  and  a73681a );
 a73686a <=( a73685a  and  a73678a );
 a73690a <=( A167  and  A169 );
 a73691a <=( (not A170)  and  a73690a );
 a73694a <=( A199  and  A166 );
 a73697a <=( (not A233)  and  A200 );
 a73698a <=( a73697a  and  a73694a );
 a73699a <=( a73698a  and  a73691a );
 a73703a <=( (not A266)  and  (not A236) );
 a73704a <=( (not A235)  and  a73703a );
 a73707a <=( (not A269)  and  (not A268) );
 a73710a <=( (not A299)  and  (not A298) );
 a73711a <=( a73710a  and  a73707a );
 a73712a <=( a73711a  and  a73704a );
 a73716a <=( A167  and  A169 );
 a73717a <=( (not A170)  and  a73716a );
 a73720a <=( A199  and  A166 );
 a73723a <=( (not A233)  and  A200 );
 a73724a <=( a73723a  and  a73720a );
 a73725a <=( a73724a  and  a73717a );
 a73729a <=( (not A266)  and  (not A236) );
 a73730a <=( (not A235)  and  a73729a );
 a73733a <=( A298  and  (not A267) );
 a73736a <=( (not A302)  and  (not A301) );
 a73737a <=( a73736a  and  a73733a );
 a73738a <=( a73737a  and  a73730a );
 a73742a <=( A167  and  A169 );
 a73743a <=( (not A170)  and  a73742a );
 a73746a <=( A199  and  A166 );
 a73749a <=( (not A233)  and  A200 );
 a73750a <=( a73749a  and  a73746a );
 a73751a <=( a73750a  and  a73743a );
 a73755a <=( (not A265)  and  (not A236) );
 a73756a <=( (not A235)  and  a73755a );
 a73759a <=( A298  and  (not A266) );
 a73762a <=( (not A302)  and  (not A301) );
 a73763a <=( a73762a  and  a73759a );
 a73764a <=( a73763a  and  a73756a );
 a73768a <=( A167  and  A169 );
 a73769a <=( (not A170)  and  a73768a );
 a73772a <=( A199  and  A166 );
 a73775a <=( (not A233)  and  A200 );
 a73776a <=( a73775a  and  a73772a );
 a73777a <=( a73776a  and  a73769a );
 a73781a <=( (not A268)  and  (not A266) );
 a73782a <=( (not A234)  and  a73781a );
 a73785a <=( A298  and  (not A269) );
 a73788a <=( (not A302)  and  (not A301) );
 a73789a <=( a73788a  and  a73785a );
 a73790a <=( a73789a  and  a73782a );
 a73794a <=( A167  and  A169 );
 a73795a <=( (not A170)  and  a73794a );
 a73798a <=( A199  and  A166 );
 a73801a <=( A232  and  A200 );
 a73802a <=( a73801a  and  a73798a );
 a73803a <=( a73802a  and  a73795a );
 a73807a <=( A235  and  A234 );
 a73808a <=( (not A233)  and  a73807a );
 a73811a <=( (not A299)  and  A298 );
 a73814a <=( A301  and  A300 );
 a73815a <=( a73814a  and  a73811a );
 a73816a <=( a73815a  and  a73808a );
 a73820a <=( A167  and  A169 );
 a73821a <=( (not A170)  and  a73820a );
 a73824a <=( A199  and  A166 );
 a73827a <=( A232  and  A200 );
 a73828a <=( a73827a  and  a73824a );
 a73829a <=( a73828a  and  a73821a );
 a73833a <=( A235  and  A234 );
 a73834a <=( (not A233)  and  a73833a );
 a73837a <=( (not A299)  and  A298 );
 a73840a <=( A302  and  A300 );
 a73841a <=( a73840a  and  a73837a );
 a73842a <=( a73841a  and  a73834a );
 a73846a <=( A167  and  A169 );
 a73847a <=( (not A170)  and  a73846a );
 a73850a <=( A199  and  A166 );
 a73853a <=( A232  and  A200 );
 a73854a <=( a73853a  and  a73850a );
 a73855a <=( a73854a  and  a73847a );
 a73859a <=( A235  and  A234 );
 a73860a <=( (not A233)  and  a73859a );
 a73863a <=( (not A266)  and  A265 );
 a73866a <=( A268  and  A267 );
 a73867a <=( a73866a  and  a73863a );
 a73868a <=( a73867a  and  a73860a );
 a73872a <=( A167  and  A169 );
 a73873a <=( (not A170)  and  a73872a );
 a73876a <=( A199  and  A166 );
 a73879a <=( A232  and  A200 );
 a73880a <=( a73879a  and  a73876a );
 a73881a <=( a73880a  and  a73873a );
 a73885a <=( A235  and  A234 );
 a73886a <=( (not A233)  and  a73885a );
 a73889a <=( (not A266)  and  A265 );
 a73892a <=( A269  and  A267 );
 a73893a <=( a73892a  and  a73889a );
 a73894a <=( a73893a  and  a73886a );
 a73898a <=( A167  and  A169 );
 a73899a <=( (not A170)  and  a73898a );
 a73902a <=( A199  and  A166 );
 a73905a <=( A232  and  A200 );
 a73906a <=( a73905a  and  a73902a );
 a73907a <=( a73906a  and  a73899a );
 a73911a <=( A236  and  A234 );
 a73912a <=( (not A233)  and  a73911a );
 a73915a <=( (not A299)  and  A298 );
 a73918a <=( A301  and  A300 );
 a73919a <=( a73918a  and  a73915a );
 a73920a <=( a73919a  and  a73912a );
 a73924a <=( A167  and  A169 );
 a73925a <=( (not A170)  and  a73924a );
 a73928a <=( A199  and  A166 );
 a73931a <=( A232  and  A200 );
 a73932a <=( a73931a  and  a73928a );
 a73933a <=( a73932a  and  a73925a );
 a73937a <=( A236  and  A234 );
 a73938a <=( (not A233)  and  a73937a );
 a73941a <=( (not A299)  and  A298 );
 a73944a <=( A302  and  A300 );
 a73945a <=( a73944a  and  a73941a );
 a73946a <=( a73945a  and  a73938a );
 a73950a <=( A167  and  A169 );
 a73951a <=( (not A170)  and  a73950a );
 a73954a <=( A199  and  A166 );
 a73957a <=( A232  and  A200 );
 a73958a <=( a73957a  and  a73954a );
 a73959a <=( a73958a  and  a73951a );
 a73963a <=( A236  and  A234 );
 a73964a <=( (not A233)  and  a73963a );
 a73967a <=( (not A266)  and  A265 );
 a73970a <=( A268  and  A267 );
 a73971a <=( a73970a  and  a73967a );
 a73972a <=( a73971a  and  a73964a );
 a73976a <=( A167  and  A169 );
 a73977a <=( (not A170)  and  a73976a );
 a73980a <=( A199  and  A166 );
 a73983a <=( A232  and  A200 );
 a73984a <=( a73983a  and  a73980a );
 a73985a <=( a73984a  and  a73977a );
 a73989a <=( A236  and  A234 );
 a73990a <=( (not A233)  and  a73989a );
 a73993a <=( (not A266)  and  A265 );
 a73996a <=( A269  and  A267 );
 a73997a <=( a73996a  and  a73993a );
 a73998a <=( a73997a  and  a73990a );
 a74002a <=( A167  and  A169 );
 a74003a <=( (not A170)  and  a74002a );
 a74006a <=( A199  and  A166 );
 a74009a <=( (not A232)  and  A200 );
 a74010a <=( a74009a  and  a74006a );
 a74011a <=( a74010a  and  a74003a );
 a74015a <=( (not A268)  and  (not A266) );
 a74016a <=( (not A233)  and  a74015a );
 a74019a <=( A298  and  (not A269) );
 a74022a <=( (not A302)  and  (not A301) );
 a74023a <=( a74022a  and  a74019a );
 a74024a <=( a74023a  and  a74016a );
 a74028a <=( A167  and  A169 );
 a74029a <=( (not A170)  and  a74028a );
 a74032a <=( (not A200)  and  A166 );
 a74035a <=( (not A203)  and  (not A202) );
 a74036a <=( a74035a  and  a74032a );
 a74037a <=( a74036a  and  a74029a );
 a74041a <=( A265  and  A233 );
 a74042a <=( A232  and  a74041a );
 a74045a <=( (not A269)  and  (not A268) );
 a74048a <=( (not A300)  and  (not A299) );
 a74049a <=( a74048a  and  a74045a );
 a74050a <=( a74049a  and  a74042a );
 a74054a <=( A167  and  A169 );
 a74055a <=( (not A170)  and  a74054a );
 a74058a <=( (not A200)  and  A166 );
 a74061a <=( (not A203)  and  (not A202) );
 a74062a <=( a74061a  and  a74058a );
 a74063a <=( a74062a  and  a74055a );
 a74067a <=( A265  and  A233 );
 a74068a <=( A232  and  a74067a );
 a74071a <=( (not A269)  and  (not A268) );
 a74074a <=( A299  and  A298 );
 a74075a <=( a74074a  and  a74071a );
 a74076a <=( a74075a  and  a74068a );
 a74080a <=( A167  and  A169 );
 a74081a <=( (not A170)  and  a74080a );
 a74084a <=( (not A200)  and  A166 );
 a74087a <=( (not A203)  and  (not A202) );
 a74088a <=( a74087a  and  a74084a );
 a74089a <=( a74088a  and  a74081a );
 a74093a <=( A265  and  A233 );
 a74094a <=( A232  and  a74093a );
 a74097a <=( (not A269)  and  (not A268) );
 a74100a <=( (not A299)  and  (not A298) );
 a74101a <=( a74100a  and  a74097a );
 a74102a <=( a74101a  and  a74094a );
 a74106a <=( A167  and  A169 );
 a74107a <=( (not A170)  and  a74106a );
 a74110a <=( (not A200)  and  A166 );
 a74113a <=( (not A203)  and  (not A202) );
 a74114a <=( a74113a  and  a74110a );
 a74115a <=( a74114a  and  a74107a );
 a74119a <=( A265  and  A233 );
 a74120a <=( A232  and  a74119a );
 a74123a <=( (not A299)  and  (not A267) );
 a74126a <=( (not A302)  and  (not A301) );
 a74127a <=( a74126a  and  a74123a );
 a74128a <=( a74127a  and  a74120a );
 a74132a <=( A167  and  A169 );
 a74133a <=( (not A170)  and  a74132a );
 a74136a <=( (not A200)  and  A166 );
 a74139a <=( (not A203)  and  (not A202) );
 a74140a <=( a74139a  and  a74136a );
 a74141a <=( a74140a  and  a74133a );
 a74145a <=( A265  and  A233 );
 a74146a <=( A232  and  a74145a );
 a74149a <=( (not A299)  and  A266 );
 a74152a <=( (not A302)  and  (not A301) );
 a74153a <=( a74152a  and  a74149a );
 a74154a <=( a74153a  and  a74146a );
 a74158a <=( A167  and  A169 );
 a74159a <=( (not A170)  and  a74158a );
 a74162a <=( (not A200)  and  A166 );
 a74165a <=( (not A203)  and  (not A202) );
 a74166a <=( a74165a  and  a74162a );
 a74167a <=( a74166a  and  a74159a );
 a74171a <=( (not A265)  and  A233 );
 a74172a <=( A232  and  a74171a );
 a74175a <=( (not A299)  and  (not A266) );
 a74178a <=( (not A302)  and  (not A301) );
 a74179a <=( a74178a  and  a74175a );
 a74180a <=( a74179a  and  a74172a );
 a74184a <=( A167  and  A169 );
 a74185a <=( (not A170)  and  a74184a );
 a74188a <=( (not A200)  and  A166 );
 a74191a <=( (not A203)  and  (not A202) );
 a74192a <=( a74191a  and  a74188a );
 a74193a <=( a74192a  and  a74185a );
 a74197a <=( (not A236)  and  (not A235) );
 a74198a <=( (not A233)  and  a74197a );
 a74201a <=( A266  and  A265 );
 a74204a <=( (not A300)  and  A298 );
 a74205a <=( a74204a  and  a74201a );
 a74206a <=( a74205a  and  a74198a );
 a74210a <=( A167  and  A169 );
 a74211a <=( (not A170)  and  a74210a );
 a74214a <=( (not A200)  and  A166 );
 a74217a <=( (not A203)  and  (not A202) );
 a74218a <=( a74217a  and  a74214a );
 a74219a <=( a74218a  and  a74211a );
 a74223a <=( (not A236)  and  (not A235) );
 a74224a <=( (not A233)  and  a74223a );
 a74227a <=( A266  and  A265 );
 a74230a <=( A299  and  A298 );
 a74231a <=( a74230a  and  a74227a );
 a74232a <=( a74231a  and  a74224a );
 a74236a <=( A167  and  A169 );
 a74237a <=( (not A170)  and  a74236a );
 a74240a <=( (not A200)  and  A166 );
 a74243a <=( (not A203)  and  (not A202) );
 a74244a <=( a74243a  and  a74240a );
 a74245a <=( a74244a  and  a74237a );
 a74249a <=( (not A236)  and  (not A235) );
 a74250a <=( (not A233)  and  a74249a );
 a74253a <=( A266  and  A265 );
 a74256a <=( (not A299)  and  (not A298) );
 a74257a <=( a74256a  and  a74253a );
 a74258a <=( a74257a  and  a74250a );
 a74262a <=( A167  and  A169 );
 a74263a <=( (not A170)  and  a74262a );
 a74266a <=( (not A200)  and  A166 );
 a74269a <=( (not A203)  and  (not A202) );
 a74270a <=( a74269a  and  a74266a );
 a74271a <=( a74270a  and  a74263a );
 a74275a <=( (not A236)  and  (not A235) );
 a74276a <=( (not A233)  and  a74275a );
 a74279a <=( (not A267)  and  (not A266) );
 a74282a <=( (not A300)  and  A298 );
 a74283a <=( a74282a  and  a74279a );
 a74284a <=( a74283a  and  a74276a );
 a74288a <=( A167  and  A169 );
 a74289a <=( (not A170)  and  a74288a );
 a74292a <=( (not A200)  and  A166 );
 a74295a <=( (not A203)  and  (not A202) );
 a74296a <=( a74295a  and  a74292a );
 a74297a <=( a74296a  and  a74289a );
 a74301a <=( (not A236)  and  (not A235) );
 a74302a <=( (not A233)  and  a74301a );
 a74305a <=( (not A267)  and  (not A266) );
 a74308a <=( A299  and  A298 );
 a74309a <=( a74308a  and  a74305a );
 a74310a <=( a74309a  and  a74302a );
 a74314a <=( A167  and  A169 );
 a74315a <=( (not A170)  and  a74314a );
 a74318a <=( (not A200)  and  A166 );
 a74321a <=( (not A203)  and  (not A202) );
 a74322a <=( a74321a  and  a74318a );
 a74323a <=( a74322a  and  a74315a );
 a74327a <=( (not A236)  and  (not A235) );
 a74328a <=( (not A233)  and  a74327a );
 a74331a <=( (not A267)  and  (not A266) );
 a74334a <=( (not A299)  and  (not A298) );
 a74335a <=( a74334a  and  a74331a );
 a74336a <=( a74335a  and  a74328a );
 a74340a <=( A167  and  A169 );
 a74341a <=( (not A170)  and  a74340a );
 a74344a <=( (not A200)  and  A166 );
 a74347a <=( (not A203)  and  (not A202) );
 a74348a <=( a74347a  and  a74344a );
 a74349a <=( a74348a  and  a74341a );
 a74353a <=( (not A236)  and  (not A235) );
 a74354a <=( (not A233)  and  a74353a );
 a74357a <=( (not A266)  and  (not A265) );
 a74360a <=( (not A300)  and  A298 );
 a74361a <=( a74360a  and  a74357a );
 a74362a <=( a74361a  and  a74354a );
 a74366a <=( A167  and  A169 );
 a74367a <=( (not A170)  and  a74366a );
 a74370a <=( (not A200)  and  A166 );
 a74373a <=( (not A203)  and  (not A202) );
 a74374a <=( a74373a  and  a74370a );
 a74375a <=( a74374a  and  a74367a );
 a74379a <=( (not A236)  and  (not A235) );
 a74380a <=( (not A233)  and  a74379a );
 a74383a <=( (not A266)  and  (not A265) );
 a74386a <=( A299  and  A298 );
 a74387a <=( a74386a  and  a74383a );
 a74388a <=( a74387a  and  a74380a );
 a74392a <=( A167  and  A169 );
 a74393a <=( (not A170)  and  a74392a );
 a74396a <=( (not A200)  and  A166 );
 a74399a <=( (not A203)  and  (not A202) );
 a74400a <=( a74399a  and  a74396a );
 a74401a <=( a74400a  and  a74393a );
 a74405a <=( (not A236)  and  (not A235) );
 a74406a <=( (not A233)  and  a74405a );
 a74409a <=( (not A266)  and  (not A265) );
 a74412a <=( (not A299)  and  (not A298) );
 a74413a <=( a74412a  and  a74409a );
 a74414a <=( a74413a  and  a74406a );
 a74418a <=( A167  and  A169 );
 a74419a <=( (not A170)  and  a74418a );
 a74422a <=( (not A200)  and  A166 );
 a74425a <=( (not A203)  and  (not A202) );
 a74426a <=( a74425a  and  a74422a );
 a74427a <=( a74426a  and  a74419a );
 a74431a <=( A265  and  (not A234) );
 a74432a <=( (not A233)  and  a74431a );
 a74435a <=( A298  and  A266 );
 a74438a <=( (not A302)  and  (not A301) );
 a74439a <=( a74438a  and  a74435a );
 a74440a <=( a74439a  and  a74432a );
 a74444a <=( A167  and  A169 );
 a74445a <=( (not A170)  and  a74444a );
 a74448a <=( (not A200)  and  A166 );
 a74451a <=( (not A203)  and  (not A202) );
 a74452a <=( a74451a  and  a74448a );
 a74453a <=( a74452a  and  a74445a );
 a74457a <=( (not A266)  and  (not A234) );
 a74458a <=( (not A233)  and  a74457a );
 a74461a <=( (not A269)  and  (not A268) );
 a74464a <=( (not A300)  and  A298 );
 a74465a <=( a74464a  and  a74461a );
 a74466a <=( a74465a  and  a74458a );
 a74470a <=( A167  and  A169 );
 a74471a <=( (not A170)  and  a74470a );
 a74474a <=( (not A200)  and  A166 );
 a74477a <=( (not A203)  and  (not A202) );
 a74478a <=( a74477a  and  a74474a );
 a74479a <=( a74478a  and  a74471a );
 a74483a <=( (not A266)  and  (not A234) );
 a74484a <=( (not A233)  and  a74483a );
 a74487a <=( (not A269)  and  (not A268) );
 a74490a <=( A299  and  A298 );
 a74491a <=( a74490a  and  a74487a );
 a74492a <=( a74491a  and  a74484a );
 a74496a <=( A167  and  A169 );
 a74497a <=( (not A170)  and  a74496a );
 a74500a <=( (not A200)  and  A166 );
 a74503a <=( (not A203)  and  (not A202) );
 a74504a <=( a74503a  and  a74500a );
 a74505a <=( a74504a  and  a74497a );
 a74509a <=( (not A266)  and  (not A234) );
 a74510a <=( (not A233)  and  a74509a );
 a74513a <=( (not A269)  and  (not A268) );
 a74516a <=( (not A299)  and  (not A298) );
 a74517a <=( a74516a  and  a74513a );
 a74518a <=( a74517a  and  a74510a );
 a74522a <=( A167  and  A169 );
 a74523a <=( (not A170)  and  a74522a );
 a74526a <=( (not A200)  and  A166 );
 a74529a <=( (not A203)  and  (not A202) );
 a74530a <=( a74529a  and  a74526a );
 a74531a <=( a74530a  and  a74523a );
 a74535a <=( (not A266)  and  (not A234) );
 a74536a <=( (not A233)  and  a74535a );
 a74539a <=( A298  and  (not A267) );
 a74542a <=( (not A302)  and  (not A301) );
 a74543a <=( a74542a  and  a74539a );
 a74544a <=( a74543a  and  a74536a );
 a74548a <=( A167  and  A169 );
 a74549a <=( (not A170)  and  a74548a );
 a74552a <=( (not A200)  and  A166 );
 a74555a <=( (not A203)  and  (not A202) );
 a74556a <=( a74555a  and  a74552a );
 a74557a <=( a74556a  and  a74549a );
 a74561a <=( (not A265)  and  (not A234) );
 a74562a <=( (not A233)  and  a74561a );
 a74565a <=( A298  and  (not A266) );
 a74568a <=( (not A302)  and  (not A301) );
 a74569a <=( a74568a  and  a74565a );
 a74570a <=( a74569a  and  a74562a );
 a74574a <=( A167  and  A169 );
 a74575a <=( (not A170)  and  a74574a );
 a74578a <=( (not A200)  and  A166 );
 a74581a <=( (not A203)  and  (not A202) );
 a74582a <=( a74581a  and  a74578a );
 a74583a <=( a74582a  and  a74575a );
 a74587a <=( A265  and  (not A233) );
 a74588a <=( (not A232)  and  a74587a );
 a74591a <=( A298  and  A266 );
 a74594a <=( (not A302)  and  (not A301) );
 a74595a <=( a74594a  and  a74591a );
 a74596a <=( a74595a  and  a74588a );
 a74600a <=( A167  and  A169 );
 a74601a <=( (not A170)  and  a74600a );
 a74604a <=( (not A200)  and  A166 );
 a74607a <=( (not A203)  and  (not A202) );
 a74608a <=( a74607a  and  a74604a );
 a74609a <=( a74608a  and  a74601a );
 a74613a <=( (not A266)  and  (not A233) );
 a74614a <=( (not A232)  and  a74613a );
 a74617a <=( (not A269)  and  (not A268) );
 a74620a <=( (not A300)  and  A298 );
 a74621a <=( a74620a  and  a74617a );
 a74622a <=( a74621a  and  a74614a );
 a74626a <=( A167  and  A169 );
 a74627a <=( (not A170)  and  a74626a );
 a74630a <=( (not A200)  and  A166 );
 a74633a <=( (not A203)  and  (not A202) );
 a74634a <=( a74633a  and  a74630a );
 a74635a <=( a74634a  and  a74627a );
 a74639a <=( (not A266)  and  (not A233) );
 a74640a <=( (not A232)  and  a74639a );
 a74643a <=( (not A269)  and  (not A268) );
 a74646a <=( A299  and  A298 );
 a74647a <=( a74646a  and  a74643a );
 a74648a <=( a74647a  and  a74640a );
 a74652a <=( A167  and  A169 );
 a74653a <=( (not A170)  and  a74652a );
 a74656a <=( (not A200)  and  A166 );
 a74659a <=( (not A203)  and  (not A202) );
 a74660a <=( a74659a  and  a74656a );
 a74661a <=( a74660a  and  a74653a );
 a74665a <=( (not A266)  and  (not A233) );
 a74666a <=( (not A232)  and  a74665a );
 a74669a <=( (not A269)  and  (not A268) );
 a74672a <=( (not A299)  and  (not A298) );
 a74673a <=( a74672a  and  a74669a );
 a74674a <=( a74673a  and  a74666a );
 a74678a <=( A167  and  A169 );
 a74679a <=( (not A170)  and  a74678a );
 a74682a <=( (not A200)  and  A166 );
 a74685a <=( (not A203)  and  (not A202) );
 a74686a <=( a74685a  and  a74682a );
 a74687a <=( a74686a  and  a74679a );
 a74691a <=( (not A266)  and  (not A233) );
 a74692a <=( (not A232)  and  a74691a );
 a74695a <=( A298  and  (not A267) );
 a74698a <=( (not A302)  and  (not A301) );
 a74699a <=( a74698a  and  a74695a );
 a74700a <=( a74699a  and  a74692a );
 a74704a <=( A167  and  A169 );
 a74705a <=( (not A170)  and  a74704a );
 a74708a <=( (not A200)  and  A166 );
 a74711a <=( (not A203)  and  (not A202) );
 a74712a <=( a74711a  and  a74708a );
 a74713a <=( a74712a  and  a74705a );
 a74717a <=( (not A265)  and  (not A233) );
 a74718a <=( (not A232)  and  a74717a );
 a74721a <=( A298  and  (not A266) );
 a74724a <=( (not A302)  and  (not A301) );
 a74725a <=( a74724a  and  a74721a );
 a74726a <=( a74725a  and  a74718a );
 a74730a <=( A167  and  A169 );
 a74731a <=( (not A170)  and  a74730a );
 a74734a <=( (not A200)  and  A166 );
 a74737a <=( A232  and  (not A201) );
 a74738a <=( a74737a  and  a74734a );
 a74739a <=( a74738a  and  a74731a );
 a74743a <=( (not A268)  and  A265 );
 a74744a <=( A233  and  a74743a );
 a74747a <=( (not A299)  and  (not A269) );
 a74750a <=( (not A302)  and  (not A301) );
 a74751a <=( a74750a  and  a74747a );
 a74752a <=( a74751a  and  a74744a );
 a74756a <=( A167  and  A169 );
 a74757a <=( (not A170)  and  a74756a );
 a74760a <=( (not A200)  and  A166 );
 a74763a <=( (not A233)  and  (not A201) );
 a74764a <=( a74763a  and  a74760a );
 a74765a <=( a74764a  and  a74757a );
 a74769a <=( A265  and  (not A236) );
 a74770a <=( (not A235)  and  a74769a );
 a74773a <=( A298  and  A266 );
 a74776a <=( (not A302)  and  (not A301) );
 a74777a <=( a74776a  and  a74773a );
 a74778a <=( a74777a  and  a74770a );
 a74782a <=( A167  and  A169 );
 a74783a <=( (not A170)  and  a74782a );
 a74786a <=( (not A200)  and  A166 );
 a74789a <=( (not A233)  and  (not A201) );
 a74790a <=( a74789a  and  a74786a );
 a74791a <=( a74790a  and  a74783a );
 a74795a <=( (not A266)  and  (not A236) );
 a74796a <=( (not A235)  and  a74795a );
 a74799a <=( (not A269)  and  (not A268) );
 a74802a <=( (not A300)  and  A298 );
 a74803a <=( a74802a  and  a74799a );
 a74804a <=( a74803a  and  a74796a );
 a74808a <=( A167  and  A169 );
 a74809a <=( (not A170)  and  a74808a );
 a74812a <=( (not A200)  and  A166 );
 a74815a <=( (not A233)  and  (not A201) );
 a74816a <=( a74815a  and  a74812a );
 a74817a <=( a74816a  and  a74809a );
 a74821a <=( (not A266)  and  (not A236) );
 a74822a <=( (not A235)  and  a74821a );
 a74825a <=( (not A269)  and  (not A268) );
 a74828a <=( A299  and  A298 );
 a74829a <=( a74828a  and  a74825a );
 a74830a <=( a74829a  and  a74822a );
 a74834a <=( A167  and  A169 );
 a74835a <=( (not A170)  and  a74834a );
 a74838a <=( (not A200)  and  A166 );
 a74841a <=( (not A233)  and  (not A201) );
 a74842a <=( a74841a  and  a74838a );
 a74843a <=( a74842a  and  a74835a );
 a74847a <=( (not A266)  and  (not A236) );
 a74848a <=( (not A235)  and  a74847a );
 a74851a <=( (not A269)  and  (not A268) );
 a74854a <=( (not A299)  and  (not A298) );
 a74855a <=( a74854a  and  a74851a );
 a74856a <=( a74855a  and  a74848a );
 a74860a <=( A167  and  A169 );
 a74861a <=( (not A170)  and  a74860a );
 a74864a <=( (not A200)  and  A166 );
 a74867a <=( (not A233)  and  (not A201) );
 a74868a <=( a74867a  and  a74864a );
 a74869a <=( a74868a  and  a74861a );
 a74873a <=( (not A266)  and  (not A236) );
 a74874a <=( (not A235)  and  a74873a );
 a74877a <=( A298  and  (not A267) );
 a74880a <=( (not A302)  and  (not A301) );
 a74881a <=( a74880a  and  a74877a );
 a74882a <=( a74881a  and  a74874a );
 a74886a <=( A167  and  A169 );
 a74887a <=( (not A170)  and  a74886a );
 a74890a <=( (not A200)  and  A166 );
 a74893a <=( (not A233)  and  (not A201) );
 a74894a <=( a74893a  and  a74890a );
 a74895a <=( a74894a  and  a74887a );
 a74899a <=( (not A265)  and  (not A236) );
 a74900a <=( (not A235)  and  a74899a );
 a74903a <=( A298  and  (not A266) );
 a74906a <=( (not A302)  and  (not A301) );
 a74907a <=( a74906a  and  a74903a );
 a74908a <=( a74907a  and  a74900a );
 a74912a <=( A167  and  A169 );
 a74913a <=( (not A170)  and  a74912a );
 a74916a <=( (not A200)  and  A166 );
 a74919a <=( (not A233)  and  (not A201) );
 a74920a <=( a74919a  and  a74916a );
 a74921a <=( a74920a  and  a74913a );
 a74925a <=( (not A268)  and  (not A266) );
 a74926a <=( (not A234)  and  a74925a );
 a74929a <=( A298  and  (not A269) );
 a74932a <=( (not A302)  and  (not A301) );
 a74933a <=( a74932a  and  a74929a );
 a74934a <=( a74933a  and  a74926a );
 a74938a <=( A167  and  A169 );
 a74939a <=( (not A170)  and  a74938a );
 a74942a <=( (not A200)  and  A166 );
 a74945a <=( A232  and  (not A201) );
 a74946a <=( a74945a  and  a74942a );
 a74947a <=( a74946a  and  a74939a );
 a74951a <=( A235  and  A234 );
 a74952a <=( (not A233)  and  a74951a );
 a74955a <=( (not A299)  and  A298 );
 a74958a <=( A301  and  A300 );
 a74959a <=( a74958a  and  a74955a );
 a74960a <=( a74959a  and  a74952a );
 a74964a <=( A167  and  A169 );
 a74965a <=( (not A170)  and  a74964a );
 a74968a <=( (not A200)  and  A166 );
 a74971a <=( A232  and  (not A201) );
 a74972a <=( a74971a  and  a74968a );
 a74973a <=( a74972a  and  a74965a );
 a74977a <=( A235  and  A234 );
 a74978a <=( (not A233)  and  a74977a );
 a74981a <=( (not A299)  and  A298 );
 a74984a <=( A302  and  A300 );
 a74985a <=( a74984a  and  a74981a );
 a74986a <=( a74985a  and  a74978a );
 a74990a <=( A167  and  A169 );
 a74991a <=( (not A170)  and  a74990a );
 a74994a <=( (not A200)  and  A166 );
 a74997a <=( A232  and  (not A201) );
 a74998a <=( a74997a  and  a74994a );
 a74999a <=( a74998a  and  a74991a );
 a75003a <=( A235  and  A234 );
 a75004a <=( (not A233)  and  a75003a );
 a75007a <=( (not A266)  and  A265 );
 a75010a <=( A268  and  A267 );
 a75011a <=( a75010a  and  a75007a );
 a75012a <=( a75011a  and  a75004a );
 a75016a <=( A167  and  A169 );
 a75017a <=( (not A170)  and  a75016a );
 a75020a <=( (not A200)  and  A166 );
 a75023a <=( A232  and  (not A201) );
 a75024a <=( a75023a  and  a75020a );
 a75025a <=( a75024a  and  a75017a );
 a75029a <=( A235  and  A234 );
 a75030a <=( (not A233)  and  a75029a );
 a75033a <=( (not A266)  and  A265 );
 a75036a <=( A269  and  A267 );
 a75037a <=( a75036a  and  a75033a );
 a75038a <=( a75037a  and  a75030a );
 a75042a <=( A167  and  A169 );
 a75043a <=( (not A170)  and  a75042a );
 a75046a <=( (not A200)  and  A166 );
 a75049a <=( A232  and  (not A201) );
 a75050a <=( a75049a  and  a75046a );
 a75051a <=( a75050a  and  a75043a );
 a75055a <=( A236  and  A234 );
 a75056a <=( (not A233)  and  a75055a );
 a75059a <=( (not A299)  and  A298 );
 a75062a <=( A301  and  A300 );
 a75063a <=( a75062a  and  a75059a );
 a75064a <=( a75063a  and  a75056a );
 a75068a <=( A167  and  A169 );
 a75069a <=( (not A170)  and  a75068a );
 a75072a <=( (not A200)  and  A166 );
 a75075a <=( A232  and  (not A201) );
 a75076a <=( a75075a  and  a75072a );
 a75077a <=( a75076a  and  a75069a );
 a75081a <=( A236  and  A234 );
 a75082a <=( (not A233)  and  a75081a );
 a75085a <=( (not A299)  and  A298 );
 a75088a <=( A302  and  A300 );
 a75089a <=( a75088a  and  a75085a );
 a75090a <=( a75089a  and  a75082a );
 a75094a <=( A167  and  A169 );
 a75095a <=( (not A170)  and  a75094a );
 a75098a <=( (not A200)  and  A166 );
 a75101a <=( A232  and  (not A201) );
 a75102a <=( a75101a  and  a75098a );
 a75103a <=( a75102a  and  a75095a );
 a75107a <=( A236  and  A234 );
 a75108a <=( (not A233)  and  a75107a );
 a75111a <=( (not A266)  and  A265 );
 a75114a <=( A268  and  A267 );
 a75115a <=( a75114a  and  a75111a );
 a75116a <=( a75115a  and  a75108a );
 a75120a <=( A167  and  A169 );
 a75121a <=( (not A170)  and  a75120a );
 a75124a <=( (not A200)  and  A166 );
 a75127a <=( A232  and  (not A201) );
 a75128a <=( a75127a  and  a75124a );
 a75129a <=( a75128a  and  a75121a );
 a75133a <=( A236  and  A234 );
 a75134a <=( (not A233)  and  a75133a );
 a75137a <=( (not A266)  and  A265 );
 a75140a <=( A269  and  A267 );
 a75141a <=( a75140a  and  a75137a );
 a75142a <=( a75141a  and  a75134a );
 a75146a <=( A167  and  A169 );
 a75147a <=( (not A170)  and  a75146a );
 a75150a <=( (not A200)  and  A166 );
 a75153a <=( (not A232)  and  (not A201) );
 a75154a <=( a75153a  and  a75150a );
 a75155a <=( a75154a  and  a75147a );
 a75159a <=( (not A268)  and  (not A266) );
 a75160a <=( (not A233)  and  a75159a );
 a75163a <=( A298  and  (not A269) );
 a75166a <=( (not A302)  and  (not A301) );
 a75167a <=( a75166a  and  a75163a );
 a75168a <=( a75167a  and  a75160a );
 a75172a <=( A167  and  A169 );
 a75173a <=( (not A170)  and  a75172a );
 a75176a <=( (not A199)  and  A166 );
 a75179a <=( A232  and  (not A200) );
 a75180a <=( a75179a  and  a75176a );
 a75181a <=( a75180a  and  a75173a );
 a75185a <=( (not A268)  and  A265 );
 a75186a <=( A233  and  a75185a );
 a75189a <=( (not A299)  and  (not A269) );
 a75192a <=( (not A302)  and  (not A301) );
 a75193a <=( a75192a  and  a75189a );
 a75194a <=( a75193a  and  a75186a );
 a75198a <=( A167  and  A169 );
 a75199a <=( (not A170)  and  a75198a );
 a75202a <=( (not A199)  and  A166 );
 a75205a <=( (not A233)  and  (not A200) );
 a75206a <=( a75205a  and  a75202a );
 a75207a <=( a75206a  and  a75199a );
 a75211a <=( A265  and  (not A236) );
 a75212a <=( (not A235)  and  a75211a );
 a75215a <=( A298  and  A266 );
 a75218a <=( (not A302)  and  (not A301) );
 a75219a <=( a75218a  and  a75215a );
 a75220a <=( a75219a  and  a75212a );
 a75224a <=( A167  and  A169 );
 a75225a <=( (not A170)  and  a75224a );
 a75228a <=( (not A199)  and  A166 );
 a75231a <=( (not A233)  and  (not A200) );
 a75232a <=( a75231a  and  a75228a );
 a75233a <=( a75232a  and  a75225a );
 a75237a <=( (not A266)  and  (not A236) );
 a75238a <=( (not A235)  and  a75237a );
 a75241a <=( (not A269)  and  (not A268) );
 a75244a <=( (not A300)  and  A298 );
 a75245a <=( a75244a  and  a75241a );
 a75246a <=( a75245a  and  a75238a );
 a75250a <=( A167  and  A169 );
 a75251a <=( (not A170)  and  a75250a );
 a75254a <=( (not A199)  and  A166 );
 a75257a <=( (not A233)  and  (not A200) );
 a75258a <=( a75257a  and  a75254a );
 a75259a <=( a75258a  and  a75251a );
 a75263a <=( (not A266)  and  (not A236) );
 a75264a <=( (not A235)  and  a75263a );
 a75267a <=( (not A269)  and  (not A268) );
 a75270a <=( A299  and  A298 );
 a75271a <=( a75270a  and  a75267a );
 a75272a <=( a75271a  and  a75264a );
 a75276a <=( A167  and  A169 );
 a75277a <=( (not A170)  and  a75276a );
 a75280a <=( (not A199)  and  A166 );
 a75283a <=( (not A233)  and  (not A200) );
 a75284a <=( a75283a  and  a75280a );
 a75285a <=( a75284a  and  a75277a );
 a75289a <=( (not A266)  and  (not A236) );
 a75290a <=( (not A235)  and  a75289a );
 a75293a <=( (not A269)  and  (not A268) );
 a75296a <=( (not A299)  and  (not A298) );
 a75297a <=( a75296a  and  a75293a );
 a75298a <=( a75297a  and  a75290a );
 a75302a <=( A167  and  A169 );
 a75303a <=( (not A170)  and  a75302a );
 a75306a <=( (not A199)  and  A166 );
 a75309a <=( (not A233)  and  (not A200) );
 a75310a <=( a75309a  and  a75306a );
 a75311a <=( a75310a  and  a75303a );
 a75315a <=( (not A266)  and  (not A236) );
 a75316a <=( (not A235)  and  a75315a );
 a75319a <=( A298  and  (not A267) );
 a75322a <=( (not A302)  and  (not A301) );
 a75323a <=( a75322a  and  a75319a );
 a75324a <=( a75323a  and  a75316a );
 a75328a <=( A167  and  A169 );
 a75329a <=( (not A170)  and  a75328a );
 a75332a <=( (not A199)  and  A166 );
 a75335a <=( (not A233)  and  (not A200) );
 a75336a <=( a75335a  and  a75332a );
 a75337a <=( a75336a  and  a75329a );
 a75341a <=( (not A265)  and  (not A236) );
 a75342a <=( (not A235)  and  a75341a );
 a75345a <=( A298  and  (not A266) );
 a75348a <=( (not A302)  and  (not A301) );
 a75349a <=( a75348a  and  a75345a );
 a75350a <=( a75349a  and  a75342a );
 a75354a <=( A167  and  A169 );
 a75355a <=( (not A170)  and  a75354a );
 a75358a <=( (not A199)  and  A166 );
 a75361a <=( (not A233)  and  (not A200) );
 a75362a <=( a75361a  and  a75358a );
 a75363a <=( a75362a  and  a75355a );
 a75367a <=( (not A268)  and  (not A266) );
 a75368a <=( (not A234)  and  a75367a );
 a75371a <=( A298  and  (not A269) );
 a75374a <=( (not A302)  and  (not A301) );
 a75375a <=( a75374a  and  a75371a );
 a75376a <=( a75375a  and  a75368a );
 a75380a <=( A167  and  A169 );
 a75381a <=( (not A170)  and  a75380a );
 a75384a <=( (not A199)  and  A166 );
 a75387a <=( A232  and  (not A200) );
 a75388a <=( a75387a  and  a75384a );
 a75389a <=( a75388a  and  a75381a );
 a75393a <=( A235  and  A234 );
 a75394a <=( (not A233)  and  a75393a );
 a75397a <=( (not A299)  and  A298 );
 a75400a <=( A301  and  A300 );
 a75401a <=( a75400a  and  a75397a );
 a75402a <=( a75401a  and  a75394a );
 a75406a <=( A167  and  A169 );
 a75407a <=( (not A170)  and  a75406a );
 a75410a <=( (not A199)  and  A166 );
 a75413a <=( A232  and  (not A200) );
 a75414a <=( a75413a  and  a75410a );
 a75415a <=( a75414a  and  a75407a );
 a75419a <=( A235  and  A234 );
 a75420a <=( (not A233)  and  a75419a );
 a75423a <=( (not A299)  and  A298 );
 a75426a <=( A302  and  A300 );
 a75427a <=( a75426a  and  a75423a );
 a75428a <=( a75427a  and  a75420a );
 a75432a <=( A167  and  A169 );
 a75433a <=( (not A170)  and  a75432a );
 a75436a <=( (not A199)  and  A166 );
 a75439a <=( A232  and  (not A200) );
 a75440a <=( a75439a  and  a75436a );
 a75441a <=( a75440a  and  a75433a );
 a75445a <=( A235  and  A234 );
 a75446a <=( (not A233)  and  a75445a );
 a75449a <=( (not A266)  and  A265 );
 a75452a <=( A268  and  A267 );
 a75453a <=( a75452a  and  a75449a );
 a75454a <=( a75453a  and  a75446a );
 a75458a <=( A167  and  A169 );
 a75459a <=( (not A170)  and  a75458a );
 a75462a <=( (not A199)  and  A166 );
 a75465a <=( A232  and  (not A200) );
 a75466a <=( a75465a  and  a75462a );
 a75467a <=( a75466a  and  a75459a );
 a75471a <=( A235  and  A234 );
 a75472a <=( (not A233)  and  a75471a );
 a75475a <=( (not A266)  and  A265 );
 a75478a <=( A269  and  A267 );
 a75479a <=( a75478a  and  a75475a );
 a75480a <=( a75479a  and  a75472a );
 a75484a <=( A167  and  A169 );
 a75485a <=( (not A170)  and  a75484a );
 a75488a <=( (not A199)  and  A166 );
 a75491a <=( A232  and  (not A200) );
 a75492a <=( a75491a  and  a75488a );
 a75493a <=( a75492a  and  a75485a );
 a75497a <=( A236  and  A234 );
 a75498a <=( (not A233)  and  a75497a );
 a75501a <=( (not A299)  and  A298 );
 a75504a <=( A301  and  A300 );
 a75505a <=( a75504a  and  a75501a );
 a75506a <=( a75505a  and  a75498a );
 a75510a <=( A167  and  A169 );
 a75511a <=( (not A170)  and  a75510a );
 a75514a <=( (not A199)  and  A166 );
 a75517a <=( A232  and  (not A200) );
 a75518a <=( a75517a  and  a75514a );
 a75519a <=( a75518a  and  a75511a );
 a75523a <=( A236  and  A234 );
 a75524a <=( (not A233)  and  a75523a );
 a75527a <=( (not A299)  and  A298 );
 a75530a <=( A302  and  A300 );
 a75531a <=( a75530a  and  a75527a );
 a75532a <=( a75531a  and  a75524a );
 a75536a <=( A167  and  A169 );
 a75537a <=( (not A170)  and  a75536a );
 a75540a <=( (not A199)  and  A166 );
 a75543a <=( A232  and  (not A200) );
 a75544a <=( a75543a  and  a75540a );
 a75545a <=( a75544a  and  a75537a );
 a75549a <=( A236  and  A234 );
 a75550a <=( (not A233)  and  a75549a );
 a75553a <=( (not A266)  and  A265 );
 a75556a <=( A268  and  A267 );
 a75557a <=( a75556a  and  a75553a );
 a75558a <=( a75557a  and  a75550a );
 a75562a <=( A167  and  A169 );
 a75563a <=( (not A170)  and  a75562a );
 a75566a <=( (not A199)  and  A166 );
 a75569a <=( A232  and  (not A200) );
 a75570a <=( a75569a  and  a75566a );
 a75571a <=( a75570a  and  a75563a );
 a75575a <=( A236  and  A234 );
 a75576a <=( (not A233)  and  a75575a );
 a75579a <=( (not A266)  and  A265 );
 a75582a <=( A269  and  A267 );
 a75583a <=( a75582a  and  a75579a );
 a75584a <=( a75583a  and  a75576a );
 a75588a <=( A167  and  A169 );
 a75589a <=( (not A170)  and  a75588a );
 a75592a <=( (not A199)  and  A166 );
 a75595a <=( (not A232)  and  (not A200) );
 a75596a <=( a75595a  and  a75592a );
 a75597a <=( a75596a  and  a75589a );
 a75601a <=( (not A268)  and  (not A266) );
 a75602a <=( (not A233)  and  a75601a );
 a75605a <=( A298  and  (not A269) );
 a75608a <=( (not A302)  and  (not A301) );
 a75609a <=( a75608a  and  a75605a );
 a75610a <=( a75609a  and  a75602a );
 a75614a <=( (not A167)  and  A169 );
 a75615a <=( (not A170)  and  a75614a );
 a75618a <=( A199  and  (not A166) );
 a75621a <=( A232  and  A200 );
 a75622a <=( a75621a  and  a75618a );
 a75623a <=( a75622a  and  a75615a );
 a75627a <=( (not A268)  and  A265 );
 a75628a <=( A233  and  a75627a );
 a75631a <=( (not A299)  and  (not A269) );
 a75634a <=( (not A302)  and  (not A301) );
 a75635a <=( a75634a  and  a75631a );
 a75636a <=( a75635a  and  a75628a );
 a75640a <=( (not A167)  and  A169 );
 a75641a <=( (not A170)  and  a75640a );
 a75644a <=( A199  and  (not A166) );
 a75647a <=( (not A233)  and  A200 );
 a75648a <=( a75647a  and  a75644a );
 a75649a <=( a75648a  and  a75641a );
 a75653a <=( A265  and  (not A236) );
 a75654a <=( (not A235)  and  a75653a );
 a75657a <=( A298  and  A266 );
 a75660a <=( (not A302)  and  (not A301) );
 a75661a <=( a75660a  and  a75657a );
 a75662a <=( a75661a  and  a75654a );
 a75666a <=( (not A167)  and  A169 );
 a75667a <=( (not A170)  and  a75666a );
 a75670a <=( A199  and  (not A166) );
 a75673a <=( (not A233)  and  A200 );
 a75674a <=( a75673a  and  a75670a );
 a75675a <=( a75674a  and  a75667a );
 a75679a <=( (not A266)  and  (not A236) );
 a75680a <=( (not A235)  and  a75679a );
 a75683a <=( (not A269)  and  (not A268) );
 a75686a <=( (not A300)  and  A298 );
 a75687a <=( a75686a  and  a75683a );
 a75688a <=( a75687a  and  a75680a );
 a75692a <=( (not A167)  and  A169 );
 a75693a <=( (not A170)  and  a75692a );
 a75696a <=( A199  and  (not A166) );
 a75699a <=( (not A233)  and  A200 );
 a75700a <=( a75699a  and  a75696a );
 a75701a <=( a75700a  and  a75693a );
 a75705a <=( (not A266)  and  (not A236) );
 a75706a <=( (not A235)  and  a75705a );
 a75709a <=( (not A269)  and  (not A268) );
 a75712a <=( A299  and  A298 );
 a75713a <=( a75712a  and  a75709a );
 a75714a <=( a75713a  and  a75706a );
 a75718a <=( (not A167)  and  A169 );
 a75719a <=( (not A170)  and  a75718a );
 a75722a <=( A199  and  (not A166) );
 a75725a <=( (not A233)  and  A200 );
 a75726a <=( a75725a  and  a75722a );
 a75727a <=( a75726a  and  a75719a );
 a75731a <=( (not A266)  and  (not A236) );
 a75732a <=( (not A235)  and  a75731a );
 a75735a <=( (not A269)  and  (not A268) );
 a75738a <=( (not A299)  and  (not A298) );
 a75739a <=( a75738a  and  a75735a );
 a75740a <=( a75739a  and  a75732a );
 a75744a <=( (not A167)  and  A169 );
 a75745a <=( (not A170)  and  a75744a );
 a75748a <=( A199  and  (not A166) );
 a75751a <=( (not A233)  and  A200 );
 a75752a <=( a75751a  and  a75748a );
 a75753a <=( a75752a  and  a75745a );
 a75757a <=( (not A266)  and  (not A236) );
 a75758a <=( (not A235)  and  a75757a );
 a75761a <=( A298  and  (not A267) );
 a75764a <=( (not A302)  and  (not A301) );
 a75765a <=( a75764a  and  a75761a );
 a75766a <=( a75765a  and  a75758a );
 a75770a <=( (not A167)  and  A169 );
 a75771a <=( (not A170)  and  a75770a );
 a75774a <=( A199  and  (not A166) );
 a75777a <=( (not A233)  and  A200 );
 a75778a <=( a75777a  and  a75774a );
 a75779a <=( a75778a  and  a75771a );
 a75783a <=( (not A265)  and  (not A236) );
 a75784a <=( (not A235)  and  a75783a );
 a75787a <=( A298  and  (not A266) );
 a75790a <=( (not A302)  and  (not A301) );
 a75791a <=( a75790a  and  a75787a );
 a75792a <=( a75791a  and  a75784a );
 a75796a <=( (not A167)  and  A169 );
 a75797a <=( (not A170)  and  a75796a );
 a75800a <=( A199  and  (not A166) );
 a75803a <=( (not A233)  and  A200 );
 a75804a <=( a75803a  and  a75800a );
 a75805a <=( a75804a  and  a75797a );
 a75809a <=( (not A268)  and  (not A266) );
 a75810a <=( (not A234)  and  a75809a );
 a75813a <=( A298  and  (not A269) );
 a75816a <=( (not A302)  and  (not A301) );
 a75817a <=( a75816a  and  a75813a );
 a75818a <=( a75817a  and  a75810a );
 a75822a <=( (not A167)  and  A169 );
 a75823a <=( (not A170)  and  a75822a );
 a75826a <=( A199  and  (not A166) );
 a75829a <=( A232  and  A200 );
 a75830a <=( a75829a  and  a75826a );
 a75831a <=( a75830a  and  a75823a );
 a75835a <=( A235  and  A234 );
 a75836a <=( (not A233)  and  a75835a );
 a75839a <=( (not A299)  and  A298 );
 a75842a <=( A301  and  A300 );
 a75843a <=( a75842a  and  a75839a );
 a75844a <=( a75843a  and  a75836a );
 a75848a <=( (not A167)  and  A169 );
 a75849a <=( (not A170)  and  a75848a );
 a75852a <=( A199  and  (not A166) );
 a75855a <=( A232  and  A200 );
 a75856a <=( a75855a  and  a75852a );
 a75857a <=( a75856a  and  a75849a );
 a75861a <=( A235  and  A234 );
 a75862a <=( (not A233)  and  a75861a );
 a75865a <=( (not A299)  and  A298 );
 a75868a <=( A302  and  A300 );
 a75869a <=( a75868a  and  a75865a );
 a75870a <=( a75869a  and  a75862a );
 a75874a <=( (not A167)  and  A169 );
 a75875a <=( (not A170)  and  a75874a );
 a75878a <=( A199  and  (not A166) );
 a75881a <=( A232  and  A200 );
 a75882a <=( a75881a  and  a75878a );
 a75883a <=( a75882a  and  a75875a );
 a75887a <=( A235  and  A234 );
 a75888a <=( (not A233)  and  a75887a );
 a75891a <=( (not A266)  and  A265 );
 a75894a <=( A268  and  A267 );
 a75895a <=( a75894a  and  a75891a );
 a75896a <=( a75895a  and  a75888a );
 a75900a <=( (not A167)  and  A169 );
 a75901a <=( (not A170)  and  a75900a );
 a75904a <=( A199  and  (not A166) );
 a75907a <=( A232  and  A200 );
 a75908a <=( a75907a  and  a75904a );
 a75909a <=( a75908a  and  a75901a );
 a75913a <=( A235  and  A234 );
 a75914a <=( (not A233)  and  a75913a );
 a75917a <=( (not A266)  and  A265 );
 a75920a <=( A269  and  A267 );
 a75921a <=( a75920a  and  a75917a );
 a75922a <=( a75921a  and  a75914a );
 a75926a <=( (not A167)  and  A169 );
 a75927a <=( (not A170)  and  a75926a );
 a75930a <=( A199  and  (not A166) );
 a75933a <=( A232  and  A200 );
 a75934a <=( a75933a  and  a75930a );
 a75935a <=( a75934a  and  a75927a );
 a75939a <=( A236  and  A234 );
 a75940a <=( (not A233)  and  a75939a );
 a75943a <=( (not A299)  and  A298 );
 a75946a <=( A301  and  A300 );
 a75947a <=( a75946a  and  a75943a );
 a75948a <=( a75947a  and  a75940a );
 a75952a <=( (not A167)  and  A169 );
 a75953a <=( (not A170)  and  a75952a );
 a75956a <=( A199  and  (not A166) );
 a75959a <=( A232  and  A200 );
 a75960a <=( a75959a  and  a75956a );
 a75961a <=( a75960a  and  a75953a );
 a75965a <=( A236  and  A234 );
 a75966a <=( (not A233)  and  a75965a );
 a75969a <=( (not A299)  and  A298 );
 a75972a <=( A302  and  A300 );
 a75973a <=( a75972a  and  a75969a );
 a75974a <=( a75973a  and  a75966a );
 a75978a <=( (not A167)  and  A169 );
 a75979a <=( (not A170)  and  a75978a );
 a75982a <=( A199  and  (not A166) );
 a75985a <=( A232  and  A200 );
 a75986a <=( a75985a  and  a75982a );
 a75987a <=( a75986a  and  a75979a );
 a75991a <=( A236  and  A234 );
 a75992a <=( (not A233)  and  a75991a );
 a75995a <=( (not A266)  and  A265 );
 a75998a <=( A268  and  A267 );
 a75999a <=( a75998a  and  a75995a );
 a76000a <=( a75999a  and  a75992a );
 a76004a <=( (not A167)  and  A169 );
 a76005a <=( (not A170)  and  a76004a );
 a76008a <=( A199  and  (not A166) );
 a76011a <=( A232  and  A200 );
 a76012a <=( a76011a  and  a76008a );
 a76013a <=( a76012a  and  a76005a );
 a76017a <=( A236  and  A234 );
 a76018a <=( (not A233)  and  a76017a );
 a76021a <=( (not A266)  and  A265 );
 a76024a <=( A269  and  A267 );
 a76025a <=( a76024a  and  a76021a );
 a76026a <=( a76025a  and  a76018a );
 a76030a <=( (not A167)  and  A169 );
 a76031a <=( (not A170)  and  a76030a );
 a76034a <=( A199  and  (not A166) );
 a76037a <=( (not A232)  and  A200 );
 a76038a <=( a76037a  and  a76034a );
 a76039a <=( a76038a  and  a76031a );
 a76043a <=( (not A268)  and  (not A266) );
 a76044a <=( (not A233)  and  a76043a );
 a76047a <=( A298  and  (not A269) );
 a76050a <=( (not A302)  and  (not A301) );
 a76051a <=( a76050a  and  a76047a );
 a76052a <=( a76051a  and  a76044a );
 a76056a <=( (not A167)  and  A169 );
 a76057a <=( (not A170)  and  a76056a );
 a76060a <=( (not A200)  and  (not A166) );
 a76063a <=( (not A203)  and  (not A202) );
 a76064a <=( a76063a  and  a76060a );
 a76065a <=( a76064a  and  a76057a );
 a76069a <=( A265  and  A233 );
 a76070a <=( A232  and  a76069a );
 a76073a <=( (not A269)  and  (not A268) );
 a76076a <=( (not A300)  and  (not A299) );
 a76077a <=( a76076a  and  a76073a );
 a76078a <=( a76077a  and  a76070a );
 a76082a <=( (not A167)  and  A169 );
 a76083a <=( (not A170)  and  a76082a );
 a76086a <=( (not A200)  and  (not A166) );
 a76089a <=( (not A203)  and  (not A202) );
 a76090a <=( a76089a  and  a76086a );
 a76091a <=( a76090a  and  a76083a );
 a76095a <=( A265  and  A233 );
 a76096a <=( A232  and  a76095a );
 a76099a <=( (not A269)  and  (not A268) );
 a76102a <=( A299  and  A298 );
 a76103a <=( a76102a  and  a76099a );
 a76104a <=( a76103a  and  a76096a );
 a76108a <=( (not A167)  and  A169 );
 a76109a <=( (not A170)  and  a76108a );
 a76112a <=( (not A200)  and  (not A166) );
 a76115a <=( (not A203)  and  (not A202) );
 a76116a <=( a76115a  and  a76112a );
 a76117a <=( a76116a  and  a76109a );
 a76121a <=( A265  and  A233 );
 a76122a <=( A232  and  a76121a );
 a76125a <=( (not A269)  and  (not A268) );
 a76128a <=( (not A299)  and  (not A298) );
 a76129a <=( a76128a  and  a76125a );
 a76130a <=( a76129a  and  a76122a );
 a76134a <=( (not A167)  and  A169 );
 a76135a <=( (not A170)  and  a76134a );
 a76138a <=( (not A200)  and  (not A166) );
 a76141a <=( (not A203)  and  (not A202) );
 a76142a <=( a76141a  and  a76138a );
 a76143a <=( a76142a  and  a76135a );
 a76147a <=( A265  and  A233 );
 a76148a <=( A232  and  a76147a );
 a76151a <=( (not A299)  and  (not A267) );
 a76154a <=( (not A302)  and  (not A301) );
 a76155a <=( a76154a  and  a76151a );
 a76156a <=( a76155a  and  a76148a );
 a76160a <=( (not A167)  and  A169 );
 a76161a <=( (not A170)  and  a76160a );
 a76164a <=( (not A200)  and  (not A166) );
 a76167a <=( (not A203)  and  (not A202) );
 a76168a <=( a76167a  and  a76164a );
 a76169a <=( a76168a  and  a76161a );
 a76173a <=( A265  and  A233 );
 a76174a <=( A232  and  a76173a );
 a76177a <=( (not A299)  and  A266 );
 a76180a <=( (not A302)  and  (not A301) );
 a76181a <=( a76180a  and  a76177a );
 a76182a <=( a76181a  and  a76174a );
 a76186a <=( (not A167)  and  A169 );
 a76187a <=( (not A170)  and  a76186a );
 a76190a <=( (not A200)  and  (not A166) );
 a76193a <=( (not A203)  and  (not A202) );
 a76194a <=( a76193a  and  a76190a );
 a76195a <=( a76194a  and  a76187a );
 a76199a <=( (not A265)  and  A233 );
 a76200a <=( A232  and  a76199a );
 a76203a <=( (not A299)  and  (not A266) );
 a76206a <=( (not A302)  and  (not A301) );
 a76207a <=( a76206a  and  a76203a );
 a76208a <=( a76207a  and  a76200a );
 a76212a <=( (not A167)  and  A169 );
 a76213a <=( (not A170)  and  a76212a );
 a76216a <=( (not A200)  and  (not A166) );
 a76219a <=( (not A203)  and  (not A202) );
 a76220a <=( a76219a  and  a76216a );
 a76221a <=( a76220a  and  a76213a );
 a76225a <=( (not A236)  and  (not A235) );
 a76226a <=( (not A233)  and  a76225a );
 a76229a <=( A266  and  A265 );
 a76232a <=( (not A300)  and  A298 );
 a76233a <=( a76232a  and  a76229a );
 a76234a <=( a76233a  and  a76226a );
 a76238a <=( (not A167)  and  A169 );
 a76239a <=( (not A170)  and  a76238a );
 a76242a <=( (not A200)  and  (not A166) );
 a76245a <=( (not A203)  and  (not A202) );
 a76246a <=( a76245a  and  a76242a );
 a76247a <=( a76246a  and  a76239a );
 a76251a <=( (not A236)  and  (not A235) );
 a76252a <=( (not A233)  and  a76251a );
 a76255a <=( A266  and  A265 );
 a76258a <=( A299  and  A298 );
 a76259a <=( a76258a  and  a76255a );
 a76260a <=( a76259a  and  a76252a );
 a76264a <=( (not A167)  and  A169 );
 a76265a <=( (not A170)  and  a76264a );
 a76268a <=( (not A200)  and  (not A166) );
 a76271a <=( (not A203)  and  (not A202) );
 a76272a <=( a76271a  and  a76268a );
 a76273a <=( a76272a  and  a76265a );
 a76277a <=( (not A236)  and  (not A235) );
 a76278a <=( (not A233)  and  a76277a );
 a76281a <=( A266  and  A265 );
 a76284a <=( (not A299)  and  (not A298) );
 a76285a <=( a76284a  and  a76281a );
 a76286a <=( a76285a  and  a76278a );
 a76290a <=( (not A167)  and  A169 );
 a76291a <=( (not A170)  and  a76290a );
 a76294a <=( (not A200)  and  (not A166) );
 a76297a <=( (not A203)  and  (not A202) );
 a76298a <=( a76297a  and  a76294a );
 a76299a <=( a76298a  and  a76291a );
 a76303a <=( (not A236)  and  (not A235) );
 a76304a <=( (not A233)  and  a76303a );
 a76307a <=( (not A267)  and  (not A266) );
 a76310a <=( (not A300)  and  A298 );
 a76311a <=( a76310a  and  a76307a );
 a76312a <=( a76311a  and  a76304a );
 a76316a <=( (not A167)  and  A169 );
 a76317a <=( (not A170)  and  a76316a );
 a76320a <=( (not A200)  and  (not A166) );
 a76323a <=( (not A203)  and  (not A202) );
 a76324a <=( a76323a  and  a76320a );
 a76325a <=( a76324a  and  a76317a );
 a76329a <=( (not A236)  and  (not A235) );
 a76330a <=( (not A233)  and  a76329a );
 a76333a <=( (not A267)  and  (not A266) );
 a76336a <=( A299  and  A298 );
 a76337a <=( a76336a  and  a76333a );
 a76338a <=( a76337a  and  a76330a );
 a76342a <=( (not A167)  and  A169 );
 a76343a <=( (not A170)  and  a76342a );
 a76346a <=( (not A200)  and  (not A166) );
 a76349a <=( (not A203)  and  (not A202) );
 a76350a <=( a76349a  and  a76346a );
 a76351a <=( a76350a  and  a76343a );
 a76355a <=( (not A236)  and  (not A235) );
 a76356a <=( (not A233)  and  a76355a );
 a76359a <=( (not A267)  and  (not A266) );
 a76362a <=( (not A299)  and  (not A298) );
 a76363a <=( a76362a  and  a76359a );
 a76364a <=( a76363a  and  a76356a );
 a76368a <=( (not A167)  and  A169 );
 a76369a <=( (not A170)  and  a76368a );
 a76372a <=( (not A200)  and  (not A166) );
 a76375a <=( (not A203)  and  (not A202) );
 a76376a <=( a76375a  and  a76372a );
 a76377a <=( a76376a  and  a76369a );
 a76381a <=( (not A236)  and  (not A235) );
 a76382a <=( (not A233)  and  a76381a );
 a76385a <=( (not A266)  and  (not A265) );
 a76388a <=( (not A300)  and  A298 );
 a76389a <=( a76388a  and  a76385a );
 a76390a <=( a76389a  and  a76382a );
 a76394a <=( (not A167)  and  A169 );
 a76395a <=( (not A170)  and  a76394a );
 a76398a <=( (not A200)  and  (not A166) );
 a76401a <=( (not A203)  and  (not A202) );
 a76402a <=( a76401a  and  a76398a );
 a76403a <=( a76402a  and  a76395a );
 a76407a <=( (not A236)  and  (not A235) );
 a76408a <=( (not A233)  and  a76407a );
 a76411a <=( (not A266)  and  (not A265) );
 a76414a <=( A299  and  A298 );
 a76415a <=( a76414a  and  a76411a );
 a76416a <=( a76415a  and  a76408a );
 a76420a <=( (not A167)  and  A169 );
 a76421a <=( (not A170)  and  a76420a );
 a76424a <=( (not A200)  and  (not A166) );
 a76427a <=( (not A203)  and  (not A202) );
 a76428a <=( a76427a  and  a76424a );
 a76429a <=( a76428a  and  a76421a );
 a76433a <=( (not A236)  and  (not A235) );
 a76434a <=( (not A233)  and  a76433a );
 a76437a <=( (not A266)  and  (not A265) );
 a76440a <=( (not A299)  and  (not A298) );
 a76441a <=( a76440a  and  a76437a );
 a76442a <=( a76441a  and  a76434a );
 a76446a <=( (not A167)  and  A169 );
 a76447a <=( (not A170)  and  a76446a );
 a76450a <=( (not A200)  and  (not A166) );
 a76453a <=( (not A203)  and  (not A202) );
 a76454a <=( a76453a  and  a76450a );
 a76455a <=( a76454a  and  a76447a );
 a76459a <=( A265  and  (not A234) );
 a76460a <=( (not A233)  and  a76459a );
 a76463a <=( A298  and  A266 );
 a76466a <=( (not A302)  and  (not A301) );
 a76467a <=( a76466a  and  a76463a );
 a76468a <=( a76467a  and  a76460a );
 a76472a <=( (not A167)  and  A169 );
 a76473a <=( (not A170)  and  a76472a );
 a76476a <=( (not A200)  and  (not A166) );
 a76479a <=( (not A203)  and  (not A202) );
 a76480a <=( a76479a  and  a76476a );
 a76481a <=( a76480a  and  a76473a );
 a76485a <=( (not A266)  and  (not A234) );
 a76486a <=( (not A233)  and  a76485a );
 a76489a <=( (not A269)  and  (not A268) );
 a76492a <=( (not A300)  and  A298 );
 a76493a <=( a76492a  and  a76489a );
 a76494a <=( a76493a  and  a76486a );
 a76498a <=( (not A167)  and  A169 );
 a76499a <=( (not A170)  and  a76498a );
 a76502a <=( (not A200)  and  (not A166) );
 a76505a <=( (not A203)  and  (not A202) );
 a76506a <=( a76505a  and  a76502a );
 a76507a <=( a76506a  and  a76499a );
 a76511a <=( (not A266)  and  (not A234) );
 a76512a <=( (not A233)  and  a76511a );
 a76515a <=( (not A269)  and  (not A268) );
 a76518a <=( A299  and  A298 );
 a76519a <=( a76518a  and  a76515a );
 a76520a <=( a76519a  and  a76512a );
 a76524a <=( (not A167)  and  A169 );
 a76525a <=( (not A170)  and  a76524a );
 a76528a <=( (not A200)  and  (not A166) );
 a76531a <=( (not A203)  and  (not A202) );
 a76532a <=( a76531a  and  a76528a );
 a76533a <=( a76532a  and  a76525a );
 a76537a <=( (not A266)  and  (not A234) );
 a76538a <=( (not A233)  and  a76537a );
 a76541a <=( (not A269)  and  (not A268) );
 a76544a <=( (not A299)  and  (not A298) );
 a76545a <=( a76544a  and  a76541a );
 a76546a <=( a76545a  and  a76538a );
 a76550a <=( (not A167)  and  A169 );
 a76551a <=( (not A170)  and  a76550a );
 a76554a <=( (not A200)  and  (not A166) );
 a76557a <=( (not A203)  and  (not A202) );
 a76558a <=( a76557a  and  a76554a );
 a76559a <=( a76558a  and  a76551a );
 a76563a <=( (not A266)  and  (not A234) );
 a76564a <=( (not A233)  and  a76563a );
 a76567a <=( A298  and  (not A267) );
 a76570a <=( (not A302)  and  (not A301) );
 a76571a <=( a76570a  and  a76567a );
 a76572a <=( a76571a  and  a76564a );
 a76576a <=( (not A167)  and  A169 );
 a76577a <=( (not A170)  and  a76576a );
 a76580a <=( (not A200)  and  (not A166) );
 a76583a <=( (not A203)  and  (not A202) );
 a76584a <=( a76583a  and  a76580a );
 a76585a <=( a76584a  and  a76577a );
 a76589a <=( (not A265)  and  (not A234) );
 a76590a <=( (not A233)  and  a76589a );
 a76593a <=( A298  and  (not A266) );
 a76596a <=( (not A302)  and  (not A301) );
 a76597a <=( a76596a  and  a76593a );
 a76598a <=( a76597a  and  a76590a );
 a76602a <=( (not A167)  and  A169 );
 a76603a <=( (not A170)  and  a76602a );
 a76606a <=( (not A200)  and  (not A166) );
 a76609a <=( (not A203)  and  (not A202) );
 a76610a <=( a76609a  and  a76606a );
 a76611a <=( a76610a  and  a76603a );
 a76615a <=( A265  and  (not A233) );
 a76616a <=( (not A232)  and  a76615a );
 a76619a <=( A298  and  A266 );
 a76622a <=( (not A302)  and  (not A301) );
 a76623a <=( a76622a  and  a76619a );
 a76624a <=( a76623a  and  a76616a );
 a76628a <=( (not A167)  and  A169 );
 a76629a <=( (not A170)  and  a76628a );
 a76632a <=( (not A200)  and  (not A166) );
 a76635a <=( (not A203)  and  (not A202) );
 a76636a <=( a76635a  and  a76632a );
 a76637a <=( a76636a  and  a76629a );
 a76641a <=( (not A266)  and  (not A233) );
 a76642a <=( (not A232)  and  a76641a );
 a76645a <=( (not A269)  and  (not A268) );
 a76648a <=( (not A300)  and  A298 );
 a76649a <=( a76648a  and  a76645a );
 a76650a <=( a76649a  and  a76642a );
 a76654a <=( (not A167)  and  A169 );
 a76655a <=( (not A170)  and  a76654a );
 a76658a <=( (not A200)  and  (not A166) );
 a76661a <=( (not A203)  and  (not A202) );
 a76662a <=( a76661a  and  a76658a );
 a76663a <=( a76662a  and  a76655a );
 a76667a <=( (not A266)  and  (not A233) );
 a76668a <=( (not A232)  and  a76667a );
 a76671a <=( (not A269)  and  (not A268) );
 a76674a <=( A299  and  A298 );
 a76675a <=( a76674a  and  a76671a );
 a76676a <=( a76675a  and  a76668a );
 a76680a <=( (not A167)  and  A169 );
 a76681a <=( (not A170)  and  a76680a );
 a76684a <=( (not A200)  and  (not A166) );
 a76687a <=( (not A203)  and  (not A202) );
 a76688a <=( a76687a  and  a76684a );
 a76689a <=( a76688a  and  a76681a );
 a76693a <=( (not A266)  and  (not A233) );
 a76694a <=( (not A232)  and  a76693a );
 a76697a <=( (not A269)  and  (not A268) );
 a76700a <=( (not A299)  and  (not A298) );
 a76701a <=( a76700a  and  a76697a );
 a76702a <=( a76701a  and  a76694a );
 a76706a <=( (not A167)  and  A169 );
 a76707a <=( (not A170)  and  a76706a );
 a76710a <=( (not A200)  and  (not A166) );
 a76713a <=( (not A203)  and  (not A202) );
 a76714a <=( a76713a  and  a76710a );
 a76715a <=( a76714a  and  a76707a );
 a76719a <=( (not A266)  and  (not A233) );
 a76720a <=( (not A232)  and  a76719a );
 a76723a <=( A298  and  (not A267) );
 a76726a <=( (not A302)  and  (not A301) );
 a76727a <=( a76726a  and  a76723a );
 a76728a <=( a76727a  and  a76720a );
 a76732a <=( (not A167)  and  A169 );
 a76733a <=( (not A170)  and  a76732a );
 a76736a <=( (not A200)  and  (not A166) );
 a76739a <=( (not A203)  and  (not A202) );
 a76740a <=( a76739a  and  a76736a );
 a76741a <=( a76740a  and  a76733a );
 a76745a <=( (not A265)  and  (not A233) );
 a76746a <=( (not A232)  and  a76745a );
 a76749a <=( A298  and  (not A266) );
 a76752a <=( (not A302)  and  (not A301) );
 a76753a <=( a76752a  and  a76749a );
 a76754a <=( a76753a  and  a76746a );
 a76758a <=( (not A167)  and  A169 );
 a76759a <=( (not A170)  and  a76758a );
 a76762a <=( (not A200)  and  (not A166) );
 a76765a <=( A232  and  (not A201) );
 a76766a <=( a76765a  and  a76762a );
 a76767a <=( a76766a  and  a76759a );
 a76771a <=( (not A268)  and  A265 );
 a76772a <=( A233  and  a76771a );
 a76775a <=( (not A299)  and  (not A269) );
 a76778a <=( (not A302)  and  (not A301) );
 a76779a <=( a76778a  and  a76775a );
 a76780a <=( a76779a  and  a76772a );
 a76784a <=( (not A167)  and  A169 );
 a76785a <=( (not A170)  and  a76784a );
 a76788a <=( (not A200)  and  (not A166) );
 a76791a <=( (not A233)  and  (not A201) );
 a76792a <=( a76791a  and  a76788a );
 a76793a <=( a76792a  and  a76785a );
 a76797a <=( A265  and  (not A236) );
 a76798a <=( (not A235)  and  a76797a );
 a76801a <=( A298  and  A266 );
 a76804a <=( (not A302)  and  (not A301) );
 a76805a <=( a76804a  and  a76801a );
 a76806a <=( a76805a  and  a76798a );
 a76810a <=( (not A167)  and  A169 );
 a76811a <=( (not A170)  and  a76810a );
 a76814a <=( (not A200)  and  (not A166) );
 a76817a <=( (not A233)  and  (not A201) );
 a76818a <=( a76817a  and  a76814a );
 a76819a <=( a76818a  and  a76811a );
 a76823a <=( (not A266)  and  (not A236) );
 a76824a <=( (not A235)  and  a76823a );
 a76827a <=( (not A269)  and  (not A268) );
 a76830a <=( (not A300)  and  A298 );
 a76831a <=( a76830a  and  a76827a );
 a76832a <=( a76831a  and  a76824a );
 a76836a <=( (not A167)  and  A169 );
 a76837a <=( (not A170)  and  a76836a );
 a76840a <=( (not A200)  and  (not A166) );
 a76843a <=( (not A233)  and  (not A201) );
 a76844a <=( a76843a  and  a76840a );
 a76845a <=( a76844a  and  a76837a );
 a76849a <=( (not A266)  and  (not A236) );
 a76850a <=( (not A235)  and  a76849a );
 a76853a <=( (not A269)  and  (not A268) );
 a76856a <=( A299  and  A298 );
 a76857a <=( a76856a  and  a76853a );
 a76858a <=( a76857a  and  a76850a );
 a76862a <=( (not A167)  and  A169 );
 a76863a <=( (not A170)  and  a76862a );
 a76866a <=( (not A200)  and  (not A166) );
 a76869a <=( (not A233)  and  (not A201) );
 a76870a <=( a76869a  and  a76866a );
 a76871a <=( a76870a  and  a76863a );
 a76875a <=( (not A266)  and  (not A236) );
 a76876a <=( (not A235)  and  a76875a );
 a76879a <=( (not A269)  and  (not A268) );
 a76882a <=( (not A299)  and  (not A298) );
 a76883a <=( a76882a  and  a76879a );
 a76884a <=( a76883a  and  a76876a );
 a76888a <=( (not A167)  and  A169 );
 a76889a <=( (not A170)  and  a76888a );
 a76892a <=( (not A200)  and  (not A166) );
 a76895a <=( (not A233)  and  (not A201) );
 a76896a <=( a76895a  and  a76892a );
 a76897a <=( a76896a  and  a76889a );
 a76901a <=( (not A266)  and  (not A236) );
 a76902a <=( (not A235)  and  a76901a );
 a76905a <=( A298  and  (not A267) );
 a76908a <=( (not A302)  and  (not A301) );
 a76909a <=( a76908a  and  a76905a );
 a76910a <=( a76909a  and  a76902a );
 a76914a <=( (not A167)  and  A169 );
 a76915a <=( (not A170)  and  a76914a );
 a76918a <=( (not A200)  and  (not A166) );
 a76921a <=( (not A233)  and  (not A201) );
 a76922a <=( a76921a  and  a76918a );
 a76923a <=( a76922a  and  a76915a );
 a76927a <=( (not A265)  and  (not A236) );
 a76928a <=( (not A235)  and  a76927a );
 a76931a <=( A298  and  (not A266) );
 a76934a <=( (not A302)  and  (not A301) );
 a76935a <=( a76934a  and  a76931a );
 a76936a <=( a76935a  and  a76928a );
 a76940a <=( (not A167)  and  A169 );
 a76941a <=( (not A170)  and  a76940a );
 a76944a <=( (not A200)  and  (not A166) );
 a76947a <=( (not A233)  and  (not A201) );
 a76948a <=( a76947a  and  a76944a );
 a76949a <=( a76948a  and  a76941a );
 a76953a <=( (not A268)  and  (not A266) );
 a76954a <=( (not A234)  and  a76953a );
 a76957a <=( A298  and  (not A269) );
 a76960a <=( (not A302)  and  (not A301) );
 a76961a <=( a76960a  and  a76957a );
 a76962a <=( a76961a  and  a76954a );
 a76966a <=( (not A167)  and  A169 );
 a76967a <=( (not A170)  and  a76966a );
 a76970a <=( (not A200)  and  (not A166) );
 a76973a <=( A232  and  (not A201) );
 a76974a <=( a76973a  and  a76970a );
 a76975a <=( a76974a  and  a76967a );
 a76979a <=( A235  and  A234 );
 a76980a <=( (not A233)  and  a76979a );
 a76983a <=( (not A299)  and  A298 );
 a76986a <=( A301  and  A300 );
 a76987a <=( a76986a  and  a76983a );
 a76988a <=( a76987a  and  a76980a );
 a76992a <=( (not A167)  and  A169 );
 a76993a <=( (not A170)  and  a76992a );
 a76996a <=( (not A200)  and  (not A166) );
 a76999a <=( A232  and  (not A201) );
 a77000a <=( a76999a  and  a76996a );
 a77001a <=( a77000a  and  a76993a );
 a77005a <=( A235  and  A234 );
 a77006a <=( (not A233)  and  a77005a );
 a77009a <=( (not A299)  and  A298 );
 a77012a <=( A302  and  A300 );
 a77013a <=( a77012a  and  a77009a );
 a77014a <=( a77013a  and  a77006a );
 a77018a <=( (not A167)  and  A169 );
 a77019a <=( (not A170)  and  a77018a );
 a77022a <=( (not A200)  and  (not A166) );
 a77025a <=( A232  and  (not A201) );
 a77026a <=( a77025a  and  a77022a );
 a77027a <=( a77026a  and  a77019a );
 a77031a <=( A235  and  A234 );
 a77032a <=( (not A233)  and  a77031a );
 a77035a <=( (not A266)  and  A265 );
 a77038a <=( A268  and  A267 );
 a77039a <=( a77038a  and  a77035a );
 a77040a <=( a77039a  and  a77032a );
 a77044a <=( (not A167)  and  A169 );
 a77045a <=( (not A170)  and  a77044a );
 a77048a <=( (not A200)  and  (not A166) );
 a77051a <=( A232  and  (not A201) );
 a77052a <=( a77051a  and  a77048a );
 a77053a <=( a77052a  and  a77045a );
 a77057a <=( A235  and  A234 );
 a77058a <=( (not A233)  and  a77057a );
 a77061a <=( (not A266)  and  A265 );
 a77064a <=( A269  and  A267 );
 a77065a <=( a77064a  and  a77061a );
 a77066a <=( a77065a  and  a77058a );
 a77070a <=( (not A167)  and  A169 );
 a77071a <=( (not A170)  and  a77070a );
 a77074a <=( (not A200)  and  (not A166) );
 a77077a <=( A232  and  (not A201) );
 a77078a <=( a77077a  and  a77074a );
 a77079a <=( a77078a  and  a77071a );
 a77083a <=( A236  and  A234 );
 a77084a <=( (not A233)  and  a77083a );
 a77087a <=( (not A299)  and  A298 );
 a77090a <=( A301  and  A300 );
 a77091a <=( a77090a  and  a77087a );
 a77092a <=( a77091a  and  a77084a );
 a77096a <=( (not A167)  and  A169 );
 a77097a <=( (not A170)  and  a77096a );
 a77100a <=( (not A200)  and  (not A166) );
 a77103a <=( A232  and  (not A201) );
 a77104a <=( a77103a  and  a77100a );
 a77105a <=( a77104a  and  a77097a );
 a77109a <=( A236  and  A234 );
 a77110a <=( (not A233)  and  a77109a );
 a77113a <=( (not A299)  and  A298 );
 a77116a <=( A302  and  A300 );
 a77117a <=( a77116a  and  a77113a );
 a77118a <=( a77117a  and  a77110a );
 a77122a <=( (not A167)  and  A169 );
 a77123a <=( (not A170)  and  a77122a );
 a77126a <=( (not A200)  and  (not A166) );
 a77129a <=( A232  and  (not A201) );
 a77130a <=( a77129a  and  a77126a );
 a77131a <=( a77130a  and  a77123a );
 a77135a <=( A236  and  A234 );
 a77136a <=( (not A233)  and  a77135a );
 a77139a <=( (not A266)  and  A265 );
 a77142a <=( A268  and  A267 );
 a77143a <=( a77142a  and  a77139a );
 a77144a <=( a77143a  and  a77136a );
 a77148a <=( (not A167)  and  A169 );
 a77149a <=( (not A170)  and  a77148a );
 a77152a <=( (not A200)  and  (not A166) );
 a77155a <=( A232  and  (not A201) );
 a77156a <=( a77155a  and  a77152a );
 a77157a <=( a77156a  and  a77149a );
 a77161a <=( A236  and  A234 );
 a77162a <=( (not A233)  and  a77161a );
 a77165a <=( (not A266)  and  A265 );
 a77168a <=( A269  and  A267 );
 a77169a <=( a77168a  and  a77165a );
 a77170a <=( a77169a  and  a77162a );
 a77174a <=( (not A167)  and  A169 );
 a77175a <=( (not A170)  and  a77174a );
 a77178a <=( (not A200)  and  (not A166) );
 a77181a <=( (not A232)  and  (not A201) );
 a77182a <=( a77181a  and  a77178a );
 a77183a <=( a77182a  and  a77175a );
 a77187a <=( (not A268)  and  (not A266) );
 a77188a <=( (not A233)  and  a77187a );
 a77191a <=( A298  and  (not A269) );
 a77194a <=( (not A302)  and  (not A301) );
 a77195a <=( a77194a  and  a77191a );
 a77196a <=( a77195a  and  a77188a );
 a77200a <=( (not A167)  and  A169 );
 a77201a <=( (not A170)  and  a77200a );
 a77204a <=( (not A199)  and  (not A166) );
 a77207a <=( A232  and  (not A200) );
 a77208a <=( a77207a  and  a77204a );
 a77209a <=( a77208a  and  a77201a );
 a77213a <=( (not A268)  and  A265 );
 a77214a <=( A233  and  a77213a );
 a77217a <=( (not A299)  and  (not A269) );
 a77220a <=( (not A302)  and  (not A301) );
 a77221a <=( a77220a  and  a77217a );
 a77222a <=( a77221a  and  a77214a );
 a77226a <=( (not A167)  and  A169 );
 a77227a <=( (not A170)  and  a77226a );
 a77230a <=( (not A199)  and  (not A166) );
 a77233a <=( (not A233)  and  (not A200) );
 a77234a <=( a77233a  and  a77230a );
 a77235a <=( a77234a  and  a77227a );
 a77239a <=( A265  and  (not A236) );
 a77240a <=( (not A235)  and  a77239a );
 a77243a <=( A298  and  A266 );
 a77246a <=( (not A302)  and  (not A301) );
 a77247a <=( a77246a  and  a77243a );
 a77248a <=( a77247a  and  a77240a );
 a77252a <=( (not A167)  and  A169 );
 a77253a <=( (not A170)  and  a77252a );
 a77256a <=( (not A199)  and  (not A166) );
 a77259a <=( (not A233)  and  (not A200) );
 a77260a <=( a77259a  and  a77256a );
 a77261a <=( a77260a  and  a77253a );
 a77265a <=( (not A266)  and  (not A236) );
 a77266a <=( (not A235)  and  a77265a );
 a77269a <=( (not A269)  and  (not A268) );
 a77272a <=( (not A300)  and  A298 );
 a77273a <=( a77272a  and  a77269a );
 a77274a <=( a77273a  and  a77266a );
 a77278a <=( (not A167)  and  A169 );
 a77279a <=( (not A170)  and  a77278a );
 a77282a <=( (not A199)  and  (not A166) );
 a77285a <=( (not A233)  and  (not A200) );
 a77286a <=( a77285a  and  a77282a );
 a77287a <=( a77286a  and  a77279a );
 a77291a <=( (not A266)  and  (not A236) );
 a77292a <=( (not A235)  and  a77291a );
 a77295a <=( (not A269)  and  (not A268) );
 a77298a <=( A299  and  A298 );
 a77299a <=( a77298a  and  a77295a );
 a77300a <=( a77299a  and  a77292a );
 a77304a <=( (not A167)  and  A169 );
 a77305a <=( (not A170)  and  a77304a );
 a77308a <=( (not A199)  and  (not A166) );
 a77311a <=( (not A233)  and  (not A200) );
 a77312a <=( a77311a  and  a77308a );
 a77313a <=( a77312a  and  a77305a );
 a77317a <=( (not A266)  and  (not A236) );
 a77318a <=( (not A235)  and  a77317a );
 a77321a <=( (not A269)  and  (not A268) );
 a77324a <=( (not A299)  and  (not A298) );
 a77325a <=( a77324a  and  a77321a );
 a77326a <=( a77325a  and  a77318a );
 a77330a <=( (not A167)  and  A169 );
 a77331a <=( (not A170)  and  a77330a );
 a77334a <=( (not A199)  and  (not A166) );
 a77337a <=( (not A233)  and  (not A200) );
 a77338a <=( a77337a  and  a77334a );
 a77339a <=( a77338a  and  a77331a );
 a77343a <=( (not A266)  and  (not A236) );
 a77344a <=( (not A235)  and  a77343a );
 a77347a <=( A298  and  (not A267) );
 a77350a <=( (not A302)  and  (not A301) );
 a77351a <=( a77350a  and  a77347a );
 a77352a <=( a77351a  and  a77344a );
 a77356a <=( (not A167)  and  A169 );
 a77357a <=( (not A170)  and  a77356a );
 a77360a <=( (not A199)  and  (not A166) );
 a77363a <=( (not A233)  and  (not A200) );
 a77364a <=( a77363a  and  a77360a );
 a77365a <=( a77364a  and  a77357a );
 a77369a <=( (not A265)  and  (not A236) );
 a77370a <=( (not A235)  and  a77369a );
 a77373a <=( A298  and  (not A266) );
 a77376a <=( (not A302)  and  (not A301) );
 a77377a <=( a77376a  and  a77373a );
 a77378a <=( a77377a  and  a77370a );
 a77382a <=( (not A167)  and  A169 );
 a77383a <=( (not A170)  and  a77382a );
 a77386a <=( (not A199)  and  (not A166) );
 a77389a <=( (not A233)  and  (not A200) );
 a77390a <=( a77389a  and  a77386a );
 a77391a <=( a77390a  and  a77383a );
 a77395a <=( (not A268)  and  (not A266) );
 a77396a <=( (not A234)  and  a77395a );
 a77399a <=( A298  and  (not A269) );
 a77402a <=( (not A302)  and  (not A301) );
 a77403a <=( a77402a  and  a77399a );
 a77404a <=( a77403a  and  a77396a );
 a77408a <=( (not A167)  and  A169 );
 a77409a <=( (not A170)  and  a77408a );
 a77412a <=( (not A199)  and  (not A166) );
 a77415a <=( A232  and  (not A200) );
 a77416a <=( a77415a  and  a77412a );
 a77417a <=( a77416a  and  a77409a );
 a77421a <=( A235  and  A234 );
 a77422a <=( (not A233)  and  a77421a );
 a77425a <=( (not A299)  and  A298 );
 a77428a <=( A301  and  A300 );
 a77429a <=( a77428a  and  a77425a );
 a77430a <=( a77429a  and  a77422a );
 a77434a <=( (not A167)  and  A169 );
 a77435a <=( (not A170)  and  a77434a );
 a77438a <=( (not A199)  and  (not A166) );
 a77441a <=( A232  and  (not A200) );
 a77442a <=( a77441a  and  a77438a );
 a77443a <=( a77442a  and  a77435a );
 a77447a <=( A235  and  A234 );
 a77448a <=( (not A233)  and  a77447a );
 a77451a <=( (not A299)  and  A298 );
 a77454a <=( A302  and  A300 );
 a77455a <=( a77454a  and  a77451a );
 a77456a <=( a77455a  and  a77448a );
 a77460a <=( (not A167)  and  A169 );
 a77461a <=( (not A170)  and  a77460a );
 a77464a <=( (not A199)  and  (not A166) );
 a77467a <=( A232  and  (not A200) );
 a77468a <=( a77467a  and  a77464a );
 a77469a <=( a77468a  and  a77461a );
 a77473a <=( A235  and  A234 );
 a77474a <=( (not A233)  and  a77473a );
 a77477a <=( (not A266)  and  A265 );
 a77480a <=( A268  and  A267 );
 a77481a <=( a77480a  and  a77477a );
 a77482a <=( a77481a  and  a77474a );
 a77486a <=( (not A167)  and  A169 );
 a77487a <=( (not A170)  and  a77486a );
 a77490a <=( (not A199)  and  (not A166) );
 a77493a <=( A232  and  (not A200) );
 a77494a <=( a77493a  and  a77490a );
 a77495a <=( a77494a  and  a77487a );
 a77499a <=( A235  and  A234 );
 a77500a <=( (not A233)  and  a77499a );
 a77503a <=( (not A266)  and  A265 );
 a77506a <=( A269  and  A267 );
 a77507a <=( a77506a  and  a77503a );
 a77508a <=( a77507a  and  a77500a );
 a77512a <=( (not A167)  and  A169 );
 a77513a <=( (not A170)  and  a77512a );
 a77516a <=( (not A199)  and  (not A166) );
 a77519a <=( A232  and  (not A200) );
 a77520a <=( a77519a  and  a77516a );
 a77521a <=( a77520a  and  a77513a );
 a77525a <=( A236  and  A234 );
 a77526a <=( (not A233)  and  a77525a );
 a77529a <=( (not A299)  and  A298 );
 a77532a <=( A301  and  A300 );
 a77533a <=( a77532a  and  a77529a );
 a77534a <=( a77533a  and  a77526a );
 a77538a <=( (not A167)  and  A169 );
 a77539a <=( (not A170)  and  a77538a );
 a77542a <=( (not A199)  and  (not A166) );
 a77545a <=( A232  and  (not A200) );
 a77546a <=( a77545a  and  a77542a );
 a77547a <=( a77546a  and  a77539a );
 a77551a <=( A236  and  A234 );
 a77552a <=( (not A233)  and  a77551a );
 a77555a <=( (not A299)  and  A298 );
 a77558a <=( A302  and  A300 );
 a77559a <=( a77558a  and  a77555a );
 a77560a <=( a77559a  and  a77552a );
 a77564a <=( (not A167)  and  A169 );
 a77565a <=( (not A170)  and  a77564a );
 a77568a <=( (not A199)  and  (not A166) );
 a77571a <=( A232  and  (not A200) );
 a77572a <=( a77571a  and  a77568a );
 a77573a <=( a77572a  and  a77565a );
 a77577a <=( A236  and  A234 );
 a77578a <=( (not A233)  and  a77577a );
 a77581a <=( (not A266)  and  A265 );
 a77584a <=( A268  and  A267 );
 a77585a <=( a77584a  and  a77581a );
 a77586a <=( a77585a  and  a77578a );
 a77590a <=( (not A167)  and  A169 );
 a77591a <=( (not A170)  and  a77590a );
 a77594a <=( (not A199)  and  (not A166) );
 a77597a <=( A232  and  (not A200) );
 a77598a <=( a77597a  and  a77594a );
 a77599a <=( a77598a  and  a77591a );
 a77603a <=( A236  and  A234 );
 a77604a <=( (not A233)  and  a77603a );
 a77607a <=( (not A266)  and  A265 );
 a77610a <=( A269  and  A267 );
 a77611a <=( a77610a  and  a77607a );
 a77612a <=( a77611a  and  a77604a );
 a77616a <=( (not A167)  and  A169 );
 a77617a <=( (not A170)  and  a77616a );
 a77620a <=( (not A199)  and  (not A166) );
 a77623a <=( (not A232)  and  (not A200) );
 a77624a <=( a77623a  and  a77620a );
 a77625a <=( a77624a  and  a77617a );
 a77629a <=( (not A268)  and  (not A266) );
 a77630a <=( (not A233)  and  a77629a );
 a77633a <=( A298  and  (not A269) );
 a77636a <=( (not A302)  and  (not A301) );
 a77637a <=( a77636a  and  a77633a );
 a77638a <=( a77637a  and  a77630a );
 a77642a <=( (not A166)  and  (not A167) );
 a77643a <=( (not A169)  and  a77642a );
 a77646a <=( A200  and  (not A199) );
 a77649a <=( (not A235)  and  (not A233) );
 a77650a <=( a77649a  and  a77646a );
 a77651a <=( a77650a  and  a77643a );
 a77655a <=( (not A268)  and  (not A266) );
 a77656a <=( (not A236)  and  a77655a );
 a77659a <=( A298  and  (not A269) );
 a77662a <=( (not A302)  and  (not A301) );
 a77663a <=( a77662a  and  a77659a );
 a77664a <=( a77663a  and  a77656a );
 a77668a <=( (not A166)  and  (not A167) );
 a77669a <=( (not A169)  and  a77668a );
 a77672a <=( (not A200)  and  A199 );
 a77675a <=( A202  and  A201 );
 a77676a <=( a77675a  and  a77672a );
 a77677a <=( a77676a  and  a77669a );
 a77681a <=( A265  and  A233 );
 a77682a <=( A232  and  a77681a );
 a77685a <=( (not A269)  and  (not A268) );
 a77688a <=( (not A300)  and  (not A299) );
 a77689a <=( a77688a  and  a77685a );
 a77690a <=( a77689a  and  a77682a );
 a77694a <=( (not A166)  and  (not A167) );
 a77695a <=( (not A169)  and  a77694a );
 a77698a <=( (not A200)  and  A199 );
 a77701a <=( A202  and  A201 );
 a77702a <=( a77701a  and  a77698a );
 a77703a <=( a77702a  and  a77695a );
 a77707a <=( A265  and  A233 );
 a77708a <=( A232  and  a77707a );
 a77711a <=( (not A269)  and  (not A268) );
 a77714a <=( A299  and  A298 );
 a77715a <=( a77714a  and  a77711a );
 a77716a <=( a77715a  and  a77708a );
 a77720a <=( (not A166)  and  (not A167) );
 a77721a <=( (not A169)  and  a77720a );
 a77724a <=( (not A200)  and  A199 );
 a77727a <=( A202  and  A201 );
 a77728a <=( a77727a  and  a77724a );
 a77729a <=( a77728a  and  a77721a );
 a77733a <=( A265  and  A233 );
 a77734a <=( A232  and  a77733a );
 a77737a <=( (not A269)  and  (not A268) );
 a77740a <=( (not A299)  and  (not A298) );
 a77741a <=( a77740a  and  a77737a );
 a77742a <=( a77741a  and  a77734a );
 a77746a <=( (not A166)  and  (not A167) );
 a77747a <=( (not A169)  and  a77746a );
 a77750a <=( (not A200)  and  A199 );
 a77753a <=( A202  and  A201 );
 a77754a <=( a77753a  and  a77750a );
 a77755a <=( a77754a  and  a77747a );
 a77759a <=( A265  and  A233 );
 a77760a <=( A232  and  a77759a );
 a77763a <=( (not A299)  and  (not A267) );
 a77766a <=( (not A302)  and  (not A301) );
 a77767a <=( a77766a  and  a77763a );
 a77768a <=( a77767a  and  a77760a );
 a77772a <=( (not A166)  and  (not A167) );
 a77773a <=( (not A169)  and  a77772a );
 a77776a <=( (not A200)  and  A199 );
 a77779a <=( A202  and  A201 );
 a77780a <=( a77779a  and  a77776a );
 a77781a <=( a77780a  and  a77773a );
 a77785a <=( A265  and  A233 );
 a77786a <=( A232  and  a77785a );
 a77789a <=( (not A299)  and  A266 );
 a77792a <=( (not A302)  and  (not A301) );
 a77793a <=( a77792a  and  a77789a );
 a77794a <=( a77793a  and  a77786a );
 a77798a <=( (not A166)  and  (not A167) );
 a77799a <=( (not A169)  and  a77798a );
 a77802a <=( (not A200)  and  A199 );
 a77805a <=( A202  and  A201 );
 a77806a <=( a77805a  and  a77802a );
 a77807a <=( a77806a  and  a77799a );
 a77811a <=( (not A265)  and  A233 );
 a77812a <=( A232  and  a77811a );
 a77815a <=( (not A299)  and  (not A266) );
 a77818a <=( (not A302)  and  (not A301) );
 a77819a <=( a77818a  and  a77815a );
 a77820a <=( a77819a  and  a77812a );
 a77824a <=( (not A166)  and  (not A167) );
 a77825a <=( (not A169)  and  a77824a );
 a77828a <=( (not A200)  and  A199 );
 a77831a <=( A202  and  A201 );
 a77832a <=( a77831a  and  a77828a );
 a77833a <=( a77832a  and  a77825a );
 a77837a <=( (not A236)  and  (not A235) );
 a77838a <=( (not A233)  and  a77837a );
 a77841a <=( A266  and  A265 );
 a77844a <=( (not A300)  and  A298 );
 a77845a <=( a77844a  and  a77841a );
 a77846a <=( a77845a  and  a77838a );
 a77850a <=( (not A166)  and  (not A167) );
 a77851a <=( (not A169)  and  a77850a );
 a77854a <=( (not A200)  and  A199 );
 a77857a <=( A202  and  A201 );
 a77858a <=( a77857a  and  a77854a );
 a77859a <=( a77858a  and  a77851a );
 a77863a <=( (not A236)  and  (not A235) );
 a77864a <=( (not A233)  and  a77863a );
 a77867a <=( A266  and  A265 );
 a77870a <=( A299  and  A298 );
 a77871a <=( a77870a  and  a77867a );
 a77872a <=( a77871a  and  a77864a );
 a77876a <=( (not A166)  and  (not A167) );
 a77877a <=( (not A169)  and  a77876a );
 a77880a <=( (not A200)  and  A199 );
 a77883a <=( A202  and  A201 );
 a77884a <=( a77883a  and  a77880a );
 a77885a <=( a77884a  and  a77877a );
 a77889a <=( (not A236)  and  (not A235) );
 a77890a <=( (not A233)  and  a77889a );
 a77893a <=( A266  and  A265 );
 a77896a <=( (not A299)  and  (not A298) );
 a77897a <=( a77896a  and  a77893a );
 a77898a <=( a77897a  and  a77890a );
 a77902a <=( (not A166)  and  (not A167) );
 a77903a <=( (not A169)  and  a77902a );
 a77906a <=( (not A200)  and  A199 );
 a77909a <=( A202  and  A201 );
 a77910a <=( a77909a  and  a77906a );
 a77911a <=( a77910a  and  a77903a );
 a77915a <=( (not A236)  and  (not A235) );
 a77916a <=( (not A233)  and  a77915a );
 a77919a <=( (not A267)  and  (not A266) );
 a77922a <=( (not A300)  and  A298 );
 a77923a <=( a77922a  and  a77919a );
 a77924a <=( a77923a  and  a77916a );
 a77928a <=( (not A166)  and  (not A167) );
 a77929a <=( (not A169)  and  a77928a );
 a77932a <=( (not A200)  and  A199 );
 a77935a <=( A202  and  A201 );
 a77936a <=( a77935a  and  a77932a );
 a77937a <=( a77936a  and  a77929a );
 a77941a <=( (not A236)  and  (not A235) );
 a77942a <=( (not A233)  and  a77941a );
 a77945a <=( (not A267)  and  (not A266) );
 a77948a <=( A299  and  A298 );
 a77949a <=( a77948a  and  a77945a );
 a77950a <=( a77949a  and  a77942a );
 a77954a <=( (not A166)  and  (not A167) );
 a77955a <=( (not A169)  and  a77954a );
 a77958a <=( (not A200)  and  A199 );
 a77961a <=( A202  and  A201 );
 a77962a <=( a77961a  and  a77958a );
 a77963a <=( a77962a  and  a77955a );
 a77967a <=( (not A236)  and  (not A235) );
 a77968a <=( (not A233)  and  a77967a );
 a77971a <=( (not A267)  and  (not A266) );
 a77974a <=( (not A299)  and  (not A298) );
 a77975a <=( a77974a  and  a77971a );
 a77976a <=( a77975a  and  a77968a );
 a77980a <=( (not A166)  and  (not A167) );
 a77981a <=( (not A169)  and  a77980a );
 a77984a <=( (not A200)  and  A199 );
 a77987a <=( A202  and  A201 );
 a77988a <=( a77987a  and  a77984a );
 a77989a <=( a77988a  and  a77981a );
 a77993a <=( (not A236)  and  (not A235) );
 a77994a <=( (not A233)  and  a77993a );
 a77997a <=( (not A266)  and  (not A265) );
 a78000a <=( (not A300)  and  A298 );
 a78001a <=( a78000a  and  a77997a );
 a78002a <=( a78001a  and  a77994a );
 a78006a <=( (not A166)  and  (not A167) );
 a78007a <=( (not A169)  and  a78006a );
 a78010a <=( (not A200)  and  A199 );
 a78013a <=( A202  and  A201 );
 a78014a <=( a78013a  and  a78010a );
 a78015a <=( a78014a  and  a78007a );
 a78019a <=( (not A236)  and  (not A235) );
 a78020a <=( (not A233)  and  a78019a );
 a78023a <=( (not A266)  and  (not A265) );
 a78026a <=( A299  and  A298 );
 a78027a <=( a78026a  and  a78023a );
 a78028a <=( a78027a  and  a78020a );
 a78032a <=( (not A166)  and  (not A167) );
 a78033a <=( (not A169)  and  a78032a );
 a78036a <=( (not A200)  and  A199 );
 a78039a <=( A202  and  A201 );
 a78040a <=( a78039a  and  a78036a );
 a78041a <=( a78040a  and  a78033a );
 a78045a <=( (not A236)  and  (not A235) );
 a78046a <=( (not A233)  and  a78045a );
 a78049a <=( (not A266)  and  (not A265) );
 a78052a <=( (not A299)  and  (not A298) );
 a78053a <=( a78052a  and  a78049a );
 a78054a <=( a78053a  and  a78046a );
 a78058a <=( (not A166)  and  (not A167) );
 a78059a <=( (not A169)  and  a78058a );
 a78062a <=( (not A200)  and  A199 );
 a78065a <=( A202  and  A201 );
 a78066a <=( a78065a  and  a78062a );
 a78067a <=( a78066a  and  a78059a );
 a78071a <=( A265  and  (not A234) );
 a78072a <=( (not A233)  and  a78071a );
 a78075a <=( A298  and  A266 );
 a78078a <=( (not A302)  and  (not A301) );
 a78079a <=( a78078a  and  a78075a );
 a78080a <=( a78079a  and  a78072a );
 a78084a <=( (not A166)  and  (not A167) );
 a78085a <=( (not A169)  and  a78084a );
 a78088a <=( (not A200)  and  A199 );
 a78091a <=( A202  and  A201 );
 a78092a <=( a78091a  and  a78088a );
 a78093a <=( a78092a  and  a78085a );
 a78097a <=( (not A266)  and  (not A234) );
 a78098a <=( (not A233)  and  a78097a );
 a78101a <=( (not A269)  and  (not A268) );
 a78104a <=( (not A300)  and  A298 );
 a78105a <=( a78104a  and  a78101a );
 a78106a <=( a78105a  and  a78098a );
 a78110a <=( (not A166)  and  (not A167) );
 a78111a <=( (not A169)  and  a78110a );
 a78114a <=( (not A200)  and  A199 );
 a78117a <=( A202  and  A201 );
 a78118a <=( a78117a  and  a78114a );
 a78119a <=( a78118a  and  a78111a );
 a78123a <=( (not A266)  and  (not A234) );
 a78124a <=( (not A233)  and  a78123a );
 a78127a <=( (not A269)  and  (not A268) );
 a78130a <=( A299  and  A298 );
 a78131a <=( a78130a  and  a78127a );
 a78132a <=( a78131a  and  a78124a );
 a78136a <=( (not A166)  and  (not A167) );
 a78137a <=( (not A169)  and  a78136a );
 a78140a <=( (not A200)  and  A199 );
 a78143a <=( A202  and  A201 );
 a78144a <=( a78143a  and  a78140a );
 a78145a <=( a78144a  and  a78137a );
 a78149a <=( (not A266)  and  (not A234) );
 a78150a <=( (not A233)  and  a78149a );
 a78153a <=( (not A269)  and  (not A268) );
 a78156a <=( (not A299)  and  (not A298) );
 a78157a <=( a78156a  and  a78153a );
 a78158a <=( a78157a  and  a78150a );
 a78162a <=( (not A166)  and  (not A167) );
 a78163a <=( (not A169)  and  a78162a );
 a78166a <=( (not A200)  and  A199 );
 a78169a <=( A202  and  A201 );
 a78170a <=( a78169a  and  a78166a );
 a78171a <=( a78170a  and  a78163a );
 a78175a <=( (not A266)  and  (not A234) );
 a78176a <=( (not A233)  and  a78175a );
 a78179a <=( A298  and  (not A267) );
 a78182a <=( (not A302)  and  (not A301) );
 a78183a <=( a78182a  and  a78179a );
 a78184a <=( a78183a  and  a78176a );
 a78188a <=( (not A166)  and  (not A167) );
 a78189a <=( (not A169)  and  a78188a );
 a78192a <=( (not A200)  and  A199 );
 a78195a <=( A202  and  A201 );
 a78196a <=( a78195a  and  a78192a );
 a78197a <=( a78196a  and  a78189a );
 a78201a <=( (not A265)  and  (not A234) );
 a78202a <=( (not A233)  and  a78201a );
 a78205a <=( A298  and  (not A266) );
 a78208a <=( (not A302)  and  (not A301) );
 a78209a <=( a78208a  and  a78205a );
 a78210a <=( a78209a  and  a78202a );
 a78214a <=( (not A166)  and  (not A167) );
 a78215a <=( (not A169)  and  a78214a );
 a78218a <=( (not A200)  and  A199 );
 a78221a <=( A202  and  A201 );
 a78222a <=( a78221a  and  a78218a );
 a78223a <=( a78222a  and  a78215a );
 a78227a <=( A265  and  (not A233) );
 a78228a <=( (not A232)  and  a78227a );
 a78231a <=( A298  and  A266 );
 a78234a <=( (not A302)  and  (not A301) );
 a78235a <=( a78234a  and  a78231a );
 a78236a <=( a78235a  and  a78228a );
 a78240a <=( (not A166)  and  (not A167) );
 a78241a <=( (not A169)  and  a78240a );
 a78244a <=( (not A200)  and  A199 );
 a78247a <=( A202  and  A201 );
 a78248a <=( a78247a  and  a78244a );
 a78249a <=( a78248a  and  a78241a );
 a78253a <=( (not A266)  and  (not A233) );
 a78254a <=( (not A232)  and  a78253a );
 a78257a <=( (not A269)  and  (not A268) );
 a78260a <=( (not A300)  and  A298 );
 a78261a <=( a78260a  and  a78257a );
 a78262a <=( a78261a  and  a78254a );
 a78266a <=( (not A166)  and  (not A167) );
 a78267a <=( (not A169)  and  a78266a );
 a78270a <=( (not A200)  and  A199 );
 a78273a <=( A202  and  A201 );
 a78274a <=( a78273a  and  a78270a );
 a78275a <=( a78274a  and  a78267a );
 a78279a <=( (not A266)  and  (not A233) );
 a78280a <=( (not A232)  and  a78279a );
 a78283a <=( (not A269)  and  (not A268) );
 a78286a <=( A299  and  A298 );
 a78287a <=( a78286a  and  a78283a );
 a78288a <=( a78287a  and  a78280a );
 a78292a <=( (not A166)  and  (not A167) );
 a78293a <=( (not A169)  and  a78292a );
 a78296a <=( (not A200)  and  A199 );
 a78299a <=( A202  and  A201 );
 a78300a <=( a78299a  and  a78296a );
 a78301a <=( a78300a  and  a78293a );
 a78305a <=( (not A266)  and  (not A233) );
 a78306a <=( (not A232)  and  a78305a );
 a78309a <=( (not A269)  and  (not A268) );
 a78312a <=( (not A299)  and  (not A298) );
 a78313a <=( a78312a  and  a78309a );
 a78314a <=( a78313a  and  a78306a );
 a78318a <=( (not A166)  and  (not A167) );
 a78319a <=( (not A169)  and  a78318a );
 a78322a <=( (not A200)  and  A199 );
 a78325a <=( A202  and  A201 );
 a78326a <=( a78325a  and  a78322a );
 a78327a <=( a78326a  and  a78319a );
 a78331a <=( (not A266)  and  (not A233) );
 a78332a <=( (not A232)  and  a78331a );
 a78335a <=( A298  and  (not A267) );
 a78338a <=( (not A302)  and  (not A301) );
 a78339a <=( a78338a  and  a78335a );
 a78340a <=( a78339a  and  a78332a );
 a78344a <=( (not A166)  and  (not A167) );
 a78345a <=( (not A169)  and  a78344a );
 a78348a <=( (not A200)  and  A199 );
 a78351a <=( A202  and  A201 );
 a78352a <=( a78351a  and  a78348a );
 a78353a <=( a78352a  and  a78345a );
 a78357a <=( (not A265)  and  (not A233) );
 a78358a <=( (not A232)  and  a78357a );
 a78361a <=( A298  and  (not A266) );
 a78364a <=( (not A302)  and  (not A301) );
 a78365a <=( a78364a  and  a78361a );
 a78366a <=( a78365a  and  a78358a );
 a78370a <=( (not A166)  and  (not A167) );
 a78371a <=( (not A169)  and  a78370a );
 a78374a <=( (not A200)  and  A199 );
 a78377a <=( A203  and  A201 );
 a78378a <=( a78377a  and  a78374a );
 a78379a <=( a78378a  and  a78371a );
 a78383a <=( A265  and  A233 );
 a78384a <=( A232  and  a78383a );
 a78387a <=( (not A269)  and  (not A268) );
 a78390a <=( (not A300)  and  (not A299) );
 a78391a <=( a78390a  and  a78387a );
 a78392a <=( a78391a  and  a78384a );
 a78396a <=( (not A166)  and  (not A167) );
 a78397a <=( (not A169)  and  a78396a );
 a78400a <=( (not A200)  and  A199 );
 a78403a <=( A203  and  A201 );
 a78404a <=( a78403a  and  a78400a );
 a78405a <=( a78404a  and  a78397a );
 a78409a <=( A265  and  A233 );
 a78410a <=( A232  and  a78409a );
 a78413a <=( (not A269)  and  (not A268) );
 a78416a <=( A299  and  A298 );
 a78417a <=( a78416a  and  a78413a );
 a78418a <=( a78417a  and  a78410a );
 a78422a <=( (not A166)  and  (not A167) );
 a78423a <=( (not A169)  and  a78422a );
 a78426a <=( (not A200)  and  A199 );
 a78429a <=( A203  and  A201 );
 a78430a <=( a78429a  and  a78426a );
 a78431a <=( a78430a  and  a78423a );
 a78435a <=( A265  and  A233 );
 a78436a <=( A232  and  a78435a );
 a78439a <=( (not A269)  and  (not A268) );
 a78442a <=( (not A299)  and  (not A298) );
 a78443a <=( a78442a  and  a78439a );
 a78444a <=( a78443a  and  a78436a );
 a78448a <=( (not A166)  and  (not A167) );
 a78449a <=( (not A169)  and  a78448a );
 a78452a <=( (not A200)  and  A199 );
 a78455a <=( A203  and  A201 );
 a78456a <=( a78455a  and  a78452a );
 a78457a <=( a78456a  and  a78449a );
 a78461a <=( A265  and  A233 );
 a78462a <=( A232  and  a78461a );
 a78465a <=( (not A299)  and  (not A267) );
 a78468a <=( (not A302)  and  (not A301) );
 a78469a <=( a78468a  and  a78465a );
 a78470a <=( a78469a  and  a78462a );
 a78474a <=( (not A166)  and  (not A167) );
 a78475a <=( (not A169)  and  a78474a );
 a78478a <=( (not A200)  and  A199 );
 a78481a <=( A203  and  A201 );
 a78482a <=( a78481a  and  a78478a );
 a78483a <=( a78482a  and  a78475a );
 a78487a <=( A265  and  A233 );
 a78488a <=( A232  and  a78487a );
 a78491a <=( (not A299)  and  A266 );
 a78494a <=( (not A302)  and  (not A301) );
 a78495a <=( a78494a  and  a78491a );
 a78496a <=( a78495a  and  a78488a );
 a78500a <=( (not A166)  and  (not A167) );
 a78501a <=( (not A169)  and  a78500a );
 a78504a <=( (not A200)  and  A199 );
 a78507a <=( A203  and  A201 );
 a78508a <=( a78507a  and  a78504a );
 a78509a <=( a78508a  and  a78501a );
 a78513a <=( (not A265)  and  A233 );
 a78514a <=( A232  and  a78513a );
 a78517a <=( (not A299)  and  (not A266) );
 a78520a <=( (not A302)  and  (not A301) );
 a78521a <=( a78520a  and  a78517a );
 a78522a <=( a78521a  and  a78514a );
 a78526a <=( (not A166)  and  (not A167) );
 a78527a <=( (not A169)  and  a78526a );
 a78530a <=( (not A200)  and  A199 );
 a78533a <=( A203  and  A201 );
 a78534a <=( a78533a  and  a78530a );
 a78535a <=( a78534a  and  a78527a );
 a78539a <=( (not A236)  and  (not A235) );
 a78540a <=( (not A233)  and  a78539a );
 a78543a <=( A266  and  A265 );
 a78546a <=( (not A300)  and  A298 );
 a78547a <=( a78546a  and  a78543a );
 a78548a <=( a78547a  and  a78540a );
 a78552a <=( (not A166)  and  (not A167) );
 a78553a <=( (not A169)  and  a78552a );
 a78556a <=( (not A200)  and  A199 );
 a78559a <=( A203  and  A201 );
 a78560a <=( a78559a  and  a78556a );
 a78561a <=( a78560a  and  a78553a );
 a78565a <=( (not A236)  and  (not A235) );
 a78566a <=( (not A233)  and  a78565a );
 a78569a <=( A266  and  A265 );
 a78572a <=( A299  and  A298 );
 a78573a <=( a78572a  and  a78569a );
 a78574a <=( a78573a  and  a78566a );
 a78578a <=( (not A166)  and  (not A167) );
 a78579a <=( (not A169)  and  a78578a );
 a78582a <=( (not A200)  and  A199 );
 a78585a <=( A203  and  A201 );
 a78586a <=( a78585a  and  a78582a );
 a78587a <=( a78586a  and  a78579a );
 a78591a <=( (not A236)  and  (not A235) );
 a78592a <=( (not A233)  and  a78591a );
 a78595a <=( A266  and  A265 );
 a78598a <=( (not A299)  and  (not A298) );
 a78599a <=( a78598a  and  a78595a );
 a78600a <=( a78599a  and  a78592a );
 a78604a <=( (not A166)  and  (not A167) );
 a78605a <=( (not A169)  and  a78604a );
 a78608a <=( (not A200)  and  A199 );
 a78611a <=( A203  and  A201 );
 a78612a <=( a78611a  and  a78608a );
 a78613a <=( a78612a  and  a78605a );
 a78617a <=( (not A236)  and  (not A235) );
 a78618a <=( (not A233)  and  a78617a );
 a78621a <=( (not A267)  and  (not A266) );
 a78624a <=( (not A300)  and  A298 );
 a78625a <=( a78624a  and  a78621a );
 a78626a <=( a78625a  and  a78618a );
 a78630a <=( (not A166)  and  (not A167) );
 a78631a <=( (not A169)  and  a78630a );
 a78634a <=( (not A200)  and  A199 );
 a78637a <=( A203  and  A201 );
 a78638a <=( a78637a  and  a78634a );
 a78639a <=( a78638a  and  a78631a );
 a78643a <=( (not A236)  and  (not A235) );
 a78644a <=( (not A233)  and  a78643a );
 a78647a <=( (not A267)  and  (not A266) );
 a78650a <=( A299  and  A298 );
 a78651a <=( a78650a  and  a78647a );
 a78652a <=( a78651a  and  a78644a );
 a78656a <=( (not A166)  and  (not A167) );
 a78657a <=( (not A169)  and  a78656a );
 a78660a <=( (not A200)  and  A199 );
 a78663a <=( A203  and  A201 );
 a78664a <=( a78663a  and  a78660a );
 a78665a <=( a78664a  and  a78657a );
 a78669a <=( (not A236)  and  (not A235) );
 a78670a <=( (not A233)  and  a78669a );
 a78673a <=( (not A267)  and  (not A266) );
 a78676a <=( (not A299)  and  (not A298) );
 a78677a <=( a78676a  and  a78673a );
 a78678a <=( a78677a  and  a78670a );
 a78682a <=( (not A166)  and  (not A167) );
 a78683a <=( (not A169)  and  a78682a );
 a78686a <=( (not A200)  and  A199 );
 a78689a <=( A203  and  A201 );
 a78690a <=( a78689a  and  a78686a );
 a78691a <=( a78690a  and  a78683a );
 a78695a <=( (not A236)  and  (not A235) );
 a78696a <=( (not A233)  and  a78695a );
 a78699a <=( (not A266)  and  (not A265) );
 a78702a <=( (not A300)  and  A298 );
 a78703a <=( a78702a  and  a78699a );
 a78704a <=( a78703a  and  a78696a );
 a78708a <=( (not A166)  and  (not A167) );
 a78709a <=( (not A169)  and  a78708a );
 a78712a <=( (not A200)  and  A199 );
 a78715a <=( A203  and  A201 );
 a78716a <=( a78715a  and  a78712a );
 a78717a <=( a78716a  and  a78709a );
 a78721a <=( (not A236)  and  (not A235) );
 a78722a <=( (not A233)  and  a78721a );
 a78725a <=( (not A266)  and  (not A265) );
 a78728a <=( A299  and  A298 );
 a78729a <=( a78728a  and  a78725a );
 a78730a <=( a78729a  and  a78722a );
 a78734a <=( (not A166)  and  (not A167) );
 a78735a <=( (not A169)  and  a78734a );
 a78738a <=( (not A200)  and  A199 );
 a78741a <=( A203  and  A201 );
 a78742a <=( a78741a  and  a78738a );
 a78743a <=( a78742a  and  a78735a );
 a78747a <=( (not A236)  and  (not A235) );
 a78748a <=( (not A233)  and  a78747a );
 a78751a <=( (not A266)  and  (not A265) );
 a78754a <=( (not A299)  and  (not A298) );
 a78755a <=( a78754a  and  a78751a );
 a78756a <=( a78755a  and  a78748a );
 a78760a <=( (not A166)  and  (not A167) );
 a78761a <=( (not A169)  and  a78760a );
 a78764a <=( (not A200)  and  A199 );
 a78767a <=( A203  and  A201 );
 a78768a <=( a78767a  and  a78764a );
 a78769a <=( a78768a  and  a78761a );
 a78773a <=( A265  and  (not A234) );
 a78774a <=( (not A233)  and  a78773a );
 a78777a <=( A298  and  A266 );
 a78780a <=( (not A302)  and  (not A301) );
 a78781a <=( a78780a  and  a78777a );
 a78782a <=( a78781a  and  a78774a );
 a78786a <=( (not A166)  and  (not A167) );
 a78787a <=( (not A169)  and  a78786a );
 a78790a <=( (not A200)  and  A199 );
 a78793a <=( A203  and  A201 );
 a78794a <=( a78793a  and  a78790a );
 a78795a <=( a78794a  and  a78787a );
 a78799a <=( (not A266)  and  (not A234) );
 a78800a <=( (not A233)  and  a78799a );
 a78803a <=( (not A269)  and  (not A268) );
 a78806a <=( (not A300)  and  A298 );
 a78807a <=( a78806a  and  a78803a );
 a78808a <=( a78807a  and  a78800a );
 a78812a <=( (not A166)  and  (not A167) );
 a78813a <=( (not A169)  and  a78812a );
 a78816a <=( (not A200)  and  A199 );
 a78819a <=( A203  and  A201 );
 a78820a <=( a78819a  and  a78816a );
 a78821a <=( a78820a  and  a78813a );
 a78825a <=( (not A266)  and  (not A234) );
 a78826a <=( (not A233)  and  a78825a );
 a78829a <=( (not A269)  and  (not A268) );
 a78832a <=( A299  and  A298 );
 a78833a <=( a78832a  and  a78829a );
 a78834a <=( a78833a  and  a78826a );
 a78838a <=( (not A166)  and  (not A167) );
 a78839a <=( (not A169)  and  a78838a );
 a78842a <=( (not A200)  and  A199 );
 a78845a <=( A203  and  A201 );
 a78846a <=( a78845a  and  a78842a );
 a78847a <=( a78846a  and  a78839a );
 a78851a <=( (not A266)  and  (not A234) );
 a78852a <=( (not A233)  and  a78851a );
 a78855a <=( (not A269)  and  (not A268) );
 a78858a <=( (not A299)  and  (not A298) );
 a78859a <=( a78858a  and  a78855a );
 a78860a <=( a78859a  and  a78852a );
 a78864a <=( (not A166)  and  (not A167) );
 a78865a <=( (not A169)  and  a78864a );
 a78868a <=( (not A200)  and  A199 );
 a78871a <=( A203  and  A201 );
 a78872a <=( a78871a  and  a78868a );
 a78873a <=( a78872a  and  a78865a );
 a78877a <=( (not A266)  and  (not A234) );
 a78878a <=( (not A233)  and  a78877a );
 a78881a <=( A298  and  (not A267) );
 a78884a <=( (not A302)  and  (not A301) );
 a78885a <=( a78884a  and  a78881a );
 a78886a <=( a78885a  and  a78878a );
 a78890a <=( (not A166)  and  (not A167) );
 a78891a <=( (not A169)  and  a78890a );
 a78894a <=( (not A200)  and  A199 );
 a78897a <=( A203  and  A201 );
 a78898a <=( a78897a  and  a78894a );
 a78899a <=( a78898a  and  a78891a );
 a78903a <=( (not A265)  and  (not A234) );
 a78904a <=( (not A233)  and  a78903a );
 a78907a <=( A298  and  (not A266) );
 a78910a <=( (not A302)  and  (not A301) );
 a78911a <=( a78910a  and  a78907a );
 a78912a <=( a78911a  and  a78904a );
 a78916a <=( (not A166)  and  (not A167) );
 a78917a <=( (not A169)  and  a78916a );
 a78920a <=( (not A200)  and  A199 );
 a78923a <=( A203  and  A201 );
 a78924a <=( a78923a  and  a78920a );
 a78925a <=( a78924a  and  a78917a );
 a78929a <=( A265  and  (not A233) );
 a78930a <=( (not A232)  and  a78929a );
 a78933a <=( A298  and  A266 );
 a78936a <=( (not A302)  and  (not A301) );
 a78937a <=( a78936a  and  a78933a );
 a78938a <=( a78937a  and  a78930a );
 a78942a <=( (not A166)  and  (not A167) );
 a78943a <=( (not A169)  and  a78942a );
 a78946a <=( (not A200)  and  A199 );
 a78949a <=( A203  and  A201 );
 a78950a <=( a78949a  and  a78946a );
 a78951a <=( a78950a  and  a78943a );
 a78955a <=( (not A266)  and  (not A233) );
 a78956a <=( (not A232)  and  a78955a );
 a78959a <=( (not A269)  and  (not A268) );
 a78962a <=( (not A300)  and  A298 );
 a78963a <=( a78962a  and  a78959a );
 a78964a <=( a78963a  and  a78956a );
 a78968a <=( (not A166)  and  (not A167) );
 a78969a <=( (not A169)  and  a78968a );
 a78972a <=( (not A200)  and  A199 );
 a78975a <=( A203  and  A201 );
 a78976a <=( a78975a  and  a78972a );
 a78977a <=( a78976a  and  a78969a );
 a78981a <=( (not A266)  and  (not A233) );
 a78982a <=( (not A232)  and  a78981a );
 a78985a <=( (not A269)  and  (not A268) );
 a78988a <=( A299  and  A298 );
 a78989a <=( a78988a  and  a78985a );
 a78990a <=( a78989a  and  a78982a );
 a78994a <=( (not A166)  and  (not A167) );
 a78995a <=( (not A169)  and  a78994a );
 a78998a <=( (not A200)  and  A199 );
 a79001a <=( A203  and  A201 );
 a79002a <=( a79001a  and  a78998a );
 a79003a <=( a79002a  and  a78995a );
 a79007a <=( (not A266)  and  (not A233) );
 a79008a <=( (not A232)  and  a79007a );
 a79011a <=( (not A269)  and  (not A268) );
 a79014a <=( (not A299)  and  (not A298) );
 a79015a <=( a79014a  and  a79011a );
 a79016a <=( a79015a  and  a79008a );
 a79020a <=( (not A166)  and  (not A167) );
 a79021a <=( (not A169)  and  a79020a );
 a79024a <=( (not A200)  and  A199 );
 a79027a <=( A203  and  A201 );
 a79028a <=( a79027a  and  a79024a );
 a79029a <=( a79028a  and  a79021a );
 a79033a <=( (not A266)  and  (not A233) );
 a79034a <=( (not A232)  and  a79033a );
 a79037a <=( A298  and  (not A267) );
 a79040a <=( (not A302)  and  (not A301) );
 a79041a <=( a79040a  and  a79037a );
 a79042a <=( a79041a  and  a79034a );
 a79046a <=( (not A166)  and  (not A167) );
 a79047a <=( (not A169)  and  a79046a );
 a79050a <=( (not A200)  and  A199 );
 a79053a <=( A203  and  A201 );
 a79054a <=( a79053a  and  a79050a );
 a79055a <=( a79054a  and  a79047a );
 a79059a <=( (not A265)  and  (not A233) );
 a79060a <=( (not A232)  and  a79059a );
 a79063a <=( A298  and  (not A266) );
 a79066a <=( (not A302)  and  (not A301) );
 a79067a <=( a79066a  and  a79063a );
 a79068a <=( a79067a  and  a79060a );
 a79072a <=( A167  and  (not A168) );
 a79073a <=( (not A169)  and  a79072a );
 a79076a <=( (not A199)  and  A166 );
 a79079a <=( A232  and  A200 );
 a79080a <=( a79079a  and  a79076a );
 a79081a <=( a79080a  and  a79073a );
 a79085a <=( (not A268)  and  A265 );
 a79086a <=( A233  and  a79085a );
 a79089a <=( (not A299)  and  (not A269) );
 a79092a <=( (not A302)  and  (not A301) );
 a79093a <=( a79092a  and  a79089a );
 a79094a <=( a79093a  and  a79086a );
 a79098a <=( A167  and  (not A168) );
 a79099a <=( (not A169)  and  a79098a );
 a79102a <=( (not A199)  and  A166 );
 a79105a <=( (not A233)  and  A200 );
 a79106a <=( a79105a  and  a79102a );
 a79107a <=( a79106a  and  a79099a );
 a79111a <=( A265  and  (not A236) );
 a79112a <=( (not A235)  and  a79111a );
 a79115a <=( A298  and  A266 );
 a79118a <=( (not A302)  and  (not A301) );
 a79119a <=( a79118a  and  a79115a );
 a79120a <=( a79119a  and  a79112a );
 a79124a <=( A167  and  (not A168) );
 a79125a <=( (not A169)  and  a79124a );
 a79128a <=( (not A199)  and  A166 );
 a79131a <=( (not A233)  and  A200 );
 a79132a <=( a79131a  and  a79128a );
 a79133a <=( a79132a  and  a79125a );
 a79137a <=( (not A266)  and  (not A236) );
 a79138a <=( (not A235)  and  a79137a );
 a79141a <=( (not A269)  and  (not A268) );
 a79144a <=( (not A300)  and  A298 );
 a79145a <=( a79144a  and  a79141a );
 a79146a <=( a79145a  and  a79138a );
 a79150a <=( A167  and  (not A168) );
 a79151a <=( (not A169)  and  a79150a );
 a79154a <=( (not A199)  and  A166 );
 a79157a <=( (not A233)  and  A200 );
 a79158a <=( a79157a  and  a79154a );
 a79159a <=( a79158a  and  a79151a );
 a79163a <=( (not A266)  and  (not A236) );
 a79164a <=( (not A235)  and  a79163a );
 a79167a <=( (not A269)  and  (not A268) );
 a79170a <=( A299  and  A298 );
 a79171a <=( a79170a  and  a79167a );
 a79172a <=( a79171a  and  a79164a );
 a79176a <=( A167  and  (not A168) );
 a79177a <=( (not A169)  and  a79176a );
 a79180a <=( (not A199)  and  A166 );
 a79183a <=( (not A233)  and  A200 );
 a79184a <=( a79183a  and  a79180a );
 a79185a <=( a79184a  and  a79177a );
 a79189a <=( (not A266)  and  (not A236) );
 a79190a <=( (not A235)  and  a79189a );
 a79193a <=( (not A269)  and  (not A268) );
 a79196a <=( (not A299)  and  (not A298) );
 a79197a <=( a79196a  and  a79193a );
 a79198a <=( a79197a  and  a79190a );
 a79202a <=( A167  and  (not A168) );
 a79203a <=( (not A169)  and  a79202a );
 a79206a <=( (not A199)  and  A166 );
 a79209a <=( (not A233)  and  A200 );
 a79210a <=( a79209a  and  a79206a );
 a79211a <=( a79210a  and  a79203a );
 a79215a <=( (not A266)  and  (not A236) );
 a79216a <=( (not A235)  and  a79215a );
 a79219a <=( A298  and  (not A267) );
 a79222a <=( (not A302)  and  (not A301) );
 a79223a <=( a79222a  and  a79219a );
 a79224a <=( a79223a  and  a79216a );
 a79228a <=( A167  and  (not A168) );
 a79229a <=( (not A169)  and  a79228a );
 a79232a <=( (not A199)  and  A166 );
 a79235a <=( (not A233)  and  A200 );
 a79236a <=( a79235a  and  a79232a );
 a79237a <=( a79236a  and  a79229a );
 a79241a <=( (not A265)  and  (not A236) );
 a79242a <=( (not A235)  and  a79241a );
 a79245a <=( A298  and  (not A266) );
 a79248a <=( (not A302)  and  (not A301) );
 a79249a <=( a79248a  and  a79245a );
 a79250a <=( a79249a  and  a79242a );
 a79254a <=( A167  and  (not A168) );
 a79255a <=( (not A169)  and  a79254a );
 a79258a <=( (not A199)  and  A166 );
 a79261a <=( (not A233)  and  A200 );
 a79262a <=( a79261a  and  a79258a );
 a79263a <=( a79262a  and  a79255a );
 a79267a <=( (not A268)  and  (not A266) );
 a79268a <=( (not A234)  and  a79267a );
 a79271a <=( A298  and  (not A269) );
 a79274a <=( (not A302)  and  (not A301) );
 a79275a <=( a79274a  and  a79271a );
 a79276a <=( a79275a  and  a79268a );
 a79280a <=( A167  and  (not A168) );
 a79281a <=( (not A169)  and  a79280a );
 a79284a <=( (not A199)  and  A166 );
 a79287a <=( A232  and  A200 );
 a79288a <=( a79287a  and  a79284a );
 a79289a <=( a79288a  and  a79281a );
 a79293a <=( A235  and  A234 );
 a79294a <=( (not A233)  and  a79293a );
 a79297a <=( (not A299)  and  A298 );
 a79300a <=( A301  and  A300 );
 a79301a <=( a79300a  and  a79297a );
 a79302a <=( a79301a  and  a79294a );
 a79306a <=( A167  and  (not A168) );
 a79307a <=( (not A169)  and  a79306a );
 a79310a <=( (not A199)  and  A166 );
 a79313a <=( A232  and  A200 );
 a79314a <=( a79313a  and  a79310a );
 a79315a <=( a79314a  and  a79307a );
 a79319a <=( A235  and  A234 );
 a79320a <=( (not A233)  and  a79319a );
 a79323a <=( (not A299)  and  A298 );
 a79326a <=( A302  and  A300 );
 a79327a <=( a79326a  and  a79323a );
 a79328a <=( a79327a  and  a79320a );
 a79332a <=( A167  and  (not A168) );
 a79333a <=( (not A169)  and  a79332a );
 a79336a <=( (not A199)  and  A166 );
 a79339a <=( A232  and  A200 );
 a79340a <=( a79339a  and  a79336a );
 a79341a <=( a79340a  and  a79333a );
 a79345a <=( A235  and  A234 );
 a79346a <=( (not A233)  and  a79345a );
 a79349a <=( (not A266)  and  A265 );
 a79352a <=( A268  and  A267 );
 a79353a <=( a79352a  and  a79349a );
 a79354a <=( a79353a  and  a79346a );
 a79358a <=( A167  and  (not A168) );
 a79359a <=( (not A169)  and  a79358a );
 a79362a <=( (not A199)  and  A166 );
 a79365a <=( A232  and  A200 );
 a79366a <=( a79365a  and  a79362a );
 a79367a <=( a79366a  and  a79359a );
 a79371a <=( A235  and  A234 );
 a79372a <=( (not A233)  and  a79371a );
 a79375a <=( (not A266)  and  A265 );
 a79378a <=( A269  and  A267 );
 a79379a <=( a79378a  and  a79375a );
 a79380a <=( a79379a  and  a79372a );
 a79384a <=( A167  and  (not A168) );
 a79385a <=( (not A169)  and  a79384a );
 a79388a <=( (not A199)  and  A166 );
 a79391a <=( A232  and  A200 );
 a79392a <=( a79391a  and  a79388a );
 a79393a <=( a79392a  and  a79385a );
 a79397a <=( A236  and  A234 );
 a79398a <=( (not A233)  and  a79397a );
 a79401a <=( (not A299)  and  A298 );
 a79404a <=( A301  and  A300 );
 a79405a <=( a79404a  and  a79401a );
 a79406a <=( a79405a  and  a79398a );
 a79410a <=( A167  and  (not A168) );
 a79411a <=( (not A169)  and  a79410a );
 a79414a <=( (not A199)  and  A166 );
 a79417a <=( A232  and  A200 );
 a79418a <=( a79417a  and  a79414a );
 a79419a <=( a79418a  and  a79411a );
 a79423a <=( A236  and  A234 );
 a79424a <=( (not A233)  and  a79423a );
 a79427a <=( (not A299)  and  A298 );
 a79430a <=( A302  and  A300 );
 a79431a <=( a79430a  and  a79427a );
 a79432a <=( a79431a  and  a79424a );
 a79436a <=( A167  and  (not A168) );
 a79437a <=( (not A169)  and  a79436a );
 a79440a <=( (not A199)  and  A166 );
 a79443a <=( A232  and  A200 );
 a79444a <=( a79443a  and  a79440a );
 a79445a <=( a79444a  and  a79437a );
 a79449a <=( A236  and  A234 );
 a79450a <=( (not A233)  and  a79449a );
 a79453a <=( (not A266)  and  A265 );
 a79456a <=( A268  and  A267 );
 a79457a <=( a79456a  and  a79453a );
 a79458a <=( a79457a  and  a79450a );
 a79462a <=( A167  and  (not A168) );
 a79463a <=( (not A169)  and  a79462a );
 a79466a <=( (not A199)  and  A166 );
 a79469a <=( A232  and  A200 );
 a79470a <=( a79469a  and  a79466a );
 a79471a <=( a79470a  and  a79463a );
 a79475a <=( A236  and  A234 );
 a79476a <=( (not A233)  and  a79475a );
 a79479a <=( (not A266)  and  A265 );
 a79482a <=( A269  and  A267 );
 a79483a <=( a79482a  and  a79479a );
 a79484a <=( a79483a  and  a79476a );
 a79488a <=( A167  and  (not A168) );
 a79489a <=( (not A169)  and  a79488a );
 a79492a <=( (not A199)  and  A166 );
 a79495a <=( (not A232)  and  A200 );
 a79496a <=( a79495a  and  a79492a );
 a79497a <=( a79496a  and  a79489a );
 a79501a <=( (not A268)  and  (not A266) );
 a79502a <=( (not A233)  and  a79501a );
 a79505a <=( A298  and  (not A269) );
 a79508a <=( (not A302)  and  (not A301) );
 a79509a <=( a79508a  and  a79505a );
 a79510a <=( a79509a  and  a79502a );
 a79514a <=( A167  and  (not A168) );
 a79515a <=( (not A169)  and  a79514a );
 a79518a <=( A199  and  A166 );
 a79521a <=( A201  and  (not A200) );
 a79522a <=( a79521a  and  a79518a );
 a79523a <=( a79522a  and  a79515a );
 a79527a <=( A233  and  A232 );
 a79528a <=( A202  and  a79527a );
 a79531a <=( (not A267)  and  A265 );
 a79534a <=( (not A300)  and  (not A299) );
 a79535a <=( a79534a  and  a79531a );
 a79536a <=( a79535a  and  a79528a );
 a79540a <=( A167  and  (not A168) );
 a79541a <=( (not A169)  and  a79540a );
 a79544a <=( A199  and  A166 );
 a79547a <=( A201  and  (not A200) );
 a79548a <=( a79547a  and  a79544a );
 a79549a <=( a79548a  and  a79541a );
 a79553a <=( A233  and  A232 );
 a79554a <=( A202  and  a79553a );
 a79557a <=( (not A267)  and  A265 );
 a79560a <=( A299  and  A298 );
 a79561a <=( a79560a  and  a79557a );
 a79562a <=( a79561a  and  a79554a );
 a79566a <=( A167  and  (not A168) );
 a79567a <=( (not A169)  and  a79566a );
 a79570a <=( A199  and  A166 );
 a79573a <=( A201  and  (not A200) );
 a79574a <=( a79573a  and  a79570a );
 a79575a <=( a79574a  and  a79567a );
 a79579a <=( A233  and  A232 );
 a79580a <=( A202  and  a79579a );
 a79583a <=( (not A267)  and  A265 );
 a79586a <=( (not A299)  and  (not A298) );
 a79587a <=( a79586a  and  a79583a );
 a79588a <=( a79587a  and  a79580a );
 a79592a <=( A167  and  (not A168) );
 a79593a <=( (not A169)  and  a79592a );
 a79596a <=( A199  and  A166 );
 a79599a <=( A201  and  (not A200) );
 a79600a <=( a79599a  and  a79596a );
 a79601a <=( a79600a  and  a79593a );
 a79605a <=( A233  and  A232 );
 a79606a <=( A202  and  a79605a );
 a79609a <=( A266  and  A265 );
 a79612a <=( (not A300)  and  (not A299) );
 a79613a <=( a79612a  and  a79609a );
 a79614a <=( a79613a  and  a79606a );
 a79618a <=( A167  and  (not A168) );
 a79619a <=( (not A169)  and  a79618a );
 a79622a <=( A199  and  A166 );
 a79625a <=( A201  and  (not A200) );
 a79626a <=( a79625a  and  a79622a );
 a79627a <=( a79626a  and  a79619a );
 a79631a <=( A233  and  A232 );
 a79632a <=( A202  and  a79631a );
 a79635a <=( A266  and  A265 );
 a79638a <=( A299  and  A298 );
 a79639a <=( a79638a  and  a79635a );
 a79640a <=( a79639a  and  a79632a );
 a79644a <=( A167  and  (not A168) );
 a79645a <=( (not A169)  and  a79644a );
 a79648a <=( A199  and  A166 );
 a79651a <=( A201  and  (not A200) );
 a79652a <=( a79651a  and  a79648a );
 a79653a <=( a79652a  and  a79645a );
 a79657a <=( A233  and  A232 );
 a79658a <=( A202  and  a79657a );
 a79661a <=( A266  and  A265 );
 a79664a <=( (not A299)  and  (not A298) );
 a79665a <=( a79664a  and  a79661a );
 a79666a <=( a79665a  and  a79658a );
 a79670a <=( A167  and  (not A168) );
 a79671a <=( (not A169)  and  a79670a );
 a79674a <=( A199  and  A166 );
 a79677a <=( A201  and  (not A200) );
 a79678a <=( a79677a  and  a79674a );
 a79679a <=( a79678a  and  a79671a );
 a79683a <=( A233  and  A232 );
 a79684a <=( A202  and  a79683a );
 a79687a <=( (not A266)  and  (not A265) );
 a79690a <=( (not A300)  and  (not A299) );
 a79691a <=( a79690a  and  a79687a );
 a79692a <=( a79691a  and  a79684a );
 a79696a <=( A167  and  (not A168) );
 a79697a <=( (not A169)  and  a79696a );
 a79700a <=( A199  and  A166 );
 a79703a <=( A201  and  (not A200) );
 a79704a <=( a79703a  and  a79700a );
 a79705a <=( a79704a  and  a79697a );
 a79709a <=( A233  and  A232 );
 a79710a <=( A202  and  a79709a );
 a79713a <=( (not A266)  and  (not A265) );
 a79716a <=( A299  and  A298 );
 a79717a <=( a79716a  and  a79713a );
 a79718a <=( a79717a  and  a79710a );
 a79722a <=( A167  and  (not A168) );
 a79723a <=( (not A169)  and  a79722a );
 a79726a <=( A199  and  A166 );
 a79729a <=( A201  and  (not A200) );
 a79730a <=( a79729a  and  a79726a );
 a79731a <=( a79730a  and  a79723a );
 a79735a <=( A233  and  A232 );
 a79736a <=( A202  and  a79735a );
 a79739a <=( (not A266)  and  (not A265) );
 a79742a <=( (not A299)  and  (not A298) );
 a79743a <=( a79742a  and  a79739a );
 a79744a <=( a79743a  and  a79736a );
 a79748a <=( A167  and  (not A168) );
 a79749a <=( (not A169)  and  a79748a );
 a79752a <=( A199  and  A166 );
 a79755a <=( A201  and  (not A200) );
 a79756a <=( a79755a  and  a79752a );
 a79757a <=( a79756a  and  a79749a );
 a79761a <=( A233  and  (not A232) );
 a79762a <=( A202  and  a79761a );
 a79765a <=( (not A299)  and  A298 );
 a79768a <=( A301  and  A300 );
 a79769a <=( a79768a  and  a79765a );
 a79770a <=( a79769a  and  a79762a );
 a79774a <=( A167  and  (not A168) );
 a79775a <=( (not A169)  and  a79774a );
 a79778a <=( A199  and  A166 );
 a79781a <=( A201  and  (not A200) );
 a79782a <=( a79781a  and  a79778a );
 a79783a <=( a79782a  and  a79775a );
 a79787a <=( A233  and  (not A232) );
 a79788a <=( A202  and  a79787a );
 a79791a <=( (not A299)  and  A298 );
 a79794a <=( A302  and  A300 );
 a79795a <=( a79794a  and  a79791a );
 a79796a <=( a79795a  and  a79788a );
 a79800a <=( A167  and  (not A168) );
 a79801a <=( (not A169)  and  a79800a );
 a79804a <=( A199  and  A166 );
 a79807a <=( A201  and  (not A200) );
 a79808a <=( a79807a  and  a79804a );
 a79809a <=( a79808a  and  a79801a );
 a79813a <=( A233  and  (not A232) );
 a79814a <=( A202  and  a79813a );
 a79817a <=( (not A266)  and  A265 );
 a79820a <=( A268  and  A267 );
 a79821a <=( a79820a  and  a79817a );
 a79822a <=( a79821a  and  a79814a );
 a79826a <=( A167  and  (not A168) );
 a79827a <=( (not A169)  and  a79826a );
 a79830a <=( A199  and  A166 );
 a79833a <=( A201  and  (not A200) );
 a79834a <=( a79833a  and  a79830a );
 a79835a <=( a79834a  and  a79827a );
 a79839a <=( A233  and  (not A232) );
 a79840a <=( A202  and  a79839a );
 a79843a <=( (not A266)  and  A265 );
 a79846a <=( A269  and  A267 );
 a79847a <=( a79846a  and  a79843a );
 a79848a <=( a79847a  and  a79840a );
 a79852a <=( A167  and  (not A168) );
 a79853a <=( (not A169)  and  a79852a );
 a79856a <=( A199  and  A166 );
 a79859a <=( A201  and  (not A200) );
 a79860a <=( a79859a  and  a79856a );
 a79861a <=( a79860a  and  a79853a );
 a79865a <=( (not A234)  and  (not A233) );
 a79866a <=( A202  and  a79865a );
 a79869a <=( A266  and  A265 );
 a79872a <=( (not A300)  and  A298 );
 a79873a <=( a79872a  and  a79869a );
 a79874a <=( a79873a  and  a79866a );
 a79878a <=( A167  and  (not A168) );
 a79879a <=( (not A169)  and  a79878a );
 a79882a <=( A199  and  A166 );
 a79885a <=( A201  and  (not A200) );
 a79886a <=( a79885a  and  a79882a );
 a79887a <=( a79886a  and  a79879a );
 a79891a <=( (not A234)  and  (not A233) );
 a79892a <=( A202  and  a79891a );
 a79895a <=( A266  and  A265 );
 a79898a <=( A299  and  A298 );
 a79899a <=( a79898a  and  a79895a );
 a79900a <=( a79899a  and  a79892a );
 a79904a <=( A167  and  (not A168) );
 a79905a <=( (not A169)  and  a79904a );
 a79908a <=( A199  and  A166 );
 a79911a <=( A201  and  (not A200) );
 a79912a <=( a79911a  and  a79908a );
 a79913a <=( a79912a  and  a79905a );
 a79917a <=( (not A234)  and  (not A233) );
 a79918a <=( A202  and  a79917a );
 a79921a <=( A266  and  A265 );
 a79924a <=( (not A299)  and  (not A298) );
 a79925a <=( a79924a  and  a79921a );
 a79926a <=( a79925a  and  a79918a );
 a79930a <=( A167  and  (not A168) );
 a79931a <=( (not A169)  and  a79930a );
 a79934a <=( A199  and  A166 );
 a79937a <=( A201  and  (not A200) );
 a79938a <=( a79937a  and  a79934a );
 a79939a <=( a79938a  and  a79931a );
 a79943a <=( (not A234)  and  (not A233) );
 a79944a <=( A202  and  a79943a );
 a79947a <=( (not A267)  and  (not A266) );
 a79950a <=( (not A300)  and  A298 );
 a79951a <=( a79950a  and  a79947a );
 a79952a <=( a79951a  and  a79944a );
 a79956a <=( A167  and  (not A168) );
 a79957a <=( (not A169)  and  a79956a );
 a79960a <=( A199  and  A166 );
 a79963a <=( A201  and  (not A200) );
 a79964a <=( a79963a  and  a79960a );
 a79965a <=( a79964a  and  a79957a );
 a79969a <=( (not A234)  and  (not A233) );
 a79970a <=( A202  and  a79969a );
 a79973a <=( (not A267)  and  (not A266) );
 a79976a <=( A299  and  A298 );
 a79977a <=( a79976a  and  a79973a );
 a79978a <=( a79977a  and  a79970a );
 a79982a <=( A167  and  (not A168) );
 a79983a <=( (not A169)  and  a79982a );
 a79986a <=( A199  and  A166 );
 a79989a <=( A201  and  (not A200) );
 a79990a <=( a79989a  and  a79986a );
 a79991a <=( a79990a  and  a79983a );
 a79995a <=( (not A234)  and  (not A233) );
 a79996a <=( A202  and  a79995a );
 a79999a <=( (not A267)  and  (not A266) );
 a80002a <=( (not A299)  and  (not A298) );
 a80003a <=( a80002a  and  a79999a );
 a80004a <=( a80003a  and  a79996a );
 a80008a <=( A167  and  (not A168) );
 a80009a <=( (not A169)  and  a80008a );
 a80012a <=( A199  and  A166 );
 a80015a <=( A201  and  (not A200) );
 a80016a <=( a80015a  and  a80012a );
 a80017a <=( a80016a  and  a80009a );
 a80021a <=( (not A234)  and  (not A233) );
 a80022a <=( A202  and  a80021a );
 a80025a <=( (not A266)  and  (not A265) );
 a80028a <=( (not A300)  and  A298 );
 a80029a <=( a80028a  and  a80025a );
 a80030a <=( a80029a  and  a80022a );
 a80034a <=( A167  and  (not A168) );
 a80035a <=( (not A169)  and  a80034a );
 a80038a <=( A199  and  A166 );
 a80041a <=( A201  and  (not A200) );
 a80042a <=( a80041a  and  a80038a );
 a80043a <=( a80042a  and  a80035a );
 a80047a <=( (not A234)  and  (not A233) );
 a80048a <=( A202  and  a80047a );
 a80051a <=( (not A266)  and  (not A265) );
 a80054a <=( A299  and  A298 );
 a80055a <=( a80054a  and  a80051a );
 a80056a <=( a80055a  and  a80048a );
 a80060a <=( A167  and  (not A168) );
 a80061a <=( (not A169)  and  a80060a );
 a80064a <=( A199  and  A166 );
 a80067a <=( A201  and  (not A200) );
 a80068a <=( a80067a  and  a80064a );
 a80069a <=( a80068a  and  a80061a );
 a80073a <=( (not A234)  and  (not A233) );
 a80074a <=( A202  and  a80073a );
 a80077a <=( (not A266)  and  (not A265) );
 a80080a <=( (not A299)  and  (not A298) );
 a80081a <=( a80080a  and  a80077a );
 a80082a <=( a80081a  and  a80074a );
 a80086a <=( A167  and  (not A168) );
 a80087a <=( (not A169)  and  a80086a );
 a80090a <=( A199  and  A166 );
 a80093a <=( A201  and  (not A200) );
 a80094a <=( a80093a  and  a80090a );
 a80095a <=( a80094a  and  a80087a );
 a80099a <=( (not A233)  and  A232 );
 a80100a <=( A202  and  a80099a );
 a80103a <=( A235  and  A234 );
 a80106a <=( A299  and  (not A298) );
 a80107a <=( a80106a  and  a80103a );
 a80108a <=( a80107a  and  a80100a );
 a80112a <=( A167  and  (not A168) );
 a80113a <=( (not A169)  and  a80112a );
 a80116a <=( A199  and  A166 );
 a80119a <=( A201  and  (not A200) );
 a80120a <=( a80119a  and  a80116a );
 a80121a <=( a80120a  and  a80113a );
 a80125a <=( (not A233)  and  A232 );
 a80126a <=( A202  and  a80125a );
 a80129a <=( A235  and  A234 );
 a80132a <=( A266  and  (not A265) );
 a80133a <=( a80132a  and  a80129a );
 a80134a <=( a80133a  and  a80126a );
 a80138a <=( A167  and  (not A168) );
 a80139a <=( (not A169)  and  a80138a );
 a80142a <=( A199  and  A166 );
 a80145a <=( A201  and  (not A200) );
 a80146a <=( a80145a  and  a80142a );
 a80147a <=( a80146a  and  a80139a );
 a80151a <=( (not A233)  and  A232 );
 a80152a <=( A202  and  a80151a );
 a80155a <=( A236  and  A234 );
 a80158a <=( A299  and  (not A298) );
 a80159a <=( a80158a  and  a80155a );
 a80160a <=( a80159a  and  a80152a );
 a80164a <=( A167  and  (not A168) );
 a80165a <=( (not A169)  and  a80164a );
 a80168a <=( A199  and  A166 );
 a80171a <=( A201  and  (not A200) );
 a80172a <=( a80171a  and  a80168a );
 a80173a <=( a80172a  and  a80165a );
 a80177a <=( (not A233)  and  A232 );
 a80178a <=( A202  and  a80177a );
 a80181a <=( A236  and  A234 );
 a80184a <=( A266  and  (not A265) );
 a80185a <=( a80184a  and  a80181a );
 a80186a <=( a80185a  and  a80178a );
 a80190a <=( A167  and  (not A168) );
 a80191a <=( (not A169)  and  a80190a );
 a80194a <=( A199  and  A166 );
 a80197a <=( A201  and  (not A200) );
 a80198a <=( a80197a  and  a80194a );
 a80199a <=( a80198a  and  a80191a );
 a80203a <=( (not A233)  and  (not A232) );
 a80204a <=( A202  and  a80203a );
 a80207a <=( A266  and  A265 );
 a80210a <=( (not A300)  and  A298 );
 a80211a <=( a80210a  and  a80207a );
 a80212a <=( a80211a  and  a80204a );
 a80216a <=( A167  and  (not A168) );
 a80217a <=( (not A169)  and  a80216a );
 a80220a <=( A199  and  A166 );
 a80223a <=( A201  and  (not A200) );
 a80224a <=( a80223a  and  a80220a );
 a80225a <=( a80224a  and  a80217a );
 a80229a <=( (not A233)  and  (not A232) );
 a80230a <=( A202  and  a80229a );
 a80233a <=( A266  and  A265 );
 a80236a <=( A299  and  A298 );
 a80237a <=( a80236a  and  a80233a );
 a80238a <=( a80237a  and  a80230a );
 a80242a <=( A167  and  (not A168) );
 a80243a <=( (not A169)  and  a80242a );
 a80246a <=( A199  and  A166 );
 a80249a <=( A201  and  (not A200) );
 a80250a <=( a80249a  and  a80246a );
 a80251a <=( a80250a  and  a80243a );
 a80255a <=( (not A233)  and  (not A232) );
 a80256a <=( A202  and  a80255a );
 a80259a <=( A266  and  A265 );
 a80262a <=( (not A299)  and  (not A298) );
 a80263a <=( a80262a  and  a80259a );
 a80264a <=( a80263a  and  a80256a );
 a80268a <=( A167  and  (not A168) );
 a80269a <=( (not A169)  and  a80268a );
 a80272a <=( A199  and  A166 );
 a80275a <=( A201  and  (not A200) );
 a80276a <=( a80275a  and  a80272a );
 a80277a <=( a80276a  and  a80269a );
 a80281a <=( (not A233)  and  (not A232) );
 a80282a <=( A202  and  a80281a );
 a80285a <=( (not A267)  and  (not A266) );
 a80288a <=( (not A300)  and  A298 );
 a80289a <=( a80288a  and  a80285a );
 a80290a <=( a80289a  and  a80282a );
 a80294a <=( A167  and  (not A168) );
 a80295a <=( (not A169)  and  a80294a );
 a80298a <=( A199  and  A166 );
 a80301a <=( A201  and  (not A200) );
 a80302a <=( a80301a  and  a80298a );
 a80303a <=( a80302a  and  a80295a );
 a80307a <=( (not A233)  and  (not A232) );
 a80308a <=( A202  and  a80307a );
 a80311a <=( (not A267)  and  (not A266) );
 a80314a <=( A299  and  A298 );
 a80315a <=( a80314a  and  a80311a );
 a80316a <=( a80315a  and  a80308a );
 a80320a <=( A167  and  (not A168) );
 a80321a <=( (not A169)  and  a80320a );
 a80324a <=( A199  and  A166 );
 a80327a <=( A201  and  (not A200) );
 a80328a <=( a80327a  and  a80324a );
 a80329a <=( a80328a  and  a80321a );
 a80333a <=( (not A233)  and  (not A232) );
 a80334a <=( A202  and  a80333a );
 a80337a <=( (not A267)  and  (not A266) );
 a80340a <=( (not A299)  and  (not A298) );
 a80341a <=( a80340a  and  a80337a );
 a80342a <=( a80341a  and  a80334a );
 a80346a <=( A167  and  (not A168) );
 a80347a <=( (not A169)  and  a80346a );
 a80350a <=( A199  and  A166 );
 a80353a <=( A201  and  (not A200) );
 a80354a <=( a80353a  and  a80350a );
 a80355a <=( a80354a  and  a80347a );
 a80359a <=( (not A233)  and  (not A232) );
 a80360a <=( A202  and  a80359a );
 a80363a <=( (not A266)  and  (not A265) );
 a80366a <=( (not A300)  and  A298 );
 a80367a <=( a80366a  and  a80363a );
 a80368a <=( a80367a  and  a80360a );
 a80372a <=( A167  and  (not A168) );
 a80373a <=( (not A169)  and  a80372a );
 a80376a <=( A199  and  A166 );
 a80379a <=( A201  and  (not A200) );
 a80380a <=( a80379a  and  a80376a );
 a80381a <=( a80380a  and  a80373a );
 a80385a <=( (not A233)  and  (not A232) );
 a80386a <=( A202  and  a80385a );
 a80389a <=( (not A266)  and  (not A265) );
 a80392a <=( A299  and  A298 );
 a80393a <=( a80392a  and  a80389a );
 a80394a <=( a80393a  and  a80386a );
 a80398a <=( A167  and  (not A168) );
 a80399a <=( (not A169)  and  a80398a );
 a80402a <=( A199  and  A166 );
 a80405a <=( A201  and  (not A200) );
 a80406a <=( a80405a  and  a80402a );
 a80407a <=( a80406a  and  a80399a );
 a80411a <=( (not A233)  and  (not A232) );
 a80412a <=( A202  and  a80411a );
 a80415a <=( (not A266)  and  (not A265) );
 a80418a <=( (not A299)  and  (not A298) );
 a80419a <=( a80418a  and  a80415a );
 a80420a <=( a80419a  and  a80412a );
 a80424a <=( A167  and  (not A168) );
 a80425a <=( (not A169)  and  a80424a );
 a80428a <=( A199  and  A166 );
 a80431a <=( A201  and  (not A200) );
 a80432a <=( a80431a  and  a80428a );
 a80433a <=( a80432a  and  a80425a );
 a80437a <=( A233  and  A232 );
 a80438a <=( A203  and  a80437a );
 a80441a <=( (not A267)  and  A265 );
 a80444a <=( (not A300)  and  (not A299) );
 a80445a <=( a80444a  and  a80441a );
 a80446a <=( a80445a  and  a80438a );
 a80450a <=( A167  and  (not A168) );
 a80451a <=( (not A169)  and  a80450a );
 a80454a <=( A199  and  A166 );
 a80457a <=( A201  and  (not A200) );
 a80458a <=( a80457a  and  a80454a );
 a80459a <=( a80458a  and  a80451a );
 a80463a <=( A233  and  A232 );
 a80464a <=( A203  and  a80463a );
 a80467a <=( (not A267)  and  A265 );
 a80470a <=( A299  and  A298 );
 a80471a <=( a80470a  and  a80467a );
 a80472a <=( a80471a  and  a80464a );
 a80476a <=( A167  and  (not A168) );
 a80477a <=( (not A169)  and  a80476a );
 a80480a <=( A199  and  A166 );
 a80483a <=( A201  and  (not A200) );
 a80484a <=( a80483a  and  a80480a );
 a80485a <=( a80484a  and  a80477a );
 a80489a <=( A233  and  A232 );
 a80490a <=( A203  and  a80489a );
 a80493a <=( (not A267)  and  A265 );
 a80496a <=( (not A299)  and  (not A298) );
 a80497a <=( a80496a  and  a80493a );
 a80498a <=( a80497a  and  a80490a );
 a80502a <=( A167  and  (not A168) );
 a80503a <=( (not A169)  and  a80502a );
 a80506a <=( A199  and  A166 );
 a80509a <=( A201  and  (not A200) );
 a80510a <=( a80509a  and  a80506a );
 a80511a <=( a80510a  and  a80503a );
 a80515a <=( A233  and  A232 );
 a80516a <=( A203  and  a80515a );
 a80519a <=( A266  and  A265 );
 a80522a <=( (not A300)  and  (not A299) );
 a80523a <=( a80522a  and  a80519a );
 a80524a <=( a80523a  and  a80516a );
 a80528a <=( A167  and  (not A168) );
 a80529a <=( (not A169)  and  a80528a );
 a80532a <=( A199  and  A166 );
 a80535a <=( A201  and  (not A200) );
 a80536a <=( a80535a  and  a80532a );
 a80537a <=( a80536a  and  a80529a );
 a80541a <=( A233  and  A232 );
 a80542a <=( A203  and  a80541a );
 a80545a <=( A266  and  A265 );
 a80548a <=( A299  and  A298 );
 a80549a <=( a80548a  and  a80545a );
 a80550a <=( a80549a  and  a80542a );
 a80554a <=( A167  and  (not A168) );
 a80555a <=( (not A169)  and  a80554a );
 a80558a <=( A199  and  A166 );
 a80561a <=( A201  and  (not A200) );
 a80562a <=( a80561a  and  a80558a );
 a80563a <=( a80562a  and  a80555a );
 a80567a <=( A233  and  A232 );
 a80568a <=( A203  and  a80567a );
 a80571a <=( A266  and  A265 );
 a80574a <=( (not A299)  and  (not A298) );
 a80575a <=( a80574a  and  a80571a );
 a80576a <=( a80575a  and  a80568a );
 a80580a <=( A167  and  (not A168) );
 a80581a <=( (not A169)  and  a80580a );
 a80584a <=( A199  and  A166 );
 a80587a <=( A201  and  (not A200) );
 a80588a <=( a80587a  and  a80584a );
 a80589a <=( a80588a  and  a80581a );
 a80593a <=( A233  and  A232 );
 a80594a <=( A203  and  a80593a );
 a80597a <=( (not A266)  and  (not A265) );
 a80600a <=( (not A300)  and  (not A299) );
 a80601a <=( a80600a  and  a80597a );
 a80602a <=( a80601a  and  a80594a );
 a80606a <=( A167  and  (not A168) );
 a80607a <=( (not A169)  and  a80606a );
 a80610a <=( A199  and  A166 );
 a80613a <=( A201  and  (not A200) );
 a80614a <=( a80613a  and  a80610a );
 a80615a <=( a80614a  and  a80607a );
 a80619a <=( A233  and  A232 );
 a80620a <=( A203  and  a80619a );
 a80623a <=( (not A266)  and  (not A265) );
 a80626a <=( A299  and  A298 );
 a80627a <=( a80626a  and  a80623a );
 a80628a <=( a80627a  and  a80620a );
 a80632a <=( A167  and  (not A168) );
 a80633a <=( (not A169)  and  a80632a );
 a80636a <=( A199  and  A166 );
 a80639a <=( A201  and  (not A200) );
 a80640a <=( a80639a  and  a80636a );
 a80641a <=( a80640a  and  a80633a );
 a80645a <=( A233  and  A232 );
 a80646a <=( A203  and  a80645a );
 a80649a <=( (not A266)  and  (not A265) );
 a80652a <=( (not A299)  and  (not A298) );
 a80653a <=( a80652a  and  a80649a );
 a80654a <=( a80653a  and  a80646a );
 a80658a <=( A167  and  (not A168) );
 a80659a <=( (not A169)  and  a80658a );
 a80662a <=( A199  and  A166 );
 a80665a <=( A201  and  (not A200) );
 a80666a <=( a80665a  and  a80662a );
 a80667a <=( a80666a  and  a80659a );
 a80671a <=( A233  and  (not A232) );
 a80672a <=( A203  and  a80671a );
 a80675a <=( (not A299)  and  A298 );
 a80678a <=( A301  and  A300 );
 a80679a <=( a80678a  and  a80675a );
 a80680a <=( a80679a  and  a80672a );
 a80684a <=( A167  and  (not A168) );
 a80685a <=( (not A169)  and  a80684a );
 a80688a <=( A199  and  A166 );
 a80691a <=( A201  and  (not A200) );
 a80692a <=( a80691a  and  a80688a );
 a80693a <=( a80692a  and  a80685a );
 a80697a <=( A233  and  (not A232) );
 a80698a <=( A203  and  a80697a );
 a80701a <=( (not A299)  and  A298 );
 a80704a <=( A302  and  A300 );
 a80705a <=( a80704a  and  a80701a );
 a80706a <=( a80705a  and  a80698a );
 a80710a <=( A167  and  (not A168) );
 a80711a <=( (not A169)  and  a80710a );
 a80714a <=( A199  and  A166 );
 a80717a <=( A201  and  (not A200) );
 a80718a <=( a80717a  and  a80714a );
 a80719a <=( a80718a  and  a80711a );
 a80723a <=( A233  and  (not A232) );
 a80724a <=( A203  and  a80723a );
 a80727a <=( (not A266)  and  A265 );
 a80730a <=( A268  and  A267 );
 a80731a <=( a80730a  and  a80727a );
 a80732a <=( a80731a  and  a80724a );
 a80736a <=( A167  and  (not A168) );
 a80737a <=( (not A169)  and  a80736a );
 a80740a <=( A199  and  A166 );
 a80743a <=( A201  and  (not A200) );
 a80744a <=( a80743a  and  a80740a );
 a80745a <=( a80744a  and  a80737a );
 a80749a <=( A233  and  (not A232) );
 a80750a <=( A203  and  a80749a );
 a80753a <=( (not A266)  and  A265 );
 a80756a <=( A269  and  A267 );
 a80757a <=( a80756a  and  a80753a );
 a80758a <=( a80757a  and  a80750a );
 a80762a <=( A167  and  (not A168) );
 a80763a <=( (not A169)  and  a80762a );
 a80766a <=( A199  and  A166 );
 a80769a <=( A201  and  (not A200) );
 a80770a <=( a80769a  and  a80766a );
 a80771a <=( a80770a  and  a80763a );
 a80775a <=( (not A234)  and  (not A233) );
 a80776a <=( A203  and  a80775a );
 a80779a <=( A266  and  A265 );
 a80782a <=( (not A300)  and  A298 );
 a80783a <=( a80782a  and  a80779a );
 a80784a <=( a80783a  and  a80776a );
 a80788a <=( A167  and  (not A168) );
 a80789a <=( (not A169)  and  a80788a );
 a80792a <=( A199  and  A166 );
 a80795a <=( A201  and  (not A200) );
 a80796a <=( a80795a  and  a80792a );
 a80797a <=( a80796a  and  a80789a );
 a80801a <=( (not A234)  and  (not A233) );
 a80802a <=( A203  and  a80801a );
 a80805a <=( A266  and  A265 );
 a80808a <=( A299  and  A298 );
 a80809a <=( a80808a  and  a80805a );
 a80810a <=( a80809a  and  a80802a );
 a80814a <=( A167  and  (not A168) );
 a80815a <=( (not A169)  and  a80814a );
 a80818a <=( A199  and  A166 );
 a80821a <=( A201  and  (not A200) );
 a80822a <=( a80821a  and  a80818a );
 a80823a <=( a80822a  and  a80815a );
 a80827a <=( (not A234)  and  (not A233) );
 a80828a <=( A203  and  a80827a );
 a80831a <=( A266  and  A265 );
 a80834a <=( (not A299)  and  (not A298) );
 a80835a <=( a80834a  and  a80831a );
 a80836a <=( a80835a  and  a80828a );
 a80840a <=( A167  and  (not A168) );
 a80841a <=( (not A169)  and  a80840a );
 a80844a <=( A199  and  A166 );
 a80847a <=( A201  and  (not A200) );
 a80848a <=( a80847a  and  a80844a );
 a80849a <=( a80848a  and  a80841a );
 a80853a <=( (not A234)  and  (not A233) );
 a80854a <=( A203  and  a80853a );
 a80857a <=( (not A267)  and  (not A266) );
 a80860a <=( (not A300)  and  A298 );
 a80861a <=( a80860a  and  a80857a );
 a80862a <=( a80861a  and  a80854a );
 a80866a <=( A167  and  (not A168) );
 a80867a <=( (not A169)  and  a80866a );
 a80870a <=( A199  and  A166 );
 a80873a <=( A201  and  (not A200) );
 a80874a <=( a80873a  and  a80870a );
 a80875a <=( a80874a  and  a80867a );
 a80879a <=( (not A234)  and  (not A233) );
 a80880a <=( A203  and  a80879a );
 a80883a <=( (not A267)  and  (not A266) );
 a80886a <=( A299  and  A298 );
 a80887a <=( a80886a  and  a80883a );
 a80888a <=( a80887a  and  a80880a );
 a80892a <=( A167  and  (not A168) );
 a80893a <=( (not A169)  and  a80892a );
 a80896a <=( A199  and  A166 );
 a80899a <=( A201  and  (not A200) );
 a80900a <=( a80899a  and  a80896a );
 a80901a <=( a80900a  and  a80893a );
 a80905a <=( (not A234)  and  (not A233) );
 a80906a <=( A203  and  a80905a );
 a80909a <=( (not A267)  and  (not A266) );
 a80912a <=( (not A299)  and  (not A298) );
 a80913a <=( a80912a  and  a80909a );
 a80914a <=( a80913a  and  a80906a );
 a80918a <=( A167  and  (not A168) );
 a80919a <=( (not A169)  and  a80918a );
 a80922a <=( A199  and  A166 );
 a80925a <=( A201  and  (not A200) );
 a80926a <=( a80925a  and  a80922a );
 a80927a <=( a80926a  and  a80919a );
 a80931a <=( (not A234)  and  (not A233) );
 a80932a <=( A203  and  a80931a );
 a80935a <=( (not A266)  and  (not A265) );
 a80938a <=( (not A300)  and  A298 );
 a80939a <=( a80938a  and  a80935a );
 a80940a <=( a80939a  and  a80932a );
 a80944a <=( A167  and  (not A168) );
 a80945a <=( (not A169)  and  a80944a );
 a80948a <=( A199  and  A166 );
 a80951a <=( A201  and  (not A200) );
 a80952a <=( a80951a  and  a80948a );
 a80953a <=( a80952a  and  a80945a );
 a80957a <=( (not A234)  and  (not A233) );
 a80958a <=( A203  and  a80957a );
 a80961a <=( (not A266)  and  (not A265) );
 a80964a <=( A299  and  A298 );
 a80965a <=( a80964a  and  a80961a );
 a80966a <=( a80965a  and  a80958a );
 a80970a <=( A167  and  (not A168) );
 a80971a <=( (not A169)  and  a80970a );
 a80974a <=( A199  and  A166 );
 a80977a <=( A201  and  (not A200) );
 a80978a <=( a80977a  and  a80974a );
 a80979a <=( a80978a  and  a80971a );
 a80983a <=( (not A234)  and  (not A233) );
 a80984a <=( A203  and  a80983a );
 a80987a <=( (not A266)  and  (not A265) );
 a80990a <=( (not A299)  and  (not A298) );
 a80991a <=( a80990a  and  a80987a );
 a80992a <=( a80991a  and  a80984a );
 a80996a <=( A167  and  (not A168) );
 a80997a <=( (not A169)  and  a80996a );
 a81000a <=( A199  and  A166 );
 a81003a <=( A201  and  (not A200) );
 a81004a <=( a81003a  and  a81000a );
 a81005a <=( a81004a  and  a80997a );
 a81009a <=( (not A233)  and  A232 );
 a81010a <=( A203  and  a81009a );
 a81013a <=( A235  and  A234 );
 a81016a <=( A299  and  (not A298) );
 a81017a <=( a81016a  and  a81013a );
 a81018a <=( a81017a  and  a81010a );
 a81022a <=( A167  and  (not A168) );
 a81023a <=( (not A169)  and  a81022a );
 a81026a <=( A199  and  A166 );
 a81029a <=( A201  and  (not A200) );
 a81030a <=( a81029a  and  a81026a );
 a81031a <=( a81030a  and  a81023a );
 a81035a <=( (not A233)  and  A232 );
 a81036a <=( A203  and  a81035a );
 a81039a <=( A235  and  A234 );
 a81042a <=( A266  and  (not A265) );
 a81043a <=( a81042a  and  a81039a );
 a81044a <=( a81043a  and  a81036a );
 a81048a <=( A167  and  (not A168) );
 a81049a <=( (not A169)  and  a81048a );
 a81052a <=( A199  and  A166 );
 a81055a <=( A201  and  (not A200) );
 a81056a <=( a81055a  and  a81052a );
 a81057a <=( a81056a  and  a81049a );
 a81061a <=( (not A233)  and  A232 );
 a81062a <=( A203  and  a81061a );
 a81065a <=( A236  and  A234 );
 a81068a <=( A299  and  (not A298) );
 a81069a <=( a81068a  and  a81065a );
 a81070a <=( a81069a  and  a81062a );
 a81074a <=( A167  and  (not A168) );
 a81075a <=( (not A169)  and  a81074a );
 a81078a <=( A199  and  A166 );
 a81081a <=( A201  and  (not A200) );
 a81082a <=( a81081a  and  a81078a );
 a81083a <=( a81082a  and  a81075a );
 a81087a <=( (not A233)  and  A232 );
 a81088a <=( A203  and  a81087a );
 a81091a <=( A236  and  A234 );
 a81094a <=( A266  and  (not A265) );
 a81095a <=( a81094a  and  a81091a );
 a81096a <=( a81095a  and  a81088a );
 a81100a <=( A167  and  (not A168) );
 a81101a <=( (not A169)  and  a81100a );
 a81104a <=( A199  and  A166 );
 a81107a <=( A201  and  (not A200) );
 a81108a <=( a81107a  and  a81104a );
 a81109a <=( a81108a  and  a81101a );
 a81113a <=( (not A233)  and  (not A232) );
 a81114a <=( A203  and  a81113a );
 a81117a <=( A266  and  A265 );
 a81120a <=( (not A300)  and  A298 );
 a81121a <=( a81120a  and  a81117a );
 a81122a <=( a81121a  and  a81114a );
 a81126a <=( A167  and  (not A168) );
 a81127a <=( (not A169)  and  a81126a );
 a81130a <=( A199  and  A166 );
 a81133a <=( A201  and  (not A200) );
 a81134a <=( a81133a  and  a81130a );
 a81135a <=( a81134a  and  a81127a );
 a81139a <=( (not A233)  and  (not A232) );
 a81140a <=( A203  and  a81139a );
 a81143a <=( A266  and  A265 );
 a81146a <=( A299  and  A298 );
 a81147a <=( a81146a  and  a81143a );
 a81148a <=( a81147a  and  a81140a );
 a81152a <=( A167  and  (not A168) );
 a81153a <=( (not A169)  and  a81152a );
 a81156a <=( A199  and  A166 );
 a81159a <=( A201  and  (not A200) );
 a81160a <=( a81159a  and  a81156a );
 a81161a <=( a81160a  and  a81153a );
 a81165a <=( (not A233)  and  (not A232) );
 a81166a <=( A203  and  a81165a );
 a81169a <=( A266  and  A265 );
 a81172a <=( (not A299)  and  (not A298) );
 a81173a <=( a81172a  and  a81169a );
 a81174a <=( a81173a  and  a81166a );
 a81178a <=( A167  and  (not A168) );
 a81179a <=( (not A169)  and  a81178a );
 a81182a <=( A199  and  A166 );
 a81185a <=( A201  and  (not A200) );
 a81186a <=( a81185a  and  a81182a );
 a81187a <=( a81186a  and  a81179a );
 a81191a <=( (not A233)  and  (not A232) );
 a81192a <=( A203  and  a81191a );
 a81195a <=( (not A267)  and  (not A266) );
 a81198a <=( (not A300)  and  A298 );
 a81199a <=( a81198a  and  a81195a );
 a81200a <=( a81199a  and  a81192a );
 a81204a <=( A167  and  (not A168) );
 a81205a <=( (not A169)  and  a81204a );
 a81208a <=( A199  and  A166 );
 a81211a <=( A201  and  (not A200) );
 a81212a <=( a81211a  and  a81208a );
 a81213a <=( a81212a  and  a81205a );
 a81217a <=( (not A233)  and  (not A232) );
 a81218a <=( A203  and  a81217a );
 a81221a <=( (not A267)  and  (not A266) );
 a81224a <=( A299  and  A298 );
 a81225a <=( a81224a  and  a81221a );
 a81226a <=( a81225a  and  a81218a );
 a81230a <=( A167  and  (not A168) );
 a81231a <=( (not A169)  and  a81230a );
 a81234a <=( A199  and  A166 );
 a81237a <=( A201  and  (not A200) );
 a81238a <=( a81237a  and  a81234a );
 a81239a <=( a81238a  and  a81231a );
 a81243a <=( (not A233)  and  (not A232) );
 a81244a <=( A203  and  a81243a );
 a81247a <=( (not A267)  and  (not A266) );
 a81250a <=( (not A299)  and  (not A298) );
 a81251a <=( a81250a  and  a81247a );
 a81252a <=( a81251a  and  a81244a );
 a81256a <=( A167  and  (not A168) );
 a81257a <=( (not A169)  and  a81256a );
 a81260a <=( A199  and  A166 );
 a81263a <=( A201  and  (not A200) );
 a81264a <=( a81263a  and  a81260a );
 a81265a <=( a81264a  and  a81257a );
 a81269a <=( (not A233)  and  (not A232) );
 a81270a <=( A203  and  a81269a );
 a81273a <=( (not A266)  and  (not A265) );
 a81276a <=( (not A300)  and  A298 );
 a81277a <=( a81276a  and  a81273a );
 a81278a <=( a81277a  and  a81270a );
 a81282a <=( A167  and  (not A168) );
 a81283a <=( (not A169)  and  a81282a );
 a81286a <=( A199  and  A166 );
 a81289a <=( A201  and  (not A200) );
 a81290a <=( a81289a  and  a81286a );
 a81291a <=( a81290a  and  a81283a );
 a81295a <=( (not A233)  and  (not A232) );
 a81296a <=( A203  and  a81295a );
 a81299a <=( (not A266)  and  (not A265) );
 a81302a <=( A299  and  A298 );
 a81303a <=( a81302a  and  a81299a );
 a81304a <=( a81303a  and  a81296a );
 a81308a <=( A167  and  (not A168) );
 a81309a <=( (not A169)  and  a81308a );
 a81312a <=( A199  and  A166 );
 a81315a <=( A201  and  (not A200) );
 a81316a <=( a81315a  and  a81312a );
 a81317a <=( a81316a  and  a81309a );
 a81321a <=( (not A233)  and  (not A232) );
 a81322a <=( A203  and  a81321a );
 a81325a <=( (not A266)  and  (not A265) );
 a81328a <=( (not A299)  and  (not A298) );
 a81329a <=( a81328a  and  a81325a );
 a81330a <=( a81329a  and  a81322a );
 a81334a <=( A167  and  (not A169) );
 a81335a <=( A170  and  a81334a );
 a81338a <=( A199  and  (not A166) );
 a81341a <=( A232  and  A200 );
 a81342a <=( a81341a  and  a81338a );
 a81343a <=( a81342a  and  a81335a );
 a81347a <=( (not A268)  and  A265 );
 a81348a <=( A233  and  a81347a );
 a81351a <=( (not A299)  and  (not A269) );
 a81354a <=( (not A302)  and  (not A301) );
 a81355a <=( a81354a  and  a81351a );
 a81356a <=( a81355a  and  a81348a );
 a81360a <=( A167  and  (not A169) );
 a81361a <=( A170  and  a81360a );
 a81364a <=( A199  and  (not A166) );
 a81367a <=( (not A233)  and  A200 );
 a81368a <=( a81367a  and  a81364a );
 a81369a <=( a81368a  and  a81361a );
 a81373a <=( A265  and  (not A236) );
 a81374a <=( (not A235)  and  a81373a );
 a81377a <=( A298  and  A266 );
 a81380a <=( (not A302)  and  (not A301) );
 a81381a <=( a81380a  and  a81377a );
 a81382a <=( a81381a  and  a81374a );
 a81386a <=( A167  and  (not A169) );
 a81387a <=( A170  and  a81386a );
 a81390a <=( A199  and  (not A166) );
 a81393a <=( (not A233)  and  A200 );
 a81394a <=( a81393a  and  a81390a );
 a81395a <=( a81394a  and  a81387a );
 a81399a <=( (not A266)  and  (not A236) );
 a81400a <=( (not A235)  and  a81399a );
 a81403a <=( (not A269)  and  (not A268) );
 a81406a <=( (not A300)  and  A298 );
 a81407a <=( a81406a  and  a81403a );
 a81408a <=( a81407a  and  a81400a );
 a81412a <=( A167  and  (not A169) );
 a81413a <=( A170  and  a81412a );
 a81416a <=( A199  and  (not A166) );
 a81419a <=( (not A233)  and  A200 );
 a81420a <=( a81419a  and  a81416a );
 a81421a <=( a81420a  and  a81413a );
 a81425a <=( (not A266)  and  (not A236) );
 a81426a <=( (not A235)  and  a81425a );
 a81429a <=( (not A269)  and  (not A268) );
 a81432a <=( A299  and  A298 );
 a81433a <=( a81432a  and  a81429a );
 a81434a <=( a81433a  and  a81426a );
 a81438a <=( A167  and  (not A169) );
 a81439a <=( A170  and  a81438a );
 a81442a <=( A199  and  (not A166) );
 a81445a <=( (not A233)  and  A200 );
 a81446a <=( a81445a  and  a81442a );
 a81447a <=( a81446a  and  a81439a );
 a81451a <=( (not A266)  and  (not A236) );
 a81452a <=( (not A235)  and  a81451a );
 a81455a <=( (not A269)  and  (not A268) );
 a81458a <=( (not A299)  and  (not A298) );
 a81459a <=( a81458a  and  a81455a );
 a81460a <=( a81459a  and  a81452a );
 a81464a <=( A167  and  (not A169) );
 a81465a <=( A170  and  a81464a );
 a81468a <=( A199  and  (not A166) );
 a81471a <=( (not A233)  and  A200 );
 a81472a <=( a81471a  and  a81468a );
 a81473a <=( a81472a  and  a81465a );
 a81477a <=( (not A266)  and  (not A236) );
 a81478a <=( (not A235)  and  a81477a );
 a81481a <=( A298  and  (not A267) );
 a81484a <=( (not A302)  and  (not A301) );
 a81485a <=( a81484a  and  a81481a );
 a81486a <=( a81485a  and  a81478a );
 a81490a <=( A167  and  (not A169) );
 a81491a <=( A170  and  a81490a );
 a81494a <=( A199  and  (not A166) );
 a81497a <=( (not A233)  and  A200 );
 a81498a <=( a81497a  and  a81494a );
 a81499a <=( a81498a  and  a81491a );
 a81503a <=( (not A265)  and  (not A236) );
 a81504a <=( (not A235)  and  a81503a );
 a81507a <=( A298  and  (not A266) );
 a81510a <=( (not A302)  and  (not A301) );
 a81511a <=( a81510a  and  a81507a );
 a81512a <=( a81511a  and  a81504a );
 a81516a <=( A167  and  (not A169) );
 a81517a <=( A170  and  a81516a );
 a81520a <=( A199  and  (not A166) );
 a81523a <=( (not A233)  and  A200 );
 a81524a <=( a81523a  and  a81520a );
 a81525a <=( a81524a  and  a81517a );
 a81529a <=( (not A268)  and  (not A266) );
 a81530a <=( (not A234)  and  a81529a );
 a81533a <=( A298  and  (not A269) );
 a81536a <=( (not A302)  and  (not A301) );
 a81537a <=( a81536a  and  a81533a );
 a81538a <=( a81537a  and  a81530a );
 a81542a <=( A167  and  (not A169) );
 a81543a <=( A170  and  a81542a );
 a81546a <=( A199  and  (not A166) );
 a81549a <=( A232  and  A200 );
 a81550a <=( a81549a  and  a81546a );
 a81551a <=( a81550a  and  a81543a );
 a81555a <=( A235  and  A234 );
 a81556a <=( (not A233)  and  a81555a );
 a81559a <=( (not A299)  and  A298 );
 a81562a <=( A301  and  A300 );
 a81563a <=( a81562a  and  a81559a );
 a81564a <=( a81563a  and  a81556a );
 a81568a <=( A167  and  (not A169) );
 a81569a <=( A170  and  a81568a );
 a81572a <=( A199  and  (not A166) );
 a81575a <=( A232  and  A200 );
 a81576a <=( a81575a  and  a81572a );
 a81577a <=( a81576a  and  a81569a );
 a81581a <=( A235  and  A234 );
 a81582a <=( (not A233)  and  a81581a );
 a81585a <=( (not A299)  and  A298 );
 a81588a <=( A302  and  A300 );
 a81589a <=( a81588a  and  a81585a );
 a81590a <=( a81589a  and  a81582a );
 a81594a <=( A167  and  (not A169) );
 a81595a <=( A170  and  a81594a );
 a81598a <=( A199  and  (not A166) );
 a81601a <=( A232  and  A200 );
 a81602a <=( a81601a  and  a81598a );
 a81603a <=( a81602a  and  a81595a );
 a81607a <=( A235  and  A234 );
 a81608a <=( (not A233)  and  a81607a );
 a81611a <=( (not A266)  and  A265 );
 a81614a <=( A268  and  A267 );
 a81615a <=( a81614a  and  a81611a );
 a81616a <=( a81615a  and  a81608a );
 a81620a <=( A167  and  (not A169) );
 a81621a <=( A170  and  a81620a );
 a81624a <=( A199  and  (not A166) );
 a81627a <=( A232  and  A200 );
 a81628a <=( a81627a  and  a81624a );
 a81629a <=( a81628a  and  a81621a );
 a81633a <=( A235  and  A234 );
 a81634a <=( (not A233)  and  a81633a );
 a81637a <=( (not A266)  and  A265 );
 a81640a <=( A269  and  A267 );
 a81641a <=( a81640a  and  a81637a );
 a81642a <=( a81641a  and  a81634a );
 a81646a <=( A167  and  (not A169) );
 a81647a <=( A170  and  a81646a );
 a81650a <=( A199  and  (not A166) );
 a81653a <=( A232  and  A200 );
 a81654a <=( a81653a  and  a81650a );
 a81655a <=( a81654a  and  a81647a );
 a81659a <=( A236  and  A234 );
 a81660a <=( (not A233)  and  a81659a );
 a81663a <=( (not A299)  and  A298 );
 a81666a <=( A301  and  A300 );
 a81667a <=( a81666a  and  a81663a );
 a81668a <=( a81667a  and  a81660a );
 a81672a <=( A167  and  (not A169) );
 a81673a <=( A170  and  a81672a );
 a81676a <=( A199  and  (not A166) );
 a81679a <=( A232  and  A200 );
 a81680a <=( a81679a  and  a81676a );
 a81681a <=( a81680a  and  a81673a );
 a81685a <=( A236  and  A234 );
 a81686a <=( (not A233)  and  a81685a );
 a81689a <=( (not A299)  and  A298 );
 a81692a <=( A302  and  A300 );
 a81693a <=( a81692a  and  a81689a );
 a81694a <=( a81693a  and  a81686a );
 a81698a <=( A167  and  (not A169) );
 a81699a <=( A170  and  a81698a );
 a81702a <=( A199  and  (not A166) );
 a81705a <=( A232  and  A200 );
 a81706a <=( a81705a  and  a81702a );
 a81707a <=( a81706a  and  a81699a );
 a81711a <=( A236  and  A234 );
 a81712a <=( (not A233)  and  a81711a );
 a81715a <=( (not A266)  and  A265 );
 a81718a <=( A268  and  A267 );
 a81719a <=( a81718a  and  a81715a );
 a81720a <=( a81719a  and  a81712a );
 a81724a <=( A167  and  (not A169) );
 a81725a <=( A170  and  a81724a );
 a81728a <=( A199  and  (not A166) );
 a81731a <=( A232  and  A200 );
 a81732a <=( a81731a  and  a81728a );
 a81733a <=( a81732a  and  a81725a );
 a81737a <=( A236  and  A234 );
 a81738a <=( (not A233)  and  a81737a );
 a81741a <=( (not A266)  and  A265 );
 a81744a <=( A269  and  A267 );
 a81745a <=( a81744a  and  a81741a );
 a81746a <=( a81745a  and  a81738a );
 a81750a <=( A167  and  (not A169) );
 a81751a <=( A170  and  a81750a );
 a81754a <=( A199  and  (not A166) );
 a81757a <=( (not A232)  and  A200 );
 a81758a <=( a81757a  and  a81754a );
 a81759a <=( a81758a  and  a81751a );
 a81763a <=( (not A268)  and  (not A266) );
 a81764a <=( (not A233)  and  a81763a );
 a81767a <=( A298  and  (not A269) );
 a81770a <=( (not A302)  and  (not A301) );
 a81771a <=( a81770a  and  a81767a );
 a81772a <=( a81771a  and  a81764a );
 a81776a <=( A167  and  (not A169) );
 a81777a <=( A170  and  a81776a );
 a81780a <=( (not A200)  and  (not A166) );
 a81783a <=( (not A203)  and  (not A202) );
 a81784a <=( a81783a  and  a81780a );
 a81785a <=( a81784a  and  a81777a );
 a81789a <=( A265  and  A233 );
 a81790a <=( A232  and  a81789a );
 a81793a <=( (not A269)  and  (not A268) );
 a81796a <=( (not A300)  and  (not A299) );
 a81797a <=( a81796a  and  a81793a );
 a81798a <=( a81797a  and  a81790a );
 a81802a <=( A167  and  (not A169) );
 a81803a <=( A170  and  a81802a );
 a81806a <=( (not A200)  and  (not A166) );
 a81809a <=( (not A203)  and  (not A202) );
 a81810a <=( a81809a  and  a81806a );
 a81811a <=( a81810a  and  a81803a );
 a81815a <=( A265  and  A233 );
 a81816a <=( A232  and  a81815a );
 a81819a <=( (not A269)  and  (not A268) );
 a81822a <=( A299  and  A298 );
 a81823a <=( a81822a  and  a81819a );
 a81824a <=( a81823a  and  a81816a );
 a81828a <=( A167  and  (not A169) );
 a81829a <=( A170  and  a81828a );
 a81832a <=( (not A200)  and  (not A166) );
 a81835a <=( (not A203)  and  (not A202) );
 a81836a <=( a81835a  and  a81832a );
 a81837a <=( a81836a  and  a81829a );
 a81841a <=( A265  and  A233 );
 a81842a <=( A232  and  a81841a );
 a81845a <=( (not A269)  and  (not A268) );
 a81848a <=( (not A299)  and  (not A298) );
 a81849a <=( a81848a  and  a81845a );
 a81850a <=( a81849a  and  a81842a );
 a81854a <=( A167  and  (not A169) );
 a81855a <=( A170  and  a81854a );
 a81858a <=( (not A200)  and  (not A166) );
 a81861a <=( (not A203)  and  (not A202) );
 a81862a <=( a81861a  and  a81858a );
 a81863a <=( a81862a  and  a81855a );
 a81867a <=( A265  and  A233 );
 a81868a <=( A232  and  a81867a );
 a81871a <=( (not A299)  and  (not A267) );
 a81874a <=( (not A302)  and  (not A301) );
 a81875a <=( a81874a  and  a81871a );
 a81876a <=( a81875a  and  a81868a );
 a81880a <=( A167  and  (not A169) );
 a81881a <=( A170  and  a81880a );
 a81884a <=( (not A200)  and  (not A166) );
 a81887a <=( (not A203)  and  (not A202) );
 a81888a <=( a81887a  and  a81884a );
 a81889a <=( a81888a  and  a81881a );
 a81893a <=( A265  and  A233 );
 a81894a <=( A232  and  a81893a );
 a81897a <=( (not A299)  and  A266 );
 a81900a <=( (not A302)  and  (not A301) );
 a81901a <=( a81900a  and  a81897a );
 a81902a <=( a81901a  and  a81894a );
 a81906a <=( A167  and  (not A169) );
 a81907a <=( A170  and  a81906a );
 a81910a <=( (not A200)  and  (not A166) );
 a81913a <=( (not A203)  and  (not A202) );
 a81914a <=( a81913a  and  a81910a );
 a81915a <=( a81914a  and  a81907a );
 a81919a <=( (not A265)  and  A233 );
 a81920a <=( A232  and  a81919a );
 a81923a <=( (not A299)  and  (not A266) );
 a81926a <=( (not A302)  and  (not A301) );
 a81927a <=( a81926a  and  a81923a );
 a81928a <=( a81927a  and  a81920a );
 a81932a <=( A167  and  (not A169) );
 a81933a <=( A170  and  a81932a );
 a81936a <=( (not A200)  and  (not A166) );
 a81939a <=( (not A203)  and  (not A202) );
 a81940a <=( a81939a  and  a81936a );
 a81941a <=( a81940a  and  a81933a );
 a81945a <=( (not A236)  and  (not A235) );
 a81946a <=( (not A233)  and  a81945a );
 a81949a <=( A266  and  A265 );
 a81952a <=( (not A300)  and  A298 );
 a81953a <=( a81952a  and  a81949a );
 a81954a <=( a81953a  and  a81946a );
 a81958a <=( A167  and  (not A169) );
 a81959a <=( A170  and  a81958a );
 a81962a <=( (not A200)  and  (not A166) );
 a81965a <=( (not A203)  and  (not A202) );
 a81966a <=( a81965a  and  a81962a );
 a81967a <=( a81966a  and  a81959a );
 a81971a <=( (not A236)  and  (not A235) );
 a81972a <=( (not A233)  and  a81971a );
 a81975a <=( A266  and  A265 );
 a81978a <=( A299  and  A298 );
 a81979a <=( a81978a  and  a81975a );
 a81980a <=( a81979a  and  a81972a );
 a81984a <=( A167  and  (not A169) );
 a81985a <=( A170  and  a81984a );
 a81988a <=( (not A200)  and  (not A166) );
 a81991a <=( (not A203)  and  (not A202) );
 a81992a <=( a81991a  and  a81988a );
 a81993a <=( a81992a  and  a81985a );
 a81997a <=( (not A236)  and  (not A235) );
 a81998a <=( (not A233)  and  a81997a );
 a82001a <=( A266  and  A265 );
 a82004a <=( (not A299)  and  (not A298) );
 a82005a <=( a82004a  and  a82001a );
 a82006a <=( a82005a  and  a81998a );
 a82010a <=( A167  and  (not A169) );
 a82011a <=( A170  and  a82010a );
 a82014a <=( (not A200)  and  (not A166) );
 a82017a <=( (not A203)  and  (not A202) );
 a82018a <=( a82017a  and  a82014a );
 a82019a <=( a82018a  and  a82011a );
 a82023a <=( (not A236)  and  (not A235) );
 a82024a <=( (not A233)  and  a82023a );
 a82027a <=( (not A267)  and  (not A266) );
 a82030a <=( (not A300)  and  A298 );
 a82031a <=( a82030a  and  a82027a );
 a82032a <=( a82031a  and  a82024a );
 a82036a <=( A167  and  (not A169) );
 a82037a <=( A170  and  a82036a );
 a82040a <=( (not A200)  and  (not A166) );
 a82043a <=( (not A203)  and  (not A202) );
 a82044a <=( a82043a  and  a82040a );
 a82045a <=( a82044a  and  a82037a );
 a82049a <=( (not A236)  and  (not A235) );
 a82050a <=( (not A233)  and  a82049a );
 a82053a <=( (not A267)  and  (not A266) );
 a82056a <=( A299  and  A298 );
 a82057a <=( a82056a  and  a82053a );
 a82058a <=( a82057a  and  a82050a );
 a82062a <=( A167  and  (not A169) );
 a82063a <=( A170  and  a82062a );
 a82066a <=( (not A200)  and  (not A166) );
 a82069a <=( (not A203)  and  (not A202) );
 a82070a <=( a82069a  and  a82066a );
 a82071a <=( a82070a  and  a82063a );
 a82075a <=( (not A236)  and  (not A235) );
 a82076a <=( (not A233)  and  a82075a );
 a82079a <=( (not A267)  and  (not A266) );
 a82082a <=( (not A299)  and  (not A298) );
 a82083a <=( a82082a  and  a82079a );
 a82084a <=( a82083a  and  a82076a );
 a82088a <=( A167  and  (not A169) );
 a82089a <=( A170  and  a82088a );
 a82092a <=( (not A200)  and  (not A166) );
 a82095a <=( (not A203)  and  (not A202) );
 a82096a <=( a82095a  and  a82092a );
 a82097a <=( a82096a  and  a82089a );
 a82101a <=( (not A236)  and  (not A235) );
 a82102a <=( (not A233)  and  a82101a );
 a82105a <=( (not A266)  and  (not A265) );
 a82108a <=( (not A300)  and  A298 );
 a82109a <=( a82108a  and  a82105a );
 a82110a <=( a82109a  and  a82102a );
 a82114a <=( A167  and  (not A169) );
 a82115a <=( A170  and  a82114a );
 a82118a <=( (not A200)  and  (not A166) );
 a82121a <=( (not A203)  and  (not A202) );
 a82122a <=( a82121a  and  a82118a );
 a82123a <=( a82122a  and  a82115a );
 a82127a <=( (not A236)  and  (not A235) );
 a82128a <=( (not A233)  and  a82127a );
 a82131a <=( (not A266)  and  (not A265) );
 a82134a <=( A299  and  A298 );
 a82135a <=( a82134a  and  a82131a );
 a82136a <=( a82135a  and  a82128a );
 a82140a <=( A167  and  (not A169) );
 a82141a <=( A170  and  a82140a );
 a82144a <=( (not A200)  and  (not A166) );
 a82147a <=( (not A203)  and  (not A202) );
 a82148a <=( a82147a  and  a82144a );
 a82149a <=( a82148a  and  a82141a );
 a82153a <=( (not A236)  and  (not A235) );
 a82154a <=( (not A233)  and  a82153a );
 a82157a <=( (not A266)  and  (not A265) );
 a82160a <=( (not A299)  and  (not A298) );
 a82161a <=( a82160a  and  a82157a );
 a82162a <=( a82161a  and  a82154a );
 a82166a <=( A167  and  (not A169) );
 a82167a <=( A170  and  a82166a );
 a82170a <=( (not A200)  and  (not A166) );
 a82173a <=( (not A203)  and  (not A202) );
 a82174a <=( a82173a  and  a82170a );
 a82175a <=( a82174a  and  a82167a );
 a82179a <=( A265  and  (not A234) );
 a82180a <=( (not A233)  and  a82179a );
 a82183a <=( A298  and  A266 );
 a82186a <=( (not A302)  and  (not A301) );
 a82187a <=( a82186a  and  a82183a );
 a82188a <=( a82187a  and  a82180a );
 a82192a <=( A167  and  (not A169) );
 a82193a <=( A170  and  a82192a );
 a82196a <=( (not A200)  and  (not A166) );
 a82199a <=( (not A203)  and  (not A202) );
 a82200a <=( a82199a  and  a82196a );
 a82201a <=( a82200a  and  a82193a );
 a82205a <=( (not A266)  and  (not A234) );
 a82206a <=( (not A233)  and  a82205a );
 a82209a <=( (not A269)  and  (not A268) );
 a82212a <=( (not A300)  and  A298 );
 a82213a <=( a82212a  and  a82209a );
 a82214a <=( a82213a  and  a82206a );
 a82218a <=( A167  and  (not A169) );
 a82219a <=( A170  and  a82218a );
 a82222a <=( (not A200)  and  (not A166) );
 a82225a <=( (not A203)  and  (not A202) );
 a82226a <=( a82225a  and  a82222a );
 a82227a <=( a82226a  and  a82219a );
 a82231a <=( (not A266)  and  (not A234) );
 a82232a <=( (not A233)  and  a82231a );
 a82235a <=( (not A269)  and  (not A268) );
 a82238a <=( A299  and  A298 );
 a82239a <=( a82238a  and  a82235a );
 a82240a <=( a82239a  and  a82232a );
 a82244a <=( A167  and  (not A169) );
 a82245a <=( A170  and  a82244a );
 a82248a <=( (not A200)  and  (not A166) );
 a82251a <=( (not A203)  and  (not A202) );
 a82252a <=( a82251a  and  a82248a );
 a82253a <=( a82252a  and  a82245a );
 a82257a <=( (not A266)  and  (not A234) );
 a82258a <=( (not A233)  and  a82257a );
 a82261a <=( (not A269)  and  (not A268) );
 a82264a <=( (not A299)  and  (not A298) );
 a82265a <=( a82264a  and  a82261a );
 a82266a <=( a82265a  and  a82258a );
 a82270a <=( A167  and  (not A169) );
 a82271a <=( A170  and  a82270a );
 a82274a <=( (not A200)  and  (not A166) );
 a82277a <=( (not A203)  and  (not A202) );
 a82278a <=( a82277a  and  a82274a );
 a82279a <=( a82278a  and  a82271a );
 a82283a <=( (not A266)  and  (not A234) );
 a82284a <=( (not A233)  and  a82283a );
 a82287a <=( A298  and  (not A267) );
 a82290a <=( (not A302)  and  (not A301) );
 a82291a <=( a82290a  and  a82287a );
 a82292a <=( a82291a  and  a82284a );
 a82296a <=( A167  and  (not A169) );
 a82297a <=( A170  and  a82296a );
 a82300a <=( (not A200)  and  (not A166) );
 a82303a <=( (not A203)  and  (not A202) );
 a82304a <=( a82303a  and  a82300a );
 a82305a <=( a82304a  and  a82297a );
 a82309a <=( (not A265)  and  (not A234) );
 a82310a <=( (not A233)  and  a82309a );
 a82313a <=( A298  and  (not A266) );
 a82316a <=( (not A302)  and  (not A301) );
 a82317a <=( a82316a  and  a82313a );
 a82318a <=( a82317a  and  a82310a );
 a82322a <=( A167  and  (not A169) );
 a82323a <=( A170  and  a82322a );
 a82326a <=( (not A200)  and  (not A166) );
 a82329a <=( (not A203)  and  (not A202) );
 a82330a <=( a82329a  and  a82326a );
 a82331a <=( a82330a  and  a82323a );
 a82335a <=( A265  and  (not A233) );
 a82336a <=( (not A232)  and  a82335a );
 a82339a <=( A298  and  A266 );
 a82342a <=( (not A302)  and  (not A301) );
 a82343a <=( a82342a  and  a82339a );
 a82344a <=( a82343a  and  a82336a );
 a82348a <=( A167  and  (not A169) );
 a82349a <=( A170  and  a82348a );
 a82352a <=( (not A200)  and  (not A166) );
 a82355a <=( (not A203)  and  (not A202) );
 a82356a <=( a82355a  and  a82352a );
 a82357a <=( a82356a  and  a82349a );
 a82361a <=( (not A266)  and  (not A233) );
 a82362a <=( (not A232)  and  a82361a );
 a82365a <=( (not A269)  and  (not A268) );
 a82368a <=( (not A300)  and  A298 );
 a82369a <=( a82368a  and  a82365a );
 a82370a <=( a82369a  and  a82362a );
 a82374a <=( A167  and  (not A169) );
 a82375a <=( A170  and  a82374a );
 a82378a <=( (not A200)  and  (not A166) );
 a82381a <=( (not A203)  and  (not A202) );
 a82382a <=( a82381a  and  a82378a );
 a82383a <=( a82382a  and  a82375a );
 a82387a <=( (not A266)  and  (not A233) );
 a82388a <=( (not A232)  and  a82387a );
 a82391a <=( (not A269)  and  (not A268) );
 a82394a <=( A299  and  A298 );
 a82395a <=( a82394a  and  a82391a );
 a82396a <=( a82395a  and  a82388a );
 a82400a <=( A167  and  (not A169) );
 a82401a <=( A170  and  a82400a );
 a82404a <=( (not A200)  and  (not A166) );
 a82407a <=( (not A203)  and  (not A202) );
 a82408a <=( a82407a  and  a82404a );
 a82409a <=( a82408a  and  a82401a );
 a82413a <=( (not A266)  and  (not A233) );
 a82414a <=( (not A232)  and  a82413a );
 a82417a <=( (not A269)  and  (not A268) );
 a82420a <=( (not A299)  and  (not A298) );
 a82421a <=( a82420a  and  a82417a );
 a82422a <=( a82421a  and  a82414a );
 a82426a <=( A167  and  (not A169) );
 a82427a <=( A170  and  a82426a );
 a82430a <=( (not A200)  and  (not A166) );
 a82433a <=( (not A203)  and  (not A202) );
 a82434a <=( a82433a  and  a82430a );
 a82435a <=( a82434a  and  a82427a );
 a82439a <=( (not A266)  and  (not A233) );
 a82440a <=( (not A232)  and  a82439a );
 a82443a <=( A298  and  (not A267) );
 a82446a <=( (not A302)  and  (not A301) );
 a82447a <=( a82446a  and  a82443a );
 a82448a <=( a82447a  and  a82440a );
 a82452a <=( A167  and  (not A169) );
 a82453a <=( A170  and  a82452a );
 a82456a <=( (not A200)  and  (not A166) );
 a82459a <=( (not A203)  and  (not A202) );
 a82460a <=( a82459a  and  a82456a );
 a82461a <=( a82460a  and  a82453a );
 a82465a <=( (not A265)  and  (not A233) );
 a82466a <=( (not A232)  and  a82465a );
 a82469a <=( A298  and  (not A266) );
 a82472a <=( (not A302)  and  (not A301) );
 a82473a <=( a82472a  and  a82469a );
 a82474a <=( a82473a  and  a82466a );
 a82478a <=( A167  and  (not A169) );
 a82479a <=( A170  and  a82478a );
 a82482a <=( (not A200)  and  (not A166) );
 a82485a <=( A232  and  (not A201) );
 a82486a <=( a82485a  and  a82482a );
 a82487a <=( a82486a  and  a82479a );
 a82491a <=( (not A268)  and  A265 );
 a82492a <=( A233  and  a82491a );
 a82495a <=( (not A299)  and  (not A269) );
 a82498a <=( (not A302)  and  (not A301) );
 a82499a <=( a82498a  and  a82495a );
 a82500a <=( a82499a  and  a82492a );
 a82504a <=( A167  and  (not A169) );
 a82505a <=( A170  and  a82504a );
 a82508a <=( (not A200)  and  (not A166) );
 a82511a <=( (not A233)  and  (not A201) );
 a82512a <=( a82511a  and  a82508a );
 a82513a <=( a82512a  and  a82505a );
 a82517a <=( A265  and  (not A236) );
 a82518a <=( (not A235)  and  a82517a );
 a82521a <=( A298  and  A266 );
 a82524a <=( (not A302)  and  (not A301) );
 a82525a <=( a82524a  and  a82521a );
 a82526a <=( a82525a  and  a82518a );
 a82530a <=( A167  and  (not A169) );
 a82531a <=( A170  and  a82530a );
 a82534a <=( (not A200)  and  (not A166) );
 a82537a <=( (not A233)  and  (not A201) );
 a82538a <=( a82537a  and  a82534a );
 a82539a <=( a82538a  and  a82531a );
 a82543a <=( (not A266)  and  (not A236) );
 a82544a <=( (not A235)  and  a82543a );
 a82547a <=( (not A269)  and  (not A268) );
 a82550a <=( (not A300)  and  A298 );
 a82551a <=( a82550a  and  a82547a );
 a82552a <=( a82551a  and  a82544a );
 a82556a <=( A167  and  (not A169) );
 a82557a <=( A170  and  a82556a );
 a82560a <=( (not A200)  and  (not A166) );
 a82563a <=( (not A233)  and  (not A201) );
 a82564a <=( a82563a  and  a82560a );
 a82565a <=( a82564a  and  a82557a );
 a82569a <=( (not A266)  and  (not A236) );
 a82570a <=( (not A235)  and  a82569a );
 a82573a <=( (not A269)  and  (not A268) );
 a82576a <=( A299  and  A298 );
 a82577a <=( a82576a  and  a82573a );
 a82578a <=( a82577a  and  a82570a );
 a82582a <=( A167  and  (not A169) );
 a82583a <=( A170  and  a82582a );
 a82586a <=( (not A200)  and  (not A166) );
 a82589a <=( (not A233)  and  (not A201) );
 a82590a <=( a82589a  and  a82586a );
 a82591a <=( a82590a  and  a82583a );
 a82595a <=( (not A266)  and  (not A236) );
 a82596a <=( (not A235)  and  a82595a );
 a82599a <=( (not A269)  and  (not A268) );
 a82602a <=( (not A299)  and  (not A298) );
 a82603a <=( a82602a  and  a82599a );
 a82604a <=( a82603a  and  a82596a );
 a82608a <=( A167  and  (not A169) );
 a82609a <=( A170  and  a82608a );
 a82612a <=( (not A200)  and  (not A166) );
 a82615a <=( (not A233)  and  (not A201) );
 a82616a <=( a82615a  and  a82612a );
 a82617a <=( a82616a  and  a82609a );
 a82621a <=( (not A266)  and  (not A236) );
 a82622a <=( (not A235)  and  a82621a );
 a82625a <=( A298  and  (not A267) );
 a82628a <=( (not A302)  and  (not A301) );
 a82629a <=( a82628a  and  a82625a );
 a82630a <=( a82629a  and  a82622a );
 a82634a <=( A167  and  (not A169) );
 a82635a <=( A170  and  a82634a );
 a82638a <=( (not A200)  and  (not A166) );
 a82641a <=( (not A233)  and  (not A201) );
 a82642a <=( a82641a  and  a82638a );
 a82643a <=( a82642a  and  a82635a );
 a82647a <=( (not A265)  and  (not A236) );
 a82648a <=( (not A235)  and  a82647a );
 a82651a <=( A298  and  (not A266) );
 a82654a <=( (not A302)  and  (not A301) );
 a82655a <=( a82654a  and  a82651a );
 a82656a <=( a82655a  and  a82648a );
 a82660a <=( A167  and  (not A169) );
 a82661a <=( A170  and  a82660a );
 a82664a <=( (not A200)  and  (not A166) );
 a82667a <=( (not A233)  and  (not A201) );
 a82668a <=( a82667a  and  a82664a );
 a82669a <=( a82668a  and  a82661a );
 a82673a <=( (not A268)  and  (not A266) );
 a82674a <=( (not A234)  and  a82673a );
 a82677a <=( A298  and  (not A269) );
 a82680a <=( (not A302)  and  (not A301) );
 a82681a <=( a82680a  and  a82677a );
 a82682a <=( a82681a  and  a82674a );
 a82686a <=( A167  and  (not A169) );
 a82687a <=( A170  and  a82686a );
 a82690a <=( (not A200)  and  (not A166) );
 a82693a <=( A232  and  (not A201) );
 a82694a <=( a82693a  and  a82690a );
 a82695a <=( a82694a  and  a82687a );
 a82699a <=( A235  and  A234 );
 a82700a <=( (not A233)  and  a82699a );
 a82703a <=( (not A299)  and  A298 );
 a82706a <=( A301  and  A300 );
 a82707a <=( a82706a  and  a82703a );
 a82708a <=( a82707a  and  a82700a );
 a82712a <=( A167  and  (not A169) );
 a82713a <=( A170  and  a82712a );
 a82716a <=( (not A200)  and  (not A166) );
 a82719a <=( A232  and  (not A201) );
 a82720a <=( a82719a  and  a82716a );
 a82721a <=( a82720a  and  a82713a );
 a82725a <=( A235  and  A234 );
 a82726a <=( (not A233)  and  a82725a );
 a82729a <=( (not A299)  and  A298 );
 a82732a <=( A302  and  A300 );
 a82733a <=( a82732a  and  a82729a );
 a82734a <=( a82733a  and  a82726a );
 a82738a <=( A167  and  (not A169) );
 a82739a <=( A170  and  a82738a );
 a82742a <=( (not A200)  and  (not A166) );
 a82745a <=( A232  and  (not A201) );
 a82746a <=( a82745a  and  a82742a );
 a82747a <=( a82746a  and  a82739a );
 a82751a <=( A235  and  A234 );
 a82752a <=( (not A233)  and  a82751a );
 a82755a <=( (not A266)  and  A265 );
 a82758a <=( A268  and  A267 );
 a82759a <=( a82758a  and  a82755a );
 a82760a <=( a82759a  and  a82752a );
 a82764a <=( A167  and  (not A169) );
 a82765a <=( A170  and  a82764a );
 a82768a <=( (not A200)  and  (not A166) );
 a82771a <=( A232  and  (not A201) );
 a82772a <=( a82771a  and  a82768a );
 a82773a <=( a82772a  and  a82765a );
 a82777a <=( A235  and  A234 );
 a82778a <=( (not A233)  and  a82777a );
 a82781a <=( (not A266)  and  A265 );
 a82784a <=( A269  and  A267 );
 a82785a <=( a82784a  and  a82781a );
 a82786a <=( a82785a  and  a82778a );
 a82790a <=( A167  and  (not A169) );
 a82791a <=( A170  and  a82790a );
 a82794a <=( (not A200)  and  (not A166) );
 a82797a <=( A232  and  (not A201) );
 a82798a <=( a82797a  and  a82794a );
 a82799a <=( a82798a  and  a82791a );
 a82803a <=( A236  and  A234 );
 a82804a <=( (not A233)  and  a82803a );
 a82807a <=( (not A299)  and  A298 );
 a82810a <=( A301  and  A300 );
 a82811a <=( a82810a  and  a82807a );
 a82812a <=( a82811a  and  a82804a );
 a82816a <=( A167  and  (not A169) );
 a82817a <=( A170  and  a82816a );
 a82820a <=( (not A200)  and  (not A166) );
 a82823a <=( A232  and  (not A201) );
 a82824a <=( a82823a  and  a82820a );
 a82825a <=( a82824a  and  a82817a );
 a82829a <=( A236  and  A234 );
 a82830a <=( (not A233)  and  a82829a );
 a82833a <=( (not A299)  and  A298 );
 a82836a <=( A302  and  A300 );
 a82837a <=( a82836a  and  a82833a );
 a82838a <=( a82837a  and  a82830a );
 a82842a <=( A167  and  (not A169) );
 a82843a <=( A170  and  a82842a );
 a82846a <=( (not A200)  and  (not A166) );
 a82849a <=( A232  and  (not A201) );
 a82850a <=( a82849a  and  a82846a );
 a82851a <=( a82850a  and  a82843a );
 a82855a <=( A236  and  A234 );
 a82856a <=( (not A233)  and  a82855a );
 a82859a <=( (not A266)  and  A265 );
 a82862a <=( A268  and  A267 );
 a82863a <=( a82862a  and  a82859a );
 a82864a <=( a82863a  and  a82856a );
 a82868a <=( A167  and  (not A169) );
 a82869a <=( A170  and  a82868a );
 a82872a <=( (not A200)  and  (not A166) );
 a82875a <=( A232  and  (not A201) );
 a82876a <=( a82875a  and  a82872a );
 a82877a <=( a82876a  and  a82869a );
 a82881a <=( A236  and  A234 );
 a82882a <=( (not A233)  and  a82881a );
 a82885a <=( (not A266)  and  A265 );
 a82888a <=( A269  and  A267 );
 a82889a <=( a82888a  and  a82885a );
 a82890a <=( a82889a  and  a82882a );
 a82894a <=( A167  and  (not A169) );
 a82895a <=( A170  and  a82894a );
 a82898a <=( (not A200)  and  (not A166) );
 a82901a <=( (not A232)  and  (not A201) );
 a82902a <=( a82901a  and  a82898a );
 a82903a <=( a82902a  and  a82895a );
 a82907a <=( (not A268)  and  (not A266) );
 a82908a <=( (not A233)  and  a82907a );
 a82911a <=( A298  and  (not A269) );
 a82914a <=( (not A302)  and  (not A301) );
 a82915a <=( a82914a  and  a82911a );
 a82916a <=( a82915a  and  a82908a );
 a82920a <=( A167  and  (not A169) );
 a82921a <=( A170  and  a82920a );
 a82924a <=( (not A199)  and  (not A166) );
 a82927a <=( A232  and  (not A200) );
 a82928a <=( a82927a  and  a82924a );
 a82929a <=( a82928a  and  a82921a );
 a82933a <=( (not A268)  and  A265 );
 a82934a <=( A233  and  a82933a );
 a82937a <=( (not A299)  and  (not A269) );
 a82940a <=( (not A302)  and  (not A301) );
 a82941a <=( a82940a  and  a82937a );
 a82942a <=( a82941a  and  a82934a );
 a82946a <=( A167  and  (not A169) );
 a82947a <=( A170  and  a82946a );
 a82950a <=( (not A199)  and  (not A166) );
 a82953a <=( (not A233)  and  (not A200) );
 a82954a <=( a82953a  and  a82950a );
 a82955a <=( a82954a  and  a82947a );
 a82959a <=( A265  and  (not A236) );
 a82960a <=( (not A235)  and  a82959a );
 a82963a <=( A298  and  A266 );
 a82966a <=( (not A302)  and  (not A301) );
 a82967a <=( a82966a  and  a82963a );
 a82968a <=( a82967a  and  a82960a );
 a82972a <=( A167  and  (not A169) );
 a82973a <=( A170  and  a82972a );
 a82976a <=( (not A199)  and  (not A166) );
 a82979a <=( (not A233)  and  (not A200) );
 a82980a <=( a82979a  and  a82976a );
 a82981a <=( a82980a  and  a82973a );
 a82985a <=( (not A266)  and  (not A236) );
 a82986a <=( (not A235)  and  a82985a );
 a82989a <=( (not A269)  and  (not A268) );
 a82992a <=( (not A300)  and  A298 );
 a82993a <=( a82992a  and  a82989a );
 a82994a <=( a82993a  and  a82986a );
 a82998a <=( A167  and  (not A169) );
 a82999a <=( A170  and  a82998a );
 a83002a <=( (not A199)  and  (not A166) );
 a83005a <=( (not A233)  and  (not A200) );
 a83006a <=( a83005a  and  a83002a );
 a83007a <=( a83006a  and  a82999a );
 a83011a <=( (not A266)  and  (not A236) );
 a83012a <=( (not A235)  and  a83011a );
 a83015a <=( (not A269)  and  (not A268) );
 a83018a <=( A299  and  A298 );
 a83019a <=( a83018a  and  a83015a );
 a83020a <=( a83019a  and  a83012a );
 a83024a <=( A167  and  (not A169) );
 a83025a <=( A170  and  a83024a );
 a83028a <=( (not A199)  and  (not A166) );
 a83031a <=( (not A233)  and  (not A200) );
 a83032a <=( a83031a  and  a83028a );
 a83033a <=( a83032a  and  a83025a );
 a83037a <=( (not A266)  and  (not A236) );
 a83038a <=( (not A235)  and  a83037a );
 a83041a <=( (not A269)  and  (not A268) );
 a83044a <=( (not A299)  and  (not A298) );
 a83045a <=( a83044a  and  a83041a );
 a83046a <=( a83045a  and  a83038a );
 a83050a <=( A167  and  (not A169) );
 a83051a <=( A170  and  a83050a );
 a83054a <=( (not A199)  and  (not A166) );
 a83057a <=( (not A233)  and  (not A200) );
 a83058a <=( a83057a  and  a83054a );
 a83059a <=( a83058a  and  a83051a );
 a83063a <=( (not A266)  and  (not A236) );
 a83064a <=( (not A235)  and  a83063a );
 a83067a <=( A298  and  (not A267) );
 a83070a <=( (not A302)  and  (not A301) );
 a83071a <=( a83070a  and  a83067a );
 a83072a <=( a83071a  and  a83064a );
 a83076a <=( A167  and  (not A169) );
 a83077a <=( A170  and  a83076a );
 a83080a <=( (not A199)  and  (not A166) );
 a83083a <=( (not A233)  and  (not A200) );
 a83084a <=( a83083a  and  a83080a );
 a83085a <=( a83084a  and  a83077a );
 a83089a <=( (not A265)  and  (not A236) );
 a83090a <=( (not A235)  and  a83089a );
 a83093a <=( A298  and  (not A266) );
 a83096a <=( (not A302)  and  (not A301) );
 a83097a <=( a83096a  and  a83093a );
 a83098a <=( a83097a  and  a83090a );
 a83102a <=( A167  and  (not A169) );
 a83103a <=( A170  and  a83102a );
 a83106a <=( (not A199)  and  (not A166) );
 a83109a <=( (not A233)  and  (not A200) );
 a83110a <=( a83109a  and  a83106a );
 a83111a <=( a83110a  and  a83103a );
 a83115a <=( (not A268)  and  (not A266) );
 a83116a <=( (not A234)  and  a83115a );
 a83119a <=( A298  and  (not A269) );
 a83122a <=( (not A302)  and  (not A301) );
 a83123a <=( a83122a  and  a83119a );
 a83124a <=( a83123a  and  a83116a );
 a83128a <=( A167  and  (not A169) );
 a83129a <=( A170  and  a83128a );
 a83132a <=( (not A199)  and  (not A166) );
 a83135a <=( A232  and  (not A200) );
 a83136a <=( a83135a  and  a83132a );
 a83137a <=( a83136a  and  a83129a );
 a83141a <=( A235  and  A234 );
 a83142a <=( (not A233)  and  a83141a );
 a83145a <=( (not A299)  and  A298 );
 a83148a <=( A301  and  A300 );
 a83149a <=( a83148a  and  a83145a );
 a83150a <=( a83149a  and  a83142a );
 a83154a <=( A167  and  (not A169) );
 a83155a <=( A170  and  a83154a );
 a83158a <=( (not A199)  and  (not A166) );
 a83161a <=( A232  and  (not A200) );
 a83162a <=( a83161a  and  a83158a );
 a83163a <=( a83162a  and  a83155a );
 a83167a <=( A235  and  A234 );
 a83168a <=( (not A233)  and  a83167a );
 a83171a <=( (not A299)  and  A298 );
 a83174a <=( A302  and  A300 );
 a83175a <=( a83174a  and  a83171a );
 a83176a <=( a83175a  and  a83168a );
 a83180a <=( A167  and  (not A169) );
 a83181a <=( A170  and  a83180a );
 a83184a <=( (not A199)  and  (not A166) );
 a83187a <=( A232  and  (not A200) );
 a83188a <=( a83187a  and  a83184a );
 a83189a <=( a83188a  and  a83181a );
 a83193a <=( A235  and  A234 );
 a83194a <=( (not A233)  and  a83193a );
 a83197a <=( (not A266)  and  A265 );
 a83200a <=( A268  and  A267 );
 a83201a <=( a83200a  and  a83197a );
 a83202a <=( a83201a  and  a83194a );
 a83206a <=( A167  and  (not A169) );
 a83207a <=( A170  and  a83206a );
 a83210a <=( (not A199)  and  (not A166) );
 a83213a <=( A232  and  (not A200) );
 a83214a <=( a83213a  and  a83210a );
 a83215a <=( a83214a  and  a83207a );
 a83219a <=( A235  and  A234 );
 a83220a <=( (not A233)  and  a83219a );
 a83223a <=( (not A266)  and  A265 );
 a83226a <=( A269  and  A267 );
 a83227a <=( a83226a  and  a83223a );
 a83228a <=( a83227a  and  a83220a );
 a83232a <=( A167  and  (not A169) );
 a83233a <=( A170  and  a83232a );
 a83236a <=( (not A199)  and  (not A166) );
 a83239a <=( A232  and  (not A200) );
 a83240a <=( a83239a  and  a83236a );
 a83241a <=( a83240a  and  a83233a );
 a83245a <=( A236  and  A234 );
 a83246a <=( (not A233)  and  a83245a );
 a83249a <=( (not A299)  and  A298 );
 a83252a <=( A301  and  A300 );
 a83253a <=( a83252a  and  a83249a );
 a83254a <=( a83253a  and  a83246a );
 a83258a <=( A167  and  (not A169) );
 a83259a <=( A170  and  a83258a );
 a83262a <=( (not A199)  and  (not A166) );
 a83265a <=( A232  and  (not A200) );
 a83266a <=( a83265a  and  a83262a );
 a83267a <=( a83266a  and  a83259a );
 a83271a <=( A236  and  A234 );
 a83272a <=( (not A233)  and  a83271a );
 a83275a <=( (not A299)  and  A298 );
 a83278a <=( A302  and  A300 );
 a83279a <=( a83278a  and  a83275a );
 a83280a <=( a83279a  and  a83272a );
 a83284a <=( A167  and  (not A169) );
 a83285a <=( A170  and  a83284a );
 a83288a <=( (not A199)  and  (not A166) );
 a83291a <=( A232  and  (not A200) );
 a83292a <=( a83291a  and  a83288a );
 a83293a <=( a83292a  and  a83285a );
 a83297a <=( A236  and  A234 );
 a83298a <=( (not A233)  and  a83297a );
 a83301a <=( (not A266)  and  A265 );
 a83304a <=( A268  and  A267 );
 a83305a <=( a83304a  and  a83301a );
 a83306a <=( a83305a  and  a83298a );
 a83310a <=( A167  and  (not A169) );
 a83311a <=( A170  and  a83310a );
 a83314a <=( (not A199)  and  (not A166) );
 a83317a <=( A232  and  (not A200) );
 a83318a <=( a83317a  and  a83314a );
 a83319a <=( a83318a  and  a83311a );
 a83323a <=( A236  and  A234 );
 a83324a <=( (not A233)  and  a83323a );
 a83327a <=( (not A266)  and  A265 );
 a83330a <=( A269  and  A267 );
 a83331a <=( a83330a  and  a83327a );
 a83332a <=( a83331a  and  a83324a );
 a83336a <=( A167  and  (not A169) );
 a83337a <=( A170  and  a83336a );
 a83340a <=( (not A199)  and  (not A166) );
 a83343a <=( (not A232)  and  (not A200) );
 a83344a <=( a83343a  and  a83340a );
 a83345a <=( a83344a  and  a83337a );
 a83349a <=( (not A268)  and  (not A266) );
 a83350a <=( (not A233)  and  a83349a );
 a83353a <=( A298  and  (not A269) );
 a83356a <=( (not A302)  and  (not A301) );
 a83357a <=( a83356a  and  a83353a );
 a83358a <=( a83357a  and  a83350a );
 a83362a <=( (not A167)  and  (not A169) );
 a83363a <=( A170  and  a83362a );
 a83366a <=( A199  and  A166 );
 a83369a <=( A232  and  A200 );
 a83370a <=( a83369a  and  a83366a );
 a83371a <=( a83370a  and  a83363a );
 a83375a <=( (not A268)  and  A265 );
 a83376a <=( A233  and  a83375a );
 a83379a <=( (not A299)  and  (not A269) );
 a83382a <=( (not A302)  and  (not A301) );
 a83383a <=( a83382a  and  a83379a );
 a83384a <=( a83383a  and  a83376a );
 a83388a <=( (not A167)  and  (not A169) );
 a83389a <=( A170  and  a83388a );
 a83392a <=( A199  and  A166 );
 a83395a <=( (not A233)  and  A200 );
 a83396a <=( a83395a  and  a83392a );
 a83397a <=( a83396a  and  a83389a );
 a83401a <=( A265  and  (not A236) );
 a83402a <=( (not A235)  and  a83401a );
 a83405a <=( A298  and  A266 );
 a83408a <=( (not A302)  and  (not A301) );
 a83409a <=( a83408a  and  a83405a );
 a83410a <=( a83409a  and  a83402a );
 a83414a <=( (not A167)  and  (not A169) );
 a83415a <=( A170  and  a83414a );
 a83418a <=( A199  and  A166 );
 a83421a <=( (not A233)  and  A200 );
 a83422a <=( a83421a  and  a83418a );
 a83423a <=( a83422a  and  a83415a );
 a83427a <=( (not A266)  and  (not A236) );
 a83428a <=( (not A235)  and  a83427a );
 a83431a <=( (not A269)  and  (not A268) );
 a83434a <=( (not A300)  and  A298 );
 a83435a <=( a83434a  and  a83431a );
 a83436a <=( a83435a  and  a83428a );
 a83440a <=( (not A167)  and  (not A169) );
 a83441a <=( A170  and  a83440a );
 a83444a <=( A199  and  A166 );
 a83447a <=( (not A233)  and  A200 );
 a83448a <=( a83447a  and  a83444a );
 a83449a <=( a83448a  and  a83441a );
 a83453a <=( (not A266)  and  (not A236) );
 a83454a <=( (not A235)  and  a83453a );
 a83457a <=( (not A269)  and  (not A268) );
 a83460a <=( A299  and  A298 );
 a83461a <=( a83460a  and  a83457a );
 a83462a <=( a83461a  and  a83454a );
 a83466a <=( (not A167)  and  (not A169) );
 a83467a <=( A170  and  a83466a );
 a83470a <=( A199  and  A166 );
 a83473a <=( (not A233)  and  A200 );
 a83474a <=( a83473a  and  a83470a );
 a83475a <=( a83474a  and  a83467a );
 a83479a <=( (not A266)  and  (not A236) );
 a83480a <=( (not A235)  and  a83479a );
 a83483a <=( (not A269)  and  (not A268) );
 a83486a <=( (not A299)  and  (not A298) );
 a83487a <=( a83486a  and  a83483a );
 a83488a <=( a83487a  and  a83480a );
 a83492a <=( (not A167)  and  (not A169) );
 a83493a <=( A170  and  a83492a );
 a83496a <=( A199  and  A166 );
 a83499a <=( (not A233)  and  A200 );
 a83500a <=( a83499a  and  a83496a );
 a83501a <=( a83500a  and  a83493a );
 a83505a <=( (not A266)  and  (not A236) );
 a83506a <=( (not A235)  and  a83505a );
 a83509a <=( A298  and  (not A267) );
 a83512a <=( (not A302)  and  (not A301) );
 a83513a <=( a83512a  and  a83509a );
 a83514a <=( a83513a  and  a83506a );
 a83518a <=( (not A167)  and  (not A169) );
 a83519a <=( A170  and  a83518a );
 a83522a <=( A199  and  A166 );
 a83525a <=( (not A233)  and  A200 );
 a83526a <=( a83525a  and  a83522a );
 a83527a <=( a83526a  and  a83519a );
 a83531a <=( (not A265)  and  (not A236) );
 a83532a <=( (not A235)  and  a83531a );
 a83535a <=( A298  and  (not A266) );
 a83538a <=( (not A302)  and  (not A301) );
 a83539a <=( a83538a  and  a83535a );
 a83540a <=( a83539a  and  a83532a );
 a83544a <=( (not A167)  and  (not A169) );
 a83545a <=( A170  and  a83544a );
 a83548a <=( A199  and  A166 );
 a83551a <=( (not A233)  and  A200 );
 a83552a <=( a83551a  and  a83548a );
 a83553a <=( a83552a  and  a83545a );
 a83557a <=( (not A268)  and  (not A266) );
 a83558a <=( (not A234)  and  a83557a );
 a83561a <=( A298  and  (not A269) );
 a83564a <=( (not A302)  and  (not A301) );
 a83565a <=( a83564a  and  a83561a );
 a83566a <=( a83565a  and  a83558a );
 a83570a <=( (not A167)  and  (not A169) );
 a83571a <=( A170  and  a83570a );
 a83574a <=( A199  and  A166 );
 a83577a <=( A232  and  A200 );
 a83578a <=( a83577a  and  a83574a );
 a83579a <=( a83578a  and  a83571a );
 a83583a <=( A235  and  A234 );
 a83584a <=( (not A233)  and  a83583a );
 a83587a <=( (not A299)  and  A298 );
 a83590a <=( A301  and  A300 );
 a83591a <=( a83590a  and  a83587a );
 a83592a <=( a83591a  and  a83584a );
 a83596a <=( (not A167)  and  (not A169) );
 a83597a <=( A170  and  a83596a );
 a83600a <=( A199  and  A166 );
 a83603a <=( A232  and  A200 );
 a83604a <=( a83603a  and  a83600a );
 a83605a <=( a83604a  and  a83597a );
 a83609a <=( A235  and  A234 );
 a83610a <=( (not A233)  and  a83609a );
 a83613a <=( (not A299)  and  A298 );
 a83616a <=( A302  and  A300 );
 a83617a <=( a83616a  and  a83613a );
 a83618a <=( a83617a  and  a83610a );
 a83622a <=( (not A167)  and  (not A169) );
 a83623a <=( A170  and  a83622a );
 a83626a <=( A199  and  A166 );
 a83629a <=( A232  and  A200 );
 a83630a <=( a83629a  and  a83626a );
 a83631a <=( a83630a  and  a83623a );
 a83635a <=( A235  and  A234 );
 a83636a <=( (not A233)  and  a83635a );
 a83639a <=( (not A266)  and  A265 );
 a83642a <=( A268  and  A267 );
 a83643a <=( a83642a  and  a83639a );
 a83644a <=( a83643a  and  a83636a );
 a83648a <=( (not A167)  and  (not A169) );
 a83649a <=( A170  and  a83648a );
 a83652a <=( A199  and  A166 );
 a83655a <=( A232  and  A200 );
 a83656a <=( a83655a  and  a83652a );
 a83657a <=( a83656a  and  a83649a );
 a83661a <=( A235  and  A234 );
 a83662a <=( (not A233)  and  a83661a );
 a83665a <=( (not A266)  and  A265 );
 a83668a <=( A269  and  A267 );
 a83669a <=( a83668a  and  a83665a );
 a83670a <=( a83669a  and  a83662a );
 a83674a <=( (not A167)  and  (not A169) );
 a83675a <=( A170  and  a83674a );
 a83678a <=( A199  and  A166 );
 a83681a <=( A232  and  A200 );
 a83682a <=( a83681a  and  a83678a );
 a83683a <=( a83682a  and  a83675a );
 a83687a <=( A236  and  A234 );
 a83688a <=( (not A233)  and  a83687a );
 a83691a <=( (not A299)  and  A298 );
 a83694a <=( A301  and  A300 );
 a83695a <=( a83694a  and  a83691a );
 a83696a <=( a83695a  and  a83688a );
 a83700a <=( (not A167)  and  (not A169) );
 a83701a <=( A170  and  a83700a );
 a83704a <=( A199  and  A166 );
 a83707a <=( A232  and  A200 );
 a83708a <=( a83707a  and  a83704a );
 a83709a <=( a83708a  and  a83701a );
 a83713a <=( A236  and  A234 );
 a83714a <=( (not A233)  and  a83713a );
 a83717a <=( (not A299)  and  A298 );
 a83720a <=( A302  and  A300 );
 a83721a <=( a83720a  and  a83717a );
 a83722a <=( a83721a  and  a83714a );
 a83726a <=( (not A167)  and  (not A169) );
 a83727a <=( A170  and  a83726a );
 a83730a <=( A199  and  A166 );
 a83733a <=( A232  and  A200 );
 a83734a <=( a83733a  and  a83730a );
 a83735a <=( a83734a  and  a83727a );
 a83739a <=( A236  and  A234 );
 a83740a <=( (not A233)  and  a83739a );
 a83743a <=( (not A266)  and  A265 );
 a83746a <=( A268  and  A267 );
 a83747a <=( a83746a  and  a83743a );
 a83748a <=( a83747a  and  a83740a );
 a83752a <=( (not A167)  and  (not A169) );
 a83753a <=( A170  and  a83752a );
 a83756a <=( A199  and  A166 );
 a83759a <=( A232  and  A200 );
 a83760a <=( a83759a  and  a83756a );
 a83761a <=( a83760a  and  a83753a );
 a83765a <=( A236  and  A234 );
 a83766a <=( (not A233)  and  a83765a );
 a83769a <=( (not A266)  and  A265 );
 a83772a <=( A269  and  A267 );
 a83773a <=( a83772a  and  a83769a );
 a83774a <=( a83773a  and  a83766a );
 a83778a <=( (not A167)  and  (not A169) );
 a83779a <=( A170  and  a83778a );
 a83782a <=( A199  and  A166 );
 a83785a <=( (not A232)  and  A200 );
 a83786a <=( a83785a  and  a83782a );
 a83787a <=( a83786a  and  a83779a );
 a83791a <=( (not A268)  and  (not A266) );
 a83792a <=( (not A233)  and  a83791a );
 a83795a <=( A298  and  (not A269) );
 a83798a <=( (not A302)  and  (not A301) );
 a83799a <=( a83798a  and  a83795a );
 a83800a <=( a83799a  and  a83792a );
 a83804a <=( (not A167)  and  (not A169) );
 a83805a <=( A170  and  a83804a );
 a83808a <=( (not A200)  and  A166 );
 a83811a <=( (not A203)  and  (not A202) );
 a83812a <=( a83811a  and  a83808a );
 a83813a <=( a83812a  and  a83805a );
 a83817a <=( A265  and  A233 );
 a83818a <=( A232  and  a83817a );
 a83821a <=( (not A269)  and  (not A268) );
 a83824a <=( (not A300)  and  (not A299) );
 a83825a <=( a83824a  and  a83821a );
 a83826a <=( a83825a  and  a83818a );
 a83830a <=( (not A167)  and  (not A169) );
 a83831a <=( A170  and  a83830a );
 a83834a <=( (not A200)  and  A166 );
 a83837a <=( (not A203)  and  (not A202) );
 a83838a <=( a83837a  and  a83834a );
 a83839a <=( a83838a  and  a83831a );
 a83843a <=( A265  and  A233 );
 a83844a <=( A232  and  a83843a );
 a83847a <=( (not A269)  and  (not A268) );
 a83850a <=( A299  and  A298 );
 a83851a <=( a83850a  and  a83847a );
 a83852a <=( a83851a  and  a83844a );
 a83856a <=( (not A167)  and  (not A169) );
 a83857a <=( A170  and  a83856a );
 a83860a <=( (not A200)  and  A166 );
 a83863a <=( (not A203)  and  (not A202) );
 a83864a <=( a83863a  and  a83860a );
 a83865a <=( a83864a  and  a83857a );
 a83869a <=( A265  and  A233 );
 a83870a <=( A232  and  a83869a );
 a83873a <=( (not A269)  and  (not A268) );
 a83876a <=( (not A299)  and  (not A298) );
 a83877a <=( a83876a  and  a83873a );
 a83878a <=( a83877a  and  a83870a );
 a83882a <=( (not A167)  and  (not A169) );
 a83883a <=( A170  and  a83882a );
 a83886a <=( (not A200)  and  A166 );
 a83889a <=( (not A203)  and  (not A202) );
 a83890a <=( a83889a  and  a83886a );
 a83891a <=( a83890a  and  a83883a );
 a83895a <=( A265  and  A233 );
 a83896a <=( A232  and  a83895a );
 a83899a <=( (not A299)  and  (not A267) );
 a83902a <=( (not A302)  and  (not A301) );
 a83903a <=( a83902a  and  a83899a );
 a83904a <=( a83903a  and  a83896a );
 a83908a <=( (not A167)  and  (not A169) );
 a83909a <=( A170  and  a83908a );
 a83912a <=( (not A200)  and  A166 );
 a83915a <=( (not A203)  and  (not A202) );
 a83916a <=( a83915a  and  a83912a );
 a83917a <=( a83916a  and  a83909a );
 a83921a <=( A265  and  A233 );
 a83922a <=( A232  and  a83921a );
 a83925a <=( (not A299)  and  A266 );
 a83928a <=( (not A302)  and  (not A301) );
 a83929a <=( a83928a  and  a83925a );
 a83930a <=( a83929a  and  a83922a );
 a83934a <=( (not A167)  and  (not A169) );
 a83935a <=( A170  and  a83934a );
 a83938a <=( (not A200)  and  A166 );
 a83941a <=( (not A203)  and  (not A202) );
 a83942a <=( a83941a  and  a83938a );
 a83943a <=( a83942a  and  a83935a );
 a83947a <=( (not A265)  and  A233 );
 a83948a <=( A232  and  a83947a );
 a83951a <=( (not A299)  and  (not A266) );
 a83954a <=( (not A302)  and  (not A301) );
 a83955a <=( a83954a  and  a83951a );
 a83956a <=( a83955a  and  a83948a );
 a83960a <=( (not A167)  and  (not A169) );
 a83961a <=( A170  and  a83960a );
 a83964a <=( (not A200)  and  A166 );
 a83967a <=( (not A203)  and  (not A202) );
 a83968a <=( a83967a  and  a83964a );
 a83969a <=( a83968a  and  a83961a );
 a83973a <=( (not A236)  and  (not A235) );
 a83974a <=( (not A233)  and  a83973a );
 a83977a <=( A266  and  A265 );
 a83980a <=( (not A300)  and  A298 );
 a83981a <=( a83980a  and  a83977a );
 a83982a <=( a83981a  and  a83974a );
 a83986a <=( (not A167)  and  (not A169) );
 a83987a <=( A170  and  a83986a );
 a83990a <=( (not A200)  and  A166 );
 a83993a <=( (not A203)  and  (not A202) );
 a83994a <=( a83993a  and  a83990a );
 a83995a <=( a83994a  and  a83987a );
 a83999a <=( (not A236)  and  (not A235) );
 a84000a <=( (not A233)  and  a83999a );
 a84003a <=( A266  and  A265 );
 a84006a <=( A299  and  A298 );
 a84007a <=( a84006a  and  a84003a );
 a84008a <=( a84007a  and  a84000a );
 a84012a <=( (not A167)  and  (not A169) );
 a84013a <=( A170  and  a84012a );
 a84016a <=( (not A200)  and  A166 );
 a84019a <=( (not A203)  and  (not A202) );
 a84020a <=( a84019a  and  a84016a );
 a84021a <=( a84020a  and  a84013a );
 a84025a <=( (not A236)  and  (not A235) );
 a84026a <=( (not A233)  and  a84025a );
 a84029a <=( A266  and  A265 );
 a84032a <=( (not A299)  and  (not A298) );
 a84033a <=( a84032a  and  a84029a );
 a84034a <=( a84033a  and  a84026a );
 a84038a <=( (not A167)  and  (not A169) );
 a84039a <=( A170  and  a84038a );
 a84042a <=( (not A200)  and  A166 );
 a84045a <=( (not A203)  and  (not A202) );
 a84046a <=( a84045a  and  a84042a );
 a84047a <=( a84046a  and  a84039a );
 a84051a <=( (not A236)  and  (not A235) );
 a84052a <=( (not A233)  and  a84051a );
 a84055a <=( (not A267)  and  (not A266) );
 a84058a <=( (not A300)  and  A298 );
 a84059a <=( a84058a  and  a84055a );
 a84060a <=( a84059a  and  a84052a );
 a84064a <=( (not A167)  and  (not A169) );
 a84065a <=( A170  and  a84064a );
 a84068a <=( (not A200)  and  A166 );
 a84071a <=( (not A203)  and  (not A202) );
 a84072a <=( a84071a  and  a84068a );
 a84073a <=( a84072a  and  a84065a );
 a84077a <=( (not A236)  and  (not A235) );
 a84078a <=( (not A233)  and  a84077a );
 a84081a <=( (not A267)  and  (not A266) );
 a84084a <=( A299  and  A298 );
 a84085a <=( a84084a  and  a84081a );
 a84086a <=( a84085a  and  a84078a );
 a84090a <=( (not A167)  and  (not A169) );
 a84091a <=( A170  and  a84090a );
 a84094a <=( (not A200)  and  A166 );
 a84097a <=( (not A203)  and  (not A202) );
 a84098a <=( a84097a  and  a84094a );
 a84099a <=( a84098a  and  a84091a );
 a84103a <=( (not A236)  and  (not A235) );
 a84104a <=( (not A233)  and  a84103a );
 a84107a <=( (not A267)  and  (not A266) );
 a84110a <=( (not A299)  and  (not A298) );
 a84111a <=( a84110a  and  a84107a );
 a84112a <=( a84111a  and  a84104a );
 a84116a <=( (not A167)  and  (not A169) );
 a84117a <=( A170  and  a84116a );
 a84120a <=( (not A200)  and  A166 );
 a84123a <=( (not A203)  and  (not A202) );
 a84124a <=( a84123a  and  a84120a );
 a84125a <=( a84124a  and  a84117a );
 a84129a <=( (not A236)  and  (not A235) );
 a84130a <=( (not A233)  and  a84129a );
 a84133a <=( (not A266)  and  (not A265) );
 a84136a <=( (not A300)  and  A298 );
 a84137a <=( a84136a  and  a84133a );
 a84138a <=( a84137a  and  a84130a );
 a84142a <=( (not A167)  and  (not A169) );
 a84143a <=( A170  and  a84142a );
 a84146a <=( (not A200)  and  A166 );
 a84149a <=( (not A203)  and  (not A202) );
 a84150a <=( a84149a  and  a84146a );
 a84151a <=( a84150a  and  a84143a );
 a84155a <=( (not A236)  and  (not A235) );
 a84156a <=( (not A233)  and  a84155a );
 a84159a <=( (not A266)  and  (not A265) );
 a84162a <=( A299  and  A298 );
 a84163a <=( a84162a  and  a84159a );
 a84164a <=( a84163a  and  a84156a );
 a84168a <=( (not A167)  and  (not A169) );
 a84169a <=( A170  and  a84168a );
 a84172a <=( (not A200)  and  A166 );
 a84175a <=( (not A203)  and  (not A202) );
 a84176a <=( a84175a  and  a84172a );
 a84177a <=( a84176a  and  a84169a );
 a84181a <=( (not A236)  and  (not A235) );
 a84182a <=( (not A233)  and  a84181a );
 a84185a <=( (not A266)  and  (not A265) );
 a84188a <=( (not A299)  and  (not A298) );
 a84189a <=( a84188a  and  a84185a );
 a84190a <=( a84189a  and  a84182a );
 a84194a <=( (not A167)  and  (not A169) );
 a84195a <=( A170  and  a84194a );
 a84198a <=( (not A200)  and  A166 );
 a84201a <=( (not A203)  and  (not A202) );
 a84202a <=( a84201a  and  a84198a );
 a84203a <=( a84202a  and  a84195a );
 a84207a <=( A265  and  (not A234) );
 a84208a <=( (not A233)  and  a84207a );
 a84211a <=( A298  and  A266 );
 a84214a <=( (not A302)  and  (not A301) );
 a84215a <=( a84214a  and  a84211a );
 a84216a <=( a84215a  and  a84208a );
 a84220a <=( (not A167)  and  (not A169) );
 a84221a <=( A170  and  a84220a );
 a84224a <=( (not A200)  and  A166 );
 a84227a <=( (not A203)  and  (not A202) );
 a84228a <=( a84227a  and  a84224a );
 a84229a <=( a84228a  and  a84221a );
 a84233a <=( (not A266)  and  (not A234) );
 a84234a <=( (not A233)  and  a84233a );
 a84237a <=( (not A269)  and  (not A268) );
 a84240a <=( (not A300)  and  A298 );
 a84241a <=( a84240a  and  a84237a );
 a84242a <=( a84241a  and  a84234a );
 a84246a <=( (not A167)  and  (not A169) );
 a84247a <=( A170  and  a84246a );
 a84250a <=( (not A200)  and  A166 );
 a84253a <=( (not A203)  and  (not A202) );
 a84254a <=( a84253a  and  a84250a );
 a84255a <=( a84254a  and  a84247a );
 a84259a <=( (not A266)  and  (not A234) );
 a84260a <=( (not A233)  and  a84259a );
 a84263a <=( (not A269)  and  (not A268) );
 a84266a <=( A299  and  A298 );
 a84267a <=( a84266a  and  a84263a );
 a84268a <=( a84267a  and  a84260a );
 a84272a <=( (not A167)  and  (not A169) );
 a84273a <=( A170  and  a84272a );
 a84276a <=( (not A200)  and  A166 );
 a84279a <=( (not A203)  and  (not A202) );
 a84280a <=( a84279a  and  a84276a );
 a84281a <=( a84280a  and  a84273a );
 a84285a <=( (not A266)  and  (not A234) );
 a84286a <=( (not A233)  and  a84285a );
 a84289a <=( (not A269)  and  (not A268) );
 a84292a <=( (not A299)  and  (not A298) );
 a84293a <=( a84292a  and  a84289a );
 a84294a <=( a84293a  and  a84286a );
 a84298a <=( (not A167)  and  (not A169) );
 a84299a <=( A170  and  a84298a );
 a84302a <=( (not A200)  and  A166 );
 a84305a <=( (not A203)  and  (not A202) );
 a84306a <=( a84305a  and  a84302a );
 a84307a <=( a84306a  and  a84299a );
 a84311a <=( (not A266)  and  (not A234) );
 a84312a <=( (not A233)  and  a84311a );
 a84315a <=( A298  and  (not A267) );
 a84318a <=( (not A302)  and  (not A301) );
 a84319a <=( a84318a  and  a84315a );
 a84320a <=( a84319a  and  a84312a );
 a84324a <=( (not A167)  and  (not A169) );
 a84325a <=( A170  and  a84324a );
 a84328a <=( (not A200)  and  A166 );
 a84331a <=( (not A203)  and  (not A202) );
 a84332a <=( a84331a  and  a84328a );
 a84333a <=( a84332a  and  a84325a );
 a84337a <=( (not A265)  and  (not A234) );
 a84338a <=( (not A233)  and  a84337a );
 a84341a <=( A298  and  (not A266) );
 a84344a <=( (not A302)  and  (not A301) );
 a84345a <=( a84344a  and  a84341a );
 a84346a <=( a84345a  and  a84338a );
 a84350a <=( (not A167)  and  (not A169) );
 a84351a <=( A170  and  a84350a );
 a84354a <=( (not A200)  and  A166 );
 a84357a <=( (not A203)  and  (not A202) );
 a84358a <=( a84357a  and  a84354a );
 a84359a <=( a84358a  and  a84351a );
 a84363a <=( A265  and  (not A233) );
 a84364a <=( (not A232)  and  a84363a );
 a84367a <=( A298  and  A266 );
 a84370a <=( (not A302)  and  (not A301) );
 a84371a <=( a84370a  and  a84367a );
 a84372a <=( a84371a  and  a84364a );
 a84376a <=( (not A167)  and  (not A169) );
 a84377a <=( A170  and  a84376a );
 a84380a <=( (not A200)  and  A166 );
 a84383a <=( (not A203)  and  (not A202) );
 a84384a <=( a84383a  and  a84380a );
 a84385a <=( a84384a  and  a84377a );
 a84389a <=( (not A266)  and  (not A233) );
 a84390a <=( (not A232)  and  a84389a );
 a84393a <=( (not A269)  and  (not A268) );
 a84396a <=( (not A300)  and  A298 );
 a84397a <=( a84396a  and  a84393a );
 a84398a <=( a84397a  and  a84390a );
 a84402a <=( (not A167)  and  (not A169) );
 a84403a <=( A170  and  a84402a );
 a84406a <=( (not A200)  and  A166 );
 a84409a <=( (not A203)  and  (not A202) );
 a84410a <=( a84409a  and  a84406a );
 a84411a <=( a84410a  and  a84403a );
 a84415a <=( (not A266)  and  (not A233) );
 a84416a <=( (not A232)  and  a84415a );
 a84419a <=( (not A269)  and  (not A268) );
 a84422a <=( A299  and  A298 );
 a84423a <=( a84422a  and  a84419a );
 a84424a <=( a84423a  and  a84416a );
 a84428a <=( (not A167)  and  (not A169) );
 a84429a <=( A170  and  a84428a );
 a84432a <=( (not A200)  and  A166 );
 a84435a <=( (not A203)  and  (not A202) );
 a84436a <=( a84435a  and  a84432a );
 a84437a <=( a84436a  and  a84429a );
 a84441a <=( (not A266)  and  (not A233) );
 a84442a <=( (not A232)  and  a84441a );
 a84445a <=( (not A269)  and  (not A268) );
 a84448a <=( (not A299)  and  (not A298) );
 a84449a <=( a84448a  and  a84445a );
 a84450a <=( a84449a  and  a84442a );
 a84454a <=( (not A167)  and  (not A169) );
 a84455a <=( A170  and  a84454a );
 a84458a <=( (not A200)  and  A166 );
 a84461a <=( (not A203)  and  (not A202) );
 a84462a <=( a84461a  and  a84458a );
 a84463a <=( a84462a  and  a84455a );
 a84467a <=( (not A266)  and  (not A233) );
 a84468a <=( (not A232)  and  a84467a );
 a84471a <=( A298  and  (not A267) );
 a84474a <=( (not A302)  and  (not A301) );
 a84475a <=( a84474a  and  a84471a );
 a84476a <=( a84475a  and  a84468a );
 a84480a <=( (not A167)  and  (not A169) );
 a84481a <=( A170  and  a84480a );
 a84484a <=( (not A200)  and  A166 );
 a84487a <=( (not A203)  and  (not A202) );
 a84488a <=( a84487a  and  a84484a );
 a84489a <=( a84488a  and  a84481a );
 a84493a <=( (not A265)  and  (not A233) );
 a84494a <=( (not A232)  and  a84493a );
 a84497a <=( A298  and  (not A266) );
 a84500a <=( (not A302)  and  (not A301) );
 a84501a <=( a84500a  and  a84497a );
 a84502a <=( a84501a  and  a84494a );
 a84506a <=( (not A167)  and  (not A169) );
 a84507a <=( A170  and  a84506a );
 a84510a <=( (not A200)  and  A166 );
 a84513a <=( A232  and  (not A201) );
 a84514a <=( a84513a  and  a84510a );
 a84515a <=( a84514a  and  a84507a );
 a84519a <=( (not A268)  and  A265 );
 a84520a <=( A233  and  a84519a );
 a84523a <=( (not A299)  and  (not A269) );
 a84526a <=( (not A302)  and  (not A301) );
 a84527a <=( a84526a  and  a84523a );
 a84528a <=( a84527a  and  a84520a );
 a84532a <=( (not A167)  and  (not A169) );
 a84533a <=( A170  and  a84532a );
 a84536a <=( (not A200)  and  A166 );
 a84539a <=( (not A233)  and  (not A201) );
 a84540a <=( a84539a  and  a84536a );
 a84541a <=( a84540a  and  a84533a );
 a84545a <=( A265  and  (not A236) );
 a84546a <=( (not A235)  and  a84545a );
 a84549a <=( A298  and  A266 );
 a84552a <=( (not A302)  and  (not A301) );
 a84553a <=( a84552a  and  a84549a );
 a84554a <=( a84553a  and  a84546a );
 a84558a <=( (not A167)  and  (not A169) );
 a84559a <=( A170  and  a84558a );
 a84562a <=( (not A200)  and  A166 );
 a84565a <=( (not A233)  and  (not A201) );
 a84566a <=( a84565a  and  a84562a );
 a84567a <=( a84566a  and  a84559a );
 a84571a <=( (not A266)  and  (not A236) );
 a84572a <=( (not A235)  and  a84571a );
 a84575a <=( (not A269)  and  (not A268) );
 a84578a <=( (not A300)  and  A298 );
 a84579a <=( a84578a  and  a84575a );
 a84580a <=( a84579a  and  a84572a );
 a84584a <=( (not A167)  and  (not A169) );
 a84585a <=( A170  and  a84584a );
 a84588a <=( (not A200)  and  A166 );
 a84591a <=( (not A233)  and  (not A201) );
 a84592a <=( a84591a  and  a84588a );
 a84593a <=( a84592a  and  a84585a );
 a84597a <=( (not A266)  and  (not A236) );
 a84598a <=( (not A235)  and  a84597a );
 a84601a <=( (not A269)  and  (not A268) );
 a84604a <=( A299  and  A298 );
 a84605a <=( a84604a  and  a84601a );
 a84606a <=( a84605a  and  a84598a );
 a84610a <=( (not A167)  and  (not A169) );
 a84611a <=( A170  and  a84610a );
 a84614a <=( (not A200)  and  A166 );
 a84617a <=( (not A233)  and  (not A201) );
 a84618a <=( a84617a  and  a84614a );
 a84619a <=( a84618a  and  a84611a );
 a84623a <=( (not A266)  and  (not A236) );
 a84624a <=( (not A235)  and  a84623a );
 a84627a <=( (not A269)  and  (not A268) );
 a84630a <=( (not A299)  and  (not A298) );
 a84631a <=( a84630a  and  a84627a );
 a84632a <=( a84631a  and  a84624a );
 a84636a <=( (not A167)  and  (not A169) );
 a84637a <=( A170  and  a84636a );
 a84640a <=( (not A200)  and  A166 );
 a84643a <=( (not A233)  and  (not A201) );
 a84644a <=( a84643a  and  a84640a );
 a84645a <=( a84644a  and  a84637a );
 a84649a <=( (not A266)  and  (not A236) );
 a84650a <=( (not A235)  and  a84649a );
 a84653a <=( A298  and  (not A267) );
 a84656a <=( (not A302)  and  (not A301) );
 a84657a <=( a84656a  and  a84653a );
 a84658a <=( a84657a  and  a84650a );
 a84662a <=( (not A167)  and  (not A169) );
 a84663a <=( A170  and  a84662a );
 a84666a <=( (not A200)  and  A166 );
 a84669a <=( (not A233)  and  (not A201) );
 a84670a <=( a84669a  and  a84666a );
 a84671a <=( a84670a  and  a84663a );
 a84675a <=( (not A265)  and  (not A236) );
 a84676a <=( (not A235)  and  a84675a );
 a84679a <=( A298  and  (not A266) );
 a84682a <=( (not A302)  and  (not A301) );
 a84683a <=( a84682a  and  a84679a );
 a84684a <=( a84683a  and  a84676a );
 a84688a <=( (not A167)  and  (not A169) );
 a84689a <=( A170  and  a84688a );
 a84692a <=( (not A200)  and  A166 );
 a84695a <=( (not A233)  and  (not A201) );
 a84696a <=( a84695a  and  a84692a );
 a84697a <=( a84696a  and  a84689a );
 a84701a <=( (not A268)  and  (not A266) );
 a84702a <=( (not A234)  and  a84701a );
 a84705a <=( A298  and  (not A269) );
 a84708a <=( (not A302)  and  (not A301) );
 a84709a <=( a84708a  and  a84705a );
 a84710a <=( a84709a  and  a84702a );
 a84714a <=( (not A167)  and  (not A169) );
 a84715a <=( A170  and  a84714a );
 a84718a <=( (not A200)  and  A166 );
 a84721a <=( A232  and  (not A201) );
 a84722a <=( a84721a  and  a84718a );
 a84723a <=( a84722a  and  a84715a );
 a84727a <=( A235  and  A234 );
 a84728a <=( (not A233)  and  a84727a );
 a84731a <=( (not A299)  and  A298 );
 a84734a <=( A301  and  A300 );
 a84735a <=( a84734a  and  a84731a );
 a84736a <=( a84735a  and  a84728a );
 a84740a <=( (not A167)  and  (not A169) );
 a84741a <=( A170  and  a84740a );
 a84744a <=( (not A200)  and  A166 );
 a84747a <=( A232  and  (not A201) );
 a84748a <=( a84747a  and  a84744a );
 a84749a <=( a84748a  and  a84741a );
 a84753a <=( A235  and  A234 );
 a84754a <=( (not A233)  and  a84753a );
 a84757a <=( (not A299)  and  A298 );
 a84760a <=( A302  and  A300 );
 a84761a <=( a84760a  and  a84757a );
 a84762a <=( a84761a  and  a84754a );
 a84766a <=( (not A167)  and  (not A169) );
 a84767a <=( A170  and  a84766a );
 a84770a <=( (not A200)  and  A166 );
 a84773a <=( A232  and  (not A201) );
 a84774a <=( a84773a  and  a84770a );
 a84775a <=( a84774a  and  a84767a );
 a84779a <=( A235  and  A234 );
 a84780a <=( (not A233)  and  a84779a );
 a84783a <=( (not A266)  and  A265 );
 a84786a <=( A268  and  A267 );
 a84787a <=( a84786a  and  a84783a );
 a84788a <=( a84787a  and  a84780a );
 a84792a <=( (not A167)  and  (not A169) );
 a84793a <=( A170  and  a84792a );
 a84796a <=( (not A200)  and  A166 );
 a84799a <=( A232  and  (not A201) );
 a84800a <=( a84799a  and  a84796a );
 a84801a <=( a84800a  and  a84793a );
 a84805a <=( A235  and  A234 );
 a84806a <=( (not A233)  and  a84805a );
 a84809a <=( (not A266)  and  A265 );
 a84812a <=( A269  and  A267 );
 a84813a <=( a84812a  and  a84809a );
 a84814a <=( a84813a  and  a84806a );
 a84818a <=( (not A167)  and  (not A169) );
 a84819a <=( A170  and  a84818a );
 a84822a <=( (not A200)  and  A166 );
 a84825a <=( A232  and  (not A201) );
 a84826a <=( a84825a  and  a84822a );
 a84827a <=( a84826a  and  a84819a );
 a84831a <=( A236  and  A234 );
 a84832a <=( (not A233)  and  a84831a );
 a84835a <=( (not A299)  and  A298 );
 a84838a <=( A301  and  A300 );
 a84839a <=( a84838a  and  a84835a );
 a84840a <=( a84839a  and  a84832a );
 a84844a <=( (not A167)  and  (not A169) );
 a84845a <=( A170  and  a84844a );
 a84848a <=( (not A200)  and  A166 );
 a84851a <=( A232  and  (not A201) );
 a84852a <=( a84851a  and  a84848a );
 a84853a <=( a84852a  and  a84845a );
 a84857a <=( A236  and  A234 );
 a84858a <=( (not A233)  and  a84857a );
 a84861a <=( (not A299)  and  A298 );
 a84864a <=( A302  and  A300 );
 a84865a <=( a84864a  and  a84861a );
 a84866a <=( a84865a  and  a84858a );
 a84870a <=( (not A167)  and  (not A169) );
 a84871a <=( A170  and  a84870a );
 a84874a <=( (not A200)  and  A166 );
 a84877a <=( A232  and  (not A201) );
 a84878a <=( a84877a  and  a84874a );
 a84879a <=( a84878a  and  a84871a );
 a84883a <=( A236  and  A234 );
 a84884a <=( (not A233)  and  a84883a );
 a84887a <=( (not A266)  and  A265 );
 a84890a <=( A268  and  A267 );
 a84891a <=( a84890a  and  a84887a );
 a84892a <=( a84891a  and  a84884a );
 a84896a <=( (not A167)  and  (not A169) );
 a84897a <=( A170  and  a84896a );
 a84900a <=( (not A200)  and  A166 );
 a84903a <=( A232  and  (not A201) );
 a84904a <=( a84903a  and  a84900a );
 a84905a <=( a84904a  and  a84897a );
 a84909a <=( A236  and  A234 );
 a84910a <=( (not A233)  and  a84909a );
 a84913a <=( (not A266)  and  A265 );
 a84916a <=( A269  and  A267 );
 a84917a <=( a84916a  and  a84913a );
 a84918a <=( a84917a  and  a84910a );
 a84922a <=( (not A167)  and  (not A169) );
 a84923a <=( A170  and  a84922a );
 a84926a <=( (not A200)  and  A166 );
 a84929a <=( (not A232)  and  (not A201) );
 a84930a <=( a84929a  and  a84926a );
 a84931a <=( a84930a  and  a84923a );
 a84935a <=( (not A268)  and  (not A266) );
 a84936a <=( (not A233)  and  a84935a );
 a84939a <=( A298  and  (not A269) );
 a84942a <=( (not A302)  and  (not A301) );
 a84943a <=( a84942a  and  a84939a );
 a84944a <=( a84943a  and  a84936a );
 a84948a <=( (not A167)  and  (not A169) );
 a84949a <=( A170  and  a84948a );
 a84952a <=( (not A199)  and  A166 );
 a84955a <=( A232  and  (not A200) );
 a84956a <=( a84955a  and  a84952a );
 a84957a <=( a84956a  and  a84949a );
 a84961a <=( (not A268)  and  A265 );
 a84962a <=( A233  and  a84961a );
 a84965a <=( (not A299)  and  (not A269) );
 a84968a <=( (not A302)  and  (not A301) );
 a84969a <=( a84968a  and  a84965a );
 a84970a <=( a84969a  and  a84962a );
 a84974a <=( (not A167)  and  (not A169) );
 a84975a <=( A170  and  a84974a );
 a84978a <=( (not A199)  and  A166 );
 a84981a <=( (not A233)  and  (not A200) );
 a84982a <=( a84981a  and  a84978a );
 a84983a <=( a84982a  and  a84975a );
 a84987a <=( A265  and  (not A236) );
 a84988a <=( (not A235)  and  a84987a );
 a84991a <=( A298  and  A266 );
 a84994a <=( (not A302)  and  (not A301) );
 a84995a <=( a84994a  and  a84991a );
 a84996a <=( a84995a  and  a84988a );
 a85000a <=( (not A167)  and  (not A169) );
 a85001a <=( A170  and  a85000a );
 a85004a <=( (not A199)  and  A166 );
 a85007a <=( (not A233)  and  (not A200) );
 a85008a <=( a85007a  and  a85004a );
 a85009a <=( a85008a  and  a85001a );
 a85013a <=( (not A266)  and  (not A236) );
 a85014a <=( (not A235)  and  a85013a );
 a85017a <=( (not A269)  and  (not A268) );
 a85020a <=( (not A300)  and  A298 );
 a85021a <=( a85020a  and  a85017a );
 a85022a <=( a85021a  and  a85014a );
 a85026a <=( (not A167)  and  (not A169) );
 a85027a <=( A170  and  a85026a );
 a85030a <=( (not A199)  and  A166 );
 a85033a <=( (not A233)  and  (not A200) );
 a85034a <=( a85033a  and  a85030a );
 a85035a <=( a85034a  and  a85027a );
 a85039a <=( (not A266)  and  (not A236) );
 a85040a <=( (not A235)  and  a85039a );
 a85043a <=( (not A269)  and  (not A268) );
 a85046a <=( A299  and  A298 );
 a85047a <=( a85046a  and  a85043a );
 a85048a <=( a85047a  and  a85040a );
 a85052a <=( (not A167)  and  (not A169) );
 a85053a <=( A170  and  a85052a );
 a85056a <=( (not A199)  and  A166 );
 a85059a <=( (not A233)  and  (not A200) );
 a85060a <=( a85059a  and  a85056a );
 a85061a <=( a85060a  and  a85053a );
 a85065a <=( (not A266)  and  (not A236) );
 a85066a <=( (not A235)  and  a85065a );
 a85069a <=( (not A269)  and  (not A268) );
 a85072a <=( (not A299)  and  (not A298) );
 a85073a <=( a85072a  and  a85069a );
 a85074a <=( a85073a  and  a85066a );
 a85078a <=( (not A167)  and  (not A169) );
 a85079a <=( A170  and  a85078a );
 a85082a <=( (not A199)  and  A166 );
 a85085a <=( (not A233)  and  (not A200) );
 a85086a <=( a85085a  and  a85082a );
 a85087a <=( a85086a  and  a85079a );
 a85091a <=( (not A266)  and  (not A236) );
 a85092a <=( (not A235)  and  a85091a );
 a85095a <=( A298  and  (not A267) );
 a85098a <=( (not A302)  and  (not A301) );
 a85099a <=( a85098a  and  a85095a );
 a85100a <=( a85099a  and  a85092a );
 a85104a <=( (not A167)  and  (not A169) );
 a85105a <=( A170  and  a85104a );
 a85108a <=( (not A199)  and  A166 );
 a85111a <=( (not A233)  and  (not A200) );
 a85112a <=( a85111a  and  a85108a );
 a85113a <=( a85112a  and  a85105a );
 a85117a <=( (not A265)  and  (not A236) );
 a85118a <=( (not A235)  and  a85117a );
 a85121a <=( A298  and  (not A266) );
 a85124a <=( (not A302)  and  (not A301) );
 a85125a <=( a85124a  and  a85121a );
 a85126a <=( a85125a  and  a85118a );
 a85130a <=( (not A167)  and  (not A169) );
 a85131a <=( A170  and  a85130a );
 a85134a <=( (not A199)  and  A166 );
 a85137a <=( (not A233)  and  (not A200) );
 a85138a <=( a85137a  and  a85134a );
 a85139a <=( a85138a  and  a85131a );
 a85143a <=( (not A268)  and  (not A266) );
 a85144a <=( (not A234)  and  a85143a );
 a85147a <=( A298  and  (not A269) );
 a85150a <=( (not A302)  and  (not A301) );
 a85151a <=( a85150a  and  a85147a );
 a85152a <=( a85151a  and  a85144a );
 a85156a <=( (not A167)  and  (not A169) );
 a85157a <=( A170  and  a85156a );
 a85160a <=( (not A199)  and  A166 );
 a85163a <=( A232  and  (not A200) );
 a85164a <=( a85163a  and  a85160a );
 a85165a <=( a85164a  and  a85157a );
 a85169a <=( A235  and  A234 );
 a85170a <=( (not A233)  and  a85169a );
 a85173a <=( (not A299)  and  A298 );
 a85176a <=( A301  and  A300 );
 a85177a <=( a85176a  and  a85173a );
 a85178a <=( a85177a  and  a85170a );
 a85182a <=( (not A167)  and  (not A169) );
 a85183a <=( A170  and  a85182a );
 a85186a <=( (not A199)  and  A166 );
 a85189a <=( A232  and  (not A200) );
 a85190a <=( a85189a  and  a85186a );
 a85191a <=( a85190a  and  a85183a );
 a85195a <=( A235  and  A234 );
 a85196a <=( (not A233)  and  a85195a );
 a85199a <=( (not A299)  and  A298 );
 a85202a <=( A302  and  A300 );
 a85203a <=( a85202a  and  a85199a );
 a85204a <=( a85203a  and  a85196a );
 a85208a <=( (not A167)  and  (not A169) );
 a85209a <=( A170  and  a85208a );
 a85212a <=( (not A199)  and  A166 );
 a85215a <=( A232  and  (not A200) );
 a85216a <=( a85215a  and  a85212a );
 a85217a <=( a85216a  and  a85209a );
 a85221a <=( A235  and  A234 );
 a85222a <=( (not A233)  and  a85221a );
 a85225a <=( (not A266)  and  A265 );
 a85228a <=( A268  and  A267 );
 a85229a <=( a85228a  and  a85225a );
 a85230a <=( a85229a  and  a85222a );
 a85234a <=( (not A167)  and  (not A169) );
 a85235a <=( A170  and  a85234a );
 a85238a <=( (not A199)  and  A166 );
 a85241a <=( A232  and  (not A200) );
 a85242a <=( a85241a  and  a85238a );
 a85243a <=( a85242a  and  a85235a );
 a85247a <=( A235  and  A234 );
 a85248a <=( (not A233)  and  a85247a );
 a85251a <=( (not A266)  and  A265 );
 a85254a <=( A269  and  A267 );
 a85255a <=( a85254a  and  a85251a );
 a85256a <=( a85255a  and  a85248a );
 a85260a <=( (not A167)  and  (not A169) );
 a85261a <=( A170  and  a85260a );
 a85264a <=( (not A199)  and  A166 );
 a85267a <=( A232  and  (not A200) );
 a85268a <=( a85267a  and  a85264a );
 a85269a <=( a85268a  and  a85261a );
 a85273a <=( A236  and  A234 );
 a85274a <=( (not A233)  and  a85273a );
 a85277a <=( (not A299)  and  A298 );
 a85280a <=( A301  and  A300 );
 a85281a <=( a85280a  and  a85277a );
 a85282a <=( a85281a  and  a85274a );
 a85286a <=( (not A167)  and  (not A169) );
 a85287a <=( A170  and  a85286a );
 a85290a <=( (not A199)  and  A166 );
 a85293a <=( A232  and  (not A200) );
 a85294a <=( a85293a  and  a85290a );
 a85295a <=( a85294a  and  a85287a );
 a85299a <=( A236  and  A234 );
 a85300a <=( (not A233)  and  a85299a );
 a85303a <=( (not A299)  and  A298 );
 a85306a <=( A302  and  A300 );
 a85307a <=( a85306a  and  a85303a );
 a85308a <=( a85307a  and  a85300a );
 a85312a <=( (not A167)  and  (not A169) );
 a85313a <=( A170  and  a85312a );
 a85316a <=( (not A199)  and  A166 );
 a85319a <=( A232  and  (not A200) );
 a85320a <=( a85319a  and  a85316a );
 a85321a <=( a85320a  and  a85313a );
 a85325a <=( A236  and  A234 );
 a85326a <=( (not A233)  and  a85325a );
 a85329a <=( (not A266)  and  A265 );
 a85332a <=( A268  and  A267 );
 a85333a <=( a85332a  and  a85329a );
 a85334a <=( a85333a  and  a85326a );
 a85338a <=( (not A167)  and  (not A169) );
 a85339a <=( A170  and  a85338a );
 a85342a <=( (not A199)  and  A166 );
 a85345a <=( A232  and  (not A200) );
 a85346a <=( a85345a  and  a85342a );
 a85347a <=( a85346a  and  a85339a );
 a85351a <=( A236  and  A234 );
 a85352a <=( (not A233)  and  a85351a );
 a85355a <=( (not A266)  and  A265 );
 a85358a <=( A269  and  A267 );
 a85359a <=( a85358a  and  a85355a );
 a85360a <=( a85359a  and  a85352a );
 a85364a <=( (not A167)  and  (not A169) );
 a85365a <=( A170  and  a85364a );
 a85368a <=( (not A199)  and  A166 );
 a85371a <=( (not A232)  and  (not A200) );
 a85372a <=( a85371a  and  a85368a );
 a85373a <=( a85372a  and  a85365a );
 a85377a <=( (not A268)  and  (not A266) );
 a85378a <=( (not A233)  and  a85377a );
 a85381a <=( A298  and  (not A269) );
 a85384a <=( (not A302)  and  (not A301) );
 a85385a <=( a85384a  and  a85381a );
 a85386a <=( a85385a  and  a85378a );
 a85390a <=( (not A168)  and  (not A169) );
 a85391a <=( (not A170)  and  a85390a );
 a85394a <=( (not A200)  and  A199 );
 a85397a <=( A202  and  A201 );
 a85398a <=( a85397a  and  a85394a );
 a85399a <=( a85398a  and  a85391a );
 a85403a <=( A265  and  A233 );
 a85404a <=( A232  and  a85403a );
 a85407a <=( (not A269)  and  (not A268) );
 a85410a <=( (not A300)  and  (not A299) );
 a85411a <=( a85410a  and  a85407a );
 a85412a <=( a85411a  and  a85404a );
 a85416a <=( (not A168)  and  (not A169) );
 a85417a <=( (not A170)  and  a85416a );
 a85420a <=( (not A200)  and  A199 );
 a85423a <=( A202  and  A201 );
 a85424a <=( a85423a  and  a85420a );
 a85425a <=( a85424a  and  a85417a );
 a85429a <=( A265  and  A233 );
 a85430a <=( A232  and  a85429a );
 a85433a <=( (not A269)  and  (not A268) );
 a85436a <=( A299  and  A298 );
 a85437a <=( a85436a  and  a85433a );
 a85438a <=( a85437a  and  a85430a );
 a85442a <=( (not A168)  and  (not A169) );
 a85443a <=( (not A170)  and  a85442a );
 a85446a <=( (not A200)  and  A199 );
 a85449a <=( A202  and  A201 );
 a85450a <=( a85449a  and  a85446a );
 a85451a <=( a85450a  and  a85443a );
 a85455a <=( A265  and  A233 );
 a85456a <=( A232  and  a85455a );
 a85459a <=( (not A269)  and  (not A268) );
 a85462a <=( (not A299)  and  (not A298) );
 a85463a <=( a85462a  and  a85459a );
 a85464a <=( a85463a  and  a85456a );
 a85468a <=( (not A168)  and  (not A169) );
 a85469a <=( (not A170)  and  a85468a );
 a85472a <=( (not A200)  and  A199 );
 a85475a <=( A202  and  A201 );
 a85476a <=( a85475a  and  a85472a );
 a85477a <=( a85476a  and  a85469a );
 a85481a <=( A265  and  A233 );
 a85482a <=( A232  and  a85481a );
 a85485a <=( (not A299)  and  (not A267) );
 a85488a <=( (not A302)  and  (not A301) );
 a85489a <=( a85488a  and  a85485a );
 a85490a <=( a85489a  and  a85482a );
 a85494a <=( (not A168)  and  (not A169) );
 a85495a <=( (not A170)  and  a85494a );
 a85498a <=( (not A200)  and  A199 );
 a85501a <=( A202  and  A201 );
 a85502a <=( a85501a  and  a85498a );
 a85503a <=( a85502a  and  a85495a );
 a85507a <=( A265  and  A233 );
 a85508a <=( A232  and  a85507a );
 a85511a <=( (not A299)  and  A266 );
 a85514a <=( (not A302)  and  (not A301) );
 a85515a <=( a85514a  and  a85511a );
 a85516a <=( a85515a  and  a85508a );
 a85520a <=( (not A168)  and  (not A169) );
 a85521a <=( (not A170)  and  a85520a );
 a85524a <=( (not A200)  and  A199 );
 a85527a <=( A202  and  A201 );
 a85528a <=( a85527a  and  a85524a );
 a85529a <=( a85528a  and  a85521a );
 a85533a <=( (not A265)  and  A233 );
 a85534a <=( A232  and  a85533a );
 a85537a <=( (not A299)  and  (not A266) );
 a85540a <=( (not A302)  and  (not A301) );
 a85541a <=( a85540a  and  a85537a );
 a85542a <=( a85541a  and  a85534a );
 a85546a <=( (not A168)  and  (not A169) );
 a85547a <=( (not A170)  and  a85546a );
 a85550a <=( (not A200)  and  A199 );
 a85553a <=( A202  and  A201 );
 a85554a <=( a85553a  and  a85550a );
 a85555a <=( a85554a  and  a85547a );
 a85559a <=( (not A236)  and  (not A235) );
 a85560a <=( (not A233)  and  a85559a );
 a85563a <=( A266  and  A265 );
 a85566a <=( (not A300)  and  A298 );
 a85567a <=( a85566a  and  a85563a );
 a85568a <=( a85567a  and  a85560a );
 a85572a <=( (not A168)  and  (not A169) );
 a85573a <=( (not A170)  and  a85572a );
 a85576a <=( (not A200)  and  A199 );
 a85579a <=( A202  and  A201 );
 a85580a <=( a85579a  and  a85576a );
 a85581a <=( a85580a  and  a85573a );
 a85585a <=( (not A236)  and  (not A235) );
 a85586a <=( (not A233)  and  a85585a );
 a85589a <=( A266  and  A265 );
 a85592a <=( A299  and  A298 );
 a85593a <=( a85592a  and  a85589a );
 a85594a <=( a85593a  and  a85586a );
 a85598a <=( (not A168)  and  (not A169) );
 a85599a <=( (not A170)  and  a85598a );
 a85602a <=( (not A200)  and  A199 );
 a85605a <=( A202  and  A201 );
 a85606a <=( a85605a  and  a85602a );
 a85607a <=( a85606a  and  a85599a );
 a85611a <=( (not A236)  and  (not A235) );
 a85612a <=( (not A233)  and  a85611a );
 a85615a <=( A266  and  A265 );
 a85618a <=( (not A299)  and  (not A298) );
 a85619a <=( a85618a  and  a85615a );
 a85620a <=( a85619a  and  a85612a );
 a85624a <=( (not A168)  and  (not A169) );
 a85625a <=( (not A170)  and  a85624a );
 a85628a <=( (not A200)  and  A199 );
 a85631a <=( A202  and  A201 );
 a85632a <=( a85631a  and  a85628a );
 a85633a <=( a85632a  and  a85625a );
 a85637a <=( (not A236)  and  (not A235) );
 a85638a <=( (not A233)  and  a85637a );
 a85641a <=( (not A267)  and  (not A266) );
 a85644a <=( (not A300)  and  A298 );
 a85645a <=( a85644a  and  a85641a );
 a85646a <=( a85645a  and  a85638a );
 a85650a <=( (not A168)  and  (not A169) );
 a85651a <=( (not A170)  and  a85650a );
 a85654a <=( (not A200)  and  A199 );
 a85657a <=( A202  and  A201 );
 a85658a <=( a85657a  and  a85654a );
 a85659a <=( a85658a  and  a85651a );
 a85663a <=( (not A236)  and  (not A235) );
 a85664a <=( (not A233)  and  a85663a );
 a85667a <=( (not A267)  and  (not A266) );
 a85670a <=( A299  and  A298 );
 a85671a <=( a85670a  and  a85667a );
 a85672a <=( a85671a  and  a85664a );
 a85676a <=( (not A168)  and  (not A169) );
 a85677a <=( (not A170)  and  a85676a );
 a85680a <=( (not A200)  and  A199 );
 a85683a <=( A202  and  A201 );
 a85684a <=( a85683a  and  a85680a );
 a85685a <=( a85684a  and  a85677a );
 a85689a <=( (not A236)  and  (not A235) );
 a85690a <=( (not A233)  and  a85689a );
 a85693a <=( (not A267)  and  (not A266) );
 a85696a <=( (not A299)  and  (not A298) );
 a85697a <=( a85696a  and  a85693a );
 a85698a <=( a85697a  and  a85690a );
 a85702a <=( (not A168)  and  (not A169) );
 a85703a <=( (not A170)  and  a85702a );
 a85706a <=( (not A200)  and  A199 );
 a85709a <=( A202  and  A201 );
 a85710a <=( a85709a  and  a85706a );
 a85711a <=( a85710a  and  a85703a );
 a85715a <=( (not A236)  and  (not A235) );
 a85716a <=( (not A233)  and  a85715a );
 a85719a <=( (not A266)  and  (not A265) );
 a85722a <=( (not A300)  and  A298 );
 a85723a <=( a85722a  and  a85719a );
 a85724a <=( a85723a  and  a85716a );
 a85728a <=( (not A168)  and  (not A169) );
 a85729a <=( (not A170)  and  a85728a );
 a85732a <=( (not A200)  and  A199 );
 a85735a <=( A202  and  A201 );
 a85736a <=( a85735a  and  a85732a );
 a85737a <=( a85736a  and  a85729a );
 a85741a <=( (not A236)  and  (not A235) );
 a85742a <=( (not A233)  and  a85741a );
 a85745a <=( (not A266)  and  (not A265) );
 a85748a <=( A299  and  A298 );
 a85749a <=( a85748a  and  a85745a );
 a85750a <=( a85749a  and  a85742a );
 a85754a <=( (not A168)  and  (not A169) );
 a85755a <=( (not A170)  and  a85754a );
 a85758a <=( (not A200)  and  A199 );
 a85761a <=( A202  and  A201 );
 a85762a <=( a85761a  and  a85758a );
 a85763a <=( a85762a  and  a85755a );
 a85767a <=( (not A236)  and  (not A235) );
 a85768a <=( (not A233)  and  a85767a );
 a85771a <=( (not A266)  and  (not A265) );
 a85774a <=( (not A299)  and  (not A298) );
 a85775a <=( a85774a  and  a85771a );
 a85776a <=( a85775a  and  a85768a );
 a85780a <=( (not A168)  and  (not A169) );
 a85781a <=( (not A170)  and  a85780a );
 a85784a <=( (not A200)  and  A199 );
 a85787a <=( A202  and  A201 );
 a85788a <=( a85787a  and  a85784a );
 a85789a <=( a85788a  and  a85781a );
 a85793a <=( A265  and  (not A234) );
 a85794a <=( (not A233)  and  a85793a );
 a85797a <=( A298  and  A266 );
 a85800a <=( (not A302)  and  (not A301) );
 a85801a <=( a85800a  and  a85797a );
 a85802a <=( a85801a  and  a85794a );
 a85806a <=( (not A168)  and  (not A169) );
 a85807a <=( (not A170)  and  a85806a );
 a85810a <=( (not A200)  and  A199 );
 a85813a <=( A202  and  A201 );
 a85814a <=( a85813a  and  a85810a );
 a85815a <=( a85814a  and  a85807a );
 a85819a <=( (not A266)  and  (not A234) );
 a85820a <=( (not A233)  and  a85819a );
 a85823a <=( (not A269)  and  (not A268) );
 a85826a <=( (not A300)  and  A298 );
 a85827a <=( a85826a  and  a85823a );
 a85828a <=( a85827a  and  a85820a );
 a85832a <=( (not A168)  and  (not A169) );
 a85833a <=( (not A170)  and  a85832a );
 a85836a <=( (not A200)  and  A199 );
 a85839a <=( A202  and  A201 );
 a85840a <=( a85839a  and  a85836a );
 a85841a <=( a85840a  and  a85833a );
 a85845a <=( (not A266)  and  (not A234) );
 a85846a <=( (not A233)  and  a85845a );
 a85849a <=( (not A269)  and  (not A268) );
 a85852a <=( A299  and  A298 );
 a85853a <=( a85852a  and  a85849a );
 a85854a <=( a85853a  and  a85846a );
 a85858a <=( (not A168)  and  (not A169) );
 a85859a <=( (not A170)  and  a85858a );
 a85862a <=( (not A200)  and  A199 );
 a85865a <=( A202  and  A201 );
 a85866a <=( a85865a  and  a85862a );
 a85867a <=( a85866a  and  a85859a );
 a85871a <=( (not A266)  and  (not A234) );
 a85872a <=( (not A233)  and  a85871a );
 a85875a <=( (not A269)  and  (not A268) );
 a85878a <=( (not A299)  and  (not A298) );
 a85879a <=( a85878a  and  a85875a );
 a85880a <=( a85879a  and  a85872a );
 a85884a <=( (not A168)  and  (not A169) );
 a85885a <=( (not A170)  and  a85884a );
 a85888a <=( (not A200)  and  A199 );
 a85891a <=( A202  and  A201 );
 a85892a <=( a85891a  and  a85888a );
 a85893a <=( a85892a  and  a85885a );
 a85897a <=( (not A266)  and  (not A234) );
 a85898a <=( (not A233)  and  a85897a );
 a85901a <=( A298  and  (not A267) );
 a85904a <=( (not A302)  and  (not A301) );
 a85905a <=( a85904a  and  a85901a );
 a85906a <=( a85905a  and  a85898a );
 a85910a <=( (not A168)  and  (not A169) );
 a85911a <=( (not A170)  and  a85910a );
 a85914a <=( (not A200)  and  A199 );
 a85917a <=( A202  and  A201 );
 a85918a <=( a85917a  and  a85914a );
 a85919a <=( a85918a  and  a85911a );
 a85923a <=( (not A265)  and  (not A234) );
 a85924a <=( (not A233)  and  a85923a );
 a85927a <=( A298  and  (not A266) );
 a85930a <=( (not A302)  and  (not A301) );
 a85931a <=( a85930a  and  a85927a );
 a85932a <=( a85931a  and  a85924a );
 a85936a <=( (not A168)  and  (not A169) );
 a85937a <=( (not A170)  and  a85936a );
 a85940a <=( (not A200)  and  A199 );
 a85943a <=( A202  and  A201 );
 a85944a <=( a85943a  and  a85940a );
 a85945a <=( a85944a  and  a85937a );
 a85949a <=( A265  and  (not A233) );
 a85950a <=( (not A232)  and  a85949a );
 a85953a <=( A298  and  A266 );
 a85956a <=( (not A302)  and  (not A301) );
 a85957a <=( a85956a  and  a85953a );
 a85958a <=( a85957a  and  a85950a );
 a85962a <=( (not A168)  and  (not A169) );
 a85963a <=( (not A170)  and  a85962a );
 a85966a <=( (not A200)  and  A199 );
 a85969a <=( A202  and  A201 );
 a85970a <=( a85969a  and  a85966a );
 a85971a <=( a85970a  and  a85963a );
 a85975a <=( (not A266)  and  (not A233) );
 a85976a <=( (not A232)  and  a85975a );
 a85979a <=( (not A269)  and  (not A268) );
 a85982a <=( (not A300)  and  A298 );
 a85983a <=( a85982a  and  a85979a );
 a85984a <=( a85983a  and  a85976a );
 a85988a <=( (not A168)  and  (not A169) );
 a85989a <=( (not A170)  and  a85988a );
 a85992a <=( (not A200)  and  A199 );
 a85995a <=( A202  and  A201 );
 a85996a <=( a85995a  and  a85992a );
 a85997a <=( a85996a  and  a85989a );
 a86001a <=( (not A266)  and  (not A233) );
 a86002a <=( (not A232)  and  a86001a );
 a86005a <=( (not A269)  and  (not A268) );
 a86008a <=( A299  and  A298 );
 a86009a <=( a86008a  and  a86005a );
 a86010a <=( a86009a  and  a86002a );
 a86014a <=( (not A168)  and  (not A169) );
 a86015a <=( (not A170)  and  a86014a );
 a86018a <=( (not A200)  and  A199 );
 a86021a <=( A202  and  A201 );
 a86022a <=( a86021a  and  a86018a );
 a86023a <=( a86022a  and  a86015a );
 a86027a <=( (not A266)  and  (not A233) );
 a86028a <=( (not A232)  and  a86027a );
 a86031a <=( (not A269)  and  (not A268) );
 a86034a <=( (not A299)  and  (not A298) );
 a86035a <=( a86034a  and  a86031a );
 a86036a <=( a86035a  and  a86028a );
 a86040a <=( (not A168)  and  (not A169) );
 a86041a <=( (not A170)  and  a86040a );
 a86044a <=( (not A200)  and  A199 );
 a86047a <=( A202  and  A201 );
 a86048a <=( a86047a  and  a86044a );
 a86049a <=( a86048a  and  a86041a );
 a86053a <=( (not A266)  and  (not A233) );
 a86054a <=( (not A232)  and  a86053a );
 a86057a <=( A298  and  (not A267) );
 a86060a <=( (not A302)  and  (not A301) );
 a86061a <=( a86060a  and  a86057a );
 a86062a <=( a86061a  and  a86054a );
 a86066a <=( (not A168)  and  (not A169) );
 a86067a <=( (not A170)  and  a86066a );
 a86070a <=( (not A200)  and  A199 );
 a86073a <=( A202  and  A201 );
 a86074a <=( a86073a  and  a86070a );
 a86075a <=( a86074a  and  a86067a );
 a86079a <=( (not A265)  and  (not A233) );
 a86080a <=( (not A232)  and  a86079a );
 a86083a <=( A298  and  (not A266) );
 a86086a <=( (not A302)  and  (not A301) );
 a86087a <=( a86086a  and  a86083a );
 a86088a <=( a86087a  and  a86080a );
 a86092a <=( (not A168)  and  (not A169) );
 a86093a <=( (not A170)  and  a86092a );
 a86096a <=( (not A200)  and  A199 );
 a86099a <=( A203  and  A201 );
 a86100a <=( a86099a  and  a86096a );
 a86101a <=( a86100a  and  a86093a );
 a86105a <=( A265  and  A233 );
 a86106a <=( A232  and  a86105a );
 a86109a <=( (not A269)  and  (not A268) );
 a86112a <=( (not A300)  and  (not A299) );
 a86113a <=( a86112a  and  a86109a );
 a86114a <=( a86113a  and  a86106a );
 a86118a <=( (not A168)  and  (not A169) );
 a86119a <=( (not A170)  and  a86118a );
 a86122a <=( (not A200)  and  A199 );
 a86125a <=( A203  and  A201 );
 a86126a <=( a86125a  and  a86122a );
 a86127a <=( a86126a  and  a86119a );
 a86131a <=( A265  and  A233 );
 a86132a <=( A232  and  a86131a );
 a86135a <=( (not A269)  and  (not A268) );
 a86138a <=( A299  and  A298 );
 a86139a <=( a86138a  and  a86135a );
 a86140a <=( a86139a  and  a86132a );
 a86144a <=( (not A168)  and  (not A169) );
 a86145a <=( (not A170)  and  a86144a );
 a86148a <=( (not A200)  and  A199 );
 a86151a <=( A203  and  A201 );
 a86152a <=( a86151a  and  a86148a );
 a86153a <=( a86152a  and  a86145a );
 a86157a <=( A265  and  A233 );
 a86158a <=( A232  and  a86157a );
 a86161a <=( (not A269)  and  (not A268) );
 a86164a <=( (not A299)  and  (not A298) );
 a86165a <=( a86164a  and  a86161a );
 a86166a <=( a86165a  and  a86158a );
 a86170a <=( (not A168)  and  (not A169) );
 a86171a <=( (not A170)  and  a86170a );
 a86174a <=( (not A200)  and  A199 );
 a86177a <=( A203  and  A201 );
 a86178a <=( a86177a  and  a86174a );
 a86179a <=( a86178a  and  a86171a );
 a86183a <=( A265  and  A233 );
 a86184a <=( A232  and  a86183a );
 a86187a <=( (not A299)  and  (not A267) );
 a86190a <=( (not A302)  and  (not A301) );
 a86191a <=( a86190a  and  a86187a );
 a86192a <=( a86191a  and  a86184a );
 a86196a <=( (not A168)  and  (not A169) );
 a86197a <=( (not A170)  and  a86196a );
 a86200a <=( (not A200)  and  A199 );
 a86203a <=( A203  and  A201 );
 a86204a <=( a86203a  and  a86200a );
 a86205a <=( a86204a  and  a86197a );
 a86209a <=( A265  and  A233 );
 a86210a <=( A232  and  a86209a );
 a86213a <=( (not A299)  and  A266 );
 a86216a <=( (not A302)  and  (not A301) );
 a86217a <=( a86216a  and  a86213a );
 a86218a <=( a86217a  and  a86210a );
 a86222a <=( (not A168)  and  (not A169) );
 a86223a <=( (not A170)  and  a86222a );
 a86226a <=( (not A200)  and  A199 );
 a86229a <=( A203  and  A201 );
 a86230a <=( a86229a  and  a86226a );
 a86231a <=( a86230a  and  a86223a );
 a86235a <=( (not A265)  and  A233 );
 a86236a <=( A232  and  a86235a );
 a86239a <=( (not A299)  and  (not A266) );
 a86242a <=( (not A302)  and  (not A301) );
 a86243a <=( a86242a  and  a86239a );
 a86244a <=( a86243a  and  a86236a );
 a86248a <=( (not A168)  and  (not A169) );
 a86249a <=( (not A170)  and  a86248a );
 a86252a <=( (not A200)  and  A199 );
 a86255a <=( A203  and  A201 );
 a86256a <=( a86255a  and  a86252a );
 a86257a <=( a86256a  and  a86249a );
 a86261a <=( (not A236)  and  (not A235) );
 a86262a <=( (not A233)  and  a86261a );
 a86265a <=( A266  and  A265 );
 a86268a <=( (not A300)  and  A298 );
 a86269a <=( a86268a  and  a86265a );
 a86270a <=( a86269a  and  a86262a );
 a86274a <=( (not A168)  and  (not A169) );
 a86275a <=( (not A170)  and  a86274a );
 a86278a <=( (not A200)  and  A199 );
 a86281a <=( A203  and  A201 );
 a86282a <=( a86281a  and  a86278a );
 a86283a <=( a86282a  and  a86275a );
 a86287a <=( (not A236)  and  (not A235) );
 a86288a <=( (not A233)  and  a86287a );
 a86291a <=( A266  and  A265 );
 a86294a <=( A299  and  A298 );
 a86295a <=( a86294a  and  a86291a );
 a86296a <=( a86295a  and  a86288a );
 a86300a <=( (not A168)  and  (not A169) );
 a86301a <=( (not A170)  and  a86300a );
 a86304a <=( (not A200)  and  A199 );
 a86307a <=( A203  and  A201 );
 a86308a <=( a86307a  and  a86304a );
 a86309a <=( a86308a  and  a86301a );
 a86313a <=( (not A236)  and  (not A235) );
 a86314a <=( (not A233)  and  a86313a );
 a86317a <=( A266  and  A265 );
 a86320a <=( (not A299)  and  (not A298) );
 a86321a <=( a86320a  and  a86317a );
 a86322a <=( a86321a  and  a86314a );
 a86326a <=( (not A168)  and  (not A169) );
 a86327a <=( (not A170)  and  a86326a );
 a86330a <=( (not A200)  and  A199 );
 a86333a <=( A203  and  A201 );
 a86334a <=( a86333a  and  a86330a );
 a86335a <=( a86334a  and  a86327a );
 a86339a <=( (not A236)  and  (not A235) );
 a86340a <=( (not A233)  and  a86339a );
 a86343a <=( (not A267)  and  (not A266) );
 a86346a <=( (not A300)  and  A298 );
 a86347a <=( a86346a  and  a86343a );
 a86348a <=( a86347a  and  a86340a );
 a86352a <=( (not A168)  and  (not A169) );
 a86353a <=( (not A170)  and  a86352a );
 a86356a <=( (not A200)  and  A199 );
 a86359a <=( A203  and  A201 );
 a86360a <=( a86359a  and  a86356a );
 a86361a <=( a86360a  and  a86353a );
 a86365a <=( (not A236)  and  (not A235) );
 a86366a <=( (not A233)  and  a86365a );
 a86369a <=( (not A267)  and  (not A266) );
 a86372a <=( A299  and  A298 );
 a86373a <=( a86372a  and  a86369a );
 a86374a <=( a86373a  and  a86366a );
 a86378a <=( (not A168)  and  (not A169) );
 a86379a <=( (not A170)  and  a86378a );
 a86382a <=( (not A200)  and  A199 );
 a86385a <=( A203  and  A201 );
 a86386a <=( a86385a  and  a86382a );
 a86387a <=( a86386a  and  a86379a );
 a86391a <=( (not A236)  and  (not A235) );
 a86392a <=( (not A233)  and  a86391a );
 a86395a <=( (not A267)  and  (not A266) );
 a86398a <=( (not A299)  and  (not A298) );
 a86399a <=( a86398a  and  a86395a );
 a86400a <=( a86399a  and  a86392a );
 a86404a <=( (not A168)  and  (not A169) );
 a86405a <=( (not A170)  and  a86404a );
 a86408a <=( (not A200)  and  A199 );
 a86411a <=( A203  and  A201 );
 a86412a <=( a86411a  and  a86408a );
 a86413a <=( a86412a  and  a86405a );
 a86417a <=( (not A236)  and  (not A235) );
 a86418a <=( (not A233)  and  a86417a );
 a86421a <=( (not A266)  and  (not A265) );
 a86424a <=( (not A300)  and  A298 );
 a86425a <=( a86424a  and  a86421a );
 a86426a <=( a86425a  and  a86418a );
 a86430a <=( (not A168)  and  (not A169) );
 a86431a <=( (not A170)  and  a86430a );
 a86434a <=( (not A200)  and  A199 );
 a86437a <=( A203  and  A201 );
 a86438a <=( a86437a  and  a86434a );
 a86439a <=( a86438a  and  a86431a );
 a86443a <=( (not A236)  and  (not A235) );
 a86444a <=( (not A233)  and  a86443a );
 a86447a <=( (not A266)  and  (not A265) );
 a86450a <=( A299  and  A298 );
 a86451a <=( a86450a  and  a86447a );
 a86452a <=( a86451a  and  a86444a );
 a86456a <=( (not A168)  and  (not A169) );
 a86457a <=( (not A170)  and  a86456a );
 a86460a <=( (not A200)  and  A199 );
 a86463a <=( A203  and  A201 );
 a86464a <=( a86463a  and  a86460a );
 a86465a <=( a86464a  and  a86457a );
 a86469a <=( (not A236)  and  (not A235) );
 a86470a <=( (not A233)  and  a86469a );
 a86473a <=( (not A266)  and  (not A265) );
 a86476a <=( (not A299)  and  (not A298) );
 a86477a <=( a86476a  and  a86473a );
 a86478a <=( a86477a  and  a86470a );
 a86482a <=( (not A168)  and  (not A169) );
 a86483a <=( (not A170)  and  a86482a );
 a86486a <=( (not A200)  and  A199 );
 a86489a <=( A203  and  A201 );
 a86490a <=( a86489a  and  a86486a );
 a86491a <=( a86490a  and  a86483a );
 a86495a <=( A265  and  (not A234) );
 a86496a <=( (not A233)  and  a86495a );
 a86499a <=( A298  and  A266 );
 a86502a <=( (not A302)  and  (not A301) );
 a86503a <=( a86502a  and  a86499a );
 a86504a <=( a86503a  and  a86496a );
 a86508a <=( (not A168)  and  (not A169) );
 a86509a <=( (not A170)  and  a86508a );
 a86512a <=( (not A200)  and  A199 );
 a86515a <=( A203  and  A201 );
 a86516a <=( a86515a  and  a86512a );
 a86517a <=( a86516a  and  a86509a );
 a86521a <=( (not A266)  and  (not A234) );
 a86522a <=( (not A233)  and  a86521a );
 a86525a <=( (not A269)  and  (not A268) );
 a86528a <=( (not A300)  and  A298 );
 a86529a <=( a86528a  and  a86525a );
 a86530a <=( a86529a  and  a86522a );
 a86534a <=( (not A168)  and  (not A169) );
 a86535a <=( (not A170)  and  a86534a );
 a86538a <=( (not A200)  and  A199 );
 a86541a <=( A203  and  A201 );
 a86542a <=( a86541a  and  a86538a );
 a86543a <=( a86542a  and  a86535a );
 a86547a <=( (not A266)  and  (not A234) );
 a86548a <=( (not A233)  and  a86547a );
 a86551a <=( (not A269)  and  (not A268) );
 a86554a <=( A299  and  A298 );
 a86555a <=( a86554a  and  a86551a );
 a86556a <=( a86555a  and  a86548a );
 a86560a <=( (not A168)  and  (not A169) );
 a86561a <=( (not A170)  and  a86560a );
 a86564a <=( (not A200)  and  A199 );
 a86567a <=( A203  and  A201 );
 a86568a <=( a86567a  and  a86564a );
 a86569a <=( a86568a  and  a86561a );
 a86573a <=( (not A266)  and  (not A234) );
 a86574a <=( (not A233)  and  a86573a );
 a86577a <=( (not A269)  and  (not A268) );
 a86580a <=( (not A299)  and  (not A298) );
 a86581a <=( a86580a  and  a86577a );
 a86582a <=( a86581a  and  a86574a );
 a86586a <=( (not A168)  and  (not A169) );
 a86587a <=( (not A170)  and  a86586a );
 a86590a <=( (not A200)  and  A199 );
 a86593a <=( A203  and  A201 );
 a86594a <=( a86593a  and  a86590a );
 a86595a <=( a86594a  and  a86587a );
 a86599a <=( (not A266)  and  (not A234) );
 a86600a <=( (not A233)  and  a86599a );
 a86603a <=( A298  and  (not A267) );
 a86606a <=( (not A302)  and  (not A301) );
 a86607a <=( a86606a  and  a86603a );
 a86608a <=( a86607a  and  a86600a );
 a86612a <=( (not A168)  and  (not A169) );
 a86613a <=( (not A170)  and  a86612a );
 a86616a <=( (not A200)  and  A199 );
 a86619a <=( A203  and  A201 );
 a86620a <=( a86619a  and  a86616a );
 a86621a <=( a86620a  and  a86613a );
 a86625a <=( (not A265)  and  (not A234) );
 a86626a <=( (not A233)  and  a86625a );
 a86629a <=( A298  and  (not A266) );
 a86632a <=( (not A302)  and  (not A301) );
 a86633a <=( a86632a  and  a86629a );
 a86634a <=( a86633a  and  a86626a );
 a86638a <=( (not A168)  and  (not A169) );
 a86639a <=( (not A170)  and  a86638a );
 a86642a <=( (not A200)  and  A199 );
 a86645a <=( A203  and  A201 );
 a86646a <=( a86645a  and  a86642a );
 a86647a <=( a86646a  and  a86639a );
 a86651a <=( A265  and  (not A233) );
 a86652a <=( (not A232)  and  a86651a );
 a86655a <=( A298  and  A266 );
 a86658a <=( (not A302)  and  (not A301) );
 a86659a <=( a86658a  and  a86655a );
 a86660a <=( a86659a  and  a86652a );
 a86664a <=( (not A168)  and  (not A169) );
 a86665a <=( (not A170)  and  a86664a );
 a86668a <=( (not A200)  and  A199 );
 a86671a <=( A203  and  A201 );
 a86672a <=( a86671a  and  a86668a );
 a86673a <=( a86672a  and  a86665a );
 a86677a <=( (not A266)  and  (not A233) );
 a86678a <=( (not A232)  and  a86677a );
 a86681a <=( (not A269)  and  (not A268) );
 a86684a <=( (not A300)  and  A298 );
 a86685a <=( a86684a  and  a86681a );
 a86686a <=( a86685a  and  a86678a );
 a86690a <=( (not A168)  and  (not A169) );
 a86691a <=( (not A170)  and  a86690a );
 a86694a <=( (not A200)  and  A199 );
 a86697a <=( A203  and  A201 );
 a86698a <=( a86697a  and  a86694a );
 a86699a <=( a86698a  and  a86691a );
 a86703a <=( (not A266)  and  (not A233) );
 a86704a <=( (not A232)  and  a86703a );
 a86707a <=( (not A269)  and  (not A268) );
 a86710a <=( A299  and  A298 );
 a86711a <=( a86710a  and  a86707a );
 a86712a <=( a86711a  and  a86704a );
 a86716a <=( (not A168)  and  (not A169) );
 a86717a <=( (not A170)  and  a86716a );
 a86720a <=( (not A200)  and  A199 );
 a86723a <=( A203  and  A201 );
 a86724a <=( a86723a  and  a86720a );
 a86725a <=( a86724a  and  a86717a );
 a86729a <=( (not A266)  and  (not A233) );
 a86730a <=( (not A232)  and  a86729a );
 a86733a <=( (not A269)  and  (not A268) );
 a86736a <=( (not A299)  and  (not A298) );
 a86737a <=( a86736a  and  a86733a );
 a86738a <=( a86737a  and  a86730a );
 a86742a <=( (not A168)  and  (not A169) );
 a86743a <=( (not A170)  and  a86742a );
 a86746a <=( (not A200)  and  A199 );
 a86749a <=( A203  and  A201 );
 a86750a <=( a86749a  and  a86746a );
 a86751a <=( a86750a  and  a86743a );
 a86755a <=( (not A266)  and  (not A233) );
 a86756a <=( (not A232)  and  a86755a );
 a86759a <=( A298  and  (not A267) );
 a86762a <=( (not A302)  and  (not A301) );
 a86763a <=( a86762a  and  a86759a );
 a86764a <=( a86763a  and  a86756a );
 a86768a <=( (not A168)  and  (not A169) );
 a86769a <=( (not A170)  and  a86768a );
 a86772a <=( (not A200)  and  A199 );
 a86775a <=( A203  and  A201 );
 a86776a <=( a86775a  and  a86772a );
 a86777a <=( a86776a  and  a86769a );
 a86781a <=( (not A265)  and  (not A233) );
 a86782a <=( (not A232)  and  a86781a );
 a86785a <=( A298  and  (not A266) );
 a86788a <=( (not A302)  and  (not A301) );
 a86789a <=( a86788a  and  a86785a );
 a86790a <=( a86789a  and  a86782a );
 a86794a <=( (not A166)  and  (not A167) );
 a86795a <=( A170  and  a86794a );
 a86798a <=( (not A200)  and  A199 );
 a86801a <=( A202  and  A201 );
 a86802a <=( a86801a  and  a86798a );
 a86803a <=( a86802a  and  a86795a );
 a86806a <=( A233  and  A232 );
 a86809a <=( (not A268)  and  A265 );
 a86810a <=( a86809a  and  a86806a );
 a86813a <=( (not A299)  and  (not A269) );
 a86816a <=( (not A302)  and  (not A301) );
 a86817a <=( a86816a  and  a86813a );
 a86818a <=( a86817a  and  a86810a );
 a86822a <=( (not A166)  and  (not A167) );
 a86823a <=( A170  and  a86822a );
 a86826a <=( (not A200)  and  A199 );
 a86829a <=( A202  and  A201 );
 a86830a <=( a86829a  and  a86826a );
 a86831a <=( a86830a  and  a86823a );
 a86834a <=( (not A235)  and  (not A233) );
 a86837a <=( A265  and  (not A236) );
 a86838a <=( a86837a  and  a86834a );
 a86841a <=( A298  and  A266 );
 a86844a <=( (not A302)  and  (not A301) );
 a86845a <=( a86844a  and  a86841a );
 a86846a <=( a86845a  and  a86838a );
 a86850a <=( (not A166)  and  (not A167) );
 a86851a <=( A170  and  a86850a );
 a86854a <=( (not A200)  and  A199 );
 a86857a <=( A202  and  A201 );
 a86858a <=( a86857a  and  a86854a );
 a86859a <=( a86858a  and  a86851a );
 a86862a <=( (not A235)  and  (not A233) );
 a86865a <=( (not A266)  and  (not A236) );
 a86866a <=( a86865a  and  a86862a );
 a86869a <=( (not A269)  and  (not A268) );
 a86872a <=( (not A300)  and  A298 );
 a86873a <=( a86872a  and  a86869a );
 a86874a <=( a86873a  and  a86866a );
 a86878a <=( (not A166)  and  (not A167) );
 a86879a <=( A170  and  a86878a );
 a86882a <=( (not A200)  and  A199 );
 a86885a <=( A202  and  A201 );
 a86886a <=( a86885a  and  a86882a );
 a86887a <=( a86886a  and  a86879a );
 a86890a <=( (not A235)  and  (not A233) );
 a86893a <=( (not A266)  and  (not A236) );
 a86894a <=( a86893a  and  a86890a );
 a86897a <=( (not A269)  and  (not A268) );
 a86900a <=( A299  and  A298 );
 a86901a <=( a86900a  and  a86897a );
 a86902a <=( a86901a  and  a86894a );
 a86906a <=( (not A166)  and  (not A167) );
 a86907a <=( A170  and  a86906a );
 a86910a <=( (not A200)  and  A199 );
 a86913a <=( A202  and  A201 );
 a86914a <=( a86913a  and  a86910a );
 a86915a <=( a86914a  and  a86907a );
 a86918a <=( (not A235)  and  (not A233) );
 a86921a <=( (not A266)  and  (not A236) );
 a86922a <=( a86921a  and  a86918a );
 a86925a <=( (not A269)  and  (not A268) );
 a86928a <=( (not A299)  and  (not A298) );
 a86929a <=( a86928a  and  a86925a );
 a86930a <=( a86929a  and  a86922a );
 a86934a <=( (not A166)  and  (not A167) );
 a86935a <=( A170  and  a86934a );
 a86938a <=( (not A200)  and  A199 );
 a86941a <=( A202  and  A201 );
 a86942a <=( a86941a  and  a86938a );
 a86943a <=( a86942a  and  a86935a );
 a86946a <=( (not A235)  and  (not A233) );
 a86949a <=( (not A266)  and  (not A236) );
 a86950a <=( a86949a  and  a86946a );
 a86953a <=( A298  and  (not A267) );
 a86956a <=( (not A302)  and  (not A301) );
 a86957a <=( a86956a  and  a86953a );
 a86958a <=( a86957a  and  a86950a );
 a86962a <=( (not A166)  and  (not A167) );
 a86963a <=( A170  and  a86962a );
 a86966a <=( (not A200)  and  A199 );
 a86969a <=( A202  and  A201 );
 a86970a <=( a86969a  and  a86966a );
 a86971a <=( a86970a  and  a86963a );
 a86974a <=( (not A235)  and  (not A233) );
 a86977a <=( (not A265)  and  (not A236) );
 a86978a <=( a86977a  and  a86974a );
 a86981a <=( A298  and  (not A266) );
 a86984a <=( (not A302)  and  (not A301) );
 a86985a <=( a86984a  and  a86981a );
 a86986a <=( a86985a  and  a86978a );
 a86990a <=( (not A166)  and  (not A167) );
 a86991a <=( A170  and  a86990a );
 a86994a <=( (not A200)  and  A199 );
 a86997a <=( A202  and  A201 );
 a86998a <=( a86997a  and  a86994a );
 a86999a <=( a86998a  and  a86991a );
 a87002a <=( (not A234)  and  (not A233) );
 a87005a <=( (not A268)  and  (not A266) );
 a87006a <=( a87005a  and  a87002a );
 a87009a <=( A298  and  (not A269) );
 a87012a <=( (not A302)  and  (not A301) );
 a87013a <=( a87012a  and  a87009a );
 a87014a <=( a87013a  and  a87006a );
 a87018a <=( (not A166)  and  (not A167) );
 a87019a <=( A170  and  a87018a );
 a87022a <=( (not A200)  and  A199 );
 a87025a <=( A202  and  A201 );
 a87026a <=( a87025a  and  a87022a );
 a87027a <=( a87026a  and  a87019a );
 a87030a <=( (not A233)  and  A232 );
 a87033a <=( A235  and  A234 );
 a87034a <=( a87033a  and  a87030a );
 a87037a <=( (not A299)  and  A298 );
 a87040a <=( A301  and  A300 );
 a87041a <=( a87040a  and  a87037a );
 a87042a <=( a87041a  and  a87034a );
 a87046a <=( (not A166)  and  (not A167) );
 a87047a <=( A170  and  a87046a );
 a87050a <=( (not A200)  and  A199 );
 a87053a <=( A202  and  A201 );
 a87054a <=( a87053a  and  a87050a );
 a87055a <=( a87054a  and  a87047a );
 a87058a <=( (not A233)  and  A232 );
 a87061a <=( A235  and  A234 );
 a87062a <=( a87061a  and  a87058a );
 a87065a <=( (not A299)  and  A298 );
 a87068a <=( A302  and  A300 );
 a87069a <=( a87068a  and  a87065a );
 a87070a <=( a87069a  and  a87062a );
 a87074a <=( (not A166)  and  (not A167) );
 a87075a <=( A170  and  a87074a );
 a87078a <=( (not A200)  and  A199 );
 a87081a <=( A202  and  A201 );
 a87082a <=( a87081a  and  a87078a );
 a87083a <=( a87082a  and  a87075a );
 a87086a <=( (not A233)  and  A232 );
 a87089a <=( A235  and  A234 );
 a87090a <=( a87089a  and  a87086a );
 a87093a <=( (not A266)  and  A265 );
 a87096a <=( A268  and  A267 );
 a87097a <=( a87096a  and  a87093a );
 a87098a <=( a87097a  and  a87090a );
 a87102a <=( (not A166)  and  (not A167) );
 a87103a <=( A170  and  a87102a );
 a87106a <=( (not A200)  and  A199 );
 a87109a <=( A202  and  A201 );
 a87110a <=( a87109a  and  a87106a );
 a87111a <=( a87110a  and  a87103a );
 a87114a <=( (not A233)  and  A232 );
 a87117a <=( A235  and  A234 );
 a87118a <=( a87117a  and  a87114a );
 a87121a <=( (not A266)  and  A265 );
 a87124a <=( A269  and  A267 );
 a87125a <=( a87124a  and  a87121a );
 a87126a <=( a87125a  and  a87118a );
 a87130a <=( (not A166)  and  (not A167) );
 a87131a <=( A170  and  a87130a );
 a87134a <=( (not A200)  and  A199 );
 a87137a <=( A202  and  A201 );
 a87138a <=( a87137a  and  a87134a );
 a87139a <=( a87138a  and  a87131a );
 a87142a <=( (not A233)  and  A232 );
 a87145a <=( A236  and  A234 );
 a87146a <=( a87145a  and  a87142a );
 a87149a <=( (not A299)  and  A298 );
 a87152a <=( A301  and  A300 );
 a87153a <=( a87152a  and  a87149a );
 a87154a <=( a87153a  and  a87146a );
 a87158a <=( (not A166)  and  (not A167) );
 a87159a <=( A170  and  a87158a );
 a87162a <=( (not A200)  and  A199 );
 a87165a <=( A202  and  A201 );
 a87166a <=( a87165a  and  a87162a );
 a87167a <=( a87166a  and  a87159a );
 a87170a <=( (not A233)  and  A232 );
 a87173a <=( A236  and  A234 );
 a87174a <=( a87173a  and  a87170a );
 a87177a <=( (not A299)  and  A298 );
 a87180a <=( A302  and  A300 );
 a87181a <=( a87180a  and  a87177a );
 a87182a <=( a87181a  and  a87174a );
 a87186a <=( (not A166)  and  (not A167) );
 a87187a <=( A170  and  a87186a );
 a87190a <=( (not A200)  and  A199 );
 a87193a <=( A202  and  A201 );
 a87194a <=( a87193a  and  a87190a );
 a87195a <=( a87194a  and  a87187a );
 a87198a <=( (not A233)  and  A232 );
 a87201a <=( A236  and  A234 );
 a87202a <=( a87201a  and  a87198a );
 a87205a <=( (not A266)  and  A265 );
 a87208a <=( A268  and  A267 );
 a87209a <=( a87208a  and  a87205a );
 a87210a <=( a87209a  and  a87202a );
 a87214a <=( (not A166)  and  (not A167) );
 a87215a <=( A170  and  a87214a );
 a87218a <=( (not A200)  and  A199 );
 a87221a <=( A202  and  A201 );
 a87222a <=( a87221a  and  a87218a );
 a87223a <=( a87222a  and  a87215a );
 a87226a <=( (not A233)  and  A232 );
 a87229a <=( A236  and  A234 );
 a87230a <=( a87229a  and  a87226a );
 a87233a <=( (not A266)  and  A265 );
 a87236a <=( A269  and  A267 );
 a87237a <=( a87236a  and  a87233a );
 a87238a <=( a87237a  and  a87230a );
 a87242a <=( (not A166)  and  (not A167) );
 a87243a <=( A170  and  a87242a );
 a87246a <=( (not A200)  and  A199 );
 a87249a <=( A202  and  A201 );
 a87250a <=( a87249a  and  a87246a );
 a87251a <=( a87250a  and  a87243a );
 a87254a <=( (not A233)  and  (not A232) );
 a87257a <=( (not A268)  and  (not A266) );
 a87258a <=( a87257a  and  a87254a );
 a87261a <=( A298  and  (not A269) );
 a87264a <=( (not A302)  and  (not A301) );
 a87265a <=( a87264a  and  a87261a );
 a87266a <=( a87265a  and  a87258a );
 a87270a <=( (not A166)  and  (not A167) );
 a87271a <=( A170  and  a87270a );
 a87274a <=( (not A200)  and  A199 );
 a87277a <=( A203  and  A201 );
 a87278a <=( a87277a  and  a87274a );
 a87279a <=( a87278a  and  a87271a );
 a87282a <=( A233  and  A232 );
 a87285a <=( (not A268)  and  A265 );
 a87286a <=( a87285a  and  a87282a );
 a87289a <=( (not A299)  and  (not A269) );
 a87292a <=( (not A302)  and  (not A301) );
 a87293a <=( a87292a  and  a87289a );
 a87294a <=( a87293a  and  a87286a );
 a87298a <=( (not A166)  and  (not A167) );
 a87299a <=( A170  and  a87298a );
 a87302a <=( (not A200)  and  A199 );
 a87305a <=( A203  and  A201 );
 a87306a <=( a87305a  and  a87302a );
 a87307a <=( a87306a  and  a87299a );
 a87310a <=( (not A235)  and  (not A233) );
 a87313a <=( A265  and  (not A236) );
 a87314a <=( a87313a  and  a87310a );
 a87317a <=( A298  and  A266 );
 a87320a <=( (not A302)  and  (not A301) );
 a87321a <=( a87320a  and  a87317a );
 a87322a <=( a87321a  and  a87314a );
 a87326a <=( (not A166)  and  (not A167) );
 a87327a <=( A170  and  a87326a );
 a87330a <=( (not A200)  and  A199 );
 a87333a <=( A203  and  A201 );
 a87334a <=( a87333a  and  a87330a );
 a87335a <=( a87334a  and  a87327a );
 a87338a <=( (not A235)  and  (not A233) );
 a87341a <=( (not A266)  and  (not A236) );
 a87342a <=( a87341a  and  a87338a );
 a87345a <=( (not A269)  and  (not A268) );
 a87348a <=( (not A300)  and  A298 );
 a87349a <=( a87348a  and  a87345a );
 a87350a <=( a87349a  and  a87342a );
 a87354a <=( (not A166)  and  (not A167) );
 a87355a <=( A170  and  a87354a );
 a87358a <=( (not A200)  and  A199 );
 a87361a <=( A203  and  A201 );
 a87362a <=( a87361a  and  a87358a );
 a87363a <=( a87362a  and  a87355a );
 a87366a <=( (not A235)  and  (not A233) );
 a87369a <=( (not A266)  and  (not A236) );
 a87370a <=( a87369a  and  a87366a );
 a87373a <=( (not A269)  and  (not A268) );
 a87376a <=( A299  and  A298 );
 a87377a <=( a87376a  and  a87373a );
 a87378a <=( a87377a  and  a87370a );
 a87382a <=( (not A166)  and  (not A167) );
 a87383a <=( A170  and  a87382a );
 a87386a <=( (not A200)  and  A199 );
 a87389a <=( A203  and  A201 );
 a87390a <=( a87389a  and  a87386a );
 a87391a <=( a87390a  and  a87383a );
 a87394a <=( (not A235)  and  (not A233) );
 a87397a <=( (not A266)  and  (not A236) );
 a87398a <=( a87397a  and  a87394a );
 a87401a <=( (not A269)  and  (not A268) );
 a87404a <=( (not A299)  and  (not A298) );
 a87405a <=( a87404a  and  a87401a );
 a87406a <=( a87405a  and  a87398a );
 a87410a <=( (not A166)  and  (not A167) );
 a87411a <=( A170  and  a87410a );
 a87414a <=( (not A200)  and  A199 );
 a87417a <=( A203  and  A201 );
 a87418a <=( a87417a  and  a87414a );
 a87419a <=( a87418a  and  a87411a );
 a87422a <=( (not A235)  and  (not A233) );
 a87425a <=( (not A266)  and  (not A236) );
 a87426a <=( a87425a  and  a87422a );
 a87429a <=( A298  and  (not A267) );
 a87432a <=( (not A302)  and  (not A301) );
 a87433a <=( a87432a  and  a87429a );
 a87434a <=( a87433a  and  a87426a );
 a87438a <=( (not A166)  and  (not A167) );
 a87439a <=( A170  and  a87438a );
 a87442a <=( (not A200)  and  A199 );
 a87445a <=( A203  and  A201 );
 a87446a <=( a87445a  and  a87442a );
 a87447a <=( a87446a  and  a87439a );
 a87450a <=( (not A235)  and  (not A233) );
 a87453a <=( (not A265)  and  (not A236) );
 a87454a <=( a87453a  and  a87450a );
 a87457a <=( A298  and  (not A266) );
 a87460a <=( (not A302)  and  (not A301) );
 a87461a <=( a87460a  and  a87457a );
 a87462a <=( a87461a  and  a87454a );
 a87466a <=( (not A166)  and  (not A167) );
 a87467a <=( A170  and  a87466a );
 a87470a <=( (not A200)  and  A199 );
 a87473a <=( A203  and  A201 );
 a87474a <=( a87473a  and  a87470a );
 a87475a <=( a87474a  and  a87467a );
 a87478a <=( (not A234)  and  (not A233) );
 a87481a <=( (not A268)  and  (not A266) );
 a87482a <=( a87481a  and  a87478a );
 a87485a <=( A298  and  (not A269) );
 a87488a <=( (not A302)  and  (not A301) );
 a87489a <=( a87488a  and  a87485a );
 a87490a <=( a87489a  and  a87482a );
 a87494a <=( (not A166)  and  (not A167) );
 a87495a <=( A170  and  a87494a );
 a87498a <=( (not A200)  and  A199 );
 a87501a <=( A203  and  A201 );
 a87502a <=( a87501a  and  a87498a );
 a87503a <=( a87502a  and  a87495a );
 a87506a <=( (not A233)  and  A232 );
 a87509a <=( A235  and  A234 );
 a87510a <=( a87509a  and  a87506a );
 a87513a <=( (not A299)  and  A298 );
 a87516a <=( A301  and  A300 );
 a87517a <=( a87516a  and  a87513a );
 a87518a <=( a87517a  and  a87510a );
 a87522a <=( (not A166)  and  (not A167) );
 a87523a <=( A170  and  a87522a );
 a87526a <=( (not A200)  and  A199 );
 a87529a <=( A203  and  A201 );
 a87530a <=( a87529a  and  a87526a );
 a87531a <=( a87530a  and  a87523a );
 a87534a <=( (not A233)  and  A232 );
 a87537a <=( A235  and  A234 );
 a87538a <=( a87537a  and  a87534a );
 a87541a <=( (not A299)  and  A298 );
 a87544a <=( A302  and  A300 );
 a87545a <=( a87544a  and  a87541a );
 a87546a <=( a87545a  and  a87538a );
 a87550a <=( (not A166)  and  (not A167) );
 a87551a <=( A170  and  a87550a );
 a87554a <=( (not A200)  and  A199 );
 a87557a <=( A203  and  A201 );
 a87558a <=( a87557a  and  a87554a );
 a87559a <=( a87558a  and  a87551a );
 a87562a <=( (not A233)  and  A232 );
 a87565a <=( A235  and  A234 );
 a87566a <=( a87565a  and  a87562a );
 a87569a <=( (not A266)  and  A265 );
 a87572a <=( A268  and  A267 );
 a87573a <=( a87572a  and  a87569a );
 a87574a <=( a87573a  and  a87566a );
 a87578a <=( (not A166)  and  (not A167) );
 a87579a <=( A170  and  a87578a );
 a87582a <=( (not A200)  and  A199 );
 a87585a <=( A203  and  A201 );
 a87586a <=( a87585a  and  a87582a );
 a87587a <=( a87586a  and  a87579a );
 a87590a <=( (not A233)  and  A232 );
 a87593a <=( A235  and  A234 );
 a87594a <=( a87593a  and  a87590a );
 a87597a <=( (not A266)  and  A265 );
 a87600a <=( A269  and  A267 );
 a87601a <=( a87600a  and  a87597a );
 a87602a <=( a87601a  and  a87594a );
 a87606a <=( (not A166)  and  (not A167) );
 a87607a <=( A170  and  a87606a );
 a87610a <=( (not A200)  and  A199 );
 a87613a <=( A203  and  A201 );
 a87614a <=( a87613a  and  a87610a );
 a87615a <=( a87614a  and  a87607a );
 a87618a <=( (not A233)  and  A232 );
 a87621a <=( A236  and  A234 );
 a87622a <=( a87621a  and  a87618a );
 a87625a <=( (not A299)  and  A298 );
 a87628a <=( A301  and  A300 );
 a87629a <=( a87628a  and  a87625a );
 a87630a <=( a87629a  and  a87622a );
 a87634a <=( (not A166)  and  (not A167) );
 a87635a <=( A170  and  a87634a );
 a87638a <=( (not A200)  and  A199 );
 a87641a <=( A203  and  A201 );
 a87642a <=( a87641a  and  a87638a );
 a87643a <=( a87642a  and  a87635a );
 a87646a <=( (not A233)  and  A232 );
 a87649a <=( A236  and  A234 );
 a87650a <=( a87649a  and  a87646a );
 a87653a <=( (not A299)  and  A298 );
 a87656a <=( A302  and  A300 );
 a87657a <=( a87656a  and  a87653a );
 a87658a <=( a87657a  and  a87650a );
 a87662a <=( (not A166)  and  (not A167) );
 a87663a <=( A170  and  a87662a );
 a87666a <=( (not A200)  and  A199 );
 a87669a <=( A203  and  A201 );
 a87670a <=( a87669a  and  a87666a );
 a87671a <=( a87670a  and  a87663a );
 a87674a <=( (not A233)  and  A232 );
 a87677a <=( A236  and  A234 );
 a87678a <=( a87677a  and  a87674a );
 a87681a <=( (not A266)  and  A265 );
 a87684a <=( A268  and  A267 );
 a87685a <=( a87684a  and  a87681a );
 a87686a <=( a87685a  and  a87678a );
 a87690a <=( (not A166)  and  (not A167) );
 a87691a <=( A170  and  a87690a );
 a87694a <=( (not A200)  and  A199 );
 a87697a <=( A203  and  A201 );
 a87698a <=( a87697a  and  a87694a );
 a87699a <=( a87698a  and  a87691a );
 a87702a <=( (not A233)  and  A232 );
 a87705a <=( A236  and  A234 );
 a87706a <=( a87705a  and  a87702a );
 a87709a <=( (not A266)  and  A265 );
 a87712a <=( A269  and  A267 );
 a87713a <=( a87712a  and  a87709a );
 a87714a <=( a87713a  and  a87706a );
 a87718a <=( (not A166)  and  (not A167) );
 a87719a <=( A170  and  a87718a );
 a87722a <=( (not A200)  and  A199 );
 a87725a <=( A203  and  A201 );
 a87726a <=( a87725a  and  a87722a );
 a87727a <=( a87726a  and  a87719a );
 a87730a <=( (not A233)  and  (not A232) );
 a87733a <=( (not A268)  and  (not A266) );
 a87734a <=( a87733a  and  a87730a );
 a87737a <=( A298  and  (not A269) );
 a87740a <=( (not A302)  and  (not A301) );
 a87741a <=( a87740a  and  a87737a );
 a87742a <=( a87741a  and  a87734a );
 a87746a <=( A167  and  (not A168) );
 a87747a <=( A170  and  a87746a );
 a87750a <=( (not A199)  and  A166 );
 a87753a <=( (not A233)  and  A200 );
 a87754a <=( a87753a  and  a87750a );
 a87755a <=( a87754a  and  a87747a );
 a87758a <=( (not A236)  and  (not A235) );
 a87761a <=( (not A268)  and  (not A266) );
 a87762a <=( a87761a  and  a87758a );
 a87765a <=( A298  and  (not A269) );
 a87768a <=( (not A302)  and  (not A301) );
 a87769a <=( a87768a  and  a87765a );
 a87770a <=( a87769a  and  a87762a );
 a87774a <=( A167  and  (not A168) );
 a87775a <=( (not A170)  and  a87774a );
 a87778a <=( (not A199)  and  (not A166) );
 a87781a <=( (not A233)  and  A200 );
 a87782a <=( a87781a  and  a87778a );
 a87783a <=( a87782a  and  a87775a );
 a87786a <=( (not A236)  and  (not A235) );
 a87789a <=( (not A268)  and  (not A266) );
 a87790a <=( a87789a  and  a87786a );
 a87793a <=( A298  and  (not A269) );
 a87796a <=( (not A302)  and  (not A301) );
 a87797a <=( a87796a  and  a87793a );
 a87798a <=( a87797a  and  a87790a );
 a87802a <=( (not A167)  and  (not A168) );
 a87803a <=( (not A170)  and  a87802a );
 a87806a <=( (not A199)  and  A166 );
 a87809a <=( (not A233)  and  A200 );
 a87810a <=( a87809a  and  a87806a );
 a87811a <=( a87810a  and  a87803a );
 a87814a <=( (not A236)  and  (not A235) );
 a87817a <=( (not A268)  and  (not A266) );
 a87818a <=( a87817a  and  a87814a );
 a87821a <=( A298  and  (not A269) );
 a87824a <=( (not A302)  and  (not A301) );
 a87825a <=( a87824a  and  a87821a );
 a87826a <=( a87825a  and  a87818a );
 a87830a <=( A167  and  (not A168) );
 a87831a <=( A169  and  a87830a );
 a87834a <=( (not A199)  and  (not A166) );
 a87837a <=( (not A233)  and  A200 );
 a87838a <=( a87837a  and  a87834a );
 a87839a <=( a87838a  and  a87831a );
 a87842a <=( (not A236)  and  (not A235) );
 a87845a <=( (not A268)  and  (not A266) );
 a87846a <=( a87845a  and  a87842a );
 a87849a <=( A298  and  (not A269) );
 a87852a <=( (not A302)  and  (not A301) );
 a87853a <=( a87852a  and  a87849a );
 a87854a <=( a87853a  and  a87846a );
 a87858a <=( A167  and  (not A168) );
 a87859a <=( A169  and  a87858a );
 a87862a <=( A199  and  (not A166) );
 a87865a <=( A201  and  (not A200) );
 a87866a <=( a87865a  and  a87862a );
 a87867a <=( a87866a  and  a87859a );
 a87870a <=( A232  and  A202 );
 a87873a <=( A265  and  A233 );
 a87874a <=( a87873a  and  a87870a );
 a87877a <=( (not A269)  and  (not A268) );
 a87880a <=( (not A300)  and  (not A299) );
 a87881a <=( a87880a  and  a87877a );
 a87882a <=( a87881a  and  a87874a );
 a87886a <=( A167  and  (not A168) );
 a87887a <=( A169  and  a87886a );
 a87890a <=( A199  and  (not A166) );
 a87893a <=( A201  and  (not A200) );
 a87894a <=( a87893a  and  a87890a );
 a87895a <=( a87894a  and  a87887a );
 a87898a <=( A232  and  A202 );
 a87901a <=( A265  and  A233 );
 a87902a <=( a87901a  and  a87898a );
 a87905a <=( (not A269)  and  (not A268) );
 a87908a <=( A299  and  A298 );
 a87909a <=( a87908a  and  a87905a );
 a87910a <=( a87909a  and  a87902a );
 a87914a <=( A167  and  (not A168) );
 a87915a <=( A169  and  a87914a );
 a87918a <=( A199  and  (not A166) );
 a87921a <=( A201  and  (not A200) );
 a87922a <=( a87921a  and  a87918a );
 a87923a <=( a87922a  and  a87915a );
 a87926a <=( A232  and  A202 );
 a87929a <=( A265  and  A233 );
 a87930a <=( a87929a  and  a87926a );
 a87933a <=( (not A269)  and  (not A268) );
 a87936a <=( (not A299)  and  (not A298) );
 a87937a <=( a87936a  and  a87933a );
 a87938a <=( a87937a  and  a87930a );
 a87942a <=( A167  and  (not A168) );
 a87943a <=( A169  and  a87942a );
 a87946a <=( A199  and  (not A166) );
 a87949a <=( A201  and  (not A200) );
 a87950a <=( a87949a  and  a87946a );
 a87951a <=( a87950a  and  a87943a );
 a87954a <=( A232  and  A202 );
 a87957a <=( A265  and  A233 );
 a87958a <=( a87957a  and  a87954a );
 a87961a <=( (not A299)  and  (not A267) );
 a87964a <=( (not A302)  and  (not A301) );
 a87965a <=( a87964a  and  a87961a );
 a87966a <=( a87965a  and  a87958a );
 a87970a <=( A167  and  (not A168) );
 a87971a <=( A169  and  a87970a );
 a87974a <=( A199  and  (not A166) );
 a87977a <=( A201  and  (not A200) );
 a87978a <=( a87977a  and  a87974a );
 a87979a <=( a87978a  and  a87971a );
 a87982a <=( A232  and  A202 );
 a87985a <=( A265  and  A233 );
 a87986a <=( a87985a  and  a87982a );
 a87989a <=( (not A299)  and  A266 );
 a87992a <=( (not A302)  and  (not A301) );
 a87993a <=( a87992a  and  a87989a );
 a87994a <=( a87993a  and  a87986a );
 a87998a <=( A167  and  (not A168) );
 a87999a <=( A169  and  a87998a );
 a88002a <=( A199  and  (not A166) );
 a88005a <=( A201  and  (not A200) );
 a88006a <=( a88005a  and  a88002a );
 a88007a <=( a88006a  and  a87999a );
 a88010a <=( A232  and  A202 );
 a88013a <=( (not A265)  and  A233 );
 a88014a <=( a88013a  and  a88010a );
 a88017a <=( (not A299)  and  (not A266) );
 a88020a <=( (not A302)  and  (not A301) );
 a88021a <=( a88020a  and  a88017a );
 a88022a <=( a88021a  and  a88014a );
 a88026a <=( A167  and  (not A168) );
 a88027a <=( A169  and  a88026a );
 a88030a <=( A199  and  (not A166) );
 a88033a <=( A201  and  (not A200) );
 a88034a <=( a88033a  and  a88030a );
 a88035a <=( a88034a  and  a88027a );
 a88038a <=( (not A233)  and  A202 );
 a88041a <=( (not A236)  and  (not A235) );
 a88042a <=( a88041a  and  a88038a );
 a88045a <=( A266  and  A265 );
 a88048a <=( (not A300)  and  A298 );
 a88049a <=( a88048a  and  a88045a );
 a88050a <=( a88049a  and  a88042a );
 a88054a <=( A167  and  (not A168) );
 a88055a <=( A169  and  a88054a );
 a88058a <=( A199  and  (not A166) );
 a88061a <=( A201  and  (not A200) );
 a88062a <=( a88061a  and  a88058a );
 a88063a <=( a88062a  and  a88055a );
 a88066a <=( (not A233)  and  A202 );
 a88069a <=( (not A236)  and  (not A235) );
 a88070a <=( a88069a  and  a88066a );
 a88073a <=( A266  and  A265 );
 a88076a <=( A299  and  A298 );
 a88077a <=( a88076a  and  a88073a );
 a88078a <=( a88077a  and  a88070a );
 a88082a <=( A167  and  (not A168) );
 a88083a <=( A169  and  a88082a );
 a88086a <=( A199  and  (not A166) );
 a88089a <=( A201  and  (not A200) );
 a88090a <=( a88089a  and  a88086a );
 a88091a <=( a88090a  and  a88083a );
 a88094a <=( (not A233)  and  A202 );
 a88097a <=( (not A236)  and  (not A235) );
 a88098a <=( a88097a  and  a88094a );
 a88101a <=( A266  and  A265 );
 a88104a <=( (not A299)  and  (not A298) );
 a88105a <=( a88104a  and  a88101a );
 a88106a <=( a88105a  and  a88098a );
 a88110a <=( A167  and  (not A168) );
 a88111a <=( A169  and  a88110a );
 a88114a <=( A199  and  (not A166) );
 a88117a <=( A201  and  (not A200) );
 a88118a <=( a88117a  and  a88114a );
 a88119a <=( a88118a  and  a88111a );
 a88122a <=( (not A233)  and  A202 );
 a88125a <=( (not A236)  and  (not A235) );
 a88126a <=( a88125a  and  a88122a );
 a88129a <=( (not A267)  and  (not A266) );
 a88132a <=( (not A300)  and  A298 );
 a88133a <=( a88132a  and  a88129a );
 a88134a <=( a88133a  and  a88126a );
 a88138a <=( A167  and  (not A168) );
 a88139a <=( A169  and  a88138a );
 a88142a <=( A199  and  (not A166) );
 a88145a <=( A201  and  (not A200) );
 a88146a <=( a88145a  and  a88142a );
 a88147a <=( a88146a  and  a88139a );
 a88150a <=( (not A233)  and  A202 );
 a88153a <=( (not A236)  and  (not A235) );
 a88154a <=( a88153a  and  a88150a );
 a88157a <=( (not A267)  and  (not A266) );
 a88160a <=( A299  and  A298 );
 a88161a <=( a88160a  and  a88157a );
 a88162a <=( a88161a  and  a88154a );
 a88166a <=( A167  and  (not A168) );
 a88167a <=( A169  and  a88166a );
 a88170a <=( A199  and  (not A166) );
 a88173a <=( A201  and  (not A200) );
 a88174a <=( a88173a  and  a88170a );
 a88175a <=( a88174a  and  a88167a );
 a88178a <=( (not A233)  and  A202 );
 a88181a <=( (not A236)  and  (not A235) );
 a88182a <=( a88181a  and  a88178a );
 a88185a <=( (not A267)  and  (not A266) );
 a88188a <=( (not A299)  and  (not A298) );
 a88189a <=( a88188a  and  a88185a );
 a88190a <=( a88189a  and  a88182a );
 a88194a <=( A167  and  (not A168) );
 a88195a <=( A169  and  a88194a );
 a88198a <=( A199  and  (not A166) );
 a88201a <=( A201  and  (not A200) );
 a88202a <=( a88201a  and  a88198a );
 a88203a <=( a88202a  and  a88195a );
 a88206a <=( (not A233)  and  A202 );
 a88209a <=( (not A236)  and  (not A235) );
 a88210a <=( a88209a  and  a88206a );
 a88213a <=( (not A266)  and  (not A265) );
 a88216a <=( (not A300)  and  A298 );
 a88217a <=( a88216a  and  a88213a );
 a88218a <=( a88217a  and  a88210a );
 a88222a <=( A167  and  (not A168) );
 a88223a <=( A169  and  a88222a );
 a88226a <=( A199  and  (not A166) );
 a88229a <=( A201  and  (not A200) );
 a88230a <=( a88229a  and  a88226a );
 a88231a <=( a88230a  and  a88223a );
 a88234a <=( (not A233)  and  A202 );
 a88237a <=( (not A236)  and  (not A235) );
 a88238a <=( a88237a  and  a88234a );
 a88241a <=( (not A266)  and  (not A265) );
 a88244a <=( A299  and  A298 );
 a88245a <=( a88244a  and  a88241a );
 a88246a <=( a88245a  and  a88238a );
 a88250a <=( A167  and  (not A168) );
 a88251a <=( A169  and  a88250a );
 a88254a <=( A199  and  (not A166) );
 a88257a <=( A201  and  (not A200) );
 a88258a <=( a88257a  and  a88254a );
 a88259a <=( a88258a  and  a88251a );
 a88262a <=( (not A233)  and  A202 );
 a88265a <=( (not A236)  and  (not A235) );
 a88266a <=( a88265a  and  a88262a );
 a88269a <=( (not A266)  and  (not A265) );
 a88272a <=( (not A299)  and  (not A298) );
 a88273a <=( a88272a  and  a88269a );
 a88274a <=( a88273a  and  a88266a );
 a88278a <=( A167  and  (not A168) );
 a88279a <=( A169  and  a88278a );
 a88282a <=( A199  and  (not A166) );
 a88285a <=( A201  and  (not A200) );
 a88286a <=( a88285a  and  a88282a );
 a88287a <=( a88286a  and  a88279a );
 a88290a <=( (not A233)  and  A202 );
 a88293a <=( A265  and  (not A234) );
 a88294a <=( a88293a  and  a88290a );
 a88297a <=( A298  and  A266 );
 a88300a <=( (not A302)  and  (not A301) );
 a88301a <=( a88300a  and  a88297a );
 a88302a <=( a88301a  and  a88294a );
 a88306a <=( A167  and  (not A168) );
 a88307a <=( A169  and  a88306a );
 a88310a <=( A199  and  (not A166) );
 a88313a <=( A201  and  (not A200) );
 a88314a <=( a88313a  and  a88310a );
 a88315a <=( a88314a  and  a88307a );
 a88318a <=( (not A233)  and  A202 );
 a88321a <=( (not A266)  and  (not A234) );
 a88322a <=( a88321a  and  a88318a );
 a88325a <=( (not A269)  and  (not A268) );
 a88328a <=( (not A300)  and  A298 );
 a88329a <=( a88328a  and  a88325a );
 a88330a <=( a88329a  and  a88322a );
 a88334a <=( A167  and  (not A168) );
 a88335a <=( A169  and  a88334a );
 a88338a <=( A199  and  (not A166) );
 a88341a <=( A201  and  (not A200) );
 a88342a <=( a88341a  and  a88338a );
 a88343a <=( a88342a  and  a88335a );
 a88346a <=( (not A233)  and  A202 );
 a88349a <=( (not A266)  and  (not A234) );
 a88350a <=( a88349a  and  a88346a );
 a88353a <=( (not A269)  and  (not A268) );
 a88356a <=( A299  and  A298 );
 a88357a <=( a88356a  and  a88353a );
 a88358a <=( a88357a  and  a88350a );
 a88362a <=( A167  and  (not A168) );
 a88363a <=( A169  and  a88362a );
 a88366a <=( A199  and  (not A166) );
 a88369a <=( A201  and  (not A200) );
 a88370a <=( a88369a  and  a88366a );
 a88371a <=( a88370a  and  a88363a );
 a88374a <=( (not A233)  and  A202 );
 a88377a <=( (not A266)  and  (not A234) );
 a88378a <=( a88377a  and  a88374a );
 a88381a <=( (not A269)  and  (not A268) );
 a88384a <=( (not A299)  and  (not A298) );
 a88385a <=( a88384a  and  a88381a );
 a88386a <=( a88385a  and  a88378a );
 a88390a <=( A167  and  (not A168) );
 a88391a <=( A169  and  a88390a );
 a88394a <=( A199  and  (not A166) );
 a88397a <=( A201  and  (not A200) );
 a88398a <=( a88397a  and  a88394a );
 a88399a <=( a88398a  and  a88391a );
 a88402a <=( (not A233)  and  A202 );
 a88405a <=( (not A266)  and  (not A234) );
 a88406a <=( a88405a  and  a88402a );
 a88409a <=( A298  and  (not A267) );
 a88412a <=( (not A302)  and  (not A301) );
 a88413a <=( a88412a  and  a88409a );
 a88414a <=( a88413a  and  a88406a );
 a88418a <=( A167  and  (not A168) );
 a88419a <=( A169  and  a88418a );
 a88422a <=( A199  and  (not A166) );
 a88425a <=( A201  and  (not A200) );
 a88426a <=( a88425a  and  a88422a );
 a88427a <=( a88426a  and  a88419a );
 a88430a <=( (not A233)  and  A202 );
 a88433a <=( (not A265)  and  (not A234) );
 a88434a <=( a88433a  and  a88430a );
 a88437a <=( A298  and  (not A266) );
 a88440a <=( (not A302)  and  (not A301) );
 a88441a <=( a88440a  and  a88437a );
 a88442a <=( a88441a  and  a88434a );
 a88446a <=( A167  and  (not A168) );
 a88447a <=( A169  and  a88446a );
 a88450a <=( A199  and  (not A166) );
 a88453a <=( A201  and  (not A200) );
 a88454a <=( a88453a  and  a88450a );
 a88455a <=( a88454a  and  a88447a );
 a88458a <=( (not A232)  and  A202 );
 a88461a <=( A265  and  (not A233) );
 a88462a <=( a88461a  and  a88458a );
 a88465a <=( A298  and  A266 );
 a88468a <=( (not A302)  and  (not A301) );
 a88469a <=( a88468a  and  a88465a );
 a88470a <=( a88469a  and  a88462a );
 a88474a <=( A167  and  (not A168) );
 a88475a <=( A169  and  a88474a );
 a88478a <=( A199  and  (not A166) );
 a88481a <=( A201  and  (not A200) );
 a88482a <=( a88481a  and  a88478a );
 a88483a <=( a88482a  and  a88475a );
 a88486a <=( (not A232)  and  A202 );
 a88489a <=( (not A266)  and  (not A233) );
 a88490a <=( a88489a  and  a88486a );
 a88493a <=( (not A269)  and  (not A268) );
 a88496a <=( (not A300)  and  A298 );
 a88497a <=( a88496a  and  a88493a );
 a88498a <=( a88497a  and  a88490a );
 a88502a <=( A167  and  (not A168) );
 a88503a <=( A169  and  a88502a );
 a88506a <=( A199  and  (not A166) );
 a88509a <=( A201  and  (not A200) );
 a88510a <=( a88509a  and  a88506a );
 a88511a <=( a88510a  and  a88503a );
 a88514a <=( (not A232)  and  A202 );
 a88517a <=( (not A266)  and  (not A233) );
 a88518a <=( a88517a  and  a88514a );
 a88521a <=( (not A269)  and  (not A268) );
 a88524a <=( A299  and  A298 );
 a88525a <=( a88524a  and  a88521a );
 a88526a <=( a88525a  and  a88518a );
 a88530a <=( A167  and  (not A168) );
 a88531a <=( A169  and  a88530a );
 a88534a <=( A199  and  (not A166) );
 a88537a <=( A201  and  (not A200) );
 a88538a <=( a88537a  and  a88534a );
 a88539a <=( a88538a  and  a88531a );
 a88542a <=( (not A232)  and  A202 );
 a88545a <=( (not A266)  and  (not A233) );
 a88546a <=( a88545a  and  a88542a );
 a88549a <=( (not A269)  and  (not A268) );
 a88552a <=( (not A299)  and  (not A298) );
 a88553a <=( a88552a  and  a88549a );
 a88554a <=( a88553a  and  a88546a );
 a88558a <=( A167  and  (not A168) );
 a88559a <=( A169  and  a88558a );
 a88562a <=( A199  and  (not A166) );
 a88565a <=( A201  and  (not A200) );
 a88566a <=( a88565a  and  a88562a );
 a88567a <=( a88566a  and  a88559a );
 a88570a <=( (not A232)  and  A202 );
 a88573a <=( (not A266)  and  (not A233) );
 a88574a <=( a88573a  and  a88570a );
 a88577a <=( A298  and  (not A267) );
 a88580a <=( (not A302)  and  (not A301) );
 a88581a <=( a88580a  and  a88577a );
 a88582a <=( a88581a  and  a88574a );
 a88586a <=( A167  and  (not A168) );
 a88587a <=( A169  and  a88586a );
 a88590a <=( A199  and  (not A166) );
 a88593a <=( A201  and  (not A200) );
 a88594a <=( a88593a  and  a88590a );
 a88595a <=( a88594a  and  a88587a );
 a88598a <=( (not A232)  and  A202 );
 a88601a <=( (not A265)  and  (not A233) );
 a88602a <=( a88601a  and  a88598a );
 a88605a <=( A298  and  (not A266) );
 a88608a <=( (not A302)  and  (not A301) );
 a88609a <=( a88608a  and  a88605a );
 a88610a <=( a88609a  and  a88602a );
 a88614a <=( A167  and  (not A168) );
 a88615a <=( A169  and  a88614a );
 a88618a <=( A199  and  (not A166) );
 a88621a <=( A201  and  (not A200) );
 a88622a <=( a88621a  and  a88618a );
 a88623a <=( a88622a  and  a88615a );
 a88626a <=( A232  and  A203 );
 a88629a <=( A265  and  A233 );
 a88630a <=( a88629a  and  a88626a );
 a88633a <=( (not A269)  and  (not A268) );
 a88636a <=( (not A300)  and  (not A299) );
 a88637a <=( a88636a  and  a88633a );
 a88638a <=( a88637a  and  a88630a );
 a88642a <=( A167  and  (not A168) );
 a88643a <=( A169  and  a88642a );
 a88646a <=( A199  and  (not A166) );
 a88649a <=( A201  and  (not A200) );
 a88650a <=( a88649a  and  a88646a );
 a88651a <=( a88650a  and  a88643a );
 a88654a <=( A232  and  A203 );
 a88657a <=( A265  and  A233 );
 a88658a <=( a88657a  and  a88654a );
 a88661a <=( (not A269)  and  (not A268) );
 a88664a <=( A299  and  A298 );
 a88665a <=( a88664a  and  a88661a );
 a88666a <=( a88665a  and  a88658a );
 a88670a <=( A167  and  (not A168) );
 a88671a <=( A169  and  a88670a );
 a88674a <=( A199  and  (not A166) );
 a88677a <=( A201  and  (not A200) );
 a88678a <=( a88677a  and  a88674a );
 a88679a <=( a88678a  and  a88671a );
 a88682a <=( A232  and  A203 );
 a88685a <=( A265  and  A233 );
 a88686a <=( a88685a  and  a88682a );
 a88689a <=( (not A269)  and  (not A268) );
 a88692a <=( (not A299)  and  (not A298) );
 a88693a <=( a88692a  and  a88689a );
 a88694a <=( a88693a  and  a88686a );
 a88698a <=( A167  and  (not A168) );
 a88699a <=( A169  and  a88698a );
 a88702a <=( A199  and  (not A166) );
 a88705a <=( A201  and  (not A200) );
 a88706a <=( a88705a  and  a88702a );
 a88707a <=( a88706a  and  a88699a );
 a88710a <=( A232  and  A203 );
 a88713a <=( A265  and  A233 );
 a88714a <=( a88713a  and  a88710a );
 a88717a <=( (not A299)  and  (not A267) );
 a88720a <=( (not A302)  and  (not A301) );
 a88721a <=( a88720a  and  a88717a );
 a88722a <=( a88721a  and  a88714a );
 a88726a <=( A167  and  (not A168) );
 a88727a <=( A169  and  a88726a );
 a88730a <=( A199  and  (not A166) );
 a88733a <=( A201  and  (not A200) );
 a88734a <=( a88733a  and  a88730a );
 a88735a <=( a88734a  and  a88727a );
 a88738a <=( A232  and  A203 );
 a88741a <=( A265  and  A233 );
 a88742a <=( a88741a  and  a88738a );
 a88745a <=( (not A299)  and  A266 );
 a88748a <=( (not A302)  and  (not A301) );
 a88749a <=( a88748a  and  a88745a );
 a88750a <=( a88749a  and  a88742a );
 a88754a <=( A167  and  (not A168) );
 a88755a <=( A169  and  a88754a );
 a88758a <=( A199  and  (not A166) );
 a88761a <=( A201  and  (not A200) );
 a88762a <=( a88761a  and  a88758a );
 a88763a <=( a88762a  and  a88755a );
 a88766a <=( A232  and  A203 );
 a88769a <=( (not A265)  and  A233 );
 a88770a <=( a88769a  and  a88766a );
 a88773a <=( (not A299)  and  (not A266) );
 a88776a <=( (not A302)  and  (not A301) );
 a88777a <=( a88776a  and  a88773a );
 a88778a <=( a88777a  and  a88770a );
 a88782a <=( A167  and  (not A168) );
 a88783a <=( A169  and  a88782a );
 a88786a <=( A199  and  (not A166) );
 a88789a <=( A201  and  (not A200) );
 a88790a <=( a88789a  and  a88786a );
 a88791a <=( a88790a  and  a88783a );
 a88794a <=( (not A233)  and  A203 );
 a88797a <=( (not A236)  and  (not A235) );
 a88798a <=( a88797a  and  a88794a );
 a88801a <=( A266  and  A265 );
 a88804a <=( (not A300)  and  A298 );
 a88805a <=( a88804a  and  a88801a );
 a88806a <=( a88805a  and  a88798a );
 a88810a <=( A167  and  (not A168) );
 a88811a <=( A169  and  a88810a );
 a88814a <=( A199  and  (not A166) );
 a88817a <=( A201  and  (not A200) );
 a88818a <=( a88817a  and  a88814a );
 a88819a <=( a88818a  and  a88811a );
 a88822a <=( (not A233)  and  A203 );
 a88825a <=( (not A236)  and  (not A235) );
 a88826a <=( a88825a  and  a88822a );
 a88829a <=( A266  and  A265 );
 a88832a <=( A299  and  A298 );
 a88833a <=( a88832a  and  a88829a );
 a88834a <=( a88833a  and  a88826a );
 a88838a <=( A167  and  (not A168) );
 a88839a <=( A169  and  a88838a );
 a88842a <=( A199  and  (not A166) );
 a88845a <=( A201  and  (not A200) );
 a88846a <=( a88845a  and  a88842a );
 a88847a <=( a88846a  and  a88839a );
 a88850a <=( (not A233)  and  A203 );
 a88853a <=( (not A236)  and  (not A235) );
 a88854a <=( a88853a  and  a88850a );
 a88857a <=( A266  and  A265 );
 a88860a <=( (not A299)  and  (not A298) );
 a88861a <=( a88860a  and  a88857a );
 a88862a <=( a88861a  and  a88854a );
 a88866a <=( A167  and  (not A168) );
 a88867a <=( A169  and  a88866a );
 a88870a <=( A199  and  (not A166) );
 a88873a <=( A201  and  (not A200) );
 a88874a <=( a88873a  and  a88870a );
 a88875a <=( a88874a  and  a88867a );
 a88878a <=( (not A233)  and  A203 );
 a88881a <=( (not A236)  and  (not A235) );
 a88882a <=( a88881a  and  a88878a );
 a88885a <=( (not A267)  and  (not A266) );
 a88888a <=( (not A300)  and  A298 );
 a88889a <=( a88888a  and  a88885a );
 a88890a <=( a88889a  and  a88882a );
 a88894a <=( A167  and  (not A168) );
 a88895a <=( A169  and  a88894a );
 a88898a <=( A199  and  (not A166) );
 a88901a <=( A201  and  (not A200) );
 a88902a <=( a88901a  and  a88898a );
 a88903a <=( a88902a  and  a88895a );
 a88906a <=( (not A233)  and  A203 );
 a88909a <=( (not A236)  and  (not A235) );
 a88910a <=( a88909a  and  a88906a );
 a88913a <=( (not A267)  and  (not A266) );
 a88916a <=( A299  and  A298 );
 a88917a <=( a88916a  and  a88913a );
 a88918a <=( a88917a  and  a88910a );
 a88922a <=( A167  and  (not A168) );
 a88923a <=( A169  and  a88922a );
 a88926a <=( A199  and  (not A166) );
 a88929a <=( A201  and  (not A200) );
 a88930a <=( a88929a  and  a88926a );
 a88931a <=( a88930a  and  a88923a );
 a88934a <=( (not A233)  and  A203 );
 a88937a <=( (not A236)  and  (not A235) );
 a88938a <=( a88937a  and  a88934a );
 a88941a <=( (not A267)  and  (not A266) );
 a88944a <=( (not A299)  and  (not A298) );
 a88945a <=( a88944a  and  a88941a );
 a88946a <=( a88945a  and  a88938a );
 a88950a <=( A167  and  (not A168) );
 a88951a <=( A169  and  a88950a );
 a88954a <=( A199  and  (not A166) );
 a88957a <=( A201  and  (not A200) );
 a88958a <=( a88957a  and  a88954a );
 a88959a <=( a88958a  and  a88951a );
 a88962a <=( (not A233)  and  A203 );
 a88965a <=( (not A236)  and  (not A235) );
 a88966a <=( a88965a  and  a88962a );
 a88969a <=( (not A266)  and  (not A265) );
 a88972a <=( (not A300)  and  A298 );
 a88973a <=( a88972a  and  a88969a );
 a88974a <=( a88973a  and  a88966a );
 a88978a <=( A167  and  (not A168) );
 a88979a <=( A169  and  a88978a );
 a88982a <=( A199  and  (not A166) );
 a88985a <=( A201  and  (not A200) );
 a88986a <=( a88985a  and  a88982a );
 a88987a <=( a88986a  and  a88979a );
 a88990a <=( (not A233)  and  A203 );
 a88993a <=( (not A236)  and  (not A235) );
 a88994a <=( a88993a  and  a88990a );
 a88997a <=( (not A266)  and  (not A265) );
 a89000a <=( A299  and  A298 );
 a89001a <=( a89000a  and  a88997a );
 a89002a <=( a89001a  and  a88994a );
 a89006a <=( A167  and  (not A168) );
 a89007a <=( A169  and  a89006a );
 a89010a <=( A199  and  (not A166) );
 a89013a <=( A201  and  (not A200) );
 a89014a <=( a89013a  and  a89010a );
 a89015a <=( a89014a  and  a89007a );
 a89018a <=( (not A233)  and  A203 );
 a89021a <=( (not A236)  and  (not A235) );
 a89022a <=( a89021a  and  a89018a );
 a89025a <=( (not A266)  and  (not A265) );
 a89028a <=( (not A299)  and  (not A298) );
 a89029a <=( a89028a  and  a89025a );
 a89030a <=( a89029a  and  a89022a );
 a89034a <=( A167  and  (not A168) );
 a89035a <=( A169  and  a89034a );
 a89038a <=( A199  and  (not A166) );
 a89041a <=( A201  and  (not A200) );
 a89042a <=( a89041a  and  a89038a );
 a89043a <=( a89042a  and  a89035a );
 a89046a <=( (not A233)  and  A203 );
 a89049a <=( A265  and  (not A234) );
 a89050a <=( a89049a  and  a89046a );
 a89053a <=( A298  and  A266 );
 a89056a <=( (not A302)  and  (not A301) );
 a89057a <=( a89056a  and  a89053a );
 a89058a <=( a89057a  and  a89050a );
 a89062a <=( A167  and  (not A168) );
 a89063a <=( A169  and  a89062a );
 a89066a <=( A199  and  (not A166) );
 a89069a <=( A201  and  (not A200) );
 a89070a <=( a89069a  and  a89066a );
 a89071a <=( a89070a  and  a89063a );
 a89074a <=( (not A233)  and  A203 );
 a89077a <=( (not A266)  and  (not A234) );
 a89078a <=( a89077a  and  a89074a );
 a89081a <=( (not A269)  and  (not A268) );
 a89084a <=( (not A300)  and  A298 );
 a89085a <=( a89084a  and  a89081a );
 a89086a <=( a89085a  and  a89078a );
 a89090a <=( A167  and  (not A168) );
 a89091a <=( A169  and  a89090a );
 a89094a <=( A199  and  (not A166) );
 a89097a <=( A201  and  (not A200) );
 a89098a <=( a89097a  and  a89094a );
 a89099a <=( a89098a  and  a89091a );
 a89102a <=( (not A233)  and  A203 );
 a89105a <=( (not A266)  and  (not A234) );
 a89106a <=( a89105a  and  a89102a );
 a89109a <=( (not A269)  and  (not A268) );
 a89112a <=( A299  and  A298 );
 a89113a <=( a89112a  and  a89109a );
 a89114a <=( a89113a  and  a89106a );
 a89118a <=( A167  and  (not A168) );
 a89119a <=( A169  and  a89118a );
 a89122a <=( A199  and  (not A166) );
 a89125a <=( A201  and  (not A200) );
 a89126a <=( a89125a  and  a89122a );
 a89127a <=( a89126a  and  a89119a );
 a89130a <=( (not A233)  and  A203 );
 a89133a <=( (not A266)  and  (not A234) );
 a89134a <=( a89133a  and  a89130a );
 a89137a <=( (not A269)  and  (not A268) );
 a89140a <=( (not A299)  and  (not A298) );
 a89141a <=( a89140a  and  a89137a );
 a89142a <=( a89141a  and  a89134a );
 a89146a <=( A167  and  (not A168) );
 a89147a <=( A169  and  a89146a );
 a89150a <=( A199  and  (not A166) );
 a89153a <=( A201  and  (not A200) );
 a89154a <=( a89153a  and  a89150a );
 a89155a <=( a89154a  and  a89147a );
 a89158a <=( (not A233)  and  A203 );
 a89161a <=( (not A266)  and  (not A234) );
 a89162a <=( a89161a  and  a89158a );
 a89165a <=( A298  and  (not A267) );
 a89168a <=( (not A302)  and  (not A301) );
 a89169a <=( a89168a  and  a89165a );
 a89170a <=( a89169a  and  a89162a );
 a89174a <=( A167  and  (not A168) );
 a89175a <=( A169  and  a89174a );
 a89178a <=( A199  and  (not A166) );
 a89181a <=( A201  and  (not A200) );
 a89182a <=( a89181a  and  a89178a );
 a89183a <=( a89182a  and  a89175a );
 a89186a <=( (not A233)  and  A203 );
 a89189a <=( (not A265)  and  (not A234) );
 a89190a <=( a89189a  and  a89186a );
 a89193a <=( A298  and  (not A266) );
 a89196a <=( (not A302)  and  (not A301) );
 a89197a <=( a89196a  and  a89193a );
 a89198a <=( a89197a  and  a89190a );
 a89202a <=( A167  and  (not A168) );
 a89203a <=( A169  and  a89202a );
 a89206a <=( A199  and  (not A166) );
 a89209a <=( A201  and  (not A200) );
 a89210a <=( a89209a  and  a89206a );
 a89211a <=( a89210a  and  a89203a );
 a89214a <=( (not A232)  and  A203 );
 a89217a <=( A265  and  (not A233) );
 a89218a <=( a89217a  and  a89214a );
 a89221a <=( A298  and  A266 );
 a89224a <=( (not A302)  and  (not A301) );
 a89225a <=( a89224a  and  a89221a );
 a89226a <=( a89225a  and  a89218a );
 a89230a <=( A167  and  (not A168) );
 a89231a <=( A169  and  a89230a );
 a89234a <=( A199  and  (not A166) );
 a89237a <=( A201  and  (not A200) );
 a89238a <=( a89237a  and  a89234a );
 a89239a <=( a89238a  and  a89231a );
 a89242a <=( (not A232)  and  A203 );
 a89245a <=( (not A266)  and  (not A233) );
 a89246a <=( a89245a  and  a89242a );
 a89249a <=( (not A269)  and  (not A268) );
 a89252a <=( (not A300)  and  A298 );
 a89253a <=( a89252a  and  a89249a );
 a89254a <=( a89253a  and  a89246a );
 a89258a <=( A167  and  (not A168) );
 a89259a <=( A169  and  a89258a );
 a89262a <=( A199  and  (not A166) );
 a89265a <=( A201  and  (not A200) );
 a89266a <=( a89265a  and  a89262a );
 a89267a <=( a89266a  and  a89259a );
 a89270a <=( (not A232)  and  A203 );
 a89273a <=( (not A266)  and  (not A233) );
 a89274a <=( a89273a  and  a89270a );
 a89277a <=( (not A269)  and  (not A268) );
 a89280a <=( A299  and  A298 );
 a89281a <=( a89280a  and  a89277a );
 a89282a <=( a89281a  and  a89274a );
 a89286a <=( A167  and  (not A168) );
 a89287a <=( A169  and  a89286a );
 a89290a <=( A199  and  (not A166) );
 a89293a <=( A201  and  (not A200) );
 a89294a <=( a89293a  and  a89290a );
 a89295a <=( a89294a  and  a89287a );
 a89298a <=( (not A232)  and  A203 );
 a89301a <=( (not A266)  and  (not A233) );
 a89302a <=( a89301a  and  a89298a );
 a89305a <=( (not A269)  and  (not A268) );
 a89308a <=( (not A299)  and  (not A298) );
 a89309a <=( a89308a  and  a89305a );
 a89310a <=( a89309a  and  a89302a );
 a89314a <=( A167  and  (not A168) );
 a89315a <=( A169  and  a89314a );
 a89318a <=( A199  and  (not A166) );
 a89321a <=( A201  and  (not A200) );
 a89322a <=( a89321a  and  a89318a );
 a89323a <=( a89322a  and  a89315a );
 a89326a <=( (not A232)  and  A203 );
 a89329a <=( (not A266)  and  (not A233) );
 a89330a <=( a89329a  and  a89326a );
 a89333a <=( A298  and  (not A267) );
 a89336a <=( (not A302)  and  (not A301) );
 a89337a <=( a89336a  and  a89333a );
 a89338a <=( a89337a  and  a89330a );
 a89342a <=( A167  and  (not A168) );
 a89343a <=( A169  and  a89342a );
 a89346a <=( A199  and  (not A166) );
 a89349a <=( A201  and  (not A200) );
 a89350a <=( a89349a  and  a89346a );
 a89351a <=( a89350a  and  a89343a );
 a89354a <=( (not A232)  and  A203 );
 a89357a <=( (not A265)  and  (not A233) );
 a89358a <=( a89357a  and  a89354a );
 a89361a <=( A298  and  (not A266) );
 a89364a <=( (not A302)  and  (not A301) );
 a89365a <=( a89364a  and  a89361a );
 a89366a <=( a89365a  and  a89358a );
 a89370a <=( (not A167)  and  (not A168) );
 a89371a <=( A169  and  a89370a );
 a89374a <=( (not A199)  and  A166 );
 a89377a <=( (not A233)  and  A200 );
 a89378a <=( a89377a  and  a89374a );
 a89379a <=( a89378a  and  a89371a );
 a89382a <=( (not A236)  and  (not A235) );
 a89385a <=( (not A268)  and  (not A266) );
 a89386a <=( a89385a  and  a89382a );
 a89389a <=( A298  and  (not A269) );
 a89392a <=( (not A302)  and  (not A301) );
 a89393a <=( a89392a  and  a89389a );
 a89394a <=( a89393a  and  a89386a );
 a89398a <=( (not A167)  and  (not A168) );
 a89399a <=( A169  and  a89398a );
 a89402a <=( A199  and  A166 );
 a89405a <=( A201  and  (not A200) );
 a89406a <=( a89405a  and  a89402a );
 a89407a <=( a89406a  and  a89399a );
 a89410a <=( A232  and  A202 );
 a89413a <=( A265  and  A233 );
 a89414a <=( a89413a  and  a89410a );
 a89417a <=( (not A269)  and  (not A268) );
 a89420a <=( (not A300)  and  (not A299) );
 a89421a <=( a89420a  and  a89417a );
 a89422a <=( a89421a  and  a89414a );
 a89426a <=( (not A167)  and  (not A168) );
 a89427a <=( A169  and  a89426a );
 a89430a <=( A199  and  A166 );
 a89433a <=( A201  and  (not A200) );
 a89434a <=( a89433a  and  a89430a );
 a89435a <=( a89434a  and  a89427a );
 a89438a <=( A232  and  A202 );
 a89441a <=( A265  and  A233 );
 a89442a <=( a89441a  and  a89438a );
 a89445a <=( (not A269)  and  (not A268) );
 a89448a <=( A299  and  A298 );
 a89449a <=( a89448a  and  a89445a );
 a89450a <=( a89449a  and  a89442a );
 a89454a <=( (not A167)  and  (not A168) );
 a89455a <=( A169  and  a89454a );
 a89458a <=( A199  and  A166 );
 a89461a <=( A201  and  (not A200) );
 a89462a <=( a89461a  and  a89458a );
 a89463a <=( a89462a  and  a89455a );
 a89466a <=( A232  and  A202 );
 a89469a <=( A265  and  A233 );
 a89470a <=( a89469a  and  a89466a );
 a89473a <=( (not A269)  and  (not A268) );
 a89476a <=( (not A299)  and  (not A298) );
 a89477a <=( a89476a  and  a89473a );
 a89478a <=( a89477a  and  a89470a );
 a89482a <=( (not A167)  and  (not A168) );
 a89483a <=( A169  and  a89482a );
 a89486a <=( A199  and  A166 );
 a89489a <=( A201  and  (not A200) );
 a89490a <=( a89489a  and  a89486a );
 a89491a <=( a89490a  and  a89483a );
 a89494a <=( A232  and  A202 );
 a89497a <=( A265  and  A233 );
 a89498a <=( a89497a  and  a89494a );
 a89501a <=( (not A299)  and  (not A267) );
 a89504a <=( (not A302)  and  (not A301) );
 a89505a <=( a89504a  and  a89501a );
 a89506a <=( a89505a  and  a89498a );
 a89510a <=( (not A167)  and  (not A168) );
 a89511a <=( A169  and  a89510a );
 a89514a <=( A199  and  A166 );
 a89517a <=( A201  and  (not A200) );
 a89518a <=( a89517a  and  a89514a );
 a89519a <=( a89518a  and  a89511a );
 a89522a <=( A232  and  A202 );
 a89525a <=( A265  and  A233 );
 a89526a <=( a89525a  and  a89522a );
 a89529a <=( (not A299)  and  A266 );
 a89532a <=( (not A302)  and  (not A301) );
 a89533a <=( a89532a  and  a89529a );
 a89534a <=( a89533a  and  a89526a );
 a89538a <=( (not A167)  and  (not A168) );
 a89539a <=( A169  and  a89538a );
 a89542a <=( A199  and  A166 );
 a89545a <=( A201  and  (not A200) );
 a89546a <=( a89545a  and  a89542a );
 a89547a <=( a89546a  and  a89539a );
 a89550a <=( A232  and  A202 );
 a89553a <=( (not A265)  and  A233 );
 a89554a <=( a89553a  and  a89550a );
 a89557a <=( (not A299)  and  (not A266) );
 a89560a <=( (not A302)  and  (not A301) );
 a89561a <=( a89560a  and  a89557a );
 a89562a <=( a89561a  and  a89554a );
 a89566a <=( (not A167)  and  (not A168) );
 a89567a <=( A169  and  a89566a );
 a89570a <=( A199  and  A166 );
 a89573a <=( A201  and  (not A200) );
 a89574a <=( a89573a  and  a89570a );
 a89575a <=( a89574a  and  a89567a );
 a89578a <=( (not A233)  and  A202 );
 a89581a <=( (not A236)  and  (not A235) );
 a89582a <=( a89581a  and  a89578a );
 a89585a <=( A266  and  A265 );
 a89588a <=( (not A300)  and  A298 );
 a89589a <=( a89588a  and  a89585a );
 a89590a <=( a89589a  and  a89582a );
 a89594a <=( (not A167)  and  (not A168) );
 a89595a <=( A169  and  a89594a );
 a89598a <=( A199  and  A166 );
 a89601a <=( A201  and  (not A200) );
 a89602a <=( a89601a  and  a89598a );
 a89603a <=( a89602a  and  a89595a );
 a89606a <=( (not A233)  and  A202 );
 a89609a <=( (not A236)  and  (not A235) );
 a89610a <=( a89609a  and  a89606a );
 a89613a <=( A266  and  A265 );
 a89616a <=( A299  and  A298 );
 a89617a <=( a89616a  and  a89613a );
 a89618a <=( a89617a  and  a89610a );
 a89622a <=( (not A167)  and  (not A168) );
 a89623a <=( A169  and  a89622a );
 a89626a <=( A199  and  A166 );
 a89629a <=( A201  and  (not A200) );
 a89630a <=( a89629a  and  a89626a );
 a89631a <=( a89630a  and  a89623a );
 a89634a <=( (not A233)  and  A202 );
 a89637a <=( (not A236)  and  (not A235) );
 a89638a <=( a89637a  and  a89634a );
 a89641a <=( A266  and  A265 );
 a89644a <=( (not A299)  and  (not A298) );
 a89645a <=( a89644a  and  a89641a );
 a89646a <=( a89645a  and  a89638a );
 a89650a <=( (not A167)  and  (not A168) );
 a89651a <=( A169  and  a89650a );
 a89654a <=( A199  and  A166 );
 a89657a <=( A201  and  (not A200) );
 a89658a <=( a89657a  and  a89654a );
 a89659a <=( a89658a  and  a89651a );
 a89662a <=( (not A233)  and  A202 );
 a89665a <=( (not A236)  and  (not A235) );
 a89666a <=( a89665a  and  a89662a );
 a89669a <=( (not A267)  and  (not A266) );
 a89672a <=( (not A300)  and  A298 );
 a89673a <=( a89672a  and  a89669a );
 a89674a <=( a89673a  and  a89666a );
 a89678a <=( (not A167)  and  (not A168) );
 a89679a <=( A169  and  a89678a );
 a89682a <=( A199  and  A166 );
 a89685a <=( A201  and  (not A200) );
 a89686a <=( a89685a  and  a89682a );
 a89687a <=( a89686a  and  a89679a );
 a89690a <=( (not A233)  and  A202 );
 a89693a <=( (not A236)  and  (not A235) );
 a89694a <=( a89693a  and  a89690a );
 a89697a <=( (not A267)  and  (not A266) );
 a89700a <=( A299  and  A298 );
 a89701a <=( a89700a  and  a89697a );
 a89702a <=( a89701a  and  a89694a );
 a89706a <=( (not A167)  and  (not A168) );
 a89707a <=( A169  and  a89706a );
 a89710a <=( A199  and  A166 );
 a89713a <=( A201  and  (not A200) );
 a89714a <=( a89713a  and  a89710a );
 a89715a <=( a89714a  and  a89707a );
 a89718a <=( (not A233)  and  A202 );
 a89721a <=( (not A236)  and  (not A235) );
 a89722a <=( a89721a  and  a89718a );
 a89725a <=( (not A267)  and  (not A266) );
 a89728a <=( (not A299)  and  (not A298) );
 a89729a <=( a89728a  and  a89725a );
 a89730a <=( a89729a  and  a89722a );
 a89734a <=( (not A167)  and  (not A168) );
 a89735a <=( A169  and  a89734a );
 a89738a <=( A199  and  A166 );
 a89741a <=( A201  and  (not A200) );
 a89742a <=( a89741a  and  a89738a );
 a89743a <=( a89742a  and  a89735a );
 a89746a <=( (not A233)  and  A202 );
 a89749a <=( (not A236)  and  (not A235) );
 a89750a <=( a89749a  and  a89746a );
 a89753a <=( (not A266)  and  (not A265) );
 a89756a <=( (not A300)  and  A298 );
 a89757a <=( a89756a  and  a89753a );
 a89758a <=( a89757a  and  a89750a );
 a89762a <=( (not A167)  and  (not A168) );
 a89763a <=( A169  and  a89762a );
 a89766a <=( A199  and  A166 );
 a89769a <=( A201  and  (not A200) );
 a89770a <=( a89769a  and  a89766a );
 a89771a <=( a89770a  and  a89763a );
 a89774a <=( (not A233)  and  A202 );
 a89777a <=( (not A236)  and  (not A235) );
 a89778a <=( a89777a  and  a89774a );
 a89781a <=( (not A266)  and  (not A265) );
 a89784a <=( A299  and  A298 );
 a89785a <=( a89784a  and  a89781a );
 a89786a <=( a89785a  and  a89778a );
 a89790a <=( (not A167)  and  (not A168) );
 a89791a <=( A169  and  a89790a );
 a89794a <=( A199  and  A166 );
 a89797a <=( A201  and  (not A200) );
 a89798a <=( a89797a  and  a89794a );
 a89799a <=( a89798a  and  a89791a );
 a89802a <=( (not A233)  and  A202 );
 a89805a <=( (not A236)  and  (not A235) );
 a89806a <=( a89805a  and  a89802a );
 a89809a <=( (not A266)  and  (not A265) );
 a89812a <=( (not A299)  and  (not A298) );
 a89813a <=( a89812a  and  a89809a );
 a89814a <=( a89813a  and  a89806a );
 a89818a <=( (not A167)  and  (not A168) );
 a89819a <=( A169  and  a89818a );
 a89822a <=( A199  and  A166 );
 a89825a <=( A201  and  (not A200) );
 a89826a <=( a89825a  and  a89822a );
 a89827a <=( a89826a  and  a89819a );
 a89830a <=( (not A233)  and  A202 );
 a89833a <=( A265  and  (not A234) );
 a89834a <=( a89833a  and  a89830a );
 a89837a <=( A298  and  A266 );
 a89840a <=( (not A302)  and  (not A301) );
 a89841a <=( a89840a  and  a89837a );
 a89842a <=( a89841a  and  a89834a );
 a89846a <=( (not A167)  and  (not A168) );
 a89847a <=( A169  and  a89846a );
 a89850a <=( A199  and  A166 );
 a89853a <=( A201  and  (not A200) );
 a89854a <=( a89853a  and  a89850a );
 a89855a <=( a89854a  and  a89847a );
 a89858a <=( (not A233)  and  A202 );
 a89861a <=( (not A266)  and  (not A234) );
 a89862a <=( a89861a  and  a89858a );
 a89865a <=( (not A269)  and  (not A268) );
 a89868a <=( (not A300)  and  A298 );
 a89869a <=( a89868a  and  a89865a );
 a89870a <=( a89869a  and  a89862a );
 a89874a <=( (not A167)  and  (not A168) );
 a89875a <=( A169  and  a89874a );
 a89878a <=( A199  and  A166 );
 a89881a <=( A201  and  (not A200) );
 a89882a <=( a89881a  and  a89878a );
 a89883a <=( a89882a  and  a89875a );
 a89886a <=( (not A233)  and  A202 );
 a89889a <=( (not A266)  and  (not A234) );
 a89890a <=( a89889a  and  a89886a );
 a89893a <=( (not A269)  and  (not A268) );
 a89896a <=( A299  and  A298 );
 a89897a <=( a89896a  and  a89893a );
 a89898a <=( a89897a  and  a89890a );
 a89902a <=( (not A167)  and  (not A168) );
 a89903a <=( A169  and  a89902a );
 a89906a <=( A199  and  A166 );
 a89909a <=( A201  and  (not A200) );
 a89910a <=( a89909a  and  a89906a );
 a89911a <=( a89910a  and  a89903a );
 a89914a <=( (not A233)  and  A202 );
 a89917a <=( (not A266)  and  (not A234) );
 a89918a <=( a89917a  and  a89914a );
 a89921a <=( (not A269)  and  (not A268) );
 a89924a <=( (not A299)  and  (not A298) );
 a89925a <=( a89924a  and  a89921a );
 a89926a <=( a89925a  and  a89918a );
 a89930a <=( (not A167)  and  (not A168) );
 a89931a <=( A169  and  a89930a );
 a89934a <=( A199  and  A166 );
 a89937a <=( A201  and  (not A200) );
 a89938a <=( a89937a  and  a89934a );
 a89939a <=( a89938a  and  a89931a );
 a89942a <=( (not A233)  and  A202 );
 a89945a <=( (not A266)  and  (not A234) );
 a89946a <=( a89945a  and  a89942a );
 a89949a <=( A298  and  (not A267) );
 a89952a <=( (not A302)  and  (not A301) );
 a89953a <=( a89952a  and  a89949a );
 a89954a <=( a89953a  and  a89946a );
 a89958a <=( (not A167)  and  (not A168) );
 a89959a <=( A169  and  a89958a );
 a89962a <=( A199  and  A166 );
 a89965a <=( A201  and  (not A200) );
 a89966a <=( a89965a  and  a89962a );
 a89967a <=( a89966a  and  a89959a );
 a89970a <=( (not A233)  and  A202 );
 a89973a <=( (not A265)  and  (not A234) );
 a89974a <=( a89973a  and  a89970a );
 a89977a <=( A298  and  (not A266) );
 a89980a <=( (not A302)  and  (not A301) );
 a89981a <=( a89980a  and  a89977a );
 a89982a <=( a89981a  and  a89974a );
 a89986a <=( (not A167)  and  (not A168) );
 a89987a <=( A169  and  a89986a );
 a89990a <=( A199  and  A166 );
 a89993a <=( A201  and  (not A200) );
 a89994a <=( a89993a  and  a89990a );
 a89995a <=( a89994a  and  a89987a );
 a89998a <=( (not A232)  and  A202 );
 a90001a <=( A265  and  (not A233) );
 a90002a <=( a90001a  and  a89998a );
 a90005a <=( A298  and  A266 );
 a90008a <=( (not A302)  and  (not A301) );
 a90009a <=( a90008a  and  a90005a );
 a90010a <=( a90009a  and  a90002a );
 a90014a <=( (not A167)  and  (not A168) );
 a90015a <=( A169  and  a90014a );
 a90018a <=( A199  and  A166 );
 a90021a <=( A201  and  (not A200) );
 a90022a <=( a90021a  and  a90018a );
 a90023a <=( a90022a  and  a90015a );
 a90026a <=( (not A232)  and  A202 );
 a90029a <=( (not A266)  and  (not A233) );
 a90030a <=( a90029a  and  a90026a );
 a90033a <=( (not A269)  and  (not A268) );
 a90036a <=( (not A300)  and  A298 );
 a90037a <=( a90036a  and  a90033a );
 a90038a <=( a90037a  and  a90030a );
 a90042a <=( (not A167)  and  (not A168) );
 a90043a <=( A169  and  a90042a );
 a90046a <=( A199  and  A166 );
 a90049a <=( A201  and  (not A200) );
 a90050a <=( a90049a  and  a90046a );
 a90051a <=( a90050a  and  a90043a );
 a90054a <=( (not A232)  and  A202 );
 a90057a <=( (not A266)  and  (not A233) );
 a90058a <=( a90057a  and  a90054a );
 a90061a <=( (not A269)  and  (not A268) );
 a90064a <=( A299  and  A298 );
 a90065a <=( a90064a  and  a90061a );
 a90066a <=( a90065a  and  a90058a );
 a90070a <=( (not A167)  and  (not A168) );
 a90071a <=( A169  and  a90070a );
 a90074a <=( A199  and  A166 );
 a90077a <=( A201  and  (not A200) );
 a90078a <=( a90077a  and  a90074a );
 a90079a <=( a90078a  and  a90071a );
 a90082a <=( (not A232)  and  A202 );
 a90085a <=( (not A266)  and  (not A233) );
 a90086a <=( a90085a  and  a90082a );
 a90089a <=( (not A269)  and  (not A268) );
 a90092a <=( (not A299)  and  (not A298) );
 a90093a <=( a90092a  and  a90089a );
 a90094a <=( a90093a  and  a90086a );
 a90098a <=( (not A167)  and  (not A168) );
 a90099a <=( A169  and  a90098a );
 a90102a <=( A199  and  A166 );
 a90105a <=( A201  and  (not A200) );
 a90106a <=( a90105a  and  a90102a );
 a90107a <=( a90106a  and  a90099a );
 a90110a <=( (not A232)  and  A202 );
 a90113a <=( (not A266)  and  (not A233) );
 a90114a <=( a90113a  and  a90110a );
 a90117a <=( A298  and  (not A267) );
 a90120a <=( (not A302)  and  (not A301) );
 a90121a <=( a90120a  and  a90117a );
 a90122a <=( a90121a  and  a90114a );
 a90126a <=( (not A167)  and  (not A168) );
 a90127a <=( A169  and  a90126a );
 a90130a <=( A199  and  A166 );
 a90133a <=( A201  and  (not A200) );
 a90134a <=( a90133a  and  a90130a );
 a90135a <=( a90134a  and  a90127a );
 a90138a <=( (not A232)  and  A202 );
 a90141a <=( (not A265)  and  (not A233) );
 a90142a <=( a90141a  and  a90138a );
 a90145a <=( A298  and  (not A266) );
 a90148a <=( (not A302)  and  (not A301) );
 a90149a <=( a90148a  and  a90145a );
 a90150a <=( a90149a  and  a90142a );
 a90154a <=( (not A167)  and  (not A168) );
 a90155a <=( A169  and  a90154a );
 a90158a <=( A199  and  A166 );
 a90161a <=( A201  and  (not A200) );
 a90162a <=( a90161a  and  a90158a );
 a90163a <=( a90162a  and  a90155a );
 a90166a <=( A232  and  A203 );
 a90169a <=( A265  and  A233 );
 a90170a <=( a90169a  and  a90166a );
 a90173a <=( (not A269)  and  (not A268) );
 a90176a <=( (not A300)  and  (not A299) );
 a90177a <=( a90176a  and  a90173a );
 a90178a <=( a90177a  and  a90170a );
 a90182a <=( (not A167)  and  (not A168) );
 a90183a <=( A169  and  a90182a );
 a90186a <=( A199  and  A166 );
 a90189a <=( A201  and  (not A200) );
 a90190a <=( a90189a  and  a90186a );
 a90191a <=( a90190a  and  a90183a );
 a90194a <=( A232  and  A203 );
 a90197a <=( A265  and  A233 );
 a90198a <=( a90197a  and  a90194a );
 a90201a <=( (not A269)  and  (not A268) );
 a90204a <=( A299  and  A298 );
 a90205a <=( a90204a  and  a90201a );
 a90206a <=( a90205a  and  a90198a );
 a90210a <=( (not A167)  and  (not A168) );
 a90211a <=( A169  and  a90210a );
 a90214a <=( A199  and  A166 );
 a90217a <=( A201  and  (not A200) );
 a90218a <=( a90217a  and  a90214a );
 a90219a <=( a90218a  and  a90211a );
 a90222a <=( A232  and  A203 );
 a90225a <=( A265  and  A233 );
 a90226a <=( a90225a  and  a90222a );
 a90229a <=( (not A269)  and  (not A268) );
 a90232a <=( (not A299)  and  (not A298) );
 a90233a <=( a90232a  and  a90229a );
 a90234a <=( a90233a  and  a90226a );
 a90238a <=( (not A167)  and  (not A168) );
 a90239a <=( A169  and  a90238a );
 a90242a <=( A199  and  A166 );
 a90245a <=( A201  and  (not A200) );
 a90246a <=( a90245a  and  a90242a );
 a90247a <=( a90246a  and  a90239a );
 a90250a <=( A232  and  A203 );
 a90253a <=( A265  and  A233 );
 a90254a <=( a90253a  and  a90250a );
 a90257a <=( (not A299)  and  (not A267) );
 a90260a <=( (not A302)  and  (not A301) );
 a90261a <=( a90260a  and  a90257a );
 a90262a <=( a90261a  and  a90254a );
 a90266a <=( (not A167)  and  (not A168) );
 a90267a <=( A169  and  a90266a );
 a90270a <=( A199  and  A166 );
 a90273a <=( A201  and  (not A200) );
 a90274a <=( a90273a  and  a90270a );
 a90275a <=( a90274a  and  a90267a );
 a90278a <=( A232  and  A203 );
 a90281a <=( A265  and  A233 );
 a90282a <=( a90281a  and  a90278a );
 a90285a <=( (not A299)  and  A266 );
 a90288a <=( (not A302)  and  (not A301) );
 a90289a <=( a90288a  and  a90285a );
 a90290a <=( a90289a  and  a90282a );
 a90294a <=( (not A167)  and  (not A168) );
 a90295a <=( A169  and  a90294a );
 a90298a <=( A199  and  A166 );
 a90301a <=( A201  and  (not A200) );
 a90302a <=( a90301a  and  a90298a );
 a90303a <=( a90302a  and  a90295a );
 a90306a <=( A232  and  A203 );
 a90309a <=( (not A265)  and  A233 );
 a90310a <=( a90309a  and  a90306a );
 a90313a <=( (not A299)  and  (not A266) );
 a90316a <=( (not A302)  and  (not A301) );
 a90317a <=( a90316a  and  a90313a );
 a90318a <=( a90317a  and  a90310a );
 a90322a <=( (not A167)  and  (not A168) );
 a90323a <=( A169  and  a90322a );
 a90326a <=( A199  and  A166 );
 a90329a <=( A201  and  (not A200) );
 a90330a <=( a90329a  and  a90326a );
 a90331a <=( a90330a  and  a90323a );
 a90334a <=( (not A233)  and  A203 );
 a90337a <=( (not A236)  and  (not A235) );
 a90338a <=( a90337a  and  a90334a );
 a90341a <=( A266  and  A265 );
 a90344a <=( (not A300)  and  A298 );
 a90345a <=( a90344a  and  a90341a );
 a90346a <=( a90345a  and  a90338a );
 a90350a <=( (not A167)  and  (not A168) );
 a90351a <=( A169  and  a90350a );
 a90354a <=( A199  and  A166 );
 a90357a <=( A201  and  (not A200) );
 a90358a <=( a90357a  and  a90354a );
 a90359a <=( a90358a  and  a90351a );
 a90362a <=( (not A233)  and  A203 );
 a90365a <=( (not A236)  and  (not A235) );
 a90366a <=( a90365a  and  a90362a );
 a90369a <=( A266  and  A265 );
 a90372a <=( A299  and  A298 );
 a90373a <=( a90372a  and  a90369a );
 a90374a <=( a90373a  and  a90366a );
 a90378a <=( (not A167)  and  (not A168) );
 a90379a <=( A169  and  a90378a );
 a90382a <=( A199  and  A166 );
 a90385a <=( A201  and  (not A200) );
 a90386a <=( a90385a  and  a90382a );
 a90387a <=( a90386a  and  a90379a );
 a90390a <=( (not A233)  and  A203 );
 a90393a <=( (not A236)  and  (not A235) );
 a90394a <=( a90393a  and  a90390a );
 a90397a <=( A266  and  A265 );
 a90400a <=( (not A299)  and  (not A298) );
 a90401a <=( a90400a  and  a90397a );
 a90402a <=( a90401a  and  a90394a );
 a90406a <=( (not A167)  and  (not A168) );
 a90407a <=( A169  and  a90406a );
 a90410a <=( A199  and  A166 );
 a90413a <=( A201  and  (not A200) );
 a90414a <=( a90413a  and  a90410a );
 a90415a <=( a90414a  and  a90407a );
 a90418a <=( (not A233)  and  A203 );
 a90421a <=( (not A236)  and  (not A235) );
 a90422a <=( a90421a  and  a90418a );
 a90425a <=( (not A267)  and  (not A266) );
 a90428a <=( (not A300)  and  A298 );
 a90429a <=( a90428a  and  a90425a );
 a90430a <=( a90429a  and  a90422a );
 a90434a <=( (not A167)  and  (not A168) );
 a90435a <=( A169  and  a90434a );
 a90438a <=( A199  and  A166 );
 a90441a <=( A201  and  (not A200) );
 a90442a <=( a90441a  and  a90438a );
 a90443a <=( a90442a  and  a90435a );
 a90446a <=( (not A233)  and  A203 );
 a90449a <=( (not A236)  and  (not A235) );
 a90450a <=( a90449a  and  a90446a );
 a90453a <=( (not A267)  and  (not A266) );
 a90456a <=( A299  and  A298 );
 a90457a <=( a90456a  and  a90453a );
 a90458a <=( a90457a  and  a90450a );
 a90462a <=( (not A167)  and  (not A168) );
 a90463a <=( A169  and  a90462a );
 a90466a <=( A199  and  A166 );
 a90469a <=( A201  and  (not A200) );
 a90470a <=( a90469a  and  a90466a );
 a90471a <=( a90470a  and  a90463a );
 a90474a <=( (not A233)  and  A203 );
 a90477a <=( (not A236)  and  (not A235) );
 a90478a <=( a90477a  and  a90474a );
 a90481a <=( (not A267)  and  (not A266) );
 a90484a <=( (not A299)  and  (not A298) );
 a90485a <=( a90484a  and  a90481a );
 a90486a <=( a90485a  and  a90478a );
 a90490a <=( (not A167)  and  (not A168) );
 a90491a <=( A169  and  a90490a );
 a90494a <=( A199  and  A166 );
 a90497a <=( A201  and  (not A200) );
 a90498a <=( a90497a  and  a90494a );
 a90499a <=( a90498a  and  a90491a );
 a90502a <=( (not A233)  and  A203 );
 a90505a <=( (not A236)  and  (not A235) );
 a90506a <=( a90505a  and  a90502a );
 a90509a <=( (not A266)  and  (not A265) );
 a90512a <=( (not A300)  and  A298 );
 a90513a <=( a90512a  and  a90509a );
 a90514a <=( a90513a  and  a90506a );
 a90518a <=( (not A167)  and  (not A168) );
 a90519a <=( A169  and  a90518a );
 a90522a <=( A199  and  A166 );
 a90525a <=( A201  and  (not A200) );
 a90526a <=( a90525a  and  a90522a );
 a90527a <=( a90526a  and  a90519a );
 a90530a <=( (not A233)  and  A203 );
 a90533a <=( (not A236)  and  (not A235) );
 a90534a <=( a90533a  and  a90530a );
 a90537a <=( (not A266)  and  (not A265) );
 a90540a <=( A299  and  A298 );
 a90541a <=( a90540a  and  a90537a );
 a90542a <=( a90541a  and  a90534a );
 a90546a <=( (not A167)  and  (not A168) );
 a90547a <=( A169  and  a90546a );
 a90550a <=( A199  and  A166 );
 a90553a <=( A201  and  (not A200) );
 a90554a <=( a90553a  and  a90550a );
 a90555a <=( a90554a  and  a90547a );
 a90558a <=( (not A233)  and  A203 );
 a90561a <=( (not A236)  and  (not A235) );
 a90562a <=( a90561a  and  a90558a );
 a90565a <=( (not A266)  and  (not A265) );
 a90568a <=( (not A299)  and  (not A298) );
 a90569a <=( a90568a  and  a90565a );
 a90570a <=( a90569a  and  a90562a );
 a90574a <=( (not A167)  and  (not A168) );
 a90575a <=( A169  and  a90574a );
 a90578a <=( A199  and  A166 );
 a90581a <=( A201  and  (not A200) );
 a90582a <=( a90581a  and  a90578a );
 a90583a <=( a90582a  and  a90575a );
 a90586a <=( (not A233)  and  A203 );
 a90589a <=( A265  and  (not A234) );
 a90590a <=( a90589a  and  a90586a );
 a90593a <=( A298  and  A266 );
 a90596a <=( (not A302)  and  (not A301) );
 a90597a <=( a90596a  and  a90593a );
 a90598a <=( a90597a  and  a90590a );
 a90602a <=( (not A167)  and  (not A168) );
 a90603a <=( A169  and  a90602a );
 a90606a <=( A199  and  A166 );
 a90609a <=( A201  and  (not A200) );
 a90610a <=( a90609a  and  a90606a );
 a90611a <=( a90610a  and  a90603a );
 a90614a <=( (not A233)  and  A203 );
 a90617a <=( (not A266)  and  (not A234) );
 a90618a <=( a90617a  and  a90614a );
 a90621a <=( (not A269)  and  (not A268) );
 a90624a <=( (not A300)  and  A298 );
 a90625a <=( a90624a  and  a90621a );
 a90626a <=( a90625a  and  a90618a );
 a90630a <=( (not A167)  and  (not A168) );
 a90631a <=( A169  and  a90630a );
 a90634a <=( A199  and  A166 );
 a90637a <=( A201  and  (not A200) );
 a90638a <=( a90637a  and  a90634a );
 a90639a <=( a90638a  and  a90631a );
 a90642a <=( (not A233)  and  A203 );
 a90645a <=( (not A266)  and  (not A234) );
 a90646a <=( a90645a  and  a90642a );
 a90649a <=( (not A269)  and  (not A268) );
 a90652a <=( A299  and  A298 );
 a90653a <=( a90652a  and  a90649a );
 a90654a <=( a90653a  and  a90646a );
 a90658a <=( (not A167)  and  (not A168) );
 a90659a <=( A169  and  a90658a );
 a90662a <=( A199  and  A166 );
 a90665a <=( A201  and  (not A200) );
 a90666a <=( a90665a  and  a90662a );
 a90667a <=( a90666a  and  a90659a );
 a90670a <=( (not A233)  and  A203 );
 a90673a <=( (not A266)  and  (not A234) );
 a90674a <=( a90673a  and  a90670a );
 a90677a <=( (not A269)  and  (not A268) );
 a90680a <=( (not A299)  and  (not A298) );
 a90681a <=( a90680a  and  a90677a );
 a90682a <=( a90681a  and  a90674a );
 a90686a <=( (not A167)  and  (not A168) );
 a90687a <=( A169  and  a90686a );
 a90690a <=( A199  and  A166 );
 a90693a <=( A201  and  (not A200) );
 a90694a <=( a90693a  and  a90690a );
 a90695a <=( a90694a  and  a90687a );
 a90698a <=( (not A233)  and  A203 );
 a90701a <=( (not A266)  and  (not A234) );
 a90702a <=( a90701a  and  a90698a );
 a90705a <=( A298  and  (not A267) );
 a90708a <=( (not A302)  and  (not A301) );
 a90709a <=( a90708a  and  a90705a );
 a90710a <=( a90709a  and  a90702a );
 a90714a <=( (not A167)  and  (not A168) );
 a90715a <=( A169  and  a90714a );
 a90718a <=( A199  and  A166 );
 a90721a <=( A201  and  (not A200) );
 a90722a <=( a90721a  and  a90718a );
 a90723a <=( a90722a  and  a90715a );
 a90726a <=( (not A233)  and  A203 );
 a90729a <=( (not A265)  and  (not A234) );
 a90730a <=( a90729a  and  a90726a );
 a90733a <=( A298  and  (not A266) );
 a90736a <=( (not A302)  and  (not A301) );
 a90737a <=( a90736a  and  a90733a );
 a90738a <=( a90737a  and  a90730a );
 a90742a <=( (not A167)  and  (not A168) );
 a90743a <=( A169  and  a90742a );
 a90746a <=( A199  and  A166 );
 a90749a <=( A201  and  (not A200) );
 a90750a <=( a90749a  and  a90746a );
 a90751a <=( a90750a  and  a90743a );
 a90754a <=( (not A232)  and  A203 );
 a90757a <=( A265  and  (not A233) );
 a90758a <=( a90757a  and  a90754a );
 a90761a <=( A298  and  A266 );
 a90764a <=( (not A302)  and  (not A301) );
 a90765a <=( a90764a  and  a90761a );
 a90766a <=( a90765a  and  a90758a );
 a90770a <=( (not A167)  and  (not A168) );
 a90771a <=( A169  and  a90770a );
 a90774a <=( A199  and  A166 );
 a90777a <=( A201  and  (not A200) );
 a90778a <=( a90777a  and  a90774a );
 a90779a <=( a90778a  and  a90771a );
 a90782a <=( (not A232)  and  A203 );
 a90785a <=( (not A266)  and  (not A233) );
 a90786a <=( a90785a  and  a90782a );
 a90789a <=( (not A269)  and  (not A268) );
 a90792a <=( (not A300)  and  A298 );
 a90793a <=( a90792a  and  a90789a );
 a90794a <=( a90793a  and  a90786a );
 a90798a <=( (not A167)  and  (not A168) );
 a90799a <=( A169  and  a90798a );
 a90802a <=( A199  and  A166 );
 a90805a <=( A201  and  (not A200) );
 a90806a <=( a90805a  and  a90802a );
 a90807a <=( a90806a  and  a90799a );
 a90810a <=( (not A232)  and  A203 );
 a90813a <=( (not A266)  and  (not A233) );
 a90814a <=( a90813a  and  a90810a );
 a90817a <=( (not A269)  and  (not A268) );
 a90820a <=( A299  and  A298 );
 a90821a <=( a90820a  and  a90817a );
 a90822a <=( a90821a  and  a90814a );
 a90826a <=( (not A167)  and  (not A168) );
 a90827a <=( A169  and  a90826a );
 a90830a <=( A199  and  A166 );
 a90833a <=( A201  and  (not A200) );
 a90834a <=( a90833a  and  a90830a );
 a90835a <=( a90834a  and  a90827a );
 a90838a <=( (not A232)  and  A203 );
 a90841a <=( (not A266)  and  (not A233) );
 a90842a <=( a90841a  and  a90838a );
 a90845a <=( (not A269)  and  (not A268) );
 a90848a <=( (not A299)  and  (not A298) );
 a90849a <=( a90848a  and  a90845a );
 a90850a <=( a90849a  and  a90842a );
 a90854a <=( (not A167)  and  (not A168) );
 a90855a <=( A169  and  a90854a );
 a90858a <=( A199  and  A166 );
 a90861a <=( A201  and  (not A200) );
 a90862a <=( a90861a  and  a90858a );
 a90863a <=( a90862a  and  a90855a );
 a90866a <=( (not A232)  and  A203 );
 a90869a <=( (not A266)  and  (not A233) );
 a90870a <=( a90869a  and  a90866a );
 a90873a <=( A298  and  (not A267) );
 a90876a <=( (not A302)  and  (not A301) );
 a90877a <=( a90876a  and  a90873a );
 a90878a <=( a90877a  and  a90870a );
 a90882a <=( (not A167)  and  (not A168) );
 a90883a <=( A169  and  a90882a );
 a90886a <=( A199  and  A166 );
 a90889a <=( A201  and  (not A200) );
 a90890a <=( a90889a  and  a90886a );
 a90891a <=( a90890a  and  a90883a );
 a90894a <=( (not A232)  and  A203 );
 a90897a <=( (not A265)  and  (not A233) );
 a90898a <=( a90897a  and  a90894a );
 a90901a <=( A298  and  (not A266) );
 a90904a <=( (not A302)  and  (not A301) );
 a90905a <=( a90904a  and  a90901a );
 a90906a <=( a90905a  and  a90898a );
 a90910a <=( (not A168)  and  A169 );
 a90911a <=( A170  and  a90910a );
 a90914a <=( (not A200)  and  A199 );
 a90917a <=( A202  and  A201 );
 a90918a <=( a90917a  and  a90914a );
 a90919a <=( a90918a  and  a90911a );
 a90922a <=( A233  and  A232 );
 a90925a <=( (not A268)  and  A265 );
 a90926a <=( a90925a  and  a90922a );
 a90929a <=( (not A299)  and  (not A269) );
 a90932a <=( (not A302)  and  (not A301) );
 a90933a <=( a90932a  and  a90929a );
 a90934a <=( a90933a  and  a90926a );
 a90938a <=( (not A168)  and  A169 );
 a90939a <=( A170  and  a90938a );
 a90942a <=( (not A200)  and  A199 );
 a90945a <=( A202  and  A201 );
 a90946a <=( a90945a  and  a90942a );
 a90947a <=( a90946a  and  a90939a );
 a90950a <=( (not A235)  and  (not A233) );
 a90953a <=( A265  and  (not A236) );
 a90954a <=( a90953a  and  a90950a );
 a90957a <=( A298  and  A266 );
 a90960a <=( (not A302)  and  (not A301) );
 a90961a <=( a90960a  and  a90957a );
 a90962a <=( a90961a  and  a90954a );
 a90966a <=( (not A168)  and  A169 );
 a90967a <=( A170  and  a90966a );
 a90970a <=( (not A200)  and  A199 );
 a90973a <=( A202  and  A201 );
 a90974a <=( a90973a  and  a90970a );
 a90975a <=( a90974a  and  a90967a );
 a90978a <=( (not A235)  and  (not A233) );
 a90981a <=( (not A266)  and  (not A236) );
 a90982a <=( a90981a  and  a90978a );
 a90985a <=( (not A269)  and  (not A268) );
 a90988a <=( (not A300)  and  A298 );
 a90989a <=( a90988a  and  a90985a );
 a90990a <=( a90989a  and  a90982a );
 a90994a <=( (not A168)  and  A169 );
 a90995a <=( A170  and  a90994a );
 a90998a <=( (not A200)  and  A199 );
 a91001a <=( A202  and  A201 );
 a91002a <=( a91001a  and  a90998a );
 a91003a <=( a91002a  and  a90995a );
 a91006a <=( (not A235)  and  (not A233) );
 a91009a <=( (not A266)  and  (not A236) );
 a91010a <=( a91009a  and  a91006a );
 a91013a <=( (not A269)  and  (not A268) );
 a91016a <=( A299  and  A298 );
 a91017a <=( a91016a  and  a91013a );
 a91018a <=( a91017a  and  a91010a );
 a91022a <=( (not A168)  and  A169 );
 a91023a <=( A170  and  a91022a );
 a91026a <=( (not A200)  and  A199 );
 a91029a <=( A202  and  A201 );
 a91030a <=( a91029a  and  a91026a );
 a91031a <=( a91030a  and  a91023a );
 a91034a <=( (not A235)  and  (not A233) );
 a91037a <=( (not A266)  and  (not A236) );
 a91038a <=( a91037a  and  a91034a );
 a91041a <=( (not A269)  and  (not A268) );
 a91044a <=( (not A299)  and  (not A298) );
 a91045a <=( a91044a  and  a91041a );
 a91046a <=( a91045a  and  a91038a );
 a91050a <=( (not A168)  and  A169 );
 a91051a <=( A170  and  a91050a );
 a91054a <=( (not A200)  and  A199 );
 a91057a <=( A202  and  A201 );
 a91058a <=( a91057a  and  a91054a );
 a91059a <=( a91058a  and  a91051a );
 a91062a <=( (not A235)  and  (not A233) );
 a91065a <=( (not A266)  and  (not A236) );
 a91066a <=( a91065a  and  a91062a );
 a91069a <=( A298  and  (not A267) );
 a91072a <=( (not A302)  and  (not A301) );
 a91073a <=( a91072a  and  a91069a );
 a91074a <=( a91073a  and  a91066a );
 a91078a <=( (not A168)  and  A169 );
 a91079a <=( A170  and  a91078a );
 a91082a <=( (not A200)  and  A199 );
 a91085a <=( A202  and  A201 );
 a91086a <=( a91085a  and  a91082a );
 a91087a <=( a91086a  and  a91079a );
 a91090a <=( (not A235)  and  (not A233) );
 a91093a <=( (not A265)  and  (not A236) );
 a91094a <=( a91093a  and  a91090a );
 a91097a <=( A298  and  (not A266) );
 a91100a <=( (not A302)  and  (not A301) );
 a91101a <=( a91100a  and  a91097a );
 a91102a <=( a91101a  and  a91094a );
 a91106a <=( (not A168)  and  A169 );
 a91107a <=( A170  and  a91106a );
 a91110a <=( (not A200)  and  A199 );
 a91113a <=( A202  and  A201 );
 a91114a <=( a91113a  and  a91110a );
 a91115a <=( a91114a  and  a91107a );
 a91118a <=( (not A234)  and  (not A233) );
 a91121a <=( (not A268)  and  (not A266) );
 a91122a <=( a91121a  and  a91118a );
 a91125a <=( A298  and  (not A269) );
 a91128a <=( (not A302)  and  (not A301) );
 a91129a <=( a91128a  and  a91125a );
 a91130a <=( a91129a  and  a91122a );
 a91134a <=( (not A168)  and  A169 );
 a91135a <=( A170  and  a91134a );
 a91138a <=( (not A200)  and  A199 );
 a91141a <=( A202  and  A201 );
 a91142a <=( a91141a  and  a91138a );
 a91143a <=( a91142a  and  a91135a );
 a91146a <=( (not A233)  and  A232 );
 a91149a <=( A235  and  A234 );
 a91150a <=( a91149a  and  a91146a );
 a91153a <=( (not A299)  and  A298 );
 a91156a <=( A301  and  A300 );
 a91157a <=( a91156a  and  a91153a );
 a91158a <=( a91157a  and  a91150a );
 a91162a <=( (not A168)  and  A169 );
 a91163a <=( A170  and  a91162a );
 a91166a <=( (not A200)  and  A199 );
 a91169a <=( A202  and  A201 );
 a91170a <=( a91169a  and  a91166a );
 a91171a <=( a91170a  and  a91163a );
 a91174a <=( (not A233)  and  A232 );
 a91177a <=( A235  and  A234 );
 a91178a <=( a91177a  and  a91174a );
 a91181a <=( (not A299)  and  A298 );
 a91184a <=( A302  and  A300 );
 a91185a <=( a91184a  and  a91181a );
 a91186a <=( a91185a  and  a91178a );
 a91190a <=( (not A168)  and  A169 );
 a91191a <=( A170  and  a91190a );
 a91194a <=( (not A200)  and  A199 );
 a91197a <=( A202  and  A201 );
 a91198a <=( a91197a  and  a91194a );
 a91199a <=( a91198a  and  a91191a );
 a91202a <=( (not A233)  and  A232 );
 a91205a <=( A235  and  A234 );
 a91206a <=( a91205a  and  a91202a );
 a91209a <=( (not A266)  and  A265 );
 a91212a <=( A268  and  A267 );
 a91213a <=( a91212a  and  a91209a );
 a91214a <=( a91213a  and  a91206a );
 a91218a <=( (not A168)  and  A169 );
 a91219a <=( A170  and  a91218a );
 a91222a <=( (not A200)  and  A199 );
 a91225a <=( A202  and  A201 );
 a91226a <=( a91225a  and  a91222a );
 a91227a <=( a91226a  and  a91219a );
 a91230a <=( (not A233)  and  A232 );
 a91233a <=( A235  and  A234 );
 a91234a <=( a91233a  and  a91230a );
 a91237a <=( (not A266)  and  A265 );
 a91240a <=( A269  and  A267 );
 a91241a <=( a91240a  and  a91237a );
 a91242a <=( a91241a  and  a91234a );
 a91246a <=( (not A168)  and  A169 );
 a91247a <=( A170  and  a91246a );
 a91250a <=( (not A200)  and  A199 );
 a91253a <=( A202  and  A201 );
 a91254a <=( a91253a  and  a91250a );
 a91255a <=( a91254a  and  a91247a );
 a91258a <=( (not A233)  and  A232 );
 a91261a <=( A236  and  A234 );
 a91262a <=( a91261a  and  a91258a );
 a91265a <=( (not A299)  and  A298 );
 a91268a <=( A301  and  A300 );
 a91269a <=( a91268a  and  a91265a );
 a91270a <=( a91269a  and  a91262a );
 a91274a <=( (not A168)  and  A169 );
 a91275a <=( A170  and  a91274a );
 a91278a <=( (not A200)  and  A199 );
 a91281a <=( A202  and  A201 );
 a91282a <=( a91281a  and  a91278a );
 a91283a <=( a91282a  and  a91275a );
 a91286a <=( (not A233)  and  A232 );
 a91289a <=( A236  and  A234 );
 a91290a <=( a91289a  and  a91286a );
 a91293a <=( (not A299)  and  A298 );
 a91296a <=( A302  and  A300 );
 a91297a <=( a91296a  and  a91293a );
 a91298a <=( a91297a  and  a91290a );
 a91302a <=( (not A168)  and  A169 );
 a91303a <=( A170  and  a91302a );
 a91306a <=( (not A200)  and  A199 );
 a91309a <=( A202  and  A201 );
 a91310a <=( a91309a  and  a91306a );
 a91311a <=( a91310a  and  a91303a );
 a91314a <=( (not A233)  and  A232 );
 a91317a <=( A236  and  A234 );
 a91318a <=( a91317a  and  a91314a );
 a91321a <=( (not A266)  and  A265 );
 a91324a <=( A268  and  A267 );
 a91325a <=( a91324a  and  a91321a );
 a91326a <=( a91325a  and  a91318a );
 a91330a <=( (not A168)  and  A169 );
 a91331a <=( A170  and  a91330a );
 a91334a <=( (not A200)  and  A199 );
 a91337a <=( A202  and  A201 );
 a91338a <=( a91337a  and  a91334a );
 a91339a <=( a91338a  and  a91331a );
 a91342a <=( (not A233)  and  A232 );
 a91345a <=( A236  and  A234 );
 a91346a <=( a91345a  and  a91342a );
 a91349a <=( (not A266)  and  A265 );
 a91352a <=( A269  and  A267 );
 a91353a <=( a91352a  and  a91349a );
 a91354a <=( a91353a  and  a91346a );
 a91358a <=( (not A168)  and  A169 );
 a91359a <=( A170  and  a91358a );
 a91362a <=( (not A200)  and  A199 );
 a91365a <=( A202  and  A201 );
 a91366a <=( a91365a  and  a91362a );
 a91367a <=( a91366a  and  a91359a );
 a91370a <=( (not A233)  and  (not A232) );
 a91373a <=( (not A268)  and  (not A266) );
 a91374a <=( a91373a  and  a91370a );
 a91377a <=( A298  and  (not A269) );
 a91380a <=( (not A302)  and  (not A301) );
 a91381a <=( a91380a  and  a91377a );
 a91382a <=( a91381a  and  a91374a );
 a91386a <=( (not A168)  and  A169 );
 a91387a <=( A170  and  a91386a );
 a91390a <=( (not A200)  and  A199 );
 a91393a <=( A203  and  A201 );
 a91394a <=( a91393a  and  a91390a );
 a91395a <=( a91394a  and  a91387a );
 a91398a <=( A233  and  A232 );
 a91401a <=( (not A268)  and  A265 );
 a91402a <=( a91401a  and  a91398a );
 a91405a <=( (not A299)  and  (not A269) );
 a91408a <=( (not A302)  and  (not A301) );
 a91409a <=( a91408a  and  a91405a );
 a91410a <=( a91409a  and  a91402a );
 a91414a <=( (not A168)  and  A169 );
 a91415a <=( A170  and  a91414a );
 a91418a <=( (not A200)  and  A199 );
 a91421a <=( A203  and  A201 );
 a91422a <=( a91421a  and  a91418a );
 a91423a <=( a91422a  and  a91415a );
 a91426a <=( (not A235)  and  (not A233) );
 a91429a <=( A265  and  (not A236) );
 a91430a <=( a91429a  and  a91426a );
 a91433a <=( A298  and  A266 );
 a91436a <=( (not A302)  and  (not A301) );
 a91437a <=( a91436a  and  a91433a );
 a91438a <=( a91437a  and  a91430a );
 a91442a <=( (not A168)  and  A169 );
 a91443a <=( A170  and  a91442a );
 a91446a <=( (not A200)  and  A199 );
 a91449a <=( A203  and  A201 );
 a91450a <=( a91449a  and  a91446a );
 a91451a <=( a91450a  and  a91443a );
 a91454a <=( (not A235)  and  (not A233) );
 a91457a <=( (not A266)  and  (not A236) );
 a91458a <=( a91457a  and  a91454a );
 a91461a <=( (not A269)  and  (not A268) );
 a91464a <=( (not A300)  and  A298 );
 a91465a <=( a91464a  and  a91461a );
 a91466a <=( a91465a  and  a91458a );
 a91470a <=( (not A168)  and  A169 );
 a91471a <=( A170  and  a91470a );
 a91474a <=( (not A200)  and  A199 );
 a91477a <=( A203  and  A201 );
 a91478a <=( a91477a  and  a91474a );
 a91479a <=( a91478a  and  a91471a );
 a91482a <=( (not A235)  and  (not A233) );
 a91485a <=( (not A266)  and  (not A236) );
 a91486a <=( a91485a  and  a91482a );
 a91489a <=( (not A269)  and  (not A268) );
 a91492a <=( A299  and  A298 );
 a91493a <=( a91492a  and  a91489a );
 a91494a <=( a91493a  and  a91486a );
 a91498a <=( (not A168)  and  A169 );
 a91499a <=( A170  and  a91498a );
 a91502a <=( (not A200)  and  A199 );
 a91505a <=( A203  and  A201 );
 a91506a <=( a91505a  and  a91502a );
 a91507a <=( a91506a  and  a91499a );
 a91510a <=( (not A235)  and  (not A233) );
 a91513a <=( (not A266)  and  (not A236) );
 a91514a <=( a91513a  and  a91510a );
 a91517a <=( (not A269)  and  (not A268) );
 a91520a <=( (not A299)  and  (not A298) );
 a91521a <=( a91520a  and  a91517a );
 a91522a <=( a91521a  and  a91514a );
 a91526a <=( (not A168)  and  A169 );
 a91527a <=( A170  and  a91526a );
 a91530a <=( (not A200)  and  A199 );
 a91533a <=( A203  and  A201 );
 a91534a <=( a91533a  and  a91530a );
 a91535a <=( a91534a  and  a91527a );
 a91538a <=( (not A235)  and  (not A233) );
 a91541a <=( (not A266)  and  (not A236) );
 a91542a <=( a91541a  and  a91538a );
 a91545a <=( A298  and  (not A267) );
 a91548a <=( (not A302)  and  (not A301) );
 a91549a <=( a91548a  and  a91545a );
 a91550a <=( a91549a  and  a91542a );
 a91554a <=( (not A168)  and  A169 );
 a91555a <=( A170  and  a91554a );
 a91558a <=( (not A200)  and  A199 );
 a91561a <=( A203  and  A201 );
 a91562a <=( a91561a  and  a91558a );
 a91563a <=( a91562a  and  a91555a );
 a91566a <=( (not A235)  and  (not A233) );
 a91569a <=( (not A265)  and  (not A236) );
 a91570a <=( a91569a  and  a91566a );
 a91573a <=( A298  and  (not A266) );
 a91576a <=( (not A302)  and  (not A301) );
 a91577a <=( a91576a  and  a91573a );
 a91578a <=( a91577a  and  a91570a );
 a91582a <=( (not A168)  and  A169 );
 a91583a <=( A170  and  a91582a );
 a91586a <=( (not A200)  and  A199 );
 a91589a <=( A203  and  A201 );
 a91590a <=( a91589a  and  a91586a );
 a91591a <=( a91590a  and  a91583a );
 a91594a <=( (not A234)  and  (not A233) );
 a91597a <=( (not A268)  and  (not A266) );
 a91598a <=( a91597a  and  a91594a );
 a91601a <=( A298  and  (not A269) );
 a91604a <=( (not A302)  and  (not A301) );
 a91605a <=( a91604a  and  a91601a );
 a91606a <=( a91605a  and  a91598a );
 a91610a <=( (not A168)  and  A169 );
 a91611a <=( A170  and  a91610a );
 a91614a <=( (not A200)  and  A199 );
 a91617a <=( A203  and  A201 );
 a91618a <=( a91617a  and  a91614a );
 a91619a <=( a91618a  and  a91611a );
 a91622a <=( (not A233)  and  A232 );
 a91625a <=( A235  and  A234 );
 a91626a <=( a91625a  and  a91622a );
 a91629a <=( (not A299)  and  A298 );
 a91632a <=( A301  and  A300 );
 a91633a <=( a91632a  and  a91629a );
 a91634a <=( a91633a  and  a91626a );
 a91638a <=( (not A168)  and  A169 );
 a91639a <=( A170  and  a91638a );
 a91642a <=( (not A200)  and  A199 );
 a91645a <=( A203  and  A201 );
 a91646a <=( a91645a  and  a91642a );
 a91647a <=( a91646a  and  a91639a );
 a91650a <=( (not A233)  and  A232 );
 a91653a <=( A235  and  A234 );
 a91654a <=( a91653a  and  a91650a );
 a91657a <=( (not A299)  and  A298 );
 a91660a <=( A302  and  A300 );
 a91661a <=( a91660a  and  a91657a );
 a91662a <=( a91661a  and  a91654a );
 a91666a <=( (not A168)  and  A169 );
 a91667a <=( A170  and  a91666a );
 a91670a <=( (not A200)  and  A199 );
 a91673a <=( A203  and  A201 );
 a91674a <=( a91673a  and  a91670a );
 a91675a <=( a91674a  and  a91667a );
 a91678a <=( (not A233)  and  A232 );
 a91681a <=( A235  and  A234 );
 a91682a <=( a91681a  and  a91678a );
 a91685a <=( (not A266)  and  A265 );
 a91688a <=( A268  and  A267 );
 a91689a <=( a91688a  and  a91685a );
 a91690a <=( a91689a  and  a91682a );
 a91694a <=( (not A168)  and  A169 );
 a91695a <=( A170  and  a91694a );
 a91698a <=( (not A200)  and  A199 );
 a91701a <=( A203  and  A201 );
 a91702a <=( a91701a  and  a91698a );
 a91703a <=( a91702a  and  a91695a );
 a91706a <=( (not A233)  and  A232 );
 a91709a <=( A235  and  A234 );
 a91710a <=( a91709a  and  a91706a );
 a91713a <=( (not A266)  and  A265 );
 a91716a <=( A269  and  A267 );
 a91717a <=( a91716a  and  a91713a );
 a91718a <=( a91717a  and  a91710a );
 a91722a <=( (not A168)  and  A169 );
 a91723a <=( A170  and  a91722a );
 a91726a <=( (not A200)  and  A199 );
 a91729a <=( A203  and  A201 );
 a91730a <=( a91729a  and  a91726a );
 a91731a <=( a91730a  and  a91723a );
 a91734a <=( (not A233)  and  A232 );
 a91737a <=( A236  and  A234 );
 a91738a <=( a91737a  and  a91734a );
 a91741a <=( (not A299)  and  A298 );
 a91744a <=( A301  and  A300 );
 a91745a <=( a91744a  and  a91741a );
 a91746a <=( a91745a  and  a91738a );
 a91750a <=( (not A168)  and  A169 );
 a91751a <=( A170  and  a91750a );
 a91754a <=( (not A200)  and  A199 );
 a91757a <=( A203  and  A201 );
 a91758a <=( a91757a  and  a91754a );
 a91759a <=( a91758a  and  a91751a );
 a91762a <=( (not A233)  and  A232 );
 a91765a <=( A236  and  A234 );
 a91766a <=( a91765a  and  a91762a );
 a91769a <=( (not A299)  and  A298 );
 a91772a <=( A302  and  A300 );
 a91773a <=( a91772a  and  a91769a );
 a91774a <=( a91773a  and  a91766a );
 a91778a <=( (not A168)  and  A169 );
 a91779a <=( A170  and  a91778a );
 a91782a <=( (not A200)  and  A199 );
 a91785a <=( A203  and  A201 );
 a91786a <=( a91785a  and  a91782a );
 a91787a <=( a91786a  and  a91779a );
 a91790a <=( (not A233)  and  A232 );
 a91793a <=( A236  and  A234 );
 a91794a <=( a91793a  and  a91790a );
 a91797a <=( (not A266)  and  A265 );
 a91800a <=( A268  and  A267 );
 a91801a <=( a91800a  and  a91797a );
 a91802a <=( a91801a  and  a91794a );
 a91806a <=( (not A168)  and  A169 );
 a91807a <=( A170  and  a91806a );
 a91810a <=( (not A200)  and  A199 );
 a91813a <=( A203  and  A201 );
 a91814a <=( a91813a  and  a91810a );
 a91815a <=( a91814a  and  a91807a );
 a91818a <=( (not A233)  and  A232 );
 a91821a <=( A236  and  A234 );
 a91822a <=( a91821a  and  a91818a );
 a91825a <=( (not A266)  and  A265 );
 a91828a <=( A269  and  A267 );
 a91829a <=( a91828a  and  a91825a );
 a91830a <=( a91829a  and  a91822a );
 a91834a <=( (not A168)  and  A169 );
 a91835a <=( A170  and  a91834a );
 a91838a <=( (not A200)  and  A199 );
 a91841a <=( A203  and  A201 );
 a91842a <=( a91841a  and  a91838a );
 a91843a <=( a91842a  and  a91835a );
 a91846a <=( (not A233)  and  (not A232) );
 a91849a <=( (not A268)  and  (not A266) );
 a91850a <=( a91849a  and  a91846a );
 a91853a <=( A298  and  (not A269) );
 a91856a <=( (not A302)  and  (not A301) );
 a91857a <=( a91856a  and  a91853a );
 a91858a <=( a91857a  and  a91850a );
 a91862a <=( A167  and  A169 );
 a91863a <=( (not A170)  and  a91862a );
 a91866a <=( A199  and  A166 );
 a91869a <=( (not A233)  and  A200 );
 a91870a <=( a91869a  and  a91866a );
 a91871a <=( a91870a  and  a91863a );
 a91874a <=( (not A236)  and  (not A235) );
 a91877a <=( (not A268)  and  (not A266) );
 a91878a <=( a91877a  and  a91874a );
 a91881a <=( A298  and  (not A269) );
 a91884a <=( (not A302)  and  (not A301) );
 a91885a <=( a91884a  and  a91881a );
 a91886a <=( a91885a  and  a91878a );
 a91890a <=( A167  and  A169 );
 a91891a <=( (not A170)  and  a91890a );
 a91894a <=( (not A200)  and  A166 );
 a91897a <=( (not A203)  and  (not A202) );
 a91898a <=( a91897a  and  a91894a );
 a91899a <=( a91898a  and  a91891a );
 a91902a <=( A233  and  A232 );
 a91905a <=( (not A268)  and  A265 );
 a91906a <=( a91905a  and  a91902a );
 a91909a <=( (not A299)  and  (not A269) );
 a91912a <=( (not A302)  and  (not A301) );
 a91913a <=( a91912a  and  a91909a );
 a91914a <=( a91913a  and  a91906a );
 a91918a <=( A167  and  A169 );
 a91919a <=( (not A170)  and  a91918a );
 a91922a <=( (not A200)  and  A166 );
 a91925a <=( (not A203)  and  (not A202) );
 a91926a <=( a91925a  and  a91922a );
 a91927a <=( a91926a  and  a91919a );
 a91930a <=( (not A235)  and  (not A233) );
 a91933a <=( A265  and  (not A236) );
 a91934a <=( a91933a  and  a91930a );
 a91937a <=( A298  and  A266 );
 a91940a <=( (not A302)  and  (not A301) );
 a91941a <=( a91940a  and  a91937a );
 a91942a <=( a91941a  and  a91934a );
 a91946a <=( A167  and  A169 );
 a91947a <=( (not A170)  and  a91946a );
 a91950a <=( (not A200)  and  A166 );
 a91953a <=( (not A203)  and  (not A202) );
 a91954a <=( a91953a  and  a91950a );
 a91955a <=( a91954a  and  a91947a );
 a91958a <=( (not A235)  and  (not A233) );
 a91961a <=( (not A266)  and  (not A236) );
 a91962a <=( a91961a  and  a91958a );
 a91965a <=( (not A269)  and  (not A268) );
 a91968a <=( (not A300)  and  A298 );
 a91969a <=( a91968a  and  a91965a );
 a91970a <=( a91969a  and  a91962a );
 a91974a <=( A167  and  A169 );
 a91975a <=( (not A170)  and  a91974a );
 a91978a <=( (not A200)  and  A166 );
 a91981a <=( (not A203)  and  (not A202) );
 a91982a <=( a91981a  and  a91978a );
 a91983a <=( a91982a  and  a91975a );
 a91986a <=( (not A235)  and  (not A233) );
 a91989a <=( (not A266)  and  (not A236) );
 a91990a <=( a91989a  and  a91986a );
 a91993a <=( (not A269)  and  (not A268) );
 a91996a <=( A299  and  A298 );
 a91997a <=( a91996a  and  a91993a );
 a91998a <=( a91997a  and  a91990a );
 a92002a <=( A167  and  A169 );
 a92003a <=( (not A170)  and  a92002a );
 a92006a <=( (not A200)  and  A166 );
 a92009a <=( (not A203)  and  (not A202) );
 a92010a <=( a92009a  and  a92006a );
 a92011a <=( a92010a  and  a92003a );
 a92014a <=( (not A235)  and  (not A233) );
 a92017a <=( (not A266)  and  (not A236) );
 a92018a <=( a92017a  and  a92014a );
 a92021a <=( (not A269)  and  (not A268) );
 a92024a <=( (not A299)  and  (not A298) );
 a92025a <=( a92024a  and  a92021a );
 a92026a <=( a92025a  and  a92018a );
 a92030a <=( A167  and  A169 );
 a92031a <=( (not A170)  and  a92030a );
 a92034a <=( (not A200)  and  A166 );
 a92037a <=( (not A203)  and  (not A202) );
 a92038a <=( a92037a  and  a92034a );
 a92039a <=( a92038a  and  a92031a );
 a92042a <=( (not A235)  and  (not A233) );
 a92045a <=( (not A266)  and  (not A236) );
 a92046a <=( a92045a  and  a92042a );
 a92049a <=( A298  and  (not A267) );
 a92052a <=( (not A302)  and  (not A301) );
 a92053a <=( a92052a  and  a92049a );
 a92054a <=( a92053a  and  a92046a );
 a92058a <=( A167  and  A169 );
 a92059a <=( (not A170)  and  a92058a );
 a92062a <=( (not A200)  and  A166 );
 a92065a <=( (not A203)  and  (not A202) );
 a92066a <=( a92065a  and  a92062a );
 a92067a <=( a92066a  and  a92059a );
 a92070a <=( (not A235)  and  (not A233) );
 a92073a <=( (not A265)  and  (not A236) );
 a92074a <=( a92073a  and  a92070a );
 a92077a <=( A298  and  (not A266) );
 a92080a <=( (not A302)  and  (not A301) );
 a92081a <=( a92080a  and  a92077a );
 a92082a <=( a92081a  and  a92074a );
 a92086a <=( A167  and  A169 );
 a92087a <=( (not A170)  and  a92086a );
 a92090a <=( (not A200)  and  A166 );
 a92093a <=( (not A203)  and  (not A202) );
 a92094a <=( a92093a  and  a92090a );
 a92095a <=( a92094a  and  a92087a );
 a92098a <=( (not A234)  and  (not A233) );
 a92101a <=( (not A268)  and  (not A266) );
 a92102a <=( a92101a  and  a92098a );
 a92105a <=( A298  and  (not A269) );
 a92108a <=( (not A302)  and  (not A301) );
 a92109a <=( a92108a  and  a92105a );
 a92110a <=( a92109a  and  a92102a );
 a92114a <=( A167  and  A169 );
 a92115a <=( (not A170)  and  a92114a );
 a92118a <=( (not A200)  and  A166 );
 a92121a <=( (not A203)  and  (not A202) );
 a92122a <=( a92121a  and  a92118a );
 a92123a <=( a92122a  and  a92115a );
 a92126a <=( (not A233)  and  A232 );
 a92129a <=( A235  and  A234 );
 a92130a <=( a92129a  and  a92126a );
 a92133a <=( (not A299)  and  A298 );
 a92136a <=( A301  and  A300 );
 a92137a <=( a92136a  and  a92133a );
 a92138a <=( a92137a  and  a92130a );
 a92142a <=( A167  and  A169 );
 a92143a <=( (not A170)  and  a92142a );
 a92146a <=( (not A200)  and  A166 );
 a92149a <=( (not A203)  and  (not A202) );
 a92150a <=( a92149a  and  a92146a );
 a92151a <=( a92150a  and  a92143a );
 a92154a <=( (not A233)  and  A232 );
 a92157a <=( A235  and  A234 );
 a92158a <=( a92157a  and  a92154a );
 a92161a <=( (not A299)  and  A298 );
 a92164a <=( A302  and  A300 );
 a92165a <=( a92164a  and  a92161a );
 a92166a <=( a92165a  and  a92158a );
 a92170a <=( A167  and  A169 );
 a92171a <=( (not A170)  and  a92170a );
 a92174a <=( (not A200)  and  A166 );
 a92177a <=( (not A203)  and  (not A202) );
 a92178a <=( a92177a  and  a92174a );
 a92179a <=( a92178a  and  a92171a );
 a92182a <=( (not A233)  and  A232 );
 a92185a <=( A235  and  A234 );
 a92186a <=( a92185a  and  a92182a );
 a92189a <=( (not A266)  and  A265 );
 a92192a <=( A268  and  A267 );
 a92193a <=( a92192a  and  a92189a );
 a92194a <=( a92193a  and  a92186a );
 a92198a <=( A167  and  A169 );
 a92199a <=( (not A170)  and  a92198a );
 a92202a <=( (not A200)  and  A166 );
 a92205a <=( (not A203)  and  (not A202) );
 a92206a <=( a92205a  and  a92202a );
 a92207a <=( a92206a  and  a92199a );
 a92210a <=( (not A233)  and  A232 );
 a92213a <=( A235  and  A234 );
 a92214a <=( a92213a  and  a92210a );
 a92217a <=( (not A266)  and  A265 );
 a92220a <=( A269  and  A267 );
 a92221a <=( a92220a  and  a92217a );
 a92222a <=( a92221a  and  a92214a );
 a92226a <=( A167  and  A169 );
 a92227a <=( (not A170)  and  a92226a );
 a92230a <=( (not A200)  and  A166 );
 a92233a <=( (not A203)  and  (not A202) );
 a92234a <=( a92233a  and  a92230a );
 a92235a <=( a92234a  and  a92227a );
 a92238a <=( (not A233)  and  A232 );
 a92241a <=( A236  and  A234 );
 a92242a <=( a92241a  and  a92238a );
 a92245a <=( (not A299)  and  A298 );
 a92248a <=( A301  and  A300 );
 a92249a <=( a92248a  and  a92245a );
 a92250a <=( a92249a  and  a92242a );
 a92254a <=( A167  and  A169 );
 a92255a <=( (not A170)  and  a92254a );
 a92258a <=( (not A200)  and  A166 );
 a92261a <=( (not A203)  and  (not A202) );
 a92262a <=( a92261a  and  a92258a );
 a92263a <=( a92262a  and  a92255a );
 a92266a <=( (not A233)  and  A232 );
 a92269a <=( A236  and  A234 );
 a92270a <=( a92269a  and  a92266a );
 a92273a <=( (not A299)  and  A298 );
 a92276a <=( A302  and  A300 );
 a92277a <=( a92276a  and  a92273a );
 a92278a <=( a92277a  and  a92270a );
 a92282a <=( A167  and  A169 );
 a92283a <=( (not A170)  and  a92282a );
 a92286a <=( (not A200)  and  A166 );
 a92289a <=( (not A203)  and  (not A202) );
 a92290a <=( a92289a  and  a92286a );
 a92291a <=( a92290a  and  a92283a );
 a92294a <=( (not A233)  and  A232 );
 a92297a <=( A236  and  A234 );
 a92298a <=( a92297a  and  a92294a );
 a92301a <=( (not A266)  and  A265 );
 a92304a <=( A268  and  A267 );
 a92305a <=( a92304a  and  a92301a );
 a92306a <=( a92305a  and  a92298a );
 a92310a <=( A167  and  A169 );
 a92311a <=( (not A170)  and  a92310a );
 a92314a <=( (not A200)  and  A166 );
 a92317a <=( (not A203)  and  (not A202) );
 a92318a <=( a92317a  and  a92314a );
 a92319a <=( a92318a  and  a92311a );
 a92322a <=( (not A233)  and  A232 );
 a92325a <=( A236  and  A234 );
 a92326a <=( a92325a  and  a92322a );
 a92329a <=( (not A266)  and  A265 );
 a92332a <=( A269  and  A267 );
 a92333a <=( a92332a  and  a92329a );
 a92334a <=( a92333a  and  a92326a );
 a92338a <=( A167  and  A169 );
 a92339a <=( (not A170)  and  a92338a );
 a92342a <=( (not A200)  and  A166 );
 a92345a <=( (not A203)  and  (not A202) );
 a92346a <=( a92345a  and  a92342a );
 a92347a <=( a92346a  and  a92339a );
 a92350a <=( (not A233)  and  (not A232) );
 a92353a <=( (not A268)  and  (not A266) );
 a92354a <=( a92353a  and  a92350a );
 a92357a <=( A298  and  (not A269) );
 a92360a <=( (not A302)  and  (not A301) );
 a92361a <=( a92360a  and  a92357a );
 a92362a <=( a92361a  and  a92354a );
 a92366a <=( A167  and  A169 );
 a92367a <=( (not A170)  and  a92366a );
 a92370a <=( (not A200)  and  A166 );
 a92373a <=( (not A233)  and  (not A201) );
 a92374a <=( a92373a  and  a92370a );
 a92375a <=( a92374a  and  a92367a );
 a92378a <=( (not A236)  and  (not A235) );
 a92381a <=( (not A268)  and  (not A266) );
 a92382a <=( a92381a  and  a92378a );
 a92385a <=( A298  and  (not A269) );
 a92388a <=( (not A302)  and  (not A301) );
 a92389a <=( a92388a  and  a92385a );
 a92390a <=( a92389a  and  a92382a );
 a92394a <=( A167  and  A169 );
 a92395a <=( (not A170)  and  a92394a );
 a92398a <=( (not A199)  and  A166 );
 a92401a <=( (not A233)  and  (not A200) );
 a92402a <=( a92401a  and  a92398a );
 a92403a <=( a92402a  and  a92395a );
 a92406a <=( (not A236)  and  (not A235) );
 a92409a <=( (not A268)  and  (not A266) );
 a92410a <=( a92409a  and  a92406a );
 a92413a <=( A298  and  (not A269) );
 a92416a <=( (not A302)  and  (not A301) );
 a92417a <=( a92416a  and  a92413a );
 a92418a <=( a92417a  and  a92410a );
 a92422a <=( (not A167)  and  A169 );
 a92423a <=( (not A170)  and  a92422a );
 a92426a <=( A199  and  (not A166) );
 a92429a <=( (not A233)  and  A200 );
 a92430a <=( a92429a  and  a92426a );
 a92431a <=( a92430a  and  a92423a );
 a92434a <=( (not A236)  and  (not A235) );
 a92437a <=( (not A268)  and  (not A266) );
 a92438a <=( a92437a  and  a92434a );
 a92441a <=( A298  and  (not A269) );
 a92444a <=( (not A302)  and  (not A301) );
 a92445a <=( a92444a  and  a92441a );
 a92446a <=( a92445a  and  a92438a );
 a92450a <=( (not A167)  and  A169 );
 a92451a <=( (not A170)  and  a92450a );
 a92454a <=( (not A200)  and  (not A166) );
 a92457a <=( (not A203)  and  (not A202) );
 a92458a <=( a92457a  and  a92454a );
 a92459a <=( a92458a  and  a92451a );
 a92462a <=( A233  and  A232 );
 a92465a <=( (not A268)  and  A265 );
 a92466a <=( a92465a  and  a92462a );
 a92469a <=( (not A299)  and  (not A269) );
 a92472a <=( (not A302)  and  (not A301) );
 a92473a <=( a92472a  and  a92469a );
 a92474a <=( a92473a  and  a92466a );
 a92478a <=( (not A167)  and  A169 );
 a92479a <=( (not A170)  and  a92478a );
 a92482a <=( (not A200)  and  (not A166) );
 a92485a <=( (not A203)  and  (not A202) );
 a92486a <=( a92485a  and  a92482a );
 a92487a <=( a92486a  and  a92479a );
 a92490a <=( (not A235)  and  (not A233) );
 a92493a <=( A265  and  (not A236) );
 a92494a <=( a92493a  and  a92490a );
 a92497a <=( A298  and  A266 );
 a92500a <=( (not A302)  and  (not A301) );
 a92501a <=( a92500a  and  a92497a );
 a92502a <=( a92501a  and  a92494a );
 a92506a <=( (not A167)  and  A169 );
 a92507a <=( (not A170)  and  a92506a );
 a92510a <=( (not A200)  and  (not A166) );
 a92513a <=( (not A203)  and  (not A202) );
 a92514a <=( a92513a  and  a92510a );
 a92515a <=( a92514a  and  a92507a );
 a92518a <=( (not A235)  and  (not A233) );
 a92521a <=( (not A266)  and  (not A236) );
 a92522a <=( a92521a  and  a92518a );
 a92525a <=( (not A269)  and  (not A268) );
 a92528a <=( (not A300)  and  A298 );
 a92529a <=( a92528a  and  a92525a );
 a92530a <=( a92529a  and  a92522a );
 a92534a <=( (not A167)  and  A169 );
 a92535a <=( (not A170)  and  a92534a );
 a92538a <=( (not A200)  and  (not A166) );
 a92541a <=( (not A203)  and  (not A202) );
 a92542a <=( a92541a  and  a92538a );
 a92543a <=( a92542a  and  a92535a );
 a92546a <=( (not A235)  and  (not A233) );
 a92549a <=( (not A266)  and  (not A236) );
 a92550a <=( a92549a  and  a92546a );
 a92553a <=( (not A269)  and  (not A268) );
 a92556a <=( A299  and  A298 );
 a92557a <=( a92556a  and  a92553a );
 a92558a <=( a92557a  and  a92550a );
 a92562a <=( (not A167)  and  A169 );
 a92563a <=( (not A170)  and  a92562a );
 a92566a <=( (not A200)  and  (not A166) );
 a92569a <=( (not A203)  and  (not A202) );
 a92570a <=( a92569a  and  a92566a );
 a92571a <=( a92570a  and  a92563a );
 a92574a <=( (not A235)  and  (not A233) );
 a92577a <=( (not A266)  and  (not A236) );
 a92578a <=( a92577a  and  a92574a );
 a92581a <=( (not A269)  and  (not A268) );
 a92584a <=( (not A299)  and  (not A298) );
 a92585a <=( a92584a  and  a92581a );
 a92586a <=( a92585a  and  a92578a );
 a92590a <=( (not A167)  and  A169 );
 a92591a <=( (not A170)  and  a92590a );
 a92594a <=( (not A200)  and  (not A166) );
 a92597a <=( (not A203)  and  (not A202) );
 a92598a <=( a92597a  and  a92594a );
 a92599a <=( a92598a  and  a92591a );
 a92602a <=( (not A235)  and  (not A233) );
 a92605a <=( (not A266)  and  (not A236) );
 a92606a <=( a92605a  and  a92602a );
 a92609a <=( A298  and  (not A267) );
 a92612a <=( (not A302)  and  (not A301) );
 a92613a <=( a92612a  and  a92609a );
 a92614a <=( a92613a  and  a92606a );
 a92618a <=( (not A167)  and  A169 );
 a92619a <=( (not A170)  and  a92618a );
 a92622a <=( (not A200)  and  (not A166) );
 a92625a <=( (not A203)  and  (not A202) );
 a92626a <=( a92625a  and  a92622a );
 a92627a <=( a92626a  and  a92619a );
 a92630a <=( (not A235)  and  (not A233) );
 a92633a <=( (not A265)  and  (not A236) );
 a92634a <=( a92633a  and  a92630a );
 a92637a <=( A298  and  (not A266) );
 a92640a <=( (not A302)  and  (not A301) );
 a92641a <=( a92640a  and  a92637a );
 a92642a <=( a92641a  and  a92634a );
 a92646a <=( (not A167)  and  A169 );
 a92647a <=( (not A170)  and  a92646a );
 a92650a <=( (not A200)  and  (not A166) );
 a92653a <=( (not A203)  and  (not A202) );
 a92654a <=( a92653a  and  a92650a );
 a92655a <=( a92654a  and  a92647a );
 a92658a <=( (not A234)  and  (not A233) );
 a92661a <=( (not A268)  and  (not A266) );
 a92662a <=( a92661a  and  a92658a );
 a92665a <=( A298  and  (not A269) );
 a92668a <=( (not A302)  and  (not A301) );
 a92669a <=( a92668a  and  a92665a );
 a92670a <=( a92669a  and  a92662a );
 a92674a <=( (not A167)  and  A169 );
 a92675a <=( (not A170)  and  a92674a );
 a92678a <=( (not A200)  and  (not A166) );
 a92681a <=( (not A203)  and  (not A202) );
 a92682a <=( a92681a  and  a92678a );
 a92683a <=( a92682a  and  a92675a );
 a92686a <=( (not A233)  and  A232 );
 a92689a <=( A235  and  A234 );
 a92690a <=( a92689a  and  a92686a );
 a92693a <=( (not A299)  and  A298 );
 a92696a <=( A301  and  A300 );
 a92697a <=( a92696a  and  a92693a );
 a92698a <=( a92697a  and  a92690a );
 a92702a <=( (not A167)  and  A169 );
 a92703a <=( (not A170)  and  a92702a );
 a92706a <=( (not A200)  and  (not A166) );
 a92709a <=( (not A203)  and  (not A202) );
 a92710a <=( a92709a  and  a92706a );
 a92711a <=( a92710a  and  a92703a );
 a92714a <=( (not A233)  and  A232 );
 a92717a <=( A235  and  A234 );
 a92718a <=( a92717a  and  a92714a );
 a92721a <=( (not A299)  and  A298 );
 a92724a <=( A302  and  A300 );
 a92725a <=( a92724a  and  a92721a );
 a92726a <=( a92725a  and  a92718a );
 a92730a <=( (not A167)  and  A169 );
 a92731a <=( (not A170)  and  a92730a );
 a92734a <=( (not A200)  and  (not A166) );
 a92737a <=( (not A203)  and  (not A202) );
 a92738a <=( a92737a  and  a92734a );
 a92739a <=( a92738a  and  a92731a );
 a92742a <=( (not A233)  and  A232 );
 a92745a <=( A235  and  A234 );
 a92746a <=( a92745a  and  a92742a );
 a92749a <=( (not A266)  and  A265 );
 a92752a <=( A268  and  A267 );
 a92753a <=( a92752a  and  a92749a );
 a92754a <=( a92753a  and  a92746a );
 a92758a <=( (not A167)  and  A169 );
 a92759a <=( (not A170)  and  a92758a );
 a92762a <=( (not A200)  and  (not A166) );
 a92765a <=( (not A203)  and  (not A202) );
 a92766a <=( a92765a  and  a92762a );
 a92767a <=( a92766a  and  a92759a );
 a92770a <=( (not A233)  and  A232 );
 a92773a <=( A235  and  A234 );
 a92774a <=( a92773a  and  a92770a );
 a92777a <=( (not A266)  and  A265 );
 a92780a <=( A269  and  A267 );
 a92781a <=( a92780a  and  a92777a );
 a92782a <=( a92781a  and  a92774a );
 a92786a <=( (not A167)  and  A169 );
 a92787a <=( (not A170)  and  a92786a );
 a92790a <=( (not A200)  and  (not A166) );
 a92793a <=( (not A203)  and  (not A202) );
 a92794a <=( a92793a  and  a92790a );
 a92795a <=( a92794a  and  a92787a );
 a92798a <=( (not A233)  and  A232 );
 a92801a <=( A236  and  A234 );
 a92802a <=( a92801a  and  a92798a );
 a92805a <=( (not A299)  and  A298 );
 a92808a <=( A301  and  A300 );
 a92809a <=( a92808a  and  a92805a );
 a92810a <=( a92809a  and  a92802a );
 a92814a <=( (not A167)  and  A169 );
 a92815a <=( (not A170)  and  a92814a );
 a92818a <=( (not A200)  and  (not A166) );
 a92821a <=( (not A203)  and  (not A202) );
 a92822a <=( a92821a  and  a92818a );
 a92823a <=( a92822a  and  a92815a );
 a92826a <=( (not A233)  and  A232 );
 a92829a <=( A236  and  A234 );
 a92830a <=( a92829a  and  a92826a );
 a92833a <=( (not A299)  and  A298 );
 a92836a <=( A302  and  A300 );
 a92837a <=( a92836a  and  a92833a );
 a92838a <=( a92837a  and  a92830a );
 a92842a <=( (not A167)  and  A169 );
 a92843a <=( (not A170)  and  a92842a );
 a92846a <=( (not A200)  and  (not A166) );
 a92849a <=( (not A203)  and  (not A202) );
 a92850a <=( a92849a  and  a92846a );
 a92851a <=( a92850a  and  a92843a );
 a92854a <=( (not A233)  and  A232 );
 a92857a <=( A236  and  A234 );
 a92858a <=( a92857a  and  a92854a );
 a92861a <=( (not A266)  and  A265 );
 a92864a <=( A268  and  A267 );
 a92865a <=( a92864a  and  a92861a );
 a92866a <=( a92865a  and  a92858a );
 a92870a <=( (not A167)  and  A169 );
 a92871a <=( (not A170)  and  a92870a );
 a92874a <=( (not A200)  and  (not A166) );
 a92877a <=( (not A203)  and  (not A202) );
 a92878a <=( a92877a  and  a92874a );
 a92879a <=( a92878a  and  a92871a );
 a92882a <=( (not A233)  and  A232 );
 a92885a <=( A236  and  A234 );
 a92886a <=( a92885a  and  a92882a );
 a92889a <=( (not A266)  and  A265 );
 a92892a <=( A269  and  A267 );
 a92893a <=( a92892a  and  a92889a );
 a92894a <=( a92893a  and  a92886a );
 a92898a <=( (not A167)  and  A169 );
 a92899a <=( (not A170)  and  a92898a );
 a92902a <=( (not A200)  and  (not A166) );
 a92905a <=( (not A203)  and  (not A202) );
 a92906a <=( a92905a  and  a92902a );
 a92907a <=( a92906a  and  a92899a );
 a92910a <=( (not A233)  and  (not A232) );
 a92913a <=( (not A268)  and  (not A266) );
 a92914a <=( a92913a  and  a92910a );
 a92917a <=( A298  and  (not A269) );
 a92920a <=( (not A302)  and  (not A301) );
 a92921a <=( a92920a  and  a92917a );
 a92922a <=( a92921a  and  a92914a );
 a92926a <=( (not A167)  and  A169 );
 a92927a <=( (not A170)  and  a92926a );
 a92930a <=( (not A200)  and  (not A166) );
 a92933a <=( (not A233)  and  (not A201) );
 a92934a <=( a92933a  and  a92930a );
 a92935a <=( a92934a  and  a92927a );
 a92938a <=( (not A236)  and  (not A235) );
 a92941a <=( (not A268)  and  (not A266) );
 a92942a <=( a92941a  and  a92938a );
 a92945a <=( A298  and  (not A269) );
 a92948a <=( (not A302)  and  (not A301) );
 a92949a <=( a92948a  and  a92945a );
 a92950a <=( a92949a  and  a92942a );
 a92954a <=( (not A167)  and  A169 );
 a92955a <=( (not A170)  and  a92954a );
 a92958a <=( (not A199)  and  (not A166) );
 a92961a <=( (not A233)  and  (not A200) );
 a92962a <=( a92961a  and  a92958a );
 a92963a <=( a92962a  and  a92955a );
 a92966a <=( (not A236)  and  (not A235) );
 a92969a <=( (not A268)  and  (not A266) );
 a92970a <=( a92969a  and  a92966a );
 a92973a <=( A298  and  (not A269) );
 a92976a <=( (not A302)  and  (not A301) );
 a92977a <=( a92976a  and  a92973a );
 a92978a <=( a92977a  and  a92970a );
 a92982a <=( (not A166)  and  (not A167) );
 a92983a <=( (not A169)  and  a92982a );
 a92986a <=( (not A200)  and  A199 );
 a92989a <=( A202  and  A201 );
 a92990a <=( a92989a  and  a92986a );
 a92991a <=( a92990a  and  a92983a );
 a92994a <=( A233  and  A232 );
 a92997a <=( (not A268)  and  A265 );
 a92998a <=( a92997a  and  a92994a );
 a93001a <=( (not A299)  and  (not A269) );
 a93004a <=( (not A302)  and  (not A301) );
 a93005a <=( a93004a  and  a93001a );
 a93006a <=( a93005a  and  a92998a );
 a93010a <=( (not A166)  and  (not A167) );
 a93011a <=( (not A169)  and  a93010a );
 a93014a <=( (not A200)  and  A199 );
 a93017a <=( A202  and  A201 );
 a93018a <=( a93017a  and  a93014a );
 a93019a <=( a93018a  and  a93011a );
 a93022a <=( (not A235)  and  (not A233) );
 a93025a <=( A265  and  (not A236) );
 a93026a <=( a93025a  and  a93022a );
 a93029a <=( A298  and  A266 );
 a93032a <=( (not A302)  and  (not A301) );
 a93033a <=( a93032a  and  a93029a );
 a93034a <=( a93033a  and  a93026a );
 a93038a <=( (not A166)  and  (not A167) );
 a93039a <=( (not A169)  and  a93038a );
 a93042a <=( (not A200)  and  A199 );
 a93045a <=( A202  and  A201 );
 a93046a <=( a93045a  and  a93042a );
 a93047a <=( a93046a  and  a93039a );
 a93050a <=( (not A235)  and  (not A233) );
 a93053a <=( (not A266)  and  (not A236) );
 a93054a <=( a93053a  and  a93050a );
 a93057a <=( (not A269)  and  (not A268) );
 a93060a <=( (not A300)  and  A298 );
 a93061a <=( a93060a  and  a93057a );
 a93062a <=( a93061a  and  a93054a );
 a93066a <=( (not A166)  and  (not A167) );
 a93067a <=( (not A169)  and  a93066a );
 a93070a <=( (not A200)  and  A199 );
 a93073a <=( A202  and  A201 );
 a93074a <=( a93073a  and  a93070a );
 a93075a <=( a93074a  and  a93067a );
 a93078a <=( (not A235)  and  (not A233) );
 a93081a <=( (not A266)  and  (not A236) );
 a93082a <=( a93081a  and  a93078a );
 a93085a <=( (not A269)  and  (not A268) );
 a93088a <=( A299  and  A298 );
 a93089a <=( a93088a  and  a93085a );
 a93090a <=( a93089a  and  a93082a );
 a93094a <=( (not A166)  and  (not A167) );
 a93095a <=( (not A169)  and  a93094a );
 a93098a <=( (not A200)  and  A199 );
 a93101a <=( A202  and  A201 );
 a93102a <=( a93101a  and  a93098a );
 a93103a <=( a93102a  and  a93095a );
 a93106a <=( (not A235)  and  (not A233) );
 a93109a <=( (not A266)  and  (not A236) );
 a93110a <=( a93109a  and  a93106a );
 a93113a <=( (not A269)  and  (not A268) );
 a93116a <=( (not A299)  and  (not A298) );
 a93117a <=( a93116a  and  a93113a );
 a93118a <=( a93117a  and  a93110a );
 a93122a <=( (not A166)  and  (not A167) );
 a93123a <=( (not A169)  and  a93122a );
 a93126a <=( (not A200)  and  A199 );
 a93129a <=( A202  and  A201 );
 a93130a <=( a93129a  and  a93126a );
 a93131a <=( a93130a  and  a93123a );
 a93134a <=( (not A235)  and  (not A233) );
 a93137a <=( (not A266)  and  (not A236) );
 a93138a <=( a93137a  and  a93134a );
 a93141a <=( A298  and  (not A267) );
 a93144a <=( (not A302)  and  (not A301) );
 a93145a <=( a93144a  and  a93141a );
 a93146a <=( a93145a  and  a93138a );
 a93150a <=( (not A166)  and  (not A167) );
 a93151a <=( (not A169)  and  a93150a );
 a93154a <=( (not A200)  and  A199 );
 a93157a <=( A202  and  A201 );
 a93158a <=( a93157a  and  a93154a );
 a93159a <=( a93158a  and  a93151a );
 a93162a <=( (not A235)  and  (not A233) );
 a93165a <=( (not A265)  and  (not A236) );
 a93166a <=( a93165a  and  a93162a );
 a93169a <=( A298  and  (not A266) );
 a93172a <=( (not A302)  and  (not A301) );
 a93173a <=( a93172a  and  a93169a );
 a93174a <=( a93173a  and  a93166a );
 a93178a <=( (not A166)  and  (not A167) );
 a93179a <=( (not A169)  and  a93178a );
 a93182a <=( (not A200)  and  A199 );
 a93185a <=( A202  and  A201 );
 a93186a <=( a93185a  and  a93182a );
 a93187a <=( a93186a  and  a93179a );
 a93190a <=( (not A234)  and  (not A233) );
 a93193a <=( (not A268)  and  (not A266) );
 a93194a <=( a93193a  and  a93190a );
 a93197a <=( A298  and  (not A269) );
 a93200a <=( (not A302)  and  (not A301) );
 a93201a <=( a93200a  and  a93197a );
 a93202a <=( a93201a  and  a93194a );
 a93206a <=( (not A166)  and  (not A167) );
 a93207a <=( (not A169)  and  a93206a );
 a93210a <=( (not A200)  and  A199 );
 a93213a <=( A202  and  A201 );
 a93214a <=( a93213a  and  a93210a );
 a93215a <=( a93214a  and  a93207a );
 a93218a <=( (not A233)  and  A232 );
 a93221a <=( A235  and  A234 );
 a93222a <=( a93221a  and  a93218a );
 a93225a <=( (not A299)  and  A298 );
 a93228a <=( A301  and  A300 );
 a93229a <=( a93228a  and  a93225a );
 a93230a <=( a93229a  and  a93222a );
 a93234a <=( (not A166)  and  (not A167) );
 a93235a <=( (not A169)  and  a93234a );
 a93238a <=( (not A200)  and  A199 );
 a93241a <=( A202  and  A201 );
 a93242a <=( a93241a  and  a93238a );
 a93243a <=( a93242a  and  a93235a );
 a93246a <=( (not A233)  and  A232 );
 a93249a <=( A235  and  A234 );
 a93250a <=( a93249a  and  a93246a );
 a93253a <=( (not A299)  and  A298 );
 a93256a <=( A302  and  A300 );
 a93257a <=( a93256a  and  a93253a );
 a93258a <=( a93257a  and  a93250a );
 a93262a <=( (not A166)  and  (not A167) );
 a93263a <=( (not A169)  and  a93262a );
 a93266a <=( (not A200)  and  A199 );
 a93269a <=( A202  and  A201 );
 a93270a <=( a93269a  and  a93266a );
 a93271a <=( a93270a  and  a93263a );
 a93274a <=( (not A233)  and  A232 );
 a93277a <=( A235  and  A234 );
 a93278a <=( a93277a  and  a93274a );
 a93281a <=( (not A266)  and  A265 );
 a93284a <=( A268  and  A267 );
 a93285a <=( a93284a  and  a93281a );
 a93286a <=( a93285a  and  a93278a );
 a93290a <=( (not A166)  and  (not A167) );
 a93291a <=( (not A169)  and  a93290a );
 a93294a <=( (not A200)  and  A199 );
 a93297a <=( A202  and  A201 );
 a93298a <=( a93297a  and  a93294a );
 a93299a <=( a93298a  and  a93291a );
 a93302a <=( (not A233)  and  A232 );
 a93305a <=( A235  and  A234 );
 a93306a <=( a93305a  and  a93302a );
 a93309a <=( (not A266)  and  A265 );
 a93312a <=( A269  and  A267 );
 a93313a <=( a93312a  and  a93309a );
 a93314a <=( a93313a  and  a93306a );
 a93318a <=( (not A166)  and  (not A167) );
 a93319a <=( (not A169)  and  a93318a );
 a93322a <=( (not A200)  and  A199 );
 a93325a <=( A202  and  A201 );
 a93326a <=( a93325a  and  a93322a );
 a93327a <=( a93326a  and  a93319a );
 a93330a <=( (not A233)  and  A232 );
 a93333a <=( A236  and  A234 );
 a93334a <=( a93333a  and  a93330a );
 a93337a <=( (not A299)  and  A298 );
 a93340a <=( A301  and  A300 );
 a93341a <=( a93340a  and  a93337a );
 a93342a <=( a93341a  and  a93334a );
 a93346a <=( (not A166)  and  (not A167) );
 a93347a <=( (not A169)  and  a93346a );
 a93350a <=( (not A200)  and  A199 );
 a93353a <=( A202  and  A201 );
 a93354a <=( a93353a  and  a93350a );
 a93355a <=( a93354a  and  a93347a );
 a93358a <=( (not A233)  and  A232 );
 a93361a <=( A236  and  A234 );
 a93362a <=( a93361a  and  a93358a );
 a93365a <=( (not A299)  and  A298 );
 a93368a <=( A302  and  A300 );
 a93369a <=( a93368a  and  a93365a );
 a93370a <=( a93369a  and  a93362a );
 a93374a <=( (not A166)  and  (not A167) );
 a93375a <=( (not A169)  and  a93374a );
 a93378a <=( (not A200)  and  A199 );
 a93381a <=( A202  and  A201 );
 a93382a <=( a93381a  and  a93378a );
 a93383a <=( a93382a  and  a93375a );
 a93386a <=( (not A233)  and  A232 );
 a93389a <=( A236  and  A234 );
 a93390a <=( a93389a  and  a93386a );
 a93393a <=( (not A266)  and  A265 );
 a93396a <=( A268  and  A267 );
 a93397a <=( a93396a  and  a93393a );
 a93398a <=( a93397a  and  a93390a );
 a93402a <=( (not A166)  and  (not A167) );
 a93403a <=( (not A169)  and  a93402a );
 a93406a <=( (not A200)  and  A199 );
 a93409a <=( A202  and  A201 );
 a93410a <=( a93409a  and  a93406a );
 a93411a <=( a93410a  and  a93403a );
 a93414a <=( (not A233)  and  A232 );
 a93417a <=( A236  and  A234 );
 a93418a <=( a93417a  and  a93414a );
 a93421a <=( (not A266)  and  A265 );
 a93424a <=( A269  and  A267 );
 a93425a <=( a93424a  and  a93421a );
 a93426a <=( a93425a  and  a93418a );
 a93430a <=( (not A166)  and  (not A167) );
 a93431a <=( (not A169)  and  a93430a );
 a93434a <=( (not A200)  and  A199 );
 a93437a <=( A202  and  A201 );
 a93438a <=( a93437a  and  a93434a );
 a93439a <=( a93438a  and  a93431a );
 a93442a <=( (not A233)  and  (not A232) );
 a93445a <=( (not A268)  and  (not A266) );
 a93446a <=( a93445a  and  a93442a );
 a93449a <=( A298  and  (not A269) );
 a93452a <=( (not A302)  and  (not A301) );
 a93453a <=( a93452a  and  a93449a );
 a93454a <=( a93453a  and  a93446a );
 a93458a <=( (not A166)  and  (not A167) );
 a93459a <=( (not A169)  and  a93458a );
 a93462a <=( (not A200)  and  A199 );
 a93465a <=( A203  and  A201 );
 a93466a <=( a93465a  and  a93462a );
 a93467a <=( a93466a  and  a93459a );
 a93470a <=( A233  and  A232 );
 a93473a <=( (not A268)  and  A265 );
 a93474a <=( a93473a  and  a93470a );
 a93477a <=( (not A299)  and  (not A269) );
 a93480a <=( (not A302)  and  (not A301) );
 a93481a <=( a93480a  and  a93477a );
 a93482a <=( a93481a  and  a93474a );
 a93486a <=( (not A166)  and  (not A167) );
 a93487a <=( (not A169)  and  a93486a );
 a93490a <=( (not A200)  and  A199 );
 a93493a <=( A203  and  A201 );
 a93494a <=( a93493a  and  a93490a );
 a93495a <=( a93494a  and  a93487a );
 a93498a <=( (not A235)  and  (not A233) );
 a93501a <=( A265  and  (not A236) );
 a93502a <=( a93501a  and  a93498a );
 a93505a <=( A298  and  A266 );
 a93508a <=( (not A302)  and  (not A301) );
 a93509a <=( a93508a  and  a93505a );
 a93510a <=( a93509a  and  a93502a );
 a93514a <=( (not A166)  and  (not A167) );
 a93515a <=( (not A169)  and  a93514a );
 a93518a <=( (not A200)  and  A199 );
 a93521a <=( A203  and  A201 );
 a93522a <=( a93521a  and  a93518a );
 a93523a <=( a93522a  and  a93515a );
 a93526a <=( (not A235)  and  (not A233) );
 a93529a <=( (not A266)  and  (not A236) );
 a93530a <=( a93529a  and  a93526a );
 a93533a <=( (not A269)  and  (not A268) );
 a93536a <=( (not A300)  and  A298 );
 a93537a <=( a93536a  and  a93533a );
 a93538a <=( a93537a  and  a93530a );
 a93542a <=( (not A166)  and  (not A167) );
 a93543a <=( (not A169)  and  a93542a );
 a93546a <=( (not A200)  and  A199 );
 a93549a <=( A203  and  A201 );
 a93550a <=( a93549a  and  a93546a );
 a93551a <=( a93550a  and  a93543a );
 a93554a <=( (not A235)  and  (not A233) );
 a93557a <=( (not A266)  and  (not A236) );
 a93558a <=( a93557a  and  a93554a );
 a93561a <=( (not A269)  and  (not A268) );
 a93564a <=( A299  and  A298 );
 a93565a <=( a93564a  and  a93561a );
 a93566a <=( a93565a  and  a93558a );
 a93570a <=( (not A166)  and  (not A167) );
 a93571a <=( (not A169)  and  a93570a );
 a93574a <=( (not A200)  and  A199 );
 a93577a <=( A203  and  A201 );
 a93578a <=( a93577a  and  a93574a );
 a93579a <=( a93578a  and  a93571a );
 a93582a <=( (not A235)  and  (not A233) );
 a93585a <=( (not A266)  and  (not A236) );
 a93586a <=( a93585a  and  a93582a );
 a93589a <=( (not A269)  and  (not A268) );
 a93592a <=( (not A299)  and  (not A298) );
 a93593a <=( a93592a  and  a93589a );
 a93594a <=( a93593a  and  a93586a );
 a93598a <=( (not A166)  and  (not A167) );
 a93599a <=( (not A169)  and  a93598a );
 a93602a <=( (not A200)  and  A199 );
 a93605a <=( A203  and  A201 );
 a93606a <=( a93605a  and  a93602a );
 a93607a <=( a93606a  and  a93599a );
 a93610a <=( (not A235)  and  (not A233) );
 a93613a <=( (not A266)  and  (not A236) );
 a93614a <=( a93613a  and  a93610a );
 a93617a <=( A298  and  (not A267) );
 a93620a <=( (not A302)  and  (not A301) );
 a93621a <=( a93620a  and  a93617a );
 a93622a <=( a93621a  and  a93614a );
 a93626a <=( (not A166)  and  (not A167) );
 a93627a <=( (not A169)  and  a93626a );
 a93630a <=( (not A200)  and  A199 );
 a93633a <=( A203  and  A201 );
 a93634a <=( a93633a  and  a93630a );
 a93635a <=( a93634a  and  a93627a );
 a93638a <=( (not A235)  and  (not A233) );
 a93641a <=( (not A265)  and  (not A236) );
 a93642a <=( a93641a  and  a93638a );
 a93645a <=( A298  and  (not A266) );
 a93648a <=( (not A302)  and  (not A301) );
 a93649a <=( a93648a  and  a93645a );
 a93650a <=( a93649a  and  a93642a );
 a93654a <=( (not A166)  and  (not A167) );
 a93655a <=( (not A169)  and  a93654a );
 a93658a <=( (not A200)  and  A199 );
 a93661a <=( A203  and  A201 );
 a93662a <=( a93661a  and  a93658a );
 a93663a <=( a93662a  and  a93655a );
 a93666a <=( (not A234)  and  (not A233) );
 a93669a <=( (not A268)  and  (not A266) );
 a93670a <=( a93669a  and  a93666a );
 a93673a <=( A298  and  (not A269) );
 a93676a <=( (not A302)  and  (not A301) );
 a93677a <=( a93676a  and  a93673a );
 a93678a <=( a93677a  and  a93670a );
 a93682a <=( (not A166)  and  (not A167) );
 a93683a <=( (not A169)  and  a93682a );
 a93686a <=( (not A200)  and  A199 );
 a93689a <=( A203  and  A201 );
 a93690a <=( a93689a  and  a93686a );
 a93691a <=( a93690a  and  a93683a );
 a93694a <=( (not A233)  and  A232 );
 a93697a <=( A235  and  A234 );
 a93698a <=( a93697a  and  a93694a );
 a93701a <=( (not A299)  and  A298 );
 a93704a <=( A301  and  A300 );
 a93705a <=( a93704a  and  a93701a );
 a93706a <=( a93705a  and  a93698a );
 a93710a <=( (not A166)  and  (not A167) );
 a93711a <=( (not A169)  and  a93710a );
 a93714a <=( (not A200)  and  A199 );
 a93717a <=( A203  and  A201 );
 a93718a <=( a93717a  and  a93714a );
 a93719a <=( a93718a  and  a93711a );
 a93722a <=( (not A233)  and  A232 );
 a93725a <=( A235  and  A234 );
 a93726a <=( a93725a  and  a93722a );
 a93729a <=( (not A299)  and  A298 );
 a93732a <=( A302  and  A300 );
 a93733a <=( a93732a  and  a93729a );
 a93734a <=( a93733a  and  a93726a );
 a93738a <=( (not A166)  and  (not A167) );
 a93739a <=( (not A169)  and  a93738a );
 a93742a <=( (not A200)  and  A199 );
 a93745a <=( A203  and  A201 );
 a93746a <=( a93745a  and  a93742a );
 a93747a <=( a93746a  and  a93739a );
 a93750a <=( (not A233)  and  A232 );
 a93753a <=( A235  and  A234 );
 a93754a <=( a93753a  and  a93750a );
 a93757a <=( (not A266)  and  A265 );
 a93760a <=( A268  and  A267 );
 a93761a <=( a93760a  and  a93757a );
 a93762a <=( a93761a  and  a93754a );
 a93766a <=( (not A166)  and  (not A167) );
 a93767a <=( (not A169)  and  a93766a );
 a93770a <=( (not A200)  and  A199 );
 a93773a <=( A203  and  A201 );
 a93774a <=( a93773a  and  a93770a );
 a93775a <=( a93774a  and  a93767a );
 a93778a <=( (not A233)  and  A232 );
 a93781a <=( A235  and  A234 );
 a93782a <=( a93781a  and  a93778a );
 a93785a <=( (not A266)  and  A265 );
 a93788a <=( A269  and  A267 );
 a93789a <=( a93788a  and  a93785a );
 a93790a <=( a93789a  and  a93782a );
 a93794a <=( (not A166)  and  (not A167) );
 a93795a <=( (not A169)  and  a93794a );
 a93798a <=( (not A200)  and  A199 );
 a93801a <=( A203  and  A201 );
 a93802a <=( a93801a  and  a93798a );
 a93803a <=( a93802a  and  a93795a );
 a93806a <=( (not A233)  and  A232 );
 a93809a <=( A236  and  A234 );
 a93810a <=( a93809a  and  a93806a );
 a93813a <=( (not A299)  and  A298 );
 a93816a <=( A301  and  A300 );
 a93817a <=( a93816a  and  a93813a );
 a93818a <=( a93817a  and  a93810a );
 a93822a <=( (not A166)  and  (not A167) );
 a93823a <=( (not A169)  and  a93822a );
 a93826a <=( (not A200)  and  A199 );
 a93829a <=( A203  and  A201 );
 a93830a <=( a93829a  and  a93826a );
 a93831a <=( a93830a  and  a93823a );
 a93834a <=( (not A233)  and  A232 );
 a93837a <=( A236  and  A234 );
 a93838a <=( a93837a  and  a93834a );
 a93841a <=( (not A299)  and  A298 );
 a93844a <=( A302  and  A300 );
 a93845a <=( a93844a  and  a93841a );
 a93846a <=( a93845a  and  a93838a );
 a93850a <=( (not A166)  and  (not A167) );
 a93851a <=( (not A169)  and  a93850a );
 a93854a <=( (not A200)  and  A199 );
 a93857a <=( A203  and  A201 );
 a93858a <=( a93857a  and  a93854a );
 a93859a <=( a93858a  and  a93851a );
 a93862a <=( (not A233)  and  A232 );
 a93865a <=( A236  and  A234 );
 a93866a <=( a93865a  and  a93862a );
 a93869a <=( (not A266)  and  A265 );
 a93872a <=( A268  and  A267 );
 a93873a <=( a93872a  and  a93869a );
 a93874a <=( a93873a  and  a93866a );
 a93878a <=( (not A166)  and  (not A167) );
 a93879a <=( (not A169)  and  a93878a );
 a93882a <=( (not A200)  and  A199 );
 a93885a <=( A203  and  A201 );
 a93886a <=( a93885a  and  a93882a );
 a93887a <=( a93886a  and  a93879a );
 a93890a <=( (not A233)  and  A232 );
 a93893a <=( A236  and  A234 );
 a93894a <=( a93893a  and  a93890a );
 a93897a <=( (not A266)  and  A265 );
 a93900a <=( A269  and  A267 );
 a93901a <=( a93900a  and  a93897a );
 a93902a <=( a93901a  and  a93894a );
 a93906a <=( (not A166)  and  (not A167) );
 a93907a <=( (not A169)  and  a93906a );
 a93910a <=( (not A200)  and  A199 );
 a93913a <=( A203  and  A201 );
 a93914a <=( a93913a  and  a93910a );
 a93915a <=( a93914a  and  a93907a );
 a93918a <=( (not A233)  and  (not A232) );
 a93921a <=( (not A268)  and  (not A266) );
 a93922a <=( a93921a  and  a93918a );
 a93925a <=( A298  and  (not A269) );
 a93928a <=( (not A302)  and  (not A301) );
 a93929a <=( a93928a  and  a93925a );
 a93930a <=( a93929a  and  a93922a );
 a93934a <=( A167  and  (not A168) );
 a93935a <=( (not A169)  and  a93934a );
 a93938a <=( (not A199)  and  A166 );
 a93941a <=( (not A233)  and  A200 );
 a93942a <=( a93941a  and  a93938a );
 a93943a <=( a93942a  and  a93935a );
 a93946a <=( (not A236)  and  (not A235) );
 a93949a <=( (not A268)  and  (not A266) );
 a93950a <=( a93949a  and  a93946a );
 a93953a <=( A298  and  (not A269) );
 a93956a <=( (not A302)  and  (not A301) );
 a93957a <=( a93956a  and  a93953a );
 a93958a <=( a93957a  and  a93950a );
 a93962a <=( A167  and  (not A168) );
 a93963a <=( (not A169)  and  a93962a );
 a93966a <=( A199  and  A166 );
 a93969a <=( A201  and  (not A200) );
 a93970a <=( a93969a  and  a93966a );
 a93971a <=( a93970a  and  a93963a );
 a93974a <=( A232  and  A202 );
 a93977a <=( A265  and  A233 );
 a93978a <=( a93977a  and  a93974a );
 a93981a <=( (not A269)  and  (not A268) );
 a93984a <=( (not A300)  and  (not A299) );
 a93985a <=( a93984a  and  a93981a );
 a93986a <=( a93985a  and  a93978a );
 a93990a <=( A167  and  (not A168) );
 a93991a <=( (not A169)  and  a93990a );
 a93994a <=( A199  and  A166 );
 a93997a <=( A201  and  (not A200) );
 a93998a <=( a93997a  and  a93994a );
 a93999a <=( a93998a  and  a93991a );
 a94002a <=( A232  and  A202 );
 a94005a <=( A265  and  A233 );
 a94006a <=( a94005a  and  a94002a );
 a94009a <=( (not A269)  and  (not A268) );
 a94012a <=( A299  and  A298 );
 a94013a <=( a94012a  and  a94009a );
 a94014a <=( a94013a  and  a94006a );
 a94018a <=( A167  and  (not A168) );
 a94019a <=( (not A169)  and  a94018a );
 a94022a <=( A199  and  A166 );
 a94025a <=( A201  and  (not A200) );
 a94026a <=( a94025a  and  a94022a );
 a94027a <=( a94026a  and  a94019a );
 a94030a <=( A232  and  A202 );
 a94033a <=( A265  and  A233 );
 a94034a <=( a94033a  and  a94030a );
 a94037a <=( (not A269)  and  (not A268) );
 a94040a <=( (not A299)  and  (not A298) );
 a94041a <=( a94040a  and  a94037a );
 a94042a <=( a94041a  and  a94034a );
 a94046a <=( A167  and  (not A168) );
 a94047a <=( (not A169)  and  a94046a );
 a94050a <=( A199  and  A166 );
 a94053a <=( A201  and  (not A200) );
 a94054a <=( a94053a  and  a94050a );
 a94055a <=( a94054a  and  a94047a );
 a94058a <=( A232  and  A202 );
 a94061a <=( A265  and  A233 );
 a94062a <=( a94061a  and  a94058a );
 a94065a <=( (not A299)  and  (not A267) );
 a94068a <=( (not A302)  and  (not A301) );
 a94069a <=( a94068a  and  a94065a );
 a94070a <=( a94069a  and  a94062a );
 a94074a <=( A167  and  (not A168) );
 a94075a <=( (not A169)  and  a94074a );
 a94078a <=( A199  and  A166 );
 a94081a <=( A201  and  (not A200) );
 a94082a <=( a94081a  and  a94078a );
 a94083a <=( a94082a  and  a94075a );
 a94086a <=( A232  and  A202 );
 a94089a <=( A265  and  A233 );
 a94090a <=( a94089a  and  a94086a );
 a94093a <=( (not A299)  and  A266 );
 a94096a <=( (not A302)  and  (not A301) );
 a94097a <=( a94096a  and  a94093a );
 a94098a <=( a94097a  and  a94090a );
 a94102a <=( A167  and  (not A168) );
 a94103a <=( (not A169)  and  a94102a );
 a94106a <=( A199  and  A166 );
 a94109a <=( A201  and  (not A200) );
 a94110a <=( a94109a  and  a94106a );
 a94111a <=( a94110a  and  a94103a );
 a94114a <=( A232  and  A202 );
 a94117a <=( (not A265)  and  A233 );
 a94118a <=( a94117a  and  a94114a );
 a94121a <=( (not A299)  and  (not A266) );
 a94124a <=( (not A302)  and  (not A301) );
 a94125a <=( a94124a  and  a94121a );
 a94126a <=( a94125a  and  a94118a );
 a94130a <=( A167  and  (not A168) );
 a94131a <=( (not A169)  and  a94130a );
 a94134a <=( A199  and  A166 );
 a94137a <=( A201  and  (not A200) );
 a94138a <=( a94137a  and  a94134a );
 a94139a <=( a94138a  and  a94131a );
 a94142a <=( (not A233)  and  A202 );
 a94145a <=( (not A236)  and  (not A235) );
 a94146a <=( a94145a  and  a94142a );
 a94149a <=( A266  and  A265 );
 a94152a <=( (not A300)  and  A298 );
 a94153a <=( a94152a  and  a94149a );
 a94154a <=( a94153a  and  a94146a );
 a94158a <=( A167  and  (not A168) );
 a94159a <=( (not A169)  and  a94158a );
 a94162a <=( A199  and  A166 );
 a94165a <=( A201  and  (not A200) );
 a94166a <=( a94165a  and  a94162a );
 a94167a <=( a94166a  and  a94159a );
 a94170a <=( (not A233)  and  A202 );
 a94173a <=( (not A236)  and  (not A235) );
 a94174a <=( a94173a  and  a94170a );
 a94177a <=( A266  and  A265 );
 a94180a <=( A299  and  A298 );
 a94181a <=( a94180a  and  a94177a );
 a94182a <=( a94181a  and  a94174a );
 a94186a <=( A167  and  (not A168) );
 a94187a <=( (not A169)  and  a94186a );
 a94190a <=( A199  and  A166 );
 a94193a <=( A201  and  (not A200) );
 a94194a <=( a94193a  and  a94190a );
 a94195a <=( a94194a  and  a94187a );
 a94198a <=( (not A233)  and  A202 );
 a94201a <=( (not A236)  and  (not A235) );
 a94202a <=( a94201a  and  a94198a );
 a94205a <=( A266  and  A265 );
 a94208a <=( (not A299)  and  (not A298) );
 a94209a <=( a94208a  and  a94205a );
 a94210a <=( a94209a  and  a94202a );
 a94214a <=( A167  and  (not A168) );
 a94215a <=( (not A169)  and  a94214a );
 a94218a <=( A199  and  A166 );
 a94221a <=( A201  and  (not A200) );
 a94222a <=( a94221a  and  a94218a );
 a94223a <=( a94222a  and  a94215a );
 a94226a <=( (not A233)  and  A202 );
 a94229a <=( (not A236)  and  (not A235) );
 a94230a <=( a94229a  and  a94226a );
 a94233a <=( (not A267)  and  (not A266) );
 a94236a <=( (not A300)  and  A298 );
 a94237a <=( a94236a  and  a94233a );
 a94238a <=( a94237a  and  a94230a );
 a94242a <=( A167  and  (not A168) );
 a94243a <=( (not A169)  and  a94242a );
 a94246a <=( A199  and  A166 );
 a94249a <=( A201  and  (not A200) );
 a94250a <=( a94249a  and  a94246a );
 a94251a <=( a94250a  and  a94243a );
 a94254a <=( (not A233)  and  A202 );
 a94257a <=( (not A236)  and  (not A235) );
 a94258a <=( a94257a  and  a94254a );
 a94261a <=( (not A267)  and  (not A266) );
 a94264a <=( A299  and  A298 );
 a94265a <=( a94264a  and  a94261a );
 a94266a <=( a94265a  and  a94258a );
 a94270a <=( A167  and  (not A168) );
 a94271a <=( (not A169)  and  a94270a );
 a94274a <=( A199  and  A166 );
 a94277a <=( A201  and  (not A200) );
 a94278a <=( a94277a  and  a94274a );
 a94279a <=( a94278a  and  a94271a );
 a94282a <=( (not A233)  and  A202 );
 a94285a <=( (not A236)  and  (not A235) );
 a94286a <=( a94285a  and  a94282a );
 a94289a <=( (not A267)  and  (not A266) );
 a94292a <=( (not A299)  and  (not A298) );
 a94293a <=( a94292a  and  a94289a );
 a94294a <=( a94293a  and  a94286a );
 a94298a <=( A167  and  (not A168) );
 a94299a <=( (not A169)  and  a94298a );
 a94302a <=( A199  and  A166 );
 a94305a <=( A201  and  (not A200) );
 a94306a <=( a94305a  and  a94302a );
 a94307a <=( a94306a  and  a94299a );
 a94310a <=( (not A233)  and  A202 );
 a94313a <=( (not A236)  and  (not A235) );
 a94314a <=( a94313a  and  a94310a );
 a94317a <=( (not A266)  and  (not A265) );
 a94320a <=( (not A300)  and  A298 );
 a94321a <=( a94320a  and  a94317a );
 a94322a <=( a94321a  and  a94314a );
 a94326a <=( A167  and  (not A168) );
 a94327a <=( (not A169)  and  a94326a );
 a94330a <=( A199  and  A166 );
 a94333a <=( A201  and  (not A200) );
 a94334a <=( a94333a  and  a94330a );
 a94335a <=( a94334a  and  a94327a );
 a94338a <=( (not A233)  and  A202 );
 a94341a <=( (not A236)  and  (not A235) );
 a94342a <=( a94341a  and  a94338a );
 a94345a <=( (not A266)  and  (not A265) );
 a94348a <=( A299  and  A298 );
 a94349a <=( a94348a  and  a94345a );
 a94350a <=( a94349a  and  a94342a );
 a94354a <=( A167  and  (not A168) );
 a94355a <=( (not A169)  and  a94354a );
 a94358a <=( A199  and  A166 );
 a94361a <=( A201  and  (not A200) );
 a94362a <=( a94361a  and  a94358a );
 a94363a <=( a94362a  and  a94355a );
 a94366a <=( (not A233)  and  A202 );
 a94369a <=( (not A236)  and  (not A235) );
 a94370a <=( a94369a  and  a94366a );
 a94373a <=( (not A266)  and  (not A265) );
 a94376a <=( (not A299)  and  (not A298) );
 a94377a <=( a94376a  and  a94373a );
 a94378a <=( a94377a  and  a94370a );
 a94382a <=( A167  and  (not A168) );
 a94383a <=( (not A169)  and  a94382a );
 a94386a <=( A199  and  A166 );
 a94389a <=( A201  and  (not A200) );
 a94390a <=( a94389a  and  a94386a );
 a94391a <=( a94390a  and  a94383a );
 a94394a <=( (not A233)  and  A202 );
 a94397a <=( A265  and  (not A234) );
 a94398a <=( a94397a  and  a94394a );
 a94401a <=( A298  and  A266 );
 a94404a <=( (not A302)  and  (not A301) );
 a94405a <=( a94404a  and  a94401a );
 a94406a <=( a94405a  and  a94398a );
 a94410a <=( A167  and  (not A168) );
 a94411a <=( (not A169)  and  a94410a );
 a94414a <=( A199  and  A166 );
 a94417a <=( A201  and  (not A200) );
 a94418a <=( a94417a  and  a94414a );
 a94419a <=( a94418a  and  a94411a );
 a94422a <=( (not A233)  and  A202 );
 a94425a <=( (not A266)  and  (not A234) );
 a94426a <=( a94425a  and  a94422a );
 a94429a <=( (not A269)  and  (not A268) );
 a94432a <=( (not A300)  and  A298 );
 a94433a <=( a94432a  and  a94429a );
 a94434a <=( a94433a  and  a94426a );
 a94438a <=( A167  and  (not A168) );
 a94439a <=( (not A169)  and  a94438a );
 a94442a <=( A199  and  A166 );
 a94445a <=( A201  and  (not A200) );
 a94446a <=( a94445a  and  a94442a );
 a94447a <=( a94446a  and  a94439a );
 a94450a <=( (not A233)  and  A202 );
 a94453a <=( (not A266)  and  (not A234) );
 a94454a <=( a94453a  and  a94450a );
 a94457a <=( (not A269)  and  (not A268) );
 a94460a <=( A299  and  A298 );
 a94461a <=( a94460a  and  a94457a );
 a94462a <=( a94461a  and  a94454a );
 a94466a <=( A167  and  (not A168) );
 a94467a <=( (not A169)  and  a94466a );
 a94470a <=( A199  and  A166 );
 a94473a <=( A201  and  (not A200) );
 a94474a <=( a94473a  and  a94470a );
 a94475a <=( a94474a  and  a94467a );
 a94478a <=( (not A233)  and  A202 );
 a94481a <=( (not A266)  and  (not A234) );
 a94482a <=( a94481a  and  a94478a );
 a94485a <=( (not A269)  and  (not A268) );
 a94488a <=( (not A299)  and  (not A298) );
 a94489a <=( a94488a  and  a94485a );
 a94490a <=( a94489a  and  a94482a );
 a94494a <=( A167  and  (not A168) );
 a94495a <=( (not A169)  and  a94494a );
 a94498a <=( A199  and  A166 );
 a94501a <=( A201  and  (not A200) );
 a94502a <=( a94501a  and  a94498a );
 a94503a <=( a94502a  and  a94495a );
 a94506a <=( (not A233)  and  A202 );
 a94509a <=( (not A266)  and  (not A234) );
 a94510a <=( a94509a  and  a94506a );
 a94513a <=( A298  and  (not A267) );
 a94516a <=( (not A302)  and  (not A301) );
 a94517a <=( a94516a  and  a94513a );
 a94518a <=( a94517a  and  a94510a );
 a94522a <=( A167  and  (not A168) );
 a94523a <=( (not A169)  and  a94522a );
 a94526a <=( A199  and  A166 );
 a94529a <=( A201  and  (not A200) );
 a94530a <=( a94529a  and  a94526a );
 a94531a <=( a94530a  and  a94523a );
 a94534a <=( (not A233)  and  A202 );
 a94537a <=( (not A265)  and  (not A234) );
 a94538a <=( a94537a  and  a94534a );
 a94541a <=( A298  and  (not A266) );
 a94544a <=( (not A302)  and  (not A301) );
 a94545a <=( a94544a  and  a94541a );
 a94546a <=( a94545a  and  a94538a );
 a94550a <=( A167  and  (not A168) );
 a94551a <=( (not A169)  and  a94550a );
 a94554a <=( A199  and  A166 );
 a94557a <=( A201  and  (not A200) );
 a94558a <=( a94557a  and  a94554a );
 a94559a <=( a94558a  and  a94551a );
 a94562a <=( (not A232)  and  A202 );
 a94565a <=( A265  and  (not A233) );
 a94566a <=( a94565a  and  a94562a );
 a94569a <=( A298  and  A266 );
 a94572a <=( (not A302)  and  (not A301) );
 a94573a <=( a94572a  and  a94569a );
 a94574a <=( a94573a  and  a94566a );
 a94578a <=( A167  and  (not A168) );
 a94579a <=( (not A169)  and  a94578a );
 a94582a <=( A199  and  A166 );
 a94585a <=( A201  and  (not A200) );
 a94586a <=( a94585a  and  a94582a );
 a94587a <=( a94586a  and  a94579a );
 a94590a <=( (not A232)  and  A202 );
 a94593a <=( (not A266)  and  (not A233) );
 a94594a <=( a94593a  and  a94590a );
 a94597a <=( (not A269)  and  (not A268) );
 a94600a <=( (not A300)  and  A298 );
 a94601a <=( a94600a  and  a94597a );
 a94602a <=( a94601a  and  a94594a );
 a94606a <=( A167  and  (not A168) );
 a94607a <=( (not A169)  and  a94606a );
 a94610a <=( A199  and  A166 );
 a94613a <=( A201  and  (not A200) );
 a94614a <=( a94613a  and  a94610a );
 a94615a <=( a94614a  and  a94607a );
 a94618a <=( (not A232)  and  A202 );
 a94621a <=( (not A266)  and  (not A233) );
 a94622a <=( a94621a  and  a94618a );
 a94625a <=( (not A269)  and  (not A268) );
 a94628a <=( A299  and  A298 );
 a94629a <=( a94628a  and  a94625a );
 a94630a <=( a94629a  and  a94622a );
 a94634a <=( A167  and  (not A168) );
 a94635a <=( (not A169)  and  a94634a );
 a94638a <=( A199  and  A166 );
 a94641a <=( A201  and  (not A200) );
 a94642a <=( a94641a  and  a94638a );
 a94643a <=( a94642a  and  a94635a );
 a94646a <=( (not A232)  and  A202 );
 a94649a <=( (not A266)  and  (not A233) );
 a94650a <=( a94649a  and  a94646a );
 a94653a <=( (not A269)  and  (not A268) );
 a94656a <=( (not A299)  and  (not A298) );
 a94657a <=( a94656a  and  a94653a );
 a94658a <=( a94657a  and  a94650a );
 a94662a <=( A167  and  (not A168) );
 a94663a <=( (not A169)  and  a94662a );
 a94666a <=( A199  and  A166 );
 a94669a <=( A201  and  (not A200) );
 a94670a <=( a94669a  and  a94666a );
 a94671a <=( a94670a  and  a94663a );
 a94674a <=( (not A232)  and  A202 );
 a94677a <=( (not A266)  and  (not A233) );
 a94678a <=( a94677a  and  a94674a );
 a94681a <=( A298  and  (not A267) );
 a94684a <=( (not A302)  and  (not A301) );
 a94685a <=( a94684a  and  a94681a );
 a94686a <=( a94685a  and  a94678a );
 a94690a <=( A167  and  (not A168) );
 a94691a <=( (not A169)  and  a94690a );
 a94694a <=( A199  and  A166 );
 a94697a <=( A201  and  (not A200) );
 a94698a <=( a94697a  and  a94694a );
 a94699a <=( a94698a  and  a94691a );
 a94702a <=( (not A232)  and  A202 );
 a94705a <=( (not A265)  and  (not A233) );
 a94706a <=( a94705a  and  a94702a );
 a94709a <=( A298  and  (not A266) );
 a94712a <=( (not A302)  and  (not A301) );
 a94713a <=( a94712a  and  a94709a );
 a94714a <=( a94713a  and  a94706a );
 a94718a <=( A167  and  (not A168) );
 a94719a <=( (not A169)  and  a94718a );
 a94722a <=( A199  and  A166 );
 a94725a <=( A201  and  (not A200) );
 a94726a <=( a94725a  and  a94722a );
 a94727a <=( a94726a  and  a94719a );
 a94730a <=( A232  and  A203 );
 a94733a <=( A265  and  A233 );
 a94734a <=( a94733a  and  a94730a );
 a94737a <=( (not A269)  and  (not A268) );
 a94740a <=( (not A300)  and  (not A299) );
 a94741a <=( a94740a  and  a94737a );
 a94742a <=( a94741a  and  a94734a );
 a94746a <=( A167  and  (not A168) );
 a94747a <=( (not A169)  and  a94746a );
 a94750a <=( A199  and  A166 );
 a94753a <=( A201  and  (not A200) );
 a94754a <=( a94753a  and  a94750a );
 a94755a <=( a94754a  and  a94747a );
 a94758a <=( A232  and  A203 );
 a94761a <=( A265  and  A233 );
 a94762a <=( a94761a  and  a94758a );
 a94765a <=( (not A269)  and  (not A268) );
 a94768a <=( A299  and  A298 );
 a94769a <=( a94768a  and  a94765a );
 a94770a <=( a94769a  and  a94762a );
 a94774a <=( A167  and  (not A168) );
 a94775a <=( (not A169)  and  a94774a );
 a94778a <=( A199  and  A166 );
 a94781a <=( A201  and  (not A200) );
 a94782a <=( a94781a  and  a94778a );
 a94783a <=( a94782a  and  a94775a );
 a94786a <=( A232  and  A203 );
 a94789a <=( A265  and  A233 );
 a94790a <=( a94789a  and  a94786a );
 a94793a <=( (not A269)  and  (not A268) );
 a94796a <=( (not A299)  and  (not A298) );
 a94797a <=( a94796a  and  a94793a );
 a94798a <=( a94797a  and  a94790a );
 a94802a <=( A167  and  (not A168) );
 a94803a <=( (not A169)  and  a94802a );
 a94806a <=( A199  and  A166 );
 a94809a <=( A201  and  (not A200) );
 a94810a <=( a94809a  and  a94806a );
 a94811a <=( a94810a  and  a94803a );
 a94814a <=( A232  and  A203 );
 a94817a <=( A265  and  A233 );
 a94818a <=( a94817a  and  a94814a );
 a94821a <=( (not A299)  and  (not A267) );
 a94824a <=( (not A302)  and  (not A301) );
 a94825a <=( a94824a  and  a94821a );
 a94826a <=( a94825a  and  a94818a );
 a94830a <=( A167  and  (not A168) );
 a94831a <=( (not A169)  and  a94830a );
 a94834a <=( A199  and  A166 );
 a94837a <=( A201  and  (not A200) );
 a94838a <=( a94837a  and  a94834a );
 a94839a <=( a94838a  and  a94831a );
 a94842a <=( A232  and  A203 );
 a94845a <=( A265  and  A233 );
 a94846a <=( a94845a  and  a94842a );
 a94849a <=( (not A299)  and  A266 );
 a94852a <=( (not A302)  and  (not A301) );
 a94853a <=( a94852a  and  a94849a );
 a94854a <=( a94853a  and  a94846a );
 a94858a <=( A167  and  (not A168) );
 a94859a <=( (not A169)  and  a94858a );
 a94862a <=( A199  and  A166 );
 a94865a <=( A201  and  (not A200) );
 a94866a <=( a94865a  and  a94862a );
 a94867a <=( a94866a  and  a94859a );
 a94870a <=( A232  and  A203 );
 a94873a <=( (not A265)  and  A233 );
 a94874a <=( a94873a  and  a94870a );
 a94877a <=( (not A299)  and  (not A266) );
 a94880a <=( (not A302)  and  (not A301) );
 a94881a <=( a94880a  and  a94877a );
 a94882a <=( a94881a  and  a94874a );
 a94886a <=( A167  and  (not A168) );
 a94887a <=( (not A169)  and  a94886a );
 a94890a <=( A199  and  A166 );
 a94893a <=( A201  and  (not A200) );
 a94894a <=( a94893a  and  a94890a );
 a94895a <=( a94894a  and  a94887a );
 a94898a <=( (not A233)  and  A203 );
 a94901a <=( (not A236)  and  (not A235) );
 a94902a <=( a94901a  and  a94898a );
 a94905a <=( A266  and  A265 );
 a94908a <=( (not A300)  and  A298 );
 a94909a <=( a94908a  and  a94905a );
 a94910a <=( a94909a  and  a94902a );
 a94914a <=( A167  and  (not A168) );
 a94915a <=( (not A169)  and  a94914a );
 a94918a <=( A199  and  A166 );
 a94921a <=( A201  and  (not A200) );
 a94922a <=( a94921a  and  a94918a );
 a94923a <=( a94922a  and  a94915a );
 a94926a <=( (not A233)  and  A203 );
 a94929a <=( (not A236)  and  (not A235) );
 a94930a <=( a94929a  and  a94926a );
 a94933a <=( A266  and  A265 );
 a94936a <=( A299  and  A298 );
 a94937a <=( a94936a  and  a94933a );
 a94938a <=( a94937a  and  a94930a );
 a94942a <=( A167  and  (not A168) );
 a94943a <=( (not A169)  and  a94942a );
 a94946a <=( A199  and  A166 );
 a94949a <=( A201  and  (not A200) );
 a94950a <=( a94949a  and  a94946a );
 a94951a <=( a94950a  and  a94943a );
 a94954a <=( (not A233)  and  A203 );
 a94957a <=( (not A236)  and  (not A235) );
 a94958a <=( a94957a  and  a94954a );
 a94961a <=( A266  and  A265 );
 a94964a <=( (not A299)  and  (not A298) );
 a94965a <=( a94964a  and  a94961a );
 a94966a <=( a94965a  and  a94958a );
 a94970a <=( A167  and  (not A168) );
 a94971a <=( (not A169)  and  a94970a );
 a94974a <=( A199  and  A166 );
 a94977a <=( A201  and  (not A200) );
 a94978a <=( a94977a  and  a94974a );
 a94979a <=( a94978a  and  a94971a );
 a94982a <=( (not A233)  and  A203 );
 a94985a <=( (not A236)  and  (not A235) );
 a94986a <=( a94985a  and  a94982a );
 a94989a <=( (not A267)  and  (not A266) );
 a94992a <=( (not A300)  and  A298 );
 a94993a <=( a94992a  and  a94989a );
 a94994a <=( a94993a  and  a94986a );
 a94998a <=( A167  and  (not A168) );
 a94999a <=( (not A169)  and  a94998a );
 a95002a <=( A199  and  A166 );
 a95005a <=( A201  and  (not A200) );
 a95006a <=( a95005a  and  a95002a );
 a95007a <=( a95006a  and  a94999a );
 a95010a <=( (not A233)  and  A203 );
 a95013a <=( (not A236)  and  (not A235) );
 a95014a <=( a95013a  and  a95010a );
 a95017a <=( (not A267)  and  (not A266) );
 a95020a <=( A299  and  A298 );
 a95021a <=( a95020a  and  a95017a );
 a95022a <=( a95021a  and  a95014a );
 a95026a <=( A167  and  (not A168) );
 a95027a <=( (not A169)  and  a95026a );
 a95030a <=( A199  and  A166 );
 a95033a <=( A201  and  (not A200) );
 a95034a <=( a95033a  and  a95030a );
 a95035a <=( a95034a  and  a95027a );
 a95038a <=( (not A233)  and  A203 );
 a95041a <=( (not A236)  and  (not A235) );
 a95042a <=( a95041a  and  a95038a );
 a95045a <=( (not A267)  and  (not A266) );
 a95048a <=( (not A299)  and  (not A298) );
 a95049a <=( a95048a  and  a95045a );
 a95050a <=( a95049a  and  a95042a );
 a95054a <=( A167  and  (not A168) );
 a95055a <=( (not A169)  and  a95054a );
 a95058a <=( A199  and  A166 );
 a95061a <=( A201  and  (not A200) );
 a95062a <=( a95061a  and  a95058a );
 a95063a <=( a95062a  and  a95055a );
 a95066a <=( (not A233)  and  A203 );
 a95069a <=( (not A236)  and  (not A235) );
 a95070a <=( a95069a  and  a95066a );
 a95073a <=( (not A266)  and  (not A265) );
 a95076a <=( (not A300)  and  A298 );
 a95077a <=( a95076a  and  a95073a );
 a95078a <=( a95077a  and  a95070a );
 a95082a <=( A167  and  (not A168) );
 a95083a <=( (not A169)  and  a95082a );
 a95086a <=( A199  and  A166 );
 a95089a <=( A201  and  (not A200) );
 a95090a <=( a95089a  and  a95086a );
 a95091a <=( a95090a  and  a95083a );
 a95094a <=( (not A233)  and  A203 );
 a95097a <=( (not A236)  and  (not A235) );
 a95098a <=( a95097a  and  a95094a );
 a95101a <=( (not A266)  and  (not A265) );
 a95104a <=( A299  and  A298 );
 a95105a <=( a95104a  and  a95101a );
 a95106a <=( a95105a  and  a95098a );
 a95110a <=( A167  and  (not A168) );
 a95111a <=( (not A169)  and  a95110a );
 a95114a <=( A199  and  A166 );
 a95117a <=( A201  and  (not A200) );
 a95118a <=( a95117a  and  a95114a );
 a95119a <=( a95118a  and  a95111a );
 a95122a <=( (not A233)  and  A203 );
 a95125a <=( (not A236)  and  (not A235) );
 a95126a <=( a95125a  and  a95122a );
 a95129a <=( (not A266)  and  (not A265) );
 a95132a <=( (not A299)  and  (not A298) );
 a95133a <=( a95132a  and  a95129a );
 a95134a <=( a95133a  and  a95126a );
 a95138a <=( A167  and  (not A168) );
 a95139a <=( (not A169)  and  a95138a );
 a95142a <=( A199  and  A166 );
 a95145a <=( A201  and  (not A200) );
 a95146a <=( a95145a  and  a95142a );
 a95147a <=( a95146a  and  a95139a );
 a95150a <=( (not A233)  and  A203 );
 a95153a <=( A265  and  (not A234) );
 a95154a <=( a95153a  and  a95150a );
 a95157a <=( A298  and  A266 );
 a95160a <=( (not A302)  and  (not A301) );
 a95161a <=( a95160a  and  a95157a );
 a95162a <=( a95161a  and  a95154a );
 a95166a <=( A167  and  (not A168) );
 a95167a <=( (not A169)  and  a95166a );
 a95170a <=( A199  and  A166 );
 a95173a <=( A201  and  (not A200) );
 a95174a <=( a95173a  and  a95170a );
 a95175a <=( a95174a  and  a95167a );
 a95178a <=( (not A233)  and  A203 );
 a95181a <=( (not A266)  and  (not A234) );
 a95182a <=( a95181a  and  a95178a );
 a95185a <=( (not A269)  and  (not A268) );
 a95188a <=( (not A300)  and  A298 );
 a95189a <=( a95188a  and  a95185a );
 a95190a <=( a95189a  and  a95182a );
 a95194a <=( A167  and  (not A168) );
 a95195a <=( (not A169)  and  a95194a );
 a95198a <=( A199  and  A166 );
 a95201a <=( A201  and  (not A200) );
 a95202a <=( a95201a  and  a95198a );
 a95203a <=( a95202a  and  a95195a );
 a95206a <=( (not A233)  and  A203 );
 a95209a <=( (not A266)  and  (not A234) );
 a95210a <=( a95209a  and  a95206a );
 a95213a <=( (not A269)  and  (not A268) );
 a95216a <=( A299  and  A298 );
 a95217a <=( a95216a  and  a95213a );
 a95218a <=( a95217a  and  a95210a );
 a95222a <=( A167  and  (not A168) );
 a95223a <=( (not A169)  and  a95222a );
 a95226a <=( A199  and  A166 );
 a95229a <=( A201  and  (not A200) );
 a95230a <=( a95229a  and  a95226a );
 a95231a <=( a95230a  and  a95223a );
 a95234a <=( (not A233)  and  A203 );
 a95237a <=( (not A266)  and  (not A234) );
 a95238a <=( a95237a  and  a95234a );
 a95241a <=( (not A269)  and  (not A268) );
 a95244a <=( (not A299)  and  (not A298) );
 a95245a <=( a95244a  and  a95241a );
 a95246a <=( a95245a  and  a95238a );
 a95250a <=( A167  and  (not A168) );
 a95251a <=( (not A169)  and  a95250a );
 a95254a <=( A199  and  A166 );
 a95257a <=( A201  and  (not A200) );
 a95258a <=( a95257a  and  a95254a );
 a95259a <=( a95258a  and  a95251a );
 a95262a <=( (not A233)  and  A203 );
 a95265a <=( (not A266)  and  (not A234) );
 a95266a <=( a95265a  and  a95262a );
 a95269a <=( A298  and  (not A267) );
 a95272a <=( (not A302)  and  (not A301) );
 a95273a <=( a95272a  and  a95269a );
 a95274a <=( a95273a  and  a95266a );
 a95278a <=( A167  and  (not A168) );
 a95279a <=( (not A169)  and  a95278a );
 a95282a <=( A199  and  A166 );
 a95285a <=( A201  and  (not A200) );
 a95286a <=( a95285a  and  a95282a );
 a95287a <=( a95286a  and  a95279a );
 a95290a <=( (not A233)  and  A203 );
 a95293a <=( (not A265)  and  (not A234) );
 a95294a <=( a95293a  and  a95290a );
 a95297a <=( A298  and  (not A266) );
 a95300a <=( (not A302)  and  (not A301) );
 a95301a <=( a95300a  and  a95297a );
 a95302a <=( a95301a  and  a95294a );
 a95306a <=( A167  and  (not A168) );
 a95307a <=( (not A169)  and  a95306a );
 a95310a <=( A199  and  A166 );
 a95313a <=( A201  and  (not A200) );
 a95314a <=( a95313a  and  a95310a );
 a95315a <=( a95314a  and  a95307a );
 a95318a <=( (not A232)  and  A203 );
 a95321a <=( A265  and  (not A233) );
 a95322a <=( a95321a  and  a95318a );
 a95325a <=( A298  and  A266 );
 a95328a <=( (not A302)  and  (not A301) );
 a95329a <=( a95328a  and  a95325a );
 a95330a <=( a95329a  and  a95322a );
 a95334a <=( A167  and  (not A168) );
 a95335a <=( (not A169)  and  a95334a );
 a95338a <=( A199  and  A166 );
 a95341a <=( A201  and  (not A200) );
 a95342a <=( a95341a  and  a95338a );
 a95343a <=( a95342a  and  a95335a );
 a95346a <=( (not A232)  and  A203 );
 a95349a <=( (not A266)  and  (not A233) );
 a95350a <=( a95349a  and  a95346a );
 a95353a <=( (not A269)  and  (not A268) );
 a95356a <=( (not A300)  and  A298 );
 a95357a <=( a95356a  and  a95353a );
 a95358a <=( a95357a  and  a95350a );
 a95362a <=( A167  and  (not A168) );
 a95363a <=( (not A169)  and  a95362a );
 a95366a <=( A199  and  A166 );
 a95369a <=( A201  and  (not A200) );
 a95370a <=( a95369a  and  a95366a );
 a95371a <=( a95370a  and  a95363a );
 a95374a <=( (not A232)  and  A203 );
 a95377a <=( (not A266)  and  (not A233) );
 a95378a <=( a95377a  and  a95374a );
 a95381a <=( (not A269)  and  (not A268) );
 a95384a <=( A299  and  A298 );
 a95385a <=( a95384a  and  a95381a );
 a95386a <=( a95385a  and  a95378a );
 a95390a <=( A167  and  (not A168) );
 a95391a <=( (not A169)  and  a95390a );
 a95394a <=( A199  and  A166 );
 a95397a <=( A201  and  (not A200) );
 a95398a <=( a95397a  and  a95394a );
 a95399a <=( a95398a  and  a95391a );
 a95402a <=( (not A232)  and  A203 );
 a95405a <=( (not A266)  and  (not A233) );
 a95406a <=( a95405a  and  a95402a );
 a95409a <=( (not A269)  and  (not A268) );
 a95412a <=( (not A299)  and  (not A298) );
 a95413a <=( a95412a  and  a95409a );
 a95414a <=( a95413a  and  a95406a );
 a95418a <=( A167  and  (not A168) );
 a95419a <=( (not A169)  and  a95418a );
 a95422a <=( A199  and  A166 );
 a95425a <=( A201  and  (not A200) );
 a95426a <=( a95425a  and  a95422a );
 a95427a <=( a95426a  and  a95419a );
 a95430a <=( (not A232)  and  A203 );
 a95433a <=( (not A266)  and  (not A233) );
 a95434a <=( a95433a  and  a95430a );
 a95437a <=( A298  and  (not A267) );
 a95440a <=( (not A302)  and  (not A301) );
 a95441a <=( a95440a  and  a95437a );
 a95442a <=( a95441a  and  a95434a );
 a95446a <=( A167  and  (not A168) );
 a95447a <=( (not A169)  and  a95446a );
 a95450a <=( A199  and  A166 );
 a95453a <=( A201  and  (not A200) );
 a95454a <=( a95453a  and  a95450a );
 a95455a <=( a95454a  and  a95447a );
 a95458a <=( (not A232)  and  A203 );
 a95461a <=( (not A265)  and  (not A233) );
 a95462a <=( a95461a  and  a95458a );
 a95465a <=( A298  and  (not A266) );
 a95468a <=( (not A302)  and  (not A301) );
 a95469a <=( a95468a  and  a95465a );
 a95470a <=( a95469a  and  a95462a );
 a95474a <=( A167  and  (not A169) );
 a95475a <=( A170  and  a95474a );
 a95478a <=( A199  and  (not A166) );
 a95481a <=( (not A233)  and  A200 );
 a95482a <=( a95481a  and  a95478a );
 a95483a <=( a95482a  and  a95475a );
 a95486a <=( (not A236)  and  (not A235) );
 a95489a <=( (not A268)  and  (not A266) );
 a95490a <=( a95489a  and  a95486a );
 a95493a <=( A298  and  (not A269) );
 a95496a <=( (not A302)  and  (not A301) );
 a95497a <=( a95496a  and  a95493a );
 a95498a <=( a95497a  and  a95490a );
 a95502a <=( A167  and  (not A169) );
 a95503a <=( A170  and  a95502a );
 a95506a <=( (not A200)  and  (not A166) );
 a95509a <=( (not A203)  and  (not A202) );
 a95510a <=( a95509a  and  a95506a );
 a95511a <=( a95510a  and  a95503a );
 a95514a <=( A233  and  A232 );
 a95517a <=( (not A268)  and  A265 );
 a95518a <=( a95517a  and  a95514a );
 a95521a <=( (not A299)  and  (not A269) );
 a95524a <=( (not A302)  and  (not A301) );
 a95525a <=( a95524a  and  a95521a );
 a95526a <=( a95525a  and  a95518a );
 a95530a <=( A167  and  (not A169) );
 a95531a <=( A170  and  a95530a );
 a95534a <=( (not A200)  and  (not A166) );
 a95537a <=( (not A203)  and  (not A202) );
 a95538a <=( a95537a  and  a95534a );
 a95539a <=( a95538a  and  a95531a );
 a95542a <=( (not A235)  and  (not A233) );
 a95545a <=( A265  and  (not A236) );
 a95546a <=( a95545a  and  a95542a );
 a95549a <=( A298  and  A266 );
 a95552a <=( (not A302)  and  (not A301) );
 a95553a <=( a95552a  and  a95549a );
 a95554a <=( a95553a  and  a95546a );
 a95558a <=( A167  and  (not A169) );
 a95559a <=( A170  and  a95558a );
 a95562a <=( (not A200)  and  (not A166) );
 a95565a <=( (not A203)  and  (not A202) );
 a95566a <=( a95565a  and  a95562a );
 a95567a <=( a95566a  and  a95559a );
 a95570a <=( (not A235)  and  (not A233) );
 a95573a <=( (not A266)  and  (not A236) );
 a95574a <=( a95573a  and  a95570a );
 a95577a <=( (not A269)  and  (not A268) );
 a95580a <=( (not A300)  and  A298 );
 a95581a <=( a95580a  and  a95577a );
 a95582a <=( a95581a  and  a95574a );
 a95586a <=( A167  and  (not A169) );
 a95587a <=( A170  and  a95586a );
 a95590a <=( (not A200)  and  (not A166) );
 a95593a <=( (not A203)  and  (not A202) );
 a95594a <=( a95593a  and  a95590a );
 a95595a <=( a95594a  and  a95587a );
 a95598a <=( (not A235)  and  (not A233) );
 a95601a <=( (not A266)  and  (not A236) );
 a95602a <=( a95601a  and  a95598a );
 a95605a <=( (not A269)  and  (not A268) );
 a95608a <=( A299  and  A298 );
 a95609a <=( a95608a  and  a95605a );
 a95610a <=( a95609a  and  a95602a );
 a95614a <=( A167  and  (not A169) );
 a95615a <=( A170  and  a95614a );
 a95618a <=( (not A200)  and  (not A166) );
 a95621a <=( (not A203)  and  (not A202) );
 a95622a <=( a95621a  and  a95618a );
 a95623a <=( a95622a  and  a95615a );
 a95626a <=( (not A235)  and  (not A233) );
 a95629a <=( (not A266)  and  (not A236) );
 a95630a <=( a95629a  and  a95626a );
 a95633a <=( (not A269)  and  (not A268) );
 a95636a <=( (not A299)  and  (not A298) );
 a95637a <=( a95636a  and  a95633a );
 a95638a <=( a95637a  and  a95630a );
 a95642a <=( A167  and  (not A169) );
 a95643a <=( A170  and  a95642a );
 a95646a <=( (not A200)  and  (not A166) );
 a95649a <=( (not A203)  and  (not A202) );
 a95650a <=( a95649a  and  a95646a );
 a95651a <=( a95650a  and  a95643a );
 a95654a <=( (not A235)  and  (not A233) );
 a95657a <=( (not A266)  and  (not A236) );
 a95658a <=( a95657a  and  a95654a );
 a95661a <=( A298  and  (not A267) );
 a95664a <=( (not A302)  and  (not A301) );
 a95665a <=( a95664a  and  a95661a );
 a95666a <=( a95665a  and  a95658a );
 a95670a <=( A167  and  (not A169) );
 a95671a <=( A170  and  a95670a );
 a95674a <=( (not A200)  and  (not A166) );
 a95677a <=( (not A203)  and  (not A202) );
 a95678a <=( a95677a  and  a95674a );
 a95679a <=( a95678a  and  a95671a );
 a95682a <=( (not A235)  and  (not A233) );
 a95685a <=( (not A265)  and  (not A236) );
 a95686a <=( a95685a  and  a95682a );
 a95689a <=( A298  and  (not A266) );
 a95692a <=( (not A302)  and  (not A301) );
 a95693a <=( a95692a  and  a95689a );
 a95694a <=( a95693a  and  a95686a );
 a95698a <=( A167  and  (not A169) );
 a95699a <=( A170  and  a95698a );
 a95702a <=( (not A200)  and  (not A166) );
 a95705a <=( (not A203)  and  (not A202) );
 a95706a <=( a95705a  and  a95702a );
 a95707a <=( a95706a  and  a95699a );
 a95710a <=( (not A234)  and  (not A233) );
 a95713a <=( (not A268)  and  (not A266) );
 a95714a <=( a95713a  and  a95710a );
 a95717a <=( A298  and  (not A269) );
 a95720a <=( (not A302)  and  (not A301) );
 a95721a <=( a95720a  and  a95717a );
 a95722a <=( a95721a  and  a95714a );
 a95726a <=( A167  and  (not A169) );
 a95727a <=( A170  and  a95726a );
 a95730a <=( (not A200)  and  (not A166) );
 a95733a <=( (not A203)  and  (not A202) );
 a95734a <=( a95733a  and  a95730a );
 a95735a <=( a95734a  and  a95727a );
 a95738a <=( (not A233)  and  A232 );
 a95741a <=( A235  and  A234 );
 a95742a <=( a95741a  and  a95738a );
 a95745a <=( (not A299)  and  A298 );
 a95748a <=( A301  and  A300 );
 a95749a <=( a95748a  and  a95745a );
 a95750a <=( a95749a  and  a95742a );
 a95754a <=( A167  and  (not A169) );
 a95755a <=( A170  and  a95754a );
 a95758a <=( (not A200)  and  (not A166) );
 a95761a <=( (not A203)  and  (not A202) );
 a95762a <=( a95761a  and  a95758a );
 a95763a <=( a95762a  and  a95755a );
 a95766a <=( (not A233)  and  A232 );
 a95769a <=( A235  and  A234 );
 a95770a <=( a95769a  and  a95766a );
 a95773a <=( (not A299)  and  A298 );
 a95776a <=( A302  and  A300 );
 a95777a <=( a95776a  and  a95773a );
 a95778a <=( a95777a  and  a95770a );
 a95782a <=( A167  and  (not A169) );
 a95783a <=( A170  and  a95782a );
 a95786a <=( (not A200)  and  (not A166) );
 a95789a <=( (not A203)  and  (not A202) );
 a95790a <=( a95789a  and  a95786a );
 a95791a <=( a95790a  and  a95783a );
 a95794a <=( (not A233)  and  A232 );
 a95797a <=( A235  and  A234 );
 a95798a <=( a95797a  and  a95794a );
 a95801a <=( (not A266)  and  A265 );
 a95804a <=( A268  and  A267 );
 a95805a <=( a95804a  and  a95801a );
 a95806a <=( a95805a  and  a95798a );
 a95810a <=( A167  and  (not A169) );
 a95811a <=( A170  and  a95810a );
 a95814a <=( (not A200)  and  (not A166) );
 a95817a <=( (not A203)  and  (not A202) );
 a95818a <=( a95817a  and  a95814a );
 a95819a <=( a95818a  and  a95811a );
 a95822a <=( (not A233)  and  A232 );
 a95825a <=( A235  and  A234 );
 a95826a <=( a95825a  and  a95822a );
 a95829a <=( (not A266)  and  A265 );
 a95832a <=( A269  and  A267 );
 a95833a <=( a95832a  and  a95829a );
 a95834a <=( a95833a  and  a95826a );
 a95838a <=( A167  and  (not A169) );
 a95839a <=( A170  and  a95838a );
 a95842a <=( (not A200)  and  (not A166) );
 a95845a <=( (not A203)  and  (not A202) );
 a95846a <=( a95845a  and  a95842a );
 a95847a <=( a95846a  and  a95839a );
 a95850a <=( (not A233)  and  A232 );
 a95853a <=( A236  and  A234 );
 a95854a <=( a95853a  and  a95850a );
 a95857a <=( (not A299)  and  A298 );
 a95860a <=( A301  and  A300 );
 a95861a <=( a95860a  and  a95857a );
 a95862a <=( a95861a  and  a95854a );
 a95866a <=( A167  and  (not A169) );
 a95867a <=( A170  and  a95866a );
 a95870a <=( (not A200)  and  (not A166) );
 a95873a <=( (not A203)  and  (not A202) );
 a95874a <=( a95873a  and  a95870a );
 a95875a <=( a95874a  and  a95867a );
 a95878a <=( (not A233)  and  A232 );
 a95881a <=( A236  and  A234 );
 a95882a <=( a95881a  and  a95878a );
 a95885a <=( (not A299)  and  A298 );
 a95888a <=( A302  and  A300 );
 a95889a <=( a95888a  and  a95885a );
 a95890a <=( a95889a  and  a95882a );
 a95894a <=( A167  and  (not A169) );
 a95895a <=( A170  and  a95894a );
 a95898a <=( (not A200)  and  (not A166) );
 a95901a <=( (not A203)  and  (not A202) );
 a95902a <=( a95901a  and  a95898a );
 a95903a <=( a95902a  and  a95895a );
 a95906a <=( (not A233)  and  A232 );
 a95909a <=( A236  and  A234 );
 a95910a <=( a95909a  and  a95906a );
 a95913a <=( (not A266)  and  A265 );
 a95916a <=( A268  and  A267 );
 a95917a <=( a95916a  and  a95913a );
 a95918a <=( a95917a  and  a95910a );
 a95922a <=( A167  and  (not A169) );
 a95923a <=( A170  and  a95922a );
 a95926a <=( (not A200)  and  (not A166) );
 a95929a <=( (not A203)  and  (not A202) );
 a95930a <=( a95929a  and  a95926a );
 a95931a <=( a95930a  and  a95923a );
 a95934a <=( (not A233)  and  A232 );
 a95937a <=( A236  and  A234 );
 a95938a <=( a95937a  and  a95934a );
 a95941a <=( (not A266)  and  A265 );
 a95944a <=( A269  and  A267 );
 a95945a <=( a95944a  and  a95941a );
 a95946a <=( a95945a  and  a95938a );
 a95950a <=( A167  and  (not A169) );
 a95951a <=( A170  and  a95950a );
 a95954a <=( (not A200)  and  (not A166) );
 a95957a <=( (not A203)  and  (not A202) );
 a95958a <=( a95957a  and  a95954a );
 a95959a <=( a95958a  and  a95951a );
 a95962a <=( (not A233)  and  (not A232) );
 a95965a <=( (not A268)  and  (not A266) );
 a95966a <=( a95965a  and  a95962a );
 a95969a <=( A298  and  (not A269) );
 a95972a <=( (not A302)  and  (not A301) );
 a95973a <=( a95972a  and  a95969a );
 a95974a <=( a95973a  and  a95966a );
 a95978a <=( A167  and  (not A169) );
 a95979a <=( A170  and  a95978a );
 a95982a <=( (not A200)  and  (not A166) );
 a95985a <=( (not A233)  and  (not A201) );
 a95986a <=( a95985a  and  a95982a );
 a95987a <=( a95986a  and  a95979a );
 a95990a <=( (not A236)  and  (not A235) );
 a95993a <=( (not A268)  and  (not A266) );
 a95994a <=( a95993a  and  a95990a );
 a95997a <=( A298  and  (not A269) );
 a96000a <=( (not A302)  and  (not A301) );
 a96001a <=( a96000a  and  a95997a );
 a96002a <=( a96001a  and  a95994a );
 a96006a <=( A167  and  (not A169) );
 a96007a <=( A170  and  a96006a );
 a96010a <=( (not A199)  and  (not A166) );
 a96013a <=( (not A233)  and  (not A200) );
 a96014a <=( a96013a  and  a96010a );
 a96015a <=( a96014a  and  a96007a );
 a96018a <=( (not A236)  and  (not A235) );
 a96021a <=( (not A268)  and  (not A266) );
 a96022a <=( a96021a  and  a96018a );
 a96025a <=( A298  and  (not A269) );
 a96028a <=( (not A302)  and  (not A301) );
 a96029a <=( a96028a  and  a96025a );
 a96030a <=( a96029a  and  a96022a );
 a96034a <=( (not A167)  and  (not A169) );
 a96035a <=( A170  and  a96034a );
 a96038a <=( A199  and  A166 );
 a96041a <=( (not A233)  and  A200 );
 a96042a <=( a96041a  and  a96038a );
 a96043a <=( a96042a  and  a96035a );
 a96046a <=( (not A236)  and  (not A235) );
 a96049a <=( (not A268)  and  (not A266) );
 a96050a <=( a96049a  and  a96046a );
 a96053a <=( A298  and  (not A269) );
 a96056a <=( (not A302)  and  (not A301) );
 a96057a <=( a96056a  and  a96053a );
 a96058a <=( a96057a  and  a96050a );
 a96062a <=( (not A167)  and  (not A169) );
 a96063a <=( A170  and  a96062a );
 a96066a <=( (not A200)  and  A166 );
 a96069a <=( (not A203)  and  (not A202) );
 a96070a <=( a96069a  and  a96066a );
 a96071a <=( a96070a  and  a96063a );
 a96074a <=( A233  and  A232 );
 a96077a <=( (not A268)  and  A265 );
 a96078a <=( a96077a  and  a96074a );
 a96081a <=( (not A299)  and  (not A269) );
 a96084a <=( (not A302)  and  (not A301) );
 a96085a <=( a96084a  and  a96081a );
 a96086a <=( a96085a  and  a96078a );
 a96090a <=( (not A167)  and  (not A169) );
 a96091a <=( A170  and  a96090a );
 a96094a <=( (not A200)  and  A166 );
 a96097a <=( (not A203)  and  (not A202) );
 a96098a <=( a96097a  and  a96094a );
 a96099a <=( a96098a  and  a96091a );
 a96102a <=( (not A235)  and  (not A233) );
 a96105a <=( A265  and  (not A236) );
 a96106a <=( a96105a  and  a96102a );
 a96109a <=( A298  and  A266 );
 a96112a <=( (not A302)  and  (not A301) );
 a96113a <=( a96112a  and  a96109a );
 a96114a <=( a96113a  and  a96106a );
 a96118a <=( (not A167)  and  (not A169) );
 a96119a <=( A170  and  a96118a );
 a96122a <=( (not A200)  and  A166 );
 a96125a <=( (not A203)  and  (not A202) );
 a96126a <=( a96125a  and  a96122a );
 a96127a <=( a96126a  and  a96119a );
 a96130a <=( (not A235)  and  (not A233) );
 a96133a <=( (not A266)  and  (not A236) );
 a96134a <=( a96133a  and  a96130a );
 a96137a <=( (not A269)  and  (not A268) );
 a96140a <=( (not A300)  and  A298 );
 a96141a <=( a96140a  and  a96137a );
 a96142a <=( a96141a  and  a96134a );
 a96146a <=( (not A167)  and  (not A169) );
 a96147a <=( A170  and  a96146a );
 a96150a <=( (not A200)  and  A166 );
 a96153a <=( (not A203)  and  (not A202) );
 a96154a <=( a96153a  and  a96150a );
 a96155a <=( a96154a  and  a96147a );
 a96158a <=( (not A235)  and  (not A233) );
 a96161a <=( (not A266)  and  (not A236) );
 a96162a <=( a96161a  and  a96158a );
 a96165a <=( (not A269)  and  (not A268) );
 a96168a <=( A299  and  A298 );
 a96169a <=( a96168a  and  a96165a );
 a96170a <=( a96169a  and  a96162a );
 a96174a <=( (not A167)  and  (not A169) );
 a96175a <=( A170  and  a96174a );
 a96178a <=( (not A200)  and  A166 );
 a96181a <=( (not A203)  and  (not A202) );
 a96182a <=( a96181a  and  a96178a );
 a96183a <=( a96182a  and  a96175a );
 a96186a <=( (not A235)  and  (not A233) );
 a96189a <=( (not A266)  and  (not A236) );
 a96190a <=( a96189a  and  a96186a );
 a96193a <=( (not A269)  and  (not A268) );
 a96196a <=( (not A299)  and  (not A298) );
 a96197a <=( a96196a  and  a96193a );
 a96198a <=( a96197a  and  a96190a );
 a96202a <=( (not A167)  and  (not A169) );
 a96203a <=( A170  and  a96202a );
 a96206a <=( (not A200)  and  A166 );
 a96209a <=( (not A203)  and  (not A202) );
 a96210a <=( a96209a  and  a96206a );
 a96211a <=( a96210a  and  a96203a );
 a96214a <=( (not A235)  and  (not A233) );
 a96217a <=( (not A266)  and  (not A236) );
 a96218a <=( a96217a  and  a96214a );
 a96221a <=( A298  and  (not A267) );
 a96224a <=( (not A302)  and  (not A301) );
 a96225a <=( a96224a  and  a96221a );
 a96226a <=( a96225a  and  a96218a );
 a96230a <=( (not A167)  and  (not A169) );
 a96231a <=( A170  and  a96230a );
 a96234a <=( (not A200)  and  A166 );
 a96237a <=( (not A203)  and  (not A202) );
 a96238a <=( a96237a  and  a96234a );
 a96239a <=( a96238a  and  a96231a );
 a96242a <=( (not A235)  and  (not A233) );
 a96245a <=( (not A265)  and  (not A236) );
 a96246a <=( a96245a  and  a96242a );
 a96249a <=( A298  and  (not A266) );
 a96252a <=( (not A302)  and  (not A301) );
 a96253a <=( a96252a  and  a96249a );
 a96254a <=( a96253a  and  a96246a );
 a96258a <=( (not A167)  and  (not A169) );
 a96259a <=( A170  and  a96258a );
 a96262a <=( (not A200)  and  A166 );
 a96265a <=( (not A203)  and  (not A202) );
 a96266a <=( a96265a  and  a96262a );
 a96267a <=( a96266a  and  a96259a );
 a96270a <=( (not A234)  and  (not A233) );
 a96273a <=( (not A268)  and  (not A266) );
 a96274a <=( a96273a  and  a96270a );
 a96277a <=( A298  and  (not A269) );
 a96280a <=( (not A302)  and  (not A301) );
 a96281a <=( a96280a  and  a96277a );
 a96282a <=( a96281a  and  a96274a );
 a96286a <=( (not A167)  and  (not A169) );
 a96287a <=( A170  and  a96286a );
 a96290a <=( (not A200)  and  A166 );
 a96293a <=( (not A203)  and  (not A202) );
 a96294a <=( a96293a  and  a96290a );
 a96295a <=( a96294a  and  a96287a );
 a96298a <=( (not A233)  and  A232 );
 a96301a <=( A235  and  A234 );
 a96302a <=( a96301a  and  a96298a );
 a96305a <=( (not A299)  and  A298 );
 a96308a <=( A301  and  A300 );
 a96309a <=( a96308a  and  a96305a );
 a96310a <=( a96309a  and  a96302a );
 a96314a <=( (not A167)  and  (not A169) );
 a96315a <=( A170  and  a96314a );
 a96318a <=( (not A200)  and  A166 );
 a96321a <=( (not A203)  and  (not A202) );
 a96322a <=( a96321a  and  a96318a );
 a96323a <=( a96322a  and  a96315a );
 a96326a <=( (not A233)  and  A232 );
 a96329a <=( A235  and  A234 );
 a96330a <=( a96329a  and  a96326a );
 a96333a <=( (not A299)  and  A298 );
 a96336a <=( A302  and  A300 );
 a96337a <=( a96336a  and  a96333a );
 a96338a <=( a96337a  and  a96330a );
 a96342a <=( (not A167)  and  (not A169) );
 a96343a <=( A170  and  a96342a );
 a96346a <=( (not A200)  and  A166 );
 a96349a <=( (not A203)  and  (not A202) );
 a96350a <=( a96349a  and  a96346a );
 a96351a <=( a96350a  and  a96343a );
 a96354a <=( (not A233)  and  A232 );
 a96357a <=( A235  and  A234 );
 a96358a <=( a96357a  and  a96354a );
 a96361a <=( (not A266)  and  A265 );
 a96364a <=( A268  and  A267 );
 a96365a <=( a96364a  and  a96361a );
 a96366a <=( a96365a  and  a96358a );
 a96370a <=( (not A167)  and  (not A169) );
 a96371a <=( A170  and  a96370a );
 a96374a <=( (not A200)  and  A166 );
 a96377a <=( (not A203)  and  (not A202) );
 a96378a <=( a96377a  and  a96374a );
 a96379a <=( a96378a  and  a96371a );
 a96382a <=( (not A233)  and  A232 );
 a96385a <=( A235  and  A234 );
 a96386a <=( a96385a  and  a96382a );
 a96389a <=( (not A266)  and  A265 );
 a96392a <=( A269  and  A267 );
 a96393a <=( a96392a  and  a96389a );
 a96394a <=( a96393a  and  a96386a );
 a96398a <=( (not A167)  and  (not A169) );
 a96399a <=( A170  and  a96398a );
 a96402a <=( (not A200)  and  A166 );
 a96405a <=( (not A203)  and  (not A202) );
 a96406a <=( a96405a  and  a96402a );
 a96407a <=( a96406a  and  a96399a );
 a96410a <=( (not A233)  and  A232 );
 a96413a <=( A236  and  A234 );
 a96414a <=( a96413a  and  a96410a );
 a96417a <=( (not A299)  and  A298 );
 a96420a <=( A301  and  A300 );
 a96421a <=( a96420a  and  a96417a );
 a96422a <=( a96421a  and  a96414a );
 a96426a <=( (not A167)  and  (not A169) );
 a96427a <=( A170  and  a96426a );
 a96430a <=( (not A200)  and  A166 );
 a96433a <=( (not A203)  and  (not A202) );
 a96434a <=( a96433a  and  a96430a );
 a96435a <=( a96434a  and  a96427a );
 a96438a <=( (not A233)  and  A232 );
 a96441a <=( A236  and  A234 );
 a96442a <=( a96441a  and  a96438a );
 a96445a <=( (not A299)  and  A298 );
 a96448a <=( A302  and  A300 );
 a96449a <=( a96448a  and  a96445a );
 a96450a <=( a96449a  and  a96442a );
 a96454a <=( (not A167)  and  (not A169) );
 a96455a <=( A170  and  a96454a );
 a96458a <=( (not A200)  and  A166 );
 a96461a <=( (not A203)  and  (not A202) );
 a96462a <=( a96461a  and  a96458a );
 a96463a <=( a96462a  and  a96455a );
 a96466a <=( (not A233)  and  A232 );
 a96469a <=( A236  and  A234 );
 a96470a <=( a96469a  and  a96466a );
 a96473a <=( (not A266)  and  A265 );
 a96476a <=( A268  and  A267 );
 a96477a <=( a96476a  and  a96473a );
 a96478a <=( a96477a  and  a96470a );
 a96482a <=( (not A167)  and  (not A169) );
 a96483a <=( A170  and  a96482a );
 a96486a <=( (not A200)  and  A166 );
 a96489a <=( (not A203)  and  (not A202) );
 a96490a <=( a96489a  and  a96486a );
 a96491a <=( a96490a  and  a96483a );
 a96494a <=( (not A233)  and  A232 );
 a96497a <=( A236  and  A234 );
 a96498a <=( a96497a  and  a96494a );
 a96501a <=( (not A266)  and  A265 );
 a96504a <=( A269  and  A267 );
 a96505a <=( a96504a  and  a96501a );
 a96506a <=( a96505a  and  a96498a );
 a96510a <=( (not A167)  and  (not A169) );
 a96511a <=( A170  and  a96510a );
 a96514a <=( (not A200)  and  A166 );
 a96517a <=( (not A203)  and  (not A202) );
 a96518a <=( a96517a  and  a96514a );
 a96519a <=( a96518a  and  a96511a );
 a96522a <=( (not A233)  and  (not A232) );
 a96525a <=( (not A268)  and  (not A266) );
 a96526a <=( a96525a  and  a96522a );
 a96529a <=( A298  and  (not A269) );
 a96532a <=( (not A302)  and  (not A301) );
 a96533a <=( a96532a  and  a96529a );
 a96534a <=( a96533a  and  a96526a );
 a96538a <=( (not A167)  and  (not A169) );
 a96539a <=( A170  and  a96538a );
 a96542a <=( (not A200)  and  A166 );
 a96545a <=( (not A233)  and  (not A201) );
 a96546a <=( a96545a  and  a96542a );
 a96547a <=( a96546a  and  a96539a );
 a96550a <=( (not A236)  and  (not A235) );
 a96553a <=( (not A268)  and  (not A266) );
 a96554a <=( a96553a  and  a96550a );
 a96557a <=( A298  and  (not A269) );
 a96560a <=( (not A302)  and  (not A301) );
 a96561a <=( a96560a  and  a96557a );
 a96562a <=( a96561a  and  a96554a );
 a96566a <=( (not A167)  and  (not A169) );
 a96567a <=( A170  and  a96566a );
 a96570a <=( (not A199)  and  A166 );
 a96573a <=( (not A233)  and  (not A200) );
 a96574a <=( a96573a  and  a96570a );
 a96575a <=( a96574a  and  a96567a );
 a96578a <=( (not A236)  and  (not A235) );
 a96581a <=( (not A268)  and  (not A266) );
 a96582a <=( a96581a  and  a96578a );
 a96585a <=( A298  and  (not A269) );
 a96588a <=( (not A302)  and  (not A301) );
 a96589a <=( a96588a  and  a96585a );
 a96590a <=( a96589a  and  a96582a );
 a96594a <=( (not A168)  and  (not A169) );
 a96595a <=( (not A170)  and  a96594a );
 a96598a <=( (not A200)  and  A199 );
 a96601a <=( A202  and  A201 );
 a96602a <=( a96601a  and  a96598a );
 a96603a <=( a96602a  and  a96595a );
 a96606a <=( A233  and  A232 );
 a96609a <=( (not A268)  and  A265 );
 a96610a <=( a96609a  and  a96606a );
 a96613a <=( (not A299)  and  (not A269) );
 a96616a <=( (not A302)  and  (not A301) );
 a96617a <=( a96616a  and  a96613a );
 a96618a <=( a96617a  and  a96610a );
 a96622a <=( (not A168)  and  (not A169) );
 a96623a <=( (not A170)  and  a96622a );
 a96626a <=( (not A200)  and  A199 );
 a96629a <=( A202  and  A201 );
 a96630a <=( a96629a  and  a96626a );
 a96631a <=( a96630a  and  a96623a );
 a96634a <=( (not A235)  and  (not A233) );
 a96637a <=( A265  and  (not A236) );
 a96638a <=( a96637a  and  a96634a );
 a96641a <=( A298  and  A266 );
 a96644a <=( (not A302)  and  (not A301) );
 a96645a <=( a96644a  and  a96641a );
 a96646a <=( a96645a  and  a96638a );
 a96650a <=( (not A168)  and  (not A169) );
 a96651a <=( (not A170)  and  a96650a );
 a96654a <=( (not A200)  and  A199 );
 a96657a <=( A202  and  A201 );
 a96658a <=( a96657a  and  a96654a );
 a96659a <=( a96658a  and  a96651a );
 a96662a <=( (not A235)  and  (not A233) );
 a96665a <=( (not A266)  and  (not A236) );
 a96666a <=( a96665a  and  a96662a );
 a96669a <=( (not A269)  and  (not A268) );
 a96672a <=( (not A300)  and  A298 );
 a96673a <=( a96672a  and  a96669a );
 a96674a <=( a96673a  and  a96666a );
 a96678a <=( (not A168)  and  (not A169) );
 a96679a <=( (not A170)  and  a96678a );
 a96682a <=( (not A200)  and  A199 );
 a96685a <=( A202  and  A201 );
 a96686a <=( a96685a  and  a96682a );
 a96687a <=( a96686a  and  a96679a );
 a96690a <=( (not A235)  and  (not A233) );
 a96693a <=( (not A266)  and  (not A236) );
 a96694a <=( a96693a  and  a96690a );
 a96697a <=( (not A269)  and  (not A268) );
 a96700a <=( A299  and  A298 );
 a96701a <=( a96700a  and  a96697a );
 a96702a <=( a96701a  and  a96694a );
 a96706a <=( (not A168)  and  (not A169) );
 a96707a <=( (not A170)  and  a96706a );
 a96710a <=( (not A200)  and  A199 );
 a96713a <=( A202  and  A201 );
 a96714a <=( a96713a  and  a96710a );
 a96715a <=( a96714a  and  a96707a );
 a96718a <=( (not A235)  and  (not A233) );
 a96721a <=( (not A266)  and  (not A236) );
 a96722a <=( a96721a  and  a96718a );
 a96725a <=( (not A269)  and  (not A268) );
 a96728a <=( (not A299)  and  (not A298) );
 a96729a <=( a96728a  and  a96725a );
 a96730a <=( a96729a  and  a96722a );
 a96734a <=( (not A168)  and  (not A169) );
 a96735a <=( (not A170)  and  a96734a );
 a96738a <=( (not A200)  and  A199 );
 a96741a <=( A202  and  A201 );
 a96742a <=( a96741a  and  a96738a );
 a96743a <=( a96742a  and  a96735a );
 a96746a <=( (not A235)  and  (not A233) );
 a96749a <=( (not A266)  and  (not A236) );
 a96750a <=( a96749a  and  a96746a );
 a96753a <=( A298  and  (not A267) );
 a96756a <=( (not A302)  and  (not A301) );
 a96757a <=( a96756a  and  a96753a );
 a96758a <=( a96757a  and  a96750a );
 a96762a <=( (not A168)  and  (not A169) );
 a96763a <=( (not A170)  and  a96762a );
 a96766a <=( (not A200)  and  A199 );
 a96769a <=( A202  and  A201 );
 a96770a <=( a96769a  and  a96766a );
 a96771a <=( a96770a  and  a96763a );
 a96774a <=( (not A235)  and  (not A233) );
 a96777a <=( (not A265)  and  (not A236) );
 a96778a <=( a96777a  and  a96774a );
 a96781a <=( A298  and  (not A266) );
 a96784a <=( (not A302)  and  (not A301) );
 a96785a <=( a96784a  and  a96781a );
 a96786a <=( a96785a  and  a96778a );
 a96790a <=( (not A168)  and  (not A169) );
 a96791a <=( (not A170)  and  a96790a );
 a96794a <=( (not A200)  and  A199 );
 a96797a <=( A202  and  A201 );
 a96798a <=( a96797a  and  a96794a );
 a96799a <=( a96798a  and  a96791a );
 a96802a <=( (not A234)  and  (not A233) );
 a96805a <=( (not A268)  and  (not A266) );
 a96806a <=( a96805a  and  a96802a );
 a96809a <=( A298  and  (not A269) );
 a96812a <=( (not A302)  and  (not A301) );
 a96813a <=( a96812a  and  a96809a );
 a96814a <=( a96813a  and  a96806a );
 a96818a <=( (not A168)  and  (not A169) );
 a96819a <=( (not A170)  and  a96818a );
 a96822a <=( (not A200)  and  A199 );
 a96825a <=( A202  and  A201 );
 a96826a <=( a96825a  and  a96822a );
 a96827a <=( a96826a  and  a96819a );
 a96830a <=( (not A233)  and  A232 );
 a96833a <=( A235  and  A234 );
 a96834a <=( a96833a  and  a96830a );
 a96837a <=( (not A299)  and  A298 );
 a96840a <=( A301  and  A300 );
 a96841a <=( a96840a  and  a96837a );
 a96842a <=( a96841a  and  a96834a );
 a96846a <=( (not A168)  and  (not A169) );
 a96847a <=( (not A170)  and  a96846a );
 a96850a <=( (not A200)  and  A199 );
 a96853a <=( A202  and  A201 );
 a96854a <=( a96853a  and  a96850a );
 a96855a <=( a96854a  and  a96847a );
 a96858a <=( (not A233)  and  A232 );
 a96861a <=( A235  and  A234 );
 a96862a <=( a96861a  and  a96858a );
 a96865a <=( (not A299)  and  A298 );
 a96868a <=( A302  and  A300 );
 a96869a <=( a96868a  and  a96865a );
 a96870a <=( a96869a  and  a96862a );
 a96874a <=( (not A168)  and  (not A169) );
 a96875a <=( (not A170)  and  a96874a );
 a96878a <=( (not A200)  and  A199 );
 a96881a <=( A202  and  A201 );
 a96882a <=( a96881a  and  a96878a );
 a96883a <=( a96882a  and  a96875a );
 a96886a <=( (not A233)  and  A232 );
 a96889a <=( A235  and  A234 );
 a96890a <=( a96889a  and  a96886a );
 a96893a <=( (not A266)  and  A265 );
 a96896a <=( A268  and  A267 );
 a96897a <=( a96896a  and  a96893a );
 a96898a <=( a96897a  and  a96890a );
 a96902a <=( (not A168)  and  (not A169) );
 a96903a <=( (not A170)  and  a96902a );
 a96906a <=( (not A200)  and  A199 );
 a96909a <=( A202  and  A201 );
 a96910a <=( a96909a  and  a96906a );
 a96911a <=( a96910a  and  a96903a );
 a96914a <=( (not A233)  and  A232 );
 a96917a <=( A235  and  A234 );
 a96918a <=( a96917a  and  a96914a );
 a96921a <=( (not A266)  and  A265 );
 a96924a <=( A269  and  A267 );
 a96925a <=( a96924a  and  a96921a );
 a96926a <=( a96925a  and  a96918a );
 a96930a <=( (not A168)  and  (not A169) );
 a96931a <=( (not A170)  and  a96930a );
 a96934a <=( (not A200)  and  A199 );
 a96937a <=( A202  and  A201 );
 a96938a <=( a96937a  and  a96934a );
 a96939a <=( a96938a  and  a96931a );
 a96942a <=( (not A233)  and  A232 );
 a96945a <=( A236  and  A234 );
 a96946a <=( a96945a  and  a96942a );
 a96949a <=( (not A299)  and  A298 );
 a96952a <=( A301  and  A300 );
 a96953a <=( a96952a  and  a96949a );
 a96954a <=( a96953a  and  a96946a );
 a96958a <=( (not A168)  and  (not A169) );
 a96959a <=( (not A170)  and  a96958a );
 a96962a <=( (not A200)  and  A199 );
 a96965a <=( A202  and  A201 );
 a96966a <=( a96965a  and  a96962a );
 a96967a <=( a96966a  and  a96959a );
 a96970a <=( (not A233)  and  A232 );
 a96973a <=( A236  and  A234 );
 a96974a <=( a96973a  and  a96970a );
 a96977a <=( (not A299)  and  A298 );
 a96980a <=( A302  and  A300 );
 a96981a <=( a96980a  and  a96977a );
 a96982a <=( a96981a  and  a96974a );
 a96986a <=( (not A168)  and  (not A169) );
 a96987a <=( (not A170)  and  a96986a );
 a96990a <=( (not A200)  and  A199 );
 a96993a <=( A202  and  A201 );
 a96994a <=( a96993a  and  a96990a );
 a96995a <=( a96994a  and  a96987a );
 a96998a <=( (not A233)  and  A232 );
 a97001a <=( A236  and  A234 );
 a97002a <=( a97001a  and  a96998a );
 a97005a <=( (not A266)  and  A265 );
 a97008a <=( A268  and  A267 );
 a97009a <=( a97008a  and  a97005a );
 a97010a <=( a97009a  and  a97002a );
 a97014a <=( (not A168)  and  (not A169) );
 a97015a <=( (not A170)  and  a97014a );
 a97018a <=( (not A200)  and  A199 );
 a97021a <=( A202  and  A201 );
 a97022a <=( a97021a  and  a97018a );
 a97023a <=( a97022a  and  a97015a );
 a97026a <=( (not A233)  and  A232 );
 a97029a <=( A236  and  A234 );
 a97030a <=( a97029a  and  a97026a );
 a97033a <=( (not A266)  and  A265 );
 a97036a <=( A269  and  A267 );
 a97037a <=( a97036a  and  a97033a );
 a97038a <=( a97037a  and  a97030a );
 a97042a <=( (not A168)  and  (not A169) );
 a97043a <=( (not A170)  and  a97042a );
 a97046a <=( (not A200)  and  A199 );
 a97049a <=( A202  and  A201 );
 a97050a <=( a97049a  and  a97046a );
 a97051a <=( a97050a  and  a97043a );
 a97054a <=( (not A233)  and  (not A232) );
 a97057a <=( (not A268)  and  (not A266) );
 a97058a <=( a97057a  and  a97054a );
 a97061a <=( A298  and  (not A269) );
 a97064a <=( (not A302)  and  (not A301) );
 a97065a <=( a97064a  and  a97061a );
 a97066a <=( a97065a  and  a97058a );
 a97070a <=( (not A168)  and  (not A169) );
 a97071a <=( (not A170)  and  a97070a );
 a97074a <=( (not A200)  and  A199 );
 a97077a <=( A203  and  A201 );
 a97078a <=( a97077a  and  a97074a );
 a97079a <=( a97078a  and  a97071a );
 a97082a <=( A233  and  A232 );
 a97085a <=( (not A268)  and  A265 );
 a97086a <=( a97085a  and  a97082a );
 a97089a <=( (not A299)  and  (not A269) );
 a97092a <=( (not A302)  and  (not A301) );
 a97093a <=( a97092a  and  a97089a );
 a97094a <=( a97093a  and  a97086a );
 a97098a <=( (not A168)  and  (not A169) );
 a97099a <=( (not A170)  and  a97098a );
 a97102a <=( (not A200)  and  A199 );
 a97105a <=( A203  and  A201 );
 a97106a <=( a97105a  and  a97102a );
 a97107a <=( a97106a  and  a97099a );
 a97110a <=( (not A235)  and  (not A233) );
 a97113a <=( A265  and  (not A236) );
 a97114a <=( a97113a  and  a97110a );
 a97117a <=( A298  and  A266 );
 a97120a <=( (not A302)  and  (not A301) );
 a97121a <=( a97120a  and  a97117a );
 a97122a <=( a97121a  and  a97114a );
 a97126a <=( (not A168)  and  (not A169) );
 a97127a <=( (not A170)  and  a97126a );
 a97130a <=( (not A200)  and  A199 );
 a97133a <=( A203  and  A201 );
 a97134a <=( a97133a  and  a97130a );
 a97135a <=( a97134a  and  a97127a );
 a97138a <=( (not A235)  and  (not A233) );
 a97141a <=( (not A266)  and  (not A236) );
 a97142a <=( a97141a  and  a97138a );
 a97145a <=( (not A269)  and  (not A268) );
 a97148a <=( (not A300)  and  A298 );
 a97149a <=( a97148a  and  a97145a );
 a97150a <=( a97149a  and  a97142a );
 a97154a <=( (not A168)  and  (not A169) );
 a97155a <=( (not A170)  and  a97154a );
 a97158a <=( (not A200)  and  A199 );
 a97161a <=( A203  and  A201 );
 a97162a <=( a97161a  and  a97158a );
 a97163a <=( a97162a  and  a97155a );
 a97166a <=( (not A235)  and  (not A233) );
 a97169a <=( (not A266)  and  (not A236) );
 a97170a <=( a97169a  and  a97166a );
 a97173a <=( (not A269)  and  (not A268) );
 a97176a <=( A299  and  A298 );
 a97177a <=( a97176a  and  a97173a );
 a97178a <=( a97177a  and  a97170a );
 a97182a <=( (not A168)  and  (not A169) );
 a97183a <=( (not A170)  and  a97182a );
 a97186a <=( (not A200)  and  A199 );
 a97189a <=( A203  and  A201 );
 a97190a <=( a97189a  and  a97186a );
 a97191a <=( a97190a  and  a97183a );
 a97194a <=( (not A235)  and  (not A233) );
 a97197a <=( (not A266)  and  (not A236) );
 a97198a <=( a97197a  and  a97194a );
 a97201a <=( (not A269)  and  (not A268) );
 a97204a <=( (not A299)  and  (not A298) );
 a97205a <=( a97204a  and  a97201a );
 a97206a <=( a97205a  and  a97198a );
 a97210a <=( (not A168)  and  (not A169) );
 a97211a <=( (not A170)  and  a97210a );
 a97214a <=( (not A200)  and  A199 );
 a97217a <=( A203  and  A201 );
 a97218a <=( a97217a  and  a97214a );
 a97219a <=( a97218a  and  a97211a );
 a97222a <=( (not A235)  and  (not A233) );
 a97225a <=( (not A266)  and  (not A236) );
 a97226a <=( a97225a  and  a97222a );
 a97229a <=( A298  and  (not A267) );
 a97232a <=( (not A302)  and  (not A301) );
 a97233a <=( a97232a  and  a97229a );
 a97234a <=( a97233a  and  a97226a );
 a97238a <=( (not A168)  and  (not A169) );
 a97239a <=( (not A170)  and  a97238a );
 a97242a <=( (not A200)  and  A199 );
 a97245a <=( A203  and  A201 );
 a97246a <=( a97245a  and  a97242a );
 a97247a <=( a97246a  and  a97239a );
 a97250a <=( (not A235)  and  (not A233) );
 a97253a <=( (not A265)  and  (not A236) );
 a97254a <=( a97253a  and  a97250a );
 a97257a <=( A298  and  (not A266) );
 a97260a <=( (not A302)  and  (not A301) );
 a97261a <=( a97260a  and  a97257a );
 a97262a <=( a97261a  and  a97254a );
 a97266a <=( (not A168)  and  (not A169) );
 a97267a <=( (not A170)  and  a97266a );
 a97270a <=( (not A200)  and  A199 );
 a97273a <=( A203  and  A201 );
 a97274a <=( a97273a  and  a97270a );
 a97275a <=( a97274a  and  a97267a );
 a97278a <=( (not A234)  and  (not A233) );
 a97281a <=( (not A268)  and  (not A266) );
 a97282a <=( a97281a  and  a97278a );
 a97285a <=( A298  and  (not A269) );
 a97288a <=( (not A302)  and  (not A301) );
 a97289a <=( a97288a  and  a97285a );
 a97290a <=( a97289a  and  a97282a );
 a97294a <=( (not A168)  and  (not A169) );
 a97295a <=( (not A170)  and  a97294a );
 a97298a <=( (not A200)  and  A199 );
 a97301a <=( A203  and  A201 );
 a97302a <=( a97301a  and  a97298a );
 a97303a <=( a97302a  and  a97295a );
 a97306a <=( (not A233)  and  A232 );
 a97309a <=( A235  and  A234 );
 a97310a <=( a97309a  and  a97306a );
 a97313a <=( (not A299)  and  A298 );
 a97316a <=( A301  and  A300 );
 a97317a <=( a97316a  and  a97313a );
 a97318a <=( a97317a  and  a97310a );
 a97322a <=( (not A168)  and  (not A169) );
 a97323a <=( (not A170)  and  a97322a );
 a97326a <=( (not A200)  and  A199 );
 a97329a <=( A203  and  A201 );
 a97330a <=( a97329a  and  a97326a );
 a97331a <=( a97330a  and  a97323a );
 a97334a <=( (not A233)  and  A232 );
 a97337a <=( A235  and  A234 );
 a97338a <=( a97337a  and  a97334a );
 a97341a <=( (not A299)  and  A298 );
 a97344a <=( A302  and  A300 );
 a97345a <=( a97344a  and  a97341a );
 a97346a <=( a97345a  and  a97338a );
 a97350a <=( (not A168)  and  (not A169) );
 a97351a <=( (not A170)  and  a97350a );
 a97354a <=( (not A200)  and  A199 );
 a97357a <=( A203  and  A201 );
 a97358a <=( a97357a  and  a97354a );
 a97359a <=( a97358a  and  a97351a );
 a97362a <=( (not A233)  and  A232 );
 a97365a <=( A235  and  A234 );
 a97366a <=( a97365a  and  a97362a );
 a97369a <=( (not A266)  and  A265 );
 a97372a <=( A268  and  A267 );
 a97373a <=( a97372a  and  a97369a );
 a97374a <=( a97373a  and  a97366a );
 a97378a <=( (not A168)  and  (not A169) );
 a97379a <=( (not A170)  and  a97378a );
 a97382a <=( (not A200)  and  A199 );
 a97385a <=( A203  and  A201 );
 a97386a <=( a97385a  and  a97382a );
 a97387a <=( a97386a  and  a97379a );
 a97390a <=( (not A233)  and  A232 );
 a97393a <=( A235  and  A234 );
 a97394a <=( a97393a  and  a97390a );
 a97397a <=( (not A266)  and  A265 );
 a97400a <=( A269  and  A267 );
 a97401a <=( a97400a  and  a97397a );
 a97402a <=( a97401a  and  a97394a );
 a97406a <=( (not A168)  and  (not A169) );
 a97407a <=( (not A170)  and  a97406a );
 a97410a <=( (not A200)  and  A199 );
 a97413a <=( A203  and  A201 );
 a97414a <=( a97413a  and  a97410a );
 a97415a <=( a97414a  and  a97407a );
 a97418a <=( (not A233)  and  A232 );
 a97421a <=( A236  and  A234 );
 a97422a <=( a97421a  and  a97418a );
 a97425a <=( (not A299)  and  A298 );
 a97428a <=( A301  and  A300 );
 a97429a <=( a97428a  and  a97425a );
 a97430a <=( a97429a  and  a97422a );
 a97434a <=( (not A168)  and  (not A169) );
 a97435a <=( (not A170)  and  a97434a );
 a97438a <=( (not A200)  and  A199 );
 a97441a <=( A203  and  A201 );
 a97442a <=( a97441a  and  a97438a );
 a97443a <=( a97442a  and  a97435a );
 a97446a <=( (not A233)  and  A232 );
 a97449a <=( A236  and  A234 );
 a97450a <=( a97449a  and  a97446a );
 a97453a <=( (not A299)  and  A298 );
 a97456a <=( A302  and  A300 );
 a97457a <=( a97456a  and  a97453a );
 a97458a <=( a97457a  and  a97450a );
 a97462a <=( (not A168)  and  (not A169) );
 a97463a <=( (not A170)  and  a97462a );
 a97466a <=( (not A200)  and  A199 );
 a97469a <=( A203  and  A201 );
 a97470a <=( a97469a  and  a97466a );
 a97471a <=( a97470a  and  a97463a );
 a97474a <=( (not A233)  and  A232 );
 a97477a <=( A236  and  A234 );
 a97478a <=( a97477a  and  a97474a );
 a97481a <=( (not A266)  and  A265 );
 a97484a <=( A268  and  A267 );
 a97485a <=( a97484a  and  a97481a );
 a97486a <=( a97485a  and  a97478a );
 a97490a <=( (not A168)  and  (not A169) );
 a97491a <=( (not A170)  and  a97490a );
 a97494a <=( (not A200)  and  A199 );
 a97497a <=( A203  and  A201 );
 a97498a <=( a97497a  and  a97494a );
 a97499a <=( a97498a  and  a97491a );
 a97502a <=( (not A233)  and  A232 );
 a97505a <=( A236  and  A234 );
 a97506a <=( a97505a  and  a97502a );
 a97509a <=( (not A266)  and  A265 );
 a97512a <=( A269  and  A267 );
 a97513a <=( a97512a  and  a97509a );
 a97514a <=( a97513a  and  a97506a );
 a97518a <=( (not A168)  and  (not A169) );
 a97519a <=( (not A170)  and  a97518a );
 a97522a <=( (not A200)  and  A199 );
 a97525a <=( A203  and  A201 );
 a97526a <=( a97525a  and  a97522a );
 a97527a <=( a97526a  and  a97519a );
 a97530a <=( (not A233)  and  (not A232) );
 a97533a <=( (not A268)  and  (not A266) );
 a97534a <=( a97533a  and  a97530a );
 a97537a <=( A298  and  (not A269) );
 a97540a <=( (not A302)  and  (not A301) );
 a97541a <=( a97540a  and  a97537a );
 a97542a <=( a97541a  and  a97534a );
 a97545a <=( (not A167)  and  A170 );
 a97548a <=( A199  and  (not A166) );
 a97549a <=( a97548a  and  a97545a );
 a97552a <=( A201  and  (not A200) );
 a97555a <=( (not A233)  and  A202 );
 a97556a <=( a97555a  and  a97552a );
 a97557a <=( a97556a  and  a97549a );
 a97560a <=( (not A236)  and  (not A235) );
 a97563a <=( (not A268)  and  (not A266) );
 a97564a <=( a97563a  and  a97560a );
 a97567a <=( A298  and  (not A269) );
 a97570a <=( (not A302)  and  (not A301) );
 a97571a <=( a97570a  and  a97567a );
 a97572a <=( a97571a  and  a97564a );
 a97575a <=( (not A167)  and  A170 );
 a97578a <=( A199  and  (not A166) );
 a97579a <=( a97578a  and  a97575a );
 a97582a <=( A201  and  (not A200) );
 a97585a <=( (not A233)  and  A203 );
 a97586a <=( a97585a  and  a97582a );
 a97587a <=( a97586a  and  a97579a );
 a97590a <=( (not A236)  and  (not A235) );
 a97593a <=( (not A268)  and  (not A266) );
 a97594a <=( a97593a  and  a97590a );
 a97597a <=( A298  and  (not A269) );
 a97600a <=( (not A302)  and  (not A301) );
 a97601a <=( a97600a  and  a97597a );
 a97602a <=( a97601a  and  a97594a );
 a97605a <=( (not A168)  and  A169 );
 a97608a <=( (not A166)  and  A167 );
 a97609a <=( a97608a  and  a97605a );
 a97612a <=( (not A200)  and  A199 );
 a97615a <=( A202  and  A201 );
 a97616a <=( a97615a  and  a97612a );
 a97617a <=( a97616a  and  a97609a );
 a97620a <=( A233  and  A232 );
 a97623a <=( (not A268)  and  A265 );
 a97624a <=( a97623a  and  a97620a );
 a97627a <=( (not A299)  and  (not A269) );
 a97630a <=( (not A302)  and  (not A301) );
 a97631a <=( a97630a  and  a97627a );
 a97632a <=( a97631a  and  a97624a );
 a97635a <=( (not A168)  and  A169 );
 a97638a <=( (not A166)  and  A167 );
 a97639a <=( a97638a  and  a97635a );
 a97642a <=( (not A200)  and  A199 );
 a97645a <=( A202  and  A201 );
 a97646a <=( a97645a  and  a97642a );
 a97647a <=( a97646a  and  a97639a );
 a97650a <=( (not A235)  and  (not A233) );
 a97653a <=( A265  and  (not A236) );
 a97654a <=( a97653a  and  a97650a );
 a97657a <=( A298  and  A266 );
 a97660a <=( (not A302)  and  (not A301) );
 a97661a <=( a97660a  and  a97657a );
 a97662a <=( a97661a  and  a97654a );
 a97665a <=( (not A168)  and  A169 );
 a97668a <=( (not A166)  and  A167 );
 a97669a <=( a97668a  and  a97665a );
 a97672a <=( (not A200)  and  A199 );
 a97675a <=( A202  and  A201 );
 a97676a <=( a97675a  and  a97672a );
 a97677a <=( a97676a  and  a97669a );
 a97680a <=( (not A235)  and  (not A233) );
 a97683a <=( (not A266)  and  (not A236) );
 a97684a <=( a97683a  and  a97680a );
 a97687a <=( (not A269)  and  (not A268) );
 a97690a <=( (not A300)  and  A298 );
 a97691a <=( a97690a  and  a97687a );
 a97692a <=( a97691a  and  a97684a );
 a97695a <=( (not A168)  and  A169 );
 a97698a <=( (not A166)  and  A167 );
 a97699a <=( a97698a  and  a97695a );
 a97702a <=( (not A200)  and  A199 );
 a97705a <=( A202  and  A201 );
 a97706a <=( a97705a  and  a97702a );
 a97707a <=( a97706a  and  a97699a );
 a97710a <=( (not A235)  and  (not A233) );
 a97713a <=( (not A266)  and  (not A236) );
 a97714a <=( a97713a  and  a97710a );
 a97717a <=( (not A269)  and  (not A268) );
 a97720a <=( A299  and  A298 );
 a97721a <=( a97720a  and  a97717a );
 a97722a <=( a97721a  and  a97714a );
 a97725a <=( (not A168)  and  A169 );
 a97728a <=( (not A166)  and  A167 );
 a97729a <=( a97728a  and  a97725a );
 a97732a <=( (not A200)  and  A199 );
 a97735a <=( A202  and  A201 );
 a97736a <=( a97735a  and  a97732a );
 a97737a <=( a97736a  and  a97729a );
 a97740a <=( (not A235)  and  (not A233) );
 a97743a <=( (not A266)  and  (not A236) );
 a97744a <=( a97743a  and  a97740a );
 a97747a <=( (not A269)  and  (not A268) );
 a97750a <=( (not A299)  and  (not A298) );
 a97751a <=( a97750a  and  a97747a );
 a97752a <=( a97751a  and  a97744a );
 a97755a <=( (not A168)  and  A169 );
 a97758a <=( (not A166)  and  A167 );
 a97759a <=( a97758a  and  a97755a );
 a97762a <=( (not A200)  and  A199 );
 a97765a <=( A202  and  A201 );
 a97766a <=( a97765a  and  a97762a );
 a97767a <=( a97766a  and  a97759a );
 a97770a <=( (not A235)  and  (not A233) );
 a97773a <=( (not A266)  and  (not A236) );
 a97774a <=( a97773a  and  a97770a );
 a97777a <=( A298  and  (not A267) );
 a97780a <=( (not A302)  and  (not A301) );
 a97781a <=( a97780a  and  a97777a );
 a97782a <=( a97781a  and  a97774a );
 a97785a <=( (not A168)  and  A169 );
 a97788a <=( (not A166)  and  A167 );
 a97789a <=( a97788a  and  a97785a );
 a97792a <=( (not A200)  and  A199 );
 a97795a <=( A202  and  A201 );
 a97796a <=( a97795a  and  a97792a );
 a97797a <=( a97796a  and  a97789a );
 a97800a <=( (not A235)  and  (not A233) );
 a97803a <=( (not A265)  and  (not A236) );
 a97804a <=( a97803a  and  a97800a );
 a97807a <=( A298  and  (not A266) );
 a97810a <=( (not A302)  and  (not A301) );
 a97811a <=( a97810a  and  a97807a );
 a97812a <=( a97811a  and  a97804a );
 a97815a <=( (not A168)  and  A169 );
 a97818a <=( (not A166)  and  A167 );
 a97819a <=( a97818a  and  a97815a );
 a97822a <=( (not A200)  and  A199 );
 a97825a <=( A202  and  A201 );
 a97826a <=( a97825a  and  a97822a );
 a97827a <=( a97826a  and  a97819a );
 a97830a <=( (not A234)  and  (not A233) );
 a97833a <=( (not A268)  and  (not A266) );
 a97834a <=( a97833a  and  a97830a );
 a97837a <=( A298  and  (not A269) );
 a97840a <=( (not A302)  and  (not A301) );
 a97841a <=( a97840a  and  a97837a );
 a97842a <=( a97841a  and  a97834a );
 a97845a <=( (not A168)  and  A169 );
 a97848a <=( (not A166)  and  A167 );
 a97849a <=( a97848a  and  a97845a );
 a97852a <=( (not A200)  and  A199 );
 a97855a <=( A202  and  A201 );
 a97856a <=( a97855a  and  a97852a );
 a97857a <=( a97856a  and  a97849a );
 a97860a <=( (not A233)  and  A232 );
 a97863a <=( A235  and  A234 );
 a97864a <=( a97863a  and  a97860a );
 a97867a <=( (not A299)  and  A298 );
 a97870a <=( A301  and  A300 );
 a97871a <=( a97870a  and  a97867a );
 a97872a <=( a97871a  and  a97864a );
 a97875a <=( (not A168)  and  A169 );
 a97878a <=( (not A166)  and  A167 );
 a97879a <=( a97878a  and  a97875a );
 a97882a <=( (not A200)  and  A199 );
 a97885a <=( A202  and  A201 );
 a97886a <=( a97885a  and  a97882a );
 a97887a <=( a97886a  and  a97879a );
 a97890a <=( (not A233)  and  A232 );
 a97893a <=( A235  and  A234 );
 a97894a <=( a97893a  and  a97890a );
 a97897a <=( (not A299)  and  A298 );
 a97900a <=( A302  and  A300 );
 a97901a <=( a97900a  and  a97897a );
 a97902a <=( a97901a  and  a97894a );
 a97905a <=( (not A168)  and  A169 );
 a97908a <=( (not A166)  and  A167 );
 a97909a <=( a97908a  and  a97905a );
 a97912a <=( (not A200)  and  A199 );
 a97915a <=( A202  and  A201 );
 a97916a <=( a97915a  and  a97912a );
 a97917a <=( a97916a  and  a97909a );
 a97920a <=( (not A233)  and  A232 );
 a97923a <=( A235  and  A234 );
 a97924a <=( a97923a  and  a97920a );
 a97927a <=( (not A266)  and  A265 );
 a97930a <=( A268  and  A267 );
 a97931a <=( a97930a  and  a97927a );
 a97932a <=( a97931a  and  a97924a );
 a97935a <=( (not A168)  and  A169 );
 a97938a <=( (not A166)  and  A167 );
 a97939a <=( a97938a  and  a97935a );
 a97942a <=( (not A200)  and  A199 );
 a97945a <=( A202  and  A201 );
 a97946a <=( a97945a  and  a97942a );
 a97947a <=( a97946a  and  a97939a );
 a97950a <=( (not A233)  and  A232 );
 a97953a <=( A235  and  A234 );
 a97954a <=( a97953a  and  a97950a );
 a97957a <=( (not A266)  and  A265 );
 a97960a <=( A269  and  A267 );
 a97961a <=( a97960a  and  a97957a );
 a97962a <=( a97961a  and  a97954a );
 a97965a <=( (not A168)  and  A169 );
 a97968a <=( (not A166)  and  A167 );
 a97969a <=( a97968a  and  a97965a );
 a97972a <=( (not A200)  and  A199 );
 a97975a <=( A202  and  A201 );
 a97976a <=( a97975a  and  a97972a );
 a97977a <=( a97976a  and  a97969a );
 a97980a <=( (not A233)  and  A232 );
 a97983a <=( A236  and  A234 );
 a97984a <=( a97983a  and  a97980a );
 a97987a <=( (not A299)  and  A298 );
 a97990a <=( A301  and  A300 );
 a97991a <=( a97990a  and  a97987a );
 a97992a <=( a97991a  and  a97984a );
 a97995a <=( (not A168)  and  A169 );
 a97998a <=( (not A166)  and  A167 );
 a97999a <=( a97998a  and  a97995a );
 a98002a <=( (not A200)  and  A199 );
 a98005a <=( A202  and  A201 );
 a98006a <=( a98005a  and  a98002a );
 a98007a <=( a98006a  and  a97999a );
 a98010a <=( (not A233)  and  A232 );
 a98013a <=( A236  and  A234 );
 a98014a <=( a98013a  and  a98010a );
 a98017a <=( (not A299)  and  A298 );
 a98020a <=( A302  and  A300 );
 a98021a <=( a98020a  and  a98017a );
 a98022a <=( a98021a  and  a98014a );
 a98025a <=( (not A168)  and  A169 );
 a98028a <=( (not A166)  and  A167 );
 a98029a <=( a98028a  and  a98025a );
 a98032a <=( (not A200)  and  A199 );
 a98035a <=( A202  and  A201 );
 a98036a <=( a98035a  and  a98032a );
 a98037a <=( a98036a  and  a98029a );
 a98040a <=( (not A233)  and  A232 );
 a98043a <=( A236  and  A234 );
 a98044a <=( a98043a  and  a98040a );
 a98047a <=( (not A266)  and  A265 );
 a98050a <=( A268  and  A267 );
 a98051a <=( a98050a  and  a98047a );
 a98052a <=( a98051a  and  a98044a );
 a98055a <=( (not A168)  and  A169 );
 a98058a <=( (not A166)  and  A167 );
 a98059a <=( a98058a  and  a98055a );
 a98062a <=( (not A200)  and  A199 );
 a98065a <=( A202  and  A201 );
 a98066a <=( a98065a  and  a98062a );
 a98067a <=( a98066a  and  a98059a );
 a98070a <=( (not A233)  and  A232 );
 a98073a <=( A236  and  A234 );
 a98074a <=( a98073a  and  a98070a );
 a98077a <=( (not A266)  and  A265 );
 a98080a <=( A269  and  A267 );
 a98081a <=( a98080a  and  a98077a );
 a98082a <=( a98081a  and  a98074a );
 a98085a <=( (not A168)  and  A169 );
 a98088a <=( (not A166)  and  A167 );
 a98089a <=( a98088a  and  a98085a );
 a98092a <=( (not A200)  and  A199 );
 a98095a <=( A202  and  A201 );
 a98096a <=( a98095a  and  a98092a );
 a98097a <=( a98096a  and  a98089a );
 a98100a <=( (not A233)  and  (not A232) );
 a98103a <=( (not A268)  and  (not A266) );
 a98104a <=( a98103a  and  a98100a );
 a98107a <=( A298  and  (not A269) );
 a98110a <=( (not A302)  and  (not A301) );
 a98111a <=( a98110a  and  a98107a );
 a98112a <=( a98111a  and  a98104a );
 a98115a <=( (not A168)  and  A169 );
 a98118a <=( (not A166)  and  A167 );
 a98119a <=( a98118a  and  a98115a );
 a98122a <=( (not A200)  and  A199 );
 a98125a <=( A203  and  A201 );
 a98126a <=( a98125a  and  a98122a );
 a98127a <=( a98126a  and  a98119a );
 a98130a <=( A233  and  A232 );
 a98133a <=( (not A268)  and  A265 );
 a98134a <=( a98133a  and  a98130a );
 a98137a <=( (not A299)  and  (not A269) );
 a98140a <=( (not A302)  and  (not A301) );
 a98141a <=( a98140a  and  a98137a );
 a98142a <=( a98141a  and  a98134a );
 a98145a <=( (not A168)  and  A169 );
 a98148a <=( (not A166)  and  A167 );
 a98149a <=( a98148a  and  a98145a );
 a98152a <=( (not A200)  and  A199 );
 a98155a <=( A203  and  A201 );
 a98156a <=( a98155a  and  a98152a );
 a98157a <=( a98156a  and  a98149a );
 a98160a <=( (not A235)  and  (not A233) );
 a98163a <=( A265  and  (not A236) );
 a98164a <=( a98163a  and  a98160a );
 a98167a <=( A298  and  A266 );
 a98170a <=( (not A302)  and  (not A301) );
 a98171a <=( a98170a  and  a98167a );
 a98172a <=( a98171a  and  a98164a );
 a98175a <=( (not A168)  and  A169 );
 a98178a <=( (not A166)  and  A167 );
 a98179a <=( a98178a  and  a98175a );
 a98182a <=( (not A200)  and  A199 );
 a98185a <=( A203  and  A201 );
 a98186a <=( a98185a  and  a98182a );
 a98187a <=( a98186a  and  a98179a );
 a98190a <=( (not A235)  and  (not A233) );
 a98193a <=( (not A266)  and  (not A236) );
 a98194a <=( a98193a  and  a98190a );
 a98197a <=( (not A269)  and  (not A268) );
 a98200a <=( (not A300)  and  A298 );
 a98201a <=( a98200a  and  a98197a );
 a98202a <=( a98201a  and  a98194a );
 a98205a <=( (not A168)  and  A169 );
 a98208a <=( (not A166)  and  A167 );
 a98209a <=( a98208a  and  a98205a );
 a98212a <=( (not A200)  and  A199 );
 a98215a <=( A203  and  A201 );
 a98216a <=( a98215a  and  a98212a );
 a98217a <=( a98216a  and  a98209a );
 a98220a <=( (not A235)  and  (not A233) );
 a98223a <=( (not A266)  and  (not A236) );
 a98224a <=( a98223a  and  a98220a );
 a98227a <=( (not A269)  and  (not A268) );
 a98230a <=( A299  and  A298 );
 a98231a <=( a98230a  and  a98227a );
 a98232a <=( a98231a  and  a98224a );
 a98235a <=( (not A168)  and  A169 );
 a98238a <=( (not A166)  and  A167 );
 a98239a <=( a98238a  and  a98235a );
 a98242a <=( (not A200)  and  A199 );
 a98245a <=( A203  and  A201 );
 a98246a <=( a98245a  and  a98242a );
 a98247a <=( a98246a  and  a98239a );
 a98250a <=( (not A235)  and  (not A233) );
 a98253a <=( (not A266)  and  (not A236) );
 a98254a <=( a98253a  and  a98250a );
 a98257a <=( (not A269)  and  (not A268) );
 a98260a <=( (not A299)  and  (not A298) );
 a98261a <=( a98260a  and  a98257a );
 a98262a <=( a98261a  and  a98254a );
 a98265a <=( (not A168)  and  A169 );
 a98268a <=( (not A166)  and  A167 );
 a98269a <=( a98268a  and  a98265a );
 a98272a <=( (not A200)  and  A199 );
 a98275a <=( A203  and  A201 );
 a98276a <=( a98275a  and  a98272a );
 a98277a <=( a98276a  and  a98269a );
 a98280a <=( (not A235)  and  (not A233) );
 a98283a <=( (not A266)  and  (not A236) );
 a98284a <=( a98283a  and  a98280a );
 a98287a <=( A298  and  (not A267) );
 a98290a <=( (not A302)  and  (not A301) );
 a98291a <=( a98290a  and  a98287a );
 a98292a <=( a98291a  and  a98284a );
 a98295a <=( (not A168)  and  A169 );
 a98298a <=( (not A166)  and  A167 );
 a98299a <=( a98298a  and  a98295a );
 a98302a <=( (not A200)  and  A199 );
 a98305a <=( A203  and  A201 );
 a98306a <=( a98305a  and  a98302a );
 a98307a <=( a98306a  and  a98299a );
 a98310a <=( (not A235)  and  (not A233) );
 a98313a <=( (not A265)  and  (not A236) );
 a98314a <=( a98313a  and  a98310a );
 a98317a <=( A298  and  (not A266) );
 a98320a <=( (not A302)  and  (not A301) );
 a98321a <=( a98320a  and  a98317a );
 a98322a <=( a98321a  and  a98314a );
 a98325a <=( (not A168)  and  A169 );
 a98328a <=( (not A166)  and  A167 );
 a98329a <=( a98328a  and  a98325a );
 a98332a <=( (not A200)  and  A199 );
 a98335a <=( A203  and  A201 );
 a98336a <=( a98335a  and  a98332a );
 a98337a <=( a98336a  and  a98329a );
 a98340a <=( (not A234)  and  (not A233) );
 a98343a <=( (not A268)  and  (not A266) );
 a98344a <=( a98343a  and  a98340a );
 a98347a <=( A298  and  (not A269) );
 a98350a <=( (not A302)  and  (not A301) );
 a98351a <=( a98350a  and  a98347a );
 a98352a <=( a98351a  and  a98344a );
 a98355a <=( (not A168)  and  A169 );
 a98358a <=( (not A166)  and  A167 );
 a98359a <=( a98358a  and  a98355a );
 a98362a <=( (not A200)  and  A199 );
 a98365a <=( A203  and  A201 );
 a98366a <=( a98365a  and  a98362a );
 a98367a <=( a98366a  and  a98359a );
 a98370a <=( (not A233)  and  A232 );
 a98373a <=( A235  and  A234 );
 a98374a <=( a98373a  and  a98370a );
 a98377a <=( (not A299)  and  A298 );
 a98380a <=( A301  and  A300 );
 a98381a <=( a98380a  and  a98377a );
 a98382a <=( a98381a  and  a98374a );
 a98385a <=( (not A168)  and  A169 );
 a98388a <=( (not A166)  and  A167 );
 a98389a <=( a98388a  and  a98385a );
 a98392a <=( (not A200)  and  A199 );
 a98395a <=( A203  and  A201 );
 a98396a <=( a98395a  and  a98392a );
 a98397a <=( a98396a  and  a98389a );
 a98400a <=( (not A233)  and  A232 );
 a98403a <=( A235  and  A234 );
 a98404a <=( a98403a  and  a98400a );
 a98407a <=( (not A299)  and  A298 );
 a98410a <=( A302  and  A300 );
 a98411a <=( a98410a  and  a98407a );
 a98412a <=( a98411a  and  a98404a );
 a98415a <=( (not A168)  and  A169 );
 a98418a <=( (not A166)  and  A167 );
 a98419a <=( a98418a  and  a98415a );
 a98422a <=( (not A200)  and  A199 );
 a98425a <=( A203  and  A201 );
 a98426a <=( a98425a  and  a98422a );
 a98427a <=( a98426a  and  a98419a );
 a98430a <=( (not A233)  and  A232 );
 a98433a <=( A235  and  A234 );
 a98434a <=( a98433a  and  a98430a );
 a98437a <=( (not A266)  and  A265 );
 a98440a <=( A268  and  A267 );
 a98441a <=( a98440a  and  a98437a );
 a98442a <=( a98441a  and  a98434a );
 a98445a <=( (not A168)  and  A169 );
 a98448a <=( (not A166)  and  A167 );
 a98449a <=( a98448a  and  a98445a );
 a98452a <=( (not A200)  and  A199 );
 a98455a <=( A203  and  A201 );
 a98456a <=( a98455a  and  a98452a );
 a98457a <=( a98456a  and  a98449a );
 a98460a <=( (not A233)  and  A232 );
 a98463a <=( A235  and  A234 );
 a98464a <=( a98463a  and  a98460a );
 a98467a <=( (not A266)  and  A265 );
 a98470a <=( A269  and  A267 );
 a98471a <=( a98470a  and  a98467a );
 a98472a <=( a98471a  and  a98464a );
 a98475a <=( (not A168)  and  A169 );
 a98478a <=( (not A166)  and  A167 );
 a98479a <=( a98478a  and  a98475a );
 a98482a <=( (not A200)  and  A199 );
 a98485a <=( A203  and  A201 );
 a98486a <=( a98485a  and  a98482a );
 a98487a <=( a98486a  and  a98479a );
 a98490a <=( (not A233)  and  A232 );
 a98493a <=( A236  and  A234 );
 a98494a <=( a98493a  and  a98490a );
 a98497a <=( (not A299)  and  A298 );
 a98500a <=( A301  and  A300 );
 a98501a <=( a98500a  and  a98497a );
 a98502a <=( a98501a  and  a98494a );
 a98505a <=( (not A168)  and  A169 );
 a98508a <=( (not A166)  and  A167 );
 a98509a <=( a98508a  and  a98505a );
 a98512a <=( (not A200)  and  A199 );
 a98515a <=( A203  and  A201 );
 a98516a <=( a98515a  and  a98512a );
 a98517a <=( a98516a  and  a98509a );
 a98520a <=( (not A233)  and  A232 );
 a98523a <=( A236  and  A234 );
 a98524a <=( a98523a  and  a98520a );
 a98527a <=( (not A299)  and  A298 );
 a98530a <=( A302  and  A300 );
 a98531a <=( a98530a  and  a98527a );
 a98532a <=( a98531a  and  a98524a );
 a98535a <=( (not A168)  and  A169 );
 a98538a <=( (not A166)  and  A167 );
 a98539a <=( a98538a  and  a98535a );
 a98542a <=( (not A200)  and  A199 );
 a98545a <=( A203  and  A201 );
 a98546a <=( a98545a  and  a98542a );
 a98547a <=( a98546a  and  a98539a );
 a98550a <=( (not A233)  and  A232 );
 a98553a <=( A236  and  A234 );
 a98554a <=( a98553a  and  a98550a );
 a98557a <=( (not A266)  and  A265 );
 a98560a <=( A268  and  A267 );
 a98561a <=( a98560a  and  a98557a );
 a98562a <=( a98561a  and  a98554a );
 a98565a <=( (not A168)  and  A169 );
 a98568a <=( (not A166)  and  A167 );
 a98569a <=( a98568a  and  a98565a );
 a98572a <=( (not A200)  and  A199 );
 a98575a <=( A203  and  A201 );
 a98576a <=( a98575a  and  a98572a );
 a98577a <=( a98576a  and  a98569a );
 a98580a <=( (not A233)  and  A232 );
 a98583a <=( A236  and  A234 );
 a98584a <=( a98583a  and  a98580a );
 a98587a <=( (not A266)  and  A265 );
 a98590a <=( A269  and  A267 );
 a98591a <=( a98590a  and  a98587a );
 a98592a <=( a98591a  and  a98584a );
 a98595a <=( (not A168)  and  A169 );
 a98598a <=( (not A166)  and  A167 );
 a98599a <=( a98598a  and  a98595a );
 a98602a <=( (not A200)  and  A199 );
 a98605a <=( A203  and  A201 );
 a98606a <=( a98605a  and  a98602a );
 a98607a <=( a98606a  and  a98599a );
 a98610a <=( (not A233)  and  (not A232) );
 a98613a <=( (not A268)  and  (not A266) );
 a98614a <=( a98613a  and  a98610a );
 a98617a <=( A298  and  (not A269) );
 a98620a <=( (not A302)  and  (not A301) );
 a98621a <=( a98620a  and  a98617a );
 a98622a <=( a98621a  and  a98614a );
 a98625a <=( (not A168)  and  A169 );
 a98628a <=( A166  and  (not A167) );
 a98629a <=( a98628a  and  a98625a );
 a98632a <=( (not A200)  and  A199 );
 a98635a <=( A202  and  A201 );
 a98636a <=( a98635a  and  a98632a );
 a98637a <=( a98636a  and  a98629a );
 a98640a <=( A233  and  A232 );
 a98643a <=( (not A268)  and  A265 );
 a98644a <=( a98643a  and  a98640a );
 a98647a <=( (not A299)  and  (not A269) );
 a98650a <=( (not A302)  and  (not A301) );
 a98651a <=( a98650a  and  a98647a );
 a98652a <=( a98651a  and  a98644a );
 a98655a <=( (not A168)  and  A169 );
 a98658a <=( A166  and  (not A167) );
 a98659a <=( a98658a  and  a98655a );
 a98662a <=( (not A200)  and  A199 );
 a98665a <=( A202  and  A201 );
 a98666a <=( a98665a  and  a98662a );
 a98667a <=( a98666a  and  a98659a );
 a98670a <=( (not A235)  and  (not A233) );
 a98673a <=( A265  and  (not A236) );
 a98674a <=( a98673a  and  a98670a );
 a98677a <=( A298  and  A266 );
 a98680a <=( (not A302)  and  (not A301) );
 a98681a <=( a98680a  and  a98677a );
 a98682a <=( a98681a  and  a98674a );
 a98685a <=( (not A168)  and  A169 );
 a98688a <=( A166  and  (not A167) );
 a98689a <=( a98688a  and  a98685a );
 a98692a <=( (not A200)  and  A199 );
 a98695a <=( A202  and  A201 );
 a98696a <=( a98695a  and  a98692a );
 a98697a <=( a98696a  and  a98689a );
 a98700a <=( (not A235)  and  (not A233) );
 a98703a <=( (not A266)  and  (not A236) );
 a98704a <=( a98703a  and  a98700a );
 a98707a <=( (not A269)  and  (not A268) );
 a98710a <=( (not A300)  and  A298 );
 a98711a <=( a98710a  and  a98707a );
 a98712a <=( a98711a  and  a98704a );
 a98715a <=( (not A168)  and  A169 );
 a98718a <=( A166  and  (not A167) );
 a98719a <=( a98718a  and  a98715a );
 a98722a <=( (not A200)  and  A199 );
 a98725a <=( A202  and  A201 );
 a98726a <=( a98725a  and  a98722a );
 a98727a <=( a98726a  and  a98719a );
 a98730a <=( (not A235)  and  (not A233) );
 a98733a <=( (not A266)  and  (not A236) );
 a98734a <=( a98733a  and  a98730a );
 a98737a <=( (not A269)  and  (not A268) );
 a98740a <=( A299  and  A298 );
 a98741a <=( a98740a  and  a98737a );
 a98742a <=( a98741a  and  a98734a );
 a98745a <=( (not A168)  and  A169 );
 a98748a <=( A166  and  (not A167) );
 a98749a <=( a98748a  and  a98745a );
 a98752a <=( (not A200)  and  A199 );
 a98755a <=( A202  and  A201 );
 a98756a <=( a98755a  and  a98752a );
 a98757a <=( a98756a  and  a98749a );
 a98760a <=( (not A235)  and  (not A233) );
 a98763a <=( (not A266)  and  (not A236) );
 a98764a <=( a98763a  and  a98760a );
 a98767a <=( (not A269)  and  (not A268) );
 a98770a <=( (not A299)  and  (not A298) );
 a98771a <=( a98770a  and  a98767a );
 a98772a <=( a98771a  and  a98764a );
 a98775a <=( (not A168)  and  A169 );
 a98778a <=( A166  and  (not A167) );
 a98779a <=( a98778a  and  a98775a );
 a98782a <=( (not A200)  and  A199 );
 a98785a <=( A202  and  A201 );
 a98786a <=( a98785a  and  a98782a );
 a98787a <=( a98786a  and  a98779a );
 a98790a <=( (not A235)  and  (not A233) );
 a98793a <=( (not A266)  and  (not A236) );
 a98794a <=( a98793a  and  a98790a );
 a98797a <=( A298  and  (not A267) );
 a98800a <=( (not A302)  and  (not A301) );
 a98801a <=( a98800a  and  a98797a );
 a98802a <=( a98801a  and  a98794a );
 a98805a <=( (not A168)  and  A169 );
 a98808a <=( A166  and  (not A167) );
 a98809a <=( a98808a  and  a98805a );
 a98812a <=( (not A200)  and  A199 );
 a98815a <=( A202  and  A201 );
 a98816a <=( a98815a  and  a98812a );
 a98817a <=( a98816a  and  a98809a );
 a98820a <=( (not A235)  and  (not A233) );
 a98823a <=( (not A265)  and  (not A236) );
 a98824a <=( a98823a  and  a98820a );
 a98827a <=( A298  and  (not A266) );
 a98830a <=( (not A302)  and  (not A301) );
 a98831a <=( a98830a  and  a98827a );
 a98832a <=( a98831a  and  a98824a );
 a98835a <=( (not A168)  and  A169 );
 a98838a <=( A166  and  (not A167) );
 a98839a <=( a98838a  and  a98835a );
 a98842a <=( (not A200)  and  A199 );
 a98845a <=( A202  and  A201 );
 a98846a <=( a98845a  and  a98842a );
 a98847a <=( a98846a  and  a98839a );
 a98850a <=( (not A234)  and  (not A233) );
 a98853a <=( (not A268)  and  (not A266) );
 a98854a <=( a98853a  and  a98850a );
 a98857a <=( A298  and  (not A269) );
 a98860a <=( (not A302)  and  (not A301) );
 a98861a <=( a98860a  and  a98857a );
 a98862a <=( a98861a  and  a98854a );
 a98865a <=( (not A168)  and  A169 );
 a98868a <=( A166  and  (not A167) );
 a98869a <=( a98868a  and  a98865a );
 a98872a <=( (not A200)  and  A199 );
 a98875a <=( A202  and  A201 );
 a98876a <=( a98875a  and  a98872a );
 a98877a <=( a98876a  and  a98869a );
 a98880a <=( (not A233)  and  A232 );
 a98883a <=( A235  and  A234 );
 a98884a <=( a98883a  and  a98880a );
 a98887a <=( (not A299)  and  A298 );
 a98890a <=( A301  and  A300 );
 a98891a <=( a98890a  and  a98887a );
 a98892a <=( a98891a  and  a98884a );
 a98895a <=( (not A168)  and  A169 );
 a98898a <=( A166  and  (not A167) );
 a98899a <=( a98898a  and  a98895a );
 a98902a <=( (not A200)  and  A199 );
 a98905a <=( A202  and  A201 );
 a98906a <=( a98905a  and  a98902a );
 a98907a <=( a98906a  and  a98899a );
 a98910a <=( (not A233)  and  A232 );
 a98913a <=( A235  and  A234 );
 a98914a <=( a98913a  and  a98910a );
 a98917a <=( (not A299)  and  A298 );
 a98920a <=( A302  and  A300 );
 a98921a <=( a98920a  and  a98917a );
 a98922a <=( a98921a  and  a98914a );
 a98925a <=( (not A168)  and  A169 );
 a98928a <=( A166  and  (not A167) );
 a98929a <=( a98928a  and  a98925a );
 a98932a <=( (not A200)  and  A199 );
 a98935a <=( A202  and  A201 );
 a98936a <=( a98935a  and  a98932a );
 a98937a <=( a98936a  and  a98929a );
 a98940a <=( (not A233)  and  A232 );
 a98943a <=( A235  and  A234 );
 a98944a <=( a98943a  and  a98940a );
 a98947a <=( (not A266)  and  A265 );
 a98950a <=( A268  and  A267 );
 a98951a <=( a98950a  and  a98947a );
 a98952a <=( a98951a  and  a98944a );
 a98955a <=( (not A168)  and  A169 );
 a98958a <=( A166  and  (not A167) );
 a98959a <=( a98958a  and  a98955a );
 a98962a <=( (not A200)  and  A199 );
 a98965a <=( A202  and  A201 );
 a98966a <=( a98965a  and  a98962a );
 a98967a <=( a98966a  and  a98959a );
 a98970a <=( (not A233)  and  A232 );
 a98973a <=( A235  and  A234 );
 a98974a <=( a98973a  and  a98970a );
 a98977a <=( (not A266)  and  A265 );
 a98980a <=( A269  and  A267 );
 a98981a <=( a98980a  and  a98977a );
 a98982a <=( a98981a  and  a98974a );
 a98985a <=( (not A168)  and  A169 );
 a98988a <=( A166  and  (not A167) );
 a98989a <=( a98988a  and  a98985a );
 a98992a <=( (not A200)  and  A199 );
 a98995a <=( A202  and  A201 );
 a98996a <=( a98995a  and  a98992a );
 a98997a <=( a98996a  and  a98989a );
 a99000a <=( (not A233)  and  A232 );
 a99003a <=( A236  and  A234 );
 a99004a <=( a99003a  and  a99000a );
 a99007a <=( (not A299)  and  A298 );
 a99010a <=( A301  and  A300 );
 a99011a <=( a99010a  and  a99007a );
 a99012a <=( a99011a  and  a99004a );
 a99015a <=( (not A168)  and  A169 );
 a99018a <=( A166  and  (not A167) );
 a99019a <=( a99018a  and  a99015a );
 a99022a <=( (not A200)  and  A199 );
 a99025a <=( A202  and  A201 );
 a99026a <=( a99025a  and  a99022a );
 a99027a <=( a99026a  and  a99019a );
 a99030a <=( (not A233)  and  A232 );
 a99033a <=( A236  and  A234 );
 a99034a <=( a99033a  and  a99030a );
 a99037a <=( (not A299)  and  A298 );
 a99040a <=( A302  and  A300 );
 a99041a <=( a99040a  and  a99037a );
 a99042a <=( a99041a  and  a99034a );
 a99045a <=( (not A168)  and  A169 );
 a99048a <=( A166  and  (not A167) );
 a99049a <=( a99048a  and  a99045a );
 a99052a <=( (not A200)  and  A199 );
 a99055a <=( A202  and  A201 );
 a99056a <=( a99055a  and  a99052a );
 a99057a <=( a99056a  and  a99049a );
 a99060a <=( (not A233)  and  A232 );
 a99063a <=( A236  and  A234 );
 a99064a <=( a99063a  and  a99060a );
 a99067a <=( (not A266)  and  A265 );
 a99070a <=( A268  and  A267 );
 a99071a <=( a99070a  and  a99067a );
 a99072a <=( a99071a  and  a99064a );
 a99075a <=( (not A168)  and  A169 );
 a99078a <=( A166  and  (not A167) );
 a99079a <=( a99078a  and  a99075a );
 a99082a <=( (not A200)  and  A199 );
 a99085a <=( A202  and  A201 );
 a99086a <=( a99085a  and  a99082a );
 a99087a <=( a99086a  and  a99079a );
 a99090a <=( (not A233)  and  A232 );
 a99093a <=( A236  and  A234 );
 a99094a <=( a99093a  and  a99090a );
 a99097a <=( (not A266)  and  A265 );
 a99100a <=( A269  and  A267 );
 a99101a <=( a99100a  and  a99097a );
 a99102a <=( a99101a  and  a99094a );
 a99105a <=( (not A168)  and  A169 );
 a99108a <=( A166  and  (not A167) );
 a99109a <=( a99108a  and  a99105a );
 a99112a <=( (not A200)  and  A199 );
 a99115a <=( A202  and  A201 );
 a99116a <=( a99115a  and  a99112a );
 a99117a <=( a99116a  and  a99109a );
 a99120a <=( (not A233)  and  (not A232) );
 a99123a <=( (not A268)  and  (not A266) );
 a99124a <=( a99123a  and  a99120a );
 a99127a <=( A298  and  (not A269) );
 a99130a <=( (not A302)  and  (not A301) );
 a99131a <=( a99130a  and  a99127a );
 a99132a <=( a99131a  and  a99124a );
 a99135a <=( (not A168)  and  A169 );
 a99138a <=( A166  and  (not A167) );
 a99139a <=( a99138a  and  a99135a );
 a99142a <=( (not A200)  and  A199 );
 a99145a <=( A203  and  A201 );
 a99146a <=( a99145a  and  a99142a );
 a99147a <=( a99146a  and  a99139a );
 a99150a <=( A233  and  A232 );
 a99153a <=( (not A268)  and  A265 );
 a99154a <=( a99153a  and  a99150a );
 a99157a <=( (not A299)  and  (not A269) );
 a99160a <=( (not A302)  and  (not A301) );
 a99161a <=( a99160a  and  a99157a );
 a99162a <=( a99161a  and  a99154a );
 a99165a <=( (not A168)  and  A169 );
 a99168a <=( A166  and  (not A167) );
 a99169a <=( a99168a  and  a99165a );
 a99172a <=( (not A200)  and  A199 );
 a99175a <=( A203  and  A201 );
 a99176a <=( a99175a  and  a99172a );
 a99177a <=( a99176a  and  a99169a );
 a99180a <=( (not A235)  and  (not A233) );
 a99183a <=( A265  and  (not A236) );
 a99184a <=( a99183a  and  a99180a );
 a99187a <=( A298  and  A266 );
 a99190a <=( (not A302)  and  (not A301) );
 a99191a <=( a99190a  and  a99187a );
 a99192a <=( a99191a  and  a99184a );
 a99195a <=( (not A168)  and  A169 );
 a99198a <=( A166  and  (not A167) );
 a99199a <=( a99198a  and  a99195a );
 a99202a <=( (not A200)  and  A199 );
 a99205a <=( A203  and  A201 );
 a99206a <=( a99205a  and  a99202a );
 a99207a <=( a99206a  and  a99199a );
 a99210a <=( (not A235)  and  (not A233) );
 a99213a <=( (not A266)  and  (not A236) );
 a99214a <=( a99213a  and  a99210a );
 a99217a <=( (not A269)  and  (not A268) );
 a99220a <=( (not A300)  and  A298 );
 a99221a <=( a99220a  and  a99217a );
 a99222a <=( a99221a  and  a99214a );
 a99225a <=( (not A168)  and  A169 );
 a99228a <=( A166  and  (not A167) );
 a99229a <=( a99228a  and  a99225a );
 a99232a <=( (not A200)  and  A199 );
 a99235a <=( A203  and  A201 );
 a99236a <=( a99235a  and  a99232a );
 a99237a <=( a99236a  and  a99229a );
 a99240a <=( (not A235)  and  (not A233) );
 a99243a <=( (not A266)  and  (not A236) );
 a99244a <=( a99243a  and  a99240a );
 a99247a <=( (not A269)  and  (not A268) );
 a99250a <=( A299  and  A298 );
 a99251a <=( a99250a  and  a99247a );
 a99252a <=( a99251a  and  a99244a );
 a99255a <=( (not A168)  and  A169 );
 a99258a <=( A166  and  (not A167) );
 a99259a <=( a99258a  and  a99255a );
 a99262a <=( (not A200)  and  A199 );
 a99265a <=( A203  and  A201 );
 a99266a <=( a99265a  and  a99262a );
 a99267a <=( a99266a  and  a99259a );
 a99270a <=( (not A235)  and  (not A233) );
 a99273a <=( (not A266)  and  (not A236) );
 a99274a <=( a99273a  and  a99270a );
 a99277a <=( (not A269)  and  (not A268) );
 a99280a <=( (not A299)  and  (not A298) );
 a99281a <=( a99280a  and  a99277a );
 a99282a <=( a99281a  and  a99274a );
 a99285a <=( (not A168)  and  A169 );
 a99288a <=( A166  and  (not A167) );
 a99289a <=( a99288a  and  a99285a );
 a99292a <=( (not A200)  and  A199 );
 a99295a <=( A203  and  A201 );
 a99296a <=( a99295a  and  a99292a );
 a99297a <=( a99296a  and  a99289a );
 a99300a <=( (not A235)  and  (not A233) );
 a99303a <=( (not A266)  and  (not A236) );
 a99304a <=( a99303a  and  a99300a );
 a99307a <=( A298  and  (not A267) );
 a99310a <=( (not A302)  and  (not A301) );
 a99311a <=( a99310a  and  a99307a );
 a99312a <=( a99311a  and  a99304a );
 a99315a <=( (not A168)  and  A169 );
 a99318a <=( A166  and  (not A167) );
 a99319a <=( a99318a  and  a99315a );
 a99322a <=( (not A200)  and  A199 );
 a99325a <=( A203  and  A201 );
 a99326a <=( a99325a  and  a99322a );
 a99327a <=( a99326a  and  a99319a );
 a99330a <=( (not A235)  and  (not A233) );
 a99333a <=( (not A265)  and  (not A236) );
 a99334a <=( a99333a  and  a99330a );
 a99337a <=( A298  and  (not A266) );
 a99340a <=( (not A302)  and  (not A301) );
 a99341a <=( a99340a  and  a99337a );
 a99342a <=( a99341a  and  a99334a );
 a99345a <=( (not A168)  and  A169 );
 a99348a <=( A166  and  (not A167) );
 a99349a <=( a99348a  and  a99345a );
 a99352a <=( (not A200)  and  A199 );
 a99355a <=( A203  and  A201 );
 a99356a <=( a99355a  and  a99352a );
 a99357a <=( a99356a  and  a99349a );
 a99360a <=( (not A234)  and  (not A233) );
 a99363a <=( (not A268)  and  (not A266) );
 a99364a <=( a99363a  and  a99360a );
 a99367a <=( A298  and  (not A269) );
 a99370a <=( (not A302)  and  (not A301) );
 a99371a <=( a99370a  and  a99367a );
 a99372a <=( a99371a  and  a99364a );
 a99375a <=( (not A168)  and  A169 );
 a99378a <=( A166  and  (not A167) );
 a99379a <=( a99378a  and  a99375a );
 a99382a <=( (not A200)  and  A199 );
 a99385a <=( A203  and  A201 );
 a99386a <=( a99385a  and  a99382a );
 a99387a <=( a99386a  and  a99379a );
 a99390a <=( (not A233)  and  A232 );
 a99393a <=( A235  and  A234 );
 a99394a <=( a99393a  and  a99390a );
 a99397a <=( (not A299)  and  A298 );
 a99400a <=( A301  and  A300 );
 a99401a <=( a99400a  and  a99397a );
 a99402a <=( a99401a  and  a99394a );
 a99405a <=( (not A168)  and  A169 );
 a99408a <=( A166  and  (not A167) );
 a99409a <=( a99408a  and  a99405a );
 a99412a <=( (not A200)  and  A199 );
 a99415a <=( A203  and  A201 );
 a99416a <=( a99415a  and  a99412a );
 a99417a <=( a99416a  and  a99409a );
 a99420a <=( (not A233)  and  A232 );
 a99423a <=( A235  and  A234 );
 a99424a <=( a99423a  and  a99420a );
 a99427a <=( (not A299)  and  A298 );
 a99430a <=( A302  and  A300 );
 a99431a <=( a99430a  and  a99427a );
 a99432a <=( a99431a  and  a99424a );
 a99435a <=( (not A168)  and  A169 );
 a99438a <=( A166  and  (not A167) );
 a99439a <=( a99438a  and  a99435a );
 a99442a <=( (not A200)  and  A199 );
 a99445a <=( A203  and  A201 );
 a99446a <=( a99445a  and  a99442a );
 a99447a <=( a99446a  and  a99439a );
 a99450a <=( (not A233)  and  A232 );
 a99453a <=( A235  and  A234 );
 a99454a <=( a99453a  and  a99450a );
 a99457a <=( (not A266)  and  A265 );
 a99460a <=( A268  and  A267 );
 a99461a <=( a99460a  and  a99457a );
 a99462a <=( a99461a  and  a99454a );
 a99465a <=( (not A168)  and  A169 );
 a99468a <=( A166  and  (not A167) );
 a99469a <=( a99468a  and  a99465a );
 a99472a <=( (not A200)  and  A199 );
 a99475a <=( A203  and  A201 );
 a99476a <=( a99475a  and  a99472a );
 a99477a <=( a99476a  and  a99469a );
 a99480a <=( (not A233)  and  A232 );
 a99483a <=( A235  and  A234 );
 a99484a <=( a99483a  and  a99480a );
 a99487a <=( (not A266)  and  A265 );
 a99490a <=( A269  and  A267 );
 a99491a <=( a99490a  and  a99487a );
 a99492a <=( a99491a  and  a99484a );
 a99495a <=( (not A168)  and  A169 );
 a99498a <=( A166  and  (not A167) );
 a99499a <=( a99498a  and  a99495a );
 a99502a <=( (not A200)  and  A199 );
 a99505a <=( A203  and  A201 );
 a99506a <=( a99505a  and  a99502a );
 a99507a <=( a99506a  and  a99499a );
 a99510a <=( (not A233)  and  A232 );
 a99513a <=( A236  and  A234 );
 a99514a <=( a99513a  and  a99510a );
 a99517a <=( (not A299)  and  A298 );
 a99520a <=( A301  and  A300 );
 a99521a <=( a99520a  and  a99517a );
 a99522a <=( a99521a  and  a99514a );
 a99525a <=( (not A168)  and  A169 );
 a99528a <=( A166  and  (not A167) );
 a99529a <=( a99528a  and  a99525a );
 a99532a <=( (not A200)  and  A199 );
 a99535a <=( A203  and  A201 );
 a99536a <=( a99535a  and  a99532a );
 a99537a <=( a99536a  and  a99529a );
 a99540a <=( (not A233)  and  A232 );
 a99543a <=( A236  and  A234 );
 a99544a <=( a99543a  and  a99540a );
 a99547a <=( (not A299)  and  A298 );
 a99550a <=( A302  and  A300 );
 a99551a <=( a99550a  and  a99547a );
 a99552a <=( a99551a  and  a99544a );
 a99555a <=( (not A168)  and  A169 );
 a99558a <=( A166  and  (not A167) );
 a99559a <=( a99558a  and  a99555a );
 a99562a <=( (not A200)  and  A199 );
 a99565a <=( A203  and  A201 );
 a99566a <=( a99565a  and  a99562a );
 a99567a <=( a99566a  and  a99559a );
 a99570a <=( (not A233)  and  A232 );
 a99573a <=( A236  and  A234 );
 a99574a <=( a99573a  and  a99570a );
 a99577a <=( (not A266)  and  A265 );
 a99580a <=( A268  and  A267 );
 a99581a <=( a99580a  and  a99577a );
 a99582a <=( a99581a  and  a99574a );
 a99585a <=( (not A168)  and  A169 );
 a99588a <=( A166  and  (not A167) );
 a99589a <=( a99588a  and  a99585a );
 a99592a <=( (not A200)  and  A199 );
 a99595a <=( A203  and  A201 );
 a99596a <=( a99595a  and  a99592a );
 a99597a <=( a99596a  and  a99589a );
 a99600a <=( (not A233)  and  A232 );
 a99603a <=( A236  and  A234 );
 a99604a <=( a99603a  and  a99600a );
 a99607a <=( (not A266)  and  A265 );
 a99610a <=( A269  and  A267 );
 a99611a <=( a99610a  and  a99607a );
 a99612a <=( a99611a  and  a99604a );
 a99615a <=( (not A168)  and  A169 );
 a99618a <=( A166  and  (not A167) );
 a99619a <=( a99618a  and  a99615a );
 a99622a <=( (not A200)  and  A199 );
 a99625a <=( A203  and  A201 );
 a99626a <=( a99625a  and  a99622a );
 a99627a <=( a99626a  and  a99619a );
 a99630a <=( (not A233)  and  (not A232) );
 a99633a <=( (not A268)  and  (not A266) );
 a99634a <=( a99633a  and  a99630a );
 a99637a <=( A298  and  (not A269) );
 a99640a <=( (not A302)  and  (not A301) );
 a99641a <=( a99640a  and  a99637a );
 a99642a <=( a99641a  and  a99634a );
 a99645a <=( A169  and  A170 );
 a99648a <=( A199  and  (not A168) );
 a99649a <=( a99648a  and  a99645a );
 a99652a <=( A201  and  (not A200) );
 a99655a <=( (not A233)  and  A202 );
 a99656a <=( a99655a  and  a99652a );
 a99657a <=( a99656a  and  a99649a );
 a99660a <=( (not A236)  and  (not A235) );
 a99663a <=( (not A268)  and  (not A266) );
 a99664a <=( a99663a  and  a99660a );
 a99667a <=( A298  and  (not A269) );
 a99670a <=( (not A302)  and  (not A301) );
 a99671a <=( a99670a  and  a99667a );
 a99672a <=( a99671a  and  a99664a );
 a99675a <=( A169  and  A170 );
 a99678a <=( A199  and  (not A168) );
 a99679a <=( a99678a  and  a99675a );
 a99682a <=( A201  and  (not A200) );
 a99685a <=( (not A233)  and  A203 );
 a99686a <=( a99685a  and  a99682a );
 a99687a <=( a99686a  and  a99679a );
 a99690a <=( (not A236)  and  (not A235) );
 a99693a <=( (not A268)  and  (not A266) );
 a99694a <=( a99693a  and  a99690a );
 a99697a <=( A298  and  (not A269) );
 a99700a <=( (not A302)  and  (not A301) );
 a99701a <=( a99700a  and  a99697a );
 a99702a <=( a99701a  and  a99694a );
 a99705a <=( A169  and  (not A170) );
 a99708a <=( A166  and  A167 );
 a99709a <=( a99708a  and  a99705a );
 a99712a <=( (not A202)  and  (not A200) );
 a99715a <=( (not A233)  and  (not A203) );
 a99716a <=( a99715a  and  a99712a );
 a99717a <=( a99716a  and  a99709a );
 a99720a <=( (not A236)  and  (not A235) );
 a99723a <=( (not A268)  and  (not A266) );
 a99724a <=( a99723a  and  a99720a );
 a99727a <=( A298  and  (not A269) );
 a99730a <=( (not A302)  and  (not A301) );
 a99731a <=( a99730a  and  a99727a );
 a99732a <=( a99731a  and  a99724a );
 a99735a <=( A169  and  (not A170) );
 a99738a <=( (not A166)  and  (not A167) );
 a99739a <=( a99738a  and  a99735a );
 a99742a <=( (not A202)  and  (not A200) );
 a99745a <=( (not A233)  and  (not A203) );
 a99746a <=( a99745a  and  a99742a );
 a99747a <=( a99746a  and  a99739a );
 a99750a <=( (not A236)  and  (not A235) );
 a99753a <=( (not A268)  and  (not A266) );
 a99754a <=( a99753a  and  a99750a );
 a99757a <=( A298  and  (not A269) );
 a99760a <=( (not A302)  and  (not A301) );
 a99761a <=( a99760a  and  a99757a );
 a99762a <=( a99761a  and  a99754a );
 a99765a <=( (not A167)  and  (not A169) );
 a99768a <=( A199  and  (not A166) );
 a99769a <=( a99768a  and  a99765a );
 a99772a <=( A201  and  (not A200) );
 a99775a <=( (not A233)  and  A202 );
 a99776a <=( a99775a  and  a99772a );
 a99777a <=( a99776a  and  a99769a );
 a99780a <=( (not A236)  and  (not A235) );
 a99783a <=( (not A268)  and  (not A266) );
 a99784a <=( a99783a  and  a99780a );
 a99787a <=( A298  and  (not A269) );
 a99790a <=( (not A302)  and  (not A301) );
 a99791a <=( a99790a  and  a99787a );
 a99792a <=( a99791a  and  a99784a );
 a99795a <=( (not A167)  and  (not A169) );
 a99798a <=( A199  and  (not A166) );
 a99799a <=( a99798a  and  a99795a );
 a99802a <=( A201  and  (not A200) );
 a99805a <=( (not A233)  and  A203 );
 a99806a <=( a99805a  and  a99802a );
 a99807a <=( a99806a  and  a99799a );
 a99810a <=( (not A236)  and  (not A235) );
 a99813a <=( (not A268)  and  (not A266) );
 a99814a <=( a99813a  and  a99810a );
 a99817a <=( A298  and  (not A269) );
 a99820a <=( (not A302)  and  (not A301) );
 a99821a <=( a99820a  and  a99817a );
 a99822a <=( a99821a  and  a99814a );
 a99825a <=( (not A168)  and  (not A169) );
 a99828a <=( A166  and  A167 );
 a99829a <=( a99828a  and  a99825a );
 a99832a <=( (not A200)  and  A199 );
 a99835a <=( A202  and  A201 );
 a99836a <=( a99835a  and  a99832a );
 a99837a <=( a99836a  and  a99829a );
 a99840a <=( A233  and  A232 );
 a99843a <=( (not A268)  and  A265 );
 a99844a <=( a99843a  and  a99840a );
 a99847a <=( (not A299)  and  (not A269) );
 a99850a <=( (not A302)  and  (not A301) );
 a99851a <=( a99850a  and  a99847a );
 a99852a <=( a99851a  and  a99844a );
 a99855a <=( (not A168)  and  (not A169) );
 a99858a <=( A166  and  A167 );
 a99859a <=( a99858a  and  a99855a );
 a99862a <=( (not A200)  and  A199 );
 a99865a <=( A202  and  A201 );
 a99866a <=( a99865a  and  a99862a );
 a99867a <=( a99866a  and  a99859a );
 a99870a <=( (not A235)  and  (not A233) );
 a99873a <=( A265  and  (not A236) );
 a99874a <=( a99873a  and  a99870a );
 a99877a <=( A298  and  A266 );
 a99880a <=( (not A302)  and  (not A301) );
 a99881a <=( a99880a  and  a99877a );
 a99882a <=( a99881a  and  a99874a );
 a99885a <=( (not A168)  and  (not A169) );
 a99888a <=( A166  and  A167 );
 a99889a <=( a99888a  and  a99885a );
 a99892a <=( (not A200)  and  A199 );
 a99895a <=( A202  and  A201 );
 a99896a <=( a99895a  and  a99892a );
 a99897a <=( a99896a  and  a99889a );
 a99900a <=( (not A235)  and  (not A233) );
 a99903a <=( (not A266)  and  (not A236) );
 a99904a <=( a99903a  and  a99900a );
 a99907a <=( (not A269)  and  (not A268) );
 a99910a <=( (not A300)  and  A298 );
 a99911a <=( a99910a  and  a99907a );
 a99912a <=( a99911a  and  a99904a );
 a99915a <=( (not A168)  and  (not A169) );
 a99918a <=( A166  and  A167 );
 a99919a <=( a99918a  and  a99915a );
 a99922a <=( (not A200)  and  A199 );
 a99925a <=( A202  and  A201 );
 a99926a <=( a99925a  and  a99922a );
 a99927a <=( a99926a  and  a99919a );
 a99930a <=( (not A235)  and  (not A233) );
 a99933a <=( (not A266)  and  (not A236) );
 a99934a <=( a99933a  and  a99930a );
 a99937a <=( (not A269)  and  (not A268) );
 a99940a <=( A299  and  A298 );
 a99941a <=( a99940a  and  a99937a );
 a99942a <=( a99941a  and  a99934a );
 a99945a <=( (not A168)  and  (not A169) );
 a99948a <=( A166  and  A167 );
 a99949a <=( a99948a  and  a99945a );
 a99952a <=( (not A200)  and  A199 );
 a99955a <=( A202  and  A201 );
 a99956a <=( a99955a  and  a99952a );
 a99957a <=( a99956a  and  a99949a );
 a99960a <=( (not A235)  and  (not A233) );
 a99963a <=( (not A266)  and  (not A236) );
 a99964a <=( a99963a  and  a99960a );
 a99967a <=( (not A269)  and  (not A268) );
 a99970a <=( (not A299)  and  (not A298) );
 a99971a <=( a99970a  and  a99967a );
 a99972a <=( a99971a  and  a99964a );
 a99975a <=( (not A168)  and  (not A169) );
 a99978a <=( A166  and  A167 );
 a99979a <=( a99978a  and  a99975a );
 a99982a <=( (not A200)  and  A199 );
 a99985a <=( A202  and  A201 );
 a99986a <=( a99985a  and  a99982a );
 a99987a <=( a99986a  and  a99979a );
 a99990a <=( (not A235)  and  (not A233) );
 a99993a <=( (not A266)  and  (not A236) );
 a99994a <=( a99993a  and  a99990a );
 a99997a <=( A298  and  (not A267) );
 a100000a <=( (not A302)  and  (not A301) );
 a100001a <=( a100000a  and  a99997a );
 a100002a <=( a100001a  and  a99994a );
 a100005a <=( (not A168)  and  (not A169) );
 a100008a <=( A166  and  A167 );
 a100009a <=( a100008a  and  a100005a );
 a100012a <=( (not A200)  and  A199 );
 a100015a <=( A202  and  A201 );
 a100016a <=( a100015a  and  a100012a );
 a100017a <=( a100016a  and  a100009a );
 a100020a <=( (not A235)  and  (not A233) );
 a100023a <=( (not A265)  and  (not A236) );
 a100024a <=( a100023a  and  a100020a );
 a100027a <=( A298  and  (not A266) );
 a100030a <=( (not A302)  and  (not A301) );
 a100031a <=( a100030a  and  a100027a );
 a100032a <=( a100031a  and  a100024a );
 a100035a <=( (not A168)  and  (not A169) );
 a100038a <=( A166  and  A167 );
 a100039a <=( a100038a  and  a100035a );
 a100042a <=( (not A200)  and  A199 );
 a100045a <=( A202  and  A201 );
 a100046a <=( a100045a  and  a100042a );
 a100047a <=( a100046a  and  a100039a );
 a100050a <=( (not A234)  and  (not A233) );
 a100053a <=( (not A268)  and  (not A266) );
 a100054a <=( a100053a  and  a100050a );
 a100057a <=( A298  and  (not A269) );
 a100060a <=( (not A302)  and  (not A301) );
 a100061a <=( a100060a  and  a100057a );
 a100062a <=( a100061a  and  a100054a );
 a100065a <=( (not A168)  and  (not A169) );
 a100068a <=( A166  and  A167 );
 a100069a <=( a100068a  and  a100065a );
 a100072a <=( (not A200)  and  A199 );
 a100075a <=( A202  and  A201 );
 a100076a <=( a100075a  and  a100072a );
 a100077a <=( a100076a  and  a100069a );
 a100080a <=( (not A233)  and  A232 );
 a100083a <=( A235  and  A234 );
 a100084a <=( a100083a  and  a100080a );
 a100087a <=( (not A299)  and  A298 );
 a100090a <=( A301  and  A300 );
 a100091a <=( a100090a  and  a100087a );
 a100092a <=( a100091a  and  a100084a );
 a100095a <=( (not A168)  and  (not A169) );
 a100098a <=( A166  and  A167 );
 a100099a <=( a100098a  and  a100095a );
 a100102a <=( (not A200)  and  A199 );
 a100105a <=( A202  and  A201 );
 a100106a <=( a100105a  and  a100102a );
 a100107a <=( a100106a  and  a100099a );
 a100110a <=( (not A233)  and  A232 );
 a100113a <=( A235  and  A234 );
 a100114a <=( a100113a  and  a100110a );
 a100117a <=( (not A299)  and  A298 );
 a100120a <=( A302  and  A300 );
 a100121a <=( a100120a  and  a100117a );
 a100122a <=( a100121a  and  a100114a );
 a100125a <=( (not A168)  and  (not A169) );
 a100128a <=( A166  and  A167 );
 a100129a <=( a100128a  and  a100125a );
 a100132a <=( (not A200)  and  A199 );
 a100135a <=( A202  and  A201 );
 a100136a <=( a100135a  and  a100132a );
 a100137a <=( a100136a  and  a100129a );
 a100140a <=( (not A233)  and  A232 );
 a100143a <=( A235  and  A234 );
 a100144a <=( a100143a  and  a100140a );
 a100147a <=( (not A266)  and  A265 );
 a100150a <=( A268  and  A267 );
 a100151a <=( a100150a  and  a100147a );
 a100152a <=( a100151a  and  a100144a );
 a100155a <=( (not A168)  and  (not A169) );
 a100158a <=( A166  and  A167 );
 a100159a <=( a100158a  and  a100155a );
 a100162a <=( (not A200)  and  A199 );
 a100165a <=( A202  and  A201 );
 a100166a <=( a100165a  and  a100162a );
 a100167a <=( a100166a  and  a100159a );
 a100170a <=( (not A233)  and  A232 );
 a100173a <=( A235  and  A234 );
 a100174a <=( a100173a  and  a100170a );
 a100177a <=( (not A266)  and  A265 );
 a100180a <=( A269  and  A267 );
 a100181a <=( a100180a  and  a100177a );
 a100182a <=( a100181a  and  a100174a );
 a100185a <=( (not A168)  and  (not A169) );
 a100188a <=( A166  and  A167 );
 a100189a <=( a100188a  and  a100185a );
 a100192a <=( (not A200)  and  A199 );
 a100195a <=( A202  and  A201 );
 a100196a <=( a100195a  and  a100192a );
 a100197a <=( a100196a  and  a100189a );
 a100200a <=( (not A233)  and  A232 );
 a100203a <=( A236  and  A234 );
 a100204a <=( a100203a  and  a100200a );
 a100207a <=( (not A299)  and  A298 );
 a100210a <=( A301  and  A300 );
 a100211a <=( a100210a  and  a100207a );
 a100212a <=( a100211a  and  a100204a );
 a100215a <=( (not A168)  and  (not A169) );
 a100218a <=( A166  and  A167 );
 a100219a <=( a100218a  and  a100215a );
 a100222a <=( (not A200)  and  A199 );
 a100225a <=( A202  and  A201 );
 a100226a <=( a100225a  and  a100222a );
 a100227a <=( a100226a  and  a100219a );
 a100230a <=( (not A233)  and  A232 );
 a100233a <=( A236  and  A234 );
 a100234a <=( a100233a  and  a100230a );
 a100237a <=( (not A299)  and  A298 );
 a100240a <=( A302  and  A300 );
 a100241a <=( a100240a  and  a100237a );
 a100242a <=( a100241a  and  a100234a );
 a100245a <=( (not A168)  and  (not A169) );
 a100248a <=( A166  and  A167 );
 a100249a <=( a100248a  and  a100245a );
 a100252a <=( (not A200)  and  A199 );
 a100255a <=( A202  and  A201 );
 a100256a <=( a100255a  and  a100252a );
 a100257a <=( a100256a  and  a100249a );
 a100260a <=( (not A233)  and  A232 );
 a100263a <=( A236  and  A234 );
 a100264a <=( a100263a  and  a100260a );
 a100267a <=( (not A266)  and  A265 );
 a100270a <=( A268  and  A267 );
 a100271a <=( a100270a  and  a100267a );
 a100272a <=( a100271a  and  a100264a );
 a100275a <=( (not A168)  and  (not A169) );
 a100278a <=( A166  and  A167 );
 a100279a <=( a100278a  and  a100275a );
 a100282a <=( (not A200)  and  A199 );
 a100285a <=( A202  and  A201 );
 a100286a <=( a100285a  and  a100282a );
 a100287a <=( a100286a  and  a100279a );
 a100290a <=( (not A233)  and  A232 );
 a100293a <=( A236  and  A234 );
 a100294a <=( a100293a  and  a100290a );
 a100297a <=( (not A266)  and  A265 );
 a100300a <=( A269  and  A267 );
 a100301a <=( a100300a  and  a100297a );
 a100302a <=( a100301a  and  a100294a );
 a100305a <=( (not A168)  and  (not A169) );
 a100308a <=( A166  and  A167 );
 a100309a <=( a100308a  and  a100305a );
 a100312a <=( (not A200)  and  A199 );
 a100315a <=( A202  and  A201 );
 a100316a <=( a100315a  and  a100312a );
 a100317a <=( a100316a  and  a100309a );
 a100320a <=( (not A233)  and  (not A232) );
 a100323a <=( (not A268)  and  (not A266) );
 a100324a <=( a100323a  and  a100320a );
 a100327a <=( A298  and  (not A269) );
 a100330a <=( (not A302)  and  (not A301) );
 a100331a <=( a100330a  and  a100327a );
 a100332a <=( a100331a  and  a100324a );
 a100335a <=( (not A168)  and  (not A169) );
 a100338a <=( A166  and  A167 );
 a100339a <=( a100338a  and  a100335a );
 a100342a <=( (not A200)  and  A199 );
 a100345a <=( A203  and  A201 );
 a100346a <=( a100345a  and  a100342a );
 a100347a <=( a100346a  and  a100339a );
 a100350a <=( A233  and  A232 );
 a100353a <=( (not A268)  and  A265 );
 a100354a <=( a100353a  and  a100350a );
 a100357a <=( (not A299)  and  (not A269) );
 a100360a <=( (not A302)  and  (not A301) );
 a100361a <=( a100360a  and  a100357a );
 a100362a <=( a100361a  and  a100354a );
 a100365a <=( (not A168)  and  (not A169) );
 a100368a <=( A166  and  A167 );
 a100369a <=( a100368a  and  a100365a );
 a100372a <=( (not A200)  and  A199 );
 a100375a <=( A203  and  A201 );
 a100376a <=( a100375a  and  a100372a );
 a100377a <=( a100376a  and  a100369a );
 a100380a <=( (not A235)  and  (not A233) );
 a100383a <=( A265  and  (not A236) );
 a100384a <=( a100383a  and  a100380a );
 a100387a <=( A298  and  A266 );
 a100390a <=( (not A302)  and  (not A301) );
 a100391a <=( a100390a  and  a100387a );
 a100392a <=( a100391a  and  a100384a );
 a100395a <=( (not A168)  and  (not A169) );
 a100398a <=( A166  and  A167 );
 a100399a <=( a100398a  and  a100395a );
 a100402a <=( (not A200)  and  A199 );
 a100405a <=( A203  and  A201 );
 a100406a <=( a100405a  and  a100402a );
 a100407a <=( a100406a  and  a100399a );
 a100410a <=( (not A235)  and  (not A233) );
 a100413a <=( (not A266)  and  (not A236) );
 a100414a <=( a100413a  and  a100410a );
 a100417a <=( (not A269)  and  (not A268) );
 a100420a <=( (not A300)  and  A298 );
 a100421a <=( a100420a  and  a100417a );
 a100422a <=( a100421a  and  a100414a );
 a100425a <=( (not A168)  and  (not A169) );
 a100428a <=( A166  and  A167 );
 a100429a <=( a100428a  and  a100425a );
 a100432a <=( (not A200)  and  A199 );
 a100435a <=( A203  and  A201 );
 a100436a <=( a100435a  and  a100432a );
 a100437a <=( a100436a  and  a100429a );
 a100440a <=( (not A235)  and  (not A233) );
 a100443a <=( (not A266)  and  (not A236) );
 a100444a <=( a100443a  and  a100440a );
 a100447a <=( (not A269)  and  (not A268) );
 a100450a <=( A299  and  A298 );
 a100451a <=( a100450a  and  a100447a );
 a100452a <=( a100451a  and  a100444a );
 a100455a <=( (not A168)  and  (not A169) );
 a100458a <=( A166  and  A167 );
 a100459a <=( a100458a  and  a100455a );
 a100462a <=( (not A200)  and  A199 );
 a100465a <=( A203  and  A201 );
 a100466a <=( a100465a  and  a100462a );
 a100467a <=( a100466a  and  a100459a );
 a100470a <=( (not A235)  and  (not A233) );
 a100473a <=( (not A266)  and  (not A236) );
 a100474a <=( a100473a  and  a100470a );
 a100477a <=( (not A269)  and  (not A268) );
 a100480a <=( (not A299)  and  (not A298) );
 a100481a <=( a100480a  and  a100477a );
 a100482a <=( a100481a  and  a100474a );
 a100485a <=( (not A168)  and  (not A169) );
 a100488a <=( A166  and  A167 );
 a100489a <=( a100488a  and  a100485a );
 a100492a <=( (not A200)  and  A199 );
 a100495a <=( A203  and  A201 );
 a100496a <=( a100495a  and  a100492a );
 a100497a <=( a100496a  and  a100489a );
 a100500a <=( (not A235)  and  (not A233) );
 a100503a <=( (not A266)  and  (not A236) );
 a100504a <=( a100503a  and  a100500a );
 a100507a <=( A298  and  (not A267) );
 a100510a <=( (not A302)  and  (not A301) );
 a100511a <=( a100510a  and  a100507a );
 a100512a <=( a100511a  and  a100504a );
 a100515a <=( (not A168)  and  (not A169) );
 a100518a <=( A166  and  A167 );
 a100519a <=( a100518a  and  a100515a );
 a100522a <=( (not A200)  and  A199 );
 a100525a <=( A203  and  A201 );
 a100526a <=( a100525a  and  a100522a );
 a100527a <=( a100526a  and  a100519a );
 a100530a <=( (not A235)  and  (not A233) );
 a100533a <=( (not A265)  and  (not A236) );
 a100534a <=( a100533a  and  a100530a );
 a100537a <=( A298  and  (not A266) );
 a100540a <=( (not A302)  and  (not A301) );
 a100541a <=( a100540a  and  a100537a );
 a100542a <=( a100541a  and  a100534a );
 a100545a <=( (not A168)  and  (not A169) );
 a100548a <=( A166  and  A167 );
 a100549a <=( a100548a  and  a100545a );
 a100552a <=( (not A200)  and  A199 );
 a100555a <=( A203  and  A201 );
 a100556a <=( a100555a  and  a100552a );
 a100557a <=( a100556a  and  a100549a );
 a100560a <=( (not A234)  and  (not A233) );
 a100563a <=( (not A268)  and  (not A266) );
 a100564a <=( a100563a  and  a100560a );
 a100567a <=( A298  and  (not A269) );
 a100570a <=( (not A302)  and  (not A301) );
 a100571a <=( a100570a  and  a100567a );
 a100572a <=( a100571a  and  a100564a );
 a100575a <=( (not A168)  and  (not A169) );
 a100578a <=( A166  and  A167 );
 a100579a <=( a100578a  and  a100575a );
 a100582a <=( (not A200)  and  A199 );
 a100585a <=( A203  and  A201 );
 a100586a <=( a100585a  and  a100582a );
 a100587a <=( a100586a  and  a100579a );
 a100590a <=( (not A233)  and  A232 );
 a100593a <=( A235  and  A234 );
 a100594a <=( a100593a  and  a100590a );
 a100597a <=( (not A299)  and  A298 );
 a100600a <=( A301  and  A300 );
 a100601a <=( a100600a  and  a100597a );
 a100602a <=( a100601a  and  a100594a );
 a100605a <=( (not A168)  and  (not A169) );
 a100608a <=( A166  and  A167 );
 a100609a <=( a100608a  and  a100605a );
 a100612a <=( (not A200)  and  A199 );
 a100615a <=( A203  and  A201 );
 a100616a <=( a100615a  and  a100612a );
 a100617a <=( a100616a  and  a100609a );
 a100620a <=( (not A233)  and  A232 );
 a100623a <=( A235  and  A234 );
 a100624a <=( a100623a  and  a100620a );
 a100627a <=( (not A299)  and  A298 );
 a100630a <=( A302  and  A300 );
 a100631a <=( a100630a  and  a100627a );
 a100632a <=( a100631a  and  a100624a );
 a100635a <=( (not A168)  and  (not A169) );
 a100638a <=( A166  and  A167 );
 a100639a <=( a100638a  and  a100635a );
 a100642a <=( (not A200)  and  A199 );
 a100645a <=( A203  and  A201 );
 a100646a <=( a100645a  and  a100642a );
 a100647a <=( a100646a  and  a100639a );
 a100650a <=( (not A233)  and  A232 );
 a100653a <=( A235  and  A234 );
 a100654a <=( a100653a  and  a100650a );
 a100657a <=( (not A266)  and  A265 );
 a100660a <=( A268  and  A267 );
 a100661a <=( a100660a  and  a100657a );
 a100662a <=( a100661a  and  a100654a );
 a100665a <=( (not A168)  and  (not A169) );
 a100668a <=( A166  and  A167 );
 a100669a <=( a100668a  and  a100665a );
 a100672a <=( (not A200)  and  A199 );
 a100675a <=( A203  and  A201 );
 a100676a <=( a100675a  and  a100672a );
 a100677a <=( a100676a  and  a100669a );
 a100680a <=( (not A233)  and  A232 );
 a100683a <=( A235  and  A234 );
 a100684a <=( a100683a  and  a100680a );
 a100687a <=( (not A266)  and  A265 );
 a100690a <=( A269  and  A267 );
 a100691a <=( a100690a  and  a100687a );
 a100692a <=( a100691a  and  a100684a );
 a100695a <=( (not A168)  and  (not A169) );
 a100698a <=( A166  and  A167 );
 a100699a <=( a100698a  and  a100695a );
 a100702a <=( (not A200)  and  A199 );
 a100705a <=( A203  and  A201 );
 a100706a <=( a100705a  and  a100702a );
 a100707a <=( a100706a  and  a100699a );
 a100710a <=( (not A233)  and  A232 );
 a100713a <=( A236  and  A234 );
 a100714a <=( a100713a  and  a100710a );
 a100717a <=( (not A299)  and  A298 );
 a100720a <=( A301  and  A300 );
 a100721a <=( a100720a  and  a100717a );
 a100722a <=( a100721a  and  a100714a );
 a100725a <=( (not A168)  and  (not A169) );
 a100728a <=( A166  and  A167 );
 a100729a <=( a100728a  and  a100725a );
 a100732a <=( (not A200)  and  A199 );
 a100735a <=( A203  and  A201 );
 a100736a <=( a100735a  and  a100732a );
 a100737a <=( a100736a  and  a100729a );
 a100740a <=( (not A233)  and  A232 );
 a100743a <=( A236  and  A234 );
 a100744a <=( a100743a  and  a100740a );
 a100747a <=( (not A299)  and  A298 );
 a100750a <=( A302  and  A300 );
 a100751a <=( a100750a  and  a100747a );
 a100752a <=( a100751a  and  a100744a );
 a100755a <=( (not A168)  and  (not A169) );
 a100758a <=( A166  and  A167 );
 a100759a <=( a100758a  and  a100755a );
 a100762a <=( (not A200)  and  A199 );
 a100765a <=( A203  and  A201 );
 a100766a <=( a100765a  and  a100762a );
 a100767a <=( a100766a  and  a100759a );
 a100770a <=( (not A233)  and  A232 );
 a100773a <=( A236  and  A234 );
 a100774a <=( a100773a  and  a100770a );
 a100777a <=( (not A266)  and  A265 );
 a100780a <=( A268  and  A267 );
 a100781a <=( a100780a  and  a100777a );
 a100782a <=( a100781a  and  a100774a );
 a100785a <=( (not A168)  and  (not A169) );
 a100788a <=( A166  and  A167 );
 a100789a <=( a100788a  and  a100785a );
 a100792a <=( (not A200)  and  A199 );
 a100795a <=( A203  and  A201 );
 a100796a <=( a100795a  and  a100792a );
 a100797a <=( a100796a  and  a100789a );
 a100800a <=( (not A233)  and  A232 );
 a100803a <=( A236  and  A234 );
 a100804a <=( a100803a  and  a100800a );
 a100807a <=( (not A266)  and  A265 );
 a100810a <=( A269  and  A267 );
 a100811a <=( a100810a  and  a100807a );
 a100812a <=( a100811a  and  a100804a );
 a100815a <=( (not A168)  and  (not A169) );
 a100818a <=( A166  and  A167 );
 a100819a <=( a100818a  and  a100815a );
 a100822a <=( (not A200)  and  A199 );
 a100825a <=( A203  and  A201 );
 a100826a <=( a100825a  and  a100822a );
 a100827a <=( a100826a  and  a100819a );
 a100830a <=( (not A233)  and  (not A232) );
 a100833a <=( (not A268)  and  (not A266) );
 a100834a <=( a100833a  and  a100830a );
 a100837a <=( A298  and  (not A269) );
 a100840a <=( (not A302)  and  (not A301) );
 a100841a <=( a100840a  and  a100837a );
 a100842a <=( a100841a  and  a100834a );
 a100845a <=( (not A169)  and  A170 );
 a100848a <=( (not A166)  and  A167 );
 a100849a <=( a100848a  and  a100845a );
 a100852a <=( (not A202)  and  (not A200) );
 a100855a <=( (not A233)  and  (not A203) );
 a100856a <=( a100855a  and  a100852a );
 a100857a <=( a100856a  and  a100849a );
 a100860a <=( (not A236)  and  (not A235) );
 a100863a <=( (not A268)  and  (not A266) );
 a100864a <=( a100863a  and  a100860a );
 a100867a <=( A298  and  (not A269) );
 a100870a <=( (not A302)  and  (not A301) );
 a100871a <=( a100870a  and  a100867a );
 a100872a <=( a100871a  and  a100864a );
 a100875a <=( (not A169)  and  A170 );
 a100878a <=( A166  and  (not A167) );
 a100879a <=( a100878a  and  a100875a );
 a100882a <=( (not A202)  and  (not A200) );
 a100885a <=( (not A233)  and  (not A203) );
 a100886a <=( a100885a  and  a100882a );
 a100887a <=( a100886a  and  a100879a );
 a100890a <=( (not A236)  and  (not A235) );
 a100893a <=( (not A268)  and  (not A266) );
 a100894a <=( a100893a  and  a100890a );
 a100897a <=( A298  and  (not A269) );
 a100900a <=( (not A302)  and  (not A301) );
 a100901a <=( a100900a  and  a100897a );
 a100902a <=( a100901a  and  a100894a );
 a100905a <=( (not A169)  and  (not A170) );
 a100908a <=( A199  and  (not A168) );
 a100909a <=( a100908a  and  a100905a );
 a100912a <=( A201  and  (not A200) );
 a100915a <=( (not A233)  and  A202 );
 a100916a <=( a100915a  and  a100912a );
 a100917a <=( a100916a  and  a100909a );
 a100920a <=( (not A236)  and  (not A235) );
 a100923a <=( (not A268)  and  (not A266) );
 a100924a <=( a100923a  and  a100920a );
 a100927a <=( A298  and  (not A269) );
 a100930a <=( (not A302)  and  (not A301) );
 a100931a <=( a100930a  and  a100927a );
 a100932a <=( a100931a  and  a100924a );
 a100935a <=( (not A169)  and  (not A170) );
 a100938a <=( A199  and  (not A168) );
 a100939a <=( a100938a  and  a100935a );
 a100942a <=( A201  and  (not A200) );
 a100945a <=( (not A233)  and  A203 );
 a100946a <=( a100945a  and  a100942a );
 a100947a <=( a100946a  and  a100939a );
 a100950a <=( (not A236)  and  (not A235) );
 a100953a <=( (not A268)  and  (not A266) );
 a100954a <=( a100953a  and  a100950a );
 a100957a <=( A298  and  (not A269) );
 a100960a <=( (not A302)  and  (not A301) );
 a100961a <=( a100960a  and  a100957a );
 a100962a <=( a100961a  and  a100954a );
 a100965a <=( (not A168)  and  A169 );
 a100968a <=( (not A166)  and  A167 );
 a100969a <=( a100968a  and  a100965a );
 a100972a <=( (not A200)  and  A199 );
 a100975a <=( A202  and  A201 );
 a100976a <=( a100975a  and  a100972a );
 a100977a <=( a100976a  and  a100969a );
 a100980a <=( (not A235)  and  (not A233) );
 a100983a <=( (not A266)  and  (not A236) );
 a100984a <=( a100983a  and  a100980a );
 a100987a <=( (not A269)  and  (not A268) );
 a100991a <=( (not A302)  and  (not A301) );
 a100992a <=( A298  and  a100991a );
 a100993a <=( a100992a  and  a100987a );
 a100994a <=( a100993a  and  a100984a );
 a100997a <=( (not A168)  and  A169 );
 a101000a <=( (not A166)  and  A167 );
 a101001a <=( a101000a  and  a100997a );
 a101004a <=( (not A200)  and  A199 );
 a101007a <=( A203  and  A201 );
 a101008a <=( a101007a  and  a101004a );
 a101009a <=( a101008a  and  a101001a );
 a101012a <=( (not A235)  and  (not A233) );
 a101015a <=( (not A266)  and  (not A236) );
 a101016a <=( a101015a  and  a101012a );
 a101019a <=( (not A269)  and  (not A268) );
 a101023a <=( (not A302)  and  (not A301) );
 a101024a <=( A298  and  a101023a );
 a101025a <=( a101024a  and  a101019a );
 a101026a <=( a101025a  and  a101016a );
 a101029a <=( (not A168)  and  A169 );
 a101032a <=( A166  and  (not A167) );
 a101033a <=( a101032a  and  a101029a );
 a101036a <=( (not A200)  and  A199 );
 a101039a <=( A202  and  A201 );
 a101040a <=( a101039a  and  a101036a );
 a101041a <=( a101040a  and  a101033a );
 a101044a <=( (not A235)  and  (not A233) );
 a101047a <=( (not A266)  and  (not A236) );
 a101048a <=( a101047a  and  a101044a );
 a101051a <=( (not A269)  and  (not A268) );
 a101055a <=( (not A302)  and  (not A301) );
 a101056a <=( A298  and  a101055a );
 a101057a <=( a101056a  and  a101051a );
 a101058a <=( a101057a  and  a101048a );
 a101061a <=( (not A168)  and  A169 );
 a101064a <=( A166  and  (not A167) );
 a101065a <=( a101064a  and  a101061a );
 a101068a <=( (not A200)  and  A199 );
 a101071a <=( A203  and  A201 );
 a101072a <=( a101071a  and  a101068a );
 a101073a <=( a101072a  and  a101065a );
 a101076a <=( (not A235)  and  (not A233) );
 a101079a <=( (not A266)  and  (not A236) );
 a101080a <=( a101079a  and  a101076a );
 a101083a <=( (not A269)  and  (not A268) );
 a101087a <=( (not A302)  and  (not A301) );
 a101088a <=( A298  and  a101087a );
 a101089a <=( a101088a  and  a101083a );
 a101090a <=( a101089a  and  a101080a );
 a101093a <=( (not A168)  and  (not A169) );
 a101096a <=( A166  and  A167 );
 a101097a <=( a101096a  and  a101093a );
 a101100a <=( (not A200)  and  A199 );
 a101103a <=( A202  and  A201 );
 a101104a <=( a101103a  and  a101100a );
 a101105a <=( a101104a  and  a101097a );
 a101108a <=( (not A235)  and  (not A233) );
 a101111a <=( (not A266)  and  (not A236) );
 a101112a <=( a101111a  and  a101108a );
 a101115a <=( (not A269)  and  (not A268) );
 a101119a <=( (not A302)  and  (not A301) );
 a101120a <=( A298  and  a101119a );
 a101121a <=( a101120a  and  a101115a );
 a101122a <=( a101121a  and  a101112a );
 a101125a <=( (not A168)  and  (not A169) );
 a101128a <=( A166  and  A167 );
 a101129a <=( a101128a  and  a101125a );
 a101132a <=( (not A200)  and  A199 );
 a101135a <=( A203  and  A201 );
 a101136a <=( a101135a  and  a101132a );
 a101137a <=( a101136a  and  a101129a );
 a101140a <=( (not A235)  and  (not A233) );
 a101143a <=( (not A266)  and  (not A236) );
 a101144a <=( a101143a  and  a101140a );
 a101147a <=( (not A269)  and  (not A268) );
 a101151a <=( (not A302)  and  (not A301) );
 a101152a <=( A298  and  a101151a );
 a101153a <=( a101152a  and  a101147a );
 a101154a <=( a101153a  and  a101144a );


end x25_6x_behav;
