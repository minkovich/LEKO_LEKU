Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_17x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A42: buffer std_logic
);
end x25_17x;

architecture x25_17x_behav of x25_17x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1756a,a1757a,a1761a,a1762a,a1763a,a1767a,a1768a,a1771a,a1774a,a1775a,a1776a,a1777a,a1781a,a1782a,a1785a,a1788a,a1789a,a1790a,a1794a,a1795a,a1798a,a1801a,a1802a,a1803a,a1804a,a1805a,a1809a,a1810a,a1814a,a1815a,a1816a,a1820a,a1821a,a1824a,a1827a,a1828a,a1829a,a1830a,a1834a,a1835a,a1838a,a1841a,a1842a,a1843a,a1847a,a1848a,a1851a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1863a,a1864a,a1868a,a1869a,a1870a,a1874a,a1875a,a1878a,a1881a,a1882a,a1883a,a1884a,a1888a,a1889a,a1892a,a1895a,a1896a,a1897a,a1901a,a1902a,a1905a,a1908a,a1909a,a1910a,a1911a,a1912a,a1916a,a1917a,a1920a,a1923a,a1924a,a1925a,a1929a,a1930a,a1933a,a1936a,a1937a,a1938a,a1939a,a1943a,a1944a,a1947a,a1950a,a1951a,a1952a,a1956a,a1957a,a1960a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1973a,a1974a,a1978a,a1979a,a1980a,a1984a,a1985a,a1988a,a1991a,a1992a,a1993a,a1994a,a1998a,a1999a,a2002a,a2005a,a2006a,a2007a,a2011a,a2012a,a2015a,a2018a,a2019a,a2020a,a2021a,a2022a,a2026a,a2027a,a2030a,a2033a,a2034a,a2035a,a2039a,a2040a,a2043a,a2046a,a2047a,a2048a,a2049a,a2053a,a2054a,a2057a,a2060a,a2061a,a2062a,a2066a,a2067a,a2070a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2082a,a2083a,a2087a,a2088a,a2089a,a2093a,a2094a,a2097a,a2100a,a2101a,a2102a,a2103a,a2107a,a2108a,a2111a,a2114a,a2115a,a2116a,a2120a,a2121a,a2124a,a2127a,a2128a,a2129a,a2130a,a2131a,a2135a,a2136a,a2139a,a2142a,a2143a,a2144a,a2148a,a2149a,a2152a,a2155a,a2156a,a2157a,a2158a,a2162a,a2163a,a2166a,a2169a,a2170a,a2171a,a2175a,a2176a,a2179a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2193a,a2194a,a2198a,a2199a,a2200a,a2204a,a2205a,a2208a,a2211a,a2212a,a2213a,a2214a,a2218a,a2219a,a2222a,a2225a,a2226a,a2227a,a2231a,a2232a,a2235a,a2238a,a2239a,a2240a,a2241a,a2242a,a2246a,a2247a,a2251a,a2252a,a2253a,a2257a,a2258a,a2261a,a2264a,a2265a,a2266a,a2267a,a2271a,a2272a,a2275a,a2278a,a2279a,a2280a,a2284a,a2285a,a2288a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2300a,a2301a,a2305a,a2306a,a2307a,a2311a,a2312a,a2315a,a2318a,a2319a,a2320a,a2321a,a2325a,a2326a,a2329a,a2332a,a2333a,a2334a,a2338a,a2339a,a2342a,a2345a,a2346a,a2347a,a2348a,a2349a,a2353a,a2354a,a2357a,a2360a,a2361a,a2362a,a2366a,a2367a,a2370a,a2373a,a2374a,a2375a,a2376a,a2380a,a2381a,a2384a,a2387a,a2388a,a2389a,a2393a,a2394a,a2397a,a2400a,a2401a,a2402a,a2403a,a2404a,a2405a,a2406a,a2410a,a2411a,a2415a,a2416a,a2417a,a2421a,a2422a,a2425a,a2428a,a2429a,a2430a,a2431a,a2435a,a2436a,a2439a,a2442a,a2443a,a2444a,a2448a,a2449a,a2452a,a2455a,a2456a,a2457a,a2458a,a2459a,a2463a,a2464a,a2467a,a2470a,a2471a,a2472a,a2476a,a2477a,a2480a,a2483a,a2484a,a2485a,a2486a,a2490a,a2491a,a2494a,a2497a,a2498a,a2499a,a2503a,a2504a,a2507a,a2510a,a2511a,a2512a,a2513a,a2514a,a2515a,a2519a,a2520a,a2524a,a2525a,a2526a,a2530a,a2531a,a2534a,a2537a,a2538a,a2539a,a2540a,a2544a,a2545a,a2548a,a2551a,a2552a,a2553a,a2557a,a2558a,a2561a,a2564a,a2565a,a2566a,a2567a,a2568a,a2572a,a2573a,a2576a,a2579a,a2580a,a2581a,a2585a,a2586a,a2589a,a2592a,a2593a,a2594a,a2595a,a2599a,a2600a,a2603a,a2606a,a2607a,a2608a,a2612a,a2613a,a2616a,a2619a,a2620a,a2621a,a2622a,a2623a,a2624a,a2625a,a2626a,a2627a,a2631a,a2632a,a2636a,a2637a,a2638a,a2642a,a2643a,a2646a,a2649a,a2650a,a2651a,a2652a,a2656a,a2657a,a2660a,a2663a,a2664a,a2665a,a2669a,a2670a,a2673a,a2676a,a2677a,a2678a,a2679a,a2680a,a2684a,a2685a,a2689a,a2690a,a2691a,a2695a,a2696a,a2699a,a2702a,a2703a,a2704a,a2705a,a2709a,a2710a,a2713a,a2716a,a2717a,a2718a,a2722a,a2723a,a2726a,a2729a,a2730a,a2731a,a2732a,a2733a,a2734a,a2738a,a2739a,a2743a,a2744a,a2745a,a2749a,a2750a,a2753a,a2756a,a2757a,a2758a,a2759a,a2763a,a2764a,a2767a,a2770a,a2771a,a2772a,a2776a,a2777a,a2780a,a2783a,a2784a,a2785a,a2786a,a2787a,a2791a,a2792a,a2795a,a2798a,a2799a,a2800a,a2804a,a2805a,a2808a,a2811a,a2812a,a2813a,a2814a,a2818a,a2819a,a2822a,a2825a,a2826a,a2827a,a2831a,a2832a,a2835a,a2838a,a2839a,a2840a,a2841a,a2842a,a2843a,a2844a,a2848a,a2849a,a2853a,a2854a,a2855a,a2859a,a2860a,a2863a,a2866a,a2867a,a2868a,a2869a,a2873a,a2874a,a2877a,a2880a,a2881a,a2882a,a2886a,a2887a,a2890a,a2893a,a2894a,a2895a,a2896a,a2897a,a2901a,a2902a,a2905a,a2908a,a2909a,a2910a,a2914a,a2915a,a2918a,a2921a,a2922a,a2923a,a2924a,a2928a,a2929a,a2932a,a2935a,a2936a,a2937a,a2941a,a2942a,a2945a,a2948a,a2949a,a2950a,a2951a,a2952a,a2953a,a2957a,a2958a,a2962a,a2963a,a2964a,a2968a,a2969a,a2972a,a2975a,a2976a,a2977a,a2978a,a2982a,a2983a,a2986a,a2989a,a2990a,a2991a,a2995a,a2996a,a2999a,a3002a,a3003a,a3004a,a3005a,a3006a,a3010a,a3011a,a3014a,a3017a,a3018a,a3019a,a3023a,a3024a,a3027a,a3030a,a3031a,a3032a,a3033a,a3037a,a3038a,a3041a,a3044a,a3045a,a3046a,a3050a,a3051a,a3054a,a3057a,a3058a,a3059a,a3060a,a3061a,a3062a,a3063a,a3064a,a3068a,a3069a,a3073a,a3074a,a3075a,a3079a,a3080a,a3083a,a3086a,a3087a,a3088a,a3089a,a3093a,a3094a,a3097a,a3100a,a3101a,a3102a,a3106a,a3107a,a3110a,a3113a,a3114a,a3115a,a3116a,a3117a,a3121a,a3122a,a3126a,a3127a,a3128a,a3132a,a3133a,a3136a,a3139a,a3140a,a3141a,a3142a,a3146a,a3147a,a3150a,a3153a,a3154a,a3155a,a3159a,a3160a,a3163a,a3166a,a3167a,a3168a,a3169a,a3170a,a3171a,a3175a,a3176a,a3180a,a3181a,a3182a,a3186a,a3187a,a3190a,a3193a,a3194a,a3195a,a3196a,a3200a,a3201a,a3204a,a3207a,a3208a,a3209a,a3213a,a3214a,a3217a,a3220a,a3221a,a3222a,a3223a,a3224a,a3228a,a3229a,a3232a,a3235a,a3236a,a3237a,a3241a,a3242a,a3245a,a3248a,a3249a,a3250a,a3251a,a3255a,a3256a,a3259a,a3262a,a3263a,a3264a,a3268a,a3269a,a3272a,a3275a,a3276a,a3277a,a3278a,a3279a,a3280a,a3281a,a3285a,a3286a,a3290a,a3291a,a3292a,a3296a,a3297a,a3300a,a3303a,a3304a,a3305a,a3306a,a3310a,a3311a,a3314a,a3317a,a3318a,a3319a,a3323a,a3324a,a3327a,a3330a,a3331a,a3332a,a3333a,a3334a,a3338a,a3339a,a3342a,a3345a,a3346a,a3347a,a3351a,a3352a,a3355a,a3358a,a3359a,a3360a,a3361a,a3365a,a3366a,a3369a,a3372a,a3373a,a3374a,a3378a,a3379a,a3382a,a3385a,a3386a,a3387a,a3388a,a3389a,a3390a,a3394a,a3395a,a3399a,a3400a,a3401a,a3405a,a3406a,a3409a,a3412a,a3413a,a3414a,a3415a,a3419a,a3420a,a3423a,a3426a,a3427a,a3428a,a3432a,a3433a,a3436a,a3439a,a3440a,a3441a,a3442a,a3443a,a3447a,a3448a,a3451a,a3454a,a3455a,a3456a,a3460a,a3461a,a3464a,a3467a,a3468a,a3469a,a3470a,a3474a,a3475a,a3478a,a3481a,a3482a,a3483a,a3487a,a3488a,a3491a,a3494a,a3495a,a3496a,a3497a,a3498a,a3499a,a3500a,a3501a,a3502a,a3503a,a3507a,a3508a,a3512a,a3513a,a3514a,a3518a,a3519a,a3522a,a3525a,a3526a,a3527a,a3528a,a3532a,a3533a,a3536a,a3539a,a3540a,a3541a,a3545a,a3546a,a3549a,a3552a,a3553a,a3554a,a3555a,a3556a,a3560a,a3561a,a3565a,a3566a,a3567a,a3571a,a3572a,a3575a,a3578a,a3579a,a3580a,a3581a,a3585a,a3586a,a3589a,a3592a,a3593a,a3594a,a3598a,a3599a,a3602a,a3605a,a3606a,a3607a,a3608a,a3609a,a3610a,a3614a,a3615a,a3619a,a3620a,a3621a,a3625a,a3626a,a3629a,a3632a,a3633a,a3634a,a3635a,a3639a,a3640a,a3643a,a3646a,a3647a,a3648a,a3652a,a3653a,a3656a,a3659a,a3660a,a3661a,a3662a,a3663a,a3667a,a3668a,a3671a,a3674a,a3675a,a3676a,a3680a,a3681a,a3684a,a3687a,a3688a,a3689a,a3690a,a3694a,a3695a,a3698a,a3701a,a3702a,a3703a,a3707a,a3708a,a3711a,a3714a,a3715a,a3716a,a3717a,a3718a,a3719a,a3720a,a3724a,a3725a,a3729a,a3730a,a3731a,a3735a,a3736a,a3739a,a3742a,a3743a,a3744a,a3745a,a3749a,a3750a,a3753a,a3756a,a3757a,a3758a,a3762a,a3763a,a3766a,a3769a,a3770a,a3771a,a3772a,a3773a,a3777a,a3778a,a3781a,a3784a,a3785a,a3786a,a3790a,a3791a,a3794a,a3797a,a3798a,a3799a,a3800a,a3804a,a3805a,a3808a,a3811a,a3812a,a3813a,a3817a,a3818a,a3821a,a3824a,a3825a,a3826a,a3827a,a3828a,a3829a,a3833a,a3834a,a3838a,a3839a,a3840a,a3844a,a3845a,a3848a,a3851a,a3852a,a3853a,a3854a,a3858a,a3859a,a3862a,a3865a,a3866a,a3867a,a3871a,a3872a,a3875a,a3878a,a3879a,a3880a,a3881a,a3882a,a3886a,a3887a,a3890a,a3893a,a3894a,a3895a,a3899a,a3900a,a3903a,a3906a,a3907a,a3908a,a3909a,a3913a,a3914a,a3917a,a3920a,a3921a,a3922a,a3926a,a3927a,a3930a,a3933a,a3934a,a3935a,a3936a,a3937a,a3938a,a3939a,a3940a,a3944a,a3945a,a3949a,a3950a,a3951a,a3955a,a3956a,a3959a,a3962a,a3963a,a3964a,a3965a,a3969a,a3970a,a3973a,a3976a,a3977a,a3978a,a3982a,a3983a,a3986a,a3989a,a3990a,a3991a,a3992a,a3993a,a3997a,a3998a,a4002a,a4003a,a4004a,a4008a,a4009a,a4012a,a4015a,a4016a,a4017a,a4018a,a4022a,a4023a,a4026a,a4029a,a4030a,a4031a,a4035a,a4036a,a4039a,a4042a,a4043a,a4044a,a4045a,a4046a,a4047a,a4051a,a4052a,a4056a,a4057a,a4058a,a4062a,a4063a,a4066a,a4069a,a4070a,a4071a,a4072a,a4076a,a4077a,a4080a,a4083a,a4084a,a4085a,a4089a,a4090a,a4093a,a4096a,a4097a,a4098a,a4099a,a4100a,a4104a,a4105a,a4108a,a4111a,a4112a,a4113a,a4117a,a4118a,a4121a,a4124a,a4125a,a4126a,a4127a,a4131a,a4132a,a4135a,a4138a,a4139a,a4140a,a4144a,a4145a,a4148a,a4151a,a4152a,a4153a,a4154a,a4155a,a4156a,a4157a,a4161a,a4162a,a4166a,a4167a,a4168a,a4172a,a4173a,a4176a,a4179a,a4180a,a4181a,a4182a,a4186a,a4187a,a4190a,a4193a,a4194a,a4195a,a4199a,a4200a,a4203a,a4206a,a4207a,a4208a,a4209a,a4210a,a4214a,a4215a,a4218a,a4221a,a4222a,a4223a,a4227a,a4228a,a4231a,a4234a,a4235a,a4236a,a4237a,a4241a,a4242a,a4245a,a4248a,a4249a,a4250a,a4254a,a4255a,a4258a,a4261a,a4262a,a4263a,a4264a,a4265a,a4266a,a4270a,a4271a,a4275a,a4276a,a4277a,a4281a,a4282a,a4285a,a4288a,a4289a,a4290a,a4291a,a4295a,a4296a,a4299a,a4302a,a4303a,a4304a,a4308a,a4309a,a4312a,a4315a,a4316a,a4317a,a4318a,a4319a,a4323a,a4324a,a4327a,a4330a,a4331a,a4332a,a4336a,a4337a,a4340a,a4343a,a4344a,a4345a,a4346a,a4350a,a4351a,a4354a,a4357a,a4358a,a4359a,a4363a,a4364a,a4367a,a4370a,a4371a,a4372a,a4373a,a4374a,a4375a,a4376a,a4377a,a4378a,a4382a,a4383a,a4387a,a4388a,a4389a,a4393a,a4394a,a4397a,a4400a,a4401a,a4402a,a4403a,a4407a,a4408a,a4411a,a4414a,a4415a,a4416a,a4420a,a4421a,a4424a,a4427a,a4428a,a4429a,a4430a,a4431a,a4435a,a4436a,a4440a,a4441a,a4442a,a4446a,a4447a,a4450a,a4453a,a4454a,a4455a,a4456a,a4460a,a4461a,a4464a,a4467a,a4468a,a4469a,a4473a,a4474a,a4477a,a4480a,a4481a,a4482a,a4483a,a4484a,a4485a,a4489a,a4490a,a4494a,a4495a,a4496a,a4500a,a4501a,a4504a,a4507a,a4508a,a4509a,a4510a,a4514a,a4515a,a4518a,a4521a,a4522a,a4523a,a4527a,a4528a,a4531a,a4534a,a4535a,a4536a,a4537a,a4538a,a4542a,a4543a,a4546a,a4549a,a4550a,a4551a,a4555a,a4556a,a4559a,a4562a,a4563a,a4564a,a4565a,a4569a,a4570a,a4573a,a4576a,a4577a,a4578a,a4582a,a4583a,a4586a,a4589a,a4590a,a4591a,a4592a,a4593a,a4594a,a4595a,a4599a,a4600a,a4604a,a4605a,a4606a,a4610a,a4611a,a4614a,a4617a,a4618a,a4619a,a4620a,a4624a,a4625a,a4628a,a4631a,a4632a,a4633a,a4637a,a4638a,a4641a,a4644a,a4645a,a4646a,a4647a,a4648a,a4652a,a4653a,a4656a,a4659a,a4660a,a4661a,a4665a,a4666a,a4669a,a4672a,a4673a,a4674a,a4675a,a4679a,a4680a,a4683a,a4686a,a4687a,a4688a,a4692a,a4693a,a4696a,a4699a,a4700a,a4701a,a4702a,a4703a,a4704a,a4708a,a4709a,a4713a,a4714a,a4715a,a4719a,a4720a,a4723a,a4726a,a4727a,a4728a,a4729a,a4733a,a4734a,a4737a,a4740a,a4741a,a4742a,a4746a,a4747a,a4750a,a4753a,a4754a,a4755a,a4756a,a4757a,a4761a,a4762a,a4765a,a4768a,a4769a,a4770a,a4774a,a4775a,a4778a,a4781a,a4782a,a4783a,a4784a,a4788a,a4789a,a4792a,a4795a,a4796a,a4797a,a4801a,a4802a,a4805a,a4808a,a4809a,a4810a,a4811a,a4812a,a4813a,a4814a,a4815a,a4819a,a4820a,a4824a,a4825a,a4826a,a4830a,a4831a,a4834a,a4837a,a4838a,a4839a,a4840a,a4844a,a4845a,a4848a,a4851a,a4852a,a4853a,a4857a,a4858a,a4861a,a4864a,a4865a,a4866a,a4867a,a4868a,a4872a,a4873a,a4877a,a4878a,a4879a,a4883a,a4884a,a4887a,a4890a,a4891a,a4892a,a4893a,a4897a,a4898a,a4901a,a4904a,a4905a,a4906a,a4910a,a4911a,a4914a,a4917a,a4918a,a4919a,a4920a,a4921a,a4922a,a4926a,a4927a,a4931a,a4932a,a4933a,a4937a,a4938a,a4941a,a4944a,a4945a,a4946a,a4947a,a4951a,a4952a,a4955a,a4958a,a4959a,a4960a,a4964a,a4965a,a4968a,a4971a,a4972a,a4973a,a4974a,a4975a,a4979a,a4980a,a4983a,a4986a,a4987a,a4988a,a4992a,a4993a,a4996a,a4999a,a5000a,a5001a,a5002a,a5006a,a5007a,a5010a,a5013a,a5014a,a5015a,a5019a,a5020a,a5023a,a5026a,a5027a,a5028a,a5029a,a5030a,a5031a,a5032a,a5036a,a5037a,a5041a,a5042a,a5043a,a5047a,a5048a,a5051a,a5054a,a5055a,a5056a,a5057a,a5061a,a5062a,a5065a,a5068a,a5069a,a5070a,a5074a,a5075a,a5078a,a5081a,a5082a,a5083a,a5084a,a5085a,a5089a,a5090a,a5093a,a5096a,a5097a,a5098a,a5102a,a5103a,a5106a,a5109a,a5110a,a5111a,a5112a,a5116a,a5117a,a5120a,a5123a,a5124a,a5125a,a5129a,a5130a,a5133a,a5136a,a5137a,a5138a,a5139a,a5140a,a5141a,a5145a,a5146a,a5150a,a5151a,a5152a,a5156a,a5157a,a5160a,a5163a,a5164a,a5165a,a5166a,a5170a,a5171a,a5174a,a5177a,a5178a,a5179a,a5183a,a5184a,a5187a,a5190a,a5191a,a5192a,a5193a,a5194a,a5198a,a5199a,a5202a,a5205a,a5206a,a5207a,a5211a,a5212a,a5215a,a5218a,a5219a,a5220a,a5221a,a5225a,a5226a,a5229a,a5232a,a5233a,a5234a,a5238a,a5239a,a5242a,a5245a,a5246a,a5247a,a5248a,a5249a,a5250a,a5251a,a5252a,a5253a,a5254a,a5257a,a5260a,a5263a,a5266a,a5269a,a5272a,a5275a,a5278a,a5281a,a5284a,a5287a,a5290a,a5293a,a5297a,a5298a,a5301a,a5305a,a5306a,a5310a,a5311a,a5315a,a5316a,a5320a,a5321a,a5325a,a5326a,a5330a,a5331a,a5335a,a5336a,a5340a,a5341a,a5345a,a5346a,a5350a,a5351a,a5355a,a5356a,a5360a,a5361a,a5365a,a5366a,a5370a,a5371a,a5375a,a5376a,a5380a,a5381a,a5385a,a5386a,a5390a,a5391a,a5395a,a5396a,a5400a,a5401a,a5405a,a5406a,a5410a,a5411a,a5415a,a5416a,a5420a,a5421a,a5425a,a5426a,a5430a,a5431a,a5434a,a5437a,a5438a,a5442a,a5443a,a5446a,a5449a,a5450a,a5454a,a5455a,a5458a,a5461a,a5462a,a5466a,a5467a,a5470a,a5473a,a5474a,a5477a,a5480a,a5481a,a5484a,a5488a,a5489a,a5490a,a5493a,a5496a,a5497a,a5500a,a5504a,a5505a,a5506a,a5509a,a5512a,a5513a,a5516a,a5520a,a5521a,a5522a,a5525a,a5528a,a5529a,a5532a,a5536a,a5537a,a5538a,a5541a,a5544a,a5545a,a5548a,a5552a,a5553a,a5554a,a5557a,a5560a,a5561a,a5564a,a5568a,a5569a,a5570a,a5573a,a5576a,a5577a,a5580a,a5584a,a5585a,a5586a,a5589a,a5592a,a5593a,a5596a,a5600a,a5601a,a5602a,a5605a,a5608a,a5609a,a5612a,a5616a,a5617a,a5618a,a5621a,a5624a,a5625a,a5628a,a5632a,a5633a,a5634a,a5637a,a5640a,a5641a,a5644a,a5648a,a5649a,a5650a,a5653a,a5656a,a5657a,a5660a,a5664a,a5665a,a5666a,a5669a,a5672a,a5673a,a5676a,a5680a,a5681a,a5682a,a5685a,a5688a,a5689a,a5692a,a5696a,a5697a,a5698a,a5701a,a5704a,a5705a,a5708a,a5712a,a5713a,a5714a,a5717a,a5720a,a5721a,a5724a,a5728a,a5729a,a5730a,a5733a,a5737a,a5738a,a5739a,a5742a,a5746a,a5747a,a5748a,a5751a,a5755a,a5756a,a5757a,a5760a,a5764a,a5765a,a5766a,a5769a,a5773a,a5774a,a5775a,a5778a,a5782a,a5783a,a5784a,a5787a,a5791a,a5792a,a5793a,a5796a,a5800a,a5801a,a5802a,a5805a,a5809a,a5810a,a5811a,a5814a,a5818a,a5819a,a5820a,a5823a,a5827a,a5828a,a5829a,a5832a,a5836a,a5837a,a5838a,a5841a,a5845a,a5846a,a5847a,a5850a,a5854a,a5855a,a5856a,a5859a,a5863a,a5864a,a5865a,a5868a,a5872a,a5873a,a5874a,a5877a,a5881a,a5882a,a5883a,a5886a,a5890a,a5891a,a5892a,a5895a,a5899a,a5900a,a5901a,a5904a,a5908a,a5909a,a5910a,a5913a,a5917a,a5918a,a5919a,a5922a,a5926a,a5927a,a5928a,a5931a,a5935a,a5936a,a5937a,a5940a,a5944a,a5945a,a5946a,a5949a,a5953a,a5954a,a5955a,a5958a,a5962a,a5963a,a5964a,a5967a,a5971a,a5972a,a5973a,a5976a,a5980a,a5981a,a5982a,a5985a,a5989a,a5990a,a5991a,a5994a,a5998a,a5999a,a6000a,a6003a,a6007a,a6008a,a6009a,a6012a,a6016a,a6017a,a6018a,a6021a,a6025a,a6026a,a6027a,a6030a,a6034a,a6035a,a6036a,a6039a,a6043a,a6044a,a6045a,a6048a,a6052a,a6053a,a6054a,a6057a,a6061a,a6062a,a6063a,a6066a,a6070a,a6071a,a6072a,a6075a,a6079a,a6080a,a6081a,a6084a,a6088a,a6089a,a6090a,a6093a,a6097a,a6098a,a6099a,a6102a,a6106a,a6107a,a6108a,a6111a,a6115a,a6116a,a6117a,a6120a,a6124a,a6125a,a6126a,a6129a,a6133a,a6134a,a6135a,a6138a,a6142a,a6143a,a6144a,a6147a,a6151a,a6152a,a6153a,a6156a,a6160a,a6161a,a6162a,a6165a,a6169a,a6170a,a6171a,a6174a,a6178a,a6179a,a6180a,a6183a,a6187a,a6188a,a6189a,a6192a,a6196a,a6197a,a6198a,a6201a,a6205a,a6206a,a6207a,a6210a,a6214a,a6215a,a6216a,a6219a,a6223a,a6224a,a6225a,a6228a,a6232a,a6233a,a6234a,a6237a,a6241a,a6242a,a6243a,a6246a,a6250a,a6251a,a6252a,a6255a,a6259a,a6260a,a6261a,a6264a,a6268a,a6269a,a6270a,a6273a,a6277a,a6278a,a6279a,a6282a,a6286a,a6287a,a6288a,a6291a,a6295a,a6296a,a6297a,a6300a,a6304a,a6305a,a6306a,a6309a,a6313a,a6314a,a6315a,a6318a,a6322a,a6323a,a6324a,a6327a,a6331a,a6332a,a6333a,a6336a,a6340a,a6341a,a6342a,a6345a,a6349a,a6350a,a6351a,a6354a,a6358a,a6359a,a6360a,a6363a,a6367a,a6368a,a6369a,a6372a,a6376a,a6377a,a6378a,a6381a,a6385a,a6386a,a6387a,a6390a,a6394a,a6395a,a6396a,a6399a,a6403a,a6404a,a6405a,a6408a,a6412a,a6413a,a6414a,a6417a,a6421a,a6422a,a6423a,a6426a,a6430a,a6431a,a6432a,a6435a,a6439a,a6440a,a6441a,a6444a,a6448a,a6449a,a6450a,a6453a,a6457a,a6458a,a6459a,a6462a,a6466a,a6467a,a6468a,a6471a,a6475a,a6476a,a6477a,a6480a,a6484a,a6485a,a6486a,a6489a,a6493a,a6494a,a6495a,a6498a,a6502a,a6503a,a6504a,a6507a,a6511a,a6512a,a6513a,a6516a,a6520a,a6521a,a6522a,a6525a,a6529a,a6530a,a6531a,a6534a,a6538a,a6539a,a6540a,a6543a,a6547a,a6548a,a6549a,a6552a,a6556a,a6557a,a6558a,a6561a,a6565a,a6566a,a6567a,a6570a,a6574a,a6575a,a6576a,a6579a,a6583a,a6584a,a6585a,a6588a,a6592a,a6593a,a6594a,a6597a,a6601a,a6602a,a6603a,a6607a,a6608a,a6612a,a6613a,a6614a,a6617a,a6621a,a6622a,a6623a,a6627a,a6628a,a6632a,a6633a,a6634a,a6637a,a6641a,a6642a,a6643a,a6647a,a6648a,a6652a,a6653a,a6654a,a6657a,a6661a,a6662a,a6663a,a6667a,a6668a,a6672a,a6673a,a6674a,a6677a,a6681a,a6682a,a6683a,a6687a,a6688a,a6692a,a6693a,a6694a,a6697a,a6701a,a6702a,a6703a,a6707a,a6708a,a6712a,a6713a,a6714a,a6717a,a6721a,a6722a,a6723a,a6727a,a6728a,a6732a,a6733a,a6734a,a6737a,a6741a,a6742a,a6743a,a6747a,a6748a,a6752a,a6753a,a6754a,a6757a,a6761a,a6762a,a6763a,a6767a,a6768a,a6772a,a6773a,a6774a,a6777a,a6781a,a6782a,a6783a,a6787a,a6788a,a6792a,a6793a,a6794a,a6797a,a6801a,a6802a,a6803a,a6807a,a6808a,a6812a,a6813a,a6814a,a6817a,a6821a,a6822a,a6823a,a6827a,a6828a,a6832a,a6833a,a6834a,a6837a,a6841a,a6842a,a6843a,a6847a,a6848a,a6852a,a6853a,a6854a,a6857a,a6861a,a6862a,a6863a,a6867a,a6868a,a6872a,a6873a,a6874a,a6877a,a6881a,a6882a,a6883a,a6887a,a6888a,a6892a,a6893a,a6894a,a6897a,a6901a,a6902a,a6903a,a6907a,a6908a,a6912a,a6913a,a6914a,a6917a,a6921a,a6922a,a6923a,a6927a,a6928a,a6932a,a6933a,a6934a,a6937a,a6941a,a6942a,a6943a,a6947a,a6948a,a6952a,a6953a,a6954a,a6957a,a6961a,a6962a,a6963a,a6967a,a6968a,a6972a,a6973a,a6974a,a6977a,a6981a,a6982a,a6983a,a6987a,a6988a,a6992a,a6993a,a6994a,a6997a,a7001a,a7002a,a7003a,a7007a,a7008a,a7012a,a7013a,a7014a,a7017a,a7021a,a7022a,a7023a,a7027a,a7028a,a7032a,a7033a,a7034a,a7037a,a7041a,a7042a,a7043a,a7047a,a7048a,a7052a,a7053a,a7054a,a7057a,a7061a,a7062a,a7063a,a7067a,a7068a,a7072a,a7073a,a7074a,a7077a,a7081a,a7082a,a7083a,a7087a,a7088a,a7092a,a7093a,a7094a,a7097a,a7101a,a7102a,a7103a,a7107a,a7108a,a7112a,a7113a,a7114a,a7117a,a7121a,a7122a,a7123a,a7127a,a7128a,a7132a,a7133a,a7134a,a7137a,a7141a,a7142a,a7143a,a7147a,a7148a,a7152a,a7153a,a7154a,a7157a,a7161a,a7162a,a7163a,a7167a,a7168a,a7172a,a7173a,a7174a,a7177a,a7181a,a7182a,a7183a,a7187a,a7188a,a7192a,a7193a,a7194a,a7197a,a7201a,a7202a,a7203a,a7207a,a7208a,a7212a,a7213a,a7214a,a7217a,a7221a,a7222a,a7223a,a7227a,a7228a,a7232a,a7233a,a7234a,a7237a,a7241a,a7242a,a7243a,a7247a,a7248a,a7252a,a7253a,a7254a,a7257a,a7261a,a7262a,a7263a,a7267a,a7268a,a7272a,a7273a,a7274a,a7277a,a7281a,a7282a,a7283a,a7287a,a7288a,a7292a,a7293a,a7294a,a7297a,a7301a,a7302a,a7303a,a7307a,a7308a,a7312a,a7313a,a7314a,a7317a,a7321a,a7322a,a7323a,a7327a,a7328a,a7332a,a7333a,a7334a,a7337a,a7341a,a7342a,a7343a,a7347a,a7348a,a7352a,a7353a,a7354a,a7357a,a7361a,a7362a,a7363a,a7367a,a7368a,a7372a,a7373a,a7374a,a7377a,a7381a,a7382a,a7383a,a7387a,a7388a,a7392a,a7393a,a7394a,a7397a,a7401a,a7402a,a7403a,a7407a,a7408a,a7412a,a7413a,a7414a,a7417a,a7421a,a7422a,a7423a,a7427a,a7428a,a7432a,a7433a,a7434a,a7437a,a7441a,a7442a,a7443a,a7447a,a7448a,a7452a,a7453a,a7454a,a7457a,a7461a,a7462a,a7463a,a7467a,a7468a,a7472a,a7473a,a7474a,a7477a,a7481a,a7482a,a7483a,a7487a,a7488a,a7492a,a7493a,a7494a,a7497a,a7501a,a7502a,a7503a,a7507a,a7508a,a7512a,a7513a,a7514a,a7517a,a7521a,a7522a,a7523a,a7527a,a7528a,a7532a,a7533a,a7534a,a7537a,a7541a,a7542a,a7543a,a7547a,a7548a,a7552a,a7553a,a7554a,a7557a,a7561a,a7562a,a7563a,a7567a,a7568a,a7572a,a7573a,a7574a,a7577a,a7581a,a7582a,a7583a,a7587a,a7588a,a7592a,a7593a,a7594a,a7597a,a7601a,a7602a,a7603a,a7607a,a7608a,a7612a,a7613a,a7614a,a7617a,a7621a,a7622a,a7623a,a7627a,a7628a,a7632a,a7633a,a7634a,a7637a,a7641a,a7642a,a7643a,a7647a,a7648a,a7652a,a7653a,a7654a,a7657a,a7661a,a7662a,a7663a,a7667a,a7668a,a7672a,a7673a,a7674a,a7677a,a7681a,a7682a,a7683a,a7687a,a7688a,a7692a,a7693a,a7694a,a7697a,a7701a,a7702a,a7703a,a7707a,a7708a,a7712a,a7713a,a7714a,a7717a,a7721a,a7722a,a7723a,a7727a,a7728a,a7732a,a7733a,a7734a,a7737a,a7741a,a7742a,a7743a,a7747a,a7748a,a7752a,a7753a,a7754a,a7757a,a7761a,a7762a,a7763a,a7767a,a7768a,a7772a,a7773a,a7774a,a7777a,a7781a,a7782a,a7783a,a7787a,a7788a,a7792a,a7793a,a7794a,a7797a,a7801a,a7802a,a7803a,a7807a,a7808a,a7812a,a7813a,a7814a,a7817a,a7821a,a7822a,a7823a,a7827a,a7828a,a7832a,a7833a,a7834a,a7837a,a7841a,a7842a,a7843a,a7847a,a7848a,a7852a,a7853a,a7854a,a7857a,a7861a,a7862a,a7863a,a7867a,a7868a,a7872a,a7873a,a7874a,a7877a,a7881a,a7882a,a7883a,a7887a,a7888a,a7892a,a7893a,a7894a,a7897a,a7901a,a7902a,a7903a,a7907a,a7908a,a7912a,a7913a,a7914a,a7917a,a7921a,a7922a,a7923a,a7927a,a7928a,a7932a,a7933a,a7934a,a7937a,a7941a,a7942a,a7943a,a7947a,a7948a,a7952a,a7953a,a7954a,a7957a,a7961a,a7962a,a7963a,a7967a,a7968a,a7972a,a7973a,a7974a,a7977a,a7981a,a7982a,a7983a,a7987a,a7988a,a7992a,a7993a,a7994a,a7997a,a8001a,a8002a,a8003a,a8007a,a8008a,a8012a,a8013a,a8014a,a8017a,a8021a,a8022a,a8023a,a8027a,a8028a,a8032a,a8033a,a8034a,a8037a,a8041a,a8042a,a8043a,a8047a,a8048a,a8052a,a8053a,a8054a,a8057a,a8061a,a8062a,a8063a,a8067a,a8068a,a8072a,a8073a,a8074a,a8077a,a8081a,a8082a,a8083a,a8087a,a8088a,a8092a,a8093a,a8094a,a8097a,a8101a,a8102a,a8103a,a8107a,a8108a,a8112a,a8113a,a8114a,a8117a,a8121a,a8122a,a8123a,a8127a,a8128a,a8132a,a8133a,a8134a,a8137a,a8141a,a8142a,a8143a,a8147a,a8148a,a8152a,a8153a,a8154a,a8157a,a8161a,a8162a,a8163a,a8167a,a8168a,a8172a,a8173a,a8174a,a8177a,a8181a,a8182a,a8183a,a8187a,a8188a,a8192a,a8193a,a8194a,a8197a,a8201a,a8202a,a8203a,a8207a,a8208a,a8212a,a8213a,a8214a,a8217a,a8221a,a8222a,a8223a,a8227a,a8228a,a8232a,a8233a,a8234a,a8237a,a8241a,a8242a,a8243a,a8247a,a8248a,a8252a,a8253a,a8254a,a8257a,a8261a,a8262a,a8263a,a8267a,a8268a,a8272a,a8273a,a8274a,a8277a,a8281a,a8282a,a8283a,a8287a,a8288a,a8292a,a8293a,a8294a,a8297a,a8301a,a8302a,a8303a,a8307a,a8308a,a8312a,a8313a,a8314a,a8317a,a8321a,a8322a,a8323a,a8327a,a8328a,a8332a,a8333a,a8334a,a8337a,a8341a,a8342a,a8343a,a8347a,a8348a,a8352a,a8353a,a8354a,a8357a,a8361a,a8362a,a8363a,a8367a,a8368a,a8372a,a8373a,a8374a,a8377a,a8381a,a8382a,a8383a,a8387a,a8388a,a8392a,a8393a,a8394a,a8397a,a8401a,a8402a,a8403a,a8407a,a8408a,a8412a,a8413a,a8414a,a8417a,a8421a,a8422a,a8423a,a8427a,a8428a,a8432a,a8433a,a8434a,a8437a,a8441a,a8442a,a8443a,a8447a,a8448a,a8452a,a8453a,a8454a,a8457a,a8461a,a8462a,a8463a,a8467a,a8468a,a8472a,a8473a,a8474a,a8477a,a8481a,a8482a,a8483a,a8487a,a8488a,a8492a,a8493a,a8494a,a8497a,a8501a,a8502a,a8503a,a8507a,a8508a,a8512a,a8513a,a8514a,a8518a,a8519a,a8523a,a8524a,a8525a,a8529a,a8530a,a8534a,a8535a,a8536a,a8540a,a8541a,a8545a,a8546a,a8547a,a8551a,a8552a,a8556a,a8557a,a8558a,a8562a,a8563a,a8567a,a8568a,a8569a,a8573a,a8574a,a8578a,a8579a,a8580a,a8584a,a8585a,a8589a,a8590a,a8591a,a8595a,a8596a,a8600a,a8601a,a8602a,a8606a,a8607a,a8611a,a8612a,a8613a,a8617a,a8618a,a8622a,a8623a,a8624a,a8628a,a8629a,a8633a,a8634a,a8635a,a8639a,a8640a,a8644a,a8645a,a8646a,a8650a,a8651a,a8655a,a8656a,a8657a,a8661a,a8662a,a8666a,a8667a,a8668a,a8672a,a8673a,a8677a,a8678a,a8679a,a8683a,a8684a,a8688a,a8689a,a8690a,a8694a,a8695a,a8699a,a8700a,a8701a,a8705a,a8706a,a8710a,a8711a,a8712a,a8716a,a8717a,a8721a,a8722a,a8723a,a8727a,a8728a,a8732a,a8733a,a8734a,a8738a,a8739a,a8743a,a8744a,a8745a,a8749a,a8750a,a8754a,a8755a,a8756a,a8760a,a8761a,a8765a,a8766a,a8767a,a8771a,a8772a,a8776a,a8777a,a8778a,a8782a,a8783a,a8787a,a8788a,a8789a,a8793a,a8794a,a8798a,a8799a,a8800a,a8804a,a8805a,a8809a,a8810a,a8811a,a8815a,a8816a,a8820a,a8821a,a8822a,a8826a,a8827a,a8831a,a8832a,a8833a,a8837a,a8838a,a8842a,a8843a,a8844a,a8848a,a8849a,a8853a,a8854a,a8855a,a8859a,a8860a,a8864a,a8865a,a8866a,a8870a,a8871a,a8875a,a8876a,a8877a,a8881a,a8882a,a8886a,a8887a,a8888a,a8892a,a8893a,a8897a,a8898a,a8899a,a8903a,a8904a,a8908a,a8909a,a8910a,a8914a,a8915a,a8919a,a8920a,a8921a,a8925a,a8926a,a8930a,a8931a,a8932a,a8936a,a8937a,a8941a,a8942a,a8943a,a8947a,a8948a,a8952a,a8953a,a8954a,a8958a,a8959a,a8963a,a8964a,a8965a,a8969a,a8970a,a8974a,a8975a,a8976a,a8980a,a8981a,a8985a,a8986a,a8987a,a8991a,a8992a,a8996a,a8997a,a8998a,a9002a,a9003a,a9007a,a9008a,a9009a,a9013a,a9014a,a9018a,a9019a,a9020a,a9024a,a9025a,a9029a,a9030a,a9031a,a9035a,a9036a,a9040a,a9041a,a9042a,a9046a,a9047a,a9051a,a9052a,a9053a,a9057a,a9058a,a9062a,a9063a,a9064a,a9068a,a9069a,a9073a,a9074a,a9075a,a9079a,a9080a,a9084a,a9085a,a9086a,a9090a,a9091a,a9095a,a9096a,a9097a,a9101a,a9102a,a9106a,a9107a,a9108a,a9112a,a9113a,a9117a,a9118a,a9119a,a9123a,a9124a,a9128a,a9129a,a9130a,a9134a,a9135a,a9139a,a9140a,a9141a,a9145a,a9146a,a9150a,a9151a,a9152a,a9156a,a9157a,a9161a,a9162a,a9163a,a9167a,a9168a,a9172a,a9173a,a9174a,a9178a,a9179a,a9183a,a9184a,a9185a,a9189a,a9190a,a9194a,a9195a,a9196a,a9200a,a9201a,a9205a,a9206a,a9207a,a9211a,a9212a,a9216a,a9217a,a9218a,a9222a,a9223a,a9227a,a9228a,a9229a,a9233a,a9234a,a9238a,a9239a,a9240a,a9244a,a9245a,a9249a,a9250a,a9251a,a9255a,a9256a,a9260a,a9261a,a9262a,a9266a,a9267a,a9271a,a9272a,a9273a,a9277a,a9278a,a9282a,a9283a,a9284a,a9288a,a9289a,a9293a,a9294a,a9295a,a9299a,a9300a,a9304a,a9305a,a9306a,a9310a,a9311a,a9315a,a9316a,a9317a,a9321a,a9322a,a9326a,a9327a,a9328a,a9332a,a9333a,a9337a,a9338a,a9339a,a9343a,a9344a,a9348a,a9349a,a9350a,a9354a,a9355a,a9359a,a9360a,a9361a,a9365a,a9366a,a9370a,a9371a,a9372a,a9376a,a9377a,a9381a,a9382a,a9383a,a9387a,a9388a,a9392a,a9393a,a9394a,a9398a,a9399a,a9403a,a9404a,a9405a,a9409a,a9410a,a9414a,a9415a,a9416a,a9420a,a9421a,a9425a,a9426a,a9427a,a9431a,a9432a,a9436a,a9437a,a9438a,a9442a,a9443a,a9447a,a9448a,a9449a,a9453a,a9454a,a9458a,a9459a,a9460a,a9464a,a9465a,a9469a,a9470a,a9471a,a9475a,a9476a,a9480a,a9481a,a9482a,a9486a,a9487a,a9491a,a9492a,a9493a,a9497a,a9498a,a9502a,a9503a,a9504a,a9508a,a9509a,a9513a,a9514a,a9515a,a9519a,a9520a,a9524a,a9525a,a9526a,a9530a,a9531a,a9535a,a9536a,a9537a,a9541a,a9542a,a9546a,a9547a,a9548a,a9552a,a9553a,a9557a,a9558a,a9559a,a9563a,a9564a,a9568a,a9569a,a9570a,a9574a,a9575a,a9579a,a9580a,a9581a,a9585a,a9586a,a9590a,a9591a,a9592a,a9596a,a9597a,a9601a,a9602a,a9603a,a9607a,a9608a,a9612a,a9613a,a9614a,a9618a,a9619a,a9623a,a9624a,a9625a,a9629a,a9630a,a9634a,a9635a,a9636a,a9640a,a9641a,a9645a,a9646a,a9647a,a9651a,a9652a,a9656a,a9657a,a9658a,a9662a,a9663a,a9667a,a9668a,a9669a,a9673a,a9674a,a9678a,a9679a,a9680a,a9684a,a9685a,a9689a,a9690a,a9691a,a9695a,a9696a,a9700a,a9701a,a9702a,a9706a,a9707a,a9711a,a9712a,a9713a,a9717a,a9718a,a9722a,a9723a,a9724a,a9728a,a9729a,a9733a,a9734a,a9735a,a9739a,a9740a,a9744a,a9745a,a9746a,a9750a,a9751a,a9755a,a9756a,a9757a,a9761a,a9762a,a9766a,a9767a,a9768a,a9772a,a9773a,a9777a,a9778a,a9779a,a9783a,a9784a,a9788a,a9789a,a9790a,a9794a,a9795a,a9799a,a9800a,a9801a,a9805a,a9806a,a9810a,a9811a,a9812a,a9816a,a9817a,a9821a,a9822a,a9823a,a9827a,a9828a,a9832a,a9833a,a9834a,a9838a,a9839a,a9843a,a9844a,a9845a,a9849a,a9850a,a9854a,a9855a,a9856a,a9860a,a9861a,a9865a,a9866a,a9867a,a9871a,a9872a,a9876a,a9877a,a9878a,a9882a,a9883a,a9887a,a9888a,a9889a,a9893a,a9894a,a9898a,a9899a,a9900a,a9904a,a9905a,a9909a,a9910a,a9911a,a9915a,a9916a,a9920a,a9921a,a9922a,a9926a,a9927a,a9931a,a9932a,a9933a,a9937a,a9938a,a9942a,a9943a,a9944a,a9948a,a9949a,a9953a,a9954a,a9955a,a9959a,a9960a,a9964a,a9965a,a9966a,a9970a,a9971a,a9975a,a9976a,a9977a,a9981a,a9982a,a9986a,a9987a,a9988a,a9992a,a9993a,a9997a,a9998a,a9999a,a10003a,a10004a,a10008a,a10009a,a10010a,a10014a,a10015a,a10019a,a10020a,a10021a,a10025a,a10026a,a10030a,a10031a,a10032a,a10036a,a10037a,a10041a,a10042a,a10043a,a10047a,a10048a,a10052a,a10053a,a10054a,a10058a,a10059a,a10063a,a10064a,a10065a,a10069a,a10070a,a10074a,a10075a,a10076a,a10080a,a10081a,a10085a,a10086a,a10087a,a10091a,a10092a,a10096a,a10097a,a10098a,a10102a,a10103a,a10107a,a10108a,a10109a,a10113a,a10114a,a10118a,a10119a,a10120a,a10124a,a10125a,a10129a,a10130a,a10131a,a10135a,a10136a,a10140a,a10141a,a10142a,a10146a,a10147a,a10151a,a10152a,a10153a,a10157a,a10158a,a10162a,a10163a,a10164a,a10168a,a10169a,a10173a,a10174a,a10175a,a10179a,a10180a,a10184a,a10185a,a10186a,a10190a,a10191a,a10195a,a10196a,a10197a,a10201a,a10202a,a10206a,a10207a,a10208a,a10212a,a10213a,a10217a,a10218a,a10219a,a10223a,a10224a,a10228a,a10229a,a10230a,a10234a,a10235a,a10239a,a10240a,a10241a,a10245a,a10246a,a10250a,a10251a,a10252a,a10256a,a10257a,a10261a,a10262a,a10263a,a10267a,a10268a,a10272a,a10273a,a10274a,a10278a,a10279a,a10283a,a10284a,a10285a,a10289a,a10290a,a10294a,a10295a,a10296a,a10300a,a10301a,a10305a,a10306a,a10307a,a10311a,a10312a,a10316a,a10317a,a10318a,a10322a,a10323a,a10327a,a10328a,a10329a,a10333a,a10334a,a10338a,a10339a,a10340a,a10344a,a10345a,a10349a,a10350a,a10351a,a10355a,a10356a,a10360a,a10361a,a10362a,a10366a,a10367a,a10371a,a10372a,a10373a,a10377a,a10378a,a10382a,a10383a,a10384a,a10388a,a10389a,a10393a,a10394a,a10395a,a10399a,a10400a,a10404a,a10405a,a10406a,a10410a,a10411a,a10415a,a10416a,a10417a,a10421a,a10422a,a10426a,a10427a,a10428a,a10432a,a10433a,a10437a,a10438a,a10439a,a10443a,a10444a,a10448a,a10449a,a10450a,a10454a,a10455a,a10459a,a10460a,a10461a,a10465a,a10466a,a10470a,a10471a,a10472a,a10476a,a10477a,a10481a,a10482a,a10483a,a10487a,a10488a,a10492a,a10493a,a10494a,a10498a,a10499a,a10503a,a10504a,a10505a,a10509a,a10510a,a10514a,a10515a,a10516a,a10520a,a10521a,a10525a,a10526a,a10527a,a10531a,a10532a,a10536a,a10537a,a10538a,a10542a,a10543a,a10547a,a10548a,a10549a,a10553a,a10554a,a10558a,a10559a,a10560a,a10564a,a10565a,a10569a,a10570a,a10571a,a10575a,a10576a,a10580a,a10581a,a10582a,a10586a,a10587a,a10591a,a10592a,a10593a,a10597a,a10598a,a10602a,a10603a,a10604a,a10608a,a10609a,a10613a,a10614a,a10615a,a10619a,a10620a,a10624a,a10625a,a10626a,a10630a,a10631a,a10635a,a10636a,a10637a,a10641a,a10642a,a10646a,a10647a,a10648a,a10652a,a10653a,a10657a,a10658a,a10659a,a10663a,a10664a,a10668a,a10669a,a10670a,a10674a,a10675a,a10679a,a10680a,a10681a,a10685a,a10686a,a10690a,a10691a,a10692a,a10696a,a10697a,a10701a,a10702a,a10703a,a10707a,a10708a,a10712a,a10713a,a10714a,a10718a,a10719a,a10723a,a10724a,a10725a,a10729a,a10730a,a10734a,a10735a,a10736a,a10740a,a10741a,a10745a,a10746a,a10747a,a10751a,a10752a,a10756a,a10757a,a10758a,a10762a,a10763a,a10767a,a10768a,a10769a,a10773a,a10774a,a10778a,a10779a,a10780a,a10784a,a10785a,a10789a,a10790a,a10791a,a10795a,a10796a,a10800a,a10801a,a10802a,a10806a,a10807a,a10811a,a10812a,a10813a,a10817a,a10818a,a10822a,a10823a,a10824a,a10828a,a10829a,a10833a,a10834a,a10835a,a10839a,a10840a,a10844a,a10845a,a10846a,a10850a,a10851a,a10855a,a10856a,a10857a,a10861a,a10862a,a10866a,a10867a,a10868a,a10872a,a10873a,a10877a,a10878a,a10879a,a10883a,a10884a,a10888a,a10889a,a10890a,a10894a,a10895a,a10899a,a10900a,a10901a,a10905a,a10906a,a10910a,a10911a,a10912a,a10916a,a10917a,a10921a,a10922a,a10923a,a10927a,a10928a,a10932a,a10933a,a10934a,a10938a,a10939a,a10943a,a10944a,a10945a,a10949a,a10950a,a10954a,a10955a,a10956a,a10960a,a10961a,a10965a,a10966a,a10967a,a10971a,a10972a,a10976a,a10977a,a10978a,a10982a,a10983a,a10987a,a10988a,a10989a,a10993a,a10994a,a10998a,a10999a,a11000a,a11004a,a11005a,a11009a,a11010a,a11011a,a11015a,a11016a,a11020a,a11021a,a11022a,a11026a,a11027a,a11031a,a11032a,a11033a,a11037a,a11038a,a11042a,a11043a,a11044a,a11048a,a11049a,a11053a,a11054a,a11055a,a11059a,a11060a,a11064a,a11065a,a11066a,a11070a,a11071a,a11075a,a11076a,a11077a,a11081a,a11082a,a11086a,a11087a,a11088a,a11092a,a11093a,a11097a,a11098a,a11099a,a11103a,a11104a,a11108a,a11109a,a11110a,a11114a,a11115a,a11119a,a11120a,a11121a,a11125a,a11126a,a11130a,a11131a,a11132a,a11136a,a11137a,a11141a,a11142a,a11143a,a11147a,a11148a,a11152a,a11153a,a11154a,a11158a,a11159a,a11163a,a11164a,a11165a,a11169a,a11170a,a11174a,a11175a,a11176a,a11180a,a11181a,a11185a,a11186a,a11187a,a11191a,a11192a,a11196a,a11197a,a11198a,a11202a,a11203a,a11207a,a11208a,a11209a,a11213a,a11214a,a11218a,a11219a,a11220a,a11224a,a11225a,a11229a,a11230a,a11231a,a11235a,a11236a,a11240a,a11241a,a11242a,a11246a,a11247a,a11251a,a11252a,a11253a,a11257a,a11258a,a11262a,a11263a,a11264a,a11268a,a11269a,a11273a,a11274a,a11275a,a11279a,a11280a,a11284a,a11285a,a11286a,a11290a,a11291a,a11295a,a11296a,a11297a,a11301a,a11302a,a11306a,a11307a,a11308a,a11312a,a11313a,a11317a,a11318a,a11319a,a11323a,a11324a,a11328a,a11329a,a11330a,a11334a,a11335a,a11339a,a11340a,a11341a,a11345a,a11346a,a11350a,a11351a,a11352a,a11356a,a11357a,a11361a,a11362a,a11363a,a11367a,a11368a,a11372a,a11373a,a11374a,a11378a,a11379a,a11383a,a11384a,a11385a,a11389a,a11390a,a11394a,a11395a,a11396a,a11400a,a11401a,a11405a,a11406a,a11407a,a11411a,a11412a,a11416a,a11417a,a11418a,a11422a,a11423a,a11427a,a11428a,a11429a,a11433a,a11434a,a11438a,a11439a,a11440a,a11444a,a11445a,a11449a,a11450a,a11451a,a11455a,a11456a,a11460a,a11461a,a11462a,a11466a,a11467a,a11471a,a11472a,a11473a,a11477a,a11478a,a11482a,a11483a,a11484a,a11488a,a11489a,a11493a,a11494a,a11495a,a11499a,a11500a,a11504a,a11505a,a11506a,a11510a,a11511a,a11515a,a11516a,a11517a,a11521a,a11522a,a11526a,a11527a,a11528a,a11532a,a11533a,a11537a,a11538a,a11539a,a11543a,a11544a,a11548a,a11549a,a11550a,a11554a,a11555a,a11559a,a11560a,a11561a,a11565a,a11566a,a11570a,a11571a,a11572a,a11576a,a11577a,a11581a,a11582a,a11583a,a11587a,a11588a,a11592a,a11593a,a11594a,a11598a,a11599a,a11603a,a11604a,a11605a,a11609a,a11610a,a11614a,a11615a,a11616a,a11620a,a11621a,a11625a,a11626a,a11627a,a11631a,a11632a,a11636a,a11637a,a11638a,a11642a,a11643a,a11647a,a11648a,a11649a,a11653a,a11654a,a11658a,a11659a,a11660a,a11664a,a11665a,a11669a,a11670a,a11671a,a11675a,a11676a,a11680a,a11681a,a11682a,a11686a,a11687a,a11691a,a11692a,a11693a,a11697a,a11698a,a11702a,a11703a,a11704a,a11708a,a11709a,a11713a,a11714a,a11715a,a11719a,a11720a,a11724a,a11725a,a11726a,a11730a,a11731a,a11735a,a11736a,a11737a,a11741a,a11742a,a11746a,a11747a,a11748a,a11752a,a11753a,a11757a,a11758a,a11759a,a11763a,a11764a,a11768a,a11769a,a11770a,a11774a,a11775a,a11779a,a11780a,a11781a,a11785a,a11786a,a11790a,a11791a,a11792a,a11796a,a11797a,a11801a,a11802a,a11803a,a11807a,a11808a,a11812a,a11813a,a11814a,a11818a,a11819a,a11823a,a11824a,a11825a,a11829a,a11830a,a11834a,a11835a,a11836a,a11840a,a11841a,a11845a,a11846a,a11847a,a11851a,a11852a,a11856a,a11857a,a11858a,a11862a,a11863a,a11867a,a11868a,a11869a,a11873a,a11874a,a11878a,a11879a,a11880a,a11884a,a11885a,a11889a,a11890a,a11891a,a11895a,a11896a,a11900a,a11901a,a11902a,a11906a,a11907a,a11911a,a11912a,a11913a,a11917a,a11918a,a11922a,a11923a,a11924a,a11928a,a11929a,a11933a,a11934a,a11935a,a11939a,a11940a,a11944a,a11945a,a11946a,a11950a,a11951a,a11955a,a11956a,a11957a,a11961a,a11962a,a11966a,a11967a,a11968a,a11972a,a11973a,a11977a,a11978a,a11979a,a11983a,a11984a,a11988a,a11989a,a11990a,a11994a,a11995a,a11999a,a12000a,a12001a,a12005a,a12006a,a12010a,a12011a,a12012a,a12016a,a12017a,a12021a,a12022a,a12023a,a12027a,a12028a,a12032a,a12033a,a12034a,a12038a,a12039a,a12043a,a12044a,a12045a,a12049a,a12050a,a12054a,a12055a,a12056a,a12060a,a12061a,a12065a,a12066a,a12067a,a12071a,a12072a,a12076a,a12077a,a12078a,a12082a,a12083a,a12087a,a12088a,a12089a,a12093a,a12094a,a12098a,a12099a,a12100a,a12104a,a12105a,a12109a,a12110a,a12111a,a12115a,a12116a,a12120a,a12121a,a12122a,a12126a,a12127a,a12131a,a12132a,a12133a,a12137a,a12138a,a12142a,a12143a,a12144a,a12148a,a12149a,a12153a,a12154a,a12155a,a12159a,a12160a,a12164a,a12165a,a12166a,a12170a,a12171a,a12175a,a12176a,a12177a,a12181a,a12182a,a12186a,a12187a,a12188a,a12192a,a12193a,a12197a,a12198a,a12199a,a12203a,a12204a,a12208a,a12209a,a12210a,a12214a,a12215a,a12219a,a12220a,a12221a,a12225a,a12226a,a12230a,a12231a,a12232a,a12236a,a12237a,a12241a,a12242a,a12243a,a12247a,a12248a,a12252a,a12253a,a12254a,a12258a,a12259a,a12263a,a12264a,a12265a,a12269a,a12270a,a12274a,a12275a,a12276a,a12280a,a12281a,a12285a,a12286a,a12287a,a12291a,a12292a,a12296a,a12297a,a12298a,a12302a,a12303a,a12307a,a12308a,a12309a,a12313a,a12314a,a12318a,a12319a,a12320a,a12324a,a12325a,a12329a,a12330a,a12331a,a12335a,a12336a,a12340a,a12341a,a12342a,a12346a,a12347a,a12351a,a12352a,a12353a,a12357a,a12358a,a12362a,a12363a,a12364a,a12368a,a12369a,a12373a,a12374a,a12375a,a12379a,a12380a,a12384a,a12385a,a12386a,a12390a,a12391a,a12395a,a12396a,a12397a,a12401a,a12402a,a12406a,a12407a,a12408a,a12412a,a12413a,a12417a,a12418a,a12419a,a12423a,a12424a,a12428a,a12429a,a12430a,a12434a,a12435a,a12439a,a12440a,a12441a,a12445a,a12446a,a12450a,a12451a,a12452a,a12456a,a12457a,a12461a,a12462a,a12463a,a12467a,a12468a,a12472a,a12473a,a12474a,a12478a,a12479a,a12483a,a12484a,a12485a,a12489a,a12490a,a12494a,a12495a,a12496a,a12500a,a12501a,a12505a,a12506a,a12507a,a12511a,a12512a,a12516a,a12517a,a12518a,a12522a,a12523a,a12527a,a12528a,a12529a,a12533a,a12534a,a12538a,a12539a,a12540a,a12544a,a12545a,a12549a,a12550a,a12551a,a12555a,a12556a,a12560a,a12561a,a12562a,a12566a,a12567a,a12571a,a12572a,a12573a,a12577a,a12578a,a12582a,a12583a,a12584a,a12588a,a12589a,a12593a,a12594a,a12595a,a12599a,a12600a,a12604a,a12605a,a12606a,a12610a,a12611a,a12615a,a12616a,a12617a,a12621a,a12622a,a12626a,a12627a,a12628a,a12632a,a12633a,a12637a,a12638a,a12639a,a12643a,a12644a,a12648a,a12649a,a12650a,a12654a,a12655a,a12659a,a12660a,a12661a,a12665a,a12666a,a12670a,a12671a,a12672a,a12676a,a12677a,a12681a,a12682a,a12683a,a12687a,a12688a,a12692a,a12693a,a12694a,a12698a,a12699a,a12703a,a12704a,a12705a,a12709a,a12710a,a12714a,a12715a,a12716a,a12720a,a12721a,a12725a,a12726a,a12727a,a12731a,a12732a,a12736a,a12737a,a12738a,a12742a,a12743a,a12747a,a12748a,a12749a,a12753a,a12754a,a12758a,a12759a,a12760a,a12764a,a12765a,a12769a,a12770a,a12771a,a12775a,a12776a,a12780a,a12781a,a12782a,a12786a,a12787a,a12791a,a12792a,a12793a,a12797a,a12798a,a12802a,a12803a,a12804a,a12808a,a12809a,a12813a,a12814a,a12815a,a12819a,a12820a,a12824a,a12825a,a12826a,a12830a,a12831a,a12835a,a12836a,a12837a,a12841a,a12842a,a12846a,a12847a,a12848a,a12852a,a12853a,a12857a,a12858a,a12859a,a12863a,a12864a,a12868a,a12869a,a12870a,a12874a,a12875a,a12879a,a12880a,a12881a,a12885a,a12886a,a12890a,a12891a,a12892a,a12896a,a12897a,a12901a,a12902a,a12903a,a12907a,a12908a,a12912a,a12913a,a12914a,a12918a,a12919a,a12923a,a12924a,a12925a,a12929a,a12930a,a12934a,a12935a,a12936a,a12940a,a12941a,a12945a,a12946a,a12947a,a12951a,a12952a,a12956a,a12957a,a12958a,a12962a,a12963a,a12967a,a12968a,a12969a,a12973a,a12974a,a12978a,a12979a,a12980a,a12984a,a12985a,a12989a,a12990a,a12991a,a12995a,a12996a,a13000a,a13001a,a13002a,a13006a,a13007a,a13011a,a13012a,a13013a,a13017a,a13018a,a13022a,a13023a,a13024a,a13028a,a13029a,a13033a,a13034a,a13035a,a13039a,a13040a,a13044a,a13045a,a13046a,a13050a,a13051a,a13055a,a13056a,a13057a,a13061a,a13062a,a13066a,a13067a,a13068a,a13072a,a13073a,a13077a,a13078a,a13079a,a13083a,a13084a,a13088a,a13089a,a13090a,a13094a,a13095a,a13099a,a13100a,a13101a,a13105a,a13106a,a13110a,a13111a,a13112a,a13116a,a13117a,a13121a,a13122a,a13123a,a13127a,a13128a,a13132a,a13133a,a13134a,a13138a,a13139a,a13143a,a13144a,a13145a,a13149a,a13150a,a13154a,a13155a,a13156a,a13160a,a13161a,a13165a,a13166a,a13167a,a13171a,a13172a,a13176a,a13177a,a13178a,a13182a,a13183a,a13187a,a13188a,a13189a,a13193a,a13194a,a13198a,a13199a,a13200a,a13204a,a13205a,a13209a,a13210a,a13211a,a13215a,a13216a,a13220a,a13221a,a13222a,a13226a,a13227a,a13231a,a13232a,a13233a,a13237a,a13238a,a13242a,a13243a,a13244a,a13248a,a13249a,a13253a,a13254a,a13255a,a13259a,a13260a,a13264a,a13265a,a13266a,a13270a,a13271a,a13275a,a13276a,a13277a,a13281a,a13282a,a13286a,a13287a,a13288a,a13292a,a13293a,a13297a,a13298a,a13299a,a13303a,a13304a,a13308a,a13309a,a13310a,a13314a,a13315a,a13319a,a13320a,a13321a,a13325a,a13326a,a13330a,a13331a,a13332a,a13336a,a13337a,a13341a,a13342a,a13343a,a13347a,a13348a,a13352a,a13353a,a13354a,a13358a,a13359a,a13363a,a13364a,a13365a,a13369a,a13370a,a13374a,a13375a,a13376a,a13380a,a13381a,a13385a,a13386a,a13387a,a13391a,a13392a,a13396a,a13397a,a13398a,a13402a,a13403a,a13407a,a13408a,a13409a,a13413a,a13414a,a13418a,a13419a,a13420a,a13424a,a13425a,a13429a,a13430a,a13431a,a13435a,a13436a,a13440a,a13441a,a13442a,a13446a,a13447a,a13451a,a13452a,a13453a,a13457a,a13458a,a13462a,a13463a,a13464a,a13468a,a13469a,a13473a,a13474a,a13475a,a13479a,a13480a,a13484a,a13485a,a13486a,a13490a,a13491a,a13495a,a13496a,a13497a,a13501a,a13502a,a13506a,a13507a,a13508a,a13512a,a13513a,a13517a,a13518a,a13519a,a13523a,a13524a,a13528a,a13529a,a13530a,a13534a,a13535a,a13539a,a13540a,a13541a,a13545a,a13546a,a13550a,a13551a,a13552a,a13556a,a13557a,a13561a,a13562a,a13563a,a13567a,a13568a,a13572a,a13573a,a13574a,a13578a,a13579a,a13583a,a13584a,a13585a,a13589a,a13590a,a13594a,a13595a,a13596a,a13600a,a13601a,a13605a,a13606a,a13607a,a13611a,a13612a,a13616a,a13617a,a13618a,a13622a,a13623a,a13627a,a13628a,a13629a,a13633a,a13634a,a13638a,a13639a,a13640a,a13644a,a13645a,a13649a,a13650a,a13651a,a13655a,a13656a,a13660a,a13661a,a13662a,a13666a,a13667a,a13671a,a13672a,a13673a,a13677a,a13678a,a13682a,a13683a,a13684a,a13688a,a13689a,a13693a,a13694a,a13695a,a13699a,a13700a,a13704a,a13705a,a13706a,a13710a,a13711a,a13715a,a13716a,a13717a,a13721a,a13722a,a13726a,a13727a,a13728a,a13732a,a13733a,a13737a,a13738a,a13739a,a13743a,a13744a,a13748a,a13749a,a13750a,a13754a,a13755a,a13759a,a13760a,a13761a,a13765a,a13766a,a13770a,a13771a,a13772a,a13776a,a13777a,a13781a,a13782a,a13783a,a13787a,a13788a,a13792a,a13793a,a13794a,a13798a,a13799a,a13803a,a13804a,a13805a,a13809a,a13810a,a13814a,a13815a,a13816a,a13820a,a13821a,a13825a,a13826a,a13827a,a13831a,a13832a,a13836a,a13837a,a13838a,a13842a,a13843a,a13847a,a13848a,a13849a,a13853a,a13854a,a13858a,a13859a,a13860a,a13864a,a13865a,a13869a,a13870a,a13871a,a13875a,a13876a,a13880a,a13881a,a13882a,a13886a,a13887a,a13891a,a13892a,a13893a,a13897a,a13898a,a13902a,a13903a,a13904a,a13908a,a13909a,a13913a,a13914a,a13915a,a13919a,a13920a,a13924a,a13925a,a13926a,a13930a,a13931a,a13935a,a13936a,a13937a,a13941a,a13942a,a13946a,a13947a,a13948a,a13952a,a13953a,a13957a,a13958a,a13959a,a13963a,a13964a,a13968a,a13969a,a13970a,a13974a,a13975a,a13979a,a13980a,a13981a,a13985a,a13986a,a13990a,a13991a,a13992a,a13996a,a13997a,a14001a,a14002a,a14003a,a14007a,a14008a,a14012a,a14013a,a14014a,a14018a,a14019a,a14023a,a14024a,a14025a,a14029a,a14030a,a14034a,a14035a,a14036a,a14040a,a14041a,a14045a,a14046a,a14047a,a14051a,a14052a,a14056a,a14057a,a14058a,a14062a,a14063a,a14067a,a14068a,a14069a,a14073a,a14074a,a14078a,a14079a,a14080a,a14084a,a14085a,a14089a,a14090a,a14091a,a14095a,a14096a,a14100a,a14101a,a14102a,a14106a,a14107a,a14111a,a14112a,a14113a,a14117a,a14118a,a14122a,a14123a,a14124a,a14128a,a14129a,a14133a,a14134a,a14135a,a14139a,a14140a,a14144a,a14145a,a14146a,a14150a,a14151a,a14155a,a14156a,a14157a,a14161a,a14162a,a14166a,a14167a,a14168a,a14172a,a14173a,a14177a,a14178a,a14179a,a14183a,a14184a,a14188a,a14189a,a14190a,a14194a,a14195a,a14199a,a14200a,a14201a,a14205a,a14206a,a14210a,a14211a,a14212a,a14216a,a14217a,a14221a,a14222a,a14223a,a14227a,a14228a,a14232a,a14233a,a14234a,a14238a,a14239a,a14243a,a14244a,a14245a,a14249a,a14250a,a14254a,a14255a,a14256a,a14260a,a14261a,a14265a,a14266a,a14267a,a14271a,a14272a,a14276a,a14277a,a14278a,a14282a,a14283a,a14287a,a14288a,a14289a,a14293a,a14294a,a14298a,a14299a,a14300a,a14304a,a14305a,a14309a,a14310a,a14311a,a14315a,a14316a,a14320a,a14321a,a14322a,a14326a,a14327a,a14331a,a14332a,a14333a,a14337a,a14338a,a14342a,a14343a,a14344a,a14348a,a14349a,a14353a,a14354a,a14355a,a14359a,a14360a,a14364a,a14365a,a14366a,a14370a,a14371a,a14375a,a14376a,a14377a,a14381a,a14382a,a14386a,a14387a,a14388a,a14392a,a14393a,a14397a,a14398a,a14399a,a14403a,a14404a,a14408a,a14409a,a14410a,a14414a,a14415a,a14419a,a14420a,a14421a,a14425a,a14426a,a14430a,a14431a,a14432a,a14436a,a14437a,a14441a,a14442a,a14443a,a14447a,a14448a,a14452a,a14453a,a14454a,a14458a,a14459a,a14463a,a14464a,a14465a,a14469a,a14470a,a14474a,a14475a,a14476a,a14480a,a14481a,a14485a,a14486a,a14487a,a14491a,a14492a,a14496a,a14497a,a14498a,a14502a,a14503a,a14507a,a14508a,a14509a,a14513a,a14514a,a14518a,a14519a,a14520a,a14524a,a14525a,a14529a,a14530a,a14531a,a14535a,a14536a,a14540a,a14541a,a14542a,a14546a,a14547a,a14551a,a14552a,a14553a,a14557a,a14558a,a14562a,a14563a,a14564a,a14568a,a14569a,a14573a,a14574a,a14575a,a14579a,a14580a,a14584a,a14585a,a14586a,a14590a,a14591a,a14595a,a14596a,a14597a,a14601a,a14602a,a14606a,a14607a,a14608a,a14612a,a14613a,a14617a,a14618a,a14619a,a14623a,a14624a,a14628a,a14629a,a14630a,a14634a,a14635a,a14639a,a14640a,a14641a,a14645a,a14646a,a14650a,a14651a,a14652a,a14656a,a14657a,a14661a,a14662a,a14663a,a14667a,a14668a,a14672a,a14673a,a14674a,a14678a,a14679a,a14683a,a14684a,a14685a,a14689a,a14690a,a14694a,a14695a,a14696a,a14700a,a14701a,a14705a,a14706a,a14707a,a14711a,a14712a,a14716a,a14717a,a14718a,a14722a,a14723a,a14727a,a14728a,a14729a,a14733a,a14734a,a14738a,a14739a,a14740a,a14744a,a14745a,a14749a,a14750a,a14751a,a14755a,a14756a,a14760a,a14761a,a14762a,a14766a,a14767a,a14771a,a14772a,a14773a,a14777a,a14778a,a14782a,a14783a,a14784a,a14788a,a14789a,a14793a,a14794a,a14795a,a14799a,a14800a,a14804a,a14805a,a14806a,a14810a,a14811a,a14815a,a14816a,a14817a,a14821a,a14822a,a14826a,a14827a,a14828a,a14832a,a14833a,a14837a,a14838a,a14839a,a14843a,a14844a,a14848a,a14849a,a14850a,a14854a,a14855a,a14859a,a14860a,a14861a,a14865a,a14866a,a14869a,a14872a,a14873a,a14874a,a14878a,a14879a,a14883a,a14884a,a14885a,a14889a,a14890a,a14893a,a14896a,a14897a,a14898a,a14902a,a14903a,a14907a,a14908a,a14909a,a14913a,a14914a,a14917a,a14920a,a14921a,a14922a,a14926a,a14927a,a14931a,a14932a,a14933a,a14937a,a14938a,a14941a,a14944a,a14945a,a14946a,a14950a,a14951a,a14955a,a14956a,a14957a,a14961a,a14962a,a14965a,a14968a,a14969a,a14970a,a14974a,a14975a,a14979a,a14980a,a14981a,a14985a,a14986a,a14989a,a14992a,a14993a,a14994a,a14998a,a14999a,a15003a,a15004a,a15005a,a15009a,a15010a,a15013a,a15016a,a15017a,a15018a,a15022a,a15023a,a15027a,a15028a,a15029a,a15033a,a15034a,a15037a,a15040a,a15041a,a15042a,a15046a,a15047a,a15051a,a15052a,a15053a,a15057a,a15058a,a15061a,a15064a,a15065a,a15066a,a15070a,a15071a,a15075a,a15076a,a15077a,a15081a,a15082a,a15085a,a15088a,a15089a,a15090a,a15094a,a15095a,a15099a,a15100a,a15101a,a15105a,a15106a,a15109a,a15112a,a15113a,a15114a,a15118a,a15119a,a15123a,a15124a,a15125a,a15129a,a15130a,a15133a,a15136a,a15137a,a15138a,a15142a,a15143a,a15147a,a15148a,a15149a,a15153a,a15154a,a15157a,a15160a,a15161a,a15162a,a15166a,a15167a,a15171a,a15172a,a15173a,a15177a,a15178a,a15181a,a15184a,a15185a,a15186a,a15190a,a15191a,a15195a,a15196a,a15197a,a15201a,a15202a,a15205a,a15208a,a15209a,a15210a,a15214a,a15215a,a15219a,a15220a,a15221a,a15225a,a15226a,a15229a,a15232a,a15233a,a15234a,a15238a,a15239a,a15243a,a15244a,a15245a,a15249a,a15250a,a15253a,a15256a,a15257a,a15258a,a15262a,a15263a,a15267a,a15268a,a15269a,a15273a,a15274a,a15277a,a15280a,a15281a,a15282a,a15286a,a15287a,a15291a,a15292a,a15293a,a15297a,a15298a,a15301a,a15304a,a15305a,a15306a,a15310a,a15311a,a15315a,a15316a,a15317a,a15321a,a15322a,a15325a,a15328a,a15329a,a15330a,a15334a,a15335a,a15339a,a15340a,a15341a,a15345a,a15346a,a15349a,a15352a,a15353a,a15354a,a15358a,a15359a,a15363a,a15364a,a15365a,a15369a,a15370a,a15373a,a15376a,a15377a,a15378a,a15382a,a15383a,a15387a,a15388a,a15389a,a15393a,a15394a,a15397a,a15400a,a15401a,a15402a,a15406a,a15407a,a15411a,a15412a,a15413a,a15417a,a15418a,a15421a,a15424a,a15425a,a15426a,a15430a,a15431a,a15435a,a15436a,a15437a,a15441a,a15442a,a15445a,a15448a,a15449a,a15450a,a15454a,a15455a,a15459a,a15460a,a15461a,a15465a,a15466a,a15469a,a15472a,a15473a,a15474a,a15478a,a15479a,a15483a,a15484a,a15485a,a15489a,a15490a,a15493a,a15496a,a15497a,a15498a,a15502a,a15503a,a15507a,a15508a,a15509a,a15513a,a15514a,a15517a,a15520a,a15521a,a15522a,a15526a,a15527a,a15531a,a15532a,a15533a,a15537a,a15538a,a15541a,a15544a,a15545a,a15546a,a15550a,a15551a,a15555a,a15556a,a15557a,a15561a,a15562a,a15565a,a15568a,a15569a,a15570a,a15574a,a15575a,a15579a,a15580a,a15581a,a15585a,a15586a,a15589a,a15592a,a15593a,a15594a,a15598a,a15599a,a15603a,a15604a,a15605a,a15609a,a15610a,a15613a,a15616a,a15617a,a15618a,a15622a,a15623a,a15627a,a15628a,a15629a,a15633a,a15634a,a15637a,a15640a,a15641a,a15642a,a15646a,a15647a,a15651a,a15652a,a15653a,a15657a,a15658a,a15661a,a15664a,a15665a,a15666a,a15670a,a15671a,a15675a,a15676a,a15677a,a15681a,a15682a,a15685a,a15688a,a15689a,a15690a,a15694a,a15695a,a15699a,a15700a,a15701a,a15705a,a15706a,a15709a,a15712a,a15713a,a15714a,a15718a,a15719a,a15723a,a15724a,a15725a,a15729a,a15730a,a15733a,a15736a,a15737a,a15738a,a15742a,a15743a,a15747a,a15748a,a15749a,a15753a,a15754a,a15757a,a15760a,a15761a,a15762a,a15766a,a15767a,a15771a,a15772a,a15773a,a15777a,a15778a,a15781a,a15784a,a15785a,a15786a,a15790a,a15791a,a15795a,a15796a,a15797a,a15801a,a15802a,a15805a,a15808a,a15809a,a15810a,a15814a,a15815a,a15819a,a15820a,a15821a,a15825a,a15826a,a15829a,a15832a,a15833a,a15834a,a15838a,a15839a,a15843a,a15844a,a15845a,a15849a,a15850a,a15853a,a15856a,a15857a,a15858a,a15862a,a15863a,a15867a,a15868a,a15869a,a15873a,a15874a,a15877a,a15880a,a15881a,a15882a,a15886a,a15887a,a15891a,a15892a,a15893a,a15897a,a15898a,a15901a,a15904a,a15905a,a15906a,a15910a,a15911a,a15915a,a15916a,a15917a,a15921a,a15922a,a15925a,a15928a,a15929a,a15930a,a15934a,a15935a,a15939a,a15940a,a15941a,a15945a,a15946a,a15949a,a15952a,a15953a,a15954a,a15958a,a15959a,a15963a,a15964a,a15965a,a15969a,a15970a,a15973a,a15976a,a15977a,a15978a,a15982a,a15983a,a15987a,a15988a,a15989a,a15993a,a15994a,a15997a,a16000a,a16001a,a16002a,a16006a,a16007a,a16011a,a16012a,a16013a,a16017a,a16018a,a16021a,a16024a,a16025a,a16026a,a16030a,a16031a,a16035a,a16036a,a16037a,a16041a,a16042a,a16045a,a16048a,a16049a,a16050a,a16054a,a16055a,a16059a,a16060a,a16061a,a16065a,a16066a,a16069a,a16072a,a16073a,a16074a,a16078a,a16079a,a16083a,a16084a,a16085a,a16089a,a16090a,a16093a,a16096a,a16097a,a16098a,a16102a,a16103a,a16107a,a16108a,a16109a,a16113a,a16114a,a16117a,a16120a,a16121a,a16122a,a16126a,a16127a,a16131a,a16132a,a16133a,a16137a,a16138a,a16141a,a16144a,a16145a,a16146a,a16150a,a16151a,a16155a,a16156a,a16157a,a16161a,a16162a,a16165a,a16168a,a16169a,a16170a,a16174a,a16175a,a16179a,a16180a,a16181a,a16185a,a16186a,a16189a,a16192a,a16193a,a16194a,a16198a,a16199a,a16203a,a16204a,a16205a,a16209a,a16210a,a16213a,a16216a,a16217a,a16218a,a16222a,a16223a,a16227a,a16228a,a16229a,a16233a,a16234a,a16237a,a16240a,a16241a,a16242a,a16246a,a16247a,a16251a,a16252a,a16253a,a16257a,a16258a,a16261a,a16264a,a16265a,a16266a,a16270a,a16271a,a16275a,a16276a,a16277a,a16281a,a16282a,a16285a,a16288a,a16289a,a16290a,a16294a,a16295a,a16299a,a16300a,a16301a,a16305a,a16306a,a16309a,a16312a,a16313a,a16314a,a16318a,a16319a,a16323a,a16324a,a16325a,a16329a,a16330a,a16333a,a16336a,a16337a,a16338a,a16342a,a16343a,a16347a,a16348a,a16349a,a16353a,a16354a,a16357a,a16360a,a16361a,a16362a,a16366a,a16367a,a16371a,a16372a,a16373a,a16377a,a16378a,a16381a,a16384a,a16385a,a16386a,a16390a,a16391a,a16395a,a16396a,a16397a,a16401a,a16402a,a16405a,a16408a,a16409a,a16410a,a16414a,a16415a,a16419a,a16420a,a16421a,a16425a,a16426a,a16429a,a16432a,a16433a,a16434a,a16438a,a16439a,a16443a,a16444a,a16445a,a16449a,a16450a,a16453a,a16456a,a16457a,a16458a,a16462a,a16463a,a16467a,a16468a,a16469a,a16473a,a16474a,a16477a,a16480a,a16481a,a16482a,a16486a,a16487a,a16491a,a16492a,a16493a,a16497a,a16498a,a16501a,a16504a,a16505a,a16506a,a16510a,a16511a,a16515a,a16516a,a16517a,a16521a,a16522a,a16525a,a16528a,a16529a,a16530a,a16534a,a16535a,a16539a,a16540a,a16541a,a16545a,a16546a,a16549a,a16552a,a16553a,a16554a,a16558a,a16559a,a16563a,a16564a,a16565a,a16569a,a16570a,a16573a,a16576a,a16577a,a16578a,a16582a,a16583a,a16587a,a16588a,a16589a,a16593a,a16594a,a16597a,a16600a,a16601a,a16602a,a16606a,a16607a,a16611a,a16612a,a16613a,a16617a,a16618a,a16621a,a16624a,a16625a,a16626a,a16630a,a16631a,a16635a,a16636a,a16637a,a16641a,a16642a,a16645a,a16648a,a16649a,a16650a,a16654a,a16655a,a16659a,a16660a,a16661a,a16665a,a16666a,a16669a,a16672a,a16673a,a16674a,a16678a,a16679a,a16683a,a16684a,a16685a,a16689a,a16690a,a16693a,a16696a,a16697a,a16698a,a16702a,a16703a,a16707a,a16708a,a16709a,a16713a,a16714a,a16717a,a16720a,a16721a,a16722a,a16726a,a16727a,a16731a,a16732a,a16733a,a16737a,a16738a,a16741a,a16744a,a16745a,a16746a,a16750a,a16751a,a16755a,a16756a,a16757a,a16761a,a16762a,a16765a,a16768a,a16769a,a16770a,a16774a,a16775a,a16779a,a16780a,a16781a,a16785a,a16786a,a16789a,a16792a,a16793a,a16794a,a16798a,a16799a,a16803a,a16804a,a16805a,a16809a,a16810a,a16813a,a16816a,a16817a,a16818a,a16822a,a16823a,a16827a,a16828a,a16829a,a16833a,a16834a,a16837a,a16840a,a16841a,a16842a,a16846a,a16847a,a16851a,a16852a,a16853a,a16857a,a16858a,a16861a,a16864a,a16865a,a16866a,a16870a,a16871a,a16875a,a16876a,a16877a,a16881a,a16882a,a16885a,a16888a,a16889a,a16890a,a16894a,a16895a,a16899a,a16900a,a16901a,a16905a,a16906a,a16909a,a16912a,a16913a,a16914a,a16918a,a16919a,a16923a,a16924a,a16925a,a16929a,a16930a,a16933a,a16936a,a16937a,a16938a,a16942a,a16943a,a16947a,a16948a,a16949a,a16953a,a16954a,a16957a,a16960a,a16961a,a16962a,a16966a,a16967a,a16971a,a16972a,a16973a,a16977a,a16978a,a16981a,a16984a,a16985a,a16986a,a16990a,a16991a,a16995a,a16996a,a16997a,a17001a,a17002a,a17005a,a17008a,a17009a,a17010a,a17014a,a17015a,a17019a,a17020a,a17021a,a17025a,a17026a,a17029a,a17032a,a17033a,a17034a,a17038a,a17039a,a17043a,a17044a,a17045a,a17049a,a17050a,a17053a,a17056a,a17057a,a17058a,a17062a,a17063a,a17067a,a17068a,a17069a,a17073a,a17074a,a17077a,a17080a,a17081a,a17082a,a17086a,a17087a,a17091a,a17092a,a17093a,a17097a,a17098a,a17101a,a17104a,a17105a,a17106a,a17110a,a17111a,a17115a,a17116a,a17117a,a17121a,a17122a,a17125a,a17128a,a17129a,a17130a,a17134a,a17135a,a17139a,a17140a,a17141a,a17145a,a17146a,a17149a,a17152a,a17153a,a17154a,a17158a,a17159a,a17163a,a17164a,a17165a,a17169a,a17170a,a17173a,a17176a,a17177a,a17178a,a17182a,a17183a,a17187a,a17188a,a17189a,a17193a,a17194a,a17197a,a17200a,a17201a,a17202a,a17206a,a17207a,a17211a,a17212a,a17213a,a17217a,a17218a,a17221a,a17224a,a17225a,a17226a,a17230a,a17231a,a17235a,a17236a,a17237a,a17241a,a17242a,a17245a,a17248a,a17249a,a17250a,a17254a,a17255a,a17259a,a17260a,a17261a,a17265a,a17266a,a17269a,a17272a,a17273a,a17274a,a17278a,a17279a,a17283a,a17284a,a17285a,a17289a,a17290a,a17293a,a17296a,a17297a,a17298a,a17302a,a17303a,a17307a,a17308a,a17309a,a17313a,a17314a,a17317a,a17320a,a17321a,a17322a,a17326a,a17327a,a17331a,a17332a,a17333a,a17337a,a17338a,a17341a,a17344a,a17345a,a17346a,a17350a,a17351a,a17355a,a17356a,a17357a,a17361a,a17362a,a17365a,a17368a,a17369a,a17370a,a17374a,a17375a,a17379a,a17380a,a17381a,a17385a,a17386a,a17389a,a17392a,a17393a,a17394a,a17398a,a17399a,a17403a,a17404a,a17405a,a17409a,a17410a,a17413a,a17416a,a17417a,a17418a,a17422a,a17423a,a17427a,a17428a,a17429a,a17433a,a17434a,a17437a,a17440a,a17441a,a17442a,a17446a,a17447a,a17451a,a17452a,a17453a,a17457a,a17458a,a17461a,a17464a,a17465a,a17466a,a17470a,a17471a,a17475a,a17476a,a17477a,a17481a,a17482a,a17485a,a17488a,a17489a,a17490a,a17494a,a17495a,a17499a,a17500a,a17501a,a17505a,a17506a,a17509a,a17512a,a17513a,a17514a,a17518a,a17519a,a17523a,a17524a,a17525a,a17529a,a17530a,a17533a,a17536a,a17537a,a17538a,a17542a,a17543a,a17547a,a17548a,a17549a,a17553a,a17554a,a17557a,a17560a,a17561a,a17562a,a17566a,a17567a,a17571a,a17572a,a17573a,a17577a,a17578a,a17581a,a17584a,a17585a,a17586a,a17590a,a17591a,a17595a,a17596a,a17597a,a17601a,a17602a,a17605a,a17608a,a17609a,a17610a,a17614a,a17615a,a17619a,a17620a,a17621a,a17625a,a17626a,a17629a,a17632a,a17633a,a17634a,a17638a,a17639a,a17643a,a17644a,a17645a,a17649a,a17650a,a17653a,a17656a,a17657a,a17658a,a17662a,a17663a,a17667a,a17668a,a17669a,a17673a,a17674a,a17677a,a17680a,a17681a,a17682a,a17686a,a17687a,a17691a,a17692a,a17693a,a17697a,a17698a,a17701a,a17704a,a17705a,a17706a,a17710a,a17711a,a17715a,a17716a,a17717a,a17721a,a17722a,a17725a,a17728a,a17729a,a17730a,a17734a,a17735a,a17739a,a17740a,a17741a,a17745a,a17746a,a17749a,a17752a,a17753a,a17754a,a17758a,a17759a,a17763a,a17764a,a17765a,a17769a,a17770a,a17773a,a17776a,a17777a,a17778a,a17782a,a17783a,a17787a,a17788a,a17789a,a17793a,a17794a,a17797a,a17800a,a17801a,a17802a,a17806a,a17807a,a17811a,a17812a,a17813a,a17817a,a17818a,a17821a,a17824a,a17825a,a17826a,a17830a,a17831a,a17835a,a17836a,a17837a,a17841a,a17842a,a17845a,a17848a,a17849a,a17850a,a17854a,a17855a,a17859a,a17860a,a17861a,a17865a,a17866a,a17869a,a17872a,a17873a,a17874a,a17878a,a17879a,a17883a,a17884a,a17885a,a17889a,a17890a,a17893a,a17896a,a17897a,a17898a,a17902a,a17903a,a17907a,a17908a,a17909a,a17913a,a17914a,a17917a,a17920a,a17921a,a17922a,a17926a,a17927a,a17931a,a17932a,a17933a,a17937a,a17938a,a17941a,a17944a,a17945a,a17946a,a17950a,a17951a,a17955a,a17956a,a17957a,a17961a,a17962a,a17965a,a17968a,a17969a,a17970a,a17974a,a17975a,a17979a,a17980a,a17981a,a17985a,a17986a,a17989a,a17992a,a17993a,a17994a,a17998a,a17999a,a18003a,a18004a,a18005a,a18009a,a18010a,a18013a,a18016a,a18017a,a18018a,a18022a,a18023a,a18027a,a18028a,a18029a,a18033a,a18034a,a18037a,a18040a,a18041a,a18042a,a18046a,a18047a,a18051a,a18052a,a18053a,a18057a,a18058a,a18061a,a18064a,a18065a,a18066a,a18070a,a18071a,a18075a,a18076a,a18077a,a18081a,a18082a,a18085a,a18088a,a18089a,a18090a,a18094a,a18095a,a18099a,a18100a,a18101a,a18105a,a18106a,a18109a,a18112a,a18113a,a18114a,a18118a,a18119a,a18123a,a18124a,a18125a,a18129a,a18130a,a18133a,a18136a,a18137a,a18138a,a18142a,a18143a,a18147a,a18148a,a18149a,a18153a,a18154a,a18157a,a18160a,a18161a,a18162a,a18166a,a18167a,a18171a,a18172a,a18173a,a18177a,a18178a,a18181a,a18184a,a18185a,a18186a,a18190a,a18191a,a18195a,a18196a,a18197a,a18201a,a18202a,a18205a,a18208a,a18209a,a18210a,a18214a,a18215a,a18219a,a18220a,a18221a,a18225a,a18226a,a18229a,a18232a,a18233a,a18234a,a18238a,a18239a,a18243a,a18244a,a18245a,a18249a,a18250a,a18253a,a18256a,a18257a,a18258a,a18262a,a18263a,a18267a,a18268a,a18269a,a18273a,a18274a,a18277a,a18280a,a18281a,a18282a,a18286a,a18287a,a18291a,a18292a,a18293a,a18297a,a18298a,a18301a,a18304a,a18305a,a18306a,a18310a,a18311a,a18315a,a18316a,a18317a,a18321a,a18322a,a18325a,a18328a,a18329a,a18330a,a18334a,a18335a,a18339a,a18340a,a18341a,a18345a,a18346a,a18349a,a18352a,a18353a,a18354a,a18358a,a18359a,a18363a,a18364a,a18365a,a18369a,a18370a,a18373a,a18376a,a18377a,a18378a,a18382a,a18383a,a18387a,a18388a,a18389a,a18393a,a18394a,a18397a,a18400a,a18401a,a18402a,a18406a,a18407a,a18411a,a18412a,a18413a,a18417a,a18418a,a18421a,a18424a,a18425a,a18426a,a18430a,a18431a,a18435a,a18436a,a18437a,a18441a,a18442a,a18445a,a18448a,a18449a,a18450a,a18454a,a18455a,a18459a,a18460a,a18461a,a18465a,a18466a,a18469a,a18472a,a18473a,a18474a,a18478a,a18479a,a18483a,a18484a,a18485a,a18489a,a18490a,a18493a,a18496a,a18497a,a18498a,a18502a,a18503a,a18507a,a18508a,a18509a,a18513a,a18514a,a18517a,a18520a,a18521a,a18522a,a18526a,a18527a,a18531a,a18532a,a18533a,a18537a,a18538a,a18541a,a18544a,a18545a,a18546a,a18550a,a18551a,a18555a,a18556a,a18557a,a18561a,a18562a,a18565a,a18568a,a18569a,a18570a,a18574a,a18575a,a18579a,a18580a,a18581a,a18585a,a18586a,a18589a,a18592a,a18593a,a18594a,a18598a,a18599a,a18603a,a18604a,a18605a,a18609a,a18610a,a18613a,a18616a,a18617a,a18618a,a18622a,a18623a,a18627a,a18628a,a18629a,a18633a,a18634a,a18637a,a18640a,a18641a,a18642a,a18646a,a18647a,a18651a,a18652a,a18653a,a18657a,a18658a,a18661a,a18664a,a18665a,a18666a,a18670a,a18671a,a18675a,a18676a,a18677a,a18681a,a18682a,a18685a,a18688a,a18689a,a18690a,a18694a,a18695a,a18699a,a18700a,a18701a,a18705a,a18706a,a18709a,a18712a,a18713a,a18714a,a18718a,a18719a,a18723a,a18724a,a18725a,a18729a,a18730a,a18733a,a18736a,a18737a,a18738a,a18742a,a18743a,a18747a,a18748a,a18749a,a18753a,a18754a,a18757a,a18760a,a18761a,a18762a,a18766a,a18767a,a18771a,a18772a,a18773a,a18777a,a18778a,a18781a,a18784a,a18785a,a18786a,a18790a,a18791a,a18795a,a18796a,a18797a,a18801a,a18802a,a18805a,a18808a,a18809a,a18810a,a18814a,a18815a,a18819a,a18820a,a18821a,a18825a,a18826a,a18829a,a18832a,a18833a,a18834a,a18838a,a18839a,a18843a,a18844a,a18845a,a18849a,a18850a,a18853a,a18856a,a18857a,a18858a,a18862a,a18863a,a18867a,a18868a,a18869a,a18873a,a18874a,a18877a,a18880a,a18881a,a18882a,a18886a,a18887a,a18891a,a18892a,a18893a,a18897a,a18898a,a18901a,a18904a,a18905a,a18906a,a18910a,a18911a,a18915a,a18916a,a18917a,a18921a,a18922a,a18925a,a18928a,a18929a,a18930a,a18934a,a18935a,a18939a,a18940a,a18941a,a18945a,a18946a,a18949a,a18952a,a18953a,a18954a,a18958a,a18959a,a18963a,a18964a,a18965a,a18969a,a18970a,a18973a,a18976a,a18977a,a18978a,a18982a,a18983a,a18987a,a18988a,a18989a,a18993a,a18994a,a18997a,a19000a,a19001a,a19002a,a19006a,a19007a,a19011a,a19012a,a19013a,a19017a,a19018a,a19021a,a19024a,a19025a,a19026a,a19030a,a19031a,a19035a,a19036a,a19037a,a19041a,a19042a,a19045a,a19048a,a19049a,a19050a,a19054a,a19055a,a19059a,a19060a,a19061a,a19065a,a19066a,a19069a,a19072a,a19073a,a19074a,a19078a,a19079a,a19083a,a19084a,a19085a,a19089a,a19090a,a19093a,a19096a,a19097a,a19098a,a19102a,a19103a,a19107a,a19108a,a19109a,a19113a,a19114a,a19117a,a19120a,a19121a,a19122a,a19126a,a19127a,a19131a,a19132a,a19133a,a19137a,a19138a,a19141a,a19144a,a19145a,a19146a,a19150a,a19151a,a19155a,a19156a,a19157a,a19161a,a19162a,a19165a,a19168a,a19169a,a19170a,a19174a,a19175a,a19179a,a19180a,a19181a,a19185a,a19186a,a19189a,a19192a,a19193a,a19194a,a19198a,a19199a,a19203a,a19204a,a19205a,a19209a,a19210a,a19213a,a19216a,a19217a,a19218a,a19222a,a19223a,a19227a,a19228a,a19229a,a19233a,a19234a,a19237a,a19240a,a19241a,a19242a,a19246a,a19247a,a19251a,a19252a,a19253a,a19257a,a19258a,a19261a,a19264a,a19265a,a19266a,a19270a,a19271a,a19275a,a19276a,a19277a,a19281a,a19282a,a19285a,a19288a,a19289a,a19290a,a19294a,a19295a,a19299a,a19300a,a19301a,a19305a,a19306a,a19309a,a19312a,a19313a,a19314a,a19318a,a19319a,a19323a,a19324a,a19325a,a19329a,a19330a,a19333a,a19336a,a19337a,a19338a,a19342a,a19343a,a19347a,a19348a,a19349a,a19353a,a19354a,a19357a,a19360a,a19361a,a19362a,a19366a,a19367a,a19371a,a19372a,a19373a,a19377a,a19378a,a19381a,a19384a,a19385a,a19386a,a19390a,a19391a,a19395a,a19396a,a19397a,a19401a,a19402a,a19405a,a19408a,a19409a,a19410a,a19414a,a19415a,a19419a,a19420a,a19421a,a19425a,a19426a,a19429a,a19432a,a19433a,a19434a,a19438a,a19439a,a19443a,a19444a,a19445a,a19449a,a19450a,a19453a,a19456a,a19457a,a19458a,a19462a,a19463a,a19466a,a19469a,a19470a,a19471a,a19475a,a19476a,a19479a,a19482a,a19483a,a19484a,a19488a,a19489a,a19492a,a19495a,a19496a,a19497a,a19501a,a19502a,a19505a,a19508a,a19509a,a19510a,a19514a,a19515a,a19518a,a19521a,a19522a,a19523a,a19527a,a19528a,a19531a,a19534a,a19535a,a19536a,a19540a,a19541a,a19544a,a19547a,a19548a,a19549a,a19553a,a19554a,a19557a,a19560a,a19561a,a19562a,a19566a,a19567a,a19570a,a19573a,a19574a,a19575a,a19579a,a19580a,a19583a,a19586a,a19587a,a19588a,a19592a,a19593a,a19596a,a19599a,a19600a,a19601a,a19605a,a19606a,a19609a,a19612a,a19613a,a19614a,a19618a,a19619a,a19622a,a19625a,a19626a,a19627a,a19631a,a19632a,a19635a,a19638a,a19639a,a19640a,a19644a,a19645a,a19648a,a19651a,a19652a,a19653a,a19657a,a19658a,a19661a,a19664a,a19665a,a19666a,a19670a,a19671a,a19674a,a19677a,a19678a,a19679a,a19683a,a19684a,a19687a,a19690a,a19691a,a19692a,a19696a,a19697a,a19700a,a19703a,a19704a,a19705a,a19709a,a19710a,a19713a,a19716a,a19717a,a19718a,a19722a,a19723a,a19726a,a19729a,a19730a,a19731a,a19735a,a19736a,a19739a,a19742a,a19743a,a19744a,a19748a,a19749a,a19752a,a19755a,a19756a,a19757a,a19761a,a19762a,a19765a,a19768a,a19769a,a19770a,a19774a,a19775a,a19778a,a19781a,a19782a,a19783a,a19787a,a19788a,a19791a,a19794a,a19795a,a19796a,a19800a,a19801a,a19804a,a19807a,a19808a,a19809a,a19813a,a19814a,a19817a,a19820a,a19821a,a19822a,a19826a,a19827a,a19830a,a19833a,a19834a,a19835a,a19839a,a19840a,a19843a,a19846a,a19847a,a19848a,a19852a,a19853a,a19856a,a19859a,a19860a,a19861a,a19865a,a19866a,a19869a,a19872a,a19873a,a19874a,a19878a,a19879a,a19882a,a19885a,a19886a,a19887a,a19891a,a19892a,a19895a,a19898a,a19899a,a19900a,a19904a,a19905a,a19908a,a19911a,a19912a,a19913a,a19917a,a19918a,a19921a,a19924a,a19925a,a19926a,a19930a,a19931a,a19934a,a19937a,a19938a,a19939a,a19943a,a19944a,a19947a,a19950a,a19951a,a19952a,a19956a,a19957a,a19960a,a19963a,a19964a,a19965a,a19969a,a19970a,a19973a,a19976a,a19977a,a19978a,a19982a,a19983a,a19986a,a19989a,a19990a,a19991a,a19995a,a19996a,a19999a,a20002a,a20003a,a20004a,a20008a,a20009a,a20012a,a20015a,a20016a,a20017a,a20021a,a20022a,a20025a,a20028a,a20029a,a20030a,a20034a,a20035a,a20038a,a20041a,a20042a,a20043a,a20047a,a20048a,a20051a,a20054a,a20055a,a20056a,a20060a,a20061a,a20064a,a20067a,a20068a,a20069a,a20073a,a20074a,a20077a,a20080a,a20081a,a20082a,a20086a,a20087a,a20090a,a20093a,a20094a,a20095a,a20099a,a20100a,a20103a,a20106a,a20107a,a20108a,a20112a,a20113a,a20116a,a20119a,a20120a,a20121a,a20125a,a20126a,a20129a,a20132a,a20133a,a20134a,a20138a,a20139a,a20142a,a20145a,a20146a,a20147a,a20151a,a20152a,a20155a,a20158a,a20159a,a20160a,a20164a,a20165a,a20168a,a20171a,a20172a,a20173a,a20177a,a20178a,a20181a,a20184a,a20185a,a20186a,a20190a,a20191a,a20194a,a20197a,a20198a,a20199a,a20203a,a20204a,a20207a,a20210a,a20211a,a20212a,a20216a,a20217a,a20220a,a20223a,a20224a,a20225a,a20229a,a20230a,a20233a,a20236a,a20237a,a20238a,a20242a,a20243a,a20246a,a20249a,a20250a,a20251a,a20255a,a20256a,a20259a,a20262a,a20263a,a20264a,a20268a,a20269a,a20272a,a20275a,a20276a,a20277a,a20281a,a20282a,a20285a,a20288a,a20289a,a20290a,a20294a,a20295a,a20298a,a20301a,a20302a,a20303a,a20307a,a20308a,a20311a,a20314a,a20315a,a20316a,a20320a,a20321a,a20324a,a20327a,a20328a,a20329a,a20333a,a20334a,a20337a,a20340a,a20341a,a20342a,a20346a,a20347a,a20350a,a20353a,a20354a,a20355a,a20359a,a20360a,a20363a,a20366a,a20367a,a20368a,a20372a,a20373a,a20376a,a20379a,a20380a,a20381a,a20385a,a20386a,a20389a,a20392a,a20393a,a20394a,a20398a,a20399a,a20402a,a20405a,a20406a,a20407a,a20411a,a20412a,a20415a,a20418a,a20419a,a20420a,a20424a,a20425a,a20428a,a20431a,a20432a,a20433a,a20437a,a20438a,a20441a,a20444a,a20445a,a20446a,a20450a,a20451a,a20454a,a20457a,a20458a,a20459a,a20463a,a20464a,a20467a,a20470a,a20471a,a20472a,a20476a,a20477a,a20480a,a20483a,a20484a,a20485a,a20489a,a20490a,a20493a,a20496a,a20497a,a20498a,a20502a,a20503a,a20506a,a20509a,a20510a,a20511a,a20515a,a20516a,a20519a,a20522a,a20523a,a20524a,a20528a,a20529a,a20532a,a20535a,a20536a,a20537a,a20541a,a20542a,a20545a,a20548a,a20549a,a20550a,a20554a,a20555a,a20558a,a20561a,a20562a,a20563a,a20567a,a20568a,a20571a,a20574a,a20575a,a20576a,a20580a,a20581a,a20584a,a20587a,a20588a,a20589a,a20593a,a20594a,a20597a,a20600a,a20601a,a20602a,a20606a,a20607a,a20610a,a20613a,a20614a,a20615a,a20619a,a20620a,a20623a,a20626a,a20627a,a20628a,a20632a,a20633a,a20636a,a20639a,a20640a,a20641a,a20645a,a20646a,a20649a,a20652a,a20653a,a20654a,a20658a,a20659a,a20662a,a20665a,a20666a,a20667a,a20671a,a20672a,a20675a,a20678a,a20679a,a20680a,a20684a,a20685a,a20688a,a20691a,a20692a,a20693a,a20697a,a20698a,a20701a,a20704a,a20705a,a20706a,a20710a,a20711a,a20714a,a20717a,a20718a,a20719a,a20723a,a20724a,a20727a,a20730a,a20731a,a20732a,a20736a,a20737a,a20740a,a20743a,a20744a,a20745a,a20749a,a20750a,a20753a,a20756a,a20757a,a20758a,a20762a,a20763a,a20766a,a20769a,a20770a,a20771a,a20775a,a20776a,a20779a,a20782a,a20783a,a20784a,a20788a,a20789a,a20792a,a20795a,a20796a,a20797a,a20801a,a20802a,a20805a,a20808a,a20809a,a20810a,a20814a,a20815a,a20818a,a20821a,a20822a,a20823a,a20827a,a20828a,a20831a,a20834a,a20835a,a20836a,a20840a,a20841a,a20844a,a20847a,a20848a,a20849a,a20853a,a20854a,a20857a,a20860a,a20861a,a20862a,a20866a,a20867a,a20870a,a20873a,a20874a,a20875a,a20879a,a20880a,a20883a,a20886a,a20887a,a20888a,a20892a,a20893a,a20896a,a20899a,a20900a,a20901a,a20905a,a20906a,a20909a,a20912a,a20913a,a20914a,a20918a,a20919a,a20922a,a20925a,a20926a,a20927a,a20931a,a20932a,a20935a,a20938a,a20939a,a20940a,a20944a,a20945a,a20948a,a20951a,a20952a,a20953a,a20957a,a20958a,a20961a,a20964a,a20965a,a20966a,a20970a,a20971a,a20974a,a20977a,a20978a,a20979a,a20983a,a20984a,a20987a,a20990a,a20991a,a20992a,a20996a,a20997a,a21000a,a21003a,a21004a,a21005a,a21009a,a21010a,a21013a,a21016a,a21017a,a21018a,a21022a,a21023a,a21026a,a21029a,a21030a,a21031a,a21035a,a21036a,a21039a,a21042a,a21043a,a21044a,a21048a,a21049a,a21052a,a21055a,a21056a,a21057a,a21061a,a21062a,a21065a,a21068a,a21069a,a21070a,a21074a,a21075a,a21078a,a21081a,a21082a,a21083a,a21087a,a21088a,a21091a,a21094a,a21095a,a21096a,a21100a,a21101a,a21104a,a21107a,a21108a,a21109a,a21113a,a21114a,a21117a,a21120a,a21121a,a21122a,a21126a,a21127a,a21130a,a21133a,a21134a,a21135a,a21139a,a21140a,a21143a,a21146a,a21147a,a21148a,a21152a,a21153a,a21156a,a21159a,a21160a,a21161a,a21165a,a21166a,a21169a,a21172a,a21173a,a21174a,a21178a,a21179a,a21182a,a21185a,a21186a,a21187a,a21191a,a21192a,a21195a,a21198a,a21199a,a21200a,a21204a,a21205a,a21208a,a21211a,a21212a,a21213a,a21217a,a21218a,a21221a,a21224a,a21225a,a21226a,a21230a,a21231a,a21234a,a21237a,a21238a,a21239a,a21243a,a21244a,a21247a,a21250a,a21251a,a21252a,a21256a,a21257a,a21260a,a21263a,a21264a,a21265a,a21269a,a21270a,a21273a,a21276a,a21277a,a21278a,a21282a,a21283a,a21286a,a21289a,a21290a,a21291a,a21295a,a21296a,a21299a,a21302a,a21303a,a21304a,a21308a,a21309a,a21312a,a21315a,a21316a,a21317a,a21321a,a21322a,a21325a,a21328a,a21329a,a21330a,a21334a,a21335a,a21338a,a21341a,a21342a,a21343a,a21347a,a21348a,a21351a,a21354a,a21355a,a21356a,a21360a,a21361a,a21364a,a21367a,a21368a,a21369a,a21373a,a21374a,a21377a,a21380a,a21381a,a21382a,a21386a,a21387a,a21390a,a21393a,a21394a,a21395a,a21399a,a21400a,a21403a,a21406a,a21407a,a21408a,a21412a,a21413a,a21416a,a21419a,a21420a,a21421a,a21425a,a21426a,a21429a,a21432a,a21433a,a21434a,a21438a,a21439a,a21442a,a21445a,a21446a,a21447a,a21451a,a21452a,a21455a,a21458a,a21459a,a21460a,a21464a,a21465a,a21468a,a21471a,a21472a,a21473a,a21477a,a21478a,a21481a,a21484a,a21485a,a21486a,a21490a,a21491a,a21494a,a21497a,a21498a,a21499a,a21503a,a21504a,a21507a,a21510a,a21511a,a21512a,a21516a,a21517a,a21520a,a21523a,a21524a,a21525a,a21529a,a21530a,a21533a,a21536a,a21537a,a21538a,a21542a,a21543a,a21546a,a21549a,a21550a,a21551a,a21555a,a21556a,a21559a,a21562a,a21563a,a21564a,a21568a,a21569a,a21572a,a21575a,a21576a,a21577a,a21581a,a21582a,a21585a,a21588a,a21589a,a21590a,a21594a,a21595a,a21598a,a21601a,a21602a,a21603a,a21607a,a21608a,a21611a,a21614a,a21615a,a21616a,a21620a,a21621a,a21624a,a21627a,a21628a,a21629a,a21633a,a21634a,a21637a,a21640a,a21641a,a21642a,a21646a,a21647a,a21650a,a21653a,a21654a,a21655a,a21659a,a21660a,a21663a,a21666a,a21667a,a21668a,a21672a,a21673a,a21676a,a21679a,a21680a,a21681a,a21685a,a21686a,a21689a,a21692a,a21693a,a21694a,a21698a,a21699a,a21702a,a21705a,a21706a,a21707a,a21711a,a21712a,a21715a,a21718a,a21719a,a21720a,a21724a,a21725a,a21728a,a21731a,a21732a,a21733a,a21737a,a21738a,a21741a,a21744a,a21745a,a21746a,a21750a,a21751a,a21754a,a21757a,a21758a,a21759a,a21763a,a21764a,a21767a,a21770a,a21771a,a21772a,a21776a,a21777a,a21780a,a21783a,a21784a,a21785a,a21789a,a21790a,a21793a,a21796a,a21797a,a21798a,a21802a,a21803a,a21806a,a21809a,a21810a,a21811a,a21815a,a21816a,a21819a,a21822a,a21823a,a21824a,a21828a,a21829a,a21832a,a21835a,a21836a,a21837a,a21841a,a21842a,a21845a,a21848a,a21849a,a21850a,a21854a,a21855a,a21858a,a21861a,a21862a,a21863a,a21867a,a21868a,a21871a,a21874a,a21875a,a21876a,a21880a,a21881a,a21884a,a21887a,a21888a,a21889a,a21893a,a21894a,a21897a,a21900a,a21901a,a21902a,a21906a,a21907a,a21910a,a21913a,a21914a,a21915a,a21919a,a21920a,a21923a,a21926a,a21927a,a21928a,a21932a,a21933a,a21936a,a21939a,a21940a,a21941a,a21945a,a21946a,a21949a,a21952a,a21953a,a21954a,a21958a,a21959a,a21962a,a21965a,a21966a,a21967a,a21971a,a21972a,a21975a,a21978a,a21979a,a21980a,a21984a,a21985a,a21988a,a21991a,a21992a,a21993a,a21997a,a21998a,a22001a,a22004a,a22005a,a22006a,a22010a,a22011a,a22014a,a22017a,a22018a,a22019a,a22023a,a22024a,a22027a,a22030a,a22031a,a22032a,a22036a,a22037a,a22040a,a22043a,a22044a,a22045a,a22049a,a22050a,a22053a,a22056a,a22057a,a22058a,a22062a,a22063a,a22066a,a22069a,a22070a,a22071a,a22075a,a22076a,a22079a,a22082a,a22083a,a22084a,a22088a,a22089a,a22092a,a22095a,a22096a,a22097a,a22101a,a22102a,a22105a,a22108a,a22109a,a22110a,a22114a,a22115a,a22118a,a22121a,a22122a,a22123a,a22127a,a22128a,a22131a,a22134a,a22135a,a22136a,a22140a,a22141a,a22144a,a22147a,a22148a,a22149a,a22153a,a22154a,a22157a,a22160a,a22161a,a22162a,a22166a,a22167a,a22170a,a22173a,a22174a,a22175a,a22179a,a22180a,a22183a,a22186a,a22187a,a22188a,a22192a,a22193a,a22196a,a22199a,a22200a,a22201a,a22205a,a22206a,a22209a,a22212a,a22213a,a22214a,a22218a,a22219a,a22222a,a22225a,a22226a,a22227a,a22231a,a22232a,a22235a,a22238a,a22239a,a22240a,a22244a,a22245a,a22248a,a22251a,a22252a,a22253a,a22257a,a22258a,a22261a,a22264a,a22265a,a22266a,a22270a,a22271a,a22274a,a22277a,a22278a,a22279a,a22283a,a22284a,a22287a,a22290a,a22291a,a22292a,a22296a,a22297a,a22300a,a22303a,a22304a,a22305a,a22309a,a22310a,a22313a,a22316a,a22317a,a22318a,a22322a,a22323a,a22326a,a22329a,a22330a,a22331a,a22335a,a22336a,a22339a,a22342a,a22343a,a22344a,a22348a,a22349a,a22352a,a22355a,a22356a,a22357a,a22361a,a22362a,a22365a,a22368a,a22369a,a22370a,a22374a,a22375a,a22378a,a22381a,a22382a,a22383a,a22387a,a22388a,a22391a,a22394a,a22395a,a22396a,a22400a,a22401a,a22404a,a22407a,a22408a,a22409a,a22413a,a22414a,a22417a,a22420a,a22421a,a22422a,a22426a,a22427a,a22430a,a22433a,a22434a,a22435a,a22439a,a22440a,a22443a,a22446a,a22447a,a22448a,a22452a,a22453a,a22456a,a22459a,a22460a,a22461a,a22465a,a22466a,a22469a,a22472a,a22473a,a22474a,a22478a,a22479a,a22482a,a22485a,a22486a,a22487a,a22491a,a22492a,a22495a,a22498a,a22499a,a22500a,a22504a,a22505a,a22508a,a22511a,a22512a,a22513a,a22517a,a22518a,a22521a,a22524a,a22525a,a22526a,a22530a,a22531a,a22534a,a22537a,a22538a,a22539a,a22543a,a22544a,a22547a,a22550a,a22551a,a22552a,a22556a,a22557a,a22560a,a22563a,a22564a,a22565a,a22569a,a22570a,a22573a,a22576a,a22577a,a22578a,a22582a,a22583a,a22586a,a22589a,a22590a,a22591a,a22595a,a22596a,a22599a,a22602a,a22603a,a22604a,a22608a,a22609a,a22612a,a22615a,a22616a,a22617a,a22621a,a22622a,a22625a,a22628a,a22629a,a22630a,a22634a,a22635a,a22638a,a22641a,a22642a,a22643a,a22647a,a22648a,a22651a,a22654a,a22655a,a22656a,a22660a,a22661a,a22664a,a22667a,a22668a,a22669a,a22673a,a22674a,a22677a,a22680a,a22681a,a22682a,a22686a,a22687a,a22690a,a22693a,a22694a,a22695a,a22699a,a22700a,a22703a,a22706a,a22707a,a22708a,a22712a,a22713a,a22716a,a22719a,a22720a,a22721a,a22725a,a22726a,a22729a,a22732a,a22733a,a22734a,a22738a,a22739a,a22742a,a22745a,a22746a,a22747a,a22751a,a22752a,a22755a,a22758a,a22759a,a22760a,a22764a,a22765a,a22768a,a22771a,a22772a,a22773a,a22777a,a22778a,a22781a,a22784a,a22785a,a22786a,a22790a,a22791a,a22794a,a22797a,a22798a,a22799a,a22803a,a22804a,a22807a,a22810a,a22811a,a22812a,a22816a,a22817a,a22820a,a22823a,a22824a,a22825a,a22829a,a22830a,a22833a,a22836a,a22837a,a22838a,a22842a,a22843a,a22846a,a22849a,a22850a,a22851a,a22855a,a22856a,a22859a,a22862a,a22863a,a22864a,a22868a,a22869a,a22872a,a22875a,a22876a,a22877a,a22881a,a22882a,a22885a,a22888a,a22889a,a22890a,a22894a,a22895a,a22898a,a22901a,a22902a,a22903a,a22907a,a22908a,a22911a,a22914a,a22915a,a22916a,a22920a,a22921a,a22924a,a22927a,a22928a,a22929a,a22933a,a22934a,a22937a,a22940a,a22941a,a22942a,a22946a,a22947a,a22950a,a22953a,a22954a,a22955a,a22959a,a22960a,a22963a,a22966a,a22967a,a22968a,a22972a,a22973a,a22976a,a22979a,a22980a,a22981a,a22985a,a22986a,a22989a,a22992a,a22993a,a22994a,a22998a,a22999a,a23002a,a23005a,a23006a,a23007a,a23011a,a23012a,a23015a,a23018a,a23019a,a23020a,a23024a,a23025a,a23028a,a23031a,a23032a,a23033a,a23037a,a23038a,a23041a,a23044a,a23045a,a23046a,a23050a,a23051a,a23054a,a23057a,a23058a,a23059a,a23063a,a23064a,a23067a,a23070a,a23071a,a23072a,a23076a,a23077a,a23080a,a23083a,a23084a,a23085a,a23089a,a23090a,a23093a,a23096a,a23097a,a23098a,a23102a,a23103a,a23106a,a23109a,a23110a,a23111a,a23115a,a23116a,a23119a,a23122a,a23123a,a23124a,a23128a,a23129a,a23132a,a23135a,a23136a,a23137a,a23141a,a23142a,a23145a,a23148a,a23149a,a23150a,a23154a,a23155a,a23158a,a23161a,a23162a,a23163a,a23167a,a23168a,a23171a,a23174a,a23175a,a23176a,a23180a,a23181a,a23184a,a23187a,a23188a,a23189a,a23193a,a23194a,a23197a,a23200a,a23201a,a23202a,a23206a,a23207a,a23210a,a23213a,a23214a,a23215a,a23219a,a23220a,a23223a,a23226a,a23227a,a23228a,a23232a,a23233a,a23236a,a23239a,a23240a,a23241a,a23245a,a23246a,a23249a,a23252a,a23253a,a23254a,a23258a,a23259a,a23262a,a23265a,a23266a,a23267a,a23271a,a23272a,a23275a,a23278a,a23279a,a23280a,a23284a,a23285a,a23288a,a23291a,a23292a,a23293a,a23297a,a23298a,a23301a,a23304a,a23305a,a23306a,a23310a,a23311a,a23314a,a23317a,a23318a,a23319a,a23323a,a23324a,a23327a,a23330a,a23331a,a23332a,a23336a,a23337a,a23340a,a23343a,a23344a,a23345a,a23349a,a23350a,a23353a,a23356a,a23357a,a23358a,a23362a,a23363a,a23366a,a23369a,a23370a,a23371a,a23375a,a23376a,a23379a,a23382a,a23383a,a23384a,a23388a,a23389a,a23392a,a23395a,a23396a,a23397a,a23401a,a23402a,a23405a,a23408a,a23409a,a23410a,a23414a,a23415a,a23418a,a23421a,a23422a,a23423a,a23427a,a23428a,a23431a,a23434a,a23435a,a23436a,a23440a,a23441a,a23444a,a23447a,a23448a,a23449a,a23453a,a23454a,a23457a,a23460a,a23461a,a23462a,a23466a,a23467a,a23470a,a23473a,a23474a,a23475a,a23479a,a23480a,a23483a,a23486a,a23487a,a23488a,a23492a,a23493a,a23496a,a23499a,a23500a,a23501a,a23505a,a23506a,a23509a,a23512a,a23513a,a23514a,a23518a,a23519a,a23522a,a23525a,a23526a,a23527a,a23531a,a23532a,a23535a,a23538a,a23539a,a23540a,a23544a,a23545a,a23548a,a23551a,a23552a,a23553a,a23557a,a23558a,a23561a,a23564a,a23565a,a23566a,a23570a,a23571a,a23574a,a23577a,a23578a,a23579a,a23583a,a23584a,a23587a,a23590a,a23591a,a23592a,a23596a,a23597a,a23600a,a23603a,a23604a,a23605a,a23609a,a23610a,a23613a,a23616a,a23617a,a23618a,a23622a,a23623a,a23626a,a23629a,a23630a,a23631a,a23635a,a23636a,a23639a,a23642a,a23643a,a23644a,a23648a,a23649a,a23652a,a23655a,a23656a,a23657a,a23661a,a23662a,a23665a,a23668a,a23669a,a23670a,a23674a,a23675a,a23678a,a23681a,a23682a,a23683a,a23687a,a23688a,a23691a,a23694a,a23695a,a23696a,a23700a,a23701a,a23704a,a23707a,a23708a,a23709a,a23713a,a23714a,a23717a,a23720a,a23721a,a23722a,a23726a,a23727a,a23730a,a23733a,a23734a,a23735a,a23739a,a23740a,a23743a,a23746a,a23747a,a23748a,a23752a,a23753a,a23756a,a23759a,a23760a,a23761a,a23765a,a23766a,a23769a,a23772a,a23773a,a23774a,a23778a,a23779a,a23782a,a23785a,a23786a,a23787a,a23791a,a23792a,a23795a,a23798a,a23799a,a23800a,a23804a,a23805a,a23808a,a23811a,a23812a,a23813a,a23817a,a23818a,a23821a,a23824a,a23825a,a23826a,a23830a,a23831a,a23834a,a23837a,a23838a,a23839a,a23843a,a23844a,a23847a,a23850a,a23851a,a23852a,a23856a,a23857a,a23860a,a23863a,a23864a,a23865a,a23869a,a23870a,a23873a,a23876a,a23877a,a23878a,a23882a,a23883a,a23886a,a23889a,a23890a,a23891a,a23895a,a23896a,a23899a,a23902a,a23903a,a23904a,a23908a,a23909a,a23912a,a23915a,a23916a,a23917a,a23921a,a23922a,a23925a,a23928a,a23929a,a23930a,a23934a,a23935a,a23938a,a23941a,a23942a,a23943a,a23947a,a23948a,a23951a,a23954a,a23955a,a23956a,a23960a,a23961a,a23964a,a23967a,a23968a,a23969a,a23973a,a23974a,a23977a,a23980a,a23981a,a23982a,a23986a,a23987a,a23990a,a23993a,a23994a,a23995a,a23999a,a24000a,a24003a,a24006a,a24007a,a24008a,a24012a,a24013a,a24016a,a24019a,a24020a,a24021a,a24025a,a24026a,a24029a,a24032a,a24033a,a24034a,a24038a,a24039a,a24042a,a24045a,a24046a,a24047a,a24051a,a24052a,a24055a,a24058a,a24059a,a24060a,a24064a,a24065a,a24068a,a24071a,a24072a,a24073a,a24077a,a24078a,a24081a,a24084a,a24085a,a24086a,a24090a,a24091a,a24094a,a24097a,a24098a,a24099a,a24103a,a24104a,a24107a,a24110a,a24111a,a24112a,a24116a,a24117a,a24120a,a24123a,a24124a,a24125a,a24129a,a24130a,a24133a,a24136a,a24137a,a24138a,a24142a,a24143a,a24146a,a24149a,a24150a,a24151a,a24155a,a24156a,a24159a,a24162a,a24163a,a24164a,a24168a,a24169a,a24172a,a24175a,a24176a,a24177a,a24181a,a24182a,a24185a,a24188a,a24189a,a24190a,a24194a,a24195a,a24198a,a24201a,a24202a,a24203a,a24207a,a24208a,a24211a,a24214a,a24215a,a24216a,a24220a,a24221a,a24224a,a24227a,a24228a,a24229a,a24233a,a24234a,a24237a,a24240a,a24241a,a24242a,a24246a,a24247a,a24250a,a24253a,a24254a,a24255a,a24259a,a24260a,a24263a,a24266a,a24267a,a24268a,a24272a,a24273a,a24276a,a24279a,a24280a,a24281a,a24285a,a24286a,a24289a,a24292a,a24293a,a24294a,a24298a,a24299a,a24302a,a24305a,a24306a,a24307a,a24311a,a24312a,a24315a,a24318a,a24319a,a24320a,a24324a,a24325a,a24328a,a24331a,a24332a,a24333a,a24337a,a24338a,a24341a,a24344a,a24345a,a24346a,a24350a,a24351a,a24354a,a24357a,a24358a,a24359a,a24363a,a24364a,a24367a,a24370a,a24371a,a24372a,a24376a,a24377a,a24380a,a24383a,a24384a,a24385a,a24389a,a24390a,a24393a,a24396a,a24397a,a24398a,a24402a,a24403a,a24406a,a24409a,a24410a,a24411a,a24415a,a24416a,a24419a,a24422a,a24423a,a24424a,a24428a,a24429a,a24432a,a24435a,a24436a,a24437a,a24441a,a24442a,a24445a,a24448a,a24449a,a24450a,a24454a,a24455a,a24458a,a24461a,a24462a,a24463a,a24467a,a24468a,a24471a,a24474a,a24475a,a24476a,a24480a,a24481a,a24484a,a24487a,a24488a,a24489a,a24493a,a24494a,a24497a,a24500a,a24501a,a24502a,a24506a,a24507a,a24510a,a24513a,a24514a,a24515a,a24519a,a24520a,a24523a,a24526a,a24527a,a24528a,a24532a,a24533a,a24536a,a24539a,a24540a,a24541a,a24545a,a24546a,a24549a,a24552a,a24553a,a24554a,a24558a,a24559a,a24562a,a24565a,a24566a,a24567a,a24571a,a24572a,a24575a,a24578a,a24579a,a24580a,a24584a,a24585a,a24588a,a24591a,a24592a,a24593a,a24597a,a24598a,a24601a,a24604a,a24605a,a24606a,a24610a,a24611a,a24614a,a24617a,a24618a,a24619a,a24623a,a24624a,a24627a,a24630a,a24631a,a24632a,a24636a,a24637a,a24640a,a24643a,a24644a,a24645a,a24649a,a24650a,a24653a,a24656a,a24657a,a24658a,a24662a,a24663a,a24666a,a24669a,a24670a,a24671a,a24675a,a24676a,a24679a,a24682a,a24683a,a24684a,a24688a,a24689a,a24692a,a24695a,a24696a,a24697a,a24701a,a24702a,a24705a,a24708a,a24709a,a24710a,a24714a,a24715a,a24718a,a24721a,a24722a,a24723a,a24727a,a24728a,a24731a,a24734a,a24735a,a24736a,a24740a,a24741a,a24744a,a24747a,a24748a,a24749a,a24753a,a24754a,a24757a,a24760a,a24761a,a24762a,a24766a,a24767a,a24770a,a24773a,a24774a,a24775a,a24779a,a24780a,a24783a,a24786a,a24787a,a24788a,a24792a,a24793a,a24796a,a24799a,a24800a,a24801a,a24805a,a24806a,a24809a,a24812a,a24813a,a24814a,a24818a,a24819a,a24822a,a24825a,a24826a,a24827a,a24831a,a24832a,a24835a,a24838a,a24839a,a24840a,a24844a,a24845a,a24848a,a24851a,a24852a,a24853a,a24857a,a24858a,a24861a,a24864a,a24865a,a24866a,a24870a,a24871a,a24874a,a24877a,a24878a,a24879a,a24883a,a24884a,a24887a,a24890a,a24891a,a24892a,a24896a,a24897a,a24900a,a24903a,a24904a,a24905a,a24909a,a24910a,a24913a,a24916a,a24917a,a24918a,a24922a,a24923a,a24926a,a24929a,a24930a,a24931a,a24935a,a24936a,a24939a,a24942a,a24943a,a24944a,a24948a,a24949a,a24952a,a24955a,a24956a,a24957a,a24961a,a24962a,a24965a,a24968a,a24969a,a24970a,a24974a,a24975a,a24978a,a24981a,a24982a,a24983a,a24987a,a24988a,a24991a,a24994a,a24995a,a24996a,a25000a,a25001a,a25004a,a25007a,a25008a,a25009a,a25013a,a25014a,a25017a,a25020a,a25021a,a25022a,a25026a,a25027a,a25030a,a25033a,a25034a,a25035a,a25039a,a25040a,a25043a,a25046a,a25047a,a25048a,a25052a,a25053a,a25056a,a25059a,a25060a,a25061a,a25065a,a25066a,a25069a,a25072a,a25073a,a25074a,a25078a,a25079a,a25082a,a25085a,a25086a,a25087a,a25091a,a25092a,a25095a,a25098a,a25099a,a25100a,a25104a,a25105a,a25108a,a25111a,a25112a,a25113a,a25117a,a25118a,a25121a,a25124a,a25125a,a25126a,a25130a,a25131a,a25134a,a25137a,a25138a,a25139a,a25143a,a25144a,a25147a,a25150a,a25151a,a25152a,a25156a,a25157a,a25160a,a25163a,a25164a,a25165a,a25169a,a25170a,a25173a,a25176a,a25177a,a25178a,a25182a,a25183a,a25186a,a25189a,a25190a,a25191a,a25195a,a25196a,a25199a,a25202a,a25203a,a25204a,a25208a,a25209a,a25212a,a25215a,a25216a,a25217a,a25221a,a25222a,a25225a,a25228a,a25229a,a25230a,a25234a,a25235a,a25238a,a25241a,a25242a,a25243a,a25247a,a25248a,a25251a,a25254a,a25255a,a25256a,a25260a,a25261a,a25264a,a25267a,a25268a,a25269a,a25273a,a25274a,a25277a,a25280a,a25281a,a25282a,a25286a,a25287a,a25290a,a25293a,a25294a,a25295a,a25299a,a25300a,a25303a,a25306a,a25307a,a25308a,a25312a,a25313a,a25316a,a25319a,a25320a,a25321a,a25325a,a25326a,a25329a,a25332a,a25333a,a25334a,a25338a,a25339a,a25342a,a25345a,a25346a,a25347a,a25351a,a25352a,a25355a,a25358a,a25359a,a25360a,a25364a,a25365a,a25368a,a25371a,a25372a,a25373a,a25377a,a25378a,a25381a,a25384a,a25385a,a25386a,a25390a,a25391a,a25394a,a25397a,a25398a,a25399a,a25403a,a25404a,a25407a,a25410a,a25411a,a25412a,a25416a,a25417a,a25420a,a25423a,a25424a,a25425a,a25429a,a25430a,a25433a,a25436a,a25437a,a25438a,a25442a,a25443a,a25446a,a25449a,a25450a,a25451a,a25455a,a25456a,a25459a,a25462a,a25463a,a25464a,a25468a,a25469a,a25472a,a25475a,a25476a,a25477a,a25481a,a25482a,a25485a,a25488a,a25489a,a25490a,a25494a,a25495a,a25498a,a25501a,a25502a,a25503a,a25507a,a25508a,a25511a,a25514a,a25515a,a25516a,a25520a,a25521a,a25524a,a25527a,a25528a,a25529a,a25533a,a25534a,a25537a,a25540a,a25541a,a25542a,a25546a,a25547a,a25550a,a25553a,a25554a,a25555a,a25559a,a25560a,a25563a,a25566a,a25567a,a25568a,a25572a,a25573a,a25576a,a25579a,a25580a,a25581a,a25585a,a25586a,a25589a,a25592a,a25593a,a25594a,a25598a,a25599a,a25602a,a25605a,a25606a,a25607a,a25611a,a25612a,a25615a,a25618a,a25619a,a25620a,a25624a,a25625a,a25628a,a25631a,a25632a,a25633a,a25637a,a25638a,a25641a,a25644a,a25645a,a25646a,a25650a,a25651a,a25654a,a25657a,a25658a,a25659a,a25663a,a25664a,a25667a,a25670a,a25671a,a25672a,a25676a,a25677a,a25680a,a25683a,a25684a,a25685a,a25689a,a25690a,a25693a,a25696a,a25697a,a25698a,a25702a,a25703a,a25706a,a25709a,a25710a,a25711a,a25715a,a25716a,a25719a,a25722a,a25723a,a25724a,a25728a,a25729a,a25732a,a25735a,a25736a,a25737a,a25741a,a25742a,a25745a,a25748a,a25749a,a25750a,a25754a,a25755a,a25758a,a25761a,a25762a,a25763a,a25767a,a25768a,a25771a,a25774a,a25775a,a25776a,a25780a,a25781a,a25784a,a25787a,a25788a,a25789a,a25793a,a25794a,a25797a,a25800a,a25801a,a25802a,a25806a,a25807a,a25810a,a25813a,a25814a,a25815a,a25819a,a25820a,a25823a,a25826a,a25827a,a25828a,a25832a,a25833a,a25836a,a25839a,a25840a,a25841a,a25845a,a25846a,a25849a,a25852a,a25853a,a25854a,a25858a,a25859a,a25862a,a25865a,a25866a,a25867a,a25871a,a25872a,a25875a,a25878a,a25879a,a25880a,a25884a,a25885a,a25888a,a25891a,a25892a,a25893a,a25897a,a25898a,a25901a,a25904a,a25905a,a25906a,a25910a,a25911a,a25914a,a25917a,a25918a,a25919a,a25923a,a25924a,a25927a,a25930a,a25931a,a25932a,a25936a,a25937a,a25940a,a25943a,a25944a,a25945a,a25949a,a25950a,a25953a,a25956a,a25957a,a25958a,a25962a,a25963a,a25966a,a25969a,a25970a,a25971a,a25975a,a25976a,a25979a,a25982a,a25983a,a25984a,a25988a,a25989a,a25992a,a25995a,a25996a,a25997a,a26001a,a26002a,a26005a,a26008a,a26009a,a26010a,a26014a,a26015a,a26018a,a26021a,a26022a,a26023a,a26027a,a26028a,a26031a,a26034a,a26035a,a26036a,a26040a,a26041a,a26044a,a26047a,a26048a,a26049a,a26053a,a26054a,a26057a,a26060a,a26061a,a26062a,a26066a,a26067a,a26070a,a26073a,a26074a,a26075a,a26079a,a26080a,a26083a,a26086a,a26087a,a26088a,a26092a,a26093a,a26096a,a26099a,a26100a,a26101a,a26105a,a26106a,a26109a,a26112a,a26113a,a26114a,a26118a,a26119a,a26122a,a26125a,a26126a,a26127a,a26131a,a26132a,a26135a,a26138a,a26139a,a26140a,a26144a,a26145a,a26148a,a26151a,a26152a,a26153a,a26157a,a26158a,a26161a,a26164a,a26165a,a26166a,a26170a,a26171a,a26174a,a26177a,a26178a,a26179a,a26183a,a26184a,a26187a,a26190a,a26191a,a26192a,a26196a,a26197a,a26200a,a26203a,a26204a,a26205a,a26209a,a26210a,a26213a,a26216a,a26217a,a26218a,a26222a,a26223a,a26226a,a26229a,a26230a,a26231a,a26235a,a26236a,a26239a,a26242a,a26243a,a26244a,a26248a,a26249a,a26252a,a26255a,a26256a,a26257a,a26261a,a26262a,a26265a,a26268a,a26269a,a26270a,a26274a,a26275a,a26278a,a26281a,a26282a,a26283a,a26287a,a26288a,a26291a,a26294a,a26295a,a26296a,a26300a,a26301a,a26304a,a26307a,a26308a,a26309a,a26313a,a26314a,a26317a,a26320a,a26321a,a26322a,a26326a,a26327a,a26330a,a26333a,a26334a,a26335a,a26339a,a26340a,a26343a,a26346a,a26347a,a26348a,a26352a,a26353a,a26356a,a26359a,a26360a,a26361a,a26365a,a26366a,a26369a,a26372a,a26373a,a26374a,a26378a,a26379a,a26382a,a26385a,a26386a,a26387a,a26391a,a26392a,a26395a,a26398a,a26399a,a26400a,a26404a,a26405a,a26408a,a26411a,a26412a,a26413a,a26417a,a26418a,a26421a,a26424a,a26425a,a26426a,a26430a,a26431a,a26434a,a26437a,a26438a,a26439a,a26443a,a26444a,a26447a,a26450a,a26451a,a26452a,a26456a,a26457a,a26460a,a26463a,a26464a,a26465a,a26469a,a26470a,a26473a,a26476a,a26477a,a26478a,a26482a,a26483a,a26486a,a26489a,a26490a,a26491a,a26495a,a26496a,a26499a,a26502a,a26503a,a26504a,a26508a,a26509a,a26512a,a26515a,a26516a,a26517a,a26521a,a26522a,a26525a,a26528a,a26529a,a26530a,a26534a,a26535a,a26538a,a26541a,a26542a,a26543a,a26547a,a26548a,a26551a,a26554a,a26555a,a26556a,a26560a,a26561a,a26564a,a26567a,a26568a,a26569a,a26573a,a26574a,a26577a,a26580a,a26581a,a26582a,a26586a,a26587a,a26590a,a26593a,a26594a,a26595a,a26599a,a26600a,a26603a,a26606a,a26607a,a26608a,a26612a,a26613a,a26616a,a26619a,a26620a,a26621a,a26625a,a26626a,a26629a,a26632a,a26633a,a26634a,a26638a,a26639a,a26642a,a26645a,a26646a,a26647a,a26651a,a26652a,a26655a,a26658a,a26659a,a26660a,a26664a,a26665a,a26668a,a26671a,a26672a,a26673a,a26677a,a26678a,a26681a,a26684a,a26685a,a26686a,a26690a,a26691a,a26694a,a26697a,a26698a,a26699a,a26703a,a26704a,a26707a,a26710a,a26711a,a26712a,a26716a,a26717a,a26720a,a26723a,a26724a,a26725a,a26729a,a26730a,a26733a,a26736a,a26737a,a26738a,a26742a,a26743a,a26746a,a26749a,a26750a,a26751a,a26755a,a26756a,a26759a,a26762a,a26763a,a26764a,a26768a,a26769a,a26772a,a26775a,a26776a,a26777a,a26781a,a26782a,a26785a,a26788a,a26789a,a26790a,a26794a,a26795a,a26798a,a26801a,a26802a,a26803a,a26807a,a26808a,a26811a,a26814a,a26815a,a26816a,a26820a,a26821a,a26824a,a26827a,a26828a,a26829a,a26833a,a26834a,a26837a,a26840a,a26841a,a26842a,a26846a,a26847a,a26850a,a26853a,a26854a,a26855a,a26859a,a26860a,a26863a,a26866a,a26867a,a26868a,a26872a,a26873a,a26876a,a26879a,a26880a,a26881a,a26885a,a26886a,a26889a,a26892a,a26893a,a26894a,a26898a,a26899a,a26902a,a26905a,a26906a,a26907a,a26911a,a26912a,a26915a,a26918a,a26919a,a26920a,a26924a,a26925a,a26928a,a26931a,a26932a,a26933a,a26937a,a26938a,a26941a,a26944a,a26945a,a26946a,a26950a,a26951a,a26954a,a26957a,a26958a,a26959a,a26963a,a26964a,a26967a,a26970a,a26971a,a26972a,a26976a,a26977a,a26980a,a26983a,a26984a,a26985a,a26989a,a26990a,a26993a,a26996a,a26997a,a26998a,a27002a,a27003a,a27006a,a27009a,a27010a,a27011a,a27015a,a27016a,a27019a,a27022a,a27023a,a27024a,a27028a,a27029a,a27032a,a27035a,a27036a,a27037a,a27041a,a27042a,a27045a,a27048a,a27049a,a27050a,a27054a,a27055a,a27058a,a27061a,a27062a,a27063a,a27067a,a27068a,a27071a,a27074a,a27075a,a27076a,a27080a,a27081a,a27084a,a27087a,a27088a,a27089a,a27093a,a27094a,a27097a,a27100a,a27101a,a27102a,a27106a,a27107a,a27110a,a27113a,a27114a,a27115a,a27119a,a27120a,a27123a,a27126a,a27127a,a27128a,a27132a,a27133a,a27136a,a27139a,a27140a,a27141a,a27145a,a27146a,a27149a,a27152a,a27153a,a27154a,a27158a,a27159a,a27162a,a27165a,a27166a,a27167a,a27171a,a27172a,a27175a,a27178a,a27179a,a27180a,a27184a,a27185a,a27188a,a27191a,a27192a,a27193a,a27197a,a27198a,a27201a,a27204a,a27205a,a27206a,a27210a,a27211a,a27214a,a27217a,a27218a,a27219a,a27223a,a27224a,a27227a,a27230a,a27231a,a27232a,a27236a,a27237a,a27240a,a27243a,a27244a,a27245a,a27249a,a27250a,a27253a,a27256a,a27257a,a27258a,a27262a,a27263a,a27266a,a27269a,a27270a,a27271a,a27275a,a27276a,a27279a,a27282a,a27283a,a27284a,a27288a,a27289a,a27292a,a27295a,a27296a,a27297a,a27301a,a27302a,a27305a,a27308a,a27309a,a27310a,a27314a,a27315a,a27318a,a27321a,a27322a,a27323a,a27327a,a27328a,a27331a,a27334a,a27335a,a27336a,a27340a,a27341a,a27344a,a27347a,a27348a,a27349a,a27353a,a27354a,a27357a,a27360a,a27361a,a27362a,a27366a,a27367a,a27370a,a27373a,a27374a,a27375a,a27379a,a27380a,a27383a,a27386a,a27387a,a27388a,a27392a,a27393a,a27396a,a27399a,a27400a,a27401a,a27405a,a27406a,a27409a,a27412a,a27413a,a27414a,a27418a,a27419a,a27422a,a27425a,a27426a,a27427a,a27431a,a27432a,a27435a,a27438a,a27439a,a27440a,a27444a,a27445a,a27448a,a27451a,a27452a,a27453a,a27457a,a27458a,a27461a,a27464a,a27465a,a27466a,a27470a,a27471a,a27474a,a27477a,a27478a,a27479a,a27483a,a27484a,a27487a,a27490a,a27491a,a27492a,a27496a,a27497a,a27500a,a27503a,a27504a,a27505a,a27509a,a27510a,a27513a,a27516a,a27517a,a27518a,a27522a,a27523a,a27526a,a27529a,a27530a,a27531a,a27535a,a27536a,a27539a,a27542a,a27543a,a27544a,a27548a,a27549a,a27552a,a27555a,a27556a,a27557a,a27561a,a27562a,a27565a,a27568a,a27569a,a27570a,a27574a,a27575a,a27578a,a27581a,a27582a,a27583a,a27587a,a27588a,a27591a,a27594a,a27595a,a27596a,a27600a,a27601a,a27604a,a27607a,a27608a,a27609a,a27613a,a27614a,a27617a,a27620a,a27621a,a27622a,a27626a,a27627a,a27630a,a27633a,a27634a,a27635a,a27639a,a27640a,a27643a,a27646a,a27647a,a27648a,a27652a,a27653a,a27656a,a27659a,a27660a,a27661a,a27665a,a27666a,a27669a,a27672a,a27673a,a27674a,a27678a,a27679a,a27682a,a27685a,a27686a,a27687a,a27691a,a27692a,a27695a,a27698a,a27699a,a27700a,a27704a,a27705a,a27708a,a27711a,a27712a,a27713a,a27717a,a27718a,a27721a,a27724a,a27725a,a27726a,a27730a,a27731a,a27734a,a27737a,a27738a,a27739a,a27743a,a27744a,a27747a,a27750a,a27751a,a27752a,a27756a,a27757a,a27760a,a27763a,a27764a,a27765a,a27769a,a27770a,a27773a,a27776a,a27777a,a27778a,a27782a,a27783a,a27786a,a27789a,a27790a,a27791a,a27795a,a27796a,a27799a,a27802a,a27803a,a27804a,a27808a,a27809a,a27812a,a27815a,a27816a,a27817a,a27821a,a27822a,a27825a,a27828a,a27829a,a27830a,a27834a,a27835a,a27838a,a27841a,a27842a,a27843a,a27847a,a27848a,a27851a,a27854a,a27855a,a27856a,a27860a,a27861a,a27864a,a27867a,a27868a,a27869a,a27873a,a27874a,a27877a,a27880a,a27881a,a27882a,a27886a,a27887a,a27890a,a27893a,a27894a,a27895a,a27899a,a27900a,a27903a,a27906a,a27907a,a27908a,a27912a,a27913a,a27916a,a27919a,a27920a,a27921a,a27925a,a27926a,a27929a,a27932a,a27933a,a27934a,a27938a,a27939a,a27942a,a27945a,a27946a,a27947a,a27951a,a27952a,a27955a,a27958a,a27959a,a27960a,a27964a,a27965a,a27968a,a27971a,a27972a,a27973a,a27977a,a27978a,a27981a,a27984a,a27985a,a27986a,a27990a,a27991a,a27994a,a27997a,a27998a,a27999a,a28003a,a28004a,a28007a,a28010a,a28011a,a28012a,a28016a,a28017a,a28020a,a28023a,a28024a,a28025a,a28029a,a28030a,a28033a,a28036a,a28037a,a28038a,a28042a,a28043a,a28046a,a28049a,a28050a,a28051a,a28055a,a28056a,a28059a,a28062a,a28063a,a28064a,a28068a,a28069a,a28072a,a28075a,a28076a,a28077a,a28081a,a28082a,a28085a,a28088a,a28089a,a28090a,a28094a,a28095a,a28098a,a28101a,a28102a,a28103a,a28107a,a28108a,a28111a,a28114a,a28115a,a28116a,a28120a,a28121a,a28124a,a28127a,a28128a,a28129a,a28133a,a28134a,a28137a,a28140a,a28141a,a28142a,a28146a,a28147a,a28150a,a28153a,a28154a,a28155a,a28159a,a28160a,a28163a,a28166a,a28167a,a28168a,a28172a,a28173a,a28176a,a28179a,a28180a,a28181a,a28185a,a28186a,a28189a,a28192a,a28193a,a28194a,a28198a,a28199a,a28202a,a28205a,a28206a,a28207a,a28211a,a28212a,a28215a,a28218a,a28219a,a28220a,a28224a,a28225a,a28228a,a28231a,a28232a,a28233a,a28237a,a28238a,a28241a,a28244a,a28245a,a28246a,a28250a,a28251a,a28254a,a28257a,a28258a,a28259a,a28263a,a28264a,a28267a,a28270a,a28271a,a28272a,a28276a,a28277a,a28280a,a28283a,a28284a,a28285a,a28289a,a28290a,a28293a,a28296a,a28297a,a28298a,a28302a,a28303a,a28306a,a28309a,a28310a,a28311a,a28315a,a28316a,a28319a,a28322a,a28323a,a28324a,a28328a,a28329a,a28332a,a28335a,a28336a,a28337a,a28341a,a28342a,a28345a,a28348a,a28349a,a28350a,a28354a,a28355a,a28358a,a28361a,a28362a,a28363a,a28367a,a28368a,a28371a,a28374a,a28375a,a28376a,a28380a,a28381a,a28384a,a28387a,a28388a,a28389a,a28393a,a28394a,a28397a,a28400a,a28401a,a28402a,a28406a,a28407a,a28410a,a28413a,a28414a,a28415a,a28419a,a28420a,a28423a,a28426a,a28427a,a28428a,a28432a,a28433a,a28436a,a28439a,a28440a,a28441a,a28445a,a28446a,a28449a,a28452a,a28453a,a28454a,a28458a,a28459a,a28462a,a28465a,a28466a,a28467a,a28471a,a28472a,a28475a,a28478a,a28479a,a28480a,a28484a,a28485a,a28488a,a28491a,a28492a,a28493a,a28497a,a28498a,a28501a,a28504a,a28505a,a28506a,a28510a,a28511a,a28514a,a28517a,a28518a,a28519a,a28523a,a28524a,a28527a,a28530a,a28531a,a28532a,a28536a,a28537a,a28540a,a28543a,a28544a,a28545a,a28549a,a28550a,a28553a,a28556a,a28557a,a28558a,a28562a,a28563a,a28566a,a28569a,a28570a,a28571a,a28575a,a28576a,a28579a,a28582a,a28583a,a28584a,a28588a,a28589a,a28592a,a28595a,a28596a,a28597a,a28601a,a28602a,a28605a,a28608a,a28609a,a28610a,a28614a,a28615a,a28618a,a28621a,a28622a,a28623a,a28627a,a28628a,a28631a,a28634a,a28635a,a28636a,a28640a,a28641a,a28644a,a28647a,a28648a,a28649a,a28653a,a28654a,a28657a,a28660a,a28661a,a28662a,a28666a,a28667a,a28670a,a28673a,a28674a,a28675a,a28679a,a28680a,a28683a,a28686a,a28687a,a28688a,a28692a,a28693a,a28696a,a28699a,a28700a,a28701a,a28705a,a28706a,a28709a,a28712a,a28713a,a28714a,a28718a,a28719a,a28722a,a28725a,a28726a,a28727a,a28731a,a28732a,a28735a,a28738a,a28739a,a28740a,a28744a,a28745a,a28748a,a28751a,a28752a,a28753a,a28757a,a28758a,a28761a,a28764a,a28765a,a28766a,a28770a,a28771a,a28774a,a28777a,a28778a,a28779a,a28783a,a28784a,a28787a,a28790a,a28791a,a28792a,a28796a,a28797a,a28800a,a28803a,a28804a,a28805a,a28809a,a28810a,a28813a,a28816a,a28817a,a28818a,a28822a,a28823a,a28826a,a28829a,a28830a,a28831a,a28835a,a28836a,a28839a,a28842a,a28843a,a28844a,a28848a,a28849a,a28852a,a28855a,a28856a,a28857a,a28861a,a28862a,a28865a,a28868a,a28869a,a28870a,a28874a,a28875a,a28878a,a28881a,a28882a,a28883a,a28887a,a28888a,a28891a,a28894a,a28895a,a28896a,a28900a,a28901a,a28904a,a28907a,a28908a,a28909a,a28913a,a28914a,a28917a,a28920a,a28921a,a28922a,a28926a,a28927a,a28930a,a28933a,a28934a,a28935a,a28939a,a28940a,a28943a,a28946a,a28947a,a28948a,a28952a,a28953a,a28956a,a28959a,a28960a,a28961a,a28965a,a28966a,a28969a,a28972a,a28973a,a28974a,a28978a,a28979a,a28982a,a28985a,a28986a,a28987a,a28991a,a28992a,a28995a,a28998a,a28999a,a29000a,a29004a,a29005a,a29008a,a29011a,a29012a,a29013a,a29017a,a29018a,a29021a,a29024a,a29025a,a29026a,a29030a,a29031a,a29034a,a29037a,a29038a,a29039a,a29043a,a29044a,a29047a,a29050a,a29051a,a29052a,a29056a,a29057a,a29060a,a29063a,a29064a,a29065a,a29069a,a29070a,a29073a,a29076a,a29077a,a29078a,a29082a,a29083a,a29086a,a29089a,a29090a,a29091a,a29095a,a29096a,a29099a,a29102a,a29103a,a29104a,a29108a,a29109a,a29112a,a29115a,a29116a,a29117a,a29121a,a29122a,a29125a,a29128a,a29129a,a29130a,a29134a,a29135a,a29138a,a29141a,a29142a,a29143a,a29147a,a29148a,a29151a,a29154a,a29155a,a29156a,a29160a,a29161a,a29164a,a29167a,a29168a,a29169a,a29173a,a29174a,a29177a,a29180a,a29181a,a29182a,a29186a,a29187a,a29190a,a29193a,a29194a,a29195a,a29199a,a29200a,a29203a,a29206a,a29207a,a29208a,a29212a,a29213a,a29216a,a29219a,a29220a,a29221a,a29225a,a29226a,a29229a,a29232a,a29233a,a29234a,a29238a,a29239a,a29242a,a29245a,a29246a,a29247a,a29251a,a29252a,a29255a,a29258a,a29259a,a29260a,a29264a,a29265a,a29268a,a29271a,a29272a,a29273a,a29277a,a29278a,a29281a,a29284a,a29285a,a29286a,a29290a,a29291a,a29294a,a29297a,a29298a,a29299a,a29303a,a29304a,a29307a,a29310a,a29311a,a29312a,a29316a,a29317a,a29320a,a29323a,a29324a,a29325a,a29329a,a29330a,a29333a,a29336a,a29337a,a29338a,a29342a,a29343a,a29346a,a29349a,a29350a,a29351a,a29355a,a29356a,a29359a,a29362a,a29363a,a29364a,a29368a,a29369a,a29372a,a29375a,a29376a,a29377a,a29381a,a29382a,a29385a,a29388a,a29389a,a29390a,a29394a,a29395a,a29398a,a29401a,a29402a,a29403a,a29407a,a29408a,a29411a,a29414a,a29415a,a29416a,a29420a,a29421a,a29424a,a29427a,a29428a,a29429a,a29433a,a29434a,a29437a,a29440a,a29441a,a29442a,a29446a,a29447a,a29450a,a29453a,a29454a,a29455a,a29459a,a29460a,a29463a,a29466a,a29467a,a29468a,a29472a,a29473a,a29476a,a29479a,a29480a,a29481a,a29485a,a29486a,a29489a,a29492a,a29493a,a29494a,a29498a,a29499a,a29502a,a29505a,a29506a,a29507a,a29511a,a29512a,a29515a,a29518a,a29519a,a29520a,a29524a,a29525a,a29528a,a29531a,a29532a,a29533a,a29537a,a29538a,a29541a,a29544a,a29545a,a29546a,a29550a,a29551a,a29554a,a29557a,a29558a,a29559a,a29563a,a29564a,a29567a,a29570a,a29571a,a29572a,a29576a,a29577a,a29580a,a29583a,a29584a,a29585a,a29589a,a29590a,a29593a,a29596a,a29597a,a29598a,a29602a,a29603a,a29606a,a29609a,a29610a,a29611a,a29615a,a29616a,a29619a,a29622a,a29623a,a29624a,a29628a,a29629a,a29632a,a29635a,a29636a,a29637a,a29641a,a29642a,a29645a,a29648a,a29649a,a29650a,a29654a,a29655a,a29658a,a29661a,a29662a,a29663a,a29667a,a29668a,a29671a,a29674a,a29675a,a29676a,a29680a,a29681a,a29684a,a29687a,a29688a,a29689a,a29693a,a29694a,a29697a,a29700a,a29701a,a29702a,a29706a,a29707a,a29710a,a29713a,a29714a,a29715a,a29719a,a29720a,a29723a,a29726a,a29727a,a29728a,a29732a,a29733a,a29736a,a29739a,a29740a,a29741a,a29745a,a29746a,a29749a,a29752a,a29753a,a29754a,a29758a,a29759a,a29762a,a29765a,a29766a,a29767a,a29771a,a29772a,a29775a,a29778a,a29779a,a29780a,a29784a,a29785a,a29788a,a29791a,a29792a,a29793a,a29797a,a29798a,a29801a,a29804a,a29805a,a29806a,a29810a,a29811a,a29814a,a29817a,a29818a,a29819a,a29823a,a29824a,a29827a,a29830a,a29831a,a29832a,a29836a,a29837a,a29840a,a29843a,a29844a,a29845a,a29849a,a29850a,a29853a,a29856a,a29857a,a29858a,a29862a,a29863a,a29866a,a29869a,a29870a,a29871a,a29875a,a29876a,a29879a,a29882a,a29883a,a29884a,a29888a,a29889a,a29892a,a29895a,a29896a,a29897a,a29901a,a29902a,a29905a,a29908a,a29909a,a29910a,a29914a,a29915a,a29918a,a29921a,a29922a,a29923a,a29927a,a29928a,a29931a,a29934a,a29935a,a29936a,a29940a,a29941a,a29944a,a29947a,a29948a,a29949a,a29953a,a29954a,a29957a,a29960a,a29961a,a29962a,a29966a,a29967a,a29970a,a29973a,a29974a,a29975a,a29979a,a29980a,a29983a,a29986a,a29987a,a29988a,a29992a,a29993a,a29996a,a29999a,a30000a,a30001a,a30005a,a30006a,a30009a,a30012a,a30013a,a30014a,a30018a,a30019a,a30022a,a30025a,a30026a,a30027a,a30031a,a30032a,a30035a,a30038a,a30039a,a30040a,a30044a,a30045a,a30048a,a30051a,a30052a,a30053a,a30057a,a30058a,a30061a,a30064a,a30065a,a30066a,a30070a,a30071a,a30074a,a30077a,a30078a,a30079a,a30083a,a30084a,a30087a,a30090a,a30091a,a30092a,a30096a,a30097a,a30100a,a30103a,a30104a,a30105a,a30109a,a30110a,a30113a,a30116a,a30117a,a30118a,a30122a,a30123a,a30126a,a30129a,a30130a,a30131a,a30135a,a30136a,a30139a,a30142a,a30143a,a30144a,a30148a,a30149a,a30152a,a30155a,a30156a,a30157a,a30161a,a30162a,a30165a,a30168a,a30169a,a30170a,a30174a,a30175a,a30178a,a30181a,a30182a,a30183a,a30187a,a30188a,a30191a,a30194a,a30195a,a30196a,a30200a,a30201a,a30204a,a30207a,a30208a,a30209a,a30213a,a30214a,a30217a,a30220a,a30221a,a30222a,a30226a,a30227a,a30230a,a30233a,a30234a,a30235a,a30239a,a30240a,a30243a,a30246a,a30247a,a30248a,a30252a,a30253a,a30256a,a30259a,a30260a,a30261a,a30265a,a30266a,a30269a,a30272a,a30273a,a30274a,a30278a,a30279a,a30282a,a30285a,a30286a,a30287a,a30291a,a30292a,a30295a,a30298a,a30299a,a30300a,a30304a,a30305a,a30308a,a30311a,a30312a,a30313a,a30317a,a30318a,a30321a,a30324a,a30325a,a30326a,a30330a,a30331a,a30334a,a30337a,a30338a,a30339a,a30343a,a30344a,a30347a,a30350a,a30351a,a30352a,a30356a,a30357a,a30360a,a30363a,a30364a,a30365a,a30369a,a30370a,a30373a,a30376a,a30377a,a30378a,a30382a,a30383a,a30386a,a30389a,a30390a,a30391a,a30395a,a30396a,a30399a,a30402a,a30403a,a30404a,a30408a,a30409a,a30412a,a30415a,a30416a,a30417a,a30421a,a30422a,a30425a,a30428a,a30429a,a30430a,a30434a,a30435a,a30438a,a30441a,a30442a,a30443a,a30447a,a30448a,a30451a,a30454a,a30455a,a30456a,a30460a,a30461a,a30464a,a30467a,a30468a,a30469a,a30473a,a30474a,a30477a,a30480a,a30481a,a30482a,a30486a,a30487a,a30490a,a30493a,a30494a,a30495a,a30499a,a30500a,a30503a,a30506a,a30507a,a30508a,a30512a,a30513a,a30516a,a30519a,a30520a,a30521a,a30525a,a30526a,a30529a,a30532a,a30533a,a30534a,a30538a,a30539a,a30542a,a30545a,a30546a,a30547a,a30551a,a30552a,a30555a,a30558a,a30559a,a30560a,a30564a,a30565a,a30568a,a30571a,a30572a,a30573a,a30577a,a30578a,a30581a,a30584a,a30585a,a30586a,a30590a,a30591a,a30594a,a30597a,a30598a,a30599a,a30603a,a30604a,a30607a,a30610a,a30611a,a30612a,a30616a,a30617a,a30620a,a30623a,a30624a,a30625a,a30629a,a30630a,a30633a,a30636a,a30637a,a30638a,a30642a,a30643a,a30646a,a30649a,a30650a,a30651a,a30655a,a30656a,a30659a,a30662a,a30663a,a30664a,a30668a,a30669a,a30672a,a30675a,a30676a,a30677a,a30681a,a30682a,a30685a,a30688a,a30689a,a30690a,a30694a,a30695a,a30698a,a30701a,a30702a,a30703a,a30707a,a30708a,a30711a,a30714a,a30715a,a30716a,a30720a,a30721a,a30724a,a30727a,a30728a,a30729a,a30733a,a30734a,a30737a,a30740a,a30741a,a30742a,a30746a,a30747a,a30750a,a30753a,a30754a,a30755a,a30759a,a30760a,a30763a,a30766a,a30767a,a30768a,a30772a,a30773a,a30776a,a30779a,a30780a,a30781a,a30785a,a30786a,a30789a,a30792a,a30793a,a30794a,a30798a,a30799a,a30802a,a30805a,a30806a,a30807a,a30811a,a30812a,a30815a,a30818a,a30819a,a30820a,a30824a,a30825a,a30828a,a30831a,a30832a,a30833a,a30837a,a30838a,a30841a,a30844a,a30845a,a30846a,a30850a,a30851a,a30854a,a30857a,a30858a,a30859a,a30863a,a30864a,a30867a,a30870a,a30871a,a30872a,a30876a,a30877a,a30880a,a30883a,a30884a,a30885a,a30889a,a30890a,a30893a,a30896a,a30897a,a30898a,a30902a,a30903a,a30906a,a30909a,a30910a,a30911a,a30915a,a30916a,a30919a,a30922a,a30923a,a30924a,a30928a,a30929a,a30932a,a30935a,a30936a,a30937a,a30941a,a30942a,a30945a,a30948a,a30949a,a30950a,a30954a,a30955a,a30958a,a30961a,a30962a,a30963a,a30967a,a30968a,a30971a,a30974a,a30975a,a30976a,a30980a,a30981a,a30984a,a30987a,a30988a,a30989a,a30993a,a30994a,a30997a,a31000a,a31001a,a31002a,a31006a,a31007a,a31010a,a31013a,a31014a,a31015a,a31019a,a31020a,a31023a,a31026a,a31027a,a31028a,a31032a,a31033a,a31036a,a31039a,a31040a,a31041a,a31045a,a31046a,a31049a,a31052a,a31053a,a31054a,a31058a,a31059a,a31062a,a31065a,a31066a,a31067a,a31071a,a31072a,a31075a,a31078a,a31079a,a31080a,a31084a,a31085a,a31088a,a31091a,a31092a,a31093a,a31097a,a31098a,a31101a,a31104a,a31105a,a31106a,a31110a,a31111a,a31114a,a31117a,a31118a,a31119a,a31123a,a31124a,a31127a,a31130a,a31131a,a31132a,a31136a,a31137a,a31140a,a31143a,a31144a,a31145a,a31149a,a31150a,a31153a,a31156a,a31157a,a31158a,a31162a,a31163a,a31166a,a31169a,a31170a,a31171a,a31175a,a31176a,a31179a,a31182a,a31183a,a31184a,a31188a,a31189a,a31192a,a31195a,a31196a,a31197a,a31201a,a31202a,a31205a,a31208a,a31209a,a31210a,a31214a,a31215a,a31218a,a31221a,a31222a,a31223a,a31227a,a31228a,a31231a,a31234a,a31235a,a31236a,a31240a,a31241a,a31244a,a31247a,a31248a,a31249a,a31253a,a31254a,a31257a,a31260a,a31261a,a31262a,a31266a,a31267a,a31270a,a31273a,a31274a,a31275a,a31279a,a31280a,a31283a,a31286a,a31287a,a31288a,a31292a,a31293a,a31296a,a31299a,a31300a,a31301a,a31305a,a31306a,a31309a,a31312a,a31313a,a31314a,a31318a,a31319a,a31322a,a31325a,a31326a,a31327a,a31331a,a31332a,a31335a,a31338a,a31339a,a31340a,a31344a,a31345a,a31348a,a31351a,a31352a,a31353a,a31357a,a31358a,a31361a,a31364a,a31365a,a31366a,a31370a,a31371a,a31374a,a31377a,a31378a,a31379a,a31383a,a31384a,a31387a,a31390a,a31391a,a31392a,a31396a,a31397a,a31400a,a31403a,a31404a,a31405a,a31409a,a31410a,a31413a,a31416a,a31417a,a31418a,a31422a,a31423a,a31426a,a31429a,a31430a,a31431a,a31435a,a31436a,a31439a,a31442a,a31443a,a31444a,a31448a,a31449a,a31452a,a31455a,a31456a,a31457a,a31461a,a31462a,a31465a,a31468a,a31469a,a31470a,a31474a,a31475a,a31478a,a31481a,a31482a,a31483a,a31487a,a31488a,a31491a,a31494a,a31495a,a31496a,a31500a,a31501a,a31504a,a31507a,a31508a,a31509a,a31513a,a31514a,a31517a,a31520a,a31521a,a31522a,a31526a,a31527a,a31530a,a31533a,a31534a,a31535a,a31539a,a31540a,a31543a,a31546a,a31547a,a31548a,a31552a,a31553a,a31556a,a31559a,a31560a,a31561a,a31565a,a31566a,a31569a,a31572a,a31573a,a31574a,a31578a,a31579a,a31582a,a31585a,a31586a,a31587a,a31591a,a31592a,a31595a,a31598a,a31599a,a31600a,a31604a,a31605a,a31608a,a31611a,a31612a,a31613a,a31617a,a31618a,a31621a,a31624a,a31625a,a31626a,a31630a,a31631a,a31634a,a31637a,a31638a,a31639a,a31643a,a31644a,a31647a,a31650a,a31651a,a31652a,a31656a,a31657a,a31660a,a31663a,a31664a,a31665a,a31669a,a31670a,a31673a,a31676a,a31677a,a31678a,a31682a,a31683a,a31686a,a31689a,a31690a,a31691a,a31695a,a31696a,a31699a,a31702a,a31703a,a31704a,a31708a,a31709a,a31712a,a31715a,a31716a,a31717a,a31721a,a31722a,a31725a,a31728a,a31729a,a31730a,a31734a,a31735a,a31738a,a31741a,a31742a,a31743a,a31747a,a31748a,a31751a,a31754a,a31755a,a31756a,a31760a,a31761a,a31764a,a31767a,a31768a,a31769a,a31773a,a31774a,a31777a,a31780a,a31781a,a31782a,a31786a,a31787a,a31790a,a31793a,a31794a,a31795a,a31799a,a31800a,a31803a,a31806a,a31807a,a31808a,a31812a,a31813a,a31816a,a31819a,a31820a,a31821a,a31825a,a31826a,a31829a,a31832a,a31833a,a31834a,a31838a,a31839a,a31842a,a31845a,a31846a,a31847a,a31851a,a31852a,a31855a,a31858a,a31859a,a31860a,a31864a,a31865a,a31868a,a31871a,a31872a,a31873a,a31877a,a31878a,a31881a,a31884a,a31885a,a31886a,a31890a,a31891a,a31894a,a31897a,a31898a,a31899a,a31903a,a31904a,a31907a,a31910a,a31911a,a31912a,a31916a,a31917a,a31920a,a31923a,a31924a,a31925a,a31929a,a31930a,a31933a,a31936a,a31937a,a31938a,a31942a,a31943a,a31946a,a31949a,a31950a,a31951a,a31955a,a31956a,a31959a,a31962a,a31963a,a31964a,a31968a,a31969a,a31972a,a31975a,a31976a,a31977a,a31981a,a31982a,a31985a,a31988a,a31989a,a31990a,a31994a,a31995a,a31998a,a32001a,a32002a,a32003a,a32007a,a32008a,a32011a,a32014a,a32015a,a32016a,a32020a,a32021a,a32024a,a32027a,a32028a,a32029a,a32033a,a32034a,a32037a,a32040a,a32041a,a32042a,a32046a,a32047a,a32050a,a32053a,a32054a,a32055a,a32059a,a32060a,a32063a,a32066a,a32067a,a32068a,a32072a,a32073a,a32076a,a32079a,a32080a,a32081a,a32085a,a32086a,a32089a,a32092a,a32093a,a32094a,a32098a,a32099a,a32102a,a32105a,a32106a,a32107a,a32111a,a32112a,a32115a,a32118a,a32119a,a32120a,a32124a,a32125a,a32128a,a32131a,a32132a,a32133a,a32137a,a32138a,a32141a,a32144a,a32145a,a32146a,a32150a,a32151a,a32154a,a32157a,a32158a,a32159a,a32163a,a32164a,a32167a,a32170a,a32171a,a32172a,a32176a,a32177a,a32180a,a32183a,a32184a,a32185a,a32189a,a32190a,a32193a,a32196a,a32197a,a32198a,a32202a,a32203a,a32206a,a32209a,a32210a,a32211a,a32215a,a32216a,a32219a,a32222a,a32223a,a32224a,a32228a,a32229a,a32232a,a32235a,a32236a,a32237a,a32241a,a32242a,a32245a,a32248a,a32249a,a32250a,a32254a,a32255a,a32258a,a32261a,a32262a,a32263a,a32267a,a32268a,a32271a,a32274a,a32275a,a32276a,a32280a,a32281a,a32284a,a32287a,a32288a,a32289a,a32293a,a32294a,a32297a,a32300a,a32301a,a32302a,a32306a,a32307a,a32310a,a32313a,a32314a,a32315a,a32319a,a32320a,a32323a,a32326a,a32327a,a32328a,a32332a,a32333a,a32336a,a32339a,a32340a,a32341a,a32345a,a32346a,a32349a,a32352a,a32353a,a32354a,a32358a,a32359a,a32362a,a32365a,a32366a,a32367a,a32371a,a32372a,a32375a,a32378a,a32379a,a32380a,a32384a,a32385a,a32388a,a32391a,a32392a,a32393a,a32397a,a32398a,a32401a,a32404a,a32405a,a32406a,a32410a,a32411a,a32414a,a32417a,a32418a,a32419a,a32423a,a32424a,a32427a,a32430a,a32431a,a32432a,a32436a,a32437a,a32440a,a32443a,a32444a,a32445a,a32449a,a32450a,a32453a,a32456a,a32457a,a32458a,a32462a,a32463a,a32466a,a32469a,a32470a,a32471a,a32475a,a32476a,a32479a,a32482a,a32483a,a32484a,a32488a,a32489a,a32492a,a32495a,a32496a,a32497a,a32501a,a32502a,a32505a,a32508a,a32509a,a32510a,a32514a,a32515a,a32518a,a32521a,a32522a,a32523a,a32527a,a32528a,a32531a,a32534a,a32535a,a32536a,a32540a,a32541a,a32544a,a32547a,a32548a,a32549a,a32553a,a32554a,a32557a,a32560a,a32561a,a32562a,a32566a,a32567a,a32570a,a32573a,a32574a,a32575a,a32579a,a32580a,a32583a,a32586a,a32587a,a32588a,a32592a,a32593a,a32596a,a32599a,a32600a,a32601a,a32605a,a32606a,a32609a,a32612a,a32613a,a32614a,a32618a,a32619a,a32622a,a32625a,a32626a,a32627a,a32631a,a32632a,a32635a,a32638a,a32639a,a32640a,a32644a,a32645a,a32648a,a32651a,a32652a,a32653a,a32657a,a32658a,a32661a,a32664a,a32665a,a32666a,a32670a,a32671a,a32674a,a32677a,a32678a,a32679a,a32683a,a32684a,a32687a,a32690a,a32691a,a32692a,a32696a,a32697a,a32700a,a32703a,a32704a,a32705a,a32709a,a32710a,a32713a,a32716a,a32717a,a32718a,a32722a,a32723a,a32726a,a32729a,a32730a,a32731a,a32735a,a32736a,a32739a,a32742a,a32743a,a32744a,a32748a,a32749a,a32752a,a32755a,a32756a,a32757a,a32761a,a32762a,a32765a,a32768a,a32769a,a32770a,a32774a,a32775a,a32778a,a32781a,a32782a,a32783a,a32787a,a32788a,a32791a,a32794a,a32795a,a32796a,a32800a,a32801a,a32804a,a32807a,a32808a,a32809a,a32813a,a32814a,a32817a,a32820a,a32821a,a32822a,a32826a,a32827a,a32830a,a32833a,a32834a,a32835a,a32839a,a32840a,a32843a,a32846a,a32847a,a32848a,a32852a,a32853a,a32856a,a32859a,a32860a,a32861a,a32865a,a32866a,a32869a,a32872a,a32873a,a32874a,a32878a,a32879a,a32882a,a32885a,a32886a,a32887a,a32891a,a32892a,a32895a,a32898a,a32899a,a32900a,a32904a,a32905a,a32908a,a32911a,a32912a,a32913a,a32917a,a32918a,a32921a,a32924a,a32925a,a32926a,a32930a,a32931a,a32934a,a32937a,a32938a,a32939a,a32943a,a32944a,a32947a,a32950a,a32951a,a32952a,a32956a,a32957a,a32960a,a32963a,a32964a,a32965a,a32969a,a32970a,a32973a,a32976a,a32977a,a32978a,a32982a,a32983a,a32986a,a32989a,a32990a,a32991a,a32995a,a32996a,a32999a,a33002a,a33003a,a33004a,a33008a,a33009a,a33012a,a33015a,a33016a,a33017a,a33021a,a33022a,a33025a,a33028a,a33029a,a33030a,a33034a,a33035a,a33038a,a33041a,a33042a,a33043a,a33047a,a33048a,a33051a,a33054a,a33055a,a33056a,a33060a,a33061a,a33064a,a33067a,a33068a,a33069a,a33073a,a33074a,a33077a,a33080a,a33081a,a33082a,a33086a,a33087a,a33090a,a33093a,a33094a,a33095a,a33099a,a33100a,a33103a,a33106a,a33107a,a33108a,a33112a,a33113a,a33116a,a33119a,a33120a,a33121a,a33125a,a33126a,a33129a,a33132a,a33133a,a33134a,a33138a,a33139a,a33142a,a33145a,a33146a,a33147a,a33151a,a33152a,a33155a,a33158a,a33159a,a33160a,a33164a,a33165a,a33168a,a33171a,a33172a,a33173a,a33177a,a33178a,a33181a,a33184a,a33185a,a33186a,a33190a,a33191a,a33194a,a33197a,a33198a,a33199a,a33203a,a33204a,a33207a,a33210a,a33211a,a33212a,a33216a,a33217a,a33220a,a33223a,a33224a,a33225a,a33229a,a33230a,a33233a,a33236a,a33237a,a33238a,a33242a,a33243a,a33246a,a33249a,a33250a,a33251a,a33255a,a33256a,a33259a,a33262a,a33263a,a33264a,a33268a,a33269a,a33272a,a33275a,a33276a,a33277a,a33281a,a33282a,a33285a,a33288a,a33289a,a33290a,a33294a,a33295a,a33298a,a33301a,a33302a,a33303a,a33307a,a33308a,a33311a,a33314a,a33315a,a33316a,a33320a,a33321a,a33324a,a33327a,a33328a,a33329a,a33333a,a33334a,a33337a,a33340a,a33341a,a33342a,a33346a,a33347a,a33350a,a33353a,a33354a,a33355a,a33359a,a33360a,a33363a,a33366a,a33367a,a33368a,a33372a,a33373a,a33376a,a33379a,a33380a,a33381a,a33385a,a33386a,a33389a,a33392a,a33393a,a33394a,a33398a,a33399a,a33402a,a33405a,a33406a,a33407a,a33411a,a33412a,a33415a,a33418a,a33419a,a33420a,a33424a,a33425a,a33428a,a33431a,a33432a,a33433a,a33437a,a33438a,a33441a,a33444a,a33445a,a33446a,a33450a,a33451a,a33454a,a33457a,a33458a,a33459a,a33463a,a33464a,a33467a,a33470a,a33471a,a33472a,a33476a,a33477a,a33480a,a33483a,a33484a,a33485a,a33489a,a33490a,a33493a,a33496a,a33497a,a33498a,a33502a,a33503a,a33506a,a33509a,a33510a,a33511a,a33515a,a33516a,a33519a,a33522a,a33523a,a33524a,a33528a,a33529a,a33532a,a33535a,a33536a,a33537a,a33541a,a33542a,a33545a,a33548a,a33549a,a33550a,a33554a,a33555a,a33558a,a33561a,a33562a,a33563a,a33567a,a33568a,a33571a,a33574a,a33575a,a33576a,a33580a,a33581a,a33584a,a33587a,a33588a,a33589a,a33593a,a33594a,a33597a,a33600a,a33601a,a33602a,a33606a,a33607a,a33610a,a33613a,a33614a,a33615a,a33619a,a33620a,a33623a,a33626a,a33627a,a33628a,a33632a,a33633a,a33636a,a33639a,a33640a,a33641a,a33645a,a33646a,a33649a,a33652a,a33653a,a33654a,a33658a,a33659a,a33662a,a33665a,a33666a,a33667a,a33671a,a33672a,a33675a,a33678a,a33679a,a33680a,a33684a,a33685a,a33688a,a33691a,a33692a,a33693a,a33697a,a33698a,a33701a,a33704a,a33705a,a33706a,a33710a,a33711a,a33714a,a33717a,a33718a,a33719a,a33723a,a33724a,a33727a,a33730a,a33731a,a33732a,a33736a,a33737a,a33740a,a33743a,a33744a,a33745a,a33749a,a33750a,a33753a,a33756a,a33757a,a33758a,a33762a,a33763a,a33766a,a33769a,a33770a,a33771a,a33775a,a33776a,a33779a,a33782a,a33783a,a33784a,a33788a,a33789a,a33792a,a33795a,a33796a,a33797a,a33801a,a33802a,a33805a,a33808a,a33809a,a33810a,a33814a,a33815a,a33818a,a33821a,a33822a,a33823a,a33827a,a33828a,a33831a,a33834a,a33835a,a33836a,a33840a,a33841a,a33844a,a33847a,a33848a,a33849a,a33853a,a33854a,a33857a,a33860a,a33861a,a33862a,a33866a,a33867a,a33870a,a33873a,a33874a,a33875a,a33879a,a33880a,a33883a,a33886a,a33887a,a33888a,a33892a,a33893a,a33896a,a33899a,a33900a,a33901a,a33905a,a33906a,a33909a,a33912a,a33913a,a33914a,a33918a,a33919a,a33922a,a33925a,a33926a,a33927a,a33931a,a33932a,a33935a,a33938a,a33939a,a33940a,a33944a,a33945a,a33948a,a33951a,a33952a,a33953a,a33957a,a33958a,a33961a,a33964a,a33965a,a33966a,a33970a,a33971a,a33974a,a33977a,a33978a,a33979a,a33983a,a33984a,a33987a,a33990a,a33991a,a33992a,a33996a,a33997a,a34000a,a34003a,a34004a,a34005a,a34009a,a34010a,a34013a,a34016a,a34017a,a34018a,a34022a,a34023a,a34026a,a34029a,a34030a,a34031a,a34035a,a34036a,a34039a,a34042a,a34043a,a34044a,a34048a,a34049a,a34052a,a34055a,a34056a,a34057a,a34061a,a34062a,a34065a,a34068a,a34069a,a34070a,a34074a,a34075a,a34078a,a34081a,a34082a,a34083a,a34087a,a34088a,a34091a,a34094a,a34095a,a34096a,a34100a,a34101a,a34104a,a34107a,a34108a,a34109a,a34113a,a34114a,a34117a,a34120a,a34121a,a34122a,a34126a,a34127a,a34130a,a34133a,a34134a,a34135a,a34139a,a34140a,a34143a,a34146a,a34147a,a34148a,a34152a,a34153a,a34156a,a34159a,a34160a,a34161a,a34165a,a34166a,a34169a,a34172a,a34173a,a34174a,a34178a,a34179a,a34182a,a34185a,a34186a,a34187a,a34191a,a34192a,a34195a,a34198a,a34199a,a34200a,a34204a,a34205a,a34208a,a34211a,a34212a,a34213a,a34217a,a34218a,a34221a,a34224a,a34225a,a34226a,a34230a,a34231a,a34234a,a34237a,a34238a,a34239a,a34243a,a34244a,a34247a,a34250a,a34251a,a34252a,a34256a,a34257a,a34260a,a34263a,a34264a,a34265a,a34269a,a34270a,a34273a,a34276a,a34277a,a34278a,a34282a,a34283a,a34286a,a34289a,a34290a,a34291a,a34295a,a34296a,a34299a,a34302a,a34303a,a34304a,a34308a,a34309a,a34312a,a34315a,a34316a,a34317a,a34321a,a34322a,a34325a,a34328a,a34329a,a34330a,a34334a,a34335a,a34338a,a34341a,a34342a,a34343a,a34347a,a34348a,a34351a,a34354a,a34355a,a34356a,a34360a,a34361a,a34364a,a34367a,a34368a,a34369a,a34373a,a34374a,a34377a,a34380a,a34381a,a34382a,a34386a,a34387a,a34390a,a34393a,a34394a,a34395a,a34399a,a34400a,a34403a,a34406a,a34407a,a34408a,a34412a,a34413a,a34416a,a34419a,a34420a,a34421a,a34425a,a34426a,a34429a,a34432a,a34433a,a34434a,a34438a,a34439a,a34442a,a34445a,a34446a,a34447a,a34450a,a34453a,a34454a,a34457a,a34460a,a34461a,a34462a,a34466a,a34467a,a34470a,a34473a,a34474a,a34475a,a34478a,a34481a,a34482a,a34485a,a34488a,a34489a,a34490a,a34494a,a34495a,a34498a,a34501a,a34502a,a34503a,a34506a,a34509a,a34510a,a34513a,a34516a,a34517a,a34518a,a34522a,a34523a,a34526a,a34529a,a34530a,a34531a,a34534a,a34537a,a34538a,a34541a,a34544a,a34545a,a34546a,a34550a,a34551a,a34554a,a34557a,a34558a,a34559a,a34562a,a34565a,a34566a,a34569a,a34572a,a34573a,a34574a,a34578a,a34579a,a34582a,a34585a,a34586a,a34587a,a34590a,a34593a,a34594a,a34597a,a34600a,a34601a,a34602a,a34606a,a34607a,a34610a,a34613a,a34614a,a34615a,a34618a,a34621a,a34622a,a34625a,a34628a,a34629a,a34630a,a34634a,a34635a,a34638a,a34641a,a34642a,a34643a,a34646a,a34649a,a34650a,a34653a,a34656a,a34657a,a34658a,a34662a,a34663a,a34666a,a34669a,a34670a,a34671a,a34674a,a34677a,a34678a,a34681a,a34684a,a34685a,a34686a,a34690a,a34691a,a34694a,a34697a,a34698a,a34699a,a34702a,a34705a,a34706a,a34709a,a34712a,a34713a,a34714a,a34718a,a34719a,a34722a,a34725a,a34726a,a34727a,a34730a,a34733a,a34734a,a34737a,a34740a,a34741a,a34742a,a34746a,a34747a,a34750a,a34753a,a34754a,a34755a,a34758a,a34761a,a34762a,a34765a,a34768a,a34769a,a34770a,a34774a,a34775a,a34778a,a34781a,a34782a,a34783a,a34786a,a34789a,a34790a,a34793a,a34796a,a34797a,a34798a,a34802a,a34803a,a34806a,a34809a,a34810a,a34811a,a34814a,a34817a,a34818a,a34821a,a34824a,a34825a,a34826a,a34830a,a34831a,a34834a,a34837a,a34838a,a34839a,a34842a,a34845a,a34846a,a34849a,a34852a,a34853a,a34854a,a34858a,a34859a,a34862a,a34865a,a34866a,a34867a,a34870a,a34873a,a34874a,a34877a,a34880a,a34881a,a34882a,a34886a,a34887a,a34890a,a34893a,a34894a,a34895a,a34898a,a34901a,a34902a,a34905a,a34908a,a34909a,a34910a,a34914a,a34915a,a34918a,a34921a,a34922a,a34923a,a34926a,a34929a,a34930a,a34933a,a34936a,a34937a,a34938a,a34942a,a34943a,a34946a,a34949a,a34950a,a34951a,a34954a,a34957a,a34958a,a34961a,a34964a,a34965a,a34966a,a34970a,a34971a,a34974a,a34977a,a34978a,a34979a,a34982a,a34985a,a34986a,a34989a,a34992a,a34993a,a34994a,a34998a,a34999a,a35002a,a35005a,a35006a,a35007a,a35010a,a35013a,a35014a,a35017a,a35020a,a35021a,a35022a,a35026a,a35027a,a35030a,a35033a,a35034a,a35035a,a35038a,a35041a,a35042a,a35045a,a35048a,a35049a,a35050a,a35054a,a35055a,a35058a,a35061a,a35062a,a35063a,a35066a,a35069a,a35070a,a35073a,a35076a,a35077a,a35078a,a35082a,a35083a,a35086a,a35089a,a35090a,a35091a,a35094a,a35097a,a35098a,a35101a,a35104a,a35105a,a35106a,a35110a,a35111a,a35114a,a35117a,a35118a,a35119a,a35122a,a35125a,a35126a,a35129a,a35132a,a35133a,a35134a,a35138a,a35139a,a35142a,a35145a,a35146a,a35147a,a35150a,a35153a,a35154a,a35157a,a35160a,a35161a,a35162a,a35166a,a35167a,a35170a,a35173a,a35174a,a35175a,a35178a,a35181a,a35182a,a35185a,a35188a,a35189a,a35190a,a35194a,a35195a,a35198a,a35201a,a35202a,a35203a,a35206a,a35209a,a35210a,a35213a,a35216a,a35217a,a35218a,a35222a,a35223a,a35226a,a35229a,a35230a,a35231a,a35234a,a35237a,a35238a,a35241a,a35244a,a35245a,a35246a,a35250a,a35251a,a35254a,a35257a,a35258a,a35259a,a35262a,a35265a,a35266a,a35269a,a35272a,a35273a,a35274a,a35278a,a35279a,a35282a,a35285a,a35286a,a35287a,a35290a,a35293a,a35294a,a35297a,a35300a,a35301a,a35302a,a35306a,a35307a,a35310a,a35313a,a35314a,a35315a,a35318a,a35321a,a35322a,a35325a,a35328a,a35329a,a35330a,a35334a,a35335a,a35338a,a35341a,a35342a,a35343a,a35346a,a35349a,a35350a,a35353a,a35356a,a35357a,a35358a,a35362a,a35363a,a35366a,a35369a,a35370a,a35371a,a35374a,a35377a,a35378a,a35381a,a35384a,a35385a,a35386a,a35390a,a35391a,a35394a,a35397a,a35398a,a35399a,a35402a,a35405a,a35406a,a35409a,a35412a,a35413a,a35414a,a35418a,a35419a,a35422a,a35425a,a35426a,a35427a,a35430a,a35433a,a35434a,a35437a,a35440a,a35441a,a35442a,a35446a,a35447a,a35450a,a35453a,a35454a,a35455a,a35458a,a35461a,a35462a,a35465a,a35468a,a35469a,a35470a,a35474a,a35475a,a35478a,a35481a,a35482a,a35483a,a35486a,a35489a,a35490a,a35493a,a35496a,a35497a,a35498a,a35502a,a35503a,a35506a,a35509a,a35510a,a35511a,a35514a,a35517a,a35518a,a35521a,a35524a,a35525a,a35526a,a35530a,a35531a,a35534a,a35537a,a35538a,a35539a,a35542a,a35545a,a35546a,a35549a,a35552a,a35553a,a35554a,a35558a,a35559a,a35562a,a35565a,a35566a,a35567a,a35570a,a35573a,a35574a,a35577a,a35580a,a35581a,a35582a,a35586a,a35587a,a35590a,a35593a,a35594a,a35595a,a35598a,a35601a,a35602a,a35605a,a35608a,a35609a,a35610a,a35614a,a35615a,a35618a,a35621a,a35622a,a35623a,a35626a,a35629a,a35630a,a35633a,a35636a,a35637a,a35638a,a35642a,a35643a,a35646a,a35649a,a35650a,a35651a,a35654a,a35657a,a35658a,a35661a,a35664a,a35665a,a35666a,a35670a,a35671a,a35674a,a35677a,a35678a,a35679a,a35682a,a35685a,a35686a,a35689a,a35692a,a35693a,a35694a,a35698a,a35699a,a35702a,a35705a,a35706a,a35707a,a35710a,a35713a,a35714a,a35717a,a35720a,a35721a,a35722a,a35726a,a35727a,a35730a,a35733a,a35734a,a35735a,a35738a,a35741a,a35742a,a35745a,a35748a,a35749a,a35750a,a35754a,a35755a,a35758a,a35761a,a35762a,a35763a,a35766a,a35769a,a35770a,a35773a,a35776a,a35777a,a35778a,a35782a,a35783a,a35786a,a35789a,a35790a,a35791a,a35794a,a35797a,a35798a,a35801a,a35804a,a35805a,a35806a,a35810a,a35811a,a35814a,a35817a,a35818a,a35819a,a35822a,a35825a,a35826a,a35829a,a35832a,a35833a,a35834a,a35838a,a35839a,a35842a,a35845a,a35846a,a35847a,a35850a,a35853a,a35854a,a35857a,a35860a,a35861a,a35862a,a35866a,a35867a,a35870a,a35873a,a35874a,a35875a,a35878a,a35881a,a35882a,a35885a,a35888a,a35889a,a35890a,a35894a,a35895a,a35898a,a35901a,a35902a,a35903a,a35906a,a35909a,a35910a,a35913a,a35916a,a35917a,a35918a,a35922a,a35923a,a35926a,a35929a,a35930a,a35931a,a35934a,a35937a,a35938a,a35941a,a35944a,a35945a,a35946a,a35950a,a35951a,a35954a,a35957a,a35958a,a35959a,a35962a,a35965a,a35966a,a35969a,a35972a,a35973a,a35974a,a35978a,a35979a,a35982a,a35985a,a35986a,a35987a,a35990a,a35993a,a35994a,a35997a,a36000a,a36001a,a36002a,a36006a,a36007a,a36010a,a36013a,a36014a,a36015a,a36018a,a36021a,a36022a,a36025a,a36028a,a36029a,a36030a,a36034a,a36035a,a36038a,a36041a,a36042a,a36043a,a36046a,a36049a,a36050a,a36053a,a36056a,a36057a,a36058a,a36062a,a36063a,a36066a,a36069a,a36070a,a36071a,a36074a,a36077a,a36078a,a36081a,a36084a,a36085a,a36086a,a36090a,a36091a,a36094a,a36097a,a36098a,a36099a,a36102a,a36105a,a36106a,a36109a,a36112a,a36113a,a36114a,a36118a,a36119a,a36122a,a36125a,a36126a,a36127a,a36130a,a36133a,a36134a,a36137a,a36140a,a36141a,a36142a,a36146a,a36147a,a36150a,a36153a,a36154a,a36155a,a36158a,a36161a,a36162a,a36165a,a36168a,a36169a,a36170a,a36174a,a36175a,a36178a,a36181a,a36182a,a36183a,a36186a,a36189a,a36190a,a36193a,a36196a,a36197a,a36198a,a36202a,a36203a,a36206a,a36209a,a36210a,a36211a,a36214a,a36217a,a36218a,a36221a,a36224a,a36225a,a36226a,a36230a,a36231a,a36234a,a36237a,a36238a,a36239a,a36242a,a36245a,a36246a,a36249a,a36252a,a36253a,a36254a,a36258a,a36259a,a36262a,a36265a,a36266a,a36267a,a36270a,a36273a,a36274a,a36277a,a36280a,a36281a,a36282a,a36286a,a36287a,a36290a,a36293a,a36294a,a36295a,a36298a,a36301a,a36302a,a36305a,a36308a,a36309a,a36310a,a36314a,a36315a,a36318a,a36321a,a36322a,a36323a,a36326a,a36329a,a36330a,a36333a,a36336a,a36337a,a36338a,a36342a,a36343a,a36346a,a36349a,a36350a,a36351a,a36354a,a36357a,a36358a,a36361a,a36364a,a36365a,a36366a,a36370a,a36371a,a36374a,a36377a,a36378a,a36379a,a36382a,a36385a,a36386a,a36389a,a36392a,a36393a,a36394a,a36398a,a36399a,a36402a,a36405a,a36406a,a36407a,a36410a,a36413a,a36414a,a36417a,a36420a,a36421a,a36422a,a36426a,a36427a,a36430a,a36433a,a36434a,a36435a,a36438a,a36441a,a36442a,a36445a,a36448a,a36449a,a36450a,a36454a,a36455a,a36458a,a36461a,a36462a,a36463a,a36466a,a36469a,a36470a,a36473a,a36476a,a36477a,a36478a,a36482a,a36483a,a36486a,a36489a,a36490a,a36491a,a36494a,a36497a,a36498a,a36501a,a36504a,a36505a,a36506a,a36510a,a36511a,a36514a,a36517a,a36518a,a36519a,a36522a,a36525a,a36526a,a36529a,a36532a,a36533a,a36534a,a36538a,a36539a,a36542a,a36545a,a36546a,a36547a,a36550a,a36553a,a36554a,a36557a,a36560a,a36561a,a36562a,a36566a,a36567a,a36570a,a36573a,a36574a,a36575a,a36578a,a36581a,a36582a,a36585a,a36588a,a36589a,a36590a,a36594a,a36595a,a36598a,a36601a,a36602a,a36603a,a36606a,a36609a,a36610a,a36613a,a36616a,a36617a,a36618a,a36622a,a36623a,a36626a,a36629a,a36630a,a36631a,a36634a,a36637a,a36638a,a36641a,a36644a,a36645a,a36646a,a36650a,a36651a,a36654a,a36657a,a36658a,a36659a,a36662a,a36665a,a36666a,a36669a,a36672a,a36673a,a36674a,a36678a,a36679a,a36682a,a36685a,a36686a,a36687a,a36690a,a36693a,a36694a,a36697a,a36700a,a36701a,a36702a,a36706a,a36707a,a36710a,a36713a,a36714a,a36715a,a36718a,a36721a,a36722a,a36725a,a36728a,a36729a,a36730a,a36734a,a36735a,a36738a,a36741a,a36742a,a36743a,a36746a,a36749a,a36750a,a36753a,a36756a,a36757a,a36758a,a36762a,a36763a,a36766a,a36769a,a36770a,a36771a,a36774a,a36777a,a36778a,a36781a,a36784a,a36785a,a36786a,a36790a,a36791a,a36794a,a36797a,a36798a,a36799a,a36802a,a36805a,a36806a,a36809a,a36812a,a36813a,a36814a,a36818a,a36819a,a36822a,a36825a,a36826a,a36827a,a36830a,a36833a,a36834a,a36837a,a36840a,a36841a,a36842a,a36846a,a36847a,a36850a,a36853a,a36854a,a36855a,a36858a,a36861a,a36862a,a36865a,a36868a,a36869a,a36870a,a36874a,a36875a,a36878a,a36881a,a36882a,a36883a,a36886a,a36889a,a36890a,a36893a,a36896a,a36897a,a36898a,a36902a,a36903a,a36906a,a36909a,a36910a,a36911a,a36914a,a36917a,a36918a,a36921a,a36924a,a36925a,a36926a,a36930a,a36931a,a36934a,a36937a,a36938a,a36939a,a36942a,a36945a,a36946a,a36949a,a36952a,a36953a,a36954a,a36958a,a36959a,a36962a,a36965a,a36966a,a36967a,a36970a,a36973a,a36974a,a36977a,a36980a,a36981a,a36982a,a36986a,a36987a,a36990a,a36993a,a36994a,a36995a,a36998a,a37001a,a37002a,a37005a,a37008a,a37009a,a37010a,a37014a,a37015a,a37018a,a37021a,a37022a,a37023a,a37026a,a37029a,a37030a,a37033a,a37036a,a37037a,a37038a,a37042a,a37043a,a37046a,a37049a,a37050a,a37051a,a37054a,a37057a,a37058a,a37061a,a37064a,a37065a,a37066a,a37070a,a37071a,a37074a,a37077a,a37078a,a37079a,a37082a,a37085a,a37086a,a37089a,a37092a,a37093a,a37094a,a37098a,a37099a,a37102a,a37105a,a37106a,a37107a,a37110a,a37113a,a37114a,a37117a,a37120a,a37121a,a37122a,a37126a,a37127a,a37130a,a37133a,a37134a,a37135a,a37138a,a37141a,a37142a,a37145a,a37148a,a37149a,a37150a,a37154a,a37155a,a37158a,a37161a,a37162a,a37163a,a37166a,a37169a,a37170a,a37173a,a37176a,a37177a,a37178a,a37182a,a37183a,a37186a,a37189a,a37190a,a37191a,a37194a,a37197a,a37198a,a37201a,a37204a,a37205a,a37206a,a37210a,a37211a,a37214a,a37217a,a37218a,a37219a,a37222a,a37225a,a37226a,a37229a,a37232a,a37233a,a37234a,a37238a,a37239a,a37242a,a37245a,a37246a,a37247a,a37250a,a37253a,a37254a,a37257a,a37260a,a37261a,a37262a,a37266a,a37267a,a37270a,a37273a,a37274a,a37275a,a37278a,a37281a,a37282a,a37285a,a37288a,a37289a,a37290a,a37294a,a37295a,a37298a,a37301a,a37302a,a37303a,a37306a,a37309a,a37310a,a37313a,a37316a,a37317a,a37318a,a37322a,a37323a,a37326a,a37329a,a37330a,a37331a,a37334a,a37337a,a37338a,a37341a,a37344a,a37345a,a37346a,a37350a,a37351a,a37354a,a37357a,a37358a,a37359a,a37362a,a37365a,a37366a,a37369a,a37372a,a37373a,a37374a,a37378a,a37379a,a37382a,a37385a,a37386a,a37387a,a37390a,a37393a,a37394a,a37397a,a37400a,a37401a,a37402a,a37406a,a37407a,a37410a,a37413a,a37414a,a37415a,a37418a,a37421a,a37422a,a37425a,a37428a,a37429a,a37430a,a37434a,a37435a,a37438a,a37441a,a37442a,a37443a,a37446a,a37449a,a37450a,a37453a,a37456a,a37457a,a37458a,a37462a,a37463a,a37466a,a37469a,a37470a,a37471a,a37474a,a37477a,a37478a,a37481a,a37484a,a37485a,a37486a,a37490a,a37491a,a37494a,a37497a,a37498a,a37499a,a37502a,a37505a,a37506a,a37509a,a37512a,a37513a,a37514a,a37518a,a37519a,a37522a,a37525a,a37526a,a37527a,a37530a,a37533a,a37534a,a37537a,a37540a,a37541a,a37542a,a37546a,a37547a,a37550a,a37553a,a37554a,a37555a,a37558a,a37561a,a37562a,a37565a,a37568a,a37569a,a37570a,a37574a,a37575a,a37578a,a37581a,a37582a,a37583a,a37586a,a37589a,a37590a,a37593a,a37596a,a37597a,a37598a,a37602a,a37603a,a37606a,a37609a,a37610a,a37611a,a37614a,a37617a,a37618a,a37621a,a37624a,a37625a,a37626a,a37630a,a37631a,a37634a,a37637a,a37638a,a37639a,a37642a,a37645a,a37646a,a37649a,a37652a,a37653a,a37654a,a37658a,a37659a,a37662a,a37665a,a37666a,a37667a,a37670a,a37673a,a37674a,a37677a,a37680a,a37681a,a37682a,a37686a,a37687a,a37690a,a37693a,a37694a,a37695a,a37698a,a37701a,a37702a,a37705a,a37708a,a37709a,a37710a,a37714a,a37715a,a37718a,a37721a,a37722a,a37723a,a37726a,a37729a,a37730a,a37733a,a37736a,a37737a,a37738a,a37742a,a37743a,a37746a,a37749a,a37750a,a37751a,a37754a,a37757a,a37758a,a37761a,a37764a,a37765a,a37766a,a37770a,a37771a,a37774a,a37777a,a37778a,a37779a,a37782a,a37785a,a37786a,a37789a,a37792a,a37793a,a37794a,a37798a,a37799a,a37802a,a37805a,a37806a,a37807a,a37810a,a37813a,a37814a,a37817a,a37820a,a37821a,a37822a,a37826a,a37827a,a37830a,a37833a,a37834a,a37835a,a37838a,a37841a,a37842a,a37845a,a37848a,a37849a,a37850a,a37854a,a37855a,a37858a,a37861a,a37862a,a37863a,a37866a,a37869a,a37870a,a37873a,a37876a,a37877a,a37878a,a37882a,a37883a,a37886a,a37889a,a37890a,a37891a,a37894a,a37897a,a37898a,a37901a,a37904a,a37905a,a37906a,a37910a,a37911a,a37914a,a37917a,a37918a,a37919a,a37922a,a37925a,a37926a,a37929a,a37932a,a37933a,a37934a,a37938a,a37939a,a37942a,a37945a,a37946a,a37947a,a37950a,a37953a,a37954a,a37957a,a37960a,a37961a,a37962a,a37966a,a37967a,a37970a,a37973a,a37974a,a37975a,a37978a,a37981a,a37982a,a37985a,a37988a,a37989a,a37990a,a37994a,a37995a,a37998a,a38001a,a38002a,a38003a,a38006a,a38009a,a38010a,a38013a,a38016a,a38017a,a38018a,a38021a,a38024a,a38025a,a38028a,a38031a,a38032a,a38033a,a38036a,a38039a,a38040a,a38043a,a38046a,a38047a,a38048a,a38051a,a38054a,a38055a,a38058a,a38061a,a38062a,a38063a,a38066a,a38069a,a38070a,a38073a,a38076a,a38077a,a38078a,a38081a,a38084a,a38085a,a38088a,a38091a,a38092a,a38093a,a38096a,a38099a,a38100a,a38103a,a38106a,a38107a,a38108a,a38111a,a38114a,a38115a,a38118a,a38121a,a38122a,a38123a,a38126a,a38129a,a38130a,a38133a,a38136a,a38137a,a38138a,a38141a,a38144a,a38145a,a38148a,a38151a,a38152a,a38153a,a38156a,a38159a,a38160a,a38163a,a38166a,a38167a,a38168a,a38171a,a38174a,a38175a,a38178a,a38181a,a38182a,a38183a,a38186a,a38189a,a38190a,a38193a,a38196a,a38197a,a38198a,a38201a,a38204a,a38205a,a38208a,a38211a,a38212a,a38213a,a38216a,a38219a,a38220a,a38223a,a38226a,a38227a,a38228a,a38231a,a38234a,a38235a,a38238a,a38241a,a38242a,a38243a,a38246a,a38249a,a38250a,a38253a,a38256a,a38257a,a38258a,a38261a,a38264a,a38265a,a38268a,a38271a,a38272a,a38273a,a38276a,a38279a,a38280a,a38283a,a38286a,a38287a,a38288a,a38291a,a38294a,a38295a,a38298a,a38301a,a38302a,a38303a,a38306a,a38309a,a38310a,a38313a,a38316a,a38317a,a38318a,a38321a,a38324a,a38325a,a38328a,a38331a,a38332a,a38333a,a38336a,a38339a,a38340a,a38343a,a38346a,a38347a,a38348a,a38351a,a38354a,a38355a,a38358a,a38361a,a38362a,a38363a,a38366a,a38369a,a38370a,a38373a,a38376a,a38377a,a38378a,a38381a,a38384a,a38385a,a38388a,a38391a,a38392a,a38393a,a38396a,a38399a,a38400a,a38403a,a38406a,a38407a,a38408a,a38411a,a38414a,a38415a,a38418a,a38421a,a38422a,a38423a,a38426a,a38429a,a38430a,a38433a,a38436a,a38437a,a38438a,a38441a,a38444a,a38445a,a38448a,a38451a,a38452a,a38453a,a38456a,a38459a,a38460a,a38463a,a38466a,a38467a,a38468a,a38471a,a38474a,a38475a,a38478a,a38481a,a38482a,a38483a,a38486a,a38489a,a38490a,a38493a,a38496a,a38497a,a38498a,a38501a,a38504a,a38505a,a38508a,a38511a,a38512a,a38513a,a38516a,a38519a,a38520a,a38523a,a38526a,a38527a,a38528a,a38531a,a38534a,a38535a,a38538a,a38541a,a38542a,a38543a,a38546a,a38549a,a38550a,a38553a,a38556a,a38557a,a38558a,a38561a,a38564a,a38565a,a38568a,a38571a,a38572a,a38573a,a38576a,a38579a,a38580a,a38583a,a38586a,a38587a,a38588a,a38591a,a38594a,a38595a,a38598a,a38601a,a38602a,a38603a,a38606a,a38609a,a38610a,a38613a,a38616a,a38617a,a38618a,a38621a,a38624a,a38625a,a38628a,a38631a,a38632a,a38633a,a38636a,a38639a,a38640a,a38643a,a38646a,a38647a,a38648a,a38651a,a38654a,a38655a,a38658a,a38661a,a38662a,a38663a,a38666a,a38669a,a38670a,a38673a,a38676a,a38677a,a38678a,a38681a,a38684a,a38685a,a38688a,a38691a,a38692a,a38693a,a38696a,a38699a,a38700a,a38703a,a38706a,a38707a,a38708a,a38711a,a38714a,a38715a,a38718a,a38721a,a38722a,a38723a,a38726a,a38729a,a38730a,a38733a,a38736a,a38737a,a38738a,a38741a,a38744a,a38745a,a38748a,a38751a,a38752a,a38753a,a38756a,a38759a,a38760a,a38763a,a38766a,a38767a,a38768a,a38771a,a38774a,a38775a,a38778a,a38781a,a38782a,a38783a,a38786a,a38789a,a38790a,a38793a,a38796a,a38797a,a38798a,a38801a,a38804a,a38805a,a38808a,a38811a,a38812a,a38813a,a38816a,a38819a,a38820a,a38823a,a38826a,a38827a,a38828a,a38831a,a38834a,a38835a,a38838a,a38841a,a38842a,a38843a,a38846a,a38849a,a38850a,a38853a,a38856a,a38857a,a38858a,a38861a,a38864a,a38865a,a38868a,a38871a,a38872a,a38873a,a38876a,a38879a,a38880a,a38883a,a38886a,a38887a,a38888a,a38891a,a38894a,a38895a,a38898a,a38901a,a38902a,a38903a,a38906a,a38909a,a38910a,a38913a,a38916a,a38917a,a38918a,a38921a,a38924a,a38925a,a38928a,a38931a,a38932a,a38933a,a38936a,a38939a,a38940a,a38943a,a38946a,a38947a,a38948a,a38951a,a38954a,a38955a,a38958a,a38961a,a38962a,a38963a,a38966a,a38969a,a38970a,a38973a,a38976a,a38977a,a38978a,a38981a,a38984a,a38985a,a38988a,a38991a,a38992a,a38993a,a38996a,a38999a,a39000a,a39003a,a39006a,a39007a,a39008a,a39011a,a39014a,a39015a,a39018a,a39021a,a39022a,a39023a,a39026a,a39029a,a39030a,a39033a,a39036a,a39037a,a39038a,a39041a,a39044a,a39045a,a39048a,a39051a,a39052a,a39053a,a39056a,a39059a,a39060a,a39063a,a39066a,a39067a,a39068a,a39071a,a39074a,a39075a,a39078a,a39081a,a39082a,a39083a,a39086a,a39089a,a39090a,a39093a,a39096a,a39097a,a39098a,a39101a,a39104a,a39105a,a39108a,a39111a,a39112a,a39113a,a39116a,a39119a,a39120a,a39123a,a39126a,a39127a,a39128a,a39131a,a39134a,a39135a,a39138a,a39141a,a39142a,a39143a,a39146a,a39149a,a39150a,a39153a,a39156a,a39157a,a39158a,a39161a,a39164a,a39165a,a39168a,a39171a,a39172a,a39173a,a39176a,a39179a,a39180a,a39183a,a39186a,a39187a,a39188a,a39191a,a39194a,a39195a,a39198a,a39201a,a39202a,a39203a,a39206a,a39209a,a39210a,a39213a,a39216a,a39217a,a39218a,a39221a,a39224a,a39225a,a39228a,a39231a,a39232a,a39233a,a39236a,a39239a,a39240a,a39243a,a39246a,a39247a,a39248a,a39251a,a39254a,a39255a,a39258a,a39261a,a39262a,a39263a,a39266a,a39269a,a39270a,a39273a,a39276a,a39277a,a39278a,a39281a,a39284a,a39285a,a39288a,a39291a,a39292a,a39293a,a39296a,a39299a,a39300a,a39303a,a39306a,a39307a,a39308a,a39311a,a39314a,a39315a,a39318a,a39321a,a39322a,a39323a,a39326a,a39329a,a39330a,a39333a,a39336a,a39337a,a39338a,a39341a,a39344a,a39345a,a39348a,a39351a,a39352a,a39353a,a39356a,a39359a,a39360a,a39363a,a39366a,a39367a,a39368a,a39371a,a39374a,a39375a,a39378a,a39381a,a39382a,a39383a,a39386a,a39389a,a39390a,a39393a,a39396a,a39397a,a39398a,a39401a,a39404a,a39405a,a39408a,a39411a,a39412a,a39413a,a39416a,a39419a,a39420a,a39423a,a39426a,a39427a,a39428a,a39431a,a39434a,a39435a,a39438a,a39441a,a39442a,a39443a,a39446a,a39449a,a39450a,a39453a,a39456a,a39457a,a39458a,a39461a,a39464a,a39465a,a39468a,a39471a,a39472a,a39473a,a39476a,a39479a,a39480a,a39483a,a39486a,a39487a,a39488a,a39491a,a39494a,a39495a,a39498a,a39501a,a39502a,a39503a,a39506a,a39509a,a39510a,a39513a,a39516a,a39517a,a39518a,a39521a,a39524a,a39525a,a39528a,a39531a,a39532a,a39533a,a39536a,a39539a,a39540a,a39543a,a39546a,a39547a,a39548a,a39551a,a39554a,a39555a,a39558a,a39561a,a39562a,a39563a,a39566a,a39569a,a39570a,a39573a,a39576a,a39577a,a39578a,a39581a,a39584a,a39585a,a39588a,a39591a,a39592a,a39593a,a39596a,a39599a,a39600a,a39603a,a39606a,a39607a,a39608a,a39611a,a39614a,a39615a,a39618a,a39621a,a39622a,a39623a,a39626a,a39629a,a39630a,a39633a,a39636a,a39637a,a39638a,a39641a,a39644a,a39645a,a39648a,a39651a,a39652a,a39653a,a39656a,a39659a,a39660a,a39663a,a39666a,a39667a,a39668a,a39671a,a39674a,a39675a,a39678a,a39681a,a39682a,a39683a,a39686a,a39689a,a39690a,a39693a,a39696a,a39697a,a39698a,a39701a,a39704a,a39705a,a39708a,a39711a,a39712a,a39713a,a39716a,a39719a,a39720a,a39723a,a39726a,a39727a,a39728a,a39731a,a39734a,a39735a,a39738a,a39741a,a39742a,a39743a,a39746a,a39749a,a39750a,a39753a,a39756a,a39757a,a39758a,a39761a,a39764a,a39765a,a39768a,a39771a,a39772a,a39773a,a39776a,a39779a,a39780a,a39783a,a39786a,a39787a,a39788a,a39791a,a39794a,a39795a,a39798a,a39801a,a39802a,a39803a,a39806a,a39809a,a39810a,a39813a,a39816a,a39817a,a39818a,a39821a,a39824a,a39825a,a39828a,a39831a,a39832a,a39833a,a39836a,a39839a,a39840a,a39843a,a39846a,a39847a,a39848a,a39851a,a39854a,a39855a,a39858a,a39861a,a39862a,a39863a,a39866a,a39869a,a39870a,a39873a,a39876a,a39877a,a39878a,a39881a,a39884a,a39885a,a39888a,a39891a,a39892a,a39893a,a39896a,a39899a,a39900a,a39903a,a39906a,a39907a,a39908a,a39911a,a39914a,a39915a,a39918a,a39921a,a39922a,a39923a,a39926a,a39929a,a39930a,a39933a,a39936a,a39937a,a39938a,a39941a,a39944a,a39945a,a39948a,a39951a,a39952a,a39953a,a39956a,a39959a,a39960a,a39963a,a39966a,a39967a,a39968a,a39971a,a39974a,a39975a,a39978a,a39981a,a39982a,a39983a,a39986a,a39989a,a39990a,a39993a,a39996a,a39997a,a39998a,a40001a,a40004a,a40005a,a40008a,a40011a,a40012a,a40013a,a40016a,a40019a,a40020a,a40023a,a40026a,a40027a,a40028a,a40031a,a40034a,a40035a,a40038a,a40041a,a40042a,a40043a,a40046a,a40049a,a40050a,a40053a,a40056a,a40057a,a40058a,a40061a,a40064a,a40065a,a40068a,a40071a,a40072a,a40073a,a40076a,a40079a,a40080a,a40083a,a40086a,a40087a,a40088a,a40091a,a40094a,a40095a,a40098a,a40101a,a40102a,a40103a,a40106a,a40109a,a40110a,a40113a,a40116a,a40117a,a40118a,a40121a,a40124a,a40125a,a40128a,a40131a,a40132a,a40133a,a40136a,a40139a,a40140a,a40143a,a40146a,a40147a,a40148a,a40151a,a40154a,a40155a,a40158a,a40161a,a40162a,a40163a,a40166a,a40169a,a40170a,a40173a,a40176a,a40177a,a40178a,a40181a,a40184a,a40185a,a40188a,a40191a,a40192a,a40193a,a40196a,a40199a,a40200a,a40203a,a40206a,a40207a,a40208a,a40211a,a40214a,a40215a,a40218a,a40221a,a40222a,a40223a,a40226a,a40229a,a40230a,a40233a,a40236a,a40237a,a40238a,a40241a,a40244a,a40245a,a40248a,a40251a,a40252a,a40253a,a40256a,a40259a,a40260a,a40263a,a40266a,a40267a,a40268a,a40271a,a40274a,a40275a,a40278a,a40281a,a40282a,a40283a,a40286a,a40289a,a40290a,a40293a,a40296a,a40297a,a40298a,a40301a,a40304a,a40305a,a40308a,a40311a,a40312a,a40313a,a40316a,a40319a,a40320a,a40323a,a40326a,a40327a,a40328a,a40331a,a40334a,a40335a,a40338a,a40341a,a40342a,a40343a,a40346a,a40349a,a40350a,a40353a,a40356a,a40357a,a40358a,a40361a,a40364a,a40365a,a40368a,a40371a,a40372a,a40373a,a40376a,a40379a,a40380a,a40383a,a40386a,a40387a,a40388a,a40391a,a40394a,a40395a,a40398a,a40401a,a40402a,a40403a,a40406a,a40409a,a40410a,a40413a,a40416a,a40417a,a40418a,a40421a,a40424a,a40425a,a40428a,a40431a,a40432a,a40433a,a40436a,a40439a,a40440a,a40443a,a40446a,a40447a,a40448a,a40451a,a40454a,a40455a,a40458a,a40461a,a40462a,a40463a,a40466a,a40469a,a40470a,a40473a,a40476a,a40477a,a40478a,a40481a,a40484a,a40485a,a40488a,a40491a,a40492a,a40493a,a40496a,a40499a,a40500a,a40503a,a40506a,a40507a,a40508a,a40511a,a40514a,a40515a,a40518a,a40521a,a40522a,a40523a,a40526a,a40529a,a40530a,a40533a,a40536a,a40537a,a40538a,a40541a,a40544a,a40545a,a40548a,a40551a,a40552a,a40553a,a40556a,a40559a,a40560a,a40563a,a40566a,a40567a,a40568a,a40571a,a40574a,a40575a,a40578a,a40581a,a40582a,a40583a,a40586a,a40589a,a40590a,a40593a,a40596a,a40597a,a40598a,a40601a,a40604a,a40605a,a40608a,a40611a,a40612a,a40613a,a40616a,a40619a,a40620a,a40623a,a40626a,a40627a,a40628a,a40631a,a40634a,a40635a,a40638a,a40641a,a40642a,a40643a,a40646a,a40649a,a40650a,a40653a,a40656a,a40657a,a40658a,a40661a,a40664a,a40665a,a40668a,a40671a,a40672a,a40673a,a40676a,a40679a,a40680a,a40683a,a40686a,a40687a,a40688a,a40691a,a40694a,a40695a,a40698a,a40701a,a40702a,a40703a,a40706a,a40709a,a40710a,a40713a,a40716a,a40717a,a40718a,a40721a,a40724a,a40725a,a40728a,a40731a,a40732a,a40733a,a40736a,a40739a,a40740a,a40743a,a40746a,a40747a,a40748a,a40751a,a40754a,a40755a,a40758a,a40761a,a40762a,a40763a,a40766a,a40769a,a40770a,a40773a,a40776a,a40777a,a40778a,a40781a,a40784a,a40785a,a40788a,a40791a,a40792a,a40793a,a40796a,a40799a,a40800a,a40803a,a40806a,a40807a,a40808a,a40811a,a40814a,a40815a,a40818a,a40821a,a40822a,a40823a,a40826a,a40829a,a40830a,a40833a,a40836a,a40837a,a40838a,a40841a,a40844a,a40845a,a40848a,a40851a,a40852a,a40853a,a40856a,a40859a,a40860a,a40863a,a40866a,a40867a,a40868a,a40871a,a40874a,a40875a,a40878a,a40881a,a40882a,a40883a,a40886a,a40889a,a40890a,a40893a,a40896a,a40897a,a40898a,a40901a,a40904a,a40905a,a40908a,a40911a,a40912a,a40913a,a40916a,a40919a,a40920a,a40923a,a40926a,a40927a,a40928a,a40931a,a40934a,a40935a,a40938a,a40941a,a40942a,a40943a,a40946a,a40949a,a40950a,a40953a,a40956a,a40957a,a40958a,a40961a,a40964a,a40965a,a40968a,a40971a,a40972a,a40973a,a40976a,a40979a,a40980a,a40983a,a40986a,a40987a,a40988a,a40991a,a40994a,a40995a,a40998a,a41001a,a41002a,a41003a,a41006a,a41009a,a41010a,a41013a,a41016a,a41017a,a41018a,a41021a,a41024a,a41025a,a41028a,a41031a,a41032a,a41033a,a41036a,a41039a,a41040a,a41043a,a41046a,a41047a,a41048a,a41051a,a41054a,a41055a,a41058a,a41061a,a41062a,a41063a,a41066a,a41069a,a41070a,a41073a,a41076a,a41077a,a41078a,a41081a,a41084a,a41085a,a41088a,a41091a,a41092a,a41093a,a41096a,a41099a,a41100a,a41103a,a41106a,a41107a,a41108a,a41111a,a41114a,a41115a,a41118a,a41121a,a41122a,a41123a,a41126a,a41129a,a41130a,a41133a,a41136a,a41137a,a41138a,a41141a,a41144a,a41145a,a41148a,a41151a,a41152a,a41153a,a41156a,a41159a,a41160a,a41163a,a41166a,a41167a,a41168a,a41171a,a41174a,a41175a,a41178a,a41181a,a41182a,a41183a,a41186a,a41189a,a41190a,a41193a,a41196a,a41197a,a41198a,a41201a,a41204a,a41205a,a41208a,a41211a,a41212a,a41213a,a41216a,a41219a,a41220a,a41223a,a41226a,a41227a,a41228a,a41231a,a41234a,a41235a,a41238a,a41241a,a41242a,a41243a,a41246a,a41249a,a41250a,a41253a,a41256a,a41257a,a41258a,a41261a,a41264a,a41265a,a41268a,a41271a,a41272a,a41273a,a41276a,a41279a,a41280a,a41283a,a41286a,a41287a,a41288a,a41291a,a41294a,a41295a,a41298a,a41301a,a41302a,a41303a,a41306a,a41309a,a41310a,a41313a,a41316a,a41317a,a41318a,a41321a,a41324a,a41325a,a41328a,a41331a,a41332a,a41333a,a41336a,a41339a,a41340a,a41343a,a41346a,a41347a,a41348a,a41351a,a41354a,a41355a,a41358a,a41361a,a41362a,a41363a,a41366a,a41369a,a41370a,a41373a,a41376a,a41377a,a41378a,a41381a,a41384a,a41385a,a41388a,a41391a,a41392a,a41393a,a41396a,a41399a,a41400a,a41403a,a41406a,a41407a,a41408a,a41411a,a41414a,a41415a,a41418a,a41421a,a41422a,a41423a,a41426a,a41429a,a41430a,a41433a,a41436a,a41437a,a41438a,a41441a,a41444a,a41445a,a41448a,a41451a,a41452a,a41453a,a41456a,a41459a,a41460a,a41463a,a41466a,a41467a,a41468a,a41471a,a41474a,a41475a,a41478a,a41481a,a41482a,a41483a,a41486a,a41489a,a41490a,a41493a,a41496a,a41497a,a41498a,a41501a,a41504a,a41505a,a41508a,a41511a,a41512a,a41513a,a41516a,a41519a,a41520a,a41523a,a41526a,a41527a,a41528a,a41531a,a41534a,a41535a,a41538a,a41541a,a41542a,a41543a,a41546a,a41549a,a41550a,a41553a,a41556a,a41557a,a41558a,a41561a,a41564a,a41565a,a41568a,a41571a,a41572a,a41573a,a41576a,a41579a,a41580a,a41583a,a41586a,a41587a,a41588a,a41591a,a41594a,a41595a,a41598a,a41601a,a41602a,a41603a,a41606a,a41609a,a41610a,a41613a,a41616a,a41617a,a41618a,a41621a,a41624a,a41625a,a41628a,a41631a,a41632a,a41633a,a41636a,a41639a,a41640a,a41643a,a41646a,a41647a,a41648a,a41651a,a41654a,a41655a,a41658a,a41661a,a41662a,a41663a,a41666a,a41669a,a41670a,a41673a,a41676a,a41677a,a41678a,a41681a,a41684a,a41685a,a41688a,a41691a,a41692a,a41693a,a41696a,a41699a,a41700a,a41703a,a41706a,a41707a,a41708a,a41711a,a41714a,a41715a,a41718a,a41721a,a41722a,a41723a,a41726a,a41729a,a41730a,a41733a,a41736a,a41737a,a41738a,a41741a,a41744a,a41745a,a41748a,a41751a,a41752a,a41753a,a41756a,a41759a,a41760a,a41763a,a41766a,a41767a,a41768a,a41771a,a41774a,a41775a,a41778a,a41781a,a41782a,a41783a,a41786a,a41789a,a41790a,a41793a,a41796a,a41797a,a41798a,a41801a,a41804a,a41805a,a41808a,a41811a,a41812a,a41813a,a41816a,a41819a,a41820a,a41823a,a41826a,a41827a,a41828a,a41831a,a41834a,a41835a,a41838a,a41841a,a41842a,a41843a,a41846a,a41849a,a41850a,a41853a,a41856a,a41857a,a41858a,a41861a,a41864a,a41865a,a41868a,a41871a,a41872a,a41873a,a41876a,a41879a,a41880a,a41883a,a41886a,a41887a,a41888a,a41891a,a41894a,a41895a,a41898a,a41901a,a41902a,a41903a,a41906a,a41909a,a41910a,a41913a,a41916a,a41917a,a41918a,a41921a,a41924a,a41925a,a41928a,a41931a,a41932a,a41933a,a41936a,a41939a,a41940a,a41943a,a41946a,a41947a,a41948a,a41951a,a41954a,a41955a,a41958a,a41961a,a41962a,a41963a,a41966a,a41969a,a41970a,a41973a,a41976a,a41977a,a41978a,a41981a,a41984a,a41985a,a41988a,a41991a,a41992a,a41993a,a41996a,a41999a,a42000a,a42003a,a42006a,a42007a,a42008a,a42011a,a42014a,a42015a,a42018a,a42021a,a42022a,a42023a,a42026a,a42029a,a42030a,a42033a,a42036a,a42037a,a42038a,a42041a,a42044a,a42045a,a42048a,a42051a,a42052a,a42053a,a42056a,a42059a,a42060a,a42063a,a42066a,a42067a,a42068a,a42071a,a42074a,a42075a,a42078a,a42081a,a42082a,a42083a,a42086a,a42089a,a42090a,a42093a,a42096a,a42097a,a42098a,a42101a,a42104a,a42105a,a42108a,a42111a,a42112a,a42113a,a42116a,a42119a,a42120a,a42123a,a42126a,a42127a,a42128a,a42131a,a42134a,a42135a,a42138a,a42141a,a42142a,a42143a,a42146a,a42149a,a42150a,a42153a,a42156a,a42157a,a42158a,a42161a,a42164a,a42165a,a42168a,a42171a,a42172a,a42173a,a42176a,a42179a,a42180a,a42183a,a42186a,a42187a,a42188a,a42191a,a42194a,a42195a,a42198a,a42201a,a42202a,a42203a,a42206a,a42209a,a42210a,a42213a,a42216a,a42217a,a42218a,a42221a,a42224a,a42225a,a42228a,a42231a,a42232a,a42233a,a42236a,a42239a,a42240a,a42243a,a42246a,a42247a,a42248a,a42251a,a42254a,a42255a,a42258a,a42261a,a42262a,a42263a,a42266a,a42269a,a42270a,a42273a,a42276a,a42277a,a42278a,a42281a,a42284a,a42285a,a42288a,a42291a,a42292a,a42293a,a42296a,a42299a,a42300a,a42303a,a42306a,a42307a,a42308a,a42311a,a42314a,a42315a,a42318a,a42321a,a42322a,a42323a,a42326a,a42329a,a42330a,a42333a,a42336a,a42337a,a42338a,a42341a,a42344a,a42345a,a42348a,a42351a,a42352a,a42353a,a42356a,a42359a,a42360a,a42363a,a42366a,a42367a,a42368a,a42371a,a42374a,a42375a,a42378a,a42381a,a42382a,a42383a,a42386a,a42389a,a42390a,a42393a,a42396a,a42397a,a42398a,a42401a,a42404a,a42405a,a42408a,a42411a,a42412a,a42413a,a42416a,a42419a,a42420a,a42423a,a42426a,a42427a,a42428a,a42431a,a42434a,a42435a,a42438a,a42441a,a42442a,a42443a,a42446a,a42449a,a42450a,a42453a,a42456a,a42457a,a42458a,a42461a,a42464a,a42465a,a42468a,a42471a,a42472a,a42473a,a42476a,a42479a,a42480a,a42483a,a42486a,a42487a,a42488a,a42491a,a42494a,a42495a,a42498a,a42501a,a42502a,a42503a,a42506a,a42509a,a42510a,a42513a,a42516a,a42517a,a42518a,a42521a,a42524a,a42525a,a42528a,a42531a,a42532a,a42533a,a42536a,a42539a,a42540a,a42543a,a42546a,a42547a,a42548a,a42551a,a42554a,a42555a,a42558a,a42561a,a42562a,a42563a,a42566a,a42569a,a42570a,a42573a,a42576a,a42577a,a42578a,a42581a,a42584a,a42585a,a42588a,a42591a,a42592a,a42593a,a42596a,a42599a,a42600a,a42603a,a42606a,a42607a,a42608a,a42611a,a42614a,a42615a,a42618a,a42621a,a42622a,a42623a,a42626a,a42629a,a42630a,a42633a,a42636a,a42637a,a42638a,a42641a,a42644a,a42645a,a42648a,a42651a,a42652a,a42653a,a42656a,a42659a,a42660a,a42663a,a42666a,a42667a,a42668a,a42671a,a42674a,a42675a,a42678a,a42681a,a42682a,a42683a,a42686a,a42689a,a42690a,a42693a,a42696a,a42697a,a42698a,a42701a,a42704a,a42705a,a42708a,a42711a,a42712a,a42713a,a42716a,a42719a,a42720a,a42723a,a42726a,a42727a,a42728a,a42731a,a42734a,a42735a,a42738a,a42741a,a42742a,a42743a,a42746a,a42749a,a42750a,a42753a,a42756a,a42757a,a42758a,a42761a,a42764a,a42765a,a42768a,a42771a,a42772a,a42773a,a42776a,a42779a,a42780a,a42783a,a42786a,a42787a,a42788a,a42791a,a42794a,a42795a,a42798a,a42801a,a42802a,a42803a,a42806a,a42809a,a42810a,a42813a,a42816a,a42817a,a42818a,a42821a,a42824a,a42825a,a42828a,a42831a,a42832a,a42833a,a42836a,a42839a,a42840a,a42843a,a42846a,a42847a,a42848a,a42851a,a42854a,a42855a,a42858a,a42861a,a42862a,a42863a,a42866a,a42869a,a42870a,a42873a,a42876a,a42877a,a42878a,a42881a,a42884a,a42885a,a42888a,a42891a,a42892a,a42893a,a42896a,a42899a,a42900a,a42903a,a42906a,a42907a,a42908a,a42911a,a42914a,a42915a,a42918a,a42921a,a42922a,a42923a,a42926a,a42929a,a42930a,a42933a,a42936a,a42937a,a42938a,a42941a,a42944a,a42945a,a42948a,a42951a,a42952a,a42953a,a42956a,a42959a,a42960a,a42963a,a42966a,a42967a,a42968a,a42971a,a42974a,a42975a,a42978a,a42981a,a42982a,a42983a,a42986a,a42989a,a42990a,a42993a,a42996a,a42997a,a42998a,a43001a,a43004a,a43005a,a43008a,a43011a,a43012a,a43013a,a43016a,a43019a,a43020a,a43023a,a43026a,a43027a,a43028a,a43031a,a43034a,a43035a,a43038a,a43041a,a43042a,a43043a,a43046a,a43049a,a43050a,a43053a,a43056a,a43057a,a43058a,a43061a,a43064a,a43065a,a43068a,a43071a,a43072a,a43073a,a43076a,a43079a,a43080a,a43083a,a43086a,a43087a,a43088a,a43091a,a43094a,a43095a,a43098a,a43101a,a43102a,a43103a,a43106a,a43109a,a43110a,a43113a,a43116a,a43117a,a43118a,a43121a,a43124a,a43125a,a43128a,a43131a,a43132a,a43133a,a43136a,a43139a,a43140a,a43143a,a43146a,a43147a,a43148a,a43151a,a43154a,a43155a,a43158a,a43161a,a43162a,a43163a,a43166a,a43169a,a43170a,a43173a,a43176a,a43177a,a43178a,a43181a,a43184a,a43185a,a43188a,a43191a,a43192a,a43193a,a43196a,a43199a,a43200a,a43203a,a43206a,a43207a,a43208a,a43211a,a43214a,a43215a,a43218a,a43221a,a43222a,a43223a,a43226a,a43229a,a43230a,a43233a,a43236a,a43237a,a43238a,a43241a,a43244a,a43245a,a43248a,a43251a,a43252a,a43253a,a43256a,a43259a,a43260a,a43263a,a43266a,a43267a,a43268a,a43271a,a43274a,a43275a,a43278a,a43281a,a43282a,a43283a,a43286a,a43289a,a43290a,a43293a,a43296a,a43297a,a43298a,a43301a,a43304a,a43305a,a43308a,a43311a,a43312a,a43313a,a43316a,a43319a,a43320a,a43323a,a43326a,a43327a,a43328a,a43331a,a43334a,a43335a,a43338a,a43341a,a43342a,a43343a,a43346a,a43349a,a43350a,a43353a,a43356a,a43357a,a43358a,a43361a,a43364a,a43365a,a43368a,a43371a,a43372a,a43373a,a43376a,a43379a,a43380a,a43383a,a43386a,a43387a,a43388a,a43391a,a43394a,a43395a,a43398a,a43401a,a43402a,a43403a,a43406a,a43409a,a43410a,a43413a,a43416a,a43417a,a43418a,a43421a,a43424a,a43425a,a43428a,a43431a,a43432a,a43433a,a43436a,a43439a,a43440a,a43443a,a43446a,a43447a,a43448a,a43451a,a43454a,a43455a,a43458a,a43461a,a43462a,a43463a,a43466a,a43469a,a43470a,a43473a,a43476a,a43477a,a43478a,a43481a,a43484a,a43485a,a43488a,a43491a,a43492a,a43493a,a43496a,a43499a,a43500a,a43503a,a43506a,a43507a,a43508a,a43511a,a43514a,a43515a,a43518a,a43521a,a43522a,a43523a,a43526a,a43529a,a43530a,a43533a,a43536a,a43537a,a43538a,a43541a,a43544a,a43545a,a43548a,a43551a,a43552a,a43553a,a43556a,a43559a,a43560a,a43563a,a43566a,a43567a,a43568a,a43571a,a43574a,a43575a,a43578a,a43581a,a43582a,a43583a,a43586a,a43589a,a43590a,a43593a,a43596a,a43597a,a43598a,a43601a,a43604a,a43605a,a43608a,a43611a,a43612a,a43613a,a43616a,a43619a,a43620a,a43623a,a43626a,a43627a,a43628a,a43631a,a43634a,a43635a,a43638a,a43641a,a43642a,a43643a,a43646a,a43649a,a43650a,a43653a,a43656a,a43657a,a43658a,a43661a,a43664a,a43665a,a43668a,a43671a,a43672a,a43673a,a43676a,a43679a,a43680a,a43683a,a43686a,a43687a,a43688a,a43691a,a43694a,a43695a,a43698a,a43701a,a43702a,a43703a,a43706a,a43709a,a43710a,a43713a,a43716a,a43717a,a43718a,a43721a,a43724a,a43725a,a43728a,a43731a,a43732a,a43733a,a43736a,a43739a,a43740a,a43743a,a43746a,a43747a,a43748a,a43751a,a43754a,a43755a,a43758a,a43761a,a43762a,a43763a,a43766a,a43769a,a43770a,a43773a,a43776a,a43777a,a43778a,a43781a,a43784a,a43785a,a43788a,a43791a,a43792a,a43793a,a43796a,a43799a,a43800a,a43803a,a43806a,a43807a,a43808a,a43811a,a43814a,a43815a,a43818a,a43821a,a43822a,a43823a,a43826a,a43829a,a43830a,a43833a,a43836a,a43837a,a43838a,a43841a,a43844a,a43845a,a43848a,a43851a,a43852a,a43853a,a43856a,a43859a,a43860a,a43863a,a43866a,a43867a,a43868a,a43871a,a43874a,a43875a,a43878a,a43881a,a43882a,a43883a,a43886a,a43889a,a43890a,a43893a,a43896a,a43897a,a43898a,a43901a,a43904a,a43905a,a43908a,a43911a,a43912a,a43913a,a43916a,a43919a,a43920a,a43923a,a43926a,a43927a,a43928a,a43931a,a43934a,a43935a,a43938a,a43941a,a43942a,a43943a,a43946a,a43949a,a43950a,a43953a,a43956a,a43957a,a43958a,a43961a,a43964a,a43965a,a43968a,a43971a,a43972a,a43973a,a43976a,a43979a,a43980a,a43983a,a43986a,a43987a,a43988a,a43991a,a43994a,a43995a,a43998a,a44001a,a44002a,a44003a,a44006a,a44009a,a44010a,a44013a,a44016a,a44017a,a44018a,a44021a,a44024a,a44025a,a44028a,a44031a,a44032a,a44033a,a44036a,a44039a,a44040a,a44043a,a44046a,a44047a,a44048a,a44051a,a44054a,a44055a,a44058a,a44061a,a44062a,a44063a,a44066a,a44069a,a44070a,a44073a,a44076a,a44077a,a44078a,a44081a,a44084a,a44085a,a44088a,a44091a,a44092a,a44093a,a44096a,a44099a,a44100a,a44103a,a44106a,a44107a,a44108a,a44111a,a44114a,a44115a,a44118a,a44121a,a44122a,a44123a,a44126a,a44129a,a44130a,a44133a,a44136a,a44137a,a44138a,a44141a,a44144a,a44145a,a44148a,a44151a,a44152a,a44153a,a44156a,a44159a,a44160a,a44163a,a44166a,a44167a,a44168a,a44171a,a44174a,a44175a,a44178a,a44181a,a44182a,a44183a,a44186a,a44189a,a44190a,a44193a,a44196a,a44197a,a44198a,a44201a,a44204a,a44205a,a44208a,a44211a,a44212a,a44213a,a44216a,a44219a,a44220a,a44223a,a44226a,a44227a,a44228a,a44231a,a44234a,a44235a,a44238a,a44241a,a44242a,a44243a,a44246a,a44249a,a44250a,a44253a,a44256a,a44257a,a44258a,a44261a,a44264a,a44265a,a44268a,a44271a,a44272a,a44273a,a44276a,a44279a,a44280a,a44283a,a44286a,a44287a,a44288a,a44291a,a44294a,a44295a,a44298a,a44301a,a44302a,a44303a,a44306a,a44309a,a44310a,a44313a,a44316a,a44317a,a44318a,a44321a,a44324a,a44325a,a44328a,a44331a,a44332a,a44333a,a44336a,a44339a,a44340a,a44343a,a44346a,a44347a,a44348a,a44351a,a44354a,a44355a,a44358a,a44361a,a44362a,a44363a,a44366a,a44369a,a44370a,a44373a,a44376a,a44377a,a44378a,a44381a,a44384a,a44385a,a44388a,a44391a,a44392a,a44393a,a44396a,a44399a,a44400a,a44403a,a44406a,a44407a,a44408a,a44411a,a44414a,a44415a,a44418a,a44421a,a44422a,a44423a,a44426a,a44429a,a44430a,a44433a,a44436a,a44437a,a44438a,a44441a,a44444a,a44445a,a44448a,a44451a,a44452a,a44453a,a44456a,a44459a,a44460a,a44463a,a44466a,a44467a,a44468a,a44471a,a44474a,a44475a,a44478a,a44481a,a44482a,a44483a,a44486a,a44489a,a44490a,a44493a,a44496a,a44497a,a44498a,a44501a,a44504a,a44505a,a44508a,a44511a,a44512a,a44513a,a44516a,a44519a,a44520a,a44523a,a44526a,a44527a,a44528a,a44531a,a44534a,a44535a,a44538a,a44541a,a44542a,a44543a,a44546a,a44549a,a44550a,a44553a,a44556a,a44557a,a44558a,a44561a,a44564a,a44565a,a44568a,a44571a,a44572a,a44573a,a44576a,a44579a,a44580a,a44583a,a44586a,a44587a,a44588a,a44591a,a44594a,a44595a,a44598a,a44601a,a44602a,a44603a,a44606a,a44609a,a44610a,a44613a,a44616a,a44617a,a44618a,a44621a,a44624a,a44625a,a44628a,a44631a,a44632a,a44633a,a44636a,a44639a,a44640a,a44643a,a44646a,a44647a,a44648a,a44651a,a44654a,a44655a,a44658a,a44661a,a44662a,a44663a,a44666a,a44669a,a44670a,a44673a,a44676a,a44677a,a44678a,a44681a,a44684a,a44685a,a44688a,a44691a,a44692a,a44693a,a44696a,a44699a,a44700a,a44703a,a44706a,a44707a,a44708a,a44711a,a44714a,a44715a,a44718a,a44721a,a44722a,a44723a,a44726a,a44729a,a44730a,a44733a,a44736a,a44737a,a44738a,a44741a,a44744a,a44745a,a44748a,a44751a,a44752a,a44753a,a44756a,a44759a,a44760a,a44763a,a44766a,a44767a,a44768a,a44771a,a44774a,a44775a,a44778a,a44781a,a44782a,a44783a,a44786a,a44789a,a44790a,a44793a,a44796a,a44797a,a44798a,a44801a,a44804a,a44805a,a44808a,a44811a,a44812a,a44813a,a44816a,a44819a,a44820a,a44823a,a44826a,a44827a,a44828a,a44831a,a44834a,a44835a,a44838a,a44841a,a44842a,a44843a,a44846a,a44849a,a44850a,a44853a,a44856a,a44857a,a44858a,a44861a,a44864a,a44865a,a44868a,a44871a,a44872a,a44873a,a44876a,a44879a,a44880a,a44883a,a44886a,a44887a,a44888a,a44891a,a44894a,a44895a,a44898a,a44901a,a44902a,a44903a,a44906a,a44909a,a44910a,a44913a,a44916a,a44917a,a44918a,a44921a,a44924a,a44925a,a44928a,a44931a,a44932a,a44933a,a44936a,a44939a,a44940a,a44943a,a44946a,a44947a,a44948a,a44951a,a44954a,a44955a,a44958a,a44961a,a44962a,a44963a,a44966a,a44969a,a44970a,a44973a,a44976a,a44977a,a44978a,a44981a,a44984a,a44985a,a44988a,a44991a,a44992a,a44993a,a44996a,a44999a,a45000a,a45003a,a45006a,a45007a,a45008a,a45011a,a45014a,a45015a,a45018a,a45021a,a45022a,a45023a,a45026a,a45029a,a45030a,a45033a,a45036a,a45037a,a45038a,a45041a,a45044a,a45045a,a45048a,a45051a,a45052a,a45053a,a45056a,a45059a,a45060a,a45063a,a45066a,a45067a,a45068a,a45071a,a45074a,a45075a,a45078a,a45081a,a45082a,a45083a,a45086a,a45089a,a45090a,a45093a,a45096a,a45097a,a45098a,a45101a,a45104a,a45105a,a45108a,a45111a,a45112a,a45113a,a45116a,a45119a,a45120a,a45123a,a45126a,a45127a,a45128a,a45131a,a45134a,a45135a,a45138a,a45141a,a45142a,a45143a,a45146a,a45149a,a45150a,a45153a,a45156a,a45157a,a45158a,a45161a,a45164a,a45165a,a45168a,a45171a,a45172a,a45173a,a45176a,a45179a,a45180a,a45183a,a45186a,a45187a,a45188a,a45191a,a45194a,a45195a,a45198a,a45201a,a45202a,a45203a,a45206a,a45209a,a45210a,a45213a,a45216a,a45217a,a45218a,a45221a,a45224a,a45225a,a45228a,a45231a,a45232a,a45233a,a45236a,a45239a,a45240a,a45243a,a45246a,a45247a,a45248a,a45251a,a45254a,a45255a,a45258a,a45261a,a45262a,a45263a,a45266a,a45269a,a45270a,a45273a,a45276a,a45277a,a45278a,a45281a,a45284a,a45285a,a45288a,a45291a,a45292a,a45293a,a45296a,a45299a,a45300a,a45303a,a45306a,a45307a,a45308a,a45311a,a45314a,a45315a,a45318a,a45321a,a45322a,a45323a,a45326a,a45329a,a45330a,a45333a,a45336a,a45337a,a45338a,a45341a,a45344a,a45345a,a45348a,a45351a,a45352a,a45353a,a45356a,a45359a,a45360a,a45363a,a45366a,a45367a,a45368a,a45371a,a45374a,a45375a,a45378a,a45381a,a45382a,a45383a,a45386a,a45389a,a45390a,a45393a,a45396a,a45397a,a45398a,a45401a,a45404a,a45405a,a45408a,a45411a,a45412a,a45413a,a45416a,a45419a,a45420a,a45423a,a45426a,a45427a,a45428a,a45431a,a45434a,a45435a,a45438a,a45441a,a45442a,a45443a,a45446a,a45449a,a45450a,a45453a,a45456a,a45457a,a45458a,a45461a,a45464a,a45465a,a45468a,a45471a,a45472a,a45473a,a45476a,a45479a,a45480a,a45483a,a45486a,a45487a,a45488a,a45491a,a45494a,a45495a,a45498a,a45501a,a45502a,a45503a,a45506a,a45509a,a45510a,a45513a,a45516a,a45517a,a45518a,a45521a,a45524a,a45525a,a45528a,a45531a,a45532a,a45533a,a45536a,a45539a,a45540a,a45543a,a45546a,a45547a,a45548a,a45551a,a45554a,a45555a,a45558a,a45561a,a45562a,a45563a,a45566a,a45569a,a45570a,a45573a,a45576a,a45577a,a45578a,a45581a,a45584a,a45585a,a45588a,a45591a,a45592a,a45593a,a45596a,a45599a,a45600a,a45603a,a45606a,a45607a,a45608a,a45611a,a45614a,a45615a,a45618a,a45621a,a45622a,a45623a,a45626a,a45629a,a45630a,a45633a,a45636a,a45637a,a45638a,a45641a,a45644a,a45645a,a45648a,a45651a,a45652a,a45653a,a45656a,a45659a,a45660a,a45663a,a45666a,a45667a,a45668a,a45671a,a45674a,a45675a,a45678a,a45681a,a45682a,a45683a,a45686a,a45689a,a45690a,a45693a,a45696a,a45697a,a45698a,a45701a,a45704a,a45705a,a45708a,a45711a,a45712a,a45713a,a45716a,a45719a,a45720a,a45723a,a45726a,a45727a,a45728a,a45731a,a45734a,a45735a,a45738a,a45741a,a45742a,a45743a,a45746a,a45749a,a45750a,a45753a,a45756a,a45757a,a45758a,a45761a,a45764a,a45765a,a45768a,a45771a,a45772a,a45773a,a45776a,a45779a,a45780a,a45783a,a45786a,a45787a,a45788a,a45791a,a45794a,a45795a,a45798a,a45801a,a45802a,a45803a,a45806a,a45809a,a45810a,a45813a,a45816a,a45817a,a45818a,a45821a,a45824a,a45825a,a45828a,a45831a,a45832a,a45833a,a45836a,a45839a,a45840a,a45843a,a45846a,a45847a,a45848a,a45851a,a45854a,a45855a,a45858a,a45861a,a45862a,a45863a,a45866a,a45869a,a45870a,a45873a,a45876a,a45877a,a45878a,a45881a,a45884a,a45885a,a45888a,a45891a,a45892a,a45893a,a45896a,a45899a,a45900a,a45903a,a45906a,a45907a,a45908a,a45911a,a45914a,a45915a,a45918a,a45921a,a45922a,a45923a,a45926a,a45929a,a45930a,a45933a,a45936a,a45937a,a45938a,a45941a,a45944a,a45945a,a45948a,a45951a,a45952a,a45953a,a45956a,a45959a,a45960a,a45963a,a45966a,a45967a,a45968a,a45971a,a45974a,a45975a,a45978a,a45981a,a45982a,a45983a,a45986a,a45989a,a45990a,a45993a,a45996a,a45997a,a45998a,a46001a,a46004a,a46005a,a46008a,a46011a,a46012a,a46013a,a46016a,a46019a,a46020a,a46023a,a46026a,a46027a,a46028a,a46031a,a46034a,a46035a,a46038a,a46041a,a46042a,a46043a,a46046a,a46049a,a46050a,a46053a,a46056a,a46057a,a46058a,a46061a,a46064a,a46065a,a46068a,a46071a,a46072a,a46073a,a46076a,a46079a,a46080a,a46083a,a46086a,a46087a,a46088a,a46091a,a46094a,a46095a,a46098a,a46101a,a46102a,a46103a,a46106a,a46109a,a46110a,a46113a,a46116a,a46117a,a46118a,a46121a,a46124a,a46125a,a46128a,a46131a,a46132a,a46133a,a46136a,a46139a,a46140a,a46143a,a46146a,a46147a,a46148a,a46151a,a46154a,a46155a,a46158a,a46161a,a46162a,a46163a,a46166a,a46169a,a46170a,a46173a,a46176a,a46177a,a46178a,a46181a,a46184a,a46185a,a46188a,a46191a,a46192a,a46193a,a46196a,a46199a,a46200a,a46203a,a46206a,a46207a,a46208a,a46211a,a46214a,a46215a,a46218a,a46221a,a46222a,a46223a,a46226a,a46229a,a46230a,a46233a,a46236a,a46237a,a46238a,a46241a,a46244a,a46245a,a46248a,a46251a,a46252a,a46253a,a46256a,a46259a,a46260a,a46263a,a46266a,a46267a,a46268a,a46271a,a46274a,a46275a,a46278a,a46281a,a46282a,a46283a,a46286a,a46289a,a46290a,a46293a,a46296a,a46297a,a46298a,a46301a,a46304a,a46305a,a46308a,a46311a,a46312a,a46313a,a46316a,a46319a,a46320a,a46323a,a46326a,a46327a,a46328a,a46331a,a46334a,a46335a,a46338a,a46341a,a46342a,a46343a,a46346a,a46349a,a46350a,a46353a,a46356a,a46357a,a46358a,a46361a,a46364a,a46365a,a46368a,a46371a,a46372a,a46373a,a46376a,a46379a,a46380a,a46383a,a46386a,a46387a,a46388a,a46391a,a46394a,a46395a,a46398a,a46401a,a46402a,a46403a,a46406a,a46409a,a46410a,a46413a,a46416a,a46417a,a46418a,a46421a,a46424a,a46425a,a46428a,a46431a,a46432a,a46433a,a46436a,a46439a,a46440a,a46443a,a46446a,a46447a,a46448a,a46451a,a46454a,a46455a,a46458a,a46461a,a46462a,a46463a,a46466a,a46469a,a46470a,a46473a,a46476a,a46477a,a46478a,a46481a,a46484a,a46485a,a46488a,a46491a,a46492a,a46493a,a46496a,a46499a,a46500a,a46503a,a46506a,a46507a,a46508a,a46511a,a46514a,a46515a,a46518a,a46521a,a46522a,a46523a,a46526a,a46529a,a46530a,a46533a,a46536a,a46537a,a46538a,a46541a,a46544a,a46545a,a46548a,a46551a,a46552a,a46553a,a46556a,a46559a,a46560a,a46563a,a46566a,a46567a,a46568a,a46571a,a46574a,a46575a,a46578a,a46581a,a46582a,a46583a,a46586a,a46589a,a46590a,a46593a,a46596a,a46597a,a46598a,a46601a,a46604a,a46605a,a46608a,a46611a,a46612a,a46613a,a46616a,a46619a,a46620a,a46623a,a46626a,a46627a,a46628a,a46631a,a46634a,a46635a,a46638a,a46641a,a46642a,a46643a,a46646a,a46649a,a46650a,a46653a,a46656a,a46657a,a46658a,a46661a,a46664a,a46665a,a46668a,a46671a,a46672a,a46673a,a46676a,a46679a,a46680a,a46683a,a46686a,a46687a,a46688a,a46691a,a46694a,a46695a,a46698a,a46701a,a46702a,a46703a,a46706a,a46709a,a46710a,a46713a,a46716a,a46717a,a46718a,a46721a,a46724a,a46725a,a46728a,a46731a,a46732a,a46733a,a46736a,a46739a,a46740a,a46743a,a46746a,a46747a,a46748a,a46751a,a46754a,a46755a,a46758a,a46761a,a46762a,a46763a,a46766a,a46769a,a46770a,a46773a,a46776a,a46777a,a46778a,a46781a,a46784a,a46785a,a46788a,a46791a,a46792a,a46793a,a46796a,a46799a,a46800a,a46803a,a46806a,a46807a,a46808a,a46811a,a46814a,a46815a,a46818a,a46821a,a46822a,a46823a,a46826a,a46829a,a46830a,a46833a,a46836a,a46837a,a46838a,a46841a,a46844a,a46845a,a46848a,a46851a,a46852a,a46853a,a46856a,a46859a,a46860a,a46863a,a46866a,a46867a,a46868a,a46871a,a46874a,a46875a,a46878a,a46881a,a46882a,a46883a,a46886a,a46889a,a46890a,a46893a,a46896a,a46897a,a46898a,a46901a,a46904a,a46905a,a46908a,a46911a,a46912a,a46913a,a46916a,a46919a,a46920a,a46923a,a46926a,a46927a,a46928a,a46931a,a46934a,a46935a,a46938a,a46941a,a46942a,a46943a,a46946a,a46949a,a46950a,a46953a,a46956a,a46957a,a46958a,a46961a,a46964a,a46965a,a46968a,a46971a,a46972a,a46973a,a46976a,a46979a,a46980a,a46983a,a46986a,a46987a,a46988a,a46991a,a46994a,a46995a,a46998a,a47001a,a47002a,a47003a,a47006a,a47009a,a47010a,a47013a,a47016a,a47017a,a47018a,a47021a,a47024a,a47025a,a47028a,a47031a,a47032a,a47033a,a47036a,a47039a,a47040a,a47043a,a47046a,a47047a,a47048a,a47051a,a47054a,a47055a,a47058a,a47061a,a47062a,a47063a,a47066a,a47069a,a47070a,a47073a,a47076a,a47077a,a47078a,a47081a,a47084a,a47085a,a47088a,a47091a,a47092a,a47093a,a47096a,a47099a,a47100a,a47103a,a47106a,a47107a,a47108a,a47111a,a47114a,a47115a,a47118a,a47121a,a47122a,a47123a,a47126a,a47129a,a47130a,a47133a,a47136a,a47137a,a47138a,a47141a,a47144a,a47145a,a47148a,a47151a,a47152a,a47153a,a47156a,a47159a,a47160a,a47163a,a47166a,a47167a,a47168a,a47171a,a47174a,a47175a,a47178a,a47181a,a47182a,a47183a,a47186a,a47189a,a47190a,a47193a,a47196a,a47197a,a47198a,a47201a,a47204a,a47205a,a47208a,a47211a,a47212a,a47213a,a47216a,a47219a,a47220a,a47223a,a47226a,a47227a,a47228a,a47231a,a47234a,a47235a,a47238a,a47241a,a47242a,a47243a,a47246a,a47249a,a47250a,a47253a,a47256a,a47257a,a47258a,a47261a,a47264a,a47265a,a47268a,a47271a,a47272a,a47273a,a47276a,a47279a,a47280a,a47283a,a47286a,a47287a,a47288a,a47291a,a47294a,a47295a,a47298a,a47301a,a47302a,a47303a,a47306a,a47309a,a47310a,a47313a,a47316a,a47317a,a47318a,a47321a,a47324a,a47325a,a47328a,a47331a,a47332a,a47333a,a47336a,a47339a,a47340a,a47343a,a47346a,a47347a,a47348a,a47351a,a47354a,a47355a,a47358a,a47361a,a47362a,a47363a,a47366a,a47369a,a47370a,a47373a,a47376a,a47377a,a47378a,a47381a,a47384a,a47385a,a47388a,a47391a,a47392a,a47393a,a47396a,a47399a,a47400a,a47403a,a47406a,a47407a,a47408a,a47411a,a47414a,a47415a,a47418a,a47421a,a47422a,a47423a,a47426a,a47429a,a47430a,a47433a,a47436a,a47437a,a47438a,a47441a,a47444a,a47445a,a47448a,a47451a,a47452a,a47453a,a47456a,a47459a,a47460a,a47463a,a47466a,a47467a,a47468a,a47471a,a47474a,a47475a,a47478a,a47481a,a47482a,a47483a,a47486a,a47489a,a47490a,a47493a,a47496a,a47497a,a47498a,a47501a,a47504a,a47505a,a47508a,a47511a,a47512a,a47513a,a47516a,a47519a,a47520a,a47523a,a47526a,a47527a,a47528a,a47531a,a47534a,a47535a,a47538a,a47541a,a47542a,a47543a,a47546a,a47549a,a47550a,a47553a,a47556a,a47557a,a47558a,a47561a,a47564a,a47565a,a47568a,a47571a,a47572a,a47573a,a47576a,a47579a,a47580a,a47583a,a47586a,a47587a,a47588a,a47591a,a47594a,a47595a,a47598a,a47601a,a47602a,a47603a,a47606a,a47609a,a47610a,a47613a,a47616a,a47617a,a47618a,a47621a,a47624a,a47625a,a47628a,a47631a,a47632a,a47633a,a47636a,a47639a,a47640a,a47643a,a47646a,a47647a,a47648a,a47651a,a47654a,a47655a,a47658a,a47661a,a47662a,a47663a,a47666a,a47669a,a47670a,a47673a,a47676a,a47677a,a47678a,a47681a,a47684a,a47685a,a47688a,a47691a,a47692a,a47693a,a47696a,a47699a,a47700a,a47703a,a47706a,a47707a,a47708a,a47711a,a47714a,a47715a,a47718a,a47721a,a47722a,a47723a,a47726a,a47729a,a47730a,a47733a,a47736a,a47737a,a47738a,a47741a,a47744a,a47745a,a47748a,a47751a,a47752a,a47753a,a47756a,a47759a,a47760a,a47763a,a47766a,a47767a,a47768a,a47771a,a47774a,a47775a,a47778a,a47781a,a47782a,a47783a,a47786a,a47789a,a47790a,a47793a,a47796a,a47797a,a47798a,a47801a,a47804a,a47805a,a47808a,a47811a,a47812a,a47813a,a47816a,a47819a,a47820a,a47823a,a47826a,a47827a,a47828a,a47831a,a47834a,a47835a,a47838a,a47841a,a47842a,a47843a,a47846a,a47849a,a47850a,a47853a,a47856a,a47857a,a47858a,a47861a,a47864a,a47865a,a47868a,a47871a,a47872a,a47873a,a47876a,a47879a,a47880a,a47883a,a47886a,a47887a,a47888a,a47891a,a47894a,a47895a,a47898a,a47901a,a47902a,a47903a,a47906a,a47909a,a47910a,a47913a,a47916a,a47917a,a47918a,a47921a,a47924a,a47925a,a47928a,a47931a,a47932a,a47933a,a47936a,a47939a,a47940a,a47943a,a47946a,a47947a,a47948a,a47951a,a47954a,a47955a,a47958a,a47961a,a47962a,a47963a,a47966a,a47969a,a47970a,a47973a,a47976a,a47977a,a47978a,a47981a,a47984a,a47985a,a47988a,a47991a,a47992a,a47993a,a47996a,a47999a,a48000a,a48003a,a48006a,a48007a,a48008a,a48011a,a48014a,a48015a,a48018a,a48021a,a48022a,a48023a,a48026a,a48029a,a48030a,a48033a,a48036a,a48037a,a48038a,a48041a,a48044a,a48045a,a48048a,a48051a,a48052a,a48053a,a48056a,a48059a,a48060a,a48063a,a48066a,a48067a,a48068a,a48071a,a48074a,a48075a,a48078a,a48081a,a48082a,a48083a,a48086a,a48089a,a48090a,a48093a,a48096a,a48097a,a48098a,a48101a,a48104a,a48105a,a48108a,a48111a,a48112a,a48113a,a48116a,a48119a,a48120a,a48123a,a48126a,a48127a,a48128a,a48131a,a48134a,a48135a,a48138a,a48141a,a48142a,a48143a,a48146a,a48149a,a48150a,a48153a,a48156a,a48157a,a48158a,a48161a,a48164a,a48165a,a48168a,a48171a,a48172a,a48173a,a48176a,a48179a,a48180a,a48183a,a48186a,a48187a,a48188a,a48191a,a48194a,a48195a,a48198a,a48201a,a48202a,a48203a,a48206a,a48209a,a48210a,a48213a,a48216a,a48217a,a48218a,a48221a,a48224a,a48225a,a48228a,a48231a,a48232a,a48233a,a48236a,a48239a,a48240a,a48243a,a48246a,a48247a,a48248a,a48251a,a48254a,a48255a,a48258a,a48261a,a48262a,a48263a,a48266a,a48269a,a48270a,a48273a,a48276a,a48277a,a48278a,a48281a,a48284a,a48285a,a48288a,a48291a,a48292a,a48293a,a48296a,a48299a,a48300a,a48303a,a48306a,a48307a,a48308a,a48311a,a48314a,a48315a,a48318a,a48321a,a48322a,a48323a,a48326a,a48329a,a48330a,a48333a,a48336a,a48337a,a48338a,a48341a,a48344a,a48345a,a48348a,a48351a,a48352a,a48353a,a48356a,a48359a,a48360a,a48363a,a48366a,a48367a,a48368a,a48371a,a48374a,a48375a,a48378a,a48381a,a48382a,a48383a,a48386a,a48389a,a48390a,a48393a,a48396a,a48397a,a48398a,a48401a,a48404a,a48405a,a48408a,a48411a,a48412a,a48413a,a48416a,a48419a,a48420a,a48423a,a48426a,a48427a,a48428a,a48431a,a48434a,a48435a,a48438a,a48441a,a48442a,a48443a,a48446a,a48449a,a48450a,a48453a,a48456a,a48457a,a48458a,a48461a,a48464a,a48465a,a48468a,a48471a,a48472a,a48473a,a48476a,a48479a,a48480a,a48483a,a48486a,a48487a,a48488a,a48491a,a48494a,a48495a,a48498a,a48501a,a48502a,a48503a,a48506a,a48509a,a48510a,a48513a,a48516a,a48517a,a48518a,a48521a,a48524a,a48525a,a48528a,a48531a,a48532a,a48533a,a48536a,a48539a,a48540a,a48543a,a48546a,a48547a,a48548a,a48551a,a48554a,a48555a,a48558a,a48561a,a48562a,a48563a,a48566a,a48569a,a48570a,a48573a,a48576a,a48577a,a48578a,a48581a,a48584a,a48585a,a48588a,a48591a,a48592a,a48593a,a48596a,a48599a,a48600a,a48603a,a48606a,a48607a,a48608a,a48611a,a48614a,a48615a,a48618a,a48621a,a48622a,a48623a,a48626a,a48629a,a48630a,a48633a,a48636a,a48637a,a48638a,a48641a,a48644a,a48645a,a48648a,a48651a,a48652a,a48653a,a48656a,a48659a,a48660a,a48663a,a48666a,a48667a,a48668a,a48671a,a48674a,a48675a,a48678a,a48681a,a48682a,a48683a,a48686a,a48689a,a48690a,a48693a,a48696a,a48697a,a48698a,a48701a,a48704a,a48705a,a48708a,a48711a,a48712a,a48713a,a48716a,a48719a,a48720a,a48723a,a48726a,a48727a,a48728a,a48731a,a48734a,a48735a,a48738a,a48741a,a48742a,a48743a,a48746a,a48749a,a48750a,a48753a,a48756a,a48757a,a48758a,a48761a,a48764a,a48765a,a48768a,a48771a,a48772a,a48773a,a48776a,a48779a,a48780a,a48783a,a48786a,a48787a,a48788a,a48791a,a48794a,a48795a,a48798a,a48801a,a48802a,a48803a,a48806a,a48809a,a48810a,a48813a,a48816a,a48817a,a48818a,a48821a,a48824a,a48825a,a48828a,a48831a,a48832a,a48833a,a48836a,a48839a,a48840a,a48843a,a48846a,a48847a,a48848a,a48851a,a48854a,a48855a,a48858a,a48861a,a48862a,a48863a,a48866a,a48869a,a48870a,a48873a,a48876a,a48877a,a48878a,a48881a,a48884a,a48885a,a48888a,a48891a,a48892a,a48893a,a48896a,a48899a,a48900a,a48903a,a48906a,a48907a,a48908a,a48911a,a48914a,a48915a,a48918a,a48921a,a48922a,a48923a,a48926a,a48929a,a48930a,a48933a,a48936a,a48937a,a48938a,a48941a,a48944a,a48945a,a48948a,a48951a,a48952a,a48953a,a48956a,a48959a,a48960a,a48963a,a48966a,a48967a,a48968a,a48971a,a48974a,a48975a,a48978a,a48981a,a48982a,a48983a,a48986a,a48989a,a48990a,a48993a,a48996a,a48997a,a48998a,a49001a,a49004a,a49005a,a49008a,a49011a,a49012a,a49013a,a49016a,a49019a,a49020a,a49023a,a49026a,a49027a,a49028a,a49031a,a49034a,a49035a,a49038a,a49041a,a49042a,a49043a,a49046a,a49049a,a49050a,a49053a,a49056a,a49057a,a49058a,a49061a,a49064a,a49065a,a49068a,a49071a,a49072a,a49073a,a49076a,a49079a,a49080a,a49083a,a49086a,a49087a,a49088a,a49091a,a49094a,a49095a,a49098a,a49101a,a49102a,a49103a,a49106a,a49109a,a49110a,a49113a,a49116a,a49117a,a49118a,a49121a,a49124a,a49125a,a49128a,a49131a,a49132a,a49133a,a49136a,a49139a,a49140a,a49143a,a49146a,a49147a,a49148a,a49151a,a49154a,a49155a,a49158a,a49161a,a49162a,a49163a,a49166a,a49169a,a49170a,a49173a,a49176a,a49177a,a49178a,a49181a,a49184a,a49185a,a49188a,a49191a,a49192a,a49193a,a49196a,a49199a,a49200a,a49203a,a49206a,a49207a,a49208a,a49211a,a49214a,a49215a,a49218a,a49221a,a49222a,a49223a,a49226a,a49229a,a49230a,a49233a,a49236a,a49237a,a49238a,a49241a,a49244a,a49245a,a49248a,a49251a,a49252a,a49253a,a49256a,a49259a,a49260a,a49263a,a49266a,a49267a,a49268a,a49271a,a49274a,a49275a,a49278a,a49281a,a49282a,a49283a,a49286a,a49289a,a49290a,a49293a,a49296a,a49297a,a49298a,a49301a,a49304a,a49305a,a49308a,a49311a,a49312a,a49313a,a49316a,a49319a,a49320a,a49323a,a49326a,a49327a,a49328a,a49331a,a49334a,a49335a,a49338a,a49341a,a49342a,a49343a,a49346a,a49349a,a49350a,a49353a,a49356a,a49357a,a49358a,a49361a,a49364a,a49365a,a49368a,a49371a,a49372a,a49373a,a49376a,a49379a,a49380a,a49383a,a49386a,a49387a,a49388a,a49391a,a49394a,a49395a,a49398a,a49401a,a49402a,a49403a,a49406a,a49409a,a49410a,a49413a,a49416a,a49417a,a49418a,a49421a,a49424a,a49425a,a49428a,a49431a,a49432a,a49433a,a49436a,a49439a,a49440a,a49443a,a49446a,a49447a,a49448a,a49451a,a49454a,a49455a,a49458a,a49461a,a49462a,a49463a,a49466a,a49469a,a49470a,a49473a,a49476a,a49477a,a49478a,a49481a,a49484a,a49485a,a49488a,a49491a,a49492a,a49493a,a49496a,a49499a,a49500a,a49503a,a49506a,a49507a,a49508a,a49511a,a49514a,a49515a,a49518a,a49521a,a49522a,a49523a,a49526a,a49529a,a49530a,a49533a,a49536a,a49537a,a49538a: std_logic;
begin

A42 <=( a5254a ) or ( a3503a );
 a1a <=( a49538a  and  a49523a );
 a2a <=( a49508a  and  a49493a );
 a3a <=( a49478a  and  a49463a );
 a4a <=( a49448a  and  a49433a );
 a5a <=( a49418a  and  a49403a );
 a6a <=( a49388a  and  a49373a );
 a7a <=( a49358a  and  a49343a );
 a8a <=( a49328a  and  a49313a );
 a9a <=( a49298a  and  a49283a );
 a10a <=( a49268a  and  a49253a );
 a11a <=( a49238a  and  a49223a );
 a12a <=( a49208a  and  a49193a );
 a13a <=( a49178a  and  a49163a );
 a14a <=( a49148a  and  a49133a );
 a15a <=( a49118a  and  a49103a );
 a16a <=( a49088a  and  a49073a );
 a17a <=( a49058a  and  a49043a );
 a18a <=( a49028a  and  a49013a );
 a19a <=( a48998a  and  a48983a );
 a20a <=( a48968a  and  a48953a );
 a21a <=( a48938a  and  a48923a );
 a22a <=( a48908a  and  a48893a );
 a23a <=( a48878a  and  a48863a );
 a24a <=( a48848a  and  a48833a );
 a25a <=( a48818a  and  a48803a );
 a26a <=( a48788a  and  a48773a );
 a27a <=( a48758a  and  a48743a );
 a28a <=( a48728a  and  a48713a );
 a29a <=( a48698a  and  a48683a );
 a30a <=( a48668a  and  a48653a );
 a31a <=( a48638a  and  a48623a );
 a32a <=( a48608a  and  a48593a );
 a33a <=( a48578a  and  a48563a );
 a34a <=( a48548a  and  a48533a );
 a35a <=( a48518a  and  a48503a );
 a36a <=( a48488a  and  a48473a );
 a37a <=( a48458a  and  a48443a );
 a38a <=( a48428a  and  a48413a );
 a39a <=( a48398a  and  a48383a );
 a40a <=( a48368a  and  a48353a );
 a41a <=( a48338a  and  a48323a );
 a42a <=( a48308a  and  a48293a );
 a43a <=( a48278a  and  a48263a );
 a44a <=( a48248a  and  a48233a );
 a45a <=( a48218a  and  a48203a );
 a46a <=( a48188a  and  a48173a );
 a47a <=( a48158a  and  a48143a );
 a48a <=( a48128a  and  a48113a );
 a49a <=( a48098a  and  a48083a );
 a50a <=( a48068a  and  a48053a );
 a51a <=( a48038a  and  a48023a );
 a52a <=( a48008a  and  a47993a );
 a53a <=( a47978a  and  a47963a );
 a54a <=( a47948a  and  a47933a );
 a55a <=( a47918a  and  a47903a );
 a56a <=( a47888a  and  a47873a );
 a57a <=( a47858a  and  a47843a );
 a58a <=( a47828a  and  a47813a );
 a59a <=( a47798a  and  a47783a );
 a60a <=( a47768a  and  a47753a );
 a61a <=( a47738a  and  a47723a );
 a62a <=( a47708a  and  a47693a );
 a63a <=( a47678a  and  a47663a );
 a64a <=( a47648a  and  a47633a );
 a65a <=( a47618a  and  a47603a );
 a66a <=( a47588a  and  a47573a );
 a67a <=( a47558a  and  a47543a );
 a68a <=( a47528a  and  a47513a );
 a69a <=( a47498a  and  a47483a );
 a70a <=( a47468a  and  a47453a );
 a71a <=( a47438a  and  a47423a );
 a72a <=( a47408a  and  a47393a );
 a73a <=( a47378a  and  a47363a );
 a74a <=( a47348a  and  a47333a );
 a75a <=( a47318a  and  a47303a );
 a76a <=( a47288a  and  a47273a );
 a77a <=( a47258a  and  a47243a );
 a78a <=( a47228a  and  a47213a );
 a79a <=( a47198a  and  a47183a );
 a80a <=( a47168a  and  a47153a );
 a81a <=( a47138a  and  a47123a );
 a82a <=( a47108a  and  a47093a );
 a83a <=( a47078a  and  a47063a );
 a84a <=( a47048a  and  a47033a );
 a85a <=( a47018a  and  a47003a );
 a86a <=( a46988a  and  a46973a );
 a87a <=( a46958a  and  a46943a );
 a88a <=( a46928a  and  a46913a );
 a89a <=( a46898a  and  a46883a );
 a90a <=( a46868a  and  a46853a );
 a91a <=( a46838a  and  a46823a );
 a92a <=( a46808a  and  a46793a );
 a93a <=( a46778a  and  a46763a );
 a94a <=( a46748a  and  a46733a );
 a95a <=( a46718a  and  a46703a );
 a96a <=( a46688a  and  a46673a );
 a97a <=( a46658a  and  a46643a );
 a98a <=( a46628a  and  a46613a );
 a99a <=( a46598a  and  a46583a );
 a100a <=( a46568a  and  a46553a );
 a101a <=( a46538a  and  a46523a );
 a102a <=( a46508a  and  a46493a );
 a103a <=( a46478a  and  a46463a );
 a104a <=( a46448a  and  a46433a );
 a105a <=( a46418a  and  a46403a );
 a106a <=( a46388a  and  a46373a );
 a107a <=( a46358a  and  a46343a );
 a108a <=( a46328a  and  a46313a );
 a109a <=( a46298a  and  a46283a );
 a110a <=( a46268a  and  a46253a );
 a111a <=( a46238a  and  a46223a );
 a112a <=( a46208a  and  a46193a );
 a113a <=( a46178a  and  a46163a );
 a114a <=( a46148a  and  a46133a );
 a115a <=( a46118a  and  a46103a );
 a116a <=( a46088a  and  a46073a );
 a117a <=( a46058a  and  a46043a );
 a118a <=( a46028a  and  a46013a );
 a119a <=( a45998a  and  a45983a );
 a120a <=( a45968a  and  a45953a );
 a121a <=( a45938a  and  a45923a );
 a122a <=( a45908a  and  a45893a );
 a123a <=( a45878a  and  a45863a );
 a124a <=( a45848a  and  a45833a );
 a125a <=( a45818a  and  a45803a );
 a126a <=( a45788a  and  a45773a );
 a127a <=( a45758a  and  a45743a );
 a128a <=( a45728a  and  a45713a );
 a129a <=( a45698a  and  a45683a );
 a130a <=( a45668a  and  a45653a );
 a131a <=( a45638a  and  a45623a );
 a132a <=( a45608a  and  a45593a );
 a133a <=( a45578a  and  a45563a );
 a134a <=( a45548a  and  a45533a );
 a135a <=( a45518a  and  a45503a );
 a136a <=( a45488a  and  a45473a );
 a137a <=( a45458a  and  a45443a );
 a138a <=( a45428a  and  a45413a );
 a139a <=( a45398a  and  a45383a );
 a140a <=( a45368a  and  a45353a );
 a141a <=( a45338a  and  a45323a );
 a142a <=( a45308a  and  a45293a );
 a143a <=( a45278a  and  a45263a );
 a144a <=( a45248a  and  a45233a );
 a145a <=( a45218a  and  a45203a );
 a146a <=( a45188a  and  a45173a );
 a147a <=( a45158a  and  a45143a );
 a148a <=( a45128a  and  a45113a );
 a149a <=( a45098a  and  a45083a );
 a150a <=( a45068a  and  a45053a );
 a151a <=( a45038a  and  a45023a );
 a152a <=( a45008a  and  a44993a );
 a153a <=( a44978a  and  a44963a );
 a154a <=( a44948a  and  a44933a );
 a155a <=( a44918a  and  a44903a );
 a156a <=( a44888a  and  a44873a );
 a157a <=( a44858a  and  a44843a );
 a158a <=( a44828a  and  a44813a );
 a159a <=( a44798a  and  a44783a );
 a160a <=( a44768a  and  a44753a );
 a161a <=( a44738a  and  a44723a );
 a162a <=( a44708a  and  a44693a );
 a163a <=( a44678a  and  a44663a );
 a164a <=( a44648a  and  a44633a );
 a165a <=( a44618a  and  a44603a );
 a166a <=( a44588a  and  a44573a );
 a167a <=( a44558a  and  a44543a );
 a168a <=( a44528a  and  a44513a );
 a169a <=( a44498a  and  a44483a );
 a170a <=( a44468a  and  a44453a );
 a171a <=( a44438a  and  a44423a );
 a172a <=( a44408a  and  a44393a );
 a173a <=( a44378a  and  a44363a );
 a174a <=( a44348a  and  a44333a );
 a175a <=( a44318a  and  a44303a );
 a176a <=( a44288a  and  a44273a );
 a177a <=( a44258a  and  a44243a );
 a178a <=( a44228a  and  a44213a );
 a179a <=( a44198a  and  a44183a );
 a180a <=( a44168a  and  a44153a );
 a181a <=( a44138a  and  a44123a );
 a182a <=( a44108a  and  a44093a );
 a183a <=( a44078a  and  a44063a );
 a184a <=( a44048a  and  a44033a );
 a185a <=( a44018a  and  a44003a );
 a186a <=( a43988a  and  a43973a );
 a187a <=( a43958a  and  a43943a );
 a188a <=( a43928a  and  a43913a );
 a189a <=( a43898a  and  a43883a );
 a190a <=( a43868a  and  a43853a );
 a191a <=( a43838a  and  a43823a );
 a192a <=( a43808a  and  a43793a );
 a193a <=( a43778a  and  a43763a );
 a194a <=( a43748a  and  a43733a );
 a195a <=( a43718a  and  a43703a );
 a196a <=( a43688a  and  a43673a );
 a197a <=( a43658a  and  a43643a );
 a198a <=( a43628a  and  a43613a );
 a199a <=( a43598a  and  a43583a );
 a200a <=( a43568a  and  a43553a );
 a201a <=( a43538a  and  a43523a );
 a202a <=( a43508a  and  a43493a );
 a203a <=( a43478a  and  a43463a );
 a204a <=( a43448a  and  a43433a );
 a205a <=( a43418a  and  a43403a );
 a206a <=( a43388a  and  a43373a );
 a207a <=( a43358a  and  a43343a );
 a208a <=( a43328a  and  a43313a );
 a209a <=( a43298a  and  a43283a );
 a210a <=( a43268a  and  a43253a );
 a211a <=( a43238a  and  a43223a );
 a212a <=( a43208a  and  a43193a );
 a213a <=( a43178a  and  a43163a );
 a214a <=( a43148a  and  a43133a );
 a215a <=( a43118a  and  a43103a );
 a216a <=( a43088a  and  a43073a );
 a217a <=( a43058a  and  a43043a );
 a218a <=( a43028a  and  a43013a );
 a219a <=( a42998a  and  a42983a );
 a220a <=( a42968a  and  a42953a );
 a221a <=( a42938a  and  a42923a );
 a222a <=( a42908a  and  a42893a );
 a223a <=( a42878a  and  a42863a );
 a224a <=( a42848a  and  a42833a );
 a225a <=( a42818a  and  a42803a );
 a226a <=( a42788a  and  a42773a );
 a227a <=( a42758a  and  a42743a );
 a228a <=( a42728a  and  a42713a );
 a229a <=( a42698a  and  a42683a );
 a230a <=( a42668a  and  a42653a );
 a231a <=( a42638a  and  a42623a );
 a232a <=( a42608a  and  a42593a );
 a233a <=( a42578a  and  a42563a );
 a234a <=( a42548a  and  a42533a );
 a235a <=( a42518a  and  a42503a );
 a236a <=( a42488a  and  a42473a );
 a237a <=( a42458a  and  a42443a );
 a238a <=( a42428a  and  a42413a );
 a239a <=( a42398a  and  a42383a );
 a240a <=( a42368a  and  a42353a );
 a241a <=( a42338a  and  a42323a );
 a242a <=( a42308a  and  a42293a );
 a243a <=( a42278a  and  a42263a );
 a244a <=( a42248a  and  a42233a );
 a245a <=( a42218a  and  a42203a );
 a246a <=( a42188a  and  a42173a );
 a247a <=( a42158a  and  a42143a );
 a248a <=( a42128a  and  a42113a );
 a249a <=( a42098a  and  a42083a );
 a250a <=( a42068a  and  a42053a );
 a251a <=( a42038a  and  a42023a );
 a252a <=( a42008a  and  a41993a );
 a253a <=( a41978a  and  a41963a );
 a254a <=( a41948a  and  a41933a );
 a255a <=( a41918a  and  a41903a );
 a256a <=( a41888a  and  a41873a );
 a257a <=( a41858a  and  a41843a );
 a258a <=( a41828a  and  a41813a );
 a259a <=( a41798a  and  a41783a );
 a260a <=( a41768a  and  a41753a );
 a261a <=( a41738a  and  a41723a );
 a262a <=( a41708a  and  a41693a );
 a263a <=( a41678a  and  a41663a );
 a264a <=( a41648a  and  a41633a );
 a265a <=( a41618a  and  a41603a );
 a266a <=( a41588a  and  a41573a );
 a267a <=( a41558a  and  a41543a );
 a268a <=( a41528a  and  a41513a );
 a269a <=( a41498a  and  a41483a );
 a270a <=( a41468a  and  a41453a );
 a271a <=( a41438a  and  a41423a );
 a272a <=( a41408a  and  a41393a );
 a273a <=( a41378a  and  a41363a );
 a274a <=( a41348a  and  a41333a );
 a275a <=( a41318a  and  a41303a );
 a276a <=( a41288a  and  a41273a );
 a277a <=( a41258a  and  a41243a );
 a278a <=( a41228a  and  a41213a );
 a279a <=( a41198a  and  a41183a );
 a280a <=( a41168a  and  a41153a );
 a281a <=( a41138a  and  a41123a );
 a282a <=( a41108a  and  a41093a );
 a283a <=( a41078a  and  a41063a );
 a284a <=( a41048a  and  a41033a );
 a285a <=( a41018a  and  a41003a );
 a286a <=( a40988a  and  a40973a );
 a287a <=( a40958a  and  a40943a );
 a288a <=( a40928a  and  a40913a );
 a289a <=( a40898a  and  a40883a );
 a290a <=( a40868a  and  a40853a );
 a291a <=( a40838a  and  a40823a );
 a292a <=( a40808a  and  a40793a );
 a293a <=( a40778a  and  a40763a );
 a294a <=( a40748a  and  a40733a );
 a295a <=( a40718a  and  a40703a );
 a296a <=( a40688a  and  a40673a );
 a297a <=( a40658a  and  a40643a );
 a298a <=( a40628a  and  a40613a );
 a299a <=( a40598a  and  a40583a );
 a300a <=( a40568a  and  a40553a );
 a301a <=( a40538a  and  a40523a );
 a302a <=( a40508a  and  a40493a );
 a303a <=( a40478a  and  a40463a );
 a304a <=( a40448a  and  a40433a );
 a305a <=( a40418a  and  a40403a );
 a306a <=( a40388a  and  a40373a );
 a307a <=( a40358a  and  a40343a );
 a308a <=( a40328a  and  a40313a );
 a309a <=( a40298a  and  a40283a );
 a310a <=( a40268a  and  a40253a );
 a311a <=( a40238a  and  a40223a );
 a312a <=( a40208a  and  a40193a );
 a313a <=( a40178a  and  a40163a );
 a314a <=( a40148a  and  a40133a );
 a315a <=( a40118a  and  a40103a );
 a316a <=( a40088a  and  a40073a );
 a317a <=( a40058a  and  a40043a );
 a318a <=( a40028a  and  a40013a );
 a319a <=( a39998a  and  a39983a );
 a320a <=( a39968a  and  a39953a );
 a321a <=( a39938a  and  a39923a );
 a322a <=( a39908a  and  a39893a );
 a323a <=( a39878a  and  a39863a );
 a324a <=( a39848a  and  a39833a );
 a325a <=( a39818a  and  a39803a );
 a326a <=( a39788a  and  a39773a );
 a327a <=( a39758a  and  a39743a );
 a328a <=( a39728a  and  a39713a );
 a329a <=( a39698a  and  a39683a );
 a330a <=( a39668a  and  a39653a );
 a331a <=( a39638a  and  a39623a );
 a332a <=( a39608a  and  a39593a );
 a333a <=( a39578a  and  a39563a );
 a334a <=( a39548a  and  a39533a );
 a335a <=( a39518a  and  a39503a );
 a336a <=( a39488a  and  a39473a );
 a337a <=( a39458a  and  a39443a );
 a338a <=( a39428a  and  a39413a );
 a339a <=( a39398a  and  a39383a );
 a340a <=( a39368a  and  a39353a );
 a341a <=( a39338a  and  a39323a );
 a342a <=( a39308a  and  a39293a );
 a343a <=( a39278a  and  a39263a );
 a344a <=( a39248a  and  a39233a );
 a345a <=( a39218a  and  a39203a );
 a346a <=( a39188a  and  a39173a );
 a347a <=( a39158a  and  a39143a );
 a348a <=( a39128a  and  a39113a );
 a349a <=( a39098a  and  a39083a );
 a350a <=( a39068a  and  a39053a );
 a351a <=( a39038a  and  a39023a );
 a352a <=( a39008a  and  a38993a );
 a353a <=( a38978a  and  a38963a );
 a354a <=( a38948a  and  a38933a );
 a355a <=( a38918a  and  a38903a );
 a356a <=( a38888a  and  a38873a );
 a357a <=( a38858a  and  a38843a );
 a358a <=( a38828a  and  a38813a );
 a359a <=( a38798a  and  a38783a );
 a360a <=( a38768a  and  a38753a );
 a361a <=( a38738a  and  a38723a );
 a362a <=( a38708a  and  a38693a );
 a363a <=( a38678a  and  a38663a );
 a364a <=( a38648a  and  a38633a );
 a365a <=( a38618a  and  a38603a );
 a366a <=( a38588a  and  a38573a );
 a367a <=( a38558a  and  a38543a );
 a368a <=( a38528a  and  a38513a );
 a369a <=( a38498a  and  a38483a );
 a370a <=( a38468a  and  a38453a );
 a371a <=( a38438a  and  a38423a );
 a372a <=( a38408a  and  a38393a );
 a373a <=( a38378a  and  a38363a );
 a374a <=( a38348a  and  a38333a );
 a375a <=( a38318a  and  a38303a );
 a376a <=( a38288a  and  a38273a );
 a377a <=( a38258a  and  a38243a );
 a378a <=( a38228a  and  a38213a );
 a379a <=( a38198a  and  a38183a );
 a380a <=( a38168a  and  a38153a );
 a381a <=( a38138a  and  a38123a );
 a382a <=( a38108a  and  a38093a );
 a383a <=( a38078a  and  a38063a );
 a384a <=( a38048a  and  a38033a );
 a385a <=( a38018a  and  a38003a );
 a386a <=( a37990a  and  a37975a );
 a387a <=( a37962a  and  a37947a );
 a388a <=( a37934a  and  a37919a );
 a389a <=( a37906a  and  a37891a );
 a390a <=( a37878a  and  a37863a );
 a391a <=( a37850a  and  a37835a );
 a392a <=( a37822a  and  a37807a );
 a393a <=( a37794a  and  a37779a );
 a394a <=( a37766a  and  a37751a );
 a395a <=( a37738a  and  a37723a );
 a396a <=( a37710a  and  a37695a );
 a397a <=( a37682a  and  a37667a );
 a398a <=( a37654a  and  a37639a );
 a399a <=( a37626a  and  a37611a );
 a400a <=( a37598a  and  a37583a );
 a401a <=( a37570a  and  a37555a );
 a402a <=( a37542a  and  a37527a );
 a403a <=( a37514a  and  a37499a );
 a404a <=( a37486a  and  a37471a );
 a405a <=( a37458a  and  a37443a );
 a406a <=( a37430a  and  a37415a );
 a407a <=( a37402a  and  a37387a );
 a408a <=( a37374a  and  a37359a );
 a409a <=( a37346a  and  a37331a );
 a410a <=( a37318a  and  a37303a );
 a411a <=( a37290a  and  a37275a );
 a412a <=( a37262a  and  a37247a );
 a413a <=( a37234a  and  a37219a );
 a414a <=( a37206a  and  a37191a );
 a415a <=( a37178a  and  a37163a );
 a416a <=( a37150a  and  a37135a );
 a417a <=( a37122a  and  a37107a );
 a418a <=( a37094a  and  a37079a );
 a419a <=( a37066a  and  a37051a );
 a420a <=( a37038a  and  a37023a );
 a421a <=( a37010a  and  a36995a );
 a422a <=( a36982a  and  a36967a );
 a423a <=( a36954a  and  a36939a );
 a424a <=( a36926a  and  a36911a );
 a425a <=( a36898a  and  a36883a );
 a426a <=( a36870a  and  a36855a );
 a427a <=( a36842a  and  a36827a );
 a428a <=( a36814a  and  a36799a );
 a429a <=( a36786a  and  a36771a );
 a430a <=( a36758a  and  a36743a );
 a431a <=( a36730a  and  a36715a );
 a432a <=( a36702a  and  a36687a );
 a433a <=( a36674a  and  a36659a );
 a434a <=( a36646a  and  a36631a );
 a435a <=( a36618a  and  a36603a );
 a436a <=( a36590a  and  a36575a );
 a437a <=( a36562a  and  a36547a );
 a438a <=( a36534a  and  a36519a );
 a439a <=( a36506a  and  a36491a );
 a440a <=( a36478a  and  a36463a );
 a441a <=( a36450a  and  a36435a );
 a442a <=( a36422a  and  a36407a );
 a443a <=( a36394a  and  a36379a );
 a444a <=( a36366a  and  a36351a );
 a445a <=( a36338a  and  a36323a );
 a446a <=( a36310a  and  a36295a );
 a447a <=( a36282a  and  a36267a );
 a448a <=( a36254a  and  a36239a );
 a449a <=( a36226a  and  a36211a );
 a450a <=( a36198a  and  a36183a );
 a451a <=( a36170a  and  a36155a );
 a452a <=( a36142a  and  a36127a );
 a453a <=( a36114a  and  a36099a );
 a454a <=( a36086a  and  a36071a );
 a455a <=( a36058a  and  a36043a );
 a456a <=( a36030a  and  a36015a );
 a457a <=( a36002a  and  a35987a );
 a458a <=( a35974a  and  a35959a );
 a459a <=( a35946a  and  a35931a );
 a460a <=( a35918a  and  a35903a );
 a461a <=( a35890a  and  a35875a );
 a462a <=( a35862a  and  a35847a );
 a463a <=( a35834a  and  a35819a );
 a464a <=( a35806a  and  a35791a );
 a465a <=( a35778a  and  a35763a );
 a466a <=( a35750a  and  a35735a );
 a467a <=( a35722a  and  a35707a );
 a468a <=( a35694a  and  a35679a );
 a469a <=( a35666a  and  a35651a );
 a470a <=( a35638a  and  a35623a );
 a471a <=( a35610a  and  a35595a );
 a472a <=( a35582a  and  a35567a );
 a473a <=( a35554a  and  a35539a );
 a474a <=( a35526a  and  a35511a );
 a475a <=( a35498a  and  a35483a );
 a476a <=( a35470a  and  a35455a );
 a477a <=( a35442a  and  a35427a );
 a478a <=( a35414a  and  a35399a );
 a479a <=( a35386a  and  a35371a );
 a480a <=( a35358a  and  a35343a );
 a481a <=( a35330a  and  a35315a );
 a482a <=( a35302a  and  a35287a );
 a483a <=( a35274a  and  a35259a );
 a484a <=( a35246a  and  a35231a );
 a485a <=( a35218a  and  a35203a );
 a486a <=( a35190a  and  a35175a );
 a487a <=( a35162a  and  a35147a );
 a488a <=( a35134a  and  a35119a );
 a489a <=( a35106a  and  a35091a );
 a490a <=( a35078a  and  a35063a );
 a491a <=( a35050a  and  a35035a );
 a492a <=( a35022a  and  a35007a );
 a493a <=( a34994a  and  a34979a );
 a494a <=( a34966a  and  a34951a );
 a495a <=( a34938a  and  a34923a );
 a496a <=( a34910a  and  a34895a );
 a497a <=( a34882a  and  a34867a );
 a498a <=( a34854a  and  a34839a );
 a499a <=( a34826a  and  a34811a );
 a500a <=( a34798a  and  a34783a );
 a501a <=( a34770a  and  a34755a );
 a502a <=( a34742a  and  a34727a );
 a503a <=( a34714a  and  a34699a );
 a504a <=( a34686a  and  a34671a );
 a505a <=( a34658a  and  a34643a );
 a506a <=( a34630a  and  a34615a );
 a507a <=( a34602a  and  a34587a );
 a508a <=( a34574a  and  a34559a );
 a509a <=( a34546a  and  a34531a );
 a510a <=( a34518a  and  a34503a );
 a511a <=( a34490a  and  a34475a );
 a512a <=( a34462a  and  a34447a );
 a513a <=( a34434a  and  a34421a );
 a514a <=( a34408a  and  a34395a );
 a515a <=( a34382a  and  a34369a );
 a516a <=( a34356a  and  a34343a );
 a517a <=( a34330a  and  a34317a );
 a518a <=( a34304a  and  a34291a );
 a519a <=( a34278a  and  a34265a );
 a520a <=( a34252a  and  a34239a );
 a521a <=( a34226a  and  a34213a );
 a522a <=( a34200a  and  a34187a );
 a523a <=( a34174a  and  a34161a );
 a524a <=( a34148a  and  a34135a );
 a525a <=( a34122a  and  a34109a );
 a526a <=( a34096a  and  a34083a );
 a527a <=( a34070a  and  a34057a );
 a528a <=( a34044a  and  a34031a );
 a529a <=( a34018a  and  a34005a );
 a530a <=( a33992a  and  a33979a );
 a531a <=( a33966a  and  a33953a );
 a532a <=( a33940a  and  a33927a );
 a533a <=( a33914a  and  a33901a );
 a534a <=( a33888a  and  a33875a );
 a535a <=( a33862a  and  a33849a );
 a536a <=( a33836a  and  a33823a );
 a537a <=( a33810a  and  a33797a );
 a538a <=( a33784a  and  a33771a );
 a539a <=( a33758a  and  a33745a );
 a540a <=( a33732a  and  a33719a );
 a541a <=( a33706a  and  a33693a );
 a542a <=( a33680a  and  a33667a );
 a543a <=( a33654a  and  a33641a );
 a544a <=( a33628a  and  a33615a );
 a545a <=( a33602a  and  a33589a );
 a546a <=( a33576a  and  a33563a );
 a547a <=( a33550a  and  a33537a );
 a548a <=( a33524a  and  a33511a );
 a549a <=( a33498a  and  a33485a );
 a550a <=( a33472a  and  a33459a );
 a551a <=( a33446a  and  a33433a );
 a552a <=( a33420a  and  a33407a );
 a553a <=( a33394a  and  a33381a );
 a554a <=( a33368a  and  a33355a );
 a555a <=( a33342a  and  a33329a );
 a556a <=( a33316a  and  a33303a );
 a557a <=( a33290a  and  a33277a );
 a558a <=( a33264a  and  a33251a );
 a559a <=( a33238a  and  a33225a );
 a560a <=( a33212a  and  a33199a );
 a561a <=( a33186a  and  a33173a );
 a562a <=( a33160a  and  a33147a );
 a563a <=( a33134a  and  a33121a );
 a564a <=( a33108a  and  a33095a );
 a565a <=( a33082a  and  a33069a );
 a566a <=( a33056a  and  a33043a );
 a567a <=( a33030a  and  a33017a );
 a568a <=( a33004a  and  a32991a );
 a569a <=( a32978a  and  a32965a );
 a570a <=( a32952a  and  a32939a );
 a571a <=( a32926a  and  a32913a );
 a572a <=( a32900a  and  a32887a );
 a573a <=( a32874a  and  a32861a );
 a574a <=( a32848a  and  a32835a );
 a575a <=( a32822a  and  a32809a );
 a576a <=( a32796a  and  a32783a );
 a577a <=( a32770a  and  a32757a );
 a578a <=( a32744a  and  a32731a );
 a579a <=( a32718a  and  a32705a );
 a580a <=( a32692a  and  a32679a );
 a581a <=( a32666a  and  a32653a );
 a582a <=( a32640a  and  a32627a );
 a583a <=( a32614a  and  a32601a );
 a584a <=( a32588a  and  a32575a );
 a585a <=( a32562a  and  a32549a );
 a586a <=( a32536a  and  a32523a );
 a587a <=( a32510a  and  a32497a );
 a588a <=( a32484a  and  a32471a );
 a589a <=( a32458a  and  a32445a );
 a590a <=( a32432a  and  a32419a );
 a591a <=( a32406a  and  a32393a );
 a592a <=( a32380a  and  a32367a );
 a593a <=( a32354a  and  a32341a );
 a594a <=( a32328a  and  a32315a );
 a595a <=( a32302a  and  a32289a );
 a596a <=( a32276a  and  a32263a );
 a597a <=( a32250a  and  a32237a );
 a598a <=( a32224a  and  a32211a );
 a599a <=( a32198a  and  a32185a );
 a600a <=( a32172a  and  a32159a );
 a601a <=( a32146a  and  a32133a );
 a602a <=( a32120a  and  a32107a );
 a603a <=( a32094a  and  a32081a );
 a604a <=( a32068a  and  a32055a );
 a605a <=( a32042a  and  a32029a );
 a606a <=( a32016a  and  a32003a );
 a607a <=( a31990a  and  a31977a );
 a608a <=( a31964a  and  a31951a );
 a609a <=( a31938a  and  a31925a );
 a610a <=( a31912a  and  a31899a );
 a611a <=( a31886a  and  a31873a );
 a612a <=( a31860a  and  a31847a );
 a613a <=( a31834a  and  a31821a );
 a614a <=( a31808a  and  a31795a );
 a615a <=( a31782a  and  a31769a );
 a616a <=( a31756a  and  a31743a );
 a617a <=( a31730a  and  a31717a );
 a618a <=( a31704a  and  a31691a );
 a619a <=( a31678a  and  a31665a );
 a620a <=( a31652a  and  a31639a );
 a621a <=( a31626a  and  a31613a );
 a622a <=( a31600a  and  a31587a );
 a623a <=( a31574a  and  a31561a );
 a624a <=( a31548a  and  a31535a );
 a625a <=( a31522a  and  a31509a );
 a626a <=( a31496a  and  a31483a );
 a627a <=( a31470a  and  a31457a );
 a628a <=( a31444a  and  a31431a );
 a629a <=( a31418a  and  a31405a );
 a630a <=( a31392a  and  a31379a );
 a631a <=( a31366a  and  a31353a );
 a632a <=( a31340a  and  a31327a );
 a633a <=( a31314a  and  a31301a );
 a634a <=( a31288a  and  a31275a );
 a635a <=( a31262a  and  a31249a );
 a636a <=( a31236a  and  a31223a );
 a637a <=( a31210a  and  a31197a );
 a638a <=( a31184a  and  a31171a );
 a639a <=( a31158a  and  a31145a );
 a640a <=( a31132a  and  a31119a );
 a641a <=( a31106a  and  a31093a );
 a642a <=( a31080a  and  a31067a );
 a643a <=( a31054a  and  a31041a );
 a644a <=( a31028a  and  a31015a );
 a645a <=( a31002a  and  a30989a );
 a646a <=( a30976a  and  a30963a );
 a647a <=( a30950a  and  a30937a );
 a648a <=( a30924a  and  a30911a );
 a649a <=( a30898a  and  a30885a );
 a650a <=( a30872a  and  a30859a );
 a651a <=( a30846a  and  a30833a );
 a652a <=( a30820a  and  a30807a );
 a653a <=( a30794a  and  a30781a );
 a654a <=( a30768a  and  a30755a );
 a655a <=( a30742a  and  a30729a );
 a656a <=( a30716a  and  a30703a );
 a657a <=( a30690a  and  a30677a );
 a658a <=( a30664a  and  a30651a );
 a659a <=( a30638a  and  a30625a );
 a660a <=( a30612a  and  a30599a );
 a661a <=( a30586a  and  a30573a );
 a662a <=( a30560a  and  a30547a );
 a663a <=( a30534a  and  a30521a );
 a664a <=( a30508a  and  a30495a );
 a665a <=( a30482a  and  a30469a );
 a666a <=( a30456a  and  a30443a );
 a667a <=( a30430a  and  a30417a );
 a668a <=( a30404a  and  a30391a );
 a669a <=( a30378a  and  a30365a );
 a670a <=( a30352a  and  a30339a );
 a671a <=( a30326a  and  a30313a );
 a672a <=( a30300a  and  a30287a );
 a673a <=( a30274a  and  a30261a );
 a674a <=( a30248a  and  a30235a );
 a675a <=( a30222a  and  a30209a );
 a676a <=( a30196a  and  a30183a );
 a677a <=( a30170a  and  a30157a );
 a678a <=( a30144a  and  a30131a );
 a679a <=( a30118a  and  a30105a );
 a680a <=( a30092a  and  a30079a );
 a681a <=( a30066a  and  a30053a );
 a682a <=( a30040a  and  a30027a );
 a683a <=( a30014a  and  a30001a );
 a684a <=( a29988a  and  a29975a );
 a685a <=( a29962a  and  a29949a );
 a686a <=( a29936a  and  a29923a );
 a687a <=( a29910a  and  a29897a );
 a688a <=( a29884a  and  a29871a );
 a689a <=( a29858a  and  a29845a );
 a690a <=( a29832a  and  a29819a );
 a691a <=( a29806a  and  a29793a );
 a692a <=( a29780a  and  a29767a );
 a693a <=( a29754a  and  a29741a );
 a694a <=( a29728a  and  a29715a );
 a695a <=( a29702a  and  a29689a );
 a696a <=( a29676a  and  a29663a );
 a697a <=( a29650a  and  a29637a );
 a698a <=( a29624a  and  a29611a );
 a699a <=( a29598a  and  a29585a );
 a700a <=( a29572a  and  a29559a );
 a701a <=( a29546a  and  a29533a );
 a702a <=( a29520a  and  a29507a );
 a703a <=( a29494a  and  a29481a );
 a704a <=( a29468a  and  a29455a );
 a705a <=( a29442a  and  a29429a );
 a706a <=( a29416a  and  a29403a );
 a707a <=( a29390a  and  a29377a );
 a708a <=( a29364a  and  a29351a );
 a709a <=( a29338a  and  a29325a );
 a710a <=( a29312a  and  a29299a );
 a711a <=( a29286a  and  a29273a );
 a712a <=( a29260a  and  a29247a );
 a713a <=( a29234a  and  a29221a );
 a714a <=( a29208a  and  a29195a );
 a715a <=( a29182a  and  a29169a );
 a716a <=( a29156a  and  a29143a );
 a717a <=( a29130a  and  a29117a );
 a718a <=( a29104a  and  a29091a );
 a719a <=( a29078a  and  a29065a );
 a720a <=( a29052a  and  a29039a );
 a721a <=( a29026a  and  a29013a );
 a722a <=( a29000a  and  a28987a );
 a723a <=( a28974a  and  a28961a );
 a724a <=( a28948a  and  a28935a );
 a725a <=( a28922a  and  a28909a );
 a726a <=( a28896a  and  a28883a );
 a727a <=( a28870a  and  a28857a );
 a728a <=( a28844a  and  a28831a );
 a729a <=( a28818a  and  a28805a );
 a730a <=( a28792a  and  a28779a );
 a731a <=( a28766a  and  a28753a );
 a732a <=( a28740a  and  a28727a );
 a733a <=( a28714a  and  a28701a );
 a734a <=( a28688a  and  a28675a );
 a735a <=( a28662a  and  a28649a );
 a736a <=( a28636a  and  a28623a );
 a737a <=( a28610a  and  a28597a );
 a738a <=( a28584a  and  a28571a );
 a739a <=( a28558a  and  a28545a );
 a740a <=( a28532a  and  a28519a );
 a741a <=( a28506a  and  a28493a );
 a742a <=( a28480a  and  a28467a );
 a743a <=( a28454a  and  a28441a );
 a744a <=( a28428a  and  a28415a );
 a745a <=( a28402a  and  a28389a );
 a746a <=( a28376a  and  a28363a );
 a747a <=( a28350a  and  a28337a );
 a748a <=( a28324a  and  a28311a );
 a749a <=( a28298a  and  a28285a );
 a750a <=( a28272a  and  a28259a );
 a751a <=( a28246a  and  a28233a );
 a752a <=( a28220a  and  a28207a );
 a753a <=( a28194a  and  a28181a );
 a754a <=( a28168a  and  a28155a );
 a755a <=( a28142a  and  a28129a );
 a756a <=( a28116a  and  a28103a );
 a757a <=( a28090a  and  a28077a );
 a758a <=( a28064a  and  a28051a );
 a759a <=( a28038a  and  a28025a );
 a760a <=( a28012a  and  a27999a );
 a761a <=( a27986a  and  a27973a );
 a762a <=( a27960a  and  a27947a );
 a763a <=( a27934a  and  a27921a );
 a764a <=( a27908a  and  a27895a );
 a765a <=( a27882a  and  a27869a );
 a766a <=( a27856a  and  a27843a );
 a767a <=( a27830a  and  a27817a );
 a768a <=( a27804a  and  a27791a );
 a769a <=( a27778a  and  a27765a );
 a770a <=( a27752a  and  a27739a );
 a771a <=( a27726a  and  a27713a );
 a772a <=( a27700a  and  a27687a );
 a773a <=( a27674a  and  a27661a );
 a774a <=( a27648a  and  a27635a );
 a775a <=( a27622a  and  a27609a );
 a776a <=( a27596a  and  a27583a );
 a777a <=( a27570a  and  a27557a );
 a778a <=( a27544a  and  a27531a );
 a779a <=( a27518a  and  a27505a );
 a780a <=( a27492a  and  a27479a );
 a781a <=( a27466a  and  a27453a );
 a782a <=( a27440a  and  a27427a );
 a783a <=( a27414a  and  a27401a );
 a784a <=( a27388a  and  a27375a );
 a785a <=( a27362a  and  a27349a );
 a786a <=( a27336a  and  a27323a );
 a787a <=( a27310a  and  a27297a );
 a788a <=( a27284a  and  a27271a );
 a789a <=( a27258a  and  a27245a );
 a790a <=( a27232a  and  a27219a );
 a791a <=( a27206a  and  a27193a );
 a792a <=( a27180a  and  a27167a );
 a793a <=( a27154a  and  a27141a );
 a794a <=( a27128a  and  a27115a );
 a795a <=( a27102a  and  a27089a );
 a796a <=( a27076a  and  a27063a );
 a797a <=( a27050a  and  a27037a );
 a798a <=( a27024a  and  a27011a );
 a799a <=( a26998a  and  a26985a );
 a800a <=( a26972a  and  a26959a );
 a801a <=( a26946a  and  a26933a );
 a802a <=( a26920a  and  a26907a );
 a803a <=( a26894a  and  a26881a );
 a804a <=( a26868a  and  a26855a );
 a805a <=( a26842a  and  a26829a );
 a806a <=( a26816a  and  a26803a );
 a807a <=( a26790a  and  a26777a );
 a808a <=( a26764a  and  a26751a );
 a809a <=( a26738a  and  a26725a );
 a810a <=( a26712a  and  a26699a );
 a811a <=( a26686a  and  a26673a );
 a812a <=( a26660a  and  a26647a );
 a813a <=( a26634a  and  a26621a );
 a814a <=( a26608a  and  a26595a );
 a815a <=( a26582a  and  a26569a );
 a816a <=( a26556a  and  a26543a );
 a817a <=( a26530a  and  a26517a );
 a818a <=( a26504a  and  a26491a );
 a819a <=( a26478a  and  a26465a );
 a820a <=( a26452a  and  a26439a );
 a821a <=( a26426a  and  a26413a );
 a822a <=( a26400a  and  a26387a );
 a823a <=( a26374a  and  a26361a );
 a824a <=( a26348a  and  a26335a );
 a825a <=( a26322a  and  a26309a );
 a826a <=( a26296a  and  a26283a );
 a827a <=( a26270a  and  a26257a );
 a828a <=( a26244a  and  a26231a );
 a829a <=( a26218a  and  a26205a );
 a830a <=( a26192a  and  a26179a );
 a831a <=( a26166a  and  a26153a );
 a832a <=( a26140a  and  a26127a );
 a833a <=( a26114a  and  a26101a );
 a834a <=( a26088a  and  a26075a );
 a835a <=( a26062a  and  a26049a );
 a836a <=( a26036a  and  a26023a );
 a837a <=( a26010a  and  a25997a );
 a838a <=( a25984a  and  a25971a );
 a839a <=( a25958a  and  a25945a );
 a840a <=( a25932a  and  a25919a );
 a841a <=( a25906a  and  a25893a );
 a842a <=( a25880a  and  a25867a );
 a843a <=( a25854a  and  a25841a );
 a844a <=( a25828a  and  a25815a );
 a845a <=( a25802a  and  a25789a );
 a846a <=( a25776a  and  a25763a );
 a847a <=( a25750a  and  a25737a );
 a848a <=( a25724a  and  a25711a );
 a849a <=( a25698a  and  a25685a );
 a850a <=( a25672a  and  a25659a );
 a851a <=( a25646a  and  a25633a );
 a852a <=( a25620a  and  a25607a );
 a853a <=( a25594a  and  a25581a );
 a854a <=( a25568a  and  a25555a );
 a855a <=( a25542a  and  a25529a );
 a856a <=( a25516a  and  a25503a );
 a857a <=( a25490a  and  a25477a );
 a858a <=( a25464a  and  a25451a );
 a859a <=( a25438a  and  a25425a );
 a860a <=( a25412a  and  a25399a );
 a861a <=( a25386a  and  a25373a );
 a862a <=( a25360a  and  a25347a );
 a863a <=( a25334a  and  a25321a );
 a864a <=( a25308a  and  a25295a );
 a865a <=( a25282a  and  a25269a );
 a866a <=( a25256a  and  a25243a );
 a867a <=( a25230a  and  a25217a );
 a868a <=( a25204a  and  a25191a );
 a869a <=( a25178a  and  a25165a );
 a870a <=( a25152a  and  a25139a );
 a871a <=( a25126a  and  a25113a );
 a872a <=( a25100a  and  a25087a );
 a873a <=( a25074a  and  a25061a );
 a874a <=( a25048a  and  a25035a );
 a875a <=( a25022a  and  a25009a );
 a876a <=( a24996a  and  a24983a );
 a877a <=( a24970a  and  a24957a );
 a878a <=( a24944a  and  a24931a );
 a879a <=( a24918a  and  a24905a );
 a880a <=( a24892a  and  a24879a );
 a881a <=( a24866a  and  a24853a );
 a882a <=( a24840a  and  a24827a );
 a883a <=( a24814a  and  a24801a );
 a884a <=( a24788a  and  a24775a );
 a885a <=( a24762a  and  a24749a );
 a886a <=( a24736a  and  a24723a );
 a887a <=( a24710a  and  a24697a );
 a888a <=( a24684a  and  a24671a );
 a889a <=( a24658a  and  a24645a );
 a890a <=( a24632a  and  a24619a );
 a891a <=( a24606a  and  a24593a );
 a892a <=( a24580a  and  a24567a );
 a893a <=( a24554a  and  a24541a );
 a894a <=( a24528a  and  a24515a );
 a895a <=( a24502a  and  a24489a );
 a896a <=( a24476a  and  a24463a );
 a897a <=( a24450a  and  a24437a );
 a898a <=( a24424a  and  a24411a );
 a899a <=( a24398a  and  a24385a );
 a900a <=( a24372a  and  a24359a );
 a901a <=( a24346a  and  a24333a );
 a902a <=( a24320a  and  a24307a );
 a903a <=( a24294a  and  a24281a );
 a904a <=( a24268a  and  a24255a );
 a905a <=( a24242a  and  a24229a );
 a906a <=( a24216a  and  a24203a );
 a907a <=( a24190a  and  a24177a );
 a908a <=( a24164a  and  a24151a );
 a909a <=( a24138a  and  a24125a );
 a910a <=( a24112a  and  a24099a );
 a911a <=( a24086a  and  a24073a );
 a912a <=( a24060a  and  a24047a );
 a913a <=( a24034a  and  a24021a );
 a914a <=( a24008a  and  a23995a );
 a915a <=( a23982a  and  a23969a );
 a916a <=( a23956a  and  a23943a );
 a917a <=( a23930a  and  a23917a );
 a918a <=( a23904a  and  a23891a );
 a919a <=( a23878a  and  a23865a );
 a920a <=( a23852a  and  a23839a );
 a921a <=( a23826a  and  a23813a );
 a922a <=( a23800a  and  a23787a );
 a923a <=( a23774a  and  a23761a );
 a924a <=( a23748a  and  a23735a );
 a925a <=( a23722a  and  a23709a );
 a926a <=( a23696a  and  a23683a );
 a927a <=( a23670a  and  a23657a );
 a928a <=( a23644a  and  a23631a );
 a929a <=( a23618a  and  a23605a );
 a930a <=( a23592a  and  a23579a );
 a931a <=( a23566a  and  a23553a );
 a932a <=( a23540a  and  a23527a );
 a933a <=( a23514a  and  a23501a );
 a934a <=( a23488a  and  a23475a );
 a935a <=( a23462a  and  a23449a );
 a936a <=( a23436a  and  a23423a );
 a937a <=( a23410a  and  a23397a );
 a938a <=( a23384a  and  a23371a );
 a939a <=( a23358a  and  a23345a );
 a940a <=( a23332a  and  a23319a );
 a941a <=( a23306a  and  a23293a );
 a942a <=( a23280a  and  a23267a );
 a943a <=( a23254a  and  a23241a );
 a944a <=( a23228a  and  a23215a );
 a945a <=( a23202a  and  a23189a );
 a946a <=( a23176a  and  a23163a );
 a947a <=( a23150a  and  a23137a );
 a948a <=( a23124a  and  a23111a );
 a949a <=( a23098a  and  a23085a );
 a950a <=( a23072a  and  a23059a );
 a951a <=( a23046a  and  a23033a );
 a952a <=( a23020a  and  a23007a );
 a953a <=( a22994a  and  a22981a );
 a954a <=( a22968a  and  a22955a );
 a955a <=( a22942a  and  a22929a );
 a956a <=( a22916a  and  a22903a );
 a957a <=( a22890a  and  a22877a );
 a958a <=( a22864a  and  a22851a );
 a959a <=( a22838a  and  a22825a );
 a960a <=( a22812a  and  a22799a );
 a961a <=( a22786a  and  a22773a );
 a962a <=( a22760a  and  a22747a );
 a963a <=( a22734a  and  a22721a );
 a964a <=( a22708a  and  a22695a );
 a965a <=( a22682a  and  a22669a );
 a966a <=( a22656a  and  a22643a );
 a967a <=( a22630a  and  a22617a );
 a968a <=( a22604a  and  a22591a );
 a969a <=( a22578a  and  a22565a );
 a970a <=( a22552a  and  a22539a );
 a971a <=( a22526a  and  a22513a );
 a972a <=( a22500a  and  a22487a );
 a973a <=( a22474a  and  a22461a );
 a974a <=( a22448a  and  a22435a );
 a975a <=( a22422a  and  a22409a );
 a976a <=( a22396a  and  a22383a );
 a977a <=( a22370a  and  a22357a );
 a978a <=( a22344a  and  a22331a );
 a979a <=( a22318a  and  a22305a );
 a980a <=( a22292a  and  a22279a );
 a981a <=( a22266a  and  a22253a );
 a982a <=( a22240a  and  a22227a );
 a983a <=( a22214a  and  a22201a );
 a984a <=( a22188a  and  a22175a );
 a985a <=( a22162a  and  a22149a );
 a986a <=( a22136a  and  a22123a );
 a987a <=( a22110a  and  a22097a );
 a988a <=( a22084a  and  a22071a );
 a989a <=( a22058a  and  a22045a );
 a990a <=( a22032a  and  a22019a );
 a991a <=( a22006a  and  a21993a );
 a992a <=( a21980a  and  a21967a );
 a993a <=( a21954a  and  a21941a );
 a994a <=( a21928a  and  a21915a );
 a995a <=( a21902a  and  a21889a );
 a996a <=( a21876a  and  a21863a );
 a997a <=( a21850a  and  a21837a );
 a998a <=( a21824a  and  a21811a );
 a999a <=( a21798a  and  a21785a );
 a1000a <=( a21772a  and  a21759a );
 a1001a <=( a21746a  and  a21733a );
 a1002a <=( a21720a  and  a21707a );
 a1003a <=( a21694a  and  a21681a );
 a1004a <=( a21668a  and  a21655a );
 a1005a <=( a21642a  and  a21629a );
 a1006a <=( a21616a  and  a21603a );
 a1007a <=( a21590a  and  a21577a );
 a1008a <=( a21564a  and  a21551a );
 a1009a <=( a21538a  and  a21525a );
 a1010a <=( a21512a  and  a21499a );
 a1011a <=( a21486a  and  a21473a );
 a1012a <=( a21460a  and  a21447a );
 a1013a <=( a21434a  and  a21421a );
 a1014a <=( a21408a  and  a21395a );
 a1015a <=( a21382a  and  a21369a );
 a1016a <=( a21356a  and  a21343a );
 a1017a <=( a21330a  and  a21317a );
 a1018a <=( a21304a  and  a21291a );
 a1019a <=( a21278a  and  a21265a );
 a1020a <=( a21252a  and  a21239a );
 a1021a <=( a21226a  and  a21213a );
 a1022a <=( a21200a  and  a21187a );
 a1023a <=( a21174a  and  a21161a );
 a1024a <=( a21148a  and  a21135a );
 a1025a <=( a21122a  and  a21109a );
 a1026a <=( a21096a  and  a21083a );
 a1027a <=( a21070a  and  a21057a );
 a1028a <=( a21044a  and  a21031a );
 a1029a <=( a21018a  and  a21005a );
 a1030a <=( a20992a  and  a20979a );
 a1031a <=( a20966a  and  a20953a );
 a1032a <=( a20940a  and  a20927a );
 a1033a <=( a20914a  and  a20901a );
 a1034a <=( a20888a  and  a20875a );
 a1035a <=( a20862a  and  a20849a );
 a1036a <=( a20836a  and  a20823a );
 a1037a <=( a20810a  and  a20797a );
 a1038a <=( a20784a  and  a20771a );
 a1039a <=( a20758a  and  a20745a );
 a1040a <=( a20732a  and  a20719a );
 a1041a <=( a20706a  and  a20693a );
 a1042a <=( a20680a  and  a20667a );
 a1043a <=( a20654a  and  a20641a );
 a1044a <=( a20628a  and  a20615a );
 a1045a <=( a20602a  and  a20589a );
 a1046a <=( a20576a  and  a20563a );
 a1047a <=( a20550a  and  a20537a );
 a1048a <=( a20524a  and  a20511a );
 a1049a <=( a20498a  and  a20485a );
 a1050a <=( a20472a  and  a20459a );
 a1051a <=( a20446a  and  a20433a );
 a1052a <=( a20420a  and  a20407a );
 a1053a <=( a20394a  and  a20381a );
 a1054a <=( a20368a  and  a20355a );
 a1055a <=( a20342a  and  a20329a );
 a1056a <=( a20316a  and  a20303a );
 a1057a <=( a20290a  and  a20277a );
 a1058a <=( a20264a  and  a20251a );
 a1059a <=( a20238a  and  a20225a );
 a1060a <=( a20212a  and  a20199a );
 a1061a <=( a20186a  and  a20173a );
 a1062a <=( a20160a  and  a20147a );
 a1063a <=( a20134a  and  a20121a );
 a1064a <=( a20108a  and  a20095a );
 a1065a <=( a20082a  and  a20069a );
 a1066a <=( a20056a  and  a20043a );
 a1067a <=( a20030a  and  a20017a );
 a1068a <=( a20004a  and  a19991a );
 a1069a <=( a19978a  and  a19965a );
 a1070a <=( a19952a  and  a19939a );
 a1071a <=( a19926a  and  a19913a );
 a1072a <=( a19900a  and  a19887a );
 a1073a <=( a19874a  and  a19861a );
 a1074a <=( a19848a  and  a19835a );
 a1075a <=( a19822a  and  a19809a );
 a1076a <=( a19796a  and  a19783a );
 a1077a <=( a19770a  and  a19757a );
 a1078a <=( a19744a  and  a19731a );
 a1079a <=( a19718a  and  a19705a );
 a1080a <=( a19692a  and  a19679a );
 a1081a <=( a19666a  and  a19653a );
 a1082a <=( a19640a  and  a19627a );
 a1083a <=( a19614a  and  a19601a );
 a1084a <=( a19588a  and  a19575a );
 a1085a <=( a19562a  and  a19549a );
 a1086a <=( a19536a  and  a19523a );
 a1087a <=( a19510a  and  a19497a );
 a1088a <=( a19484a  and  a19471a );
 a1089a <=( a19458a  and  a19445a );
 a1090a <=( a19434a  and  a19421a );
 a1091a <=( a19410a  and  a19397a );
 a1092a <=( a19386a  and  a19373a );
 a1093a <=( a19362a  and  a19349a );
 a1094a <=( a19338a  and  a19325a );
 a1095a <=( a19314a  and  a19301a );
 a1096a <=( a19290a  and  a19277a );
 a1097a <=( a19266a  and  a19253a );
 a1098a <=( a19242a  and  a19229a );
 a1099a <=( a19218a  and  a19205a );
 a1100a <=( a19194a  and  a19181a );
 a1101a <=( a19170a  and  a19157a );
 a1102a <=( a19146a  and  a19133a );
 a1103a <=( a19122a  and  a19109a );
 a1104a <=( a19098a  and  a19085a );
 a1105a <=( a19074a  and  a19061a );
 a1106a <=( a19050a  and  a19037a );
 a1107a <=( a19026a  and  a19013a );
 a1108a <=( a19002a  and  a18989a );
 a1109a <=( a18978a  and  a18965a );
 a1110a <=( a18954a  and  a18941a );
 a1111a <=( a18930a  and  a18917a );
 a1112a <=( a18906a  and  a18893a );
 a1113a <=( a18882a  and  a18869a );
 a1114a <=( a18858a  and  a18845a );
 a1115a <=( a18834a  and  a18821a );
 a1116a <=( a18810a  and  a18797a );
 a1117a <=( a18786a  and  a18773a );
 a1118a <=( a18762a  and  a18749a );
 a1119a <=( a18738a  and  a18725a );
 a1120a <=( a18714a  and  a18701a );
 a1121a <=( a18690a  and  a18677a );
 a1122a <=( a18666a  and  a18653a );
 a1123a <=( a18642a  and  a18629a );
 a1124a <=( a18618a  and  a18605a );
 a1125a <=( a18594a  and  a18581a );
 a1126a <=( a18570a  and  a18557a );
 a1127a <=( a18546a  and  a18533a );
 a1128a <=( a18522a  and  a18509a );
 a1129a <=( a18498a  and  a18485a );
 a1130a <=( a18474a  and  a18461a );
 a1131a <=( a18450a  and  a18437a );
 a1132a <=( a18426a  and  a18413a );
 a1133a <=( a18402a  and  a18389a );
 a1134a <=( a18378a  and  a18365a );
 a1135a <=( a18354a  and  a18341a );
 a1136a <=( a18330a  and  a18317a );
 a1137a <=( a18306a  and  a18293a );
 a1138a <=( a18282a  and  a18269a );
 a1139a <=( a18258a  and  a18245a );
 a1140a <=( a18234a  and  a18221a );
 a1141a <=( a18210a  and  a18197a );
 a1142a <=( a18186a  and  a18173a );
 a1143a <=( a18162a  and  a18149a );
 a1144a <=( a18138a  and  a18125a );
 a1145a <=( a18114a  and  a18101a );
 a1146a <=( a18090a  and  a18077a );
 a1147a <=( a18066a  and  a18053a );
 a1148a <=( a18042a  and  a18029a );
 a1149a <=( a18018a  and  a18005a );
 a1150a <=( a17994a  and  a17981a );
 a1151a <=( a17970a  and  a17957a );
 a1152a <=( a17946a  and  a17933a );
 a1153a <=( a17922a  and  a17909a );
 a1154a <=( a17898a  and  a17885a );
 a1155a <=( a17874a  and  a17861a );
 a1156a <=( a17850a  and  a17837a );
 a1157a <=( a17826a  and  a17813a );
 a1158a <=( a17802a  and  a17789a );
 a1159a <=( a17778a  and  a17765a );
 a1160a <=( a17754a  and  a17741a );
 a1161a <=( a17730a  and  a17717a );
 a1162a <=( a17706a  and  a17693a );
 a1163a <=( a17682a  and  a17669a );
 a1164a <=( a17658a  and  a17645a );
 a1165a <=( a17634a  and  a17621a );
 a1166a <=( a17610a  and  a17597a );
 a1167a <=( a17586a  and  a17573a );
 a1168a <=( a17562a  and  a17549a );
 a1169a <=( a17538a  and  a17525a );
 a1170a <=( a17514a  and  a17501a );
 a1171a <=( a17490a  and  a17477a );
 a1172a <=( a17466a  and  a17453a );
 a1173a <=( a17442a  and  a17429a );
 a1174a <=( a17418a  and  a17405a );
 a1175a <=( a17394a  and  a17381a );
 a1176a <=( a17370a  and  a17357a );
 a1177a <=( a17346a  and  a17333a );
 a1178a <=( a17322a  and  a17309a );
 a1179a <=( a17298a  and  a17285a );
 a1180a <=( a17274a  and  a17261a );
 a1181a <=( a17250a  and  a17237a );
 a1182a <=( a17226a  and  a17213a );
 a1183a <=( a17202a  and  a17189a );
 a1184a <=( a17178a  and  a17165a );
 a1185a <=( a17154a  and  a17141a );
 a1186a <=( a17130a  and  a17117a );
 a1187a <=( a17106a  and  a17093a );
 a1188a <=( a17082a  and  a17069a );
 a1189a <=( a17058a  and  a17045a );
 a1190a <=( a17034a  and  a17021a );
 a1191a <=( a17010a  and  a16997a );
 a1192a <=( a16986a  and  a16973a );
 a1193a <=( a16962a  and  a16949a );
 a1194a <=( a16938a  and  a16925a );
 a1195a <=( a16914a  and  a16901a );
 a1196a <=( a16890a  and  a16877a );
 a1197a <=( a16866a  and  a16853a );
 a1198a <=( a16842a  and  a16829a );
 a1199a <=( a16818a  and  a16805a );
 a1200a <=( a16794a  and  a16781a );
 a1201a <=( a16770a  and  a16757a );
 a1202a <=( a16746a  and  a16733a );
 a1203a <=( a16722a  and  a16709a );
 a1204a <=( a16698a  and  a16685a );
 a1205a <=( a16674a  and  a16661a );
 a1206a <=( a16650a  and  a16637a );
 a1207a <=( a16626a  and  a16613a );
 a1208a <=( a16602a  and  a16589a );
 a1209a <=( a16578a  and  a16565a );
 a1210a <=( a16554a  and  a16541a );
 a1211a <=( a16530a  and  a16517a );
 a1212a <=( a16506a  and  a16493a );
 a1213a <=( a16482a  and  a16469a );
 a1214a <=( a16458a  and  a16445a );
 a1215a <=( a16434a  and  a16421a );
 a1216a <=( a16410a  and  a16397a );
 a1217a <=( a16386a  and  a16373a );
 a1218a <=( a16362a  and  a16349a );
 a1219a <=( a16338a  and  a16325a );
 a1220a <=( a16314a  and  a16301a );
 a1221a <=( a16290a  and  a16277a );
 a1222a <=( a16266a  and  a16253a );
 a1223a <=( a16242a  and  a16229a );
 a1224a <=( a16218a  and  a16205a );
 a1225a <=( a16194a  and  a16181a );
 a1226a <=( a16170a  and  a16157a );
 a1227a <=( a16146a  and  a16133a );
 a1228a <=( a16122a  and  a16109a );
 a1229a <=( a16098a  and  a16085a );
 a1230a <=( a16074a  and  a16061a );
 a1231a <=( a16050a  and  a16037a );
 a1232a <=( a16026a  and  a16013a );
 a1233a <=( a16002a  and  a15989a );
 a1234a <=( a15978a  and  a15965a );
 a1235a <=( a15954a  and  a15941a );
 a1236a <=( a15930a  and  a15917a );
 a1237a <=( a15906a  and  a15893a );
 a1238a <=( a15882a  and  a15869a );
 a1239a <=( a15858a  and  a15845a );
 a1240a <=( a15834a  and  a15821a );
 a1241a <=( a15810a  and  a15797a );
 a1242a <=( a15786a  and  a15773a );
 a1243a <=( a15762a  and  a15749a );
 a1244a <=( a15738a  and  a15725a );
 a1245a <=( a15714a  and  a15701a );
 a1246a <=( a15690a  and  a15677a );
 a1247a <=( a15666a  and  a15653a );
 a1248a <=( a15642a  and  a15629a );
 a1249a <=( a15618a  and  a15605a );
 a1250a <=( a15594a  and  a15581a );
 a1251a <=( a15570a  and  a15557a );
 a1252a <=( a15546a  and  a15533a );
 a1253a <=( a15522a  and  a15509a );
 a1254a <=( a15498a  and  a15485a );
 a1255a <=( a15474a  and  a15461a );
 a1256a <=( a15450a  and  a15437a );
 a1257a <=( a15426a  and  a15413a );
 a1258a <=( a15402a  and  a15389a );
 a1259a <=( a15378a  and  a15365a );
 a1260a <=( a15354a  and  a15341a );
 a1261a <=( a15330a  and  a15317a );
 a1262a <=( a15306a  and  a15293a );
 a1263a <=( a15282a  and  a15269a );
 a1264a <=( a15258a  and  a15245a );
 a1265a <=( a15234a  and  a15221a );
 a1266a <=( a15210a  and  a15197a );
 a1267a <=( a15186a  and  a15173a );
 a1268a <=( a15162a  and  a15149a );
 a1269a <=( a15138a  and  a15125a );
 a1270a <=( a15114a  and  a15101a );
 a1271a <=( a15090a  and  a15077a );
 a1272a <=( a15066a  and  a15053a );
 a1273a <=( a15042a  and  a15029a );
 a1274a <=( a15018a  and  a15005a );
 a1275a <=( a14994a  and  a14981a );
 a1276a <=( a14970a  and  a14957a );
 a1277a <=( a14946a  and  a14933a );
 a1278a <=( a14922a  and  a14909a );
 a1279a <=( a14898a  and  a14885a );
 a1280a <=( a14874a  and  a14861a );
 a1281a <=( a14850a  and  a14839a );
 a1282a <=( a14828a  and  a14817a );
 a1283a <=( a14806a  and  a14795a );
 a1284a <=( a14784a  and  a14773a );
 a1285a <=( a14762a  and  a14751a );
 a1286a <=( a14740a  and  a14729a );
 a1287a <=( a14718a  and  a14707a );
 a1288a <=( a14696a  and  a14685a );
 a1289a <=( a14674a  and  a14663a );
 a1290a <=( a14652a  and  a14641a );
 a1291a <=( a14630a  and  a14619a );
 a1292a <=( a14608a  and  a14597a );
 a1293a <=( a14586a  and  a14575a );
 a1294a <=( a14564a  and  a14553a );
 a1295a <=( a14542a  and  a14531a );
 a1296a <=( a14520a  and  a14509a );
 a1297a <=( a14498a  and  a14487a );
 a1298a <=( a14476a  and  a14465a );
 a1299a <=( a14454a  and  a14443a );
 a1300a <=( a14432a  and  a14421a );
 a1301a <=( a14410a  and  a14399a );
 a1302a <=( a14388a  and  a14377a );
 a1303a <=( a14366a  and  a14355a );
 a1304a <=( a14344a  and  a14333a );
 a1305a <=( a14322a  and  a14311a );
 a1306a <=( a14300a  and  a14289a );
 a1307a <=( a14278a  and  a14267a );
 a1308a <=( a14256a  and  a14245a );
 a1309a <=( a14234a  and  a14223a );
 a1310a <=( a14212a  and  a14201a );
 a1311a <=( a14190a  and  a14179a );
 a1312a <=( a14168a  and  a14157a );
 a1313a <=( a14146a  and  a14135a );
 a1314a <=( a14124a  and  a14113a );
 a1315a <=( a14102a  and  a14091a );
 a1316a <=( a14080a  and  a14069a );
 a1317a <=( a14058a  and  a14047a );
 a1318a <=( a14036a  and  a14025a );
 a1319a <=( a14014a  and  a14003a );
 a1320a <=( a13992a  and  a13981a );
 a1321a <=( a13970a  and  a13959a );
 a1322a <=( a13948a  and  a13937a );
 a1323a <=( a13926a  and  a13915a );
 a1324a <=( a13904a  and  a13893a );
 a1325a <=( a13882a  and  a13871a );
 a1326a <=( a13860a  and  a13849a );
 a1327a <=( a13838a  and  a13827a );
 a1328a <=( a13816a  and  a13805a );
 a1329a <=( a13794a  and  a13783a );
 a1330a <=( a13772a  and  a13761a );
 a1331a <=( a13750a  and  a13739a );
 a1332a <=( a13728a  and  a13717a );
 a1333a <=( a13706a  and  a13695a );
 a1334a <=( a13684a  and  a13673a );
 a1335a <=( a13662a  and  a13651a );
 a1336a <=( a13640a  and  a13629a );
 a1337a <=( a13618a  and  a13607a );
 a1338a <=( a13596a  and  a13585a );
 a1339a <=( a13574a  and  a13563a );
 a1340a <=( a13552a  and  a13541a );
 a1341a <=( a13530a  and  a13519a );
 a1342a <=( a13508a  and  a13497a );
 a1343a <=( a13486a  and  a13475a );
 a1344a <=( a13464a  and  a13453a );
 a1345a <=( a13442a  and  a13431a );
 a1346a <=( a13420a  and  a13409a );
 a1347a <=( a13398a  and  a13387a );
 a1348a <=( a13376a  and  a13365a );
 a1349a <=( a13354a  and  a13343a );
 a1350a <=( a13332a  and  a13321a );
 a1351a <=( a13310a  and  a13299a );
 a1352a <=( a13288a  and  a13277a );
 a1353a <=( a13266a  and  a13255a );
 a1354a <=( a13244a  and  a13233a );
 a1355a <=( a13222a  and  a13211a );
 a1356a <=( a13200a  and  a13189a );
 a1357a <=( a13178a  and  a13167a );
 a1358a <=( a13156a  and  a13145a );
 a1359a <=( a13134a  and  a13123a );
 a1360a <=( a13112a  and  a13101a );
 a1361a <=( a13090a  and  a13079a );
 a1362a <=( a13068a  and  a13057a );
 a1363a <=( a13046a  and  a13035a );
 a1364a <=( a13024a  and  a13013a );
 a1365a <=( a13002a  and  a12991a );
 a1366a <=( a12980a  and  a12969a );
 a1367a <=( a12958a  and  a12947a );
 a1368a <=( a12936a  and  a12925a );
 a1369a <=( a12914a  and  a12903a );
 a1370a <=( a12892a  and  a12881a );
 a1371a <=( a12870a  and  a12859a );
 a1372a <=( a12848a  and  a12837a );
 a1373a <=( a12826a  and  a12815a );
 a1374a <=( a12804a  and  a12793a );
 a1375a <=( a12782a  and  a12771a );
 a1376a <=( a12760a  and  a12749a );
 a1377a <=( a12738a  and  a12727a );
 a1378a <=( a12716a  and  a12705a );
 a1379a <=( a12694a  and  a12683a );
 a1380a <=( a12672a  and  a12661a );
 a1381a <=( a12650a  and  a12639a );
 a1382a <=( a12628a  and  a12617a );
 a1383a <=( a12606a  and  a12595a );
 a1384a <=( a12584a  and  a12573a );
 a1385a <=( a12562a  and  a12551a );
 a1386a <=( a12540a  and  a12529a );
 a1387a <=( a12518a  and  a12507a );
 a1388a <=( a12496a  and  a12485a );
 a1389a <=( a12474a  and  a12463a );
 a1390a <=( a12452a  and  a12441a );
 a1391a <=( a12430a  and  a12419a );
 a1392a <=( a12408a  and  a12397a );
 a1393a <=( a12386a  and  a12375a );
 a1394a <=( a12364a  and  a12353a );
 a1395a <=( a12342a  and  a12331a );
 a1396a <=( a12320a  and  a12309a );
 a1397a <=( a12298a  and  a12287a );
 a1398a <=( a12276a  and  a12265a );
 a1399a <=( a12254a  and  a12243a );
 a1400a <=( a12232a  and  a12221a );
 a1401a <=( a12210a  and  a12199a );
 a1402a <=( a12188a  and  a12177a );
 a1403a <=( a12166a  and  a12155a );
 a1404a <=( a12144a  and  a12133a );
 a1405a <=( a12122a  and  a12111a );
 a1406a <=( a12100a  and  a12089a );
 a1407a <=( a12078a  and  a12067a );
 a1408a <=( a12056a  and  a12045a );
 a1409a <=( a12034a  and  a12023a );
 a1410a <=( a12012a  and  a12001a );
 a1411a <=( a11990a  and  a11979a );
 a1412a <=( a11968a  and  a11957a );
 a1413a <=( a11946a  and  a11935a );
 a1414a <=( a11924a  and  a11913a );
 a1415a <=( a11902a  and  a11891a );
 a1416a <=( a11880a  and  a11869a );
 a1417a <=( a11858a  and  a11847a );
 a1418a <=( a11836a  and  a11825a );
 a1419a <=( a11814a  and  a11803a );
 a1420a <=( a11792a  and  a11781a );
 a1421a <=( a11770a  and  a11759a );
 a1422a <=( a11748a  and  a11737a );
 a1423a <=( a11726a  and  a11715a );
 a1424a <=( a11704a  and  a11693a );
 a1425a <=( a11682a  and  a11671a );
 a1426a <=( a11660a  and  a11649a );
 a1427a <=( a11638a  and  a11627a );
 a1428a <=( a11616a  and  a11605a );
 a1429a <=( a11594a  and  a11583a );
 a1430a <=( a11572a  and  a11561a );
 a1431a <=( a11550a  and  a11539a );
 a1432a <=( a11528a  and  a11517a );
 a1433a <=( a11506a  and  a11495a );
 a1434a <=( a11484a  and  a11473a );
 a1435a <=( a11462a  and  a11451a );
 a1436a <=( a11440a  and  a11429a );
 a1437a <=( a11418a  and  a11407a );
 a1438a <=( a11396a  and  a11385a );
 a1439a <=( a11374a  and  a11363a );
 a1440a <=( a11352a  and  a11341a );
 a1441a <=( a11330a  and  a11319a );
 a1442a <=( a11308a  and  a11297a );
 a1443a <=( a11286a  and  a11275a );
 a1444a <=( a11264a  and  a11253a );
 a1445a <=( a11242a  and  a11231a );
 a1446a <=( a11220a  and  a11209a );
 a1447a <=( a11198a  and  a11187a );
 a1448a <=( a11176a  and  a11165a );
 a1449a <=( a11154a  and  a11143a );
 a1450a <=( a11132a  and  a11121a );
 a1451a <=( a11110a  and  a11099a );
 a1452a <=( a11088a  and  a11077a );
 a1453a <=( a11066a  and  a11055a );
 a1454a <=( a11044a  and  a11033a );
 a1455a <=( a11022a  and  a11011a );
 a1456a <=( a11000a  and  a10989a );
 a1457a <=( a10978a  and  a10967a );
 a1458a <=( a10956a  and  a10945a );
 a1459a <=( a10934a  and  a10923a );
 a1460a <=( a10912a  and  a10901a );
 a1461a <=( a10890a  and  a10879a );
 a1462a <=( a10868a  and  a10857a );
 a1463a <=( a10846a  and  a10835a );
 a1464a <=( a10824a  and  a10813a );
 a1465a <=( a10802a  and  a10791a );
 a1466a <=( a10780a  and  a10769a );
 a1467a <=( a10758a  and  a10747a );
 a1468a <=( a10736a  and  a10725a );
 a1469a <=( a10714a  and  a10703a );
 a1470a <=( a10692a  and  a10681a );
 a1471a <=( a10670a  and  a10659a );
 a1472a <=( a10648a  and  a10637a );
 a1473a <=( a10626a  and  a10615a );
 a1474a <=( a10604a  and  a10593a );
 a1475a <=( a10582a  and  a10571a );
 a1476a <=( a10560a  and  a10549a );
 a1477a <=( a10538a  and  a10527a );
 a1478a <=( a10516a  and  a10505a );
 a1479a <=( a10494a  and  a10483a );
 a1480a <=( a10472a  and  a10461a );
 a1481a <=( a10450a  and  a10439a );
 a1482a <=( a10428a  and  a10417a );
 a1483a <=( a10406a  and  a10395a );
 a1484a <=( a10384a  and  a10373a );
 a1485a <=( a10362a  and  a10351a );
 a1486a <=( a10340a  and  a10329a );
 a1487a <=( a10318a  and  a10307a );
 a1488a <=( a10296a  and  a10285a );
 a1489a <=( a10274a  and  a10263a );
 a1490a <=( a10252a  and  a10241a );
 a1491a <=( a10230a  and  a10219a );
 a1492a <=( a10208a  and  a10197a );
 a1493a <=( a10186a  and  a10175a );
 a1494a <=( a10164a  and  a10153a );
 a1495a <=( a10142a  and  a10131a );
 a1496a <=( a10120a  and  a10109a );
 a1497a <=( a10098a  and  a10087a );
 a1498a <=( a10076a  and  a10065a );
 a1499a <=( a10054a  and  a10043a );
 a1500a <=( a10032a  and  a10021a );
 a1501a <=( a10010a  and  a9999a );
 a1502a <=( a9988a  and  a9977a );
 a1503a <=( a9966a  and  a9955a );
 a1504a <=( a9944a  and  a9933a );
 a1505a <=( a9922a  and  a9911a );
 a1506a <=( a9900a  and  a9889a );
 a1507a <=( a9878a  and  a9867a );
 a1508a <=( a9856a  and  a9845a );
 a1509a <=( a9834a  and  a9823a );
 a1510a <=( a9812a  and  a9801a );
 a1511a <=( a9790a  and  a9779a );
 a1512a <=( a9768a  and  a9757a );
 a1513a <=( a9746a  and  a9735a );
 a1514a <=( a9724a  and  a9713a );
 a1515a <=( a9702a  and  a9691a );
 a1516a <=( a9680a  and  a9669a );
 a1517a <=( a9658a  and  a9647a );
 a1518a <=( a9636a  and  a9625a );
 a1519a <=( a9614a  and  a9603a );
 a1520a <=( a9592a  and  a9581a );
 a1521a <=( a9570a  and  a9559a );
 a1522a <=( a9548a  and  a9537a );
 a1523a <=( a9526a  and  a9515a );
 a1524a <=( a9504a  and  a9493a );
 a1525a <=( a9482a  and  a9471a );
 a1526a <=( a9460a  and  a9449a );
 a1527a <=( a9438a  and  a9427a );
 a1528a <=( a9416a  and  a9405a );
 a1529a <=( a9394a  and  a9383a );
 a1530a <=( a9372a  and  a9361a );
 a1531a <=( a9350a  and  a9339a );
 a1532a <=( a9328a  and  a9317a );
 a1533a <=( a9306a  and  a9295a );
 a1534a <=( a9284a  and  a9273a );
 a1535a <=( a9262a  and  a9251a );
 a1536a <=( a9240a  and  a9229a );
 a1537a <=( a9218a  and  a9207a );
 a1538a <=( a9196a  and  a9185a );
 a1539a <=( a9174a  and  a9163a );
 a1540a <=( a9152a  and  a9141a );
 a1541a <=( a9130a  and  a9119a );
 a1542a <=( a9108a  and  a9097a );
 a1543a <=( a9086a  and  a9075a );
 a1544a <=( a9064a  and  a9053a );
 a1545a <=( a9042a  and  a9031a );
 a1546a <=( a9020a  and  a9009a );
 a1547a <=( a8998a  and  a8987a );
 a1548a <=( a8976a  and  a8965a );
 a1549a <=( a8954a  and  a8943a );
 a1550a <=( a8932a  and  a8921a );
 a1551a <=( a8910a  and  a8899a );
 a1552a <=( a8888a  and  a8877a );
 a1553a <=( a8866a  and  a8855a );
 a1554a <=( a8844a  and  a8833a );
 a1555a <=( a8822a  and  a8811a );
 a1556a <=( a8800a  and  a8789a );
 a1557a <=( a8778a  and  a8767a );
 a1558a <=( a8756a  and  a8745a );
 a1559a <=( a8734a  and  a8723a );
 a1560a <=( a8712a  and  a8701a );
 a1561a <=( a8690a  and  a8679a );
 a1562a <=( a8668a  and  a8657a );
 a1563a <=( a8646a  and  a8635a );
 a1564a <=( a8624a  and  a8613a );
 a1565a <=( a8602a  and  a8591a );
 a1566a <=( a8580a  and  a8569a );
 a1567a <=( a8558a  and  a8547a );
 a1568a <=( a8536a  and  a8525a );
 a1569a <=( a8514a  and  a8503a );
 a1570a <=( a8494a  and  a8483a );
 a1571a <=( a8474a  and  a8463a );
 a1572a <=( a8454a  and  a8443a );
 a1573a <=( a8434a  and  a8423a );
 a1574a <=( a8414a  and  a8403a );
 a1575a <=( a8394a  and  a8383a );
 a1576a <=( a8374a  and  a8363a );
 a1577a <=( a8354a  and  a8343a );
 a1578a <=( a8334a  and  a8323a );
 a1579a <=( a8314a  and  a8303a );
 a1580a <=( a8294a  and  a8283a );
 a1581a <=( a8274a  and  a8263a );
 a1582a <=( a8254a  and  a8243a );
 a1583a <=( a8234a  and  a8223a );
 a1584a <=( a8214a  and  a8203a );
 a1585a <=( a8194a  and  a8183a );
 a1586a <=( a8174a  and  a8163a );
 a1587a <=( a8154a  and  a8143a );
 a1588a <=( a8134a  and  a8123a );
 a1589a <=( a8114a  and  a8103a );
 a1590a <=( a8094a  and  a8083a );
 a1591a <=( a8074a  and  a8063a );
 a1592a <=( a8054a  and  a8043a );
 a1593a <=( a8034a  and  a8023a );
 a1594a <=( a8014a  and  a8003a );
 a1595a <=( a7994a  and  a7983a );
 a1596a <=( a7974a  and  a7963a );
 a1597a <=( a7954a  and  a7943a );
 a1598a <=( a7934a  and  a7923a );
 a1599a <=( a7914a  and  a7903a );
 a1600a <=( a7894a  and  a7883a );
 a1601a <=( a7874a  and  a7863a );
 a1602a <=( a7854a  and  a7843a );
 a1603a <=( a7834a  and  a7823a );
 a1604a <=( a7814a  and  a7803a );
 a1605a <=( a7794a  and  a7783a );
 a1606a <=( a7774a  and  a7763a );
 a1607a <=( a7754a  and  a7743a );
 a1608a <=( a7734a  and  a7723a );
 a1609a <=( a7714a  and  a7703a );
 a1610a <=( a7694a  and  a7683a );
 a1611a <=( a7674a  and  a7663a );
 a1612a <=( a7654a  and  a7643a );
 a1613a <=( a7634a  and  a7623a );
 a1614a <=( a7614a  and  a7603a );
 a1615a <=( a7594a  and  a7583a );
 a1616a <=( a7574a  and  a7563a );
 a1617a <=( a7554a  and  a7543a );
 a1618a <=( a7534a  and  a7523a );
 a1619a <=( a7514a  and  a7503a );
 a1620a <=( a7494a  and  a7483a );
 a1621a <=( a7474a  and  a7463a );
 a1622a <=( a7454a  and  a7443a );
 a1623a <=( a7434a  and  a7423a );
 a1624a <=( a7414a  and  a7403a );
 a1625a <=( a7394a  and  a7383a );
 a1626a <=( a7374a  and  a7363a );
 a1627a <=( a7354a  and  a7343a );
 a1628a <=( a7334a  and  a7323a );
 a1629a <=( a7314a  and  a7303a );
 a1630a <=( a7294a  and  a7283a );
 a1631a <=( a7274a  and  a7263a );
 a1632a <=( a7254a  and  a7243a );
 a1633a <=( a7234a  and  a7223a );
 a1634a <=( a7214a  and  a7203a );
 a1635a <=( a7194a  and  a7183a );
 a1636a <=( a7174a  and  a7163a );
 a1637a <=( a7154a  and  a7143a );
 a1638a <=( a7134a  and  a7123a );
 a1639a <=( a7114a  and  a7103a );
 a1640a <=( a7094a  and  a7083a );
 a1641a <=( a7074a  and  a7063a );
 a1642a <=( a7054a  and  a7043a );
 a1643a <=( a7034a  and  a7023a );
 a1644a <=( a7014a  and  a7003a );
 a1645a <=( a6994a  and  a6983a );
 a1646a <=( a6974a  and  a6963a );
 a1647a <=( a6954a  and  a6943a );
 a1648a <=( a6934a  and  a6923a );
 a1649a <=( a6914a  and  a6903a );
 a1650a <=( a6894a  and  a6883a );
 a1651a <=( a6874a  and  a6863a );
 a1652a <=( a6854a  and  a6843a );
 a1653a <=( a6834a  and  a6823a );
 a1654a <=( a6814a  and  a6803a );
 a1655a <=( a6794a  and  a6783a );
 a1656a <=( a6774a  and  a6763a );
 a1657a <=( a6754a  and  a6743a );
 a1658a <=( a6734a  and  a6723a );
 a1659a <=( a6714a  and  a6703a );
 a1660a <=( a6694a  and  a6683a );
 a1661a <=( a6674a  and  a6663a );
 a1662a <=( a6654a  and  a6643a );
 a1663a <=( a6634a  and  a6623a );
 a1664a <=( a6614a  and  a6603a );
 a1665a <=( a6594a  and  a6585a );
 a1666a <=( a6576a  and  a6567a );
 a1667a <=( a6558a  and  a6549a );
 a1668a <=( a6540a  and  a6531a );
 a1669a <=( a6522a  and  a6513a );
 a1670a <=( a6504a  and  a6495a );
 a1671a <=( a6486a  and  a6477a );
 a1672a <=( a6468a  and  a6459a );
 a1673a <=( a6450a  and  a6441a );
 a1674a <=( a6432a  and  a6423a );
 a1675a <=( a6414a  and  a6405a );
 a1676a <=( a6396a  and  a6387a );
 a1677a <=( a6378a  and  a6369a );
 a1678a <=( a6360a  and  a6351a );
 a1679a <=( a6342a  and  a6333a );
 a1680a <=( a6324a  and  a6315a );
 a1681a <=( a6306a  and  a6297a );
 a1682a <=( a6288a  and  a6279a );
 a1683a <=( a6270a  and  a6261a );
 a1684a <=( a6252a  and  a6243a );
 a1685a <=( a6234a  and  a6225a );
 a1686a <=( a6216a  and  a6207a );
 a1687a <=( a6198a  and  a6189a );
 a1688a <=( a6180a  and  a6171a );
 a1689a <=( a6162a  and  a6153a );
 a1690a <=( a6144a  and  a6135a );
 a1691a <=( a6126a  and  a6117a );
 a1692a <=( a6108a  and  a6099a );
 a1693a <=( a6090a  and  a6081a );
 a1694a <=( a6072a  and  a6063a );
 a1695a <=( a6054a  and  a6045a );
 a1696a <=( a6036a  and  a6027a );
 a1697a <=( a6018a  and  a6009a );
 a1698a <=( a6000a  and  a5991a );
 a1699a <=( a5982a  and  a5973a );
 a1700a <=( a5964a  and  a5955a );
 a1701a <=( a5946a  and  a5937a );
 a1702a <=( a5928a  and  a5919a );
 a1703a <=( a5910a  and  a5901a );
 a1704a <=( a5892a  and  a5883a );
 a1705a <=( a5874a  and  a5865a );
 a1706a <=( a5856a  and  a5847a );
 a1707a <=( a5838a  and  a5829a );
 a1708a <=( a5820a  and  a5811a );
 a1709a <=( a5802a  and  a5793a );
 a1710a <=( a5784a  and  a5775a );
 a1711a <=( a5766a  and  a5757a );
 a1712a <=( a5748a  and  a5739a );
 a1713a <=( a5730a  and  a5721a );
 a1714a <=( a5714a  and  a5705a );
 a1715a <=( a5698a  and  a5689a );
 a1716a <=( a5682a  and  a5673a );
 a1717a <=( a5666a  and  a5657a );
 a1718a <=( a5650a  and  a5641a );
 a1719a <=( a5634a  and  a5625a );
 a1720a <=( a5618a  and  a5609a );
 a1721a <=( a5602a  and  a5593a );
 a1722a <=( a5586a  and  a5577a );
 a1723a <=( a5570a  and  a5561a );
 a1724a <=( a5554a  and  a5545a );
 a1725a <=( a5538a  and  a5529a );
 a1726a <=( a5522a  and  a5513a );
 a1727a <=( a5506a  and  a5497a );
 a1728a <=( a5490a  and  a5481a );
 a1729a <=( a5474a  and  a5467a );
 a1730a <=( a5462a  and  a5455a );
 a1731a <=( a5450a  and  a5443a );
 a1732a <=( a5438a  and  a5431a );
 a1733a <=( a5426a  and  a5421a );
 a1734a <=( a5416a  and  a5411a );
 a1735a <=( a5406a  and  a5401a );
 a1736a <=( a5396a  and  a5391a );
 a1737a <=( a5386a  and  a5381a );
 a1738a <=( a5376a  and  a5371a );
 a1739a <=( a5366a  and  a5361a );
 a1740a <=( a5356a  and  a5351a );
 a1741a <=( a5346a  and  a5341a );
 a1742a <=( a5336a  and  a5331a );
 a1743a <=( a5326a  and  a5321a );
 a1744a <=( a5316a  and  a5311a );
 a1745a <=( a5306a  and  a5301a );
 a1746a <=( a5298a  and  a5293a );
 a1747a <=( a5290a  and  a5287a );
 a1748a <=( a5284a  and  a5281a );
 a1749a <=( a5278a  and  a5275a );
 a1750a <=( a5272a  and  a5269a );
 a1751a <=( a5266a  and  a5263a );
 a1752a <=( a5260a  and  a5257a );
 a1756a <=( a1750a ) or ( a1751a );
 a1757a <=( a1752a ) or ( a1756a );
 a1761a <=( a1747a ) or ( a1748a );
 a1762a <=( a1749a ) or ( a1761a );
 a1763a <=( a1762a ) or ( a1757a );
 a1767a <=( a1744a ) or ( a1745a );
 a1768a <=( a1746a ) or ( a1767a );
 a1771a <=( a1742a ) or ( a1743a );
 a1774a <=( a1740a ) or ( a1741a );
 a1775a <=( a1774a ) or ( a1771a );
 a1776a <=( a1775a ) or ( a1768a );
 a1777a <=( a1776a ) or ( a1763a );
 a1781a <=( a1737a ) or ( a1738a );
 a1782a <=( a1739a ) or ( a1781a );
 a1785a <=( a1735a ) or ( a1736a );
 a1788a <=( a1733a ) or ( a1734a );
 a1789a <=( a1788a ) or ( a1785a );
 a1790a <=( a1789a ) or ( a1782a );
 a1794a <=( a1730a ) or ( a1731a );
 a1795a <=( a1732a ) or ( a1794a );
 a1798a <=( a1728a ) or ( a1729a );
 a1801a <=( a1726a ) or ( a1727a );
 a1802a <=( a1801a ) or ( a1798a );
 a1803a <=( a1802a ) or ( a1795a );
 a1804a <=( a1803a ) or ( a1790a );
 a1805a <=( a1804a ) or ( a1777a );
 a1809a <=( a1723a ) or ( a1724a );
 a1810a <=( a1725a ) or ( a1809a );
 a1814a <=( a1720a ) or ( a1721a );
 a1815a <=( a1722a ) or ( a1814a );
 a1816a <=( a1815a ) or ( a1810a );
 a1820a <=( a1717a ) or ( a1718a );
 a1821a <=( a1719a ) or ( a1820a );
 a1824a <=( a1715a ) or ( a1716a );
 a1827a <=( a1713a ) or ( a1714a );
 a1828a <=( a1827a ) or ( a1824a );
 a1829a <=( a1828a ) or ( a1821a );
 a1830a <=( a1829a ) or ( a1816a );
 a1834a <=( a1710a ) or ( a1711a );
 a1835a <=( a1712a ) or ( a1834a );
 a1838a <=( a1708a ) or ( a1709a );
 a1841a <=( a1706a ) or ( a1707a );
 a1842a <=( a1841a ) or ( a1838a );
 a1843a <=( a1842a ) or ( a1835a );
 a1847a <=( a1703a ) or ( a1704a );
 a1848a <=( a1705a ) or ( a1847a );
 a1851a <=( a1701a ) or ( a1702a );
 a1854a <=( a1699a ) or ( a1700a );
 a1855a <=( a1854a ) or ( a1851a );
 a1856a <=( a1855a ) or ( a1848a );
 a1857a <=( a1856a ) or ( a1843a );
 a1858a <=( a1857a ) or ( a1830a );
 a1859a <=( a1858a ) or ( a1805a );
 a1863a <=( a1696a ) or ( a1697a );
 a1864a <=( a1698a ) or ( a1863a );
 a1868a <=( a1693a ) or ( a1694a );
 a1869a <=( a1695a ) or ( a1868a );
 a1870a <=( a1869a ) or ( a1864a );
 a1874a <=( a1690a ) or ( a1691a );
 a1875a <=( a1692a ) or ( a1874a );
 a1878a <=( a1688a ) or ( a1689a );
 a1881a <=( a1686a ) or ( a1687a );
 a1882a <=( a1881a ) or ( a1878a );
 a1883a <=( a1882a ) or ( a1875a );
 a1884a <=( a1883a ) or ( a1870a );
 a1888a <=( a1683a ) or ( a1684a );
 a1889a <=( a1685a ) or ( a1888a );
 a1892a <=( a1681a ) or ( a1682a );
 a1895a <=( a1679a ) or ( a1680a );
 a1896a <=( a1895a ) or ( a1892a );
 a1897a <=( a1896a ) or ( a1889a );
 a1901a <=( a1676a ) or ( a1677a );
 a1902a <=( a1678a ) or ( a1901a );
 a1905a <=( a1674a ) or ( a1675a );
 a1908a <=( a1672a ) or ( a1673a );
 a1909a <=( a1908a ) or ( a1905a );
 a1910a <=( a1909a ) or ( a1902a );
 a1911a <=( a1910a ) or ( a1897a );
 a1912a <=( a1911a ) or ( a1884a );
 a1916a <=( a1669a ) or ( a1670a );
 a1917a <=( a1671a ) or ( a1916a );
 a1920a <=( a1667a ) or ( a1668a );
 a1923a <=( a1665a ) or ( a1666a );
 a1924a <=( a1923a ) or ( a1920a );
 a1925a <=( a1924a ) or ( a1917a );
 a1929a <=( a1662a ) or ( a1663a );
 a1930a <=( a1664a ) or ( a1929a );
 a1933a <=( a1660a ) or ( a1661a );
 a1936a <=( a1658a ) or ( a1659a );
 a1937a <=( a1936a ) or ( a1933a );
 a1938a <=( a1937a ) or ( a1930a );
 a1939a <=( a1938a ) or ( a1925a );
 a1943a <=( a1655a ) or ( a1656a );
 a1944a <=( a1657a ) or ( a1943a );
 a1947a <=( a1653a ) or ( a1654a );
 a1950a <=( a1651a ) or ( a1652a );
 a1951a <=( a1950a ) or ( a1947a );
 a1952a <=( a1951a ) or ( a1944a );
 a1956a <=( a1648a ) or ( a1649a );
 a1957a <=( a1650a ) or ( a1956a );
 a1960a <=( a1646a ) or ( a1647a );
 a1963a <=( a1644a ) or ( a1645a );
 a1964a <=( a1963a ) or ( a1960a );
 a1965a <=( a1964a ) or ( a1957a );
 a1966a <=( a1965a ) or ( a1952a );
 a1967a <=( a1966a ) or ( a1939a );
 a1968a <=( a1967a ) or ( a1912a );
 a1969a <=( a1968a ) or ( a1859a );
 a1973a <=( a1641a ) or ( a1642a );
 a1974a <=( a1643a ) or ( a1973a );
 a1978a <=( a1638a ) or ( a1639a );
 a1979a <=( a1640a ) or ( a1978a );
 a1980a <=( a1979a ) or ( a1974a );
 a1984a <=( a1635a ) or ( a1636a );
 a1985a <=( a1637a ) or ( a1984a );
 a1988a <=( a1633a ) or ( a1634a );
 a1991a <=( a1631a ) or ( a1632a );
 a1992a <=( a1991a ) or ( a1988a );
 a1993a <=( a1992a ) or ( a1985a );
 a1994a <=( a1993a ) or ( a1980a );
 a1998a <=( a1628a ) or ( a1629a );
 a1999a <=( a1630a ) or ( a1998a );
 a2002a <=( a1626a ) or ( a1627a );
 a2005a <=( a1624a ) or ( a1625a );
 a2006a <=( a2005a ) or ( a2002a );
 a2007a <=( a2006a ) or ( a1999a );
 a2011a <=( a1621a ) or ( a1622a );
 a2012a <=( a1623a ) or ( a2011a );
 a2015a <=( a1619a ) or ( a1620a );
 a2018a <=( a1617a ) or ( a1618a );
 a2019a <=( a2018a ) or ( a2015a );
 a2020a <=( a2019a ) or ( a2012a );
 a2021a <=( a2020a ) or ( a2007a );
 a2022a <=( a2021a ) or ( a1994a );
 a2026a <=( a1614a ) or ( a1615a );
 a2027a <=( a1616a ) or ( a2026a );
 a2030a <=( a1612a ) or ( a1613a );
 a2033a <=( a1610a ) or ( a1611a );
 a2034a <=( a2033a ) or ( a2030a );
 a2035a <=( a2034a ) or ( a2027a );
 a2039a <=( a1607a ) or ( a1608a );
 a2040a <=( a1609a ) or ( a2039a );
 a2043a <=( a1605a ) or ( a1606a );
 a2046a <=( a1603a ) or ( a1604a );
 a2047a <=( a2046a ) or ( a2043a );
 a2048a <=( a2047a ) or ( a2040a );
 a2049a <=( a2048a ) or ( a2035a );
 a2053a <=( a1600a ) or ( a1601a );
 a2054a <=( a1602a ) or ( a2053a );
 a2057a <=( a1598a ) or ( a1599a );
 a2060a <=( a1596a ) or ( a1597a );
 a2061a <=( a2060a ) or ( a2057a );
 a2062a <=( a2061a ) or ( a2054a );
 a2066a <=( a1593a ) or ( a1594a );
 a2067a <=( a1595a ) or ( a2066a );
 a2070a <=( a1591a ) or ( a1592a );
 a2073a <=( a1589a ) or ( a1590a );
 a2074a <=( a2073a ) or ( a2070a );
 a2075a <=( a2074a ) or ( a2067a );
 a2076a <=( a2075a ) or ( a2062a );
 a2077a <=( a2076a ) or ( a2049a );
 a2078a <=( a2077a ) or ( a2022a );
 a2082a <=( a1586a ) or ( a1587a );
 a2083a <=( a1588a ) or ( a2082a );
 a2087a <=( a1583a ) or ( a1584a );
 a2088a <=( a1585a ) or ( a2087a );
 a2089a <=( a2088a ) or ( a2083a );
 a2093a <=( a1580a ) or ( a1581a );
 a2094a <=( a1582a ) or ( a2093a );
 a2097a <=( a1578a ) or ( a1579a );
 a2100a <=( a1576a ) or ( a1577a );
 a2101a <=( a2100a ) or ( a2097a );
 a2102a <=( a2101a ) or ( a2094a );
 a2103a <=( a2102a ) or ( a2089a );
 a2107a <=( a1573a ) or ( a1574a );
 a2108a <=( a1575a ) or ( a2107a );
 a2111a <=( a1571a ) or ( a1572a );
 a2114a <=( a1569a ) or ( a1570a );
 a2115a <=( a2114a ) or ( a2111a );
 a2116a <=( a2115a ) or ( a2108a );
 a2120a <=( a1566a ) or ( a1567a );
 a2121a <=( a1568a ) or ( a2120a );
 a2124a <=( a1564a ) or ( a1565a );
 a2127a <=( a1562a ) or ( a1563a );
 a2128a <=( a2127a ) or ( a2124a );
 a2129a <=( a2128a ) or ( a2121a );
 a2130a <=( a2129a ) or ( a2116a );
 a2131a <=( a2130a ) or ( a2103a );
 a2135a <=( a1559a ) or ( a1560a );
 a2136a <=( a1561a ) or ( a2135a );
 a2139a <=( a1557a ) or ( a1558a );
 a2142a <=( a1555a ) or ( a1556a );
 a2143a <=( a2142a ) or ( a2139a );
 a2144a <=( a2143a ) or ( a2136a );
 a2148a <=( a1552a ) or ( a1553a );
 a2149a <=( a1554a ) or ( a2148a );
 a2152a <=( a1550a ) or ( a1551a );
 a2155a <=( a1548a ) or ( a1549a );
 a2156a <=( a2155a ) or ( a2152a );
 a2157a <=( a2156a ) or ( a2149a );
 a2158a <=( a2157a ) or ( a2144a );
 a2162a <=( a1545a ) or ( a1546a );
 a2163a <=( a1547a ) or ( a2162a );
 a2166a <=( a1543a ) or ( a1544a );
 a2169a <=( a1541a ) or ( a1542a );
 a2170a <=( a2169a ) or ( a2166a );
 a2171a <=( a2170a ) or ( a2163a );
 a2175a <=( a1538a ) or ( a1539a );
 a2176a <=( a1540a ) or ( a2175a );
 a2179a <=( a1536a ) or ( a1537a );
 a2182a <=( a1534a ) or ( a1535a );
 a2183a <=( a2182a ) or ( a2179a );
 a2184a <=( a2183a ) or ( a2176a );
 a2185a <=( a2184a ) or ( a2171a );
 a2186a <=( a2185a ) or ( a2158a );
 a2187a <=( a2186a ) or ( a2131a );
 a2188a <=( a2187a ) or ( a2078a );
 a2189a <=( a2188a ) or ( a1969a );
 a2193a <=( a1531a ) or ( a1532a );
 a2194a <=( a1533a ) or ( a2193a );
 a2198a <=( a1528a ) or ( a1529a );
 a2199a <=( a1530a ) or ( a2198a );
 a2200a <=( a2199a ) or ( a2194a );
 a2204a <=( a1525a ) or ( a1526a );
 a2205a <=( a1527a ) or ( a2204a );
 a2208a <=( a1523a ) or ( a1524a );
 a2211a <=( a1521a ) or ( a1522a );
 a2212a <=( a2211a ) or ( a2208a );
 a2213a <=( a2212a ) or ( a2205a );
 a2214a <=( a2213a ) or ( a2200a );
 a2218a <=( a1518a ) or ( a1519a );
 a2219a <=( a1520a ) or ( a2218a );
 a2222a <=( a1516a ) or ( a1517a );
 a2225a <=( a1514a ) or ( a1515a );
 a2226a <=( a2225a ) or ( a2222a );
 a2227a <=( a2226a ) or ( a2219a );
 a2231a <=( a1511a ) or ( a1512a );
 a2232a <=( a1513a ) or ( a2231a );
 a2235a <=( a1509a ) or ( a1510a );
 a2238a <=( a1507a ) or ( a1508a );
 a2239a <=( a2238a ) or ( a2235a );
 a2240a <=( a2239a ) or ( a2232a );
 a2241a <=( a2240a ) or ( a2227a );
 a2242a <=( a2241a ) or ( a2214a );
 a2246a <=( a1504a ) or ( a1505a );
 a2247a <=( a1506a ) or ( a2246a );
 a2251a <=( a1501a ) or ( a1502a );
 a2252a <=( a1503a ) or ( a2251a );
 a2253a <=( a2252a ) or ( a2247a );
 a2257a <=( a1498a ) or ( a1499a );
 a2258a <=( a1500a ) or ( a2257a );
 a2261a <=( a1496a ) or ( a1497a );
 a2264a <=( a1494a ) or ( a1495a );
 a2265a <=( a2264a ) or ( a2261a );
 a2266a <=( a2265a ) or ( a2258a );
 a2267a <=( a2266a ) or ( a2253a );
 a2271a <=( a1491a ) or ( a1492a );
 a2272a <=( a1493a ) or ( a2271a );
 a2275a <=( a1489a ) or ( a1490a );
 a2278a <=( a1487a ) or ( a1488a );
 a2279a <=( a2278a ) or ( a2275a );
 a2280a <=( a2279a ) or ( a2272a );
 a2284a <=( a1484a ) or ( a1485a );
 a2285a <=( a1486a ) or ( a2284a );
 a2288a <=( a1482a ) or ( a1483a );
 a2291a <=( a1480a ) or ( a1481a );
 a2292a <=( a2291a ) or ( a2288a );
 a2293a <=( a2292a ) or ( a2285a );
 a2294a <=( a2293a ) or ( a2280a );
 a2295a <=( a2294a ) or ( a2267a );
 a2296a <=( a2295a ) or ( a2242a );
 a2300a <=( a1477a ) or ( a1478a );
 a2301a <=( a1479a ) or ( a2300a );
 a2305a <=( a1474a ) or ( a1475a );
 a2306a <=( a1476a ) or ( a2305a );
 a2307a <=( a2306a ) or ( a2301a );
 a2311a <=( a1471a ) or ( a1472a );
 a2312a <=( a1473a ) or ( a2311a );
 a2315a <=( a1469a ) or ( a1470a );
 a2318a <=( a1467a ) or ( a1468a );
 a2319a <=( a2318a ) or ( a2315a );
 a2320a <=( a2319a ) or ( a2312a );
 a2321a <=( a2320a ) or ( a2307a );
 a2325a <=( a1464a ) or ( a1465a );
 a2326a <=( a1466a ) or ( a2325a );
 a2329a <=( a1462a ) or ( a1463a );
 a2332a <=( a1460a ) or ( a1461a );
 a2333a <=( a2332a ) or ( a2329a );
 a2334a <=( a2333a ) or ( a2326a );
 a2338a <=( a1457a ) or ( a1458a );
 a2339a <=( a1459a ) or ( a2338a );
 a2342a <=( a1455a ) or ( a1456a );
 a2345a <=( a1453a ) or ( a1454a );
 a2346a <=( a2345a ) or ( a2342a );
 a2347a <=( a2346a ) or ( a2339a );
 a2348a <=( a2347a ) or ( a2334a );
 a2349a <=( a2348a ) or ( a2321a );
 a2353a <=( a1450a ) or ( a1451a );
 a2354a <=( a1452a ) or ( a2353a );
 a2357a <=( a1448a ) or ( a1449a );
 a2360a <=( a1446a ) or ( a1447a );
 a2361a <=( a2360a ) or ( a2357a );
 a2362a <=( a2361a ) or ( a2354a );
 a2366a <=( a1443a ) or ( a1444a );
 a2367a <=( a1445a ) or ( a2366a );
 a2370a <=( a1441a ) or ( a1442a );
 a2373a <=( a1439a ) or ( a1440a );
 a2374a <=( a2373a ) or ( a2370a );
 a2375a <=( a2374a ) or ( a2367a );
 a2376a <=( a2375a ) or ( a2362a );
 a2380a <=( a1436a ) or ( a1437a );
 a2381a <=( a1438a ) or ( a2380a );
 a2384a <=( a1434a ) or ( a1435a );
 a2387a <=( a1432a ) or ( a1433a );
 a2388a <=( a2387a ) or ( a2384a );
 a2389a <=( a2388a ) or ( a2381a );
 a2393a <=( a1429a ) or ( a1430a );
 a2394a <=( a1431a ) or ( a2393a );
 a2397a <=( a1427a ) or ( a1428a );
 a2400a <=( a1425a ) or ( a1426a );
 a2401a <=( a2400a ) or ( a2397a );
 a2402a <=( a2401a ) or ( a2394a );
 a2403a <=( a2402a ) or ( a2389a );
 a2404a <=( a2403a ) or ( a2376a );
 a2405a <=( a2404a ) or ( a2349a );
 a2406a <=( a2405a ) or ( a2296a );
 a2410a <=( a1422a ) or ( a1423a );
 a2411a <=( a1424a ) or ( a2410a );
 a2415a <=( a1419a ) or ( a1420a );
 a2416a <=( a1421a ) or ( a2415a );
 a2417a <=( a2416a ) or ( a2411a );
 a2421a <=( a1416a ) or ( a1417a );
 a2422a <=( a1418a ) or ( a2421a );
 a2425a <=( a1414a ) or ( a1415a );
 a2428a <=( a1412a ) or ( a1413a );
 a2429a <=( a2428a ) or ( a2425a );
 a2430a <=( a2429a ) or ( a2422a );
 a2431a <=( a2430a ) or ( a2417a );
 a2435a <=( a1409a ) or ( a1410a );
 a2436a <=( a1411a ) or ( a2435a );
 a2439a <=( a1407a ) or ( a1408a );
 a2442a <=( a1405a ) or ( a1406a );
 a2443a <=( a2442a ) or ( a2439a );
 a2444a <=( a2443a ) or ( a2436a );
 a2448a <=( a1402a ) or ( a1403a );
 a2449a <=( a1404a ) or ( a2448a );
 a2452a <=( a1400a ) or ( a1401a );
 a2455a <=( a1398a ) or ( a1399a );
 a2456a <=( a2455a ) or ( a2452a );
 a2457a <=( a2456a ) or ( a2449a );
 a2458a <=( a2457a ) or ( a2444a );
 a2459a <=( a2458a ) or ( a2431a );
 a2463a <=( a1395a ) or ( a1396a );
 a2464a <=( a1397a ) or ( a2463a );
 a2467a <=( a1393a ) or ( a1394a );
 a2470a <=( a1391a ) or ( a1392a );
 a2471a <=( a2470a ) or ( a2467a );
 a2472a <=( a2471a ) or ( a2464a );
 a2476a <=( a1388a ) or ( a1389a );
 a2477a <=( a1390a ) or ( a2476a );
 a2480a <=( a1386a ) or ( a1387a );
 a2483a <=( a1384a ) or ( a1385a );
 a2484a <=( a2483a ) or ( a2480a );
 a2485a <=( a2484a ) or ( a2477a );
 a2486a <=( a2485a ) or ( a2472a );
 a2490a <=( a1381a ) or ( a1382a );
 a2491a <=( a1383a ) or ( a2490a );
 a2494a <=( a1379a ) or ( a1380a );
 a2497a <=( a1377a ) or ( a1378a );
 a2498a <=( a2497a ) or ( a2494a );
 a2499a <=( a2498a ) or ( a2491a );
 a2503a <=( a1374a ) or ( a1375a );
 a2504a <=( a1376a ) or ( a2503a );
 a2507a <=( a1372a ) or ( a1373a );
 a2510a <=( a1370a ) or ( a1371a );
 a2511a <=( a2510a ) or ( a2507a );
 a2512a <=( a2511a ) or ( a2504a );
 a2513a <=( a2512a ) or ( a2499a );
 a2514a <=( a2513a ) or ( a2486a );
 a2515a <=( a2514a ) or ( a2459a );
 a2519a <=( a1367a ) or ( a1368a );
 a2520a <=( a1369a ) or ( a2519a );
 a2524a <=( a1364a ) or ( a1365a );
 a2525a <=( a1366a ) or ( a2524a );
 a2526a <=( a2525a ) or ( a2520a );
 a2530a <=( a1361a ) or ( a1362a );
 a2531a <=( a1363a ) or ( a2530a );
 a2534a <=( a1359a ) or ( a1360a );
 a2537a <=( a1357a ) or ( a1358a );
 a2538a <=( a2537a ) or ( a2534a );
 a2539a <=( a2538a ) or ( a2531a );
 a2540a <=( a2539a ) or ( a2526a );
 a2544a <=( a1354a ) or ( a1355a );
 a2545a <=( a1356a ) or ( a2544a );
 a2548a <=( a1352a ) or ( a1353a );
 a2551a <=( a1350a ) or ( a1351a );
 a2552a <=( a2551a ) or ( a2548a );
 a2553a <=( a2552a ) or ( a2545a );
 a2557a <=( a1347a ) or ( a1348a );
 a2558a <=( a1349a ) or ( a2557a );
 a2561a <=( a1345a ) or ( a1346a );
 a2564a <=( a1343a ) or ( a1344a );
 a2565a <=( a2564a ) or ( a2561a );
 a2566a <=( a2565a ) or ( a2558a );
 a2567a <=( a2566a ) or ( a2553a );
 a2568a <=( a2567a ) or ( a2540a );
 a2572a <=( a1340a ) or ( a1341a );
 a2573a <=( a1342a ) or ( a2572a );
 a2576a <=( a1338a ) or ( a1339a );
 a2579a <=( a1336a ) or ( a1337a );
 a2580a <=( a2579a ) or ( a2576a );
 a2581a <=( a2580a ) or ( a2573a );
 a2585a <=( a1333a ) or ( a1334a );
 a2586a <=( a1335a ) or ( a2585a );
 a2589a <=( a1331a ) or ( a1332a );
 a2592a <=( a1329a ) or ( a1330a );
 a2593a <=( a2592a ) or ( a2589a );
 a2594a <=( a2593a ) or ( a2586a );
 a2595a <=( a2594a ) or ( a2581a );
 a2599a <=( a1326a ) or ( a1327a );
 a2600a <=( a1328a ) or ( a2599a );
 a2603a <=( a1324a ) or ( a1325a );
 a2606a <=( a1322a ) or ( a1323a );
 a2607a <=( a2606a ) or ( a2603a );
 a2608a <=( a2607a ) or ( a2600a );
 a2612a <=( a1319a ) or ( a1320a );
 a2613a <=( a1321a ) or ( a2612a );
 a2616a <=( a1317a ) or ( a1318a );
 a2619a <=( a1315a ) or ( a1316a );
 a2620a <=( a2619a ) or ( a2616a );
 a2621a <=( a2620a ) or ( a2613a );
 a2622a <=( a2621a ) or ( a2608a );
 a2623a <=( a2622a ) or ( a2595a );
 a2624a <=( a2623a ) or ( a2568a );
 a2625a <=( a2624a ) or ( a2515a );
 a2626a <=( a2625a ) or ( a2406a );
 a2627a <=( a2626a ) or ( a2189a );
 a2631a <=( a1312a ) or ( a1313a );
 a2632a <=( a1314a ) or ( a2631a );
 a2636a <=( a1309a ) or ( a1310a );
 a2637a <=( a1311a ) or ( a2636a );
 a2638a <=( a2637a ) or ( a2632a );
 a2642a <=( a1306a ) or ( a1307a );
 a2643a <=( a1308a ) or ( a2642a );
 a2646a <=( a1304a ) or ( a1305a );
 a2649a <=( a1302a ) or ( a1303a );
 a2650a <=( a2649a ) or ( a2646a );
 a2651a <=( a2650a ) or ( a2643a );
 a2652a <=( a2651a ) or ( a2638a );
 a2656a <=( a1299a ) or ( a1300a );
 a2657a <=( a1301a ) or ( a2656a );
 a2660a <=( a1297a ) or ( a1298a );
 a2663a <=( a1295a ) or ( a1296a );
 a2664a <=( a2663a ) or ( a2660a );
 a2665a <=( a2664a ) or ( a2657a );
 a2669a <=( a1292a ) or ( a1293a );
 a2670a <=( a1294a ) or ( a2669a );
 a2673a <=( a1290a ) or ( a1291a );
 a2676a <=( a1288a ) or ( a1289a );
 a2677a <=( a2676a ) or ( a2673a );
 a2678a <=( a2677a ) or ( a2670a );
 a2679a <=( a2678a ) or ( a2665a );
 a2680a <=( a2679a ) or ( a2652a );
 a2684a <=( a1285a ) or ( a1286a );
 a2685a <=( a1287a ) or ( a2684a );
 a2689a <=( a1282a ) or ( a1283a );
 a2690a <=( a1284a ) or ( a2689a );
 a2691a <=( a2690a ) or ( a2685a );
 a2695a <=( a1279a ) or ( a1280a );
 a2696a <=( a1281a ) or ( a2695a );
 a2699a <=( a1277a ) or ( a1278a );
 a2702a <=( a1275a ) or ( a1276a );
 a2703a <=( a2702a ) or ( a2699a );
 a2704a <=( a2703a ) or ( a2696a );
 a2705a <=( a2704a ) or ( a2691a );
 a2709a <=( a1272a ) or ( a1273a );
 a2710a <=( a1274a ) or ( a2709a );
 a2713a <=( a1270a ) or ( a1271a );
 a2716a <=( a1268a ) or ( a1269a );
 a2717a <=( a2716a ) or ( a2713a );
 a2718a <=( a2717a ) or ( a2710a );
 a2722a <=( a1265a ) or ( a1266a );
 a2723a <=( a1267a ) or ( a2722a );
 a2726a <=( a1263a ) or ( a1264a );
 a2729a <=( a1261a ) or ( a1262a );
 a2730a <=( a2729a ) or ( a2726a );
 a2731a <=( a2730a ) or ( a2723a );
 a2732a <=( a2731a ) or ( a2718a );
 a2733a <=( a2732a ) or ( a2705a );
 a2734a <=( a2733a ) or ( a2680a );
 a2738a <=( a1258a ) or ( a1259a );
 a2739a <=( a1260a ) or ( a2738a );
 a2743a <=( a1255a ) or ( a1256a );
 a2744a <=( a1257a ) or ( a2743a );
 a2745a <=( a2744a ) or ( a2739a );
 a2749a <=( a1252a ) or ( a1253a );
 a2750a <=( a1254a ) or ( a2749a );
 a2753a <=( a1250a ) or ( a1251a );
 a2756a <=( a1248a ) or ( a1249a );
 a2757a <=( a2756a ) or ( a2753a );
 a2758a <=( a2757a ) or ( a2750a );
 a2759a <=( a2758a ) or ( a2745a );
 a2763a <=( a1245a ) or ( a1246a );
 a2764a <=( a1247a ) or ( a2763a );
 a2767a <=( a1243a ) or ( a1244a );
 a2770a <=( a1241a ) or ( a1242a );
 a2771a <=( a2770a ) or ( a2767a );
 a2772a <=( a2771a ) or ( a2764a );
 a2776a <=( a1238a ) or ( a1239a );
 a2777a <=( a1240a ) or ( a2776a );
 a2780a <=( a1236a ) or ( a1237a );
 a2783a <=( a1234a ) or ( a1235a );
 a2784a <=( a2783a ) or ( a2780a );
 a2785a <=( a2784a ) or ( a2777a );
 a2786a <=( a2785a ) or ( a2772a );
 a2787a <=( a2786a ) or ( a2759a );
 a2791a <=( a1231a ) or ( a1232a );
 a2792a <=( a1233a ) or ( a2791a );
 a2795a <=( a1229a ) or ( a1230a );
 a2798a <=( a1227a ) or ( a1228a );
 a2799a <=( a2798a ) or ( a2795a );
 a2800a <=( a2799a ) or ( a2792a );
 a2804a <=( a1224a ) or ( a1225a );
 a2805a <=( a1226a ) or ( a2804a );
 a2808a <=( a1222a ) or ( a1223a );
 a2811a <=( a1220a ) or ( a1221a );
 a2812a <=( a2811a ) or ( a2808a );
 a2813a <=( a2812a ) or ( a2805a );
 a2814a <=( a2813a ) or ( a2800a );
 a2818a <=( a1217a ) or ( a1218a );
 a2819a <=( a1219a ) or ( a2818a );
 a2822a <=( a1215a ) or ( a1216a );
 a2825a <=( a1213a ) or ( a1214a );
 a2826a <=( a2825a ) or ( a2822a );
 a2827a <=( a2826a ) or ( a2819a );
 a2831a <=( a1210a ) or ( a1211a );
 a2832a <=( a1212a ) or ( a2831a );
 a2835a <=( a1208a ) or ( a1209a );
 a2838a <=( a1206a ) or ( a1207a );
 a2839a <=( a2838a ) or ( a2835a );
 a2840a <=( a2839a ) or ( a2832a );
 a2841a <=( a2840a ) or ( a2827a );
 a2842a <=( a2841a ) or ( a2814a );
 a2843a <=( a2842a ) or ( a2787a );
 a2844a <=( a2843a ) or ( a2734a );
 a2848a <=( a1203a ) or ( a1204a );
 a2849a <=( a1205a ) or ( a2848a );
 a2853a <=( a1200a ) or ( a1201a );
 a2854a <=( a1202a ) or ( a2853a );
 a2855a <=( a2854a ) or ( a2849a );
 a2859a <=( a1197a ) or ( a1198a );
 a2860a <=( a1199a ) or ( a2859a );
 a2863a <=( a1195a ) or ( a1196a );
 a2866a <=( a1193a ) or ( a1194a );
 a2867a <=( a2866a ) or ( a2863a );
 a2868a <=( a2867a ) or ( a2860a );
 a2869a <=( a2868a ) or ( a2855a );
 a2873a <=( a1190a ) or ( a1191a );
 a2874a <=( a1192a ) or ( a2873a );
 a2877a <=( a1188a ) or ( a1189a );
 a2880a <=( a1186a ) or ( a1187a );
 a2881a <=( a2880a ) or ( a2877a );
 a2882a <=( a2881a ) or ( a2874a );
 a2886a <=( a1183a ) or ( a1184a );
 a2887a <=( a1185a ) or ( a2886a );
 a2890a <=( a1181a ) or ( a1182a );
 a2893a <=( a1179a ) or ( a1180a );
 a2894a <=( a2893a ) or ( a2890a );
 a2895a <=( a2894a ) or ( a2887a );
 a2896a <=( a2895a ) or ( a2882a );
 a2897a <=( a2896a ) or ( a2869a );
 a2901a <=( a1176a ) or ( a1177a );
 a2902a <=( a1178a ) or ( a2901a );
 a2905a <=( a1174a ) or ( a1175a );
 a2908a <=( a1172a ) or ( a1173a );
 a2909a <=( a2908a ) or ( a2905a );
 a2910a <=( a2909a ) or ( a2902a );
 a2914a <=( a1169a ) or ( a1170a );
 a2915a <=( a1171a ) or ( a2914a );
 a2918a <=( a1167a ) or ( a1168a );
 a2921a <=( a1165a ) or ( a1166a );
 a2922a <=( a2921a ) or ( a2918a );
 a2923a <=( a2922a ) or ( a2915a );
 a2924a <=( a2923a ) or ( a2910a );
 a2928a <=( a1162a ) or ( a1163a );
 a2929a <=( a1164a ) or ( a2928a );
 a2932a <=( a1160a ) or ( a1161a );
 a2935a <=( a1158a ) or ( a1159a );
 a2936a <=( a2935a ) or ( a2932a );
 a2937a <=( a2936a ) or ( a2929a );
 a2941a <=( a1155a ) or ( a1156a );
 a2942a <=( a1157a ) or ( a2941a );
 a2945a <=( a1153a ) or ( a1154a );
 a2948a <=( a1151a ) or ( a1152a );
 a2949a <=( a2948a ) or ( a2945a );
 a2950a <=( a2949a ) or ( a2942a );
 a2951a <=( a2950a ) or ( a2937a );
 a2952a <=( a2951a ) or ( a2924a );
 a2953a <=( a2952a ) or ( a2897a );
 a2957a <=( a1148a ) or ( a1149a );
 a2958a <=( a1150a ) or ( a2957a );
 a2962a <=( a1145a ) or ( a1146a );
 a2963a <=( a1147a ) or ( a2962a );
 a2964a <=( a2963a ) or ( a2958a );
 a2968a <=( a1142a ) or ( a1143a );
 a2969a <=( a1144a ) or ( a2968a );
 a2972a <=( a1140a ) or ( a1141a );
 a2975a <=( a1138a ) or ( a1139a );
 a2976a <=( a2975a ) or ( a2972a );
 a2977a <=( a2976a ) or ( a2969a );
 a2978a <=( a2977a ) or ( a2964a );
 a2982a <=( a1135a ) or ( a1136a );
 a2983a <=( a1137a ) or ( a2982a );
 a2986a <=( a1133a ) or ( a1134a );
 a2989a <=( a1131a ) or ( a1132a );
 a2990a <=( a2989a ) or ( a2986a );
 a2991a <=( a2990a ) or ( a2983a );
 a2995a <=( a1128a ) or ( a1129a );
 a2996a <=( a1130a ) or ( a2995a );
 a2999a <=( a1126a ) or ( a1127a );
 a3002a <=( a1124a ) or ( a1125a );
 a3003a <=( a3002a ) or ( a2999a );
 a3004a <=( a3003a ) or ( a2996a );
 a3005a <=( a3004a ) or ( a2991a );
 a3006a <=( a3005a ) or ( a2978a );
 a3010a <=( a1121a ) or ( a1122a );
 a3011a <=( a1123a ) or ( a3010a );
 a3014a <=( a1119a ) or ( a1120a );
 a3017a <=( a1117a ) or ( a1118a );
 a3018a <=( a3017a ) or ( a3014a );
 a3019a <=( a3018a ) or ( a3011a );
 a3023a <=( a1114a ) or ( a1115a );
 a3024a <=( a1116a ) or ( a3023a );
 a3027a <=( a1112a ) or ( a1113a );
 a3030a <=( a1110a ) or ( a1111a );
 a3031a <=( a3030a ) or ( a3027a );
 a3032a <=( a3031a ) or ( a3024a );
 a3033a <=( a3032a ) or ( a3019a );
 a3037a <=( a1107a ) or ( a1108a );
 a3038a <=( a1109a ) or ( a3037a );
 a3041a <=( a1105a ) or ( a1106a );
 a3044a <=( a1103a ) or ( a1104a );
 a3045a <=( a3044a ) or ( a3041a );
 a3046a <=( a3045a ) or ( a3038a );
 a3050a <=( a1100a ) or ( a1101a );
 a3051a <=( a1102a ) or ( a3050a );
 a3054a <=( a1098a ) or ( a1099a );
 a3057a <=( a1096a ) or ( a1097a );
 a3058a <=( a3057a ) or ( a3054a );
 a3059a <=( a3058a ) or ( a3051a );
 a3060a <=( a3059a ) or ( a3046a );
 a3061a <=( a3060a ) or ( a3033a );
 a3062a <=( a3061a ) or ( a3006a );
 a3063a <=( a3062a ) or ( a2953a );
 a3064a <=( a3063a ) or ( a2844a );
 a3068a <=( a1093a ) or ( a1094a );
 a3069a <=( a1095a ) or ( a3068a );
 a3073a <=( a1090a ) or ( a1091a );
 a3074a <=( a1092a ) or ( a3073a );
 a3075a <=( a3074a ) or ( a3069a );
 a3079a <=( a1087a ) or ( a1088a );
 a3080a <=( a1089a ) or ( a3079a );
 a3083a <=( a1085a ) or ( a1086a );
 a3086a <=( a1083a ) or ( a1084a );
 a3087a <=( a3086a ) or ( a3083a );
 a3088a <=( a3087a ) or ( a3080a );
 a3089a <=( a3088a ) or ( a3075a );
 a3093a <=( a1080a ) or ( a1081a );
 a3094a <=( a1082a ) or ( a3093a );
 a3097a <=( a1078a ) or ( a1079a );
 a3100a <=( a1076a ) or ( a1077a );
 a3101a <=( a3100a ) or ( a3097a );
 a3102a <=( a3101a ) or ( a3094a );
 a3106a <=( a1073a ) or ( a1074a );
 a3107a <=( a1075a ) or ( a3106a );
 a3110a <=( a1071a ) or ( a1072a );
 a3113a <=( a1069a ) or ( a1070a );
 a3114a <=( a3113a ) or ( a3110a );
 a3115a <=( a3114a ) or ( a3107a );
 a3116a <=( a3115a ) or ( a3102a );
 a3117a <=( a3116a ) or ( a3089a );
 a3121a <=( a1066a ) or ( a1067a );
 a3122a <=( a1068a ) or ( a3121a );
 a3126a <=( a1063a ) or ( a1064a );
 a3127a <=( a1065a ) or ( a3126a );
 a3128a <=( a3127a ) or ( a3122a );
 a3132a <=( a1060a ) or ( a1061a );
 a3133a <=( a1062a ) or ( a3132a );
 a3136a <=( a1058a ) or ( a1059a );
 a3139a <=( a1056a ) or ( a1057a );
 a3140a <=( a3139a ) or ( a3136a );
 a3141a <=( a3140a ) or ( a3133a );
 a3142a <=( a3141a ) or ( a3128a );
 a3146a <=( a1053a ) or ( a1054a );
 a3147a <=( a1055a ) or ( a3146a );
 a3150a <=( a1051a ) or ( a1052a );
 a3153a <=( a1049a ) or ( a1050a );
 a3154a <=( a3153a ) or ( a3150a );
 a3155a <=( a3154a ) or ( a3147a );
 a3159a <=( a1046a ) or ( a1047a );
 a3160a <=( a1048a ) or ( a3159a );
 a3163a <=( a1044a ) or ( a1045a );
 a3166a <=( a1042a ) or ( a1043a );
 a3167a <=( a3166a ) or ( a3163a );
 a3168a <=( a3167a ) or ( a3160a );
 a3169a <=( a3168a ) or ( a3155a );
 a3170a <=( a3169a ) or ( a3142a );
 a3171a <=( a3170a ) or ( a3117a );
 a3175a <=( a1039a ) or ( a1040a );
 a3176a <=( a1041a ) or ( a3175a );
 a3180a <=( a1036a ) or ( a1037a );
 a3181a <=( a1038a ) or ( a3180a );
 a3182a <=( a3181a ) or ( a3176a );
 a3186a <=( a1033a ) or ( a1034a );
 a3187a <=( a1035a ) or ( a3186a );
 a3190a <=( a1031a ) or ( a1032a );
 a3193a <=( a1029a ) or ( a1030a );
 a3194a <=( a3193a ) or ( a3190a );
 a3195a <=( a3194a ) or ( a3187a );
 a3196a <=( a3195a ) or ( a3182a );
 a3200a <=( a1026a ) or ( a1027a );
 a3201a <=( a1028a ) or ( a3200a );
 a3204a <=( a1024a ) or ( a1025a );
 a3207a <=( a1022a ) or ( a1023a );
 a3208a <=( a3207a ) or ( a3204a );
 a3209a <=( a3208a ) or ( a3201a );
 a3213a <=( a1019a ) or ( a1020a );
 a3214a <=( a1021a ) or ( a3213a );
 a3217a <=( a1017a ) or ( a1018a );
 a3220a <=( a1015a ) or ( a1016a );
 a3221a <=( a3220a ) or ( a3217a );
 a3222a <=( a3221a ) or ( a3214a );
 a3223a <=( a3222a ) or ( a3209a );
 a3224a <=( a3223a ) or ( a3196a );
 a3228a <=( a1012a ) or ( a1013a );
 a3229a <=( a1014a ) or ( a3228a );
 a3232a <=( a1010a ) or ( a1011a );
 a3235a <=( a1008a ) or ( a1009a );
 a3236a <=( a3235a ) or ( a3232a );
 a3237a <=( a3236a ) or ( a3229a );
 a3241a <=( a1005a ) or ( a1006a );
 a3242a <=( a1007a ) or ( a3241a );
 a3245a <=( a1003a ) or ( a1004a );
 a3248a <=( a1001a ) or ( a1002a );
 a3249a <=( a3248a ) or ( a3245a );
 a3250a <=( a3249a ) or ( a3242a );
 a3251a <=( a3250a ) or ( a3237a );
 a3255a <=( a998a ) or ( a999a );
 a3256a <=( a1000a ) or ( a3255a );
 a3259a <=( a996a ) or ( a997a );
 a3262a <=( a994a ) or ( a995a );
 a3263a <=( a3262a ) or ( a3259a );
 a3264a <=( a3263a ) or ( a3256a );
 a3268a <=( a991a ) or ( a992a );
 a3269a <=( a993a ) or ( a3268a );
 a3272a <=( a989a ) or ( a990a );
 a3275a <=( a987a ) or ( a988a );
 a3276a <=( a3275a ) or ( a3272a );
 a3277a <=( a3276a ) or ( a3269a );
 a3278a <=( a3277a ) or ( a3264a );
 a3279a <=( a3278a ) or ( a3251a );
 a3280a <=( a3279a ) or ( a3224a );
 a3281a <=( a3280a ) or ( a3171a );
 a3285a <=( a984a ) or ( a985a );
 a3286a <=( a986a ) or ( a3285a );
 a3290a <=( a981a ) or ( a982a );
 a3291a <=( a983a ) or ( a3290a );
 a3292a <=( a3291a ) or ( a3286a );
 a3296a <=( a978a ) or ( a979a );
 a3297a <=( a980a ) or ( a3296a );
 a3300a <=( a976a ) or ( a977a );
 a3303a <=( a974a ) or ( a975a );
 a3304a <=( a3303a ) or ( a3300a );
 a3305a <=( a3304a ) or ( a3297a );
 a3306a <=( a3305a ) or ( a3292a );
 a3310a <=( a971a ) or ( a972a );
 a3311a <=( a973a ) or ( a3310a );
 a3314a <=( a969a ) or ( a970a );
 a3317a <=( a967a ) or ( a968a );
 a3318a <=( a3317a ) or ( a3314a );
 a3319a <=( a3318a ) or ( a3311a );
 a3323a <=( a964a ) or ( a965a );
 a3324a <=( a966a ) or ( a3323a );
 a3327a <=( a962a ) or ( a963a );
 a3330a <=( a960a ) or ( a961a );
 a3331a <=( a3330a ) or ( a3327a );
 a3332a <=( a3331a ) or ( a3324a );
 a3333a <=( a3332a ) or ( a3319a );
 a3334a <=( a3333a ) or ( a3306a );
 a3338a <=( a957a ) or ( a958a );
 a3339a <=( a959a ) or ( a3338a );
 a3342a <=( a955a ) or ( a956a );
 a3345a <=( a953a ) or ( a954a );
 a3346a <=( a3345a ) or ( a3342a );
 a3347a <=( a3346a ) or ( a3339a );
 a3351a <=( a950a ) or ( a951a );
 a3352a <=( a952a ) or ( a3351a );
 a3355a <=( a948a ) or ( a949a );
 a3358a <=( a946a ) or ( a947a );
 a3359a <=( a3358a ) or ( a3355a );
 a3360a <=( a3359a ) or ( a3352a );
 a3361a <=( a3360a ) or ( a3347a );
 a3365a <=( a943a ) or ( a944a );
 a3366a <=( a945a ) or ( a3365a );
 a3369a <=( a941a ) or ( a942a );
 a3372a <=( a939a ) or ( a940a );
 a3373a <=( a3372a ) or ( a3369a );
 a3374a <=( a3373a ) or ( a3366a );
 a3378a <=( a936a ) or ( a937a );
 a3379a <=( a938a ) or ( a3378a );
 a3382a <=( a934a ) or ( a935a );
 a3385a <=( a932a ) or ( a933a );
 a3386a <=( a3385a ) or ( a3382a );
 a3387a <=( a3386a ) or ( a3379a );
 a3388a <=( a3387a ) or ( a3374a );
 a3389a <=( a3388a ) or ( a3361a );
 a3390a <=( a3389a ) or ( a3334a );
 a3394a <=( a929a ) or ( a930a );
 a3395a <=( a931a ) or ( a3394a );
 a3399a <=( a926a ) or ( a927a );
 a3400a <=( a928a ) or ( a3399a );
 a3401a <=( a3400a ) or ( a3395a );
 a3405a <=( a923a ) or ( a924a );
 a3406a <=( a925a ) or ( a3405a );
 a3409a <=( a921a ) or ( a922a );
 a3412a <=( a919a ) or ( a920a );
 a3413a <=( a3412a ) or ( a3409a );
 a3414a <=( a3413a ) or ( a3406a );
 a3415a <=( a3414a ) or ( a3401a );
 a3419a <=( a916a ) or ( a917a );
 a3420a <=( a918a ) or ( a3419a );
 a3423a <=( a914a ) or ( a915a );
 a3426a <=( a912a ) or ( a913a );
 a3427a <=( a3426a ) or ( a3423a );
 a3428a <=( a3427a ) or ( a3420a );
 a3432a <=( a909a ) or ( a910a );
 a3433a <=( a911a ) or ( a3432a );
 a3436a <=( a907a ) or ( a908a );
 a3439a <=( a905a ) or ( a906a );
 a3440a <=( a3439a ) or ( a3436a );
 a3441a <=( a3440a ) or ( a3433a );
 a3442a <=( a3441a ) or ( a3428a );
 a3443a <=( a3442a ) or ( a3415a );
 a3447a <=( a902a ) or ( a903a );
 a3448a <=( a904a ) or ( a3447a );
 a3451a <=( a900a ) or ( a901a );
 a3454a <=( a898a ) or ( a899a );
 a3455a <=( a3454a ) or ( a3451a );
 a3456a <=( a3455a ) or ( a3448a );
 a3460a <=( a895a ) or ( a896a );
 a3461a <=( a897a ) or ( a3460a );
 a3464a <=( a893a ) or ( a894a );
 a3467a <=( a891a ) or ( a892a );
 a3468a <=( a3467a ) or ( a3464a );
 a3469a <=( a3468a ) or ( a3461a );
 a3470a <=( a3469a ) or ( a3456a );
 a3474a <=( a888a ) or ( a889a );
 a3475a <=( a890a ) or ( a3474a );
 a3478a <=( a886a ) or ( a887a );
 a3481a <=( a884a ) or ( a885a );
 a3482a <=( a3481a ) or ( a3478a );
 a3483a <=( a3482a ) or ( a3475a );
 a3487a <=( a881a ) or ( a882a );
 a3488a <=( a883a ) or ( a3487a );
 a3491a <=( a879a ) or ( a880a );
 a3494a <=( a877a ) or ( a878a );
 a3495a <=( a3494a ) or ( a3491a );
 a3496a <=( a3495a ) or ( a3488a );
 a3497a <=( a3496a ) or ( a3483a );
 a3498a <=( a3497a ) or ( a3470a );
 a3499a <=( a3498a ) or ( a3443a );
 a3500a <=( a3499a ) or ( a3390a );
 a3501a <=( a3500a ) or ( a3281a );
 a3502a <=( a3501a ) or ( a3064a );
 a3503a <=( a3502a ) or ( a2627a );
 a3507a <=( a874a ) or ( a875a );
 a3508a <=( a876a ) or ( a3507a );
 a3512a <=( a871a ) or ( a872a );
 a3513a <=( a873a ) or ( a3512a );
 a3514a <=( a3513a ) or ( a3508a );
 a3518a <=( a868a ) or ( a869a );
 a3519a <=( a870a ) or ( a3518a );
 a3522a <=( a866a ) or ( a867a );
 a3525a <=( a864a ) or ( a865a );
 a3526a <=( a3525a ) or ( a3522a );
 a3527a <=( a3526a ) or ( a3519a );
 a3528a <=( a3527a ) or ( a3514a );
 a3532a <=( a861a ) or ( a862a );
 a3533a <=( a863a ) or ( a3532a );
 a3536a <=( a859a ) or ( a860a );
 a3539a <=( a857a ) or ( a858a );
 a3540a <=( a3539a ) or ( a3536a );
 a3541a <=( a3540a ) or ( a3533a );
 a3545a <=( a854a ) or ( a855a );
 a3546a <=( a856a ) or ( a3545a );
 a3549a <=( a852a ) or ( a853a );
 a3552a <=( a850a ) or ( a851a );
 a3553a <=( a3552a ) or ( a3549a );
 a3554a <=( a3553a ) or ( a3546a );
 a3555a <=( a3554a ) or ( a3541a );
 a3556a <=( a3555a ) or ( a3528a );
 a3560a <=( a847a ) or ( a848a );
 a3561a <=( a849a ) or ( a3560a );
 a3565a <=( a844a ) or ( a845a );
 a3566a <=( a846a ) or ( a3565a );
 a3567a <=( a3566a ) or ( a3561a );
 a3571a <=( a841a ) or ( a842a );
 a3572a <=( a843a ) or ( a3571a );
 a3575a <=( a839a ) or ( a840a );
 a3578a <=( a837a ) or ( a838a );
 a3579a <=( a3578a ) or ( a3575a );
 a3580a <=( a3579a ) or ( a3572a );
 a3581a <=( a3580a ) or ( a3567a );
 a3585a <=( a834a ) or ( a835a );
 a3586a <=( a836a ) or ( a3585a );
 a3589a <=( a832a ) or ( a833a );
 a3592a <=( a830a ) or ( a831a );
 a3593a <=( a3592a ) or ( a3589a );
 a3594a <=( a3593a ) or ( a3586a );
 a3598a <=( a827a ) or ( a828a );
 a3599a <=( a829a ) or ( a3598a );
 a3602a <=( a825a ) or ( a826a );
 a3605a <=( a823a ) or ( a824a );
 a3606a <=( a3605a ) or ( a3602a );
 a3607a <=( a3606a ) or ( a3599a );
 a3608a <=( a3607a ) or ( a3594a );
 a3609a <=( a3608a ) or ( a3581a );
 a3610a <=( a3609a ) or ( a3556a );
 a3614a <=( a820a ) or ( a821a );
 a3615a <=( a822a ) or ( a3614a );
 a3619a <=( a817a ) or ( a818a );
 a3620a <=( a819a ) or ( a3619a );
 a3621a <=( a3620a ) or ( a3615a );
 a3625a <=( a814a ) or ( a815a );
 a3626a <=( a816a ) or ( a3625a );
 a3629a <=( a812a ) or ( a813a );
 a3632a <=( a810a ) or ( a811a );
 a3633a <=( a3632a ) or ( a3629a );
 a3634a <=( a3633a ) or ( a3626a );
 a3635a <=( a3634a ) or ( a3621a );
 a3639a <=( a807a ) or ( a808a );
 a3640a <=( a809a ) or ( a3639a );
 a3643a <=( a805a ) or ( a806a );
 a3646a <=( a803a ) or ( a804a );
 a3647a <=( a3646a ) or ( a3643a );
 a3648a <=( a3647a ) or ( a3640a );
 a3652a <=( a800a ) or ( a801a );
 a3653a <=( a802a ) or ( a3652a );
 a3656a <=( a798a ) or ( a799a );
 a3659a <=( a796a ) or ( a797a );
 a3660a <=( a3659a ) or ( a3656a );
 a3661a <=( a3660a ) or ( a3653a );
 a3662a <=( a3661a ) or ( a3648a );
 a3663a <=( a3662a ) or ( a3635a );
 a3667a <=( a793a ) or ( a794a );
 a3668a <=( a795a ) or ( a3667a );
 a3671a <=( a791a ) or ( a792a );
 a3674a <=( a789a ) or ( a790a );
 a3675a <=( a3674a ) or ( a3671a );
 a3676a <=( a3675a ) or ( a3668a );
 a3680a <=( a786a ) or ( a787a );
 a3681a <=( a788a ) or ( a3680a );
 a3684a <=( a784a ) or ( a785a );
 a3687a <=( a782a ) or ( a783a );
 a3688a <=( a3687a ) or ( a3684a );
 a3689a <=( a3688a ) or ( a3681a );
 a3690a <=( a3689a ) or ( a3676a );
 a3694a <=( a779a ) or ( a780a );
 a3695a <=( a781a ) or ( a3694a );
 a3698a <=( a777a ) or ( a778a );
 a3701a <=( a775a ) or ( a776a );
 a3702a <=( a3701a ) or ( a3698a );
 a3703a <=( a3702a ) or ( a3695a );
 a3707a <=( a772a ) or ( a773a );
 a3708a <=( a774a ) or ( a3707a );
 a3711a <=( a770a ) or ( a771a );
 a3714a <=( a768a ) or ( a769a );
 a3715a <=( a3714a ) or ( a3711a );
 a3716a <=( a3715a ) or ( a3708a );
 a3717a <=( a3716a ) or ( a3703a );
 a3718a <=( a3717a ) or ( a3690a );
 a3719a <=( a3718a ) or ( a3663a );
 a3720a <=( a3719a ) or ( a3610a );
 a3724a <=( a765a ) or ( a766a );
 a3725a <=( a767a ) or ( a3724a );
 a3729a <=( a762a ) or ( a763a );
 a3730a <=( a764a ) or ( a3729a );
 a3731a <=( a3730a ) or ( a3725a );
 a3735a <=( a759a ) or ( a760a );
 a3736a <=( a761a ) or ( a3735a );
 a3739a <=( a757a ) or ( a758a );
 a3742a <=( a755a ) or ( a756a );
 a3743a <=( a3742a ) or ( a3739a );
 a3744a <=( a3743a ) or ( a3736a );
 a3745a <=( a3744a ) or ( a3731a );
 a3749a <=( a752a ) or ( a753a );
 a3750a <=( a754a ) or ( a3749a );
 a3753a <=( a750a ) or ( a751a );
 a3756a <=( a748a ) or ( a749a );
 a3757a <=( a3756a ) or ( a3753a );
 a3758a <=( a3757a ) or ( a3750a );
 a3762a <=( a745a ) or ( a746a );
 a3763a <=( a747a ) or ( a3762a );
 a3766a <=( a743a ) or ( a744a );
 a3769a <=( a741a ) or ( a742a );
 a3770a <=( a3769a ) or ( a3766a );
 a3771a <=( a3770a ) or ( a3763a );
 a3772a <=( a3771a ) or ( a3758a );
 a3773a <=( a3772a ) or ( a3745a );
 a3777a <=( a738a ) or ( a739a );
 a3778a <=( a740a ) or ( a3777a );
 a3781a <=( a736a ) or ( a737a );
 a3784a <=( a734a ) or ( a735a );
 a3785a <=( a3784a ) or ( a3781a );
 a3786a <=( a3785a ) or ( a3778a );
 a3790a <=( a731a ) or ( a732a );
 a3791a <=( a733a ) or ( a3790a );
 a3794a <=( a729a ) or ( a730a );
 a3797a <=( a727a ) or ( a728a );
 a3798a <=( a3797a ) or ( a3794a );
 a3799a <=( a3798a ) or ( a3791a );
 a3800a <=( a3799a ) or ( a3786a );
 a3804a <=( a724a ) or ( a725a );
 a3805a <=( a726a ) or ( a3804a );
 a3808a <=( a722a ) or ( a723a );
 a3811a <=( a720a ) or ( a721a );
 a3812a <=( a3811a ) or ( a3808a );
 a3813a <=( a3812a ) or ( a3805a );
 a3817a <=( a717a ) or ( a718a );
 a3818a <=( a719a ) or ( a3817a );
 a3821a <=( a715a ) or ( a716a );
 a3824a <=( a713a ) or ( a714a );
 a3825a <=( a3824a ) or ( a3821a );
 a3826a <=( a3825a ) or ( a3818a );
 a3827a <=( a3826a ) or ( a3813a );
 a3828a <=( a3827a ) or ( a3800a );
 a3829a <=( a3828a ) or ( a3773a );
 a3833a <=( a710a ) or ( a711a );
 a3834a <=( a712a ) or ( a3833a );
 a3838a <=( a707a ) or ( a708a );
 a3839a <=( a709a ) or ( a3838a );
 a3840a <=( a3839a ) or ( a3834a );
 a3844a <=( a704a ) or ( a705a );
 a3845a <=( a706a ) or ( a3844a );
 a3848a <=( a702a ) or ( a703a );
 a3851a <=( a700a ) or ( a701a );
 a3852a <=( a3851a ) or ( a3848a );
 a3853a <=( a3852a ) or ( a3845a );
 a3854a <=( a3853a ) or ( a3840a );
 a3858a <=( a697a ) or ( a698a );
 a3859a <=( a699a ) or ( a3858a );
 a3862a <=( a695a ) or ( a696a );
 a3865a <=( a693a ) or ( a694a );
 a3866a <=( a3865a ) or ( a3862a );
 a3867a <=( a3866a ) or ( a3859a );
 a3871a <=( a690a ) or ( a691a );
 a3872a <=( a692a ) or ( a3871a );
 a3875a <=( a688a ) or ( a689a );
 a3878a <=( a686a ) or ( a687a );
 a3879a <=( a3878a ) or ( a3875a );
 a3880a <=( a3879a ) or ( a3872a );
 a3881a <=( a3880a ) or ( a3867a );
 a3882a <=( a3881a ) or ( a3854a );
 a3886a <=( a683a ) or ( a684a );
 a3887a <=( a685a ) or ( a3886a );
 a3890a <=( a681a ) or ( a682a );
 a3893a <=( a679a ) or ( a680a );
 a3894a <=( a3893a ) or ( a3890a );
 a3895a <=( a3894a ) or ( a3887a );
 a3899a <=( a676a ) or ( a677a );
 a3900a <=( a678a ) or ( a3899a );
 a3903a <=( a674a ) or ( a675a );
 a3906a <=( a672a ) or ( a673a );
 a3907a <=( a3906a ) or ( a3903a );
 a3908a <=( a3907a ) or ( a3900a );
 a3909a <=( a3908a ) or ( a3895a );
 a3913a <=( a669a ) or ( a670a );
 a3914a <=( a671a ) or ( a3913a );
 a3917a <=( a667a ) or ( a668a );
 a3920a <=( a665a ) or ( a666a );
 a3921a <=( a3920a ) or ( a3917a );
 a3922a <=( a3921a ) or ( a3914a );
 a3926a <=( a662a ) or ( a663a );
 a3927a <=( a664a ) or ( a3926a );
 a3930a <=( a660a ) or ( a661a );
 a3933a <=( a658a ) or ( a659a );
 a3934a <=( a3933a ) or ( a3930a );
 a3935a <=( a3934a ) or ( a3927a );
 a3936a <=( a3935a ) or ( a3922a );
 a3937a <=( a3936a ) or ( a3909a );
 a3938a <=( a3937a ) or ( a3882a );
 a3939a <=( a3938a ) or ( a3829a );
 a3940a <=( a3939a ) or ( a3720a );
 a3944a <=( a655a ) or ( a656a );
 a3945a <=( a657a ) or ( a3944a );
 a3949a <=( a652a ) or ( a653a );
 a3950a <=( a654a ) or ( a3949a );
 a3951a <=( a3950a ) or ( a3945a );
 a3955a <=( a649a ) or ( a650a );
 a3956a <=( a651a ) or ( a3955a );
 a3959a <=( a647a ) or ( a648a );
 a3962a <=( a645a ) or ( a646a );
 a3963a <=( a3962a ) or ( a3959a );
 a3964a <=( a3963a ) or ( a3956a );
 a3965a <=( a3964a ) or ( a3951a );
 a3969a <=( a642a ) or ( a643a );
 a3970a <=( a644a ) or ( a3969a );
 a3973a <=( a640a ) or ( a641a );
 a3976a <=( a638a ) or ( a639a );
 a3977a <=( a3976a ) or ( a3973a );
 a3978a <=( a3977a ) or ( a3970a );
 a3982a <=( a635a ) or ( a636a );
 a3983a <=( a637a ) or ( a3982a );
 a3986a <=( a633a ) or ( a634a );
 a3989a <=( a631a ) or ( a632a );
 a3990a <=( a3989a ) or ( a3986a );
 a3991a <=( a3990a ) or ( a3983a );
 a3992a <=( a3991a ) or ( a3978a );
 a3993a <=( a3992a ) or ( a3965a );
 a3997a <=( a628a ) or ( a629a );
 a3998a <=( a630a ) or ( a3997a );
 a4002a <=( a625a ) or ( a626a );
 a4003a <=( a627a ) or ( a4002a );
 a4004a <=( a4003a ) or ( a3998a );
 a4008a <=( a622a ) or ( a623a );
 a4009a <=( a624a ) or ( a4008a );
 a4012a <=( a620a ) or ( a621a );
 a4015a <=( a618a ) or ( a619a );
 a4016a <=( a4015a ) or ( a4012a );
 a4017a <=( a4016a ) or ( a4009a );
 a4018a <=( a4017a ) or ( a4004a );
 a4022a <=( a615a ) or ( a616a );
 a4023a <=( a617a ) or ( a4022a );
 a4026a <=( a613a ) or ( a614a );
 a4029a <=( a611a ) or ( a612a );
 a4030a <=( a4029a ) or ( a4026a );
 a4031a <=( a4030a ) or ( a4023a );
 a4035a <=( a608a ) or ( a609a );
 a4036a <=( a610a ) or ( a4035a );
 a4039a <=( a606a ) or ( a607a );
 a4042a <=( a604a ) or ( a605a );
 a4043a <=( a4042a ) or ( a4039a );
 a4044a <=( a4043a ) or ( a4036a );
 a4045a <=( a4044a ) or ( a4031a );
 a4046a <=( a4045a ) or ( a4018a );
 a4047a <=( a4046a ) or ( a3993a );
 a4051a <=( a601a ) or ( a602a );
 a4052a <=( a603a ) or ( a4051a );
 a4056a <=( a598a ) or ( a599a );
 a4057a <=( a600a ) or ( a4056a );
 a4058a <=( a4057a ) or ( a4052a );
 a4062a <=( a595a ) or ( a596a );
 a4063a <=( a597a ) or ( a4062a );
 a4066a <=( a593a ) or ( a594a );
 a4069a <=( a591a ) or ( a592a );
 a4070a <=( a4069a ) or ( a4066a );
 a4071a <=( a4070a ) or ( a4063a );
 a4072a <=( a4071a ) or ( a4058a );
 a4076a <=( a588a ) or ( a589a );
 a4077a <=( a590a ) or ( a4076a );
 a4080a <=( a586a ) or ( a587a );
 a4083a <=( a584a ) or ( a585a );
 a4084a <=( a4083a ) or ( a4080a );
 a4085a <=( a4084a ) or ( a4077a );
 a4089a <=( a581a ) or ( a582a );
 a4090a <=( a583a ) or ( a4089a );
 a4093a <=( a579a ) or ( a580a );
 a4096a <=( a577a ) or ( a578a );
 a4097a <=( a4096a ) or ( a4093a );
 a4098a <=( a4097a ) or ( a4090a );
 a4099a <=( a4098a ) or ( a4085a );
 a4100a <=( a4099a ) or ( a4072a );
 a4104a <=( a574a ) or ( a575a );
 a4105a <=( a576a ) or ( a4104a );
 a4108a <=( a572a ) or ( a573a );
 a4111a <=( a570a ) or ( a571a );
 a4112a <=( a4111a ) or ( a4108a );
 a4113a <=( a4112a ) or ( a4105a );
 a4117a <=( a567a ) or ( a568a );
 a4118a <=( a569a ) or ( a4117a );
 a4121a <=( a565a ) or ( a566a );
 a4124a <=( a563a ) or ( a564a );
 a4125a <=( a4124a ) or ( a4121a );
 a4126a <=( a4125a ) or ( a4118a );
 a4127a <=( a4126a ) or ( a4113a );
 a4131a <=( a560a ) or ( a561a );
 a4132a <=( a562a ) or ( a4131a );
 a4135a <=( a558a ) or ( a559a );
 a4138a <=( a556a ) or ( a557a );
 a4139a <=( a4138a ) or ( a4135a );
 a4140a <=( a4139a ) or ( a4132a );
 a4144a <=( a553a ) or ( a554a );
 a4145a <=( a555a ) or ( a4144a );
 a4148a <=( a551a ) or ( a552a );
 a4151a <=( a549a ) or ( a550a );
 a4152a <=( a4151a ) or ( a4148a );
 a4153a <=( a4152a ) or ( a4145a );
 a4154a <=( a4153a ) or ( a4140a );
 a4155a <=( a4154a ) or ( a4127a );
 a4156a <=( a4155a ) or ( a4100a );
 a4157a <=( a4156a ) or ( a4047a );
 a4161a <=( a546a ) or ( a547a );
 a4162a <=( a548a ) or ( a4161a );
 a4166a <=( a543a ) or ( a544a );
 a4167a <=( a545a ) or ( a4166a );
 a4168a <=( a4167a ) or ( a4162a );
 a4172a <=( a540a ) or ( a541a );
 a4173a <=( a542a ) or ( a4172a );
 a4176a <=( a538a ) or ( a539a );
 a4179a <=( a536a ) or ( a537a );
 a4180a <=( a4179a ) or ( a4176a );
 a4181a <=( a4180a ) or ( a4173a );
 a4182a <=( a4181a ) or ( a4168a );
 a4186a <=( a533a ) or ( a534a );
 a4187a <=( a535a ) or ( a4186a );
 a4190a <=( a531a ) or ( a532a );
 a4193a <=( a529a ) or ( a530a );
 a4194a <=( a4193a ) or ( a4190a );
 a4195a <=( a4194a ) or ( a4187a );
 a4199a <=( a526a ) or ( a527a );
 a4200a <=( a528a ) or ( a4199a );
 a4203a <=( a524a ) or ( a525a );
 a4206a <=( a522a ) or ( a523a );
 a4207a <=( a4206a ) or ( a4203a );
 a4208a <=( a4207a ) or ( a4200a );
 a4209a <=( a4208a ) or ( a4195a );
 a4210a <=( a4209a ) or ( a4182a );
 a4214a <=( a519a ) or ( a520a );
 a4215a <=( a521a ) or ( a4214a );
 a4218a <=( a517a ) or ( a518a );
 a4221a <=( a515a ) or ( a516a );
 a4222a <=( a4221a ) or ( a4218a );
 a4223a <=( a4222a ) or ( a4215a );
 a4227a <=( a512a ) or ( a513a );
 a4228a <=( a514a ) or ( a4227a );
 a4231a <=( a510a ) or ( a511a );
 a4234a <=( a508a ) or ( a509a );
 a4235a <=( a4234a ) or ( a4231a );
 a4236a <=( a4235a ) or ( a4228a );
 a4237a <=( a4236a ) or ( a4223a );
 a4241a <=( a505a ) or ( a506a );
 a4242a <=( a507a ) or ( a4241a );
 a4245a <=( a503a ) or ( a504a );
 a4248a <=( a501a ) or ( a502a );
 a4249a <=( a4248a ) or ( a4245a );
 a4250a <=( a4249a ) or ( a4242a );
 a4254a <=( a498a ) or ( a499a );
 a4255a <=( a500a ) or ( a4254a );
 a4258a <=( a496a ) or ( a497a );
 a4261a <=( a494a ) or ( a495a );
 a4262a <=( a4261a ) or ( a4258a );
 a4263a <=( a4262a ) or ( a4255a );
 a4264a <=( a4263a ) or ( a4250a );
 a4265a <=( a4264a ) or ( a4237a );
 a4266a <=( a4265a ) or ( a4210a );
 a4270a <=( a491a ) or ( a492a );
 a4271a <=( a493a ) or ( a4270a );
 a4275a <=( a488a ) or ( a489a );
 a4276a <=( a490a ) or ( a4275a );
 a4277a <=( a4276a ) or ( a4271a );
 a4281a <=( a485a ) or ( a486a );
 a4282a <=( a487a ) or ( a4281a );
 a4285a <=( a483a ) or ( a484a );
 a4288a <=( a481a ) or ( a482a );
 a4289a <=( a4288a ) or ( a4285a );
 a4290a <=( a4289a ) or ( a4282a );
 a4291a <=( a4290a ) or ( a4277a );
 a4295a <=( a478a ) or ( a479a );
 a4296a <=( a480a ) or ( a4295a );
 a4299a <=( a476a ) or ( a477a );
 a4302a <=( a474a ) or ( a475a );
 a4303a <=( a4302a ) or ( a4299a );
 a4304a <=( a4303a ) or ( a4296a );
 a4308a <=( a471a ) or ( a472a );
 a4309a <=( a473a ) or ( a4308a );
 a4312a <=( a469a ) or ( a470a );
 a4315a <=( a467a ) or ( a468a );
 a4316a <=( a4315a ) or ( a4312a );
 a4317a <=( a4316a ) or ( a4309a );
 a4318a <=( a4317a ) or ( a4304a );
 a4319a <=( a4318a ) or ( a4291a );
 a4323a <=( a464a ) or ( a465a );
 a4324a <=( a466a ) or ( a4323a );
 a4327a <=( a462a ) or ( a463a );
 a4330a <=( a460a ) or ( a461a );
 a4331a <=( a4330a ) or ( a4327a );
 a4332a <=( a4331a ) or ( a4324a );
 a4336a <=( a457a ) or ( a458a );
 a4337a <=( a459a ) or ( a4336a );
 a4340a <=( a455a ) or ( a456a );
 a4343a <=( a453a ) or ( a454a );
 a4344a <=( a4343a ) or ( a4340a );
 a4345a <=( a4344a ) or ( a4337a );
 a4346a <=( a4345a ) or ( a4332a );
 a4350a <=( a450a ) or ( a451a );
 a4351a <=( a452a ) or ( a4350a );
 a4354a <=( a448a ) or ( a449a );
 a4357a <=( a446a ) or ( a447a );
 a4358a <=( a4357a ) or ( a4354a );
 a4359a <=( a4358a ) or ( a4351a );
 a4363a <=( a443a ) or ( a444a );
 a4364a <=( a445a ) or ( a4363a );
 a4367a <=( a441a ) or ( a442a );
 a4370a <=( a439a ) or ( a440a );
 a4371a <=( a4370a ) or ( a4367a );
 a4372a <=( a4371a ) or ( a4364a );
 a4373a <=( a4372a ) or ( a4359a );
 a4374a <=( a4373a ) or ( a4346a );
 a4375a <=( a4374a ) or ( a4319a );
 a4376a <=( a4375a ) or ( a4266a );
 a4377a <=( a4376a ) or ( a4157a );
 a4378a <=( a4377a ) or ( a3940a );
 a4382a <=( a436a ) or ( a437a );
 a4383a <=( a438a ) or ( a4382a );
 a4387a <=( a433a ) or ( a434a );
 a4388a <=( a435a ) or ( a4387a );
 a4389a <=( a4388a ) or ( a4383a );
 a4393a <=( a430a ) or ( a431a );
 a4394a <=( a432a ) or ( a4393a );
 a4397a <=( a428a ) or ( a429a );
 a4400a <=( a426a ) or ( a427a );
 a4401a <=( a4400a ) or ( a4397a );
 a4402a <=( a4401a ) or ( a4394a );
 a4403a <=( a4402a ) or ( a4389a );
 a4407a <=( a423a ) or ( a424a );
 a4408a <=( a425a ) or ( a4407a );
 a4411a <=( a421a ) or ( a422a );
 a4414a <=( a419a ) or ( a420a );
 a4415a <=( a4414a ) or ( a4411a );
 a4416a <=( a4415a ) or ( a4408a );
 a4420a <=( a416a ) or ( a417a );
 a4421a <=( a418a ) or ( a4420a );
 a4424a <=( a414a ) or ( a415a );
 a4427a <=( a412a ) or ( a413a );
 a4428a <=( a4427a ) or ( a4424a );
 a4429a <=( a4428a ) or ( a4421a );
 a4430a <=( a4429a ) or ( a4416a );
 a4431a <=( a4430a ) or ( a4403a );
 a4435a <=( a409a ) or ( a410a );
 a4436a <=( a411a ) or ( a4435a );
 a4440a <=( a406a ) or ( a407a );
 a4441a <=( a408a ) or ( a4440a );
 a4442a <=( a4441a ) or ( a4436a );
 a4446a <=( a403a ) or ( a404a );
 a4447a <=( a405a ) or ( a4446a );
 a4450a <=( a401a ) or ( a402a );
 a4453a <=( a399a ) or ( a400a );
 a4454a <=( a4453a ) or ( a4450a );
 a4455a <=( a4454a ) or ( a4447a );
 a4456a <=( a4455a ) or ( a4442a );
 a4460a <=( a396a ) or ( a397a );
 a4461a <=( a398a ) or ( a4460a );
 a4464a <=( a394a ) or ( a395a );
 a4467a <=( a392a ) or ( a393a );
 a4468a <=( a4467a ) or ( a4464a );
 a4469a <=( a4468a ) or ( a4461a );
 a4473a <=( a389a ) or ( a390a );
 a4474a <=( a391a ) or ( a4473a );
 a4477a <=( a387a ) or ( a388a );
 a4480a <=( a385a ) or ( a386a );
 a4481a <=( a4480a ) or ( a4477a );
 a4482a <=( a4481a ) or ( a4474a );
 a4483a <=( a4482a ) or ( a4469a );
 a4484a <=( a4483a ) or ( a4456a );
 a4485a <=( a4484a ) or ( a4431a );
 a4489a <=( a382a ) or ( a383a );
 a4490a <=( a384a ) or ( a4489a );
 a4494a <=( a379a ) or ( a380a );
 a4495a <=( a381a ) or ( a4494a );
 a4496a <=( a4495a ) or ( a4490a );
 a4500a <=( a376a ) or ( a377a );
 a4501a <=( a378a ) or ( a4500a );
 a4504a <=( a374a ) or ( a375a );
 a4507a <=( a372a ) or ( a373a );
 a4508a <=( a4507a ) or ( a4504a );
 a4509a <=( a4508a ) or ( a4501a );
 a4510a <=( a4509a ) or ( a4496a );
 a4514a <=( a369a ) or ( a370a );
 a4515a <=( a371a ) or ( a4514a );
 a4518a <=( a367a ) or ( a368a );
 a4521a <=( a365a ) or ( a366a );
 a4522a <=( a4521a ) or ( a4518a );
 a4523a <=( a4522a ) or ( a4515a );
 a4527a <=( a362a ) or ( a363a );
 a4528a <=( a364a ) or ( a4527a );
 a4531a <=( a360a ) or ( a361a );
 a4534a <=( a358a ) or ( a359a );
 a4535a <=( a4534a ) or ( a4531a );
 a4536a <=( a4535a ) or ( a4528a );
 a4537a <=( a4536a ) or ( a4523a );
 a4538a <=( a4537a ) or ( a4510a );
 a4542a <=( a355a ) or ( a356a );
 a4543a <=( a357a ) or ( a4542a );
 a4546a <=( a353a ) or ( a354a );
 a4549a <=( a351a ) or ( a352a );
 a4550a <=( a4549a ) or ( a4546a );
 a4551a <=( a4550a ) or ( a4543a );
 a4555a <=( a348a ) or ( a349a );
 a4556a <=( a350a ) or ( a4555a );
 a4559a <=( a346a ) or ( a347a );
 a4562a <=( a344a ) or ( a345a );
 a4563a <=( a4562a ) or ( a4559a );
 a4564a <=( a4563a ) or ( a4556a );
 a4565a <=( a4564a ) or ( a4551a );
 a4569a <=( a341a ) or ( a342a );
 a4570a <=( a343a ) or ( a4569a );
 a4573a <=( a339a ) or ( a340a );
 a4576a <=( a337a ) or ( a338a );
 a4577a <=( a4576a ) or ( a4573a );
 a4578a <=( a4577a ) or ( a4570a );
 a4582a <=( a334a ) or ( a335a );
 a4583a <=( a336a ) or ( a4582a );
 a4586a <=( a332a ) or ( a333a );
 a4589a <=( a330a ) or ( a331a );
 a4590a <=( a4589a ) or ( a4586a );
 a4591a <=( a4590a ) or ( a4583a );
 a4592a <=( a4591a ) or ( a4578a );
 a4593a <=( a4592a ) or ( a4565a );
 a4594a <=( a4593a ) or ( a4538a );
 a4595a <=( a4594a ) or ( a4485a );
 a4599a <=( a327a ) or ( a328a );
 a4600a <=( a329a ) or ( a4599a );
 a4604a <=( a324a ) or ( a325a );
 a4605a <=( a326a ) or ( a4604a );
 a4606a <=( a4605a ) or ( a4600a );
 a4610a <=( a321a ) or ( a322a );
 a4611a <=( a323a ) or ( a4610a );
 a4614a <=( a319a ) or ( a320a );
 a4617a <=( a317a ) or ( a318a );
 a4618a <=( a4617a ) or ( a4614a );
 a4619a <=( a4618a ) or ( a4611a );
 a4620a <=( a4619a ) or ( a4606a );
 a4624a <=( a314a ) or ( a315a );
 a4625a <=( a316a ) or ( a4624a );
 a4628a <=( a312a ) or ( a313a );
 a4631a <=( a310a ) or ( a311a );
 a4632a <=( a4631a ) or ( a4628a );
 a4633a <=( a4632a ) or ( a4625a );
 a4637a <=( a307a ) or ( a308a );
 a4638a <=( a309a ) or ( a4637a );
 a4641a <=( a305a ) or ( a306a );
 a4644a <=( a303a ) or ( a304a );
 a4645a <=( a4644a ) or ( a4641a );
 a4646a <=( a4645a ) or ( a4638a );
 a4647a <=( a4646a ) or ( a4633a );
 a4648a <=( a4647a ) or ( a4620a );
 a4652a <=( a300a ) or ( a301a );
 a4653a <=( a302a ) or ( a4652a );
 a4656a <=( a298a ) or ( a299a );
 a4659a <=( a296a ) or ( a297a );
 a4660a <=( a4659a ) or ( a4656a );
 a4661a <=( a4660a ) or ( a4653a );
 a4665a <=( a293a ) or ( a294a );
 a4666a <=( a295a ) or ( a4665a );
 a4669a <=( a291a ) or ( a292a );
 a4672a <=( a289a ) or ( a290a );
 a4673a <=( a4672a ) or ( a4669a );
 a4674a <=( a4673a ) or ( a4666a );
 a4675a <=( a4674a ) or ( a4661a );
 a4679a <=( a286a ) or ( a287a );
 a4680a <=( a288a ) or ( a4679a );
 a4683a <=( a284a ) or ( a285a );
 a4686a <=( a282a ) or ( a283a );
 a4687a <=( a4686a ) or ( a4683a );
 a4688a <=( a4687a ) or ( a4680a );
 a4692a <=( a279a ) or ( a280a );
 a4693a <=( a281a ) or ( a4692a );
 a4696a <=( a277a ) or ( a278a );
 a4699a <=( a275a ) or ( a276a );
 a4700a <=( a4699a ) or ( a4696a );
 a4701a <=( a4700a ) or ( a4693a );
 a4702a <=( a4701a ) or ( a4688a );
 a4703a <=( a4702a ) or ( a4675a );
 a4704a <=( a4703a ) or ( a4648a );
 a4708a <=( a272a ) or ( a273a );
 a4709a <=( a274a ) or ( a4708a );
 a4713a <=( a269a ) or ( a270a );
 a4714a <=( a271a ) or ( a4713a );
 a4715a <=( a4714a ) or ( a4709a );
 a4719a <=( a266a ) or ( a267a );
 a4720a <=( a268a ) or ( a4719a );
 a4723a <=( a264a ) or ( a265a );
 a4726a <=( a262a ) or ( a263a );
 a4727a <=( a4726a ) or ( a4723a );
 a4728a <=( a4727a ) or ( a4720a );
 a4729a <=( a4728a ) or ( a4715a );
 a4733a <=( a259a ) or ( a260a );
 a4734a <=( a261a ) or ( a4733a );
 a4737a <=( a257a ) or ( a258a );
 a4740a <=( a255a ) or ( a256a );
 a4741a <=( a4740a ) or ( a4737a );
 a4742a <=( a4741a ) or ( a4734a );
 a4746a <=( a252a ) or ( a253a );
 a4747a <=( a254a ) or ( a4746a );
 a4750a <=( a250a ) or ( a251a );
 a4753a <=( a248a ) or ( a249a );
 a4754a <=( a4753a ) or ( a4750a );
 a4755a <=( a4754a ) or ( a4747a );
 a4756a <=( a4755a ) or ( a4742a );
 a4757a <=( a4756a ) or ( a4729a );
 a4761a <=( a245a ) or ( a246a );
 a4762a <=( a247a ) or ( a4761a );
 a4765a <=( a243a ) or ( a244a );
 a4768a <=( a241a ) or ( a242a );
 a4769a <=( a4768a ) or ( a4765a );
 a4770a <=( a4769a ) or ( a4762a );
 a4774a <=( a238a ) or ( a239a );
 a4775a <=( a240a ) or ( a4774a );
 a4778a <=( a236a ) or ( a237a );
 a4781a <=( a234a ) or ( a235a );
 a4782a <=( a4781a ) or ( a4778a );
 a4783a <=( a4782a ) or ( a4775a );
 a4784a <=( a4783a ) or ( a4770a );
 a4788a <=( a231a ) or ( a232a );
 a4789a <=( a233a ) or ( a4788a );
 a4792a <=( a229a ) or ( a230a );
 a4795a <=( a227a ) or ( a228a );
 a4796a <=( a4795a ) or ( a4792a );
 a4797a <=( a4796a ) or ( a4789a );
 a4801a <=( a224a ) or ( a225a );
 a4802a <=( a226a ) or ( a4801a );
 a4805a <=( a222a ) or ( a223a );
 a4808a <=( a220a ) or ( a221a );
 a4809a <=( a4808a ) or ( a4805a );
 a4810a <=( a4809a ) or ( a4802a );
 a4811a <=( a4810a ) or ( a4797a );
 a4812a <=( a4811a ) or ( a4784a );
 a4813a <=( a4812a ) or ( a4757a );
 a4814a <=( a4813a ) or ( a4704a );
 a4815a <=( a4814a ) or ( a4595a );
 a4819a <=( a217a ) or ( a218a );
 a4820a <=( a219a ) or ( a4819a );
 a4824a <=( a214a ) or ( a215a );
 a4825a <=( a216a ) or ( a4824a );
 a4826a <=( a4825a ) or ( a4820a );
 a4830a <=( a211a ) or ( a212a );
 a4831a <=( a213a ) or ( a4830a );
 a4834a <=( a209a ) or ( a210a );
 a4837a <=( a207a ) or ( a208a );
 a4838a <=( a4837a ) or ( a4834a );
 a4839a <=( a4838a ) or ( a4831a );
 a4840a <=( a4839a ) or ( a4826a );
 a4844a <=( a204a ) or ( a205a );
 a4845a <=( a206a ) or ( a4844a );
 a4848a <=( a202a ) or ( a203a );
 a4851a <=( a200a ) or ( a201a );
 a4852a <=( a4851a ) or ( a4848a );
 a4853a <=( a4852a ) or ( a4845a );
 a4857a <=( a197a ) or ( a198a );
 a4858a <=( a199a ) or ( a4857a );
 a4861a <=( a195a ) or ( a196a );
 a4864a <=( a193a ) or ( a194a );
 a4865a <=( a4864a ) or ( a4861a );
 a4866a <=( a4865a ) or ( a4858a );
 a4867a <=( a4866a ) or ( a4853a );
 a4868a <=( a4867a ) or ( a4840a );
 a4872a <=( a190a ) or ( a191a );
 a4873a <=( a192a ) or ( a4872a );
 a4877a <=( a187a ) or ( a188a );
 a4878a <=( a189a ) or ( a4877a );
 a4879a <=( a4878a ) or ( a4873a );
 a4883a <=( a184a ) or ( a185a );
 a4884a <=( a186a ) or ( a4883a );
 a4887a <=( a182a ) or ( a183a );
 a4890a <=( a180a ) or ( a181a );
 a4891a <=( a4890a ) or ( a4887a );
 a4892a <=( a4891a ) or ( a4884a );
 a4893a <=( a4892a ) or ( a4879a );
 a4897a <=( a177a ) or ( a178a );
 a4898a <=( a179a ) or ( a4897a );
 a4901a <=( a175a ) or ( a176a );
 a4904a <=( a173a ) or ( a174a );
 a4905a <=( a4904a ) or ( a4901a );
 a4906a <=( a4905a ) or ( a4898a );
 a4910a <=( a170a ) or ( a171a );
 a4911a <=( a172a ) or ( a4910a );
 a4914a <=( a168a ) or ( a169a );
 a4917a <=( a166a ) or ( a167a );
 a4918a <=( a4917a ) or ( a4914a );
 a4919a <=( a4918a ) or ( a4911a );
 a4920a <=( a4919a ) or ( a4906a );
 a4921a <=( a4920a ) or ( a4893a );
 a4922a <=( a4921a ) or ( a4868a );
 a4926a <=( a163a ) or ( a164a );
 a4927a <=( a165a ) or ( a4926a );
 a4931a <=( a160a ) or ( a161a );
 a4932a <=( a162a ) or ( a4931a );
 a4933a <=( a4932a ) or ( a4927a );
 a4937a <=( a157a ) or ( a158a );
 a4938a <=( a159a ) or ( a4937a );
 a4941a <=( a155a ) or ( a156a );
 a4944a <=( a153a ) or ( a154a );
 a4945a <=( a4944a ) or ( a4941a );
 a4946a <=( a4945a ) or ( a4938a );
 a4947a <=( a4946a ) or ( a4933a );
 a4951a <=( a150a ) or ( a151a );
 a4952a <=( a152a ) or ( a4951a );
 a4955a <=( a148a ) or ( a149a );
 a4958a <=( a146a ) or ( a147a );
 a4959a <=( a4958a ) or ( a4955a );
 a4960a <=( a4959a ) or ( a4952a );
 a4964a <=( a143a ) or ( a144a );
 a4965a <=( a145a ) or ( a4964a );
 a4968a <=( a141a ) or ( a142a );
 a4971a <=( a139a ) or ( a140a );
 a4972a <=( a4971a ) or ( a4968a );
 a4973a <=( a4972a ) or ( a4965a );
 a4974a <=( a4973a ) or ( a4960a );
 a4975a <=( a4974a ) or ( a4947a );
 a4979a <=( a136a ) or ( a137a );
 a4980a <=( a138a ) or ( a4979a );
 a4983a <=( a134a ) or ( a135a );
 a4986a <=( a132a ) or ( a133a );
 a4987a <=( a4986a ) or ( a4983a );
 a4988a <=( a4987a ) or ( a4980a );
 a4992a <=( a129a ) or ( a130a );
 a4993a <=( a131a ) or ( a4992a );
 a4996a <=( a127a ) or ( a128a );
 a4999a <=( a125a ) or ( a126a );
 a5000a <=( a4999a ) or ( a4996a );
 a5001a <=( a5000a ) or ( a4993a );
 a5002a <=( a5001a ) or ( a4988a );
 a5006a <=( a122a ) or ( a123a );
 a5007a <=( a124a ) or ( a5006a );
 a5010a <=( a120a ) or ( a121a );
 a5013a <=( a118a ) or ( a119a );
 a5014a <=( a5013a ) or ( a5010a );
 a5015a <=( a5014a ) or ( a5007a );
 a5019a <=( a115a ) or ( a116a );
 a5020a <=( a117a ) or ( a5019a );
 a5023a <=( a113a ) or ( a114a );
 a5026a <=( a111a ) or ( a112a );
 a5027a <=( a5026a ) or ( a5023a );
 a5028a <=( a5027a ) or ( a5020a );
 a5029a <=( a5028a ) or ( a5015a );
 a5030a <=( a5029a ) or ( a5002a );
 a5031a <=( a5030a ) or ( a4975a );
 a5032a <=( a5031a ) or ( a4922a );
 a5036a <=( a108a ) or ( a109a );
 a5037a <=( a110a ) or ( a5036a );
 a5041a <=( a105a ) or ( a106a );
 a5042a <=( a107a ) or ( a5041a );
 a5043a <=( a5042a ) or ( a5037a );
 a5047a <=( a102a ) or ( a103a );
 a5048a <=( a104a ) or ( a5047a );
 a5051a <=( a100a ) or ( a101a );
 a5054a <=( a98a ) or ( a99a );
 a5055a <=( a5054a ) or ( a5051a );
 a5056a <=( a5055a ) or ( a5048a );
 a5057a <=( a5056a ) or ( a5043a );
 a5061a <=( a95a ) or ( a96a );
 a5062a <=( a97a ) or ( a5061a );
 a5065a <=( a93a ) or ( a94a );
 a5068a <=( a91a ) or ( a92a );
 a5069a <=( a5068a ) or ( a5065a );
 a5070a <=( a5069a ) or ( a5062a );
 a5074a <=( a88a ) or ( a89a );
 a5075a <=( a90a ) or ( a5074a );
 a5078a <=( a86a ) or ( a87a );
 a5081a <=( a84a ) or ( a85a );
 a5082a <=( a5081a ) or ( a5078a );
 a5083a <=( a5082a ) or ( a5075a );
 a5084a <=( a5083a ) or ( a5070a );
 a5085a <=( a5084a ) or ( a5057a );
 a5089a <=( a81a ) or ( a82a );
 a5090a <=( a83a ) or ( a5089a );
 a5093a <=( a79a ) or ( a80a );
 a5096a <=( a77a ) or ( a78a );
 a5097a <=( a5096a ) or ( a5093a );
 a5098a <=( a5097a ) or ( a5090a );
 a5102a <=( a74a ) or ( a75a );
 a5103a <=( a76a ) or ( a5102a );
 a5106a <=( a72a ) or ( a73a );
 a5109a <=( a70a ) or ( a71a );
 a5110a <=( a5109a ) or ( a5106a );
 a5111a <=( a5110a ) or ( a5103a );
 a5112a <=( a5111a ) or ( a5098a );
 a5116a <=( a67a ) or ( a68a );
 a5117a <=( a69a ) or ( a5116a );
 a5120a <=( a65a ) or ( a66a );
 a5123a <=( a63a ) or ( a64a );
 a5124a <=( a5123a ) or ( a5120a );
 a5125a <=( a5124a ) or ( a5117a );
 a5129a <=( a60a ) or ( a61a );
 a5130a <=( a62a ) or ( a5129a );
 a5133a <=( a58a ) or ( a59a );
 a5136a <=( a56a ) or ( a57a );
 a5137a <=( a5136a ) or ( a5133a );
 a5138a <=( a5137a ) or ( a5130a );
 a5139a <=( a5138a ) or ( a5125a );
 a5140a <=( a5139a ) or ( a5112a );
 a5141a <=( a5140a ) or ( a5085a );
 a5145a <=( a53a ) or ( a54a );
 a5146a <=( a55a ) or ( a5145a );
 a5150a <=( a50a ) or ( a51a );
 a5151a <=( a52a ) or ( a5150a );
 a5152a <=( a5151a ) or ( a5146a );
 a5156a <=( a47a ) or ( a48a );
 a5157a <=( a49a ) or ( a5156a );
 a5160a <=( a45a ) or ( a46a );
 a5163a <=( a43a ) or ( a44a );
 a5164a <=( a5163a ) or ( a5160a );
 a5165a <=( a5164a ) or ( a5157a );
 a5166a <=( a5165a ) or ( a5152a );
 a5170a <=( a40a ) or ( a41a );
 a5171a <=( a42a ) or ( a5170a );
 a5174a <=( a38a ) or ( a39a );
 a5177a <=( a36a ) or ( a37a );
 a5178a <=( a5177a ) or ( a5174a );
 a5179a <=( a5178a ) or ( a5171a );
 a5183a <=( a33a ) or ( a34a );
 a5184a <=( a35a ) or ( a5183a );
 a5187a <=( a31a ) or ( a32a );
 a5190a <=( a29a ) or ( a30a );
 a5191a <=( a5190a ) or ( a5187a );
 a5192a <=( a5191a ) or ( a5184a );
 a5193a <=( a5192a ) or ( a5179a );
 a5194a <=( a5193a ) or ( a5166a );
 a5198a <=( a26a ) or ( a27a );
 a5199a <=( a28a ) or ( a5198a );
 a5202a <=( a24a ) or ( a25a );
 a5205a <=( a22a ) or ( a23a );
 a5206a <=( a5205a ) or ( a5202a );
 a5207a <=( a5206a ) or ( a5199a );
 a5211a <=( a19a ) or ( a20a );
 a5212a <=( a21a ) or ( a5211a );
 a5215a <=( a17a ) or ( a18a );
 a5218a <=( a15a ) or ( a16a );
 a5219a <=( a5218a ) or ( a5215a );
 a5220a <=( a5219a ) or ( a5212a );
 a5221a <=( a5220a ) or ( a5207a );
 a5225a <=( a12a ) or ( a13a );
 a5226a <=( a14a ) or ( a5225a );
 a5229a <=( a10a ) or ( a11a );
 a5232a <=( a8a ) or ( a9a );
 a5233a <=( a5232a ) or ( a5229a );
 a5234a <=( a5233a ) or ( a5226a );
 a5238a <=( a5a ) or ( a6a );
 a5239a <=( a7a ) or ( a5238a );
 a5242a <=( a3a ) or ( a4a );
 a5245a <=( a1a ) or ( a2a );
 a5246a <=( a5245a ) or ( a5242a );
 a5247a <=( a5246a ) or ( a5239a );
 a5248a <=( a5247a ) or ( a5234a );
 a5249a <=( a5248a ) or ( a5221a );
 a5250a <=( a5249a ) or ( a5194a );
 a5251a <=( a5250a ) or ( a5141a );
 a5252a <=( a5251a ) or ( a5032a );
 a5253a <=( a5252a ) or ( a4815a );
 a5254a <=( a5253a ) or ( a4378a );
 a5257a <=( A166  and  A167 );
 a5260a <=( A201  and  A199 );
 a5263a <=( A166  and  A167 );
 a5266a <=( A201  and  A200 );
 a5269a <=( (not A166)  and  (not A167) );
 a5272a <=( A201  and  A199 );
 a5275a <=( (not A166)  and  (not A167) );
 a5278a <=( A201  and  A200 );
 a5281a <=( (not A167)  and  (not A168) );
 a5284a <=( A201  and  A199 );
 a5287a <=( (not A167)  and  (not A168) );
 a5290a <=( A201  and  A200 );
 a5293a <=( (not A169)  and  (not A170) );
 a5297a <=( A201  and  A199 );
 a5298a <=( (not A167)  and  a5297a );
 a5301a <=( (not A169)  and  (not A170) );
 a5305a <=( A201  and  A200 );
 a5306a <=( (not A167)  and  a5305a );
 a5310a <=( A199  and  A166 );
 a5311a <=( A167  and  a5310a );
 a5315a <=( (not A203)  and  A202 );
 a5316a <=( A200  and  a5315a );
 a5320a <=( (not A199)  and  A166 );
 a5321a <=( A167  and  a5320a );
 a5325a <=( A203  and  (not A202) );
 a5326a <=( A200  and  a5325a );
 a5330a <=( A199  and  A166 );
 a5331a <=( A167  and  a5330a );
 a5335a <=( A203  and  (not A202) );
 a5336a <=( (not A200)  and  a5335a );
 a5340a <=( (not A199)  and  A166 );
 a5341a <=( A167  and  a5340a );
 a5345a <=( (not A203)  and  A202 );
 a5346a <=( (not A200)  and  a5345a );
 a5350a <=( A199  and  (not A166) );
 a5351a <=( (not A167)  and  a5350a );
 a5355a <=( (not A203)  and  A202 );
 a5356a <=( A200  and  a5355a );
 a5360a <=( (not A199)  and  (not A166) );
 a5361a <=( (not A167)  and  a5360a );
 a5365a <=( A203  and  (not A202) );
 a5366a <=( A200  and  a5365a );
 a5370a <=( A199  and  (not A166) );
 a5371a <=( (not A167)  and  a5370a );
 a5375a <=( A203  and  (not A202) );
 a5376a <=( (not A200)  and  a5375a );
 a5380a <=( (not A199)  and  (not A166) );
 a5381a <=( (not A167)  and  a5380a );
 a5385a <=( (not A203)  and  A202 );
 a5386a <=( (not A200)  and  a5385a );
 a5390a <=( A199  and  (not A167) );
 a5391a <=( (not A168)  and  a5390a );
 a5395a <=( (not A203)  and  A202 );
 a5396a <=( A200  and  a5395a );
 a5400a <=( (not A199)  and  (not A167) );
 a5401a <=( (not A168)  and  a5400a );
 a5405a <=( A203  and  (not A202) );
 a5406a <=( A200  and  a5405a );
 a5410a <=( A199  and  (not A167) );
 a5411a <=( (not A168)  and  a5410a );
 a5415a <=( A203  and  (not A202) );
 a5416a <=( (not A200)  and  a5415a );
 a5420a <=( (not A199)  and  (not A167) );
 a5421a <=( (not A168)  and  a5420a );
 a5425a <=( (not A203)  and  A202 );
 a5426a <=( (not A200)  and  a5425a );
 a5430a <=( (not A167)  and  (not A169) );
 a5431a <=( (not A170)  and  a5430a );
 a5434a <=( A200  and  A199 );
 a5437a <=( (not A203)  and  A202 );
 a5438a <=( a5437a  and  a5434a );
 a5442a <=( (not A167)  and  (not A169) );
 a5443a <=( (not A170)  and  a5442a );
 a5446a <=( A200  and  (not A199) );
 a5449a <=( A203  and  (not A202) );
 a5450a <=( a5449a  and  a5446a );
 a5454a <=( (not A167)  and  (not A169) );
 a5455a <=( (not A170)  and  a5454a );
 a5458a <=( (not A200)  and  A199 );
 a5461a <=( A203  and  (not A202) );
 a5462a <=( a5461a  and  a5458a );
 a5466a <=( (not A167)  and  (not A169) );
 a5467a <=( (not A170)  and  a5466a );
 a5470a <=( (not A200)  and  (not A199) );
 a5473a <=( (not A203)  and  A202 );
 a5474a <=( a5473a  and  a5470a );
 a5477a <=( (not A166)  and  A167 );
 a5480a <=( (not A200)  and  (not A199) );
 a5481a <=( a5480a  and  a5477a );
 a5484a <=( A232  and  (not A202) );
 a5488a <=( A300  and  A299 );
 a5489a <=( A234  and  a5488a );
 a5490a <=( a5489a  and  a5484a );
 a5493a <=( (not A166)  and  A167 );
 a5496a <=( (not A200)  and  (not A199) );
 a5497a <=( a5496a  and  a5493a );
 a5500a <=( A232  and  (not A202) );
 a5504a <=( A300  and  A298 );
 a5505a <=( A234  and  a5504a );
 a5506a <=( a5505a  and  a5500a );
 a5509a <=( (not A166)  and  A167 );
 a5512a <=( (not A200)  and  (not A199) );
 a5513a <=( a5512a  and  a5509a );
 a5516a <=( A232  and  (not A202) );
 a5520a <=( A267  and  A265 );
 a5521a <=( A234  and  a5520a );
 a5522a <=( a5521a  and  a5516a );
 a5525a <=( (not A166)  and  A167 );
 a5528a <=( (not A200)  and  (not A199) );
 a5529a <=( a5528a  and  a5525a );
 a5532a <=( A232  and  (not A202) );
 a5536a <=( A267  and  A266 );
 a5537a <=( A234  and  a5536a );
 a5538a <=( a5537a  and  a5532a );
 a5541a <=( (not A166)  and  A167 );
 a5544a <=( (not A200)  and  (not A199) );
 a5545a <=( a5544a  and  a5541a );
 a5548a <=( A233  and  (not A202) );
 a5552a <=( A300  and  A299 );
 a5553a <=( A234  and  a5552a );
 a5554a <=( a5553a  and  a5548a );
 a5557a <=( (not A166)  and  A167 );
 a5560a <=( (not A200)  and  (not A199) );
 a5561a <=( a5560a  and  a5557a );
 a5564a <=( A233  and  (not A202) );
 a5568a <=( A300  and  A298 );
 a5569a <=( A234  and  a5568a );
 a5570a <=( a5569a  and  a5564a );
 a5573a <=( (not A166)  and  A167 );
 a5576a <=( (not A200)  and  (not A199) );
 a5577a <=( a5576a  and  a5573a );
 a5580a <=( A233  and  (not A202) );
 a5584a <=( A267  and  A265 );
 a5585a <=( A234  and  a5584a );
 a5586a <=( a5585a  and  a5580a );
 a5589a <=( (not A166)  and  A167 );
 a5592a <=( (not A200)  and  (not A199) );
 a5593a <=( a5592a  and  a5589a );
 a5596a <=( A233  and  (not A202) );
 a5600a <=( A267  and  A266 );
 a5601a <=( A234  and  a5600a );
 a5602a <=( a5601a  and  a5596a );
 a5605a <=( (not A166)  and  A167 );
 a5608a <=( (not A200)  and  (not A199) );
 a5609a <=( a5608a  and  a5605a );
 a5612a <=( A232  and  A203 );
 a5616a <=( A300  and  A299 );
 a5617a <=( A234  and  a5616a );
 a5618a <=( a5617a  and  a5612a );
 a5621a <=( (not A166)  and  A167 );
 a5624a <=( (not A200)  and  (not A199) );
 a5625a <=( a5624a  and  a5621a );
 a5628a <=( A232  and  A203 );
 a5632a <=( A300  and  A298 );
 a5633a <=( A234  and  a5632a );
 a5634a <=( a5633a  and  a5628a );
 a5637a <=( (not A166)  and  A167 );
 a5640a <=( (not A200)  and  (not A199) );
 a5641a <=( a5640a  and  a5637a );
 a5644a <=( A232  and  A203 );
 a5648a <=( A267  and  A265 );
 a5649a <=( A234  and  a5648a );
 a5650a <=( a5649a  and  a5644a );
 a5653a <=( (not A166)  and  A167 );
 a5656a <=( (not A200)  and  (not A199) );
 a5657a <=( a5656a  and  a5653a );
 a5660a <=( A232  and  A203 );
 a5664a <=( A267  and  A266 );
 a5665a <=( A234  and  a5664a );
 a5666a <=( a5665a  and  a5660a );
 a5669a <=( (not A166)  and  A167 );
 a5672a <=( (not A200)  and  (not A199) );
 a5673a <=( a5672a  and  a5669a );
 a5676a <=( A233  and  A203 );
 a5680a <=( A300  and  A299 );
 a5681a <=( A234  and  a5680a );
 a5682a <=( a5681a  and  a5676a );
 a5685a <=( (not A166)  and  A167 );
 a5688a <=( (not A200)  and  (not A199) );
 a5689a <=( a5688a  and  a5685a );
 a5692a <=( A233  and  A203 );
 a5696a <=( A300  and  A298 );
 a5697a <=( A234  and  a5696a );
 a5698a <=( a5697a  and  a5692a );
 a5701a <=( (not A166)  and  A167 );
 a5704a <=( (not A200)  and  (not A199) );
 a5705a <=( a5704a  and  a5701a );
 a5708a <=( A233  and  A203 );
 a5712a <=( A267  and  A265 );
 a5713a <=( A234  and  a5712a );
 a5714a <=( a5713a  and  a5708a );
 a5717a <=( (not A166)  and  A167 );
 a5720a <=( (not A200)  and  (not A199) );
 a5721a <=( a5720a  and  a5717a );
 a5724a <=( A233  and  A203 );
 a5728a <=( A267  and  A266 );
 a5729a <=( A234  and  a5728a );
 a5730a <=( a5729a  and  a5724a );
 a5733a <=( (not A166)  and  A167 );
 a5737a <=( (not A201)  and  A200 );
 a5738a <=( A199  and  a5737a );
 a5739a <=( a5738a  and  a5733a );
 a5742a <=( A232  and  (not A202) );
 a5746a <=( A300  and  A299 );
 a5747a <=( A234  and  a5746a );
 a5748a <=( a5747a  and  a5742a );
 a5751a <=( (not A166)  and  A167 );
 a5755a <=( (not A201)  and  A200 );
 a5756a <=( A199  and  a5755a );
 a5757a <=( a5756a  and  a5751a );
 a5760a <=( A232  and  (not A202) );
 a5764a <=( A300  and  A298 );
 a5765a <=( A234  and  a5764a );
 a5766a <=( a5765a  and  a5760a );
 a5769a <=( (not A166)  and  A167 );
 a5773a <=( (not A201)  and  A200 );
 a5774a <=( A199  and  a5773a );
 a5775a <=( a5774a  and  a5769a );
 a5778a <=( A232  and  (not A202) );
 a5782a <=( A267  and  A265 );
 a5783a <=( A234  and  a5782a );
 a5784a <=( a5783a  and  a5778a );
 a5787a <=( (not A166)  and  A167 );
 a5791a <=( (not A201)  and  A200 );
 a5792a <=( A199  and  a5791a );
 a5793a <=( a5792a  and  a5787a );
 a5796a <=( A232  and  (not A202) );
 a5800a <=( A267  and  A266 );
 a5801a <=( A234  and  a5800a );
 a5802a <=( a5801a  and  a5796a );
 a5805a <=( (not A166)  and  A167 );
 a5809a <=( (not A201)  and  A200 );
 a5810a <=( A199  and  a5809a );
 a5811a <=( a5810a  and  a5805a );
 a5814a <=( A233  and  (not A202) );
 a5818a <=( A300  and  A299 );
 a5819a <=( A234  and  a5818a );
 a5820a <=( a5819a  and  a5814a );
 a5823a <=( (not A166)  and  A167 );
 a5827a <=( (not A201)  and  A200 );
 a5828a <=( A199  and  a5827a );
 a5829a <=( a5828a  and  a5823a );
 a5832a <=( A233  and  (not A202) );
 a5836a <=( A300  and  A298 );
 a5837a <=( A234  and  a5836a );
 a5838a <=( a5837a  and  a5832a );
 a5841a <=( (not A166)  and  A167 );
 a5845a <=( (not A201)  and  A200 );
 a5846a <=( A199  and  a5845a );
 a5847a <=( a5846a  and  a5841a );
 a5850a <=( A233  and  (not A202) );
 a5854a <=( A267  and  A265 );
 a5855a <=( A234  and  a5854a );
 a5856a <=( a5855a  and  a5850a );
 a5859a <=( (not A166)  and  A167 );
 a5863a <=( (not A201)  and  A200 );
 a5864a <=( A199  and  a5863a );
 a5865a <=( a5864a  and  a5859a );
 a5868a <=( A233  and  (not A202) );
 a5872a <=( A267  and  A266 );
 a5873a <=( A234  and  a5872a );
 a5874a <=( a5873a  and  a5868a );
 a5877a <=( (not A166)  and  A167 );
 a5881a <=( (not A201)  and  A200 );
 a5882a <=( A199  and  a5881a );
 a5883a <=( a5882a  and  a5877a );
 a5886a <=( A232  and  A203 );
 a5890a <=( A300  and  A299 );
 a5891a <=( A234  and  a5890a );
 a5892a <=( a5891a  and  a5886a );
 a5895a <=( (not A166)  and  A167 );
 a5899a <=( (not A201)  and  A200 );
 a5900a <=( A199  and  a5899a );
 a5901a <=( a5900a  and  a5895a );
 a5904a <=( A232  and  A203 );
 a5908a <=( A300  and  A298 );
 a5909a <=( A234  and  a5908a );
 a5910a <=( a5909a  and  a5904a );
 a5913a <=( (not A166)  and  A167 );
 a5917a <=( (not A201)  and  A200 );
 a5918a <=( A199  and  a5917a );
 a5919a <=( a5918a  and  a5913a );
 a5922a <=( A232  and  A203 );
 a5926a <=( A267  and  A265 );
 a5927a <=( A234  and  a5926a );
 a5928a <=( a5927a  and  a5922a );
 a5931a <=( (not A166)  and  A167 );
 a5935a <=( (not A201)  and  A200 );
 a5936a <=( A199  and  a5935a );
 a5937a <=( a5936a  and  a5931a );
 a5940a <=( A232  and  A203 );
 a5944a <=( A267  and  A266 );
 a5945a <=( A234  and  a5944a );
 a5946a <=( a5945a  and  a5940a );
 a5949a <=( (not A166)  and  A167 );
 a5953a <=( (not A201)  and  A200 );
 a5954a <=( A199  and  a5953a );
 a5955a <=( a5954a  and  a5949a );
 a5958a <=( A233  and  A203 );
 a5962a <=( A300  and  A299 );
 a5963a <=( A234  and  a5962a );
 a5964a <=( a5963a  and  a5958a );
 a5967a <=( (not A166)  and  A167 );
 a5971a <=( (not A201)  and  A200 );
 a5972a <=( A199  and  a5971a );
 a5973a <=( a5972a  and  a5967a );
 a5976a <=( A233  and  A203 );
 a5980a <=( A300  and  A298 );
 a5981a <=( A234  and  a5980a );
 a5982a <=( a5981a  and  a5976a );
 a5985a <=( (not A166)  and  A167 );
 a5989a <=( (not A201)  and  A200 );
 a5990a <=( A199  and  a5989a );
 a5991a <=( a5990a  and  a5985a );
 a5994a <=( A233  and  A203 );
 a5998a <=( A267  and  A265 );
 a5999a <=( A234  and  a5998a );
 a6000a <=( a5999a  and  a5994a );
 a6003a <=( (not A166)  and  A167 );
 a6007a <=( (not A201)  and  A200 );
 a6008a <=( A199  and  a6007a );
 a6009a <=( a6008a  and  a6003a );
 a6012a <=( A233  and  A203 );
 a6016a <=( A267  and  A266 );
 a6017a <=( A234  and  a6016a );
 a6018a <=( a6017a  and  a6012a );
 a6021a <=( (not A166)  and  A167 );
 a6025a <=( (not A201)  and  A200 );
 a6026a <=( (not A199)  and  a6025a );
 a6027a <=( a6026a  and  a6021a );
 a6030a <=( A232  and  A202 );
 a6034a <=( A300  and  A299 );
 a6035a <=( A234  and  a6034a );
 a6036a <=( a6035a  and  a6030a );
 a6039a <=( (not A166)  and  A167 );
 a6043a <=( (not A201)  and  A200 );
 a6044a <=( (not A199)  and  a6043a );
 a6045a <=( a6044a  and  a6039a );
 a6048a <=( A232  and  A202 );
 a6052a <=( A300  and  A298 );
 a6053a <=( A234  and  a6052a );
 a6054a <=( a6053a  and  a6048a );
 a6057a <=( (not A166)  and  A167 );
 a6061a <=( (not A201)  and  A200 );
 a6062a <=( (not A199)  and  a6061a );
 a6063a <=( a6062a  and  a6057a );
 a6066a <=( A232  and  A202 );
 a6070a <=( A267  and  A265 );
 a6071a <=( A234  and  a6070a );
 a6072a <=( a6071a  and  a6066a );
 a6075a <=( (not A166)  and  A167 );
 a6079a <=( (not A201)  and  A200 );
 a6080a <=( (not A199)  and  a6079a );
 a6081a <=( a6080a  and  a6075a );
 a6084a <=( A232  and  A202 );
 a6088a <=( A267  and  A266 );
 a6089a <=( A234  and  a6088a );
 a6090a <=( a6089a  and  a6084a );
 a6093a <=( (not A166)  and  A167 );
 a6097a <=( (not A201)  and  A200 );
 a6098a <=( (not A199)  and  a6097a );
 a6099a <=( a6098a  and  a6093a );
 a6102a <=( A233  and  A202 );
 a6106a <=( A300  and  A299 );
 a6107a <=( A234  and  a6106a );
 a6108a <=( a6107a  and  a6102a );
 a6111a <=( (not A166)  and  A167 );
 a6115a <=( (not A201)  and  A200 );
 a6116a <=( (not A199)  and  a6115a );
 a6117a <=( a6116a  and  a6111a );
 a6120a <=( A233  and  A202 );
 a6124a <=( A300  and  A298 );
 a6125a <=( A234  and  a6124a );
 a6126a <=( a6125a  and  a6120a );
 a6129a <=( (not A166)  and  A167 );
 a6133a <=( (not A201)  and  A200 );
 a6134a <=( (not A199)  and  a6133a );
 a6135a <=( a6134a  and  a6129a );
 a6138a <=( A233  and  A202 );
 a6142a <=( A267  and  A265 );
 a6143a <=( A234  and  a6142a );
 a6144a <=( a6143a  and  a6138a );
 a6147a <=( (not A166)  and  A167 );
 a6151a <=( (not A201)  and  A200 );
 a6152a <=( (not A199)  and  a6151a );
 a6153a <=( a6152a  and  a6147a );
 a6156a <=( A233  and  A202 );
 a6160a <=( A267  and  A266 );
 a6161a <=( A234  and  a6160a );
 a6162a <=( a6161a  and  a6156a );
 a6165a <=( (not A166)  and  A167 );
 a6169a <=( (not A201)  and  A200 );
 a6170a <=( (not A199)  and  a6169a );
 a6171a <=( a6170a  and  a6165a );
 a6174a <=( A232  and  (not A203) );
 a6178a <=( A300  and  A299 );
 a6179a <=( A234  and  a6178a );
 a6180a <=( a6179a  and  a6174a );
 a6183a <=( (not A166)  and  A167 );
 a6187a <=( (not A201)  and  A200 );
 a6188a <=( (not A199)  and  a6187a );
 a6189a <=( a6188a  and  a6183a );
 a6192a <=( A232  and  (not A203) );
 a6196a <=( A300  and  A298 );
 a6197a <=( A234  and  a6196a );
 a6198a <=( a6197a  and  a6192a );
 a6201a <=( (not A166)  and  A167 );
 a6205a <=( (not A201)  and  A200 );
 a6206a <=( (not A199)  and  a6205a );
 a6207a <=( a6206a  and  a6201a );
 a6210a <=( A232  and  (not A203) );
 a6214a <=( A267  and  A265 );
 a6215a <=( A234  and  a6214a );
 a6216a <=( a6215a  and  a6210a );
 a6219a <=( (not A166)  and  A167 );
 a6223a <=( (not A201)  and  A200 );
 a6224a <=( (not A199)  and  a6223a );
 a6225a <=( a6224a  and  a6219a );
 a6228a <=( A232  and  (not A203) );
 a6232a <=( A267  and  A266 );
 a6233a <=( A234  and  a6232a );
 a6234a <=( a6233a  and  a6228a );
 a6237a <=( (not A166)  and  A167 );
 a6241a <=( (not A201)  and  A200 );
 a6242a <=( (not A199)  and  a6241a );
 a6243a <=( a6242a  and  a6237a );
 a6246a <=( A233  and  (not A203) );
 a6250a <=( A300  and  A299 );
 a6251a <=( A234  and  a6250a );
 a6252a <=( a6251a  and  a6246a );
 a6255a <=( (not A166)  and  A167 );
 a6259a <=( (not A201)  and  A200 );
 a6260a <=( (not A199)  and  a6259a );
 a6261a <=( a6260a  and  a6255a );
 a6264a <=( A233  and  (not A203) );
 a6268a <=( A300  and  A298 );
 a6269a <=( A234  and  a6268a );
 a6270a <=( a6269a  and  a6264a );
 a6273a <=( (not A166)  and  A167 );
 a6277a <=( (not A201)  and  A200 );
 a6278a <=( (not A199)  and  a6277a );
 a6279a <=( a6278a  and  a6273a );
 a6282a <=( A233  and  (not A203) );
 a6286a <=( A267  and  A265 );
 a6287a <=( A234  and  a6286a );
 a6288a <=( a6287a  and  a6282a );
 a6291a <=( (not A166)  and  A167 );
 a6295a <=( (not A201)  and  A200 );
 a6296a <=( (not A199)  and  a6295a );
 a6297a <=( a6296a  and  a6291a );
 a6300a <=( A233  and  (not A203) );
 a6304a <=( A267  and  A266 );
 a6305a <=( A234  and  a6304a );
 a6306a <=( a6305a  and  a6300a );
 a6309a <=( (not A166)  and  A167 );
 a6313a <=( (not A201)  and  (not A200) );
 a6314a <=( A199  and  a6313a );
 a6315a <=( a6314a  and  a6309a );
 a6318a <=( A232  and  A202 );
 a6322a <=( A300  and  A299 );
 a6323a <=( A234  and  a6322a );
 a6324a <=( a6323a  and  a6318a );
 a6327a <=( (not A166)  and  A167 );
 a6331a <=( (not A201)  and  (not A200) );
 a6332a <=( A199  and  a6331a );
 a6333a <=( a6332a  and  a6327a );
 a6336a <=( A232  and  A202 );
 a6340a <=( A300  and  A298 );
 a6341a <=( A234  and  a6340a );
 a6342a <=( a6341a  and  a6336a );
 a6345a <=( (not A166)  and  A167 );
 a6349a <=( (not A201)  and  (not A200) );
 a6350a <=( A199  and  a6349a );
 a6351a <=( a6350a  and  a6345a );
 a6354a <=( A232  and  A202 );
 a6358a <=( A267  and  A265 );
 a6359a <=( A234  and  a6358a );
 a6360a <=( a6359a  and  a6354a );
 a6363a <=( (not A166)  and  A167 );
 a6367a <=( (not A201)  and  (not A200) );
 a6368a <=( A199  and  a6367a );
 a6369a <=( a6368a  and  a6363a );
 a6372a <=( A232  and  A202 );
 a6376a <=( A267  and  A266 );
 a6377a <=( A234  and  a6376a );
 a6378a <=( a6377a  and  a6372a );
 a6381a <=( (not A166)  and  A167 );
 a6385a <=( (not A201)  and  (not A200) );
 a6386a <=( A199  and  a6385a );
 a6387a <=( a6386a  and  a6381a );
 a6390a <=( A233  and  A202 );
 a6394a <=( A300  and  A299 );
 a6395a <=( A234  and  a6394a );
 a6396a <=( a6395a  and  a6390a );
 a6399a <=( (not A166)  and  A167 );
 a6403a <=( (not A201)  and  (not A200) );
 a6404a <=( A199  and  a6403a );
 a6405a <=( a6404a  and  a6399a );
 a6408a <=( A233  and  A202 );
 a6412a <=( A300  and  A298 );
 a6413a <=( A234  and  a6412a );
 a6414a <=( a6413a  and  a6408a );
 a6417a <=( (not A166)  and  A167 );
 a6421a <=( (not A201)  and  (not A200) );
 a6422a <=( A199  and  a6421a );
 a6423a <=( a6422a  and  a6417a );
 a6426a <=( A233  and  A202 );
 a6430a <=( A267  and  A265 );
 a6431a <=( A234  and  a6430a );
 a6432a <=( a6431a  and  a6426a );
 a6435a <=( (not A166)  and  A167 );
 a6439a <=( (not A201)  and  (not A200) );
 a6440a <=( A199  and  a6439a );
 a6441a <=( a6440a  and  a6435a );
 a6444a <=( A233  and  A202 );
 a6448a <=( A267  and  A266 );
 a6449a <=( A234  and  a6448a );
 a6450a <=( a6449a  and  a6444a );
 a6453a <=( (not A166)  and  A167 );
 a6457a <=( (not A201)  and  (not A200) );
 a6458a <=( A199  and  a6457a );
 a6459a <=( a6458a  and  a6453a );
 a6462a <=( A232  and  (not A203) );
 a6466a <=( A300  and  A299 );
 a6467a <=( A234  and  a6466a );
 a6468a <=( a6467a  and  a6462a );
 a6471a <=( (not A166)  and  A167 );
 a6475a <=( (not A201)  and  (not A200) );
 a6476a <=( A199  and  a6475a );
 a6477a <=( a6476a  and  a6471a );
 a6480a <=( A232  and  (not A203) );
 a6484a <=( A300  and  A298 );
 a6485a <=( A234  and  a6484a );
 a6486a <=( a6485a  and  a6480a );
 a6489a <=( (not A166)  and  A167 );
 a6493a <=( (not A201)  and  (not A200) );
 a6494a <=( A199  and  a6493a );
 a6495a <=( a6494a  and  a6489a );
 a6498a <=( A232  and  (not A203) );
 a6502a <=( A267  and  A265 );
 a6503a <=( A234  and  a6502a );
 a6504a <=( a6503a  and  a6498a );
 a6507a <=( (not A166)  and  A167 );
 a6511a <=( (not A201)  and  (not A200) );
 a6512a <=( A199  and  a6511a );
 a6513a <=( a6512a  and  a6507a );
 a6516a <=( A232  and  (not A203) );
 a6520a <=( A267  and  A266 );
 a6521a <=( A234  and  a6520a );
 a6522a <=( a6521a  and  a6516a );
 a6525a <=( (not A166)  and  A167 );
 a6529a <=( (not A201)  and  (not A200) );
 a6530a <=( A199  and  a6529a );
 a6531a <=( a6530a  and  a6525a );
 a6534a <=( A233  and  (not A203) );
 a6538a <=( A300  and  A299 );
 a6539a <=( A234  and  a6538a );
 a6540a <=( a6539a  and  a6534a );
 a6543a <=( (not A166)  and  A167 );
 a6547a <=( (not A201)  and  (not A200) );
 a6548a <=( A199  and  a6547a );
 a6549a <=( a6548a  and  a6543a );
 a6552a <=( A233  and  (not A203) );
 a6556a <=( A300  and  A298 );
 a6557a <=( A234  and  a6556a );
 a6558a <=( a6557a  and  a6552a );
 a6561a <=( (not A166)  and  A167 );
 a6565a <=( (not A201)  and  (not A200) );
 a6566a <=( A199  and  a6565a );
 a6567a <=( a6566a  and  a6561a );
 a6570a <=( A233  and  (not A203) );
 a6574a <=( A267  and  A265 );
 a6575a <=( A234  and  a6574a );
 a6576a <=( a6575a  and  a6570a );
 a6579a <=( (not A166)  and  A167 );
 a6583a <=( (not A201)  and  (not A200) );
 a6584a <=( A199  and  a6583a );
 a6585a <=( a6584a  and  a6579a );
 a6588a <=( A233  and  (not A203) );
 a6592a <=( A267  and  A266 );
 a6593a <=( A234  and  a6592a );
 a6594a <=( a6593a  and  a6588a );
 a6597a <=( (not A166)  and  A167 );
 a6601a <=( (not A202)  and  (not A200) );
 a6602a <=( (not A199)  and  a6601a );
 a6603a <=( a6602a  and  a6597a );
 a6607a <=( A298  and  A234 );
 a6608a <=( A232  and  a6607a );
 a6612a <=( (not A302)  and  A301 );
 a6613a <=( A299  and  a6612a );
 a6614a <=( a6613a  and  a6608a );
 a6617a <=( (not A166)  and  A167 );
 a6621a <=( (not A202)  and  (not A200) );
 a6622a <=( (not A199)  and  a6621a );
 a6623a <=( a6622a  and  a6617a );
 a6627a <=( A298  and  A234 );
 a6628a <=( A232  and  a6627a );
 a6632a <=( A302  and  (not A301) );
 a6633a <=( (not A299)  and  a6632a );
 a6634a <=( a6633a  and  a6628a );
 a6637a <=( (not A166)  and  A167 );
 a6641a <=( (not A202)  and  (not A200) );
 a6642a <=( (not A199)  and  a6641a );
 a6643a <=( a6642a  and  a6637a );
 a6647a <=( (not A298)  and  A234 );
 a6648a <=( A232  and  a6647a );
 a6652a <=( A302  and  (not A301) );
 a6653a <=( A299  and  a6652a );
 a6654a <=( a6653a  and  a6648a );
 a6657a <=( (not A166)  and  A167 );
 a6661a <=( (not A202)  and  (not A200) );
 a6662a <=( (not A199)  and  a6661a );
 a6663a <=( a6662a  and  a6657a );
 a6667a <=( (not A298)  and  A234 );
 a6668a <=( A232  and  a6667a );
 a6672a <=( (not A302)  and  A301 );
 a6673a <=( (not A299)  and  a6672a );
 a6674a <=( a6673a  and  a6668a );
 a6677a <=( (not A166)  and  A167 );
 a6681a <=( (not A202)  and  (not A200) );
 a6682a <=( (not A199)  and  a6681a );
 a6683a <=( a6682a  and  a6677a );
 a6687a <=( A265  and  A234 );
 a6688a <=( A232  and  a6687a );
 a6692a <=( (not A269)  and  A268 );
 a6693a <=( A266  and  a6692a );
 a6694a <=( a6693a  and  a6688a );
 a6697a <=( (not A166)  and  A167 );
 a6701a <=( (not A202)  and  (not A200) );
 a6702a <=( (not A199)  and  a6701a );
 a6703a <=( a6702a  and  a6697a );
 a6707a <=( (not A265)  and  A234 );
 a6708a <=( A232  and  a6707a );
 a6712a <=( A269  and  (not A268) );
 a6713a <=( A266  and  a6712a );
 a6714a <=( a6713a  and  a6708a );
 a6717a <=( (not A166)  and  A167 );
 a6721a <=( (not A202)  and  (not A200) );
 a6722a <=( (not A199)  and  a6721a );
 a6723a <=( a6722a  and  a6717a );
 a6727a <=( A265  and  A234 );
 a6728a <=( A232  and  a6727a );
 a6732a <=( A269  and  (not A268) );
 a6733a <=( (not A266)  and  a6732a );
 a6734a <=( a6733a  and  a6728a );
 a6737a <=( (not A166)  and  A167 );
 a6741a <=( (not A202)  and  (not A200) );
 a6742a <=( (not A199)  and  a6741a );
 a6743a <=( a6742a  and  a6737a );
 a6747a <=( (not A265)  and  A234 );
 a6748a <=( A232  and  a6747a );
 a6752a <=( (not A269)  and  A268 );
 a6753a <=( (not A266)  and  a6752a );
 a6754a <=( a6753a  and  a6748a );
 a6757a <=( (not A166)  and  A167 );
 a6761a <=( (not A202)  and  (not A200) );
 a6762a <=( (not A199)  and  a6761a );
 a6763a <=( a6762a  and  a6757a );
 a6767a <=( A298  and  A234 );
 a6768a <=( A233  and  a6767a );
 a6772a <=( (not A302)  and  A301 );
 a6773a <=( A299  and  a6772a );
 a6774a <=( a6773a  and  a6768a );
 a6777a <=( (not A166)  and  A167 );
 a6781a <=( (not A202)  and  (not A200) );
 a6782a <=( (not A199)  and  a6781a );
 a6783a <=( a6782a  and  a6777a );
 a6787a <=( A298  and  A234 );
 a6788a <=( A233  and  a6787a );
 a6792a <=( A302  and  (not A301) );
 a6793a <=( (not A299)  and  a6792a );
 a6794a <=( a6793a  and  a6788a );
 a6797a <=( (not A166)  and  A167 );
 a6801a <=( (not A202)  and  (not A200) );
 a6802a <=( (not A199)  and  a6801a );
 a6803a <=( a6802a  and  a6797a );
 a6807a <=( (not A298)  and  A234 );
 a6808a <=( A233  and  a6807a );
 a6812a <=( A302  and  (not A301) );
 a6813a <=( A299  and  a6812a );
 a6814a <=( a6813a  and  a6808a );
 a6817a <=( (not A166)  and  A167 );
 a6821a <=( (not A202)  and  (not A200) );
 a6822a <=( (not A199)  and  a6821a );
 a6823a <=( a6822a  and  a6817a );
 a6827a <=( (not A298)  and  A234 );
 a6828a <=( A233  and  a6827a );
 a6832a <=( (not A302)  and  A301 );
 a6833a <=( (not A299)  and  a6832a );
 a6834a <=( a6833a  and  a6828a );
 a6837a <=( (not A166)  and  A167 );
 a6841a <=( (not A202)  and  (not A200) );
 a6842a <=( (not A199)  and  a6841a );
 a6843a <=( a6842a  and  a6837a );
 a6847a <=( A265  and  A234 );
 a6848a <=( A233  and  a6847a );
 a6852a <=( (not A269)  and  A268 );
 a6853a <=( A266  and  a6852a );
 a6854a <=( a6853a  and  a6848a );
 a6857a <=( (not A166)  and  A167 );
 a6861a <=( (not A202)  and  (not A200) );
 a6862a <=( (not A199)  and  a6861a );
 a6863a <=( a6862a  and  a6857a );
 a6867a <=( (not A265)  and  A234 );
 a6868a <=( A233  and  a6867a );
 a6872a <=( A269  and  (not A268) );
 a6873a <=( A266  and  a6872a );
 a6874a <=( a6873a  and  a6868a );
 a6877a <=( (not A166)  and  A167 );
 a6881a <=( (not A202)  and  (not A200) );
 a6882a <=( (not A199)  and  a6881a );
 a6883a <=( a6882a  and  a6877a );
 a6887a <=( A265  and  A234 );
 a6888a <=( A233  and  a6887a );
 a6892a <=( A269  and  (not A268) );
 a6893a <=( (not A266)  and  a6892a );
 a6894a <=( a6893a  and  a6888a );
 a6897a <=( (not A166)  and  A167 );
 a6901a <=( (not A202)  and  (not A200) );
 a6902a <=( (not A199)  and  a6901a );
 a6903a <=( a6902a  and  a6897a );
 a6907a <=( (not A265)  and  A234 );
 a6908a <=( A233  and  a6907a );
 a6912a <=( (not A269)  and  A268 );
 a6913a <=( (not A266)  and  a6912a );
 a6914a <=( a6913a  and  a6908a );
 a6917a <=( (not A166)  and  A167 );
 a6921a <=( (not A202)  and  (not A200) );
 a6922a <=( (not A199)  and  a6921a );
 a6923a <=( a6922a  and  a6917a );
 a6927a <=( A235  and  A233 );
 a6928a <=( A232  and  a6927a );
 a6932a <=( A300  and  A299 );
 a6933a <=( (not A236)  and  a6932a );
 a6934a <=( a6933a  and  a6928a );
 a6937a <=( (not A166)  and  A167 );
 a6941a <=( (not A202)  and  (not A200) );
 a6942a <=( (not A199)  and  a6941a );
 a6943a <=( a6942a  and  a6937a );
 a6947a <=( A235  and  A233 );
 a6948a <=( A232  and  a6947a );
 a6952a <=( A300  and  A298 );
 a6953a <=( (not A236)  and  a6952a );
 a6954a <=( a6953a  and  a6948a );
 a6957a <=( (not A166)  and  A167 );
 a6961a <=( (not A202)  and  (not A200) );
 a6962a <=( (not A199)  and  a6961a );
 a6963a <=( a6962a  and  a6957a );
 a6967a <=( A235  and  A233 );
 a6968a <=( A232  and  a6967a );
 a6972a <=( A267  and  A265 );
 a6973a <=( (not A236)  and  a6972a );
 a6974a <=( a6973a  and  a6968a );
 a6977a <=( (not A166)  and  A167 );
 a6981a <=( (not A202)  and  (not A200) );
 a6982a <=( (not A199)  and  a6981a );
 a6983a <=( a6982a  and  a6977a );
 a6987a <=( A235  and  A233 );
 a6988a <=( A232  and  a6987a );
 a6992a <=( A267  and  A266 );
 a6993a <=( (not A236)  and  a6992a );
 a6994a <=( a6993a  and  a6988a );
 a6997a <=( (not A166)  and  A167 );
 a7001a <=( (not A202)  and  (not A200) );
 a7002a <=( (not A199)  and  a7001a );
 a7003a <=( a7002a  and  a6997a );
 a7007a <=( (not A235)  and  A233 );
 a7008a <=( (not A232)  and  a7007a );
 a7012a <=( A300  and  A299 );
 a7013a <=( A236  and  a7012a );
 a7014a <=( a7013a  and  a7008a );
 a7017a <=( (not A166)  and  A167 );
 a7021a <=( (not A202)  and  (not A200) );
 a7022a <=( (not A199)  and  a7021a );
 a7023a <=( a7022a  and  a7017a );
 a7027a <=( (not A235)  and  A233 );
 a7028a <=( (not A232)  and  a7027a );
 a7032a <=( A300  and  A298 );
 a7033a <=( A236  and  a7032a );
 a7034a <=( a7033a  and  a7028a );
 a7037a <=( (not A166)  and  A167 );
 a7041a <=( (not A202)  and  (not A200) );
 a7042a <=( (not A199)  and  a7041a );
 a7043a <=( a7042a  and  a7037a );
 a7047a <=( (not A235)  and  A233 );
 a7048a <=( (not A232)  and  a7047a );
 a7052a <=( A267  and  A265 );
 a7053a <=( A236  and  a7052a );
 a7054a <=( a7053a  and  a7048a );
 a7057a <=( (not A166)  and  A167 );
 a7061a <=( (not A202)  and  (not A200) );
 a7062a <=( (not A199)  and  a7061a );
 a7063a <=( a7062a  and  a7057a );
 a7067a <=( (not A235)  and  A233 );
 a7068a <=( (not A232)  and  a7067a );
 a7072a <=( A267  and  A266 );
 a7073a <=( A236  and  a7072a );
 a7074a <=( a7073a  and  a7068a );
 a7077a <=( (not A166)  and  A167 );
 a7081a <=( (not A202)  and  (not A200) );
 a7082a <=( (not A199)  and  a7081a );
 a7083a <=( a7082a  and  a7077a );
 a7087a <=( (not A235)  and  (not A233) );
 a7088a <=( A232  and  a7087a );
 a7092a <=( A300  and  A299 );
 a7093a <=( A236  and  a7092a );
 a7094a <=( a7093a  and  a7088a );
 a7097a <=( (not A166)  and  A167 );
 a7101a <=( (not A202)  and  (not A200) );
 a7102a <=( (not A199)  and  a7101a );
 a7103a <=( a7102a  and  a7097a );
 a7107a <=( (not A235)  and  (not A233) );
 a7108a <=( A232  and  a7107a );
 a7112a <=( A300  and  A298 );
 a7113a <=( A236  and  a7112a );
 a7114a <=( a7113a  and  a7108a );
 a7117a <=( (not A166)  and  A167 );
 a7121a <=( (not A202)  and  (not A200) );
 a7122a <=( (not A199)  and  a7121a );
 a7123a <=( a7122a  and  a7117a );
 a7127a <=( (not A235)  and  (not A233) );
 a7128a <=( A232  and  a7127a );
 a7132a <=( A267  and  A265 );
 a7133a <=( A236  and  a7132a );
 a7134a <=( a7133a  and  a7128a );
 a7137a <=( (not A166)  and  A167 );
 a7141a <=( (not A202)  and  (not A200) );
 a7142a <=( (not A199)  and  a7141a );
 a7143a <=( a7142a  and  a7137a );
 a7147a <=( (not A235)  and  (not A233) );
 a7148a <=( A232  and  a7147a );
 a7152a <=( A267  and  A266 );
 a7153a <=( A236  and  a7152a );
 a7154a <=( a7153a  and  a7148a );
 a7157a <=( (not A166)  and  A167 );
 a7161a <=( (not A202)  and  (not A200) );
 a7162a <=( (not A199)  and  a7161a );
 a7163a <=( a7162a  and  a7157a );
 a7167a <=( A235  and  (not A233) );
 a7168a <=( (not A232)  and  a7167a );
 a7172a <=( A300  and  A299 );
 a7173a <=( (not A236)  and  a7172a );
 a7174a <=( a7173a  and  a7168a );
 a7177a <=( (not A166)  and  A167 );
 a7181a <=( (not A202)  and  (not A200) );
 a7182a <=( (not A199)  and  a7181a );
 a7183a <=( a7182a  and  a7177a );
 a7187a <=( A235  and  (not A233) );
 a7188a <=( (not A232)  and  a7187a );
 a7192a <=( A300  and  A298 );
 a7193a <=( (not A236)  and  a7192a );
 a7194a <=( a7193a  and  a7188a );
 a7197a <=( (not A166)  and  A167 );
 a7201a <=( (not A202)  and  (not A200) );
 a7202a <=( (not A199)  and  a7201a );
 a7203a <=( a7202a  and  a7197a );
 a7207a <=( A235  and  (not A233) );
 a7208a <=( (not A232)  and  a7207a );
 a7212a <=( A267  and  A265 );
 a7213a <=( (not A236)  and  a7212a );
 a7214a <=( a7213a  and  a7208a );
 a7217a <=( (not A166)  and  A167 );
 a7221a <=( (not A202)  and  (not A200) );
 a7222a <=( (not A199)  and  a7221a );
 a7223a <=( a7222a  and  a7217a );
 a7227a <=( A235  and  (not A233) );
 a7228a <=( (not A232)  and  a7227a );
 a7232a <=( A267  and  A266 );
 a7233a <=( (not A236)  and  a7232a );
 a7234a <=( a7233a  and  a7228a );
 a7237a <=( (not A166)  and  A167 );
 a7241a <=( A203  and  (not A200) );
 a7242a <=( (not A199)  and  a7241a );
 a7243a <=( a7242a  and  a7237a );
 a7247a <=( A298  and  A234 );
 a7248a <=( A232  and  a7247a );
 a7252a <=( (not A302)  and  A301 );
 a7253a <=( A299  and  a7252a );
 a7254a <=( a7253a  and  a7248a );
 a7257a <=( (not A166)  and  A167 );
 a7261a <=( A203  and  (not A200) );
 a7262a <=( (not A199)  and  a7261a );
 a7263a <=( a7262a  and  a7257a );
 a7267a <=( A298  and  A234 );
 a7268a <=( A232  and  a7267a );
 a7272a <=( A302  and  (not A301) );
 a7273a <=( (not A299)  and  a7272a );
 a7274a <=( a7273a  and  a7268a );
 a7277a <=( (not A166)  and  A167 );
 a7281a <=( A203  and  (not A200) );
 a7282a <=( (not A199)  and  a7281a );
 a7283a <=( a7282a  and  a7277a );
 a7287a <=( (not A298)  and  A234 );
 a7288a <=( A232  and  a7287a );
 a7292a <=( A302  and  (not A301) );
 a7293a <=( A299  and  a7292a );
 a7294a <=( a7293a  and  a7288a );
 a7297a <=( (not A166)  and  A167 );
 a7301a <=( A203  and  (not A200) );
 a7302a <=( (not A199)  and  a7301a );
 a7303a <=( a7302a  and  a7297a );
 a7307a <=( (not A298)  and  A234 );
 a7308a <=( A232  and  a7307a );
 a7312a <=( (not A302)  and  A301 );
 a7313a <=( (not A299)  and  a7312a );
 a7314a <=( a7313a  and  a7308a );
 a7317a <=( (not A166)  and  A167 );
 a7321a <=( A203  and  (not A200) );
 a7322a <=( (not A199)  and  a7321a );
 a7323a <=( a7322a  and  a7317a );
 a7327a <=( A265  and  A234 );
 a7328a <=( A232  and  a7327a );
 a7332a <=( (not A269)  and  A268 );
 a7333a <=( A266  and  a7332a );
 a7334a <=( a7333a  and  a7328a );
 a7337a <=( (not A166)  and  A167 );
 a7341a <=( A203  and  (not A200) );
 a7342a <=( (not A199)  and  a7341a );
 a7343a <=( a7342a  and  a7337a );
 a7347a <=( (not A265)  and  A234 );
 a7348a <=( A232  and  a7347a );
 a7352a <=( A269  and  (not A268) );
 a7353a <=( A266  and  a7352a );
 a7354a <=( a7353a  and  a7348a );
 a7357a <=( (not A166)  and  A167 );
 a7361a <=( A203  and  (not A200) );
 a7362a <=( (not A199)  and  a7361a );
 a7363a <=( a7362a  and  a7357a );
 a7367a <=( A265  and  A234 );
 a7368a <=( A232  and  a7367a );
 a7372a <=( A269  and  (not A268) );
 a7373a <=( (not A266)  and  a7372a );
 a7374a <=( a7373a  and  a7368a );
 a7377a <=( (not A166)  and  A167 );
 a7381a <=( A203  and  (not A200) );
 a7382a <=( (not A199)  and  a7381a );
 a7383a <=( a7382a  and  a7377a );
 a7387a <=( (not A265)  and  A234 );
 a7388a <=( A232  and  a7387a );
 a7392a <=( (not A269)  and  A268 );
 a7393a <=( (not A266)  and  a7392a );
 a7394a <=( a7393a  and  a7388a );
 a7397a <=( (not A166)  and  A167 );
 a7401a <=( A203  and  (not A200) );
 a7402a <=( (not A199)  and  a7401a );
 a7403a <=( a7402a  and  a7397a );
 a7407a <=( A298  and  A234 );
 a7408a <=( A233  and  a7407a );
 a7412a <=( (not A302)  and  A301 );
 a7413a <=( A299  and  a7412a );
 a7414a <=( a7413a  and  a7408a );
 a7417a <=( (not A166)  and  A167 );
 a7421a <=( A203  and  (not A200) );
 a7422a <=( (not A199)  and  a7421a );
 a7423a <=( a7422a  and  a7417a );
 a7427a <=( A298  and  A234 );
 a7428a <=( A233  and  a7427a );
 a7432a <=( A302  and  (not A301) );
 a7433a <=( (not A299)  and  a7432a );
 a7434a <=( a7433a  and  a7428a );
 a7437a <=( (not A166)  and  A167 );
 a7441a <=( A203  and  (not A200) );
 a7442a <=( (not A199)  and  a7441a );
 a7443a <=( a7442a  and  a7437a );
 a7447a <=( (not A298)  and  A234 );
 a7448a <=( A233  and  a7447a );
 a7452a <=( A302  and  (not A301) );
 a7453a <=( A299  and  a7452a );
 a7454a <=( a7453a  and  a7448a );
 a7457a <=( (not A166)  and  A167 );
 a7461a <=( A203  and  (not A200) );
 a7462a <=( (not A199)  and  a7461a );
 a7463a <=( a7462a  and  a7457a );
 a7467a <=( (not A298)  and  A234 );
 a7468a <=( A233  and  a7467a );
 a7472a <=( (not A302)  and  A301 );
 a7473a <=( (not A299)  and  a7472a );
 a7474a <=( a7473a  and  a7468a );
 a7477a <=( (not A166)  and  A167 );
 a7481a <=( A203  and  (not A200) );
 a7482a <=( (not A199)  and  a7481a );
 a7483a <=( a7482a  and  a7477a );
 a7487a <=( A265  and  A234 );
 a7488a <=( A233  and  a7487a );
 a7492a <=( (not A269)  and  A268 );
 a7493a <=( A266  and  a7492a );
 a7494a <=( a7493a  and  a7488a );
 a7497a <=( (not A166)  and  A167 );
 a7501a <=( A203  and  (not A200) );
 a7502a <=( (not A199)  and  a7501a );
 a7503a <=( a7502a  and  a7497a );
 a7507a <=( (not A265)  and  A234 );
 a7508a <=( A233  and  a7507a );
 a7512a <=( A269  and  (not A268) );
 a7513a <=( A266  and  a7512a );
 a7514a <=( a7513a  and  a7508a );
 a7517a <=( (not A166)  and  A167 );
 a7521a <=( A203  and  (not A200) );
 a7522a <=( (not A199)  and  a7521a );
 a7523a <=( a7522a  and  a7517a );
 a7527a <=( A265  and  A234 );
 a7528a <=( A233  and  a7527a );
 a7532a <=( A269  and  (not A268) );
 a7533a <=( (not A266)  and  a7532a );
 a7534a <=( a7533a  and  a7528a );
 a7537a <=( (not A166)  and  A167 );
 a7541a <=( A203  and  (not A200) );
 a7542a <=( (not A199)  and  a7541a );
 a7543a <=( a7542a  and  a7537a );
 a7547a <=( (not A265)  and  A234 );
 a7548a <=( A233  and  a7547a );
 a7552a <=( (not A269)  and  A268 );
 a7553a <=( (not A266)  and  a7552a );
 a7554a <=( a7553a  and  a7548a );
 a7557a <=( (not A166)  and  A167 );
 a7561a <=( A203  and  (not A200) );
 a7562a <=( (not A199)  and  a7561a );
 a7563a <=( a7562a  and  a7557a );
 a7567a <=( A235  and  A233 );
 a7568a <=( A232  and  a7567a );
 a7572a <=( A300  and  A299 );
 a7573a <=( (not A236)  and  a7572a );
 a7574a <=( a7573a  and  a7568a );
 a7577a <=( (not A166)  and  A167 );
 a7581a <=( A203  and  (not A200) );
 a7582a <=( (not A199)  and  a7581a );
 a7583a <=( a7582a  and  a7577a );
 a7587a <=( A235  and  A233 );
 a7588a <=( A232  and  a7587a );
 a7592a <=( A300  and  A298 );
 a7593a <=( (not A236)  and  a7592a );
 a7594a <=( a7593a  and  a7588a );
 a7597a <=( (not A166)  and  A167 );
 a7601a <=( A203  and  (not A200) );
 a7602a <=( (not A199)  and  a7601a );
 a7603a <=( a7602a  and  a7597a );
 a7607a <=( A235  and  A233 );
 a7608a <=( A232  and  a7607a );
 a7612a <=( A267  and  A265 );
 a7613a <=( (not A236)  and  a7612a );
 a7614a <=( a7613a  and  a7608a );
 a7617a <=( (not A166)  and  A167 );
 a7621a <=( A203  and  (not A200) );
 a7622a <=( (not A199)  and  a7621a );
 a7623a <=( a7622a  and  a7617a );
 a7627a <=( A235  and  A233 );
 a7628a <=( A232  and  a7627a );
 a7632a <=( A267  and  A266 );
 a7633a <=( (not A236)  and  a7632a );
 a7634a <=( a7633a  and  a7628a );
 a7637a <=( (not A166)  and  A167 );
 a7641a <=( A203  and  (not A200) );
 a7642a <=( (not A199)  and  a7641a );
 a7643a <=( a7642a  and  a7637a );
 a7647a <=( (not A235)  and  A233 );
 a7648a <=( (not A232)  and  a7647a );
 a7652a <=( A300  and  A299 );
 a7653a <=( A236  and  a7652a );
 a7654a <=( a7653a  and  a7648a );
 a7657a <=( (not A166)  and  A167 );
 a7661a <=( A203  and  (not A200) );
 a7662a <=( (not A199)  and  a7661a );
 a7663a <=( a7662a  and  a7657a );
 a7667a <=( (not A235)  and  A233 );
 a7668a <=( (not A232)  and  a7667a );
 a7672a <=( A300  and  A298 );
 a7673a <=( A236  and  a7672a );
 a7674a <=( a7673a  and  a7668a );
 a7677a <=( (not A166)  and  A167 );
 a7681a <=( A203  and  (not A200) );
 a7682a <=( (not A199)  and  a7681a );
 a7683a <=( a7682a  and  a7677a );
 a7687a <=( (not A235)  and  A233 );
 a7688a <=( (not A232)  and  a7687a );
 a7692a <=( A267  and  A265 );
 a7693a <=( A236  and  a7692a );
 a7694a <=( a7693a  and  a7688a );
 a7697a <=( (not A166)  and  A167 );
 a7701a <=( A203  and  (not A200) );
 a7702a <=( (not A199)  and  a7701a );
 a7703a <=( a7702a  and  a7697a );
 a7707a <=( (not A235)  and  A233 );
 a7708a <=( (not A232)  and  a7707a );
 a7712a <=( A267  and  A266 );
 a7713a <=( A236  and  a7712a );
 a7714a <=( a7713a  and  a7708a );
 a7717a <=( (not A166)  and  A167 );
 a7721a <=( A203  and  (not A200) );
 a7722a <=( (not A199)  and  a7721a );
 a7723a <=( a7722a  and  a7717a );
 a7727a <=( (not A235)  and  (not A233) );
 a7728a <=( A232  and  a7727a );
 a7732a <=( A300  and  A299 );
 a7733a <=( A236  and  a7732a );
 a7734a <=( a7733a  and  a7728a );
 a7737a <=( (not A166)  and  A167 );
 a7741a <=( A203  and  (not A200) );
 a7742a <=( (not A199)  and  a7741a );
 a7743a <=( a7742a  and  a7737a );
 a7747a <=( (not A235)  and  (not A233) );
 a7748a <=( A232  and  a7747a );
 a7752a <=( A300  and  A298 );
 a7753a <=( A236  and  a7752a );
 a7754a <=( a7753a  and  a7748a );
 a7757a <=( (not A166)  and  A167 );
 a7761a <=( A203  and  (not A200) );
 a7762a <=( (not A199)  and  a7761a );
 a7763a <=( a7762a  and  a7757a );
 a7767a <=( (not A235)  and  (not A233) );
 a7768a <=( A232  and  a7767a );
 a7772a <=( A267  and  A265 );
 a7773a <=( A236  and  a7772a );
 a7774a <=( a7773a  and  a7768a );
 a7777a <=( (not A166)  and  A167 );
 a7781a <=( A203  and  (not A200) );
 a7782a <=( (not A199)  and  a7781a );
 a7783a <=( a7782a  and  a7777a );
 a7787a <=( (not A235)  and  (not A233) );
 a7788a <=( A232  and  a7787a );
 a7792a <=( A267  and  A266 );
 a7793a <=( A236  and  a7792a );
 a7794a <=( a7793a  and  a7788a );
 a7797a <=( (not A166)  and  A167 );
 a7801a <=( A203  and  (not A200) );
 a7802a <=( (not A199)  and  a7801a );
 a7803a <=( a7802a  and  a7797a );
 a7807a <=( A235  and  (not A233) );
 a7808a <=( (not A232)  and  a7807a );
 a7812a <=( A300  and  A299 );
 a7813a <=( (not A236)  and  a7812a );
 a7814a <=( a7813a  and  a7808a );
 a7817a <=( (not A166)  and  A167 );
 a7821a <=( A203  and  (not A200) );
 a7822a <=( (not A199)  and  a7821a );
 a7823a <=( a7822a  and  a7817a );
 a7827a <=( A235  and  (not A233) );
 a7828a <=( (not A232)  and  a7827a );
 a7832a <=( A300  and  A298 );
 a7833a <=( (not A236)  and  a7832a );
 a7834a <=( a7833a  and  a7828a );
 a7837a <=( (not A166)  and  A167 );
 a7841a <=( A203  and  (not A200) );
 a7842a <=( (not A199)  and  a7841a );
 a7843a <=( a7842a  and  a7837a );
 a7847a <=( A235  and  (not A233) );
 a7848a <=( (not A232)  and  a7847a );
 a7852a <=( A267  and  A265 );
 a7853a <=( (not A236)  and  a7852a );
 a7854a <=( a7853a  and  a7848a );
 a7857a <=( (not A166)  and  A167 );
 a7861a <=( A203  and  (not A200) );
 a7862a <=( (not A199)  and  a7861a );
 a7863a <=( a7862a  and  a7857a );
 a7867a <=( A235  and  (not A233) );
 a7868a <=( (not A232)  and  a7867a );
 a7872a <=( A267  and  A266 );
 a7873a <=( (not A236)  and  a7872a );
 a7874a <=( a7873a  and  a7868a );
 a7877a <=( A168  and  A170 );
 a7881a <=( (not A199)  and  A166 );
 a7882a <=( (not A167)  and  a7881a );
 a7883a <=( a7882a  and  a7877a );
 a7887a <=( A232  and  (not A202) );
 a7888a <=( (not A200)  and  a7887a );
 a7892a <=( A300  and  A299 );
 a7893a <=( A234  and  a7892a );
 a7894a <=( a7893a  and  a7888a );
 a7897a <=( A168  and  A170 );
 a7901a <=( (not A199)  and  A166 );
 a7902a <=( (not A167)  and  a7901a );
 a7903a <=( a7902a  and  a7897a );
 a7907a <=( A232  and  (not A202) );
 a7908a <=( (not A200)  and  a7907a );
 a7912a <=( A300  and  A298 );
 a7913a <=( A234  and  a7912a );
 a7914a <=( a7913a  and  a7908a );
 a7917a <=( A168  and  A170 );
 a7921a <=( (not A199)  and  A166 );
 a7922a <=( (not A167)  and  a7921a );
 a7923a <=( a7922a  and  a7917a );
 a7927a <=( A232  and  (not A202) );
 a7928a <=( (not A200)  and  a7927a );
 a7932a <=( A267  and  A265 );
 a7933a <=( A234  and  a7932a );
 a7934a <=( a7933a  and  a7928a );
 a7937a <=( A168  and  A170 );
 a7941a <=( (not A199)  and  A166 );
 a7942a <=( (not A167)  and  a7941a );
 a7943a <=( a7942a  and  a7937a );
 a7947a <=( A232  and  (not A202) );
 a7948a <=( (not A200)  and  a7947a );
 a7952a <=( A267  and  A266 );
 a7953a <=( A234  and  a7952a );
 a7954a <=( a7953a  and  a7948a );
 a7957a <=( A168  and  A170 );
 a7961a <=( (not A199)  and  A166 );
 a7962a <=( (not A167)  and  a7961a );
 a7963a <=( a7962a  and  a7957a );
 a7967a <=( A233  and  (not A202) );
 a7968a <=( (not A200)  and  a7967a );
 a7972a <=( A300  and  A299 );
 a7973a <=( A234  and  a7972a );
 a7974a <=( a7973a  and  a7968a );
 a7977a <=( A168  and  A170 );
 a7981a <=( (not A199)  and  A166 );
 a7982a <=( (not A167)  and  a7981a );
 a7983a <=( a7982a  and  a7977a );
 a7987a <=( A233  and  (not A202) );
 a7988a <=( (not A200)  and  a7987a );
 a7992a <=( A300  and  A298 );
 a7993a <=( A234  and  a7992a );
 a7994a <=( a7993a  and  a7988a );
 a7997a <=( A168  and  A170 );
 a8001a <=( (not A199)  and  A166 );
 a8002a <=( (not A167)  and  a8001a );
 a8003a <=( a8002a  and  a7997a );
 a8007a <=( A233  and  (not A202) );
 a8008a <=( (not A200)  and  a8007a );
 a8012a <=( A267  and  A265 );
 a8013a <=( A234  and  a8012a );
 a8014a <=( a8013a  and  a8008a );
 a8017a <=( A168  and  A170 );
 a8021a <=( (not A199)  and  A166 );
 a8022a <=( (not A167)  and  a8021a );
 a8023a <=( a8022a  and  a8017a );
 a8027a <=( A233  and  (not A202) );
 a8028a <=( (not A200)  and  a8027a );
 a8032a <=( A267  and  A266 );
 a8033a <=( A234  and  a8032a );
 a8034a <=( a8033a  and  a8028a );
 a8037a <=( A168  and  A170 );
 a8041a <=( (not A199)  and  A166 );
 a8042a <=( (not A167)  and  a8041a );
 a8043a <=( a8042a  and  a8037a );
 a8047a <=( A232  and  A203 );
 a8048a <=( (not A200)  and  a8047a );
 a8052a <=( A300  and  A299 );
 a8053a <=( A234  and  a8052a );
 a8054a <=( a8053a  and  a8048a );
 a8057a <=( A168  and  A170 );
 a8061a <=( (not A199)  and  A166 );
 a8062a <=( (not A167)  and  a8061a );
 a8063a <=( a8062a  and  a8057a );
 a8067a <=( A232  and  A203 );
 a8068a <=( (not A200)  and  a8067a );
 a8072a <=( A300  and  A298 );
 a8073a <=( A234  and  a8072a );
 a8074a <=( a8073a  and  a8068a );
 a8077a <=( A168  and  A170 );
 a8081a <=( (not A199)  and  A166 );
 a8082a <=( (not A167)  and  a8081a );
 a8083a <=( a8082a  and  a8077a );
 a8087a <=( A232  and  A203 );
 a8088a <=( (not A200)  and  a8087a );
 a8092a <=( A267  and  A265 );
 a8093a <=( A234  and  a8092a );
 a8094a <=( a8093a  and  a8088a );
 a8097a <=( A168  and  A170 );
 a8101a <=( (not A199)  and  A166 );
 a8102a <=( (not A167)  and  a8101a );
 a8103a <=( a8102a  and  a8097a );
 a8107a <=( A232  and  A203 );
 a8108a <=( (not A200)  and  a8107a );
 a8112a <=( A267  and  A266 );
 a8113a <=( A234  and  a8112a );
 a8114a <=( a8113a  and  a8108a );
 a8117a <=( A168  and  A170 );
 a8121a <=( (not A199)  and  A166 );
 a8122a <=( (not A167)  and  a8121a );
 a8123a <=( a8122a  and  a8117a );
 a8127a <=( A233  and  A203 );
 a8128a <=( (not A200)  and  a8127a );
 a8132a <=( A300  and  A299 );
 a8133a <=( A234  and  a8132a );
 a8134a <=( a8133a  and  a8128a );
 a8137a <=( A168  and  A170 );
 a8141a <=( (not A199)  and  A166 );
 a8142a <=( (not A167)  and  a8141a );
 a8143a <=( a8142a  and  a8137a );
 a8147a <=( A233  and  A203 );
 a8148a <=( (not A200)  and  a8147a );
 a8152a <=( A300  and  A298 );
 a8153a <=( A234  and  a8152a );
 a8154a <=( a8153a  and  a8148a );
 a8157a <=( A168  and  A170 );
 a8161a <=( (not A199)  and  A166 );
 a8162a <=( (not A167)  and  a8161a );
 a8163a <=( a8162a  and  a8157a );
 a8167a <=( A233  and  A203 );
 a8168a <=( (not A200)  and  a8167a );
 a8172a <=( A267  and  A265 );
 a8173a <=( A234  and  a8172a );
 a8174a <=( a8173a  and  a8168a );
 a8177a <=( A168  and  A170 );
 a8181a <=( (not A199)  and  A166 );
 a8182a <=( (not A167)  and  a8181a );
 a8183a <=( a8182a  and  a8177a );
 a8187a <=( A233  and  A203 );
 a8188a <=( (not A200)  and  a8187a );
 a8192a <=( A267  and  A266 );
 a8193a <=( A234  and  a8192a );
 a8194a <=( a8193a  and  a8188a );
 a8197a <=( A168  and  A169 );
 a8201a <=( (not A199)  and  A166 );
 a8202a <=( (not A167)  and  a8201a );
 a8203a <=( a8202a  and  a8197a );
 a8207a <=( A232  and  (not A202) );
 a8208a <=( (not A200)  and  a8207a );
 a8212a <=( A300  and  A299 );
 a8213a <=( A234  and  a8212a );
 a8214a <=( a8213a  and  a8208a );
 a8217a <=( A168  and  A169 );
 a8221a <=( (not A199)  and  A166 );
 a8222a <=( (not A167)  and  a8221a );
 a8223a <=( a8222a  and  a8217a );
 a8227a <=( A232  and  (not A202) );
 a8228a <=( (not A200)  and  a8227a );
 a8232a <=( A300  and  A298 );
 a8233a <=( A234  and  a8232a );
 a8234a <=( a8233a  and  a8228a );
 a8237a <=( A168  and  A169 );
 a8241a <=( (not A199)  and  A166 );
 a8242a <=( (not A167)  and  a8241a );
 a8243a <=( a8242a  and  a8237a );
 a8247a <=( A232  and  (not A202) );
 a8248a <=( (not A200)  and  a8247a );
 a8252a <=( A267  and  A265 );
 a8253a <=( A234  and  a8252a );
 a8254a <=( a8253a  and  a8248a );
 a8257a <=( A168  and  A169 );
 a8261a <=( (not A199)  and  A166 );
 a8262a <=( (not A167)  and  a8261a );
 a8263a <=( a8262a  and  a8257a );
 a8267a <=( A232  and  (not A202) );
 a8268a <=( (not A200)  and  a8267a );
 a8272a <=( A267  and  A266 );
 a8273a <=( A234  and  a8272a );
 a8274a <=( a8273a  and  a8268a );
 a8277a <=( A168  and  A169 );
 a8281a <=( (not A199)  and  A166 );
 a8282a <=( (not A167)  and  a8281a );
 a8283a <=( a8282a  and  a8277a );
 a8287a <=( A233  and  (not A202) );
 a8288a <=( (not A200)  and  a8287a );
 a8292a <=( A300  and  A299 );
 a8293a <=( A234  and  a8292a );
 a8294a <=( a8293a  and  a8288a );
 a8297a <=( A168  and  A169 );
 a8301a <=( (not A199)  and  A166 );
 a8302a <=( (not A167)  and  a8301a );
 a8303a <=( a8302a  and  a8297a );
 a8307a <=( A233  and  (not A202) );
 a8308a <=( (not A200)  and  a8307a );
 a8312a <=( A300  and  A298 );
 a8313a <=( A234  and  a8312a );
 a8314a <=( a8313a  and  a8308a );
 a8317a <=( A168  and  A169 );
 a8321a <=( (not A199)  and  A166 );
 a8322a <=( (not A167)  and  a8321a );
 a8323a <=( a8322a  and  a8317a );
 a8327a <=( A233  and  (not A202) );
 a8328a <=( (not A200)  and  a8327a );
 a8332a <=( A267  and  A265 );
 a8333a <=( A234  and  a8332a );
 a8334a <=( a8333a  and  a8328a );
 a8337a <=( A168  and  A169 );
 a8341a <=( (not A199)  and  A166 );
 a8342a <=( (not A167)  and  a8341a );
 a8343a <=( a8342a  and  a8337a );
 a8347a <=( A233  and  (not A202) );
 a8348a <=( (not A200)  and  a8347a );
 a8352a <=( A267  and  A266 );
 a8353a <=( A234  and  a8352a );
 a8354a <=( a8353a  and  a8348a );
 a8357a <=( A168  and  A169 );
 a8361a <=( (not A199)  and  A166 );
 a8362a <=( (not A167)  and  a8361a );
 a8363a <=( a8362a  and  a8357a );
 a8367a <=( A232  and  A203 );
 a8368a <=( (not A200)  and  a8367a );
 a8372a <=( A300  and  A299 );
 a8373a <=( A234  and  a8372a );
 a8374a <=( a8373a  and  a8368a );
 a8377a <=( A168  and  A169 );
 a8381a <=( (not A199)  and  A166 );
 a8382a <=( (not A167)  and  a8381a );
 a8383a <=( a8382a  and  a8377a );
 a8387a <=( A232  and  A203 );
 a8388a <=( (not A200)  and  a8387a );
 a8392a <=( A300  and  A298 );
 a8393a <=( A234  and  a8392a );
 a8394a <=( a8393a  and  a8388a );
 a8397a <=( A168  and  A169 );
 a8401a <=( (not A199)  and  A166 );
 a8402a <=( (not A167)  and  a8401a );
 a8403a <=( a8402a  and  a8397a );
 a8407a <=( A232  and  A203 );
 a8408a <=( (not A200)  and  a8407a );
 a8412a <=( A267  and  A265 );
 a8413a <=( A234  and  a8412a );
 a8414a <=( a8413a  and  a8408a );
 a8417a <=( A168  and  A169 );
 a8421a <=( (not A199)  and  A166 );
 a8422a <=( (not A167)  and  a8421a );
 a8423a <=( a8422a  and  a8417a );
 a8427a <=( A232  and  A203 );
 a8428a <=( (not A200)  and  a8427a );
 a8432a <=( A267  and  A266 );
 a8433a <=( A234  and  a8432a );
 a8434a <=( a8433a  and  a8428a );
 a8437a <=( A168  and  A169 );
 a8441a <=( (not A199)  and  A166 );
 a8442a <=( (not A167)  and  a8441a );
 a8443a <=( a8442a  and  a8437a );
 a8447a <=( A233  and  A203 );
 a8448a <=( (not A200)  and  a8447a );
 a8452a <=( A300  and  A299 );
 a8453a <=( A234  and  a8452a );
 a8454a <=( a8453a  and  a8448a );
 a8457a <=( A168  and  A169 );
 a8461a <=( (not A199)  and  A166 );
 a8462a <=( (not A167)  and  a8461a );
 a8463a <=( a8462a  and  a8457a );
 a8467a <=( A233  and  A203 );
 a8468a <=( (not A200)  and  a8467a );
 a8472a <=( A300  and  A298 );
 a8473a <=( A234  and  a8472a );
 a8474a <=( a8473a  and  a8468a );
 a8477a <=( A168  and  A169 );
 a8481a <=( (not A199)  and  A166 );
 a8482a <=( (not A167)  and  a8481a );
 a8483a <=( a8482a  and  a8477a );
 a8487a <=( A233  and  A203 );
 a8488a <=( (not A200)  and  a8487a );
 a8492a <=( A267  and  A265 );
 a8493a <=( A234  and  a8492a );
 a8494a <=( a8493a  and  a8488a );
 a8497a <=( A168  and  A169 );
 a8501a <=( (not A199)  and  A166 );
 a8502a <=( (not A167)  and  a8501a );
 a8503a <=( a8502a  and  a8497a );
 a8507a <=( A233  and  A203 );
 a8508a <=( (not A200)  and  a8507a );
 a8512a <=( A267  and  A266 );
 a8513a <=( A234  and  a8512a );
 a8514a <=( a8513a  and  a8508a );
 a8518a <=( A199  and  (not A166) );
 a8519a <=( A167  and  a8518a );
 a8523a <=( (not A202)  and  (not A201) );
 a8524a <=( A200  and  a8523a );
 a8525a <=( a8524a  and  a8519a );
 a8529a <=( A298  and  A234 );
 a8530a <=( A232  and  a8529a );
 a8534a <=( (not A302)  and  A301 );
 a8535a <=( A299  and  a8534a );
 a8536a <=( a8535a  and  a8530a );
 a8540a <=( A199  and  (not A166) );
 a8541a <=( A167  and  a8540a );
 a8545a <=( (not A202)  and  (not A201) );
 a8546a <=( A200  and  a8545a );
 a8547a <=( a8546a  and  a8541a );
 a8551a <=( A298  and  A234 );
 a8552a <=( A232  and  a8551a );
 a8556a <=( A302  and  (not A301) );
 a8557a <=( (not A299)  and  a8556a );
 a8558a <=( a8557a  and  a8552a );
 a8562a <=( A199  and  (not A166) );
 a8563a <=( A167  and  a8562a );
 a8567a <=( (not A202)  and  (not A201) );
 a8568a <=( A200  and  a8567a );
 a8569a <=( a8568a  and  a8563a );
 a8573a <=( (not A298)  and  A234 );
 a8574a <=( A232  and  a8573a );
 a8578a <=( A302  and  (not A301) );
 a8579a <=( A299  and  a8578a );
 a8580a <=( a8579a  and  a8574a );
 a8584a <=( A199  and  (not A166) );
 a8585a <=( A167  and  a8584a );
 a8589a <=( (not A202)  and  (not A201) );
 a8590a <=( A200  and  a8589a );
 a8591a <=( a8590a  and  a8585a );
 a8595a <=( (not A298)  and  A234 );
 a8596a <=( A232  and  a8595a );
 a8600a <=( (not A302)  and  A301 );
 a8601a <=( (not A299)  and  a8600a );
 a8602a <=( a8601a  and  a8596a );
 a8606a <=( A199  and  (not A166) );
 a8607a <=( A167  and  a8606a );
 a8611a <=( (not A202)  and  (not A201) );
 a8612a <=( A200  and  a8611a );
 a8613a <=( a8612a  and  a8607a );
 a8617a <=( A265  and  A234 );
 a8618a <=( A232  and  a8617a );
 a8622a <=( (not A269)  and  A268 );
 a8623a <=( A266  and  a8622a );
 a8624a <=( a8623a  and  a8618a );
 a8628a <=( A199  and  (not A166) );
 a8629a <=( A167  and  a8628a );
 a8633a <=( (not A202)  and  (not A201) );
 a8634a <=( A200  and  a8633a );
 a8635a <=( a8634a  and  a8629a );
 a8639a <=( (not A265)  and  A234 );
 a8640a <=( A232  and  a8639a );
 a8644a <=( A269  and  (not A268) );
 a8645a <=( A266  and  a8644a );
 a8646a <=( a8645a  and  a8640a );
 a8650a <=( A199  and  (not A166) );
 a8651a <=( A167  and  a8650a );
 a8655a <=( (not A202)  and  (not A201) );
 a8656a <=( A200  and  a8655a );
 a8657a <=( a8656a  and  a8651a );
 a8661a <=( A265  and  A234 );
 a8662a <=( A232  and  a8661a );
 a8666a <=( A269  and  (not A268) );
 a8667a <=( (not A266)  and  a8666a );
 a8668a <=( a8667a  and  a8662a );
 a8672a <=( A199  and  (not A166) );
 a8673a <=( A167  and  a8672a );
 a8677a <=( (not A202)  and  (not A201) );
 a8678a <=( A200  and  a8677a );
 a8679a <=( a8678a  and  a8673a );
 a8683a <=( (not A265)  and  A234 );
 a8684a <=( A232  and  a8683a );
 a8688a <=( (not A269)  and  A268 );
 a8689a <=( (not A266)  and  a8688a );
 a8690a <=( a8689a  and  a8684a );
 a8694a <=( A199  and  (not A166) );
 a8695a <=( A167  and  a8694a );
 a8699a <=( (not A202)  and  (not A201) );
 a8700a <=( A200  and  a8699a );
 a8701a <=( a8700a  and  a8695a );
 a8705a <=( A298  and  A234 );
 a8706a <=( A233  and  a8705a );
 a8710a <=( (not A302)  and  A301 );
 a8711a <=( A299  and  a8710a );
 a8712a <=( a8711a  and  a8706a );
 a8716a <=( A199  and  (not A166) );
 a8717a <=( A167  and  a8716a );
 a8721a <=( (not A202)  and  (not A201) );
 a8722a <=( A200  and  a8721a );
 a8723a <=( a8722a  and  a8717a );
 a8727a <=( A298  and  A234 );
 a8728a <=( A233  and  a8727a );
 a8732a <=( A302  and  (not A301) );
 a8733a <=( (not A299)  and  a8732a );
 a8734a <=( a8733a  and  a8728a );
 a8738a <=( A199  and  (not A166) );
 a8739a <=( A167  and  a8738a );
 a8743a <=( (not A202)  and  (not A201) );
 a8744a <=( A200  and  a8743a );
 a8745a <=( a8744a  and  a8739a );
 a8749a <=( (not A298)  and  A234 );
 a8750a <=( A233  and  a8749a );
 a8754a <=( A302  and  (not A301) );
 a8755a <=( A299  and  a8754a );
 a8756a <=( a8755a  and  a8750a );
 a8760a <=( A199  and  (not A166) );
 a8761a <=( A167  and  a8760a );
 a8765a <=( (not A202)  and  (not A201) );
 a8766a <=( A200  and  a8765a );
 a8767a <=( a8766a  and  a8761a );
 a8771a <=( (not A298)  and  A234 );
 a8772a <=( A233  and  a8771a );
 a8776a <=( (not A302)  and  A301 );
 a8777a <=( (not A299)  and  a8776a );
 a8778a <=( a8777a  and  a8772a );
 a8782a <=( A199  and  (not A166) );
 a8783a <=( A167  and  a8782a );
 a8787a <=( (not A202)  and  (not A201) );
 a8788a <=( A200  and  a8787a );
 a8789a <=( a8788a  and  a8783a );
 a8793a <=( A265  and  A234 );
 a8794a <=( A233  and  a8793a );
 a8798a <=( (not A269)  and  A268 );
 a8799a <=( A266  and  a8798a );
 a8800a <=( a8799a  and  a8794a );
 a8804a <=( A199  and  (not A166) );
 a8805a <=( A167  and  a8804a );
 a8809a <=( (not A202)  and  (not A201) );
 a8810a <=( A200  and  a8809a );
 a8811a <=( a8810a  and  a8805a );
 a8815a <=( (not A265)  and  A234 );
 a8816a <=( A233  and  a8815a );
 a8820a <=( A269  and  (not A268) );
 a8821a <=( A266  and  a8820a );
 a8822a <=( a8821a  and  a8816a );
 a8826a <=( A199  and  (not A166) );
 a8827a <=( A167  and  a8826a );
 a8831a <=( (not A202)  and  (not A201) );
 a8832a <=( A200  and  a8831a );
 a8833a <=( a8832a  and  a8827a );
 a8837a <=( A265  and  A234 );
 a8838a <=( A233  and  a8837a );
 a8842a <=( A269  and  (not A268) );
 a8843a <=( (not A266)  and  a8842a );
 a8844a <=( a8843a  and  a8838a );
 a8848a <=( A199  and  (not A166) );
 a8849a <=( A167  and  a8848a );
 a8853a <=( (not A202)  and  (not A201) );
 a8854a <=( A200  and  a8853a );
 a8855a <=( a8854a  and  a8849a );
 a8859a <=( (not A265)  and  A234 );
 a8860a <=( A233  and  a8859a );
 a8864a <=( (not A269)  and  A268 );
 a8865a <=( (not A266)  and  a8864a );
 a8866a <=( a8865a  and  a8860a );
 a8870a <=( A199  and  (not A166) );
 a8871a <=( A167  and  a8870a );
 a8875a <=( (not A202)  and  (not A201) );
 a8876a <=( A200  and  a8875a );
 a8877a <=( a8876a  and  a8871a );
 a8881a <=( A235  and  A233 );
 a8882a <=( A232  and  a8881a );
 a8886a <=( A300  and  A299 );
 a8887a <=( (not A236)  and  a8886a );
 a8888a <=( a8887a  and  a8882a );
 a8892a <=( A199  and  (not A166) );
 a8893a <=( A167  and  a8892a );
 a8897a <=( (not A202)  and  (not A201) );
 a8898a <=( A200  and  a8897a );
 a8899a <=( a8898a  and  a8893a );
 a8903a <=( A235  and  A233 );
 a8904a <=( A232  and  a8903a );
 a8908a <=( A300  and  A298 );
 a8909a <=( (not A236)  and  a8908a );
 a8910a <=( a8909a  and  a8904a );
 a8914a <=( A199  and  (not A166) );
 a8915a <=( A167  and  a8914a );
 a8919a <=( (not A202)  and  (not A201) );
 a8920a <=( A200  and  a8919a );
 a8921a <=( a8920a  and  a8915a );
 a8925a <=( A235  and  A233 );
 a8926a <=( A232  and  a8925a );
 a8930a <=( A267  and  A265 );
 a8931a <=( (not A236)  and  a8930a );
 a8932a <=( a8931a  and  a8926a );
 a8936a <=( A199  and  (not A166) );
 a8937a <=( A167  and  a8936a );
 a8941a <=( (not A202)  and  (not A201) );
 a8942a <=( A200  and  a8941a );
 a8943a <=( a8942a  and  a8937a );
 a8947a <=( A235  and  A233 );
 a8948a <=( A232  and  a8947a );
 a8952a <=( A267  and  A266 );
 a8953a <=( (not A236)  and  a8952a );
 a8954a <=( a8953a  and  a8948a );
 a8958a <=( A199  and  (not A166) );
 a8959a <=( A167  and  a8958a );
 a8963a <=( (not A202)  and  (not A201) );
 a8964a <=( A200  and  a8963a );
 a8965a <=( a8964a  and  a8959a );
 a8969a <=( (not A235)  and  A233 );
 a8970a <=( (not A232)  and  a8969a );
 a8974a <=( A300  and  A299 );
 a8975a <=( A236  and  a8974a );
 a8976a <=( a8975a  and  a8970a );
 a8980a <=( A199  and  (not A166) );
 a8981a <=( A167  and  a8980a );
 a8985a <=( (not A202)  and  (not A201) );
 a8986a <=( A200  and  a8985a );
 a8987a <=( a8986a  and  a8981a );
 a8991a <=( (not A235)  and  A233 );
 a8992a <=( (not A232)  and  a8991a );
 a8996a <=( A300  and  A298 );
 a8997a <=( A236  and  a8996a );
 a8998a <=( a8997a  and  a8992a );
 a9002a <=( A199  and  (not A166) );
 a9003a <=( A167  and  a9002a );
 a9007a <=( (not A202)  and  (not A201) );
 a9008a <=( A200  and  a9007a );
 a9009a <=( a9008a  and  a9003a );
 a9013a <=( (not A235)  and  A233 );
 a9014a <=( (not A232)  and  a9013a );
 a9018a <=( A267  and  A265 );
 a9019a <=( A236  and  a9018a );
 a9020a <=( a9019a  and  a9014a );
 a9024a <=( A199  and  (not A166) );
 a9025a <=( A167  and  a9024a );
 a9029a <=( (not A202)  and  (not A201) );
 a9030a <=( A200  and  a9029a );
 a9031a <=( a9030a  and  a9025a );
 a9035a <=( (not A235)  and  A233 );
 a9036a <=( (not A232)  and  a9035a );
 a9040a <=( A267  and  A266 );
 a9041a <=( A236  and  a9040a );
 a9042a <=( a9041a  and  a9036a );
 a9046a <=( A199  and  (not A166) );
 a9047a <=( A167  and  a9046a );
 a9051a <=( (not A202)  and  (not A201) );
 a9052a <=( A200  and  a9051a );
 a9053a <=( a9052a  and  a9047a );
 a9057a <=( (not A235)  and  (not A233) );
 a9058a <=( A232  and  a9057a );
 a9062a <=( A300  and  A299 );
 a9063a <=( A236  and  a9062a );
 a9064a <=( a9063a  and  a9058a );
 a9068a <=( A199  and  (not A166) );
 a9069a <=( A167  and  a9068a );
 a9073a <=( (not A202)  and  (not A201) );
 a9074a <=( A200  and  a9073a );
 a9075a <=( a9074a  and  a9069a );
 a9079a <=( (not A235)  and  (not A233) );
 a9080a <=( A232  and  a9079a );
 a9084a <=( A300  and  A298 );
 a9085a <=( A236  and  a9084a );
 a9086a <=( a9085a  and  a9080a );
 a9090a <=( A199  and  (not A166) );
 a9091a <=( A167  and  a9090a );
 a9095a <=( (not A202)  and  (not A201) );
 a9096a <=( A200  and  a9095a );
 a9097a <=( a9096a  and  a9091a );
 a9101a <=( (not A235)  and  (not A233) );
 a9102a <=( A232  and  a9101a );
 a9106a <=( A267  and  A265 );
 a9107a <=( A236  and  a9106a );
 a9108a <=( a9107a  and  a9102a );
 a9112a <=( A199  and  (not A166) );
 a9113a <=( A167  and  a9112a );
 a9117a <=( (not A202)  and  (not A201) );
 a9118a <=( A200  and  a9117a );
 a9119a <=( a9118a  and  a9113a );
 a9123a <=( (not A235)  and  (not A233) );
 a9124a <=( A232  and  a9123a );
 a9128a <=( A267  and  A266 );
 a9129a <=( A236  and  a9128a );
 a9130a <=( a9129a  and  a9124a );
 a9134a <=( A199  and  (not A166) );
 a9135a <=( A167  and  a9134a );
 a9139a <=( (not A202)  and  (not A201) );
 a9140a <=( A200  and  a9139a );
 a9141a <=( a9140a  and  a9135a );
 a9145a <=( A235  and  (not A233) );
 a9146a <=( (not A232)  and  a9145a );
 a9150a <=( A300  and  A299 );
 a9151a <=( (not A236)  and  a9150a );
 a9152a <=( a9151a  and  a9146a );
 a9156a <=( A199  and  (not A166) );
 a9157a <=( A167  and  a9156a );
 a9161a <=( (not A202)  and  (not A201) );
 a9162a <=( A200  and  a9161a );
 a9163a <=( a9162a  and  a9157a );
 a9167a <=( A235  and  (not A233) );
 a9168a <=( (not A232)  and  a9167a );
 a9172a <=( A300  and  A298 );
 a9173a <=( (not A236)  and  a9172a );
 a9174a <=( a9173a  and  a9168a );
 a9178a <=( A199  and  (not A166) );
 a9179a <=( A167  and  a9178a );
 a9183a <=( (not A202)  and  (not A201) );
 a9184a <=( A200  and  a9183a );
 a9185a <=( a9184a  and  a9179a );
 a9189a <=( A235  and  (not A233) );
 a9190a <=( (not A232)  and  a9189a );
 a9194a <=( A267  and  A265 );
 a9195a <=( (not A236)  and  a9194a );
 a9196a <=( a9195a  and  a9190a );
 a9200a <=( A199  and  (not A166) );
 a9201a <=( A167  and  a9200a );
 a9205a <=( (not A202)  and  (not A201) );
 a9206a <=( A200  and  a9205a );
 a9207a <=( a9206a  and  a9201a );
 a9211a <=( A235  and  (not A233) );
 a9212a <=( (not A232)  and  a9211a );
 a9216a <=( A267  and  A266 );
 a9217a <=( (not A236)  and  a9216a );
 a9218a <=( a9217a  and  a9212a );
 a9222a <=( A199  and  (not A166) );
 a9223a <=( A167  and  a9222a );
 a9227a <=( A203  and  (not A201) );
 a9228a <=( A200  and  a9227a );
 a9229a <=( a9228a  and  a9223a );
 a9233a <=( A298  and  A234 );
 a9234a <=( A232  and  a9233a );
 a9238a <=( (not A302)  and  A301 );
 a9239a <=( A299  and  a9238a );
 a9240a <=( a9239a  and  a9234a );
 a9244a <=( A199  and  (not A166) );
 a9245a <=( A167  and  a9244a );
 a9249a <=( A203  and  (not A201) );
 a9250a <=( A200  and  a9249a );
 a9251a <=( a9250a  and  a9245a );
 a9255a <=( A298  and  A234 );
 a9256a <=( A232  and  a9255a );
 a9260a <=( A302  and  (not A301) );
 a9261a <=( (not A299)  and  a9260a );
 a9262a <=( a9261a  and  a9256a );
 a9266a <=( A199  and  (not A166) );
 a9267a <=( A167  and  a9266a );
 a9271a <=( A203  and  (not A201) );
 a9272a <=( A200  and  a9271a );
 a9273a <=( a9272a  and  a9267a );
 a9277a <=( (not A298)  and  A234 );
 a9278a <=( A232  and  a9277a );
 a9282a <=( A302  and  (not A301) );
 a9283a <=( A299  and  a9282a );
 a9284a <=( a9283a  and  a9278a );
 a9288a <=( A199  and  (not A166) );
 a9289a <=( A167  and  a9288a );
 a9293a <=( A203  and  (not A201) );
 a9294a <=( A200  and  a9293a );
 a9295a <=( a9294a  and  a9289a );
 a9299a <=( (not A298)  and  A234 );
 a9300a <=( A232  and  a9299a );
 a9304a <=( (not A302)  and  A301 );
 a9305a <=( (not A299)  and  a9304a );
 a9306a <=( a9305a  and  a9300a );
 a9310a <=( A199  and  (not A166) );
 a9311a <=( A167  and  a9310a );
 a9315a <=( A203  and  (not A201) );
 a9316a <=( A200  and  a9315a );
 a9317a <=( a9316a  and  a9311a );
 a9321a <=( A265  and  A234 );
 a9322a <=( A232  and  a9321a );
 a9326a <=( (not A269)  and  A268 );
 a9327a <=( A266  and  a9326a );
 a9328a <=( a9327a  and  a9322a );
 a9332a <=( A199  and  (not A166) );
 a9333a <=( A167  and  a9332a );
 a9337a <=( A203  and  (not A201) );
 a9338a <=( A200  and  a9337a );
 a9339a <=( a9338a  and  a9333a );
 a9343a <=( (not A265)  and  A234 );
 a9344a <=( A232  and  a9343a );
 a9348a <=( A269  and  (not A268) );
 a9349a <=( A266  and  a9348a );
 a9350a <=( a9349a  and  a9344a );
 a9354a <=( A199  and  (not A166) );
 a9355a <=( A167  and  a9354a );
 a9359a <=( A203  and  (not A201) );
 a9360a <=( A200  and  a9359a );
 a9361a <=( a9360a  and  a9355a );
 a9365a <=( A265  and  A234 );
 a9366a <=( A232  and  a9365a );
 a9370a <=( A269  and  (not A268) );
 a9371a <=( (not A266)  and  a9370a );
 a9372a <=( a9371a  and  a9366a );
 a9376a <=( A199  and  (not A166) );
 a9377a <=( A167  and  a9376a );
 a9381a <=( A203  and  (not A201) );
 a9382a <=( A200  and  a9381a );
 a9383a <=( a9382a  and  a9377a );
 a9387a <=( (not A265)  and  A234 );
 a9388a <=( A232  and  a9387a );
 a9392a <=( (not A269)  and  A268 );
 a9393a <=( (not A266)  and  a9392a );
 a9394a <=( a9393a  and  a9388a );
 a9398a <=( A199  and  (not A166) );
 a9399a <=( A167  and  a9398a );
 a9403a <=( A203  and  (not A201) );
 a9404a <=( A200  and  a9403a );
 a9405a <=( a9404a  and  a9399a );
 a9409a <=( A298  and  A234 );
 a9410a <=( A233  and  a9409a );
 a9414a <=( (not A302)  and  A301 );
 a9415a <=( A299  and  a9414a );
 a9416a <=( a9415a  and  a9410a );
 a9420a <=( A199  and  (not A166) );
 a9421a <=( A167  and  a9420a );
 a9425a <=( A203  and  (not A201) );
 a9426a <=( A200  and  a9425a );
 a9427a <=( a9426a  and  a9421a );
 a9431a <=( A298  and  A234 );
 a9432a <=( A233  and  a9431a );
 a9436a <=( A302  and  (not A301) );
 a9437a <=( (not A299)  and  a9436a );
 a9438a <=( a9437a  and  a9432a );
 a9442a <=( A199  and  (not A166) );
 a9443a <=( A167  and  a9442a );
 a9447a <=( A203  and  (not A201) );
 a9448a <=( A200  and  a9447a );
 a9449a <=( a9448a  and  a9443a );
 a9453a <=( (not A298)  and  A234 );
 a9454a <=( A233  and  a9453a );
 a9458a <=( A302  and  (not A301) );
 a9459a <=( A299  and  a9458a );
 a9460a <=( a9459a  and  a9454a );
 a9464a <=( A199  and  (not A166) );
 a9465a <=( A167  and  a9464a );
 a9469a <=( A203  and  (not A201) );
 a9470a <=( A200  and  a9469a );
 a9471a <=( a9470a  and  a9465a );
 a9475a <=( (not A298)  and  A234 );
 a9476a <=( A233  and  a9475a );
 a9480a <=( (not A302)  and  A301 );
 a9481a <=( (not A299)  and  a9480a );
 a9482a <=( a9481a  and  a9476a );
 a9486a <=( A199  and  (not A166) );
 a9487a <=( A167  and  a9486a );
 a9491a <=( A203  and  (not A201) );
 a9492a <=( A200  and  a9491a );
 a9493a <=( a9492a  and  a9487a );
 a9497a <=( A265  and  A234 );
 a9498a <=( A233  and  a9497a );
 a9502a <=( (not A269)  and  A268 );
 a9503a <=( A266  and  a9502a );
 a9504a <=( a9503a  and  a9498a );
 a9508a <=( A199  and  (not A166) );
 a9509a <=( A167  and  a9508a );
 a9513a <=( A203  and  (not A201) );
 a9514a <=( A200  and  a9513a );
 a9515a <=( a9514a  and  a9509a );
 a9519a <=( (not A265)  and  A234 );
 a9520a <=( A233  and  a9519a );
 a9524a <=( A269  and  (not A268) );
 a9525a <=( A266  and  a9524a );
 a9526a <=( a9525a  and  a9520a );
 a9530a <=( A199  and  (not A166) );
 a9531a <=( A167  and  a9530a );
 a9535a <=( A203  and  (not A201) );
 a9536a <=( A200  and  a9535a );
 a9537a <=( a9536a  and  a9531a );
 a9541a <=( A265  and  A234 );
 a9542a <=( A233  and  a9541a );
 a9546a <=( A269  and  (not A268) );
 a9547a <=( (not A266)  and  a9546a );
 a9548a <=( a9547a  and  a9542a );
 a9552a <=( A199  and  (not A166) );
 a9553a <=( A167  and  a9552a );
 a9557a <=( A203  and  (not A201) );
 a9558a <=( A200  and  a9557a );
 a9559a <=( a9558a  and  a9553a );
 a9563a <=( (not A265)  and  A234 );
 a9564a <=( A233  and  a9563a );
 a9568a <=( (not A269)  and  A268 );
 a9569a <=( (not A266)  and  a9568a );
 a9570a <=( a9569a  and  a9564a );
 a9574a <=( A199  and  (not A166) );
 a9575a <=( A167  and  a9574a );
 a9579a <=( A203  and  (not A201) );
 a9580a <=( A200  and  a9579a );
 a9581a <=( a9580a  and  a9575a );
 a9585a <=( A235  and  A233 );
 a9586a <=( A232  and  a9585a );
 a9590a <=( A300  and  A299 );
 a9591a <=( (not A236)  and  a9590a );
 a9592a <=( a9591a  and  a9586a );
 a9596a <=( A199  and  (not A166) );
 a9597a <=( A167  and  a9596a );
 a9601a <=( A203  and  (not A201) );
 a9602a <=( A200  and  a9601a );
 a9603a <=( a9602a  and  a9597a );
 a9607a <=( A235  and  A233 );
 a9608a <=( A232  and  a9607a );
 a9612a <=( A300  and  A298 );
 a9613a <=( (not A236)  and  a9612a );
 a9614a <=( a9613a  and  a9608a );
 a9618a <=( A199  and  (not A166) );
 a9619a <=( A167  and  a9618a );
 a9623a <=( A203  and  (not A201) );
 a9624a <=( A200  and  a9623a );
 a9625a <=( a9624a  and  a9619a );
 a9629a <=( A235  and  A233 );
 a9630a <=( A232  and  a9629a );
 a9634a <=( A267  and  A265 );
 a9635a <=( (not A236)  and  a9634a );
 a9636a <=( a9635a  and  a9630a );
 a9640a <=( A199  and  (not A166) );
 a9641a <=( A167  and  a9640a );
 a9645a <=( A203  and  (not A201) );
 a9646a <=( A200  and  a9645a );
 a9647a <=( a9646a  and  a9641a );
 a9651a <=( A235  and  A233 );
 a9652a <=( A232  and  a9651a );
 a9656a <=( A267  and  A266 );
 a9657a <=( (not A236)  and  a9656a );
 a9658a <=( a9657a  and  a9652a );
 a9662a <=( A199  and  (not A166) );
 a9663a <=( A167  and  a9662a );
 a9667a <=( A203  and  (not A201) );
 a9668a <=( A200  and  a9667a );
 a9669a <=( a9668a  and  a9663a );
 a9673a <=( (not A235)  and  A233 );
 a9674a <=( (not A232)  and  a9673a );
 a9678a <=( A300  and  A299 );
 a9679a <=( A236  and  a9678a );
 a9680a <=( a9679a  and  a9674a );
 a9684a <=( A199  and  (not A166) );
 a9685a <=( A167  and  a9684a );
 a9689a <=( A203  and  (not A201) );
 a9690a <=( A200  and  a9689a );
 a9691a <=( a9690a  and  a9685a );
 a9695a <=( (not A235)  and  A233 );
 a9696a <=( (not A232)  and  a9695a );
 a9700a <=( A300  and  A298 );
 a9701a <=( A236  and  a9700a );
 a9702a <=( a9701a  and  a9696a );
 a9706a <=( A199  and  (not A166) );
 a9707a <=( A167  and  a9706a );
 a9711a <=( A203  and  (not A201) );
 a9712a <=( A200  and  a9711a );
 a9713a <=( a9712a  and  a9707a );
 a9717a <=( (not A235)  and  A233 );
 a9718a <=( (not A232)  and  a9717a );
 a9722a <=( A267  and  A265 );
 a9723a <=( A236  and  a9722a );
 a9724a <=( a9723a  and  a9718a );
 a9728a <=( A199  and  (not A166) );
 a9729a <=( A167  and  a9728a );
 a9733a <=( A203  and  (not A201) );
 a9734a <=( A200  and  a9733a );
 a9735a <=( a9734a  and  a9729a );
 a9739a <=( (not A235)  and  A233 );
 a9740a <=( (not A232)  and  a9739a );
 a9744a <=( A267  and  A266 );
 a9745a <=( A236  and  a9744a );
 a9746a <=( a9745a  and  a9740a );
 a9750a <=( A199  and  (not A166) );
 a9751a <=( A167  and  a9750a );
 a9755a <=( A203  and  (not A201) );
 a9756a <=( A200  and  a9755a );
 a9757a <=( a9756a  and  a9751a );
 a9761a <=( (not A235)  and  (not A233) );
 a9762a <=( A232  and  a9761a );
 a9766a <=( A300  and  A299 );
 a9767a <=( A236  and  a9766a );
 a9768a <=( a9767a  and  a9762a );
 a9772a <=( A199  and  (not A166) );
 a9773a <=( A167  and  a9772a );
 a9777a <=( A203  and  (not A201) );
 a9778a <=( A200  and  a9777a );
 a9779a <=( a9778a  and  a9773a );
 a9783a <=( (not A235)  and  (not A233) );
 a9784a <=( A232  and  a9783a );
 a9788a <=( A300  and  A298 );
 a9789a <=( A236  and  a9788a );
 a9790a <=( a9789a  and  a9784a );
 a9794a <=( A199  and  (not A166) );
 a9795a <=( A167  and  a9794a );
 a9799a <=( A203  and  (not A201) );
 a9800a <=( A200  and  a9799a );
 a9801a <=( a9800a  and  a9795a );
 a9805a <=( (not A235)  and  (not A233) );
 a9806a <=( A232  and  a9805a );
 a9810a <=( A267  and  A265 );
 a9811a <=( A236  and  a9810a );
 a9812a <=( a9811a  and  a9806a );
 a9816a <=( A199  and  (not A166) );
 a9817a <=( A167  and  a9816a );
 a9821a <=( A203  and  (not A201) );
 a9822a <=( A200  and  a9821a );
 a9823a <=( a9822a  and  a9817a );
 a9827a <=( (not A235)  and  (not A233) );
 a9828a <=( A232  and  a9827a );
 a9832a <=( A267  and  A266 );
 a9833a <=( A236  and  a9832a );
 a9834a <=( a9833a  and  a9828a );
 a9838a <=( A199  and  (not A166) );
 a9839a <=( A167  and  a9838a );
 a9843a <=( A203  and  (not A201) );
 a9844a <=( A200  and  a9843a );
 a9845a <=( a9844a  and  a9839a );
 a9849a <=( A235  and  (not A233) );
 a9850a <=( (not A232)  and  a9849a );
 a9854a <=( A300  and  A299 );
 a9855a <=( (not A236)  and  a9854a );
 a9856a <=( a9855a  and  a9850a );
 a9860a <=( A199  and  (not A166) );
 a9861a <=( A167  and  a9860a );
 a9865a <=( A203  and  (not A201) );
 a9866a <=( A200  and  a9865a );
 a9867a <=( a9866a  and  a9861a );
 a9871a <=( A235  and  (not A233) );
 a9872a <=( (not A232)  and  a9871a );
 a9876a <=( A300  and  A298 );
 a9877a <=( (not A236)  and  a9876a );
 a9878a <=( a9877a  and  a9872a );
 a9882a <=( A199  and  (not A166) );
 a9883a <=( A167  and  a9882a );
 a9887a <=( A203  and  (not A201) );
 a9888a <=( A200  and  a9887a );
 a9889a <=( a9888a  and  a9883a );
 a9893a <=( A235  and  (not A233) );
 a9894a <=( (not A232)  and  a9893a );
 a9898a <=( A267  and  A265 );
 a9899a <=( (not A236)  and  a9898a );
 a9900a <=( a9899a  and  a9894a );
 a9904a <=( A199  and  (not A166) );
 a9905a <=( A167  and  a9904a );
 a9909a <=( A203  and  (not A201) );
 a9910a <=( A200  and  a9909a );
 a9911a <=( a9910a  and  a9905a );
 a9915a <=( A235  and  (not A233) );
 a9916a <=( (not A232)  and  a9915a );
 a9920a <=( A267  and  A266 );
 a9921a <=( (not A236)  and  a9920a );
 a9922a <=( a9921a  and  a9916a );
 a9926a <=( (not A199)  and  (not A166) );
 a9927a <=( A167  and  a9926a );
 a9931a <=( A202  and  (not A201) );
 a9932a <=( A200  and  a9931a );
 a9933a <=( a9932a  and  a9927a );
 a9937a <=( A298  and  A234 );
 a9938a <=( A232  and  a9937a );
 a9942a <=( (not A302)  and  A301 );
 a9943a <=( A299  and  a9942a );
 a9944a <=( a9943a  and  a9938a );
 a9948a <=( (not A199)  and  (not A166) );
 a9949a <=( A167  and  a9948a );
 a9953a <=( A202  and  (not A201) );
 a9954a <=( A200  and  a9953a );
 a9955a <=( a9954a  and  a9949a );
 a9959a <=( A298  and  A234 );
 a9960a <=( A232  and  a9959a );
 a9964a <=( A302  and  (not A301) );
 a9965a <=( (not A299)  and  a9964a );
 a9966a <=( a9965a  and  a9960a );
 a9970a <=( (not A199)  and  (not A166) );
 a9971a <=( A167  and  a9970a );
 a9975a <=( A202  and  (not A201) );
 a9976a <=( A200  and  a9975a );
 a9977a <=( a9976a  and  a9971a );
 a9981a <=( (not A298)  and  A234 );
 a9982a <=( A232  and  a9981a );
 a9986a <=( A302  and  (not A301) );
 a9987a <=( A299  and  a9986a );
 a9988a <=( a9987a  and  a9982a );
 a9992a <=( (not A199)  and  (not A166) );
 a9993a <=( A167  and  a9992a );
 a9997a <=( A202  and  (not A201) );
 a9998a <=( A200  and  a9997a );
 a9999a <=( a9998a  and  a9993a );
 a10003a <=( (not A298)  and  A234 );
 a10004a <=( A232  and  a10003a );
 a10008a <=( (not A302)  and  A301 );
 a10009a <=( (not A299)  and  a10008a );
 a10010a <=( a10009a  and  a10004a );
 a10014a <=( (not A199)  and  (not A166) );
 a10015a <=( A167  and  a10014a );
 a10019a <=( A202  and  (not A201) );
 a10020a <=( A200  and  a10019a );
 a10021a <=( a10020a  and  a10015a );
 a10025a <=( A265  and  A234 );
 a10026a <=( A232  and  a10025a );
 a10030a <=( (not A269)  and  A268 );
 a10031a <=( A266  and  a10030a );
 a10032a <=( a10031a  and  a10026a );
 a10036a <=( (not A199)  and  (not A166) );
 a10037a <=( A167  and  a10036a );
 a10041a <=( A202  and  (not A201) );
 a10042a <=( A200  and  a10041a );
 a10043a <=( a10042a  and  a10037a );
 a10047a <=( (not A265)  and  A234 );
 a10048a <=( A232  and  a10047a );
 a10052a <=( A269  and  (not A268) );
 a10053a <=( A266  and  a10052a );
 a10054a <=( a10053a  and  a10048a );
 a10058a <=( (not A199)  and  (not A166) );
 a10059a <=( A167  and  a10058a );
 a10063a <=( A202  and  (not A201) );
 a10064a <=( A200  and  a10063a );
 a10065a <=( a10064a  and  a10059a );
 a10069a <=( A265  and  A234 );
 a10070a <=( A232  and  a10069a );
 a10074a <=( A269  and  (not A268) );
 a10075a <=( (not A266)  and  a10074a );
 a10076a <=( a10075a  and  a10070a );
 a10080a <=( (not A199)  and  (not A166) );
 a10081a <=( A167  and  a10080a );
 a10085a <=( A202  and  (not A201) );
 a10086a <=( A200  and  a10085a );
 a10087a <=( a10086a  and  a10081a );
 a10091a <=( (not A265)  and  A234 );
 a10092a <=( A232  and  a10091a );
 a10096a <=( (not A269)  and  A268 );
 a10097a <=( (not A266)  and  a10096a );
 a10098a <=( a10097a  and  a10092a );
 a10102a <=( (not A199)  and  (not A166) );
 a10103a <=( A167  and  a10102a );
 a10107a <=( A202  and  (not A201) );
 a10108a <=( A200  and  a10107a );
 a10109a <=( a10108a  and  a10103a );
 a10113a <=( A298  and  A234 );
 a10114a <=( A233  and  a10113a );
 a10118a <=( (not A302)  and  A301 );
 a10119a <=( A299  and  a10118a );
 a10120a <=( a10119a  and  a10114a );
 a10124a <=( (not A199)  and  (not A166) );
 a10125a <=( A167  and  a10124a );
 a10129a <=( A202  and  (not A201) );
 a10130a <=( A200  and  a10129a );
 a10131a <=( a10130a  and  a10125a );
 a10135a <=( A298  and  A234 );
 a10136a <=( A233  and  a10135a );
 a10140a <=( A302  and  (not A301) );
 a10141a <=( (not A299)  and  a10140a );
 a10142a <=( a10141a  and  a10136a );
 a10146a <=( (not A199)  and  (not A166) );
 a10147a <=( A167  and  a10146a );
 a10151a <=( A202  and  (not A201) );
 a10152a <=( A200  and  a10151a );
 a10153a <=( a10152a  and  a10147a );
 a10157a <=( (not A298)  and  A234 );
 a10158a <=( A233  and  a10157a );
 a10162a <=( A302  and  (not A301) );
 a10163a <=( A299  and  a10162a );
 a10164a <=( a10163a  and  a10158a );
 a10168a <=( (not A199)  and  (not A166) );
 a10169a <=( A167  and  a10168a );
 a10173a <=( A202  and  (not A201) );
 a10174a <=( A200  and  a10173a );
 a10175a <=( a10174a  and  a10169a );
 a10179a <=( (not A298)  and  A234 );
 a10180a <=( A233  and  a10179a );
 a10184a <=( (not A302)  and  A301 );
 a10185a <=( (not A299)  and  a10184a );
 a10186a <=( a10185a  and  a10180a );
 a10190a <=( (not A199)  and  (not A166) );
 a10191a <=( A167  and  a10190a );
 a10195a <=( A202  and  (not A201) );
 a10196a <=( A200  and  a10195a );
 a10197a <=( a10196a  and  a10191a );
 a10201a <=( A265  and  A234 );
 a10202a <=( A233  and  a10201a );
 a10206a <=( (not A269)  and  A268 );
 a10207a <=( A266  and  a10206a );
 a10208a <=( a10207a  and  a10202a );
 a10212a <=( (not A199)  and  (not A166) );
 a10213a <=( A167  and  a10212a );
 a10217a <=( A202  and  (not A201) );
 a10218a <=( A200  and  a10217a );
 a10219a <=( a10218a  and  a10213a );
 a10223a <=( (not A265)  and  A234 );
 a10224a <=( A233  and  a10223a );
 a10228a <=( A269  and  (not A268) );
 a10229a <=( A266  and  a10228a );
 a10230a <=( a10229a  and  a10224a );
 a10234a <=( (not A199)  and  (not A166) );
 a10235a <=( A167  and  a10234a );
 a10239a <=( A202  and  (not A201) );
 a10240a <=( A200  and  a10239a );
 a10241a <=( a10240a  and  a10235a );
 a10245a <=( A265  and  A234 );
 a10246a <=( A233  and  a10245a );
 a10250a <=( A269  and  (not A268) );
 a10251a <=( (not A266)  and  a10250a );
 a10252a <=( a10251a  and  a10246a );
 a10256a <=( (not A199)  and  (not A166) );
 a10257a <=( A167  and  a10256a );
 a10261a <=( A202  and  (not A201) );
 a10262a <=( A200  and  a10261a );
 a10263a <=( a10262a  and  a10257a );
 a10267a <=( (not A265)  and  A234 );
 a10268a <=( A233  and  a10267a );
 a10272a <=( (not A269)  and  A268 );
 a10273a <=( (not A266)  and  a10272a );
 a10274a <=( a10273a  and  a10268a );
 a10278a <=( (not A199)  and  (not A166) );
 a10279a <=( A167  and  a10278a );
 a10283a <=( A202  and  (not A201) );
 a10284a <=( A200  and  a10283a );
 a10285a <=( a10284a  and  a10279a );
 a10289a <=( A235  and  A233 );
 a10290a <=( A232  and  a10289a );
 a10294a <=( A300  and  A299 );
 a10295a <=( (not A236)  and  a10294a );
 a10296a <=( a10295a  and  a10290a );
 a10300a <=( (not A199)  and  (not A166) );
 a10301a <=( A167  and  a10300a );
 a10305a <=( A202  and  (not A201) );
 a10306a <=( A200  and  a10305a );
 a10307a <=( a10306a  and  a10301a );
 a10311a <=( A235  and  A233 );
 a10312a <=( A232  and  a10311a );
 a10316a <=( A300  and  A298 );
 a10317a <=( (not A236)  and  a10316a );
 a10318a <=( a10317a  and  a10312a );
 a10322a <=( (not A199)  and  (not A166) );
 a10323a <=( A167  and  a10322a );
 a10327a <=( A202  and  (not A201) );
 a10328a <=( A200  and  a10327a );
 a10329a <=( a10328a  and  a10323a );
 a10333a <=( A235  and  A233 );
 a10334a <=( A232  and  a10333a );
 a10338a <=( A267  and  A265 );
 a10339a <=( (not A236)  and  a10338a );
 a10340a <=( a10339a  and  a10334a );
 a10344a <=( (not A199)  and  (not A166) );
 a10345a <=( A167  and  a10344a );
 a10349a <=( A202  and  (not A201) );
 a10350a <=( A200  and  a10349a );
 a10351a <=( a10350a  and  a10345a );
 a10355a <=( A235  and  A233 );
 a10356a <=( A232  and  a10355a );
 a10360a <=( A267  and  A266 );
 a10361a <=( (not A236)  and  a10360a );
 a10362a <=( a10361a  and  a10356a );
 a10366a <=( (not A199)  and  (not A166) );
 a10367a <=( A167  and  a10366a );
 a10371a <=( A202  and  (not A201) );
 a10372a <=( A200  and  a10371a );
 a10373a <=( a10372a  and  a10367a );
 a10377a <=( (not A235)  and  A233 );
 a10378a <=( (not A232)  and  a10377a );
 a10382a <=( A300  and  A299 );
 a10383a <=( A236  and  a10382a );
 a10384a <=( a10383a  and  a10378a );
 a10388a <=( (not A199)  and  (not A166) );
 a10389a <=( A167  and  a10388a );
 a10393a <=( A202  and  (not A201) );
 a10394a <=( A200  and  a10393a );
 a10395a <=( a10394a  and  a10389a );
 a10399a <=( (not A235)  and  A233 );
 a10400a <=( (not A232)  and  a10399a );
 a10404a <=( A300  and  A298 );
 a10405a <=( A236  and  a10404a );
 a10406a <=( a10405a  and  a10400a );
 a10410a <=( (not A199)  and  (not A166) );
 a10411a <=( A167  and  a10410a );
 a10415a <=( A202  and  (not A201) );
 a10416a <=( A200  and  a10415a );
 a10417a <=( a10416a  and  a10411a );
 a10421a <=( (not A235)  and  A233 );
 a10422a <=( (not A232)  and  a10421a );
 a10426a <=( A267  and  A265 );
 a10427a <=( A236  and  a10426a );
 a10428a <=( a10427a  and  a10422a );
 a10432a <=( (not A199)  and  (not A166) );
 a10433a <=( A167  and  a10432a );
 a10437a <=( A202  and  (not A201) );
 a10438a <=( A200  and  a10437a );
 a10439a <=( a10438a  and  a10433a );
 a10443a <=( (not A235)  and  A233 );
 a10444a <=( (not A232)  and  a10443a );
 a10448a <=( A267  and  A266 );
 a10449a <=( A236  and  a10448a );
 a10450a <=( a10449a  and  a10444a );
 a10454a <=( (not A199)  and  (not A166) );
 a10455a <=( A167  and  a10454a );
 a10459a <=( A202  and  (not A201) );
 a10460a <=( A200  and  a10459a );
 a10461a <=( a10460a  and  a10455a );
 a10465a <=( (not A235)  and  (not A233) );
 a10466a <=( A232  and  a10465a );
 a10470a <=( A300  and  A299 );
 a10471a <=( A236  and  a10470a );
 a10472a <=( a10471a  and  a10466a );
 a10476a <=( (not A199)  and  (not A166) );
 a10477a <=( A167  and  a10476a );
 a10481a <=( A202  and  (not A201) );
 a10482a <=( A200  and  a10481a );
 a10483a <=( a10482a  and  a10477a );
 a10487a <=( (not A235)  and  (not A233) );
 a10488a <=( A232  and  a10487a );
 a10492a <=( A300  and  A298 );
 a10493a <=( A236  and  a10492a );
 a10494a <=( a10493a  and  a10488a );
 a10498a <=( (not A199)  and  (not A166) );
 a10499a <=( A167  and  a10498a );
 a10503a <=( A202  and  (not A201) );
 a10504a <=( A200  and  a10503a );
 a10505a <=( a10504a  and  a10499a );
 a10509a <=( (not A235)  and  (not A233) );
 a10510a <=( A232  and  a10509a );
 a10514a <=( A267  and  A265 );
 a10515a <=( A236  and  a10514a );
 a10516a <=( a10515a  and  a10510a );
 a10520a <=( (not A199)  and  (not A166) );
 a10521a <=( A167  and  a10520a );
 a10525a <=( A202  and  (not A201) );
 a10526a <=( A200  and  a10525a );
 a10527a <=( a10526a  and  a10521a );
 a10531a <=( (not A235)  and  (not A233) );
 a10532a <=( A232  and  a10531a );
 a10536a <=( A267  and  A266 );
 a10537a <=( A236  and  a10536a );
 a10538a <=( a10537a  and  a10532a );
 a10542a <=( (not A199)  and  (not A166) );
 a10543a <=( A167  and  a10542a );
 a10547a <=( A202  and  (not A201) );
 a10548a <=( A200  and  a10547a );
 a10549a <=( a10548a  and  a10543a );
 a10553a <=( A235  and  (not A233) );
 a10554a <=( (not A232)  and  a10553a );
 a10558a <=( A300  and  A299 );
 a10559a <=( (not A236)  and  a10558a );
 a10560a <=( a10559a  and  a10554a );
 a10564a <=( (not A199)  and  (not A166) );
 a10565a <=( A167  and  a10564a );
 a10569a <=( A202  and  (not A201) );
 a10570a <=( A200  and  a10569a );
 a10571a <=( a10570a  and  a10565a );
 a10575a <=( A235  and  (not A233) );
 a10576a <=( (not A232)  and  a10575a );
 a10580a <=( A300  and  A298 );
 a10581a <=( (not A236)  and  a10580a );
 a10582a <=( a10581a  and  a10576a );
 a10586a <=( (not A199)  and  (not A166) );
 a10587a <=( A167  and  a10586a );
 a10591a <=( A202  and  (not A201) );
 a10592a <=( A200  and  a10591a );
 a10593a <=( a10592a  and  a10587a );
 a10597a <=( A235  and  (not A233) );
 a10598a <=( (not A232)  and  a10597a );
 a10602a <=( A267  and  A265 );
 a10603a <=( (not A236)  and  a10602a );
 a10604a <=( a10603a  and  a10598a );
 a10608a <=( (not A199)  and  (not A166) );
 a10609a <=( A167  and  a10608a );
 a10613a <=( A202  and  (not A201) );
 a10614a <=( A200  and  a10613a );
 a10615a <=( a10614a  and  a10609a );
 a10619a <=( A235  and  (not A233) );
 a10620a <=( (not A232)  and  a10619a );
 a10624a <=( A267  and  A266 );
 a10625a <=( (not A236)  and  a10624a );
 a10626a <=( a10625a  and  a10620a );
 a10630a <=( (not A199)  and  (not A166) );
 a10631a <=( A167  and  a10630a );
 a10635a <=( (not A203)  and  (not A201) );
 a10636a <=( A200  and  a10635a );
 a10637a <=( a10636a  and  a10631a );
 a10641a <=( A298  and  A234 );
 a10642a <=( A232  and  a10641a );
 a10646a <=( (not A302)  and  A301 );
 a10647a <=( A299  and  a10646a );
 a10648a <=( a10647a  and  a10642a );
 a10652a <=( (not A199)  and  (not A166) );
 a10653a <=( A167  and  a10652a );
 a10657a <=( (not A203)  and  (not A201) );
 a10658a <=( A200  and  a10657a );
 a10659a <=( a10658a  and  a10653a );
 a10663a <=( A298  and  A234 );
 a10664a <=( A232  and  a10663a );
 a10668a <=( A302  and  (not A301) );
 a10669a <=( (not A299)  and  a10668a );
 a10670a <=( a10669a  and  a10664a );
 a10674a <=( (not A199)  and  (not A166) );
 a10675a <=( A167  and  a10674a );
 a10679a <=( (not A203)  and  (not A201) );
 a10680a <=( A200  and  a10679a );
 a10681a <=( a10680a  and  a10675a );
 a10685a <=( (not A298)  and  A234 );
 a10686a <=( A232  and  a10685a );
 a10690a <=( A302  and  (not A301) );
 a10691a <=( A299  and  a10690a );
 a10692a <=( a10691a  and  a10686a );
 a10696a <=( (not A199)  and  (not A166) );
 a10697a <=( A167  and  a10696a );
 a10701a <=( (not A203)  and  (not A201) );
 a10702a <=( A200  and  a10701a );
 a10703a <=( a10702a  and  a10697a );
 a10707a <=( (not A298)  and  A234 );
 a10708a <=( A232  and  a10707a );
 a10712a <=( (not A302)  and  A301 );
 a10713a <=( (not A299)  and  a10712a );
 a10714a <=( a10713a  and  a10708a );
 a10718a <=( (not A199)  and  (not A166) );
 a10719a <=( A167  and  a10718a );
 a10723a <=( (not A203)  and  (not A201) );
 a10724a <=( A200  and  a10723a );
 a10725a <=( a10724a  and  a10719a );
 a10729a <=( A265  and  A234 );
 a10730a <=( A232  and  a10729a );
 a10734a <=( (not A269)  and  A268 );
 a10735a <=( A266  and  a10734a );
 a10736a <=( a10735a  and  a10730a );
 a10740a <=( (not A199)  and  (not A166) );
 a10741a <=( A167  and  a10740a );
 a10745a <=( (not A203)  and  (not A201) );
 a10746a <=( A200  and  a10745a );
 a10747a <=( a10746a  and  a10741a );
 a10751a <=( (not A265)  and  A234 );
 a10752a <=( A232  and  a10751a );
 a10756a <=( A269  and  (not A268) );
 a10757a <=( A266  and  a10756a );
 a10758a <=( a10757a  and  a10752a );
 a10762a <=( (not A199)  and  (not A166) );
 a10763a <=( A167  and  a10762a );
 a10767a <=( (not A203)  and  (not A201) );
 a10768a <=( A200  and  a10767a );
 a10769a <=( a10768a  and  a10763a );
 a10773a <=( A265  and  A234 );
 a10774a <=( A232  and  a10773a );
 a10778a <=( A269  and  (not A268) );
 a10779a <=( (not A266)  and  a10778a );
 a10780a <=( a10779a  and  a10774a );
 a10784a <=( (not A199)  and  (not A166) );
 a10785a <=( A167  and  a10784a );
 a10789a <=( (not A203)  and  (not A201) );
 a10790a <=( A200  and  a10789a );
 a10791a <=( a10790a  and  a10785a );
 a10795a <=( (not A265)  and  A234 );
 a10796a <=( A232  and  a10795a );
 a10800a <=( (not A269)  and  A268 );
 a10801a <=( (not A266)  and  a10800a );
 a10802a <=( a10801a  and  a10796a );
 a10806a <=( (not A199)  and  (not A166) );
 a10807a <=( A167  and  a10806a );
 a10811a <=( (not A203)  and  (not A201) );
 a10812a <=( A200  and  a10811a );
 a10813a <=( a10812a  and  a10807a );
 a10817a <=( A298  and  A234 );
 a10818a <=( A233  and  a10817a );
 a10822a <=( (not A302)  and  A301 );
 a10823a <=( A299  and  a10822a );
 a10824a <=( a10823a  and  a10818a );
 a10828a <=( (not A199)  and  (not A166) );
 a10829a <=( A167  and  a10828a );
 a10833a <=( (not A203)  and  (not A201) );
 a10834a <=( A200  and  a10833a );
 a10835a <=( a10834a  and  a10829a );
 a10839a <=( A298  and  A234 );
 a10840a <=( A233  and  a10839a );
 a10844a <=( A302  and  (not A301) );
 a10845a <=( (not A299)  and  a10844a );
 a10846a <=( a10845a  and  a10840a );
 a10850a <=( (not A199)  and  (not A166) );
 a10851a <=( A167  and  a10850a );
 a10855a <=( (not A203)  and  (not A201) );
 a10856a <=( A200  and  a10855a );
 a10857a <=( a10856a  and  a10851a );
 a10861a <=( (not A298)  and  A234 );
 a10862a <=( A233  and  a10861a );
 a10866a <=( A302  and  (not A301) );
 a10867a <=( A299  and  a10866a );
 a10868a <=( a10867a  and  a10862a );
 a10872a <=( (not A199)  and  (not A166) );
 a10873a <=( A167  and  a10872a );
 a10877a <=( (not A203)  and  (not A201) );
 a10878a <=( A200  and  a10877a );
 a10879a <=( a10878a  and  a10873a );
 a10883a <=( (not A298)  and  A234 );
 a10884a <=( A233  and  a10883a );
 a10888a <=( (not A302)  and  A301 );
 a10889a <=( (not A299)  and  a10888a );
 a10890a <=( a10889a  and  a10884a );
 a10894a <=( (not A199)  and  (not A166) );
 a10895a <=( A167  and  a10894a );
 a10899a <=( (not A203)  and  (not A201) );
 a10900a <=( A200  and  a10899a );
 a10901a <=( a10900a  and  a10895a );
 a10905a <=( A265  and  A234 );
 a10906a <=( A233  and  a10905a );
 a10910a <=( (not A269)  and  A268 );
 a10911a <=( A266  and  a10910a );
 a10912a <=( a10911a  and  a10906a );
 a10916a <=( (not A199)  and  (not A166) );
 a10917a <=( A167  and  a10916a );
 a10921a <=( (not A203)  and  (not A201) );
 a10922a <=( A200  and  a10921a );
 a10923a <=( a10922a  and  a10917a );
 a10927a <=( (not A265)  and  A234 );
 a10928a <=( A233  and  a10927a );
 a10932a <=( A269  and  (not A268) );
 a10933a <=( A266  and  a10932a );
 a10934a <=( a10933a  and  a10928a );
 a10938a <=( (not A199)  and  (not A166) );
 a10939a <=( A167  and  a10938a );
 a10943a <=( (not A203)  and  (not A201) );
 a10944a <=( A200  and  a10943a );
 a10945a <=( a10944a  and  a10939a );
 a10949a <=( A265  and  A234 );
 a10950a <=( A233  and  a10949a );
 a10954a <=( A269  and  (not A268) );
 a10955a <=( (not A266)  and  a10954a );
 a10956a <=( a10955a  and  a10950a );
 a10960a <=( (not A199)  and  (not A166) );
 a10961a <=( A167  and  a10960a );
 a10965a <=( (not A203)  and  (not A201) );
 a10966a <=( A200  and  a10965a );
 a10967a <=( a10966a  and  a10961a );
 a10971a <=( (not A265)  and  A234 );
 a10972a <=( A233  and  a10971a );
 a10976a <=( (not A269)  and  A268 );
 a10977a <=( (not A266)  and  a10976a );
 a10978a <=( a10977a  and  a10972a );
 a10982a <=( (not A199)  and  (not A166) );
 a10983a <=( A167  and  a10982a );
 a10987a <=( (not A203)  and  (not A201) );
 a10988a <=( A200  and  a10987a );
 a10989a <=( a10988a  and  a10983a );
 a10993a <=( A235  and  A233 );
 a10994a <=( A232  and  a10993a );
 a10998a <=( A300  and  A299 );
 a10999a <=( (not A236)  and  a10998a );
 a11000a <=( a10999a  and  a10994a );
 a11004a <=( (not A199)  and  (not A166) );
 a11005a <=( A167  and  a11004a );
 a11009a <=( (not A203)  and  (not A201) );
 a11010a <=( A200  and  a11009a );
 a11011a <=( a11010a  and  a11005a );
 a11015a <=( A235  and  A233 );
 a11016a <=( A232  and  a11015a );
 a11020a <=( A300  and  A298 );
 a11021a <=( (not A236)  and  a11020a );
 a11022a <=( a11021a  and  a11016a );
 a11026a <=( (not A199)  and  (not A166) );
 a11027a <=( A167  and  a11026a );
 a11031a <=( (not A203)  and  (not A201) );
 a11032a <=( A200  and  a11031a );
 a11033a <=( a11032a  and  a11027a );
 a11037a <=( A235  and  A233 );
 a11038a <=( A232  and  a11037a );
 a11042a <=( A267  and  A265 );
 a11043a <=( (not A236)  and  a11042a );
 a11044a <=( a11043a  and  a11038a );
 a11048a <=( (not A199)  and  (not A166) );
 a11049a <=( A167  and  a11048a );
 a11053a <=( (not A203)  and  (not A201) );
 a11054a <=( A200  and  a11053a );
 a11055a <=( a11054a  and  a11049a );
 a11059a <=( A235  and  A233 );
 a11060a <=( A232  and  a11059a );
 a11064a <=( A267  and  A266 );
 a11065a <=( (not A236)  and  a11064a );
 a11066a <=( a11065a  and  a11060a );
 a11070a <=( (not A199)  and  (not A166) );
 a11071a <=( A167  and  a11070a );
 a11075a <=( (not A203)  and  (not A201) );
 a11076a <=( A200  and  a11075a );
 a11077a <=( a11076a  and  a11071a );
 a11081a <=( (not A235)  and  A233 );
 a11082a <=( (not A232)  and  a11081a );
 a11086a <=( A300  and  A299 );
 a11087a <=( A236  and  a11086a );
 a11088a <=( a11087a  and  a11082a );
 a11092a <=( (not A199)  and  (not A166) );
 a11093a <=( A167  and  a11092a );
 a11097a <=( (not A203)  and  (not A201) );
 a11098a <=( A200  and  a11097a );
 a11099a <=( a11098a  and  a11093a );
 a11103a <=( (not A235)  and  A233 );
 a11104a <=( (not A232)  and  a11103a );
 a11108a <=( A300  and  A298 );
 a11109a <=( A236  and  a11108a );
 a11110a <=( a11109a  and  a11104a );
 a11114a <=( (not A199)  and  (not A166) );
 a11115a <=( A167  and  a11114a );
 a11119a <=( (not A203)  and  (not A201) );
 a11120a <=( A200  and  a11119a );
 a11121a <=( a11120a  and  a11115a );
 a11125a <=( (not A235)  and  A233 );
 a11126a <=( (not A232)  and  a11125a );
 a11130a <=( A267  and  A265 );
 a11131a <=( A236  and  a11130a );
 a11132a <=( a11131a  and  a11126a );
 a11136a <=( (not A199)  and  (not A166) );
 a11137a <=( A167  and  a11136a );
 a11141a <=( (not A203)  and  (not A201) );
 a11142a <=( A200  and  a11141a );
 a11143a <=( a11142a  and  a11137a );
 a11147a <=( (not A235)  and  A233 );
 a11148a <=( (not A232)  and  a11147a );
 a11152a <=( A267  and  A266 );
 a11153a <=( A236  and  a11152a );
 a11154a <=( a11153a  and  a11148a );
 a11158a <=( (not A199)  and  (not A166) );
 a11159a <=( A167  and  a11158a );
 a11163a <=( (not A203)  and  (not A201) );
 a11164a <=( A200  and  a11163a );
 a11165a <=( a11164a  and  a11159a );
 a11169a <=( (not A235)  and  (not A233) );
 a11170a <=( A232  and  a11169a );
 a11174a <=( A300  and  A299 );
 a11175a <=( A236  and  a11174a );
 a11176a <=( a11175a  and  a11170a );
 a11180a <=( (not A199)  and  (not A166) );
 a11181a <=( A167  and  a11180a );
 a11185a <=( (not A203)  and  (not A201) );
 a11186a <=( A200  and  a11185a );
 a11187a <=( a11186a  and  a11181a );
 a11191a <=( (not A235)  and  (not A233) );
 a11192a <=( A232  and  a11191a );
 a11196a <=( A300  and  A298 );
 a11197a <=( A236  and  a11196a );
 a11198a <=( a11197a  and  a11192a );
 a11202a <=( (not A199)  and  (not A166) );
 a11203a <=( A167  and  a11202a );
 a11207a <=( (not A203)  and  (not A201) );
 a11208a <=( A200  and  a11207a );
 a11209a <=( a11208a  and  a11203a );
 a11213a <=( (not A235)  and  (not A233) );
 a11214a <=( A232  and  a11213a );
 a11218a <=( A267  and  A265 );
 a11219a <=( A236  and  a11218a );
 a11220a <=( a11219a  and  a11214a );
 a11224a <=( (not A199)  and  (not A166) );
 a11225a <=( A167  and  a11224a );
 a11229a <=( (not A203)  and  (not A201) );
 a11230a <=( A200  and  a11229a );
 a11231a <=( a11230a  and  a11225a );
 a11235a <=( (not A235)  and  (not A233) );
 a11236a <=( A232  and  a11235a );
 a11240a <=( A267  and  A266 );
 a11241a <=( A236  and  a11240a );
 a11242a <=( a11241a  and  a11236a );
 a11246a <=( (not A199)  and  (not A166) );
 a11247a <=( A167  and  a11246a );
 a11251a <=( (not A203)  and  (not A201) );
 a11252a <=( A200  and  a11251a );
 a11253a <=( a11252a  and  a11247a );
 a11257a <=( A235  and  (not A233) );
 a11258a <=( (not A232)  and  a11257a );
 a11262a <=( A300  and  A299 );
 a11263a <=( (not A236)  and  a11262a );
 a11264a <=( a11263a  and  a11258a );
 a11268a <=( (not A199)  and  (not A166) );
 a11269a <=( A167  and  a11268a );
 a11273a <=( (not A203)  and  (not A201) );
 a11274a <=( A200  and  a11273a );
 a11275a <=( a11274a  and  a11269a );
 a11279a <=( A235  and  (not A233) );
 a11280a <=( (not A232)  and  a11279a );
 a11284a <=( A300  and  A298 );
 a11285a <=( (not A236)  and  a11284a );
 a11286a <=( a11285a  and  a11280a );
 a11290a <=( (not A199)  and  (not A166) );
 a11291a <=( A167  and  a11290a );
 a11295a <=( (not A203)  and  (not A201) );
 a11296a <=( A200  and  a11295a );
 a11297a <=( a11296a  and  a11291a );
 a11301a <=( A235  and  (not A233) );
 a11302a <=( (not A232)  and  a11301a );
 a11306a <=( A267  and  A265 );
 a11307a <=( (not A236)  and  a11306a );
 a11308a <=( a11307a  and  a11302a );
 a11312a <=( (not A199)  and  (not A166) );
 a11313a <=( A167  and  a11312a );
 a11317a <=( (not A203)  and  (not A201) );
 a11318a <=( A200  and  a11317a );
 a11319a <=( a11318a  and  a11313a );
 a11323a <=( A235  and  (not A233) );
 a11324a <=( (not A232)  and  a11323a );
 a11328a <=( A267  and  A266 );
 a11329a <=( (not A236)  and  a11328a );
 a11330a <=( a11329a  and  a11324a );
 a11334a <=( A199  and  (not A166) );
 a11335a <=( A167  and  a11334a );
 a11339a <=( A202  and  (not A201) );
 a11340a <=( (not A200)  and  a11339a );
 a11341a <=( a11340a  and  a11335a );
 a11345a <=( A298  and  A234 );
 a11346a <=( A232  and  a11345a );
 a11350a <=( (not A302)  and  A301 );
 a11351a <=( A299  and  a11350a );
 a11352a <=( a11351a  and  a11346a );
 a11356a <=( A199  and  (not A166) );
 a11357a <=( A167  and  a11356a );
 a11361a <=( A202  and  (not A201) );
 a11362a <=( (not A200)  and  a11361a );
 a11363a <=( a11362a  and  a11357a );
 a11367a <=( A298  and  A234 );
 a11368a <=( A232  and  a11367a );
 a11372a <=( A302  and  (not A301) );
 a11373a <=( (not A299)  and  a11372a );
 a11374a <=( a11373a  and  a11368a );
 a11378a <=( A199  and  (not A166) );
 a11379a <=( A167  and  a11378a );
 a11383a <=( A202  and  (not A201) );
 a11384a <=( (not A200)  and  a11383a );
 a11385a <=( a11384a  and  a11379a );
 a11389a <=( (not A298)  and  A234 );
 a11390a <=( A232  and  a11389a );
 a11394a <=( A302  and  (not A301) );
 a11395a <=( A299  and  a11394a );
 a11396a <=( a11395a  and  a11390a );
 a11400a <=( A199  and  (not A166) );
 a11401a <=( A167  and  a11400a );
 a11405a <=( A202  and  (not A201) );
 a11406a <=( (not A200)  and  a11405a );
 a11407a <=( a11406a  and  a11401a );
 a11411a <=( (not A298)  and  A234 );
 a11412a <=( A232  and  a11411a );
 a11416a <=( (not A302)  and  A301 );
 a11417a <=( (not A299)  and  a11416a );
 a11418a <=( a11417a  and  a11412a );
 a11422a <=( A199  and  (not A166) );
 a11423a <=( A167  and  a11422a );
 a11427a <=( A202  and  (not A201) );
 a11428a <=( (not A200)  and  a11427a );
 a11429a <=( a11428a  and  a11423a );
 a11433a <=( A265  and  A234 );
 a11434a <=( A232  and  a11433a );
 a11438a <=( (not A269)  and  A268 );
 a11439a <=( A266  and  a11438a );
 a11440a <=( a11439a  and  a11434a );
 a11444a <=( A199  and  (not A166) );
 a11445a <=( A167  and  a11444a );
 a11449a <=( A202  and  (not A201) );
 a11450a <=( (not A200)  and  a11449a );
 a11451a <=( a11450a  and  a11445a );
 a11455a <=( (not A265)  and  A234 );
 a11456a <=( A232  and  a11455a );
 a11460a <=( A269  and  (not A268) );
 a11461a <=( A266  and  a11460a );
 a11462a <=( a11461a  and  a11456a );
 a11466a <=( A199  and  (not A166) );
 a11467a <=( A167  and  a11466a );
 a11471a <=( A202  and  (not A201) );
 a11472a <=( (not A200)  and  a11471a );
 a11473a <=( a11472a  and  a11467a );
 a11477a <=( A265  and  A234 );
 a11478a <=( A232  and  a11477a );
 a11482a <=( A269  and  (not A268) );
 a11483a <=( (not A266)  and  a11482a );
 a11484a <=( a11483a  and  a11478a );
 a11488a <=( A199  and  (not A166) );
 a11489a <=( A167  and  a11488a );
 a11493a <=( A202  and  (not A201) );
 a11494a <=( (not A200)  and  a11493a );
 a11495a <=( a11494a  and  a11489a );
 a11499a <=( (not A265)  and  A234 );
 a11500a <=( A232  and  a11499a );
 a11504a <=( (not A269)  and  A268 );
 a11505a <=( (not A266)  and  a11504a );
 a11506a <=( a11505a  and  a11500a );
 a11510a <=( A199  and  (not A166) );
 a11511a <=( A167  and  a11510a );
 a11515a <=( A202  and  (not A201) );
 a11516a <=( (not A200)  and  a11515a );
 a11517a <=( a11516a  and  a11511a );
 a11521a <=( A298  and  A234 );
 a11522a <=( A233  and  a11521a );
 a11526a <=( (not A302)  and  A301 );
 a11527a <=( A299  and  a11526a );
 a11528a <=( a11527a  and  a11522a );
 a11532a <=( A199  and  (not A166) );
 a11533a <=( A167  and  a11532a );
 a11537a <=( A202  and  (not A201) );
 a11538a <=( (not A200)  and  a11537a );
 a11539a <=( a11538a  and  a11533a );
 a11543a <=( A298  and  A234 );
 a11544a <=( A233  and  a11543a );
 a11548a <=( A302  and  (not A301) );
 a11549a <=( (not A299)  and  a11548a );
 a11550a <=( a11549a  and  a11544a );
 a11554a <=( A199  and  (not A166) );
 a11555a <=( A167  and  a11554a );
 a11559a <=( A202  and  (not A201) );
 a11560a <=( (not A200)  and  a11559a );
 a11561a <=( a11560a  and  a11555a );
 a11565a <=( (not A298)  and  A234 );
 a11566a <=( A233  and  a11565a );
 a11570a <=( A302  and  (not A301) );
 a11571a <=( A299  and  a11570a );
 a11572a <=( a11571a  and  a11566a );
 a11576a <=( A199  and  (not A166) );
 a11577a <=( A167  and  a11576a );
 a11581a <=( A202  and  (not A201) );
 a11582a <=( (not A200)  and  a11581a );
 a11583a <=( a11582a  and  a11577a );
 a11587a <=( (not A298)  and  A234 );
 a11588a <=( A233  and  a11587a );
 a11592a <=( (not A302)  and  A301 );
 a11593a <=( (not A299)  and  a11592a );
 a11594a <=( a11593a  and  a11588a );
 a11598a <=( A199  and  (not A166) );
 a11599a <=( A167  and  a11598a );
 a11603a <=( A202  and  (not A201) );
 a11604a <=( (not A200)  and  a11603a );
 a11605a <=( a11604a  and  a11599a );
 a11609a <=( A265  and  A234 );
 a11610a <=( A233  and  a11609a );
 a11614a <=( (not A269)  and  A268 );
 a11615a <=( A266  and  a11614a );
 a11616a <=( a11615a  and  a11610a );
 a11620a <=( A199  and  (not A166) );
 a11621a <=( A167  and  a11620a );
 a11625a <=( A202  and  (not A201) );
 a11626a <=( (not A200)  and  a11625a );
 a11627a <=( a11626a  and  a11621a );
 a11631a <=( (not A265)  and  A234 );
 a11632a <=( A233  and  a11631a );
 a11636a <=( A269  and  (not A268) );
 a11637a <=( A266  and  a11636a );
 a11638a <=( a11637a  and  a11632a );
 a11642a <=( A199  and  (not A166) );
 a11643a <=( A167  and  a11642a );
 a11647a <=( A202  and  (not A201) );
 a11648a <=( (not A200)  and  a11647a );
 a11649a <=( a11648a  and  a11643a );
 a11653a <=( A265  and  A234 );
 a11654a <=( A233  and  a11653a );
 a11658a <=( A269  and  (not A268) );
 a11659a <=( (not A266)  and  a11658a );
 a11660a <=( a11659a  and  a11654a );
 a11664a <=( A199  and  (not A166) );
 a11665a <=( A167  and  a11664a );
 a11669a <=( A202  and  (not A201) );
 a11670a <=( (not A200)  and  a11669a );
 a11671a <=( a11670a  and  a11665a );
 a11675a <=( (not A265)  and  A234 );
 a11676a <=( A233  and  a11675a );
 a11680a <=( (not A269)  and  A268 );
 a11681a <=( (not A266)  and  a11680a );
 a11682a <=( a11681a  and  a11676a );
 a11686a <=( A199  and  (not A166) );
 a11687a <=( A167  and  a11686a );
 a11691a <=( A202  and  (not A201) );
 a11692a <=( (not A200)  and  a11691a );
 a11693a <=( a11692a  and  a11687a );
 a11697a <=( A235  and  A233 );
 a11698a <=( A232  and  a11697a );
 a11702a <=( A300  and  A299 );
 a11703a <=( (not A236)  and  a11702a );
 a11704a <=( a11703a  and  a11698a );
 a11708a <=( A199  and  (not A166) );
 a11709a <=( A167  and  a11708a );
 a11713a <=( A202  and  (not A201) );
 a11714a <=( (not A200)  and  a11713a );
 a11715a <=( a11714a  and  a11709a );
 a11719a <=( A235  and  A233 );
 a11720a <=( A232  and  a11719a );
 a11724a <=( A300  and  A298 );
 a11725a <=( (not A236)  and  a11724a );
 a11726a <=( a11725a  and  a11720a );
 a11730a <=( A199  and  (not A166) );
 a11731a <=( A167  and  a11730a );
 a11735a <=( A202  and  (not A201) );
 a11736a <=( (not A200)  and  a11735a );
 a11737a <=( a11736a  and  a11731a );
 a11741a <=( A235  and  A233 );
 a11742a <=( A232  and  a11741a );
 a11746a <=( A267  and  A265 );
 a11747a <=( (not A236)  and  a11746a );
 a11748a <=( a11747a  and  a11742a );
 a11752a <=( A199  and  (not A166) );
 a11753a <=( A167  and  a11752a );
 a11757a <=( A202  and  (not A201) );
 a11758a <=( (not A200)  and  a11757a );
 a11759a <=( a11758a  and  a11753a );
 a11763a <=( A235  and  A233 );
 a11764a <=( A232  and  a11763a );
 a11768a <=( A267  and  A266 );
 a11769a <=( (not A236)  and  a11768a );
 a11770a <=( a11769a  and  a11764a );
 a11774a <=( A199  and  (not A166) );
 a11775a <=( A167  and  a11774a );
 a11779a <=( A202  and  (not A201) );
 a11780a <=( (not A200)  and  a11779a );
 a11781a <=( a11780a  and  a11775a );
 a11785a <=( (not A235)  and  A233 );
 a11786a <=( (not A232)  and  a11785a );
 a11790a <=( A300  and  A299 );
 a11791a <=( A236  and  a11790a );
 a11792a <=( a11791a  and  a11786a );
 a11796a <=( A199  and  (not A166) );
 a11797a <=( A167  and  a11796a );
 a11801a <=( A202  and  (not A201) );
 a11802a <=( (not A200)  and  a11801a );
 a11803a <=( a11802a  and  a11797a );
 a11807a <=( (not A235)  and  A233 );
 a11808a <=( (not A232)  and  a11807a );
 a11812a <=( A300  and  A298 );
 a11813a <=( A236  and  a11812a );
 a11814a <=( a11813a  and  a11808a );
 a11818a <=( A199  and  (not A166) );
 a11819a <=( A167  and  a11818a );
 a11823a <=( A202  and  (not A201) );
 a11824a <=( (not A200)  and  a11823a );
 a11825a <=( a11824a  and  a11819a );
 a11829a <=( (not A235)  and  A233 );
 a11830a <=( (not A232)  and  a11829a );
 a11834a <=( A267  and  A265 );
 a11835a <=( A236  and  a11834a );
 a11836a <=( a11835a  and  a11830a );
 a11840a <=( A199  and  (not A166) );
 a11841a <=( A167  and  a11840a );
 a11845a <=( A202  and  (not A201) );
 a11846a <=( (not A200)  and  a11845a );
 a11847a <=( a11846a  and  a11841a );
 a11851a <=( (not A235)  and  A233 );
 a11852a <=( (not A232)  and  a11851a );
 a11856a <=( A267  and  A266 );
 a11857a <=( A236  and  a11856a );
 a11858a <=( a11857a  and  a11852a );
 a11862a <=( A199  and  (not A166) );
 a11863a <=( A167  and  a11862a );
 a11867a <=( A202  and  (not A201) );
 a11868a <=( (not A200)  and  a11867a );
 a11869a <=( a11868a  and  a11863a );
 a11873a <=( (not A235)  and  (not A233) );
 a11874a <=( A232  and  a11873a );
 a11878a <=( A300  and  A299 );
 a11879a <=( A236  and  a11878a );
 a11880a <=( a11879a  and  a11874a );
 a11884a <=( A199  and  (not A166) );
 a11885a <=( A167  and  a11884a );
 a11889a <=( A202  and  (not A201) );
 a11890a <=( (not A200)  and  a11889a );
 a11891a <=( a11890a  and  a11885a );
 a11895a <=( (not A235)  and  (not A233) );
 a11896a <=( A232  and  a11895a );
 a11900a <=( A300  and  A298 );
 a11901a <=( A236  and  a11900a );
 a11902a <=( a11901a  and  a11896a );
 a11906a <=( A199  and  (not A166) );
 a11907a <=( A167  and  a11906a );
 a11911a <=( A202  and  (not A201) );
 a11912a <=( (not A200)  and  a11911a );
 a11913a <=( a11912a  and  a11907a );
 a11917a <=( (not A235)  and  (not A233) );
 a11918a <=( A232  and  a11917a );
 a11922a <=( A267  and  A265 );
 a11923a <=( A236  and  a11922a );
 a11924a <=( a11923a  and  a11918a );
 a11928a <=( A199  and  (not A166) );
 a11929a <=( A167  and  a11928a );
 a11933a <=( A202  and  (not A201) );
 a11934a <=( (not A200)  and  a11933a );
 a11935a <=( a11934a  and  a11929a );
 a11939a <=( (not A235)  and  (not A233) );
 a11940a <=( A232  and  a11939a );
 a11944a <=( A267  and  A266 );
 a11945a <=( A236  and  a11944a );
 a11946a <=( a11945a  and  a11940a );
 a11950a <=( A199  and  (not A166) );
 a11951a <=( A167  and  a11950a );
 a11955a <=( A202  and  (not A201) );
 a11956a <=( (not A200)  and  a11955a );
 a11957a <=( a11956a  and  a11951a );
 a11961a <=( A235  and  (not A233) );
 a11962a <=( (not A232)  and  a11961a );
 a11966a <=( A300  and  A299 );
 a11967a <=( (not A236)  and  a11966a );
 a11968a <=( a11967a  and  a11962a );
 a11972a <=( A199  and  (not A166) );
 a11973a <=( A167  and  a11972a );
 a11977a <=( A202  and  (not A201) );
 a11978a <=( (not A200)  and  a11977a );
 a11979a <=( a11978a  and  a11973a );
 a11983a <=( A235  and  (not A233) );
 a11984a <=( (not A232)  and  a11983a );
 a11988a <=( A300  and  A298 );
 a11989a <=( (not A236)  and  a11988a );
 a11990a <=( a11989a  and  a11984a );
 a11994a <=( A199  and  (not A166) );
 a11995a <=( A167  and  a11994a );
 a11999a <=( A202  and  (not A201) );
 a12000a <=( (not A200)  and  a11999a );
 a12001a <=( a12000a  and  a11995a );
 a12005a <=( A235  and  (not A233) );
 a12006a <=( (not A232)  and  a12005a );
 a12010a <=( A267  and  A265 );
 a12011a <=( (not A236)  and  a12010a );
 a12012a <=( a12011a  and  a12006a );
 a12016a <=( A199  and  (not A166) );
 a12017a <=( A167  and  a12016a );
 a12021a <=( A202  and  (not A201) );
 a12022a <=( (not A200)  and  a12021a );
 a12023a <=( a12022a  and  a12017a );
 a12027a <=( A235  and  (not A233) );
 a12028a <=( (not A232)  and  a12027a );
 a12032a <=( A267  and  A266 );
 a12033a <=( (not A236)  and  a12032a );
 a12034a <=( a12033a  and  a12028a );
 a12038a <=( A199  and  (not A166) );
 a12039a <=( A167  and  a12038a );
 a12043a <=( (not A203)  and  (not A201) );
 a12044a <=( (not A200)  and  a12043a );
 a12045a <=( a12044a  and  a12039a );
 a12049a <=( A298  and  A234 );
 a12050a <=( A232  and  a12049a );
 a12054a <=( (not A302)  and  A301 );
 a12055a <=( A299  and  a12054a );
 a12056a <=( a12055a  and  a12050a );
 a12060a <=( A199  and  (not A166) );
 a12061a <=( A167  and  a12060a );
 a12065a <=( (not A203)  and  (not A201) );
 a12066a <=( (not A200)  and  a12065a );
 a12067a <=( a12066a  and  a12061a );
 a12071a <=( A298  and  A234 );
 a12072a <=( A232  and  a12071a );
 a12076a <=( A302  and  (not A301) );
 a12077a <=( (not A299)  and  a12076a );
 a12078a <=( a12077a  and  a12072a );
 a12082a <=( A199  and  (not A166) );
 a12083a <=( A167  and  a12082a );
 a12087a <=( (not A203)  and  (not A201) );
 a12088a <=( (not A200)  and  a12087a );
 a12089a <=( a12088a  and  a12083a );
 a12093a <=( (not A298)  and  A234 );
 a12094a <=( A232  and  a12093a );
 a12098a <=( A302  and  (not A301) );
 a12099a <=( A299  and  a12098a );
 a12100a <=( a12099a  and  a12094a );
 a12104a <=( A199  and  (not A166) );
 a12105a <=( A167  and  a12104a );
 a12109a <=( (not A203)  and  (not A201) );
 a12110a <=( (not A200)  and  a12109a );
 a12111a <=( a12110a  and  a12105a );
 a12115a <=( (not A298)  and  A234 );
 a12116a <=( A232  and  a12115a );
 a12120a <=( (not A302)  and  A301 );
 a12121a <=( (not A299)  and  a12120a );
 a12122a <=( a12121a  and  a12116a );
 a12126a <=( A199  and  (not A166) );
 a12127a <=( A167  and  a12126a );
 a12131a <=( (not A203)  and  (not A201) );
 a12132a <=( (not A200)  and  a12131a );
 a12133a <=( a12132a  and  a12127a );
 a12137a <=( A265  and  A234 );
 a12138a <=( A232  and  a12137a );
 a12142a <=( (not A269)  and  A268 );
 a12143a <=( A266  and  a12142a );
 a12144a <=( a12143a  and  a12138a );
 a12148a <=( A199  and  (not A166) );
 a12149a <=( A167  and  a12148a );
 a12153a <=( (not A203)  and  (not A201) );
 a12154a <=( (not A200)  and  a12153a );
 a12155a <=( a12154a  and  a12149a );
 a12159a <=( (not A265)  and  A234 );
 a12160a <=( A232  and  a12159a );
 a12164a <=( A269  and  (not A268) );
 a12165a <=( A266  and  a12164a );
 a12166a <=( a12165a  and  a12160a );
 a12170a <=( A199  and  (not A166) );
 a12171a <=( A167  and  a12170a );
 a12175a <=( (not A203)  and  (not A201) );
 a12176a <=( (not A200)  and  a12175a );
 a12177a <=( a12176a  and  a12171a );
 a12181a <=( A265  and  A234 );
 a12182a <=( A232  and  a12181a );
 a12186a <=( A269  and  (not A268) );
 a12187a <=( (not A266)  and  a12186a );
 a12188a <=( a12187a  and  a12182a );
 a12192a <=( A199  and  (not A166) );
 a12193a <=( A167  and  a12192a );
 a12197a <=( (not A203)  and  (not A201) );
 a12198a <=( (not A200)  and  a12197a );
 a12199a <=( a12198a  and  a12193a );
 a12203a <=( (not A265)  and  A234 );
 a12204a <=( A232  and  a12203a );
 a12208a <=( (not A269)  and  A268 );
 a12209a <=( (not A266)  and  a12208a );
 a12210a <=( a12209a  and  a12204a );
 a12214a <=( A199  and  (not A166) );
 a12215a <=( A167  and  a12214a );
 a12219a <=( (not A203)  and  (not A201) );
 a12220a <=( (not A200)  and  a12219a );
 a12221a <=( a12220a  and  a12215a );
 a12225a <=( A298  and  A234 );
 a12226a <=( A233  and  a12225a );
 a12230a <=( (not A302)  and  A301 );
 a12231a <=( A299  and  a12230a );
 a12232a <=( a12231a  and  a12226a );
 a12236a <=( A199  and  (not A166) );
 a12237a <=( A167  and  a12236a );
 a12241a <=( (not A203)  and  (not A201) );
 a12242a <=( (not A200)  and  a12241a );
 a12243a <=( a12242a  and  a12237a );
 a12247a <=( A298  and  A234 );
 a12248a <=( A233  and  a12247a );
 a12252a <=( A302  and  (not A301) );
 a12253a <=( (not A299)  and  a12252a );
 a12254a <=( a12253a  and  a12248a );
 a12258a <=( A199  and  (not A166) );
 a12259a <=( A167  and  a12258a );
 a12263a <=( (not A203)  and  (not A201) );
 a12264a <=( (not A200)  and  a12263a );
 a12265a <=( a12264a  and  a12259a );
 a12269a <=( (not A298)  and  A234 );
 a12270a <=( A233  and  a12269a );
 a12274a <=( A302  and  (not A301) );
 a12275a <=( A299  and  a12274a );
 a12276a <=( a12275a  and  a12270a );
 a12280a <=( A199  and  (not A166) );
 a12281a <=( A167  and  a12280a );
 a12285a <=( (not A203)  and  (not A201) );
 a12286a <=( (not A200)  and  a12285a );
 a12287a <=( a12286a  and  a12281a );
 a12291a <=( (not A298)  and  A234 );
 a12292a <=( A233  and  a12291a );
 a12296a <=( (not A302)  and  A301 );
 a12297a <=( (not A299)  and  a12296a );
 a12298a <=( a12297a  and  a12292a );
 a12302a <=( A199  and  (not A166) );
 a12303a <=( A167  and  a12302a );
 a12307a <=( (not A203)  and  (not A201) );
 a12308a <=( (not A200)  and  a12307a );
 a12309a <=( a12308a  and  a12303a );
 a12313a <=( A265  and  A234 );
 a12314a <=( A233  and  a12313a );
 a12318a <=( (not A269)  and  A268 );
 a12319a <=( A266  and  a12318a );
 a12320a <=( a12319a  and  a12314a );
 a12324a <=( A199  and  (not A166) );
 a12325a <=( A167  and  a12324a );
 a12329a <=( (not A203)  and  (not A201) );
 a12330a <=( (not A200)  and  a12329a );
 a12331a <=( a12330a  and  a12325a );
 a12335a <=( (not A265)  and  A234 );
 a12336a <=( A233  and  a12335a );
 a12340a <=( A269  and  (not A268) );
 a12341a <=( A266  and  a12340a );
 a12342a <=( a12341a  and  a12336a );
 a12346a <=( A199  and  (not A166) );
 a12347a <=( A167  and  a12346a );
 a12351a <=( (not A203)  and  (not A201) );
 a12352a <=( (not A200)  and  a12351a );
 a12353a <=( a12352a  and  a12347a );
 a12357a <=( A265  and  A234 );
 a12358a <=( A233  and  a12357a );
 a12362a <=( A269  and  (not A268) );
 a12363a <=( (not A266)  and  a12362a );
 a12364a <=( a12363a  and  a12358a );
 a12368a <=( A199  and  (not A166) );
 a12369a <=( A167  and  a12368a );
 a12373a <=( (not A203)  and  (not A201) );
 a12374a <=( (not A200)  and  a12373a );
 a12375a <=( a12374a  and  a12369a );
 a12379a <=( (not A265)  and  A234 );
 a12380a <=( A233  and  a12379a );
 a12384a <=( (not A269)  and  A268 );
 a12385a <=( (not A266)  and  a12384a );
 a12386a <=( a12385a  and  a12380a );
 a12390a <=( A199  and  (not A166) );
 a12391a <=( A167  and  a12390a );
 a12395a <=( (not A203)  and  (not A201) );
 a12396a <=( (not A200)  and  a12395a );
 a12397a <=( a12396a  and  a12391a );
 a12401a <=( A235  and  A233 );
 a12402a <=( A232  and  a12401a );
 a12406a <=( A300  and  A299 );
 a12407a <=( (not A236)  and  a12406a );
 a12408a <=( a12407a  and  a12402a );
 a12412a <=( A199  and  (not A166) );
 a12413a <=( A167  and  a12412a );
 a12417a <=( (not A203)  and  (not A201) );
 a12418a <=( (not A200)  and  a12417a );
 a12419a <=( a12418a  and  a12413a );
 a12423a <=( A235  and  A233 );
 a12424a <=( A232  and  a12423a );
 a12428a <=( A300  and  A298 );
 a12429a <=( (not A236)  and  a12428a );
 a12430a <=( a12429a  and  a12424a );
 a12434a <=( A199  and  (not A166) );
 a12435a <=( A167  and  a12434a );
 a12439a <=( (not A203)  and  (not A201) );
 a12440a <=( (not A200)  and  a12439a );
 a12441a <=( a12440a  and  a12435a );
 a12445a <=( A235  and  A233 );
 a12446a <=( A232  and  a12445a );
 a12450a <=( A267  and  A265 );
 a12451a <=( (not A236)  and  a12450a );
 a12452a <=( a12451a  and  a12446a );
 a12456a <=( A199  and  (not A166) );
 a12457a <=( A167  and  a12456a );
 a12461a <=( (not A203)  and  (not A201) );
 a12462a <=( (not A200)  and  a12461a );
 a12463a <=( a12462a  and  a12457a );
 a12467a <=( A235  and  A233 );
 a12468a <=( A232  and  a12467a );
 a12472a <=( A267  and  A266 );
 a12473a <=( (not A236)  and  a12472a );
 a12474a <=( a12473a  and  a12468a );
 a12478a <=( A199  and  (not A166) );
 a12479a <=( A167  and  a12478a );
 a12483a <=( (not A203)  and  (not A201) );
 a12484a <=( (not A200)  and  a12483a );
 a12485a <=( a12484a  and  a12479a );
 a12489a <=( (not A235)  and  A233 );
 a12490a <=( (not A232)  and  a12489a );
 a12494a <=( A300  and  A299 );
 a12495a <=( A236  and  a12494a );
 a12496a <=( a12495a  and  a12490a );
 a12500a <=( A199  and  (not A166) );
 a12501a <=( A167  and  a12500a );
 a12505a <=( (not A203)  and  (not A201) );
 a12506a <=( (not A200)  and  a12505a );
 a12507a <=( a12506a  and  a12501a );
 a12511a <=( (not A235)  and  A233 );
 a12512a <=( (not A232)  and  a12511a );
 a12516a <=( A300  and  A298 );
 a12517a <=( A236  and  a12516a );
 a12518a <=( a12517a  and  a12512a );
 a12522a <=( A199  and  (not A166) );
 a12523a <=( A167  and  a12522a );
 a12527a <=( (not A203)  and  (not A201) );
 a12528a <=( (not A200)  and  a12527a );
 a12529a <=( a12528a  and  a12523a );
 a12533a <=( (not A235)  and  A233 );
 a12534a <=( (not A232)  and  a12533a );
 a12538a <=( A267  and  A265 );
 a12539a <=( A236  and  a12538a );
 a12540a <=( a12539a  and  a12534a );
 a12544a <=( A199  and  (not A166) );
 a12545a <=( A167  and  a12544a );
 a12549a <=( (not A203)  and  (not A201) );
 a12550a <=( (not A200)  and  a12549a );
 a12551a <=( a12550a  and  a12545a );
 a12555a <=( (not A235)  and  A233 );
 a12556a <=( (not A232)  and  a12555a );
 a12560a <=( A267  and  A266 );
 a12561a <=( A236  and  a12560a );
 a12562a <=( a12561a  and  a12556a );
 a12566a <=( A199  and  (not A166) );
 a12567a <=( A167  and  a12566a );
 a12571a <=( (not A203)  and  (not A201) );
 a12572a <=( (not A200)  and  a12571a );
 a12573a <=( a12572a  and  a12567a );
 a12577a <=( (not A235)  and  (not A233) );
 a12578a <=( A232  and  a12577a );
 a12582a <=( A300  and  A299 );
 a12583a <=( A236  and  a12582a );
 a12584a <=( a12583a  and  a12578a );
 a12588a <=( A199  and  (not A166) );
 a12589a <=( A167  and  a12588a );
 a12593a <=( (not A203)  and  (not A201) );
 a12594a <=( (not A200)  and  a12593a );
 a12595a <=( a12594a  and  a12589a );
 a12599a <=( (not A235)  and  (not A233) );
 a12600a <=( A232  and  a12599a );
 a12604a <=( A300  and  A298 );
 a12605a <=( A236  and  a12604a );
 a12606a <=( a12605a  and  a12600a );
 a12610a <=( A199  and  (not A166) );
 a12611a <=( A167  and  a12610a );
 a12615a <=( (not A203)  and  (not A201) );
 a12616a <=( (not A200)  and  a12615a );
 a12617a <=( a12616a  and  a12611a );
 a12621a <=( (not A235)  and  (not A233) );
 a12622a <=( A232  and  a12621a );
 a12626a <=( A267  and  A265 );
 a12627a <=( A236  and  a12626a );
 a12628a <=( a12627a  and  a12622a );
 a12632a <=( A199  and  (not A166) );
 a12633a <=( A167  and  a12632a );
 a12637a <=( (not A203)  and  (not A201) );
 a12638a <=( (not A200)  and  a12637a );
 a12639a <=( a12638a  and  a12633a );
 a12643a <=( (not A235)  and  (not A233) );
 a12644a <=( A232  and  a12643a );
 a12648a <=( A267  and  A266 );
 a12649a <=( A236  and  a12648a );
 a12650a <=( a12649a  and  a12644a );
 a12654a <=( A199  and  (not A166) );
 a12655a <=( A167  and  a12654a );
 a12659a <=( (not A203)  and  (not A201) );
 a12660a <=( (not A200)  and  a12659a );
 a12661a <=( a12660a  and  a12655a );
 a12665a <=( A235  and  (not A233) );
 a12666a <=( (not A232)  and  a12665a );
 a12670a <=( A300  and  A299 );
 a12671a <=( (not A236)  and  a12670a );
 a12672a <=( a12671a  and  a12666a );
 a12676a <=( A199  and  (not A166) );
 a12677a <=( A167  and  a12676a );
 a12681a <=( (not A203)  and  (not A201) );
 a12682a <=( (not A200)  and  a12681a );
 a12683a <=( a12682a  and  a12677a );
 a12687a <=( A235  and  (not A233) );
 a12688a <=( (not A232)  and  a12687a );
 a12692a <=( A300  and  A298 );
 a12693a <=( (not A236)  and  a12692a );
 a12694a <=( a12693a  and  a12688a );
 a12698a <=( A199  and  (not A166) );
 a12699a <=( A167  and  a12698a );
 a12703a <=( (not A203)  and  (not A201) );
 a12704a <=( (not A200)  and  a12703a );
 a12705a <=( a12704a  and  a12699a );
 a12709a <=( A235  and  (not A233) );
 a12710a <=( (not A232)  and  a12709a );
 a12714a <=( A267  and  A265 );
 a12715a <=( (not A236)  and  a12714a );
 a12716a <=( a12715a  and  a12710a );
 a12720a <=( A199  and  (not A166) );
 a12721a <=( A167  and  a12720a );
 a12725a <=( (not A203)  and  (not A201) );
 a12726a <=( (not A200)  and  a12725a );
 a12727a <=( a12726a  and  a12721a );
 a12731a <=( A235  and  (not A233) );
 a12732a <=( (not A232)  and  a12731a );
 a12736a <=( A267  and  A266 );
 a12737a <=( (not A236)  and  a12736a );
 a12738a <=( a12737a  and  a12732a );
 a12742a <=( (not A167)  and  A168 );
 a12743a <=( A170  and  a12742a );
 a12747a <=( A200  and  A199 );
 a12748a <=( A166  and  a12747a );
 a12749a <=( a12748a  and  a12743a );
 a12753a <=( A232  and  (not A202) );
 a12754a <=( (not A201)  and  a12753a );
 a12758a <=( A300  and  A299 );
 a12759a <=( A234  and  a12758a );
 a12760a <=( a12759a  and  a12754a );
 a12764a <=( (not A167)  and  A168 );
 a12765a <=( A170  and  a12764a );
 a12769a <=( A200  and  A199 );
 a12770a <=( A166  and  a12769a );
 a12771a <=( a12770a  and  a12765a );
 a12775a <=( A232  and  (not A202) );
 a12776a <=( (not A201)  and  a12775a );
 a12780a <=( A300  and  A298 );
 a12781a <=( A234  and  a12780a );
 a12782a <=( a12781a  and  a12776a );
 a12786a <=( (not A167)  and  A168 );
 a12787a <=( A170  and  a12786a );
 a12791a <=( A200  and  A199 );
 a12792a <=( A166  and  a12791a );
 a12793a <=( a12792a  and  a12787a );
 a12797a <=( A232  and  (not A202) );
 a12798a <=( (not A201)  and  a12797a );
 a12802a <=( A267  and  A265 );
 a12803a <=( A234  and  a12802a );
 a12804a <=( a12803a  and  a12798a );
 a12808a <=( (not A167)  and  A168 );
 a12809a <=( A170  and  a12808a );
 a12813a <=( A200  and  A199 );
 a12814a <=( A166  and  a12813a );
 a12815a <=( a12814a  and  a12809a );
 a12819a <=( A232  and  (not A202) );
 a12820a <=( (not A201)  and  a12819a );
 a12824a <=( A267  and  A266 );
 a12825a <=( A234  and  a12824a );
 a12826a <=( a12825a  and  a12820a );
 a12830a <=( (not A167)  and  A168 );
 a12831a <=( A170  and  a12830a );
 a12835a <=( A200  and  A199 );
 a12836a <=( A166  and  a12835a );
 a12837a <=( a12836a  and  a12831a );
 a12841a <=( A233  and  (not A202) );
 a12842a <=( (not A201)  and  a12841a );
 a12846a <=( A300  and  A299 );
 a12847a <=( A234  and  a12846a );
 a12848a <=( a12847a  and  a12842a );
 a12852a <=( (not A167)  and  A168 );
 a12853a <=( A170  and  a12852a );
 a12857a <=( A200  and  A199 );
 a12858a <=( A166  and  a12857a );
 a12859a <=( a12858a  and  a12853a );
 a12863a <=( A233  and  (not A202) );
 a12864a <=( (not A201)  and  a12863a );
 a12868a <=( A300  and  A298 );
 a12869a <=( A234  and  a12868a );
 a12870a <=( a12869a  and  a12864a );
 a12874a <=( (not A167)  and  A168 );
 a12875a <=( A170  and  a12874a );
 a12879a <=( A200  and  A199 );
 a12880a <=( A166  and  a12879a );
 a12881a <=( a12880a  and  a12875a );
 a12885a <=( A233  and  (not A202) );
 a12886a <=( (not A201)  and  a12885a );
 a12890a <=( A267  and  A265 );
 a12891a <=( A234  and  a12890a );
 a12892a <=( a12891a  and  a12886a );
 a12896a <=( (not A167)  and  A168 );
 a12897a <=( A170  and  a12896a );
 a12901a <=( A200  and  A199 );
 a12902a <=( A166  and  a12901a );
 a12903a <=( a12902a  and  a12897a );
 a12907a <=( A233  and  (not A202) );
 a12908a <=( (not A201)  and  a12907a );
 a12912a <=( A267  and  A266 );
 a12913a <=( A234  and  a12912a );
 a12914a <=( a12913a  and  a12908a );
 a12918a <=( (not A167)  and  A168 );
 a12919a <=( A170  and  a12918a );
 a12923a <=( A200  and  A199 );
 a12924a <=( A166  and  a12923a );
 a12925a <=( a12924a  and  a12919a );
 a12929a <=( A232  and  A203 );
 a12930a <=( (not A201)  and  a12929a );
 a12934a <=( A300  and  A299 );
 a12935a <=( A234  and  a12934a );
 a12936a <=( a12935a  and  a12930a );
 a12940a <=( (not A167)  and  A168 );
 a12941a <=( A170  and  a12940a );
 a12945a <=( A200  and  A199 );
 a12946a <=( A166  and  a12945a );
 a12947a <=( a12946a  and  a12941a );
 a12951a <=( A232  and  A203 );
 a12952a <=( (not A201)  and  a12951a );
 a12956a <=( A300  and  A298 );
 a12957a <=( A234  and  a12956a );
 a12958a <=( a12957a  and  a12952a );
 a12962a <=( (not A167)  and  A168 );
 a12963a <=( A170  and  a12962a );
 a12967a <=( A200  and  A199 );
 a12968a <=( A166  and  a12967a );
 a12969a <=( a12968a  and  a12963a );
 a12973a <=( A232  and  A203 );
 a12974a <=( (not A201)  and  a12973a );
 a12978a <=( A267  and  A265 );
 a12979a <=( A234  and  a12978a );
 a12980a <=( a12979a  and  a12974a );
 a12984a <=( (not A167)  and  A168 );
 a12985a <=( A170  and  a12984a );
 a12989a <=( A200  and  A199 );
 a12990a <=( A166  and  a12989a );
 a12991a <=( a12990a  and  a12985a );
 a12995a <=( A232  and  A203 );
 a12996a <=( (not A201)  and  a12995a );
 a13000a <=( A267  and  A266 );
 a13001a <=( A234  and  a13000a );
 a13002a <=( a13001a  and  a12996a );
 a13006a <=( (not A167)  and  A168 );
 a13007a <=( A170  and  a13006a );
 a13011a <=( A200  and  A199 );
 a13012a <=( A166  and  a13011a );
 a13013a <=( a13012a  and  a13007a );
 a13017a <=( A233  and  A203 );
 a13018a <=( (not A201)  and  a13017a );
 a13022a <=( A300  and  A299 );
 a13023a <=( A234  and  a13022a );
 a13024a <=( a13023a  and  a13018a );
 a13028a <=( (not A167)  and  A168 );
 a13029a <=( A170  and  a13028a );
 a13033a <=( A200  and  A199 );
 a13034a <=( A166  and  a13033a );
 a13035a <=( a13034a  and  a13029a );
 a13039a <=( A233  and  A203 );
 a13040a <=( (not A201)  and  a13039a );
 a13044a <=( A300  and  A298 );
 a13045a <=( A234  and  a13044a );
 a13046a <=( a13045a  and  a13040a );
 a13050a <=( (not A167)  and  A168 );
 a13051a <=( A170  and  a13050a );
 a13055a <=( A200  and  A199 );
 a13056a <=( A166  and  a13055a );
 a13057a <=( a13056a  and  a13051a );
 a13061a <=( A233  and  A203 );
 a13062a <=( (not A201)  and  a13061a );
 a13066a <=( A267  and  A265 );
 a13067a <=( A234  and  a13066a );
 a13068a <=( a13067a  and  a13062a );
 a13072a <=( (not A167)  and  A168 );
 a13073a <=( A170  and  a13072a );
 a13077a <=( A200  and  A199 );
 a13078a <=( A166  and  a13077a );
 a13079a <=( a13078a  and  a13073a );
 a13083a <=( A233  and  A203 );
 a13084a <=( (not A201)  and  a13083a );
 a13088a <=( A267  and  A266 );
 a13089a <=( A234  and  a13088a );
 a13090a <=( a13089a  and  a13084a );
 a13094a <=( (not A167)  and  A168 );
 a13095a <=( A170  and  a13094a );
 a13099a <=( A200  and  (not A199) );
 a13100a <=( A166  and  a13099a );
 a13101a <=( a13100a  and  a13095a );
 a13105a <=( A232  and  A202 );
 a13106a <=( (not A201)  and  a13105a );
 a13110a <=( A300  and  A299 );
 a13111a <=( A234  and  a13110a );
 a13112a <=( a13111a  and  a13106a );
 a13116a <=( (not A167)  and  A168 );
 a13117a <=( A170  and  a13116a );
 a13121a <=( A200  and  (not A199) );
 a13122a <=( A166  and  a13121a );
 a13123a <=( a13122a  and  a13117a );
 a13127a <=( A232  and  A202 );
 a13128a <=( (not A201)  and  a13127a );
 a13132a <=( A300  and  A298 );
 a13133a <=( A234  and  a13132a );
 a13134a <=( a13133a  and  a13128a );
 a13138a <=( (not A167)  and  A168 );
 a13139a <=( A170  and  a13138a );
 a13143a <=( A200  and  (not A199) );
 a13144a <=( A166  and  a13143a );
 a13145a <=( a13144a  and  a13139a );
 a13149a <=( A232  and  A202 );
 a13150a <=( (not A201)  and  a13149a );
 a13154a <=( A267  and  A265 );
 a13155a <=( A234  and  a13154a );
 a13156a <=( a13155a  and  a13150a );
 a13160a <=( (not A167)  and  A168 );
 a13161a <=( A170  and  a13160a );
 a13165a <=( A200  and  (not A199) );
 a13166a <=( A166  and  a13165a );
 a13167a <=( a13166a  and  a13161a );
 a13171a <=( A232  and  A202 );
 a13172a <=( (not A201)  and  a13171a );
 a13176a <=( A267  and  A266 );
 a13177a <=( A234  and  a13176a );
 a13178a <=( a13177a  and  a13172a );
 a13182a <=( (not A167)  and  A168 );
 a13183a <=( A170  and  a13182a );
 a13187a <=( A200  and  (not A199) );
 a13188a <=( A166  and  a13187a );
 a13189a <=( a13188a  and  a13183a );
 a13193a <=( A233  and  A202 );
 a13194a <=( (not A201)  and  a13193a );
 a13198a <=( A300  and  A299 );
 a13199a <=( A234  and  a13198a );
 a13200a <=( a13199a  and  a13194a );
 a13204a <=( (not A167)  and  A168 );
 a13205a <=( A170  and  a13204a );
 a13209a <=( A200  and  (not A199) );
 a13210a <=( A166  and  a13209a );
 a13211a <=( a13210a  and  a13205a );
 a13215a <=( A233  and  A202 );
 a13216a <=( (not A201)  and  a13215a );
 a13220a <=( A300  and  A298 );
 a13221a <=( A234  and  a13220a );
 a13222a <=( a13221a  and  a13216a );
 a13226a <=( (not A167)  and  A168 );
 a13227a <=( A170  and  a13226a );
 a13231a <=( A200  and  (not A199) );
 a13232a <=( A166  and  a13231a );
 a13233a <=( a13232a  and  a13227a );
 a13237a <=( A233  and  A202 );
 a13238a <=( (not A201)  and  a13237a );
 a13242a <=( A267  and  A265 );
 a13243a <=( A234  and  a13242a );
 a13244a <=( a13243a  and  a13238a );
 a13248a <=( (not A167)  and  A168 );
 a13249a <=( A170  and  a13248a );
 a13253a <=( A200  and  (not A199) );
 a13254a <=( A166  and  a13253a );
 a13255a <=( a13254a  and  a13249a );
 a13259a <=( A233  and  A202 );
 a13260a <=( (not A201)  and  a13259a );
 a13264a <=( A267  and  A266 );
 a13265a <=( A234  and  a13264a );
 a13266a <=( a13265a  and  a13260a );
 a13270a <=( (not A167)  and  A168 );
 a13271a <=( A170  and  a13270a );
 a13275a <=( A200  and  (not A199) );
 a13276a <=( A166  and  a13275a );
 a13277a <=( a13276a  and  a13271a );
 a13281a <=( A232  and  (not A203) );
 a13282a <=( (not A201)  and  a13281a );
 a13286a <=( A300  and  A299 );
 a13287a <=( A234  and  a13286a );
 a13288a <=( a13287a  and  a13282a );
 a13292a <=( (not A167)  and  A168 );
 a13293a <=( A170  and  a13292a );
 a13297a <=( A200  and  (not A199) );
 a13298a <=( A166  and  a13297a );
 a13299a <=( a13298a  and  a13293a );
 a13303a <=( A232  and  (not A203) );
 a13304a <=( (not A201)  and  a13303a );
 a13308a <=( A300  and  A298 );
 a13309a <=( A234  and  a13308a );
 a13310a <=( a13309a  and  a13304a );
 a13314a <=( (not A167)  and  A168 );
 a13315a <=( A170  and  a13314a );
 a13319a <=( A200  and  (not A199) );
 a13320a <=( A166  and  a13319a );
 a13321a <=( a13320a  and  a13315a );
 a13325a <=( A232  and  (not A203) );
 a13326a <=( (not A201)  and  a13325a );
 a13330a <=( A267  and  A265 );
 a13331a <=( A234  and  a13330a );
 a13332a <=( a13331a  and  a13326a );
 a13336a <=( (not A167)  and  A168 );
 a13337a <=( A170  and  a13336a );
 a13341a <=( A200  and  (not A199) );
 a13342a <=( A166  and  a13341a );
 a13343a <=( a13342a  and  a13337a );
 a13347a <=( A232  and  (not A203) );
 a13348a <=( (not A201)  and  a13347a );
 a13352a <=( A267  and  A266 );
 a13353a <=( A234  and  a13352a );
 a13354a <=( a13353a  and  a13348a );
 a13358a <=( (not A167)  and  A168 );
 a13359a <=( A170  and  a13358a );
 a13363a <=( A200  and  (not A199) );
 a13364a <=( A166  and  a13363a );
 a13365a <=( a13364a  and  a13359a );
 a13369a <=( A233  and  (not A203) );
 a13370a <=( (not A201)  and  a13369a );
 a13374a <=( A300  and  A299 );
 a13375a <=( A234  and  a13374a );
 a13376a <=( a13375a  and  a13370a );
 a13380a <=( (not A167)  and  A168 );
 a13381a <=( A170  and  a13380a );
 a13385a <=( A200  and  (not A199) );
 a13386a <=( A166  and  a13385a );
 a13387a <=( a13386a  and  a13381a );
 a13391a <=( A233  and  (not A203) );
 a13392a <=( (not A201)  and  a13391a );
 a13396a <=( A300  and  A298 );
 a13397a <=( A234  and  a13396a );
 a13398a <=( a13397a  and  a13392a );
 a13402a <=( (not A167)  and  A168 );
 a13403a <=( A170  and  a13402a );
 a13407a <=( A200  and  (not A199) );
 a13408a <=( A166  and  a13407a );
 a13409a <=( a13408a  and  a13403a );
 a13413a <=( A233  and  (not A203) );
 a13414a <=( (not A201)  and  a13413a );
 a13418a <=( A267  and  A265 );
 a13419a <=( A234  and  a13418a );
 a13420a <=( a13419a  and  a13414a );
 a13424a <=( (not A167)  and  A168 );
 a13425a <=( A170  and  a13424a );
 a13429a <=( A200  and  (not A199) );
 a13430a <=( A166  and  a13429a );
 a13431a <=( a13430a  and  a13425a );
 a13435a <=( A233  and  (not A203) );
 a13436a <=( (not A201)  and  a13435a );
 a13440a <=( A267  and  A266 );
 a13441a <=( A234  and  a13440a );
 a13442a <=( a13441a  and  a13436a );
 a13446a <=( (not A167)  and  A168 );
 a13447a <=( A170  and  a13446a );
 a13451a <=( (not A200)  and  A199 );
 a13452a <=( A166  and  a13451a );
 a13453a <=( a13452a  and  a13447a );
 a13457a <=( A232  and  A202 );
 a13458a <=( (not A201)  and  a13457a );
 a13462a <=( A300  and  A299 );
 a13463a <=( A234  and  a13462a );
 a13464a <=( a13463a  and  a13458a );
 a13468a <=( (not A167)  and  A168 );
 a13469a <=( A170  and  a13468a );
 a13473a <=( (not A200)  and  A199 );
 a13474a <=( A166  and  a13473a );
 a13475a <=( a13474a  and  a13469a );
 a13479a <=( A232  and  A202 );
 a13480a <=( (not A201)  and  a13479a );
 a13484a <=( A300  and  A298 );
 a13485a <=( A234  and  a13484a );
 a13486a <=( a13485a  and  a13480a );
 a13490a <=( (not A167)  and  A168 );
 a13491a <=( A170  and  a13490a );
 a13495a <=( (not A200)  and  A199 );
 a13496a <=( A166  and  a13495a );
 a13497a <=( a13496a  and  a13491a );
 a13501a <=( A232  and  A202 );
 a13502a <=( (not A201)  and  a13501a );
 a13506a <=( A267  and  A265 );
 a13507a <=( A234  and  a13506a );
 a13508a <=( a13507a  and  a13502a );
 a13512a <=( (not A167)  and  A168 );
 a13513a <=( A170  and  a13512a );
 a13517a <=( (not A200)  and  A199 );
 a13518a <=( A166  and  a13517a );
 a13519a <=( a13518a  and  a13513a );
 a13523a <=( A232  and  A202 );
 a13524a <=( (not A201)  and  a13523a );
 a13528a <=( A267  and  A266 );
 a13529a <=( A234  and  a13528a );
 a13530a <=( a13529a  and  a13524a );
 a13534a <=( (not A167)  and  A168 );
 a13535a <=( A170  and  a13534a );
 a13539a <=( (not A200)  and  A199 );
 a13540a <=( A166  and  a13539a );
 a13541a <=( a13540a  and  a13535a );
 a13545a <=( A233  and  A202 );
 a13546a <=( (not A201)  and  a13545a );
 a13550a <=( A300  and  A299 );
 a13551a <=( A234  and  a13550a );
 a13552a <=( a13551a  and  a13546a );
 a13556a <=( (not A167)  and  A168 );
 a13557a <=( A170  and  a13556a );
 a13561a <=( (not A200)  and  A199 );
 a13562a <=( A166  and  a13561a );
 a13563a <=( a13562a  and  a13557a );
 a13567a <=( A233  and  A202 );
 a13568a <=( (not A201)  and  a13567a );
 a13572a <=( A300  and  A298 );
 a13573a <=( A234  and  a13572a );
 a13574a <=( a13573a  and  a13568a );
 a13578a <=( (not A167)  and  A168 );
 a13579a <=( A170  and  a13578a );
 a13583a <=( (not A200)  and  A199 );
 a13584a <=( A166  and  a13583a );
 a13585a <=( a13584a  and  a13579a );
 a13589a <=( A233  and  A202 );
 a13590a <=( (not A201)  and  a13589a );
 a13594a <=( A267  and  A265 );
 a13595a <=( A234  and  a13594a );
 a13596a <=( a13595a  and  a13590a );
 a13600a <=( (not A167)  and  A168 );
 a13601a <=( A170  and  a13600a );
 a13605a <=( (not A200)  and  A199 );
 a13606a <=( A166  and  a13605a );
 a13607a <=( a13606a  and  a13601a );
 a13611a <=( A233  and  A202 );
 a13612a <=( (not A201)  and  a13611a );
 a13616a <=( A267  and  A266 );
 a13617a <=( A234  and  a13616a );
 a13618a <=( a13617a  and  a13612a );
 a13622a <=( (not A167)  and  A168 );
 a13623a <=( A170  and  a13622a );
 a13627a <=( (not A200)  and  A199 );
 a13628a <=( A166  and  a13627a );
 a13629a <=( a13628a  and  a13623a );
 a13633a <=( A232  and  (not A203) );
 a13634a <=( (not A201)  and  a13633a );
 a13638a <=( A300  and  A299 );
 a13639a <=( A234  and  a13638a );
 a13640a <=( a13639a  and  a13634a );
 a13644a <=( (not A167)  and  A168 );
 a13645a <=( A170  and  a13644a );
 a13649a <=( (not A200)  and  A199 );
 a13650a <=( A166  and  a13649a );
 a13651a <=( a13650a  and  a13645a );
 a13655a <=( A232  and  (not A203) );
 a13656a <=( (not A201)  and  a13655a );
 a13660a <=( A300  and  A298 );
 a13661a <=( A234  and  a13660a );
 a13662a <=( a13661a  and  a13656a );
 a13666a <=( (not A167)  and  A168 );
 a13667a <=( A170  and  a13666a );
 a13671a <=( (not A200)  and  A199 );
 a13672a <=( A166  and  a13671a );
 a13673a <=( a13672a  and  a13667a );
 a13677a <=( A232  and  (not A203) );
 a13678a <=( (not A201)  and  a13677a );
 a13682a <=( A267  and  A265 );
 a13683a <=( A234  and  a13682a );
 a13684a <=( a13683a  and  a13678a );
 a13688a <=( (not A167)  and  A168 );
 a13689a <=( A170  and  a13688a );
 a13693a <=( (not A200)  and  A199 );
 a13694a <=( A166  and  a13693a );
 a13695a <=( a13694a  and  a13689a );
 a13699a <=( A232  and  (not A203) );
 a13700a <=( (not A201)  and  a13699a );
 a13704a <=( A267  and  A266 );
 a13705a <=( A234  and  a13704a );
 a13706a <=( a13705a  and  a13700a );
 a13710a <=( (not A167)  and  A168 );
 a13711a <=( A170  and  a13710a );
 a13715a <=( (not A200)  and  A199 );
 a13716a <=( A166  and  a13715a );
 a13717a <=( a13716a  and  a13711a );
 a13721a <=( A233  and  (not A203) );
 a13722a <=( (not A201)  and  a13721a );
 a13726a <=( A300  and  A299 );
 a13727a <=( A234  and  a13726a );
 a13728a <=( a13727a  and  a13722a );
 a13732a <=( (not A167)  and  A168 );
 a13733a <=( A170  and  a13732a );
 a13737a <=( (not A200)  and  A199 );
 a13738a <=( A166  and  a13737a );
 a13739a <=( a13738a  and  a13733a );
 a13743a <=( A233  and  (not A203) );
 a13744a <=( (not A201)  and  a13743a );
 a13748a <=( A300  and  A298 );
 a13749a <=( A234  and  a13748a );
 a13750a <=( a13749a  and  a13744a );
 a13754a <=( (not A167)  and  A168 );
 a13755a <=( A170  and  a13754a );
 a13759a <=( (not A200)  and  A199 );
 a13760a <=( A166  and  a13759a );
 a13761a <=( a13760a  and  a13755a );
 a13765a <=( A233  and  (not A203) );
 a13766a <=( (not A201)  and  a13765a );
 a13770a <=( A267  and  A265 );
 a13771a <=( A234  and  a13770a );
 a13772a <=( a13771a  and  a13766a );
 a13776a <=( (not A167)  and  A168 );
 a13777a <=( A170  and  a13776a );
 a13781a <=( (not A200)  and  A199 );
 a13782a <=( A166  and  a13781a );
 a13783a <=( a13782a  and  a13777a );
 a13787a <=( A233  and  (not A203) );
 a13788a <=( (not A201)  and  a13787a );
 a13792a <=( A267  and  A266 );
 a13793a <=( A234  and  a13792a );
 a13794a <=( a13793a  and  a13788a );
 a13798a <=( (not A167)  and  A168 );
 a13799a <=( A169  and  a13798a );
 a13803a <=( A200  and  A199 );
 a13804a <=( A166  and  a13803a );
 a13805a <=( a13804a  and  a13799a );
 a13809a <=( A232  and  (not A202) );
 a13810a <=( (not A201)  and  a13809a );
 a13814a <=( A300  and  A299 );
 a13815a <=( A234  and  a13814a );
 a13816a <=( a13815a  and  a13810a );
 a13820a <=( (not A167)  and  A168 );
 a13821a <=( A169  and  a13820a );
 a13825a <=( A200  and  A199 );
 a13826a <=( A166  and  a13825a );
 a13827a <=( a13826a  and  a13821a );
 a13831a <=( A232  and  (not A202) );
 a13832a <=( (not A201)  and  a13831a );
 a13836a <=( A300  and  A298 );
 a13837a <=( A234  and  a13836a );
 a13838a <=( a13837a  and  a13832a );
 a13842a <=( (not A167)  and  A168 );
 a13843a <=( A169  and  a13842a );
 a13847a <=( A200  and  A199 );
 a13848a <=( A166  and  a13847a );
 a13849a <=( a13848a  and  a13843a );
 a13853a <=( A232  and  (not A202) );
 a13854a <=( (not A201)  and  a13853a );
 a13858a <=( A267  and  A265 );
 a13859a <=( A234  and  a13858a );
 a13860a <=( a13859a  and  a13854a );
 a13864a <=( (not A167)  and  A168 );
 a13865a <=( A169  and  a13864a );
 a13869a <=( A200  and  A199 );
 a13870a <=( A166  and  a13869a );
 a13871a <=( a13870a  and  a13865a );
 a13875a <=( A232  and  (not A202) );
 a13876a <=( (not A201)  and  a13875a );
 a13880a <=( A267  and  A266 );
 a13881a <=( A234  and  a13880a );
 a13882a <=( a13881a  and  a13876a );
 a13886a <=( (not A167)  and  A168 );
 a13887a <=( A169  and  a13886a );
 a13891a <=( A200  and  A199 );
 a13892a <=( A166  and  a13891a );
 a13893a <=( a13892a  and  a13887a );
 a13897a <=( A233  and  (not A202) );
 a13898a <=( (not A201)  and  a13897a );
 a13902a <=( A300  and  A299 );
 a13903a <=( A234  and  a13902a );
 a13904a <=( a13903a  and  a13898a );
 a13908a <=( (not A167)  and  A168 );
 a13909a <=( A169  and  a13908a );
 a13913a <=( A200  and  A199 );
 a13914a <=( A166  and  a13913a );
 a13915a <=( a13914a  and  a13909a );
 a13919a <=( A233  and  (not A202) );
 a13920a <=( (not A201)  and  a13919a );
 a13924a <=( A300  and  A298 );
 a13925a <=( A234  and  a13924a );
 a13926a <=( a13925a  and  a13920a );
 a13930a <=( (not A167)  and  A168 );
 a13931a <=( A169  and  a13930a );
 a13935a <=( A200  and  A199 );
 a13936a <=( A166  and  a13935a );
 a13937a <=( a13936a  and  a13931a );
 a13941a <=( A233  and  (not A202) );
 a13942a <=( (not A201)  and  a13941a );
 a13946a <=( A267  and  A265 );
 a13947a <=( A234  and  a13946a );
 a13948a <=( a13947a  and  a13942a );
 a13952a <=( (not A167)  and  A168 );
 a13953a <=( A169  and  a13952a );
 a13957a <=( A200  and  A199 );
 a13958a <=( A166  and  a13957a );
 a13959a <=( a13958a  and  a13953a );
 a13963a <=( A233  and  (not A202) );
 a13964a <=( (not A201)  and  a13963a );
 a13968a <=( A267  and  A266 );
 a13969a <=( A234  and  a13968a );
 a13970a <=( a13969a  and  a13964a );
 a13974a <=( (not A167)  and  A168 );
 a13975a <=( A169  and  a13974a );
 a13979a <=( A200  and  A199 );
 a13980a <=( A166  and  a13979a );
 a13981a <=( a13980a  and  a13975a );
 a13985a <=( A232  and  A203 );
 a13986a <=( (not A201)  and  a13985a );
 a13990a <=( A300  and  A299 );
 a13991a <=( A234  and  a13990a );
 a13992a <=( a13991a  and  a13986a );
 a13996a <=( (not A167)  and  A168 );
 a13997a <=( A169  and  a13996a );
 a14001a <=( A200  and  A199 );
 a14002a <=( A166  and  a14001a );
 a14003a <=( a14002a  and  a13997a );
 a14007a <=( A232  and  A203 );
 a14008a <=( (not A201)  and  a14007a );
 a14012a <=( A300  and  A298 );
 a14013a <=( A234  and  a14012a );
 a14014a <=( a14013a  and  a14008a );
 a14018a <=( (not A167)  and  A168 );
 a14019a <=( A169  and  a14018a );
 a14023a <=( A200  and  A199 );
 a14024a <=( A166  and  a14023a );
 a14025a <=( a14024a  and  a14019a );
 a14029a <=( A232  and  A203 );
 a14030a <=( (not A201)  and  a14029a );
 a14034a <=( A267  and  A265 );
 a14035a <=( A234  and  a14034a );
 a14036a <=( a14035a  and  a14030a );
 a14040a <=( (not A167)  and  A168 );
 a14041a <=( A169  and  a14040a );
 a14045a <=( A200  and  A199 );
 a14046a <=( A166  and  a14045a );
 a14047a <=( a14046a  and  a14041a );
 a14051a <=( A232  and  A203 );
 a14052a <=( (not A201)  and  a14051a );
 a14056a <=( A267  and  A266 );
 a14057a <=( A234  and  a14056a );
 a14058a <=( a14057a  and  a14052a );
 a14062a <=( (not A167)  and  A168 );
 a14063a <=( A169  and  a14062a );
 a14067a <=( A200  and  A199 );
 a14068a <=( A166  and  a14067a );
 a14069a <=( a14068a  and  a14063a );
 a14073a <=( A233  and  A203 );
 a14074a <=( (not A201)  and  a14073a );
 a14078a <=( A300  and  A299 );
 a14079a <=( A234  and  a14078a );
 a14080a <=( a14079a  and  a14074a );
 a14084a <=( (not A167)  and  A168 );
 a14085a <=( A169  and  a14084a );
 a14089a <=( A200  and  A199 );
 a14090a <=( A166  and  a14089a );
 a14091a <=( a14090a  and  a14085a );
 a14095a <=( A233  and  A203 );
 a14096a <=( (not A201)  and  a14095a );
 a14100a <=( A300  and  A298 );
 a14101a <=( A234  and  a14100a );
 a14102a <=( a14101a  and  a14096a );
 a14106a <=( (not A167)  and  A168 );
 a14107a <=( A169  and  a14106a );
 a14111a <=( A200  and  A199 );
 a14112a <=( A166  and  a14111a );
 a14113a <=( a14112a  and  a14107a );
 a14117a <=( A233  and  A203 );
 a14118a <=( (not A201)  and  a14117a );
 a14122a <=( A267  and  A265 );
 a14123a <=( A234  and  a14122a );
 a14124a <=( a14123a  and  a14118a );
 a14128a <=( (not A167)  and  A168 );
 a14129a <=( A169  and  a14128a );
 a14133a <=( A200  and  A199 );
 a14134a <=( A166  and  a14133a );
 a14135a <=( a14134a  and  a14129a );
 a14139a <=( A233  and  A203 );
 a14140a <=( (not A201)  and  a14139a );
 a14144a <=( A267  and  A266 );
 a14145a <=( A234  and  a14144a );
 a14146a <=( a14145a  and  a14140a );
 a14150a <=( (not A167)  and  A168 );
 a14151a <=( A169  and  a14150a );
 a14155a <=( A200  and  (not A199) );
 a14156a <=( A166  and  a14155a );
 a14157a <=( a14156a  and  a14151a );
 a14161a <=( A232  and  A202 );
 a14162a <=( (not A201)  and  a14161a );
 a14166a <=( A300  and  A299 );
 a14167a <=( A234  and  a14166a );
 a14168a <=( a14167a  and  a14162a );
 a14172a <=( (not A167)  and  A168 );
 a14173a <=( A169  and  a14172a );
 a14177a <=( A200  and  (not A199) );
 a14178a <=( A166  and  a14177a );
 a14179a <=( a14178a  and  a14173a );
 a14183a <=( A232  and  A202 );
 a14184a <=( (not A201)  and  a14183a );
 a14188a <=( A300  and  A298 );
 a14189a <=( A234  and  a14188a );
 a14190a <=( a14189a  and  a14184a );
 a14194a <=( (not A167)  and  A168 );
 a14195a <=( A169  and  a14194a );
 a14199a <=( A200  and  (not A199) );
 a14200a <=( A166  and  a14199a );
 a14201a <=( a14200a  and  a14195a );
 a14205a <=( A232  and  A202 );
 a14206a <=( (not A201)  and  a14205a );
 a14210a <=( A267  and  A265 );
 a14211a <=( A234  and  a14210a );
 a14212a <=( a14211a  and  a14206a );
 a14216a <=( (not A167)  and  A168 );
 a14217a <=( A169  and  a14216a );
 a14221a <=( A200  and  (not A199) );
 a14222a <=( A166  and  a14221a );
 a14223a <=( a14222a  and  a14217a );
 a14227a <=( A232  and  A202 );
 a14228a <=( (not A201)  and  a14227a );
 a14232a <=( A267  and  A266 );
 a14233a <=( A234  and  a14232a );
 a14234a <=( a14233a  and  a14228a );
 a14238a <=( (not A167)  and  A168 );
 a14239a <=( A169  and  a14238a );
 a14243a <=( A200  and  (not A199) );
 a14244a <=( A166  and  a14243a );
 a14245a <=( a14244a  and  a14239a );
 a14249a <=( A233  and  A202 );
 a14250a <=( (not A201)  and  a14249a );
 a14254a <=( A300  and  A299 );
 a14255a <=( A234  and  a14254a );
 a14256a <=( a14255a  and  a14250a );
 a14260a <=( (not A167)  and  A168 );
 a14261a <=( A169  and  a14260a );
 a14265a <=( A200  and  (not A199) );
 a14266a <=( A166  and  a14265a );
 a14267a <=( a14266a  and  a14261a );
 a14271a <=( A233  and  A202 );
 a14272a <=( (not A201)  and  a14271a );
 a14276a <=( A300  and  A298 );
 a14277a <=( A234  and  a14276a );
 a14278a <=( a14277a  and  a14272a );
 a14282a <=( (not A167)  and  A168 );
 a14283a <=( A169  and  a14282a );
 a14287a <=( A200  and  (not A199) );
 a14288a <=( A166  and  a14287a );
 a14289a <=( a14288a  and  a14283a );
 a14293a <=( A233  and  A202 );
 a14294a <=( (not A201)  and  a14293a );
 a14298a <=( A267  and  A265 );
 a14299a <=( A234  and  a14298a );
 a14300a <=( a14299a  and  a14294a );
 a14304a <=( (not A167)  and  A168 );
 a14305a <=( A169  and  a14304a );
 a14309a <=( A200  and  (not A199) );
 a14310a <=( A166  and  a14309a );
 a14311a <=( a14310a  and  a14305a );
 a14315a <=( A233  and  A202 );
 a14316a <=( (not A201)  and  a14315a );
 a14320a <=( A267  and  A266 );
 a14321a <=( A234  and  a14320a );
 a14322a <=( a14321a  and  a14316a );
 a14326a <=( (not A167)  and  A168 );
 a14327a <=( A169  and  a14326a );
 a14331a <=( A200  and  (not A199) );
 a14332a <=( A166  and  a14331a );
 a14333a <=( a14332a  and  a14327a );
 a14337a <=( A232  and  (not A203) );
 a14338a <=( (not A201)  and  a14337a );
 a14342a <=( A300  and  A299 );
 a14343a <=( A234  and  a14342a );
 a14344a <=( a14343a  and  a14338a );
 a14348a <=( (not A167)  and  A168 );
 a14349a <=( A169  and  a14348a );
 a14353a <=( A200  and  (not A199) );
 a14354a <=( A166  and  a14353a );
 a14355a <=( a14354a  and  a14349a );
 a14359a <=( A232  and  (not A203) );
 a14360a <=( (not A201)  and  a14359a );
 a14364a <=( A300  and  A298 );
 a14365a <=( A234  and  a14364a );
 a14366a <=( a14365a  and  a14360a );
 a14370a <=( (not A167)  and  A168 );
 a14371a <=( A169  and  a14370a );
 a14375a <=( A200  and  (not A199) );
 a14376a <=( A166  and  a14375a );
 a14377a <=( a14376a  and  a14371a );
 a14381a <=( A232  and  (not A203) );
 a14382a <=( (not A201)  and  a14381a );
 a14386a <=( A267  and  A265 );
 a14387a <=( A234  and  a14386a );
 a14388a <=( a14387a  and  a14382a );
 a14392a <=( (not A167)  and  A168 );
 a14393a <=( A169  and  a14392a );
 a14397a <=( A200  and  (not A199) );
 a14398a <=( A166  and  a14397a );
 a14399a <=( a14398a  and  a14393a );
 a14403a <=( A232  and  (not A203) );
 a14404a <=( (not A201)  and  a14403a );
 a14408a <=( A267  and  A266 );
 a14409a <=( A234  and  a14408a );
 a14410a <=( a14409a  and  a14404a );
 a14414a <=( (not A167)  and  A168 );
 a14415a <=( A169  and  a14414a );
 a14419a <=( A200  and  (not A199) );
 a14420a <=( A166  and  a14419a );
 a14421a <=( a14420a  and  a14415a );
 a14425a <=( A233  and  (not A203) );
 a14426a <=( (not A201)  and  a14425a );
 a14430a <=( A300  and  A299 );
 a14431a <=( A234  and  a14430a );
 a14432a <=( a14431a  and  a14426a );
 a14436a <=( (not A167)  and  A168 );
 a14437a <=( A169  and  a14436a );
 a14441a <=( A200  and  (not A199) );
 a14442a <=( A166  and  a14441a );
 a14443a <=( a14442a  and  a14437a );
 a14447a <=( A233  and  (not A203) );
 a14448a <=( (not A201)  and  a14447a );
 a14452a <=( A300  and  A298 );
 a14453a <=( A234  and  a14452a );
 a14454a <=( a14453a  and  a14448a );
 a14458a <=( (not A167)  and  A168 );
 a14459a <=( A169  and  a14458a );
 a14463a <=( A200  and  (not A199) );
 a14464a <=( A166  and  a14463a );
 a14465a <=( a14464a  and  a14459a );
 a14469a <=( A233  and  (not A203) );
 a14470a <=( (not A201)  and  a14469a );
 a14474a <=( A267  and  A265 );
 a14475a <=( A234  and  a14474a );
 a14476a <=( a14475a  and  a14470a );
 a14480a <=( (not A167)  and  A168 );
 a14481a <=( A169  and  a14480a );
 a14485a <=( A200  and  (not A199) );
 a14486a <=( A166  and  a14485a );
 a14487a <=( a14486a  and  a14481a );
 a14491a <=( A233  and  (not A203) );
 a14492a <=( (not A201)  and  a14491a );
 a14496a <=( A267  and  A266 );
 a14497a <=( A234  and  a14496a );
 a14498a <=( a14497a  and  a14492a );
 a14502a <=( (not A167)  and  A168 );
 a14503a <=( A169  and  a14502a );
 a14507a <=( (not A200)  and  A199 );
 a14508a <=( A166  and  a14507a );
 a14509a <=( a14508a  and  a14503a );
 a14513a <=( A232  and  A202 );
 a14514a <=( (not A201)  and  a14513a );
 a14518a <=( A300  and  A299 );
 a14519a <=( A234  and  a14518a );
 a14520a <=( a14519a  and  a14514a );
 a14524a <=( (not A167)  and  A168 );
 a14525a <=( A169  and  a14524a );
 a14529a <=( (not A200)  and  A199 );
 a14530a <=( A166  and  a14529a );
 a14531a <=( a14530a  and  a14525a );
 a14535a <=( A232  and  A202 );
 a14536a <=( (not A201)  and  a14535a );
 a14540a <=( A300  and  A298 );
 a14541a <=( A234  and  a14540a );
 a14542a <=( a14541a  and  a14536a );
 a14546a <=( (not A167)  and  A168 );
 a14547a <=( A169  and  a14546a );
 a14551a <=( (not A200)  and  A199 );
 a14552a <=( A166  and  a14551a );
 a14553a <=( a14552a  and  a14547a );
 a14557a <=( A232  and  A202 );
 a14558a <=( (not A201)  and  a14557a );
 a14562a <=( A267  and  A265 );
 a14563a <=( A234  and  a14562a );
 a14564a <=( a14563a  and  a14558a );
 a14568a <=( (not A167)  and  A168 );
 a14569a <=( A169  and  a14568a );
 a14573a <=( (not A200)  and  A199 );
 a14574a <=( A166  and  a14573a );
 a14575a <=( a14574a  and  a14569a );
 a14579a <=( A232  and  A202 );
 a14580a <=( (not A201)  and  a14579a );
 a14584a <=( A267  and  A266 );
 a14585a <=( A234  and  a14584a );
 a14586a <=( a14585a  and  a14580a );
 a14590a <=( (not A167)  and  A168 );
 a14591a <=( A169  and  a14590a );
 a14595a <=( (not A200)  and  A199 );
 a14596a <=( A166  and  a14595a );
 a14597a <=( a14596a  and  a14591a );
 a14601a <=( A233  and  A202 );
 a14602a <=( (not A201)  and  a14601a );
 a14606a <=( A300  and  A299 );
 a14607a <=( A234  and  a14606a );
 a14608a <=( a14607a  and  a14602a );
 a14612a <=( (not A167)  and  A168 );
 a14613a <=( A169  and  a14612a );
 a14617a <=( (not A200)  and  A199 );
 a14618a <=( A166  and  a14617a );
 a14619a <=( a14618a  and  a14613a );
 a14623a <=( A233  and  A202 );
 a14624a <=( (not A201)  and  a14623a );
 a14628a <=( A300  and  A298 );
 a14629a <=( A234  and  a14628a );
 a14630a <=( a14629a  and  a14624a );
 a14634a <=( (not A167)  and  A168 );
 a14635a <=( A169  and  a14634a );
 a14639a <=( (not A200)  and  A199 );
 a14640a <=( A166  and  a14639a );
 a14641a <=( a14640a  and  a14635a );
 a14645a <=( A233  and  A202 );
 a14646a <=( (not A201)  and  a14645a );
 a14650a <=( A267  and  A265 );
 a14651a <=( A234  and  a14650a );
 a14652a <=( a14651a  and  a14646a );
 a14656a <=( (not A167)  and  A168 );
 a14657a <=( A169  and  a14656a );
 a14661a <=( (not A200)  and  A199 );
 a14662a <=( A166  and  a14661a );
 a14663a <=( a14662a  and  a14657a );
 a14667a <=( A233  and  A202 );
 a14668a <=( (not A201)  and  a14667a );
 a14672a <=( A267  and  A266 );
 a14673a <=( A234  and  a14672a );
 a14674a <=( a14673a  and  a14668a );
 a14678a <=( (not A167)  and  A168 );
 a14679a <=( A169  and  a14678a );
 a14683a <=( (not A200)  and  A199 );
 a14684a <=( A166  and  a14683a );
 a14685a <=( a14684a  and  a14679a );
 a14689a <=( A232  and  (not A203) );
 a14690a <=( (not A201)  and  a14689a );
 a14694a <=( A300  and  A299 );
 a14695a <=( A234  and  a14694a );
 a14696a <=( a14695a  and  a14690a );
 a14700a <=( (not A167)  and  A168 );
 a14701a <=( A169  and  a14700a );
 a14705a <=( (not A200)  and  A199 );
 a14706a <=( A166  and  a14705a );
 a14707a <=( a14706a  and  a14701a );
 a14711a <=( A232  and  (not A203) );
 a14712a <=( (not A201)  and  a14711a );
 a14716a <=( A300  and  A298 );
 a14717a <=( A234  and  a14716a );
 a14718a <=( a14717a  and  a14712a );
 a14722a <=( (not A167)  and  A168 );
 a14723a <=( A169  and  a14722a );
 a14727a <=( (not A200)  and  A199 );
 a14728a <=( A166  and  a14727a );
 a14729a <=( a14728a  and  a14723a );
 a14733a <=( A232  and  (not A203) );
 a14734a <=( (not A201)  and  a14733a );
 a14738a <=( A267  and  A265 );
 a14739a <=( A234  and  a14738a );
 a14740a <=( a14739a  and  a14734a );
 a14744a <=( (not A167)  and  A168 );
 a14745a <=( A169  and  a14744a );
 a14749a <=( (not A200)  and  A199 );
 a14750a <=( A166  and  a14749a );
 a14751a <=( a14750a  and  a14745a );
 a14755a <=( A232  and  (not A203) );
 a14756a <=( (not A201)  and  a14755a );
 a14760a <=( A267  and  A266 );
 a14761a <=( A234  and  a14760a );
 a14762a <=( a14761a  and  a14756a );
 a14766a <=( (not A167)  and  A168 );
 a14767a <=( A169  and  a14766a );
 a14771a <=( (not A200)  and  A199 );
 a14772a <=( A166  and  a14771a );
 a14773a <=( a14772a  and  a14767a );
 a14777a <=( A233  and  (not A203) );
 a14778a <=( (not A201)  and  a14777a );
 a14782a <=( A300  and  A299 );
 a14783a <=( A234  and  a14782a );
 a14784a <=( a14783a  and  a14778a );
 a14788a <=( (not A167)  and  A168 );
 a14789a <=( A169  and  a14788a );
 a14793a <=( (not A200)  and  A199 );
 a14794a <=( A166  and  a14793a );
 a14795a <=( a14794a  and  a14789a );
 a14799a <=( A233  and  (not A203) );
 a14800a <=( (not A201)  and  a14799a );
 a14804a <=( A300  and  A298 );
 a14805a <=( A234  and  a14804a );
 a14806a <=( a14805a  and  a14800a );
 a14810a <=( (not A167)  and  A168 );
 a14811a <=( A169  and  a14810a );
 a14815a <=( (not A200)  and  A199 );
 a14816a <=( A166  and  a14815a );
 a14817a <=( a14816a  and  a14811a );
 a14821a <=( A233  and  (not A203) );
 a14822a <=( (not A201)  and  a14821a );
 a14826a <=( A267  and  A265 );
 a14827a <=( A234  and  a14826a );
 a14828a <=( a14827a  and  a14822a );
 a14832a <=( (not A167)  and  A168 );
 a14833a <=( A169  and  a14832a );
 a14837a <=( (not A200)  and  A199 );
 a14838a <=( A166  and  a14837a );
 a14839a <=( a14838a  and  a14833a );
 a14843a <=( A233  and  (not A203) );
 a14844a <=( (not A201)  and  a14843a );
 a14848a <=( A267  and  A266 );
 a14849a <=( A234  and  a14848a );
 a14850a <=( a14849a  and  a14844a );
 a14854a <=( (not A199)  and  (not A166) );
 a14855a <=( A167  and  a14854a );
 a14859a <=( A232  and  (not A202) );
 a14860a <=( (not A200)  and  a14859a );
 a14861a <=( a14860a  and  a14855a );
 a14865a <=( (not A236)  and  A235 );
 a14866a <=( A233  and  a14865a );
 a14869a <=( A299  and  A298 );
 a14872a <=( (not A302)  and  A301 );
 a14873a <=( a14872a  and  a14869a );
 a14874a <=( a14873a  and  a14866a );
 a14878a <=( (not A199)  and  (not A166) );
 a14879a <=( A167  and  a14878a );
 a14883a <=( A232  and  (not A202) );
 a14884a <=( (not A200)  and  a14883a );
 a14885a <=( a14884a  and  a14879a );
 a14889a <=( (not A236)  and  A235 );
 a14890a <=( A233  and  a14889a );
 a14893a <=( (not A299)  and  A298 );
 a14896a <=( A302  and  (not A301) );
 a14897a <=( a14896a  and  a14893a );
 a14898a <=( a14897a  and  a14890a );
 a14902a <=( (not A199)  and  (not A166) );
 a14903a <=( A167  and  a14902a );
 a14907a <=( A232  and  (not A202) );
 a14908a <=( (not A200)  and  a14907a );
 a14909a <=( a14908a  and  a14903a );
 a14913a <=( (not A236)  and  A235 );
 a14914a <=( A233  and  a14913a );
 a14917a <=( A299  and  (not A298) );
 a14920a <=( A302  and  (not A301) );
 a14921a <=( a14920a  and  a14917a );
 a14922a <=( a14921a  and  a14914a );
 a14926a <=( (not A199)  and  (not A166) );
 a14927a <=( A167  and  a14926a );
 a14931a <=( A232  and  (not A202) );
 a14932a <=( (not A200)  and  a14931a );
 a14933a <=( a14932a  and  a14927a );
 a14937a <=( (not A236)  and  A235 );
 a14938a <=( A233  and  a14937a );
 a14941a <=( (not A299)  and  (not A298) );
 a14944a <=( (not A302)  and  A301 );
 a14945a <=( a14944a  and  a14941a );
 a14946a <=( a14945a  and  a14938a );
 a14950a <=( (not A199)  and  (not A166) );
 a14951a <=( A167  and  a14950a );
 a14955a <=( A232  and  (not A202) );
 a14956a <=( (not A200)  and  a14955a );
 a14957a <=( a14956a  and  a14951a );
 a14961a <=( (not A236)  and  A235 );
 a14962a <=( A233  and  a14961a );
 a14965a <=( A266  and  A265 );
 a14968a <=( (not A269)  and  A268 );
 a14969a <=( a14968a  and  a14965a );
 a14970a <=( a14969a  and  a14962a );
 a14974a <=( (not A199)  and  (not A166) );
 a14975a <=( A167  and  a14974a );
 a14979a <=( A232  and  (not A202) );
 a14980a <=( (not A200)  and  a14979a );
 a14981a <=( a14980a  and  a14975a );
 a14985a <=( (not A236)  and  A235 );
 a14986a <=( A233  and  a14985a );
 a14989a <=( A266  and  (not A265) );
 a14992a <=( A269  and  (not A268) );
 a14993a <=( a14992a  and  a14989a );
 a14994a <=( a14993a  and  a14986a );
 a14998a <=( (not A199)  and  (not A166) );
 a14999a <=( A167  and  a14998a );
 a15003a <=( A232  and  (not A202) );
 a15004a <=( (not A200)  and  a15003a );
 a15005a <=( a15004a  and  a14999a );
 a15009a <=( (not A236)  and  A235 );
 a15010a <=( A233  and  a15009a );
 a15013a <=( (not A266)  and  A265 );
 a15016a <=( A269  and  (not A268) );
 a15017a <=( a15016a  and  a15013a );
 a15018a <=( a15017a  and  a15010a );
 a15022a <=( (not A199)  and  (not A166) );
 a15023a <=( A167  and  a15022a );
 a15027a <=( A232  and  (not A202) );
 a15028a <=( (not A200)  and  a15027a );
 a15029a <=( a15028a  and  a15023a );
 a15033a <=( (not A236)  and  A235 );
 a15034a <=( A233  and  a15033a );
 a15037a <=( (not A266)  and  (not A265) );
 a15040a <=( (not A269)  and  A268 );
 a15041a <=( a15040a  and  a15037a );
 a15042a <=( a15041a  and  a15034a );
 a15046a <=( (not A199)  and  (not A166) );
 a15047a <=( A167  and  a15046a );
 a15051a <=( (not A232)  and  (not A202) );
 a15052a <=( (not A200)  and  a15051a );
 a15053a <=( a15052a  and  a15047a );
 a15057a <=( A236  and  (not A235) );
 a15058a <=( A233  and  a15057a );
 a15061a <=( A299  and  A298 );
 a15064a <=( (not A302)  and  A301 );
 a15065a <=( a15064a  and  a15061a );
 a15066a <=( a15065a  and  a15058a );
 a15070a <=( (not A199)  and  (not A166) );
 a15071a <=( A167  and  a15070a );
 a15075a <=( (not A232)  and  (not A202) );
 a15076a <=( (not A200)  and  a15075a );
 a15077a <=( a15076a  and  a15071a );
 a15081a <=( A236  and  (not A235) );
 a15082a <=( A233  and  a15081a );
 a15085a <=( (not A299)  and  A298 );
 a15088a <=( A302  and  (not A301) );
 a15089a <=( a15088a  and  a15085a );
 a15090a <=( a15089a  and  a15082a );
 a15094a <=( (not A199)  and  (not A166) );
 a15095a <=( A167  and  a15094a );
 a15099a <=( (not A232)  and  (not A202) );
 a15100a <=( (not A200)  and  a15099a );
 a15101a <=( a15100a  and  a15095a );
 a15105a <=( A236  and  (not A235) );
 a15106a <=( A233  and  a15105a );
 a15109a <=( A299  and  (not A298) );
 a15112a <=( A302  and  (not A301) );
 a15113a <=( a15112a  and  a15109a );
 a15114a <=( a15113a  and  a15106a );
 a15118a <=( (not A199)  and  (not A166) );
 a15119a <=( A167  and  a15118a );
 a15123a <=( (not A232)  and  (not A202) );
 a15124a <=( (not A200)  and  a15123a );
 a15125a <=( a15124a  and  a15119a );
 a15129a <=( A236  and  (not A235) );
 a15130a <=( A233  and  a15129a );
 a15133a <=( (not A299)  and  (not A298) );
 a15136a <=( (not A302)  and  A301 );
 a15137a <=( a15136a  and  a15133a );
 a15138a <=( a15137a  and  a15130a );
 a15142a <=( (not A199)  and  (not A166) );
 a15143a <=( A167  and  a15142a );
 a15147a <=( (not A232)  and  (not A202) );
 a15148a <=( (not A200)  and  a15147a );
 a15149a <=( a15148a  and  a15143a );
 a15153a <=( A236  and  (not A235) );
 a15154a <=( A233  and  a15153a );
 a15157a <=( A266  and  A265 );
 a15160a <=( (not A269)  and  A268 );
 a15161a <=( a15160a  and  a15157a );
 a15162a <=( a15161a  and  a15154a );
 a15166a <=( (not A199)  and  (not A166) );
 a15167a <=( A167  and  a15166a );
 a15171a <=( (not A232)  and  (not A202) );
 a15172a <=( (not A200)  and  a15171a );
 a15173a <=( a15172a  and  a15167a );
 a15177a <=( A236  and  (not A235) );
 a15178a <=( A233  and  a15177a );
 a15181a <=( A266  and  (not A265) );
 a15184a <=( A269  and  (not A268) );
 a15185a <=( a15184a  and  a15181a );
 a15186a <=( a15185a  and  a15178a );
 a15190a <=( (not A199)  and  (not A166) );
 a15191a <=( A167  and  a15190a );
 a15195a <=( (not A232)  and  (not A202) );
 a15196a <=( (not A200)  and  a15195a );
 a15197a <=( a15196a  and  a15191a );
 a15201a <=( A236  and  (not A235) );
 a15202a <=( A233  and  a15201a );
 a15205a <=( (not A266)  and  A265 );
 a15208a <=( A269  and  (not A268) );
 a15209a <=( a15208a  and  a15205a );
 a15210a <=( a15209a  and  a15202a );
 a15214a <=( (not A199)  and  (not A166) );
 a15215a <=( A167  and  a15214a );
 a15219a <=( (not A232)  and  (not A202) );
 a15220a <=( (not A200)  and  a15219a );
 a15221a <=( a15220a  and  a15215a );
 a15225a <=( A236  and  (not A235) );
 a15226a <=( A233  and  a15225a );
 a15229a <=( (not A266)  and  (not A265) );
 a15232a <=( (not A269)  and  A268 );
 a15233a <=( a15232a  and  a15229a );
 a15234a <=( a15233a  and  a15226a );
 a15238a <=( (not A199)  and  (not A166) );
 a15239a <=( A167  and  a15238a );
 a15243a <=( A232  and  (not A202) );
 a15244a <=( (not A200)  and  a15243a );
 a15245a <=( a15244a  and  a15239a );
 a15249a <=( A236  and  (not A235) );
 a15250a <=( (not A233)  and  a15249a );
 a15253a <=( A299  and  A298 );
 a15256a <=( (not A302)  and  A301 );
 a15257a <=( a15256a  and  a15253a );
 a15258a <=( a15257a  and  a15250a );
 a15262a <=( (not A199)  and  (not A166) );
 a15263a <=( A167  and  a15262a );
 a15267a <=( A232  and  (not A202) );
 a15268a <=( (not A200)  and  a15267a );
 a15269a <=( a15268a  and  a15263a );
 a15273a <=( A236  and  (not A235) );
 a15274a <=( (not A233)  and  a15273a );
 a15277a <=( (not A299)  and  A298 );
 a15280a <=( A302  and  (not A301) );
 a15281a <=( a15280a  and  a15277a );
 a15282a <=( a15281a  and  a15274a );
 a15286a <=( (not A199)  and  (not A166) );
 a15287a <=( A167  and  a15286a );
 a15291a <=( A232  and  (not A202) );
 a15292a <=( (not A200)  and  a15291a );
 a15293a <=( a15292a  and  a15287a );
 a15297a <=( A236  and  (not A235) );
 a15298a <=( (not A233)  and  a15297a );
 a15301a <=( A299  and  (not A298) );
 a15304a <=( A302  and  (not A301) );
 a15305a <=( a15304a  and  a15301a );
 a15306a <=( a15305a  and  a15298a );
 a15310a <=( (not A199)  and  (not A166) );
 a15311a <=( A167  and  a15310a );
 a15315a <=( A232  and  (not A202) );
 a15316a <=( (not A200)  and  a15315a );
 a15317a <=( a15316a  and  a15311a );
 a15321a <=( A236  and  (not A235) );
 a15322a <=( (not A233)  and  a15321a );
 a15325a <=( (not A299)  and  (not A298) );
 a15328a <=( (not A302)  and  A301 );
 a15329a <=( a15328a  and  a15325a );
 a15330a <=( a15329a  and  a15322a );
 a15334a <=( (not A199)  and  (not A166) );
 a15335a <=( A167  and  a15334a );
 a15339a <=( A232  and  (not A202) );
 a15340a <=( (not A200)  and  a15339a );
 a15341a <=( a15340a  and  a15335a );
 a15345a <=( A236  and  (not A235) );
 a15346a <=( (not A233)  and  a15345a );
 a15349a <=( A266  and  A265 );
 a15352a <=( (not A269)  and  A268 );
 a15353a <=( a15352a  and  a15349a );
 a15354a <=( a15353a  and  a15346a );
 a15358a <=( (not A199)  and  (not A166) );
 a15359a <=( A167  and  a15358a );
 a15363a <=( A232  and  (not A202) );
 a15364a <=( (not A200)  and  a15363a );
 a15365a <=( a15364a  and  a15359a );
 a15369a <=( A236  and  (not A235) );
 a15370a <=( (not A233)  and  a15369a );
 a15373a <=( A266  and  (not A265) );
 a15376a <=( A269  and  (not A268) );
 a15377a <=( a15376a  and  a15373a );
 a15378a <=( a15377a  and  a15370a );
 a15382a <=( (not A199)  and  (not A166) );
 a15383a <=( A167  and  a15382a );
 a15387a <=( A232  and  (not A202) );
 a15388a <=( (not A200)  and  a15387a );
 a15389a <=( a15388a  and  a15383a );
 a15393a <=( A236  and  (not A235) );
 a15394a <=( (not A233)  and  a15393a );
 a15397a <=( (not A266)  and  A265 );
 a15400a <=( A269  and  (not A268) );
 a15401a <=( a15400a  and  a15397a );
 a15402a <=( a15401a  and  a15394a );
 a15406a <=( (not A199)  and  (not A166) );
 a15407a <=( A167  and  a15406a );
 a15411a <=( A232  and  (not A202) );
 a15412a <=( (not A200)  and  a15411a );
 a15413a <=( a15412a  and  a15407a );
 a15417a <=( A236  and  (not A235) );
 a15418a <=( (not A233)  and  a15417a );
 a15421a <=( (not A266)  and  (not A265) );
 a15424a <=( (not A269)  and  A268 );
 a15425a <=( a15424a  and  a15421a );
 a15426a <=( a15425a  and  a15418a );
 a15430a <=( (not A199)  and  (not A166) );
 a15431a <=( A167  and  a15430a );
 a15435a <=( (not A232)  and  (not A202) );
 a15436a <=( (not A200)  and  a15435a );
 a15437a <=( a15436a  and  a15431a );
 a15441a <=( (not A236)  and  A235 );
 a15442a <=( (not A233)  and  a15441a );
 a15445a <=( A299  and  A298 );
 a15448a <=( (not A302)  and  A301 );
 a15449a <=( a15448a  and  a15445a );
 a15450a <=( a15449a  and  a15442a );
 a15454a <=( (not A199)  and  (not A166) );
 a15455a <=( A167  and  a15454a );
 a15459a <=( (not A232)  and  (not A202) );
 a15460a <=( (not A200)  and  a15459a );
 a15461a <=( a15460a  and  a15455a );
 a15465a <=( (not A236)  and  A235 );
 a15466a <=( (not A233)  and  a15465a );
 a15469a <=( (not A299)  and  A298 );
 a15472a <=( A302  and  (not A301) );
 a15473a <=( a15472a  and  a15469a );
 a15474a <=( a15473a  and  a15466a );
 a15478a <=( (not A199)  and  (not A166) );
 a15479a <=( A167  and  a15478a );
 a15483a <=( (not A232)  and  (not A202) );
 a15484a <=( (not A200)  and  a15483a );
 a15485a <=( a15484a  and  a15479a );
 a15489a <=( (not A236)  and  A235 );
 a15490a <=( (not A233)  and  a15489a );
 a15493a <=( A299  and  (not A298) );
 a15496a <=( A302  and  (not A301) );
 a15497a <=( a15496a  and  a15493a );
 a15498a <=( a15497a  and  a15490a );
 a15502a <=( (not A199)  and  (not A166) );
 a15503a <=( A167  and  a15502a );
 a15507a <=( (not A232)  and  (not A202) );
 a15508a <=( (not A200)  and  a15507a );
 a15509a <=( a15508a  and  a15503a );
 a15513a <=( (not A236)  and  A235 );
 a15514a <=( (not A233)  and  a15513a );
 a15517a <=( (not A299)  and  (not A298) );
 a15520a <=( (not A302)  and  A301 );
 a15521a <=( a15520a  and  a15517a );
 a15522a <=( a15521a  and  a15514a );
 a15526a <=( (not A199)  and  (not A166) );
 a15527a <=( A167  and  a15526a );
 a15531a <=( (not A232)  and  (not A202) );
 a15532a <=( (not A200)  and  a15531a );
 a15533a <=( a15532a  and  a15527a );
 a15537a <=( (not A236)  and  A235 );
 a15538a <=( (not A233)  and  a15537a );
 a15541a <=( A266  and  A265 );
 a15544a <=( (not A269)  and  A268 );
 a15545a <=( a15544a  and  a15541a );
 a15546a <=( a15545a  and  a15538a );
 a15550a <=( (not A199)  and  (not A166) );
 a15551a <=( A167  and  a15550a );
 a15555a <=( (not A232)  and  (not A202) );
 a15556a <=( (not A200)  and  a15555a );
 a15557a <=( a15556a  and  a15551a );
 a15561a <=( (not A236)  and  A235 );
 a15562a <=( (not A233)  and  a15561a );
 a15565a <=( A266  and  (not A265) );
 a15568a <=( A269  and  (not A268) );
 a15569a <=( a15568a  and  a15565a );
 a15570a <=( a15569a  and  a15562a );
 a15574a <=( (not A199)  and  (not A166) );
 a15575a <=( A167  and  a15574a );
 a15579a <=( (not A232)  and  (not A202) );
 a15580a <=( (not A200)  and  a15579a );
 a15581a <=( a15580a  and  a15575a );
 a15585a <=( (not A236)  and  A235 );
 a15586a <=( (not A233)  and  a15585a );
 a15589a <=( (not A266)  and  A265 );
 a15592a <=( A269  and  (not A268) );
 a15593a <=( a15592a  and  a15589a );
 a15594a <=( a15593a  and  a15586a );
 a15598a <=( (not A199)  and  (not A166) );
 a15599a <=( A167  and  a15598a );
 a15603a <=( (not A232)  and  (not A202) );
 a15604a <=( (not A200)  and  a15603a );
 a15605a <=( a15604a  and  a15599a );
 a15609a <=( (not A236)  and  A235 );
 a15610a <=( (not A233)  and  a15609a );
 a15613a <=( (not A266)  and  (not A265) );
 a15616a <=( (not A269)  and  A268 );
 a15617a <=( a15616a  and  a15613a );
 a15618a <=( a15617a  and  a15610a );
 a15622a <=( (not A199)  and  (not A166) );
 a15623a <=( A167  and  a15622a );
 a15627a <=( A232  and  A203 );
 a15628a <=( (not A200)  and  a15627a );
 a15629a <=( a15628a  and  a15623a );
 a15633a <=( (not A236)  and  A235 );
 a15634a <=( A233  and  a15633a );
 a15637a <=( A299  and  A298 );
 a15640a <=( (not A302)  and  A301 );
 a15641a <=( a15640a  and  a15637a );
 a15642a <=( a15641a  and  a15634a );
 a15646a <=( (not A199)  and  (not A166) );
 a15647a <=( A167  and  a15646a );
 a15651a <=( A232  and  A203 );
 a15652a <=( (not A200)  and  a15651a );
 a15653a <=( a15652a  and  a15647a );
 a15657a <=( (not A236)  and  A235 );
 a15658a <=( A233  and  a15657a );
 a15661a <=( (not A299)  and  A298 );
 a15664a <=( A302  and  (not A301) );
 a15665a <=( a15664a  and  a15661a );
 a15666a <=( a15665a  and  a15658a );
 a15670a <=( (not A199)  and  (not A166) );
 a15671a <=( A167  and  a15670a );
 a15675a <=( A232  and  A203 );
 a15676a <=( (not A200)  and  a15675a );
 a15677a <=( a15676a  and  a15671a );
 a15681a <=( (not A236)  and  A235 );
 a15682a <=( A233  and  a15681a );
 a15685a <=( A299  and  (not A298) );
 a15688a <=( A302  and  (not A301) );
 a15689a <=( a15688a  and  a15685a );
 a15690a <=( a15689a  and  a15682a );
 a15694a <=( (not A199)  and  (not A166) );
 a15695a <=( A167  and  a15694a );
 a15699a <=( A232  and  A203 );
 a15700a <=( (not A200)  and  a15699a );
 a15701a <=( a15700a  and  a15695a );
 a15705a <=( (not A236)  and  A235 );
 a15706a <=( A233  and  a15705a );
 a15709a <=( (not A299)  and  (not A298) );
 a15712a <=( (not A302)  and  A301 );
 a15713a <=( a15712a  and  a15709a );
 a15714a <=( a15713a  and  a15706a );
 a15718a <=( (not A199)  and  (not A166) );
 a15719a <=( A167  and  a15718a );
 a15723a <=( A232  and  A203 );
 a15724a <=( (not A200)  and  a15723a );
 a15725a <=( a15724a  and  a15719a );
 a15729a <=( (not A236)  and  A235 );
 a15730a <=( A233  and  a15729a );
 a15733a <=( A266  and  A265 );
 a15736a <=( (not A269)  and  A268 );
 a15737a <=( a15736a  and  a15733a );
 a15738a <=( a15737a  and  a15730a );
 a15742a <=( (not A199)  and  (not A166) );
 a15743a <=( A167  and  a15742a );
 a15747a <=( A232  and  A203 );
 a15748a <=( (not A200)  and  a15747a );
 a15749a <=( a15748a  and  a15743a );
 a15753a <=( (not A236)  and  A235 );
 a15754a <=( A233  and  a15753a );
 a15757a <=( A266  and  (not A265) );
 a15760a <=( A269  and  (not A268) );
 a15761a <=( a15760a  and  a15757a );
 a15762a <=( a15761a  and  a15754a );
 a15766a <=( (not A199)  and  (not A166) );
 a15767a <=( A167  and  a15766a );
 a15771a <=( A232  and  A203 );
 a15772a <=( (not A200)  and  a15771a );
 a15773a <=( a15772a  and  a15767a );
 a15777a <=( (not A236)  and  A235 );
 a15778a <=( A233  and  a15777a );
 a15781a <=( (not A266)  and  A265 );
 a15784a <=( A269  and  (not A268) );
 a15785a <=( a15784a  and  a15781a );
 a15786a <=( a15785a  and  a15778a );
 a15790a <=( (not A199)  and  (not A166) );
 a15791a <=( A167  and  a15790a );
 a15795a <=( A232  and  A203 );
 a15796a <=( (not A200)  and  a15795a );
 a15797a <=( a15796a  and  a15791a );
 a15801a <=( (not A236)  and  A235 );
 a15802a <=( A233  and  a15801a );
 a15805a <=( (not A266)  and  (not A265) );
 a15808a <=( (not A269)  and  A268 );
 a15809a <=( a15808a  and  a15805a );
 a15810a <=( a15809a  and  a15802a );
 a15814a <=( (not A199)  and  (not A166) );
 a15815a <=( A167  and  a15814a );
 a15819a <=( (not A232)  and  A203 );
 a15820a <=( (not A200)  and  a15819a );
 a15821a <=( a15820a  and  a15815a );
 a15825a <=( A236  and  (not A235) );
 a15826a <=( A233  and  a15825a );
 a15829a <=( A299  and  A298 );
 a15832a <=( (not A302)  and  A301 );
 a15833a <=( a15832a  and  a15829a );
 a15834a <=( a15833a  and  a15826a );
 a15838a <=( (not A199)  and  (not A166) );
 a15839a <=( A167  and  a15838a );
 a15843a <=( (not A232)  and  A203 );
 a15844a <=( (not A200)  and  a15843a );
 a15845a <=( a15844a  and  a15839a );
 a15849a <=( A236  and  (not A235) );
 a15850a <=( A233  and  a15849a );
 a15853a <=( (not A299)  and  A298 );
 a15856a <=( A302  and  (not A301) );
 a15857a <=( a15856a  and  a15853a );
 a15858a <=( a15857a  and  a15850a );
 a15862a <=( (not A199)  and  (not A166) );
 a15863a <=( A167  and  a15862a );
 a15867a <=( (not A232)  and  A203 );
 a15868a <=( (not A200)  and  a15867a );
 a15869a <=( a15868a  and  a15863a );
 a15873a <=( A236  and  (not A235) );
 a15874a <=( A233  and  a15873a );
 a15877a <=( A299  and  (not A298) );
 a15880a <=( A302  and  (not A301) );
 a15881a <=( a15880a  and  a15877a );
 a15882a <=( a15881a  and  a15874a );
 a15886a <=( (not A199)  and  (not A166) );
 a15887a <=( A167  and  a15886a );
 a15891a <=( (not A232)  and  A203 );
 a15892a <=( (not A200)  and  a15891a );
 a15893a <=( a15892a  and  a15887a );
 a15897a <=( A236  and  (not A235) );
 a15898a <=( A233  and  a15897a );
 a15901a <=( (not A299)  and  (not A298) );
 a15904a <=( (not A302)  and  A301 );
 a15905a <=( a15904a  and  a15901a );
 a15906a <=( a15905a  and  a15898a );
 a15910a <=( (not A199)  and  (not A166) );
 a15911a <=( A167  and  a15910a );
 a15915a <=( (not A232)  and  A203 );
 a15916a <=( (not A200)  and  a15915a );
 a15917a <=( a15916a  and  a15911a );
 a15921a <=( A236  and  (not A235) );
 a15922a <=( A233  and  a15921a );
 a15925a <=( A266  and  A265 );
 a15928a <=( (not A269)  and  A268 );
 a15929a <=( a15928a  and  a15925a );
 a15930a <=( a15929a  and  a15922a );
 a15934a <=( (not A199)  and  (not A166) );
 a15935a <=( A167  and  a15934a );
 a15939a <=( (not A232)  and  A203 );
 a15940a <=( (not A200)  and  a15939a );
 a15941a <=( a15940a  and  a15935a );
 a15945a <=( A236  and  (not A235) );
 a15946a <=( A233  and  a15945a );
 a15949a <=( A266  and  (not A265) );
 a15952a <=( A269  and  (not A268) );
 a15953a <=( a15952a  and  a15949a );
 a15954a <=( a15953a  and  a15946a );
 a15958a <=( (not A199)  and  (not A166) );
 a15959a <=( A167  and  a15958a );
 a15963a <=( (not A232)  and  A203 );
 a15964a <=( (not A200)  and  a15963a );
 a15965a <=( a15964a  and  a15959a );
 a15969a <=( A236  and  (not A235) );
 a15970a <=( A233  and  a15969a );
 a15973a <=( (not A266)  and  A265 );
 a15976a <=( A269  and  (not A268) );
 a15977a <=( a15976a  and  a15973a );
 a15978a <=( a15977a  and  a15970a );
 a15982a <=( (not A199)  and  (not A166) );
 a15983a <=( A167  and  a15982a );
 a15987a <=( (not A232)  and  A203 );
 a15988a <=( (not A200)  and  a15987a );
 a15989a <=( a15988a  and  a15983a );
 a15993a <=( A236  and  (not A235) );
 a15994a <=( A233  and  a15993a );
 a15997a <=( (not A266)  and  (not A265) );
 a16000a <=( (not A269)  and  A268 );
 a16001a <=( a16000a  and  a15997a );
 a16002a <=( a16001a  and  a15994a );
 a16006a <=( (not A199)  and  (not A166) );
 a16007a <=( A167  and  a16006a );
 a16011a <=( A232  and  A203 );
 a16012a <=( (not A200)  and  a16011a );
 a16013a <=( a16012a  and  a16007a );
 a16017a <=( A236  and  (not A235) );
 a16018a <=( (not A233)  and  a16017a );
 a16021a <=( A299  and  A298 );
 a16024a <=( (not A302)  and  A301 );
 a16025a <=( a16024a  and  a16021a );
 a16026a <=( a16025a  and  a16018a );
 a16030a <=( (not A199)  and  (not A166) );
 a16031a <=( A167  and  a16030a );
 a16035a <=( A232  and  A203 );
 a16036a <=( (not A200)  and  a16035a );
 a16037a <=( a16036a  and  a16031a );
 a16041a <=( A236  and  (not A235) );
 a16042a <=( (not A233)  and  a16041a );
 a16045a <=( (not A299)  and  A298 );
 a16048a <=( A302  and  (not A301) );
 a16049a <=( a16048a  and  a16045a );
 a16050a <=( a16049a  and  a16042a );
 a16054a <=( (not A199)  and  (not A166) );
 a16055a <=( A167  and  a16054a );
 a16059a <=( A232  and  A203 );
 a16060a <=( (not A200)  and  a16059a );
 a16061a <=( a16060a  and  a16055a );
 a16065a <=( A236  and  (not A235) );
 a16066a <=( (not A233)  and  a16065a );
 a16069a <=( A299  and  (not A298) );
 a16072a <=( A302  and  (not A301) );
 a16073a <=( a16072a  and  a16069a );
 a16074a <=( a16073a  and  a16066a );
 a16078a <=( (not A199)  and  (not A166) );
 a16079a <=( A167  and  a16078a );
 a16083a <=( A232  and  A203 );
 a16084a <=( (not A200)  and  a16083a );
 a16085a <=( a16084a  and  a16079a );
 a16089a <=( A236  and  (not A235) );
 a16090a <=( (not A233)  and  a16089a );
 a16093a <=( (not A299)  and  (not A298) );
 a16096a <=( (not A302)  and  A301 );
 a16097a <=( a16096a  and  a16093a );
 a16098a <=( a16097a  and  a16090a );
 a16102a <=( (not A199)  and  (not A166) );
 a16103a <=( A167  and  a16102a );
 a16107a <=( A232  and  A203 );
 a16108a <=( (not A200)  and  a16107a );
 a16109a <=( a16108a  and  a16103a );
 a16113a <=( A236  and  (not A235) );
 a16114a <=( (not A233)  and  a16113a );
 a16117a <=( A266  and  A265 );
 a16120a <=( (not A269)  and  A268 );
 a16121a <=( a16120a  and  a16117a );
 a16122a <=( a16121a  and  a16114a );
 a16126a <=( (not A199)  and  (not A166) );
 a16127a <=( A167  and  a16126a );
 a16131a <=( A232  and  A203 );
 a16132a <=( (not A200)  and  a16131a );
 a16133a <=( a16132a  and  a16127a );
 a16137a <=( A236  and  (not A235) );
 a16138a <=( (not A233)  and  a16137a );
 a16141a <=( A266  and  (not A265) );
 a16144a <=( A269  and  (not A268) );
 a16145a <=( a16144a  and  a16141a );
 a16146a <=( a16145a  and  a16138a );
 a16150a <=( (not A199)  and  (not A166) );
 a16151a <=( A167  and  a16150a );
 a16155a <=( A232  and  A203 );
 a16156a <=( (not A200)  and  a16155a );
 a16157a <=( a16156a  and  a16151a );
 a16161a <=( A236  and  (not A235) );
 a16162a <=( (not A233)  and  a16161a );
 a16165a <=( (not A266)  and  A265 );
 a16168a <=( A269  and  (not A268) );
 a16169a <=( a16168a  and  a16165a );
 a16170a <=( a16169a  and  a16162a );
 a16174a <=( (not A199)  and  (not A166) );
 a16175a <=( A167  and  a16174a );
 a16179a <=( A232  and  A203 );
 a16180a <=( (not A200)  and  a16179a );
 a16181a <=( a16180a  and  a16175a );
 a16185a <=( A236  and  (not A235) );
 a16186a <=( (not A233)  and  a16185a );
 a16189a <=( (not A266)  and  (not A265) );
 a16192a <=( (not A269)  and  A268 );
 a16193a <=( a16192a  and  a16189a );
 a16194a <=( a16193a  and  a16186a );
 a16198a <=( (not A199)  and  (not A166) );
 a16199a <=( A167  and  a16198a );
 a16203a <=( (not A232)  and  A203 );
 a16204a <=( (not A200)  and  a16203a );
 a16205a <=( a16204a  and  a16199a );
 a16209a <=( (not A236)  and  A235 );
 a16210a <=( (not A233)  and  a16209a );
 a16213a <=( A299  and  A298 );
 a16216a <=( (not A302)  and  A301 );
 a16217a <=( a16216a  and  a16213a );
 a16218a <=( a16217a  and  a16210a );
 a16222a <=( (not A199)  and  (not A166) );
 a16223a <=( A167  and  a16222a );
 a16227a <=( (not A232)  and  A203 );
 a16228a <=( (not A200)  and  a16227a );
 a16229a <=( a16228a  and  a16223a );
 a16233a <=( (not A236)  and  A235 );
 a16234a <=( (not A233)  and  a16233a );
 a16237a <=( (not A299)  and  A298 );
 a16240a <=( A302  and  (not A301) );
 a16241a <=( a16240a  and  a16237a );
 a16242a <=( a16241a  and  a16234a );
 a16246a <=( (not A199)  and  (not A166) );
 a16247a <=( A167  and  a16246a );
 a16251a <=( (not A232)  and  A203 );
 a16252a <=( (not A200)  and  a16251a );
 a16253a <=( a16252a  and  a16247a );
 a16257a <=( (not A236)  and  A235 );
 a16258a <=( (not A233)  and  a16257a );
 a16261a <=( A299  and  (not A298) );
 a16264a <=( A302  and  (not A301) );
 a16265a <=( a16264a  and  a16261a );
 a16266a <=( a16265a  and  a16258a );
 a16270a <=( (not A199)  and  (not A166) );
 a16271a <=( A167  and  a16270a );
 a16275a <=( (not A232)  and  A203 );
 a16276a <=( (not A200)  and  a16275a );
 a16277a <=( a16276a  and  a16271a );
 a16281a <=( (not A236)  and  A235 );
 a16282a <=( (not A233)  and  a16281a );
 a16285a <=( (not A299)  and  (not A298) );
 a16288a <=( (not A302)  and  A301 );
 a16289a <=( a16288a  and  a16285a );
 a16290a <=( a16289a  and  a16282a );
 a16294a <=( (not A199)  and  (not A166) );
 a16295a <=( A167  and  a16294a );
 a16299a <=( (not A232)  and  A203 );
 a16300a <=( (not A200)  and  a16299a );
 a16301a <=( a16300a  and  a16295a );
 a16305a <=( (not A236)  and  A235 );
 a16306a <=( (not A233)  and  a16305a );
 a16309a <=( A266  and  A265 );
 a16312a <=( (not A269)  and  A268 );
 a16313a <=( a16312a  and  a16309a );
 a16314a <=( a16313a  and  a16306a );
 a16318a <=( (not A199)  and  (not A166) );
 a16319a <=( A167  and  a16318a );
 a16323a <=( (not A232)  and  A203 );
 a16324a <=( (not A200)  and  a16323a );
 a16325a <=( a16324a  and  a16319a );
 a16329a <=( (not A236)  and  A235 );
 a16330a <=( (not A233)  and  a16329a );
 a16333a <=( A266  and  (not A265) );
 a16336a <=( A269  and  (not A268) );
 a16337a <=( a16336a  and  a16333a );
 a16338a <=( a16337a  and  a16330a );
 a16342a <=( (not A199)  and  (not A166) );
 a16343a <=( A167  and  a16342a );
 a16347a <=( (not A232)  and  A203 );
 a16348a <=( (not A200)  and  a16347a );
 a16349a <=( a16348a  and  a16343a );
 a16353a <=( (not A236)  and  A235 );
 a16354a <=( (not A233)  and  a16353a );
 a16357a <=( (not A266)  and  A265 );
 a16360a <=( A269  and  (not A268) );
 a16361a <=( a16360a  and  a16357a );
 a16362a <=( a16361a  and  a16354a );
 a16366a <=( (not A199)  and  (not A166) );
 a16367a <=( A167  and  a16366a );
 a16371a <=( (not A232)  and  A203 );
 a16372a <=( (not A200)  and  a16371a );
 a16373a <=( a16372a  and  a16367a );
 a16377a <=( (not A236)  and  A235 );
 a16378a <=( (not A233)  and  a16377a );
 a16381a <=( (not A266)  and  (not A265) );
 a16384a <=( (not A269)  and  A268 );
 a16385a <=( a16384a  and  a16381a );
 a16386a <=( a16385a  and  a16378a );
 a16390a <=( (not A167)  and  A168 );
 a16391a <=( A170  and  a16390a );
 a16395a <=( (not A200)  and  (not A199) );
 a16396a <=( A166  and  a16395a );
 a16397a <=( a16396a  and  a16391a );
 a16401a <=( A234  and  A232 );
 a16402a <=( (not A202)  and  a16401a );
 a16405a <=( A299  and  A298 );
 a16408a <=( (not A302)  and  A301 );
 a16409a <=( a16408a  and  a16405a );
 a16410a <=( a16409a  and  a16402a );
 a16414a <=( (not A167)  and  A168 );
 a16415a <=( A170  and  a16414a );
 a16419a <=( (not A200)  and  (not A199) );
 a16420a <=( A166  and  a16419a );
 a16421a <=( a16420a  and  a16415a );
 a16425a <=( A234  and  A232 );
 a16426a <=( (not A202)  and  a16425a );
 a16429a <=( (not A299)  and  A298 );
 a16432a <=( A302  and  (not A301) );
 a16433a <=( a16432a  and  a16429a );
 a16434a <=( a16433a  and  a16426a );
 a16438a <=( (not A167)  and  A168 );
 a16439a <=( A170  and  a16438a );
 a16443a <=( (not A200)  and  (not A199) );
 a16444a <=( A166  and  a16443a );
 a16445a <=( a16444a  and  a16439a );
 a16449a <=( A234  and  A232 );
 a16450a <=( (not A202)  and  a16449a );
 a16453a <=( A299  and  (not A298) );
 a16456a <=( A302  and  (not A301) );
 a16457a <=( a16456a  and  a16453a );
 a16458a <=( a16457a  and  a16450a );
 a16462a <=( (not A167)  and  A168 );
 a16463a <=( A170  and  a16462a );
 a16467a <=( (not A200)  and  (not A199) );
 a16468a <=( A166  and  a16467a );
 a16469a <=( a16468a  and  a16463a );
 a16473a <=( A234  and  A232 );
 a16474a <=( (not A202)  and  a16473a );
 a16477a <=( (not A299)  and  (not A298) );
 a16480a <=( (not A302)  and  A301 );
 a16481a <=( a16480a  and  a16477a );
 a16482a <=( a16481a  and  a16474a );
 a16486a <=( (not A167)  and  A168 );
 a16487a <=( A170  and  a16486a );
 a16491a <=( (not A200)  and  (not A199) );
 a16492a <=( A166  and  a16491a );
 a16493a <=( a16492a  and  a16487a );
 a16497a <=( A234  and  A232 );
 a16498a <=( (not A202)  and  a16497a );
 a16501a <=( A266  and  A265 );
 a16504a <=( (not A269)  and  A268 );
 a16505a <=( a16504a  and  a16501a );
 a16506a <=( a16505a  and  a16498a );
 a16510a <=( (not A167)  and  A168 );
 a16511a <=( A170  and  a16510a );
 a16515a <=( (not A200)  and  (not A199) );
 a16516a <=( A166  and  a16515a );
 a16517a <=( a16516a  and  a16511a );
 a16521a <=( A234  and  A232 );
 a16522a <=( (not A202)  and  a16521a );
 a16525a <=( A266  and  (not A265) );
 a16528a <=( A269  and  (not A268) );
 a16529a <=( a16528a  and  a16525a );
 a16530a <=( a16529a  and  a16522a );
 a16534a <=( (not A167)  and  A168 );
 a16535a <=( A170  and  a16534a );
 a16539a <=( (not A200)  and  (not A199) );
 a16540a <=( A166  and  a16539a );
 a16541a <=( a16540a  and  a16535a );
 a16545a <=( A234  and  A232 );
 a16546a <=( (not A202)  and  a16545a );
 a16549a <=( (not A266)  and  A265 );
 a16552a <=( A269  and  (not A268) );
 a16553a <=( a16552a  and  a16549a );
 a16554a <=( a16553a  and  a16546a );
 a16558a <=( (not A167)  and  A168 );
 a16559a <=( A170  and  a16558a );
 a16563a <=( (not A200)  and  (not A199) );
 a16564a <=( A166  and  a16563a );
 a16565a <=( a16564a  and  a16559a );
 a16569a <=( A234  and  A232 );
 a16570a <=( (not A202)  and  a16569a );
 a16573a <=( (not A266)  and  (not A265) );
 a16576a <=( (not A269)  and  A268 );
 a16577a <=( a16576a  and  a16573a );
 a16578a <=( a16577a  and  a16570a );
 a16582a <=( (not A167)  and  A168 );
 a16583a <=( A170  and  a16582a );
 a16587a <=( (not A200)  and  (not A199) );
 a16588a <=( A166  and  a16587a );
 a16589a <=( a16588a  and  a16583a );
 a16593a <=( A234  and  A233 );
 a16594a <=( (not A202)  and  a16593a );
 a16597a <=( A299  and  A298 );
 a16600a <=( (not A302)  and  A301 );
 a16601a <=( a16600a  and  a16597a );
 a16602a <=( a16601a  and  a16594a );
 a16606a <=( (not A167)  and  A168 );
 a16607a <=( A170  and  a16606a );
 a16611a <=( (not A200)  and  (not A199) );
 a16612a <=( A166  and  a16611a );
 a16613a <=( a16612a  and  a16607a );
 a16617a <=( A234  and  A233 );
 a16618a <=( (not A202)  and  a16617a );
 a16621a <=( (not A299)  and  A298 );
 a16624a <=( A302  and  (not A301) );
 a16625a <=( a16624a  and  a16621a );
 a16626a <=( a16625a  and  a16618a );
 a16630a <=( (not A167)  and  A168 );
 a16631a <=( A170  and  a16630a );
 a16635a <=( (not A200)  and  (not A199) );
 a16636a <=( A166  and  a16635a );
 a16637a <=( a16636a  and  a16631a );
 a16641a <=( A234  and  A233 );
 a16642a <=( (not A202)  and  a16641a );
 a16645a <=( A299  and  (not A298) );
 a16648a <=( A302  and  (not A301) );
 a16649a <=( a16648a  and  a16645a );
 a16650a <=( a16649a  and  a16642a );
 a16654a <=( (not A167)  and  A168 );
 a16655a <=( A170  and  a16654a );
 a16659a <=( (not A200)  and  (not A199) );
 a16660a <=( A166  and  a16659a );
 a16661a <=( a16660a  and  a16655a );
 a16665a <=( A234  and  A233 );
 a16666a <=( (not A202)  and  a16665a );
 a16669a <=( (not A299)  and  (not A298) );
 a16672a <=( (not A302)  and  A301 );
 a16673a <=( a16672a  and  a16669a );
 a16674a <=( a16673a  and  a16666a );
 a16678a <=( (not A167)  and  A168 );
 a16679a <=( A170  and  a16678a );
 a16683a <=( (not A200)  and  (not A199) );
 a16684a <=( A166  and  a16683a );
 a16685a <=( a16684a  and  a16679a );
 a16689a <=( A234  and  A233 );
 a16690a <=( (not A202)  and  a16689a );
 a16693a <=( A266  and  A265 );
 a16696a <=( (not A269)  and  A268 );
 a16697a <=( a16696a  and  a16693a );
 a16698a <=( a16697a  and  a16690a );
 a16702a <=( (not A167)  and  A168 );
 a16703a <=( A170  and  a16702a );
 a16707a <=( (not A200)  and  (not A199) );
 a16708a <=( A166  and  a16707a );
 a16709a <=( a16708a  and  a16703a );
 a16713a <=( A234  and  A233 );
 a16714a <=( (not A202)  and  a16713a );
 a16717a <=( A266  and  (not A265) );
 a16720a <=( A269  and  (not A268) );
 a16721a <=( a16720a  and  a16717a );
 a16722a <=( a16721a  and  a16714a );
 a16726a <=( (not A167)  and  A168 );
 a16727a <=( A170  and  a16726a );
 a16731a <=( (not A200)  and  (not A199) );
 a16732a <=( A166  and  a16731a );
 a16733a <=( a16732a  and  a16727a );
 a16737a <=( A234  and  A233 );
 a16738a <=( (not A202)  and  a16737a );
 a16741a <=( (not A266)  and  A265 );
 a16744a <=( A269  and  (not A268) );
 a16745a <=( a16744a  and  a16741a );
 a16746a <=( a16745a  and  a16738a );
 a16750a <=( (not A167)  and  A168 );
 a16751a <=( A170  and  a16750a );
 a16755a <=( (not A200)  and  (not A199) );
 a16756a <=( A166  and  a16755a );
 a16757a <=( a16756a  and  a16751a );
 a16761a <=( A234  and  A233 );
 a16762a <=( (not A202)  and  a16761a );
 a16765a <=( (not A266)  and  (not A265) );
 a16768a <=( (not A269)  and  A268 );
 a16769a <=( a16768a  and  a16765a );
 a16770a <=( a16769a  and  a16762a );
 a16774a <=( (not A167)  and  A168 );
 a16775a <=( A170  and  a16774a );
 a16779a <=( (not A200)  and  (not A199) );
 a16780a <=( A166  and  a16779a );
 a16781a <=( a16780a  and  a16775a );
 a16785a <=( A233  and  A232 );
 a16786a <=( (not A202)  and  a16785a );
 a16789a <=( (not A236)  and  A235 );
 a16792a <=( A300  and  A299 );
 a16793a <=( a16792a  and  a16789a );
 a16794a <=( a16793a  and  a16786a );
 a16798a <=( (not A167)  and  A168 );
 a16799a <=( A170  and  a16798a );
 a16803a <=( (not A200)  and  (not A199) );
 a16804a <=( A166  and  a16803a );
 a16805a <=( a16804a  and  a16799a );
 a16809a <=( A233  and  A232 );
 a16810a <=( (not A202)  and  a16809a );
 a16813a <=( (not A236)  and  A235 );
 a16816a <=( A300  and  A298 );
 a16817a <=( a16816a  and  a16813a );
 a16818a <=( a16817a  and  a16810a );
 a16822a <=( (not A167)  and  A168 );
 a16823a <=( A170  and  a16822a );
 a16827a <=( (not A200)  and  (not A199) );
 a16828a <=( A166  and  a16827a );
 a16829a <=( a16828a  and  a16823a );
 a16833a <=( A233  and  A232 );
 a16834a <=( (not A202)  and  a16833a );
 a16837a <=( (not A236)  and  A235 );
 a16840a <=( A267  and  A265 );
 a16841a <=( a16840a  and  a16837a );
 a16842a <=( a16841a  and  a16834a );
 a16846a <=( (not A167)  and  A168 );
 a16847a <=( A170  and  a16846a );
 a16851a <=( (not A200)  and  (not A199) );
 a16852a <=( A166  and  a16851a );
 a16853a <=( a16852a  and  a16847a );
 a16857a <=( A233  and  A232 );
 a16858a <=( (not A202)  and  a16857a );
 a16861a <=( (not A236)  and  A235 );
 a16864a <=( A267  and  A266 );
 a16865a <=( a16864a  and  a16861a );
 a16866a <=( a16865a  and  a16858a );
 a16870a <=( (not A167)  and  A168 );
 a16871a <=( A170  and  a16870a );
 a16875a <=( (not A200)  and  (not A199) );
 a16876a <=( A166  and  a16875a );
 a16877a <=( a16876a  and  a16871a );
 a16881a <=( A233  and  (not A232) );
 a16882a <=( (not A202)  and  a16881a );
 a16885a <=( A236  and  (not A235) );
 a16888a <=( A300  and  A299 );
 a16889a <=( a16888a  and  a16885a );
 a16890a <=( a16889a  and  a16882a );
 a16894a <=( (not A167)  and  A168 );
 a16895a <=( A170  and  a16894a );
 a16899a <=( (not A200)  and  (not A199) );
 a16900a <=( A166  and  a16899a );
 a16901a <=( a16900a  and  a16895a );
 a16905a <=( A233  and  (not A232) );
 a16906a <=( (not A202)  and  a16905a );
 a16909a <=( A236  and  (not A235) );
 a16912a <=( A300  and  A298 );
 a16913a <=( a16912a  and  a16909a );
 a16914a <=( a16913a  and  a16906a );
 a16918a <=( (not A167)  and  A168 );
 a16919a <=( A170  and  a16918a );
 a16923a <=( (not A200)  and  (not A199) );
 a16924a <=( A166  and  a16923a );
 a16925a <=( a16924a  and  a16919a );
 a16929a <=( A233  and  (not A232) );
 a16930a <=( (not A202)  and  a16929a );
 a16933a <=( A236  and  (not A235) );
 a16936a <=( A267  and  A265 );
 a16937a <=( a16936a  and  a16933a );
 a16938a <=( a16937a  and  a16930a );
 a16942a <=( (not A167)  and  A168 );
 a16943a <=( A170  and  a16942a );
 a16947a <=( (not A200)  and  (not A199) );
 a16948a <=( A166  and  a16947a );
 a16949a <=( a16948a  and  a16943a );
 a16953a <=( A233  and  (not A232) );
 a16954a <=( (not A202)  and  a16953a );
 a16957a <=( A236  and  (not A235) );
 a16960a <=( A267  and  A266 );
 a16961a <=( a16960a  and  a16957a );
 a16962a <=( a16961a  and  a16954a );
 a16966a <=( (not A167)  and  A168 );
 a16967a <=( A170  and  a16966a );
 a16971a <=( (not A200)  and  (not A199) );
 a16972a <=( A166  and  a16971a );
 a16973a <=( a16972a  and  a16967a );
 a16977a <=( (not A233)  and  A232 );
 a16978a <=( (not A202)  and  a16977a );
 a16981a <=( A236  and  (not A235) );
 a16984a <=( A300  and  A299 );
 a16985a <=( a16984a  and  a16981a );
 a16986a <=( a16985a  and  a16978a );
 a16990a <=( (not A167)  and  A168 );
 a16991a <=( A170  and  a16990a );
 a16995a <=( (not A200)  and  (not A199) );
 a16996a <=( A166  and  a16995a );
 a16997a <=( a16996a  and  a16991a );
 a17001a <=( (not A233)  and  A232 );
 a17002a <=( (not A202)  and  a17001a );
 a17005a <=( A236  and  (not A235) );
 a17008a <=( A300  and  A298 );
 a17009a <=( a17008a  and  a17005a );
 a17010a <=( a17009a  and  a17002a );
 a17014a <=( (not A167)  and  A168 );
 a17015a <=( A170  and  a17014a );
 a17019a <=( (not A200)  and  (not A199) );
 a17020a <=( A166  and  a17019a );
 a17021a <=( a17020a  and  a17015a );
 a17025a <=( (not A233)  and  A232 );
 a17026a <=( (not A202)  and  a17025a );
 a17029a <=( A236  and  (not A235) );
 a17032a <=( A267  and  A265 );
 a17033a <=( a17032a  and  a17029a );
 a17034a <=( a17033a  and  a17026a );
 a17038a <=( (not A167)  and  A168 );
 a17039a <=( A170  and  a17038a );
 a17043a <=( (not A200)  and  (not A199) );
 a17044a <=( A166  and  a17043a );
 a17045a <=( a17044a  and  a17039a );
 a17049a <=( (not A233)  and  A232 );
 a17050a <=( (not A202)  and  a17049a );
 a17053a <=( A236  and  (not A235) );
 a17056a <=( A267  and  A266 );
 a17057a <=( a17056a  and  a17053a );
 a17058a <=( a17057a  and  a17050a );
 a17062a <=( (not A167)  and  A168 );
 a17063a <=( A170  and  a17062a );
 a17067a <=( (not A200)  and  (not A199) );
 a17068a <=( A166  and  a17067a );
 a17069a <=( a17068a  and  a17063a );
 a17073a <=( (not A233)  and  (not A232) );
 a17074a <=( (not A202)  and  a17073a );
 a17077a <=( (not A236)  and  A235 );
 a17080a <=( A300  and  A299 );
 a17081a <=( a17080a  and  a17077a );
 a17082a <=( a17081a  and  a17074a );
 a17086a <=( (not A167)  and  A168 );
 a17087a <=( A170  and  a17086a );
 a17091a <=( (not A200)  and  (not A199) );
 a17092a <=( A166  and  a17091a );
 a17093a <=( a17092a  and  a17087a );
 a17097a <=( (not A233)  and  (not A232) );
 a17098a <=( (not A202)  and  a17097a );
 a17101a <=( (not A236)  and  A235 );
 a17104a <=( A300  and  A298 );
 a17105a <=( a17104a  and  a17101a );
 a17106a <=( a17105a  and  a17098a );
 a17110a <=( (not A167)  and  A168 );
 a17111a <=( A170  and  a17110a );
 a17115a <=( (not A200)  and  (not A199) );
 a17116a <=( A166  and  a17115a );
 a17117a <=( a17116a  and  a17111a );
 a17121a <=( (not A233)  and  (not A232) );
 a17122a <=( (not A202)  and  a17121a );
 a17125a <=( (not A236)  and  A235 );
 a17128a <=( A267  and  A265 );
 a17129a <=( a17128a  and  a17125a );
 a17130a <=( a17129a  and  a17122a );
 a17134a <=( (not A167)  and  A168 );
 a17135a <=( A170  and  a17134a );
 a17139a <=( (not A200)  and  (not A199) );
 a17140a <=( A166  and  a17139a );
 a17141a <=( a17140a  and  a17135a );
 a17145a <=( (not A233)  and  (not A232) );
 a17146a <=( (not A202)  and  a17145a );
 a17149a <=( (not A236)  and  A235 );
 a17152a <=( A267  and  A266 );
 a17153a <=( a17152a  and  a17149a );
 a17154a <=( a17153a  and  a17146a );
 a17158a <=( (not A167)  and  A168 );
 a17159a <=( A170  and  a17158a );
 a17163a <=( (not A200)  and  (not A199) );
 a17164a <=( A166  and  a17163a );
 a17165a <=( a17164a  and  a17159a );
 a17169a <=( A234  and  A232 );
 a17170a <=( A203  and  a17169a );
 a17173a <=( A299  and  A298 );
 a17176a <=( (not A302)  and  A301 );
 a17177a <=( a17176a  and  a17173a );
 a17178a <=( a17177a  and  a17170a );
 a17182a <=( (not A167)  and  A168 );
 a17183a <=( A170  and  a17182a );
 a17187a <=( (not A200)  and  (not A199) );
 a17188a <=( A166  and  a17187a );
 a17189a <=( a17188a  and  a17183a );
 a17193a <=( A234  and  A232 );
 a17194a <=( A203  and  a17193a );
 a17197a <=( (not A299)  and  A298 );
 a17200a <=( A302  and  (not A301) );
 a17201a <=( a17200a  and  a17197a );
 a17202a <=( a17201a  and  a17194a );
 a17206a <=( (not A167)  and  A168 );
 a17207a <=( A170  and  a17206a );
 a17211a <=( (not A200)  and  (not A199) );
 a17212a <=( A166  and  a17211a );
 a17213a <=( a17212a  and  a17207a );
 a17217a <=( A234  and  A232 );
 a17218a <=( A203  and  a17217a );
 a17221a <=( A299  and  (not A298) );
 a17224a <=( A302  and  (not A301) );
 a17225a <=( a17224a  and  a17221a );
 a17226a <=( a17225a  and  a17218a );
 a17230a <=( (not A167)  and  A168 );
 a17231a <=( A170  and  a17230a );
 a17235a <=( (not A200)  and  (not A199) );
 a17236a <=( A166  and  a17235a );
 a17237a <=( a17236a  and  a17231a );
 a17241a <=( A234  and  A232 );
 a17242a <=( A203  and  a17241a );
 a17245a <=( (not A299)  and  (not A298) );
 a17248a <=( (not A302)  and  A301 );
 a17249a <=( a17248a  and  a17245a );
 a17250a <=( a17249a  and  a17242a );
 a17254a <=( (not A167)  and  A168 );
 a17255a <=( A170  and  a17254a );
 a17259a <=( (not A200)  and  (not A199) );
 a17260a <=( A166  and  a17259a );
 a17261a <=( a17260a  and  a17255a );
 a17265a <=( A234  and  A232 );
 a17266a <=( A203  and  a17265a );
 a17269a <=( A266  and  A265 );
 a17272a <=( (not A269)  and  A268 );
 a17273a <=( a17272a  and  a17269a );
 a17274a <=( a17273a  and  a17266a );
 a17278a <=( (not A167)  and  A168 );
 a17279a <=( A170  and  a17278a );
 a17283a <=( (not A200)  and  (not A199) );
 a17284a <=( A166  and  a17283a );
 a17285a <=( a17284a  and  a17279a );
 a17289a <=( A234  and  A232 );
 a17290a <=( A203  and  a17289a );
 a17293a <=( A266  and  (not A265) );
 a17296a <=( A269  and  (not A268) );
 a17297a <=( a17296a  and  a17293a );
 a17298a <=( a17297a  and  a17290a );
 a17302a <=( (not A167)  and  A168 );
 a17303a <=( A170  and  a17302a );
 a17307a <=( (not A200)  and  (not A199) );
 a17308a <=( A166  and  a17307a );
 a17309a <=( a17308a  and  a17303a );
 a17313a <=( A234  and  A232 );
 a17314a <=( A203  and  a17313a );
 a17317a <=( (not A266)  and  A265 );
 a17320a <=( A269  and  (not A268) );
 a17321a <=( a17320a  and  a17317a );
 a17322a <=( a17321a  and  a17314a );
 a17326a <=( (not A167)  and  A168 );
 a17327a <=( A170  and  a17326a );
 a17331a <=( (not A200)  and  (not A199) );
 a17332a <=( A166  and  a17331a );
 a17333a <=( a17332a  and  a17327a );
 a17337a <=( A234  and  A232 );
 a17338a <=( A203  and  a17337a );
 a17341a <=( (not A266)  and  (not A265) );
 a17344a <=( (not A269)  and  A268 );
 a17345a <=( a17344a  and  a17341a );
 a17346a <=( a17345a  and  a17338a );
 a17350a <=( (not A167)  and  A168 );
 a17351a <=( A170  and  a17350a );
 a17355a <=( (not A200)  and  (not A199) );
 a17356a <=( A166  and  a17355a );
 a17357a <=( a17356a  and  a17351a );
 a17361a <=( A234  and  A233 );
 a17362a <=( A203  and  a17361a );
 a17365a <=( A299  and  A298 );
 a17368a <=( (not A302)  and  A301 );
 a17369a <=( a17368a  and  a17365a );
 a17370a <=( a17369a  and  a17362a );
 a17374a <=( (not A167)  and  A168 );
 a17375a <=( A170  and  a17374a );
 a17379a <=( (not A200)  and  (not A199) );
 a17380a <=( A166  and  a17379a );
 a17381a <=( a17380a  and  a17375a );
 a17385a <=( A234  and  A233 );
 a17386a <=( A203  and  a17385a );
 a17389a <=( (not A299)  and  A298 );
 a17392a <=( A302  and  (not A301) );
 a17393a <=( a17392a  and  a17389a );
 a17394a <=( a17393a  and  a17386a );
 a17398a <=( (not A167)  and  A168 );
 a17399a <=( A170  and  a17398a );
 a17403a <=( (not A200)  and  (not A199) );
 a17404a <=( A166  and  a17403a );
 a17405a <=( a17404a  and  a17399a );
 a17409a <=( A234  and  A233 );
 a17410a <=( A203  and  a17409a );
 a17413a <=( A299  and  (not A298) );
 a17416a <=( A302  and  (not A301) );
 a17417a <=( a17416a  and  a17413a );
 a17418a <=( a17417a  and  a17410a );
 a17422a <=( (not A167)  and  A168 );
 a17423a <=( A170  and  a17422a );
 a17427a <=( (not A200)  and  (not A199) );
 a17428a <=( A166  and  a17427a );
 a17429a <=( a17428a  and  a17423a );
 a17433a <=( A234  and  A233 );
 a17434a <=( A203  and  a17433a );
 a17437a <=( (not A299)  and  (not A298) );
 a17440a <=( (not A302)  and  A301 );
 a17441a <=( a17440a  and  a17437a );
 a17442a <=( a17441a  and  a17434a );
 a17446a <=( (not A167)  and  A168 );
 a17447a <=( A170  and  a17446a );
 a17451a <=( (not A200)  and  (not A199) );
 a17452a <=( A166  and  a17451a );
 a17453a <=( a17452a  and  a17447a );
 a17457a <=( A234  and  A233 );
 a17458a <=( A203  and  a17457a );
 a17461a <=( A266  and  A265 );
 a17464a <=( (not A269)  and  A268 );
 a17465a <=( a17464a  and  a17461a );
 a17466a <=( a17465a  and  a17458a );
 a17470a <=( (not A167)  and  A168 );
 a17471a <=( A170  and  a17470a );
 a17475a <=( (not A200)  and  (not A199) );
 a17476a <=( A166  and  a17475a );
 a17477a <=( a17476a  and  a17471a );
 a17481a <=( A234  and  A233 );
 a17482a <=( A203  and  a17481a );
 a17485a <=( A266  and  (not A265) );
 a17488a <=( A269  and  (not A268) );
 a17489a <=( a17488a  and  a17485a );
 a17490a <=( a17489a  and  a17482a );
 a17494a <=( (not A167)  and  A168 );
 a17495a <=( A170  and  a17494a );
 a17499a <=( (not A200)  and  (not A199) );
 a17500a <=( A166  and  a17499a );
 a17501a <=( a17500a  and  a17495a );
 a17505a <=( A234  and  A233 );
 a17506a <=( A203  and  a17505a );
 a17509a <=( (not A266)  and  A265 );
 a17512a <=( A269  and  (not A268) );
 a17513a <=( a17512a  and  a17509a );
 a17514a <=( a17513a  and  a17506a );
 a17518a <=( (not A167)  and  A168 );
 a17519a <=( A170  and  a17518a );
 a17523a <=( (not A200)  and  (not A199) );
 a17524a <=( A166  and  a17523a );
 a17525a <=( a17524a  and  a17519a );
 a17529a <=( A234  and  A233 );
 a17530a <=( A203  and  a17529a );
 a17533a <=( (not A266)  and  (not A265) );
 a17536a <=( (not A269)  and  A268 );
 a17537a <=( a17536a  and  a17533a );
 a17538a <=( a17537a  and  a17530a );
 a17542a <=( (not A167)  and  A168 );
 a17543a <=( A170  and  a17542a );
 a17547a <=( (not A200)  and  (not A199) );
 a17548a <=( A166  and  a17547a );
 a17549a <=( a17548a  and  a17543a );
 a17553a <=( A233  and  A232 );
 a17554a <=( A203  and  a17553a );
 a17557a <=( (not A236)  and  A235 );
 a17560a <=( A300  and  A299 );
 a17561a <=( a17560a  and  a17557a );
 a17562a <=( a17561a  and  a17554a );
 a17566a <=( (not A167)  and  A168 );
 a17567a <=( A170  and  a17566a );
 a17571a <=( (not A200)  and  (not A199) );
 a17572a <=( A166  and  a17571a );
 a17573a <=( a17572a  and  a17567a );
 a17577a <=( A233  and  A232 );
 a17578a <=( A203  and  a17577a );
 a17581a <=( (not A236)  and  A235 );
 a17584a <=( A300  and  A298 );
 a17585a <=( a17584a  and  a17581a );
 a17586a <=( a17585a  and  a17578a );
 a17590a <=( (not A167)  and  A168 );
 a17591a <=( A170  and  a17590a );
 a17595a <=( (not A200)  and  (not A199) );
 a17596a <=( A166  and  a17595a );
 a17597a <=( a17596a  and  a17591a );
 a17601a <=( A233  and  A232 );
 a17602a <=( A203  and  a17601a );
 a17605a <=( (not A236)  and  A235 );
 a17608a <=( A267  and  A265 );
 a17609a <=( a17608a  and  a17605a );
 a17610a <=( a17609a  and  a17602a );
 a17614a <=( (not A167)  and  A168 );
 a17615a <=( A170  and  a17614a );
 a17619a <=( (not A200)  and  (not A199) );
 a17620a <=( A166  and  a17619a );
 a17621a <=( a17620a  and  a17615a );
 a17625a <=( A233  and  A232 );
 a17626a <=( A203  and  a17625a );
 a17629a <=( (not A236)  and  A235 );
 a17632a <=( A267  and  A266 );
 a17633a <=( a17632a  and  a17629a );
 a17634a <=( a17633a  and  a17626a );
 a17638a <=( (not A167)  and  A168 );
 a17639a <=( A170  and  a17638a );
 a17643a <=( (not A200)  and  (not A199) );
 a17644a <=( A166  and  a17643a );
 a17645a <=( a17644a  and  a17639a );
 a17649a <=( A233  and  (not A232) );
 a17650a <=( A203  and  a17649a );
 a17653a <=( A236  and  (not A235) );
 a17656a <=( A300  and  A299 );
 a17657a <=( a17656a  and  a17653a );
 a17658a <=( a17657a  and  a17650a );
 a17662a <=( (not A167)  and  A168 );
 a17663a <=( A170  and  a17662a );
 a17667a <=( (not A200)  and  (not A199) );
 a17668a <=( A166  and  a17667a );
 a17669a <=( a17668a  and  a17663a );
 a17673a <=( A233  and  (not A232) );
 a17674a <=( A203  and  a17673a );
 a17677a <=( A236  and  (not A235) );
 a17680a <=( A300  and  A298 );
 a17681a <=( a17680a  and  a17677a );
 a17682a <=( a17681a  and  a17674a );
 a17686a <=( (not A167)  and  A168 );
 a17687a <=( A170  and  a17686a );
 a17691a <=( (not A200)  and  (not A199) );
 a17692a <=( A166  and  a17691a );
 a17693a <=( a17692a  and  a17687a );
 a17697a <=( A233  and  (not A232) );
 a17698a <=( A203  and  a17697a );
 a17701a <=( A236  and  (not A235) );
 a17704a <=( A267  and  A265 );
 a17705a <=( a17704a  and  a17701a );
 a17706a <=( a17705a  and  a17698a );
 a17710a <=( (not A167)  and  A168 );
 a17711a <=( A170  and  a17710a );
 a17715a <=( (not A200)  and  (not A199) );
 a17716a <=( A166  and  a17715a );
 a17717a <=( a17716a  and  a17711a );
 a17721a <=( A233  and  (not A232) );
 a17722a <=( A203  and  a17721a );
 a17725a <=( A236  and  (not A235) );
 a17728a <=( A267  and  A266 );
 a17729a <=( a17728a  and  a17725a );
 a17730a <=( a17729a  and  a17722a );
 a17734a <=( (not A167)  and  A168 );
 a17735a <=( A170  and  a17734a );
 a17739a <=( (not A200)  and  (not A199) );
 a17740a <=( A166  and  a17739a );
 a17741a <=( a17740a  and  a17735a );
 a17745a <=( (not A233)  and  A232 );
 a17746a <=( A203  and  a17745a );
 a17749a <=( A236  and  (not A235) );
 a17752a <=( A300  and  A299 );
 a17753a <=( a17752a  and  a17749a );
 a17754a <=( a17753a  and  a17746a );
 a17758a <=( (not A167)  and  A168 );
 a17759a <=( A170  and  a17758a );
 a17763a <=( (not A200)  and  (not A199) );
 a17764a <=( A166  and  a17763a );
 a17765a <=( a17764a  and  a17759a );
 a17769a <=( (not A233)  and  A232 );
 a17770a <=( A203  and  a17769a );
 a17773a <=( A236  and  (not A235) );
 a17776a <=( A300  and  A298 );
 a17777a <=( a17776a  and  a17773a );
 a17778a <=( a17777a  and  a17770a );
 a17782a <=( (not A167)  and  A168 );
 a17783a <=( A170  and  a17782a );
 a17787a <=( (not A200)  and  (not A199) );
 a17788a <=( A166  and  a17787a );
 a17789a <=( a17788a  and  a17783a );
 a17793a <=( (not A233)  and  A232 );
 a17794a <=( A203  and  a17793a );
 a17797a <=( A236  and  (not A235) );
 a17800a <=( A267  and  A265 );
 a17801a <=( a17800a  and  a17797a );
 a17802a <=( a17801a  and  a17794a );
 a17806a <=( (not A167)  and  A168 );
 a17807a <=( A170  and  a17806a );
 a17811a <=( (not A200)  and  (not A199) );
 a17812a <=( A166  and  a17811a );
 a17813a <=( a17812a  and  a17807a );
 a17817a <=( (not A233)  and  A232 );
 a17818a <=( A203  and  a17817a );
 a17821a <=( A236  and  (not A235) );
 a17824a <=( A267  and  A266 );
 a17825a <=( a17824a  and  a17821a );
 a17826a <=( a17825a  and  a17818a );
 a17830a <=( (not A167)  and  A168 );
 a17831a <=( A170  and  a17830a );
 a17835a <=( (not A200)  and  (not A199) );
 a17836a <=( A166  and  a17835a );
 a17837a <=( a17836a  and  a17831a );
 a17841a <=( (not A233)  and  (not A232) );
 a17842a <=( A203  and  a17841a );
 a17845a <=( (not A236)  and  A235 );
 a17848a <=( A300  and  A299 );
 a17849a <=( a17848a  and  a17845a );
 a17850a <=( a17849a  and  a17842a );
 a17854a <=( (not A167)  and  A168 );
 a17855a <=( A170  and  a17854a );
 a17859a <=( (not A200)  and  (not A199) );
 a17860a <=( A166  and  a17859a );
 a17861a <=( a17860a  and  a17855a );
 a17865a <=( (not A233)  and  (not A232) );
 a17866a <=( A203  and  a17865a );
 a17869a <=( (not A236)  and  A235 );
 a17872a <=( A300  and  A298 );
 a17873a <=( a17872a  and  a17869a );
 a17874a <=( a17873a  and  a17866a );
 a17878a <=( (not A167)  and  A168 );
 a17879a <=( A170  and  a17878a );
 a17883a <=( (not A200)  and  (not A199) );
 a17884a <=( A166  and  a17883a );
 a17885a <=( a17884a  and  a17879a );
 a17889a <=( (not A233)  and  (not A232) );
 a17890a <=( A203  and  a17889a );
 a17893a <=( (not A236)  and  A235 );
 a17896a <=( A267  and  A265 );
 a17897a <=( a17896a  and  a17893a );
 a17898a <=( a17897a  and  a17890a );
 a17902a <=( (not A167)  and  A168 );
 a17903a <=( A170  and  a17902a );
 a17907a <=( (not A200)  and  (not A199) );
 a17908a <=( A166  and  a17907a );
 a17909a <=( a17908a  and  a17903a );
 a17913a <=( (not A233)  and  (not A232) );
 a17914a <=( A203  and  a17913a );
 a17917a <=( (not A236)  and  A235 );
 a17920a <=( A267  and  A266 );
 a17921a <=( a17920a  and  a17917a );
 a17922a <=( a17921a  and  a17914a );
 a17926a <=( (not A167)  and  A168 );
 a17927a <=( A169  and  a17926a );
 a17931a <=( (not A200)  and  (not A199) );
 a17932a <=( A166  and  a17931a );
 a17933a <=( a17932a  and  a17927a );
 a17937a <=( A234  and  A232 );
 a17938a <=( (not A202)  and  a17937a );
 a17941a <=( A299  and  A298 );
 a17944a <=( (not A302)  and  A301 );
 a17945a <=( a17944a  and  a17941a );
 a17946a <=( a17945a  and  a17938a );
 a17950a <=( (not A167)  and  A168 );
 a17951a <=( A169  and  a17950a );
 a17955a <=( (not A200)  and  (not A199) );
 a17956a <=( A166  and  a17955a );
 a17957a <=( a17956a  and  a17951a );
 a17961a <=( A234  and  A232 );
 a17962a <=( (not A202)  and  a17961a );
 a17965a <=( (not A299)  and  A298 );
 a17968a <=( A302  and  (not A301) );
 a17969a <=( a17968a  and  a17965a );
 a17970a <=( a17969a  and  a17962a );
 a17974a <=( (not A167)  and  A168 );
 a17975a <=( A169  and  a17974a );
 a17979a <=( (not A200)  and  (not A199) );
 a17980a <=( A166  and  a17979a );
 a17981a <=( a17980a  and  a17975a );
 a17985a <=( A234  and  A232 );
 a17986a <=( (not A202)  and  a17985a );
 a17989a <=( A299  and  (not A298) );
 a17992a <=( A302  and  (not A301) );
 a17993a <=( a17992a  and  a17989a );
 a17994a <=( a17993a  and  a17986a );
 a17998a <=( (not A167)  and  A168 );
 a17999a <=( A169  and  a17998a );
 a18003a <=( (not A200)  and  (not A199) );
 a18004a <=( A166  and  a18003a );
 a18005a <=( a18004a  and  a17999a );
 a18009a <=( A234  and  A232 );
 a18010a <=( (not A202)  and  a18009a );
 a18013a <=( (not A299)  and  (not A298) );
 a18016a <=( (not A302)  and  A301 );
 a18017a <=( a18016a  and  a18013a );
 a18018a <=( a18017a  and  a18010a );
 a18022a <=( (not A167)  and  A168 );
 a18023a <=( A169  and  a18022a );
 a18027a <=( (not A200)  and  (not A199) );
 a18028a <=( A166  and  a18027a );
 a18029a <=( a18028a  and  a18023a );
 a18033a <=( A234  and  A232 );
 a18034a <=( (not A202)  and  a18033a );
 a18037a <=( A266  and  A265 );
 a18040a <=( (not A269)  and  A268 );
 a18041a <=( a18040a  and  a18037a );
 a18042a <=( a18041a  and  a18034a );
 a18046a <=( (not A167)  and  A168 );
 a18047a <=( A169  and  a18046a );
 a18051a <=( (not A200)  and  (not A199) );
 a18052a <=( A166  and  a18051a );
 a18053a <=( a18052a  and  a18047a );
 a18057a <=( A234  and  A232 );
 a18058a <=( (not A202)  and  a18057a );
 a18061a <=( A266  and  (not A265) );
 a18064a <=( A269  and  (not A268) );
 a18065a <=( a18064a  and  a18061a );
 a18066a <=( a18065a  and  a18058a );
 a18070a <=( (not A167)  and  A168 );
 a18071a <=( A169  and  a18070a );
 a18075a <=( (not A200)  and  (not A199) );
 a18076a <=( A166  and  a18075a );
 a18077a <=( a18076a  and  a18071a );
 a18081a <=( A234  and  A232 );
 a18082a <=( (not A202)  and  a18081a );
 a18085a <=( (not A266)  and  A265 );
 a18088a <=( A269  and  (not A268) );
 a18089a <=( a18088a  and  a18085a );
 a18090a <=( a18089a  and  a18082a );
 a18094a <=( (not A167)  and  A168 );
 a18095a <=( A169  and  a18094a );
 a18099a <=( (not A200)  and  (not A199) );
 a18100a <=( A166  and  a18099a );
 a18101a <=( a18100a  and  a18095a );
 a18105a <=( A234  and  A232 );
 a18106a <=( (not A202)  and  a18105a );
 a18109a <=( (not A266)  and  (not A265) );
 a18112a <=( (not A269)  and  A268 );
 a18113a <=( a18112a  and  a18109a );
 a18114a <=( a18113a  and  a18106a );
 a18118a <=( (not A167)  and  A168 );
 a18119a <=( A169  and  a18118a );
 a18123a <=( (not A200)  and  (not A199) );
 a18124a <=( A166  and  a18123a );
 a18125a <=( a18124a  and  a18119a );
 a18129a <=( A234  and  A233 );
 a18130a <=( (not A202)  and  a18129a );
 a18133a <=( A299  and  A298 );
 a18136a <=( (not A302)  and  A301 );
 a18137a <=( a18136a  and  a18133a );
 a18138a <=( a18137a  and  a18130a );
 a18142a <=( (not A167)  and  A168 );
 a18143a <=( A169  and  a18142a );
 a18147a <=( (not A200)  and  (not A199) );
 a18148a <=( A166  and  a18147a );
 a18149a <=( a18148a  and  a18143a );
 a18153a <=( A234  and  A233 );
 a18154a <=( (not A202)  and  a18153a );
 a18157a <=( (not A299)  and  A298 );
 a18160a <=( A302  and  (not A301) );
 a18161a <=( a18160a  and  a18157a );
 a18162a <=( a18161a  and  a18154a );
 a18166a <=( (not A167)  and  A168 );
 a18167a <=( A169  and  a18166a );
 a18171a <=( (not A200)  and  (not A199) );
 a18172a <=( A166  and  a18171a );
 a18173a <=( a18172a  and  a18167a );
 a18177a <=( A234  and  A233 );
 a18178a <=( (not A202)  and  a18177a );
 a18181a <=( A299  and  (not A298) );
 a18184a <=( A302  and  (not A301) );
 a18185a <=( a18184a  and  a18181a );
 a18186a <=( a18185a  and  a18178a );
 a18190a <=( (not A167)  and  A168 );
 a18191a <=( A169  and  a18190a );
 a18195a <=( (not A200)  and  (not A199) );
 a18196a <=( A166  and  a18195a );
 a18197a <=( a18196a  and  a18191a );
 a18201a <=( A234  and  A233 );
 a18202a <=( (not A202)  and  a18201a );
 a18205a <=( (not A299)  and  (not A298) );
 a18208a <=( (not A302)  and  A301 );
 a18209a <=( a18208a  and  a18205a );
 a18210a <=( a18209a  and  a18202a );
 a18214a <=( (not A167)  and  A168 );
 a18215a <=( A169  and  a18214a );
 a18219a <=( (not A200)  and  (not A199) );
 a18220a <=( A166  and  a18219a );
 a18221a <=( a18220a  and  a18215a );
 a18225a <=( A234  and  A233 );
 a18226a <=( (not A202)  and  a18225a );
 a18229a <=( A266  and  A265 );
 a18232a <=( (not A269)  and  A268 );
 a18233a <=( a18232a  and  a18229a );
 a18234a <=( a18233a  and  a18226a );
 a18238a <=( (not A167)  and  A168 );
 a18239a <=( A169  and  a18238a );
 a18243a <=( (not A200)  and  (not A199) );
 a18244a <=( A166  and  a18243a );
 a18245a <=( a18244a  and  a18239a );
 a18249a <=( A234  and  A233 );
 a18250a <=( (not A202)  and  a18249a );
 a18253a <=( A266  and  (not A265) );
 a18256a <=( A269  and  (not A268) );
 a18257a <=( a18256a  and  a18253a );
 a18258a <=( a18257a  and  a18250a );
 a18262a <=( (not A167)  and  A168 );
 a18263a <=( A169  and  a18262a );
 a18267a <=( (not A200)  and  (not A199) );
 a18268a <=( A166  and  a18267a );
 a18269a <=( a18268a  and  a18263a );
 a18273a <=( A234  and  A233 );
 a18274a <=( (not A202)  and  a18273a );
 a18277a <=( (not A266)  and  A265 );
 a18280a <=( A269  and  (not A268) );
 a18281a <=( a18280a  and  a18277a );
 a18282a <=( a18281a  and  a18274a );
 a18286a <=( (not A167)  and  A168 );
 a18287a <=( A169  and  a18286a );
 a18291a <=( (not A200)  and  (not A199) );
 a18292a <=( A166  and  a18291a );
 a18293a <=( a18292a  and  a18287a );
 a18297a <=( A234  and  A233 );
 a18298a <=( (not A202)  and  a18297a );
 a18301a <=( (not A266)  and  (not A265) );
 a18304a <=( (not A269)  and  A268 );
 a18305a <=( a18304a  and  a18301a );
 a18306a <=( a18305a  and  a18298a );
 a18310a <=( (not A167)  and  A168 );
 a18311a <=( A169  and  a18310a );
 a18315a <=( (not A200)  and  (not A199) );
 a18316a <=( A166  and  a18315a );
 a18317a <=( a18316a  and  a18311a );
 a18321a <=( A233  and  A232 );
 a18322a <=( (not A202)  and  a18321a );
 a18325a <=( (not A236)  and  A235 );
 a18328a <=( A300  and  A299 );
 a18329a <=( a18328a  and  a18325a );
 a18330a <=( a18329a  and  a18322a );
 a18334a <=( (not A167)  and  A168 );
 a18335a <=( A169  and  a18334a );
 a18339a <=( (not A200)  and  (not A199) );
 a18340a <=( A166  and  a18339a );
 a18341a <=( a18340a  and  a18335a );
 a18345a <=( A233  and  A232 );
 a18346a <=( (not A202)  and  a18345a );
 a18349a <=( (not A236)  and  A235 );
 a18352a <=( A300  and  A298 );
 a18353a <=( a18352a  and  a18349a );
 a18354a <=( a18353a  and  a18346a );
 a18358a <=( (not A167)  and  A168 );
 a18359a <=( A169  and  a18358a );
 a18363a <=( (not A200)  and  (not A199) );
 a18364a <=( A166  and  a18363a );
 a18365a <=( a18364a  and  a18359a );
 a18369a <=( A233  and  A232 );
 a18370a <=( (not A202)  and  a18369a );
 a18373a <=( (not A236)  and  A235 );
 a18376a <=( A267  and  A265 );
 a18377a <=( a18376a  and  a18373a );
 a18378a <=( a18377a  and  a18370a );
 a18382a <=( (not A167)  and  A168 );
 a18383a <=( A169  and  a18382a );
 a18387a <=( (not A200)  and  (not A199) );
 a18388a <=( A166  and  a18387a );
 a18389a <=( a18388a  and  a18383a );
 a18393a <=( A233  and  A232 );
 a18394a <=( (not A202)  and  a18393a );
 a18397a <=( (not A236)  and  A235 );
 a18400a <=( A267  and  A266 );
 a18401a <=( a18400a  and  a18397a );
 a18402a <=( a18401a  and  a18394a );
 a18406a <=( (not A167)  and  A168 );
 a18407a <=( A169  and  a18406a );
 a18411a <=( (not A200)  and  (not A199) );
 a18412a <=( A166  and  a18411a );
 a18413a <=( a18412a  and  a18407a );
 a18417a <=( A233  and  (not A232) );
 a18418a <=( (not A202)  and  a18417a );
 a18421a <=( A236  and  (not A235) );
 a18424a <=( A300  and  A299 );
 a18425a <=( a18424a  and  a18421a );
 a18426a <=( a18425a  and  a18418a );
 a18430a <=( (not A167)  and  A168 );
 a18431a <=( A169  and  a18430a );
 a18435a <=( (not A200)  and  (not A199) );
 a18436a <=( A166  and  a18435a );
 a18437a <=( a18436a  and  a18431a );
 a18441a <=( A233  and  (not A232) );
 a18442a <=( (not A202)  and  a18441a );
 a18445a <=( A236  and  (not A235) );
 a18448a <=( A300  and  A298 );
 a18449a <=( a18448a  and  a18445a );
 a18450a <=( a18449a  and  a18442a );
 a18454a <=( (not A167)  and  A168 );
 a18455a <=( A169  and  a18454a );
 a18459a <=( (not A200)  and  (not A199) );
 a18460a <=( A166  and  a18459a );
 a18461a <=( a18460a  and  a18455a );
 a18465a <=( A233  and  (not A232) );
 a18466a <=( (not A202)  and  a18465a );
 a18469a <=( A236  and  (not A235) );
 a18472a <=( A267  and  A265 );
 a18473a <=( a18472a  and  a18469a );
 a18474a <=( a18473a  and  a18466a );
 a18478a <=( (not A167)  and  A168 );
 a18479a <=( A169  and  a18478a );
 a18483a <=( (not A200)  and  (not A199) );
 a18484a <=( A166  and  a18483a );
 a18485a <=( a18484a  and  a18479a );
 a18489a <=( A233  and  (not A232) );
 a18490a <=( (not A202)  and  a18489a );
 a18493a <=( A236  and  (not A235) );
 a18496a <=( A267  and  A266 );
 a18497a <=( a18496a  and  a18493a );
 a18498a <=( a18497a  and  a18490a );
 a18502a <=( (not A167)  and  A168 );
 a18503a <=( A169  and  a18502a );
 a18507a <=( (not A200)  and  (not A199) );
 a18508a <=( A166  and  a18507a );
 a18509a <=( a18508a  and  a18503a );
 a18513a <=( (not A233)  and  A232 );
 a18514a <=( (not A202)  and  a18513a );
 a18517a <=( A236  and  (not A235) );
 a18520a <=( A300  and  A299 );
 a18521a <=( a18520a  and  a18517a );
 a18522a <=( a18521a  and  a18514a );
 a18526a <=( (not A167)  and  A168 );
 a18527a <=( A169  and  a18526a );
 a18531a <=( (not A200)  and  (not A199) );
 a18532a <=( A166  and  a18531a );
 a18533a <=( a18532a  and  a18527a );
 a18537a <=( (not A233)  and  A232 );
 a18538a <=( (not A202)  and  a18537a );
 a18541a <=( A236  and  (not A235) );
 a18544a <=( A300  and  A298 );
 a18545a <=( a18544a  and  a18541a );
 a18546a <=( a18545a  and  a18538a );
 a18550a <=( (not A167)  and  A168 );
 a18551a <=( A169  and  a18550a );
 a18555a <=( (not A200)  and  (not A199) );
 a18556a <=( A166  and  a18555a );
 a18557a <=( a18556a  and  a18551a );
 a18561a <=( (not A233)  and  A232 );
 a18562a <=( (not A202)  and  a18561a );
 a18565a <=( A236  and  (not A235) );
 a18568a <=( A267  and  A265 );
 a18569a <=( a18568a  and  a18565a );
 a18570a <=( a18569a  and  a18562a );
 a18574a <=( (not A167)  and  A168 );
 a18575a <=( A169  and  a18574a );
 a18579a <=( (not A200)  and  (not A199) );
 a18580a <=( A166  and  a18579a );
 a18581a <=( a18580a  and  a18575a );
 a18585a <=( (not A233)  and  A232 );
 a18586a <=( (not A202)  and  a18585a );
 a18589a <=( A236  and  (not A235) );
 a18592a <=( A267  and  A266 );
 a18593a <=( a18592a  and  a18589a );
 a18594a <=( a18593a  and  a18586a );
 a18598a <=( (not A167)  and  A168 );
 a18599a <=( A169  and  a18598a );
 a18603a <=( (not A200)  and  (not A199) );
 a18604a <=( A166  and  a18603a );
 a18605a <=( a18604a  and  a18599a );
 a18609a <=( (not A233)  and  (not A232) );
 a18610a <=( (not A202)  and  a18609a );
 a18613a <=( (not A236)  and  A235 );
 a18616a <=( A300  and  A299 );
 a18617a <=( a18616a  and  a18613a );
 a18618a <=( a18617a  and  a18610a );
 a18622a <=( (not A167)  and  A168 );
 a18623a <=( A169  and  a18622a );
 a18627a <=( (not A200)  and  (not A199) );
 a18628a <=( A166  and  a18627a );
 a18629a <=( a18628a  and  a18623a );
 a18633a <=( (not A233)  and  (not A232) );
 a18634a <=( (not A202)  and  a18633a );
 a18637a <=( (not A236)  and  A235 );
 a18640a <=( A300  and  A298 );
 a18641a <=( a18640a  and  a18637a );
 a18642a <=( a18641a  and  a18634a );
 a18646a <=( (not A167)  and  A168 );
 a18647a <=( A169  and  a18646a );
 a18651a <=( (not A200)  and  (not A199) );
 a18652a <=( A166  and  a18651a );
 a18653a <=( a18652a  and  a18647a );
 a18657a <=( (not A233)  and  (not A232) );
 a18658a <=( (not A202)  and  a18657a );
 a18661a <=( (not A236)  and  A235 );
 a18664a <=( A267  and  A265 );
 a18665a <=( a18664a  and  a18661a );
 a18666a <=( a18665a  and  a18658a );
 a18670a <=( (not A167)  and  A168 );
 a18671a <=( A169  and  a18670a );
 a18675a <=( (not A200)  and  (not A199) );
 a18676a <=( A166  and  a18675a );
 a18677a <=( a18676a  and  a18671a );
 a18681a <=( (not A233)  and  (not A232) );
 a18682a <=( (not A202)  and  a18681a );
 a18685a <=( (not A236)  and  A235 );
 a18688a <=( A267  and  A266 );
 a18689a <=( a18688a  and  a18685a );
 a18690a <=( a18689a  and  a18682a );
 a18694a <=( (not A167)  and  A168 );
 a18695a <=( A169  and  a18694a );
 a18699a <=( (not A200)  and  (not A199) );
 a18700a <=( A166  and  a18699a );
 a18701a <=( a18700a  and  a18695a );
 a18705a <=( A234  and  A232 );
 a18706a <=( A203  and  a18705a );
 a18709a <=( A299  and  A298 );
 a18712a <=( (not A302)  and  A301 );
 a18713a <=( a18712a  and  a18709a );
 a18714a <=( a18713a  and  a18706a );
 a18718a <=( (not A167)  and  A168 );
 a18719a <=( A169  and  a18718a );
 a18723a <=( (not A200)  and  (not A199) );
 a18724a <=( A166  and  a18723a );
 a18725a <=( a18724a  and  a18719a );
 a18729a <=( A234  and  A232 );
 a18730a <=( A203  and  a18729a );
 a18733a <=( (not A299)  and  A298 );
 a18736a <=( A302  and  (not A301) );
 a18737a <=( a18736a  and  a18733a );
 a18738a <=( a18737a  and  a18730a );
 a18742a <=( (not A167)  and  A168 );
 a18743a <=( A169  and  a18742a );
 a18747a <=( (not A200)  and  (not A199) );
 a18748a <=( A166  and  a18747a );
 a18749a <=( a18748a  and  a18743a );
 a18753a <=( A234  and  A232 );
 a18754a <=( A203  and  a18753a );
 a18757a <=( A299  and  (not A298) );
 a18760a <=( A302  and  (not A301) );
 a18761a <=( a18760a  and  a18757a );
 a18762a <=( a18761a  and  a18754a );
 a18766a <=( (not A167)  and  A168 );
 a18767a <=( A169  and  a18766a );
 a18771a <=( (not A200)  and  (not A199) );
 a18772a <=( A166  and  a18771a );
 a18773a <=( a18772a  and  a18767a );
 a18777a <=( A234  and  A232 );
 a18778a <=( A203  and  a18777a );
 a18781a <=( (not A299)  and  (not A298) );
 a18784a <=( (not A302)  and  A301 );
 a18785a <=( a18784a  and  a18781a );
 a18786a <=( a18785a  and  a18778a );
 a18790a <=( (not A167)  and  A168 );
 a18791a <=( A169  and  a18790a );
 a18795a <=( (not A200)  and  (not A199) );
 a18796a <=( A166  and  a18795a );
 a18797a <=( a18796a  and  a18791a );
 a18801a <=( A234  and  A232 );
 a18802a <=( A203  and  a18801a );
 a18805a <=( A266  and  A265 );
 a18808a <=( (not A269)  and  A268 );
 a18809a <=( a18808a  and  a18805a );
 a18810a <=( a18809a  and  a18802a );
 a18814a <=( (not A167)  and  A168 );
 a18815a <=( A169  and  a18814a );
 a18819a <=( (not A200)  and  (not A199) );
 a18820a <=( A166  and  a18819a );
 a18821a <=( a18820a  and  a18815a );
 a18825a <=( A234  and  A232 );
 a18826a <=( A203  and  a18825a );
 a18829a <=( A266  and  (not A265) );
 a18832a <=( A269  and  (not A268) );
 a18833a <=( a18832a  and  a18829a );
 a18834a <=( a18833a  and  a18826a );
 a18838a <=( (not A167)  and  A168 );
 a18839a <=( A169  and  a18838a );
 a18843a <=( (not A200)  and  (not A199) );
 a18844a <=( A166  and  a18843a );
 a18845a <=( a18844a  and  a18839a );
 a18849a <=( A234  and  A232 );
 a18850a <=( A203  and  a18849a );
 a18853a <=( (not A266)  and  A265 );
 a18856a <=( A269  and  (not A268) );
 a18857a <=( a18856a  and  a18853a );
 a18858a <=( a18857a  and  a18850a );
 a18862a <=( (not A167)  and  A168 );
 a18863a <=( A169  and  a18862a );
 a18867a <=( (not A200)  and  (not A199) );
 a18868a <=( A166  and  a18867a );
 a18869a <=( a18868a  and  a18863a );
 a18873a <=( A234  and  A232 );
 a18874a <=( A203  and  a18873a );
 a18877a <=( (not A266)  and  (not A265) );
 a18880a <=( (not A269)  and  A268 );
 a18881a <=( a18880a  and  a18877a );
 a18882a <=( a18881a  and  a18874a );
 a18886a <=( (not A167)  and  A168 );
 a18887a <=( A169  and  a18886a );
 a18891a <=( (not A200)  and  (not A199) );
 a18892a <=( A166  and  a18891a );
 a18893a <=( a18892a  and  a18887a );
 a18897a <=( A234  and  A233 );
 a18898a <=( A203  and  a18897a );
 a18901a <=( A299  and  A298 );
 a18904a <=( (not A302)  and  A301 );
 a18905a <=( a18904a  and  a18901a );
 a18906a <=( a18905a  and  a18898a );
 a18910a <=( (not A167)  and  A168 );
 a18911a <=( A169  and  a18910a );
 a18915a <=( (not A200)  and  (not A199) );
 a18916a <=( A166  and  a18915a );
 a18917a <=( a18916a  and  a18911a );
 a18921a <=( A234  and  A233 );
 a18922a <=( A203  and  a18921a );
 a18925a <=( (not A299)  and  A298 );
 a18928a <=( A302  and  (not A301) );
 a18929a <=( a18928a  and  a18925a );
 a18930a <=( a18929a  and  a18922a );
 a18934a <=( (not A167)  and  A168 );
 a18935a <=( A169  and  a18934a );
 a18939a <=( (not A200)  and  (not A199) );
 a18940a <=( A166  and  a18939a );
 a18941a <=( a18940a  and  a18935a );
 a18945a <=( A234  and  A233 );
 a18946a <=( A203  and  a18945a );
 a18949a <=( A299  and  (not A298) );
 a18952a <=( A302  and  (not A301) );
 a18953a <=( a18952a  and  a18949a );
 a18954a <=( a18953a  and  a18946a );
 a18958a <=( (not A167)  and  A168 );
 a18959a <=( A169  and  a18958a );
 a18963a <=( (not A200)  and  (not A199) );
 a18964a <=( A166  and  a18963a );
 a18965a <=( a18964a  and  a18959a );
 a18969a <=( A234  and  A233 );
 a18970a <=( A203  and  a18969a );
 a18973a <=( (not A299)  and  (not A298) );
 a18976a <=( (not A302)  and  A301 );
 a18977a <=( a18976a  and  a18973a );
 a18978a <=( a18977a  and  a18970a );
 a18982a <=( (not A167)  and  A168 );
 a18983a <=( A169  and  a18982a );
 a18987a <=( (not A200)  and  (not A199) );
 a18988a <=( A166  and  a18987a );
 a18989a <=( a18988a  and  a18983a );
 a18993a <=( A234  and  A233 );
 a18994a <=( A203  and  a18993a );
 a18997a <=( A266  and  A265 );
 a19000a <=( (not A269)  and  A268 );
 a19001a <=( a19000a  and  a18997a );
 a19002a <=( a19001a  and  a18994a );
 a19006a <=( (not A167)  and  A168 );
 a19007a <=( A169  and  a19006a );
 a19011a <=( (not A200)  and  (not A199) );
 a19012a <=( A166  and  a19011a );
 a19013a <=( a19012a  and  a19007a );
 a19017a <=( A234  and  A233 );
 a19018a <=( A203  and  a19017a );
 a19021a <=( A266  and  (not A265) );
 a19024a <=( A269  and  (not A268) );
 a19025a <=( a19024a  and  a19021a );
 a19026a <=( a19025a  and  a19018a );
 a19030a <=( (not A167)  and  A168 );
 a19031a <=( A169  and  a19030a );
 a19035a <=( (not A200)  and  (not A199) );
 a19036a <=( A166  and  a19035a );
 a19037a <=( a19036a  and  a19031a );
 a19041a <=( A234  and  A233 );
 a19042a <=( A203  and  a19041a );
 a19045a <=( (not A266)  and  A265 );
 a19048a <=( A269  and  (not A268) );
 a19049a <=( a19048a  and  a19045a );
 a19050a <=( a19049a  and  a19042a );
 a19054a <=( (not A167)  and  A168 );
 a19055a <=( A169  and  a19054a );
 a19059a <=( (not A200)  and  (not A199) );
 a19060a <=( A166  and  a19059a );
 a19061a <=( a19060a  and  a19055a );
 a19065a <=( A234  and  A233 );
 a19066a <=( A203  and  a19065a );
 a19069a <=( (not A266)  and  (not A265) );
 a19072a <=( (not A269)  and  A268 );
 a19073a <=( a19072a  and  a19069a );
 a19074a <=( a19073a  and  a19066a );
 a19078a <=( (not A167)  and  A168 );
 a19079a <=( A169  and  a19078a );
 a19083a <=( (not A200)  and  (not A199) );
 a19084a <=( A166  and  a19083a );
 a19085a <=( a19084a  and  a19079a );
 a19089a <=( A233  and  A232 );
 a19090a <=( A203  and  a19089a );
 a19093a <=( (not A236)  and  A235 );
 a19096a <=( A300  and  A299 );
 a19097a <=( a19096a  and  a19093a );
 a19098a <=( a19097a  and  a19090a );
 a19102a <=( (not A167)  and  A168 );
 a19103a <=( A169  and  a19102a );
 a19107a <=( (not A200)  and  (not A199) );
 a19108a <=( A166  and  a19107a );
 a19109a <=( a19108a  and  a19103a );
 a19113a <=( A233  and  A232 );
 a19114a <=( A203  and  a19113a );
 a19117a <=( (not A236)  and  A235 );
 a19120a <=( A300  and  A298 );
 a19121a <=( a19120a  and  a19117a );
 a19122a <=( a19121a  and  a19114a );
 a19126a <=( (not A167)  and  A168 );
 a19127a <=( A169  and  a19126a );
 a19131a <=( (not A200)  and  (not A199) );
 a19132a <=( A166  and  a19131a );
 a19133a <=( a19132a  and  a19127a );
 a19137a <=( A233  and  A232 );
 a19138a <=( A203  and  a19137a );
 a19141a <=( (not A236)  and  A235 );
 a19144a <=( A267  and  A265 );
 a19145a <=( a19144a  and  a19141a );
 a19146a <=( a19145a  and  a19138a );
 a19150a <=( (not A167)  and  A168 );
 a19151a <=( A169  and  a19150a );
 a19155a <=( (not A200)  and  (not A199) );
 a19156a <=( A166  and  a19155a );
 a19157a <=( a19156a  and  a19151a );
 a19161a <=( A233  and  A232 );
 a19162a <=( A203  and  a19161a );
 a19165a <=( (not A236)  and  A235 );
 a19168a <=( A267  and  A266 );
 a19169a <=( a19168a  and  a19165a );
 a19170a <=( a19169a  and  a19162a );
 a19174a <=( (not A167)  and  A168 );
 a19175a <=( A169  and  a19174a );
 a19179a <=( (not A200)  and  (not A199) );
 a19180a <=( A166  and  a19179a );
 a19181a <=( a19180a  and  a19175a );
 a19185a <=( A233  and  (not A232) );
 a19186a <=( A203  and  a19185a );
 a19189a <=( A236  and  (not A235) );
 a19192a <=( A300  and  A299 );
 a19193a <=( a19192a  and  a19189a );
 a19194a <=( a19193a  and  a19186a );
 a19198a <=( (not A167)  and  A168 );
 a19199a <=( A169  and  a19198a );
 a19203a <=( (not A200)  and  (not A199) );
 a19204a <=( A166  and  a19203a );
 a19205a <=( a19204a  and  a19199a );
 a19209a <=( A233  and  (not A232) );
 a19210a <=( A203  and  a19209a );
 a19213a <=( A236  and  (not A235) );
 a19216a <=( A300  and  A298 );
 a19217a <=( a19216a  and  a19213a );
 a19218a <=( a19217a  and  a19210a );
 a19222a <=( (not A167)  and  A168 );
 a19223a <=( A169  and  a19222a );
 a19227a <=( (not A200)  and  (not A199) );
 a19228a <=( A166  and  a19227a );
 a19229a <=( a19228a  and  a19223a );
 a19233a <=( A233  and  (not A232) );
 a19234a <=( A203  and  a19233a );
 a19237a <=( A236  and  (not A235) );
 a19240a <=( A267  and  A265 );
 a19241a <=( a19240a  and  a19237a );
 a19242a <=( a19241a  and  a19234a );
 a19246a <=( (not A167)  and  A168 );
 a19247a <=( A169  and  a19246a );
 a19251a <=( (not A200)  and  (not A199) );
 a19252a <=( A166  and  a19251a );
 a19253a <=( a19252a  and  a19247a );
 a19257a <=( A233  and  (not A232) );
 a19258a <=( A203  and  a19257a );
 a19261a <=( A236  and  (not A235) );
 a19264a <=( A267  and  A266 );
 a19265a <=( a19264a  and  a19261a );
 a19266a <=( a19265a  and  a19258a );
 a19270a <=( (not A167)  and  A168 );
 a19271a <=( A169  and  a19270a );
 a19275a <=( (not A200)  and  (not A199) );
 a19276a <=( A166  and  a19275a );
 a19277a <=( a19276a  and  a19271a );
 a19281a <=( (not A233)  and  A232 );
 a19282a <=( A203  and  a19281a );
 a19285a <=( A236  and  (not A235) );
 a19288a <=( A300  and  A299 );
 a19289a <=( a19288a  and  a19285a );
 a19290a <=( a19289a  and  a19282a );
 a19294a <=( (not A167)  and  A168 );
 a19295a <=( A169  and  a19294a );
 a19299a <=( (not A200)  and  (not A199) );
 a19300a <=( A166  and  a19299a );
 a19301a <=( a19300a  and  a19295a );
 a19305a <=( (not A233)  and  A232 );
 a19306a <=( A203  and  a19305a );
 a19309a <=( A236  and  (not A235) );
 a19312a <=( A300  and  A298 );
 a19313a <=( a19312a  and  a19309a );
 a19314a <=( a19313a  and  a19306a );
 a19318a <=( (not A167)  and  A168 );
 a19319a <=( A169  and  a19318a );
 a19323a <=( (not A200)  and  (not A199) );
 a19324a <=( A166  and  a19323a );
 a19325a <=( a19324a  and  a19319a );
 a19329a <=( (not A233)  and  A232 );
 a19330a <=( A203  and  a19329a );
 a19333a <=( A236  and  (not A235) );
 a19336a <=( A267  and  A265 );
 a19337a <=( a19336a  and  a19333a );
 a19338a <=( a19337a  and  a19330a );
 a19342a <=( (not A167)  and  A168 );
 a19343a <=( A169  and  a19342a );
 a19347a <=( (not A200)  and  (not A199) );
 a19348a <=( A166  and  a19347a );
 a19349a <=( a19348a  and  a19343a );
 a19353a <=( (not A233)  and  A232 );
 a19354a <=( A203  and  a19353a );
 a19357a <=( A236  and  (not A235) );
 a19360a <=( A267  and  A266 );
 a19361a <=( a19360a  and  a19357a );
 a19362a <=( a19361a  and  a19354a );
 a19366a <=( (not A167)  and  A168 );
 a19367a <=( A169  and  a19366a );
 a19371a <=( (not A200)  and  (not A199) );
 a19372a <=( A166  and  a19371a );
 a19373a <=( a19372a  and  a19367a );
 a19377a <=( (not A233)  and  (not A232) );
 a19378a <=( A203  and  a19377a );
 a19381a <=( (not A236)  and  A235 );
 a19384a <=( A300  and  A299 );
 a19385a <=( a19384a  and  a19381a );
 a19386a <=( a19385a  and  a19378a );
 a19390a <=( (not A167)  and  A168 );
 a19391a <=( A169  and  a19390a );
 a19395a <=( (not A200)  and  (not A199) );
 a19396a <=( A166  and  a19395a );
 a19397a <=( a19396a  and  a19391a );
 a19401a <=( (not A233)  and  (not A232) );
 a19402a <=( A203  and  a19401a );
 a19405a <=( (not A236)  and  A235 );
 a19408a <=( A300  and  A298 );
 a19409a <=( a19408a  and  a19405a );
 a19410a <=( a19409a  and  a19402a );
 a19414a <=( (not A167)  and  A168 );
 a19415a <=( A169  and  a19414a );
 a19419a <=( (not A200)  and  (not A199) );
 a19420a <=( A166  and  a19419a );
 a19421a <=( a19420a  and  a19415a );
 a19425a <=( (not A233)  and  (not A232) );
 a19426a <=( A203  and  a19425a );
 a19429a <=( (not A236)  and  A235 );
 a19432a <=( A267  and  A265 );
 a19433a <=( a19432a  and  a19429a );
 a19434a <=( a19433a  and  a19426a );
 a19438a <=( (not A167)  and  A168 );
 a19439a <=( A169  and  a19438a );
 a19443a <=( (not A200)  and  (not A199) );
 a19444a <=( A166  and  a19443a );
 a19445a <=( a19444a  and  a19439a );
 a19449a <=( (not A233)  and  (not A232) );
 a19450a <=( A203  and  a19449a );
 a19453a <=( (not A236)  and  A235 );
 a19456a <=( A267  and  A266 );
 a19457a <=( a19456a  and  a19453a );
 a19458a <=( a19457a  and  a19450a );
 a19462a <=( A199  and  (not A166) );
 a19463a <=( A167  and  a19462a );
 a19466a <=( (not A201)  and  A200 );
 a19469a <=( A232  and  (not A202) );
 a19470a <=( a19469a  and  a19466a );
 a19471a <=( a19470a  and  a19463a );
 a19475a <=( (not A236)  and  A235 );
 a19476a <=( A233  and  a19475a );
 a19479a <=( A299  and  A298 );
 a19482a <=( (not A302)  and  A301 );
 a19483a <=( a19482a  and  a19479a );
 a19484a <=( a19483a  and  a19476a );
 a19488a <=( A199  and  (not A166) );
 a19489a <=( A167  and  a19488a );
 a19492a <=( (not A201)  and  A200 );
 a19495a <=( A232  and  (not A202) );
 a19496a <=( a19495a  and  a19492a );
 a19497a <=( a19496a  and  a19489a );
 a19501a <=( (not A236)  and  A235 );
 a19502a <=( A233  and  a19501a );
 a19505a <=( (not A299)  and  A298 );
 a19508a <=( A302  and  (not A301) );
 a19509a <=( a19508a  and  a19505a );
 a19510a <=( a19509a  and  a19502a );
 a19514a <=( A199  and  (not A166) );
 a19515a <=( A167  and  a19514a );
 a19518a <=( (not A201)  and  A200 );
 a19521a <=( A232  and  (not A202) );
 a19522a <=( a19521a  and  a19518a );
 a19523a <=( a19522a  and  a19515a );
 a19527a <=( (not A236)  and  A235 );
 a19528a <=( A233  and  a19527a );
 a19531a <=( A299  and  (not A298) );
 a19534a <=( A302  and  (not A301) );
 a19535a <=( a19534a  and  a19531a );
 a19536a <=( a19535a  and  a19528a );
 a19540a <=( A199  and  (not A166) );
 a19541a <=( A167  and  a19540a );
 a19544a <=( (not A201)  and  A200 );
 a19547a <=( A232  and  (not A202) );
 a19548a <=( a19547a  and  a19544a );
 a19549a <=( a19548a  and  a19541a );
 a19553a <=( (not A236)  and  A235 );
 a19554a <=( A233  and  a19553a );
 a19557a <=( (not A299)  and  (not A298) );
 a19560a <=( (not A302)  and  A301 );
 a19561a <=( a19560a  and  a19557a );
 a19562a <=( a19561a  and  a19554a );
 a19566a <=( A199  and  (not A166) );
 a19567a <=( A167  and  a19566a );
 a19570a <=( (not A201)  and  A200 );
 a19573a <=( A232  and  (not A202) );
 a19574a <=( a19573a  and  a19570a );
 a19575a <=( a19574a  and  a19567a );
 a19579a <=( (not A236)  and  A235 );
 a19580a <=( A233  and  a19579a );
 a19583a <=( A266  and  A265 );
 a19586a <=( (not A269)  and  A268 );
 a19587a <=( a19586a  and  a19583a );
 a19588a <=( a19587a  and  a19580a );
 a19592a <=( A199  and  (not A166) );
 a19593a <=( A167  and  a19592a );
 a19596a <=( (not A201)  and  A200 );
 a19599a <=( A232  and  (not A202) );
 a19600a <=( a19599a  and  a19596a );
 a19601a <=( a19600a  and  a19593a );
 a19605a <=( (not A236)  and  A235 );
 a19606a <=( A233  and  a19605a );
 a19609a <=( A266  and  (not A265) );
 a19612a <=( A269  and  (not A268) );
 a19613a <=( a19612a  and  a19609a );
 a19614a <=( a19613a  and  a19606a );
 a19618a <=( A199  and  (not A166) );
 a19619a <=( A167  and  a19618a );
 a19622a <=( (not A201)  and  A200 );
 a19625a <=( A232  and  (not A202) );
 a19626a <=( a19625a  and  a19622a );
 a19627a <=( a19626a  and  a19619a );
 a19631a <=( (not A236)  and  A235 );
 a19632a <=( A233  and  a19631a );
 a19635a <=( (not A266)  and  A265 );
 a19638a <=( A269  and  (not A268) );
 a19639a <=( a19638a  and  a19635a );
 a19640a <=( a19639a  and  a19632a );
 a19644a <=( A199  and  (not A166) );
 a19645a <=( A167  and  a19644a );
 a19648a <=( (not A201)  and  A200 );
 a19651a <=( A232  and  (not A202) );
 a19652a <=( a19651a  and  a19648a );
 a19653a <=( a19652a  and  a19645a );
 a19657a <=( (not A236)  and  A235 );
 a19658a <=( A233  and  a19657a );
 a19661a <=( (not A266)  and  (not A265) );
 a19664a <=( (not A269)  and  A268 );
 a19665a <=( a19664a  and  a19661a );
 a19666a <=( a19665a  and  a19658a );
 a19670a <=( A199  and  (not A166) );
 a19671a <=( A167  and  a19670a );
 a19674a <=( (not A201)  and  A200 );
 a19677a <=( (not A232)  and  (not A202) );
 a19678a <=( a19677a  and  a19674a );
 a19679a <=( a19678a  and  a19671a );
 a19683a <=( A236  and  (not A235) );
 a19684a <=( A233  and  a19683a );
 a19687a <=( A299  and  A298 );
 a19690a <=( (not A302)  and  A301 );
 a19691a <=( a19690a  and  a19687a );
 a19692a <=( a19691a  and  a19684a );
 a19696a <=( A199  and  (not A166) );
 a19697a <=( A167  and  a19696a );
 a19700a <=( (not A201)  and  A200 );
 a19703a <=( (not A232)  and  (not A202) );
 a19704a <=( a19703a  and  a19700a );
 a19705a <=( a19704a  and  a19697a );
 a19709a <=( A236  and  (not A235) );
 a19710a <=( A233  and  a19709a );
 a19713a <=( (not A299)  and  A298 );
 a19716a <=( A302  and  (not A301) );
 a19717a <=( a19716a  and  a19713a );
 a19718a <=( a19717a  and  a19710a );
 a19722a <=( A199  and  (not A166) );
 a19723a <=( A167  and  a19722a );
 a19726a <=( (not A201)  and  A200 );
 a19729a <=( (not A232)  and  (not A202) );
 a19730a <=( a19729a  and  a19726a );
 a19731a <=( a19730a  and  a19723a );
 a19735a <=( A236  and  (not A235) );
 a19736a <=( A233  and  a19735a );
 a19739a <=( A299  and  (not A298) );
 a19742a <=( A302  and  (not A301) );
 a19743a <=( a19742a  and  a19739a );
 a19744a <=( a19743a  and  a19736a );
 a19748a <=( A199  and  (not A166) );
 a19749a <=( A167  and  a19748a );
 a19752a <=( (not A201)  and  A200 );
 a19755a <=( (not A232)  and  (not A202) );
 a19756a <=( a19755a  and  a19752a );
 a19757a <=( a19756a  and  a19749a );
 a19761a <=( A236  and  (not A235) );
 a19762a <=( A233  and  a19761a );
 a19765a <=( (not A299)  and  (not A298) );
 a19768a <=( (not A302)  and  A301 );
 a19769a <=( a19768a  and  a19765a );
 a19770a <=( a19769a  and  a19762a );
 a19774a <=( A199  and  (not A166) );
 a19775a <=( A167  and  a19774a );
 a19778a <=( (not A201)  and  A200 );
 a19781a <=( (not A232)  and  (not A202) );
 a19782a <=( a19781a  and  a19778a );
 a19783a <=( a19782a  and  a19775a );
 a19787a <=( A236  and  (not A235) );
 a19788a <=( A233  and  a19787a );
 a19791a <=( A266  and  A265 );
 a19794a <=( (not A269)  and  A268 );
 a19795a <=( a19794a  and  a19791a );
 a19796a <=( a19795a  and  a19788a );
 a19800a <=( A199  and  (not A166) );
 a19801a <=( A167  and  a19800a );
 a19804a <=( (not A201)  and  A200 );
 a19807a <=( (not A232)  and  (not A202) );
 a19808a <=( a19807a  and  a19804a );
 a19809a <=( a19808a  and  a19801a );
 a19813a <=( A236  and  (not A235) );
 a19814a <=( A233  and  a19813a );
 a19817a <=( A266  and  (not A265) );
 a19820a <=( A269  and  (not A268) );
 a19821a <=( a19820a  and  a19817a );
 a19822a <=( a19821a  and  a19814a );
 a19826a <=( A199  and  (not A166) );
 a19827a <=( A167  and  a19826a );
 a19830a <=( (not A201)  and  A200 );
 a19833a <=( (not A232)  and  (not A202) );
 a19834a <=( a19833a  and  a19830a );
 a19835a <=( a19834a  and  a19827a );
 a19839a <=( A236  and  (not A235) );
 a19840a <=( A233  and  a19839a );
 a19843a <=( (not A266)  and  A265 );
 a19846a <=( A269  and  (not A268) );
 a19847a <=( a19846a  and  a19843a );
 a19848a <=( a19847a  and  a19840a );
 a19852a <=( A199  and  (not A166) );
 a19853a <=( A167  and  a19852a );
 a19856a <=( (not A201)  and  A200 );
 a19859a <=( (not A232)  and  (not A202) );
 a19860a <=( a19859a  and  a19856a );
 a19861a <=( a19860a  and  a19853a );
 a19865a <=( A236  and  (not A235) );
 a19866a <=( A233  and  a19865a );
 a19869a <=( (not A266)  and  (not A265) );
 a19872a <=( (not A269)  and  A268 );
 a19873a <=( a19872a  and  a19869a );
 a19874a <=( a19873a  and  a19866a );
 a19878a <=( A199  and  (not A166) );
 a19879a <=( A167  and  a19878a );
 a19882a <=( (not A201)  and  A200 );
 a19885a <=( A232  and  (not A202) );
 a19886a <=( a19885a  and  a19882a );
 a19887a <=( a19886a  and  a19879a );
 a19891a <=( A236  and  (not A235) );
 a19892a <=( (not A233)  and  a19891a );
 a19895a <=( A299  and  A298 );
 a19898a <=( (not A302)  and  A301 );
 a19899a <=( a19898a  and  a19895a );
 a19900a <=( a19899a  and  a19892a );
 a19904a <=( A199  and  (not A166) );
 a19905a <=( A167  and  a19904a );
 a19908a <=( (not A201)  and  A200 );
 a19911a <=( A232  and  (not A202) );
 a19912a <=( a19911a  and  a19908a );
 a19913a <=( a19912a  and  a19905a );
 a19917a <=( A236  and  (not A235) );
 a19918a <=( (not A233)  and  a19917a );
 a19921a <=( (not A299)  and  A298 );
 a19924a <=( A302  and  (not A301) );
 a19925a <=( a19924a  and  a19921a );
 a19926a <=( a19925a  and  a19918a );
 a19930a <=( A199  and  (not A166) );
 a19931a <=( A167  and  a19930a );
 a19934a <=( (not A201)  and  A200 );
 a19937a <=( A232  and  (not A202) );
 a19938a <=( a19937a  and  a19934a );
 a19939a <=( a19938a  and  a19931a );
 a19943a <=( A236  and  (not A235) );
 a19944a <=( (not A233)  and  a19943a );
 a19947a <=( A299  and  (not A298) );
 a19950a <=( A302  and  (not A301) );
 a19951a <=( a19950a  and  a19947a );
 a19952a <=( a19951a  and  a19944a );
 a19956a <=( A199  and  (not A166) );
 a19957a <=( A167  and  a19956a );
 a19960a <=( (not A201)  and  A200 );
 a19963a <=( A232  and  (not A202) );
 a19964a <=( a19963a  and  a19960a );
 a19965a <=( a19964a  and  a19957a );
 a19969a <=( A236  and  (not A235) );
 a19970a <=( (not A233)  and  a19969a );
 a19973a <=( (not A299)  and  (not A298) );
 a19976a <=( (not A302)  and  A301 );
 a19977a <=( a19976a  and  a19973a );
 a19978a <=( a19977a  and  a19970a );
 a19982a <=( A199  and  (not A166) );
 a19983a <=( A167  and  a19982a );
 a19986a <=( (not A201)  and  A200 );
 a19989a <=( A232  and  (not A202) );
 a19990a <=( a19989a  and  a19986a );
 a19991a <=( a19990a  and  a19983a );
 a19995a <=( A236  and  (not A235) );
 a19996a <=( (not A233)  and  a19995a );
 a19999a <=( A266  and  A265 );
 a20002a <=( (not A269)  and  A268 );
 a20003a <=( a20002a  and  a19999a );
 a20004a <=( a20003a  and  a19996a );
 a20008a <=( A199  and  (not A166) );
 a20009a <=( A167  and  a20008a );
 a20012a <=( (not A201)  and  A200 );
 a20015a <=( A232  and  (not A202) );
 a20016a <=( a20015a  and  a20012a );
 a20017a <=( a20016a  and  a20009a );
 a20021a <=( A236  and  (not A235) );
 a20022a <=( (not A233)  and  a20021a );
 a20025a <=( A266  and  (not A265) );
 a20028a <=( A269  and  (not A268) );
 a20029a <=( a20028a  and  a20025a );
 a20030a <=( a20029a  and  a20022a );
 a20034a <=( A199  and  (not A166) );
 a20035a <=( A167  and  a20034a );
 a20038a <=( (not A201)  and  A200 );
 a20041a <=( A232  and  (not A202) );
 a20042a <=( a20041a  and  a20038a );
 a20043a <=( a20042a  and  a20035a );
 a20047a <=( A236  and  (not A235) );
 a20048a <=( (not A233)  and  a20047a );
 a20051a <=( (not A266)  and  A265 );
 a20054a <=( A269  and  (not A268) );
 a20055a <=( a20054a  and  a20051a );
 a20056a <=( a20055a  and  a20048a );
 a20060a <=( A199  and  (not A166) );
 a20061a <=( A167  and  a20060a );
 a20064a <=( (not A201)  and  A200 );
 a20067a <=( A232  and  (not A202) );
 a20068a <=( a20067a  and  a20064a );
 a20069a <=( a20068a  and  a20061a );
 a20073a <=( A236  and  (not A235) );
 a20074a <=( (not A233)  and  a20073a );
 a20077a <=( (not A266)  and  (not A265) );
 a20080a <=( (not A269)  and  A268 );
 a20081a <=( a20080a  and  a20077a );
 a20082a <=( a20081a  and  a20074a );
 a20086a <=( A199  and  (not A166) );
 a20087a <=( A167  and  a20086a );
 a20090a <=( (not A201)  and  A200 );
 a20093a <=( (not A232)  and  (not A202) );
 a20094a <=( a20093a  and  a20090a );
 a20095a <=( a20094a  and  a20087a );
 a20099a <=( (not A236)  and  A235 );
 a20100a <=( (not A233)  and  a20099a );
 a20103a <=( A299  and  A298 );
 a20106a <=( (not A302)  and  A301 );
 a20107a <=( a20106a  and  a20103a );
 a20108a <=( a20107a  and  a20100a );
 a20112a <=( A199  and  (not A166) );
 a20113a <=( A167  and  a20112a );
 a20116a <=( (not A201)  and  A200 );
 a20119a <=( (not A232)  and  (not A202) );
 a20120a <=( a20119a  and  a20116a );
 a20121a <=( a20120a  and  a20113a );
 a20125a <=( (not A236)  and  A235 );
 a20126a <=( (not A233)  and  a20125a );
 a20129a <=( (not A299)  and  A298 );
 a20132a <=( A302  and  (not A301) );
 a20133a <=( a20132a  and  a20129a );
 a20134a <=( a20133a  and  a20126a );
 a20138a <=( A199  and  (not A166) );
 a20139a <=( A167  and  a20138a );
 a20142a <=( (not A201)  and  A200 );
 a20145a <=( (not A232)  and  (not A202) );
 a20146a <=( a20145a  and  a20142a );
 a20147a <=( a20146a  and  a20139a );
 a20151a <=( (not A236)  and  A235 );
 a20152a <=( (not A233)  and  a20151a );
 a20155a <=( A299  and  (not A298) );
 a20158a <=( A302  and  (not A301) );
 a20159a <=( a20158a  and  a20155a );
 a20160a <=( a20159a  and  a20152a );
 a20164a <=( A199  and  (not A166) );
 a20165a <=( A167  and  a20164a );
 a20168a <=( (not A201)  and  A200 );
 a20171a <=( (not A232)  and  (not A202) );
 a20172a <=( a20171a  and  a20168a );
 a20173a <=( a20172a  and  a20165a );
 a20177a <=( (not A236)  and  A235 );
 a20178a <=( (not A233)  and  a20177a );
 a20181a <=( (not A299)  and  (not A298) );
 a20184a <=( (not A302)  and  A301 );
 a20185a <=( a20184a  and  a20181a );
 a20186a <=( a20185a  and  a20178a );
 a20190a <=( A199  and  (not A166) );
 a20191a <=( A167  and  a20190a );
 a20194a <=( (not A201)  and  A200 );
 a20197a <=( (not A232)  and  (not A202) );
 a20198a <=( a20197a  and  a20194a );
 a20199a <=( a20198a  and  a20191a );
 a20203a <=( (not A236)  and  A235 );
 a20204a <=( (not A233)  and  a20203a );
 a20207a <=( A266  and  A265 );
 a20210a <=( (not A269)  and  A268 );
 a20211a <=( a20210a  and  a20207a );
 a20212a <=( a20211a  and  a20204a );
 a20216a <=( A199  and  (not A166) );
 a20217a <=( A167  and  a20216a );
 a20220a <=( (not A201)  and  A200 );
 a20223a <=( (not A232)  and  (not A202) );
 a20224a <=( a20223a  and  a20220a );
 a20225a <=( a20224a  and  a20217a );
 a20229a <=( (not A236)  and  A235 );
 a20230a <=( (not A233)  and  a20229a );
 a20233a <=( A266  and  (not A265) );
 a20236a <=( A269  and  (not A268) );
 a20237a <=( a20236a  and  a20233a );
 a20238a <=( a20237a  and  a20230a );
 a20242a <=( A199  and  (not A166) );
 a20243a <=( A167  and  a20242a );
 a20246a <=( (not A201)  and  A200 );
 a20249a <=( (not A232)  and  (not A202) );
 a20250a <=( a20249a  and  a20246a );
 a20251a <=( a20250a  and  a20243a );
 a20255a <=( (not A236)  and  A235 );
 a20256a <=( (not A233)  and  a20255a );
 a20259a <=( (not A266)  and  A265 );
 a20262a <=( A269  and  (not A268) );
 a20263a <=( a20262a  and  a20259a );
 a20264a <=( a20263a  and  a20256a );
 a20268a <=( A199  and  (not A166) );
 a20269a <=( A167  and  a20268a );
 a20272a <=( (not A201)  and  A200 );
 a20275a <=( (not A232)  and  (not A202) );
 a20276a <=( a20275a  and  a20272a );
 a20277a <=( a20276a  and  a20269a );
 a20281a <=( (not A236)  and  A235 );
 a20282a <=( (not A233)  and  a20281a );
 a20285a <=( (not A266)  and  (not A265) );
 a20288a <=( (not A269)  and  A268 );
 a20289a <=( a20288a  and  a20285a );
 a20290a <=( a20289a  and  a20282a );
 a20294a <=( A199  and  (not A166) );
 a20295a <=( A167  and  a20294a );
 a20298a <=( (not A201)  and  A200 );
 a20301a <=( A232  and  A203 );
 a20302a <=( a20301a  and  a20298a );
 a20303a <=( a20302a  and  a20295a );
 a20307a <=( (not A236)  and  A235 );
 a20308a <=( A233  and  a20307a );
 a20311a <=( A299  and  A298 );
 a20314a <=( (not A302)  and  A301 );
 a20315a <=( a20314a  and  a20311a );
 a20316a <=( a20315a  and  a20308a );
 a20320a <=( A199  and  (not A166) );
 a20321a <=( A167  and  a20320a );
 a20324a <=( (not A201)  and  A200 );
 a20327a <=( A232  and  A203 );
 a20328a <=( a20327a  and  a20324a );
 a20329a <=( a20328a  and  a20321a );
 a20333a <=( (not A236)  and  A235 );
 a20334a <=( A233  and  a20333a );
 a20337a <=( (not A299)  and  A298 );
 a20340a <=( A302  and  (not A301) );
 a20341a <=( a20340a  and  a20337a );
 a20342a <=( a20341a  and  a20334a );
 a20346a <=( A199  and  (not A166) );
 a20347a <=( A167  and  a20346a );
 a20350a <=( (not A201)  and  A200 );
 a20353a <=( A232  and  A203 );
 a20354a <=( a20353a  and  a20350a );
 a20355a <=( a20354a  and  a20347a );
 a20359a <=( (not A236)  and  A235 );
 a20360a <=( A233  and  a20359a );
 a20363a <=( A299  and  (not A298) );
 a20366a <=( A302  and  (not A301) );
 a20367a <=( a20366a  and  a20363a );
 a20368a <=( a20367a  and  a20360a );
 a20372a <=( A199  and  (not A166) );
 a20373a <=( A167  and  a20372a );
 a20376a <=( (not A201)  and  A200 );
 a20379a <=( A232  and  A203 );
 a20380a <=( a20379a  and  a20376a );
 a20381a <=( a20380a  and  a20373a );
 a20385a <=( (not A236)  and  A235 );
 a20386a <=( A233  and  a20385a );
 a20389a <=( (not A299)  and  (not A298) );
 a20392a <=( (not A302)  and  A301 );
 a20393a <=( a20392a  and  a20389a );
 a20394a <=( a20393a  and  a20386a );
 a20398a <=( A199  and  (not A166) );
 a20399a <=( A167  and  a20398a );
 a20402a <=( (not A201)  and  A200 );
 a20405a <=( A232  and  A203 );
 a20406a <=( a20405a  and  a20402a );
 a20407a <=( a20406a  and  a20399a );
 a20411a <=( (not A236)  and  A235 );
 a20412a <=( A233  and  a20411a );
 a20415a <=( A266  and  A265 );
 a20418a <=( (not A269)  and  A268 );
 a20419a <=( a20418a  and  a20415a );
 a20420a <=( a20419a  and  a20412a );
 a20424a <=( A199  and  (not A166) );
 a20425a <=( A167  and  a20424a );
 a20428a <=( (not A201)  and  A200 );
 a20431a <=( A232  and  A203 );
 a20432a <=( a20431a  and  a20428a );
 a20433a <=( a20432a  and  a20425a );
 a20437a <=( (not A236)  and  A235 );
 a20438a <=( A233  and  a20437a );
 a20441a <=( A266  and  (not A265) );
 a20444a <=( A269  and  (not A268) );
 a20445a <=( a20444a  and  a20441a );
 a20446a <=( a20445a  and  a20438a );
 a20450a <=( A199  and  (not A166) );
 a20451a <=( A167  and  a20450a );
 a20454a <=( (not A201)  and  A200 );
 a20457a <=( A232  and  A203 );
 a20458a <=( a20457a  and  a20454a );
 a20459a <=( a20458a  and  a20451a );
 a20463a <=( (not A236)  and  A235 );
 a20464a <=( A233  and  a20463a );
 a20467a <=( (not A266)  and  A265 );
 a20470a <=( A269  and  (not A268) );
 a20471a <=( a20470a  and  a20467a );
 a20472a <=( a20471a  and  a20464a );
 a20476a <=( A199  and  (not A166) );
 a20477a <=( A167  and  a20476a );
 a20480a <=( (not A201)  and  A200 );
 a20483a <=( A232  and  A203 );
 a20484a <=( a20483a  and  a20480a );
 a20485a <=( a20484a  and  a20477a );
 a20489a <=( (not A236)  and  A235 );
 a20490a <=( A233  and  a20489a );
 a20493a <=( (not A266)  and  (not A265) );
 a20496a <=( (not A269)  and  A268 );
 a20497a <=( a20496a  and  a20493a );
 a20498a <=( a20497a  and  a20490a );
 a20502a <=( A199  and  (not A166) );
 a20503a <=( A167  and  a20502a );
 a20506a <=( (not A201)  and  A200 );
 a20509a <=( (not A232)  and  A203 );
 a20510a <=( a20509a  and  a20506a );
 a20511a <=( a20510a  and  a20503a );
 a20515a <=( A236  and  (not A235) );
 a20516a <=( A233  and  a20515a );
 a20519a <=( A299  and  A298 );
 a20522a <=( (not A302)  and  A301 );
 a20523a <=( a20522a  and  a20519a );
 a20524a <=( a20523a  and  a20516a );
 a20528a <=( A199  and  (not A166) );
 a20529a <=( A167  and  a20528a );
 a20532a <=( (not A201)  and  A200 );
 a20535a <=( (not A232)  and  A203 );
 a20536a <=( a20535a  and  a20532a );
 a20537a <=( a20536a  and  a20529a );
 a20541a <=( A236  and  (not A235) );
 a20542a <=( A233  and  a20541a );
 a20545a <=( (not A299)  and  A298 );
 a20548a <=( A302  and  (not A301) );
 a20549a <=( a20548a  and  a20545a );
 a20550a <=( a20549a  and  a20542a );
 a20554a <=( A199  and  (not A166) );
 a20555a <=( A167  and  a20554a );
 a20558a <=( (not A201)  and  A200 );
 a20561a <=( (not A232)  and  A203 );
 a20562a <=( a20561a  and  a20558a );
 a20563a <=( a20562a  and  a20555a );
 a20567a <=( A236  and  (not A235) );
 a20568a <=( A233  and  a20567a );
 a20571a <=( A299  and  (not A298) );
 a20574a <=( A302  and  (not A301) );
 a20575a <=( a20574a  and  a20571a );
 a20576a <=( a20575a  and  a20568a );
 a20580a <=( A199  and  (not A166) );
 a20581a <=( A167  and  a20580a );
 a20584a <=( (not A201)  and  A200 );
 a20587a <=( (not A232)  and  A203 );
 a20588a <=( a20587a  and  a20584a );
 a20589a <=( a20588a  and  a20581a );
 a20593a <=( A236  and  (not A235) );
 a20594a <=( A233  and  a20593a );
 a20597a <=( (not A299)  and  (not A298) );
 a20600a <=( (not A302)  and  A301 );
 a20601a <=( a20600a  and  a20597a );
 a20602a <=( a20601a  and  a20594a );
 a20606a <=( A199  and  (not A166) );
 a20607a <=( A167  and  a20606a );
 a20610a <=( (not A201)  and  A200 );
 a20613a <=( (not A232)  and  A203 );
 a20614a <=( a20613a  and  a20610a );
 a20615a <=( a20614a  and  a20607a );
 a20619a <=( A236  and  (not A235) );
 a20620a <=( A233  and  a20619a );
 a20623a <=( A266  and  A265 );
 a20626a <=( (not A269)  and  A268 );
 a20627a <=( a20626a  and  a20623a );
 a20628a <=( a20627a  and  a20620a );
 a20632a <=( A199  and  (not A166) );
 a20633a <=( A167  and  a20632a );
 a20636a <=( (not A201)  and  A200 );
 a20639a <=( (not A232)  and  A203 );
 a20640a <=( a20639a  and  a20636a );
 a20641a <=( a20640a  and  a20633a );
 a20645a <=( A236  and  (not A235) );
 a20646a <=( A233  and  a20645a );
 a20649a <=( A266  and  (not A265) );
 a20652a <=( A269  and  (not A268) );
 a20653a <=( a20652a  and  a20649a );
 a20654a <=( a20653a  and  a20646a );
 a20658a <=( A199  and  (not A166) );
 a20659a <=( A167  and  a20658a );
 a20662a <=( (not A201)  and  A200 );
 a20665a <=( (not A232)  and  A203 );
 a20666a <=( a20665a  and  a20662a );
 a20667a <=( a20666a  and  a20659a );
 a20671a <=( A236  and  (not A235) );
 a20672a <=( A233  and  a20671a );
 a20675a <=( (not A266)  and  A265 );
 a20678a <=( A269  and  (not A268) );
 a20679a <=( a20678a  and  a20675a );
 a20680a <=( a20679a  and  a20672a );
 a20684a <=( A199  and  (not A166) );
 a20685a <=( A167  and  a20684a );
 a20688a <=( (not A201)  and  A200 );
 a20691a <=( (not A232)  and  A203 );
 a20692a <=( a20691a  and  a20688a );
 a20693a <=( a20692a  and  a20685a );
 a20697a <=( A236  and  (not A235) );
 a20698a <=( A233  and  a20697a );
 a20701a <=( (not A266)  and  (not A265) );
 a20704a <=( (not A269)  and  A268 );
 a20705a <=( a20704a  and  a20701a );
 a20706a <=( a20705a  and  a20698a );
 a20710a <=( A199  and  (not A166) );
 a20711a <=( A167  and  a20710a );
 a20714a <=( (not A201)  and  A200 );
 a20717a <=( A232  and  A203 );
 a20718a <=( a20717a  and  a20714a );
 a20719a <=( a20718a  and  a20711a );
 a20723a <=( A236  and  (not A235) );
 a20724a <=( (not A233)  and  a20723a );
 a20727a <=( A299  and  A298 );
 a20730a <=( (not A302)  and  A301 );
 a20731a <=( a20730a  and  a20727a );
 a20732a <=( a20731a  and  a20724a );
 a20736a <=( A199  and  (not A166) );
 a20737a <=( A167  and  a20736a );
 a20740a <=( (not A201)  and  A200 );
 a20743a <=( A232  and  A203 );
 a20744a <=( a20743a  and  a20740a );
 a20745a <=( a20744a  and  a20737a );
 a20749a <=( A236  and  (not A235) );
 a20750a <=( (not A233)  and  a20749a );
 a20753a <=( (not A299)  and  A298 );
 a20756a <=( A302  and  (not A301) );
 a20757a <=( a20756a  and  a20753a );
 a20758a <=( a20757a  and  a20750a );
 a20762a <=( A199  and  (not A166) );
 a20763a <=( A167  and  a20762a );
 a20766a <=( (not A201)  and  A200 );
 a20769a <=( A232  and  A203 );
 a20770a <=( a20769a  and  a20766a );
 a20771a <=( a20770a  and  a20763a );
 a20775a <=( A236  and  (not A235) );
 a20776a <=( (not A233)  and  a20775a );
 a20779a <=( A299  and  (not A298) );
 a20782a <=( A302  and  (not A301) );
 a20783a <=( a20782a  and  a20779a );
 a20784a <=( a20783a  and  a20776a );
 a20788a <=( A199  and  (not A166) );
 a20789a <=( A167  and  a20788a );
 a20792a <=( (not A201)  and  A200 );
 a20795a <=( A232  and  A203 );
 a20796a <=( a20795a  and  a20792a );
 a20797a <=( a20796a  and  a20789a );
 a20801a <=( A236  and  (not A235) );
 a20802a <=( (not A233)  and  a20801a );
 a20805a <=( (not A299)  and  (not A298) );
 a20808a <=( (not A302)  and  A301 );
 a20809a <=( a20808a  and  a20805a );
 a20810a <=( a20809a  and  a20802a );
 a20814a <=( A199  and  (not A166) );
 a20815a <=( A167  and  a20814a );
 a20818a <=( (not A201)  and  A200 );
 a20821a <=( A232  and  A203 );
 a20822a <=( a20821a  and  a20818a );
 a20823a <=( a20822a  and  a20815a );
 a20827a <=( A236  and  (not A235) );
 a20828a <=( (not A233)  and  a20827a );
 a20831a <=( A266  and  A265 );
 a20834a <=( (not A269)  and  A268 );
 a20835a <=( a20834a  and  a20831a );
 a20836a <=( a20835a  and  a20828a );
 a20840a <=( A199  and  (not A166) );
 a20841a <=( A167  and  a20840a );
 a20844a <=( (not A201)  and  A200 );
 a20847a <=( A232  and  A203 );
 a20848a <=( a20847a  and  a20844a );
 a20849a <=( a20848a  and  a20841a );
 a20853a <=( A236  and  (not A235) );
 a20854a <=( (not A233)  and  a20853a );
 a20857a <=( A266  and  (not A265) );
 a20860a <=( A269  and  (not A268) );
 a20861a <=( a20860a  and  a20857a );
 a20862a <=( a20861a  and  a20854a );
 a20866a <=( A199  and  (not A166) );
 a20867a <=( A167  and  a20866a );
 a20870a <=( (not A201)  and  A200 );
 a20873a <=( A232  and  A203 );
 a20874a <=( a20873a  and  a20870a );
 a20875a <=( a20874a  and  a20867a );
 a20879a <=( A236  and  (not A235) );
 a20880a <=( (not A233)  and  a20879a );
 a20883a <=( (not A266)  and  A265 );
 a20886a <=( A269  and  (not A268) );
 a20887a <=( a20886a  and  a20883a );
 a20888a <=( a20887a  and  a20880a );
 a20892a <=( A199  and  (not A166) );
 a20893a <=( A167  and  a20892a );
 a20896a <=( (not A201)  and  A200 );
 a20899a <=( A232  and  A203 );
 a20900a <=( a20899a  and  a20896a );
 a20901a <=( a20900a  and  a20893a );
 a20905a <=( A236  and  (not A235) );
 a20906a <=( (not A233)  and  a20905a );
 a20909a <=( (not A266)  and  (not A265) );
 a20912a <=( (not A269)  and  A268 );
 a20913a <=( a20912a  and  a20909a );
 a20914a <=( a20913a  and  a20906a );
 a20918a <=( A199  and  (not A166) );
 a20919a <=( A167  and  a20918a );
 a20922a <=( (not A201)  and  A200 );
 a20925a <=( (not A232)  and  A203 );
 a20926a <=( a20925a  and  a20922a );
 a20927a <=( a20926a  and  a20919a );
 a20931a <=( (not A236)  and  A235 );
 a20932a <=( (not A233)  and  a20931a );
 a20935a <=( A299  and  A298 );
 a20938a <=( (not A302)  and  A301 );
 a20939a <=( a20938a  and  a20935a );
 a20940a <=( a20939a  and  a20932a );
 a20944a <=( A199  and  (not A166) );
 a20945a <=( A167  and  a20944a );
 a20948a <=( (not A201)  and  A200 );
 a20951a <=( (not A232)  and  A203 );
 a20952a <=( a20951a  and  a20948a );
 a20953a <=( a20952a  and  a20945a );
 a20957a <=( (not A236)  and  A235 );
 a20958a <=( (not A233)  and  a20957a );
 a20961a <=( (not A299)  and  A298 );
 a20964a <=( A302  and  (not A301) );
 a20965a <=( a20964a  and  a20961a );
 a20966a <=( a20965a  and  a20958a );
 a20970a <=( A199  and  (not A166) );
 a20971a <=( A167  and  a20970a );
 a20974a <=( (not A201)  and  A200 );
 a20977a <=( (not A232)  and  A203 );
 a20978a <=( a20977a  and  a20974a );
 a20979a <=( a20978a  and  a20971a );
 a20983a <=( (not A236)  and  A235 );
 a20984a <=( (not A233)  and  a20983a );
 a20987a <=( A299  and  (not A298) );
 a20990a <=( A302  and  (not A301) );
 a20991a <=( a20990a  and  a20987a );
 a20992a <=( a20991a  and  a20984a );
 a20996a <=( A199  and  (not A166) );
 a20997a <=( A167  and  a20996a );
 a21000a <=( (not A201)  and  A200 );
 a21003a <=( (not A232)  and  A203 );
 a21004a <=( a21003a  and  a21000a );
 a21005a <=( a21004a  and  a20997a );
 a21009a <=( (not A236)  and  A235 );
 a21010a <=( (not A233)  and  a21009a );
 a21013a <=( (not A299)  and  (not A298) );
 a21016a <=( (not A302)  and  A301 );
 a21017a <=( a21016a  and  a21013a );
 a21018a <=( a21017a  and  a21010a );
 a21022a <=( A199  and  (not A166) );
 a21023a <=( A167  and  a21022a );
 a21026a <=( (not A201)  and  A200 );
 a21029a <=( (not A232)  and  A203 );
 a21030a <=( a21029a  and  a21026a );
 a21031a <=( a21030a  and  a21023a );
 a21035a <=( (not A236)  and  A235 );
 a21036a <=( (not A233)  and  a21035a );
 a21039a <=( A266  and  A265 );
 a21042a <=( (not A269)  and  A268 );
 a21043a <=( a21042a  and  a21039a );
 a21044a <=( a21043a  and  a21036a );
 a21048a <=( A199  and  (not A166) );
 a21049a <=( A167  and  a21048a );
 a21052a <=( (not A201)  and  A200 );
 a21055a <=( (not A232)  and  A203 );
 a21056a <=( a21055a  and  a21052a );
 a21057a <=( a21056a  and  a21049a );
 a21061a <=( (not A236)  and  A235 );
 a21062a <=( (not A233)  and  a21061a );
 a21065a <=( A266  and  (not A265) );
 a21068a <=( A269  and  (not A268) );
 a21069a <=( a21068a  and  a21065a );
 a21070a <=( a21069a  and  a21062a );
 a21074a <=( A199  and  (not A166) );
 a21075a <=( A167  and  a21074a );
 a21078a <=( (not A201)  and  A200 );
 a21081a <=( (not A232)  and  A203 );
 a21082a <=( a21081a  and  a21078a );
 a21083a <=( a21082a  and  a21075a );
 a21087a <=( (not A236)  and  A235 );
 a21088a <=( (not A233)  and  a21087a );
 a21091a <=( (not A266)  and  A265 );
 a21094a <=( A269  and  (not A268) );
 a21095a <=( a21094a  and  a21091a );
 a21096a <=( a21095a  and  a21088a );
 a21100a <=( A199  and  (not A166) );
 a21101a <=( A167  and  a21100a );
 a21104a <=( (not A201)  and  A200 );
 a21107a <=( (not A232)  and  A203 );
 a21108a <=( a21107a  and  a21104a );
 a21109a <=( a21108a  and  a21101a );
 a21113a <=( (not A236)  and  A235 );
 a21114a <=( (not A233)  and  a21113a );
 a21117a <=( (not A266)  and  (not A265) );
 a21120a <=( (not A269)  and  A268 );
 a21121a <=( a21120a  and  a21117a );
 a21122a <=( a21121a  and  a21114a );
 a21126a <=( (not A199)  and  (not A166) );
 a21127a <=( A167  and  a21126a );
 a21130a <=( (not A201)  and  A200 );
 a21133a <=( A232  and  A202 );
 a21134a <=( a21133a  and  a21130a );
 a21135a <=( a21134a  and  a21127a );
 a21139a <=( (not A236)  and  A235 );
 a21140a <=( A233  and  a21139a );
 a21143a <=( A299  and  A298 );
 a21146a <=( (not A302)  and  A301 );
 a21147a <=( a21146a  and  a21143a );
 a21148a <=( a21147a  and  a21140a );
 a21152a <=( (not A199)  and  (not A166) );
 a21153a <=( A167  and  a21152a );
 a21156a <=( (not A201)  and  A200 );
 a21159a <=( A232  and  A202 );
 a21160a <=( a21159a  and  a21156a );
 a21161a <=( a21160a  and  a21153a );
 a21165a <=( (not A236)  and  A235 );
 a21166a <=( A233  and  a21165a );
 a21169a <=( (not A299)  and  A298 );
 a21172a <=( A302  and  (not A301) );
 a21173a <=( a21172a  and  a21169a );
 a21174a <=( a21173a  and  a21166a );
 a21178a <=( (not A199)  and  (not A166) );
 a21179a <=( A167  and  a21178a );
 a21182a <=( (not A201)  and  A200 );
 a21185a <=( A232  and  A202 );
 a21186a <=( a21185a  and  a21182a );
 a21187a <=( a21186a  and  a21179a );
 a21191a <=( (not A236)  and  A235 );
 a21192a <=( A233  and  a21191a );
 a21195a <=( A299  and  (not A298) );
 a21198a <=( A302  and  (not A301) );
 a21199a <=( a21198a  and  a21195a );
 a21200a <=( a21199a  and  a21192a );
 a21204a <=( (not A199)  and  (not A166) );
 a21205a <=( A167  and  a21204a );
 a21208a <=( (not A201)  and  A200 );
 a21211a <=( A232  and  A202 );
 a21212a <=( a21211a  and  a21208a );
 a21213a <=( a21212a  and  a21205a );
 a21217a <=( (not A236)  and  A235 );
 a21218a <=( A233  and  a21217a );
 a21221a <=( (not A299)  and  (not A298) );
 a21224a <=( (not A302)  and  A301 );
 a21225a <=( a21224a  and  a21221a );
 a21226a <=( a21225a  and  a21218a );
 a21230a <=( (not A199)  and  (not A166) );
 a21231a <=( A167  and  a21230a );
 a21234a <=( (not A201)  and  A200 );
 a21237a <=( A232  and  A202 );
 a21238a <=( a21237a  and  a21234a );
 a21239a <=( a21238a  and  a21231a );
 a21243a <=( (not A236)  and  A235 );
 a21244a <=( A233  and  a21243a );
 a21247a <=( A266  and  A265 );
 a21250a <=( (not A269)  and  A268 );
 a21251a <=( a21250a  and  a21247a );
 a21252a <=( a21251a  and  a21244a );
 a21256a <=( (not A199)  and  (not A166) );
 a21257a <=( A167  and  a21256a );
 a21260a <=( (not A201)  and  A200 );
 a21263a <=( A232  and  A202 );
 a21264a <=( a21263a  and  a21260a );
 a21265a <=( a21264a  and  a21257a );
 a21269a <=( (not A236)  and  A235 );
 a21270a <=( A233  and  a21269a );
 a21273a <=( A266  and  (not A265) );
 a21276a <=( A269  and  (not A268) );
 a21277a <=( a21276a  and  a21273a );
 a21278a <=( a21277a  and  a21270a );
 a21282a <=( (not A199)  and  (not A166) );
 a21283a <=( A167  and  a21282a );
 a21286a <=( (not A201)  and  A200 );
 a21289a <=( A232  and  A202 );
 a21290a <=( a21289a  and  a21286a );
 a21291a <=( a21290a  and  a21283a );
 a21295a <=( (not A236)  and  A235 );
 a21296a <=( A233  and  a21295a );
 a21299a <=( (not A266)  and  A265 );
 a21302a <=( A269  and  (not A268) );
 a21303a <=( a21302a  and  a21299a );
 a21304a <=( a21303a  and  a21296a );
 a21308a <=( (not A199)  and  (not A166) );
 a21309a <=( A167  and  a21308a );
 a21312a <=( (not A201)  and  A200 );
 a21315a <=( A232  and  A202 );
 a21316a <=( a21315a  and  a21312a );
 a21317a <=( a21316a  and  a21309a );
 a21321a <=( (not A236)  and  A235 );
 a21322a <=( A233  and  a21321a );
 a21325a <=( (not A266)  and  (not A265) );
 a21328a <=( (not A269)  and  A268 );
 a21329a <=( a21328a  and  a21325a );
 a21330a <=( a21329a  and  a21322a );
 a21334a <=( (not A199)  and  (not A166) );
 a21335a <=( A167  and  a21334a );
 a21338a <=( (not A201)  and  A200 );
 a21341a <=( (not A232)  and  A202 );
 a21342a <=( a21341a  and  a21338a );
 a21343a <=( a21342a  and  a21335a );
 a21347a <=( A236  and  (not A235) );
 a21348a <=( A233  and  a21347a );
 a21351a <=( A299  and  A298 );
 a21354a <=( (not A302)  and  A301 );
 a21355a <=( a21354a  and  a21351a );
 a21356a <=( a21355a  and  a21348a );
 a21360a <=( (not A199)  and  (not A166) );
 a21361a <=( A167  and  a21360a );
 a21364a <=( (not A201)  and  A200 );
 a21367a <=( (not A232)  and  A202 );
 a21368a <=( a21367a  and  a21364a );
 a21369a <=( a21368a  and  a21361a );
 a21373a <=( A236  and  (not A235) );
 a21374a <=( A233  and  a21373a );
 a21377a <=( (not A299)  and  A298 );
 a21380a <=( A302  and  (not A301) );
 a21381a <=( a21380a  and  a21377a );
 a21382a <=( a21381a  and  a21374a );
 a21386a <=( (not A199)  and  (not A166) );
 a21387a <=( A167  and  a21386a );
 a21390a <=( (not A201)  and  A200 );
 a21393a <=( (not A232)  and  A202 );
 a21394a <=( a21393a  and  a21390a );
 a21395a <=( a21394a  and  a21387a );
 a21399a <=( A236  and  (not A235) );
 a21400a <=( A233  and  a21399a );
 a21403a <=( A299  and  (not A298) );
 a21406a <=( A302  and  (not A301) );
 a21407a <=( a21406a  and  a21403a );
 a21408a <=( a21407a  and  a21400a );
 a21412a <=( (not A199)  and  (not A166) );
 a21413a <=( A167  and  a21412a );
 a21416a <=( (not A201)  and  A200 );
 a21419a <=( (not A232)  and  A202 );
 a21420a <=( a21419a  and  a21416a );
 a21421a <=( a21420a  and  a21413a );
 a21425a <=( A236  and  (not A235) );
 a21426a <=( A233  and  a21425a );
 a21429a <=( (not A299)  and  (not A298) );
 a21432a <=( (not A302)  and  A301 );
 a21433a <=( a21432a  and  a21429a );
 a21434a <=( a21433a  and  a21426a );
 a21438a <=( (not A199)  and  (not A166) );
 a21439a <=( A167  and  a21438a );
 a21442a <=( (not A201)  and  A200 );
 a21445a <=( (not A232)  and  A202 );
 a21446a <=( a21445a  and  a21442a );
 a21447a <=( a21446a  and  a21439a );
 a21451a <=( A236  and  (not A235) );
 a21452a <=( A233  and  a21451a );
 a21455a <=( A266  and  A265 );
 a21458a <=( (not A269)  and  A268 );
 a21459a <=( a21458a  and  a21455a );
 a21460a <=( a21459a  and  a21452a );
 a21464a <=( (not A199)  and  (not A166) );
 a21465a <=( A167  and  a21464a );
 a21468a <=( (not A201)  and  A200 );
 a21471a <=( (not A232)  and  A202 );
 a21472a <=( a21471a  and  a21468a );
 a21473a <=( a21472a  and  a21465a );
 a21477a <=( A236  and  (not A235) );
 a21478a <=( A233  and  a21477a );
 a21481a <=( A266  and  (not A265) );
 a21484a <=( A269  and  (not A268) );
 a21485a <=( a21484a  and  a21481a );
 a21486a <=( a21485a  and  a21478a );
 a21490a <=( (not A199)  and  (not A166) );
 a21491a <=( A167  and  a21490a );
 a21494a <=( (not A201)  and  A200 );
 a21497a <=( (not A232)  and  A202 );
 a21498a <=( a21497a  and  a21494a );
 a21499a <=( a21498a  and  a21491a );
 a21503a <=( A236  and  (not A235) );
 a21504a <=( A233  and  a21503a );
 a21507a <=( (not A266)  and  A265 );
 a21510a <=( A269  and  (not A268) );
 a21511a <=( a21510a  and  a21507a );
 a21512a <=( a21511a  and  a21504a );
 a21516a <=( (not A199)  and  (not A166) );
 a21517a <=( A167  and  a21516a );
 a21520a <=( (not A201)  and  A200 );
 a21523a <=( (not A232)  and  A202 );
 a21524a <=( a21523a  and  a21520a );
 a21525a <=( a21524a  and  a21517a );
 a21529a <=( A236  and  (not A235) );
 a21530a <=( A233  and  a21529a );
 a21533a <=( (not A266)  and  (not A265) );
 a21536a <=( (not A269)  and  A268 );
 a21537a <=( a21536a  and  a21533a );
 a21538a <=( a21537a  and  a21530a );
 a21542a <=( (not A199)  and  (not A166) );
 a21543a <=( A167  and  a21542a );
 a21546a <=( (not A201)  and  A200 );
 a21549a <=( A232  and  A202 );
 a21550a <=( a21549a  and  a21546a );
 a21551a <=( a21550a  and  a21543a );
 a21555a <=( A236  and  (not A235) );
 a21556a <=( (not A233)  and  a21555a );
 a21559a <=( A299  and  A298 );
 a21562a <=( (not A302)  and  A301 );
 a21563a <=( a21562a  and  a21559a );
 a21564a <=( a21563a  and  a21556a );
 a21568a <=( (not A199)  and  (not A166) );
 a21569a <=( A167  and  a21568a );
 a21572a <=( (not A201)  and  A200 );
 a21575a <=( A232  and  A202 );
 a21576a <=( a21575a  and  a21572a );
 a21577a <=( a21576a  and  a21569a );
 a21581a <=( A236  and  (not A235) );
 a21582a <=( (not A233)  and  a21581a );
 a21585a <=( (not A299)  and  A298 );
 a21588a <=( A302  and  (not A301) );
 a21589a <=( a21588a  and  a21585a );
 a21590a <=( a21589a  and  a21582a );
 a21594a <=( (not A199)  and  (not A166) );
 a21595a <=( A167  and  a21594a );
 a21598a <=( (not A201)  and  A200 );
 a21601a <=( A232  and  A202 );
 a21602a <=( a21601a  and  a21598a );
 a21603a <=( a21602a  and  a21595a );
 a21607a <=( A236  and  (not A235) );
 a21608a <=( (not A233)  and  a21607a );
 a21611a <=( A299  and  (not A298) );
 a21614a <=( A302  and  (not A301) );
 a21615a <=( a21614a  and  a21611a );
 a21616a <=( a21615a  and  a21608a );
 a21620a <=( (not A199)  and  (not A166) );
 a21621a <=( A167  and  a21620a );
 a21624a <=( (not A201)  and  A200 );
 a21627a <=( A232  and  A202 );
 a21628a <=( a21627a  and  a21624a );
 a21629a <=( a21628a  and  a21621a );
 a21633a <=( A236  and  (not A235) );
 a21634a <=( (not A233)  and  a21633a );
 a21637a <=( (not A299)  and  (not A298) );
 a21640a <=( (not A302)  and  A301 );
 a21641a <=( a21640a  and  a21637a );
 a21642a <=( a21641a  and  a21634a );
 a21646a <=( (not A199)  and  (not A166) );
 a21647a <=( A167  and  a21646a );
 a21650a <=( (not A201)  and  A200 );
 a21653a <=( A232  and  A202 );
 a21654a <=( a21653a  and  a21650a );
 a21655a <=( a21654a  and  a21647a );
 a21659a <=( A236  and  (not A235) );
 a21660a <=( (not A233)  and  a21659a );
 a21663a <=( A266  and  A265 );
 a21666a <=( (not A269)  and  A268 );
 a21667a <=( a21666a  and  a21663a );
 a21668a <=( a21667a  and  a21660a );
 a21672a <=( (not A199)  and  (not A166) );
 a21673a <=( A167  and  a21672a );
 a21676a <=( (not A201)  and  A200 );
 a21679a <=( A232  and  A202 );
 a21680a <=( a21679a  and  a21676a );
 a21681a <=( a21680a  and  a21673a );
 a21685a <=( A236  and  (not A235) );
 a21686a <=( (not A233)  and  a21685a );
 a21689a <=( A266  and  (not A265) );
 a21692a <=( A269  and  (not A268) );
 a21693a <=( a21692a  and  a21689a );
 a21694a <=( a21693a  and  a21686a );
 a21698a <=( (not A199)  and  (not A166) );
 a21699a <=( A167  and  a21698a );
 a21702a <=( (not A201)  and  A200 );
 a21705a <=( A232  and  A202 );
 a21706a <=( a21705a  and  a21702a );
 a21707a <=( a21706a  and  a21699a );
 a21711a <=( A236  and  (not A235) );
 a21712a <=( (not A233)  and  a21711a );
 a21715a <=( (not A266)  and  A265 );
 a21718a <=( A269  and  (not A268) );
 a21719a <=( a21718a  and  a21715a );
 a21720a <=( a21719a  and  a21712a );
 a21724a <=( (not A199)  and  (not A166) );
 a21725a <=( A167  and  a21724a );
 a21728a <=( (not A201)  and  A200 );
 a21731a <=( A232  and  A202 );
 a21732a <=( a21731a  and  a21728a );
 a21733a <=( a21732a  and  a21725a );
 a21737a <=( A236  and  (not A235) );
 a21738a <=( (not A233)  and  a21737a );
 a21741a <=( (not A266)  and  (not A265) );
 a21744a <=( (not A269)  and  A268 );
 a21745a <=( a21744a  and  a21741a );
 a21746a <=( a21745a  and  a21738a );
 a21750a <=( (not A199)  and  (not A166) );
 a21751a <=( A167  and  a21750a );
 a21754a <=( (not A201)  and  A200 );
 a21757a <=( (not A232)  and  A202 );
 a21758a <=( a21757a  and  a21754a );
 a21759a <=( a21758a  and  a21751a );
 a21763a <=( (not A236)  and  A235 );
 a21764a <=( (not A233)  and  a21763a );
 a21767a <=( A299  and  A298 );
 a21770a <=( (not A302)  and  A301 );
 a21771a <=( a21770a  and  a21767a );
 a21772a <=( a21771a  and  a21764a );
 a21776a <=( (not A199)  and  (not A166) );
 a21777a <=( A167  and  a21776a );
 a21780a <=( (not A201)  and  A200 );
 a21783a <=( (not A232)  and  A202 );
 a21784a <=( a21783a  and  a21780a );
 a21785a <=( a21784a  and  a21777a );
 a21789a <=( (not A236)  and  A235 );
 a21790a <=( (not A233)  and  a21789a );
 a21793a <=( (not A299)  and  A298 );
 a21796a <=( A302  and  (not A301) );
 a21797a <=( a21796a  and  a21793a );
 a21798a <=( a21797a  and  a21790a );
 a21802a <=( (not A199)  and  (not A166) );
 a21803a <=( A167  and  a21802a );
 a21806a <=( (not A201)  and  A200 );
 a21809a <=( (not A232)  and  A202 );
 a21810a <=( a21809a  and  a21806a );
 a21811a <=( a21810a  and  a21803a );
 a21815a <=( (not A236)  and  A235 );
 a21816a <=( (not A233)  and  a21815a );
 a21819a <=( A299  and  (not A298) );
 a21822a <=( A302  and  (not A301) );
 a21823a <=( a21822a  and  a21819a );
 a21824a <=( a21823a  and  a21816a );
 a21828a <=( (not A199)  and  (not A166) );
 a21829a <=( A167  and  a21828a );
 a21832a <=( (not A201)  and  A200 );
 a21835a <=( (not A232)  and  A202 );
 a21836a <=( a21835a  and  a21832a );
 a21837a <=( a21836a  and  a21829a );
 a21841a <=( (not A236)  and  A235 );
 a21842a <=( (not A233)  and  a21841a );
 a21845a <=( (not A299)  and  (not A298) );
 a21848a <=( (not A302)  and  A301 );
 a21849a <=( a21848a  and  a21845a );
 a21850a <=( a21849a  and  a21842a );
 a21854a <=( (not A199)  and  (not A166) );
 a21855a <=( A167  and  a21854a );
 a21858a <=( (not A201)  and  A200 );
 a21861a <=( (not A232)  and  A202 );
 a21862a <=( a21861a  and  a21858a );
 a21863a <=( a21862a  and  a21855a );
 a21867a <=( (not A236)  and  A235 );
 a21868a <=( (not A233)  and  a21867a );
 a21871a <=( A266  and  A265 );
 a21874a <=( (not A269)  and  A268 );
 a21875a <=( a21874a  and  a21871a );
 a21876a <=( a21875a  and  a21868a );
 a21880a <=( (not A199)  and  (not A166) );
 a21881a <=( A167  and  a21880a );
 a21884a <=( (not A201)  and  A200 );
 a21887a <=( (not A232)  and  A202 );
 a21888a <=( a21887a  and  a21884a );
 a21889a <=( a21888a  and  a21881a );
 a21893a <=( (not A236)  and  A235 );
 a21894a <=( (not A233)  and  a21893a );
 a21897a <=( A266  and  (not A265) );
 a21900a <=( A269  and  (not A268) );
 a21901a <=( a21900a  and  a21897a );
 a21902a <=( a21901a  and  a21894a );
 a21906a <=( (not A199)  and  (not A166) );
 a21907a <=( A167  and  a21906a );
 a21910a <=( (not A201)  and  A200 );
 a21913a <=( (not A232)  and  A202 );
 a21914a <=( a21913a  and  a21910a );
 a21915a <=( a21914a  and  a21907a );
 a21919a <=( (not A236)  and  A235 );
 a21920a <=( (not A233)  and  a21919a );
 a21923a <=( (not A266)  and  A265 );
 a21926a <=( A269  and  (not A268) );
 a21927a <=( a21926a  and  a21923a );
 a21928a <=( a21927a  and  a21920a );
 a21932a <=( (not A199)  and  (not A166) );
 a21933a <=( A167  and  a21932a );
 a21936a <=( (not A201)  and  A200 );
 a21939a <=( (not A232)  and  A202 );
 a21940a <=( a21939a  and  a21936a );
 a21941a <=( a21940a  and  a21933a );
 a21945a <=( (not A236)  and  A235 );
 a21946a <=( (not A233)  and  a21945a );
 a21949a <=( (not A266)  and  (not A265) );
 a21952a <=( (not A269)  and  A268 );
 a21953a <=( a21952a  and  a21949a );
 a21954a <=( a21953a  and  a21946a );
 a21958a <=( (not A199)  and  (not A166) );
 a21959a <=( A167  and  a21958a );
 a21962a <=( (not A201)  and  A200 );
 a21965a <=( A232  and  (not A203) );
 a21966a <=( a21965a  and  a21962a );
 a21967a <=( a21966a  and  a21959a );
 a21971a <=( (not A236)  and  A235 );
 a21972a <=( A233  and  a21971a );
 a21975a <=( A299  and  A298 );
 a21978a <=( (not A302)  and  A301 );
 a21979a <=( a21978a  and  a21975a );
 a21980a <=( a21979a  and  a21972a );
 a21984a <=( (not A199)  and  (not A166) );
 a21985a <=( A167  and  a21984a );
 a21988a <=( (not A201)  and  A200 );
 a21991a <=( A232  and  (not A203) );
 a21992a <=( a21991a  and  a21988a );
 a21993a <=( a21992a  and  a21985a );
 a21997a <=( (not A236)  and  A235 );
 a21998a <=( A233  and  a21997a );
 a22001a <=( (not A299)  and  A298 );
 a22004a <=( A302  and  (not A301) );
 a22005a <=( a22004a  and  a22001a );
 a22006a <=( a22005a  and  a21998a );
 a22010a <=( (not A199)  and  (not A166) );
 a22011a <=( A167  and  a22010a );
 a22014a <=( (not A201)  and  A200 );
 a22017a <=( A232  and  (not A203) );
 a22018a <=( a22017a  and  a22014a );
 a22019a <=( a22018a  and  a22011a );
 a22023a <=( (not A236)  and  A235 );
 a22024a <=( A233  and  a22023a );
 a22027a <=( A299  and  (not A298) );
 a22030a <=( A302  and  (not A301) );
 a22031a <=( a22030a  and  a22027a );
 a22032a <=( a22031a  and  a22024a );
 a22036a <=( (not A199)  and  (not A166) );
 a22037a <=( A167  and  a22036a );
 a22040a <=( (not A201)  and  A200 );
 a22043a <=( A232  and  (not A203) );
 a22044a <=( a22043a  and  a22040a );
 a22045a <=( a22044a  and  a22037a );
 a22049a <=( (not A236)  and  A235 );
 a22050a <=( A233  and  a22049a );
 a22053a <=( (not A299)  and  (not A298) );
 a22056a <=( (not A302)  and  A301 );
 a22057a <=( a22056a  and  a22053a );
 a22058a <=( a22057a  and  a22050a );
 a22062a <=( (not A199)  and  (not A166) );
 a22063a <=( A167  and  a22062a );
 a22066a <=( (not A201)  and  A200 );
 a22069a <=( A232  and  (not A203) );
 a22070a <=( a22069a  and  a22066a );
 a22071a <=( a22070a  and  a22063a );
 a22075a <=( (not A236)  and  A235 );
 a22076a <=( A233  and  a22075a );
 a22079a <=( A266  and  A265 );
 a22082a <=( (not A269)  and  A268 );
 a22083a <=( a22082a  and  a22079a );
 a22084a <=( a22083a  and  a22076a );
 a22088a <=( (not A199)  and  (not A166) );
 a22089a <=( A167  and  a22088a );
 a22092a <=( (not A201)  and  A200 );
 a22095a <=( A232  and  (not A203) );
 a22096a <=( a22095a  and  a22092a );
 a22097a <=( a22096a  and  a22089a );
 a22101a <=( (not A236)  and  A235 );
 a22102a <=( A233  and  a22101a );
 a22105a <=( A266  and  (not A265) );
 a22108a <=( A269  and  (not A268) );
 a22109a <=( a22108a  and  a22105a );
 a22110a <=( a22109a  and  a22102a );
 a22114a <=( (not A199)  and  (not A166) );
 a22115a <=( A167  and  a22114a );
 a22118a <=( (not A201)  and  A200 );
 a22121a <=( A232  and  (not A203) );
 a22122a <=( a22121a  and  a22118a );
 a22123a <=( a22122a  and  a22115a );
 a22127a <=( (not A236)  and  A235 );
 a22128a <=( A233  and  a22127a );
 a22131a <=( (not A266)  and  A265 );
 a22134a <=( A269  and  (not A268) );
 a22135a <=( a22134a  and  a22131a );
 a22136a <=( a22135a  and  a22128a );
 a22140a <=( (not A199)  and  (not A166) );
 a22141a <=( A167  and  a22140a );
 a22144a <=( (not A201)  and  A200 );
 a22147a <=( A232  and  (not A203) );
 a22148a <=( a22147a  and  a22144a );
 a22149a <=( a22148a  and  a22141a );
 a22153a <=( (not A236)  and  A235 );
 a22154a <=( A233  and  a22153a );
 a22157a <=( (not A266)  and  (not A265) );
 a22160a <=( (not A269)  and  A268 );
 a22161a <=( a22160a  and  a22157a );
 a22162a <=( a22161a  and  a22154a );
 a22166a <=( (not A199)  and  (not A166) );
 a22167a <=( A167  and  a22166a );
 a22170a <=( (not A201)  and  A200 );
 a22173a <=( (not A232)  and  (not A203) );
 a22174a <=( a22173a  and  a22170a );
 a22175a <=( a22174a  and  a22167a );
 a22179a <=( A236  and  (not A235) );
 a22180a <=( A233  and  a22179a );
 a22183a <=( A299  and  A298 );
 a22186a <=( (not A302)  and  A301 );
 a22187a <=( a22186a  and  a22183a );
 a22188a <=( a22187a  and  a22180a );
 a22192a <=( (not A199)  and  (not A166) );
 a22193a <=( A167  and  a22192a );
 a22196a <=( (not A201)  and  A200 );
 a22199a <=( (not A232)  and  (not A203) );
 a22200a <=( a22199a  and  a22196a );
 a22201a <=( a22200a  and  a22193a );
 a22205a <=( A236  and  (not A235) );
 a22206a <=( A233  and  a22205a );
 a22209a <=( (not A299)  and  A298 );
 a22212a <=( A302  and  (not A301) );
 a22213a <=( a22212a  and  a22209a );
 a22214a <=( a22213a  and  a22206a );
 a22218a <=( (not A199)  and  (not A166) );
 a22219a <=( A167  and  a22218a );
 a22222a <=( (not A201)  and  A200 );
 a22225a <=( (not A232)  and  (not A203) );
 a22226a <=( a22225a  and  a22222a );
 a22227a <=( a22226a  and  a22219a );
 a22231a <=( A236  and  (not A235) );
 a22232a <=( A233  and  a22231a );
 a22235a <=( A299  and  (not A298) );
 a22238a <=( A302  and  (not A301) );
 a22239a <=( a22238a  and  a22235a );
 a22240a <=( a22239a  and  a22232a );
 a22244a <=( (not A199)  and  (not A166) );
 a22245a <=( A167  and  a22244a );
 a22248a <=( (not A201)  and  A200 );
 a22251a <=( (not A232)  and  (not A203) );
 a22252a <=( a22251a  and  a22248a );
 a22253a <=( a22252a  and  a22245a );
 a22257a <=( A236  and  (not A235) );
 a22258a <=( A233  and  a22257a );
 a22261a <=( (not A299)  and  (not A298) );
 a22264a <=( (not A302)  and  A301 );
 a22265a <=( a22264a  and  a22261a );
 a22266a <=( a22265a  and  a22258a );
 a22270a <=( (not A199)  and  (not A166) );
 a22271a <=( A167  and  a22270a );
 a22274a <=( (not A201)  and  A200 );
 a22277a <=( (not A232)  and  (not A203) );
 a22278a <=( a22277a  and  a22274a );
 a22279a <=( a22278a  and  a22271a );
 a22283a <=( A236  and  (not A235) );
 a22284a <=( A233  and  a22283a );
 a22287a <=( A266  and  A265 );
 a22290a <=( (not A269)  and  A268 );
 a22291a <=( a22290a  and  a22287a );
 a22292a <=( a22291a  and  a22284a );
 a22296a <=( (not A199)  and  (not A166) );
 a22297a <=( A167  and  a22296a );
 a22300a <=( (not A201)  and  A200 );
 a22303a <=( (not A232)  and  (not A203) );
 a22304a <=( a22303a  and  a22300a );
 a22305a <=( a22304a  and  a22297a );
 a22309a <=( A236  and  (not A235) );
 a22310a <=( A233  and  a22309a );
 a22313a <=( A266  and  (not A265) );
 a22316a <=( A269  and  (not A268) );
 a22317a <=( a22316a  and  a22313a );
 a22318a <=( a22317a  and  a22310a );
 a22322a <=( (not A199)  and  (not A166) );
 a22323a <=( A167  and  a22322a );
 a22326a <=( (not A201)  and  A200 );
 a22329a <=( (not A232)  and  (not A203) );
 a22330a <=( a22329a  and  a22326a );
 a22331a <=( a22330a  and  a22323a );
 a22335a <=( A236  and  (not A235) );
 a22336a <=( A233  and  a22335a );
 a22339a <=( (not A266)  and  A265 );
 a22342a <=( A269  and  (not A268) );
 a22343a <=( a22342a  and  a22339a );
 a22344a <=( a22343a  and  a22336a );
 a22348a <=( (not A199)  and  (not A166) );
 a22349a <=( A167  and  a22348a );
 a22352a <=( (not A201)  and  A200 );
 a22355a <=( (not A232)  and  (not A203) );
 a22356a <=( a22355a  and  a22352a );
 a22357a <=( a22356a  and  a22349a );
 a22361a <=( A236  and  (not A235) );
 a22362a <=( A233  and  a22361a );
 a22365a <=( (not A266)  and  (not A265) );
 a22368a <=( (not A269)  and  A268 );
 a22369a <=( a22368a  and  a22365a );
 a22370a <=( a22369a  and  a22362a );
 a22374a <=( (not A199)  and  (not A166) );
 a22375a <=( A167  and  a22374a );
 a22378a <=( (not A201)  and  A200 );
 a22381a <=( A232  and  (not A203) );
 a22382a <=( a22381a  and  a22378a );
 a22383a <=( a22382a  and  a22375a );
 a22387a <=( A236  and  (not A235) );
 a22388a <=( (not A233)  and  a22387a );
 a22391a <=( A299  and  A298 );
 a22394a <=( (not A302)  and  A301 );
 a22395a <=( a22394a  and  a22391a );
 a22396a <=( a22395a  and  a22388a );
 a22400a <=( (not A199)  and  (not A166) );
 a22401a <=( A167  and  a22400a );
 a22404a <=( (not A201)  and  A200 );
 a22407a <=( A232  and  (not A203) );
 a22408a <=( a22407a  and  a22404a );
 a22409a <=( a22408a  and  a22401a );
 a22413a <=( A236  and  (not A235) );
 a22414a <=( (not A233)  and  a22413a );
 a22417a <=( (not A299)  and  A298 );
 a22420a <=( A302  and  (not A301) );
 a22421a <=( a22420a  and  a22417a );
 a22422a <=( a22421a  and  a22414a );
 a22426a <=( (not A199)  and  (not A166) );
 a22427a <=( A167  and  a22426a );
 a22430a <=( (not A201)  and  A200 );
 a22433a <=( A232  and  (not A203) );
 a22434a <=( a22433a  and  a22430a );
 a22435a <=( a22434a  and  a22427a );
 a22439a <=( A236  and  (not A235) );
 a22440a <=( (not A233)  and  a22439a );
 a22443a <=( A299  and  (not A298) );
 a22446a <=( A302  and  (not A301) );
 a22447a <=( a22446a  and  a22443a );
 a22448a <=( a22447a  and  a22440a );
 a22452a <=( (not A199)  and  (not A166) );
 a22453a <=( A167  and  a22452a );
 a22456a <=( (not A201)  and  A200 );
 a22459a <=( A232  and  (not A203) );
 a22460a <=( a22459a  and  a22456a );
 a22461a <=( a22460a  and  a22453a );
 a22465a <=( A236  and  (not A235) );
 a22466a <=( (not A233)  and  a22465a );
 a22469a <=( (not A299)  and  (not A298) );
 a22472a <=( (not A302)  and  A301 );
 a22473a <=( a22472a  and  a22469a );
 a22474a <=( a22473a  and  a22466a );
 a22478a <=( (not A199)  and  (not A166) );
 a22479a <=( A167  and  a22478a );
 a22482a <=( (not A201)  and  A200 );
 a22485a <=( A232  and  (not A203) );
 a22486a <=( a22485a  and  a22482a );
 a22487a <=( a22486a  and  a22479a );
 a22491a <=( A236  and  (not A235) );
 a22492a <=( (not A233)  and  a22491a );
 a22495a <=( A266  and  A265 );
 a22498a <=( (not A269)  and  A268 );
 a22499a <=( a22498a  and  a22495a );
 a22500a <=( a22499a  and  a22492a );
 a22504a <=( (not A199)  and  (not A166) );
 a22505a <=( A167  and  a22504a );
 a22508a <=( (not A201)  and  A200 );
 a22511a <=( A232  and  (not A203) );
 a22512a <=( a22511a  and  a22508a );
 a22513a <=( a22512a  and  a22505a );
 a22517a <=( A236  and  (not A235) );
 a22518a <=( (not A233)  and  a22517a );
 a22521a <=( A266  and  (not A265) );
 a22524a <=( A269  and  (not A268) );
 a22525a <=( a22524a  and  a22521a );
 a22526a <=( a22525a  and  a22518a );
 a22530a <=( (not A199)  and  (not A166) );
 a22531a <=( A167  and  a22530a );
 a22534a <=( (not A201)  and  A200 );
 a22537a <=( A232  and  (not A203) );
 a22538a <=( a22537a  and  a22534a );
 a22539a <=( a22538a  and  a22531a );
 a22543a <=( A236  and  (not A235) );
 a22544a <=( (not A233)  and  a22543a );
 a22547a <=( (not A266)  and  A265 );
 a22550a <=( A269  and  (not A268) );
 a22551a <=( a22550a  and  a22547a );
 a22552a <=( a22551a  and  a22544a );
 a22556a <=( (not A199)  and  (not A166) );
 a22557a <=( A167  and  a22556a );
 a22560a <=( (not A201)  and  A200 );
 a22563a <=( A232  and  (not A203) );
 a22564a <=( a22563a  and  a22560a );
 a22565a <=( a22564a  and  a22557a );
 a22569a <=( A236  and  (not A235) );
 a22570a <=( (not A233)  and  a22569a );
 a22573a <=( (not A266)  and  (not A265) );
 a22576a <=( (not A269)  and  A268 );
 a22577a <=( a22576a  and  a22573a );
 a22578a <=( a22577a  and  a22570a );
 a22582a <=( (not A199)  and  (not A166) );
 a22583a <=( A167  and  a22582a );
 a22586a <=( (not A201)  and  A200 );
 a22589a <=( (not A232)  and  (not A203) );
 a22590a <=( a22589a  and  a22586a );
 a22591a <=( a22590a  and  a22583a );
 a22595a <=( (not A236)  and  A235 );
 a22596a <=( (not A233)  and  a22595a );
 a22599a <=( A299  and  A298 );
 a22602a <=( (not A302)  and  A301 );
 a22603a <=( a22602a  and  a22599a );
 a22604a <=( a22603a  and  a22596a );
 a22608a <=( (not A199)  and  (not A166) );
 a22609a <=( A167  and  a22608a );
 a22612a <=( (not A201)  and  A200 );
 a22615a <=( (not A232)  and  (not A203) );
 a22616a <=( a22615a  and  a22612a );
 a22617a <=( a22616a  and  a22609a );
 a22621a <=( (not A236)  and  A235 );
 a22622a <=( (not A233)  and  a22621a );
 a22625a <=( (not A299)  and  A298 );
 a22628a <=( A302  and  (not A301) );
 a22629a <=( a22628a  and  a22625a );
 a22630a <=( a22629a  and  a22622a );
 a22634a <=( (not A199)  and  (not A166) );
 a22635a <=( A167  and  a22634a );
 a22638a <=( (not A201)  and  A200 );
 a22641a <=( (not A232)  and  (not A203) );
 a22642a <=( a22641a  and  a22638a );
 a22643a <=( a22642a  and  a22635a );
 a22647a <=( (not A236)  and  A235 );
 a22648a <=( (not A233)  and  a22647a );
 a22651a <=( A299  and  (not A298) );
 a22654a <=( A302  and  (not A301) );
 a22655a <=( a22654a  and  a22651a );
 a22656a <=( a22655a  and  a22648a );
 a22660a <=( (not A199)  and  (not A166) );
 a22661a <=( A167  and  a22660a );
 a22664a <=( (not A201)  and  A200 );
 a22667a <=( (not A232)  and  (not A203) );
 a22668a <=( a22667a  and  a22664a );
 a22669a <=( a22668a  and  a22661a );
 a22673a <=( (not A236)  and  A235 );
 a22674a <=( (not A233)  and  a22673a );
 a22677a <=( (not A299)  and  (not A298) );
 a22680a <=( (not A302)  and  A301 );
 a22681a <=( a22680a  and  a22677a );
 a22682a <=( a22681a  and  a22674a );
 a22686a <=( (not A199)  and  (not A166) );
 a22687a <=( A167  and  a22686a );
 a22690a <=( (not A201)  and  A200 );
 a22693a <=( (not A232)  and  (not A203) );
 a22694a <=( a22693a  and  a22690a );
 a22695a <=( a22694a  and  a22687a );
 a22699a <=( (not A236)  and  A235 );
 a22700a <=( (not A233)  and  a22699a );
 a22703a <=( A266  and  A265 );
 a22706a <=( (not A269)  and  A268 );
 a22707a <=( a22706a  and  a22703a );
 a22708a <=( a22707a  and  a22700a );
 a22712a <=( (not A199)  and  (not A166) );
 a22713a <=( A167  and  a22712a );
 a22716a <=( (not A201)  and  A200 );
 a22719a <=( (not A232)  and  (not A203) );
 a22720a <=( a22719a  and  a22716a );
 a22721a <=( a22720a  and  a22713a );
 a22725a <=( (not A236)  and  A235 );
 a22726a <=( (not A233)  and  a22725a );
 a22729a <=( A266  and  (not A265) );
 a22732a <=( A269  and  (not A268) );
 a22733a <=( a22732a  and  a22729a );
 a22734a <=( a22733a  and  a22726a );
 a22738a <=( (not A199)  and  (not A166) );
 a22739a <=( A167  and  a22738a );
 a22742a <=( (not A201)  and  A200 );
 a22745a <=( (not A232)  and  (not A203) );
 a22746a <=( a22745a  and  a22742a );
 a22747a <=( a22746a  and  a22739a );
 a22751a <=( (not A236)  and  A235 );
 a22752a <=( (not A233)  and  a22751a );
 a22755a <=( (not A266)  and  A265 );
 a22758a <=( A269  and  (not A268) );
 a22759a <=( a22758a  and  a22755a );
 a22760a <=( a22759a  and  a22752a );
 a22764a <=( (not A199)  and  (not A166) );
 a22765a <=( A167  and  a22764a );
 a22768a <=( (not A201)  and  A200 );
 a22771a <=( (not A232)  and  (not A203) );
 a22772a <=( a22771a  and  a22768a );
 a22773a <=( a22772a  and  a22765a );
 a22777a <=( (not A236)  and  A235 );
 a22778a <=( (not A233)  and  a22777a );
 a22781a <=( (not A266)  and  (not A265) );
 a22784a <=( (not A269)  and  A268 );
 a22785a <=( a22784a  and  a22781a );
 a22786a <=( a22785a  and  a22778a );
 a22790a <=( A199  and  (not A166) );
 a22791a <=( A167  and  a22790a );
 a22794a <=( (not A201)  and  (not A200) );
 a22797a <=( A232  and  A202 );
 a22798a <=( a22797a  and  a22794a );
 a22799a <=( a22798a  and  a22791a );
 a22803a <=( (not A236)  and  A235 );
 a22804a <=( A233  and  a22803a );
 a22807a <=( A299  and  A298 );
 a22810a <=( (not A302)  and  A301 );
 a22811a <=( a22810a  and  a22807a );
 a22812a <=( a22811a  and  a22804a );
 a22816a <=( A199  and  (not A166) );
 a22817a <=( A167  and  a22816a );
 a22820a <=( (not A201)  and  (not A200) );
 a22823a <=( A232  and  A202 );
 a22824a <=( a22823a  and  a22820a );
 a22825a <=( a22824a  and  a22817a );
 a22829a <=( (not A236)  and  A235 );
 a22830a <=( A233  and  a22829a );
 a22833a <=( (not A299)  and  A298 );
 a22836a <=( A302  and  (not A301) );
 a22837a <=( a22836a  and  a22833a );
 a22838a <=( a22837a  and  a22830a );
 a22842a <=( A199  and  (not A166) );
 a22843a <=( A167  and  a22842a );
 a22846a <=( (not A201)  and  (not A200) );
 a22849a <=( A232  and  A202 );
 a22850a <=( a22849a  and  a22846a );
 a22851a <=( a22850a  and  a22843a );
 a22855a <=( (not A236)  and  A235 );
 a22856a <=( A233  and  a22855a );
 a22859a <=( A299  and  (not A298) );
 a22862a <=( A302  and  (not A301) );
 a22863a <=( a22862a  and  a22859a );
 a22864a <=( a22863a  and  a22856a );
 a22868a <=( A199  and  (not A166) );
 a22869a <=( A167  and  a22868a );
 a22872a <=( (not A201)  and  (not A200) );
 a22875a <=( A232  and  A202 );
 a22876a <=( a22875a  and  a22872a );
 a22877a <=( a22876a  and  a22869a );
 a22881a <=( (not A236)  and  A235 );
 a22882a <=( A233  and  a22881a );
 a22885a <=( (not A299)  and  (not A298) );
 a22888a <=( (not A302)  and  A301 );
 a22889a <=( a22888a  and  a22885a );
 a22890a <=( a22889a  and  a22882a );
 a22894a <=( A199  and  (not A166) );
 a22895a <=( A167  and  a22894a );
 a22898a <=( (not A201)  and  (not A200) );
 a22901a <=( A232  and  A202 );
 a22902a <=( a22901a  and  a22898a );
 a22903a <=( a22902a  and  a22895a );
 a22907a <=( (not A236)  and  A235 );
 a22908a <=( A233  and  a22907a );
 a22911a <=( A266  and  A265 );
 a22914a <=( (not A269)  and  A268 );
 a22915a <=( a22914a  and  a22911a );
 a22916a <=( a22915a  and  a22908a );
 a22920a <=( A199  and  (not A166) );
 a22921a <=( A167  and  a22920a );
 a22924a <=( (not A201)  and  (not A200) );
 a22927a <=( A232  and  A202 );
 a22928a <=( a22927a  and  a22924a );
 a22929a <=( a22928a  and  a22921a );
 a22933a <=( (not A236)  and  A235 );
 a22934a <=( A233  and  a22933a );
 a22937a <=( A266  and  (not A265) );
 a22940a <=( A269  and  (not A268) );
 a22941a <=( a22940a  and  a22937a );
 a22942a <=( a22941a  and  a22934a );
 a22946a <=( A199  and  (not A166) );
 a22947a <=( A167  and  a22946a );
 a22950a <=( (not A201)  and  (not A200) );
 a22953a <=( A232  and  A202 );
 a22954a <=( a22953a  and  a22950a );
 a22955a <=( a22954a  and  a22947a );
 a22959a <=( (not A236)  and  A235 );
 a22960a <=( A233  and  a22959a );
 a22963a <=( (not A266)  and  A265 );
 a22966a <=( A269  and  (not A268) );
 a22967a <=( a22966a  and  a22963a );
 a22968a <=( a22967a  and  a22960a );
 a22972a <=( A199  and  (not A166) );
 a22973a <=( A167  and  a22972a );
 a22976a <=( (not A201)  and  (not A200) );
 a22979a <=( A232  and  A202 );
 a22980a <=( a22979a  and  a22976a );
 a22981a <=( a22980a  and  a22973a );
 a22985a <=( (not A236)  and  A235 );
 a22986a <=( A233  and  a22985a );
 a22989a <=( (not A266)  and  (not A265) );
 a22992a <=( (not A269)  and  A268 );
 a22993a <=( a22992a  and  a22989a );
 a22994a <=( a22993a  and  a22986a );
 a22998a <=( A199  and  (not A166) );
 a22999a <=( A167  and  a22998a );
 a23002a <=( (not A201)  and  (not A200) );
 a23005a <=( (not A232)  and  A202 );
 a23006a <=( a23005a  and  a23002a );
 a23007a <=( a23006a  and  a22999a );
 a23011a <=( A236  and  (not A235) );
 a23012a <=( A233  and  a23011a );
 a23015a <=( A299  and  A298 );
 a23018a <=( (not A302)  and  A301 );
 a23019a <=( a23018a  and  a23015a );
 a23020a <=( a23019a  and  a23012a );
 a23024a <=( A199  and  (not A166) );
 a23025a <=( A167  and  a23024a );
 a23028a <=( (not A201)  and  (not A200) );
 a23031a <=( (not A232)  and  A202 );
 a23032a <=( a23031a  and  a23028a );
 a23033a <=( a23032a  and  a23025a );
 a23037a <=( A236  and  (not A235) );
 a23038a <=( A233  and  a23037a );
 a23041a <=( (not A299)  and  A298 );
 a23044a <=( A302  and  (not A301) );
 a23045a <=( a23044a  and  a23041a );
 a23046a <=( a23045a  and  a23038a );
 a23050a <=( A199  and  (not A166) );
 a23051a <=( A167  and  a23050a );
 a23054a <=( (not A201)  and  (not A200) );
 a23057a <=( (not A232)  and  A202 );
 a23058a <=( a23057a  and  a23054a );
 a23059a <=( a23058a  and  a23051a );
 a23063a <=( A236  and  (not A235) );
 a23064a <=( A233  and  a23063a );
 a23067a <=( A299  and  (not A298) );
 a23070a <=( A302  and  (not A301) );
 a23071a <=( a23070a  and  a23067a );
 a23072a <=( a23071a  and  a23064a );
 a23076a <=( A199  and  (not A166) );
 a23077a <=( A167  and  a23076a );
 a23080a <=( (not A201)  and  (not A200) );
 a23083a <=( (not A232)  and  A202 );
 a23084a <=( a23083a  and  a23080a );
 a23085a <=( a23084a  and  a23077a );
 a23089a <=( A236  and  (not A235) );
 a23090a <=( A233  and  a23089a );
 a23093a <=( (not A299)  and  (not A298) );
 a23096a <=( (not A302)  and  A301 );
 a23097a <=( a23096a  and  a23093a );
 a23098a <=( a23097a  and  a23090a );
 a23102a <=( A199  and  (not A166) );
 a23103a <=( A167  and  a23102a );
 a23106a <=( (not A201)  and  (not A200) );
 a23109a <=( (not A232)  and  A202 );
 a23110a <=( a23109a  and  a23106a );
 a23111a <=( a23110a  and  a23103a );
 a23115a <=( A236  and  (not A235) );
 a23116a <=( A233  and  a23115a );
 a23119a <=( A266  and  A265 );
 a23122a <=( (not A269)  and  A268 );
 a23123a <=( a23122a  and  a23119a );
 a23124a <=( a23123a  and  a23116a );
 a23128a <=( A199  and  (not A166) );
 a23129a <=( A167  and  a23128a );
 a23132a <=( (not A201)  and  (not A200) );
 a23135a <=( (not A232)  and  A202 );
 a23136a <=( a23135a  and  a23132a );
 a23137a <=( a23136a  and  a23129a );
 a23141a <=( A236  and  (not A235) );
 a23142a <=( A233  and  a23141a );
 a23145a <=( A266  and  (not A265) );
 a23148a <=( A269  and  (not A268) );
 a23149a <=( a23148a  and  a23145a );
 a23150a <=( a23149a  and  a23142a );
 a23154a <=( A199  and  (not A166) );
 a23155a <=( A167  and  a23154a );
 a23158a <=( (not A201)  and  (not A200) );
 a23161a <=( (not A232)  and  A202 );
 a23162a <=( a23161a  and  a23158a );
 a23163a <=( a23162a  and  a23155a );
 a23167a <=( A236  and  (not A235) );
 a23168a <=( A233  and  a23167a );
 a23171a <=( (not A266)  and  A265 );
 a23174a <=( A269  and  (not A268) );
 a23175a <=( a23174a  and  a23171a );
 a23176a <=( a23175a  and  a23168a );
 a23180a <=( A199  and  (not A166) );
 a23181a <=( A167  and  a23180a );
 a23184a <=( (not A201)  and  (not A200) );
 a23187a <=( (not A232)  and  A202 );
 a23188a <=( a23187a  and  a23184a );
 a23189a <=( a23188a  and  a23181a );
 a23193a <=( A236  and  (not A235) );
 a23194a <=( A233  and  a23193a );
 a23197a <=( (not A266)  and  (not A265) );
 a23200a <=( (not A269)  and  A268 );
 a23201a <=( a23200a  and  a23197a );
 a23202a <=( a23201a  and  a23194a );
 a23206a <=( A199  and  (not A166) );
 a23207a <=( A167  and  a23206a );
 a23210a <=( (not A201)  and  (not A200) );
 a23213a <=( A232  and  A202 );
 a23214a <=( a23213a  and  a23210a );
 a23215a <=( a23214a  and  a23207a );
 a23219a <=( A236  and  (not A235) );
 a23220a <=( (not A233)  and  a23219a );
 a23223a <=( A299  and  A298 );
 a23226a <=( (not A302)  and  A301 );
 a23227a <=( a23226a  and  a23223a );
 a23228a <=( a23227a  and  a23220a );
 a23232a <=( A199  and  (not A166) );
 a23233a <=( A167  and  a23232a );
 a23236a <=( (not A201)  and  (not A200) );
 a23239a <=( A232  and  A202 );
 a23240a <=( a23239a  and  a23236a );
 a23241a <=( a23240a  and  a23233a );
 a23245a <=( A236  and  (not A235) );
 a23246a <=( (not A233)  and  a23245a );
 a23249a <=( (not A299)  and  A298 );
 a23252a <=( A302  and  (not A301) );
 a23253a <=( a23252a  and  a23249a );
 a23254a <=( a23253a  and  a23246a );
 a23258a <=( A199  and  (not A166) );
 a23259a <=( A167  and  a23258a );
 a23262a <=( (not A201)  and  (not A200) );
 a23265a <=( A232  and  A202 );
 a23266a <=( a23265a  and  a23262a );
 a23267a <=( a23266a  and  a23259a );
 a23271a <=( A236  and  (not A235) );
 a23272a <=( (not A233)  and  a23271a );
 a23275a <=( A299  and  (not A298) );
 a23278a <=( A302  and  (not A301) );
 a23279a <=( a23278a  and  a23275a );
 a23280a <=( a23279a  and  a23272a );
 a23284a <=( A199  and  (not A166) );
 a23285a <=( A167  and  a23284a );
 a23288a <=( (not A201)  and  (not A200) );
 a23291a <=( A232  and  A202 );
 a23292a <=( a23291a  and  a23288a );
 a23293a <=( a23292a  and  a23285a );
 a23297a <=( A236  and  (not A235) );
 a23298a <=( (not A233)  and  a23297a );
 a23301a <=( (not A299)  and  (not A298) );
 a23304a <=( (not A302)  and  A301 );
 a23305a <=( a23304a  and  a23301a );
 a23306a <=( a23305a  and  a23298a );
 a23310a <=( A199  and  (not A166) );
 a23311a <=( A167  and  a23310a );
 a23314a <=( (not A201)  and  (not A200) );
 a23317a <=( A232  and  A202 );
 a23318a <=( a23317a  and  a23314a );
 a23319a <=( a23318a  and  a23311a );
 a23323a <=( A236  and  (not A235) );
 a23324a <=( (not A233)  and  a23323a );
 a23327a <=( A266  and  A265 );
 a23330a <=( (not A269)  and  A268 );
 a23331a <=( a23330a  and  a23327a );
 a23332a <=( a23331a  and  a23324a );
 a23336a <=( A199  and  (not A166) );
 a23337a <=( A167  and  a23336a );
 a23340a <=( (not A201)  and  (not A200) );
 a23343a <=( A232  and  A202 );
 a23344a <=( a23343a  and  a23340a );
 a23345a <=( a23344a  and  a23337a );
 a23349a <=( A236  and  (not A235) );
 a23350a <=( (not A233)  and  a23349a );
 a23353a <=( A266  and  (not A265) );
 a23356a <=( A269  and  (not A268) );
 a23357a <=( a23356a  and  a23353a );
 a23358a <=( a23357a  and  a23350a );
 a23362a <=( A199  and  (not A166) );
 a23363a <=( A167  and  a23362a );
 a23366a <=( (not A201)  and  (not A200) );
 a23369a <=( A232  and  A202 );
 a23370a <=( a23369a  and  a23366a );
 a23371a <=( a23370a  and  a23363a );
 a23375a <=( A236  and  (not A235) );
 a23376a <=( (not A233)  and  a23375a );
 a23379a <=( (not A266)  and  A265 );
 a23382a <=( A269  and  (not A268) );
 a23383a <=( a23382a  and  a23379a );
 a23384a <=( a23383a  and  a23376a );
 a23388a <=( A199  and  (not A166) );
 a23389a <=( A167  and  a23388a );
 a23392a <=( (not A201)  and  (not A200) );
 a23395a <=( A232  and  A202 );
 a23396a <=( a23395a  and  a23392a );
 a23397a <=( a23396a  and  a23389a );
 a23401a <=( A236  and  (not A235) );
 a23402a <=( (not A233)  and  a23401a );
 a23405a <=( (not A266)  and  (not A265) );
 a23408a <=( (not A269)  and  A268 );
 a23409a <=( a23408a  and  a23405a );
 a23410a <=( a23409a  and  a23402a );
 a23414a <=( A199  and  (not A166) );
 a23415a <=( A167  and  a23414a );
 a23418a <=( (not A201)  and  (not A200) );
 a23421a <=( (not A232)  and  A202 );
 a23422a <=( a23421a  and  a23418a );
 a23423a <=( a23422a  and  a23415a );
 a23427a <=( (not A236)  and  A235 );
 a23428a <=( (not A233)  and  a23427a );
 a23431a <=( A299  and  A298 );
 a23434a <=( (not A302)  and  A301 );
 a23435a <=( a23434a  and  a23431a );
 a23436a <=( a23435a  and  a23428a );
 a23440a <=( A199  and  (not A166) );
 a23441a <=( A167  and  a23440a );
 a23444a <=( (not A201)  and  (not A200) );
 a23447a <=( (not A232)  and  A202 );
 a23448a <=( a23447a  and  a23444a );
 a23449a <=( a23448a  and  a23441a );
 a23453a <=( (not A236)  and  A235 );
 a23454a <=( (not A233)  and  a23453a );
 a23457a <=( (not A299)  and  A298 );
 a23460a <=( A302  and  (not A301) );
 a23461a <=( a23460a  and  a23457a );
 a23462a <=( a23461a  and  a23454a );
 a23466a <=( A199  and  (not A166) );
 a23467a <=( A167  and  a23466a );
 a23470a <=( (not A201)  and  (not A200) );
 a23473a <=( (not A232)  and  A202 );
 a23474a <=( a23473a  and  a23470a );
 a23475a <=( a23474a  and  a23467a );
 a23479a <=( (not A236)  and  A235 );
 a23480a <=( (not A233)  and  a23479a );
 a23483a <=( A299  and  (not A298) );
 a23486a <=( A302  and  (not A301) );
 a23487a <=( a23486a  and  a23483a );
 a23488a <=( a23487a  and  a23480a );
 a23492a <=( A199  and  (not A166) );
 a23493a <=( A167  and  a23492a );
 a23496a <=( (not A201)  and  (not A200) );
 a23499a <=( (not A232)  and  A202 );
 a23500a <=( a23499a  and  a23496a );
 a23501a <=( a23500a  and  a23493a );
 a23505a <=( (not A236)  and  A235 );
 a23506a <=( (not A233)  and  a23505a );
 a23509a <=( (not A299)  and  (not A298) );
 a23512a <=( (not A302)  and  A301 );
 a23513a <=( a23512a  and  a23509a );
 a23514a <=( a23513a  and  a23506a );
 a23518a <=( A199  and  (not A166) );
 a23519a <=( A167  and  a23518a );
 a23522a <=( (not A201)  and  (not A200) );
 a23525a <=( (not A232)  and  A202 );
 a23526a <=( a23525a  and  a23522a );
 a23527a <=( a23526a  and  a23519a );
 a23531a <=( (not A236)  and  A235 );
 a23532a <=( (not A233)  and  a23531a );
 a23535a <=( A266  and  A265 );
 a23538a <=( (not A269)  and  A268 );
 a23539a <=( a23538a  and  a23535a );
 a23540a <=( a23539a  and  a23532a );
 a23544a <=( A199  and  (not A166) );
 a23545a <=( A167  and  a23544a );
 a23548a <=( (not A201)  and  (not A200) );
 a23551a <=( (not A232)  and  A202 );
 a23552a <=( a23551a  and  a23548a );
 a23553a <=( a23552a  and  a23545a );
 a23557a <=( (not A236)  and  A235 );
 a23558a <=( (not A233)  and  a23557a );
 a23561a <=( A266  and  (not A265) );
 a23564a <=( A269  and  (not A268) );
 a23565a <=( a23564a  and  a23561a );
 a23566a <=( a23565a  and  a23558a );
 a23570a <=( A199  and  (not A166) );
 a23571a <=( A167  and  a23570a );
 a23574a <=( (not A201)  and  (not A200) );
 a23577a <=( (not A232)  and  A202 );
 a23578a <=( a23577a  and  a23574a );
 a23579a <=( a23578a  and  a23571a );
 a23583a <=( (not A236)  and  A235 );
 a23584a <=( (not A233)  and  a23583a );
 a23587a <=( (not A266)  and  A265 );
 a23590a <=( A269  and  (not A268) );
 a23591a <=( a23590a  and  a23587a );
 a23592a <=( a23591a  and  a23584a );
 a23596a <=( A199  and  (not A166) );
 a23597a <=( A167  and  a23596a );
 a23600a <=( (not A201)  and  (not A200) );
 a23603a <=( (not A232)  and  A202 );
 a23604a <=( a23603a  and  a23600a );
 a23605a <=( a23604a  and  a23597a );
 a23609a <=( (not A236)  and  A235 );
 a23610a <=( (not A233)  and  a23609a );
 a23613a <=( (not A266)  and  (not A265) );
 a23616a <=( (not A269)  and  A268 );
 a23617a <=( a23616a  and  a23613a );
 a23618a <=( a23617a  and  a23610a );
 a23622a <=( A199  and  (not A166) );
 a23623a <=( A167  and  a23622a );
 a23626a <=( (not A201)  and  (not A200) );
 a23629a <=( A232  and  (not A203) );
 a23630a <=( a23629a  and  a23626a );
 a23631a <=( a23630a  and  a23623a );
 a23635a <=( (not A236)  and  A235 );
 a23636a <=( A233  and  a23635a );
 a23639a <=( A299  and  A298 );
 a23642a <=( (not A302)  and  A301 );
 a23643a <=( a23642a  and  a23639a );
 a23644a <=( a23643a  and  a23636a );
 a23648a <=( A199  and  (not A166) );
 a23649a <=( A167  and  a23648a );
 a23652a <=( (not A201)  and  (not A200) );
 a23655a <=( A232  and  (not A203) );
 a23656a <=( a23655a  and  a23652a );
 a23657a <=( a23656a  and  a23649a );
 a23661a <=( (not A236)  and  A235 );
 a23662a <=( A233  and  a23661a );
 a23665a <=( (not A299)  and  A298 );
 a23668a <=( A302  and  (not A301) );
 a23669a <=( a23668a  and  a23665a );
 a23670a <=( a23669a  and  a23662a );
 a23674a <=( A199  and  (not A166) );
 a23675a <=( A167  and  a23674a );
 a23678a <=( (not A201)  and  (not A200) );
 a23681a <=( A232  and  (not A203) );
 a23682a <=( a23681a  and  a23678a );
 a23683a <=( a23682a  and  a23675a );
 a23687a <=( (not A236)  and  A235 );
 a23688a <=( A233  and  a23687a );
 a23691a <=( A299  and  (not A298) );
 a23694a <=( A302  and  (not A301) );
 a23695a <=( a23694a  and  a23691a );
 a23696a <=( a23695a  and  a23688a );
 a23700a <=( A199  and  (not A166) );
 a23701a <=( A167  and  a23700a );
 a23704a <=( (not A201)  and  (not A200) );
 a23707a <=( A232  and  (not A203) );
 a23708a <=( a23707a  and  a23704a );
 a23709a <=( a23708a  and  a23701a );
 a23713a <=( (not A236)  and  A235 );
 a23714a <=( A233  and  a23713a );
 a23717a <=( (not A299)  and  (not A298) );
 a23720a <=( (not A302)  and  A301 );
 a23721a <=( a23720a  and  a23717a );
 a23722a <=( a23721a  and  a23714a );
 a23726a <=( A199  and  (not A166) );
 a23727a <=( A167  and  a23726a );
 a23730a <=( (not A201)  and  (not A200) );
 a23733a <=( A232  and  (not A203) );
 a23734a <=( a23733a  and  a23730a );
 a23735a <=( a23734a  and  a23727a );
 a23739a <=( (not A236)  and  A235 );
 a23740a <=( A233  and  a23739a );
 a23743a <=( A266  and  A265 );
 a23746a <=( (not A269)  and  A268 );
 a23747a <=( a23746a  and  a23743a );
 a23748a <=( a23747a  and  a23740a );
 a23752a <=( A199  and  (not A166) );
 a23753a <=( A167  and  a23752a );
 a23756a <=( (not A201)  and  (not A200) );
 a23759a <=( A232  and  (not A203) );
 a23760a <=( a23759a  and  a23756a );
 a23761a <=( a23760a  and  a23753a );
 a23765a <=( (not A236)  and  A235 );
 a23766a <=( A233  and  a23765a );
 a23769a <=( A266  and  (not A265) );
 a23772a <=( A269  and  (not A268) );
 a23773a <=( a23772a  and  a23769a );
 a23774a <=( a23773a  and  a23766a );
 a23778a <=( A199  and  (not A166) );
 a23779a <=( A167  and  a23778a );
 a23782a <=( (not A201)  and  (not A200) );
 a23785a <=( A232  and  (not A203) );
 a23786a <=( a23785a  and  a23782a );
 a23787a <=( a23786a  and  a23779a );
 a23791a <=( (not A236)  and  A235 );
 a23792a <=( A233  and  a23791a );
 a23795a <=( (not A266)  and  A265 );
 a23798a <=( A269  and  (not A268) );
 a23799a <=( a23798a  and  a23795a );
 a23800a <=( a23799a  and  a23792a );
 a23804a <=( A199  and  (not A166) );
 a23805a <=( A167  and  a23804a );
 a23808a <=( (not A201)  and  (not A200) );
 a23811a <=( A232  and  (not A203) );
 a23812a <=( a23811a  and  a23808a );
 a23813a <=( a23812a  and  a23805a );
 a23817a <=( (not A236)  and  A235 );
 a23818a <=( A233  and  a23817a );
 a23821a <=( (not A266)  and  (not A265) );
 a23824a <=( (not A269)  and  A268 );
 a23825a <=( a23824a  and  a23821a );
 a23826a <=( a23825a  and  a23818a );
 a23830a <=( A199  and  (not A166) );
 a23831a <=( A167  and  a23830a );
 a23834a <=( (not A201)  and  (not A200) );
 a23837a <=( (not A232)  and  (not A203) );
 a23838a <=( a23837a  and  a23834a );
 a23839a <=( a23838a  and  a23831a );
 a23843a <=( A236  and  (not A235) );
 a23844a <=( A233  and  a23843a );
 a23847a <=( A299  and  A298 );
 a23850a <=( (not A302)  and  A301 );
 a23851a <=( a23850a  and  a23847a );
 a23852a <=( a23851a  and  a23844a );
 a23856a <=( A199  and  (not A166) );
 a23857a <=( A167  and  a23856a );
 a23860a <=( (not A201)  and  (not A200) );
 a23863a <=( (not A232)  and  (not A203) );
 a23864a <=( a23863a  and  a23860a );
 a23865a <=( a23864a  and  a23857a );
 a23869a <=( A236  and  (not A235) );
 a23870a <=( A233  and  a23869a );
 a23873a <=( (not A299)  and  A298 );
 a23876a <=( A302  and  (not A301) );
 a23877a <=( a23876a  and  a23873a );
 a23878a <=( a23877a  and  a23870a );
 a23882a <=( A199  and  (not A166) );
 a23883a <=( A167  and  a23882a );
 a23886a <=( (not A201)  and  (not A200) );
 a23889a <=( (not A232)  and  (not A203) );
 a23890a <=( a23889a  and  a23886a );
 a23891a <=( a23890a  and  a23883a );
 a23895a <=( A236  and  (not A235) );
 a23896a <=( A233  and  a23895a );
 a23899a <=( A299  and  (not A298) );
 a23902a <=( A302  and  (not A301) );
 a23903a <=( a23902a  and  a23899a );
 a23904a <=( a23903a  and  a23896a );
 a23908a <=( A199  and  (not A166) );
 a23909a <=( A167  and  a23908a );
 a23912a <=( (not A201)  and  (not A200) );
 a23915a <=( (not A232)  and  (not A203) );
 a23916a <=( a23915a  and  a23912a );
 a23917a <=( a23916a  and  a23909a );
 a23921a <=( A236  and  (not A235) );
 a23922a <=( A233  and  a23921a );
 a23925a <=( (not A299)  and  (not A298) );
 a23928a <=( (not A302)  and  A301 );
 a23929a <=( a23928a  and  a23925a );
 a23930a <=( a23929a  and  a23922a );
 a23934a <=( A199  and  (not A166) );
 a23935a <=( A167  and  a23934a );
 a23938a <=( (not A201)  and  (not A200) );
 a23941a <=( (not A232)  and  (not A203) );
 a23942a <=( a23941a  and  a23938a );
 a23943a <=( a23942a  and  a23935a );
 a23947a <=( A236  and  (not A235) );
 a23948a <=( A233  and  a23947a );
 a23951a <=( A266  and  A265 );
 a23954a <=( (not A269)  and  A268 );
 a23955a <=( a23954a  and  a23951a );
 a23956a <=( a23955a  and  a23948a );
 a23960a <=( A199  and  (not A166) );
 a23961a <=( A167  and  a23960a );
 a23964a <=( (not A201)  and  (not A200) );
 a23967a <=( (not A232)  and  (not A203) );
 a23968a <=( a23967a  and  a23964a );
 a23969a <=( a23968a  and  a23961a );
 a23973a <=( A236  and  (not A235) );
 a23974a <=( A233  and  a23973a );
 a23977a <=( A266  and  (not A265) );
 a23980a <=( A269  and  (not A268) );
 a23981a <=( a23980a  and  a23977a );
 a23982a <=( a23981a  and  a23974a );
 a23986a <=( A199  and  (not A166) );
 a23987a <=( A167  and  a23986a );
 a23990a <=( (not A201)  and  (not A200) );
 a23993a <=( (not A232)  and  (not A203) );
 a23994a <=( a23993a  and  a23990a );
 a23995a <=( a23994a  and  a23987a );
 a23999a <=( A236  and  (not A235) );
 a24000a <=( A233  and  a23999a );
 a24003a <=( (not A266)  and  A265 );
 a24006a <=( A269  and  (not A268) );
 a24007a <=( a24006a  and  a24003a );
 a24008a <=( a24007a  and  a24000a );
 a24012a <=( A199  and  (not A166) );
 a24013a <=( A167  and  a24012a );
 a24016a <=( (not A201)  and  (not A200) );
 a24019a <=( (not A232)  and  (not A203) );
 a24020a <=( a24019a  and  a24016a );
 a24021a <=( a24020a  and  a24013a );
 a24025a <=( A236  and  (not A235) );
 a24026a <=( A233  and  a24025a );
 a24029a <=( (not A266)  and  (not A265) );
 a24032a <=( (not A269)  and  A268 );
 a24033a <=( a24032a  and  a24029a );
 a24034a <=( a24033a  and  a24026a );
 a24038a <=( A199  and  (not A166) );
 a24039a <=( A167  and  a24038a );
 a24042a <=( (not A201)  and  (not A200) );
 a24045a <=( A232  and  (not A203) );
 a24046a <=( a24045a  and  a24042a );
 a24047a <=( a24046a  and  a24039a );
 a24051a <=( A236  and  (not A235) );
 a24052a <=( (not A233)  and  a24051a );
 a24055a <=( A299  and  A298 );
 a24058a <=( (not A302)  and  A301 );
 a24059a <=( a24058a  and  a24055a );
 a24060a <=( a24059a  and  a24052a );
 a24064a <=( A199  and  (not A166) );
 a24065a <=( A167  and  a24064a );
 a24068a <=( (not A201)  and  (not A200) );
 a24071a <=( A232  and  (not A203) );
 a24072a <=( a24071a  and  a24068a );
 a24073a <=( a24072a  and  a24065a );
 a24077a <=( A236  and  (not A235) );
 a24078a <=( (not A233)  and  a24077a );
 a24081a <=( (not A299)  and  A298 );
 a24084a <=( A302  and  (not A301) );
 a24085a <=( a24084a  and  a24081a );
 a24086a <=( a24085a  and  a24078a );
 a24090a <=( A199  and  (not A166) );
 a24091a <=( A167  and  a24090a );
 a24094a <=( (not A201)  and  (not A200) );
 a24097a <=( A232  and  (not A203) );
 a24098a <=( a24097a  and  a24094a );
 a24099a <=( a24098a  and  a24091a );
 a24103a <=( A236  and  (not A235) );
 a24104a <=( (not A233)  and  a24103a );
 a24107a <=( A299  and  (not A298) );
 a24110a <=( A302  and  (not A301) );
 a24111a <=( a24110a  and  a24107a );
 a24112a <=( a24111a  and  a24104a );
 a24116a <=( A199  and  (not A166) );
 a24117a <=( A167  and  a24116a );
 a24120a <=( (not A201)  and  (not A200) );
 a24123a <=( A232  and  (not A203) );
 a24124a <=( a24123a  and  a24120a );
 a24125a <=( a24124a  and  a24117a );
 a24129a <=( A236  and  (not A235) );
 a24130a <=( (not A233)  and  a24129a );
 a24133a <=( (not A299)  and  (not A298) );
 a24136a <=( (not A302)  and  A301 );
 a24137a <=( a24136a  and  a24133a );
 a24138a <=( a24137a  and  a24130a );
 a24142a <=( A199  and  (not A166) );
 a24143a <=( A167  and  a24142a );
 a24146a <=( (not A201)  and  (not A200) );
 a24149a <=( A232  and  (not A203) );
 a24150a <=( a24149a  and  a24146a );
 a24151a <=( a24150a  and  a24143a );
 a24155a <=( A236  and  (not A235) );
 a24156a <=( (not A233)  and  a24155a );
 a24159a <=( A266  and  A265 );
 a24162a <=( (not A269)  and  A268 );
 a24163a <=( a24162a  and  a24159a );
 a24164a <=( a24163a  and  a24156a );
 a24168a <=( A199  and  (not A166) );
 a24169a <=( A167  and  a24168a );
 a24172a <=( (not A201)  and  (not A200) );
 a24175a <=( A232  and  (not A203) );
 a24176a <=( a24175a  and  a24172a );
 a24177a <=( a24176a  and  a24169a );
 a24181a <=( A236  and  (not A235) );
 a24182a <=( (not A233)  and  a24181a );
 a24185a <=( A266  and  (not A265) );
 a24188a <=( A269  and  (not A268) );
 a24189a <=( a24188a  and  a24185a );
 a24190a <=( a24189a  and  a24182a );
 a24194a <=( A199  and  (not A166) );
 a24195a <=( A167  and  a24194a );
 a24198a <=( (not A201)  and  (not A200) );
 a24201a <=( A232  and  (not A203) );
 a24202a <=( a24201a  and  a24198a );
 a24203a <=( a24202a  and  a24195a );
 a24207a <=( A236  and  (not A235) );
 a24208a <=( (not A233)  and  a24207a );
 a24211a <=( (not A266)  and  A265 );
 a24214a <=( A269  and  (not A268) );
 a24215a <=( a24214a  and  a24211a );
 a24216a <=( a24215a  and  a24208a );
 a24220a <=( A199  and  (not A166) );
 a24221a <=( A167  and  a24220a );
 a24224a <=( (not A201)  and  (not A200) );
 a24227a <=( A232  and  (not A203) );
 a24228a <=( a24227a  and  a24224a );
 a24229a <=( a24228a  and  a24221a );
 a24233a <=( A236  and  (not A235) );
 a24234a <=( (not A233)  and  a24233a );
 a24237a <=( (not A266)  and  (not A265) );
 a24240a <=( (not A269)  and  A268 );
 a24241a <=( a24240a  and  a24237a );
 a24242a <=( a24241a  and  a24234a );
 a24246a <=( A199  and  (not A166) );
 a24247a <=( A167  and  a24246a );
 a24250a <=( (not A201)  and  (not A200) );
 a24253a <=( (not A232)  and  (not A203) );
 a24254a <=( a24253a  and  a24250a );
 a24255a <=( a24254a  and  a24247a );
 a24259a <=( (not A236)  and  A235 );
 a24260a <=( (not A233)  and  a24259a );
 a24263a <=( A299  and  A298 );
 a24266a <=( (not A302)  and  A301 );
 a24267a <=( a24266a  and  a24263a );
 a24268a <=( a24267a  and  a24260a );
 a24272a <=( A199  and  (not A166) );
 a24273a <=( A167  and  a24272a );
 a24276a <=( (not A201)  and  (not A200) );
 a24279a <=( (not A232)  and  (not A203) );
 a24280a <=( a24279a  and  a24276a );
 a24281a <=( a24280a  and  a24273a );
 a24285a <=( (not A236)  and  A235 );
 a24286a <=( (not A233)  and  a24285a );
 a24289a <=( (not A299)  and  A298 );
 a24292a <=( A302  and  (not A301) );
 a24293a <=( a24292a  and  a24289a );
 a24294a <=( a24293a  and  a24286a );
 a24298a <=( A199  and  (not A166) );
 a24299a <=( A167  and  a24298a );
 a24302a <=( (not A201)  and  (not A200) );
 a24305a <=( (not A232)  and  (not A203) );
 a24306a <=( a24305a  and  a24302a );
 a24307a <=( a24306a  and  a24299a );
 a24311a <=( (not A236)  and  A235 );
 a24312a <=( (not A233)  and  a24311a );
 a24315a <=( A299  and  (not A298) );
 a24318a <=( A302  and  (not A301) );
 a24319a <=( a24318a  and  a24315a );
 a24320a <=( a24319a  and  a24312a );
 a24324a <=( A199  and  (not A166) );
 a24325a <=( A167  and  a24324a );
 a24328a <=( (not A201)  and  (not A200) );
 a24331a <=( (not A232)  and  (not A203) );
 a24332a <=( a24331a  and  a24328a );
 a24333a <=( a24332a  and  a24325a );
 a24337a <=( (not A236)  and  A235 );
 a24338a <=( (not A233)  and  a24337a );
 a24341a <=( (not A299)  and  (not A298) );
 a24344a <=( (not A302)  and  A301 );
 a24345a <=( a24344a  and  a24341a );
 a24346a <=( a24345a  and  a24338a );
 a24350a <=( A199  and  (not A166) );
 a24351a <=( A167  and  a24350a );
 a24354a <=( (not A201)  and  (not A200) );
 a24357a <=( (not A232)  and  (not A203) );
 a24358a <=( a24357a  and  a24354a );
 a24359a <=( a24358a  and  a24351a );
 a24363a <=( (not A236)  and  A235 );
 a24364a <=( (not A233)  and  a24363a );
 a24367a <=( A266  and  A265 );
 a24370a <=( (not A269)  and  A268 );
 a24371a <=( a24370a  and  a24367a );
 a24372a <=( a24371a  and  a24364a );
 a24376a <=( A199  and  (not A166) );
 a24377a <=( A167  and  a24376a );
 a24380a <=( (not A201)  and  (not A200) );
 a24383a <=( (not A232)  and  (not A203) );
 a24384a <=( a24383a  and  a24380a );
 a24385a <=( a24384a  and  a24377a );
 a24389a <=( (not A236)  and  A235 );
 a24390a <=( (not A233)  and  a24389a );
 a24393a <=( A266  and  (not A265) );
 a24396a <=( A269  and  (not A268) );
 a24397a <=( a24396a  and  a24393a );
 a24398a <=( a24397a  and  a24390a );
 a24402a <=( A199  and  (not A166) );
 a24403a <=( A167  and  a24402a );
 a24406a <=( (not A201)  and  (not A200) );
 a24409a <=( (not A232)  and  (not A203) );
 a24410a <=( a24409a  and  a24406a );
 a24411a <=( a24410a  and  a24403a );
 a24415a <=( (not A236)  and  A235 );
 a24416a <=( (not A233)  and  a24415a );
 a24419a <=( (not A266)  and  A265 );
 a24422a <=( A269  and  (not A268) );
 a24423a <=( a24422a  and  a24419a );
 a24424a <=( a24423a  and  a24416a );
 a24428a <=( A199  and  (not A166) );
 a24429a <=( A167  and  a24428a );
 a24432a <=( (not A201)  and  (not A200) );
 a24435a <=( (not A232)  and  (not A203) );
 a24436a <=( a24435a  and  a24432a );
 a24437a <=( a24436a  and  a24429a );
 a24441a <=( (not A236)  and  A235 );
 a24442a <=( (not A233)  and  a24441a );
 a24445a <=( (not A266)  and  (not A265) );
 a24448a <=( (not A269)  and  A268 );
 a24449a <=( a24448a  and  a24445a );
 a24450a <=( a24449a  and  a24442a );
 a24454a <=( (not A167)  and  A168 );
 a24455a <=( A170  and  a24454a );
 a24458a <=( A199  and  A166 );
 a24461a <=( (not A201)  and  A200 );
 a24462a <=( a24461a  and  a24458a );
 a24463a <=( a24462a  and  a24455a );
 a24467a <=( A234  and  A232 );
 a24468a <=( (not A202)  and  a24467a );
 a24471a <=( A299  and  A298 );
 a24474a <=( (not A302)  and  A301 );
 a24475a <=( a24474a  and  a24471a );
 a24476a <=( a24475a  and  a24468a );
 a24480a <=( (not A167)  and  A168 );
 a24481a <=( A170  and  a24480a );
 a24484a <=( A199  and  A166 );
 a24487a <=( (not A201)  and  A200 );
 a24488a <=( a24487a  and  a24484a );
 a24489a <=( a24488a  and  a24481a );
 a24493a <=( A234  and  A232 );
 a24494a <=( (not A202)  and  a24493a );
 a24497a <=( (not A299)  and  A298 );
 a24500a <=( A302  and  (not A301) );
 a24501a <=( a24500a  and  a24497a );
 a24502a <=( a24501a  and  a24494a );
 a24506a <=( (not A167)  and  A168 );
 a24507a <=( A170  and  a24506a );
 a24510a <=( A199  and  A166 );
 a24513a <=( (not A201)  and  A200 );
 a24514a <=( a24513a  and  a24510a );
 a24515a <=( a24514a  and  a24507a );
 a24519a <=( A234  and  A232 );
 a24520a <=( (not A202)  and  a24519a );
 a24523a <=( A299  and  (not A298) );
 a24526a <=( A302  and  (not A301) );
 a24527a <=( a24526a  and  a24523a );
 a24528a <=( a24527a  and  a24520a );
 a24532a <=( (not A167)  and  A168 );
 a24533a <=( A170  and  a24532a );
 a24536a <=( A199  and  A166 );
 a24539a <=( (not A201)  and  A200 );
 a24540a <=( a24539a  and  a24536a );
 a24541a <=( a24540a  and  a24533a );
 a24545a <=( A234  and  A232 );
 a24546a <=( (not A202)  and  a24545a );
 a24549a <=( (not A299)  and  (not A298) );
 a24552a <=( (not A302)  and  A301 );
 a24553a <=( a24552a  and  a24549a );
 a24554a <=( a24553a  and  a24546a );
 a24558a <=( (not A167)  and  A168 );
 a24559a <=( A170  and  a24558a );
 a24562a <=( A199  and  A166 );
 a24565a <=( (not A201)  and  A200 );
 a24566a <=( a24565a  and  a24562a );
 a24567a <=( a24566a  and  a24559a );
 a24571a <=( A234  and  A232 );
 a24572a <=( (not A202)  and  a24571a );
 a24575a <=( A266  and  A265 );
 a24578a <=( (not A269)  and  A268 );
 a24579a <=( a24578a  and  a24575a );
 a24580a <=( a24579a  and  a24572a );
 a24584a <=( (not A167)  and  A168 );
 a24585a <=( A170  and  a24584a );
 a24588a <=( A199  and  A166 );
 a24591a <=( (not A201)  and  A200 );
 a24592a <=( a24591a  and  a24588a );
 a24593a <=( a24592a  and  a24585a );
 a24597a <=( A234  and  A232 );
 a24598a <=( (not A202)  and  a24597a );
 a24601a <=( A266  and  (not A265) );
 a24604a <=( A269  and  (not A268) );
 a24605a <=( a24604a  and  a24601a );
 a24606a <=( a24605a  and  a24598a );
 a24610a <=( (not A167)  and  A168 );
 a24611a <=( A170  and  a24610a );
 a24614a <=( A199  and  A166 );
 a24617a <=( (not A201)  and  A200 );
 a24618a <=( a24617a  and  a24614a );
 a24619a <=( a24618a  and  a24611a );
 a24623a <=( A234  and  A232 );
 a24624a <=( (not A202)  and  a24623a );
 a24627a <=( (not A266)  and  A265 );
 a24630a <=( A269  and  (not A268) );
 a24631a <=( a24630a  and  a24627a );
 a24632a <=( a24631a  and  a24624a );
 a24636a <=( (not A167)  and  A168 );
 a24637a <=( A170  and  a24636a );
 a24640a <=( A199  and  A166 );
 a24643a <=( (not A201)  and  A200 );
 a24644a <=( a24643a  and  a24640a );
 a24645a <=( a24644a  and  a24637a );
 a24649a <=( A234  and  A232 );
 a24650a <=( (not A202)  and  a24649a );
 a24653a <=( (not A266)  and  (not A265) );
 a24656a <=( (not A269)  and  A268 );
 a24657a <=( a24656a  and  a24653a );
 a24658a <=( a24657a  and  a24650a );
 a24662a <=( (not A167)  and  A168 );
 a24663a <=( A170  and  a24662a );
 a24666a <=( A199  and  A166 );
 a24669a <=( (not A201)  and  A200 );
 a24670a <=( a24669a  and  a24666a );
 a24671a <=( a24670a  and  a24663a );
 a24675a <=( A234  and  A233 );
 a24676a <=( (not A202)  and  a24675a );
 a24679a <=( A299  and  A298 );
 a24682a <=( (not A302)  and  A301 );
 a24683a <=( a24682a  and  a24679a );
 a24684a <=( a24683a  and  a24676a );
 a24688a <=( (not A167)  and  A168 );
 a24689a <=( A170  and  a24688a );
 a24692a <=( A199  and  A166 );
 a24695a <=( (not A201)  and  A200 );
 a24696a <=( a24695a  and  a24692a );
 a24697a <=( a24696a  and  a24689a );
 a24701a <=( A234  and  A233 );
 a24702a <=( (not A202)  and  a24701a );
 a24705a <=( (not A299)  and  A298 );
 a24708a <=( A302  and  (not A301) );
 a24709a <=( a24708a  and  a24705a );
 a24710a <=( a24709a  and  a24702a );
 a24714a <=( (not A167)  and  A168 );
 a24715a <=( A170  and  a24714a );
 a24718a <=( A199  and  A166 );
 a24721a <=( (not A201)  and  A200 );
 a24722a <=( a24721a  and  a24718a );
 a24723a <=( a24722a  and  a24715a );
 a24727a <=( A234  and  A233 );
 a24728a <=( (not A202)  and  a24727a );
 a24731a <=( A299  and  (not A298) );
 a24734a <=( A302  and  (not A301) );
 a24735a <=( a24734a  and  a24731a );
 a24736a <=( a24735a  and  a24728a );
 a24740a <=( (not A167)  and  A168 );
 a24741a <=( A170  and  a24740a );
 a24744a <=( A199  and  A166 );
 a24747a <=( (not A201)  and  A200 );
 a24748a <=( a24747a  and  a24744a );
 a24749a <=( a24748a  and  a24741a );
 a24753a <=( A234  and  A233 );
 a24754a <=( (not A202)  and  a24753a );
 a24757a <=( (not A299)  and  (not A298) );
 a24760a <=( (not A302)  and  A301 );
 a24761a <=( a24760a  and  a24757a );
 a24762a <=( a24761a  and  a24754a );
 a24766a <=( (not A167)  and  A168 );
 a24767a <=( A170  and  a24766a );
 a24770a <=( A199  and  A166 );
 a24773a <=( (not A201)  and  A200 );
 a24774a <=( a24773a  and  a24770a );
 a24775a <=( a24774a  and  a24767a );
 a24779a <=( A234  and  A233 );
 a24780a <=( (not A202)  and  a24779a );
 a24783a <=( A266  and  A265 );
 a24786a <=( (not A269)  and  A268 );
 a24787a <=( a24786a  and  a24783a );
 a24788a <=( a24787a  and  a24780a );
 a24792a <=( (not A167)  and  A168 );
 a24793a <=( A170  and  a24792a );
 a24796a <=( A199  and  A166 );
 a24799a <=( (not A201)  and  A200 );
 a24800a <=( a24799a  and  a24796a );
 a24801a <=( a24800a  and  a24793a );
 a24805a <=( A234  and  A233 );
 a24806a <=( (not A202)  and  a24805a );
 a24809a <=( A266  and  (not A265) );
 a24812a <=( A269  and  (not A268) );
 a24813a <=( a24812a  and  a24809a );
 a24814a <=( a24813a  and  a24806a );
 a24818a <=( (not A167)  and  A168 );
 a24819a <=( A170  and  a24818a );
 a24822a <=( A199  and  A166 );
 a24825a <=( (not A201)  and  A200 );
 a24826a <=( a24825a  and  a24822a );
 a24827a <=( a24826a  and  a24819a );
 a24831a <=( A234  and  A233 );
 a24832a <=( (not A202)  and  a24831a );
 a24835a <=( (not A266)  and  A265 );
 a24838a <=( A269  and  (not A268) );
 a24839a <=( a24838a  and  a24835a );
 a24840a <=( a24839a  and  a24832a );
 a24844a <=( (not A167)  and  A168 );
 a24845a <=( A170  and  a24844a );
 a24848a <=( A199  and  A166 );
 a24851a <=( (not A201)  and  A200 );
 a24852a <=( a24851a  and  a24848a );
 a24853a <=( a24852a  and  a24845a );
 a24857a <=( A234  and  A233 );
 a24858a <=( (not A202)  and  a24857a );
 a24861a <=( (not A266)  and  (not A265) );
 a24864a <=( (not A269)  and  A268 );
 a24865a <=( a24864a  and  a24861a );
 a24866a <=( a24865a  and  a24858a );
 a24870a <=( (not A167)  and  A168 );
 a24871a <=( A170  and  a24870a );
 a24874a <=( A199  and  A166 );
 a24877a <=( (not A201)  and  A200 );
 a24878a <=( a24877a  and  a24874a );
 a24879a <=( a24878a  and  a24871a );
 a24883a <=( A233  and  A232 );
 a24884a <=( (not A202)  and  a24883a );
 a24887a <=( (not A236)  and  A235 );
 a24890a <=( A300  and  A299 );
 a24891a <=( a24890a  and  a24887a );
 a24892a <=( a24891a  and  a24884a );
 a24896a <=( (not A167)  and  A168 );
 a24897a <=( A170  and  a24896a );
 a24900a <=( A199  and  A166 );
 a24903a <=( (not A201)  and  A200 );
 a24904a <=( a24903a  and  a24900a );
 a24905a <=( a24904a  and  a24897a );
 a24909a <=( A233  and  A232 );
 a24910a <=( (not A202)  and  a24909a );
 a24913a <=( (not A236)  and  A235 );
 a24916a <=( A300  and  A298 );
 a24917a <=( a24916a  and  a24913a );
 a24918a <=( a24917a  and  a24910a );
 a24922a <=( (not A167)  and  A168 );
 a24923a <=( A170  and  a24922a );
 a24926a <=( A199  and  A166 );
 a24929a <=( (not A201)  and  A200 );
 a24930a <=( a24929a  and  a24926a );
 a24931a <=( a24930a  and  a24923a );
 a24935a <=( A233  and  A232 );
 a24936a <=( (not A202)  and  a24935a );
 a24939a <=( (not A236)  and  A235 );
 a24942a <=( A267  and  A265 );
 a24943a <=( a24942a  and  a24939a );
 a24944a <=( a24943a  and  a24936a );
 a24948a <=( (not A167)  and  A168 );
 a24949a <=( A170  and  a24948a );
 a24952a <=( A199  and  A166 );
 a24955a <=( (not A201)  and  A200 );
 a24956a <=( a24955a  and  a24952a );
 a24957a <=( a24956a  and  a24949a );
 a24961a <=( A233  and  A232 );
 a24962a <=( (not A202)  and  a24961a );
 a24965a <=( (not A236)  and  A235 );
 a24968a <=( A267  and  A266 );
 a24969a <=( a24968a  and  a24965a );
 a24970a <=( a24969a  and  a24962a );
 a24974a <=( (not A167)  and  A168 );
 a24975a <=( A170  and  a24974a );
 a24978a <=( A199  and  A166 );
 a24981a <=( (not A201)  and  A200 );
 a24982a <=( a24981a  and  a24978a );
 a24983a <=( a24982a  and  a24975a );
 a24987a <=( A233  and  (not A232) );
 a24988a <=( (not A202)  and  a24987a );
 a24991a <=( A236  and  (not A235) );
 a24994a <=( A300  and  A299 );
 a24995a <=( a24994a  and  a24991a );
 a24996a <=( a24995a  and  a24988a );
 a25000a <=( (not A167)  and  A168 );
 a25001a <=( A170  and  a25000a );
 a25004a <=( A199  and  A166 );
 a25007a <=( (not A201)  and  A200 );
 a25008a <=( a25007a  and  a25004a );
 a25009a <=( a25008a  and  a25001a );
 a25013a <=( A233  and  (not A232) );
 a25014a <=( (not A202)  and  a25013a );
 a25017a <=( A236  and  (not A235) );
 a25020a <=( A300  and  A298 );
 a25021a <=( a25020a  and  a25017a );
 a25022a <=( a25021a  and  a25014a );
 a25026a <=( (not A167)  and  A168 );
 a25027a <=( A170  and  a25026a );
 a25030a <=( A199  and  A166 );
 a25033a <=( (not A201)  and  A200 );
 a25034a <=( a25033a  and  a25030a );
 a25035a <=( a25034a  and  a25027a );
 a25039a <=( A233  and  (not A232) );
 a25040a <=( (not A202)  and  a25039a );
 a25043a <=( A236  and  (not A235) );
 a25046a <=( A267  and  A265 );
 a25047a <=( a25046a  and  a25043a );
 a25048a <=( a25047a  and  a25040a );
 a25052a <=( (not A167)  and  A168 );
 a25053a <=( A170  and  a25052a );
 a25056a <=( A199  and  A166 );
 a25059a <=( (not A201)  and  A200 );
 a25060a <=( a25059a  and  a25056a );
 a25061a <=( a25060a  and  a25053a );
 a25065a <=( A233  and  (not A232) );
 a25066a <=( (not A202)  and  a25065a );
 a25069a <=( A236  and  (not A235) );
 a25072a <=( A267  and  A266 );
 a25073a <=( a25072a  and  a25069a );
 a25074a <=( a25073a  and  a25066a );
 a25078a <=( (not A167)  and  A168 );
 a25079a <=( A170  and  a25078a );
 a25082a <=( A199  and  A166 );
 a25085a <=( (not A201)  and  A200 );
 a25086a <=( a25085a  and  a25082a );
 a25087a <=( a25086a  and  a25079a );
 a25091a <=( (not A233)  and  A232 );
 a25092a <=( (not A202)  and  a25091a );
 a25095a <=( A236  and  (not A235) );
 a25098a <=( A300  and  A299 );
 a25099a <=( a25098a  and  a25095a );
 a25100a <=( a25099a  and  a25092a );
 a25104a <=( (not A167)  and  A168 );
 a25105a <=( A170  and  a25104a );
 a25108a <=( A199  and  A166 );
 a25111a <=( (not A201)  and  A200 );
 a25112a <=( a25111a  and  a25108a );
 a25113a <=( a25112a  and  a25105a );
 a25117a <=( (not A233)  and  A232 );
 a25118a <=( (not A202)  and  a25117a );
 a25121a <=( A236  and  (not A235) );
 a25124a <=( A300  and  A298 );
 a25125a <=( a25124a  and  a25121a );
 a25126a <=( a25125a  and  a25118a );
 a25130a <=( (not A167)  and  A168 );
 a25131a <=( A170  and  a25130a );
 a25134a <=( A199  and  A166 );
 a25137a <=( (not A201)  and  A200 );
 a25138a <=( a25137a  and  a25134a );
 a25139a <=( a25138a  and  a25131a );
 a25143a <=( (not A233)  and  A232 );
 a25144a <=( (not A202)  and  a25143a );
 a25147a <=( A236  and  (not A235) );
 a25150a <=( A267  and  A265 );
 a25151a <=( a25150a  and  a25147a );
 a25152a <=( a25151a  and  a25144a );
 a25156a <=( (not A167)  and  A168 );
 a25157a <=( A170  and  a25156a );
 a25160a <=( A199  and  A166 );
 a25163a <=( (not A201)  and  A200 );
 a25164a <=( a25163a  and  a25160a );
 a25165a <=( a25164a  and  a25157a );
 a25169a <=( (not A233)  and  A232 );
 a25170a <=( (not A202)  and  a25169a );
 a25173a <=( A236  and  (not A235) );
 a25176a <=( A267  and  A266 );
 a25177a <=( a25176a  and  a25173a );
 a25178a <=( a25177a  and  a25170a );
 a25182a <=( (not A167)  and  A168 );
 a25183a <=( A170  and  a25182a );
 a25186a <=( A199  and  A166 );
 a25189a <=( (not A201)  and  A200 );
 a25190a <=( a25189a  and  a25186a );
 a25191a <=( a25190a  and  a25183a );
 a25195a <=( (not A233)  and  (not A232) );
 a25196a <=( (not A202)  and  a25195a );
 a25199a <=( (not A236)  and  A235 );
 a25202a <=( A300  and  A299 );
 a25203a <=( a25202a  and  a25199a );
 a25204a <=( a25203a  and  a25196a );
 a25208a <=( (not A167)  and  A168 );
 a25209a <=( A170  and  a25208a );
 a25212a <=( A199  and  A166 );
 a25215a <=( (not A201)  and  A200 );
 a25216a <=( a25215a  and  a25212a );
 a25217a <=( a25216a  and  a25209a );
 a25221a <=( (not A233)  and  (not A232) );
 a25222a <=( (not A202)  and  a25221a );
 a25225a <=( (not A236)  and  A235 );
 a25228a <=( A300  and  A298 );
 a25229a <=( a25228a  and  a25225a );
 a25230a <=( a25229a  and  a25222a );
 a25234a <=( (not A167)  and  A168 );
 a25235a <=( A170  and  a25234a );
 a25238a <=( A199  and  A166 );
 a25241a <=( (not A201)  and  A200 );
 a25242a <=( a25241a  and  a25238a );
 a25243a <=( a25242a  and  a25235a );
 a25247a <=( (not A233)  and  (not A232) );
 a25248a <=( (not A202)  and  a25247a );
 a25251a <=( (not A236)  and  A235 );
 a25254a <=( A267  and  A265 );
 a25255a <=( a25254a  and  a25251a );
 a25256a <=( a25255a  and  a25248a );
 a25260a <=( (not A167)  and  A168 );
 a25261a <=( A170  and  a25260a );
 a25264a <=( A199  and  A166 );
 a25267a <=( (not A201)  and  A200 );
 a25268a <=( a25267a  and  a25264a );
 a25269a <=( a25268a  and  a25261a );
 a25273a <=( (not A233)  and  (not A232) );
 a25274a <=( (not A202)  and  a25273a );
 a25277a <=( (not A236)  and  A235 );
 a25280a <=( A267  and  A266 );
 a25281a <=( a25280a  and  a25277a );
 a25282a <=( a25281a  and  a25274a );
 a25286a <=( (not A167)  and  A168 );
 a25287a <=( A170  and  a25286a );
 a25290a <=( A199  and  A166 );
 a25293a <=( (not A201)  and  A200 );
 a25294a <=( a25293a  and  a25290a );
 a25295a <=( a25294a  and  a25287a );
 a25299a <=( A234  and  A232 );
 a25300a <=( A203  and  a25299a );
 a25303a <=( A299  and  A298 );
 a25306a <=( (not A302)  and  A301 );
 a25307a <=( a25306a  and  a25303a );
 a25308a <=( a25307a  and  a25300a );
 a25312a <=( (not A167)  and  A168 );
 a25313a <=( A170  and  a25312a );
 a25316a <=( A199  and  A166 );
 a25319a <=( (not A201)  and  A200 );
 a25320a <=( a25319a  and  a25316a );
 a25321a <=( a25320a  and  a25313a );
 a25325a <=( A234  and  A232 );
 a25326a <=( A203  and  a25325a );
 a25329a <=( (not A299)  and  A298 );
 a25332a <=( A302  and  (not A301) );
 a25333a <=( a25332a  and  a25329a );
 a25334a <=( a25333a  and  a25326a );
 a25338a <=( (not A167)  and  A168 );
 a25339a <=( A170  and  a25338a );
 a25342a <=( A199  and  A166 );
 a25345a <=( (not A201)  and  A200 );
 a25346a <=( a25345a  and  a25342a );
 a25347a <=( a25346a  and  a25339a );
 a25351a <=( A234  and  A232 );
 a25352a <=( A203  and  a25351a );
 a25355a <=( A299  and  (not A298) );
 a25358a <=( A302  and  (not A301) );
 a25359a <=( a25358a  and  a25355a );
 a25360a <=( a25359a  and  a25352a );
 a25364a <=( (not A167)  and  A168 );
 a25365a <=( A170  and  a25364a );
 a25368a <=( A199  and  A166 );
 a25371a <=( (not A201)  and  A200 );
 a25372a <=( a25371a  and  a25368a );
 a25373a <=( a25372a  and  a25365a );
 a25377a <=( A234  and  A232 );
 a25378a <=( A203  and  a25377a );
 a25381a <=( (not A299)  and  (not A298) );
 a25384a <=( (not A302)  and  A301 );
 a25385a <=( a25384a  and  a25381a );
 a25386a <=( a25385a  and  a25378a );
 a25390a <=( (not A167)  and  A168 );
 a25391a <=( A170  and  a25390a );
 a25394a <=( A199  and  A166 );
 a25397a <=( (not A201)  and  A200 );
 a25398a <=( a25397a  and  a25394a );
 a25399a <=( a25398a  and  a25391a );
 a25403a <=( A234  and  A232 );
 a25404a <=( A203  and  a25403a );
 a25407a <=( A266  and  A265 );
 a25410a <=( (not A269)  and  A268 );
 a25411a <=( a25410a  and  a25407a );
 a25412a <=( a25411a  and  a25404a );
 a25416a <=( (not A167)  and  A168 );
 a25417a <=( A170  and  a25416a );
 a25420a <=( A199  and  A166 );
 a25423a <=( (not A201)  and  A200 );
 a25424a <=( a25423a  and  a25420a );
 a25425a <=( a25424a  and  a25417a );
 a25429a <=( A234  and  A232 );
 a25430a <=( A203  and  a25429a );
 a25433a <=( A266  and  (not A265) );
 a25436a <=( A269  and  (not A268) );
 a25437a <=( a25436a  and  a25433a );
 a25438a <=( a25437a  and  a25430a );
 a25442a <=( (not A167)  and  A168 );
 a25443a <=( A170  and  a25442a );
 a25446a <=( A199  and  A166 );
 a25449a <=( (not A201)  and  A200 );
 a25450a <=( a25449a  and  a25446a );
 a25451a <=( a25450a  and  a25443a );
 a25455a <=( A234  and  A232 );
 a25456a <=( A203  and  a25455a );
 a25459a <=( (not A266)  and  A265 );
 a25462a <=( A269  and  (not A268) );
 a25463a <=( a25462a  and  a25459a );
 a25464a <=( a25463a  and  a25456a );
 a25468a <=( (not A167)  and  A168 );
 a25469a <=( A170  and  a25468a );
 a25472a <=( A199  and  A166 );
 a25475a <=( (not A201)  and  A200 );
 a25476a <=( a25475a  and  a25472a );
 a25477a <=( a25476a  and  a25469a );
 a25481a <=( A234  and  A232 );
 a25482a <=( A203  and  a25481a );
 a25485a <=( (not A266)  and  (not A265) );
 a25488a <=( (not A269)  and  A268 );
 a25489a <=( a25488a  and  a25485a );
 a25490a <=( a25489a  and  a25482a );
 a25494a <=( (not A167)  and  A168 );
 a25495a <=( A170  and  a25494a );
 a25498a <=( A199  and  A166 );
 a25501a <=( (not A201)  and  A200 );
 a25502a <=( a25501a  and  a25498a );
 a25503a <=( a25502a  and  a25495a );
 a25507a <=( A234  and  A233 );
 a25508a <=( A203  and  a25507a );
 a25511a <=( A299  and  A298 );
 a25514a <=( (not A302)  and  A301 );
 a25515a <=( a25514a  and  a25511a );
 a25516a <=( a25515a  and  a25508a );
 a25520a <=( (not A167)  and  A168 );
 a25521a <=( A170  and  a25520a );
 a25524a <=( A199  and  A166 );
 a25527a <=( (not A201)  and  A200 );
 a25528a <=( a25527a  and  a25524a );
 a25529a <=( a25528a  and  a25521a );
 a25533a <=( A234  and  A233 );
 a25534a <=( A203  and  a25533a );
 a25537a <=( (not A299)  and  A298 );
 a25540a <=( A302  and  (not A301) );
 a25541a <=( a25540a  and  a25537a );
 a25542a <=( a25541a  and  a25534a );
 a25546a <=( (not A167)  and  A168 );
 a25547a <=( A170  and  a25546a );
 a25550a <=( A199  and  A166 );
 a25553a <=( (not A201)  and  A200 );
 a25554a <=( a25553a  and  a25550a );
 a25555a <=( a25554a  and  a25547a );
 a25559a <=( A234  and  A233 );
 a25560a <=( A203  and  a25559a );
 a25563a <=( A299  and  (not A298) );
 a25566a <=( A302  and  (not A301) );
 a25567a <=( a25566a  and  a25563a );
 a25568a <=( a25567a  and  a25560a );
 a25572a <=( (not A167)  and  A168 );
 a25573a <=( A170  and  a25572a );
 a25576a <=( A199  and  A166 );
 a25579a <=( (not A201)  and  A200 );
 a25580a <=( a25579a  and  a25576a );
 a25581a <=( a25580a  and  a25573a );
 a25585a <=( A234  and  A233 );
 a25586a <=( A203  and  a25585a );
 a25589a <=( (not A299)  and  (not A298) );
 a25592a <=( (not A302)  and  A301 );
 a25593a <=( a25592a  and  a25589a );
 a25594a <=( a25593a  and  a25586a );
 a25598a <=( (not A167)  and  A168 );
 a25599a <=( A170  and  a25598a );
 a25602a <=( A199  and  A166 );
 a25605a <=( (not A201)  and  A200 );
 a25606a <=( a25605a  and  a25602a );
 a25607a <=( a25606a  and  a25599a );
 a25611a <=( A234  and  A233 );
 a25612a <=( A203  and  a25611a );
 a25615a <=( A266  and  A265 );
 a25618a <=( (not A269)  and  A268 );
 a25619a <=( a25618a  and  a25615a );
 a25620a <=( a25619a  and  a25612a );
 a25624a <=( (not A167)  and  A168 );
 a25625a <=( A170  and  a25624a );
 a25628a <=( A199  and  A166 );
 a25631a <=( (not A201)  and  A200 );
 a25632a <=( a25631a  and  a25628a );
 a25633a <=( a25632a  and  a25625a );
 a25637a <=( A234  and  A233 );
 a25638a <=( A203  and  a25637a );
 a25641a <=( A266  and  (not A265) );
 a25644a <=( A269  and  (not A268) );
 a25645a <=( a25644a  and  a25641a );
 a25646a <=( a25645a  and  a25638a );
 a25650a <=( (not A167)  and  A168 );
 a25651a <=( A170  and  a25650a );
 a25654a <=( A199  and  A166 );
 a25657a <=( (not A201)  and  A200 );
 a25658a <=( a25657a  and  a25654a );
 a25659a <=( a25658a  and  a25651a );
 a25663a <=( A234  and  A233 );
 a25664a <=( A203  and  a25663a );
 a25667a <=( (not A266)  and  A265 );
 a25670a <=( A269  and  (not A268) );
 a25671a <=( a25670a  and  a25667a );
 a25672a <=( a25671a  and  a25664a );
 a25676a <=( (not A167)  and  A168 );
 a25677a <=( A170  and  a25676a );
 a25680a <=( A199  and  A166 );
 a25683a <=( (not A201)  and  A200 );
 a25684a <=( a25683a  and  a25680a );
 a25685a <=( a25684a  and  a25677a );
 a25689a <=( A234  and  A233 );
 a25690a <=( A203  and  a25689a );
 a25693a <=( (not A266)  and  (not A265) );
 a25696a <=( (not A269)  and  A268 );
 a25697a <=( a25696a  and  a25693a );
 a25698a <=( a25697a  and  a25690a );
 a25702a <=( (not A167)  and  A168 );
 a25703a <=( A170  and  a25702a );
 a25706a <=( A199  and  A166 );
 a25709a <=( (not A201)  and  A200 );
 a25710a <=( a25709a  and  a25706a );
 a25711a <=( a25710a  and  a25703a );
 a25715a <=( A233  and  A232 );
 a25716a <=( A203  and  a25715a );
 a25719a <=( (not A236)  and  A235 );
 a25722a <=( A300  and  A299 );
 a25723a <=( a25722a  and  a25719a );
 a25724a <=( a25723a  and  a25716a );
 a25728a <=( (not A167)  and  A168 );
 a25729a <=( A170  and  a25728a );
 a25732a <=( A199  and  A166 );
 a25735a <=( (not A201)  and  A200 );
 a25736a <=( a25735a  and  a25732a );
 a25737a <=( a25736a  and  a25729a );
 a25741a <=( A233  and  A232 );
 a25742a <=( A203  and  a25741a );
 a25745a <=( (not A236)  and  A235 );
 a25748a <=( A300  and  A298 );
 a25749a <=( a25748a  and  a25745a );
 a25750a <=( a25749a  and  a25742a );
 a25754a <=( (not A167)  and  A168 );
 a25755a <=( A170  and  a25754a );
 a25758a <=( A199  and  A166 );
 a25761a <=( (not A201)  and  A200 );
 a25762a <=( a25761a  and  a25758a );
 a25763a <=( a25762a  and  a25755a );
 a25767a <=( A233  and  A232 );
 a25768a <=( A203  and  a25767a );
 a25771a <=( (not A236)  and  A235 );
 a25774a <=( A267  and  A265 );
 a25775a <=( a25774a  and  a25771a );
 a25776a <=( a25775a  and  a25768a );
 a25780a <=( (not A167)  and  A168 );
 a25781a <=( A170  and  a25780a );
 a25784a <=( A199  and  A166 );
 a25787a <=( (not A201)  and  A200 );
 a25788a <=( a25787a  and  a25784a );
 a25789a <=( a25788a  and  a25781a );
 a25793a <=( A233  and  A232 );
 a25794a <=( A203  and  a25793a );
 a25797a <=( (not A236)  and  A235 );
 a25800a <=( A267  and  A266 );
 a25801a <=( a25800a  and  a25797a );
 a25802a <=( a25801a  and  a25794a );
 a25806a <=( (not A167)  and  A168 );
 a25807a <=( A170  and  a25806a );
 a25810a <=( A199  and  A166 );
 a25813a <=( (not A201)  and  A200 );
 a25814a <=( a25813a  and  a25810a );
 a25815a <=( a25814a  and  a25807a );
 a25819a <=( A233  and  (not A232) );
 a25820a <=( A203  and  a25819a );
 a25823a <=( A236  and  (not A235) );
 a25826a <=( A300  and  A299 );
 a25827a <=( a25826a  and  a25823a );
 a25828a <=( a25827a  and  a25820a );
 a25832a <=( (not A167)  and  A168 );
 a25833a <=( A170  and  a25832a );
 a25836a <=( A199  and  A166 );
 a25839a <=( (not A201)  and  A200 );
 a25840a <=( a25839a  and  a25836a );
 a25841a <=( a25840a  and  a25833a );
 a25845a <=( A233  and  (not A232) );
 a25846a <=( A203  and  a25845a );
 a25849a <=( A236  and  (not A235) );
 a25852a <=( A300  and  A298 );
 a25853a <=( a25852a  and  a25849a );
 a25854a <=( a25853a  and  a25846a );
 a25858a <=( (not A167)  and  A168 );
 a25859a <=( A170  and  a25858a );
 a25862a <=( A199  and  A166 );
 a25865a <=( (not A201)  and  A200 );
 a25866a <=( a25865a  and  a25862a );
 a25867a <=( a25866a  and  a25859a );
 a25871a <=( A233  and  (not A232) );
 a25872a <=( A203  and  a25871a );
 a25875a <=( A236  and  (not A235) );
 a25878a <=( A267  and  A265 );
 a25879a <=( a25878a  and  a25875a );
 a25880a <=( a25879a  and  a25872a );
 a25884a <=( (not A167)  and  A168 );
 a25885a <=( A170  and  a25884a );
 a25888a <=( A199  and  A166 );
 a25891a <=( (not A201)  and  A200 );
 a25892a <=( a25891a  and  a25888a );
 a25893a <=( a25892a  and  a25885a );
 a25897a <=( A233  and  (not A232) );
 a25898a <=( A203  and  a25897a );
 a25901a <=( A236  and  (not A235) );
 a25904a <=( A267  and  A266 );
 a25905a <=( a25904a  and  a25901a );
 a25906a <=( a25905a  and  a25898a );
 a25910a <=( (not A167)  and  A168 );
 a25911a <=( A170  and  a25910a );
 a25914a <=( A199  and  A166 );
 a25917a <=( (not A201)  and  A200 );
 a25918a <=( a25917a  and  a25914a );
 a25919a <=( a25918a  and  a25911a );
 a25923a <=( (not A233)  and  A232 );
 a25924a <=( A203  and  a25923a );
 a25927a <=( A236  and  (not A235) );
 a25930a <=( A300  and  A299 );
 a25931a <=( a25930a  and  a25927a );
 a25932a <=( a25931a  and  a25924a );
 a25936a <=( (not A167)  and  A168 );
 a25937a <=( A170  and  a25936a );
 a25940a <=( A199  and  A166 );
 a25943a <=( (not A201)  and  A200 );
 a25944a <=( a25943a  and  a25940a );
 a25945a <=( a25944a  and  a25937a );
 a25949a <=( (not A233)  and  A232 );
 a25950a <=( A203  and  a25949a );
 a25953a <=( A236  and  (not A235) );
 a25956a <=( A300  and  A298 );
 a25957a <=( a25956a  and  a25953a );
 a25958a <=( a25957a  and  a25950a );
 a25962a <=( (not A167)  and  A168 );
 a25963a <=( A170  and  a25962a );
 a25966a <=( A199  and  A166 );
 a25969a <=( (not A201)  and  A200 );
 a25970a <=( a25969a  and  a25966a );
 a25971a <=( a25970a  and  a25963a );
 a25975a <=( (not A233)  and  A232 );
 a25976a <=( A203  and  a25975a );
 a25979a <=( A236  and  (not A235) );
 a25982a <=( A267  and  A265 );
 a25983a <=( a25982a  and  a25979a );
 a25984a <=( a25983a  and  a25976a );
 a25988a <=( (not A167)  and  A168 );
 a25989a <=( A170  and  a25988a );
 a25992a <=( A199  and  A166 );
 a25995a <=( (not A201)  and  A200 );
 a25996a <=( a25995a  and  a25992a );
 a25997a <=( a25996a  and  a25989a );
 a26001a <=( (not A233)  and  A232 );
 a26002a <=( A203  and  a26001a );
 a26005a <=( A236  and  (not A235) );
 a26008a <=( A267  and  A266 );
 a26009a <=( a26008a  and  a26005a );
 a26010a <=( a26009a  and  a26002a );
 a26014a <=( (not A167)  and  A168 );
 a26015a <=( A170  and  a26014a );
 a26018a <=( A199  and  A166 );
 a26021a <=( (not A201)  and  A200 );
 a26022a <=( a26021a  and  a26018a );
 a26023a <=( a26022a  and  a26015a );
 a26027a <=( (not A233)  and  (not A232) );
 a26028a <=( A203  and  a26027a );
 a26031a <=( (not A236)  and  A235 );
 a26034a <=( A300  and  A299 );
 a26035a <=( a26034a  and  a26031a );
 a26036a <=( a26035a  and  a26028a );
 a26040a <=( (not A167)  and  A168 );
 a26041a <=( A170  and  a26040a );
 a26044a <=( A199  and  A166 );
 a26047a <=( (not A201)  and  A200 );
 a26048a <=( a26047a  and  a26044a );
 a26049a <=( a26048a  and  a26041a );
 a26053a <=( (not A233)  and  (not A232) );
 a26054a <=( A203  and  a26053a );
 a26057a <=( (not A236)  and  A235 );
 a26060a <=( A300  and  A298 );
 a26061a <=( a26060a  and  a26057a );
 a26062a <=( a26061a  and  a26054a );
 a26066a <=( (not A167)  and  A168 );
 a26067a <=( A170  and  a26066a );
 a26070a <=( A199  and  A166 );
 a26073a <=( (not A201)  and  A200 );
 a26074a <=( a26073a  and  a26070a );
 a26075a <=( a26074a  and  a26067a );
 a26079a <=( (not A233)  and  (not A232) );
 a26080a <=( A203  and  a26079a );
 a26083a <=( (not A236)  and  A235 );
 a26086a <=( A267  and  A265 );
 a26087a <=( a26086a  and  a26083a );
 a26088a <=( a26087a  and  a26080a );
 a26092a <=( (not A167)  and  A168 );
 a26093a <=( A170  and  a26092a );
 a26096a <=( A199  and  A166 );
 a26099a <=( (not A201)  and  A200 );
 a26100a <=( a26099a  and  a26096a );
 a26101a <=( a26100a  and  a26093a );
 a26105a <=( (not A233)  and  (not A232) );
 a26106a <=( A203  and  a26105a );
 a26109a <=( (not A236)  and  A235 );
 a26112a <=( A267  and  A266 );
 a26113a <=( a26112a  and  a26109a );
 a26114a <=( a26113a  and  a26106a );
 a26118a <=( (not A167)  and  A168 );
 a26119a <=( A170  and  a26118a );
 a26122a <=( (not A199)  and  A166 );
 a26125a <=( (not A201)  and  A200 );
 a26126a <=( a26125a  and  a26122a );
 a26127a <=( a26126a  and  a26119a );
 a26131a <=( A234  and  A232 );
 a26132a <=( A202  and  a26131a );
 a26135a <=( A299  and  A298 );
 a26138a <=( (not A302)  and  A301 );
 a26139a <=( a26138a  and  a26135a );
 a26140a <=( a26139a  and  a26132a );
 a26144a <=( (not A167)  and  A168 );
 a26145a <=( A170  and  a26144a );
 a26148a <=( (not A199)  and  A166 );
 a26151a <=( (not A201)  and  A200 );
 a26152a <=( a26151a  and  a26148a );
 a26153a <=( a26152a  and  a26145a );
 a26157a <=( A234  and  A232 );
 a26158a <=( A202  and  a26157a );
 a26161a <=( (not A299)  and  A298 );
 a26164a <=( A302  and  (not A301) );
 a26165a <=( a26164a  and  a26161a );
 a26166a <=( a26165a  and  a26158a );
 a26170a <=( (not A167)  and  A168 );
 a26171a <=( A170  and  a26170a );
 a26174a <=( (not A199)  and  A166 );
 a26177a <=( (not A201)  and  A200 );
 a26178a <=( a26177a  and  a26174a );
 a26179a <=( a26178a  and  a26171a );
 a26183a <=( A234  and  A232 );
 a26184a <=( A202  and  a26183a );
 a26187a <=( A299  and  (not A298) );
 a26190a <=( A302  and  (not A301) );
 a26191a <=( a26190a  and  a26187a );
 a26192a <=( a26191a  and  a26184a );
 a26196a <=( (not A167)  and  A168 );
 a26197a <=( A170  and  a26196a );
 a26200a <=( (not A199)  and  A166 );
 a26203a <=( (not A201)  and  A200 );
 a26204a <=( a26203a  and  a26200a );
 a26205a <=( a26204a  and  a26197a );
 a26209a <=( A234  and  A232 );
 a26210a <=( A202  and  a26209a );
 a26213a <=( (not A299)  and  (not A298) );
 a26216a <=( (not A302)  and  A301 );
 a26217a <=( a26216a  and  a26213a );
 a26218a <=( a26217a  and  a26210a );
 a26222a <=( (not A167)  and  A168 );
 a26223a <=( A170  and  a26222a );
 a26226a <=( (not A199)  and  A166 );
 a26229a <=( (not A201)  and  A200 );
 a26230a <=( a26229a  and  a26226a );
 a26231a <=( a26230a  and  a26223a );
 a26235a <=( A234  and  A232 );
 a26236a <=( A202  and  a26235a );
 a26239a <=( A266  and  A265 );
 a26242a <=( (not A269)  and  A268 );
 a26243a <=( a26242a  and  a26239a );
 a26244a <=( a26243a  and  a26236a );
 a26248a <=( (not A167)  and  A168 );
 a26249a <=( A170  and  a26248a );
 a26252a <=( (not A199)  and  A166 );
 a26255a <=( (not A201)  and  A200 );
 a26256a <=( a26255a  and  a26252a );
 a26257a <=( a26256a  and  a26249a );
 a26261a <=( A234  and  A232 );
 a26262a <=( A202  and  a26261a );
 a26265a <=( A266  and  (not A265) );
 a26268a <=( A269  and  (not A268) );
 a26269a <=( a26268a  and  a26265a );
 a26270a <=( a26269a  and  a26262a );
 a26274a <=( (not A167)  and  A168 );
 a26275a <=( A170  and  a26274a );
 a26278a <=( (not A199)  and  A166 );
 a26281a <=( (not A201)  and  A200 );
 a26282a <=( a26281a  and  a26278a );
 a26283a <=( a26282a  and  a26275a );
 a26287a <=( A234  and  A232 );
 a26288a <=( A202  and  a26287a );
 a26291a <=( (not A266)  and  A265 );
 a26294a <=( A269  and  (not A268) );
 a26295a <=( a26294a  and  a26291a );
 a26296a <=( a26295a  and  a26288a );
 a26300a <=( (not A167)  and  A168 );
 a26301a <=( A170  and  a26300a );
 a26304a <=( (not A199)  and  A166 );
 a26307a <=( (not A201)  and  A200 );
 a26308a <=( a26307a  and  a26304a );
 a26309a <=( a26308a  and  a26301a );
 a26313a <=( A234  and  A232 );
 a26314a <=( A202  and  a26313a );
 a26317a <=( (not A266)  and  (not A265) );
 a26320a <=( (not A269)  and  A268 );
 a26321a <=( a26320a  and  a26317a );
 a26322a <=( a26321a  and  a26314a );
 a26326a <=( (not A167)  and  A168 );
 a26327a <=( A170  and  a26326a );
 a26330a <=( (not A199)  and  A166 );
 a26333a <=( (not A201)  and  A200 );
 a26334a <=( a26333a  and  a26330a );
 a26335a <=( a26334a  and  a26327a );
 a26339a <=( A234  and  A233 );
 a26340a <=( A202  and  a26339a );
 a26343a <=( A299  and  A298 );
 a26346a <=( (not A302)  and  A301 );
 a26347a <=( a26346a  and  a26343a );
 a26348a <=( a26347a  and  a26340a );
 a26352a <=( (not A167)  and  A168 );
 a26353a <=( A170  and  a26352a );
 a26356a <=( (not A199)  and  A166 );
 a26359a <=( (not A201)  and  A200 );
 a26360a <=( a26359a  and  a26356a );
 a26361a <=( a26360a  and  a26353a );
 a26365a <=( A234  and  A233 );
 a26366a <=( A202  and  a26365a );
 a26369a <=( (not A299)  and  A298 );
 a26372a <=( A302  and  (not A301) );
 a26373a <=( a26372a  and  a26369a );
 a26374a <=( a26373a  and  a26366a );
 a26378a <=( (not A167)  and  A168 );
 a26379a <=( A170  and  a26378a );
 a26382a <=( (not A199)  and  A166 );
 a26385a <=( (not A201)  and  A200 );
 a26386a <=( a26385a  and  a26382a );
 a26387a <=( a26386a  and  a26379a );
 a26391a <=( A234  and  A233 );
 a26392a <=( A202  and  a26391a );
 a26395a <=( A299  and  (not A298) );
 a26398a <=( A302  and  (not A301) );
 a26399a <=( a26398a  and  a26395a );
 a26400a <=( a26399a  and  a26392a );
 a26404a <=( (not A167)  and  A168 );
 a26405a <=( A170  and  a26404a );
 a26408a <=( (not A199)  and  A166 );
 a26411a <=( (not A201)  and  A200 );
 a26412a <=( a26411a  and  a26408a );
 a26413a <=( a26412a  and  a26405a );
 a26417a <=( A234  and  A233 );
 a26418a <=( A202  and  a26417a );
 a26421a <=( (not A299)  and  (not A298) );
 a26424a <=( (not A302)  and  A301 );
 a26425a <=( a26424a  and  a26421a );
 a26426a <=( a26425a  and  a26418a );
 a26430a <=( (not A167)  and  A168 );
 a26431a <=( A170  and  a26430a );
 a26434a <=( (not A199)  and  A166 );
 a26437a <=( (not A201)  and  A200 );
 a26438a <=( a26437a  and  a26434a );
 a26439a <=( a26438a  and  a26431a );
 a26443a <=( A234  and  A233 );
 a26444a <=( A202  and  a26443a );
 a26447a <=( A266  and  A265 );
 a26450a <=( (not A269)  and  A268 );
 a26451a <=( a26450a  and  a26447a );
 a26452a <=( a26451a  and  a26444a );
 a26456a <=( (not A167)  and  A168 );
 a26457a <=( A170  and  a26456a );
 a26460a <=( (not A199)  and  A166 );
 a26463a <=( (not A201)  and  A200 );
 a26464a <=( a26463a  and  a26460a );
 a26465a <=( a26464a  and  a26457a );
 a26469a <=( A234  and  A233 );
 a26470a <=( A202  and  a26469a );
 a26473a <=( A266  and  (not A265) );
 a26476a <=( A269  and  (not A268) );
 a26477a <=( a26476a  and  a26473a );
 a26478a <=( a26477a  and  a26470a );
 a26482a <=( (not A167)  and  A168 );
 a26483a <=( A170  and  a26482a );
 a26486a <=( (not A199)  and  A166 );
 a26489a <=( (not A201)  and  A200 );
 a26490a <=( a26489a  and  a26486a );
 a26491a <=( a26490a  and  a26483a );
 a26495a <=( A234  and  A233 );
 a26496a <=( A202  and  a26495a );
 a26499a <=( (not A266)  and  A265 );
 a26502a <=( A269  and  (not A268) );
 a26503a <=( a26502a  and  a26499a );
 a26504a <=( a26503a  and  a26496a );
 a26508a <=( (not A167)  and  A168 );
 a26509a <=( A170  and  a26508a );
 a26512a <=( (not A199)  and  A166 );
 a26515a <=( (not A201)  and  A200 );
 a26516a <=( a26515a  and  a26512a );
 a26517a <=( a26516a  and  a26509a );
 a26521a <=( A234  and  A233 );
 a26522a <=( A202  and  a26521a );
 a26525a <=( (not A266)  and  (not A265) );
 a26528a <=( (not A269)  and  A268 );
 a26529a <=( a26528a  and  a26525a );
 a26530a <=( a26529a  and  a26522a );
 a26534a <=( (not A167)  and  A168 );
 a26535a <=( A170  and  a26534a );
 a26538a <=( (not A199)  and  A166 );
 a26541a <=( (not A201)  and  A200 );
 a26542a <=( a26541a  and  a26538a );
 a26543a <=( a26542a  and  a26535a );
 a26547a <=( A233  and  A232 );
 a26548a <=( A202  and  a26547a );
 a26551a <=( (not A236)  and  A235 );
 a26554a <=( A300  and  A299 );
 a26555a <=( a26554a  and  a26551a );
 a26556a <=( a26555a  and  a26548a );
 a26560a <=( (not A167)  and  A168 );
 a26561a <=( A170  and  a26560a );
 a26564a <=( (not A199)  and  A166 );
 a26567a <=( (not A201)  and  A200 );
 a26568a <=( a26567a  and  a26564a );
 a26569a <=( a26568a  and  a26561a );
 a26573a <=( A233  and  A232 );
 a26574a <=( A202  and  a26573a );
 a26577a <=( (not A236)  and  A235 );
 a26580a <=( A300  and  A298 );
 a26581a <=( a26580a  and  a26577a );
 a26582a <=( a26581a  and  a26574a );
 a26586a <=( (not A167)  and  A168 );
 a26587a <=( A170  and  a26586a );
 a26590a <=( (not A199)  and  A166 );
 a26593a <=( (not A201)  and  A200 );
 a26594a <=( a26593a  and  a26590a );
 a26595a <=( a26594a  and  a26587a );
 a26599a <=( A233  and  A232 );
 a26600a <=( A202  and  a26599a );
 a26603a <=( (not A236)  and  A235 );
 a26606a <=( A267  and  A265 );
 a26607a <=( a26606a  and  a26603a );
 a26608a <=( a26607a  and  a26600a );
 a26612a <=( (not A167)  and  A168 );
 a26613a <=( A170  and  a26612a );
 a26616a <=( (not A199)  and  A166 );
 a26619a <=( (not A201)  and  A200 );
 a26620a <=( a26619a  and  a26616a );
 a26621a <=( a26620a  and  a26613a );
 a26625a <=( A233  and  A232 );
 a26626a <=( A202  and  a26625a );
 a26629a <=( (not A236)  and  A235 );
 a26632a <=( A267  and  A266 );
 a26633a <=( a26632a  and  a26629a );
 a26634a <=( a26633a  and  a26626a );
 a26638a <=( (not A167)  and  A168 );
 a26639a <=( A170  and  a26638a );
 a26642a <=( (not A199)  and  A166 );
 a26645a <=( (not A201)  and  A200 );
 a26646a <=( a26645a  and  a26642a );
 a26647a <=( a26646a  and  a26639a );
 a26651a <=( A233  and  (not A232) );
 a26652a <=( A202  and  a26651a );
 a26655a <=( A236  and  (not A235) );
 a26658a <=( A300  and  A299 );
 a26659a <=( a26658a  and  a26655a );
 a26660a <=( a26659a  and  a26652a );
 a26664a <=( (not A167)  and  A168 );
 a26665a <=( A170  and  a26664a );
 a26668a <=( (not A199)  and  A166 );
 a26671a <=( (not A201)  and  A200 );
 a26672a <=( a26671a  and  a26668a );
 a26673a <=( a26672a  and  a26665a );
 a26677a <=( A233  and  (not A232) );
 a26678a <=( A202  and  a26677a );
 a26681a <=( A236  and  (not A235) );
 a26684a <=( A300  and  A298 );
 a26685a <=( a26684a  and  a26681a );
 a26686a <=( a26685a  and  a26678a );
 a26690a <=( (not A167)  and  A168 );
 a26691a <=( A170  and  a26690a );
 a26694a <=( (not A199)  and  A166 );
 a26697a <=( (not A201)  and  A200 );
 a26698a <=( a26697a  and  a26694a );
 a26699a <=( a26698a  and  a26691a );
 a26703a <=( A233  and  (not A232) );
 a26704a <=( A202  and  a26703a );
 a26707a <=( A236  and  (not A235) );
 a26710a <=( A267  and  A265 );
 a26711a <=( a26710a  and  a26707a );
 a26712a <=( a26711a  and  a26704a );
 a26716a <=( (not A167)  and  A168 );
 a26717a <=( A170  and  a26716a );
 a26720a <=( (not A199)  and  A166 );
 a26723a <=( (not A201)  and  A200 );
 a26724a <=( a26723a  and  a26720a );
 a26725a <=( a26724a  and  a26717a );
 a26729a <=( A233  and  (not A232) );
 a26730a <=( A202  and  a26729a );
 a26733a <=( A236  and  (not A235) );
 a26736a <=( A267  and  A266 );
 a26737a <=( a26736a  and  a26733a );
 a26738a <=( a26737a  and  a26730a );
 a26742a <=( (not A167)  and  A168 );
 a26743a <=( A170  and  a26742a );
 a26746a <=( (not A199)  and  A166 );
 a26749a <=( (not A201)  and  A200 );
 a26750a <=( a26749a  and  a26746a );
 a26751a <=( a26750a  and  a26743a );
 a26755a <=( (not A233)  and  A232 );
 a26756a <=( A202  and  a26755a );
 a26759a <=( A236  and  (not A235) );
 a26762a <=( A300  and  A299 );
 a26763a <=( a26762a  and  a26759a );
 a26764a <=( a26763a  and  a26756a );
 a26768a <=( (not A167)  and  A168 );
 a26769a <=( A170  and  a26768a );
 a26772a <=( (not A199)  and  A166 );
 a26775a <=( (not A201)  and  A200 );
 a26776a <=( a26775a  and  a26772a );
 a26777a <=( a26776a  and  a26769a );
 a26781a <=( (not A233)  and  A232 );
 a26782a <=( A202  and  a26781a );
 a26785a <=( A236  and  (not A235) );
 a26788a <=( A300  and  A298 );
 a26789a <=( a26788a  and  a26785a );
 a26790a <=( a26789a  and  a26782a );
 a26794a <=( (not A167)  and  A168 );
 a26795a <=( A170  and  a26794a );
 a26798a <=( (not A199)  and  A166 );
 a26801a <=( (not A201)  and  A200 );
 a26802a <=( a26801a  and  a26798a );
 a26803a <=( a26802a  and  a26795a );
 a26807a <=( (not A233)  and  A232 );
 a26808a <=( A202  and  a26807a );
 a26811a <=( A236  and  (not A235) );
 a26814a <=( A267  and  A265 );
 a26815a <=( a26814a  and  a26811a );
 a26816a <=( a26815a  and  a26808a );
 a26820a <=( (not A167)  and  A168 );
 a26821a <=( A170  and  a26820a );
 a26824a <=( (not A199)  and  A166 );
 a26827a <=( (not A201)  and  A200 );
 a26828a <=( a26827a  and  a26824a );
 a26829a <=( a26828a  and  a26821a );
 a26833a <=( (not A233)  and  A232 );
 a26834a <=( A202  and  a26833a );
 a26837a <=( A236  and  (not A235) );
 a26840a <=( A267  and  A266 );
 a26841a <=( a26840a  and  a26837a );
 a26842a <=( a26841a  and  a26834a );
 a26846a <=( (not A167)  and  A168 );
 a26847a <=( A170  and  a26846a );
 a26850a <=( (not A199)  and  A166 );
 a26853a <=( (not A201)  and  A200 );
 a26854a <=( a26853a  and  a26850a );
 a26855a <=( a26854a  and  a26847a );
 a26859a <=( (not A233)  and  (not A232) );
 a26860a <=( A202  and  a26859a );
 a26863a <=( (not A236)  and  A235 );
 a26866a <=( A300  and  A299 );
 a26867a <=( a26866a  and  a26863a );
 a26868a <=( a26867a  and  a26860a );
 a26872a <=( (not A167)  and  A168 );
 a26873a <=( A170  and  a26872a );
 a26876a <=( (not A199)  and  A166 );
 a26879a <=( (not A201)  and  A200 );
 a26880a <=( a26879a  and  a26876a );
 a26881a <=( a26880a  and  a26873a );
 a26885a <=( (not A233)  and  (not A232) );
 a26886a <=( A202  and  a26885a );
 a26889a <=( (not A236)  and  A235 );
 a26892a <=( A300  and  A298 );
 a26893a <=( a26892a  and  a26889a );
 a26894a <=( a26893a  and  a26886a );
 a26898a <=( (not A167)  and  A168 );
 a26899a <=( A170  and  a26898a );
 a26902a <=( (not A199)  and  A166 );
 a26905a <=( (not A201)  and  A200 );
 a26906a <=( a26905a  and  a26902a );
 a26907a <=( a26906a  and  a26899a );
 a26911a <=( (not A233)  and  (not A232) );
 a26912a <=( A202  and  a26911a );
 a26915a <=( (not A236)  and  A235 );
 a26918a <=( A267  and  A265 );
 a26919a <=( a26918a  and  a26915a );
 a26920a <=( a26919a  and  a26912a );
 a26924a <=( (not A167)  and  A168 );
 a26925a <=( A170  and  a26924a );
 a26928a <=( (not A199)  and  A166 );
 a26931a <=( (not A201)  and  A200 );
 a26932a <=( a26931a  and  a26928a );
 a26933a <=( a26932a  and  a26925a );
 a26937a <=( (not A233)  and  (not A232) );
 a26938a <=( A202  and  a26937a );
 a26941a <=( (not A236)  and  A235 );
 a26944a <=( A267  and  A266 );
 a26945a <=( a26944a  and  a26941a );
 a26946a <=( a26945a  and  a26938a );
 a26950a <=( (not A167)  and  A168 );
 a26951a <=( A170  and  a26950a );
 a26954a <=( (not A199)  and  A166 );
 a26957a <=( (not A201)  and  A200 );
 a26958a <=( a26957a  and  a26954a );
 a26959a <=( a26958a  and  a26951a );
 a26963a <=( A234  and  A232 );
 a26964a <=( (not A203)  and  a26963a );
 a26967a <=( A299  and  A298 );
 a26970a <=( (not A302)  and  A301 );
 a26971a <=( a26970a  and  a26967a );
 a26972a <=( a26971a  and  a26964a );
 a26976a <=( (not A167)  and  A168 );
 a26977a <=( A170  and  a26976a );
 a26980a <=( (not A199)  and  A166 );
 a26983a <=( (not A201)  and  A200 );
 a26984a <=( a26983a  and  a26980a );
 a26985a <=( a26984a  and  a26977a );
 a26989a <=( A234  and  A232 );
 a26990a <=( (not A203)  and  a26989a );
 a26993a <=( (not A299)  and  A298 );
 a26996a <=( A302  and  (not A301) );
 a26997a <=( a26996a  and  a26993a );
 a26998a <=( a26997a  and  a26990a );
 a27002a <=( (not A167)  and  A168 );
 a27003a <=( A170  and  a27002a );
 a27006a <=( (not A199)  and  A166 );
 a27009a <=( (not A201)  and  A200 );
 a27010a <=( a27009a  and  a27006a );
 a27011a <=( a27010a  and  a27003a );
 a27015a <=( A234  and  A232 );
 a27016a <=( (not A203)  and  a27015a );
 a27019a <=( A299  and  (not A298) );
 a27022a <=( A302  and  (not A301) );
 a27023a <=( a27022a  and  a27019a );
 a27024a <=( a27023a  and  a27016a );
 a27028a <=( (not A167)  and  A168 );
 a27029a <=( A170  and  a27028a );
 a27032a <=( (not A199)  and  A166 );
 a27035a <=( (not A201)  and  A200 );
 a27036a <=( a27035a  and  a27032a );
 a27037a <=( a27036a  and  a27029a );
 a27041a <=( A234  and  A232 );
 a27042a <=( (not A203)  and  a27041a );
 a27045a <=( (not A299)  and  (not A298) );
 a27048a <=( (not A302)  and  A301 );
 a27049a <=( a27048a  and  a27045a );
 a27050a <=( a27049a  and  a27042a );
 a27054a <=( (not A167)  and  A168 );
 a27055a <=( A170  and  a27054a );
 a27058a <=( (not A199)  and  A166 );
 a27061a <=( (not A201)  and  A200 );
 a27062a <=( a27061a  and  a27058a );
 a27063a <=( a27062a  and  a27055a );
 a27067a <=( A234  and  A232 );
 a27068a <=( (not A203)  and  a27067a );
 a27071a <=( A266  and  A265 );
 a27074a <=( (not A269)  and  A268 );
 a27075a <=( a27074a  and  a27071a );
 a27076a <=( a27075a  and  a27068a );
 a27080a <=( (not A167)  and  A168 );
 a27081a <=( A170  and  a27080a );
 a27084a <=( (not A199)  and  A166 );
 a27087a <=( (not A201)  and  A200 );
 a27088a <=( a27087a  and  a27084a );
 a27089a <=( a27088a  and  a27081a );
 a27093a <=( A234  and  A232 );
 a27094a <=( (not A203)  and  a27093a );
 a27097a <=( A266  and  (not A265) );
 a27100a <=( A269  and  (not A268) );
 a27101a <=( a27100a  and  a27097a );
 a27102a <=( a27101a  and  a27094a );
 a27106a <=( (not A167)  and  A168 );
 a27107a <=( A170  and  a27106a );
 a27110a <=( (not A199)  and  A166 );
 a27113a <=( (not A201)  and  A200 );
 a27114a <=( a27113a  and  a27110a );
 a27115a <=( a27114a  and  a27107a );
 a27119a <=( A234  and  A232 );
 a27120a <=( (not A203)  and  a27119a );
 a27123a <=( (not A266)  and  A265 );
 a27126a <=( A269  and  (not A268) );
 a27127a <=( a27126a  and  a27123a );
 a27128a <=( a27127a  and  a27120a );
 a27132a <=( (not A167)  and  A168 );
 a27133a <=( A170  and  a27132a );
 a27136a <=( (not A199)  and  A166 );
 a27139a <=( (not A201)  and  A200 );
 a27140a <=( a27139a  and  a27136a );
 a27141a <=( a27140a  and  a27133a );
 a27145a <=( A234  and  A232 );
 a27146a <=( (not A203)  and  a27145a );
 a27149a <=( (not A266)  and  (not A265) );
 a27152a <=( (not A269)  and  A268 );
 a27153a <=( a27152a  and  a27149a );
 a27154a <=( a27153a  and  a27146a );
 a27158a <=( (not A167)  and  A168 );
 a27159a <=( A170  and  a27158a );
 a27162a <=( (not A199)  and  A166 );
 a27165a <=( (not A201)  and  A200 );
 a27166a <=( a27165a  and  a27162a );
 a27167a <=( a27166a  and  a27159a );
 a27171a <=( A234  and  A233 );
 a27172a <=( (not A203)  and  a27171a );
 a27175a <=( A299  and  A298 );
 a27178a <=( (not A302)  and  A301 );
 a27179a <=( a27178a  and  a27175a );
 a27180a <=( a27179a  and  a27172a );
 a27184a <=( (not A167)  and  A168 );
 a27185a <=( A170  and  a27184a );
 a27188a <=( (not A199)  and  A166 );
 a27191a <=( (not A201)  and  A200 );
 a27192a <=( a27191a  and  a27188a );
 a27193a <=( a27192a  and  a27185a );
 a27197a <=( A234  and  A233 );
 a27198a <=( (not A203)  and  a27197a );
 a27201a <=( (not A299)  and  A298 );
 a27204a <=( A302  and  (not A301) );
 a27205a <=( a27204a  and  a27201a );
 a27206a <=( a27205a  and  a27198a );
 a27210a <=( (not A167)  and  A168 );
 a27211a <=( A170  and  a27210a );
 a27214a <=( (not A199)  and  A166 );
 a27217a <=( (not A201)  and  A200 );
 a27218a <=( a27217a  and  a27214a );
 a27219a <=( a27218a  and  a27211a );
 a27223a <=( A234  and  A233 );
 a27224a <=( (not A203)  and  a27223a );
 a27227a <=( A299  and  (not A298) );
 a27230a <=( A302  and  (not A301) );
 a27231a <=( a27230a  and  a27227a );
 a27232a <=( a27231a  and  a27224a );
 a27236a <=( (not A167)  and  A168 );
 a27237a <=( A170  and  a27236a );
 a27240a <=( (not A199)  and  A166 );
 a27243a <=( (not A201)  and  A200 );
 a27244a <=( a27243a  and  a27240a );
 a27245a <=( a27244a  and  a27237a );
 a27249a <=( A234  and  A233 );
 a27250a <=( (not A203)  and  a27249a );
 a27253a <=( (not A299)  and  (not A298) );
 a27256a <=( (not A302)  and  A301 );
 a27257a <=( a27256a  and  a27253a );
 a27258a <=( a27257a  and  a27250a );
 a27262a <=( (not A167)  and  A168 );
 a27263a <=( A170  and  a27262a );
 a27266a <=( (not A199)  and  A166 );
 a27269a <=( (not A201)  and  A200 );
 a27270a <=( a27269a  and  a27266a );
 a27271a <=( a27270a  and  a27263a );
 a27275a <=( A234  and  A233 );
 a27276a <=( (not A203)  and  a27275a );
 a27279a <=( A266  and  A265 );
 a27282a <=( (not A269)  and  A268 );
 a27283a <=( a27282a  and  a27279a );
 a27284a <=( a27283a  and  a27276a );
 a27288a <=( (not A167)  and  A168 );
 a27289a <=( A170  and  a27288a );
 a27292a <=( (not A199)  and  A166 );
 a27295a <=( (not A201)  and  A200 );
 a27296a <=( a27295a  and  a27292a );
 a27297a <=( a27296a  and  a27289a );
 a27301a <=( A234  and  A233 );
 a27302a <=( (not A203)  and  a27301a );
 a27305a <=( A266  and  (not A265) );
 a27308a <=( A269  and  (not A268) );
 a27309a <=( a27308a  and  a27305a );
 a27310a <=( a27309a  and  a27302a );
 a27314a <=( (not A167)  and  A168 );
 a27315a <=( A170  and  a27314a );
 a27318a <=( (not A199)  and  A166 );
 a27321a <=( (not A201)  and  A200 );
 a27322a <=( a27321a  and  a27318a );
 a27323a <=( a27322a  and  a27315a );
 a27327a <=( A234  and  A233 );
 a27328a <=( (not A203)  and  a27327a );
 a27331a <=( (not A266)  and  A265 );
 a27334a <=( A269  and  (not A268) );
 a27335a <=( a27334a  and  a27331a );
 a27336a <=( a27335a  and  a27328a );
 a27340a <=( (not A167)  and  A168 );
 a27341a <=( A170  and  a27340a );
 a27344a <=( (not A199)  and  A166 );
 a27347a <=( (not A201)  and  A200 );
 a27348a <=( a27347a  and  a27344a );
 a27349a <=( a27348a  and  a27341a );
 a27353a <=( A234  and  A233 );
 a27354a <=( (not A203)  and  a27353a );
 a27357a <=( (not A266)  and  (not A265) );
 a27360a <=( (not A269)  and  A268 );
 a27361a <=( a27360a  and  a27357a );
 a27362a <=( a27361a  and  a27354a );
 a27366a <=( (not A167)  and  A168 );
 a27367a <=( A170  and  a27366a );
 a27370a <=( (not A199)  and  A166 );
 a27373a <=( (not A201)  and  A200 );
 a27374a <=( a27373a  and  a27370a );
 a27375a <=( a27374a  and  a27367a );
 a27379a <=( A233  and  A232 );
 a27380a <=( (not A203)  and  a27379a );
 a27383a <=( (not A236)  and  A235 );
 a27386a <=( A300  and  A299 );
 a27387a <=( a27386a  and  a27383a );
 a27388a <=( a27387a  and  a27380a );
 a27392a <=( (not A167)  and  A168 );
 a27393a <=( A170  and  a27392a );
 a27396a <=( (not A199)  and  A166 );
 a27399a <=( (not A201)  and  A200 );
 a27400a <=( a27399a  and  a27396a );
 a27401a <=( a27400a  and  a27393a );
 a27405a <=( A233  and  A232 );
 a27406a <=( (not A203)  and  a27405a );
 a27409a <=( (not A236)  and  A235 );
 a27412a <=( A300  and  A298 );
 a27413a <=( a27412a  and  a27409a );
 a27414a <=( a27413a  and  a27406a );
 a27418a <=( (not A167)  and  A168 );
 a27419a <=( A170  and  a27418a );
 a27422a <=( (not A199)  and  A166 );
 a27425a <=( (not A201)  and  A200 );
 a27426a <=( a27425a  and  a27422a );
 a27427a <=( a27426a  and  a27419a );
 a27431a <=( A233  and  A232 );
 a27432a <=( (not A203)  and  a27431a );
 a27435a <=( (not A236)  and  A235 );
 a27438a <=( A267  and  A265 );
 a27439a <=( a27438a  and  a27435a );
 a27440a <=( a27439a  and  a27432a );
 a27444a <=( (not A167)  and  A168 );
 a27445a <=( A170  and  a27444a );
 a27448a <=( (not A199)  and  A166 );
 a27451a <=( (not A201)  and  A200 );
 a27452a <=( a27451a  and  a27448a );
 a27453a <=( a27452a  and  a27445a );
 a27457a <=( A233  and  A232 );
 a27458a <=( (not A203)  and  a27457a );
 a27461a <=( (not A236)  and  A235 );
 a27464a <=( A267  and  A266 );
 a27465a <=( a27464a  and  a27461a );
 a27466a <=( a27465a  and  a27458a );
 a27470a <=( (not A167)  and  A168 );
 a27471a <=( A170  and  a27470a );
 a27474a <=( (not A199)  and  A166 );
 a27477a <=( (not A201)  and  A200 );
 a27478a <=( a27477a  and  a27474a );
 a27479a <=( a27478a  and  a27471a );
 a27483a <=( A233  and  (not A232) );
 a27484a <=( (not A203)  and  a27483a );
 a27487a <=( A236  and  (not A235) );
 a27490a <=( A300  and  A299 );
 a27491a <=( a27490a  and  a27487a );
 a27492a <=( a27491a  and  a27484a );
 a27496a <=( (not A167)  and  A168 );
 a27497a <=( A170  and  a27496a );
 a27500a <=( (not A199)  and  A166 );
 a27503a <=( (not A201)  and  A200 );
 a27504a <=( a27503a  and  a27500a );
 a27505a <=( a27504a  and  a27497a );
 a27509a <=( A233  and  (not A232) );
 a27510a <=( (not A203)  and  a27509a );
 a27513a <=( A236  and  (not A235) );
 a27516a <=( A300  and  A298 );
 a27517a <=( a27516a  and  a27513a );
 a27518a <=( a27517a  and  a27510a );
 a27522a <=( (not A167)  and  A168 );
 a27523a <=( A170  and  a27522a );
 a27526a <=( (not A199)  and  A166 );
 a27529a <=( (not A201)  and  A200 );
 a27530a <=( a27529a  and  a27526a );
 a27531a <=( a27530a  and  a27523a );
 a27535a <=( A233  and  (not A232) );
 a27536a <=( (not A203)  and  a27535a );
 a27539a <=( A236  and  (not A235) );
 a27542a <=( A267  and  A265 );
 a27543a <=( a27542a  and  a27539a );
 a27544a <=( a27543a  and  a27536a );
 a27548a <=( (not A167)  and  A168 );
 a27549a <=( A170  and  a27548a );
 a27552a <=( (not A199)  and  A166 );
 a27555a <=( (not A201)  and  A200 );
 a27556a <=( a27555a  and  a27552a );
 a27557a <=( a27556a  and  a27549a );
 a27561a <=( A233  and  (not A232) );
 a27562a <=( (not A203)  and  a27561a );
 a27565a <=( A236  and  (not A235) );
 a27568a <=( A267  and  A266 );
 a27569a <=( a27568a  and  a27565a );
 a27570a <=( a27569a  and  a27562a );
 a27574a <=( (not A167)  and  A168 );
 a27575a <=( A170  and  a27574a );
 a27578a <=( (not A199)  and  A166 );
 a27581a <=( (not A201)  and  A200 );
 a27582a <=( a27581a  and  a27578a );
 a27583a <=( a27582a  and  a27575a );
 a27587a <=( (not A233)  and  A232 );
 a27588a <=( (not A203)  and  a27587a );
 a27591a <=( A236  and  (not A235) );
 a27594a <=( A300  and  A299 );
 a27595a <=( a27594a  and  a27591a );
 a27596a <=( a27595a  and  a27588a );
 a27600a <=( (not A167)  and  A168 );
 a27601a <=( A170  and  a27600a );
 a27604a <=( (not A199)  and  A166 );
 a27607a <=( (not A201)  and  A200 );
 a27608a <=( a27607a  and  a27604a );
 a27609a <=( a27608a  and  a27601a );
 a27613a <=( (not A233)  and  A232 );
 a27614a <=( (not A203)  and  a27613a );
 a27617a <=( A236  and  (not A235) );
 a27620a <=( A300  and  A298 );
 a27621a <=( a27620a  and  a27617a );
 a27622a <=( a27621a  and  a27614a );
 a27626a <=( (not A167)  and  A168 );
 a27627a <=( A170  and  a27626a );
 a27630a <=( (not A199)  and  A166 );
 a27633a <=( (not A201)  and  A200 );
 a27634a <=( a27633a  and  a27630a );
 a27635a <=( a27634a  and  a27627a );
 a27639a <=( (not A233)  and  A232 );
 a27640a <=( (not A203)  and  a27639a );
 a27643a <=( A236  and  (not A235) );
 a27646a <=( A267  and  A265 );
 a27647a <=( a27646a  and  a27643a );
 a27648a <=( a27647a  and  a27640a );
 a27652a <=( (not A167)  and  A168 );
 a27653a <=( A170  and  a27652a );
 a27656a <=( (not A199)  and  A166 );
 a27659a <=( (not A201)  and  A200 );
 a27660a <=( a27659a  and  a27656a );
 a27661a <=( a27660a  and  a27653a );
 a27665a <=( (not A233)  and  A232 );
 a27666a <=( (not A203)  and  a27665a );
 a27669a <=( A236  and  (not A235) );
 a27672a <=( A267  and  A266 );
 a27673a <=( a27672a  and  a27669a );
 a27674a <=( a27673a  and  a27666a );
 a27678a <=( (not A167)  and  A168 );
 a27679a <=( A170  and  a27678a );
 a27682a <=( (not A199)  and  A166 );
 a27685a <=( (not A201)  and  A200 );
 a27686a <=( a27685a  and  a27682a );
 a27687a <=( a27686a  and  a27679a );
 a27691a <=( (not A233)  and  (not A232) );
 a27692a <=( (not A203)  and  a27691a );
 a27695a <=( (not A236)  and  A235 );
 a27698a <=( A300  and  A299 );
 a27699a <=( a27698a  and  a27695a );
 a27700a <=( a27699a  and  a27692a );
 a27704a <=( (not A167)  and  A168 );
 a27705a <=( A170  and  a27704a );
 a27708a <=( (not A199)  and  A166 );
 a27711a <=( (not A201)  and  A200 );
 a27712a <=( a27711a  and  a27708a );
 a27713a <=( a27712a  and  a27705a );
 a27717a <=( (not A233)  and  (not A232) );
 a27718a <=( (not A203)  and  a27717a );
 a27721a <=( (not A236)  and  A235 );
 a27724a <=( A300  and  A298 );
 a27725a <=( a27724a  and  a27721a );
 a27726a <=( a27725a  and  a27718a );
 a27730a <=( (not A167)  and  A168 );
 a27731a <=( A170  and  a27730a );
 a27734a <=( (not A199)  and  A166 );
 a27737a <=( (not A201)  and  A200 );
 a27738a <=( a27737a  and  a27734a );
 a27739a <=( a27738a  and  a27731a );
 a27743a <=( (not A233)  and  (not A232) );
 a27744a <=( (not A203)  and  a27743a );
 a27747a <=( (not A236)  and  A235 );
 a27750a <=( A267  and  A265 );
 a27751a <=( a27750a  and  a27747a );
 a27752a <=( a27751a  and  a27744a );
 a27756a <=( (not A167)  and  A168 );
 a27757a <=( A170  and  a27756a );
 a27760a <=( (not A199)  and  A166 );
 a27763a <=( (not A201)  and  A200 );
 a27764a <=( a27763a  and  a27760a );
 a27765a <=( a27764a  and  a27757a );
 a27769a <=( (not A233)  and  (not A232) );
 a27770a <=( (not A203)  and  a27769a );
 a27773a <=( (not A236)  and  A235 );
 a27776a <=( A267  and  A266 );
 a27777a <=( a27776a  and  a27773a );
 a27778a <=( a27777a  and  a27770a );
 a27782a <=( (not A167)  and  A168 );
 a27783a <=( A170  and  a27782a );
 a27786a <=( A199  and  A166 );
 a27789a <=( (not A201)  and  (not A200) );
 a27790a <=( a27789a  and  a27786a );
 a27791a <=( a27790a  and  a27783a );
 a27795a <=( A234  and  A232 );
 a27796a <=( A202  and  a27795a );
 a27799a <=( A299  and  A298 );
 a27802a <=( (not A302)  and  A301 );
 a27803a <=( a27802a  and  a27799a );
 a27804a <=( a27803a  and  a27796a );
 a27808a <=( (not A167)  and  A168 );
 a27809a <=( A170  and  a27808a );
 a27812a <=( A199  and  A166 );
 a27815a <=( (not A201)  and  (not A200) );
 a27816a <=( a27815a  and  a27812a );
 a27817a <=( a27816a  and  a27809a );
 a27821a <=( A234  and  A232 );
 a27822a <=( A202  and  a27821a );
 a27825a <=( (not A299)  and  A298 );
 a27828a <=( A302  and  (not A301) );
 a27829a <=( a27828a  and  a27825a );
 a27830a <=( a27829a  and  a27822a );
 a27834a <=( (not A167)  and  A168 );
 a27835a <=( A170  and  a27834a );
 a27838a <=( A199  and  A166 );
 a27841a <=( (not A201)  and  (not A200) );
 a27842a <=( a27841a  and  a27838a );
 a27843a <=( a27842a  and  a27835a );
 a27847a <=( A234  and  A232 );
 a27848a <=( A202  and  a27847a );
 a27851a <=( A299  and  (not A298) );
 a27854a <=( A302  and  (not A301) );
 a27855a <=( a27854a  and  a27851a );
 a27856a <=( a27855a  and  a27848a );
 a27860a <=( (not A167)  and  A168 );
 a27861a <=( A170  and  a27860a );
 a27864a <=( A199  and  A166 );
 a27867a <=( (not A201)  and  (not A200) );
 a27868a <=( a27867a  and  a27864a );
 a27869a <=( a27868a  and  a27861a );
 a27873a <=( A234  and  A232 );
 a27874a <=( A202  and  a27873a );
 a27877a <=( (not A299)  and  (not A298) );
 a27880a <=( (not A302)  and  A301 );
 a27881a <=( a27880a  and  a27877a );
 a27882a <=( a27881a  and  a27874a );
 a27886a <=( (not A167)  and  A168 );
 a27887a <=( A170  and  a27886a );
 a27890a <=( A199  and  A166 );
 a27893a <=( (not A201)  and  (not A200) );
 a27894a <=( a27893a  and  a27890a );
 a27895a <=( a27894a  and  a27887a );
 a27899a <=( A234  and  A232 );
 a27900a <=( A202  and  a27899a );
 a27903a <=( A266  and  A265 );
 a27906a <=( (not A269)  and  A268 );
 a27907a <=( a27906a  and  a27903a );
 a27908a <=( a27907a  and  a27900a );
 a27912a <=( (not A167)  and  A168 );
 a27913a <=( A170  and  a27912a );
 a27916a <=( A199  and  A166 );
 a27919a <=( (not A201)  and  (not A200) );
 a27920a <=( a27919a  and  a27916a );
 a27921a <=( a27920a  and  a27913a );
 a27925a <=( A234  and  A232 );
 a27926a <=( A202  and  a27925a );
 a27929a <=( A266  and  (not A265) );
 a27932a <=( A269  and  (not A268) );
 a27933a <=( a27932a  and  a27929a );
 a27934a <=( a27933a  and  a27926a );
 a27938a <=( (not A167)  and  A168 );
 a27939a <=( A170  and  a27938a );
 a27942a <=( A199  and  A166 );
 a27945a <=( (not A201)  and  (not A200) );
 a27946a <=( a27945a  and  a27942a );
 a27947a <=( a27946a  and  a27939a );
 a27951a <=( A234  and  A232 );
 a27952a <=( A202  and  a27951a );
 a27955a <=( (not A266)  and  A265 );
 a27958a <=( A269  and  (not A268) );
 a27959a <=( a27958a  and  a27955a );
 a27960a <=( a27959a  and  a27952a );
 a27964a <=( (not A167)  and  A168 );
 a27965a <=( A170  and  a27964a );
 a27968a <=( A199  and  A166 );
 a27971a <=( (not A201)  and  (not A200) );
 a27972a <=( a27971a  and  a27968a );
 a27973a <=( a27972a  and  a27965a );
 a27977a <=( A234  and  A232 );
 a27978a <=( A202  and  a27977a );
 a27981a <=( (not A266)  and  (not A265) );
 a27984a <=( (not A269)  and  A268 );
 a27985a <=( a27984a  and  a27981a );
 a27986a <=( a27985a  and  a27978a );
 a27990a <=( (not A167)  and  A168 );
 a27991a <=( A170  and  a27990a );
 a27994a <=( A199  and  A166 );
 a27997a <=( (not A201)  and  (not A200) );
 a27998a <=( a27997a  and  a27994a );
 a27999a <=( a27998a  and  a27991a );
 a28003a <=( A234  and  A233 );
 a28004a <=( A202  and  a28003a );
 a28007a <=( A299  and  A298 );
 a28010a <=( (not A302)  and  A301 );
 a28011a <=( a28010a  and  a28007a );
 a28012a <=( a28011a  and  a28004a );
 a28016a <=( (not A167)  and  A168 );
 a28017a <=( A170  and  a28016a );
 a28020a <=( A199  and  A166 );
 a28023a <=( (not A201)  and  (not A200) );
 a28024a <=( a28023a  and  a28020a );
 a28025a <=( a28024a  and  a28017a );
 a28029a <=( A234  and  A233 );
 a28030a <=( A202  and  a28029a );
 a28033a <=( (not A299)  and  A298 );
 a28036a <=( A302  and  (not A301) );
 a28037a <=( a28036a  and  a28033a );
 a28038a <=( a28037a  and  a28030a );
 a28042a <=( (not A167)  and  A168 );
 a28043a <=( A170  and  a28042a );
 a28046a <=( A199  and  A166 );
 a28049a <=( (not A201)  and  (not A200) );
 a28050a <=( a28049a  and  a28046a );
 a28051a <=( a28050a  and  a28043a );
 a28055a <=( A234  and  A233 );
 a28056a <=( A202  and  a28055a );
 a28059a <=( A299  and  (not A298) );
 a28062a <=( A302  and  (not A301) );
 a28063a <=( a28062a  and  a28059a );
 a28064a <=( a28063a  and  a28056a );
 a28068a <=( (not A167)  and  A168 );
 a28069a <=( A170  and  a28068a );
 a28072a <=( A199  and  A166 );
 a28075a <=( (not A201)  and  (not A200) );
 a28076a <=( a28075a  and  a28072a );
 a28077a <=( a28076a  and  a28069a );
 a28081a <=( A234  and  A233 );
 a28082a <=( A202  and  a28081a );
 a28085a <=( (not A299)  and  (not A298) );
 a28088a <=( (not A302)  and  A301 );
 a28089a <=( a28088a  and  a28085a );
 a28090a <=( a28089a  and  a28082a );
 a28094a <=( (not A167)  and  A168 );
 a28095a <=( A170  and  a28094a );
 a28098a <=( A199  and  A166 );
 a28101a <=( (not A201)  and  (not A200) );
 a28102a <=( a28101a  and  a28098a );
 a28103a <=( a28102a  and  a28095a );
 a28107a <=( A234  and  A233 );
 a28108a <=( A202  and  a28107a );
 a28111a <=( A266  and  A265 );
 a28114a <=( (not A269)  and  A268 );
 a28115a <=( a28114a  and  a28111a );
 a28116a <=( a28115a  and  a28108a );
 a28120a <=( (not A167)  and  A168 );
 a28121a <=( A170  and  a28120a );
 a28124a <=( A199  and  A166 );
 a28127a <=( (not A201)  and  (not A200) );
 a28128a <=( a28127a  and  a28124a );
 a28129a <=( a28128a  and  a28121a );
 a28133a <=( A234  and  A233 );
 a28134a <=( A202  and  a28133a );
 a28137a <=( A266  and  (not A265) );
 a28140a <=( A269  and  (not A268) );
 a28141a <=( a28140a  and  a28137a );
 a28142a <=( a28141a  and  a28134a );
 a28146a <=( (not A167)  and  A168 );
 a28147a <=( A170  and  a28146a );
 a28150a <=( A199  and  A166 );
 a28153a <=( (not A201)  and  (not A200) );
 a28154a <=( a28153a  and  a28150a );
 a28155a <=( a28154a  and  a28147a );
 a28159a <=( A234  and  A233 );
 a28160a <=( A202  and  a28159a );
 a28163a <=( (not A266)  and  A265 );
 a28166a <=( A269  and  (not A268) );
 a28167a <=( a28166a  and  a28163a );
 a28168a <=( a28167a  and  a28160a );
 a28172a <=( (not A167)  and  A168 );
 a28173a <=( A170  and  a28172a );
 a28176a <=( A199  and  A166 );
 a28179a <=( (not A201)  and  (not A200) );
 a28180a <=( a28179a  and  a28176a );
 a28181a <=( a28180a  and  a28173a );
 a28185a <=( A234  and  A233 );
 a28186a <=( A202  and  a28185a );
 a28189a <=( (not A266)  and  (not A265) );
 a28192a <=( (not A269)  and  A268 );
 a28193a <=( a28192a  and  a28189a );
 a28194a <=( a28193a  and  a28186a );
 a28198a <=( (not A167)  and  A168 );
 a28199a <=( A170  and  a28198a );
 a28202a <=( A199  and  A166 );
 a28205a <=( (not A201)  and  (not A200) );
 a28206a <=( a28205a  and  a28202a );
 a28207a <=( a28206a  and  a28199a );
 a28211a <=( A233  and  A232 );
 a28212a <=( A202  and  a28211a );
 a28215a <=( (not A236)  and  A235 );
 a28218a <=( A300  and  A299 );
 a28219a <=( a28218a  and  a28215a );
 a28220a <=( a28219a  and  a28212a );
 a28224a <=( (not A167)  and  A168 );
 a28225a <=( A170  and  a28224a );
 a28228a <=( A199  and  A166 );
 a28231a <=( (not A201)  and  (not A200) );
 a28232a <=( a28231a  and  a28228a );
 a28233a <=( a28232a  and  a28225a );
 a28237a <=( A233  and  A232 );
 a28238a <=( A202  and  a28237a );
 a28241a <=( (not A236)  and  A235 );
 a28244a <=( A300  and  A298 );
 a28245a <=( a28244a  and  a28241a );
 a28246a <=( a28245a  and  a28238a );
 a28250a <=( (not A167)  and  A168 );
 a28251a <=( A170  and  a28250a );
 a28254a <=( A199  and  A166 );
 a28257a <=( (not A201)  and  (not A200) );
 a28258a <=( a28257a  and  a28254a );
 a28259a <=( a28258a  and  a28251a );
 a28263a <=( A233  and  A232 );
 a28264a <=( A202  and  a28263a );
 a28267a <=( (not A236)  and  A235 );
 a28270a <=( A267  and  A265 );
 a28271a <=( a28270a  and  a28267a );
 a28272a <=( a28271a  and  a28264a );
 a28276a <=( (not A167)  and  A168 );
 a28277a <=( A170  and  a28276a );
 a28280a <=( A199  and  A166 );
 a28283a <=( (not A201)  and  (not A200) );
 a28284a <=( a28283a  and  a28280a );
 a28285a <=( a28284a  and  a28277a );
 a28289a <=( A233  and  A232 );
 a28290a <=( A202  and  a28289a );
 a28293a <=( (not A236)  and  A235 );
 a28296a <=( A267  and  A266 );
 a28297a <=( a28296a  and  a28293a );
 a28298a <=( a28297a  and  a28290a );
 a28302a <=( (not A167)  and  A168 );
 a28303a <=( A170  and  a28302a );
 a28306a <=( A199  and  A166 );
 a28309a <=( (not A201)  and  (not A200) );
 a28310a <=( a28309a  and  a28306a );
 a28311a <=( a28310a  and  a28303a );
 a28315a <=( A233  and  (not A232) );
 a28316a <=( A202  and  a28315a );
 a28319a <=( A236  and  (not A235) );
 a28322a <=( A300  and  A299 );
 a28323a <=( a28322a  and  a28319a );
 a28324a <=( a28323a  and  a28316a );
 a28328a <=( (not A167)  and  A168 );
 a28329a <=( A170  and  a28328a );
 a28332a <=( A199  and  A166 );
 a28335a <=( (not A201)  and  (not A200) );
 a28336a <=( a28335a  and  a28332a );
 a28337a <=( a28336a  and  a28329a );
 a28341a <=( A233  and  (not A232) );
 a28342a <=( A202  and  a28341a );
 a28345a <=( A236  and  (not A235) );
 a28348a <=( A300  and  A298 );
 a28349a <=( a28348a  and  a28345a );
 a28350a <=( a28349a  and  a28342a );
 a28354a <=( (not A167)  and  A168 );
 a28355a <=( A170  and  a28354a );
 a28358a <=( A199  and  A166 );
 a28361a <=( (not A201)  and  (not A200) );
 a28362a <=( a28361a  and  a28358a );
 a28363a <=( a28362a  and  a28355a );
 a28367a <=( A233  and  (not A232) );
 a28368a <=( A202  and  a28367a );
 a28371a <=( A236  and  (not A235) );
 a28374a <=( A267  and  A265 );
 a28375a <=( a28374a  and  a28371a );
 a28376a <=( a28375a  and  a28368a );
 a28380a <=( (not A167)  and  A168 );
 a28381a <=( A170  and  a28380a );
 a28384a <=( A199  and  A166 );
 a28387a <=( (not A201)  and  (not A200) );
 a28388a <=( a28387a  and  a28384a );
 a28389a <=( a28388a  and  a28381a );
 a28393a <=( A233  and  (not A232) );
 a28394a <=( A202  and  a28393a );
 a28397a <=( A236  and  (not A235) );
 a28400a <=( A267  and  A266 );
 a28401a <=( a28400a  and  a28397a );
 a28402a <=( a28401a  and  a28394a );
 a28406a <=( (not A167)  and  A168 );
 a28407a <=( A170  and  a28406a );
 a28410a <=( A199  and  A166 );
 a28413a <=( (not A201)  and  (not A200) );
 a28414a <=( a28413a  and  a28410a );
 a28415a <=( a28414a  and  a28407a );
 a28419a <=( (not A233)  and  A232 );
 a28420a <=( A202  and  a28419a );
 a28423a <=( A236  and  (not A235) );
 a28426a <=( A300  and  A299 );
 a28427a <=( a28426a  and  a28423a );
 a28428a <=( a28427a  and  a28420a );
 a28432a <=( (not A167)  and  A168 );
 a28433a <=( A170  and  a28432a );
 a28436a <=( A199  and  A166 );
 a28439a <=( (not A201)  and  (not A200) );
 a28440a <=( a28439a  and  a28436a );
 a28441a <=( a28440a  and  a28433a );
 a28445a <=( (not A233)  and  A232 );
 a28446a <=( A202  and  a28445a );
 a28449a <=( A236  and  (not A235) );
 a28452a <=( A300  and  A298 );
 a28453a <=( a28452a  and  a28449a );
 a28454a <=( a28453a  and  a28446a );
 a28458a <=( (not A167)  and  A168 );
 a28459a <=( A170  and  a28458a );
 a28462a <=( A199  and  A166 );
 a28465a <=( (not A201)  and  (not A200) );
 a28466a <=( a28465a  and  a28462a );
 a28467a <=( a28466a  and  a28459a );
 a28471a <=( (not A233)  and  A232 );
 a28472a <=( A202  and  a28471a );
 a28475a <=( A236  and  (not A235) );
 a28478a <=( A267  and  A265 );
 a28479a <=( a28478a  and  a28475a );
 a28480a <=( a28479a  and  a28472a );
 a28484a <=( (not A167)  and  A168 );
 a28485a <=( A170  and  a28484a );
 a28488a <=( A199  and  A166 );
 a28491a <=( (not A201)  and  (not A200) );
 a28492a <=( a28491a  and  a28488a );
 a28493a <=( a28492a  and  a28485a );
 a28497a <=( (not A233)  and  A232 );
 a28498a <=( A202  and  a28497a );
 a28501a <=( A236  and  (not A235) );
 a28504a <=( A267  and  A266 );
 a28505a <=( a28504a  and  a28501a );
 a28506a <=( a28505a  and  a28498a );
 a28510a <=( (not A167)  and  A168 );
 a28511a <=( A170  and  a28510a );
 a28514a <=( A199  and  A166 );
 a28517a <=( (not A201)  and  (not A200) );
 a28518a <=( a28517a  and  a28514a );
 a28519a <=( a28518a  and  a28511a );
 a28523a <=( (not A233)  and  (not A232) );
 a28524a <=( A202  and  a28523a );
 a28527a <=( (not A236)  and  A235 );
 a28530a <=( A300  and  A299 );
 a28531a <=( a28530a  and  a28527a );
 a28532a <=( a28531a  and  a28524a );
 a28536a <=( (not A167)  and  A168 );
 a28537a <=( A170  and  a28536a );
 a28540a <=( A199  and  A166 );
 a28543a <=( (not A201)  and  (not A200) );
 a28544a <=( a28543a  and  a28540a );
 a28545a <=( a28544a  and  a28537a );
 a28549a <=( (not A233)  and  (not A232) );
 a28550a <=( A202  and  a28549a );
 a28553a <=( (not A236)  and  A235 );
 a28556a <=( A300  and  A298 );
 a28557a <=( a28556a  and  a28553a );
 a28558a <=( a28557a  and  a28550a );
 a28562a <=( (not A167)  and  A168 );
 a28563a <=( A170  and  a28562a );
 a28566a <=( A199  and  A166 );
 a28569a <=( (not A201)  and  (not A200) );
 a28570a <=( a28569a  and  a28566a );
 a28571a <=( a28570a  and  a28563a );
 a28575a <=( (not A233)  and  (not A232) );
 a28576a <=( A202  and  a28575a );
 a28579a <=( (not A236)  and  A235 );
 a28582a <=( A267  and  A265 );
 a28583a <=( a28582a  and  a28579a );
 a28584a <=( a28583a  and  a28576a );
 a28588a <=( (not A167)  and  A168 );
 a28589a <=( A170  and  a28588a );
 a28592a <=( A199  and  A166 );
 a28595a <=( (not A201)  and  (not A200) );
 a28596a <=( a28595a  and  a28592a );
 a28597a <=( a28596a  and  a28589a );
 a28601a <=( (not A233)  and  (not A232) );
 a28602a <=( A202  and  a28601a );
 a28605a <=( (not A236)  and  A235 );
 a28608a <=( A267  and  A266 );
 a28609a <=( a28608a  and  a28605a );
 a28610a <=( a28609a  and  a28602a );
 a28614a <=( (not A167)  and  A168 );
 a28615a <=( A170  and  a28614a );
 a28618a <=( A199  and  A166 );
 a28621a <=( (not A201)  and  (not A200) );
 a28622a <=( a28621a  and  a28618a );
 a28623a <=( a28622a  and  a28615a );
 a28627a <=( A234  and  A232 );
 a28628a <=( (not A203)  and  a28627a );
 a28631a <=( A299  and  A298 );
 a28634a <=( (not A302)  and  A301 );
 a28635a <=( a28634a  and  a28631a );
 a28636a <=( a28635a  and  a28628a );
 a28640a <=( (not A167)  and  A168 );
 a28641a <=( A170  and  a28640a );
 a28644a <=( A199  and  A166 );
 a28647a <=( (not A201)  and  (not A200) );
 a28648a <=( a28647a  and  a28644a );
 a28649a <=( a28648a  and  a28641a );
 a28653a <=( A234  and  A232 );
 a28654a <=( (not A203)  and  a28653a );
 a28657a <=( (not A299)  and  A298 );
 a28660a <=( A302  and  (not A301) );
 a28661a <=( a28660a  and  a28657a );
 a28662a <=( a28661a  and  a28654a );
 a28666a <=( (not A167)  and  A168 );
 a28667a <=( A170  and  a28666a );
 a28670a <=( A199  and  A166 );
 a28673a <=( (not A201)  and  (not A200) );
 a28674a <=( a28673a  and  a28670a );
 a28675a <=( a28674a  and  a28667a );
 a28679a <=( A234  and  A232 );
 a28680a <=( (not A203)  and  a28679a );
 a28683a <=( A299  and  (not A298) );
 a28686a <=( A302  and  (not A301) );
 a28687a <=( a28686a  and  a28683a );
 a28688a <=( a28687a  and  a28680a );
 a28692a <=( (not A167)  and  A168 );
 a28693a <=( A170  and  a28692a );
 a28696a <=( A199  and  A166 );
 a28699a <=( (not A201)  and  (not A200) );
 a28700a <=( a28699a  and  a28696a );
 a28701a <=( a28700a  and  a28693a );
 a28705a <=( A234  and  A232 );
 a28706a <=( (not A203)  and  a28705a );
 a28709a <=( (not A299)  and  (not A298) );
 a28712a <=( (not A302)  and  A301 );
 a28713a <=( a28712a  and  a28709a );
 a28714a <=( a28713a  and  a28706a );
 a28718a <=( (not A167)  and  A168 );
 a28719a <=( A170  and  a28718a );
 a28722a <=( A199  and  A166 );
 a28725a <=( (not A201)  and  (not A200) );
 a28726a <=( a28725a  and  a28722a );
 a28727a <=( a28726a  and  a28719a );
 a28731a <=( A234  and  A232 );
 a28732a <=( (not A203)  and  a28731a );
 a28735a <=( A266  and  A265 );
 a28738a <=( (not A269)  and  A268 );
 a28739a <=( a28738a  and  a28735a );
 a28740a <=( a28739a  and  a28732a );
 a28744a <=( (not A167)  and  A168 );
 a28745a <=( A170  and  a28744a );
 a28748a <=( A199  and  A166 );
 a28751a <=( (not A201)  and  (not A200) );
 a28752a <=( a28751a  and  a28748a );
 a28753a <=( a28752a  and  a28745a );
 a28757a <=( A234  and  A232 );
 a28758a <=( (not A203)  and  a28757a );
 a28761a <=( A266  and  (not A265) );
 a28764a <=( A269  and  (not A268) );
 a28765a <=( a28764a  and  a28761a );
 a28766a <=( a28765a  and  a28758a );
 a28770a <=( (not A167)  and  A168 );
 a28771a <=( A170  and  a28770a );
 a28774a <=( A199  and  A166 );
 a28777a <=( (not A201)  and  (not A200) );
 a28778a <=( a28777a  and  a28774a );
 a28779a <=( a28778a  and  a28771a );
 a28783a <=( A234  and  A232 );
 a28784a <=( (not A203)  and  a28783a );
 a28787a <=( (not A266)  and  A265 );
 a28790a <=( A269  and  (not A268) );
 a28791a <=( a28790a  and  a28787a );
 a28792a <=( a28791a  and  a28784a );
 a28796a <=( (not A167)  and  A168 );
 a28797a <=( A170  and  a28796a );
 a28800a <=( A199  and  A166 );
 a28803a <=( (not A201)  and  (not A200) );
 a28804a <=( a28803a  and  a28800a );
 a28805a <=( a28804a  and  a28797a );
 a28809a <=( A234  and  A232 );
 a28810a <=( (not A203)  and  a28809a );
 a28813a <=( (not A266)  and  (not A265) );
 a28816a <=( (not A269)  and  A268 );
 a28817a <=( a28816a  and  a28813a );
 a28818a <=( a28817a  and  a28810a );
 a28822a <=( (not A167)  and  A168 );
 a28823a <=( A170  and  a28822a );
 a28826a <=( A199  and  A166 );
 a28829a <=( (not A201)  and  (not A200) );
 a28830a <=( a28829a  and  a28826a );
 a28831a <=( a28830a  and  a28823a );
 a28835a <=( A234  and  A233 );
 a28836a <=( (not A203)  and  a28835a );
 a28839a <=( A299  and  A298 );
 a28842a <=( (not A302)  and  A301 );
 a28843a <=( a28842a  and  a28839a );
 a28844a <=( a28843a  and  a28836a );
 a28848a <=( (not A167)  and  A168 );
 a28849a <=( A170  and  a28848a );
 a28852a <=( A199  and  A166 );
 a28855a <=( (not A201)  and  (not A200) );
 a28856a <=( a28855a  and  a28852a );
 a28857a <=( a28856a  and  a28849a );
 a28861a <=( A234  and  A233 );
 a28862a <=( (not A203)  and  a28861a );
 a28865a <=( (not A299)  and  A298 );
 a28868a <=( A302  and  (not A301) );
 a28869a <=( a28868a  and  a28865a );
 a28870a <=( a28869a  and  a28862a );
 a28874a <=( (not A167)  and  A168 );
 a28875a <=( A170  and  a28874a );
 a28878a <=( A199  and  A166 );
 a28881a <=( (not A201)  and  (not A200) );
 a28882a <=( a28881a  and  a28878a );
 a28883a <=( a28882a  and  a28875a );
 a28887a <=( A234  and  A233 );
 a28888a <=( (not A203)  and  a28887a );
 a28891a <=( A299  and  (not A298) );
 a28894a <=( A302  and  (not A301) );
 a28895a <=( a28894a  and  a28891a );
 a28896a <=( a28895a  and  a28888a );
 a28900a <=( (not A167)  and  A168 );
 a28901a <=( A170  and  a28900a );
 a28904a <=( A199  and  A166 );
 a28907a <=( (not A201)  and  (not A200) );
 a28908a <=( a28907a  and  a28904a );
 a28909a <=( a28908a  and  a28901a );
 a28913a <=( A234  and  A233 );
 a28914a <=( (not A203)  and  a28913a );
 a28917a <=( (not A299)  and  (not A298) );
 a28920a <=( (not A302)  and  A301 );
 a28921a <=( a28920a  and  a28917a );
 a28922a <=( a28921a  and  a28914a );
 a28926a <=( (not A167)  and  A168 );
 a28927a <=( A170  and  a28926a );
 a28930a <=( A199  and  A166 );
 a28933a <=( (not A201)  and  (not A200) );
 a28934a <=( a28933a  and  a28930a );
 a28935a <=( a28934a  and  a28927a );
 a28939a <=( A234  and  A233 );
 a28940a <=( (not A203)  and  a28939a );
 a28943a <=( A266  and  A265 );
 a28946a <=( (not A269)  and  A268 );
 a28947a <=( a28946a  and  a28943a );
 a28948a <=( a28947a  and  a28940a );
 a28952a <=( (not A167)  and  A168 );
 a28953a <=( A170  and  a28952a );
 a28956a <=( A199  and  A166 );
 a28959a <=( (not A201)  and  (not A200) );
 a28960a <=( a28959a  and  a28956a );
 a28961a <=( a28960a  and  a28953a );
 a28965a <=( A234  and  A233 );
 a28966a <=( (not A203)  and  a28965a );
 a28969a <=( A266  and  (not A265) );
 a28972a <=( A269  and  (not A268) );
 a28973a <=( a28972a  and  a28969a );
 a28974a <=( a28973a  and  a28966a );
 a28978a <=( (not A167)  and  A168 );
 a28979a <=( A170  and  a28978a );
 a28982a <=( A199  and  A166 );
 a28985a <=( (not A201)  and  (not A200) );
 a28986a <=( a28985a  and  a28982a );
 a28987a <=( a28986a  and  a28979a );
 a28991a <=( A234  and  A233 );
 a28992a <=( (not A203)  and  a28991a );
 a28995a <=( (not A266)  and  A265 );
 a28998a <=( A269  and  (not A268) );
 a28999a <=( a28998a  and  a28995a );
 a29000a <=( a28999a  and  a28992a );
 a29004a <=( (not A167)  and  A168 );
 a29005a <=( A170  and  a29004a );
 a29008a <=( A199  and  A166 );
 a29011a <=( (not A201)  and  (not A200) );
 a29012a <=( a29011a  and  a29008a );
 a29013a <=( a29012a  and  a29005a );
 a29017a <=( A234  and  A233 );
 a29018a <=( (not A203)  and  a29017a );
 a29021a <=( (not A266)  and  (not A265) );
 a29024a <=( (not A269)  and  A268 );
 a29025a <=( a29024a  and  a29021a );
 a29026a <=( a29025a  and  a29018a );
 a29030a <=( (not A167)  and  A168 );
 a29031a <=( A170  and  a29030a );
 a29034a <=( A199  and  A166 );
 a29037a <=( (not A201)  and  (not A200) );
 a29038a <=( a29037a  and  a29034a );
 a29039a <=( a29038a  and  a29031a );
 a29043a <=( A233  and  A232 );
 a29044a <=( (not A203)  and  a29043a );
 a29047a <=( (not A236)  and  A235 );
 a29050a <=( A300  and  A299 );
 a29051a <=( a29050a  and  a29047a );
 a29052a <=( a29051a  and  a29044a );
 a29056a <=( (not A167)  and  A168 );
 a29057a <=( A170  and  a29056a );
 a29060a <=( A199  and  A166 );
 a29063a <=( (not A201)  and  (not A200) );
 a29064a <=( a29063a  and  a29060a );
 a29065a <=( a29064a  and  a29057a );
 a29069a <=( A233  and  A232 );
 a29070a <=( (not A203)  and  a29069a );
 a29073a <=( (not A236)  and  A235 );
 a29076a <=( A300  and  A298 );
 a29077a <=( a29076a  and  a29073a );
 a29078a <=( a29077a  and  a29070a );
 a29082a <=( (not A167)  and  A168 );
 a29083a <=( A170  and  a29082a );
 a29086a <=( A199  and  A166 );
 a29089a <=( (not A201)  and  (not A200) );
 a29090a <=( a29089a  and  a29086a );
 a29091a <=( a29090a  and  a29083a );
 a29095a <=( A233  and  A232 );
 a29096a <=( (not A203)  and  a29095a );
 a29099a <=( (not A236)  and  A235 );
 a29102a <=( A267  and  A265 );
 a29103a <=( a29102a  and  a29099a );
 a29104a <=( a29103a  and  a29096a );
 a29108a <=( (not A167)  and  A168 );
 a29109a <=( A170  and  a29108a );
 a29112a <=( A199  and  A166 );
 a29115a <=( (not A201)  and  (not A200) );
 a29116a <=( a29115a  and  a29112a );
 a29117a <=( a29116a  and  a29109a );
 a29121a <=( A233  and  A232 );
 a29122a <=( (not A203)  and  a29121a );
 a29125a <=( (not A236)  and  A235 );
 a29128a <=( A267  and  A266 );
 a29129a <=( a29128a  and  a29125a );
 a29130a <=( a29129a  and  a29122a );
 a29134a <=( (not A167)  and  A168 );
 a29135a <=( A170  and  a29134a );
 a29138a <=( A199  and  A166 );
 a29141a <=( (not A201)  and  (not A200) );
 a29142a <=( a29141a  and  a29138a );
 a29143a <=( a29142a  and  a29135a );
 a29147a <=( A233  and  (not A232) );
 a29148a <=( (not A203)  and  a29147a );
 a29151a <=( A236  and  (not A235) );
 a29154a <=( A300  and  A299 );
 a29155a <=( a29154a  and  a29151a );
 a29156a <=( a29155a  and  a29148a );
 a29160a <=( (not A167)  and  A168 );
 a29161a <=( A170  and  a29160a );
 a29164a <=( A199  and  A166 );
 a29167a <=( (not A201)  and  (not A200) );
 a29168a <=( a29167a  and  a29164a );
 a29169a <=( a29168a  and  a29161a );
 a29173a <=( A233  and  (not A232) );
 a29174a <=( (not A203)  and  a29173a );
 a29177a <=( A236  and  (not A235) );
 a29180a <=( A300  and  A298 );
 a29181a <=( a29180a  and  a29177a );
 a29182a <=( a29181a  and  a29174a );
 a29186a <=( (not A167)  and  A168 );
 a29187a <=( A170  and  a29186a );
 a29190a <=( A199  and  A166 );
 a29193a <=( (not A201)  and  (not A200) );
 a29194a <=( a29193a  and  a29190a );
 a29195a <=( a29194a  and  a29187a );
 a29199a <=( A233  and  (not A232) );
 a29200a <=( (not A203)  and  a29199a );
 a29203a <=( A236  and  (not A235) );
 a29206a <=( A267  and  A265 );
 a29207a <=( a29206a  and  a29203a );
 a29208a <=( a29207a  and  a29200a );
 a29212a <=( (not A167)  and  A168 );
 a29213a <=( A170  and  a29212a );
 a29216a <=( A199  and  A166 );
 a29219a <=( (not A201)  and  (not A200) );
 a29220a <=( a29219a  and  a29216a );
 a29221a <=( a29220a  and  a29213a );
 a29225a <=( A233  and  (not A232) );
 a29226a <=( (not A203)  and  a29225a );
 a29229a <=( A236  and  (not A235) );
 a29232a <=( A267  and  A266 );
 a29233a <=( a29232a  and  a29229a );
 a29234a <=( a29233a  and  a29226a );
 a29238a <=( (not A167)  and  A168 );
 a29239a <=( A170  and  a29238a );
 a29242a <=( A199  and  A166 );
 a29245a <=( (not A201)  and  (not A200) );
 a29246a <=( a29245a  and  a29242a );
 a29247a <=( a29246a  and  a29239a );
 a29251a <=( (not A233)  and  A232 );
 a29252a <=( (not A203)  and  a29251a );
 a29255a <=( A236  and  (not A235) );
 a29258a <=( A300  and  A299 );
 a29259a <=( a29258a  and  a29255a );
 a29260a <=( a29259a  and  a29252a );
 a29264a <=( (not A167)  and  A168 );
 a29265a <=( A170  and  a29264a );
 a29268a <=( A199  and  A166 );
 a29271a <=( (not A201)  and  (not A200) );
 a29272a <=( a29271a  and  a29268a );
 a29273a <=( a29272a  and  a29265a );
 a29277a <=( (not A233)  and  A232 );
 a29278a <=( (not A203)  and  a29277a );
 a29281a <=( A236  and  (not A235) );
 a29284a <=( A300  and  A298 );
 a29285a <=( a29284a  and  a29281a );
 a29286a <=( a29285a  and  a29278a );
 a29290a <=( (not A167)  and  A168 );
 a29291a <=( A170  and  a29290a );
 a29294a <=( A199  and  A166 );
 a29297a <=( (not A201)  and  (not A200) );
 a29298a <=( a29297a  and  a29294a );
 a29299a <=( a29298a  and  a29291a );
 a29303a <=( (not A233)  and  A232 );
 a29304a <=( (not A203)  and  a29303a );
 a29307a <=( A236  and  (not A235) );
 a29310a <=( A267  and  A265 );
 a29311a <=( a29310a  and  a29307a );
 a29312a <=( a29311a  and  a29304a );
 a29316a <=( (not A167)  and  A168 );
 a29317a <=( A170  and  a29316a );
 a29320a <=( A199  and  A166 );
 a29323a <=( (not A201)  and  (not A200) );
 a29324a <=( a29323a  and  a29320a );
 a29325a <=( a29324a  and  a29317a );
 a29329a <=( (not A233)  and  A232 );
 a29330a <=( (not A203)  and  a29329a );
 a29333a <=( A236  and  (not A235) );
 a29336a <=( A267  and  A266 );
 a29337a <=( a29336a  and  a29333a );
 a29338a <=( a29337a  and  a29330a );
 a29342a <=( (not A167)  and  A168 );
 a29343a <=( A170  and  a29342a );
 a29346a <=( A199  and  A166 );
 a29349a <=( (not A201)  and  (not A200) );
 a29350a <=( a29349a  and  a29346a );
 a29351a <=( a29350a  and  a29343a );
 a29355a <=( (not A233)  and  (not A232) );
 a29356a <=( (not A203)  and  a29355a );
 a29359a <=( (not A236)  and  A235 );
 a29362a <=( A300  and  A299 );
 a29363a <=( a29362a  and  a29359a );
 a29364a <=( a29363a  and  a29356a );
 a29368a <=( (not A167)  and  A168 );
 a29369a <=( A170  and  a29368a );
 a29372a <=( A199  and  A166 );
 a29375a <=( (not A201)  and  (not A200) );
 a29376a <=( a29375a  and  a29372a );
 a29377a <=( a29376a  and  a29369a );
 a29381a <=( (not A233)  and  (not A232) );
 a29382a <=( (not A203)  and  a29381a );
 a29385a <=( (not A236)  and  A235 );
 a29388a <=( A300  and  A298 );
 a29389a <=( a29388a  and  a29385a );
 a29390a <=( a29389a  and  a29382a );
 a29394a <=( (not A167)  and  A168 );
 a29395a <=( A170  and  a29394a );
 a29398a <=( A199  and  A166 );
 a29401a <=( (not A201)  and  (not A200) );
 a29402a <=( a29401a  and  a29398a );
 a29403a <=( a29402a  and  a29395a );
 a29407a <=( (not A233)  and  (not A232) );
 a29408a <=( (not A203)  and  a29407a );
 a29411a <=( (not A236)  and  A235 );
 a29414a <=( A267  and  A265 );
 a29415a <=( a29414a  and  a29411a );
 a29416a <=( a29415a  and  a29408a );
 a29420a <=( (not A167)  and  A168 );
 a29421a <=( A170  and  a29420a );
 a29424a <=( A199  and  A166 );
 a29427a <=( (not A201)  and  (not A200) );
 a29428a <=( a29427a  and  a29424a );
 a29429a <=( a29428a  and  a29421a );
 a29433a <=( (not A233)  and  (not A232) );
 a29434a <=( (not A203)  and  a29433a );
 a29437a <=( (not A236)  and  A235 );
 a29440a <=( A267  and  A266 );
 a29441a <=( a29440a  and  a29437a );
 a29442a <=( a29441a  and  a29434a );
 a29446a <=( (not A167)  and  A168 );
 a29447a <=( A169  and  a29446a );
 a29450a <=( A199  and  A166 );
 a29453a <=( (not A201)  and  A200 );
 a29454a <=( a29453a  and  a29450a );
 a29455a <=( a29454a  and  a29447a );
 a29459a <=( A234  and  A232 );
 a29460a <=( (not A202)  and  a29459a );
 a29463a <=( A299  and  A298 );
 a29466a <=( (not A302)  and  A301 );
 a29467a <=( a29466a  and  a29463a );
 a29468a <=( a29467a  and  a29460a );
 a29472a <=( (not A167)  and  A168 );
 a29473a <=( A169  and  a29472a );
 a29476a <=( A199  and  A166 );
 a29479a <=( (not A201)  and  A200 );
 a29480a <=( a29479a  and  a29476a );
 a29481a <=( a29480a  and  a29473a );
 a29485a <=( A234  and  A232 );
 a29486a <=( (not A202)  and  a29485a );
 a29489a <=( (not A299)  and  A298 );
 a29492a <=( A302  and  (not A301) );
 a29493a <=( a29492a  and  a29489a );
 a29494a <=( a29493a  and  a29486a );
 a29498a <=( (not A167)  and  A168 );
 a29499a <=( A169  and  a29498a );
 a29502a <=( A199  and  A166 );
 a29505a <=( (not A201)  and  A200 );
 a29506a <=( a29505a  and  a29502a );
 a29507a <=( a29506a  and  a29499a );
 a29511a <=( A234  and  A232 );
 a29512a <=( (not A202)  and  a29511a );
 a29515a <=( A299  and  (not A298) );
 a29518a <=( A302  and  (not A301) );
 a29519a <=( a29518a  and  a29515a );
 a29520a <=( a29519a  and  a29512a );
 a29524a <=( (not A167)  and  A168 );
 a29525a <=( A169  and  a29524a );
 a29528a <=( A199  and  A166 );
 a29531a <=( (not A201)  and  A200 );
 a29532a <=( a29531a  and  a29528a );
 a29533a <=( a29532a  and  a29525a );
 a29537a <=( A234  and  A232 );
 a29538a <=( (not A202)  and  a29537a );
 a29541a <=( (not A299)  and  (not A298) );
 a29544a <=( (not A302)  and  A301 );
 a29545a <=( a29544a  and  a29541a );
 a29546a <=( a29545a  and  a29538a );
 a29550a <=( (not A167)  and  A168 );
 a29551a <=( A169  and  a29550a );
 a29554a <=( A199  and  A166 );
 a29557a <=( (not A201)  and  A200 );
 a29558a <=( a29557a  and  a29554a );
 a29559a <=( a29558a  and  a29551a );
 a29563a <=( A234  and  A232 );
 a29564a <=( (not A202)  and  a29563a );
 a29567a <=( A266  and  A265 );
 a29570a <=( (not A269)  and  A268 );
 a29571a <=( a29570a  and  a29567a );
 a29572a <=( a29571a  and  a29564a );
 a29576a <=( (not A167)  and  A168 );
 a29577a <=( A169  and  a29576a );
 a29580a <=( A199  and  A166 );
 a29583a <=( (not A201)  and  A200 );
 a29584a <=( a29583a  and  a29580a );
 a29585a <=( a29584a  and  a29577a );
 a29589a <=( A234  and  A232 );
 a29590a <=( (not A202)  and  a29589a );
 a29593a <=( A266  and  (not A265) );
 a29596a <=( A269  and  (not A268) );
 a29597a <=( a29596a  and  a29593a );
 a29598a <=( a29597a  and  a29590a );
 a29602a <=( (not A167)  and  A168 );
 a29603a <=( A169  and  a29602a );
 a29606a <=( A199  and  A166 );
 a29609a <=( (not A201)  and  A200 );
 a29610a <=( a29609a  and  a29606a );
 a29611a <=( a29610a  and  a29603a );
 a29615a <=( A234  and  A232 );
 a29616a <=( (not A202)  and  a29615a );
 a29619a <=( (not A266)  and  A265 );
 a29622a <=( A269  and  (not A268) );
 a29623a <=( a29622a  and  a29619a );
 a29624a <=( a29623a  and  a29616a );
 a29628a <=( (not A167)  and  A168 );
 a29629a <=( A169  and  a29628a );
 a29632a <=( A199  and  A166 );
 a29635a <=( (not A201)  and  A200 );
 a29636a <=( a29635a  and  a29632a );
 a29637a <=( a29636a  and  a29629a );
 a29641a <=( A234  and  A232 );
 a29642a <=( (not A202)  and  a29641a );
 a29645a <=( (not A266)  and  (not A265) );
 a29648a <=( (not A269)  and  A268 );
 a29649a <=( a29648a  and  a29645a );
 a29650a <=( a29649a  and  a29642a );
 a29654a <=( (not A167)  and  A168 );
 a29655a <=( A169  and  a29654a );
 a29658a <=( A199  and  A166 );
 a29661a <=( (not A201)  and  A200 );
 a29662a <=( a29661a  and  a29658a );
 a29663a <=( a29662a  and  a29655a );
 a29667a <=( A234  and  A233 );
 a29668a <=( (not A202)  and  a29667a );
 a29671a <=( A299  and  A298 );
 a29674a <=( (not A302)  and  A301 );
 a29675a <=( a29674a  and  a29671a );
 a29676a <=( a29675a  and  a29668a );
 a29680a <=( (not A167)  and  A168 );
 a29681a <=( A169  and  a29680a );
 a29684a <=( A199  and  A166 );
 a29687a <=( (not A201)  and  A200 );
 a29688a <=( a29687a  and  a29684a );
 a29689a <=( a29688a  and  a29681a );
 a29693a <=( A234  and  A233 );
 a29694a <=( (not A202)  and  a29693a );
 a29697a <=( (not A299)  and  A298 );
 a29700a <=( A302  and  (not A301) );
 a29701a <=( a29700a  and  a29697a );
 a29702a <=( a29701a  and  a29694a );
 a29706a <=( (not A167)  and  A168 );
 a29707a <=( A169  and  a29706a );
 a29710a <=( A199  and  A166 );
 a29713a <=( (not A201)  and  A200 );
 a29714a <=( a29713a  and  a29710a );
 a29715a <=( a29714a  and  a29707a );
 a29719a <=( A234  and  A233 );
 a29720a <=( (not A202)  and  a29719a );
 a29723a <=( A299  and  (not A298) );
 a29726a <=( A302  and  (not A301) );
 a29727a <=( a29726a  and  a29723a );
 a29728a <=( a29727a  and  a29720a );
 a29732a <=( (not A167)  and  A168 );
 a29733a <=( A169  and  a29732a );
 a29736a <=( A199  and  A166 );
 a29739a <=( (not A201)  and  A200 );
 a29740a <=( a29739a  and  a29736a );
 a29741a <=( a29740a  and  a29733a );
 a29745a <=( A234  and  A233 );
 a29746a <=( (not A202)  and  a29745a );
 a29749a <=( (not A299)  and  (not A298) );
 a29752a <=( (not A302)  and  A301 );
 a29753a <=( a29752a  and  a29749a );
 a29754a <=( a29753a  and  a29746a );
 a29758a <=( (not A167)  and  A168 );
 a29759a <=( A169  and  a29758a );
 a29762a <=( A199  and  A166 );
 a29765a <=( (not A201)  and  A200 );
 a29766a <=( a29765a  and  a29762a );
 a29767a <=( a29766a  and  a29759a );
 a29771a <=( A234  and  A233 );
 a29772a <=( (not A202)  and  a29771a );
 a29775a <=( A266  and  A265 );
 a29778a <=( (not A269)  and  A268 );
 a29779a <=( a29778a  and  a29775a );
 a29780a <=( a29779a  and  a29772a );
 a29784a <=( (not A167)  and  A168 );
 a29785a <=( A169  and  a29784a );
 a29788a <=( A199  and  A166 );
 a29791a <=( (not A201)  and  A200 );
 a29792a <=( a29791a  and  a29788a );
 a29793a <=( a29792a  and  a29785a );
 a29797a <=( A234  and  A233 );
 a29798a <=( (not A202)  and  a29797a );
 a29801a <=( A266  and  (not A265) );
 a29804a <=( A269  and  (not A268) );
 a29805a <=( a29804a  and  a29801a );
 a29806a <=( a29805a  and  a29798a );
 a29810a <=( (not A167)  and  A168 );
 a29811a <=( A169  and  a29810a );
 a29814a <=( A199  and  A166 );
 a29817a <=( (not A201)  and  A200 );
 a29818a <=( a29817a  and  a29814a );
 a29819a <=( a29818a  and  a29811a );
 a29823a <=( A234  and  A233 );
 a29824a <=( (not A202)  and  a29823a );
 a29827a <=( (not A266)  and  A265 );
 a29830a <=( A269  and  (not A268) );
 a29831a <=( a29830a  and  a29827a );
 a29832a <=( a29831a  and  a29824a );
 a29836a <=( (not A167)  and  A168 );
 a29837a <=( A169  and  a29836a );
 a29840a <=( A199  and  A166 );
 a29843a <=( (not A201)  and  A200 );
 a29844a <=( a29843a  and  a29840a );
 a29845a <=( a29844a  and  a29837a );
 a29849a <=( A234  and  A233 );
 a29850a <=( (not A202)  and  a29849a );
 a29853a <=( (not A266)  and  (not A265) );
 a29856a <=( (not A269)  and  A268 );
 a29857a <=( a29856a  and  a29853a );
 a29858a <=( a29857a  and  a29850a );
 a29862a <=( (not A167)  and  A168 );
 a29863a <=( A169  and  a29862a );
 a29866a <=( A199  and  A166 );
 a29869a <=( (not A201)  and  A200 );
 a29870a <=( a29869a  and  a29866a );
 a29871a <=( a29870a  and  a29863a );
 a29875a <=( A233  and  A232 );
 a29876a <=( (not A202)  and  a29875a );
 a29879a <=( (not A236)  and  A235 );
 a29882a <=( A300  and  A299 );
 a29883a <=( a29882a  and  a29879a );
 a29884a <=( a29883a  and  a29876a );
 a29888a <=( (not A167)  and  A168 );
 a29889a <=( A169  and  a29888a );
 a29892a <=( A199  and  A166 );
 a29895a <=( (not A201)  and  A200 );
 a29896a <=( a29895a  and  a29892a );
 a29897a <=( a29896a  and  a29889a );
 a29901a <=( A233  and  A232 );
 a29902a <=( (not A202)  and  a29901a );
 a29905a <=( (not A236)  and  A235 );
 a29908a <=( A300  and  A298 );
 a29909a <=( a29908a  and  a29905a );
 a29910a <=( a29909a  and  a29902a );
 a29914a <=( (not A167)  and  A168 );
 a29915a <=( A169  and  a29914a );
 a29918a <=( A199  and  A166 );
 a29921a <=( (not A201)  and  A200 );
 a29922a <=( a29921a  and  a29918a );
 a29923a <=( a29922a  and  a29915a );
 a29927a <=( A233  and  A232 );
 a29928a <=( (not A202)  and  a29927a );
 a29931a <=( (not A236)  and  A235 );
 a29934a <=( A267  and  A265 );
 a29935a <=( a29934a  and  a29931a );
 a29936a <=( a29935a  and  a29928a );
 a29940a <=( (not A167)  and  A168 );
 a29941a <=( A169  and  a29940a );
 a29944a <=( A199  and  A166 );
 a29947a <=( (not A201)  and  A200 );
 a29948a <=( a29947a  and  a29944a );
 a29949a <=( a29948a  and  a29941a );
 a29953a <=( A233  and  A232 );
 a29954a <=( (not A202)  and  a29953a );
 a29957a <=( (not A236)  and  A235 );
 a29960a <=( A267  and  A266 );
 a29961a <=( a29960a  and  a29957a );
 a29962a <=( a29961a  and  a29954a );
 a29966a <=( (not A167)  and  A168 );
 a29967a <=( A169  and  a29966a );
 a29970a <=( A199  and  A166 );
 a29973a <=( (not A201)  and  A200 );
 a29974a <=( a29973a  and  a29970a );
 a29975a <=( a29974a  and  a29967a );
 a29979a <=( A233  and  (not A232) );
 a29980a <=( (not A202)  and  a29979a );
 a29983a <=( A236  and  (not A235) );
 a29986a <=( A300  and  A299 );
 a29987a <=( a29986a  and  a29983a );
 a29988a <=( a29987a  and  a29980a );
 a29992a <=( (not A167)  and  A168 );
 a29993a <=( A169  and  a29992a );
 a29996a <=( A199  and  A166 );
 a29999a <=( (not A201)  and  A200 );
 a30000a <=( a29999a  and  a29996a );
 a30001a <=( a30000a  and  a29993a );
 a30005a <=( A233  and  (not A232) );
 a30006a <=( (not A202)  and  a30005a );
 a30009a <=( A236  and  (not A235) );
 a30012a <=( A300  and  A298 );
 a30013a <=( a30012a  and  a30009a );
 a30014a <=( a30013a  and  a30006a );
 a30018a <=( (not A167)  and  A168 );
 a30019a <=( A169  and  a30018a );
 a30022a <=( A199  and  A166 );
 a30025a <=( (not A201)  and  A200 );
 a30026a <=( a30025a  and  a30022a );
 a30027a <=( a30026a  and  a30019a );
 a30031a <=( A233  and  (not A232) );
 a30032a <=( (not A202)  and  a30031a );
 a30035a <=( A236  and  (not A235) );
 a30038a <=( A267  and  A265 );
 a30039a <=( a30038a  and  a30035a );
 a30040a <=( a30039a  and  a30032a );
 a30044a <=( (not A167)  and  A168 );
 a30045a <=( A169  and  a30044a );
 a30048a <=( A199  and  A166 );
 a30051a <=( (not A201)  and  A200 );
 a30052a <=( a30051a  and  a30048a );
 a30053a <=( a30052a  and  a30045a );
 a30057a <=( A233  and  (not A232) );
 a30058a <=( (not A202)  and  a30057a );
 a30061a <=( A236  and  (not A235) );
 a30064a <=( A267  and  A266 );
 a30065a <=( a30064a  and  a30061a );
 a30066a <=( a30065a  and  a30058a );
 a30070a <=( (not A167)  and  A168 );
 a30071a <=( A169  and  a30070a );
 a30074a <=( A199  and  A166 );
 a30077a <=( (not A201)  and  A200 );
 a30078a <=( a30077a  and  a30074a );
 a30079a <=( a30078a  and  a30071a );
 a30083a <=( (not A233)  and  A232 );
 a30084a <=( (not A202)  and  a30083a );
 a30087a <=( A236  and  (not A235) );
 a30090a <=( A300  and  A299 );
 a30091a <=( a30090a  and  a30087a );
 a30092a <=( a30091a  and  a30084a );
 a30096a <=( (not A167)  and  A168 );
 a30097a <=( A169  and  a30096a );
 a30100a <=( A199  and  A166 );
 a30103a <=( (not A201)  and  A200 );
 a30104a <=( a30103a  and  a30100a );
 a30105a <=( a30104a  and  a30097a );
 a30109a <=( (not A233)  and  A232 );
 a30110a <=( (not A202)  and  a30109a );
 a30113a <=( A236  and  (not A235) );
 a30116a <=( A300  and  A298 );
 a30117a <=( a30116a  and  a30113a );
 a30118a <=( a30117a  and  a30110a );
 a30122a <=( (not A167)  and  A168 );
 a30123a <=( A169  and  a30122a );
 a30126a <=( A199  and  A166 );
 a30129a <=( (not A201)  and  A200 );
 a30130a <=( a30129a  and  a30126a );
 a30131a <=( a30130a  and  a30123a );
 a30135a <=( (not A233)  and  A232 );
 a30136a <=( (not A202)  and  a30135a );
 a30139a <=( A236  and  (not A235) );
 a30142a <=( A267  and  A265 );
 a30143a <=( a30142a  and  a30139a );
 a30144a <=( a30143a  and  a30136a );
 a30148a <=( (not A167)  and  A168 );
 a30149a <=( A169  and  a30148a );
 a30152a <=( A199  and  A166 );
 a30155a <=( (not A201)  and  A200 );
 a30156a <=( a30155a  and  a30152a );
 a30157a <=( a30156a  and  a30149a );
 a30161a <=( (not A233)  and  A232 );
 a30162a <=( (not A202)  and  a30161a );
 a30165a <=( A236  and  (not A235) );
 a30168a <=( A267  and  A266 );
 a30169a <=( a30168a  and  a30165a );
 a30170a <=( a30169a  and  a30162a );
 a30174a <=( (not A167)  and  A168 );
 a30175a <=( A169  and  a30174a );
 a30178a <=( A199  and  A166 );
 a30181a <=( (not A201)  and  A200 );
 a30182a <=( a30181a  and  a30178a );
 a30183a <=( a30182a  and  a30175a );
 a30187a <=( (not A233)  and  (not A232) );
 a30188a <=( (not A202)  and  a30187a );
 a30191a <=( (not A236)  and  A235 );
 a30194a <=( A300  and  A299 );
 a30195a <=( a30194a  and  a30191a );
 a30196a <=( a30195a  and  a30188a );
 a30200a <=( (not A167)  and  A168 );
 a30201a <=( A169  and  a30200a );
 a30204a <=( A199  and  A166 );
 a30207a <=( (not A201)  and  A200 );
 a30208a <=( a30207a  and  a30204a );
 a30209a <=( a30208a  and  a30201a );
 a30213a <=( (not A233)  and  (not A232) );
 a30214a <=( (not A202)  and  a30213a );
 a30217a <=( (not A236)  and  A235 );
 a30220a <=( A300  and  A298 );
 a30221a <=( a30220a  and  a30217a );
 a30222a <=( a30221a  and  a30214a );
 a30226a <=( (not A167)  and  A168 );
 a30227a <=( A169  and  a30226a );
 a30230a <=( A199  and  A166 );
 a30233a <=( (not A201)  and  A200 );
 a30234a <=( a30233a  and  a30230a );
 a30235a <=( a30234a  and  a30227a );
 a30239a <=( (not A233)  and  (not A232) );
 a30240a <=( (not A202)  and  a30239a );
 a30243a <=( (not A236)  and  A235 );
 a30246a <=( A267  and  A265 );
 a30247a <=( a30246a  and  a30243a );
 a30248a <=( a30247a  and  a30240a );
 a30252a <=( (not A167)  and  A168 );
 a30253a <=( A169  and  a30252a );
 a30256a <=( A199  and  A166 );
 a30259a <=( (not A201)  and  A200 );
 a30260a <=( a30259a  and  a30256a );
 a30261a <=( a30260a  and  a30253a );
 a30265a <=( (not A233)  and  (not A232) );
 a30266a <=( (not A202)  and  a30265a );
 a30269a <=( (not A236)  and  A235 );
 a30272a <=( A267  and  A266 );
 a30273a <=( a30272a  and  a30269a );
 a30274a <=( a30273a  and  a30266a );
 a30278a <=( (not A167)  and  A168 );
 a30279a <=( A169  and  a30278a );
 a30282a <=( A199  and  A166 );
 a30285a <=( (not A201)  and  A200 );
 a30286a <=( a30285a  and  a30282a );
 a30287a <=( a30286a  and  a30279a );
 a30291a <=( A234  and  A232 );
 a30292a <=( A203  and  a30291a );
 a30295a <=( A299  and  A298 );
 a30298a <=( (not A302)  and  A301 );
 a30299a <=( a30298a  and  a30295a );
 a30300a <=( a30299a  and  a30292a );
 a30304a <=( (not A167)  and  A168 );
 a30305a <=( A169  and  a30304a );
 a30308a <=( A199  and  A166 );
 a30311a <=( (not A201)  and  A200 );
 a30312a <=( a30311a  and  a30308a );
 a30313a <=( a30312a  and  a30305a );
 a30317a <=( A234  and  A232 );
 a30318a <=( A203  and  a30317a );
 a30321a <=( (not A299)  and  A298 );
 a30324a <=( A302  and  (not A301) );
 a30325a <=( a30324a  and  a30321a );
 a30326a <=( a30325a  and  a30318a );
 a30330a <=( (not A167)  and  A168 );
 a30331a <=( A169  and  a30330a );
 a30334a <=( A199  and  A166 );
 a30337a <=( (not A201)  and  A200 );
 a30338a <=( a30337a  and  a30334a );
 a30339a <=( a30338a  and  a30331a );
 a30343a <=( A234  and  A232 );
 a30344a <=( A203  and  a30343a );
 a30347a <=( A299  and  (not A298) );
 a30350a <=( A302  and  (not A301) );
 a30351a <=( a30350a  and  a30347a );
 a30352a <=( a30351a  and  a30344a );
 a30356a <=( (not A167)  and  A168 );
 a30357a <=( A169  and  a30356a );
 a30360a <=( A199  and  A166 );
 a30363a <=( (not A201)  and  A200 );
 a30364a <=( a30363a  and  a30360a );
 a30365a <=( a30364a  and  a30357a );
 a30369a <=( A234  and  A232 );
 a30370a <=( A203  and  a30369a );
 a30373a <=( (not A299)  and  (not A298) );
 a30376a <=( (not A302)  and  A301 );
 a30377a <=( a30376a  and  a30373a );
 a30378a <=( a30377a  and  a30370a );
 a30382a <=( (not A167)  and  A168 );
 a30383a <=( A169  and  a30382a );
 a30386a <=( A199  and  A166 );
 a30389a <=( (not A201)  and  A200 );
 a30390a <=( a30389a  and  a30386a );
 a30391a <=( a30390a  and  a30383a );
 a30395a <=( A234  and  A232 );
 a30396a <=( A203  and  a30395a );
 a30399a <=( A266  and  A265 );
 a30402a <=( (not A269)  and  A268 );
 a30403a <=( a30402a  and  a30399a );
 a30404a <=( a30403a  and  a30396a );
 a30408a <=( (not A167)  and  A168 );
 a30409a <=( A169  and  a30408a );
 a30412a <=( A199  and  A166 );
 a30415a <=( (not A201)  and  A200 );
 a30416a <=( a30415a  and  a30412a );
 a30417a <=( a30416a  and  a30409a );
 a30421a <=( A234  and  A232 );
 a30422a <=( A203  and  a30421a );
 a30425a <=( A266  and  (not A265) );
 a30428a <=( A269  and  (not A268) );
 a30429a <=( a30428a  and  a30425a );
 a30430a <=( a30429a  and  a30422a );
 a30434a <=( (not A167)  and  A168 );
 a30435a <=( A169  and  a30434a );
 a30438a <=( A199  and  A166 );
 a30441a <=( (not A201)  and  A200 );
 a30442a <=( a30441a  and  a30438a );
 a30443a <=( a30442a  and  a30435a );
 a30447a <=( A234  and  A232 );
 a30448a <=( A203  and  a30447a );
 a30451a <=( (not A266)  and  A265 );
 a30454a <=( A269  and  (not A268) );
 a30455a <=( a30454a  and  a30451a );
 a30456a <=( a30455a  and  a30448a );
 a30460a <=( (not A167)  and  A168 );
 a30461a <=( A169  and  a30460a );
 a30464a <=( A199  and  A166 );
 a30467a <=( (not A201)  and  A200 );
 a30468a <=( a30467a  and  a30464a );
 a30469a <=( a30468a  and  a30461a );
 a30473a <=( A234  and  A232 );
 a30474a <=( A203  and  a30473a );
 a30477a <=( (not A266)  and  (not A265) );
 a30480a <=( (not A269)  and  A268 );
 a30481a <=( a30480a  and  a30477a );
 a30482a <=( a30481a  and  a30474a );
 a30486a <=( (not A167)  and  A168 );
 a30487a <=( A169  and  a30486a );
 a30490a <=( A199  and  A166 );
 a30493a <=( (not A201)  and  A200 );
 a30494a <=( a30493a  and  a30490a );
 a30495a <=( a30494a  and  a30487a );
 a30499a <=( A234  and  A233 );
 a30500a <=( A203  and  a30499a );
 a30503a <=( A299  and  A298 );
 a30506a <=( (not A302)  and  A301 );
 a30507a <=( a30506a  and  a30503a );
 a30508a <=( a30507a  and  a30500a );
 a30512a <=( (not A167)  and  A168 );
 a30513a <=( A169  and  a30512a );
 a30516a <=( A199  and  A166 );
 a30519a <=( (not A201)  and  A200 );
 a30520a <=( a30519a  and  a30516a );
 a30521a <=( a30520a  and  a30513a );
 a30525a <=( A234  and  A233 );
 a30526a <=( A203  and  a30525a );
 a30529a <=( (not A299)  and  A298 );
 a30532a <=( A302  and  (not A301) );
 a30533a <=( a30532a  and  a30529a );
 a30534a <=( a30533a  and  a30526a );
 a30538a <=( (not A167)  and  A168 );
 a30539a <=( A169  and  a30538a );
 a30542a <=( A199  and  A166 );
 a30545a <=( (not A201)  and  A200 );
 a30546a <=( a30545a  and  a30542a );
 a30547a <=( a30546a  and  a30539a );
 a30551a <=( A234  and  A233 );
 a30552a <=( A203  and  a30551a );
 a30555a <=( A299  and  (not A298) );
 a30558a <=( A302  and  (not A301) );
 a30559a <=( a30558a  and  a30555a );
 a30560a <=( a30559a  and  a30552a );
 a30564a <=( (not A167)  and  A168 );
 a30565a <=( A169  and  a30564a );
 a30568a <=( A199  and  A166 );
 a30571a <=( (not A201)  and  A200 );
 a30572a <=( a30571a  and  a30568a );
 a30573a <=( a30572a  and  a30565a );
 a30577a <=( A234  and  A233 );
 a30578a <=( A203  and  a30577a );
 a30581a <=( (not A299)  and  (not A298) );
 a30584a <=( (not A302)  and  A301 );
 a30585a <=( a30584a  and  a30581a );
 a30586a <=( a30585a  and  a30578a );
 a30590a <=( (not A167)  and  A168 );
 a30591a <=( A169  and  a30590a );
 a30594a <=( A199  and  A166 );
 a30597a <=( (not A201)  and  A200 );
 a30598a <=( a30597a  and  a30594a );
 a30599a <=( a30598a  and  a30591a );
 a30603a <=( A234  and  A233 );
 a30604a <=( A203  and  a30603a );
 a30607a <=( A266  and  A265 );
 a30610a <=( (not A269)  and  A268 );
 a30611a <=( a30610a  and  a30607a );
 a30612a <=( a30611a  and  a30604a );
 a30616a <=( (not A167)  and  A168 );
 a30617a <=( A169  and  a30616a );
 a30620a <=( A199  and  A166 );
 a30623a <=( (not A201)  and  A200 );
 a30624a <=( a30623a  and  a30620a );
 a30625a <=( a30624a  and  a30617a );
 a30629a <=( A234  and  A233 );
 a30630a <=( A203  and  a30629a );
 a30633a <=( A266  and  (not A265) );
 a30636a <=( A269  and  (not A268) );
 a30637a <=( a30636a  and  a30633a );
 a30638a <=( a30637a  and  a30630a );
 a30642a <=( (not A167)  and  A168 );
 a30643a <=( A169  and  a30642a );
 a30646a <=( A199  and  A166 );
 a30649a <=( (not A201)  and  A200 );
 a30650a <=( a30649a  and  a30646a );
 a30651a <=( a30650a  and  a30643a );
 a30655a <=( A234  and  A233 );
 a30656a <=( A203  and  a30655a );
 a30659a <=( (not A266)  and  A265 );
 a30662a <=( A269  and  (not A268) );
 a30663a <=( a30662a  and  a30659a );
 a30664a <=( a30663a  and  a30656a );
 a30668a <=( (not A167)  and  A168 );
 a30669a <=( A169  and  a30668a );
 a30672a <=( A199  and  A166 );
 a30675a <=( (not A201)  and  A200 );
 a30676a <=( a30675a  and  a30672a );
 a30677a <=( a30676a  and  a30669a );
 a30681a <=( A234  and  A233 );
 a30682a <=( A203  and  a30681a );
 a30685a <=( (not A266)  and  (not A265) );
 a30688a <=( (not A269)  and  A268 );
 a30689a <=( a30688a  and  a30685a );
 a30690a <=( a30689a  and  a30682a );
 a30694a <=( (not A167)  and  A168 );
 a30695a <=( A169  and  a30694a );
 a30698a <=( A199  and  A166 );
 a30701a <=( (not A201)  and  A200 );
 a30702a <=( a30701a  and  a30698a );
 a30703a <=( a30702a  and  a30695a );
 a30707a <=( A233  and  A232 );
 a30708a <=( A203  and  a30707a );
 a30711a <=( (not A236)  and  A235 );
 a30714a <=( A300  and  A299 );
 a30715a <=( a30714a  and  a30711a );
 a30716a <=( a30715a  and  a30708a );
 a30720a <=( (not A167)  and  A168 );
 a30721a <=( A169  and  a30720a );
 a30724a <=( A199  and  A166 );
 a30727a <=( (not A201)  and  A200 );
 a30728a <=( a30727a  and  a30724a );
 a30729a <=( a30728a  and  a30721a );
 a30733a <=( A233  and  A232 );
 a30734a <=( A203  and  a30733a );
 a30737a <=( (not A236)  and  A235 );
 a30740a <=( A300  and  A298 );
 a30741a <=( a30740a  and  a30737a );
 a30742a <=( a30741a  and  a30734a );
 a30746a <=( (not A167)  and  A168 );
 a30747a <=( A169  and  a30746a );
 a30750a <=( A199  and  A166 );
 a30753a <=( (not A201)  and  A200 );
 a30754a <=( a30753a  and  a30750a );
 a30755a <=( a30754a  and  a30747a );
 a30759a <=( A233  and  A232 );
 a30760a <=( A203  and  a30759a );
 a30763a <=( (not A236)  and  A235 );
 a30766a <=( A267  and  A265 );
 a30767a <=( a30766a  and  a30763a );
 a30768a <=( a30767a  and  a30760a );
 a30772a <=( (not A167)  and  A168 );
 a30773a <=( A169  and  a30772a );
 a30776a <=( A199  and  A166 );
 a30779a <=( (not A201)  and  A200 );
 a30780a <=( a30779a  and  a30776a );
 a30781a <=( a30780a  and  a30773a );
 a30785a <=( A233  and  A232 );
 a30786a <=( A203  and  a30785a );
 a30789a <=( (not A236)  and  A235 );
 a30792a <=( A267  and  A266 );
 a30793a <=( a30792a  and  a30789a );
 a30794a <=( a30793a  and  a30786a );
 a30798a <=( (not A167)  and  A168 );
 a30799a <=( A169  and  a30798a );
 a30802a <=( A199  and  A166 );
 a30805a <=( (not A201)  and  A200 );
 a30806a <=( a30805a  and  a30802a );
 a30807a <=( a30806a  and  a30799a );
 a30811a <=( A233  and  (not A232) );
 a30812a <=( A203  and  a30811a );
 a30815a <=( A236  and  (not A235) );
 a30818a <=( A300  and  A299 );
 a30819a <=( a30818a  and  a30815a );
 a30820a <=( a30819a  and  a30812a );
 a30824a <=( (not A167)  and  A168 );
 a30825a <=( A169  and  a30824a );
 a30828a <=( A199  and  A166 );
 a30831a <=( (not A201)  and  A200 );
 a30832a <=( a30831a  and  a30828a );
 a30833a <=( a30832a  and  a30825a );
 a30837a <=( A233  and  (not A232) );
 a30838a <=( A203  and  a30837a );
 a30841a <=( A236  and  (not A235) );
 a30844a <=( A300  and  A298 );
 a30845a <=( a30844a  and  a30841a );
 a30846a <=( a30845a  and  a30838a );
 a30850a <=( (not A167)  and  A168 );
 a30851a <=( A169  and  a30850a );
 a30854a <=( A199  and  A166 );
 a30857a <=( (not A201)  and  A200 );
 a30858a <=( a30857a  and  a30854a );
 a30859a <=( a30858a  and  a30851a );
 a30863a <=( A233  and  (not A232) );
 a30864a <=( A203  and  a30863a );
 a30867a <=( A236  and  (not A235) );
 a30870a <=( A267  and  A265 );
 a30871a <=( a30870a  and  a30867a );
 a30872a <=( a30871a  and  a30864a );
 a30876a <=( (not A167)  and  A168 );
 a30877a <=( A169  and  a30876a );
 a30880a <=( A199  and  A166 );
 a30883a <=( (not A201)  and  A200 );
 a30884a <=( a30883a  and  a30880a );
 a30885a <=( a30884a  and  a30877a );
 a30889a <=( A233  and  (not A232) );
 a30890a <=( A203  and  a30889a );
 a30893a <=( A236  and  (not A235) );
 a30896a <=( A267  and  A266 );
 a30897a <=( a30896a  and  a30893a );
 a30898a <=( a30897a  and  a30890a );
 a30902a <=( (not A167)  and  A168 );
 a30903a <=( A169  and  a30902a );
 a30906a <=( A199  and  A166 );
 a30909a <=( (not A201)  and  A200 );
 a30910a <=( a30909a  and  a30906a );
 a30911a <=( a30910a  and  a30903a );
 a30915a <=( (not A233)  and  A232 );
 a30916a <=( A203  and  a30915a );
 a30919a <=( A236  and  (not A235) );
 a30922a <=( A300  and  A299 );
 a30923a <=( a30922a  and  a30919a );
 a30924a <=( a30923a  and  a30916a );
 a30928a <=( (not A167)  and  A168 );
 a30929a <=( A169  and  a30928a );
 a30932a <=( A199  and  A166 );
 a30935a <=( (not A201)  and  A200 );
 a30936a <=( a30935a  and  a30932a );
 a30937a <=( a30936a  and  a30929a );
 a30941a <=( (not A233)  and  A232 );
 a30942a <=( A203  and  a30941a );
 a30945a <=( A236  and  (not A235) );
 a30948a <=( A300  and  A298 );
 a30949a <=( a30948a  and  a30945a );
 a30950a <=( a30949a  and  a30942a );
 a30954a <=( (not A167)  and  A168 );
 a30955a <=( A169  and  a30954a );
 a30958a <=( A199  and  A166 );
 a30961a <=( (not A201)  and  A200 );
 a30962a <=( a30961a  and  a30958a );
 a30963a <=( a30962a  and  a30955a );
 a30967a <=( (not A233)  and  A232 );
 a30968a <=( A203  and  a30967a );
 a30971a <=( A236  and  (not A235) );
 a30974a <=( A267  and  A265 );
 a30975a <=( a30974a  and  a30971a );
 a30976a <=( a30975a  and  a30968a );
 a30980a <=( (not A167)  and  A168 );
 a30981a <=( A169  and  a30980a );
 a30984a <=( A199  and  A166 );
 a30987a <=( (not A201)  and  A200 );
 a30988a <=( a30987a  and  a30984a );
 a30989a <=( a30988a  and  a30981a );
 a30993a <=( (not A233)  and  A232 );
 a30994a <=( A203  and  a30993a );
 a30997a <=( A236  and  (not A235) );
 a31000a <=( A267  and  A266 );
 a31001a <=( a31000a  and  a30997a );
 a31002a <=( a31001a  and  a30994a );
 a31006a <=( (not A167)  and  A168 );
 a31007a <=( A169  and  a31006a );
 a31010a <=( A199  and  A166 );
 a31013a <=( (not A201)  and  A200 );
 a31014a <=( a31013a  and  a31010a );
 a31015a <=( a31014a  and  a31007a );
 a31019a <=( (not A233)  and  (not A232) );
 a31020a <=( A203  and  a31019a );
 a31023a <=( (not A236)  and  A235 );
 a31026a <=( A300  and  A299 );
 a31027a <=( a31026a  and  a31023a );
 a31028a <=( a31027a  and  a31020a );
 a31032a <=( (not A167)  and  A168 );
 a31033a <=( A169  and  a31032a );
 a31036a <=( A199  and  A166 );
 a31039a <=( (not A201)  and  A200 );
 a31040a <=( a31039a  and  a31036a );
 a31041a <=( a31040a  and  a31033a );
 a31045a <=( (not A233)  and  (not A232) );
 a31046a <=( A203  and  a31045a );
 a31049a <=( (not A236)  and  A235 );
 a31052a <=( A300  and  A298 );
 a31053a <=( a31052a  and  a31049a );
 a31054a <=( a31053a  and  a31046a );
 a31058a <=( (not A167)  and  A168 );
 a31059a <=( A169  and  a31058a );
 a31062a <=( A199  and  A166 );
 a31065a <=( (not A201)  and  A200 );
 a31066a <=( a31065a  and  a31062a );
 a31067a <=( a31066a  and  a31059a );
 a31071a <=( (not A233)  and  (not A232) );
 a31072a <=( A203  and  a31071a );
 a31075a <=( (not A236)  and  A235 );
 a31078a <=( A267  and  A265 );
 a31079a <=( a31078a  and  a31075a );
 a31080a <=( a31079a  and  a31072a );
 a31084a <=( (not A167)  and  A168 );
 a31085a <=( A169  and  a31084a );
 a31088a <=( A199  and  A166 );
 a31091a <=( (not A201)  and  A200 );
 a31092a <=( a31091a  and  a31088a );
 a31093a <=( a31092a  and  a31085a );
 a31097a <=( (not A233)  and  (not A232) );
 a31098a <=( A203  and  a31097a );
 a31101a <=( (not A236)  and  A235 );
 a31104a <=( A267  and  A266 );
 a31105a <=( a31104a  and  a31101a );
 a31106a <=( a31105a  and  a31098a );
 a31110a <=( (not A167)  and  A168 );
 a31111a <=( A169  and  a31110a );
 a31114a <=( (not A199)  and  A166 );
 a31117a <=( (not A201)  and  A200 );
 a31118a <=( a31117a  and  a31114a );
 a31119a <=( a31118a  and  a31111a );
 a31123a <=( A234  and  A232 );
 a31124a <=( A202  and  a31123a );
 a31127a <=( A299  and  A298 );
 a31130a <=( (not A302)  and  A301 );
 a31131a <=( a31130a  and  a31127a );
 a31132a <=( a31131a  and  a31124a );
 a31136a <=( (not A167)  and  A168 );
 a31137a <=( A169  and  a31136a );
 a31140a <=( (not A199)  and  A166 );
 a31143a <=( (not A201)  and  A200 );
 a31144a <=( a31143a  and  a31140a );
 a31145a <=( a31144a  and  a31137a );
 a31149a <=( A234  and  A232 );
 a31150a <=( A202  and  a31149a );
 a31153a <=( (not A299)  and  A298 );
 a31156a <=( A302  and  (not A301) );
 a31157a <=( a31156a  and  a31153a );
 a31158a <=( a31157a  and  a31150a );
 a31162a <=( (not A167)  and  A168 );
 a31163a <=( A169  and  a31162a );
 a31166a <=( (not A199)  and  A166 );
 a31169a <=( (not A201)  and  A200 );
 a31170a <=( a31169a  and  a31166a );
 a31171a <=( a31170a  and  a31163a );
 a31175a <=( A234  and  A232 );
 a31176a <=( A202  and  a31175a );
 a31179a <=( A299  and  (not A298) );
 a31182a <=( A302  and  (not A301) );
 a31183a <=( a31182a  and  a31179a );
 a31184a <=( a31183a  and  a31176a );
 a31188a <=( (not A167)  and  A168 );
 a31189a <=( A169  and  a31188a );
 a31192a <=( (not A199)  and  A166 );
 a31195a <=( (not A201)  and  A200 );
 a31196a <=( a31195a  and  a31192a );
 a31197a <=( a31196a  and  a31189a );
 a31201a <=( A234  and  A232 );
 a31202a <=( A202  and  a31201a );
 a31205a <=( (not A299)  and  (not A298) );
 a31208a <=( (not A302)  and  A301 );
 a31209a <=( a31208a  and  a31205a );
 a31210a <=( a31209a  and  a31202a );
 a31214a <=( (not A167)  and  A168 );
 a31215a <=( A169  and  a31214a );
 a31218a <=( (not A199)  and  A166 );
 a31221a <=( (not A201)  and  A200 );
 a31222a <=( a31221a  and  a31218a );
 a31223a <=( a31222a  and  a31215a );
 a31227a <=( A234  and  A232 );
 a31228a <=( A202  and  a31227a );
 a31231a <=( A266  and  A265 );
 a31234a <=( (not A269)  and  A268 );
 a31235a <=( a31234a  and  a31231a );
 a31236a <=( a31235a  and  a31228a );
 a31240a <=( (not A167)  and  A168 );
 a31241a <=( A169  and  a31240a );
 a31244a <=( (not A199)  and  A166 );
 a31247a <=( (not A201)  and  A200 );
 a31248a <=( a31247a  and  a31244a );
 a31249a <=( a31248a  and  a31241a );
 a31253a <=( A234  and  A232 );
 a31254a <=( A202  and  a31253a );
 a31257a <=( A266  and  (not A265) );
 a31260a <=( A269  and  (not A268) );
 a31261a <=( a31260a  and  a31257a );
 a31262a <=( a31261a  and  a31254a );
 a31266a <=( (not A167)  and  A168 );
 a31267a <=( A169  and  a31266a );
 a31270a <=( (not A199)  and  A166 );
 a31273a <=( (not A201)  and  A200 );
 a31274a <=( a31273a  and  a31270a );
 a31275a <=( a31274a  and  a31267a );
 a31279a <=( A234  and  A232 );
 a31280a <=( A202  and  a31279a );
 a31283a <=( (not A266)  and  A265 );
 a31286a <=( A269  and  (not A268) );
 a31287a <=( a31286a  and  a31283a );
 a31288a <=( a31287a  and  a31280a );
 a31292a <=( (not A167)  and  A168 );
 a31293a <=( A169  and  a31292a );
 a31296a <=( (not A199)  and  A166 );
 a31299a <=( (not A201)  and  A200 );
 a31300a <=( a31299a  and  a31296a );
 a31301a <=( a31300a  and  a31293a );
 a31305a <=( A234  and  A232 );
 a31306a <=( A202  and  a31305a );
 a31309a <=( (not A266)  and  (not A265) );
 a31312a <=( (not A269)  and  A268 );
 a31313a <=( a31312a  and  a31309a );
 a31314a <=( a31313a  and  a31306a );
 a31318a <=( (not A167)  and  A168 );
 a31319a <=( A169  and  a31318a );
 a31322a <=( (not A199)  and  A166 );
 a31325a <=( (not A201)  and  A200 );
 a31326a <=( a31325a  and  a31322a );
 a31327a <=( a31326a  and  a31319a );
 a31331a <=( A234  and  A233 );
 a31332a <=( A202  and  a31331a );
 a31335a <=( A299  and  A298 );
 a31338a <=( (not A302)  and  A301 );
 a31339a <=( a31338a  and  a31335a );
 a31340a <=( a31339a  and  a31332a );
 a31344a <=( (not A167)  and  A168 );
 a31345a <=( A169  and  a31344a );
 a31348a <=( (not A199)  and  A166 );
 a31351a <=( (not A201)  and  A200 );
 a31352a <=( a31351a  and  a31348a );
 a31353a <=( a31352a  and  a31345a );
 a31357a <=( A234  and  A233 );
 a31358a <=( A202  and  a31357a );
 a31361a <=( (not A299)  and  A298 );
 a31364a <=( A302  and  (not A301) );
 a31365a <=( a31364a  and  a31361a );
 a31366a <=( a31365a  and  a31358a );
 a31370a <=( (not A167)  and  A168 );
 a31371a <=( A169  and  a31370a );
 a31374a <=( (not A199)  and  A166 );
 a31377a <=( (not A201)  and  A200 );
 a31378a <=( a31377a  and  a31374a );
 a31379a <=( a31378a  and  a31371a );
 a31383a <=( A234  and  A233 );
 a31384a <=( A202  and  a31383a );
 a31387a <=( A299  and  (not A298) );
 a31390a <=( A302  and  (not A301) );
 a31391a <=( a31390a  and  a31387a );
 a31392a <=( a31391a  and  a31384a );
 a31396a <=( (not A167)  and  A168 );
 a31397a <=( A169  and  a31396a );
 a31400a <=( (not A199)  and  A166 );
 a31403a <=( (not A201)  and  A200 );
 a31404a <=( a31403a  and  a31400a );
 a31405a <=( a31404a  and  a31397a );
 a31409a <=( A234  and  A233 );
 a31410a <=( A202  and  a31409a );
 a31413a <=( (not A299)  and  (not A298) );
 a31416a <=( (not A302)  and  A301 );
 a31417a <=( a31416a  and  a31413a );
 a31418a <=( a31417a  and  a31410a );
 a31422a <=( (not A167)  and  A168 );
 a31423a <=( A169  and  a31422a );
 a31426a <=( (not A199)  and  A166 );
 a31429a <=( (not A201)  and  A200 );
 a31430a <=( a31429a  and  a31426a );
 a31431a <=( a31430a  and  a31423a );
 a31435a <=( A234  and  A233 );
 a31436a <=( A202  and  a31435a );
 a31439a <=( A266  and  A265 );
 a31442a <=( (not A269)  and  A268 );
 a31443a <=( a31442a  and  a31439a );
 a31444a <=( a31443a  and  a31436a );
 a31448a <=( (not A167)  and  A168 );
 a31449a <=( A169  and  a31448a );
 a31452a <=( (not A199)  and  A166 );
 a31455a <=( (not A201)  and  A200 );
 a31456a <=( a31455a  and  a31452a );
 a31457a <=( a31456a  and  a31449a );
 a31461a <=( A234  and  A233 );
 a31462a <=( A202  and  a31461a );
 a31465a <=( A266  and  (not A265) );
 a31468a <=( A269  and  (not A268) );
 a31469a <=( a31468a  and  a31465a );
 a31470a <=( a31469a  and  a31462a );
 a31474a <=( (not A167)  and  A168 );
 a31475a <=( A169  and  a31474a );
 a31478a <=( (not A199)  and  A166 );
 a31481a <=( (not A201)  and  A200 );
 a31482a <=( a31481a  and  a31478a );
 a31483a <=( a31482a  and  a31475a );
 a31487a <=( A234  and  A233 );
 a31488a <=( A202  and  a31487a );
 a31491a <=( (not A266)  and  A265 );
 a31494a <=( A269  and  (not A268) );
 a31495a <=( a31494a  and  a31491a );
 a31496a <=( a31495a  and  a31488a );
 a31500a <=( (not A167)  and  A168 );
 a31501a <=( A169  and  a31500a );
 a31504a <=( (not A199)  and  A166 );
 a31507a <=( (not A201)  and  A200 );
 a31508a <=( a31507a  and  a31504a );
 a31509a <=( a31508a  and  a31501a );
 a31513a <=( A234  and  A233 );
 a31514a <=( A202  and  a31513a );
 a31517a <=( (not A266)  and  (not A265) );
 a31520a <=( (not A269)  and  A268 );
 a31521a <=( a31520a  and  a31517a );
 a31522a <=( a31521a  and  a31514a );
 a31526a <=( (not A167)  and  A168 );
 a31527a <=( A169  and  a31526a );
 a31530a <=( (not A199)  and  A166 );
 a31533a <=( (not A201)  and  A200 );
 a31534a <=( a31533a  and  a31530a );
 a31535a <=( a31534a  and  a31527a );
 a31539a <=( A233  and  A232 );
 a31540a <=( A202  and  a31539a );
 a31543a <=( (not A236)  and  A235 );
 a31546a <=( A300  and  A299 );
 a31547a <=( a31546a  and  a31543a );
 a31548a <=( a31547a  and  a31540a );
 a31552a <=( (not A167)  and  A168 );
 a31553a <=( A169  and  a31552a );
 a31556a <=( (not A199)  and  A166 );
 a31559a <=( (not A201)  and  A200 );
 a31560a <=( a31559a  and  a31556a );
 a31561a <=( a31560a  and  a31553a );
 a31565a <=( A233  and  A232 );
 a31566a <=( A202  and  a31565a );
 a31569a <=( (not A236)  and  A235 );
 a31572a <=( A300  and  A298 );
 a31573a <=( a31572a  and  a31569a );
 a31574a <=( a31573a  and  a31566a );
 a31578a <=( (not A167)  and  A168 );
 a31579a <=( A169  and  a31578a );
 a31582a <=( (not A199)  and  A166 );
 a31585a <=( (not A201)  and  A200 );
 a31586a <=( a31585a  and  a31582a );
 a31587a <=( a31586a  and  a31579a );
 a31591a <=( A233  and  A232 );
 a31592a <=( A202  and  a31591a );
 a31595a <=( (not A236)  and  A235 );
 a31598a <=( A267  and  A265 );
 a31599a <=( a31598a  and  a31595a );
 a31600a <=( a31599a  and  a31592a );
 a31604a <=( (not A167)  and  A168 );
 a31605a <=( A169  and  a31604a );
 a31608a <=( (not A199)  and  A166 );
 a31611a <=( (not A201)  and  A200 );
 a31612a <=( a31611a  and  a31608a );
 a31613a <=( a31612a  and  a31605a );
 a31617a <=( A233  and  A232 );
 a31618a <=( A202  and  a31617a );
 a31621a <=( (not A236)  and  A235 );
 a31624a <=( A267  and  A266 );
 a31625a <=( a31624a  and  a31621a );
 a31626a <=( a31625a  and  a31618a );
 a31630a <=( (not A167)  and  A168 );
 a31631a <=( A169  and  a31630a );
 a31634a <=( (not A199)  and  A166 );
 a31637a <=( (not A201)  and  A200 );
 a31638a <=( a31637a  and  a31634a );
 a31639a <=( a31638a  and  a31631a );
 a31643a <=( A233  and  (not A232) );
 a31644a <=( A202  and  a31643a );
 a31647a <=( A236  and  (not A235) );
 a31650a <=( A300  and  A299 );
 a31651a <=( a31650a  and  a31647a );
 a31652a <=( a31651a  and  a31644a );
 a31656a <=( (not A167)  and  A168 );
 a31657a <=( A169  and  a31656a );
 a31660a <=( (not A199)  and  A166 );
 a31663a <=( (not A201)  and  A200 );
 a31664a <=( a31663a  and  a31660a );
 a31665a <=( a31664a  and  a31657a );
 a31669a <=( A233  and  (not A232) );
 a31670a <=( A202  and  a31669a );
 a31673a <=( A236  and  (not A235) );
 a31676a <=( A300  and  A298 );
 a31677a <=( a31676a  and  a31673a );
 a31678a <=( a31677a  and  a31670a );
 a31682a <=( (not A167)  and  A168 );
 a31683a <=( A169  and  a31682a );
 a31686a <=( (not A199)  and  A166 );
 a31689a <=( (not A201)  and  A200 );
 a31690a <=( a31689a  and  a31686a );
 a31691a <=( a31690a  and  a31683a );
 a31695a <=( A233  and  (not A232) );
 a31696a <=( A202  and  a31695a );
 a31699a <=( A236  and  (not A235) );
 a31702a <=( A267  and  A265 );
 a31703a <=( a31702a  and  a31699a );
 a31704a <=( a31703a  and  a31696a );
 a31708a <=( (not A167)  and  A168 );
 a31709a <=( A169  and  a31708a );
 a31712a <=( (not A199)  and  A166 );
 a31715a <=( (not A201)  and  A200 );
 a31716a <=( a31715a  and  a31712a );
 a31717a <=( a31716a  and  a31709a );
 a31721a <=( A233  and  (not A232) );
 a31722a <=( A202  and  a31721a );
 a31725a <=( A236  and  (not A235) );
 a31728a <=( A267  and  A266 );
 a31729a <=( a31728a  and  a31725a );
 a31730a <=( a31729a  and  a31722a );
 a31734a <=( (not A167)  and  A168 );
 a31735a <=( A169  and  a31734a );
 a31738a <=( (not A199)  and  A166 );
 a31741a <=( (not A201)  and  A200 );
 a31742a <=( a31741a  and  a31738a );
 a31743a <=( a31742a  and  a31735a );
 a31747a <=( (not A233)  and  A232 );
 a31748a <=( A202  and  a31747a );
 a31751a <=( A236  and  (not A235) );
 a31754a <=( A300  and  A299 );
 a31755a <=( a31754a  and  a31751a );
 a31756a <=( a31755a  and  a31748a );
 a31760a <=( (not A167)  and  A168 );
 a31761a <=( A169  and  a31760a );
 a31764a <=( (not A199)  and  A166 );
 a31767a <=( (not A201)  and  A200 );
 a31768a <=( a31767a  and  a31764a );
 a31769a <=( a31768a  and  a31761a );
 a31773a <=( (not A233)  and  A232 );
 a31774a <=( A202  and  a31773a );
 a31777a <=( A236  and  (not A235) );
 a31780a <=( A300  and  A298 );
 a31781a <=( a31780a  and  a31777a );
 a31782a <=( a31781a  and  a31774a );
 a31786a <=( (not A167)  and  A168 );
 a31787a <=( A169  and  a31786a );
 a31790a <=( (not A199)  and  A166 );
 a31793a <=( (not A201)  and  A200 );
 a31794a <=( a31793a  and  a31790a );
 a31795a <=( a31794a  and  a31787a );
 a31799a <=( (not A233)  and  A232 );
 a31800a <=( A202  and  a31799a );
 a31803a <=( A236  and  (not A235) );
 a31806a <=( A267  and  A265 );
 a31807a <=( a31806a  and  a31803a );
 a31808a <=( a31807a  and  a31800a );
 a31812a <=( (not A167)  and  A168 );
 a31813a <=( A169  and  a31812a );
 a31816a <=( (not A199)  and  A166 );
 a31819a <=( (not A201)  and  A200 );
 a31820a <=( a31819a  and  a31816a );
 a31821a <=( a31820a  and  a31813a );
 a31825a <=( (not A233)  and  A232 );
 a31826a <=( A202  and  a31825a );
 a31829a <=( A236  and  (not A235) );
 a31832a <=( A267  and  A266 );
 a31833a <=( a31832a  and  a31829a );
 a31834a <=( a31833a  and  a31826a );
 a31838a <=( (not A167)  and  A168 );
 a31839a <=( A169  and  a31838a );
 a31842a <=( (not A199)  and  A166 );
 a31845a <=( (not A201)  and  A200 );
 a31846a <=( a31845a  and  a31842a );
 a31847a <=( a31846a  and  a31839a );
 a31851a <=( (not A233)  and  (not A232) );
 a31852a <=( A202  and  a31851a );
 a31855a <=( (not A236)  and  A235 );
 a31858a <=( A300  and  A299 );
 a31859a <=( a31858a  and  a31855a );
 a31860a <=( a31859a  and  a31852a );
 a31864a <=( (not A167)  and  A168 );
 a31865a <=( A169  and  a31864a );
 a31868a <=( (not A199)  and  A166 );
 a31871a <=( (not A201)  and  A200 );
 a31872a <=( a31871a  and  a31868a );
 a31873a <=( a31872a  and  a31865a );
 a31877a <=( (not A233)  and  (not A232) );
 a31878a <=( A202  and  a31877a );
 a31881a <=( (not A236)  and  A235 );
 a31884a <=( A300  and  A298 );
 a31885a <=( a31884a  and  a31881a );
 a31886a <=( a31885a  and  a31878a );
 a31890a <=( (not A167)  and  A168 );
 a31891a <=( A169  and  a31890a );
 a31894a <=( (not A199)  and  A166 );
 a31897a <=( (not A201)  and  A200 );
 a31898a <=( a31897a  and  a31894a );
 a31899a <=( a31898a  and  a31891a );
 a31903a <=( (not A233)  and  (not A232) );
 a31904a <=( A202  and  a31903a );
 a31907a <=( (not A236)  and  A235 );
 a31910a <=( A267  and  A265 );
 a31911a <=( a31910a  and  a31907a );
 a31912a <=( a31911a  and  a31904a );
 a31916a <=( (not A167)  and  A168 );
 a31917a <=( A169  and  a31916a );
 a31920a <=( (not A199)  and  A166 );
 a31923a <=( (not A201)  and  A200 );
 a31924a <=( a31923a  and  a31920a );
 a31925a <=( a31924a  and  a31917a );
 a31929a <=( (not A233)  and  (not A232) );
 a31930a <=( A202  and  a31929a );
 a31933a <=( (not A236)  and  A235 );
 a31936a <=( A267  and  A266 );
 a31937a <=( a31936a  and  a31933a );
 a31938a <=( a31937a  and  a31930a );
 a31942a <=( (not A167)  and  A168 );
 a31943a <=( A169  and  a31942a );
 a31946a <=( (not A199)  and  A166 );
 a31949a <=( (not A201)  and  A200 );
 a31950a <=( a31949a  and  a31946a );
 a31951a <=( a31950a  and  a31943a );
 a31955a <=( A234  and  A232 );
 a31956a <=( (not A203)  and  a31955a );
 a31959a <=( A299  and  A298 );
 a31962a <=( (not A302)  and  A301 );
 a31963a <=( a31962a  and  a31959a );
 a31964a <=( a31963a  and  a31956a );
 a31968a <=( (not A167)  and  A168 );
 a31969a <=( A169  and  a31968a );
 a31972a <=( (not A199)  and  A166 );
 a31975a <=( (not A201)  and  A200 );
 a31976a <=( a31975a  and  a31972a );
 a31977a <=( a31976a  and  a31969a );
 a31981a <=( A234  and  A232 );
 a31982a <=( (not A203)  and  a31981a );
 a31985a <=( (not A299)  and  A298 );
 a31988a <=( A302  and  (not A301) );
 a31989a <=( a31988a  and  a31985a );
 a31990a <=( a31989a  and  a31982a );
 a31994a <=( (not A167)  and  A168 );
 a31995a <=( A169  and  a31994a );
 a31998a <=( (not A199)  and  A166 );
 a32001a <=( (not A201)  and  A200 );
 a32002a <=( a32001a  and  a31998a );
 a32003a <=( a32002a  and  a31995a );
 a32007a <=( A234  and  A232 );
 a32008a <=( (not A203)  and  a32007a );
 a32011a <=( A299  and  (not A298) );
 a32014a <=( A302  and  (not A301) );
 a32015a <=( a32014a  and  a32011a );
 a32016a <=( a32015a  and  a32008a );
 a32020a <=( (not A167)  and  A168 );
 a32021a <=( A169  and  a32020a );
 a32024a <=( (not A199)  and  A166 );
 a32027a <=( (not A201)  and  A200 );
 a32028a <=( a32027a  and  a32024a );
 a32029a <=( a32028a  and  a32021a );
 a32033a <=( A234  and  A232 );
 a32034a <=( (not A203)  and  a32033a );
 a32037a <=( (not A299)  and  (not A298) );
 a32040a <=( (not A302)  and  A301 );
 a32041a <=( a32040a  and  a32037a );
 a32042a <=( a32041a  and  a32034a );
 a32046a <=( (not A167)  and  A168 );
 a32047a <=( A169  and  a32046a );
 a32050a <=( (not A199)  and  A166 );
 a32053a <=( (not A201)  and  A200 );
 a32054a <=( a32053a  and  a32050a );
 a32055a <=( a32054a  and  a32047a );
 a32059a <=( A234  and  A232 );
 a32060a <=( (not A203)  and  a32059a );
 a32063a <=( A266  and  A265 );
 a32066a <=( (not A269)  and  A268 );
 a32067a <=( a32066a  and  a32063a );
 a32068a <=( a32067a  and  a32060a );
 a32072a <=( (not A167)  and  A168 );
 a32073a <=( A169  and  a32072a );
 a32076a <=( (not A199)  and  A166 );
 a32079a <=( (not A201)  and  A200 );
 a32080a <=( a32079a  and  a32076a );
 a32081a <=( a32080a  and  a32073a );
 a32085a <=( A234  and  A232 );
 a32086a <=( (not A203)  and  a32085a );
 a32089a <=( A266  and  (not A265) );
 a32092a <=( A269  and  (not A268) );
 a32093a <=( a32092a  and  a32089a );
 a32094a <=( a32093a  and  a32086a );
 a32098a <=( (not A167)  and  A168 );
 a32099a <=( A169  and  a32098a );
 a32102a <=( (not A199)  and  A166 );
 a32105a <=( (not A201)  and  A200 );
 a32106a <=( a32105a  and  a32102a );
 a32107a <=( a32106a  and  a32099a );
 a32111a <=( A234  and  A232 );
 a32112a <=( (not A203)  and  a32111a );
 a32115a <=( (not A266)  and  A265 );
 a32118a <=( A269  and  (not A268) );
 a32119a <=( a32118a  and  a32115a );
 a32120a <=( a32119a  and  a32112a );
 a32124a <=( (not A167)  and  A168 );
 a32125a <=( A169  and  a32124a );
 a32128a <=( (not A199)  and  A166 );
 a32131a <=( (not A201)  and  A200 );
 a32132a <=( a32131a  and  a32128a );
 a32133a <=( a32132a  and  a32125a );
 a32137a <=( A234  and  A232 );
 a32138a <=( (not A203)  and  a32137a );
 a32141a <=( (not A266)  and  (not A265) );
 a32144a <=( (not A269)  and  A268 );
 a32145a <=( a32144a  and  a32141a );
 a32146a <=( a32145a  and  a32138a );
 a32150a <=( (not A167)  and  A168 );
 a32151a <=( A169  and  a32150a );
 a32154a <=( (not A199)  and  A166 );
 a32157a <=( (not A201)  and  A200 );
 a32158a <=( a32157a  and  a32154a );
 a32159a <=( a32158a  and  a32151a );
 a32163a <=( A234  and  A233 );
 a32164a <=( (not A203)  and  a32163a );
 a32167a <=( A299  and  A298 );
 a32170a <=( (not A302)  and  A301 );
 a32171a <=( a32170a  and  a32167a );
 a32172a <=( a32171a  and  a32164a );
 a32176a <=( (not A167)  and  A168 );
 a32177a <=( A169  and  a32176a );
 a32180a <=( (not A199)  and  A166 );
 a32183a <=( (not A201)  and  A200 );
 a32184a <=( a32183a  and  a32180a );
 a32185a <=( a32184a  and  a32177a );
 a32189a <=( A234  and  A233 );
 a32190a <=( (not A203)  and  a32189a );
 a32193a <=( (not A299)  and  A298 );
 a32196a <=( A302  and  (not A301) );
 a32197a <=( a32196a  and  a32193a );
 a32198a <=( a32197a  and  a32190a );
 a32202a <=( (not A167)  and  A168 );
 a32203a <=( A169  and  a32202a );
 a32206a <=( (not A199)  and  A166 );
 a32209a <=( (not A201)  and  A200 );
 a32210a <=( a32209a  and  a32206a );
 a32211a <=( a32210a  and  a32203a );
 a32215a <=( A234  and  A233 );
 a32216a <=( (not A203)  and  a32215a );
 a32219a <=( A299  and  (not A298) );
 a32222a <=( A302  and  (not A301) );
 a32223a <=( a32222a  and  a32219a );
 a32224a <=( a32223a  and  a32216a );
 a32228a <=( (not A167)  and  A168 );
 a32229a <=( A169  and  a32228a );
 a32232a <=( (not A199)  and  A166 );
 a32235a <=( (not A201)  and  A200 );
 a32236a <=( a32235a  and  a32232a );
 a32237a <=( a32236a  and  a32229a );
 a32241a <=( A234  and  A233 );
 a32242a <=( (not A203)  and  a32241a );
 a32245a <=( (not A299)  and  (not A298) );
 a32248a <=( (not A302)  and  A301 );
 a32249a <=( a32248a  and  a32245a );
 a32250a <=( a32249a  and  a32242a );
 a32254a <=( (not A167)  and  A168 );
 a32255a <=( A169  and  a32254a );
 a32258a <=( (not A199)  and  A166 );
 a32261a <=( (not A201)  and  A200 );
 a32262a <=( a32261a  and  a32258a );
 a32263a <=( a32262a  and  a32255a );
 a32267a <=( A234  and  A233 );
 a32268a <=( (not A203)  and  a32267a );
 a32271a <=( A266  and  A265 );
 a32274a <=( (not A269)  and  A268 );
 a32275a <=( a32274a  and  a32271a );
 a32276a <=( a32275a  and  a32268a );
 a32280a <=( (not A167)  and  A168 );
 a32281a <=( A169  and  a32280a );
 a32284a <=( (not A199)  and  A166 );
 a32287a <=( (not A201)  and  A200 );
 a32288a <=( a32287a  and  a32284a );
 a32289a <=( a32288a  and  a32281a );
 a32293a <=( A234  and  A233 );
 a32294a <=( (not A203)  and  a32293a );
 a32297a <=( A266  and  (not A265) );
 a32300a <=( A269  and  (not A268) );
 a32301a <=( a32300a  and  a32297a );
 a32302a <=( a32301a  and  a32294a );
 a32306a <=( (not A167)  and  A168 );
 a32307a <=( A169  and  a32306a );
 a32310a <=( (not A199)  and  A166 );
 a32313a <=( (not A201)  and  A200 );
 a32314a <=( a32313a  and  a32310a );
 a32315a <=( a32314a  and  a32307a );
 a32319a <=( A234  and  A233 );
 a32320a <=( (not A203)  and  a32319a );
 a32323a <=( (not A266)  and  A265 );
 a32326a <=( A269  and  (not A268) );
 a32327a <=( a32326a  and  a32323a );
 a32328a <=( a32327a  and  a32320a );
 a32332a <=( (not A167)  and  A168 );
 a32333a <=( A169  and  a32332a );
 a32336a <=( (not A199)  and  A166 );
 a32339a <=( (not A201)  and  A200 );
 a32340a <=( a32339a  and  a32336a );
 a32341a <=( a32340a  and  a32333a );
 a32345a <=( A234  and  A233 );
 a32346a <=( (not A203)  and  a32345a );
 a32349a <=( (not A266)  and  (not A265) );
 a32352a <=( (not A269)  and  A268 );
 a32353a <=( a32352a  and  a32349a );
 a32354a <=( a32353a  and  a32346a );
 a32358a <=( (not A167)  and  A168 );
 a32359a <=( A169  and  a32358a );
 a32362a <=( (not A199)  and  A166 );
 a32365a <=( (not A201)  and  A200 );
 a32366a <=( a32365a  and  a32362a );
 a32367a <=( a32366a  and  a32359a );
 a32371a <=( A233  and  A232 );
 a32372a <=( (not A203)  and  a32371a );
 a32375a <=( (not A236)  and  A235 );
 a32378a <=( A300  and  A299 );
 a32379a <=( a32378a  and  a32375a );
 a32380a <=( a32379a  and  a32372a );
 a32384a <=( (not A167)  and  A168 );
 a32385a <=( A169  and  a32384a );
 a32388a <=( (not A199)  and  A166 );
 a32391a <=( (not A201)  and  A200 );
 a32392a <=( a32391a  and  a32388a );
 a32393a <=( a32392a  and  a32385a );
 a32397a <=( A233  and  A232 );
 a32398a <=( (not A203)  and  a32397a );
 a32401a <=( (not A236)  and  A235 );
 a32404a <=( A300  and  A298 );
 a32405a <=( a32404a  and  a32401a );
 a32406a <=( a32405a  and  a32398a );
 a32410a <=( (not A167)  and  A168 );
 a32411a <=( A169  and  a32410a );
 a32414a <=( (not A199)  and  A166 );
 a32417a <=( (not A201)  and  A200 );
 a32418a <=( a32417a  and  a32414a );
 a32419a <=( a32418a  and  a32411a );
 a32423a <=( A233  and  A232 );
 a32424a <=( (not A203)  and  a32423a );
 a32427a <=( (not A236)  and  A235 );
 a32430a <=( A267  and  A265 );
 a32431a <=( a32430a  and  a32427a );
 a32432a <=( a32431a  and  a32424a );
 a32436a <=( (not A167)  and  A168 );
 a32437a <=( A169  and  a32436a );
 a32440a <=( (not A199)  and  A166 );
 a32443a <=( (not A201)  and  A200 );
 a32444a <=( a32443a  and  a32440a );
 a32445a <=( a32444a  and  a32437a );
 a32449a <=( A233  and  A232 );
 a32450a <=( (not A203)  and  a32449a );
 a32453a <=( (not A236)  and  A235 );
 a32456a <=( A267  and  A266 );
 a32457a <=( a32456a  and  a32453a );
 a32458a <=( a32457a  and  a32450a );
 a32462a <=( (not A167)  and  A168 );
 a32463a <=( A169  and  a32462a );
 a32466a <=( (not A199)  and  A166 );
 a32469a <=( (not A201)  and  A200 );
 a32470a <=( a32469a  and  a32466a );
 a32471a <=( a32470a  and  a32463a );
 a32475a <=( A233  and  (not A232) );
 a32476a <=( (not A203)  and  a32475a );
 a32479a <=( A236  and  (not A235) );
 a32482a <=( A300  and  A299 );
 a32483a <=( a32482a  and  a32479a );
 a32484a <=( a32483a  and  a32476a );
 a32488a <=( (not A167)  and  A168 );
 a32489a <=( A169  and  a32488a );
 a32492a <=( (not A199)  and  A166 );
 a32495a <=( (not A201)  and  A200 );
 a32496a <=( a32495a  and  a32492a );
 a32497a <=( a32496a  and  a32489a );
 a32501a <=( A233  and  (not A232) );
 a32502a <=( (not A203)  and  a32501a );
 a32505a <=( A236  and  (not A235) );
 a32508a <=( A300  and  A298 );
 a32509a <=( a32508a  and  a32505a );
 a32510a <=( a32509a  and  a32502a );
 a32514a <=( (not A167)  and  A168 );
 a32515a <=( A169  and  a32514a );
 a32518a <=( (not A199)  and  A166 );
 a32521a <=( (not A201)  and  A200 );
 a32522a <=( a32521a  and  a32518a );
 a32523a <=( a32522a  and  a32515a );
 a32527a <=( A233  and  (not A232) );
 a32528a <=( (not A203)  and  a32527a );
 a32531a <=( A236  and  (not A235) );
 a32534a <=( A267  and  A265 );
 a32535a <=( a32534a  and  a32531a );
 a32536a <=( a32535a  and  a32528a );
 a32540a <=( (not A167)  and  A168 );
 a32541a <=( A169  and  a32540a );
 a32544a <=( (not A199)  and  A166 );
 a32547a <=( (not A201)  and  A200 );
 a32548a <=( a32547a  and  a32544a );
 a32549a <=( a32548a  and  a32541a );
 a32553a <=( A233  and  (not A232) );
 a32554a <=( (not A203)  and  a32553a );
 a32557a <=( A236  and  (not A235) );
 a32560a <=( A267  and  A266 );
 a32561a <=( a32560a  and  a32557a );
 a32562a <=( a32561a  and  a32554a );
 a32566a <=( (not A167)  and  A168 );
 a32567a <=( A169  and  a32566a );
 a32570a <=( (not A199)  and  A166 );
 a32573a <=( (not A201)  and  A200 );
 a32574a <=( a32573a  and  a32570a );
 a32575a <=( a32574a  and  a32567a );
 a32579a <=( (not A233)  and  A232 );
 a32580a <=( (not A203)  and  a32579a );
 a32583a <=( A236  and  (not A235) );
 a32586a <=( A300  and  A299 );
 a32587a <=( a32586a  and  a32583a );
 a32588a <=( a32587a  and  a32580a );
 a32592a <=( (not A167)  and  A168 );
 a32593a <=( A169  and  a32592a );
 a32596a <=( (not A199)  and  A166 );
 a32599a <=( (not A201)  and  A200 );
 a32600a <=( a32599a  and  a32596a );
 a32601a <=( a32600a  and  a32593a );
 a32605a <=( (not A233)  and  A232 );
 a32606a <=( (not A203)  and  a32605a );
 a32609a <=( A236  and  (not A235) );
 a32612a <=( A300  and  A298 );
 a32613a <=( a32612a  and  a32609a );
 a32614a <=( a32613a  and  a32606a );
 a32618a <=( (not A167)  and  A168 );
 a32619a <=( A169  and  a32618a );
 a32622a <=( (not A199)  and  A166 );
 a32625a <=( (not A201)  and  A200 );
 a32626a <=( a32625a  and  a32622a );
 a32627a <=( a32626a  and  a32619a );
 a32631a <=( (not A233)  and  A232 );
 a32632a <=( (not A203)  and  a32631a );
 a32635a <=( A236  and  (not A235) );
 a32638a <=( A267  and  A265 );
 a32639a <=( a32638a  and  a32635a );
 a32640a <=( a32639a  and  a32632a );
 a32644a <=( (not A167)  and  A168 );
 a32645a <=( A169  and  a32644a );
 a32648a <=( (not A199)  and  A166 );
 a32651a <=( (not A201)  and  A200 );
 a32652a <=( a32651a  and  a32648a );
 a32653a <=( a32652a  and  a32645a );
 a32657a <=( (not A233)  and  A232 );
 a32658a <=( (not A203)  and  a32657a );
 a32661a <=( A236  and  (not A235) );
 a32664a <=( A267  and  A266 );
 a32665a <=( a32664a  and  a32661a );
 a32666a <=( a32665a  and  a32658a );
 a32670a <=( (not A167)  and  A168 );
 a32671a <=( A169  and  a32670a );
 a32674a <=( (not A199)  and  A166 );
 a32677a <=( (not A201)  and  A200 );
 a32678a <=( a32677a  and  a32674a );
 a32679a <=( a32678a  and  a32671a );
 a32683a <=( (not A233)  and  (not A232) );
 a32684a <=( (not A203)  and  a32683a );
 a32687a <=( (not A236)  and  A235 );
 a32690a <=( A300  and  A299 );
 a32691a <=( a32690a  and  a32687a );
 a32692a <=( a32691a  and  a32684a );
 a32696a <=( (not A167)  and  A168 );
 a32697a <=( A169  and  a32696a );
 a32700a <=( (not A199)  and  A166 );
 a32703a <=( (not A201)  and  A200 );
 a32704a <=( a32703a  and  a32700a );
 a32705a <=( a32704a  and  a32697a );
 a32709a <=( (not A233)  and  (not A232) );
 a32710a <=( (not A203)  and  a32709a );
 a32713a <=( (not A236)  and  A235 );
 a32716a <=( A300  and  A298 );
 a32717a <=( a32716a  and  a32713a );
 a32718a <=( a32717a  and  a32710a );
 a32722a <=( (not A167)  and  A168 );
 a32723a <=( A169  and  a32722a );
 a32726a <=( (not A199)  and  A166 );
 a32729a <=( (not A201)  and  A200 );
 a32730a <=( a32729a  and  a32726a );
 a32731a <=( a32730a  and  a32723a );
 a32735a <=( (not A233)  and  (not A232) );
 a32736a <=( (not A203)  and  a32735a );
 a32739a <=( (not A236)  and  A235 );
 a32742a <=( A267  and  A265 );
 a32743a <=( a32742a  and  a32739a );
 a32744a <=( a32743a  and  a32736a );
 a32748a <=( (not A167)  and  A168 );
 a32749a <=( A169  and  a32748a );
 a32752a <=( (not A199)  and  A166 );
 a32755a <=( (not A201)  and  A200 );
 a32756a <=( a32755a  and  a32752a );
 a32757a <=( a32756a  and  a32749a );
 a32761a <=( (not A233)  and  (not A232) );
 a32762a <=( (not A203)  and  a32761a );
 a32765a <=( (not A236)  and  A235 );
 a32768a <=( A267  and  A266 );
 a32769a <=( a32768a  and  a32765a );
 a32770a <=( a32769a  and  a32762a );
 a32774a <=( (not A167)  and  A168 );
 a32775a <=( A169  and  a32774a );
 a32778a <=( A199  and  A166 );
 a32781a <=( (not A201)  and  (not A200) );
 a32782a <=( a32781a  and  a32778a );
 a32783a <=( a32782a  and  a32775a );
 a32787a <=( A234  and  A232 );
 a32788a <=( A202  and  a32787a );
 a32791a <=( A299  and  A298 );
 a32794a <=( (not A302)  and  A301 );
 a32795a <=( a32794a  and  a32791a );
 a32796a <=( a32795a  and  a32788a );
 a32800a <=( (not A167)  and  A168 );
 a32801a <=( A169  and  a32800a );
 a32804a <=( A199  and  A166 );
 a32807a <=( (not A201)  and  (not A200) );
 a32808a <=( a32807a  and  a32804a );
 a32809a <=( a32808a  and  a32801a );
 a32813a <=( A234  and  A232 );
 a32814a <=( A202  and  a32813a );
 a32817a <=( (not A299)  and  A298 );
 a32820a <=( A302  and  (not A301) );
 a32821a <=( a32820a  and  a32817a );
 a32822a <=( a32821a  and  a32814a );
 a32826a <=( (not A167)  and  A168 );
 a32827a <=( A169  and  a32826a );
 a32830a <=( A199  and  A166 );
 a32833a <=( (not A201)  and  (not A200) );
 a32834a <=( a32833a  and  a32830a );
 a32835a <=( a32834a  and  a32827a );
 a32839a <=( A234  and  A232 );
 a32840a <=( A202  and  a32839a );
 a32843a <=( A299  and  (not A298) );
 a32846a <=( A302  and  (not A301) );
 a32847a <=( a32846a  and  a32843a );
 a32848a <=( a32847a  and  a32840a );
 a32852a <=( (not A167)  and  A168 );
 a32853a <=( A169  and  a32852a );
 a32856a <=( A199  and  A166 );
 a32859a <=( (not A201)  and  (not A200) );
 a32860a <=( a32859a  and  a32856a );
 a32861a <=( a32860a  and  a32853a );
 a32865a <=( A234  and  A232 );
 a32866a <=( A202  and  a32865a );
 a32869a <=( (not A299)  and  (not A298) );
 a32872a <=( (not A302)  and  A301 );
 a32873a <=( a32872a  and  a32869a );
 a32874a <=( a32873a  and  a32866a );
 a32878a <=( (not A167)  and  A168 );
 a32879a <=( A169  and  a32878a );
 a32882a <=( A199  and  A166 );
 a32885a <=( (not A201)  and  (not A200) );
 a32886a <=( a32885a  and  a32882a );
 a32887a <=( a32886a  and  a32879a );
 a32891a <=( A234  and  A232 );
 a32892a <=( A202  and  a32891a );
 a32895a <=( A266  and  A265 );
 a32898a <=( (not A269)  and  A268 );
 a32899a <=( a32898a  and  a32895a );
 a32900a <=( a32899a  and  a32892a );
 a32904a <=( (not A167)  and  A168 );
 a32905a <=( A169  and  a32904a );
 a32908a <=( A199  and  A166 );
 a32911a <=( (not A201)  and  (not A200) );
 a32912a <=( a32911a  and  a32908a );
 a32913a <=( a32912a  and  a32905a );
 a32917a <=( A234  and  A232 );
 a32918a <=( A202  and  a32917a );
 a32921a <=( A266  and  (not A265) );
 a32924a <=( A269  and  (not A268) );
 a32925a <=( a32924a  and  a32921a );
 a32926a <=( a32925a  and  a32918a );
 a32930a <=( (not A167)  and  A168 );
 a32931a <=( A169  and  a32930a );
 a32934a <=( A199  and  A166 );
 a32937a <=( (not A201)  and  (not A200) );
 a32938a <=( a32937a  and  a32934a );
 a32939a <=( a32938a  and  a32931a );
 a32943a <=( A234  and  A232 );
 a32944a <=( A202  and  a32943a );
 a32947a <=( (not A266)  and  A265 );
 a32950a <=( A269  and  (not A268) );
 a32951a <=( a32950a  and  a32947a );
 a32952a <=( a32951a  and  a32944a );
 a32956a <=( (not A167)  and  A168 );
 a32957a <=( A169  and  a32956a );
 a32960a <=( A199  and  A166 );
 a32963a <=( (not A201)  and  (not A200) );
 a32964a <=( a32963a  and  a32960a );
 a32965a <=( a32964a  and  a32957a );
 a32969a <=( A234  and  A232 );
 a32970a <=( A202  and  a32969a );
 a32973a <=( (not A266)  and  (not A265) );
 a32976a <=( (not A269)  and  A268 );
 a32977a <=( a32976a  and  a32973a );
 a32978a <=( a32977a  and  a32970a );
 a32982a <=( (not A167)  and  A168 );
 a32983a <=( A169  and  a32982a );
 a32986a <=( A199  and  A166 );
 a32989a <=( (not A201)  and  (not A200) );
 a32990a <=( a32989a  and  a32986a );
 a32991a <=( a32990a  and  a32983a );
 a32995a <=( A234  and  A233 );
 a32996a <=( A202  and  a32995a );
 a32999a <=( A299  and  A298 );
 a33002a <=( (not A302)  and  A301 );
 a33003a <=( a33002a  and  a32999a );
 a33004a <=( a33003a  and  a32996a );
 a33008a <=( (not A167)  and  A168 );
 a33009a <=( A169  and  a33008a );
 a33012a <=( A199  and  A166 );
 a33015a <=( (not A201)  and  (not A200) );
 a33016a <=( a33015a  and  a33012a );
 a33017a <=( a33016a  and  a33009a );
 a33021a <=( A234  and  A233 );
 a33022a <=( A202  and  a33021a );
 a33025a <=( (not A299)  and  A298 );
 a33028a <=( A302  and  (not A301) );
 a33029a <=( a33028a  and  a33025a );
 a33030a <=( a33029a  and  a33022a );
 a33034a <=( (not A167)  and  A168 );
 a33035a <=( A169  and  a33034a );
 a33038a <=( A199  and  A166 );
 a33041a <=( (not A201)  and  (not A200) );
 a33042a <=( a33041a  and  a33038a );
 a33043a <=( a33042a  and  a33035a );
 a33047a <=( A234  and  A233 );
 a33048a <=( A202  and  a33047a );
 a33051a <=( A299  and  (not A298) );
 a33054a <=( A302  and  (not A301) );
 a33055a <=( a33054a  and  a33051a );
 a33056a <=( a33055a  and  a33048a );
 a33060a <=( (not A167)  and  A168 );
 a33061a <=( A169  and  a33060a );
 a33064a <=( A199  and  A166 );
 a33067a <=( (not A201)  and  (not A200) );
 a33068a <=( a33067a  and  a33064a );
 a33069a <=( a33068a  and  a33061a );
 a33073a <=( A234  and  A233 );
 a33074a <=( A202  and  a33073a );
 a33077a <=( (not A299)  and  (not A298) );
 a33080a <=( (not A302)  and  A301 );
 a33081a <=( a33080a  and  a33077a );
 a33082a <=( a33081a  and  a33074a );
 a33086a <=( (not A167)  and  A168 );
 a33087a <=( A169  and  a33086a );
 a33090a <=( A199  and  A166 );
 a33093a <=( (not A201)  and  (not A200) );
 a33094a <=( a33093a  and  a33090a );
 a33095a <=( a33094a  and  a33087a );
 a33099a <=( A234  and  A233 );
 a33100a <=( A202  and  a33099a );
 a33103a <=( A266  and  A265 );
 a33106a <=( (not A269)  and  A268 );
 a33107a <=( a33106a  and  a33103a );
 a33108a <=( a33107a  and  a33100a );
 a33112a <=( (not A167)  and  A168 );
 a33113a <=( A169  and  a33112a );
 a33116a <=( A199  and  A166 );
 a33119a <=( (not A201)  and  (not A200) );
 a33120a <=( a33119a  and  a33116a );
 a33121a <=( a33120a  and  a33113a );
 a33125a <=( A234  and  A233 );
 a33126a <=( A202  and  a33125a );
 a33129a <=( A266  and  (not A265) );
 a33132a <=( A269  and  (not A268) );
 a33133a <=( a33132a  and  a33129a );
 a33134a <=( a33133a  and  a33126a );
 a33138a <=( (not A167)  and  A168 );
 a33139a <=( A169  and  a33138a );
 a33142a <=( A199  and  A166 );
 a33145a <=( (not A201)  and  (not A200) );
 a33146a <=( a33145a  and  a33142a );
 a33147a <=( a33146a  and  a33139a );
 a33151a <=( A234  and  A233 );
 a33152a <=( A202  and  a33151a );
 a33155a <=( (not A266)  and  A265 );
 a33158a <=( A269  and  (not A268) );
 a33159a <=( a33158a  and  a33155a );
 a33160a <=( a33159a  and  a33152a );
 a33164a <=( (not A167)  and  A168 );
 a33165a <=( A169  and  a33164a );
 a33168a <=( A199  and  A166 );
 a33171a <=( (not A201)  and  (not A200) );
 a33172a <=( a33171a  and  a33168a );
 a33173a <=( a33172a  and  a33165a );
 a33177a <=( A234  and  A233 );
 a33178a <=( A202  and  a33177a );
 a33181a <=( (not A266)  and  (not A265) );
 a33184a <=( (not A269)  and  A268 );
 a33185a <=( a33184a  and  a33181a );
 a33186a <=( a33185a  and  a33178a );
 a33190a <=( (not A167)  and  A168 );
 a33191a <=( A169  and  a33190a );
 a33194a <=( A199  and  A166 );
 a33197a <=( (not A201)  and  (not A200) );
 a33198a <=( a33197a  and  a33194a );
 a33199a <=( a33198a  and  a33191a );
 a33203a <=( A233  and  A232 );
 a33204a <=( A202  and  a33203a );
 a33207a <=( (not A236)  and  A235 );
 a33210a <=( A300  and  A299 );
 a33211a <=( a33210a  and  a33207a );
 a33212a <=( a33211a  and  a33204a );
 a33216a <=( (not A167)  and  A168 );
 a33217a <=( A169  and  a33216a );
 a33220a <=( A199  and  A166 );
 a33223a <=( (not A201)  and  (not A200) );
 a33224a <=( a33223a  and  a33220a );
 a33225a <=( a33224a  and  a33217a );
 a33229a <=( A233  and  A232 );
 a33230a <=( A202  and  a33229a );
 a33233a <=( (not A236)  and  A235 );
 a33236a <=( A300  and  A298 );
 a33237a <=( a33236a  and  a33233a );
 a33238a <=( a33237a  and  a33230a );
 a33242a <=( (not A167)  and  A168 );
 a33243a <=( A169  and  a33242a );
 a33246a <=( A199  and  A166 );
 a33249a <=( (not A201)  and  (not A200) );
 a33250a <=( a33249a  and  a33246a );
 a33251a <=( a33250a  and  a33243a );
 a33255a <=( A233  and  A232 );
 a33256a <=( A202  and  a33255a );
 a33259a <=( (not A236)  and  A235 );
 a33262a <=( A267  and  A265 );
 a33263a <=( a33262a  and  a33259a );
 a33264a <=( a33263a  and  a33256a );
 a33268a <=( (not A167)  and  A168 );
 a33269a <=( A169  and  a33268a );
 a33272a <=( A199  and  A166 );
 a33275a <=( (not A201)  and  (not A200) );
 a33276a <=( a33275a  and  a33272a );
 a33277a <=( a33276a  and  a33269a );
 a33281a <=( A233  and  A232 );
 a33282a <=( A202  and  a33281a );
 a33285a <=( (not A236)  and  A235 );
 a33288a <=( A267  and  A266 );
 a33289a <=( a33288a  and  a33285a );
 a33290a <=( a33289a  and  a33282a );
 a33294a <=( (not A167)  and  A168 );
 a33295a <=( A169  and  a33294a );
 a33298a <=( A199  and  A166 );
 a33301a <=( (not A201)  and  (not A200) );
 a33302a <=( a33301a  and  a33298a );
 a33303a <=( a33302a  and  a33295a );
 a33307a <=( A233  and  (not A232) );
 a33308a <=( A202  and  a33307a );
 a33311a <=( A236  and  (not A235) );
 a33314a <=( A300  and  A299 );
 a33315a <=( a33314a  and  a33311a );
 a33316a <=( a33315a  and  a33308a );
 a33320a <=( (not A167)  and  A168 );
 a33321a <=( A169  and  a33320a );
 a33324a <=( A199  and  A166 );
 a33327a <=( (not A201)  and  (not A200) );
 a33328a <=( a33327a  and  a33324a );
 a33329a <=( a33328a  and  a33321a );
 a33333a <=( A233  and  (not A232) );
 a33334a <=( A202  and  a33333a );
 a33337a <=( A236  and  (not A235) );
 a33340a <=( A300  and  A298 );
 a33341a <=( a33340a  and  a33337a );
 a33342a <=( a33341a  and  a33334a );
 a33346a <=( (not A167)  and  A168 );
 a33347a <=( A169  and  a33346a );
 a33350a <=( A199  and  A166 );
 a33353a <=( (not A201)  and  (not A200) );
 a33354a <=( a33353a  and  a33350a );
 a33355a <=( a33354a  and  a33347a );
 a33359a <=( A233  and  (not A232) );
 a33360a <=( A202  and  a33359a );
 a33363a <=( A236  and  (not A235) );
 a33366a <=( A267  and  A265 );
 a33367a <=( a33366a  and  a33363a );
 a33368a <=( a33367a  and  a33360a );
 a33372a <=( (not A167)  and  A168 );
 a33373a <=( A169  and  a33372a );
 a33376a <=( A199  and  A166 );
 a33379a <=( (not A201)  and  (not A200) );
 a33380a <=( a33379a  and  a33376a );
 a33381a <=( a33380a  and  a33373a );
 a33385a <=( A233  and  (not A232) );
 a33386a <=( A202  and  a33385a );
 a33389a <=( A236  and  (not A235) );
 a33392a <=( A267  and  A266 );
 a33393a <=( a33392a  and  a33389a );
 a33394a <=( a33393a  and  a33386a );
 a33398a <=( (not A167)  and  A168 );
 a33399a <=( A169  and  a33398a );
 a33402a <=( A199  and  A166 );
 a33405a <=( (not A201)  and  (not A200) );
 a33406a <=( a33405a  and  a33402a );
 a33407a <=( a33406a  and  a33399a );
 a33411a <=( (not A233)  and  A232 );
 a33412a <=( A202  and  a33411a );
 a33415a <=( A236  and  (not A235) );
 a33418a <=( A300  and  A299 );
 a33419a <=( a33418a  and  a33415a );
 a33420a <=( a33419a  and  a33412a );
 a33424a <=( (not A167)  and  A168 );
 a33425a <=( A169  and  a33424a );
 a33428a <=( A199  and  A166 );
 a33431a <=( (not A201)  and  (not A200) );
 a33432a <=( a33431a  and  a33428a );
 a33433a <=( a33432a  and  a33425a );
 a33437a <=( (not A233)  and  A232 );
 a33438a <=( A202  and  a33437a );
 a33441a <=( A236  and  (not A235) );
 a33444a <=( A300  and  A298 );
 a33445a <=( a33444a  and  a33441a );
 a33446a <=( a33445a  and  a33438a );
 a33450a <=( (not A167)  and  A168 );
 a33451a <=( A169  and  a33450a );
 a33454a <=( A199  and  A166 );
 a33457a <=( (not A201)  and  (not A200) );
 a33458a <=( a33457a  and  a33454a );
 a33459a <=( a33458a  and  a33451a );
 a33463a <=( (not A233)  and  A232 );
 a33464a <=( A202  and  a33463a );
 a33467a <=( A236  and  (not A235) );
 a33470a <=( A267  and  A265 );
 a33471a <=( a33470a  and  a33467a );
 a33472a <=( a33471a  and  a33464a );
 a33476a <=( (not A167)  and  A168 );
 a33477a <=( A169  and  a33476a );
 a33480a <=( A199  and  A166 );
 a33483a <=( (not A201)  and  (not A200) );
 a33484a <=( a33483a  and  a33480a );
 a33485a <=( a33484a  and  a33477a );
 a33489a <=( (not A233)  and  A232 );
 a33490a <=( A202  and  a33489a );
 a33493a <=( A236  and  (not A235) );
 a33496a <=( A267  and  A266 );
 a33497a <=( a33496a  and  a33493a );
 a33498a <=( a33497a  and  a33490a );
 a33502a <=( (not A167)  and  A168 );
 a33503a <=( A169  and  a33502a );
 a33506a <=( A199  and  A166 );
 a33509a <=( (not A201)  and  (not A200) );
 a33510a <=( a33509a  and  a33506a );
 a33511a <=( a33510a  and  a33503a );
 a33515a <=( (not A233)  and  (not A232) );
 a33516a <=( A202  and  a33515a );
 a33519a <=( (not A236)  and  A235 );
 a33522a <=( A300  and  A299 );
 a33523a <=( a33522a  and  a33519a );
 a33524a <=( a33523a  and  a33516a );
 a33528a <=( (not A167)  and  A168 );
 a33529a <=( A169  and  a33528a );
 a33532a <=( A199  and  A166 );
 a33535a <=( (not A201)  and  (not A200) );
 a33536a <=( a33535a  and  a33532a );
 a33537a <=( a33536a  and  a33529a );
 a33541a <=( (not A233)  and  (not A232) );
 a33542a <=( A202  and  a33541a );
 a33545a <=( (not A236)  and  A235 );
 a33548a <=( A300  and  A298 );
 a33549a <=( a33548a  and  a33545a );
 a33550a <=( a33549a  and  a33542a );
 a33554a <=( (not A167)  and  A168 );
 a33555a <=( A169  and  a33554a );
 a33558a <=( A199  and  A166 );
 a33561a <=( (not A201)  and  (not A200) );
 a33562a <=( a33561a  and  a33558a );
 a33563a <=( a33562a  and  a33555a );
 a33567a <=( (not A233)  and  (not A232) );
 a33568a <=( A202  and  a33567a );
 a33571a <=( (not A236)  and  A235 );
 a33574a <=( A267  and  A265 );
 a33575a <=( a33574a  and  a33571a );
 a33576a <=( a33575a  and  a33568a );
 a33580a <=( (not A167)  and  A168 );
 a33581a <=( A169  and  a33580a );
 a33584a <=( A199  and  A166 );
 a33587a <=( (not A201)  and  (not A200) );
 a33588a <=( a33587a  and  a33584a );
 a33589a <=( a33588a  and  a33581a );
 a33593a <=( (not A233)  and  (not A232) );
 a33594a <=( A202  and  a33593a );
 a33597a <=( (not A236)  and  A235 );
 a33600a <=( A267  and  A266 );
 a33601a <=( a33600a  and  a33597a );
 a33602a <=( a33601a  and  a33594a );
 a33606a <=( (not A167)  and  A168 );
 a33607a <=( A169  and  a33606a );
 a33610a <=( A199  and  A166 );
 a33613a <=( (not A201)  and  (not A200) );
 a33614a <=( a33613a  and  a33610a );
 a33615a <=( a33614a  and  a33607a );
 a33619a <=( A234  and  A232 );
 a33620a <=( (not A203)  and  a33619a );
 a33623a <=( A299  and  A298 );
 a33626a <=( (not A302)  and  A301 );
 a33627a <=( a33626a  and  a33623a );
 a33628a <=( a33627a  and  a33620a );
 a33632a <=( (not A167)  and  A168 );
 a33633a <=( A169  and  a33632a );
 a33636a <=( A199  and  A166 );
 a33639a <=( (not A201)  and  (not A200) );
 a33640a <=( a33639a  and  a33636a );
 a33641a <=( a33640a  and  a33633a );
 a33645a <=( A234  and  A232 );
 a33646a <=( (not A203)  and  a33645a );
 a33649a <=( (not A299)  and  A298 );
 a33652a <=( A302  and  (not A301) );
 a33653a <=( a33652a  and  a33649a );
 a33654a <=( a33653a  and  a33646a );
 a33658a <=( (not A167)  and  A168 );
 a33659a <=( A169  and  a33658a );
 a33662a <=( A199  and  A166 );
 a33665a <=( (not A201)  and  (not A200) );
 a33666a <=( a33665a  and  a33662a );
 a33667a <=( a33666a  and  a33659a );
 a33671a <=( A234  and  A232 );
 a33672a <=( (not A203)  and  a33671a );
 a33675a <=( A299  and  (not A298) );
 a33678a <=( A302  and  (not A301) );
 a33679a <=( a33678a  and  a33675a );
 a33680a <=( a33679a  and  a33672a );
 a33684a <=( (not A167)  and  A168 );
 a33685a <=( A169  and  a33684a );
 a33688a <=( A199  and  A166 );
 a33691a <=( (not A201)  and  (not A200) );
 a33692a <=( a33691a  and  a33688a );
 a33693a <=( a33692a  and  a33685a );
 a33697a <=( A234  and  A232 );
 a33698a <=( (not A203)  and  a33697a );
 a33701a <=( (not A299)  and  (not A298) );
 a33704a <=( (not A302)  and  A301 );
 a33705a <=( a33704a  and  a33701a );
 a33706a <=( a33705a  and  a33698a );
 a33710a <=( (not A167)  and  A168 );
 a33711a <=( A169  and  a33710a );
 a33714a <=( A199  and  A166 );
 a33717a <=( (not A201)  and  (not A200) );
 a33718a <=( a33717a  and  a33714a );
 a33719a <=( a33718a  and  a33711a );
 a33723a <=( A234  and  A232 );
 a33724a <=( (not A203)  and  a33723a );
 a33727a <=( A266  and  A265 );
 a33730a <=( (not A269)  and  A268 );
 a33731a <=( a33730a  and  a33727a );
 a33732a <=( a33731a  and  a33724a );
 a33736a <=( (not A167)  and  A168 );
 a33737a <=( A169  and  a33736a );
 a33740a <=( A199  and  A166 );
 a33743a <=( (not A201)  and  (not A200) );
 a33744a <=( a33743a  and  a33740a );
 a33745a <=( a33744a  and  a33737a );
 a33749a <=( A234  and  A232 );
 a33750a <=( (not A203)  and  a33749a );
 a33753a <=( A266  and  (not A265) );
 a33756a <=( A269  and  (not A268) );
 a33757a <=( a33756a  and  a33753a );
 a33758a <=( a33757a  and  a33750a );
 a33762a <=( (not A167)  and  A168 );
 a33763a <=( A169  and  a33762a );
 a33766a <=( A199  and  A166 );
 a33769a <=( (not A201)  and  (not A200) );
 a33770a <=( a33769a  and  a33766a );
 a33771a <=( a33770a  and  a33763a );
 a33775a <=( A234  and  A232 );
 a33776a <=( (not A203)  and  a33775a );
 a33779a <=( (not A266)  and  A265 );
 a33782a <=( A269  and  (not A268) );
 a33783a <=( a33782a  and  a33779a );
 a33784a <=( a33783a  and  a33776a );
 a33788a <=( (not A167)  and  A168 );
 a33789a <=( A169  and  a33788a );
 a33792a <=( A199  and  A166 );
 a33795a <=( (not A201)  and  (not A200) );
 a33796a <=( a33795a  and  a33792a );
 a33797a <=( a33796a  and  a33789a );
 a33801a <=( A234  and  A232 );
 a33802a <=( (not A203)  and  a33801a );
 a33805a <=( (not A266)  and  (not A265) );
 a33808a <=( (not A269)  and  A268 );
 a33809a <=( a33808a  and  a33805a );
 a33810a <=( a33809a  and  a33802a );
 a33814a <=( (not A167)  and  A168 );
 a33815a <=( A169  and  a33814a );
 a33818a <=( A199  and  A166 );
 a33821a <=( (not A201)  and  (not A200) );
 a33822a <=( a33821a  and  a33818a );
 a33823a <=( a33822a  and  a33815a );
 a33827a <=( A234  and  A233 );
 a33828a <=( (not A203)  and  a33827a );
 a33831a <=( A299  and  A298 );
 a33834a <=( (not A302)  and  A301 );
 a33835a <=( a33834a  and  a33831a );
 a33836a <=( a33835a  and  a33828a );
 a33840a <=( (not A167)  and  A168 );
 a33841a <=( A169  and  a33840a );
 a33844a <=( A199  and  A166 );
 a33847a <=( (not A201)  and  (not A200) );
 a33848a <=( a33847a  and  a33844a );
 a33849a <=( a33848a  and  a33841a );
 a33853a <=( A234  and  A233 );
 a33854a <=( (not A203)  and  a33853a );
 a33857a <=( (not A299)  and  A298 );
 a33860a <=( A302  and  (not A301) );
 a33861a <=( a33860a  and  a33857a );
 a33862a <=( a33861a  and  a33854a );
 a33866a <=( (not A167)  and  A168 );
 a33867a <=( A169  and  a33866a );
 a33870a <=( A199  and  A166 );
 a33873a <=( (not A201)  and  (not A200) );
 a33874a <=( a33873a  and  a33870a );
 a33875a <=( a33874a  and  a33867a );
 a33879a <=( A234  and  A233 );
 a33880a <=( (not A203)  and  a33879a );
 a33883a <=( A299  and  (not A298) );
 a33886a <=( A302  and  (not A301) );
 a33887a <=( a33886a  and  a33883a );
 a33888a <=( a33887a  and  a33880a );
 a33892a <=( (not A167)  and  A168 );
 a33893a <=( A169  and  a33892a );
 a33896a <=( A199  and  A166 );
 a33899a <=( (not A201)  and  (not A200) );
 a33900a <=( a33899a  and  a33896a );
 a33901a <=( a33900a  and  a33893a );
 a33905a <=( A234  and  A233 );
 a33906a <=( (not A203)  and  a33905a );
 a33909a <=( (not A299)  and  (not A298) );
 a33912a <=( (not A302)  and  A301 );
 a33913a <=( a33912a  and  a33909a );
 a33914a <=( a33913a  and  a33906a );
 a33918a <=( (not A167)  and  A168 );
 a33919a <=( A169  and  a33918a );
 a33922a <=( A199  and  A166 );
 a33925a <=( (not A201)  and  (not A200) );
 a33926a <=( a33925a  and  a33922a );
 a33927a <=( a33926a  and  a33919a );
 a33931a <=( A234  and  A233 );
 a33932a <=( (not A203)  and  a33931a );
 a33935a <=( A266  and  A265 );
 a33938a <=( (not A269)  and  A268 );
 a33939a <=( a33938a  and  a33935a );
 a33940a <=( a33939a  and  a33932a );
 a33944a <=( (not A167)  and  A168 );
 a33945a <=( A169  and  a33944a );
 a33948a <=( A199  and  A166 );
 a33951a <=( (not A201)  and  (not A200) );
 a33952a <=( a33951a  and  a33948a );
 a33953a <=( a33952a  and  a33945a );
 a33957a <=( A234  and  A233 );
 a33958a <=( (not A203)  and  a33957a );
 a33961a <=( A266  and  (not A265) );
 a33964a <=( A269  and  (not A268) );
 a33965a <=( a33964a  and  a33961a );
 a33966a <=( a33965a  and  a33958a );
 a33970a <=( (not A167)  and  A168 );
 a33971a <=( A169  and  a33970a );
 a33974a <=( A199  and  A166 );
 a33977a <=( (not A201)  and  (not A200) );
 a33978a <=( a33977a  and  a33974a );
 a33979a <=( a33978a  and  a33971a );
 a33983a <=( A234  and  A233 );
 a33984a <=( (not A203)  and  a33983a );
 a33987a <=( (not A266)  and  A265 );
 a33990a <=( A269  and  (not A268) );
 a33991a <=( a33990a  and  a33987a );
 a33992a <=( a33991a  and  a33984a );
 a33996a <=( (not A167)  and  A168 );
 a33997a <=( A169  and  a33996a );
 a34000a <=( A199  and  A166 );
 a34003a <=( (not A201)  and  (not A200) );
 a34004a <=( a34003a  and  a34000a );
 a34005a <=( a34004a  and  a33997a );
 a34009a <=( A234  and  A233 );
 a34010a <=( (not A203)  and  a34009a );
 a34013a <=( (not A266)  and  (not A265) );
 a34016a <=( (not A269)  and  A268 );
 a34017a <=( a34016a  and  a34013a );
 a34018a <=( a34017a  and  a34010a );
 a34022a <=( (not A167)  and  A168 );
 a34023a <=( A169  and  a34022a );
 a34026a <=( A199  and  A166 );
 a34029a <=( (not A201)  and  (not A200) );
 a34030a <=( a34029a  and  a34026a );
 a34031a <=( a34030a  and  a34023a );
 a34035a <=( A233  and  A232 );
 a34036a <=( (not A203)  and  a34035a );
 a34039a <=( (not A236)  and  A235 );
 a34042a <=( A300  and  A299 );
 a34043a <=( a34042a  and  a34039a );
 a34044a <=( a34043a  and  a34036a );
 a34048a <=( (not A167)  and  A168 );
 a34049a <=( A169  and  a34048a );
 a34052a <=( A199  and  A166 );
 a34055a <=( (not A201)  and  (not A200) );
 a34056a <=( a34055a  and  a34052a );
 a34057a <=( a34056a  and  a34049a );
 a34061a <=( A233  and  A232 );
 a34062a <=( (not A203)  and  a34061a );
 a34065a <=( (not A236)  and  A235 );
 a34068a <=( A300  and  A298 );
 a34069a <=( a34068a  and  a34065a );
 a34070a <=( a34069a  and  a34062a );
 a34074a <=( (not A167)  and  A168 );
 a34075a <=( A169  and  a34074a );
 a34078a <=( A199  and  A166 );
 a34081a <=( (not A201)  and  (not A200) );
 a34082a <=( a34081a  and  a34078a );
 a34083a <=( a34082a  and  a34075a );
 a34087a <=( A233  and  A232 );
 a34088a <=( (not A203)  and  a34087a );
 a34091a <=( (not A236)  and  A235 );
 a34094a <=( A267  and  A265 );
 a34095a <=( a34094a  and  a34091a );
 a34096a <=( a34095a  and  a34088a );
 a34100a <=( (not A167)  and  A168 );
 a34101a <=( A169  and  a34100a );
 a34104a <=( A199  and  A166 );
 a34107a <=( (not A201)  and  (not A200) );
 a34108a <=( a34107a  and  a34104a );
 a34109a <=( a34108a  and  a34101a );
 a34113a <=( A233  and  A232 );
 a34114a <=( (not A203)  and  a34113a );
 a34117a <=( (not A236)  and  A235 );
 a34120a <=( A267  and  A266 );
 a34121a <=( a34120a  and  a34117a );
 a34122a <=( a34121a  and  a34114a );
 a34126a <=( (not A167)  and  A168 );
 a34127a <=( A169  and  a34126a );
 a34130a <=( A199  and  A166 );
 a34133a <=( (not A201)  and  (not A200) );
 a34134a <=( a34133a  and  a34130a );
 a34135a <=( a34134a  and  a34127a );
 a34139a <=( A233  and  (not A232) );
 a34140a <=( (not A203)  and  a34139a );
 a34143a <=( A236  and  (not A235) );
 a34146a <=( A300  and  A299 );
 a34147a <=( a34146a  and  a34143a );
 a34148a <=( a34147a  and  a34140a );
 a34152a <=( (not A167)  and  A168 );
 a34153a <=( A169  and  a34152a );
 a34156a <=( A199  and  A166 );
 a34159a <=( (not A201)  and  (not A200) );
 a34160a <=( a34159a  and  a34156a );
 a34161a <=( a34160a  and  a34153a );
 a34165a <=( A233  and  (not A232) );
 a34166a <=( (not A203)  and  a34165a );
 a34169a <=( A236  and  (not A235) );
 a34172a <=( A300  and  A298 );
 a34173a <=( a34172a  and  a34169a );
 a34174a <=( a34173a  and  a34166a );
 a34178a <=( (not A167)  and  A168 );
 a34179a <=( A169  and  a34178a );
 a34182a <=( A199  and  A166 );
 a34185a <=( (not A201)  and  (not A200) );
 a34186a <=( a34185a  and  a34182a );
 a34187a <=( a34186a  and  a34179a );
 a34191a <=( A233  and  (not A232) );
 a34192a <=( (not A203)  and  a34191a );
 a34195a <=( A236  and  (not A235) );
 a34198a <=( A267  and  A265 );
 a34199a <=( a34198a  and  a34195a );
 a34200a <=( a34199a  and  a34192a );
 a34204a <=( (not A167)  and  A168 );
 a34205a <=( A169  and  a34204a );
 a34208a <=( A199  and  A166 );
 a34211a <=( (not A201)  and  (not A200) );
 a34212a <=( a34211a  and  a34208a );
 a34213a <=( a34212a  and  a34205a );
 a34217a <=( A233  and  (not A232) );
 a34218a <=( (not A203)  and  a34217a );
 a34221a <=( A236  and  (not A235) );
 a34224a <=( A267  and  A266 );
 a34225a <=( a34224a  and  a34221a );
 a34226a <=( a34225a  and  a34218a );
 a34230a <=( (not A167)  and  A168 );
 a34231a <=( A169  and  a34230a );
 a34234a <=( A199  and  A166 );
 a34237a <=( (not A201)  and  (not A200) );
 a34238a <=( a34237a  and  a34234a );
 a34239a <=( a34238a  and  a34231a );
 a34243a <=( (not A233)  and  A232 );
 a34244a <=( (not A203)  and  a34243a );
 a34247a <=( A236  and  (not A235) );
 a34250a <=( A300  and  A299 );
 a34251a <=( a34250a  and  a34247a );
 a34252a <=( a34251a  and  a34244a );
 a34256a <=( (not A167)  and  A168 );
 a34257a <=( A169  and  a34256a );
 a34260a <=( A199  and  A166 );
 a34263a <=( (not A201)  and  (not A200) );
 a34264a <=( a34263a  and  a34260a );
 a34265a <=( a34264a  and  a34257a );
 a34269a <=( (not A233)  and  A232 );
 a34270a <=( (not A203)  and  a34269a );
 a34273a <=( A236  and  (not A235) );
 a34276a <=( A300  and  A298 );
 a34277a <=( a34276a  and  a34273a );
 a34278a <=( a34277a  and  a34270a );
 a34282a <=( (not A167)  and  A168 );
 a34283a <=( A169  and  a34282a );
 a34286a <=( A199  and  A166 );
 a34289a <=( (not A201)  and  (not A200) );
 a34290a <=( a34289a  and  a34286a );
 a34291a <=( a34290a  and  a34283a );
 a34295a <=( (not A233)  and  A232 );
 a34296a <=( (not A203)  and  a34295a );
 a34299a <=( A236  and  (not A235) );
 a34302a <=( A267  and  A265 );
 a34303a <=( a34302a  and  a34299a );
 a34304a <=( a34303a  and  a34296a );
 a34308a <=( (not A167)  and  A168 );
 a34309a <=( A169  and  a34308a );
 a34312a <=( A199  and  A166 );
 a34315a <=( (not A201)  and  (not A200) );
 a34316a <=( a34315a  and  a34312a );
 a34317a <=( a34316a  and  a34309a );
 a34321a <=( (not A233)  and  A232 );
 a34322a <=( (not A203)  and  a34321a );
 a34325a <=( A236  and  (not A235) );
 a34328a <=( A267  and  A266 );
 a34329a <=( a34328a  and  a34325a );
 a34330a <=( a34329a  and  a34322a );
 a34334a <=( (not A167)  and  A168 );
 a34335a <=( A169  and  a34334a );
 a34338a <=( A199  and  A166 );
 a34341a <=( (not A201)  and  (not A200) );
 a34342a <=( a34341a  and  a34338a );
 a34343a <=( a34342a  and  a34335a );
 a34347a <=( (not A233)  and  (not A232) );
 a34348a <=( (not A203)  and  a34347a );
 a34351a <=( (not A236)  and  A235 );
 a34354a <=( A300  and  A299 );
 a34355a <=( a34354a  and  a34351a );
 a34356a <=( a34355a  and  a34348a );
 a34360a <=( (not A167)  and  A168 );
 a34361a <=( A169  and  a34360a );
 a34364a <=( A199  and  A166 );
 a34367a <=( (not A201)  and  (not A200) );
 a34368a <=( a34367a  and  a34364a );
 a34369a <=( a34368a  and  a34361a );
 a34373a <=( (not A233)  and  (not A232) );
 a34374a <=( (not A203)  and  a34373a );
 a34377a <=( (not A236)  and  A235 );
 a34380a <=( A300  and  A298 );
 a34381a <=( a34380a  and  a34377a );
 a34382a <=( a34381a  and  a34374a );
 a34386a <=( (not A167)  and  A168 );
 a34387a <=( A169  and  a34386a );
 a34390a <=( A199  and  A166 );
 a34393a <=( (not A201)  and  (not A200) );
 a34394a <=( a34393a  and  a34390a );
 a34395a <=( a34394a  and  a34387a );
 a34399a <=( (not A233)  and  (not A232) );
 a34400a <=( (not A203)  and  a34399a );
 a34403a <=( (not A236)  and  A235 );
 a34406a <=( A267  and  A265 );
 a34407a <=( a34406a  and  a34403a );
 a34408a <=( a34407a  and  a34400a );
 a34412a <=( (not A167)  and  A168 );
 a34413a <=( A169  and  a34412a );
 a34416a <=( A199  and  A166 );
 a34419a <=( (not A201)  and  (not A200) );
 a34420a <=( a34419a  and  a34416a );
 a34421a <=( a34420a  and  a34413a );
 a34425a <=( (not A233)  and  (not A232) );
 a34426a <=( (not A203)  and  a34425a );
 a34429a <=( (not A236)  and  A235 );
 a34432a <=( A267  and  A266 );
 a34433a <=( a34432a  and  a34429a );
 a34434a <=( a34433a  and  a34426a );
 a34438a <=( (not A167)  and  A168 );
 a34439a <=( A170  and  a34438a );
 a34442a <=( (not A199)  and  A166 );
 a34445a <=( (not A202)  and  (not A200) );
 a34446a <=( a34445a  and  a34442a );
 a34447a <=( a34446a  and  a34439a );
 a34450a <=( A233  and  A232 );
 a34453a <=( (not A236)  and  A235 );
 a34454a <=( a34453a  and  a34450a );
 a34457a <=( A299  and  A298 );
 a34460a <=( (not A302)  and  A301 );
 a34461a <=( a34460a  and  a34457a );
 a34462a <=( a34461a  and  a34454a );
 a34466a <=( (not A167)  and  A168 );
 a34467a <=( A170  and  a34466a );
 a34470a <=( (not A199)  and  A166 );
 a34473a <=( (not A202)  and  (not A200) );
 a34474a <=( a34473a  and  a34470a );
 a34475a <=( a34474a  and  a34467a );
 a34478a <=( A233  and  A232 );
 a34481a <=( (not A236)  and  A235 );
 a34482a <=( a34481a  and  a34478a );
 a34485a <=( (not A299)  and  A298 );
 a34488a <=( A302  and  (not A301) );
 a34489a <=( a34488a  and  a34485a );
 a34490a <=( a34489a  and  a34482a );
 a34494a <=( (not A167)  and  A168 );
 a34495a <=( A170  and  a34494a );
 a34498a <=( (not A199)  and  A166 );
 a34501a <=( (not A202)  and  (not A200) );
 a34502a <=( a34501a  and  a34498a );
 a34503a <=( a34502a  and  a34495a );
 a34506a <=( A233  and  A232 );
 a34509a <=( (not A236)  and  A235 );
 a34510a <=( a34509a  and  a34506a );
 a34513a <=( A299  and  (not A298) );
 a34516a <=( A302  and  (not A301) );
 a34517a <=( a34516a  and  a34513a );
 a34518a <=( a34517a  and  a34510a );
 a34522a <=( (not A167)  and  A168 );
 a34523a <=( A170  and  a34522a );
 a34526a <=( (not A199)  and  A166 );
 a34529a <=( (not A202)  and  (not A200) );
 a34530a <=( a34529a  and  a34526a );
 a34531a <=( a34530a  and  a34523a );
 a34534a <=( A233  and  A232 );
 a34537a <=( (not A236)  and  A235 );
 a34538a <=( a34537a  and  a34534a );
 a34541a <=( (not A299)  and  (not A298) );
 a34544a <=( (not A302)  and  A301 );
 a34545a <=( a34544a  and  a34541a );
 a34546a <=( a34545a  and  a34538a );
 a34550a <=( (not A167)  and  A168 );
 a34551a <=( A170  and  a34550a );
 a34554a <=( (not A199)  and  A166 );
 a34557a <=( (not A202)  and  (not A200) );
 a34558a <=( a34557a  and  a34554a );
 a34559a <=( a34558a  and  a34551a );
 a34562a <=( A233  and  A232 );
 a34565a <=( (not A236)  and  A235 );
 a34566a <=( a34565a  and  a34562a );
 a34569a <=( A266  and  A265 );
 a34572a <=( (not A269)  and  A268 );
 a34573a <=( a34572a  and  a34569a );
 a34574a <=( a34573a  and  a34566a );
 a34578a <=( (not A167)  and  A168 );
 a34579a <=( A170  and  a34578a );
 a34582a <=( (not A199)  and  A166 );
 a34585a <=( (not A202)  and  (not A200) );
 a34586a <=( a34585a  and  a34582a );
 a34587a <=( a34586a  and  a34579a );
 a34590a <=( A233  and  A232 );
 a34593a <=( (not A236)  and  A235 );
 a34594a <=( a34593a  and  a34590a );
 a34597a <=( A266  and  (not A265) );
 a34600a <=( A269  and  (not A268) );
 a34601a <=( a34600a  and  a34597a );
 a34602a <=( a34601a  and  a34594a );
 a34606a <=( (not A167)  and  A168 );
 a34607a <=( A170  and  a34606a );
 a34610a <=( (not A199)  and  A166 );
 a34613a <=( (not A202)  and  (not A200) );
 a34614a <=( a34613a  and  a34610a );
 a34615a <=( a34614a  and  a34607a );
 a34618a <=( A233  and  A232 );
 a34621a <=( (not A236)  and  A235 );
 a34622a <=( a34621a  and  a34618a );
 a34625a <=( (not A266)  and  A265 );
 a34628a <=( A269  and  (not A268) );
 a34629a <=( a34628a  and  a34625a );
 a34630a <=( a34629a  and  a34622a );
 a34634a <=( (not A167)  and  A168 );
 a34635a <=( A170  and  a34634a );
 a34638a <=( (not A199)  and  A166 );
 a34641a <=( (not A202)  and  (not A200) );
 a34642a <=( a34641a  and  a34638a );
 a34643a <=( a34642a  and  a34635a );
 a34646a <=( A233  and  A232 );
 a34649a <=( (not A236)  and  A235 );
 a34650a <=( a34649a  and  a34646a );
 a34653a <=( (not A266)  and  (not A265) );
 a34656a <=( (not A269)  and  A268 );
 a34657a <=( a34656a  and  a34653a );
 a34658a <=( a34657a  and  a34650a );
 a34662a <=( (not A167)  and  A168 );
 a34663a <=( A170  and  a34662a );
 a34666a <=( (not A199)  and  A166 );
 a34669a <=( (not A202)  and  (not A200) );
 a34670a <=( a34669a  and  a34666a );
 a34671a <=( a34670a  and  a34663a );
 a34674a <=( A233  and  (not A232) );
 a34677a <=( A236  and  (not A235) );
 a34678a <=( a34677a  and  a34674a );
 a34681a <=( A299  and  A298 );
 a34684a <=( (not A302)  and  A301 );
 a34685a <=( a34684a  and  a34681a );
 a34686a <=( a34685a  and  a34678a );
 a34690a <=( (not A167)  and  A168 );
 a34691a <=( A170  and  a34690a );
 a34694a <=( (not A199)  and  A166 );
 a34697a <=( (not A202)  and  (not A200) );
 a34698a <=( a34697a  and  a34694a );
 a34699a <=( a34698a  and  a34691a );
 a34702a <=( A233  and  (not A232) );
 a34705a <=( A236  and  (not A235) );
 a34706a <=( a34705a  and  a34702a );
 a34709a <=( (not A299)  and  A298 );
 a34712a <=( A302  and  (not A301) );
 a34713a <=( a34712a  and  a34709a );
 a34714a <=( a34713a  and  a34706a );
 a34718a <=( (not A167)  and  A168 );
 a34719a <=( A170  and  a34718a );
 a34722a <=( (not A199)  and  A166 );
 a34725a <=( (not A202)  and  (not A200) );
 a34726a <=( a34725a  and  a34722a );
 a34727a <=( a34726a  and  a34719a );
 a34730a <=( A233  and  (not A232) );
 a34733a <=( A236  and  (not A235) );
 a34734a <=( a34733a  and  a34730a );
 a34737a <=( A299  and  (not A298) );
 a34740a <=( A302  and  (not A301) );
 a34741a <=( a34740a  and  a34737a );
 a34742a <=( a34741a  and  a34734a );
 a34746a <=( (not A167)  and  A168 );
 a34747a <=( A170  and  a34746a );
 a34750a <=( (not A199)  and  A166 );
 a34753a <=( (not A202)  and  (not A200) );
 a34754a <=( a34753a  and  a34750a );
 a34755a <=( a34754a  and  a34747a );
 a34758a <=( A233  and  (not A232) );
 a34761a <=( A236  and  (not A235) );
 a34762a <=( a34761a  and  a34758a );
 a34765a <=( (not A299)  and  (not A298) );
 a34768a <=( (not A302)  and  A301 );
 a34769a <=( a34768a  and  a34765a );
 a34770a <=( a34769a  and  a34762a );
 a34774a <=( (not A167)  and  A168 );
 a34775a <=( A170  and  a34774a );
 a34778a <=( (not A199)  and  A166 );
 a34781a <=( (not A202)  and  (not A200) );
 a34782a <=( a34781a  and  a34778a );
 a34783a <=( a34782a  and  a34775a );
 a34786a <=( A233  and  (not A232) );
 a34789a <=( A236  and  (not A235) );
 a34790a <=( a34789a  and  a34786a );
 a34793a <=( A266  and  A265 );
 a34796a <=( (not A269)  and  A268 );
 a34797a <=( a34796a  and  a34793a );
 a34798a <=( a34797a  and  a34790a );
 a34802a <=( (not A167)  and  A168 );
 a34803a <=( A170  and  a34802a );
 a34806a <=( (not A199)  and  A166 );
 a34809a <=( (not A202)  and  (not A200) );
 a34810a <=( a34809a  and  a34806a );
 a34811a <=( a34810a  and  a34803a );
 a34814a <=( A233  and  (not A232) );
 a34817a <=( A236  and  (not A235) );
 a34818a <=( a34817a  and  a34814a );
 a34821a <=( A266  and  (not A265) );
 a34824a <=( A269  and  (not A268) );
 a34825a <=( a34824a  and  a34821a );
 a34826a <=( a34825a  and  a34818a );
 a34830a <=( (not A167)  and  A168 );
 a34831a <=( A170  and  a34830a );
 a34834a <=( (not A199)  and  A166 );
 a34837a <=( (not A202)  and  (not A200) );
 a34838a <=( a34837a  and  a34834a );
 a34839a <=( a34838a  and  a34831a );
 a34842a <=( A233  and  (not A232) );
 a34845a <=( A236  and  (not A235) );
 a34846a <=( a34845a  and  a34842a );
 a34849a <=( (not A266)  and  A265 );
 a34852a <=( A269  and  (not A268) );
 a34853a <=( a34852a  and  a34849a );
 a34854a <=( a34853a  and  a34846a );
 a34858a <=( (not A167)  and  A168 );
 a34859a <=( A170  and  a34858a );
 a34862a <=( (not A199)  and  A166 );
 a34865a <=( (not A202)  and  (not A200) );
 a34866a <=( a34865a  and  a34862a );
 a34867a <=( a34866a  and  a34859a );
 a34870a <=( A233  and  (not A232) );
 a34873a <=( A236  and  (not A235) );
 a34874a <=( a34873a  and  a34870a );
 a34877a <=( (not A266)  and  (not A265) );
 a34880a <=( (not A269)  and  A268 );
 a34881a <=( a34880a  and  a34877a );
 a34882a <=( a34881a  and  a34874a );
 a34886a <=( (not A167)  and  A168 );
 a34887a <=( A170  and  a34886a );
 a34890a <=( (not A199)  and  A166 );
 a34893a <=( (not A202)  and  (not A200) );
 a34894a <=( a34893a  and  a34890a );
 a34895a <=( a34894a  and  a34887a );
 a34898a <=( (not A233)  and  A232 );
 a34901a <=( A236  and  (not A235) );
 a34902a <=( a34901a  and  a34898a );
 a34905a <=( A299  and  A298 );
 a34908a <=( (not A302)  and  A301 );
 a34909a <=( a34908a  and  a34905a );
 a34910a <=( a34909a  and  a34902a );
 a34914a <=( (not A167)  and  A168 );
 a34915a <=( A170  and  a34914a );
 a34918a <=( (not A199)  and  A166 );
 a34921a <=( (not A202)  and  (not A200) );
 a34922a <=( a34921a  and  a34918a );
 a34923a <=( a34922a  and  a34915a );
 a34926a <=( (not A233)  and  A232 );
 a34929a <=( A236  and  (not A235) );
 a34930a <=( a34929a  and  a34926a );
 a34933a <=( (not A299)  and  A298 );
 a34936a <=( A302  and  (not A301) );
 a34937a <=( a34936a  and  a34933a );
 a34938a <=( a34937a  and  a34930a );
 a34942a <=( (not A167)  and  A168 );
 a34943a <=( A170  and  a34942a );
 a34946a <=( (not A199)  and  A166 );
 a34949a <=( (not A202)  and  (not A200) );
 a34950a <=( a34949a  and  a34946a );
 a34951a <=( a34950a  and  a34943a );
 a34954a <=( (not A233)  and  A232 );
 a34957a <=( A236  and  (not A235) );
 a34958a <=( a34957a  and  a34954a );
 a34961a <=( A299  and  (not A298) );
 a34964a <=( A302  and  (not A301) );
 a34965a <=( a34964a  and  a34961a );
 a34966a <=( a34965a  and  a34958a );
 a34970a <=( (not A167)  and  A168 );
 a34971a <=( A170  and  a34970a );
 a34974a <=( (not A199)  and  A166 );
 a34977a <=( (not A202)  and  (not A200) );
 a34978a <=( a34977a  and  a34974a );
 a34979a <=( a34978a  and  a34971a );
 a34982a <=( (not A233)  and  A232 );
 a34985a <=( A236  and  (not A235) );
 a34986a <=( a34985a  and  a34982a );
 a34989a <=( (not A299)  and  (not A298) );
 a34992a <=( (not A302)  and  A301 );
 a34993a <=( a34992a  and  a34989a );
 a34994a <=( a34993a  and  a34986a );
 a34998a <=( (not A167)  and  A168 );
 a34999a <=( A170  and  a34998a );
 a35002a <=( (not A199)  and  A166 );
 a35005a <=( (not A202)  and  (not A200) );
 a35006a <=( a35005a  and  a35002a );
 a35007a <=( a35006a  and  a34999a );
 a35010a <=( (not A233)  and  A232 );
 a35013a <=( A236  and  (not A235) );
 a35014a <=( a35013a  and  a35010a );
 a35017a <=( A266  and  A265 );
 a35020a <=( (not A269)  and  A268 );
 a35021a <=( a35020a  and  a35017a );
 a35022a <=( a35021a  and  a35014a );
 a35026a <=( (not A167)  and  A168 );
 a35027a <=( A170  and  a35026a );
 a35030a <=( (not A199)  and  A166 );
 a35033a <=( (not A202)  and  (not A200) );
 a35034a <=( a35033a  and  a35030a );
 a35035a <=( a35034a  and  a35027a );
 a35038a <=( (not A233)  and  A232 );
 a35041a <=( A236  and  (not A235) );
 a35042a <=( a35041a  and  a35038a );
 a35045a <=( A266  and  (not A265) );
 a35048a <=( A269  and  (not A268) );
 a35049a <=( a35048a  and  a35045a );
 a35050a <=( a35049a  and  a35042a );
 a35054a <=( (not A167)  and  A168 );
 a35055a <=( A170  and  a35054a );
 a35058a <=( (not A199)  and  A166 );
 a35061a <=( (not A202)  and  (not A200) );
 a35062a <=( a35061a  and  a35058a );
 a35063a <=( a35062a  and  a35055a );
 a35066a <=( (not A233)  and  A232 );
 a35069a <=( A236  and  (not A235) );
 a35070a <=( a35069a  and  a35066a );
 a35073a <=( (not A266)  and  A265 );
 a35076a <=( A269  and  (not A268) );
 a35077a <=( a35076a  and  a35073a );
 a35078a <=( a35077a  and  a35070a );
 a35082a <=( (not A167)  and  A168 );
 a35083a <=( A170  and  a35082a );
 a35086a <=( (not A199)  and  A166 );
 a35089a <=( (not A202)  and  (not A200) );
 a35090a <=( a35089a  and  a35086a );
 a35091a <=( a35090a  and  a35083a );
 a35094a <=( (not A233)  and  A232 );
 a35097a <=( A236  and  (not A235) );
 a35098a <=( a35097a  and  a35094a );
 a35101a <=( (not A266)  and  (not A265) );
 a35104a <=( (not A269)  and  A268 );
 a35105a <=( a35104a  and  a35101a );
 a35106a <=( a35105a  and  a35098a );
 a35110a <=( (not A167)  and  A168 );
 a35111a <=( A170  and  a35110a );
 a35114a <=( (not A199)  and  A166 );
 a35117a <=( (not A202)  and  (not A200) );
 a35118a <=( a35117a  and  a35114a );
 a35119a <=( a35118a  and  a35111a );
 a35122a <=( (not A233)  and  (not A232) );
 a35125a <=( (not A236)  and  A235 );
 a35126a <=( a35125a  and  a35122a );
 a35129a <=( A299  and  A298 );
 a35132a <=( (not A302)  and  A301 );
 a35133a <=( a35132a  and  a35129a );
 a35134a <=( a35133a  and  a35126a );
 a35138a <=( (not A167)  and  A168 );
 a35139a <=( A170  and  a35138a );
 a35142a <=( (not A199)  and  A166 );
 a35145a <=( (not A202)  and  (not A200) );
 a35146a <=( a35145a  and  a35142a );
 a35147a <=( a35146a  and  a35139a );
 a35150a <=( (not A233)  and  (not A232) );
 a35153a <=( (not A236)  and  A235 );
 a35154a <=( a35153a  and  a35150a );
 a35157a <=( (not A299)  and  A298 );
 a35160a <=( A302  and  (not A301) );
 a35161a <=( a35160a  and  a35157a );
 a35162a <=( a35161a  and  a35154a );
 a35166a <=( (not A167)  and  A168 );
 a35167a <=( A170  and  a35166a );
 a35170a <=( (not A199)  and  A166 );
 a35173a <=( (not A202)  and  (not A200) );
 a35174a <=( a35173a  and  a35170a );
 a35175a <=( a35174a  and  a35167a );
 a35178a <=( (not A233)  and  (not A232) );
 a35181a <=( (not A236)  and  A235 );
 a35182a <=( a35181a  and  a35178a );
 a35185a <=( A299  and  (not A298) );
 a35188a <=( A302  and  (not A301) );
 a35189a <=( a35188a  and  a35185a );
 a35190a <=( a35189a  and  a35182a );
 a35194a <=( (not A167)  and  A168 );
 a35195a <=( A170  and  a35194a );
 a35198a <=( (not A199)  and  A166 );
 a35201a <=( (not A202)  and  (not A200) );
 a35202a <=( a35201a  and  a35198a );
 a35203a <=( a35202a  and  a35195a );
 a35206a <=( (not A233)  and  (not A232) );
 a35209a <=( (not A236)  and  A235 );
 a35210a <=( a35209a  and  a35206a );
 a35213a <=( (not A299)  and  (not A298) );
 a35216a <=( (not A302)  and  A301 );
 a35217a <=( a35216a  and  a35213a );
 a35218a <=( a35217a  and  a35210a );
 a35222a <=( (not A167)  and  A168 );
 a35223a <=( A170  and  a35222a );
 a35226a <=( (not A199)  and  A166 );
 a35229a <=( (not A202)  and  (not A200) );
 a35230a <=( a35229a  and  a35226a );
 a35231a <=( a35230a  and  a35223a );
 a35234a <=( (not A233)  and  (not A232) );
 a35237a <=( (not A236)  and  A235 );
 a35238a <=( a35237a  and  a35234a );
 a35241a <=( A266  and  A265 );
 a35244a <=( (not A269)  and  A268 );
 a35245a <=( a35244a  and  a35241a );
 a35246a <=( a35245a  and  a35238a );
 a35250a <=( (not A167)  and  A168 );
 a35251a <=( A170  and  a35250a );
 a35254a <=( (not A199)  and  A166 );
 a35257a <=( (not A202)  and  (not A200) );
 a35258a <=( a35257a  and  a35254a );
 a35259a <=( a35258a  and  a35251a );
 a35262a <=( (not A233)  and  (not A232) );
 a35265a <=( (not A236)  and  A235 );
 a35266a <=( a35265a  and  a35262a );
 a35269a <=( A266  and  (not A265) );
 a35272a <=( A269  and  (not A268) );
 a35273a <=( a35272a  and  a35269a );
 a35274a <=( a35273a  and  a35266a );
 a35278a <=( (not A167)  and  A168 );
 a35279a <=( A170  and  a35278a );
 a35282a <=( (not A199)  and  A166 );
 a35285a <=( (not A202)  and  (not A200) );
 a35286a <=( a35285a  and  a35282a );
 a35287a <=( a35286a  and  a35279a );
 a35290a <=( (not A233)  and  (not A232) );
 a35293a <=( (not A236)  and  A235 );
 a35294a <=( a35293a  and  a35290a );
 a35297a <=( (not A266)  and  A265 );
 a35300a <=( A269  and  (not A268) );
 a35301a <=( a35300a  and  a35297a );
 a35302a <=( a35301a  and  a35294a );
 a35306a <=( (not A167)  and  A168 );
 a35307a <=( A170  and  a35306a );
 a35310a <=( (not A199)  and  A166 );
 a35313a <=( (not A202)  and  (not A200) );
 a35314a <=( a35313a  and  a35310a );
 a35315a <=( a35314a  and  a35307a );
 a35318a <=( (not A233)  and  (not A232) );
 a35321a <=( (not A236)  and  A235 );
 a35322a <=( a35321a  and  a35318a );
 a35325a <=( (not A266)  and  (not A265) );
 a35328a <=( (not A269)  and  A268 );
 a35329a <=( a35328a  and  a35325a );
 a35330a <=( a35329a  and  a35322a );
 a35334a <=( (not A167)  and  A168 );
 a35335a <=( A170  and  a35334a );
 a35338a <=( (not A199)  and  A166 );
 a35341a <=( A203  and  (not A200) );
 a35342a <=( a35341a  and  a35338a );
 a35343a <=( a35342a  and  a35335a );
 a35346a <=( A233  and  A232 );
 a35349a <=( (not A236)  and  A235 );
 a35350a <=( a35349a  and  a35346a );
 a35353a <=( A299  and  A298 );
 a35356a <=( (not A302)  and  A301 );
 a35357a <=( a35356a  and  a35353a );
 a35358a <=( a35357a  and  a35350a );
 a35362a <=( (not A167)  and  A168 );
 a35363a <=( A170  and  a35362a );
 a35366a <=( (not A199)  and  A166 );
 a35369a <=( A203  and  (not A200) );
 a35370a <=( a35369a  and  a35366a );
 a35371a <=( a35370a  and  a35363a );
 a35374a <=( A233  and  A232 );
 a35377a <=( (not A236)  and  A235 );
 a35378a <=( a35377a  and  a35374a );
 a35381a <=( (not A299)  and  A298 );
 a35384a <=( A302  and  (not A301) );
 a35385a <=( a35384a  and  a35381a );
 a35386a <=( a35385a  and  a35378a );
 a35390a <=( (not A167)  and  A168 );
 a35391a <=( A170  and  a35390a );
 a35394a <=( (not A199)  and  A166 );
 a35397a <=( A203  and  (not A200) );
 a35398a <=( a35397a  and  a35394a );
 a35399a <=( a35398a  and  a35391a );
 a35402a <=( A233  and  A232 );
 a35405a <=( (not A236)  and  A235 );
 a35406a <=( a35405a  and  a35402a );
 a35409a <=( A299  and  (not A298) );
 a35412a <=( A302  and  (not A301) );
 a35413a <=( a35412a  and  a35409a );
 a35414a <=( a35413a  and  a35406a );
 a35418a <=( (not A167)  and  A168 );
 a35419a <=( A170  and  a35418a );
 a35422a <=( (not A199)  and  A166 );
 a35425a <=( A203  and  (not A200) );
 a35426a <=( a35425a  and  a35422a );
 a35427a <=( a35426a  and  a35419a );
 a35430a <=( A233  and  A232 );
 a35433a <=( (not A236)  and  A235 );
 a35434a <=( a35433a  and  a35430a );
 a35437a <=( (not A299)  and  (not A298) );
 a35440a <=( (not A302)  and  A301 );
 a35441a <=( a35440a  and  a35437a );
 a35442a <=( a35441a  and  a35434a );
 a35446a <=( (not A167)  and  A168 );
 a35447a <=( A170  and  a35446a );
 a35450a <=( (not A199)  and  A166 );
 a35453a <=( A203  and  (not A200) );
 a35454a <=( a35453a  and  a35450a );
 a35455a <=( a35454a  and  a35447a );
 a35458a <=( A233  and  A232 );
 a35461a <=( (not A236)  and  A235 );
 a35462a <=( a35461a  and  a35458a );
 a35465a <=( A266  and  A265 );
 a35468a <=( (not A269)  and  A268 );
 a35469a <=( a35468a  and  a35465a );
 a35470a <=( a35469a  and  a35462a );
 a35474a <=( (not A167)  and  A168 );
 a35475a <=( A170  and  a35474a );
 a35478a <=( (not A199)  and  A166 );
 a35481a <=( A203  and  (not A200) );
 a35482a <=( a35481a  and  a35478a );
 a35483a <=( a35482a  and  a35475a );
 a35486a <=( A233  and  A232 );
 a35489a <=( (not A236)  and  A235 );
 a35490a <=( a35489a  and  a35486a );
 a35493a <=( A266  and  (not A265) );
 a35496a <=( A269  and  (not A268) );
 a35497a <=( a35496a  and  a35493a );
 a35498a <=( a35497a  and  a35490a );
 a35502a <=( (not A167)  and  A168 );
 a35503a <=( A170  and  a35502a );
 a35506a <=( (not A199)  and  A166 );
 a35509a <=( A203  and  (not A200) );
 a35510a <=( a35509a  and  a35506a );
 a35511a <=( a35510a  and  a35503a );
 a35514a <=( A233  and  A232 );
 a35517a <=( (not A236)  and  A235 );
 a35518a <=( a35517a  and  a35514a );
 a35521a <=( (not A266)  and  A265 );
 a35524a <=( A269  and  (not A268) );
 a35525a <=( a35524a  and  a35521a );
 a35526a <=( a35525a  and  a35518a );
 a35530a <=( (not A167)  and  A168 );
 a35531a <=( A170  and  a35530a );
 a35534a <=( (not A199)  and  A166 );
 a35537a <=( A203  and  (not A200) );
 a35538a <=( a35537a  and  a35534a );
 a35539a <=( a35538a  and  a35531a );
 a35542a <=( A233  and  A232 );
 a35545a <=( (not A236)  and  A235 );
 a35546a <=( a35545a  and  a35542a );
 a35549a <=( (not A266)  and  (not A265) );
 a35552a <=( (not A269)  and  A268 );
 a35553a <=( a35552a  and  a35549a );
 a35554a <=( a35553a  and  a35546a );
 a35558a <=( (not A167)  and  A168 );
 a35559a <=( A170  and  a35558a );
 a35562a <=( (not A199)  and  A166 );
 a35565a <=( A203  and  (not A200) );
 a35566a <=( a35565a  and  a35562a );
 a35567a <=( a35566a  and  a35559a );
 a35570a <=( A233  and  (not A232) );
 a35573a <=( A236  and  (not A235) );
 a35574a <=( a35573a  and  a35570a );
 a35577a <=( A299  and  A298 );
 a35580a <=( (not A302)  and  A301 );
 a35581a <=( a35580a  and  a35577a );
 a35582a <=( a35581a  and  a35574a );
 a35586a <=( (not A167)  and  A168 );
 a35587a <=( A170  and  a35586a );
 a35590a <=( (not A199)  and  A166 );
 a35593a <=( A203  and  (not A200) );
 a35594a <=( a35593a  and  a35590a );
 a35595a <=( a35594a  and  a35587a );
 a35598a <=( A233  and  (not A232) );
 a35601a <=( A236  and  (not A235) );
 a35602a <=( a35601a  and  a35598a );
 a35605a <=( (not A299)  and  A298 );
 a35608a <=( A302  and  (not A301) );
 a35609a <=( a35608a  and  a35605a );
 a35610a <=( a35609a  and  a35602a );
 a35614a <=( (not A167)  and  A168 );
 a35615a <=( A170  and  a35614a );
 a35618a <=( (not A199)  and  A166 );
 a35621a <=( A203  and  (not A200) );
 a35622a <=( a35621a  and  a35618a );
 a35623a <=( a35622a  and  a35615a );
 a35626a <=( A233  and  (not A232) );
 a35629a <=( A236  and  (not A235) );
 a35630a <=( a35629a  and  a35626a );
 a35633a <=( A299  and  (not A298) );
 a35636a <=( A302  and  (not A301) );
 a35637a <=( a35636a  and  a35633a );
 a35638a <=( a35637a  and  a35630a );
 a35642a <=( (not A167)  and  A168 );
 a35643a <=( A170  and  a35642a );
 a35646a <=( (not A199)  and  A166 );
 a35649a <=( A203  and  (not A200) );
 a35650a <=( a35649a  and  a35646a );
 a35651a <=( a35650a  and  a35643a );
 a35654a <=( A233  and  (not A232) );
 a35657a <=( A236  and  (not A235) );
 a35658a <=( a35657a  and  a35654a );
 a35661a <=( (not A299)  and  (not A298) );
 a35664a <=( (not A302)  and  A301 );
 a35665a <=( a35664a  and  a35661a );
 a35666a <=( a35665a  and  a35658a );
 a35670a <=( (not A167)  and  A168 );
 a35671a <=( A170  and  a35670a );
 a35674a <=( (not A199)  and  A166 );
 a35677a <=( A203  and  (not A200) );
 a35678a <=( a35677a  and  a35674a );
 a35679a <=( a35678a  and  a35671a );
 a35682a <=( A233  and  (not A232) );
 a35685a <=( A236  and  (not A235) );
 a35686a <=( a35685a  and  a35682a );
 a35689a <=( A266  and  A265 );
 a35692a <=( (not A269)  and  A268 );
 a35693a <=( a35692a  and  a35689a );
 a35694a <=( a35693a  and  a35686a );
 a35698a <=( (not A167)  and  A168 );
 a35699a <=( A170  and  a35698a );
 a35702a <=( (not A199)  and  A166 );
 a35705a <=( A203  and  (not A200) );
 a35706a <=( a35705a  and  a35702a );
 a35707a <=( a35706a  and  a35699a );
 a35710a <=( A233  and  (not A232) );
 a35713a <=( A236  and  (not A235) );
 a35714a <=( a35713a  and  a35710a );
 a35717a <=( A266  and  (not A265) );
 a35720a <=( A269  and  (not A268) );
 a35721a <=( a35720a  and  a35717a );
 a35722a <=( a35721a  and  a35714a );
 a35726a <=( (not A167)  and  A168 );
 a35727a <=( A170  and  a35726a );
 a35730a <=( (not A199)  and  A166 );
 a35733a <=( A203  and  (not A200) );
 a35734a <=( a35733a  and  a35730a );
 a35735a <=( a35734a  and  a35727a );
 a35738a <=( A233  and  (not A232) );
 a35741a <=( A236  and  (not A235) );
 a35742a <=( a35741a  and  a35738a );
 a35745a <=( (not A266)  and  A265 );
 a35748a <=( A269  and  (not A268) );
 a35749a <=( a35748a  and  a35745a );
 a35750a <=( a35749a  and  a35742a );
 a35754a <=( (not A167)  and  A168 );
 a35755a <=( A170  and  a35754a );
 a35758a <=( (not A199)  and  A166 );
 a35761a <=( A203  and  (not A200) );
 a35762a <=( a35761a  and  a35758a );
 a35763a <=( a35762a  and  a35755a );
 a35766a <=( A233  and  (not A232) );
 a35769a <=( A236  and  (not A235) );
 a35770a <=( a35769a  and  a35766a );
 a35773a <=( (not A266)  and  (not A265) );
 a35776a <=( (not A269)  and  A268 );
 a35777a <=( a35776a  and  a35773a );
 a35778a <=( a35777a  and  a35770a );
 a35782a <=( (not A167)  and  A168 );
 a35783a <=( A170  and  a35782a );
 a35786a <=( (not A199)  and  A166 );
 a35789a <=( A203  and  (not A200) );
 a35790a <=( a35789a  and  a35786a );
 a35791a <=( a35790a  and  a35783a );
 a35794a <=( (not A233)  and  A232 );
 a35797a <=( A236  and  (not A235) );
 a35798a <=( a35797a  and  a35794a );
 a35801a <=( A299  and  A298 );
 a35804a <=( (not A302)  and  A301 );
 a35805a <=( a35804a  and  a35801a );
 a35806a <=( a35805a  and  a35798a );
 a35810a <=( (not A167)  and  A168 );
 a35811a <=( A170  and  a35810a );
 a35814a <=( (not A199)  and  A166 );
 a35817a <=( A203  and  (not A200) );
 a35818a <=( a35817a  and  a35814a );
 a35819a <=( a35818a  and  a35811a );
 a35822a <=( (not A233)  and  A232 );
 a35825a <=( A236  and  (not A235) );
 a35826a <=( a35825a  and  a35822a );
 a35829a <=( (not A299)  and  A298 );
 a35832a <=( A302  and  (not A301) );
 a35833a <=( a35832a  and  a35829a );
 a35834a <=( a35833a  and  a35826a );
 a35838a <=( (not A167)  and  A168 );
 a35839a <=( A170  and  a35838a );
 a35842a <=( (not A199)  and  A166 );
 a35845a <=( A203  and  (not A200) );
 a35846a <=( a35845a  and  a35842a );
 a35847a <=( a35846a  and  a35839a );
 a35850a <=( (not A233)  and  A232 );
 a35853a <=( A236  and  (not A235) );
 a35854a <=( a35853a  and  a35850a );
 a35857a <=( A299  and  (not A298) );
 a35860a <=( A302  and  (not A301) );
 a35861a <=( a35860a  and  a35857a );
 a35862a <=( a35861a  and  a35854a );
 a35866a <=( (not A167)  and  A168 );
 a35867a <=( A170  and  a35866a );
 a35870a <=( (not A199)  and  A166 );
 a35873a <=( A203  and  (not A200) );
 a35874a <=( a35873a  and  a35870a );
 a35875a <=( a35874a  and  a35867a );
 a35878a <=( (not A233)  and  A232 );
 a35881a <=( A236  and  (not A235) );
 a35882a <=( a35881a  and  a35878a );
 a35885a <=( (not A299)  and  (not A298) );
 a35888a <=( (not A302)  and  A301 );
 a35889a <=( a35888a  and  a35885a );
 a35890a <=( a35889a  and  a35882a );
 a35894a <=( (not A167)  and  A168 );
 a35895a <=( A170  and  a35894a );
 a35898a <=( (not A199)  and  A166 );
 a35901a <=( A203  and  (not A200) );
 a35902a <=( a35901a  and  a35898a );
 a35903a <=( a35902a  and  a35895a );
 a35906a <=( (not A233)  and  A232 );
 a35909a <=( A236  and  (not A235) );
 a35910a <=( a35909a  and  a35906a );
 a35913a <=( A266  and  A265 );
 a35916a <=( (not A269)  and  A268 );
 a35917a <=( a35916a  and  a35913a );
 a35918a <=( a35917a  and  a35910a );
 a35922a <=( (not A167)  and  A168 );
 a35923a <=( A170  and  a35922a );
 a35926a <=( (not A199)  and  A166 );
 a35929a <=( A203  and  (not A200) );
 a35930a <=( a35929a  and  a35926a );
 a35931a <=( a35930a  and  a35923a );
 a35934a <=( (not A233)  and  A232 );
 a35937a <=( A236  and  (not A235) );
 a35938a <=( a35937a  and  a35934a );
 a35941a <=( A266  and  (not A265) );
 a35944a <=( A269  and  (not A268) );
 a35945a <=( a35944a  and  a35941a );
 a35946a <=( a35945a  and  a35938a );
 a35950a <=( (not A167)  and  A168 );
 a35951a <=( A170  and  a35950a );
 a35954a <=( (not A199)  and  A166 );
 a35957a <=( A203  and  (not A200) );
 a35958a <=( a35957a  and  a35954a );
 a35959a <=( a35958a  and  a35951a );
 a35962a <=( (not A233)  and  A232 );
 a35965a <=( A236  and  (not A235) );
 a35966a <=( a35965a  and  a35962a );
 a35969a <=( (not A266)  and  A265 );
 a35972a <=( A269  and  (not A268) );
 a35973a <=( a35972a  and  a35969a );
 a35974a <=( a35973a  and  a35966a );
 a35978a <=( (not A167)  and  A168 );
 a35979a <=( A170  and  a35978a );
 a35982a <=( (not A199)  and  A166 );
 a35985a <=( A203  and  (not A200) );
 a35986a <=( a35985a  and  a35982a );
 a35987a <=( a35986a  and  a35979a );
 a35990a <=( (not A233)  and  A232 );
 a35993a <=( A236  and  (not A235) );
 a35994a <=( a35993a  and  a35990a );
 a35997a <=( (not A266)  and  (not A265) );
 a36000a <=( (not A269)  and  A268 );
 a36001a <=( a36000a  and  a35997a );
 a36002a <=( a36001a  and  a35994a );
 a36006a <=( (not A167)  and  A168 );
 a36007a <=( A170  and  a36006a );
 a36010a <=( (not A199)  and  A166 );
 a36013a <=( A203  and  (not A200) );
 a36014a <=( a36013a  and  a36010a );
 a36015a <=( a36014a  and  a36007a );
 a36018a <=( (not A233)  and  (not A232) );
 a36021a <=( (not A236)  and  A235 );
 a36022a <=( a36021a  and  a36018a );
 a36025a <=( A299  and  A298 );
 a36028a <=( (not A302)  and  A301 );
 a36029a <=( a36028a  and  a36025a );
 a36030a <=( a36029a  and  a36022a );
 a36034a <=( (not A167)  and  A168 );
 a36035a <=( A170  and  a36034a );
 a36038a <=( (not A199)  and  A166 );
 a36041a <=( A203  and  (not A200) );
 a36042a <=( a36041a  and  a36038a );
 a36043a <=( a36042a  and  a36035a );
 a36046a <=( (not A233)  and  (not A232) );
 a36049a <=( (not A236)  and  A235 );
 a36050a <=( a36049a  and  a36046a );
 a36053a <=( (not A299)  and  A298 );
 a36056a <=( A302  and  (not A301) );
 a36057a <=( a36056a  and  a36053a );
 a36058a <=( a36057a  and  a36050a );
 a36062a <=( (not A167)  and  A168 );
 a36063a <=( A170  and  a36062a );
 a36066a <=( (not A199)  and  A166 );
 a36069a <=( A203  and  (not A200) );
 a36070a <=( a36069a  and  a36066a );
 a36071a <=( a36070a  and  a36063a );
 a36074a <=( (not A233)  and  (not A232) );
 a36077a <=( (not A236)  and  A235 );
 a36078a <=( a36077a  and  a36074a );
 a36081a <=( A299  and  (not A298) );
 a36084a <=( A302  and  (not A301) );
 a36085a <=( a36084a  and  a36081a );
 a36086a <=( a36085a  and  a36078a );
 a36090a <=( (not A167)  and  A168 );
 a36091a <=( A170  and  a36090a );
 a36094a <=( (not A199)  and  A166 );
 a36097a <=( A203  and  (not A200) );
 a36098a <=( a36097a  and  a36094a );
 a36099a <=( a36098a  and  a36091a );
 a36102a <=( (not A233)  and  (not A232) );
 a36105a <=( (not A236)  and  A235 );
 a36106a <=( a36105a  and  a36102a );
 a36109a <=( (not A299)  and  (not A298) );
 a36112a <=( (not A302)  and  A301 );
 a36113a <=( a36112a  and  a36109a );
 a36114a <=( a36113a  and  a36106a );
 a36118a <=( (not A167)  and  A168 );
 a36119a <=( A170  and  a36118a );
 a36122a <=( (not A199)  and  A166 );
 a36125a <=( A203  and  (not A200) );
 a36126a <=( a36125a  and  a36122a );
 a36127a <=( a36126a  and  a36119a );
 a36130a <=( (not A233)  and  (not A232) );
 a36133a <=( (not A236)  and  A235 );
 a36134a <=( a36133a  and  a36130a );
 a36137a <=( A266  and  A265 );
 a36140a <=( (not A269)  and  A268 );
 a36141a <=( a36140a  and  a36137a );
 a36142a <=( a36141a  and  a36134a );
 a36146a <=( (not A167)  and  A168 );
 a36147a <=( A170  and  a36146a );
 a36150a <=( (not A199)  and  A166 );
 a36153a <=( A203  and  (not A200) );
 a36154a <=( a36153a  and  a36150a );
 a36155a <=( a36154a  and  a36147a );
 a36158a <=( (not A233)  and  (not A232) );
 a36161a <=( (not A236)  and  A235 );
 a36162a <=( a36161a  and  a36158a );
 a36165a <=( A266  and  (not A265) );
 a36168a <=( A269  and  (not A268) );
 a36169a <=( a36168a  and  a36165a );
 a36170a <=( a36169a  and  a36162a );
 a36174a <=( (not A167)  and  A168 );
 a36175a <=( A170  and  a36174a );
 a36178a <=( (not A199)  and  A166 );
 a36181a <=( A203  and  (not A200) );
 a36182a <=( a36181a  and  a36178a );
 a36183a <=( a36182a  and  a36175a );
 a36186a <=( (not A233)  and  (not A232) );
 a36189a <=( (not A236)  and  A235 );
 a36190a <=( a36189a  and  a36186a );
 a36193a <=( (not A266)  and  A265 );
 a36196a <=( A269  and  (not A268) );
 a36197a <=( a36196a  and  a36193a );
 a36198a <=( a36197a  and  a36190a );
 a36202a <=( (not A167)  and  A168 );
 a36203a <=( A170  and  a36202a );
 a36206a <=( (not A199)  and  A166 );
 a36209a <=( A203  and  (not A200) );
 a36210a <=( a36209a  and  a36206a );
 a36211a <=( a36210a  and  a36203a );
 a36214a <=( (not A233)  and  (not A232) );
 a36217a <=( (not A236)  and  A235 );
 a36218a <=( a36217a  and  a36214a );
 a36221a <=( (not A266)  and  (not A265) );
 a36224a <=( (not A269)  and  A268 );
 a36225a <=( a36224a  and  a36221a );
 a36226a <=( a36225a  and  a36218a );
 a36230a <=( (not A167)  and  A168 );
 a36231a <=( A169  and  a36230a );
 a36234a <=( (not A199)  and  A166 );
 a36237a <=( (not A202)  and  (not A200) );
 a36238a <=( a36237a  and  a36234a );
 a36239a <=( a36238a  and  a36231a );
 a36242a <=( A233  and  A232 );
 a36245a <=( (not A236)  and  A235 );
 a36246a <=( a36245a  and  a36242a );
 a36249a <=( A299  and  A298 );
 a36252a <=( (not A302)  and  A301 );
 a36253a <=( a36252a  and  a36249a );
 a36254a <=( a36253a  and  a36246a );
 a36258a <=( (not A167)  and  A168 );
 a36259a <=( A169  and  a36258a );
 a36262a <=( (not A199)  and  A166 );
 a36265a <=( (not A202)  and  (not A200) );
 a36266a <=( a36265a  and  a36262a );
 a36267a <=( a36266a  and  a36259a );
 a36270a <=( A233  and  A232 );
 a36273a <=( (not A236)  and  A235 );
 a36274a <=( a36273a  and  a36270a );
 a36277a <=( (not A299)  and  A298 );
 a36280a <=( A302  and  (not A301) );
 a36281a <=( a36280a  and  a36277a );
 a36282a <=( a36281a  and  a36274a );
 a36286a <=( (not A167)  and  A168 );
 a36287a <=( A169  and  a36286a );
 a36290a <=( (not A199)  and  A166 );
 a36293a <=( (not A202)  and  (not A200) );
 a36294a <=( a36293a  and  a36290a );
 a36295a <=( a36294a  and  a36287a );
 a36298a <=( A233  and  A232 );
 a36301a <=( (not A236)  and  A235 );
 a36302a <=( a36301a  and  a36298a );
 a36305a <=( A299  and  (not A298) );
 a36308a <=( A302  and  (not A301) );
 a36309a <=( a36308a  and  a36305a );
 a36310a <=( a36309a  and  a36302a );
 a36314a <=( (not A167)  and  A168 );
 a36315a <=( A169  and  a36314a );
 a36318a <=( (not A199)  and  A166 );
 a36321a <=( (not A202)  and  (not A200) );
 a36322a <=( a36321a  and  a36318a );
 a36323a <=( a36322a  and  a36315a );
 a36326a <=( A233  and  A232 );
 a36329a <=( (not A236)  and  A235 );
 a36330a <=( a36329a  and  a36326a );
 a36333a <=( (not A299)  and  (not A298) );
 a36336a <=( (not A302)  and  A301 );
 a36337a <=( a36336a  and  a36333a );
 a36338a <=( a36337a  and  a36330a );
 a36342a <=( (not A167)  and  A168 );
 a36343a <=( A169  and  a36342a );
 a36346a <=( (not A199)  and  A166 );
 a36349a <=( (not A202)  and  (not A200) );
 a36350a <=( a36349a  and  a36346a );
 a36351a <=( a36350a  and  a36343a );
 a36354a <=( A233  and  A232 );
 a36357a <=( (not A236)  and  A235 );
 a36358a <=( a36357a  and  a36354a );
 a36361a <=( A266  and  A265 );
 a36364a <=( (not A269)  and  A268 );
 a36365a <=( a36364a  and  a36361a );
 a36366a <=( a36365a  and  a36358a );
 a36370a <=( (not A167)  and  A168 );
 a36371a <=( A169  and  a36370a );
 a36374a <=( (not A199)  and  A166 );
 a36377a <=( (not A202)  and  (not A200) );
 a36378a <=( a36377a  and  a36374a );
 a36379a <=( a36378a  and  a36371a );
 a36382a <=( A233  and  A232 );
 a36385a <=( (not A236)  and  A235 );
 a36386a <=( a36385a  and  a36382a );
 a36389a <=( A266  and  (not A265) );
 a36392a <=( A269  and  (not A268) );
 a36393a <=( a36392a  and  a36389a );
 a36394a <=( a36393a  and  a36386a );
 a36398a <=( (not A167)  and  A168 );
 a36399a <=( A169  and  a36398a );
 a36402a <=( (not A199)  and  A166 );
 a36405a <=( (not A202)  and  (not A200) );
 a36406a <=( a36405a  and  a36402a );
 a36407a <=( a36406a  and  a36399a );
 a36410a <=( A233  and  A232 );
 a36413a <=( (not A236)  and  A235 );
 a36414a <=( a36413a  and  a36410a );
 a36417a <=( (not A266)  and  A265 );
 a36420a <=( A269  and  (not A268) );
 a36421a <=( a36420a  and  a36417a );
 a36422a <=( a36421a  and  a36414a );
 a36426a <=( (not A167)  and  A168 );
 a36427a <=( A169  and  a36426a );
 a36430a <=( (not A199)  and  A166 );
 a36433a <=( (not A202)  and  (not A200) );
 a36434a <=( a36433a  and  a36430a );
 a36435a <=( a36434a  and  a36427a );
 a36438a <=( A233  and  A232 );
 a36441a <=( (not A236)  and  A235 );
 a36442a <=( a36441a  and  a36438a );
 a36445a <=( (not A266)  and  (not A265) );
 a36448a <=( (not A269)  and  A268 );
 a36449a <=( a36448a  and  a36445a );
 a36450a <=( a36449a  and  a36442a );
 a36454a <=( (not A167)  and  A168 );
 a36455a <=( A169  and  a36454a );
 a36458a <=( (not A199)  and  A166 );
 a36461a <=( (not A202)  and  (not A200) );
 a36462a <=( a36461a  and  a36458a );
 a36463a <=( a36462a  and  a36455a );
 a36466a <=( A233  and  (not A232) );
 a36469a <=( A236  and  (not A235) );
 a36470a <=( a36469a  and  a36466a );
 a36473a <=( A299  and  A298 );
 a36476a <=( (not A302)  and  A301 );
 a36477a <=( a36476a  and  a36473a );
 a36478a <=( a36477a  and  a36470a );
 a36482a <=( (not A167)  and  A168 );
 a36483a <=( A169  and  a36482a );
 a36486a <=( (not A199)  and  A166 );
 a36489a <=( (not A202)  and  (not A200) );
 a36490a <=( a36489a  and  a36486a );
 a36491a <=( a36490a  and  a36483a );
 a36494a <=( A233  and  (not A232) );
 a36497a <=( A236  and  (not A235) );
 a36498a <=( a36497a  and  a36494a );
 a36501a <=( (not A299)  and  A298 );
 a36504a <=( A302  and  (not A301) );
 a36505a <=( a36504a  and  a36501a );
 a36506a <=( a36505a  and  a36498a );
 a36510a <=( (not A167)  and  A168 );
 a36511a <=( A169  and  a36510a );
 a36514a <=( (not A199)  and  A166 );
 a36517a <=( (not A202)  and  (not A200) );
 a36518a <=( a36517a  and  a36514a );
 a36519a <=( a36518a  and  a36511a );
 a36522a <=( A233  and  (not A232) );
 a36525a <=( A236  and  (not A235) );
 a36526a <=( a36525a  and  a36522a );
 a36529a <=( A299  and  (not A298) );
 a36532a <=( A302  and  (not A301) );
 a36533a <=( a36532a  and  a36529a );
 a36534a <=( a36533a  and  a36526a );
 a36538a <=( (not A167)  and  A168 );
 a36539a <=( A169  and  a36538a );
 a36542a <=( (not A199)  and  A166 );
 a36545a <=( (not A202)  and  (not A200) );
 a36546a <=( a36545a  and  a36542a );
 a36547a <=( a36546a  and  a36539a );
 a36550a <=( A233  and  (not A232) );
 a36553a <=( A236  and  (not A235) );
 a36554a <=( a36553a  and  a36550a );
 a36557a <=( (not A299)  and  (not A298) );
 a36560a <=( (not A302)  and  A301 );
 a36561a <=( a36560a  and  a36557a );
 a36562a <=( a36561a  and  a36554a );
 a36566a <=( (not A167)  and  A168 );
 a36567a <=( A169  and  a36566a );
 a36570a <=( (not A199)  and  A166 );
 a36573a <=( (not A202)  and  (not A200) );
 a36574a <=( a36573a  and  a36570a );
 a36575a <=( a36574a  and  a36567a );
 a36578a <=( A233  and  (not A232) );
 a36581a <=( A236  and  (not A235) );
 a36582a <=( a36581a  and  a36578a );
 a36585a <=( A266  and  A265 );
 a36588a <=( (not A269)  and  A268 );
 a36589a <=( a36588a  and  a36585a );
 a36590a <=( a36589a  and  a36582a );
 a36594a <=( (not A167)  and  A168 );
 a36595a <=( A169  and  a36594a );
 a36598a <=( (not A199)  and  A166 );
 a36601a <=( (not A202)  and  (not A200) );
 a36602a <=( a36601a  and  a36598a );
 a36603a <=( a36602a  and  a36595a );
 a36606a <=( A233  and  (not A232) );
 a36609a <=( A236  and  (not A235) );
 a36610a <=( a36609a  and  a36606a );
 a36613a <=( A266  and  (not A265) );
 a36616a <=( A269  and  (not A268) );
 a36617a <=( a36616a  and  a36613a );
 a36618a <=( a36617a  and  a36610a );
 a36622a <=( (not A167)  and  A168 );
 a36623a <=( A169  and  a36622a );
 a36626a <=( (not A199)  and  A166 );
 a36629a <=( (not A202)  and  (not A200) );
 a36630a <=( a36629a  and  a36626a );
 a36631a <=( a36630a  and  a36623a );
 a36634a <=( A233  and  (not A232) );
 a36637a <=( A236  and  (not A235) );
 a36638a <=( a36637a  and  a36634a );
 a36641a <=( (not A266)  and  A265 );
 a36644a <=( A269  and  (not A268) );
 a36645a <=( a36644a  and  a36641a );
 a36646a <=( a36645a  and  a36638a );
 a36650a <=( (not A167)  and  A168 );
 a36651a <=( A169  and  a36650a );
 a36654a <=( (not A199)  and  A166 );
 a36657a <=( (not A202)  and  (not A200) );
 a36658a <=( a36657a  and  a36654a );
 a36659a <=( a36658a  and  a36651a );
 a36662a <=( A233  and  (not A232) );
 a36665a <=( A236  and  (not A235) );
 a36666a <=( a36665a  and  a36662a );
 a36669a <=( (not A266)  and  (not A265) );
 a36672a <=( (not A269)  and  A268 );
 a36673a <=( a36672a  and  a36669a );
 a36674a <=( a36673a  and  a36666a );
 a36678a <=( (not A167)  and  A168 );
 a36679a <=( A169  and  a36678a );
 a36682a <=( (not A199)  and  A166 );
 a36685a <=( (not A202)  and  (not A200) );
 a36686a <=( a36685a  and  a36682a );
 a36687a <=( a36686a  and  a36679a );
 a36690a <=( (not A233)  and  A232 );
 a36693a <=( A236  and  (not A235) );
 a36694a <=( a36693a  and  a36690a );
 a36697a <=( A299  and  A298 );
 a36700a <=( (not A302)  and  A301 );
 a36701a <=( a36700a  and  a36697a );
 a36702a <=( a36701a  and  a36694a );
 a36706a <=( (not A167)  and  A168 );
 a36707a <=( A169  and  a36706a );
 a36710a <=( (not A199)  and  A166 );
 a36713a <=( (not A202)  and  (not A200) );
 a36714a <=( a36713a  and  a36710a );
 a36715a <=( a36714a  and  a36707a );
 a36718a <=( (not A233)  and  A232 );
 a36721a <=( A236  and  (not A235) );
 a36722a <=( a36721a  and  a36718a );
 a36725a <=( (not A299)  and  A298 );
 a36728a <=( A302  and  (not A301) );
 a36729a <=( a36728a  and  a36725a );
 a36730a <=( a36729a  and  a36722a );
 a36734a <=( (not A167)  and  A168 );
 a36735a <=( A169  and  a36734a );
 a36738a <=( (not A199)  and  A166 );
 a36741a <=( (not A202)  and  (not A200) );
 a36742a <=( a36741a  and  a36738a );
 a36743a <=( a36742a  and  a36735a );
 a36746a <=( (not A233)  and  A232 );
 a36749a <=( A236  and  (not A235) );
 a36750a <=( a36749a  and  a36746a );
 a36753a <=( A299  and  (not A298) );
 a36756a <=( A302  and  (not A301) );
 a36757a <=( a36756a  and  a36753a );
 a36758a <=( a36757a  and  a36750a );
 a36762a <=( (not A167)  and  A168 );
 a36763a <=( A169  and  a36762a );
 a36766a <=( (not A199)  and  A166 );
 a36769a <=( (not A202)  and  (not A200) );
 a36770a <=( a36769a  and  a36766a );
 a36771a <=( a36770a  and  a36763a );
 a36774a <=( (not A233)  and  A232 );
 a36777a <=( A236  and  (not A235) );
 a36778a <=( a36777a  and  a36774a );
 a36781a <=( (not A299)  and  (not A298) );
 a36784a <=( (not A302)  and  A301 );
 a36785a <=( a36784a  and  a36781a );
 a36786a <=( a36785a  and  a36778a );
 a36790a <=( (not A167)  and  A168 );
 a36791a <=( A169  and  a36790a );
 a36794a <=( (not A199)  and  A166 );
 a36797a <=( (not A202)  and  (not A200) );
 a36798a <=( a36797a  and  a36794a );
 a36799a <=( a36798a  and  a36791a );
 a36802a <=( (not A233)  and  A232 );
 a36805a <=( A236  and  (not A235) );
 a36806a <=( a36805a  and  a36802a );
 a36809a <=( A266  and  A265 );
 a36812a <=( (not A269)  and  A268 );
 a36813a <=( a36812a  and  a36809a );
 a36814a <=( a36813a  and  a36806a );
 a36818a <=( (not A167)  and  A168 );
 a36819a <=( A169  and  a36818a );
 a36822a <=( (not A199)  and  A166 );
 a36825a <=( (not A202)  and  (not A200) );
 a36826a <=( a36825a  and  a36822a );
 a36827a <=( a36826a  and  a36819a );
 a36830a <=( (not A233)  and  A232 );
 a36833a <=( A236  and  (not A235) );
 a36834a <=( a36833a  and  a36830a );
 a36837a <=( A266  and  (not A265) );
 a36840a <=( A269  and  (not A268) );
 a36841a <=( a36840a  and  a36837a );
 a36842a <=( a36841a  and  a36834a );
 a36846a <=( (not A167)  and  A168 );
 a36847a <=( A169  and  a36846a );
 a36850a <=( (not A199)  and  A166 );
 a36853a <=( (not A202)  and  (not A200) );
 a36854a <=( a36853a  and  a36850a );
 a36855a <=( a36854a  and  a36847a );
 a36858a <=( (not A233)  and  A232 );
 a36861a <=( A236  and  (not A235) );
 a36862a <=( a36861a  and  a36858a );
 a36865a <=( (not A266)  and  A265 );
 a36868a <=( A269  and  (not A268) );
 a36869a <=( a36868a  and  a36865a );
 a36870a <=( a36869a  and  a36862a );
 a36874a <=( (not A167)  and  A168 );
 a36875a <=( A169  and  a36874a );
 a36878a <=( (not A199)  and  A166 );
 a36881a <=( (not A202)  and  (not A200) );
 a36882a <=( a36881a  and  a36878a );
 a36883a <=( a36882a  and  a36875a );
 a36886a <=( (not A233)  and  A232 );
 a36889a <=( A236  and  (not A235) );
 a36890a <=( a36889a  and  a36886a );
 a36893a <=( (not A266)  and  (not A265) );
 a36896a <=( (not A269)  and  A268 );
 a36897a <=( a36896a  and  a36893a );
 a36898a <=( a36897a  and  a36890a );
 a36902a <=( (not A167)  and  A168 );
 a36903a <=( A169  and  a36902a );
 a36906a <=( (not A199)  and  A166 );
 a36909a <=( (not A202)  and  (not A200) );
 a36910a <=( a36909a  and  a36906a );
 a36911a <=( a36910a  and  a36903a );
 a36914a <=( (not A233)  and  (not A232) );
 a36917a <=( (not A236)  and  A235 );
 a36918a <=( a36917a  and  a36914a );
 a36921a <=( A299  and  A298 );
 a36924a <=( (not A302)  and  A301 );
 a36925a <=( a36924a  and  a36921a );
 a36926a <=( a36925a  and  a36918a );
 a36930a <=( (not A167)  and  A168 );
 a36931a <=( A169  and  a36930a );
 a36934a <=( (not A199)  and  A166 );
 a36937a <=( (not A202)  and  (not A200) );
 a36938a <=( a36937a  and  a36934a );
 a36939a <=( a36938a  and  a36931a );
 a36942a <=( (not A233)  and  (not A232) );
 a36945a <=( (not A236)  and  A235 );
 a36946a <=( a36945a  and  a36942a );
 a36949a <=( (not A299)  and  A298 );
 a36952a <=( A302  and  (not A301) );
 a36953a <=( a36952a  and  a36949a );
 a36954a <=( a36953a  and  a36946a );
 a36958a <=( (not A167)  and  A168 );
 a36959a <=( A169  and  a36958a );
 a36962a <=( (not A199)  and  A166 );
 a36965a <=( (not A202)  and  (not A200) );
 a36966a <=( a36965a  and  a36962a );
 a36967a <=( a36966a  and  a36959a );
 a36970a <=( (not A233)  and  (not A232) );
 a36973a <=( (not A236)  and  A235 );
 a36974a <=( a36973a  and  a36970a );
 a36977a <=( A299  and  (not A298) );
 a36980a <=( A302  and  (not A301) );
 a36981a <=( a36980a  and  a36977a );
 a36982a <=( a36981a  and  a36974a );
 a36986a <=( (not A167)  and  A168 );
 a36987a <=( A169  and  a36986a );
 a36990a <=( (not A199)  and  A166 );
 a36993a <=( (not A202)  and  (not A200) );
 a36994a <=( a36993a  and  a36990a );
 a36995a <=( a36994a  and  a36987a );
 a36998a <=( (not A233)  and  (not A232) );
 a37001a <=( (not A236)  and  A235 );
 a37002a <=( a37001a  and  a36998a );
 a37005a <=( (not A299)  and  (not A298) );
 a37008a <=( (not A302)  and  A301 );
 a37009a <=( a37008a  and  a37005a );
 a37010a <=( a37009a  and  a37002a );
 a37014a <=( (not A167)  and  A168 );
 a37015a <=( A169  and  a37014a );
 a37018a <=( (not A199)  and  A166 );
 a37021a <=( (not A202)  and  (not A200) );
 a37022a <=( a37021a  and  a37018a );
 a37023a <=( a37022a  and  a37015a );
 a37026a <=( (not A233)  and  (not A232) );
 a37029a <=( (not A236)  and  A235 );
 a37030a <=( a37029a  and  a37026a );
 a37033a <=( A266  and  A265 );
 a37036a <=( (not A269)  and  A268 );
 a37037a <=( a37036a  and  a37033a );
 a37038a <=( a37037a  and  a37030a );
 a37042a <=( (not A167)  and  A168 );
 a37043a <=( A169  and  a37042a );
 a37046a <=( (not A199)  and  A166 );
 a37049a <=( (not A202)  and  (not A200) );
 a37050a <=( a37049a  and  a37046a );
 a37051a <=( a37050a  and  a37043a );
 a37054a <=( (not A233)  and  (not A232) );
 a37057a <=( (not A236)  and  A235 );
 a37058a <=( a37057a  and  a37054a );
 a37061a <=( A266  and  (not A265) );
 a37064a <=( A269  and  (not A268) );
 a37065a <=( a37064a  and  a37061a );
 a37066a <=( a37065a  and  a37058a );
 a37070a <=( (not A167)  and  A168 );
 a37071a <=( A169  and  a37070a );
 a37074a <=( (not A199)  and  A166 );
 a37077a <=( (not A202)  and  (not A200) );
 a37078a <=( a37077a  and  a37074a );
 a37079a <=( a37078a  and  a37071a );
 a37082a <=( (not A233)  and  (not A232) );
 a37085a <=( (not A236)  and  A235 );
 a37086a <=( a37085a  and  a37082a );
 a37089a <=( (not A266)  and  A265 );
 a37092a <=( A269  and  (not A268) );
 a37093a <=( a37092a  and  a37089a );
 a37094a <=( a37093a  and  a37086a );
 a37098a <=( (not A167)  and  A168 );
 a37099a <=( A169  and  a37098a );
 a37102a <=( (not A199)  and  A166 );
 a37105a <=( (not A202)  and  (not A200) );
 a37106a <=( a37105a  and  a37102a );
 a37107a <=( a37106a  and  a37099a );
 a37110a <=( (not A233)  and  (not A232) );
 a37113a <=( (not A236)  and  A235 );
 a37114a <=( a37113a  and  a37110a );
 a37117a <=( (not A266)  and  (not A265) );
 a37120a <=( (not A269)  and  A268 );
 a37121a <=( a37120a  and  a37117a );
 a37122a <=( a37121a  and  a37114a );
 a37126a <=( (not A167)  and  A168 );
 a37127a <=( A169  and  a37126a );
 a37130a <=( (not A199)  and  A166 );
 a37133a <=( A203  and  (not A200) );
 a37134a <=( a37133a  and  a37130a );
 a37135a <=( a37134a  and  a37127a );
 a37138a <=( A233  and  A232 );
 a37141a <=( (not A236)  and  A235 );
 a37142a <=( a37141a  and  a37138a );
 a37145a <=( A299  and  A298 );
 a37148a <=( (not A302)  and  A301 );
 a37149a <=( a37148a  and  a37145a );
 a37150a <=( a37149a  and  a37142a );
 a37154a <=( (not A167)  and  A168 );
 a37155a <=( A169  and  a37154a );
 a37158a <=( (not A199)  and  A166 );
 a37161a <=( A203  and  (not A200) );
 a37162a <=( a37161a  and  a37158a );
 a37163a <=( a37162a  and  a37155a );
 a37166a <=( A233  and  A232 );
 a37169a <=( (not A236)  and  A235 );
 a37170a <=( a37169a  and  a37166a );
 a37173a <=( (not A299)  and  A298 );
 a37176a <=( A302  and  (not A301) );
 a37177a <=( a37176a  and  a37173a );
 a37178a <=( a37177a  and  a37170a );
 a37182a <=( (not A167)  and  A168 );
 a37183a <=( A169  and  a37182a );
 a37186a <=( (not A199)  and  A166 );
 a37189a <=( A203  and  (not A200) );
 a37190a <=( a37189a  and  a37186a );
 a37191a <=( a37190a  and  a37183a );
 a37194a <=( A233  and  A232 );
 a37197a <=( (not A236)  and  A235 );
 a37198a <=( a37197a  and  a37194a );
 a37201a <=( A299  and  (not A298) );
 a37204a <=( A302  and  (not A301) );
 a37205a <=( a37204a  and  a37201a );
 a37206a <=( a37205a  and  a37198a );
 a37210a <=( (not A167)  and  A168 );
 a37211a <=( A169  and  a37210a );
 a37214a <=( (not A199)  and  A166 );
 a37217a <=( A203  and  (not A200) );
 a37218a <=( a37217a  and  a37214a );
 a37219a <=( a37218a  and  a37211a );
 a37222a <=( A233  and  A232 );
 a37225a <=( (not A236)  and  A235 );
 a37226a <=( a37225a  and  a37222a );
 a37229a <=( (not A299)  and  (not A298) );
 a37232a <=( (not A302)  and  A301 );
 a37233a <=( a37232a  and  a37229a );
 a37234a <=( a37233a  and  a37226a );
 a37238a <=( (not A167)  and  A168 );
 a37239a <=( A169  and  a37238a );
 a37242a <=( (not A199)  and  A166 );
 a37245a <=( A203  and  (not A200) );
 a37246a <=( a37245a  and  a37242a );
 a37247a <=( a37246a  and  a37239a );
 a37250a <=( A233  and  A232 );
 a37253a <=( (not A236)  and  A235 );
 a37254a <=( a37253a  and  a37250a );
 a37257a <=( A266  and  A265 );
 a37260a <=( (not A269)  and  A268 );
 a37261a <=( a37260a  and  a37257a );
 a37262a <=( a37261a  and  a37254a );
 a37266a <=( (not A167)  and  A168 );
 a37267a <=( A169  and  a37266a );
 a37270a <=( (not A199)  and  A166 );
 a37273a <=( A203  and  (not A200) );
 a37274a <=( a37273a  and  a37270a );
 a37275a <=( a37274a  and  a37267a );
 a37278a <=( A233  and  A232 );
 a37281a <=( (not A236)  and  A235 );
 a37282a <=( a37281a  and  a37278a );
 a37285a <=( A266  and  (not A265) );
 a37288a <=( A269  and  (not A268) );
 a37289a <=( a37288a  and  a37285a );
 a37290a <=( a37289a  and  a37282a );
 a37294a <=( (not A167)  and  A168 );
 a37295a <=( A169  and  a37294a );
 a37298a <=( (not A199)  and  A166 );
 a37301a <=( A203  and  (not A200) );
 a37302a <=( a37301a  and  a37298a );
 a37303a <=( a37302a  and  a37295a );
 a37306a <=( A233  and  A232 );
 a37309a <=( (not A236)  and  A235 );
 a37310a <=( a37309a  and  a37306a );
 a37313a <=( (not A266)  and  A265 );
 a37316a <=( A269  and  (not A268) );
 a37317a <=( a37316a  and  a37313a );
 a37318a <=( a37317a  and  a37310a );
 a37322a <=( (not A167)  and  A168 );
 a37323a <=( A169  and  a37322a );
 a37326a <=( (not A199)  and  A166 );
 a37329a <=( A203  and  (not A200) );
 a37330a <=( a37329a  and  a37326a );
 a37331a <=( a37330a  and  a37323a );
 a37334a <=( A233  and  A232 );
 a37337a <=( (not A236)  and  A235 );
 a37338a <=( a37337a  and  a37334a );
 a37341a <=( (not A266)  and  (not A265) );
 a37344a <=( (not A269)  and  A268 );
 a37345a <=( a37344a  and  a37341a );
 a37346a <=( a37345a  and  a37338a );
 a37350a <=( (not A167)  and  A168 );
 a37351a <=( A169  and  a37350a );
 a37354a <=( (not A199)  and  A166 );
 a37357a <=( A203  and  (not A200) );
 a37358a <=( a37357a  and  a37354a );
 a37359a <=( a37358a  and  a37351a );
 a37362a <=( A233  and  (not A232) );
 a37365a <=( A236  and  (not A235) );
 a37366a <=( a37365a  and  a37362a );
 a37369a <=( A299  and  A298 );
 a37372a <=( (not A302)  and  A301 );
 a37373a <=( a37372a  and  a37369a );
 a37374a <=( a37373a  and  a37366a );
 a37378a <=( (not A167)  and  A168 );
 a37379a <=( A169  and  a37378a );
 a37382a <=( (not A199)  and  A166 );
 a37385a <=( A203  and  (not A200) );
 a37386a <=( a37385a  and  a37382a );
 a37387a <=( a37386a  and  a37379a );
 a37390a <=( A233  and  (not A232) );
 a37393a <=( A236  and  (not A235) );
 a37394a <=( a37393a  and  a37390a );
 a37397a <=( (not A299)  and  A298 );
 a37400a <=( A302  and  (not A301) );
 a37401a <=( a37400a  and  a37397a );
 a37402a <=( a37401a  and  a37394a );
 a37406a <=( (not A167)  and  A168 );
 a37407a <=( A169  and  a37406a );
 a37410a <=( (not A199)  and  A166 );
 a37413a <=( A203  and  (not A200) );
 a37414a <=( a37413a  and  a37410a );
 a37415a <=( a37414a  and  a37407a );
 a37418a <=( A233  and  (not A232) );
 a37421a <=( A236  and  (not A235) );
 a37422a <=( a37421a  and  a37418a );
 a37425a <=( A299  and  (not A298) );
 a37428a <=( A302  and  (not A301) );
 a37429a <=( a37428a  and  a37425a );
 a37430a <=( a37429a  and  a37422a );
 a37434a <=( (not A167)  and  A168 );
 a37435a <=( A169  and  a37434a );
 a37438a <=( (not A199)  and  A166 );
 a37441a <=( A203  and  (not A200) );
 a37442a <=( a37441a  and  a37438a );
 a37443a <=( a37442a  and  a37435a );
 a37446a <=( A233  and  (not A232) );
 a37449a <=( A236  and  (not A235) );
 a37450a <=( a37449a  and  a37446a );
 a37453a <=( (not A299)  and  (not A298) );
 a37456a <=( (not A302)  and  A301 );
 a37457a <=( a37456a  and  a37453a );
 a37458a <=( a37457a  and  a37450a );
 a37462a <=( (not A167)  and  A168 );
 a37463a <=( A169  and  a37462a );
 a37466a <=( (not A199)  and  A166 );
 a37469a <=( A203  and  (not A200) );
 a37470a <=( a37469a  and  a37466a );
 a37471a <=( a37470a  and  a37463a );
 a37474a <=( A233  and  (not A232) );
 a37477a <=( A236  and  (not A235) );
 a37478a <=( a37477a  and  a37474a );
 a37481a <=( A266  and  A265 );
 a37484a <=( (not A269)  and  A268 );
 a37485a <=( a37484a  and  a37481a );
 a37486a <=( a37485a  and  a37478a );
 a37490a <=( (not A167)  and  A168 );
 a37491a <=( A169  and  a37490a );
 a37494a <=( (not A199)  and  A166 );
 a37497a <=( A203  and  (not A200) );
 a37498a <=( a37497a  and  a37494a );
 a37499a <=( a37498a  and  a37491a );
 a37502a <=( A233  and  (not A232) );
 a37505a <=( A236  and  (not A235) );
 a37506a <=( a37505a  and  a37502a );
 a37509a <=( A266  and  (not A265) );
 a37512a <=( A269  and  (not A268) );
 a37513a <=( a37512a  and  a37509a );
 a37514a <=( a37513a  and  a37506a );
 a37518a <=( (not A167)  and  A168 );
 a37519a <=( A169  and  a37518a );
 a37522a <=( (not A199)  and  A166 );
 a37525a <=( A203  and  (not A200) );
 a37526a <=( a37525a  and  a37522a );
 a37527a <=( a37526a  and  a37519a );
 a37530a <=( A233  and  (not A232) );
 a37533a <=( A236  and  (not A235) );
 a37534a <=( a37533a  and  a37530a );
 a37537a <=( (not A266)  and  A265 );
 a37540a <=( A269  and  (not A268) );
 a37541a <=( a37540a  and  a37537a );
 a37542a <=( a37541a  and  a37534a );
 a37546a <=( (not A167)  and  A168 );
 a37547a <=( A169  and  a37546a );
 a37550a <=( (not A199)  and  A166 );
 a37553a <=( A203  and  (not A200) );
 a37554a <=( a37553a  and  a37550a );
 a37555a <=( a37554a  and  a37547a );
 a37558a <=( A233  and  (not A232) );
 a37561a <=( A236  and  (not A235) );
 a37562a <=( a37561a  and  a37558a );
 a37565a <=( (not A266)  and  (not A265) );
 a37568a <=( (not A269)  and  A268 );
 a37569a <=( a37568a  and  a37565a );
 a37570a <=( a37569a  and  a37562a );
 a37574a <=( (not A167)  and  A168 );
 a37575a <=( A169  and  a37574a );
 a37578a <=( (not A199)  and  A166 );
 a37581a <=( A203  and  (not A200) );
 a37582a <=( a37581a  and  a37578a );
 a37583a <=( a37582a  and  a37575a );
 a37586a <=( (not A233)  and  A232 );
 a37589a <=( A236  and  (not A235) );
 a37590a <=( a37589a  and  a37586a );
 a37593a <=( A299  and  A298 );
 a37596a <=( (not A302)  and  A301 );
 a37597a <=( a37596a  and  a37593a );
 a37598a <=( a37597a  and  a37590a );
 a37602a <=( (not A167)  and  A168 );
 a37603a <=( A169  and  a37602a );
 a37606a <=( (not A199)  and  A166 );
 a37609a <=( A203  and  (not A200) );
 a37610a <=( a37609a  and  a37606a );
 a37611a <=( a37610a  and  a37603a );
 a37614a <=( (not A233)  and  A232 );
 a37617a <=( A236  and  (not A235) );
 a37618a <=( a37617a  and  a37614a );
 a37621a <=( (not A299)  and  A298 );
 a37624a <=( A302  and  (not A301) );
 a37625a <=( a37624a  and  a37621a );
 a37626a <=( a37625a  and  a37618a );
 a37630a <=( (not A167)  and  A168 );
 a37631a <=( A169  and  a37630a );
 a37634a <=( (not A199)  and  A166 );
 a37637a <=( A203  and  (not A200) );
 a37638a <=( a37637a  and  a37634a );
 a37639a <=( a37638a  and  a37631a );
 a37642a <=( (not A233)  and  A232 );
 a37645a <=( A236  and  (not A235) );
 a37646a <=( a37645a  and  a37642a );
 a37649a <=( A299  and  (not A298) );
 a37652a <=( A302  and  (not A301) );
 a37653a <=( a37652a  and  a37649a );
 a37654a <=( a37653a  and  a37646a );
 a37658a <=( (not A167)  and  A168 );
 a37659a <=( A169  and  a37658a );
 a37662a <=( (not A199)  and  A166 );
 a37665a <=( A203  and  (not A200) );
 a37666a <=( a37665a  and  a37662a );
 a37667a <=( a37666a  and  a37659a );
 a37670a <=( (not A233)  and  A232 );
 a37673a <=( A236  and  (not A235) );
 a37674a <=( a37673a  and  a37670a );
 a37677a <=( (not A299)  and  (not A298) );
 a37680a <=( (not A302)  and  A301 );
 a37681a <=( a37680a  and  a37677a );
 a37682a <=( a37681a  and  a37674a );
 a37686a <=( (not A167)  and  A168 );
 a37687a <=( A169  and  a37686a );
 a37690a <=( (not A199)  and  A166 );
 a37693a <=( A203  and  (not A200) );
 a37694a <=( a37693a  and  a37690a );
 a37695a <=( a37694a  and  a37687a );
 a37698a <=( (not A233)  and  A232 );
 a37701a <=( A236  and  (not A235) );
 a37702a <=( a37701a  and  a37698a );
 a37705a <=( A266  and  A265 );
 a37708a <=( (not A269)  and  A268 );
 a37709a <=( a37708a  and  a37705a );
 a37710a <=( a37709a  and  a37702a );
 a37714a <=( (not A167)  and  A168 );
 a37715a <=( A169  and  a37714a );
 a37718a <=( (not A199)  and  A166 );
 a37721a <=( A203  and  (not A200) );
 a37722a <=( a37721a  and  a37718a );
 a37723a <=( a37722a  and  a37715a );
 a37726a <=( (not A233)  and  A232 );
 a37729a <=( A236  and  (not A235) );
 a37730a <=( a37729a  and  a37726a );
 a37733a <=( A266  and  (not A265) );
 a37736a <=( A269  and  (not A268) );
 a37737a <=( a37736a  and  a37733a );
 a37738a <=( a37737a  and  a37730a );
 a37742a <=( (not A167)  and  A168 );
 a37743a <=( A169  and  a37742a );
 a37746a <=( (not A199)  and  A166 );
 a37749a <=( A203  and  (not A200) );
 a37750a <=( a37749a  and  a37746a );
 a37751a <=( a37750a  and  a37743a );
 a37754a <=( (not A233)  and  A232 );
 a37757a <=( A236  and  (not A235) );
 a37758a <=( a37757a  and  a37754a );
 a37761a <=( (not A266)  and  A265 );
 a37764a <=( A269  and  (not A268) );
 a37765a <=( a37764a  and  a37761a );
 a37766a <=( a37765a  and  a37758a );
 a37770a <=( (not A167)  and  A168 );
 a37771a <=( A169  and  a37770a );
 a37774a <=( (not A199)  and  A166 );
 a37777a <=( A203  and  (not A200) );
 a37778a <=( a37777a  and  a37774a );
 a37779a <=( a37778a  and  a37771a );
 a37782a <=( (not A233)  and  A232 );
 a37785a <=( A236  and  (not A235) );
 a37786a <=( a37785a  and  a37782a );
 a37789a <=( (not A266)  and  (not A265) );
 a37792a <=( (not A269)  and  A268 );
 a37793a <=( a37792a  and  a37789a );
 a37794a <=( a37793a  and  a37786a );
 a37798a <=( (not A167)  and  A168 );
 a37799a <=( A169  and  a37798a );
 a37802a <=( (not A199)  and  A166 );
 a37805a <=( A203  and  (not A200) );
 a37806a <=( a37805a  and  a37802a );
 a37807a <=( a37806a  and  a37799a );
 a37810a <=( (not A233)  and  (not A232) );
 a37813a <=( (not A236)  and  A235 );
 a37814a <=( a37813a  and  a37810a );
 a37817a <=( A299  and  A298 );
 a37820a <=( (not A302)  and  A301 );
 a37821a <=( a37820a  and  a37817a );
 a37822a <=( a37821a  and  a37814a );
 a37826a <=( (not A167)  and  A168 );
 a37827a <=( A169  and  a37826a );
 a37830a <=( (not A199)  and  A166 );
 a37833a <=( A203  and  (not A200) );
 a37834a <=( a37833a  and  a37830a );
 a37835a <=( a37834a  and  a37827a );
 a37838a <=( (not A233)  and  (not A232) );
 a37841a <=( (not A236)  and  A235 );
 a37842a <=( a37841a  and  a37838a );
 a37845a <=( (not A299)  and  A298 );
 a37848a <=( A302  and  (not A301) );
 a37849a <=( a37848a  and  a37845a );
 a37850a <=( a37849a  and  a37842a );
 a37854a <=( (not A167)  and  A168 );
 a37855a <=( A169  and  a37854a );
 a37858a <=( (not A199)  and  A166 );
 a37861a <=( A203  and  (not A200) );
 a37862a <=( a37861a  and  a37858a );
 a37863a <=( a37862a  and  a37855a );
 a37866a <=( (not A233)  and  (not A232) );
 a37869a <=( (not A236)  and  A235 );
 a37870a <=( a37869a  and  a37866a );
 a37873a <=( A299  and  (not A298) );
 a37876a <=( A302  and  (not A301) );
 a37877a <=( a37876a  and  a37873a );
 a37878a <=( a37877a  and  a37870a );
 a37882a <=( (not A167)  and  A168 );
 a37883a <=( A169  and  a37882a );
 a37886a <=( (not A199)  and  A166 );
 a37889a <=( A203  and  (not A200) );
 a37890a <=( a37889a  and  a37886a );
 a37891a <=( a37890a  and  a37883a );
 a37894a <=( (not A233)  and  (not A232) );
 a37897a <=( (not A236)  and  A235 );
 a37898a <=( a37897a  and  a37894a );
 a37901a <=( (not A299)  and  (not A298) );
 a37904a <=( (not A302)  and  A301 );
 a37905a <=( a37904a  and  a37901a );
 a37906a <=( a37905a  and  a37898a );
 a37910a <=( (not A167)  and  A168 );
 a37911a <=( A169  and  a37910a );
 a37914a <=( (not A199)  and  A166 );
 a37917a <=( A203  and  (not A200) );
 a37918a <=( a37917a  and  a37914a );
 a37919a <=( a37918a  and  a37911a );
 a37922a <=( (not A233)  and  (not A232) );
 a37925a <=( (not A236)  and  A235 );
 a37926a <=( a37925a  and  a37922a );
 a37929a <=( A266  and  A265 );
 a37932a <=( (not A269)  and  A268 );
 a37933a <=( a37932a  and  a37929a );
 a37934a <=( a37933a  and  a37926a );
 a37938a <=( (not A167)  and  A168 );
 a37939a <=( A169  and  a37938a );
 a37942a <=( (not A199)  and  A166 );
 a37945a <=( A203  and  (not A200) );
 a37946a <=( a37945a  and  a37942a );
 a37947a <=( a37946a  and  a37939a );
 a37950a <=( (not A233)  and  (not A232) );
 a37953a <=( (not A236)  and  A235 );
 a37954a <=( a37953a  and  a37950a );
 a37957a <=( A266  and  (not A265) );
 a37960a <=( A269  and  (not A268) );
 a37961a <=( a37960a  and  a37957a );
 a37962a <=( a37961a  and  a37954a );
 a37966a <=( (not A167)  and  A168 );
 a37967a <=( A169  and  a37966a );
 a37970a <=( (not A199)  and  A166 );
 a37973a <=( A203  and  (not A200) );
 a37974a <=( a37973a  and  a37970a );
 a37975a <=( a37974a  and  a37967a );
 a37978a <=( (not A233)  and  (not A232) );
 a37981a <=( (not A236)  and  A235 );
 a37982a <=( a37981a  and  a37978a );
 a37985a <=( (not A266)  and  A265 );
 a37988a <=( A269  and  (not A268) );
 a37989a <=( a37988a  and  a37985a );
 a37990a <=( a37989a  and  a37982a );
 a37994a <=( (not A167)  and  A168 );
 a37995a <=( A169  and  a37994a );
 a37998a <=( (not A199)  and  A166 );
 a38001a <=( A203  and  (not A200) );
 a38002a <=( a38001a  and  a37998a );
 a38003a <=( a38002a  and  a37995a );
 a38006a <=( (not A233)  and  (not A232) );
 a38009a <=( (not A236)  and  A235 );
 a38010a <=( a38009a  and  a38006a );
 a38013a <=( (not A266)  and  (not A265) );
 a38016a <=( (not A269)  and  A268 );
 a38017a <=( a38016a  and  a38013a );
 a38018a <=( a38017a  and  a38010a );
 a38021a <=( A168  and  A170 );
 a38024a <=( A166  and  (not A167) );
 a38025a <=( a38024a  and  a38021a );
 a38028a <=( A200  and  A199 );
 a38031a <=( (not A202)  and  (not A201) );
 a38032a <=( a38031a  and  a38028a );
 a38033a <=( a38032a  and  a38025a );
 a38036a <=( A233  and  A232 );
 a38039a <=( (not A236)  and  A235 );
 a38040a <=( a38039a  and  a38036a );
 a38043a <=( A299  and  A298 );
 a38046a <=( (not A302)  and  A301 );
 a38047a <=( a38046a  and  a38043a );
 a38048a <=( a38047a  and  a38040a );
 a38051a <=( A168  and  A170 );
 a38054a <=( A166  and  (not A167) );
 a38055a <=( a38054a  and  a38051a );
 a38058a <=( A200  and  A199 );
 a38061a <=( (not A202)  and  (not A201) );
 a38062a <=( a38061a  and  a38058a );
 a38063a <=( a38062a  and  a38055a );
 a38066a <=( A233  and  A232 );
 a38069a <=( (not A236)  and  A235 );
 a38070a <=( a38069a  and  a38066a );
 a38073a <=( (not A299)  and  A298 );
 a38076a <=( A302  and  (not A301) );
 a38077a <=( a38076a  and  a38073a );
 a38078a <=( a38077a  and  a38070a );
 a38081a <=( A168  and  A170 );
 a38084a <=( A166  and  (not A167) );
 a38085a <=( a38084a  and  a38081a );
 a38088a <=( A200  and  A199 );
 a38091a <=( (not A202)  and  (not A201) );
 a38092a <=( a38091a  and  a38088a );
 a38093a <=( a38092a  and  a38085a );
 a38096a <=( A233  and  A232 );
 a38099a <=( (not A236)  and  A235 );
 a38100a <=( a38099a  and  a38096a );
 a38103a <=( A299  and  (not A298) );
 a38106a <=( A302  and  (not A301) );
 a38107a <=( a38106a  and  a38103a );
 a38108a <=( a38107a  and  a38100a );
 a38111a <=( A168  and  A170 );
 a38114a <=( A166  and  (not A167) );
 a38115a <=( a38114a  and  a38111a );
 a38118a <=( A200  and  A199 );
 a38121a <=( (not A202)  and  (not A201) );
 a38122a <=( a38121a  and  a38118a );
 a38123a <=( a38122a  and  a38115a );
 a38126a <=( A233  and  A232 );
 a38129a <=( (not A236)  and  A235 );
 a38130a <=( a38129a  and  a38126a );
 a38133a <=( (not A299)  and  (not A298) );
 a38136a <=( (not A302)  and  A301 );
 a38137a <=( a38136a  and  a38133a );
 a38138a <=( a38137a  and  a38130a );
 a38141a <=( A168  and  A170 );
 a38144a <=( A166  and  (not A167) );
 a38145a <=( a38144a  and  a38141a );
 a38148a <=( A200  and  A199 );
 a38151a <=( (not A202)  and  (not A201) );
 a38152a <=( a38151a  and  a38148a );
 a38153a <=( a38152a  and  a38145a );
 a38156a <=( A233  and  A232 );
 a38159a <=( (not A236)  and  A235 );
 a38160a <=( a38159a  and  a38156a );
 a38163a <=( A266  and  A265 );
 a38166a <=( (not A269)  and  A268 );
 a38167a <=( a38166a  and  a38163a );
 a38168a <=( a38167a  and  a38160a );
 a38171a <=( A168  and  A170 );
 a38174a <=( A166  and  (not A167) );
 a38175a <=( a38174a  and  a38171a );
 a38178a <=( A200  and  A199 );
 a38181a <=( (not A202)  and  (not A201) );
 a38182a <=( a38181a  and  a38178a );
 a38183a <=( a38182a  and  a38175a );
 a38186a <=( A233  and  A232 );
 a38189a <=( (not A236)  and  A235 );
 a38190a <=( a38189a  and  a38186a );
 a38193a <=( A266  and  (not A265) );
 a38196a <=( A269  and  (not A268) );
 a38197a <=( a38196a  and  a38193a );
 a38198a <=( a38197a  and  a38190a );
 a38201a <=( A168  and  A170 );
 a38204a <=( A166  and  (not A167) );
 a38205a <=( a38204a  and  a38201a );
 a38208a <=( A200  and  A199 );
 a38211a <=( (not A202)  and  (not A201) );
 a38212a <=( a38211a  and  a38208a );
 a38213a <=( a38212a  and  a38205a );
 a38216a <=( A233  and  A232 );
 a38219a <=( (not A236)  and  A235 );
 a38220a <=( a38219a  and  a38216a );
 a38223a <=( (not A266)  and  A265 );
 a38226a <=( A269  and  (not A268) );
 a38227a <=( a38226a  and  a38223a );
 a38228a <=( a38227a  and  a38220a );
 a38231a <=( A168  and  A170 );
 a38234a <=( A166  and  (not A167) );
 a38235a <=( a38234a  and  a38231a );
 a38238a <=( A200  and  A199 );
 a38241a <=( (not A202)  and  (not A201) );
 a38242a <=( a38241a  and  a38238a );
 a38243a <=( a38242a  and  a38235a );
 a38246a <=( A233  and  A232 );
 a38249a <=( (not A236)  and  A235 );
 a38250a <=( a38249a  and  a38246a );
 a38253a <=( (not A266)  and  (not A265) );
 a38256a <=( (not A269)  and  A268 );
 a38257a <=( a38256a  and  a38253a );
 a38258a <=( a38257a  and  a38250a );
 a38261a <=( A168  and  A170 );
 a38264a <=( A166  and  (not A167) );
 a38265a <=( a38264a  and  a38261a );
 a38268a <=( A200  and  A199 );
 a38271a <=( (not A202)  and  (not A201) );
 a38272a <=( a38271a  and  a38268a );
 a38273a <=( a38272a  and  a38265a );
 a38276a <=( A233  and  (not A232) );
 a38279a <=( A236  and  (not A235) );
 a38280a <=( a38279a  and  a38276a );
 a38283a <=( A299  and  A298 );
 a38286a <=( (not A302)  and  A301 );
 a38287a <=( a38286a  and  a38283a );
 a38288a <=( a38287a  and  a38280a );
 a38291a <=( A168  and  A170 );
 a38294a <=( A166  and  (not A167) );
 a38295a <=( a38294a  and  a38291a );
 a38298a <=( A200  and  A199 );
 a38301a <=( (not A202)  and  (not A201) );
 a38302a <=( a38301a  and  a38298a );
 a38303a <=( a38302a  and  a38295a );
 a38306a <=( A233  and  (not A232) );
 a38309a <=( A236  and  (not A235) );
 a38310a <=( a38309a  and  a38306a );
 a38313a <=( (not A299)  and  A298 );
 a38316a <=( A302  and  (not A301) );
 a38317a <=( a38316a  and  a38313a );
 a38318a <=( a38317a  and  a38310a );
 a38321a <=( A168  and  A170 );
 a38324a <=( A166  and  (not A167) );
 a38325a <=( a38324a  and  a38321a );
 a38328a <=( A200  and  A199 );
 a38331a <=( (not A202)  and  (not A201) );
 a38332a <=( a38331a  and  a38328a );
 a38333a <=( a38332a  and  a38325a );
 a38336a <=( A233  and  (not A232) );
 a38339a <=( A236  and  (not A235) );
 a38340a <=( a38339a  and  a38336a );
 a38343a <=( A299  and  (not A298) );
 a38346a <=( A302  and  (not A301) );
 a38347a <=( a38346a  and  a38343a );
 a38348a <=( a38347a  and  a38340a );
 a38351a <=( A168  and  A170 );
 a38354a <=( A166  and  (not A167) );
 a38355a <=( a38354a  and  a38351a );
 a38358a <=( A200  and  A199 );
 a38361a <=( (not A202)  and  (not A201) );
 a38362a <=( a38361a  and  a38358a );
 a38363a <=( a38362a  and  a38355a );
 a38366a <=( A233  and  (not A232) );
 a38369a <=( A236  and  (not A235) );
 a38370a <=( a38369a  and  a38366a );
 a38373a <=( (not A299)  and  (not A298) );
 a38376a <=( (not A302)  and  A301 );
 a38377a <=( a38376a  and  a38373a );
 a38378a <=( a38377a  and  a38370a );
 a38381a <=( A168  and  A170 );
 a38384a <=( A166  and  (not A167) );
 a38385a <=( a38384a  and  a38381a );
 a38388a <=( A200  and  A199 );
 a38391a <=( (not A202)  and  (not A201) );
 a38392a <=( a38391a  and  a38388a );
 a38393a <=( a38392a  and  a38385a );
 a38396a <=( A233  and  (not A232) );
 a38399a <=( A236  and  (not A235) );
 a38400a <=( a38399a  and  a38396a );
 a38403a <=( A266  and  A265 );
 a38406a <=( (not A269)  and  A268 );
 a38407a <=( a38406a  and  a38403a );
 a38408a <=( a38407a  and  a38400a );
 a38411a <=( A168  and  A170 );
 a38414a <=( A166  and  (not A167) );
 a38415a <=( a38414a  and  a38411a );
 a38418a <=( A200  and  A199 );
 a38421a <=( (not A202)  and  (not A201) );
 a38422a <=( a38421a  and  a38418a );
 a38423a <=( a38422a  and  a38415a );
 a38426a <=( A233  and  (not A232) );
 a38429a <=( A236  and  (not A235) );
 a38430a <=( a38429a  and  a38426a );
 a38433a <=( A266  and  (not A265) );
 a38436a <=( A269  and  (not A268) );
 a38437a <=( a38436a  and  a38433a );
 a38438a <=( a38437a  and  a38430a );
 a38441a <=( A168  and  A170 );
 a38444a <=( A166  and  (not A167) );
 a38445a <=( a38444a  and  a38441a );
 a38448a <=( A200  and  A199 );
 a38451a <=( (not A202)  and  (not A201) );
 a38452a <=( a38451a  and  a38448a );
 a38453a <=( a38452a  and  a38445a );
 a38456a <=( A233  and  (not A232) );
 a38459a <=( A236  and  (not A235) );
 a38460a <=( a38459a  and  a38456a );
 a38463a <=( (not A266)  and  A265 );
 a38466a <=( A269  and  (not A268) );
 a38467a <=( a38466a  and  a38463a );
 a38468a <=( a38467a  and  a38460a );
 a38471a <=( A168  and  A170 );
 a38474a <=( A166  and  (not A167) );
 a38475a <=( a38474a  and  a38471a );
 a38478a <=( A200  and  A199 );
 a38481a <=( (not A202)  and  (not A201) );
 a38482a <=( a38481a  and  a38478a );
 a38483a <=( a38482a  and  a38475a );
 a38486a <=( A233  and  (not A232) );
 a38489a <=( A236  and  (not A235) );
 a38490a <=( a38489a  and  a38486a );
 a38493a <=( (not A266)  and  (not A265) );
 a38496a <=( (not A269)  and  A268 );
 a38497a <=( a38496a  and  a38493a );
 a38498a <=( a38497a  and  a38490a );
 a38501a <=( A168  and  A170 );
 a38504a <=( A166  and  (not A167) );
 a38505a <=( a38504a  and  a38501a );
 a38508a <=( A200  and  A199 );
 a38511a <=( (not A202)  and  (not A201) );
 a38512a <=( a38511a  and  a38508a );
 a38513a <=( a38512a  and  a38505a );
 a38516a <=( (not A233)  and  A232 );
 a38519a <=( A236  and  (not A235) );
 a38520a <=( a38519a  and  a38516a );
 a38523a <=( A299  and  A298 );
 a38526a <=( (not A302)  and  A301 );
 a38527a <=( a38526a  and  a38523a );
 a38528a <=( a38527a  and  a38520a );
 a38531a <=( A168  and  A170 );
 a38534a <=( A166  and  (not A167) );
 a38535a <=( a38534a  and  a38531a );
 a38538a <=( A200  and  A199 );
 a38541a <=( (not A202)  and  (not A201) );
 a38542a <=( a38541a  and  a38538a );
 a38543a <=( a38542a  and  a38535a );
 a38546a <=( (not A233)  and  A232 );
 a38549a <=( A236  and  (not A235) );
 a38550a <=( a38549a  and  a38546a );
 a38553a <=( (not A299)  and  A298 );
 a38556a <=( A302  and  (not A301) );
 a38557a <=( a38556a  and  a38553a );
 a38558a <=( a38557a  and  a38550a );
 a38561a <=( A168  and  A170 );
 a38564a <=( A166  and  (not A167) );
 a38565a <=( a38564a  and  a38561a );
 a38568a <=( A200  and  A199 );
 a38571a <=( (not A202)  and  (not A201) );
 a38572a <=( a38571a  and  a38568a );
 a38573a <=( a38572a  and  a38565a );
 a38576a <=( (not A233)  and  A232 );
 a38579a <=( A236  and  (not A235) );
 a38580a <=( a38579a  and  a38576a );
 a38583a <=( A299  and  (not A298) );
 a38586a <=( A302  and  (not A301) );
 a38587a <=( a38586a  and  a38583a );
 a38588a <=( a38587a  and  a38580a );
 a38591a <=( A168  and  A170 );
 a38594a <=( A166  and  (not A167) );
 a38595a <=( a38594a  and  a38591a );
 a38598a <=( A200  and  A199 );
 a38601a <=( (not A202)  and  (not A201) );
 a38602a <=( a38601a  and  a38598a );
 a38603a <=( a38602a  and  a38595a );
 a38606a <=( (not A233)  and  A232 );
 a38609a <=( A236  and  (not A235) );
 a38610a <=( a38609a  and  a38606a );
 a38613a <=( (not A299)  and  (not A298) );
 a38616a <=( (not A302)  and  A301 );
 a38617a <=( a38616a  and  a38613a );
 a38618a <=( a38617a  and  a38610a );
 a38621a <=( A168  and  A170 );
 a38624a <=( A166  and  (not A167) );
 a38625a <=( a38624a  and  a38621a );
 a38628a <=( A200  and  A199 );
 a38631a <=( (not A202)  and  (not A201) );
 a38632a <=( a38631a  and  a38628a );
 a38633a <=( a38632a  and  a38625a );
 a38636a <=( (not A233)  and  A232 );
 a38639a <=( A236  and  (not A235) );
 a38640a <=( a38639a  and  a38636a );
 a38643a <=( A266  and  A265 );
 a38646a <=( (not A269)  and  A268 );
 a38647a <=( a38646a  and  a38643a );
 a38648a <=( a38647a  and  a38640a );
 a38651a <=( A168  and  A170 );
 a38654a <=( A166  and  (not A167) );
 a38655a <=( a38654a  and  a38651a );
 a38658a <=( A200  and  A199 );
 a38661a <=( (not A202)  and  (not A201) );
 a38662a <=( a38661a  and  a38658a );
 a38663a <=( a38662a  and  a38655a );
 a38666a <=( (not A233)  and  A232 );
 a38669a <=( A236  and  (not A235) );
 a38670a <=( a38669a  and  a38666a );
 a38673a <=( A266  and  (not A265) );
 a38676a <=( A269  and  (not A268) );
 a38677a <=( a38676a  and  a38673a );
 a38678a <=( a38677a  and  a38670a );
 a38681a <=( A168  and  A170 );
 a38684a <=( A166  and  (not A167) );
 a38685a <=( a38684a  and  a38681a );
 a38688a <=( A200  and  A199 );
 a38691a <=( (not A202)  and  (not A201) );
 a38692a <=( a38691a  and  a38688a );
 a38693a <=( a38692a  and  a38685a );
 a38696a <=( (not A233)  and  A232 );
 a38699a <=( A236  and  (not A235) );
 a38700a <=( a38699a  and  a38696a );
 a38703a <=( (not A266)  and  A265 );
 a38706a <=( A269  and  (not A268) );
 a38707a <=( a38706a  and  a38703a );
 a38708a <=( a38707a  and  a38700a );
 a38711a <=( A168  and  A170 );
 a38714a <=( A166  and  (not A167) );
 a38715a <=( a38714a  and  a38711a );
 a38718a <=( A200  and  A199 );
 a38721a <=( (not A202)  and  (not A201) );
 a38722a <=( a38721a  and  a38718a );
 a38723a <=( a38722a  and  a38715a );
 a38726a <=( (not A233)  and  A232 );
 a38729a <=( A236  and  (not A235) );
 a38730a <=( a38729a  and  a38726a );
 a38733a <=( (not A266)  and  (not A265) );
 a38736a <=( (not A269)  and  A268 );
 a38737a <=( a38736a  and  a38733a );
 a38738a <=( a38737a  and  a38730a );
 a38741a <=( A168  and  A170 );
 a38744a <=( A166  and  (not A167) );
 a38745a <=( a38744a  and  a38741a );
 a38748a <=( A200  and  A199 );
 a38751a <=( (not A202)  and  (not A201) );
 a38752a <=( a38751a  and  a38748a );
 a38753a <=( a38752a  and  a38745a );
 a38756a <=( (not A233)  and  (not A232) );
 a38759a <=( (not A236)  and  A235 );
 a38760a <=( a38759a  and  a38756a );
 a38763a <=( A299  and  A298 );
 a38766a <=( (not A302)  and  A301 );
 a38767a <=( a38766a  and  a38763a );
 a38768a <=( a38767a  and  a38760a );
 a38771a <=( A168  and  A170 );
 a38774a <=( A166  and  (not A167) );
 a38775a <=( a38774a  and  a38771a );
 a38778a <=( A200  and  A199 );
 a38781a <=( (not A202)  and  (not A201) );
 a38782a <=( a38781a  and  a38778a );
 a38783a <=( a38782a  and  a38775a );
 a38786a <=( (not A233)  and  (not A232) );
 a38789a <=( (not A236)  and  A235 );
 a38790a <=( a38789a  and  a38786a );
 a38793a <=( (not A299)  and  A298 );
 a38796a <=( A302  and  (not A301) );
 a38797a <=( a38796a  and  a38793a );
 a38798a <=( a38797a  and  a38790a );
 a38801a <=( A168  and  A170 );
 a38804a <=( A166  and  (not A167) );
 a38805a <=( a38804a  and  a38801a );
 a38808a <=( A200  and  A199 );
 a38811a <=( (not A202)  and  (not A201) );
 a38812a <=( a38811a  and  a38808a );
 a38813a <=( a38812a  and  a38805a );
 a38816a <=( (not A233)  and  (not A232) );
 a38819a <=( (not A236)  and  A235 );
 a38820a <=( a38819a  and  a38816a );
 a38823a <=( A299  and  (not A298) );
 a38826a <=( A302  and  (not A301) );
 a38827a <=( a38826a  and  a38823a );
 a38828a <=( a38827a  and  a38820a );
 a38831a <=( A168  and  A170 );
 a38834a <=( A166  and  (not A167) );
 a38835a <=( a38834a  and  a38831a );
 a38838a <=( A200  and  A199 );
 a38841a <=( (not A202)  and  (not A201) );
 a38842a <=( a38841a  and  a38838a );
 a38843a <=( a38842a  and  a38835a );
 a38846a <=( (not A233)  and  (not A232) );
 a38849a <=( (not A236)  and  A235 );
 a38850a <=( a38849a  and  a38846a );
 a38853a <=( (not A299)  and  (not A298) );
 a38856a <=( (not A302)  and  A301 );
 a38857a <=( a38856a  and  a38853a );
 a38858a <=( a38857a  and  a38850a );
 a38861a <=( A168  and  A170 );
 a38864a <=( A166  and  (not A167) );
 a38865a <=( a38864a  and  a38861a );
 a38868a <=( A200  and  A199 );
 a38871a <=( (not A202)  and  (not A201) );
 a38872a <=( a38871a  and  a38868a );
 a38873a <=( a38872a  and  a38865a );
 a38876a <=( (not A233)  and  (not A232) );
 a38879a <=( (not A236)  and  A235 );
 a38880a <=( a38879a  and  a38876a );
 a38883a <=( A266  and  A265 );
 a38886a <=( (not A269)  and  A268 );
 a38887a <=( a38886a  and  a38883a );
 a38888a <=( a38887a  and  a38880a );
 a38891a <=( A168  and  A170 );
 a38894a <=( A166  and  (not A167) );
 a38895a <=( a38894a  and  a38891a );
 a38898a <=( A200  and  A199 );
 a38901a <=( (not A202)  and  (not A201) );
 a38902a <=( a38901a  and  a38898a );
 a38903a <=( a38902a  and  a38895a );
 a38906a <=( (not A233)  and  (not A232) );
 a38909a <=( (not A236)  and  A235 );
 a38910a <=( a38909a  and  a38906a );
 a38913a <=( A266  and  (not A265) );
 a38916a <=( A269  and  (not A268) );
 a38917a <=( a38916a  and  a38913a );
 a38918a <=( a38917a  and  a38910a );
 a38921a <=( A168  and  A170 );
 a38924a <=( A166  and  (not A167) );
 a38925a <=( a38924a  and  a38921a );
 a38928a <=( A200  and  A199 );
 a38931a <=( (not A202)  and  (not A201) );
 a38932a <=( a38931a  and  a38928a );
 a38933a <=( a38932a  and  a38925a );
 a38936a <=( (not A233)  and  (not A232) );
 a38939a <=( (not A236)  and  A235 );
 a38940a <=( a38939a  and  a38936a );
 a38943a <=( (not A266)  and  A265 );
 a38946a <=( A269  and  (not A268) );
 a38947a <=( a38946a  and  a38943a );
 a38948a <=( a38947a  and  a38940a );
 a38951a <=( A168  and  A170 );
 a38954a <=( A166  and  (not A167) );
 a38955a <=( a38954a  and  a38951a );
 a38958a <=( A200  and  A199 );
 a38961a <=( (not A202)  and  (not A201) );
 a38962a <=( a38961a  and  a38958a );
 a38963a <=( a38962a  and  a38955a );
 a38966a <=( (not A233)  and  (not A232) );
 a38969a <=( (not A236)  and  A235 );
 a38970a <=( a38969a  and  a38966a );
 a38973a <=( (not A266)  and  (not A265) );
 a38976a <=( (not A269)  and  A268 );
 a38977a <=( a38976a  and  a38973a );
 a38978a <=( a38977a  and  a38970a );
 a38981a <=( A168  and  A170 );
 a38984a <=( A166  and  (not A167) );
 a38985a <=( a38984a  and  a38981a );
 a38988a <=( A200  and  A199 );
 a38991a <=( A203  and  (not A201) );
 a38992a <=( a38991a  and  a38988a );
 a38993a <=( a38992a  and  a38985a );
 a38996a <=( A233  and  A232 );
 a38999a <=( (not A236)  and  A235 );
 a39000a <=( a38999a  and  a38996a );
 a39003a <=( A299  and  A298 );
 a39006a <=( (not A302)  and  A301 );
 a39007a <=( a39006a  and  a39003a );
 a39008a <=( a39007a  and  a39000a );
 a39011a <=( A168  and  A170 );
 a39014a <=( A166  and  (not A167) );
 a39015a <=( a39014a  and  a39011a );
 a39018a <=( A200  and  A199 );
 a39021a <=( A203  and  (not A201) );
 a39022a <=( a39021a  and  a39018a );
 a39023a <=( a39022a  and  a39015a );
 a39026a <=( A233  and  A232 );
 a39029a <=( (not A236)  and  A235 );
 a39030a <=( a39029a  and  a39026a );
 a39033a <=( (not A299)  and  A298 );
 a39036a <=( A302  and  (not A301) );
 a39037a <=( a39036a  and  a39033a );
 a39038a <=( a39037a  and  a39030a );
 a39041a <=( A168  and  A170 );
 a39044a <=( A166  and  (not A167) );
 a39045a <=( a39044a  and  a39041a );
 a39048a <=( A200  and  A199 );
 a39051a <=( A203  and  (not A201) );
 a39052a <=( a39051a  and  a39048a );
 a39053a <=( a39052a  and  a39045a );
 a39056a <=( A233  and  A232 );
 a39059a <=( (not A236)  and  A235 );
 a39060a <=( a39059a  and  a39056a );
 a39063a <=( A299  and  (not A298) );
 a39066a <=( A302  and  (not A301) );
 a39067a <=( a39066a  and  a39063a );
 a39068a <=( a39067a  and  a39060a );
 a39071a <=( A168  and  A170 );
 a39074a <=( A166  and  (not A167) );
 a39075a <=( a39074a  and  a39071a );
 a39078a <=( A200  and  A199 );
 a39081a <=( A203  and  (not A201) );
 a39082a <=( a39081a  and  a39078a );
 a39083a <=( a39082a  and  a39075a );
 a39086a <=( A233  and  A232 );
 a39089a <=( (not A236)  and  A235 );
 a39090a <=( a39089a  and  a39086a );
 a39093a <=( (not A299)  and  (not A298) );
 a39096a <=( (not A302)  and  A301 );
 a39097a <=( a39096a  and  a39093a );
 a39098a <=( a39097a  and  a39090a );
 a39101a <=( A168  and  A170 );
 a39104a <=( A166  and  (not A167) );
 a39105a <=( a39104a  and  a39101a );
 a39108a <=( A200  and  A199 );
 a39111a <=( A203  and  (not A201) );
 a39112a <=( a39111a  and  a39108a );
 a39113a <=( a39112a  and  a39105a );
 a39116a <=( A233  and  A232 );
 a39119a <=( (not A236)  and  A235 );
 a39120a <=( a39119a  and  a39116a );
 a39123a <=( A266  and  A265 );
 a39126a <=( (not A269)  and  A268 );
 a39127a <=( a39126a  and  a39123a );
 a39128a <=( a39127a  and  a39120a );
 a39131a <=( A168  and  A170 );
 a39134a <=( A166  and  (not A167) );
 a39135a <=( a39134a  and  a39131a );
 a39138a <=( A200  and  A199 );
 a39141a <=( A203  and  (not A201) );
 a39142a <=( a39141a  and  a39138a );
 a39143a <=( a39142a  and  a39135a );
 a39146a <=( A233  and  A232 );
 a39149a <=( (not A236)  and  A235 );
 a39150a <=( a39149a  and  a39146a );
 a39153a <=( A266  and  (not A265) );
 a39156a <=( A269  and  (not A268) );
 a39157a <=( a39156a  and  a39153a );
 a39158a <=( a39157a  and  a39150a );
 a39161a <=( A168  and  A170 );
 a39164a <=( A166  and  (not A167) );
 a39165a <=( a39164a  and  a39161a );
 a39168a <=( A200  and  A199 );
 a39171a <=( A203  and  (not A201) );
 a39172a <=( a39171a  and  a39168a );
 a39173a <=( a39172a  and  a39165a );
 a39176a <=( A233  and  A232 );
 a39179a <=( (not A236)  and  A235 );
 a39180a <=( a39179a  and  a39176a );
 a39183a <=( (not A266)  and  A265 );
 a39186a <=( A269  and  (not A268) );
 a39187a <=( a39186a  and  a39183a );
 a39188a <=( a39187a  and  a39180a );
 a39191a <=( A168  and  A170 );
 a39194a <=( A166  and  (not A167) );
 a39195a <=( a39194a  and  a39191a );
 a39198a <=( A200  and  A199 );
 a39201a <=( A203  and  (not A201) );
 a39202a <=( a39201a  and  a39198a );
 a39203a <=( a39202a  and  a39195a );
 a39206a <=( A233  and  A232 );
 a39209a <=( (not A236)  and  A235 );
 a39210a <=( a39209a  and  a39206a );
 a39213a <=( (not A266)  and  (not A265) );
 a39216a <=( (not A269)  and  A268 );
 a39217a <=( a39216a  and  a39213a );
 a39218a <=( a39217a  and  a39210a );
 a39221a <=( A168  and  A170 );
 a39224a <=( A166  and  (not A167) );
 a39225a <=( a39224a  and  a39221a );
 a39228a <=( A200  and  A199 );
 a39231a <=( A203  and  (not A201) );
 a39232a <=( a39231a  and  a39228a );
 a39233a <=( a39232a  and  a39225a );
 a39236a <=( A233  and  (not A232) );
 a39239a <=( A236  and  (not A235) );
 a39240a <=( a39239a  and  a39236a );
 a39243a <=( A299  and  A298 );
 a39246a <=( (not A302)  and  A301 );
 a39247a <=( a39246a  and  a39243a );
 a39248a <=( a39247a  and  a39240a );
 a39251a <=( A168  and  A170 );
 a39254a <=( A166  and  (not A167) );
 a39255a <=( a39254a  and  a39251a );
 a39258a <=( A200  and  A199 );
 a39261a <=( A203  and  (not A201) );
 a39262a <=( a39261a  and  a39258a );
 a39263a <=( a39262a  and  a39255a );
 a39266a <=( A233  and  (not A232) );
 a39269a <=( A236  and  (not A235) );
 a39270a <=( a39269a  and  a39266a );
 a39273a <=( (not A299)  and  A298 );
 a39276a <=( A302  and  (not A301) );
 a39277a <=( a39276a  and  a39273a );
 a39278a <=( a39277a  and  a39270a );
 a39281a <=( A168  and  A170 );
 a39284a <=( A166  and  (not A167) );
 a39285a <=( a39284a  and  a39281a );
 a39288a <=( A200  and  A199 );
 a39291a <=( A203  and  (not A201) );
 a39292a <=( a39291a  and  a39288a );
 a39293a <=( a39292a  and  a39285a );
 a39296a <=( A233  and  (not A232) );
 a39299a <=( A236  and  (not A235) );
 a39300a <=( a39299a  and  a39296a );
 a39303a <=( A299  and  (not A298) );
 a39306a <=( A302  and  (not A301) );
 a39307a <=( a39306a  and  a39303a );
 a39308a <=( a39307a  and  a39300a );
 a39311a <=( A168  and  A170 );
 a39314a <=( A166  and  (not A167) );
 a39315a <=( a39314a  and  a39311a );
 a39318a <=( A200  and  A199 );
 a39321a <=( A203  and  (not A201) );
 a39322a <=( a39321a  and  a39318a );
 a39323a <=( a39322a  and  a39315a );
 a39326a <=( A233  and  (not A232) );
 a39329a <=( A236  and  (not A235) );
 a39330a <=( a39329a  and  a39326a );
 a39333a <=( (not A299)  and  (not A298) );
 a39336a <=( (not A302)  and  A301 );
 a39337a <=( a39336a  and  a39333a );
 a39338a <=( a39337a  and  a39330a );
 a39341a <=( A168  and  A170 );
 a39344a <=( A166  and  (not A167) );
 a39345a <=( a39344a  and  a39341a );
 a39348a <=( A200  and  A199 );
 a39351a <=( A203  and  (not A201) );
 a39352a <=( a39351a  and  a39348a );
 a39353a <=( a39352a  and  a39345a );
 a39356a <=( A233  and  (not A232) );
 a39359a <=( A236  and  (not A235) );
 a39360a <=( a39359a  and  a39356a );
 a39363a <=( A266  and  A265 );
 a39366a <=( (not A269)  and  A268 );
 a39367a <=( a39366a  and  a39363a );
 a39368a <=( a39367a  and  a39360a );
 a39371a <=( A168  and  A170 );
 a39374a <=( A166  and  (not A167) );
 a39375a <=( a39374a  and  a39371a );
 a39378a <=( A200  and  A199 );
 a39381a <=( A203  and  (not A201) );
 a39382a <=( a39381a  and  a39378a );
 a39383a <=( a39382a  and  a39375a );
 a39386a <=( A233  and  (not A232) );
 a39389a <=( A236  and  (not A235) );
 a39390a <=( a39389a  and  a39386a );
 a39393a <=( A266  and  (not A265) );
 a39396a <=( A269  and  (not A268) );
 a39397a <=( a39396a  and  a39393a );
 a39398a <=( a39397a  and  a39390a );
 a39401a <=( A168  and  A170 );
 a39404a <=( A166  and  (not A167) );
 a39405a <=( a39404a  and  a39401a );
 a39408a <=( A200  and  A199 );
 a39411a <=( A203  and  (not A201) );
 a39412a <=( a39411a  and  a39408a );
 a39413a <=( a39412a  and  a39405a );
 a39416a <=( A233  and  (not A232) );
 a39419a <=( A236  and  (not A235) );
 a39420a <=( a39419a  and  a39416a );
 a39423a <=( (not A266)  and  A265 );
 a39426a <=( A269  and  (not A268) );
 a39427a <=( a39426a  and  a39423a );
 a39428a <=( a39427a  and  a39420a );
 a39431a <=( A168  and  A170 );
 a39434a <=( A166  and  (not A167) );
 a39435a <=( a39434a  and  a39431a );
 a39438a <=( A200  and  A199 );
 a39441a <=( A203  and  (not A201) );
 a39442a <=( a39441a  and  a39438a );
 a39443a <=( a39442a  and  a39435a );
 a39446a <=( A233  and  (not A232) );
 a39449a <=( A236  and  (not A235) );
 a39450a <=( a39449a  and  a39446a );
 a39453a <=( (not A266)  and  (not A265) );
 a39456a <=( (not A269)  and  A268 );
 a39457a <=( a39456a  and  a39453a );
 a39458a <=( a39457a  and  a39450a );
 a39461a <=( A168  and  A170 );
 a39464a <=( A166  and  (not A167) );
 a39465a <=( a39464a  and  a39461a );
 a39468a <=( A200  and  A199 );
 a39471a <=( A203  and  (not A201) );
 a39472a <=( a39471a  and  a39468a );
 a39473a <=( a39472a  and  a39465a );
 a39476a <=( (not A233)  and  A232 );
 a39479a <=( A236  and  (not A235) );
 a39480a <=( a39479a  and  a39476a );
 a39483a <=( A299  and  A298 );
 a39486a <=( (not A302)  and  A301 );
 a39487a <=( a39486a  and  a39483a );
 a39488a <=( a39487a  and  a39480a );
 a39491a <=( A168  and  A170 );
 a39494a <=( A166  and  (not A167) );
 a39495a <=( a39494a  and  a39491a );
 a39498a <=( A200  and  A199 );
 a39501a <=( A203  and  (not A201) );
 a39502a <=( a39501a  and  a39498a );
 a39503a <=( a39502a  and  a39495a );
 a39506a <=( (not A233)  and  A232 );
 a39509a <=( A236  and  (not A235) );
 a39510a <=( a39509a  and  a39506a );
 a39513a <=( (not A299)  and  A298 );
 a39516a <=( A302  and  (not A301) );
 a39517a <=( a39516a  and  a39513a );
 a39518a <=( a39517a  and  a39510a );
 a39521a <=( A168  and  A170 );
 a39524a <=( A166  and  (not A167) );
 a39525a <=( a39524a  and  a39521a );
 a39528a <=( A200  and  A199 );
 a39531a <=( A203  and  (not A201) );
 a39532a <=( a39531a  and  a39528a );
 a39533a <=( a39532a  and  a39525a );
 a39536a <=( (not A233)  and  A232 );
 a39539a <=( A236  and  (not A235) );
 a39540a <=( a39539a  and  a39536a );
 a39543a <=( A299  and  (not A298) );
 a39546a <=( A302  and  (not A301) );
 a39547a <=( a39546a  and  a39543a );
 a39548a <=( a39547a  and  a39540a );
 a39551a <=( A168  and  A170 );
 a39554a <=( A166  and  (not A167) );
 a39555a <=( a39554a  and  a39551a );
 a39558a <=( A200  and  A199 );
 a39561a <=( A203  and  (not A201) );
 a39562a <=( a39561a  and  a39558a );
 a39563a <=( a39562a  and  a39555a );
 a39566a <=( (not A233)  and  A232 );
 a39569a <=( A236  and  (not A235) );
 a39570a <=( a39569a  and  a39566a );
 a39573a <=( (not A299)  and  (not A298) );
 a39576a <=( (not A302)  and  A301 );
 a39577a <=( a39576a  and  a39573a );
 a39578a <=( a39577a  and  a39570a );
 a39581a <=( A168  and  A170 );
 a39584a <=( A166  and  (not A167) );
 a39585a <=( a39584a  and  a39581a );
 a39588a <=( A200  and  A199 );
 a39591a <=( A203  and  (not A201) );
 a39592a <=( a39591a  and  a39588a );
 a39593a <=( a39592a  and  a39585a );
 a39596a <=( (not A233)  and  A232 );
 a39599a <=( A236  and  (not A235) );
 a39600a <=( a39599a  and  a39596a );
 a39603a <=( A266  and  A265 );
 a39606a <=( (not A269)  and  A268 );
 a39607a <=( a39606a  and  a39603a );
 a39608a <=( a39607a  and  a39600a );
 a39611a <=( A168  and  A170 );
 a39614a <=( A166  and  (not A167) );
 a39615a <=( a39614a  and  a39611a );
 a39618a <=( A200  and  A199 );
 a39621a <=( A203  and  (not A201) );
 a39622a <=( a39621a  and  a39618a );
 a39623a <=( a39622a  and  a39615a );
 a39626a <=( (not A233)  and  A232 );
 a39629a <=( A236  and  (not A235) );
 a39630a <=( a39629a  and  a39626a );
 a39633a <=( A266  and  (not A265) );
 a39636a <=( A269  and  (not A268) );
 a39637a <=( a39636a  and  a39633a );
 a39638a <=( a39637a  and  a39630a );
 a39641a <=( A168  and  A170 );
 a39644a <=( A166  and  (not A167) );
 a39645a <=( a39644a  and  a39641a );
 a39648a <=( A200  and  A199 );
 a39651a <=( A203  and  (not A201) );
 a39652a <=( a39651a  and  a39648a );
 a39653a <=( a39652a  and  a39645a );
 a39656a <=( (not A233)  and  A232 );
 a39659a <=( A236  and  (not A235) );
 a39660a <=( a39659a  and  a39656a );
 a39663a <=( (not A266)  and  A265 );
 a39666a <=( A269  and  (not A268) );
 a39667a <=( a39666a  and  a39663a );
 a39668a <=( a39667a  and  a39660a );
 a39671a <=( A168  and  A170 );
 a39674a <=( A166  and  (not A167) );
 a39675a <=( a39674a  and  a39671a );
 a39678a <=( A200  and  A199 );
 a39681a <=( A203  and  (not A201) );
 a39682a <=( a39681a  and  a39678a );
 a39683a <=( a39682a  and  a39675a );
 a39686a <=( (not A233)  and  A232 );
 a39689a <=( A236  and  (not A235) );
 a39690a <=( a39689a  and  a39686a );
 a39693a <=( (not A266)  and  (not A265) );
 a39696a <=( (not A269)  and  A268 );
 a39697a <=( a39696a  and  a39693a );
 a39698a <=( a39697a  and  a39690a );
 a39701a <=( A168  and  A170 );
 a39704a <=( A166  and  (not A167) );
 a39705a <=( a39704a  and  a39701a );
 a39708a <=( A200  and  A199 );
 a39711a <=( A203  and  (not A201) );
 a39712a <=( a39711a  and  a39708a );
 a39713a <=( a39712a  and  a39705a );
 a39716a <=( (not A233)  and  (not A232) );
 a39719a <=( (not A236)  and  A235 );
 a39720a <=( a39719a  and  a39716a );
 a39723a <=( A299  and  A298 );
 a39726a <=( (not A302)  and  A301 );
 a39727a <=( a39726a  and  a39723a );
 a39728a <=( a39727a  and  a39720a );
 a39731a <=( A168  and  A170 );
 a39734a <=( A166  and  (not A167) );
 a39735a <=( a39734a  and  a39731a );
 a39738a <=( A200  and  A199 );
 a39741a <=( A203  and  (not A201) );
 a39742a <=( a39741a  and  a39738a );
 a39743a <=( a39742a  and  a39735a );
 a39746a <=( (not A233)  and  (not A232) );
 a39749a <=( (not A236)  and  A235 );
 a39750a <=( a39749a  and  a39746a );
 a39753a <=( (not A299)  and  A298 );
 a39756a <=( A302  and  (not A301) );
 a39757a <=( a39756a  and  a39753a );
 a39758a <=( a39757a  and  a39750a );
 a39761a <=( A168  and  A170 );
 a39764a <=( A166  and  (not A167) );
 a39765a <=( a39764a  and  a39761a );
 a39768a <=( A200  and  A199 );
 a39771a <=( A203  and  (not A201) );
 a39772a <=( a39771a  and  a39768a );
 a39773a <=( a39772a  and  a39765a );
 a39776a <=( (not A233)  and  (not A232) );
 a39779a <=( (not A236)  and  A235 );
 a39780a <=( a39779a  and  a39776a );
 a39783a <=( A299  and  (not A298) );
 a39786a <=( A302  and  (not A301) );
 a39787a <=( a39786a  and  a39783a );
 a39788a <=( a39787a  and  a39780a );
 a39791a <=( A168  and  A170 );
 a39794a <=( A166  and  (not A167) );
 a39795a <=( a39794a  and  a39791a );
 a39798a <=( A200  and  A199 );
 a39801a <=( A203  and  (not A201) );
 a39802a <=( a39801a  and  a39798a );
 a39803a <=( a39802a  and  a39795a );
 a39806a <=( (not A233)  and  (not A232) );
 a39809a <=( (not A236)  and  A235 );
 a39810a <=( a39809a  and  a39806a );
 a39813a <=( (not A299)  and  (not A298) );
 a39816a <=( (not A302)  and  A301 );
 a39817a <=( a39816a  and  a39813a );
 a39818a <=( a39817a  and  a39810a );
 a39821a <=( A168  and  A170 );
 a39824a <=( A166  and  (not A167) );
 a39825a <=( a39824a  and  a39821a );
 a39828a <=( A200  and  A199 );
 a39831a <=( A203  and  (not A201) );
 a39832a <=( a39831a  and  a39828a );
 a39833a <=( a39832a  and  a39825a );
 a39836a <=( (not A233)  and  (not A232) );
 a39839a <=( (not A236)  and  A235 );
 a39840a <=( a39839a  and  a39836a );
 a39843a <=( A266  and  A265 );
 a39846a <=( (not A269)  and  A268 );
 a39847a <=( a39846a  and  a39843a );
 a39848a <=( a39847a  and  a39840a );
 a39851a <=( A168  and  A170 );
 a39854a <=( A166  and  (not A167) );
 a39855a <=( a39854a  and  a39851a );
 a39858a <=( A200  and  A199 );
 a39861a <=( A203  and  (not A201) );
 a39862a <=( a39861a  and  a39858a );
 a39863a <=( a39862a  and  a39855a );
 a39866a <=( (not A233)  and  (not A232) );
 a39869a <=( (not A236)  and  A235 );
 a39870a <=( a39869a  and  a39866a );
 a39873a <=( A266  and  (not A265) );
 a39876a <=( A269  and  (not A268) );
 a39877a <=( a39876a  and  a39873a );
 a39878a <=( a39877a  and  a39870a );
 a39881a <=( A168  and  A170 );
 a39884a <=( A166  and  (not A167) );
 a39885a <=( a39884a  and  a39881a );
 a39888a <=( A200  and  A199 );
 a39891a <=( A203  and  (not A201) );
 a39892a <=( a39891a  and  a39888a );
 a39893a <=( a39892a  and  a39885a );
 a39896a <=( (not A233)  and  (not A232) );
 a39899a <=( (not A236)  and  A235 );
 a39900a <=( a39899a  and  a39896a );
 a39903a <=( (not A266)  and  A265 );
 a39906a <=( A269  and  (not A268) );
 a39907a <=( a39906a  and  a39903a );
 a39908a <=( a39907a  and  a39900a );
 a39911a <=( A168  and  A170 );
 a39914a <=( A166  and  (not A167) );
 a39915a <=( a39914a  and  a39911a );
 a39918a <=( A200  and  A199 );
 a39921a <=( A203  and  (not A201) );
 a39922a <=( a39921a  and  a39918a );
 a39923a <=( a39922a  and  a39915a );
 a39926a <=( (not A233)  and  (not A232) );
 a39929a <=( (not A236)  and  A235 );
 a39930a <=( a39929a  and  a39926a );
 a39933a <=( (not A266)  and  (not A265) );
 a39936a <=( (not A269)  and  A268 );
 a39937a <=( a39936a  and  a39933a );
 a39938a <=( a39937a  and  a39930a );
 a39941a <=( A168  and  A170 );
 a39944a <=( A166  and  (not A167) );
 a39945a <=( a39944a  and  a39941a );
 a39948a <=( A200  and  (not A199) );
 a39951a <=( A202  and  (not A201) );
 a39952a <=( a39951a  and  a39948a );
 a39953a <=( a39952a  and  a39945a );
 a39956a <=( A233  and  A232 );
 a39959a <=( (not A236)  and  A235 );
 a39960a <=( a39959a  and  a39956a );
 a39963a <=( A299  and  A298 );
 a39966a <=( (not A302)  and  A301 );
 a39967a <=( a39966a  and  a39963a );
 a39968a <=( a39967a  and  a39960a );
 a39971a <=( A168  and  A170 );
 a39974a <=( A166  and  (not A167) );
 a39975a <=( a39974a  and  a39971a );
 a39978a <=( A200  and  (not A199) );
 a39981a <=( A202  and  (not A201) );
 a39982a <=( a39981a  and  a39978a );
 a39983a <=( a39982a  and  a39975a );
 a39986a <=( A233  and  A232 );
 a39989a <=( (not A236)  and  A235 );
 a39990a <=( a39989a  and  a39986a );
 a39993a <=( (not A299)  and  A298 );
 a39996a <=( A302  and  (not A301) );
 a39997a <=( a39996a  and  a39993a );
 a39998a <=( a39997a  and  a39990a );
 a40001a <=( A168  and  A170 );
 a40004a <=( A166  and  (not A167) );
 a40005a <=( a40004a  and  a40001a );
 a40008a <=( A200  and  (not A199) );
 a40011a <=( A202  and  (not A201) );
 a40012a <=( a40011a  and  a40008a );
 a40013a <=( a40012a  and  a40005a );
 a40016a <=( A233  and  A232 );
 a40019a <=( (not A236)  and  A235 );
 a40020a <=( a40019a  and  a40016a );
 a40023a <=( A299  and  (not A298) );
 a40026a <=( A302  and  (not A301) );
 a40027a <=( a40026a  and  a40023a );
 a40028a <=( a40027a  and  a40020a );
 a40031a <=( A168  and  A170 );
 a40034a <=( A166  and  (not A167) );
 a40035a <=( a40034a  and  a40031a );
 a40038a <=( A200  and  (not A199) );
 a40041a <=( A202  and  (not A201) );
 a40042a <=( a40041a  and  a40038a );
 a40043a <=( a40042a  and  a40035a );
 a40046a <=( A233  and  A232 );
 a40049a <=( (not A236)  and  A235 );
 a40050a <=( a40049a  and  a40046a );
 a40053a <=( (not A299)  and  (not A298) );
 a40056a <=( (not A302)  and  A301 );
 a40057a <=( a40056a  and  a40053a );
 a40058a <=( a40057a  and  a40050a );
 a40061a <=( A168  and  A170 );
 a40064a <=( A166  and  (not A167) );
 a40065a <=( a40064a  and  a40061a );
 a40068a <=( A200  and  (not A199) );
 a40071a <=( A202  and  (not A201) );
 a40072a <=( a40071a  and  a40068a );
 a40073a <=( a40072a  and  a40065a );
 a40076a <=( A233  and  A232 );
 a40079a <=( (not A236)  and  A235 );
 a40080a <=( a40079a  and  a40076a );
 a40083a <=( A266  and  A265 );
 a40086a <=( (not A269)  and  A268 );
 a40087a <=( a40086a  and  a40083a );
 a40088a <=( a40087a  and  a40080a );
 a40091a <=( A168  and  A170 );
 a40094a <=( A166  and  (not A167) );
 a40095a <=( a40094a  and  a40091a );
 a40098a <=( A200  and  (not A199) );
 a40101a <=( A202  and  (not A201) );
 a40102a <=( a40101a  and  a40098a );
 a40103a <=( a40102a  and  a40095a );
 a40106a <=( A233  and  A232 );
 a40109a <=( (not A236)  and  A235 );
 a40110a <=( a40109a  and  a40106a );
 a40113a <=( A266  and  (not A265) );
 a40116a <=( A269  and  (not A268) );
 a40117a <=( a40116a  and  a40113a );
 a40118a <=( a40117a  and  a40110a );
 a40121a <=( A168  and  A170 );
 a40124a <=( A166  and  (not A167) );
 a40125a <=( a40124a  and  a40121a );
 a40128a <=( A200  and  (not A199) );
 a40131a <=( A202  and  (not A201) );
 a40132a <=( a40131a  and  a40128a );
 a40133a <=( a40132a  and  a40125a );
 a40136a <=( A233  and  A232 );
 a40139a <=( (not A236)  and  A235 );
 a40140a <=( a40139a  and  a40136a );
 a40143a <=( (not A266)  and  A265 );
 a40146a <=( A269  and  (not A268) );
 a40147a <=( a40146a  and  a40143a );
 a40148a <=( a40147a  and  a40140a );
 a40151a <=( A168  and  A170 );
 a40154a <=( A166  and  (not A167) );
 a40155a <=( a40154a  and  a40151a );
 a40158a <=( A200  and  (not A199) );
 a40161a <=( A202  and  (not A201) );
 a40162a <=( a40161a  and  a40158a );
 a40163a <=( a40162a  and  a40155a );
 a40166a <=( A233  and  A232 );
 a40169a <=( (not A236)  and  A235 );
 a40170a <=( a40169a  and  a40166a );
 a40173a <=( (not A266)  and  (not A265) );
 a40176a <=( (not A269)  and  A268 );
 a40177a <=( a40176a  and  a40173a );
 a40178a <=( a40177a  and  a40170a );
 a40181a <=( A168  and  A170 );
 a40184a <=( A166  and  (not A167) );
 a40185a <=( a40184a  and  a40181a );
 a40188a <=( A200  and  (not A199) );
 a40191a <=( A202  and  (not A201) );
 a40192a <=( a40191a  and  a40188a );
 a40193a <=( a40192a  and  a40185a );
 a40196a <=( A233  and  (not A232) );
 a40199a <=( A236  and  (not A235) );
 a40200a <=( a40199a  and  a40196a );
 a40203a <=( A299  and  A298 );
 a40206a <=( (not A302)  and  A301 );
 a40207a <=( a40206a  and  a40203a );
 a40208a <=( a40207a  and  a40200a );
 a40211a <=( A168  and  A170 );
 a40214a <=( A166  and  (not A167) );
 a40215a <=( a40214a  and  a40211a );
 a40218a <=( A200  and  (not A199) );
 a40221a <=( A202  and  (not A201) );
 a40222a <=( a40221a  and  a40218a );
 a40223a <=( a40222a  and  a40215a );
 a40226a <=( A233  and  (not A232) );
 a40229a <=( A236  and  (not A235) );
 a40230a <=( a40229a  and  a40226a );
 a40233a <=( (not A299)  and  A298 );
 a40236a <=( A302  and  (not A301) );
 a40237a <=( a40236a  and  a40233a );
 a40238a <=( a40237a  and  a40230a );
 a40241a <=( A168  and  A170 );
 a40244a <=( A166  and  (not A167) );
 a40245a <=( a40244a  and  a40241a );
 a40248a <=( A200  and  (not A199) );
 a40251a <=( A202  and  (not A201) );
 a40252a <=( a40251a  and  a40248a );
 a40253a <=( a40252a  and  a40245a );
 a40256a <=( A233  and  (not A232) );
 a40259a <=( A236  and  (not A235) );
 a40260a <=( a40259a  and  a40256a );
 a40263a <=( A299  and  (not A298) );
 a40266a <=( A302  and  (not A301) );
 a40267a <=( a40266a  and  a40263a );
 a40268a <=( a40267a  and  a40260a );
 a40271a <=( A168  and  A170 );
 a40274a <=( A166  and  (not A167) );
 a40275a <=( a40274a  and  a40271a );
 a40278a <=( A200  and  (not A199) );
 a40281a <=( A202  and  (not A201) );
 a40282a <=( a40281a  and  a40278a );
 a40283a <=( a40282a  and  a40275a );
 a40286a <=( A233  and  (not A232) );
 a40289a <=( A236  and  (not A235) );
 a40290a <=( a40289a  and  a40286a );
 a40293a <=( (not A299)  and  (not A298) );
 a40296a <=( (not A302)  and  A301 );
 a40297a <=( a40296a  and  a40293a );
 a40298a <=( a40297a  and  a40290a );
 a40301a <=( A168  and  A170 );
 a40304a <=( A166  and  (not A167) );
 a40305a <=( a40304a  and  a40301a );
 a40308a <=( A200  and  (not A199) );
 a40311a <=( A202  and  (not A201) );
 a40312a <=( a40311a  and  a40308a );
 a40313a <=( a40312a  and  a40305a );
 a40316a <=( A233  and  (not A232) );
 a40319a <=( A236  and  (not A235) );
 a40320a <=( a40319a  and  a40316a );
 a40323a <=( A266  and  A265 );
 a40326a <=( (not A269)  and  A268 );
 a40327a <=( a40326a  and  a40323a );
 a40328a <=( a40327a  and  a40320a );
 a40331a <=( A168  and  A170 );
 a40334a <=( A166  and  (not A167) );
 a40335a <=( a40334a  and  a40331a );
 a40338a <=( A200  and  (not A199) );
 a40341a <=( A202  and  (not A201) );
 a40342a <=( a40341a  and  a40338a );
 a40343a <=( a40342a  and  a40335a );
 a40346a <=( A233  and  (not A232) );
 a40349a <=( A236  and  (not A235) );
 a40350a <=( a40349a  and  a40346a );
 a40353a <=( A266  and  (not A265) );
 a40356a <=( A269  and  (not A268) );
 a40357a <=( a40356a  and  a40353a );
 a40358a <=( a40357a  and  a40350a );
 a40361a <=( A168  and  A170 );
 a40364a <=( A166  and  (not A167) );
 a40365a <=( a40364a  and  a40361a );
 a40368a <=( A200  and  (not A199) );
 a40371a <=( A202  and  (not A201) );
 a40372a <=( a40371a  and  a40368a );
 a40373a <=( a40372a  and  a40365a );
 a40376a <=( A233  and  (not A232) );
 a40379a <=( A236  and  (not A235) );
 a40380a <=( a40379a  and  a40376a );
 a40383a <=( (not A266)  and  A265 );
 a40386a <=( A269  and  (not A268) );
 a40387a <=( a40386a  and  a40383a );
 a40388a <=( a40387a  and  a40380a );
 a40391a <=( A168  and  A170 );
 a40394a <=( A166  and  (not A167) );
 a40395a <=( a40394a  and  a40391a );
 a40398a <=( A200  and  (not A199) );
 a40401a <=( A202  and  (not A201) );
 a40402a <=( a40401a  and  a40398a );
 a40403a <=( a40402a  and  a40395a );
 a40406a <=( A233  and  (not A232) );
 a40409a <=( A236  and  (not A235) );
 a40410a <=( a40409a  and  a40406a );
 a40413a <=( (not A266)  and  (not A265) );
 a40416a <=( (not A269)  and  A268 );
 a40417a <=( a40416a  and  a40413a );
 a40418a <=( a40417a  and  a40410a );
 a40421a <=( A168  and  A170 );
 a40424a <=( A166  and  (not A167) );
 a40425a <=( a40424a  and  a40421a );
 a40428a <=( A200  and  (not A199) );
 a40431a <=( A202  and  (not A201) );
 a40432a <=( a40431a  and  a40428a );
 a40433a <=( a40432a  and  a40425a );
 a40436a <=( (not A233)  and  A232 );
 a40439a <=( A236  and  (not A235) );
 a40440a <=( a40439a  and  a40436a );
 a40443a <=( A299  and  A298 );
 a40446a <=( (not A302)  and  A301 );
 a40447a <=( a40446a  and  a40443a );
 a40448a <=( a40447a  and  a40440a );
 a40451a <=( A168  and  A170 );
 a40454a <=( A166  and  (not A167) );
 a40455a <=( a40454a  and  a40451a );
 a40458a <=( A200  and  (not A199) );
 a40461a <=( A202  and  (not A201) );
 a40462a <=( a40461a  and  a40458a );
 a40463a <=( a40462a  and  a40455a );
 a40466a <=( (not A233)  and  A232 );
 a40469a <=( A236  and  (not A235) );
 a40470a <=( a40469a  and  a40466a );
 a40473a <=( (not A299)  and  A298 );
 a40476a <=( A302  and  (not A301) );
 a40477a <=( a40476a  and  a40473a );
 a40478a <=( a40477a  and  a40470a );
 a40481a <=( A168  and  A170 );
 a40484a <=( A166  and  (not A167) );
 a40485a <=( a40484a  and  a40481a );
 a40488a <=( A200  and  (not A199) );
 a40491a <=( A202  and  (not A201) );
 a40492a <=( a40491a  and  a40488a );
 a40493a <=( a40492a  and  a40485a );
 a40496a <=( (not A233)  and  A232 );
 a40499a <=( A236  and  (not A235) );
 a40500a <=( a40499a  and  a40496a );
 a40503a <=( A299  and  (not A298) );
 a40506a <=( A302  and  (not A301) );
 a40507a <=( a40506a  and  a40503a );
 a40508a <=( a40507a  and  a40500a );
 a40511a <=( A168  and  A170 );
 a40514a <=( A166  and  (not A167) );
 a40515a <=( a40514a  and  a40511a );
 a40518a <=( A200  and  (not A199) );
 a40521a <=( A202  and  (not A201) );
 a40522a <=( a40521a  and  a40518a );
 a40523a <=( a40522a  and  a40515a );
 a40526a <=( (not A233)  and  A232 );
 a40529a <=( A236  and  (not A235) );
 a40530a <=( a40529a  and  a40526a );
 a40533a <=( (not A299)  and  (not A298) );
 a40536a <=( (not A302)  and  A301 );
 a40537a <=( a40536a  and  a40533a );
 a40538a <=( a40537a  and  a40530a );
 a40541a <=( A168  and  A170 );
 a40544a <=( A166  and  (not A167) );
 a40545a <=( a40544a  and  a40541a );
 a40548a <=( A200  and  (not A199) );
 a40551a <=( A202  and  (not A201) );
 a40552a <=( a40551a  and  a40548a );
 a40553a <=( a40552a  and  a40545a );
 a40556a <=( (not A233)  and  A232 );
 a40559a <=( A236  and  (not A235) );
 a40560a <=( a40559a  and  a40556a );
 a40563a <=( A266  and  A265 );
 a40566a <=( (not A269)  and  A268 );
 a40567a <=( a40566a  and  a40563a );
 a40568a <=( a40567a  and  a40560a );
 a40571a <=( A168  and  A170 );
 a40574a <=( A166  and  (not A167) );
 a40575a <=( a40574a  and  a40571a );
 a40578a <=( A200  and  (not A199) );
 a40581a <=( A202  and  (not A201) );
 a40582a <=( a40581a  and  a40578a );
 a40583a <=( a40582a  and  a40575a );
 a40586a <=( (not A233)  and  A232 );
 a40589a <=( A236  and  (not A235) );
 a40590a <=( a40589a  and  a40586a );
 a40593a <=( A266  and  (not A265) );
 a40596a <=( A269  and  (not A268) );
 a40597a <=( a40596a  and  a40593a );
 a40598a <=( a40597a  and  a40590a );
 a40601a <=( A168  and  A170 );
 a40604a <=( A166  and  (not A167) );
 a40605a <=( a40604a  and  a40601a );
 a40608a <=( A200  and  (not A199) );
 a40611a <=( A202  and  (not A201) );
 a40612a <=( a40611a  and  a40608a );
 a40613a <=( a40612a  and  a40605a );
 a40616a <=( (not A233)  and  A232 );
 a40619a <=( A236  and  (not A235) );
 a40620a <=( a40619a  and  a40616a );
 a40623a <=( (not A266)  and  A265 );
 a40626a <=( A269  and  (not A268) );
 a40627a <=( a40626a  and  a40623a );
 a40628a <=( a40627a  and  a40620a );
 a40631a <=( A168  and  A170 );
 a40634a <=( A166  and  (not A167) );
 a40635a <=( a40634a  and  a40631a );
 a40638a <=( A200  and  (not A199) );
 a40641a <=( A202  and  (not A201) );
 a40642a <=( a40641a  and  a40638a );
 a40643a <=( a40642a  and  a40635a );
 a40646a <=( (not A233)  and  A232 );
 a40649a <=( A236  and  (not A235) );
 a40650a <=( a40649a  and  a40646a );
 a40653a <=( (not A266)  and  (not A265) );
 a40656a <=( (not A269)  and  A268 );
 a40657a <=( a40656a  and  a40653a );
 a40658a <=( a40657a  and  a40650a );
 a40661a <=( A168  and  A170 );
 a40664a <=( A166  and  (not A167) );
 a40665a <=( a40664a  and  a40661a );
 a40668a <=( A200  and  (not A199) );
 a40671a <=( A202  and  (not A201) );
 a40672a <=( a40671a  and  a40668a );
 a40673a <=( a40672a  and  a40665a );
 a40676a <=( (not A233)  and  (not A232) );
 a40679a <=( (not A236)  and  A235 );
 a40680a <=( a40679a  and  a40676a );
 a40683a <=( A299  and  A298 );
 a40686a <=( (not A302)  and  A301 );
 a40687a <=( a40686a  and  a40683a );
 a40688a <=( a40687a  and  a40680a );
 a40691a <=( A168  and  A170 );
 a40694a <=( A166  and  (not A167) );
 a40695a <=( a40694a  and  a40691a );
 a40698a <=( A200  and  (not A199) );
 a40701a <=( A202  and  (not A201) );
 a40702a <=( a40701a  and  a40698a );
 a40703a <=( a40702a  and  a40695a );
 a40706a <=( (not A233)  and  (not A232) );
 a40709a <=( (not A236)  and  A235 );
 a40710a <=( a40709a  and  a40706a );
 a40713a <=( (not A299)  and  A298 );
 a40716a <=( A302  and  (not A301) );
 a40717a <=( a40716a  and  a40713a );
 a40718a <=( a40717a  and  a40710a );
 a40721a <=( A168  and  A170 );
 a40724a <=( A166  and  (not A167) );
 a40725a <=( a40724a  and  a40721a );
 a40728a <=( A200  and  (not A199) );
 a40731a <=( A202  and  (not A201) );
 a40732a <=( a40731a  and  a40728a );
 a40733a <=( a40732a  and  a40725a );
 a40736a <=( (not A233)  and  (not A232) );
 a40739a <=( (not A236)  and  A235 );
 a40740a <=( a40739a  and  a40736a );
 a40743a <=( A299  and  (not A298) );
 a40746a <=( A302  and  (not A301) );
 a40747a <=( a40746a  and  a40743a );
 a40748a <=( a40747a  and  a40740a );
 a40751a <=( A168  and  A170 );
 a40754a <=( A166  and  (not A167) );
 a40755a <=( a40754a  and  a40751a );
 a40758a <=( A200  and  (not A199) );
 a40761a <=( A202  and  (not A201) );
 a40762a <=( a40761a  and  a40758a );
 a40763a <=( a40762a  and  a40755a );
 a40766a <=( (not A233)  and  (not A232) );
 a40769a <=( (not A236)  and  A235 );
 a40770a <=( a40769a  and  a40766a );
 a40773a <=( (not A299)  and  (not A298) );
 a40776a <=( (not A302)  and  A301 );
 a40777a <=( a40776a  and  a40773a );
 a40778a <=( a40777a  and  a40770a );
 a40781a <=( A168  and  A170 );
 a40784a <=( A166  and  (not A167) );
 a40785a <=( a40784a  and  a40781a );
 a40788a <=( A200  and  (not A199) );
 a40791a <=( A202  and  (not A201) );
 a40792a <=( a40791a  and  a40788a );
 a40793a <=( a40792a  and  a40785a );
 a40796a <=( (not A233)  and  (not A232) );
 a40799a <=( (not A236)  and  A235 );
 a40800a <=( a40799a  and  a40796a );
 a40803a <=( A266  and  A265 );
 a40806a <=( (not A269)  and  A268 );
 a40807a <=( a40806a  and  a40803a );
 a40808a <=( a40807a  and  a40800a );
 a40811a <=( A168  and  A170 );
 a40814a <=( A166  and  (not A167) );
 a40815a <=( a40814a  and  a40811a );
 a40818a <=( A200  and  (not A199) );
 a40821a <=( A202  and  (not A201) );
 a40822a <=( a40821a  and  a40818a );
 a40823a <=( a40822a  and  a40815a );
 a40826a <=( (not A233)  and  (not A232) );
 a40829a <=( (not A236)  and  A235 );
 a40830a <=( a40829a  and  a40826a );
 a40833a <=( A266  and  (not A265) );
 a40836a <=( A269  and  (not A268) );
 a40837a <=( a40836a  and  a40833a );
 a40838a <=( a40837a  and  a40830a );
 a40841a <=( A168  and  A170 );
 a40844a <=( A166  and  (not A167) );
 a40845a <=( a40844a  and  a40841a );
 a40848a <=( A200  and  (not A199) );
 a40851a <=( A202  and  (not A201) );
 a40852a <=( a40851a  and  a40848a );
 a40853a <=( a40852a  and  a40845a );
 a40856a <=( (not A233)  and  (not A232) );
 a40859a <=( (not A236)  and  A235 );
 a40860a <=( a40859a  and  a40856a );
 a40863a <=( (not A266)  and  A265 );
 a40866a <=( A269  and  (not A268) );
 a40867a <=( a40866a  and  a40863a );
 a40868a <=( a40867a  and  a40860a );
 a40871a <=( A168  and  A170 );
 a40874a <=( A166  and  (not A167) );
 a40875a <=( a40874a  and  a40871a );
 a40878a <=( A200  and  (not A199) );
 a40881a <=( A202  and  (not A201) );
 a40882a <=( a40881a  and  a40878a );
 a40883a <=( a40882a  and  a40875a );
 a40886a <=( (not A233)  and  (not A232) );
 a40889a <=( (not A236)  and  A235 );
 a40890a <=( a40889a  and  a40886a );
 a40893a <=( (not A266)  and  (not A265) );
 a40896a <=( (not A269)  and  A268 );
 a40897a <=( a40896a  and  a40893a );
 a40898a <=( a40897a  and  a40890a );
 a40901a <=( A168  and  A170 );
 a40904a <=( A166  and  (not A167) );
 a40905a <=( a40904a  and  a40901a );
 a40908a <=( A200  and  (not A199) );
 a40911a <=( (not A203)  and  (not A201) );
 a40912a <=( a40911a  and  a40908a );
 a40913a <=( a40912a  and  a40905a );
 a40916a <=( A233  and  A232 );
 a40919a <=( (not A236)  and  A235 );
 a40920a <=( a40919a  and  a40916a );
 a40923a <=( A299  and  A298 );
 a40926a <=( (not A302)  and  A301 );
 a40927a <=( a40926a  and  a40923a );
 a40928a <=( a40927a  and  a40920a );
 a40931a <=( A168  and  A170 );
 a40934a <=( A166  and  (not A167) );
 a40935a <=( a40934a  and  a40931a );
 a40938a <=( A200  and  (not A199) );
 a40941a <=( (not A203)  and  (not A201) );
 a40942a <=( a40941a  and  a40938a );
 a40943a <=( a40942a  and  a40935a );
 a40946a <=( A233  and  A232 );
 a40949a <=( (not A236)  and  A235 );
 a40950a <=( a40949a  and  a40946a );
 a40953a <=( (not A299)  and  A298 );
 a40956a <=( A302  and  (not A301) );
 a40957a <=( a40956a  and  a40953a );
 a40958a <=( a40957a  and  a40950a );
 a40961a <=( A168  and  A170 );
 a40964a <=( A166  and  (not A167) );
 a40965a <=( a40964a  and  a40961a );
 a40968a <=( A200  and  (not A199) );
 a40971a <=( (not A203)  and  (not A201) );
 a40972a <=( a40971a  and  a40968a );
 a40973a <=( a40972a  and  a40965a );
 a40976a <=( A233  and  A232 );
 a40979a <=( (not A236)  and  A235 );
 a40980a <=( a40979a  and  a40976a );
 a40983a <=( A299  and  (not A298) );
 a40986a <=( A302  and  (not A301) );
 a40987a <=( a40986a  and  a40983a );
 a40988a <=( a40987a  and  a40980a );
 a40991a <=( A168  and  A170 );
 a40994a <=( A166  and  (not A167) );
 a40995a <=( a40994a  and  a40991a );
 a40998a <=( A200  and  (not A199) );
 a41001a <=( (not A203)  and  (not A201) );
 a41002a <=( a41001a  and  a40998a );
 a41003a <=( a41002a  and  a40995a );
 a41006a <=( A233  and  A232 );
 a41009a <=( (not A236)  and  A235 );
 a41010a <=( a41009a  and  a41006a );
 a41013a <=( (not A299)  and  (not A298) );
 a41016a <=( (not A302)  and  A301 );
 a41017a <=( a41016a  and  a41013a );
 a41018a <=( a41017a  and  a41010a );
 a41021a <=( A168  and  A170 );
 a41024a <=( A166  and  (not A167) );
 a41025a <=( a41024a  and  a41021a );
 a41028a <=( A200  and  (not A199) );
 a41031a <=( (not A203)  and  (not A201) );
 a41032a <=( a41031a  and  a41028a );
 a41033a <=( a41032a  and  a41025a );
 a41036a <=( A233  and  A232 );
 a41039a <=( (not A236)  and  A235 );
 a41040a <=( a41039a  and  a41036a );
 a41043a <=( A266  and  A265 );
 a41046a <=( (not A269)  and  A268 );
 a41047a <=( a41046a  and  a41043a );
 a41048a <=( a41047a  and  a41040a );
 a41051a <=( A168  and  A170 );
 a41054a <=( A166  and  (not A167) );
 a41055a <=( a41054a  and  a41051a );
 a41058a <=( A200  and  (not A199) );
 a41061a <=( (not A203)  and  (not A201) );
 a41062a <=( a41061a  and  a41058a );
 a41063a <=( a41062a  and  a41055a );
 a41066a <=( A233  and  A232 );
 a41069a <=( (not A236)  and  A235 );
 a41070a <=( a41069a  and  a41066a );
 a41073a <=( A266  and  (not A265) );
 a41076a <=( A269  and  (not A268) );
 a41077a <=( a41076a  and  a41073a );
 a41078a <=( a41077a  and  a41070a );
 a41081a <=( A168  and  A170 );
 a41084a <=( A166  and  (not A167) );
 a41085a <=( a41084a  and  a41081a );
 a41088a <=( A200  and  (not A199) );
 a41091a <=( (not A203)  and  (not A201) );
 a41092a <=( a41091a  and  a41088a );
 a41093a <=( a41092a  and  a41085a );
 a41096a <=( A233  and  A232 );
 a41099a <=( (not A236)  and  A235 );
 a41100a <=( a41099a  and  a41096a );
 a41103a <=( (not A266)  and  A265 );
 a41106a <=( A269  and  (not A268) );
 a41107a <=( a41106a  and  a41103a );
 a41108a <=( a41107a  and  a41100a );
 a41111a <=( A168  and  A170 );
 a41114a <=( A166  and  (not A167) );
 a41115a <=( a41114a  and  a41111a );
 a41118a <=( A200  and  (not A199) );
 a41121a <=( (not A203)  and  (not A201) );
 a41122a <=( a41121a  and  a41118a );
 a41123a <=( a41122a  and  a41115a );
 a41126a <=( A233  and  A232 );
 a41129a <=( (not A236)  and  A235 );
 a41130a <=( a41129a  and  a41126a );
 a41133a <=( (not A266)  and  (not A265) );
 a41136a <=( (not A269)  and  A268 );
 a41137a <=( a41136a  and  a41133a );
 a41138a <=( a41137a  and  a41130a );
 a41141a <=( A168  and  A170 );
 a41144a <=( A166  and  (not A167) );
 a41145a <=( a41144a  and  a41141a );
 a41148a <=( A200  and  (not A199) );
 a41151a <=( (not A203)  and  (not A201) );
 a41152a <=( a41151a  and  a41148a );
 a41153a <=( a41152a  and  a41145a );
 a41156a <=( A233  and  (not A232) );
 a41159a <=( A236  and  (not A235) );
 a41160a <=( a41159a  and  a41156a );
 a41163a <=( A299  and  A298 );
 a41166a <=( (not A302)  and  A301 );
 a41167a <=( a41166a  and  a41163a );
 a41168a <=( a41167a  and  a41160a );
 a41171a <=( A168  and  A170 );
 a41174a <=( A166  and  (not A167) );
 a41175a <=( a41174a  and  a41171a );
 a41178a <=( A200  and  (not A199) );
 a41181a <=( (not A203)  and  (not A201) );
 a41182a <=( a41181a  and  a41178a );
 a41183a <=( a41182a  and  a41175a );
 a41186a <=( A233  and  (not A232) );
 a41189a <=( A236  and  (not A235) );
 a41190a <=( a41189a  and  a41186a );
 a41193a <=( (not A299)  and  A298 );
 a41196a <=( A302  and  (not A301) );
 a41197a <=( a41196a  and  a41193a );
 a41198a <=( a41197a  and  a41190a );
 a41201a <=( A168  and  A170 );
 a41204a <=( A166  and  (not A167) );
 a41205a <=( a41204a  and  a41201a );
 a41208a <=( A200  and  (not A199) );
 a41211a <=( (not A203)  and  (not A201) );
 a41212a <=( a41211a  and  a41208a );
 a41213a <=( a41212a  and  a41205a );
 a41216a <=( A233  and  (not A232) );
 a41219a <=( A236  and  (not A235) );
 a41220a <=( a41219a  and  a41216a );
 a41223a <=( A299  and  (not A298) );
 a41226a <=( A302  and  (not A301) );
 a41227a <=( a41226a  and  a41223a );
 a41228a <=( a41227a  and  a41220a );
 a41231a <=( A168  and  A170 );
 a41234a <=( A166  and  (not A167) );
 a41235a <=( a41234a  and  a41231a );
 a41238a <=( A200  and  (not A199) );
 a41241a <=( (not A203)  and  (not A201) );
 a41242a <=( a41241a  and  a41238a );
 a41243a <=( a41242a  and  a41235a );
 a41246a <=( A233  and  (not A232) );
 a41249a <=( A236  and  (not A235) );
 a41250a <=( a41249a  and  a41246a );
 a41253a <=( (not A299)  and  (not A298) );
 a41256a <=( (not A302)  and  A301 );
 a41257a <=( a41256a  and  a41253a );
 a41258a <=( a41257a  and  a41250a );
 a41261a <=( A168  and  A170 );
 a41264a <=( A166  and  (not A167) );
 a41265a <=( a41264a  and  a41261a );
 a41268a <=( A200  and  (not A199) );
 a41271a <=( (not A203)  and  (not A201) );
 a41272a <=( a41271a  and  a41268a );
 a41273a <=( a41272a  and  a41265a );
 a41276a <=( A233  and  (not A232) );
 a41279a <=( A236  and  (not A235) );
 a41280a <=( a41279a  and  a41276a );
 a41283a <=( A266  and  A265 );
 a41286a <=( (not A269)  and  A268 );
 a41287a <=( a41286a  and  a41283a );
 a41288a <=( a41287a  and  a41280a );
 a41291a <=( A168  and  A170 );
 a41294a <=( A166  and  (not A167) );
 a41295a <=( a41294a  and  a41291a );
 a41298a <=( A200  and  (not A199) );
 a41301a <=( (not A203)  and  (not A201) );
 a41302a <=( a41301a  and  a41298a );
 a41303a <=( a41302a  and  a41295a );
 a41306a <=( A233  and  (not A232) );
 a41309a <=( A236  and  (not A235) );
 a41310a <=( a41309a  and  a41306a );
 a41313a <=( A266  and  (not A265) );
 a41316a <=( A269  and  (not A268) );
 a41317a <=( a41316a  and  a41313a );
 a41318a <=( a41317a  and  a41310a );
 a41321a <=( A168  and  A170 );
 a41324a <=( A166  and  (not A167) );
 a41325a <=( a41324a  and  a41321a );
 a41328a <=( A200  and  (not A199) );
 a41331a <=( (not A203)  and  (not A201) );
 a41332a <=( a41331a  and  a41328a );
 a41333a <=( a41332a  and  a41325a );
 a41336a <=( A233  and  (not A232) );
 a41339a <=( A236  and  (not A235) );
 a41340a <=( a41339a  and  a41336a );
 a41343a <=( (not A266)  and  A265 );
 a41346a <=( A269  and  (not A268) );
 a41347a <=( a41346a  and  a41343a );
 a41348a <=( a41347a  and  a41340a );
 a41351a <=( A168  and  A170 );
 a41354a <=( A166  and  (not A167) );
 a41355a <=( a41354a  and  a41351a );
 a41358a <=( A200  and  (not A199) );
 a41361a <=( (not A203)  and  (not A201) );
 a41362a <=( a41361a  and  a41358a );
 a41363a <=( a41362a  and  a41355a );
 a41366a <=( A233  and  (not A232) );
 a41369a <=( A236  and  (not A235) );
 a41370a <=( a41369a  and  a41366a );
 a41373a <=( (not A266)  and  (not A265) );
 a41376a <=( (not A269)  and  A268 );
 a41377a <=( a41376a  and  a41373a );
 a41378a <=( a41377a  and  a41370a );
 a41381a <=( A168  and  A170 );
 a41384a <=( A166  and  (not A167) );
 a41385a <=( a41384a  and  a41381a );
 a41388a <=( A200  and  (not A199) );
 a41391a <=( (not A203)  and  (not A201) );
 a41392a <=( a41391a  and  a41388a );
 a41393a <=( a41392a  and  a41385a );
 a41396a <=( (not A233)  and  A232 );
 a41399a <=( A236  and  (not A235) );
 a41400a <=( a41399a  and  a41396a );
 a41403a <=( A299  and  A298 );
 a41406a <=( (not A302)  and  A301 );
 a41407a <=( a41406a  and  a41403a );
 a41408a <=( a41407a  and  a41400a );
 a41411a <=( A168  and  A170 );
 a41414a <=( A166  and  (not A167) );
 a41415a <=( a41414a  and  a41411a );
 a41418a <=( A200  and  (not A199) );
 a41421a <=( (not A203)  and  (not A201) );
 a41422a <=( a41421a  and  a41418a );
 a41423a <=( a41422a  and  a41415a );
 a41426a <=( (not A233)  and  A232 );
 a41429a <=( A236  and  (not A235) );
 a41430a <=( a41429a  and  a41426a );
 a41433a <=( (not A299)  and  A298 );
 a41436a <=( A302  and  (not A301) );
 a41437a <=( a41436a  and  a41433a );
 a41438a <=( a41437a  and  a41430a );
 a41441a <=( A168  and  A170 );
 a41444a <=( A166  and  (not A167) );
 a41445a <=( a41444a  and  a41441a );
 a41448a <=( A200  and  (not A199) );
 a41451a <=( (not A203)  and  (not A201) );
 a41452a <=( a41451a  and  a41448a );
 a41453a <=( a41452a  and  a41445a );
 a41456a <=( (not A233)  and  A232 );
 a41459a <=( A236  and  (not A235) );
 a41460a <=( a41459a  and  a41456a );
 a41463a <=( A299  and  (not A298) );
 a41466a <=( A302  and  (not A301) );
 a41467a <=( a41466a  and  a41463a );
 a41468a <=( a41467a  and  a41460a );
 a41471a <=( A168  and  A170 );
 a41474a <=( A166  and  (not A167) );
 a41475a <=( a41474a  and  a41471a );
 a41478a <=( A200  and  (not A199) );
 a41481a <=( (not A203)  and  (not A201) );
 a41482a <=( a41481a  and  a41478a );
 a41483a <=( a41482a  and  a41475a );
 a41486a <=( (not A233)  and  A232 );
 a41489a <=( A236  and  (not A235) );
 a41490a <=( a41489a  and  a41486a );
 a41493a <=( (not A299)  and  (not A298) );
 a41496a <=( (not A302)  and  A301 );
 a41497a <=( a41496a  and  a41493a );
 a41498a <=( a41497a  and  a41490a );
 a41501a <=( A168  and  A170 );
 a41504a <=( A166  and  (not A167) );
 a41505a <=( a41504a  and  a41501a );
 a41508a <=( A200  and  (not A199) );
 a41511a <=( (not A203)  and  (not A201) );
 a41512a <=( a41511a  and  a41508a );
 a41513a <=( a41512a  and  a41505a );
 a41516a <=( (not A233)  and  A232 );
 a41519a <=( A236  and  (not A235) );
 a41520a <=( a41519a  and  a41516a );
 a41523a <=( A266  and  A265 );
 a41526a <=( (not A269)  and  A268 );
 a41527a <=( a41526a  and  a41523a );
 a41528a <=( a41527a  and  a41520a );
 a41531a <=( A168  and  A170 );
 a41534a <=( A166  and  (not A167) );
 a41535a <=( a41534a  and  a41531a );
 a41538a <=( A200  and  (not A199) );
 a41541a <=( (not A203)  and  (not A201) );
 a41542a <=( a41541a  and  a41538a );
 a41543a <=( a41542a  and  a41535a );
 a41546a <=( (not A233)  and  A232 );
 a41549a <=( A236  and  (not A235) );
 a41550a <=( a41549a  and  a41546a );
 a41553a <=( A266  and  (not A265) );
 a41556a <=( A269  and  (not A268) );
 a41557a <=( a41556a  and  a41553a );
 a41558a <=( a41557a  and  a41550a );
 a41561a <=( A168  and  A170 );
 a41564a <=( A166  and  (not A167) );
 a41565a <=( a41564a  and  a41561a );
 a41568a <=( A200  and  (not A199) );
 a41571a <=( (not A203)  and  (not A201) );
 a41572a <=( a41571a  and  a41568a );
 a41573a <=( a41572a  and  a41565a );
 a41576a <=( (not A233)  and  A232 );
 a41579a <=( A236  and  (not A235) );
 a41580a <=( a41579a  and  a41576a );
 a41583a <=( (not A266)  and  A265 );
 a41586a <=( A269  and  (not A268) );
 a41587a <=( a41586a  and  a41583a );
 a41588a <=( a41587a  and  a41580a );
 a41591a <=( A168  and  A170 );
 a41594a <=( A166  and  (not A167) );
 a41595a <=( a41594a  and  a41591a );
 a41598a <=( A200  and  (not A199) );
 a41601a <=( (not A203)  and  (not A201) );
 a41602a <=( a41601a  and  a41598a );
 a41603a <=( a41602a  and  a41595a );
 a41606a <=( (not A233)  and  A232 );
 a41609a <=( A236  and  (not A235) );
 a41610a <=( a41609a  and  a41606a );
 a41613a <=( (not A266)  and  (not A265) );
 a41616a <=( (not A269)  and  A268 );
 a41617a <=( a41616a  and  a41613a );
 a41618a <=( a41617a  and  a41610a );
 a41621a <=( A168  and  A170 );
 a41624a <=( A166  and  (not A167) );
 a41625a <=( a41624a  and  a41621a );
 a41628a <=( A200  and  (not A199) );
 a41631a <=( (not A203)  and  (not A201) );
 a41632a <=( a41631a  and  a41628a );
 a41633a <=( a41632a  and  a41625a );
 a41636a <=( (not A233)  and  (not A232) );
 a41639a <=( (not A236)  and  A235 );
 a41640a <=( a41639a  and  a41636a );
 a41643a <=( A299  and  A298 );
 a41646a <=( (not A302)  and  A301 );
 a41647a <=( a41646a  and  a41643a );
 a41648a <=( a41647a  and  a41640a );
 a41651a <=( A168  and  A170 );
 a41654a <=( A166  and  (not A167) );
 a41655a <=( a41654a  and  a41651a );
 a41658a <=( A200  and  (not A199) );
 a41661a <=( (not A203)  and  (not A201) );
 a41662a <=( a41661a  and  a41658a );
 a41663a <=( a41662a  and  a41655a );
 a41666a <=( (not A233)  and  (not A232) );
 a41669a <=( (not A236)  and  A235 );
 a41670a <=( a41669a  and  a41666a );
 a41673a <=( (not A299)  and  A298 );
 a41676a <=( A302  and  (not A301) );
 a41677a <=( a41676a  and  a41673a );
 a41678a <=( a41677a  and  a41670a );
 a41681a <=( A168  and  A170 );
 a41684a <=( A166  and  (not A167) );
 a41685a <=( a41684a  and  a41681a );
 a41688a <=( A200  and  (not A199) );
 a41691a <=( (not A203)  and  (not A201) );
 a41692a <=( a41691a  and  a41688a );
 a41693a <=( a41692a  and  a41685a );
 a41696a <=( (not A233)  and  (not A232) );
 a41699a <=( (not A236)  and  A235 );
 a41700a <=( a41699a  and  a41696a );
 a41703a <=( A299  and  (not A298) );
 a41706a <=( A302  and  (not A301) );
 a41707a <=( a41706a  and  a41703a );
 a41708a <=( a41707a  and  a41700a );
 a41711a <=( A168  and  A170 );
 a41714a <=( A166  and  (not A167) );
 a41715a <=( a41714a  and  a41711a );
 a41718a <=( A200  and  (not A199) );
 a41721a <=( (not A203)  and  (not A201) );
 a41722a <=( a41721a  and  a41718a );
 a41723a <=( a41722a  and  a41715a );
 a41726a <=( (not A233)  and  (not A232) );
 a41729a <=( (not A236)  and  A235 );
 a41730a <=( a41729a  and  a41726a );
 a41733a <=( (not A299)  and  (not A298) );
 a41736a <=( (not A302)  and  A301 );
 a41737a <=( a41736a  and  a41733a );
 a41738a <=( a41737a  and  a41730a );
 a41741a <=( A168  and  A170 );
 a41744a <=( A166  and  (not A167) );
 a41745a <=( a41744a  and  a41741a );
 a41748a <=( A200  and  (not A199) );
 a41751a <=( (not A203)  and  (not A201) );
 a41752a <=( a41751a  and  a41748a );
 a41753a <=( a41752a  and  a41745a );
 a41756a <=( (not A233)  and  (not A232) );
 a41759a <=( (not A236)  and  A235 );
 a41760a <=( a41759a  and  a41756a );
 a41763a <=( A266  and  A265 );
 a41766a <=( (not A269)  and  A268 );
 a41767a <=( a41766a  and  a41763a );
 a41768a <=( a41767a  and  a41760a );
 a41771a <=( A168  and  A170 );
 a41774a <=( A166  and  (not A167) );
 a41775a <=( a41774a  and  a41771a );
 a41778a <=( A200  and  (not A199) );
 a41781a <=( (not A203)  and  (not A201) );
 a41782a <=( a41781a  and  a41778a );
 a41783a <=( a41782a  and  a41775a );
 a41786a <=( (not A233)  and  (not A232) );
 a41789a <=( (not A236)  and  A235 );
 a41790a <=( a41789a  and  a41786a );
 a41793a <=( A266  and  (not A265) );
 a41796a <=( A269  and  (not A268) );
 a41797a <=( a41796a  and  a41793a );
 a41798a <=( a41797a  and  a41790a );
 a41801a <=( A168  and  A170 );
 a41804a <=( A166  and  (not A167) );
 a41805a <=( a41804a  and  a41801a );
 a41808a <=( A200  and  (not A199) );
 a41811a <=( (not A203)  and  (not A201) );
 a41812a <=( a41811a  and  a41808a );
 a41813a <=( a41812a  and  a41805a );
 a41816a <=( (not A233)  and  (not A232) );
 a41819a <=( (not A236)  and  A235 );
 a41820a <=( a41819a  and  a41816a );
 a41823a <=( (not A266)  and  A265 );
 a41826a <=( A269  and  (not A268) );
 a41827a <=( a41826a  and  a41823a );
 a41828a <=( a41827a  and  a41820a );
 a41831a <=( A168  and  A170 );
 a41834a <=( A166  and  (not A167) );
 a41835a <=( a41834a  and  a41831a );
 a41838a <=( A200  and  (not A199) );
 a41841a <=( (not A203)  and  (not A201) );
 a41842a <=( a41841a  and  a41838a );
 a41843a <=( a41842a  and  a41835a );
 a41846a <=( (not A233)  and  (not A232) );
 a41849a <=( (not A236)  and  A235 );
 a41850a <=( a41849a  and  a41846a );
 a41853a <=( (not A266)  and  (not A265) );
 a41856a <=( (not A269)  and  A268 );
 a41857a <=( a41856a  and  a41853a );
 a41858a <=( a41857a  and  a41850a );
 a41861a <=( A168  and  A170 );
 a41864a <=( A166  and  (not A167) );
 a41865a <=( a41864a  and  a41861a );
 a41868a <=( (not A200)  and  A199 );
 a41871a <=( A202  and  (not A201) );
 a41872a <=( a41871a  and  a41868a );
 a41873a <=( a41872a  and  a41865a );
 a41876a <=( A233  and  A232 );
 a41879a <=( (not A236)  and  A235 );
 a41880a <=( a41879a  and  a41876a );
 a41883a <=( A299  and  A298 );
 a41886a <=( (not A302)  and  A301 );
 a41887a <=( a41886a  and  a41883a );
 a41888a <=( a41887a  and  a41880a );
 a41891a <=( A168  and  A170 );
 a41894a <=( A166  and  (not A167) );
 a41895a <=( a41894a  and  a41891a );
 a41898a <=( (not A200)  and  A199 );
 a41901a <=( A202  and  (not A201) );
 a41902a <=( a41901a  and  a41898a );
 a41903a <=( a41902a  and  a41895a );
 a41906a <=( A233  and  A232 );
 a41909a <=( (not A236)  and  A235 );
 a41910a <=( a41909a  and  a41906a );
 a41913a <=( (not A299)  and  A298 );
 a41916a <=( A302  and  (not A301) );
 a41917a <=( a41916a  and  a41913a );
 a41918a <=( a41917a  and  a41910a );
 a41921a <=( A168  and  A170 );
 a41924a <=( A166  and  (not A167) );
 a41925a <=( a41924a  and  a41921a );
 a41928a <=( (not A200)  and  A199 );
 a41931a <=( A202  and  (not A201) );
 a41932a <=( a41931a  and  a41928a );
 a41933a <=( a41932a  and  a41925a );
 a41936a <=( A233  and  A232 );
 a41939a <=( (not A236)  and  A235 );
 a41940a <=( a41939a  and  a41936a );
 a41943a <=( A299  and  (not A298) );
 a41946a <=( A302  and  (not A301) );
 a41947a <=( a41946a  and  a41943a );
 a41948a <=( a41947a  and  a41940a );
 a41951a <=( A168  and  A170 );
 a41954a <=( A166  and  (not A167) );
 a41955a <=( a41954a  and  a41951a );
 a41958a <=( (not A200)  and  A199 );
 a41961a <=( A202  and  (not A201) );
 a41962a <=( a41961a  and  a41958a );
 a41963a <=( a41962a  and  a41955a );
 a41966a <=( A233  and  A232 );
 a41969a <=( (not A236)  and  A235 );
 a41970a <=( a41969a  and  a41966a );
 a41973a <=( (not A299)  and  (not A298) );
 a41976a <=( (not A302)  and  A301 );
 a41977a <=( a41976a  and  a41973a );
 a41978a <=( a41977a  and  a41970a );
 a41981a <=( A168  and  A170 );
 a41984a <=( A166  and  (not A167) );
 a41985a <=( a41984a  and  a41981a );
 a41988a <=( (not A200)  and  A199 );
 a41991a <=( A202  and  (not A201) );
 a41992a <=( a41991a  and  a41988a );
 a41993a <=( a41992a  and  a41985a );
 a41996a <=( A233  and  A232 );
 a41999a <=( (not A236)  and  A235 );
 a42000a <=( a41999a  and  a41996a );
 a42003a <=( A266  and  A265 );
 a42006a <=( (not A269)  and  A268 );
 a42007a <=( a42006a  and  a42003a );
 a42008a <=( a42007a  and  a42000a );
 a42011a <=( A168  and  A170 );
 a42014a <=( A166  and  (not A167) );
 a42015a <=( a42014a  and  a42011a );
 a42018a <=( (not A200)  and  A199 );
 a42021a <=( A202  and  (not A201) );
 a42022a <=( a42021a  and  a42018a );
 a42023a <=( a42022a  and  a42015a );
 a42026a <=( A233  and  A232 );
 a42029a <=( (not A236)  and  A235 );
 a42030a <=( a42029a  and  a42026a );
 a42033a <=( A266  and  (not A265) );
 a42036a <=( A269  and  (not A268) );
 a42037a <=( a42036a  and  a42033a );
 a42038a <=( a42037a  and  a42030a );
 a42041a <=( A168  and  A170 );
 a42044a <=( A166  and  (not A167) );
 a42045a <=( a42044a  and  a42041a );
 a42048a <=( (not A200)  and  A199 );
 a42051a <=( A202  and  (not A201) );
 a42052a <=( a42051a  and  a42048a );
 a42053a <=( a42052a  and  a42045a );
 a42056a <=( A233  and  A232 );
 a42059a <=( (not A236)  and  A235 );
 a42060a <=( a42059a  and  a42056a );
 a42063a <=( (not A266)  and  A265 );
 a42066a <=( A269  and  (not A268) );
 a42067a <=( a42066a  and  a42063a );
 a42068a <=( a42067a  and  a42060a );
 a42071a <=( A168  and  A170 );
 a42074a <=( A166  and  (not A167) );
 a42075a <=( a42074a  and  a42071a );
 a42078a <=( (not A200)  and  A199 );
 a42081a <=( A202  and  (not A201) );
 a42082a <=( a42081a  and  a42078a );
 a42083a <=( a42082a  and  a42075a );
 a42086a <=( A233  and  A232 );
 a42089a <=( (not A236)  and  A235 );
 a42090a <=( a42089a  and  a42086a );
 a42093a <=( (not A266)  and  (not A265) );
 a42096a <=( (not A269)  and  A268 );
 a42097a <=( a42096a  and  a42093a );
 a42098a <=( a42097a  and  a42090a );
 a42101a <=( A168  and  A170 );
 a42104a <=( A166  and  (not A167) );
 a42105a <=( a42104a  and  a42101a );
 a42108a <=( (not A200)  and  A199 );
 a42111a <=( A202  and  (not A201) );
 a42112a <=( a42111a  and  a42108a );
 a42113a <=( a42112a  and  a42105a );
 a42116a <=( A233  and  (not A232) );
 a42119a <=( A236  and  (not A235) );
 a42120a <=( a42119a  and  a42116a );
 a42123a <=( A299  and  A298 );
 a42126a <=( (not A302)  and  A301 );
 a42127a <=( a42126a  and  a42123a );
 a42128a <=( a42127a  and  a42120a );
 a42131a <=( A168  and  A170 );
 a42134a <=( A166  and  (not A167) );
 a42135a <=( a42134a  and  a42131a );
 a42138a <=( (not A200)  and  A199 );
 a42141a <=( A202  and  (not A201) );
 a42142a <=( a42141a  and  a42138a );
 a42143a <=( a42142a  and  a42135a );
 a42146a <=( A233  and  (not A232) );
 a42149a <=( A236  and  (not A235) );
 a42150a <=( a42149a  and  a42146a );
 a42153a <=( (not A299)  and  A298 );
 a42156a <=( A302  and  (not A301) );
 a42157a <=( a42156a  and  a42153a );
 a42158a <=( a42157a  and  a42150a );
 a42161a <=( A168  and  A170 );
 a42164a <=( A166  and  (not A167) );
 a42165a <=( a42164a  and  a42161a );
 a42168a <=( (not A200)  and  A199 );
 a42171a <=( A202  and  (not A201) );
 a42172a <=( a42171a  and  a42168a );
 a42173a <=( a42172a  and  a42165a );
 a42176a <=( A233  and  (not A232) );
 a42179a <=( A236  and  (not A235) );
 a42180a <=( a42179a  and  a42176a );
 a42183a <=( A299  and  (not A298) );
 a42186a <=( A302  and  (not A301) );
 a42187a <=( a42186a  and  a42183a );
 a42188a <=( a42187a  and  a42180a );
 a42191a <=( A168  and  A170 );
 a42194a <=( A166  and  (not A167) );
 a42195a <=( a42194a  and  a42191a );
 a42198a <=( (not A200)  and  A199 );
 a42201a <=( A202  and  (not A201) );
 a42202a <=( a42201a  and  a42198a );
 a42203a <=( a42202a  and  a42195a );
 a42206a <=( A233  and  (not A232) );
 a42209a <=( A236  and  (not A235) );
 a42210a <=( a42209a  and  a42206a );
 a42213a <=( (not A299)  and  (not A298) );
 a42216a <=( (not A302)  and  A301 );
 a42217a <=( a42216a  and  a42213a );
 a42218a <=( a42217a  and  a42210a );
 a42221a <=( A168  and  A170 );
 a42224a <=( A166  and  (not A167) );
 a42225a <=( a42224a  and  a42221a );
 a42228a <=( (not A200)  and  A199 );
 a42231a <=( A202  and  (not A201) );
 a42232a <=( a42231a  and  a42228a );
 a42233a <=( a42232a  and  a42225a );
 a42236a <=( A233  and  (not A232) );
 a42239a <=( A236  and  (not A235) );
 a42240a <=( a42239a  and  a42236a );
 a42243a <=( A266  and  A265 );
 a42246a <=( (not A269)  and  A268 );
 a42247a <=( a42246a  and  a42243a );
 a42248a <=( a42247a  and  a42240a );
 a42251a <=( A168  and  A170 );
 a42254a <=( A166  and  (not A167) );
 a42255a <=( a42254a  and  a42251a );
 a42258a <=( (not A200)  and  A199 );
 a42261a <=( A202  and  (not A201) );
 a42262a <=( a42261a  and  a42258a );
 a42263a <=( a42262a  and  a42255a );
 a42266a <=( A233  and  (not A232) );
 a42269a <=( A236  and  (not A235) );
 a42270a <=( a42269a  and  a42266a );
 a42273a <=( A266  and  (not A265) );
 a42276a <=( A269  and  (not A268) );
 a42277a <=( a42276a  and  a42273a );
 a42278a <=( a42277a  and  a42270a );
 a42281a <=( A168  and  A170 );
 a42284a <=( A166  and  (not A167) );
 a42285a <=( a42284a  and  a42281a );
 a42288a <=( (not A200)  and  A199 );
 a42291a <=( A202  and  (not A201) );
 a42292a <=( a42291a  and  a42288a );
 a42293a <=( a42292a  and  a42285a );
 a42296a <=( A233  and  (not A232) );
 a42299a <=( A236  and  (not A235) );
 a42300a <=( a42299a  and  a42296a );
 a42303a <=( (not A266)  and  A265 );
 a42306a <=( A269  and  (not A268) );
 a42307a <=( a42306a  and  a42303a );
 a42308a <=( a42307a  and  a42300a );
 a42311a <=( A168  and  A170 );
 a42314a <=( A166  and  (not A167) );
 a42315a <=( a42314a  and  a42311a );
 a42318a <=( (not A200)  and  A199 );
 a42321a <=( A202  and  (not A201) );
 a42322a <=( a42321a  and  a42318a );
 a42323a <=( a42322a  and  a42315a );
 a42326a <=( A233  and  (not A232) );
 a42329a <=( A236  and  (not A235) );
 a42330a <=( a42329a  and  a42326a );
 a42333a <=( (not A266)  and  (not A265) );
 a42336a <=( (not A269)  and  A268 );
 a42337a <=( a42336a  and  a42333a );
 a42338a <=( a42337a  and  a42330a );
 a42341a <=( A168  and  A170 );
 a42344a <=( A166  and  (not A167) );
 a42345a <=( a42344a  and  a42341a );
 a42348a <=( (not A200)  and  A199 );
 a42351a <=( A202  and  (not A201) );
 a42352a <=( a42351a  and  a42348a );
 a42353a <=( a42352a  and  a42345a );
 a42356a <=( (not A233)  and  A232 );
 a42359a <=( A236  and  (not A235) );
 a42360a <=( a42359a  and  a42356a );
 a42363a <=( A299  and  A298 );
 a42366a <=( (not A302)  and  A301 );
 a42367a <=( a42366a  and  a42363a );
 a42368a <=( a42367a  and  a42360a );
 a42371a <=( A168  and  A170 );
 a42374a <=( A166  and  (not A167) );
 a42375a <=( a42374a  and  a42371a );
 a42378a <=( (not A200)  and  A199 );
 a42381a <=( A202  and  (not A201) );
 a42382a <=( a42381a  and  a42378a );
 a42383a <=( a42382a  and  a42375a );
 a42386a <=( (not A233)  and  A232 );
 a42389a <=( A236  and  (not A235) );
 a42390a <=( a42389a  and  a42386a );
 a42393a <=( (not A299)  and  A298 );
 a42396a <=( A302  and  (not A301) );
 a42397a <=( a42396a  and  a42393a );
 a42398a <=( a42397a  and  a42390a );
 a42401a <=( A168  and  A170 );
 a42404a <=( A166  and  (not A167) );
 a42405a <=( a42404a  and  a42401a );
 a42408a <=( (not A200)  and  A199 );
 a42411a <=( A202  and  (not A201) );
 a42412a <=( a42411a  and  a42408a );
 a42413a <=( a42412a  and  a42405a );
 a42416a <=( (not A233)  and  A232 );
 a42419a <=( A236  and  (not A235) );
 a42420a <=( a42419a  and  a42416a );
 a42423a <=( A299  and  (not A298) );
 a42426a <=( A302  and  (not A301) );
 a42427a <=( a42426a  and  a42423a );
 a42428a <=( a42427a  and  a42420a );
 a42431a <=( A168  and  A170 );
 a42434a <=( A166  and  (not A167) );
 a42435a <=( a42434a  and  a42431a );
 a42438a <=( (not A200)  and  A199 );
 a42441a <=( A202  and  (not A201) );
 a42442a <=( a42441a  and  a42438a );
 a42443a <=( a42442a  and  a42435a );
 a42446a <=( (not A233)  and  A232 );
 a42449a <=( A236  and  (not A235) );
 a42450a <=( a42449a  and  a42446a );
 a42453a <=( (not A299)  and  (not A298) );
 a42456a <=( (not A302)  and  A301 );
 a42457a <=( a42456a  and  a42453a );
 a42458a <=( a42457a  and  a42450a );
 a42461a <=( A168  and  A170 );
 a42464a <=( A166  and  (not A167) );
 a42465a <=( a42464a  and  a42461a );
 a42468a <=( (not A200)  and  A199 );
 a42471a <=( A202  and  (not A201) );
 a42472a <=( a42471a  and  a42468a );
 a42473a <=( a42472a  and  a42465a );
 a42476a <=( (not A233)  and  A232 );
 a42479a <=( A236  and  (not A235) );
 a42480a <=( a42479a  and  a42476a );
 a42483a <=( A266  and  A265 );
 a42486a <=( (not A269)  and  A268 );
 a42487a <=( a42486a  and  a42483a );
 a42488a <=( a42487a  and  a42480a );
 a42491a <=( A168  and  A170 );
 a42494a <=( A166  and  (not A167) );
 a42495a <=( a42494a  and  a42491a );
 a42498a <=( (not A200)  and  A199 );
 a42501a <=( A202  and  (not A201) );
 a42502a <=( a42501a  and  a42498a );
 a42503a <=( a42502a  and  a42495a );
 a42506a <=( (not A233)  and  A232 );
 a42509a <=( A236  and  (not A235) );
 a42510a <=( a42509a  and  a42506a );
 a42513a <=( A266  and  (not A265) );
 a42516a <=( A269  and  (not A268) );
 a42517a <=( a42516a  and  a42513a );
 a42518a <=( a42517a  and  a42510a );
 a42521a <=( A168  and  A170 );
 a42524a <=( A166  and  (not A167) );
 a42525a <=( a42524a  and  a42521a );
 a42528a <=( (not A200)  and  A199 );
 a42531a <=( A202  and  (not A201) );
 a42532a <=( a42531a  and  a42528a );
 a42533a <=( a42532a  and  a42525a );
 a42536a <=( (not A233)  and  A232 );
 a42539a <=( A236  and  (not A235) );
 a42540a <=( a42539a  and  a42536a );
 a42543a <=( (not A266)  and  A265 );
 a42546a <=( A269  and  (not A268) );
 a42547a <=( a42546a  and  a42543a );
 a42548a <=( a42547a  and  a42540a );
 a42551a <=( A168  and  A170 );
 a42554a <=( A166  and  (not A167) );
 a42555a <=( a42554a  and  a42551a );
 a42558a <=( (not A200)  and  A199 );
 a42561a <=( A202  and  (not A201) );
 a42562a <=( a42561a  and  a42558a );
 a42563a <=( a42562a  and  a42555a );
 a42566a <=( (not A233)  and  A232 );
 a42569a <=( A236  and  (not A235) );
 a42570a <=( a42569a  and  a42566a );
 a42573a <=( (not A266)  and  (not A265) );
 a42576a <=( (not A269)  and  A268 );
 a42577a <=( a42576a  and  a42573a );
 a42578a <=( a42577a  and  a42570a );
 a42581a <=( A168  and  A170 );
 a42584a <=( A166  and  (not A167) );
 a42585a <=( a42584a  and  a42581a );
 a42588a <=( (not A200)  and  A199 );
 a42591a <=( A202  and  (not A201) );
 a42592a <=( a42591a  and  a42588a );
 a42593a <=( a42592a  and  a42585a );
 a42596a <=( (not A233)  and  (not A232) );
 a42599a <=( (not A236)  and  A235 );
 a42600a <=( a42599a  and  a42596a );
 a42603a <=( A299  and  A298 );
 a42606a <=( (not A302)  and  A301 );
 a42607a <=( a42606a  and  a42603a );
 a42608a <=( a42607a  and  a42600a );
 a42611a <=( A168  and  A170 );
 a42614a <=( A166  and  (not A167) );
 a42615a <=( a42614a  and  a42611a );
 a42618a <=( (not A200)  and  A199 );
 a42621a <=( A202  and  (not A201) );
 a42622a <=( a42621a  and  a42618a );
 a42623a <=( a42622a  and  a42615a );
 a42626a <=( (not A233)  and  (not A232) );
 a42629a <=( (not A236)  and  A235 );
 a42630a <=( a42629a  and  a42626a );
 a42633a <=( (not A299)  and  A298 );
 a42636a <=( A302  and  (not A301) );
 a42637a <=( a42636a  and  a42633a );
 a42638a <=( a42637a  and  a42630a );
 a42641a <=( A168  and  A170 );
 a42644a <=( A166  and  (not A167) );
 a42645a <=( a42644a  and  a42641a );
 a42648a <=( (not A200)  and  A199 );
 a42651a <=( A202  and  (not A201) );
 a42652a <=( a42651a  and  a42648a );
 a42653a <=( a42652a  and  a42645a );
 a42656a <=( (not A233)  and  (not A232) );
 a42659a <=( (not A236)  and  A235 );
 a42660a <=( a42659a  and  a42656a );
 a42663a <=( A299  and  (not A298) );
 a42666a <=( A302  and  (not A301) );
 a42667a <=( a42666a  and  a42663a );
 a42668a <=( a42667a  and  a42660a );
 a42671a <=( A168  and  A170 );
 a42674a <=( A166  and  (not A167) );
 a42675a <=( a42674a  and  a42671a );
 a42678a <=( (not A200)  and  A199 );
 a42681a <=( A202  and  (not A201) );
 a42682a <=( a42681a  and  a42678a );
 a42683a <=( a42682a  and  a42675a );
 a42686a <=( (not A233)  and  (not A232) );
 a42689a <=( (not A236)  and  A235 );
 a42690a <=( a42689a  and  a42686a );
 a42693a <=( (not A299)  and  (not A298) );
 a42696a <=( (not A302)  and  A301 );
 a42697a <=( a42696a  and  a42693a );
 a42698a <=( a42697a  and  a42690a );
 a42701a <=( A168  and  A170 );
 a42704a <=( A166  and  (not A167) );
 a42705a <=( a42704a  and  a42701a );
 a42708a <=( (not A200)  and  A199 );
 a42711a <=( A202  and  (not A201) );
 a42712a <=( a42711a  and  a42708a );
 a42713a <=( a42712a  and  a42705a );
 a42716a <=( (not A233)  and  (not A232) );
 a42719a <=( (not A236)  and  A235 );
 a42720a <=( a42719a  and  a42716a );
 a42723a <=( A266  and  A265 );
 a42726a <=( (not A269)  and  A268 );
 a42727a <=( a42726a  and  a42723a );
 a42728a <=( a42727a  and  a42720a );
 a42731a <=( A168  and  A170 );
 a42734a <=( A166  and  (not A167) );
 a42735a <=( a42734a  and  a42731a );
 a42738a <=( (not A200)  and  A199 );
 a42741a <=( A202  and  (not A201) );
 a42742a <=( a42741a  and  a42738a );
 a42743a <=( a42742a  and  a42735a );
 a42746a <=( (not A233)  and  (not A232) );
 a42749a <=( (not A236)  and  A235 );
 a42750a <=( a42749a  and  a42746a );
 a42753a <=( A266  and  (not A265) );
 a42756a <=( A269  and  (not A268) );
 a42757a <=( a42756a  and  a42753a );
 a42758a <=( a42757a  and  a42750a );
 a42761a <=( A168  and  A170 );
 a42764a <=( A166  and  (not A167) );
 a42765a <=( a42764a  and  a42761a );
 a42768a <=( (not A200)  and  A199 );
 a42771a <=( A202  and  (not A201) );
 a42772a <=( a42771a  and  a42768a );
 a42773a <=( a42772a  and  a42765a );
 a42776a <=( (not A233)  and  (not A232) );
 a42779a <=( (not A236)  and  A235 );
 a42780a <=( a42779a  and  a42776a );
 a42783a <=( (not A266)  and  A265 );
 a42786a <=( A269  and  (not A268) );
 a42787a <=( a42786a  and  a42783a );
 a42788a <=( a42787a  and  a42780a );
 a42791a <=( A168  and  A170 );
 a42794a <=( A166  and  (not A167) );
 a42795a <=( a42794a  and  a42791a );
 a42798a <=( (not A200)  and  A199 );
 a42801a <=( A202  and  (not A201) );
 a42802a <=( a42801a  and  a42798a );
 a42803a <=( a42802a  and  a42795a );
 a42806a <=( (not A233)  and  (not A232) );
 a42809a <=( (not A236)  and  A235 );
 a42810a <=( a42809a  and  a42806a );
 a42813a <=( (not A266)  and  (not A265) );
 a42816a <=( (not A269)  and  A268 );
 a42817a <=( a42816a  and  a42813a );
 a42818a <=( a42817a  and  a42810a );
 a42821a <=( A168  and  A170 );
 a42824a <=( A166  and  (not A167) );
 a42825a <=( a42824a  and  a42821a );
 a42828a <=( (not A200)  and  A199 );
 a42831a <=( (not A203)  and  (not A201) );
 a42832a <=( a42831a  and  a42828a );
 a42833a <=( a42832a  and  a42825a );
 a42836a <=( A233  and  A232 );
 a42839a <=( (not A236)  and  A235 );
 a42840a <=( a42839a  and  a42836a );
 a42843a <=( A299  and  A298 );
 a42846a <=( (not A302)  and  A301 );
 a42847a <=( a42846a  and  a42843a );
 a42848a <=( a42847a  and  a42840a );
 a42851a <=( A168  and  A170 );
 a42854a <=( A166  and  (not A167) );
 a42855a <=( a42854a  and  a42851a );
 a42858a <=( (not A200)  and  A199 );
 a42861a <=( (not A203)  and  (not A201) );
 a42862a <=( a42861a  and  a42858a );
 a42863a <=( a42862a  and  a42855a );
 a42866a <=( A233  and  A232 );
 a42869a <=( (not A236)  and  A235 );
 a42870a <=( a42869a  and  a42866a );
 a42873a <=( (not A299)  and  A298 );
 a42876a <=( A302  and  (not A301) );
 a42877a <=( a42876a  and  a42873a );
 a42878a <=( a42877a  and  a42870a );
 a42881a <=( A168  and  A170 );
 a42884a <=( A166  and  (not A167) );
 a42885a <=( a42884a  and  a42881a );
 a42888a <=( (not A200)  and  A199 );
 a42891a <=( (not A203)  and  (not A201) );
 a42892a <=( a42891a  and  a42888a );
 a42893a <=( a42892a  and  a42885a );
 a42896a <=( A233  and  A232 );
 a42899a <=( (not A236)  and  A235 );
 a42900a <=( a42899a  and  a42896a );
 a42903a <=( A299  and  (not A298) );
 a42906a <=( A302  and  (not A301) );
 a42907a <=( a42906a  and  a42903a );
 a42908a <=( a42907a  and  a42900a );
 a42911a <=( A168  and  A170 );
 a42914a <=( A166  and  (not A167) );
 a42915a <=( a42914a  and  a42911a );
 a42918a <=( (not A200)  and  A199 );
 a42921a <=( (not A203)  and  (not A201) );
 a42922a <=( a42921a  and  a42918a );
 a42923a <=( a42922a  and  a42915a );
 a42926a <=( A233  and  A232 );
 a42929a <=( (not A236)  and  A235 );
 a42930a <=( a42929a  and  a42926a );
 a42933a <=( (not A299)  and  (not A298) );
 a42936a <=( (not A302)  and  A301 );
 a42937a <=( a42936a  and  a42933a );
 a42938a <=( a42937a  and  a42930a );
 a42941a <=( A168  and  A170 );
 a42944a <=( A166  and  (not A167) );
 a42945a <=( a42944a  and  a42941a );
 a42948a <=( (not A200)  and  A199 );
 a42951a <=( (not A203)  and  (not A201) );
 a42952a <=( a42951a  and  a42948a );
 a42953a <=( a42952a  and  a42945a );
 a42956a <=( A233  and  A232 );
 a42959a <=( (not A236)  and  A235 );
 a42960a <=( a42959a  and  a42956a );
 a42963a <=( A266  and  A265 );
 a42966a <=( (not A269)  and  A268 );
 a42967a <=( a42966a  and  a42963a );
 a42968a <=( a42967a  and  a42960a );
 a42971a <=( A168  and  A170 );
 a42974a <=( A166  and  (not A167) );
 a42975a <=( a42974a  and  a42971a );
 a42978a <=( (not A200)  and  A199 );
 a42981a <=( (not A203)  and  (not A201) );
 a42982a <=( a42981a  and  a42978a );
 a42983a <=( a42982a  and  a42975a );
 a42986a <=( A233  and  A232 );
 a42989a <=( (not A236)  and  A235 );
 a42990a <=( a42989a  and  a42986a );
 a42993a <=( A266  and  (not A265) );
 a42996a <=( A269  and  (not A268) );
 a42997a <=( a42996a  and  a42993a );
 a42998a <=( a42997a  and  a42990a );
 a43001a <=( A168  and  A170 );
 a43004a <=( A166  and  (not A167) );
 a43005a <=( a43004a  and  a43001a );
 a43008a <=( (not A200)  and  A199 );
 a43011a <=( (not A203)  and  (not A201) );
 a43012a <=( a43011a  and  a43008a );
 a43013a <=( a43012a  and  a43005a );
 a43016a <=( A233  and  A232 );
 a43019a <=( (not A236)  and  A235 );
 a43020a <=( a43019a  and  a43016a );
 a43023a <=( (not A266)  and  A265 );
 a43026a <=( A269  and  (not A268) );
 a43027a <=( a43026a  and  a43023a );
 a43028a <=( a43027a  and  a43020a );
 a43031a <=( A168  and  A170 );
 a43034a <=( A166  and  (not A167) );
 a43035a <=( a43034a  and  a43031a );
 a43038a <=( (not A200)  and  A199 );
 a43041a <=( (not A203)  and  (not A201) );
 a43042a <=( a43041a  and  a43038a );
 a43043a <=( a43042a  and  a43035a );
 a43046a <=( A233  and  A232 );
 a43049a <=( (not A236)  and  A235 );
 a43050a <=( a43049a  and  a43046a );
 a43053a <=( (not A266)  and  (not A265) );
 a43056a <=( (not A269)  and  A268 );
 a43057a <=( a43056a  and  a43053a );
 a43058a <=( a43057a  and  a43050a );
 a43061a <=( A168  and  A170 );
 a43064a <=( A166  and  (not A167) );
 a43065a <=( a43064a  and  a43061a );
 a43068a <=( (not A200)  and  A199 );
 a43071a <=( (not A203)  and  (not A201) );
 a43072a <=( a43071a  and  a43068a );
 a43073a <=( a43072a  and  a43065a );
 a43076a <=( A233  and  (not A232) );
 a43079a <=( A236  and  (not A235) );
 a43080a <=( a43079a  and  a43076a );
 a43083a <=( A299  and  A298 );
 a43086a <=( (not A302)  and  A301 );
 a43087a <=( a43086a  and  a43083a );
 a43088a <=( a43087a  and  a43080a );
 a43091a <=( A168  and  A170 );
 a43094a <=( A166  and  (not A167) );
 a43095a <=( a43094a  and  a43091a );
 a43098a <=( (not A200)  and  A199 );
 a43101a <=( (not A203)  and  (not A201) );
 a43102a <=( a43101a  and  a43098a );
 a43103a <=( a43102a  and  a43095a );
 a43106a <=( A233  and  (not A232) );
 a43109a <=( A236  and  (not A235) );
 a43110a <=( a43109a  and  a43106a );
 a43113a <=( (not A299)  and  A298 );
 a43116a <=( A302  and  (not A301) );
 a43117a <=( a43116a  and  a43113a );
 a43118a <=( a43117a  and  a43110a );
 a43121a <=( A168  and  A170 );
 a43124a <=( A166  and  (not A167) );
 a43125a <=( a43124a  and  a43121a );
 a43128a <=( (not A200)  and  A199 );
 a43131a <=( (not A203)  and  (not A201) );
 a43132a <=( a43131a  and  a43128a );
 a43133a <=( a43132a  and  a43125a );
 a43136a <=( A233  and  (not A232) );
 a43139a <=( A236  and  (not A235) );
 a43140a <=( a43139a  and  a43136a );
 a43143a <=( A299  and  (not A298) );
 a43146a <=( A302  and  (not A301) );
 a43147a <=( a43146a  and  a43143a );
 a43148a <=( a43147a  and  a43140a );
 a43151a <=( A168  and  A170 );
 a43154a <=( A166  and  (not A167) );
 a43155a <=( a43154a  and  a43151a );
 a43158a <=( (not A200)  and  A199 );
 a43161a <=( (not A203)  and  (not A201) );
 a43162a <=( a43161a  and  a43158a );
 a43163a <=( a43162a  and  a43155a );
 a43166a <=( A233  and  (not A232) );
 a43169a <=( A236  and  (not A235) );
 a43170a <=( a43169a  and  a43166a );
 a43173a <=( (not A299)  and  (not A298) );
 a43176a <=( (not A302)  and  A301 );
 a43177a <=( a43176a  and  a43173a );
 a43178a <=( a43177a  and  a43170a );
 a43181a <=( A168  and  A170 );
 a43184a <=( A166  and  (not A167) );
 a43185a <=( a43184a  and  a43181a );
 a43188a <=( (not A200)  and  A199 );
 a43191a <=( (not A203)  and  (not A201) );
 a43192a <=( a43191a  and  a43188a );
 a43193a <=( a43192a  and  a43185a );
 a43196a <=( A233  and  (not A232) );
 a43199a <=( A236  and  (not A235) );
 a43200a <=( a43199a  and  a43196a );
 a43203a <=( A266  and  A265 );
 a43206a <=( (not A269)  and  A268 );
 a43207a <=( a43206a  and  a43203a );
 a43208a <=( a43207a  and  a43200a );
 a43211a <=( A168  and  A170 );
 a43214a <=( A166  and  (not A167) );
 a43215a <=( a43214a  and  a43211a );
 a43218a <=( (not A200)  and  A199 );
 a43221a <=( (not A203)  and  (not A201) );
 a43222a <=( a43221a  and  a43218a );
 a43223a <=( a43222a  and  a43215a );
 a43226a <=( A233  and  (not A232) );
 a43229a <=( A236  and  (not A235) );
 a43230a <=( a43229a  and  a43226a );
 a43233a <=( A266  and  (not A265) );
 a43236a <=( A269  and  (not A268) );
 a43237a <=( a43236a  and  a43233a );
 a43238a <=( a43237a  and  a43230a );
 a43241a <=( A168  and  A170 );
 a43244a <=( A166  and  (not A167) );
 a43245a <=( a43244a  and  a43241a );
 a43248a <=( (not A200)  and  A199 );
 a43251a <=( (not A203)  and  (not A201) );
 a43252a <=( a43251a  and  a43248a );
 a43253a <=( a43252a  and  a43245a );
 a43256a <=( A233  and  (not A232) );
 a43259a <=( A236  and  (not A235) );
 a43260a <=( a43259a  and  a43256a );
 a43263a <=( (not A266)  and  A265 );
 a43266a <=( A269  and  (not A268) );
 a43267a <=( a43266a  and  a43263a );
 a43268a <=( a43267a  and  a43260a );
 a43271a <=( A168  and  A170 );
 a43274a <=( A166  and  (not A167) );
 a43275a <=( a43274a  and  a43271a );
 a43278a <=( (not A200)  and  A199 );
 a43281a <=( (not A203)  and  (not A201) );
 a43282a <=( a43281a  and  a43278a );
 a43283a <=( a43282a  and  a43275a );
 a43286a <=( A233  and  (not A232) );
 a43289a <=( A236  and  (not A235) );
 a43290a <=( a43289a  and  a43286a );
 a43293a <=( (not A266)  and  (not A265) );
 a43296a <=( (not A269)  and  A268 );
 a43297a <=( a43296a  and  a43293a );
 a43298a <=( a43297a  and  a43290a );
 a43301a <=( A168  and  A170 );
 a43304a <=( A166  and  (not A167) );
 a43305a <=( a43304a  and  a43301a );
 a43308a <=( (not A200)  and  A199 );
 a43311a <=( (not A203)  and  (not A201) );
 a43312a <=( a43311a  and  a43308a );
 a43313a <=( a43312a  and  a43305a );
 a43316a <=( (not A233)  and  A232 );
 a43319a <=( A236  and  (not A235) );
 a43320a <=( a43319a  and  a43316a );
 a43323a <=( A299  and  A298 );
 a43326a <=( (not A302)  and  A301 );
 a43327a <=( a43326a  and  a43323a );
 a43328a <=( a43327a  and  a43320a );
 a43331a <=( A168  and  A170 );
 a43334a <=( A166  and  (not A167) );
 a43335a <=( a43334a  and  a43331a );
 a43338a <=( (not A200)  and  A199 );
 a43341a <=( (not A203)  and  (not A201) );
 a43342a <=( a43341a  and  a43338a );
 a43343a <=( a43342a  and  a43335a );
 a43346a <=( (not A233)  and  A232 );
 a43349a <=( A236  and  (not A235) );
 a43350a <=( a43349a  and  a43346a );
 a43353a <=( (not A299)  and  A298 );
 a43356a <=( A302  and  (not A301) );
 a43357a <=( a43356a  and  a43353a );
 a43358a <=( a43357a  and  a43350a );
 a43361a <=( A168  and  A170 );
 a43364a <=( A166  and  (not A167) );
 a43365a <=( a43364a  and  a43361a );
 a43368a <=( (not A200)  and  A199 );
 a43371a <=( (not A203)  and  (not A201) );
 a43372a <=( a43371a  and  a43368a );
 a43373a <=( a43372a  and  a43365a );
 a43376a <=( (not A233)  and  A232 );
 a43379a <=( A236  and  (not A235) );
 a43380a <=( a43379a  and  a43376a );
 a43383a <=( A299  and  (not A298) );
 a43386a <=( A302  and  (not A301) );
 a43387a <=( a43386a  and  a43383a );
 a43388a <=( a43387a  and  a43380a );
 a43391a <=( A168  and  A170 );
 a43394a <=( A166  and  (not A167) );
 a43395a <=( a43394a  and  a43391a );
 a43398a <=( (not A200)  and  A199 );
 a43401a <=( (not A203)  and  (not A201) );
 a43402a <=( a43401a  and  a43398a );
 a43403a <=( a43402a  and  a43395a );
 a43406a <=( (not A233)  and  A232 );
 a43409a <=( A236  and  (not A235) );
 a43410a <=( a43409a  and  a43406a );
 a43413a <=( (not A299)  and  (not A298) );
 a43416a <=( (not A302)  and  A301 );
 a43417a <=( a43416a  and  a43413a );
 a43418a <=( a43417a  and  a43410a );
 a43421a <=( A168  and  A170 );
 a43424a <=( A166  and  (not A167) );
 a43425a <=( a43424a  and  a43421a );
 a43428a <=( (not A200)  and  A199 );
 a43431a <=( (not A203)  and  (not A201) );
 a43432a <=( a43431a  and  a43428a );
 a43433a <=( a43432a  and  a43425a );
 a43436a <=( (not A233)  and  A232 );
 a43439a <=( A236  and  (not A235) );
 a43440a <=( a43439a  and  a43436a );
 a43443a <=( A266  and  A265 );
 a43446a <=( (not A269)  and  A268 );
 a43447a <=( a43446a  and  a43443a );
 a43448a <=( a43447a  and  a43440a );
 a43451a <=( A168  and  A170 );
 a43454a <=( A166  and  (not A167) );
 a43455a <=( a43454a  and  a43451a );
 a43458a <=( (not A200)  and  A199 );
 a43461a <=( (not A203)  and  (not A201) );
 a43462a <=( a43461a  and  a43458a );
 a43463a <=( a43462a  and  a43455a );
 a43466a <=( (not A233)  and  A232 );
 a43469a <=( A236  and  (not A235) );
 a43470a <=( a43469a  and  a43466a );
 a43473a <=( A266  and  (not A265) );
 a43476a <=( A269  and  (not A268) );
 a43477a <=( a43476a  and  a43473a );
 a43478a <=( a43477a  and  a43470a );
 a43481a <=( A168  and  A170 );
 a43484a <=( A166  and  (not A167) );
 a43485a <=( a43484a  and  a43481a );
 a43488a <=( (not A200)  and  A199 );
 a43491a <=( (not A203)  and  (not A201) );
 a43492a <=( a43491a  and  a43488a );
 a43493a <=( a43492a  and  a43485a );
 a43496a <=( (not A233)  and  A232 );
 a43499a <=( A236  and  (not A235) );
 a43500a <=( a43499a  and  a43496a );
 a43503a <=( (not A266)  and  A265 );
 a43506a <=( A269  and  (not A268) );
 a43507a <=( a43506a  and  a43503a );
 a43508a <=( a43507a  and  a43500a );
 a43511a <=( A168  and  A170 );
 a43514a <=( A166  and  (not A167) );
 a43515a <=( a43514a  and  a43511a );
 a43518a <=( (not A200)  and  A199 );
 a43521a <=( (not A203)  and  (not A201) );
 a43522a <=( a43521a  and  a43518a );
 a43523a <=( a43522a  and  a43515a );
 a43526a <=( (not A233)  and  A232 );
 a43529a <=( A236  and  (not A235) );
 a43530a <=( a43529a  and  a43526a );
 a43533a <=( (not A266)  and  (not A265) );
 a43536a <=( (not A269)  and  A268 );
 a43537a <=( a43536a  and  a43533a );
 a43538a <=( a43537a  and  a43530a );
 a43541a <=( A168  and  A170 );
 a43544a <=( A166  and  (not A167) );
 a43545a <=( a43544a  and  a43541a );
 a43548a <=( (not A200)  and  A199 );
 a43551a <=( (not A203)  and  (not A201) );
 a43552a <=( a43551a  and  a43548a );
 a43553a <=( a43552a  and  a43545a );
 a43556a <=( (not A233)  and  (not A232) );
 a43559a <=( (not A236)  and  A235 );
 a43560a <=( a43559a  and  a43556a );
 a43563a <=( A299  and  A298 );
 a43566a <=( (not A302)  and  A301 );
 a43567a <=( a43566a  and  a43563a );
 a43568a <=( a43567a  and  a43560a );
 a43571a <=( A168  and  A170 );
 a43574a <=( A166  and  (not A167) );
 a43575a <=( a43574a  and  a43571a );
 a43578a <=( (not A200)  and  A199 );
 a43581a <=( (not A203)  and  (not A201) );
 a43582a <=( a43581a  and  a43578a );
 a43583a <=( a43582a  and  a43575a );
 a43586a <=( (not A233)  and  (not A232) );
 a43589a <=( (not A236)  and  A235 );
 a43590a <=( a43589a  and  a43586a );
 a43593a <=( (not A299)  and  A298 );
 a43596a <=( A302  and  (not A301) );
 a43597a <=( a43596a  and  a43593a );
 a43598a <=( a43597a  and  a43590a );
 a43601a <=( A168  and  A170 );
 a43604a <=( A166  and  (not A167) );
 a43605a <=( a43604a  and  a43601a );
 a43608a <=( (not A200)  and  A199 );
 a43611a <=( (not A203)  and  (not A201) );
 a43612a <=( a43611a  and  a43608a );
 a43613a <=( a43612a  and  a43605a );
 a43616a <=( (not A233)  and  (not A232) );
 a43619a <=( (not A236)  and  A235 );
 a43620a <=( a43619a  and  a43616a );
 a43623a <=( A299  and  (not A298) );
 a43626a <=( A302  and  (not A301) );
 a43627a <=( a43626a  and  a43623a );
 a43628a <=( a43627a  and  a43620a );
 a43631a <=( A168  and  A170 );
 a43634a <=( A166  and  (not A167) );
 a43635a <=( a43634a  and  a43631a );
 a43638a <=( (not A200)  and  A199 );
 a43641a <=( (not A203)  and  (not A201) );
 a43642a <=( a43641a  and  a43638a );
 a43643a <=( a43642a  and  a43635a );
 a43646a <=( (not A233)  and  (not A232) );
 a43649a <=( (not A236)  and  A235 );
 a43650a <=( a43649a  and  a43646a );
 a43653a <=( (not A299)  and  (not A298) );
 a43656a <=( (not A302)  and  A301 );
 a43657a <=( a43656a  and  a43653a );
 a43658a <=( a43657a  and  a43650a );
 a43661a <=( A168  and  A170 );
 a43664a <=( A166  and  (not A167) );
 a43665a <=( a43664a  and  a43661a );
 a43668a <=( (not A200)  and  A199 );
 a43671a <=( (not A203)  and  (not A201) );
 a43672a <=( a43671a  and  a43668a );
 a43673a <=( a43672a  and  a43665a );
 a43676a <=( (not A233)  and  (not A232) );
 a43679a <=( (not A236)  and  A235 );
 a43680a <=( a43679a  and  a43676a );
 a43683a <=( A266  and  A265 );
 a43686a <=( (not A269)  and  A268 );
 a43687a <=( a43686a  and  a43683a );
 a43688a <=( a43687a  and  a43680a );
 a43691a <=( A168  and  A170 );
 a43694a <=( A166  and  (not A167) );
 a43695a <=( a43694a  and  a43691a );
 a43698a <=( (not A200)  and  A199 );
 a43701a <=( (not A203)  and  (not A201) );
 a43702a <=( a43701a  and  a43698a );
 a43703a <=( a43702a  and  a43695a );
 a43706a <=( (not A233)  and  (not A232) );
 a43709a <=( (not A236)  and  A235 );
 a43710a <=( a43709a  and  a43706a );
 a43713a <=( A266  and  (not A265) );
 a43716a <=( A269  and  (not A268) );
 a43717a <=( a43716a  and  a43713a );
 a43718a <=( a43717a  and  a43710a );
 a43721a <=( A168  and  A170 );
 a43724a <=( A166  and  (not A167) );
 a43725a <=( a43724a  and  a43721a );
 a43728a <=( (not A200)  and  A199 );
 a43731a <=( (not A203)  and  (not A201) );
 a43732a <=( a43731a  and  a43728a );
 a43733a <=( a43732a  and  a43725a );
 a43736a <=( (not A233)  and  (not A232) );
 a43739a <=( (not A236)  and  A235 );
 a43740a <=( a43739a  and  a43736a );
 a43743a <=( (not A266)  and  A265 );
 a43746a <=( A269  and  (not A268) );
 a43747a <=( a43746a  and  a43743a );
 a43748a <=( a43747a  and  a43740a );
 a43751a <=( A168  and  A170 );
 a43754a <=( A166  and  (not A167) );
 a43755a <=( a43754a  and  a43751a );
 a43758a <=( (not A200)  and  A199 );
 a43761a <=( (not A203)  and  (not A201) );
 a43762a <=( a43761a  and  a43758a );
 a43763a <=( a43762a  and  a43755a );
 a43766a <=( (not A233)  and  (not A232) );
 a43769a <=( (not A236)  and  A235 );
 a43770a <=( a43769a  and  a43766a );
 a43773a <=( (not A266)  and  (not A265) );
 a43776a <=( (not A269)  and  A268 );
 a43777a <=( a43776a  and  a43773a );
 a43778a <=( a43777a  and  a43770a );
 a43781a <=( A168  and  A169 );
 a43784a <=( A166  and  (not A167) );
 a43785a <=( a43784a  and  a43781a );
 a43788a <=( A200  and  A199 );
 a43791a <=( (not A202)  and  (not A201) );
 a43792a <=( a43791a  and  a43788a );
 a43793a <=( a43792a  and  a43785a );
 a43796a <=( A233  and  A232 );
 a43799a <=( (not A236)  and  A235 );
 a43800a <=( a43799a  and  a43796a );
 a43803a <=( A299  and  A298 );
 a43806a <=( (not A302)  and  A301 );
 a43807a <=( a43806a  and  a43803a );
 a43808a <=( a43807a  and  a43800a );
 a43811a <=( A168  and  A169 );
 a43814a <=( A166  and  (not A167) );
 a43815a <=( a43814a  and  a43811a );
 a43818a <=( A200  and  A199 );
 a43821a <=( (not A202)  and  (not A201) );
 a43822a <=( a43821a  and  a43818a );
 a43823a <=( a43822a  and  a43815a );
 a43826a <=( A233  and  A232 );
 a43829a <=( (not A236)  and  A235 );
 a43830a <=( a43829a  and  a43826a );
 a43833a <=( (not A299)  and  A298 );
 a43836a <=( A302  and  (not A301) );
 a43837a <=( a43836a  and  a43833a );
 a43838a <=( a43837a  and  a43830a );
 a43841a <=( A168  and  A169 );
 a43844a <=( A166  and  (not A167) );
 a43845a <=( a43844a  and  a43841a );
 a43848a <=( A200  and  A199 );
 a43851a <=( (not A202)  and  (not A201) );
 a43852a <=( a43851a  and  a43848a );
 a43853a <=( a43852a  and  a43845a );
 a43856a <=( A233  and  A232 );
 a43859a <=( (not A236)  and  A235 );
 a43860a <=( a43859a  and  a43856a );
 a43863a <=( A299  and  (not A298) );
 a43866a <=( A302  and  (not A301) );
 a43867a <=( a43866a  and  a43863a );
 a43868a <=( a43867a  and  a43860a );
 a43871a <=( A168  and  A169 );
 a43874a <=( A166  and  (not A167) );
 a43875a <=( a43874a  and  a43871a );
 a43878a <=( A200  and  A199 );
 a43881a <=( (not A202)  and  (not A201) );
 a43882a <=( a43881a  and  a43878a );
 a43883a <=( a43882a  and  a43875a );
 a43886a <=( A233  and  A232 );
 a43889a <=( (not A236)  and  A235 );
 a43890a <=( a43889a  and  a43886a );
 a43893a <=( (not A299)  and  (not A298) );
 a43896a <=( (not A302)  and  A301 );
 a43897a <=( a43896a  and  a43893a );
 a43898a <=( a43897a  and  a43890a );
 a43901a <=( A168  and  A169 );
 a43904a <=( A166  and  (not A167) );
 a43905a <=( a43904a  and  a43901a );
 a43908a <=( A200  and  A199 );
 a43911a <=( (not A202)  and  (not A201) );
 a43912a <=( a43911a  and  a43908a );
 a43913a <=( a43912a  and  a43905a );
 a43916a <=( A233  and  A232 );
 a43919a <=( (not A236)  and  A235 );
 a43920a <=( a43919a  and  a43916a );
 a43923a <=( A266  and  A265 );
 a43926a <=( (not A269)  and  A268 );
 a43927a <=( a43926a  and  a43923a );
 a43928a <=( a43927a  and  a43920a );
 a43931a <=( A168  and  A169 );
 a43934a <=( A166  and  (not A167) );
 a43935a <=( a43934a  and  a43931a );
 a43938a <=( A200  and  A199 );
 a43941a <=( (not A202)  and  (not A201) );
 a43942a <=( a43941a  and  a43938a );
 a43943a <=( a43942a  and  a43935a );
 a43946a <=( A233  and  A232 );
 a43949a <=( (not A236)  and  A235 );
 a43950a <=( a43949a  and  a43946a );
 a43953a <=( A266  and  (not A265) );
 a43956a <=( A269  and  (not A268) );
 a43957a <=( a43956a  and  a43953a );
 a43958a <=( a43957a  and  a43950a );
 a43961a <=( A168  and  A169 );
 a43964a <=( A166  and  (not A167) );
 a43965a <=( a43964a  and  a43961a );
 a43968a <=( A200  and  A199 );
 a43971a <=( (not A202)  and  (not A201) );
 a43972a <=( a43971a  and  a43968a );
 a43973a <=( a43972a  and  a43965a );
 a43976a <=( A233  and  A232 );
 a43979a <=( (not A236)  and  A235 );
 a43980a <=( a43979a  and  a43976a );
 a43983a <=( (not A266)  and  A265 );
 a43986a <=( A269  and  (not A268) );
 a43987a <=( a43986a  and  a43983a );
 a43988a <=( a43987a  and  a43980a );
 a43991a <=( A168  and  A169 );
 a43994a <=( A166  and  (not A167) );
 a43995a <=( a43994a  and  a43991a );
 a43998a <=( A200  and  A199 );
 a44001a <=( (not A202)  and  (not A201) );
 a44002a <=( a44001a  and  a43998a );
 a44003a <=( a44002a  and  a43995a );
 a44006a <=( A233  and  A232 );
 a44009a <=( (not A236)  and  A235 );
 a44010a <=( a44009a  and  a44006a );
 a44013a <=( (not A266)  and  (not A265) );
 a44016a <=( (not A269)  and  A268 );
 a44017a <=( a44016a  and  a44013a );
 a44018a <=( a44017a  and  a44010a );
 a44021a <=( A168  and  A169 );
 a44024a <=( A166  and  (not A167) );
 a44025a <=( a44024a  and  a44021a );
 a44028a <=( A200  and  A199 );
 a44031a <=( (not A202)  and  (not A201) );
 a44032a <=( a44031a  and  a44028a );
 a44033a <=( a44032a  and  a44025a );
 a44036a <=( A233  and  (not A232) );
 a44039a <=( A236  and  (not A235) );
 a44040a <=( a44039a  and  a44036a );
 a44043a <=( A299  and  A298 );
 a44046a <=( (not A302)  and  A301 );
 a44047a <=( a44046a  and  a44043a );
 a44048a <=( a44047a  and  a44040a );
 a44051a <=( A168  and  A169 );
 a44054a <=( A166  and  (not A167) );
 a44055a <=( a44054a  and  a44051a );
 a44058a <=( A200  and  A199 );
 a44061a <=( (not A202)  and  (not A201) );
 a44062a <=( a44061a  and  a44058a );
 a44063a <=( a44062a  and  a44055a );
 a44066a <=( A233  and  (not A232) );
 a44069a <=( A236  and  (not A235) );
 a44070a <=( a44069a  and  a44066a );
 a44073a <=( (not A299)  and  A298 );
 a44076a <=( A302  and  (not A301) );
 a44077a <=( a44076a  and  a44073a );
 a44078a <=( a44077a  and  a44070a );
 a44081a <=( A168  and  A169 );
 a44084a <=( A166  and  (not A167) );
 a44085a <=( a44084a  and  a44081a );
 a44088a <=( A200  and  A199 );
 a44091a <=( (not A202)  and  (not A201) );
 a44092a <=( a44091a  and  a44088a );
 a44093a <=( a44092a  and  a44085a );
 a44096a <=( A233  and  (not A232) );
 a44099a <=( A236  and  (not A235) );
 a44100a <=( a44099a  and  a44096a );
 a44103a <=( A299  and  (not A298) );
 a44106a <=( A302  and  (not A301) );
 a44107a <=( a44106a  and  a44103a );
 a44108a <=( a44107a  and  a44100a );
 a44111a <=( A168  and  A169 );
 a44114a <=( A166  and  (not A167) );
 a44115a <=( a44114a  and  a44111a );
 a44118a <=( A200  and  A199 );
 a44121a <=( (not A202)  and  (not A201) );
 a44122a <=( a44121a  and  a44118a );
 a44123a <=( a44122a  and  a44115a );
 a44126a <=( A233  and  (not A232) );
 a44129a <=( A236  and  (not A235) );
 a44130a <=( a44129a  and  a44126a );
 a44133a <=( (not A299)  and  (not A298) );
 a44136a <=( (not A302)  and  A301 );
 a44137a <=( a44136a  and  a44133a );
 a44138a <=( a44137a  and  a44130a );
 a44141a <=( A168  and  A169 );
 a44144a <=( A166  and  (not A167) );
 a44145a <=( a44144a  and  a44141a );
 a44148a <=( A200  and  A199 );
 a44151a <=( (not A202)  and  (not A201) );
 a44152a <=( a44151a  and  a44148a );
 a44153a <=( a44152a  and  a44145a );
 a44156a <=( A233  and  (not A232) );
 a44159a <=( A236  and  (not A235) );
 a44160a <=( a44159a  and  a44156a );
 a44163a <=( A266  and  A265 );
 a44166a <=( (not A269)  and  A268 );
 a44167a <=( a44166a  and  a44163a );
 a44168a <=( a44167a  and  a44160a );
 a44171a <=( A168  and  A169 );
 a44174a <=( A166  and  (not A167) );
 a44175a <=( a44174a  and  a44171a );
 a44178a <=( A200  and  A199 );
 a44181a <=( (not A202)  and  (not A201) );
 a44182a <=( a44181a  and  a44178a );
 a44183a <=( a44182a  and  a44175a );
 a44186a <=( A233  and  (not A232) );
 a44189a <=( A236  and  (not A235) );
 a44190a <=( a44189a  and  a44186a );
 a44193a <=( A266  and  (not A265) );
 a44196a <=( A269  and  (not A268) );
 a44197a <=( a44196a  and  a44193a );
 a44198a <=( a44197a  and  a44190a );
 a44201a <=( A168  and  A169 );
 a44204a <=( A166  and  (not A167) );
 a44205a <=( a44204a  and  a44201a );
 a44208a <=( A200  and  A199 );
 a44211a <=( (not A202)  and  (not A201) );
 a44212a <=( a44211a  and  a44208a );
 a44213a <=( a44212a  and  a44205a );
 a44216a <=( A233  and  (not A232) );
 a44219a <=( A236  and  (not A235) );
 a44220a <=( a44219a  and  a44216a );
 a44223a <=( (not A266)  and  A265 );
 a44226a <=( A269  and  (not A268) );
 a44227a <=( a44226a  and  a44223a );
 a44228a <=( a44227a  and  a44220a );
 a44231a <=( A168  and  A169 );
 a44234a <=( A166  and  (not A167) );
 a44235a <=( a44234a  and  a44231a );
 a44238a <=( A200  and  A199 );
 a44241a <=( (not A202)  and  (not A201) );
 a44242a <=( a44241a  and  a44238a );
 a44243a <=( a44242a  and  a44235a );
 a44246a <=( A233  and  (not A232) );
 a44249a <=( A236  and  (not A235) );
 a44250a <=( a44249a  and  a44246a );
 a44253a <=( (not A266)  and  (not A265) );
 a44256a <=( (not A269)  and  A268 );
 a44257a <=( a44256a  and  a44253a );
 a44258a <=( a44257a  and  a44250a );
 a44261a <=( A168  and  A169 );
 a44264a <=( A166  and  (not A167) );
 a44265a <=( a44264a  and  a44261a );
 a44268a <=( A200  and  A199 );
 a44271a <=( (not A202)  and  (not A201) );
 a44272a <=( a44271a  and  a44268a );
 a44273a <=( a44272a  and  a44265a );
 a44276a <=( (not A233)  and  A232 );
 a44279a <=( A236  and  (not A235) );
 a44280a <=( a44279a  and  a44276a );
 a44283a <=( A299  and  A298 );
 a44286a <=( (not A302)  and  A301 );
 a44287a <=( a44286a  and  a44283a );
 a44288a <=( a44287a  and  a44280a );
 a44291a <=( A168  and  A169 );
 a44294a <=( A166  and  (not A167) );
 a44295a <=( a44294a  and  a44291a );
 a44298a <=( A200  and  A199 );
 a44301a <=( (not A202)  and  (not A201) );
 a44302a <=( a44301a  and  a44298a );
 a44303a <=( a44302a  and  a44295a );
 a44306a <=( (not A233)  and  A232 );
 a44309a <=( A236  and  (not A235) );
 a44310a <=( a44309a  and  a44306a );
 a44313a <=( (not A299)  and  A298 );
 a44316a <=( A302  and  (not A301) );
 a44317a <=( a44316a  and  a44313a );
 a44318a <=( a44317a  and  a44310a );
 a44321a <=( A168  and  A169 );
 a44324a <=( A166  and  (not A167) );
 a44325a <=( a44324a  and  a44321a );
 a44328a <=( A200  and  A199 );
 a44331a <=( (not A202)  and  (not A201) );
 a44332a <=( a44331a  and  a44328a );
 a44333a <=( a44332a  and  a44325a );
 a44336a <=( (not A233)  and  A232 );
 a44339a <=( A236  and  (not A235) );
 a44340a <=( a44339a  and  a44336a );
 a44343a <=( A299  and  (not A298) );
 a44346a <=( A302  and  (not A301) );
 a44347a <=( a44346a  and  a44343a );
 a44348a <=( a44347a  and  a44340a );
 a44351a <=( A168  and  A169 );
 a44354a <=( A166  and  (not A167) );
 a44355a <=( a44354a  and  a44351a );
 a44358a <=( A200  and  A199 );
 a44361a <=( (not A202)  and  (not A201) );
 a44362a <=( a44361a  and  a44358a );
 a44363a <=( a44362a  and  a44355a );
 a44366a <=( (not A233)  and  A232 );
 a44369a <=( A236  and  (not A235) );
 a44370a <=( a44369a  and  a44366a );
 a44373a <=( (not A299)  and  (not A298) );
 a44376a <=( (not A302)  and  A301 );
 a44377a <=( a44376a  and  a44373a );
 a44378a <=( a44377a  and  a44370a );
 a44381a <=( A168  and  A169 );
 a44384a <=( A166  and  (not A167) );
 a44385a <=( a44384a  and  a44381a );
 a44388a <=( A200  and  A199 );
 a44391a <=( (not A202)  and  (not A201) );
 a44392a <=( a44391a  and  a44388a );
 a44393a <=( a44392a  and  a44385a );
 a44396a <=( (not A233)  and  A232 );
 a44399a <=( A236  and  (not A235) );
 a44400a <=( a44399a  and  a44396a );
 a44403a <=( A266  and  A265 );
 a44406a <=( (not A269)  and  A268 );
 a44407a <=( a44406a  and  a44403a );
 a44408a <=( a44407a  and  a44400a );
 a44411a <=( A168  and  A169 );
 a44414a <=( A166  and  (not A167) );
 a44415a <=( a44414a  and  a44411a );
 a44418a <=( A200  and  A199 );
 a44421a <=( (not A202)  and  (not A201) );
 a44422a <=( a44421a  and  a44418a );
 a44423a <=( a44422a  and  a44415a );
 a44426a <=( (not A233)  and  A232 );
 a44429a <=( A236  and  (not A235) );
 a44430a <=( a44429a  and  a44426a );
 a44433a <=( A266  and  (not A265) );
 a44436a <=( A269  and  (not A268) );
 a44437a <=( a44436a  and  a44433a );
 a44438a <=( a44437a  and  a44430a );
 a44441a <=( A168  and  A169 );
 a44444a <=( A166  and  (not A167) );
 a44445a <=( a44444a  and  a44441a );
 a44448a <=( A200  and  A199 );
 a44451a <=( (not A202)  and  (not A201) );
 a44452a <=( a44451a  and  a44448a );
 a44453a <=( a44452a  and  a44445a );
 a44456a <=( (not A233)  and  A232 );
 a44459a <=( A236  and  (not A235) );
 a44460a <=( a44459a  and  a44456a );
 a44463a <=( (not A266)  and  A265 );
 a44466a <=( A269  and  (not A268) );
 a44467a <=( a44466a  and  a44463a );
 a44468a <=( a44467a  and  a44460a );
 a44471a <=( A168  and  A169 );
 a44474a <=( A166  and  (not A167) );
 a44475a <=( a44474a  and  a44471a );
 a44478a <=( A200  and  A199 );
 a44481a <=( (not A202)  and  (not A201) );
 a44482a <=( a44481a  and  a44478a );
 a44483a <=( a44482a  and  a44475a );
 a44486a <=( (not A233)  and  A232 );
 a44489a <=( A236  and  (not A235) );
 a44490a <=( a44489a  and  a44486a );
 a44493a <=( (not A266)  and  (not A265) );
 a44496a <=( (not A269)  and  A268 );
 a44497a <=( a44496a  and  a44493a );
 a44498a <=( a44497a  and  a44490a );
 a44501a <=( A168  and  A169 );
 a44504a <=( A166  and  (not A167) );
 a44505a <=( a44504a  and  a44501a );
 a44508a <=( A200  and  A199 );
 a44511a <=( (not A202)  and  (not A201) );
 a44512a <=( a44511a  and  a44508a );
 a44513a <=( a44512a  and  a44505a );
 a44516a <=( (not A233)  and  (not A232) );
 a44519a <=( (not A236)  and  A235 );
 a44520a <=( a44519a  and  a44516a );
 a44523a <=( A299  and  A298 );
 a44526a <=( (not A302)  and  A301 );
 a44527a <=( a44526a  and  a44523a );
 a44528a <=( a44527a  and  a44520a );
 a44531a <=( A168  and  A169 );
 a44534a <=( A166  and  (not A167) );
 a44535a <=( a44534a  and  a44531a );
 a44538a <=( A200  and  A199 );
 a44541a <=( (not A202)  and  (not A201) );
 a44542a <=( a44541a  and  a44538a );
 a44543a <=( a44542a  and  a44535a );
 a44546a <=( (not A233)  and  (not A232) );
 a44549a <=( (not A236)  and  A235 );
 a44550a <=( a44549a  and  a44546a );
 a44553a <=( (not A299)  and  A298 );
 a44556a <=( A302  and  (not A301) );
 a44557a <=( a44556a  and  a44553a );
 a44558a <=( a44557a  and  a44550a );
 a44561a <=( A168  and  A169 );
 a44564a <=( A166  and  (not A167) );
 a44565a <=( a44564a  and  a44561a );
 a44568a <=( A200  and  A199 );
 a44571a <=( (not A202)  and  (not A201) );
 a44572a <=( a44571a  and  a44568a );
 a44573a <=( a44572a  and  a44565a );
 a44576a <=( (not A233)  and  (not A232) );
 a44579a <=( (not A236)  and  A235 );
 a44580a <=( a44579a  and  a44576a );
 a44583a <=( A299  and  (not A298) );
 a44586a <=( A302  and  (not A301) );
 a44587a <=( a44586a  and  a44583a );
 a44588a <=( a44587a  and  a44580a );
 a44591a <=( A168  and  A169 );
 a44594a <=( A166  and  (not A167) );
 a44595a <=( a44594a  and  a44591a );
 a44598a <=( A200  and  A199 );
 a44601a <=( (not A202)  and  (not A201) );
 a44602a <=( a44601a  and  a44598a );
 a44603a <=( a44602a  and  a44595a );
 a44606a <=( (not A233)  and  (not A232) );
 a44609a <=( (not A236)  and  A235 );
 a44610a <=( a44609a  and  a44606a );
 a44613a <=( (not A299)  and  (not A298) );
 a44616a <=( (not A302)  and  A301 );
 a44617a <=( a44616a  and  a44613a );
 a44618a <=( a44617a  and  a44610a );
 a44621a <=( A168  and  A169 );
 a44624a <=( A166  and  (not A167) );
 a44625a <=( a44624a  and  a44621a );
 a44628a <=( A200  and  A199 );
 a44631a <=( (not A202)  and  (not A201) );
 a44632a <=( a44631a  and  a44628a );
 a44633a <=( a44632a  and  a44625a );
 a44636a <=( (not A233)  and  (not A232) );
 a44639a <=( (not A236)  and  A235 );
 a44640a <=( a44639a  and  a44636a );
 a44643a <=( A266  and  A265 );
 a44646a <=( (not A269)  and  A268 );
 a44647a <=( a44646a  and  a44643a );
 a44648a <=( a44647a  and  a44640a );
 a44651a <=( A168  and  A169 );
 a44654a <=( A166  and  (not A167) );
 a44655a <=( a44654a  and  a44651a );
 a44658a <=( A200  and  A199 );
 a44661a <=( (not A202)  and  (not A201) );
 a44662a <=( a44661a  and  a44658a );
 a44663a <=( a44662a  and  a44655a );
 a44666a <=( (not A233)  and  (not A232) );
 a44669a <=( (not A236)  and  A235 );
 a44670a <=( a44669a  and  a44666a );
 a44673a <=( A266  and  (not A265) );
 a44676a <=( A269  and  (not A268) );
 a44677a <=( a44676a  and  a44673a );
 a44678a <=( a44677a  and  a44670a );
 a44681a <=( A168  and  A169 );
 a44684a <=( A166  and  (not A167) );
 a44685a <=( a44684a  and  a44681a );
 a44688a <=( A200  and  A199 );
 a44691a <=( (not A202)  and  (not A201) );
 a44692a <=( a44691a  and  a44688a );
 a44693a <=( a44692a  and  a44685a );
 a44696a <=( (not A233)  and  (not A232) );
 a44699a <=( (not A236)  and  A235 );
 a44700a <=( a44699a  and  a44696a );
 a44703a <=( (not A266)  and  A265 );
 a44706a <=( A269  and  (not A268) );
 a44707a <=( a44706a  and  a44703a );
 a44708a <=( a44707a  and  a44700a );
 a44711a <=( A168  and  A169 );
 a44714a <=( A166  and  (not A167) );
 a44715a <=( a44714a  and  a44711a );
 a44718a <=( A200  and  A199 );
 a44721a <=( (not A202)  and  (not A201) );
 a44722a <=( a44721a  and  a44718a );
 a44723a <=( a44722a  and  a44715a );
 a44726a <=( (not A233)  and  (not A232) );
 a44729a <=( (not A236)  and  A235 );
 a44730a <=( a44729a  and  a44726a );
 a44733a <=( (not A266)  and  (not A265) );
 a44736a <=( (not A269)  and  A268 );
 a44737a <=( a44736a  and  a44733a );
 a44738a <=( a44737a  and  a44730a );
 a44741a <=( A168  and  A169 );
 a44744a <=( A166  and  (not A167) );
 a44745a <=( a44744a  and  a44741a );
 a44748a <=( A200  and  A199 );
 a44751a <=( A203  and  (not A201) );
 a44752a <=( a44751a  and  a44748a );
 a44753a <=( a44752a  and  a44745a );
 a44756a <=( A233  and  A232 );
 a44759a <=( (not A236)  and  A235 );
 a44760a <=( a44759a  and  a44756a );
 a44763a <=( A299  and  A298 );
 a44766a <=( (not A302)  and  A301 );
 a44767a <=( a44766a  and  a44763a );
 a44768a <=( a44767a  and  a44760a );
 a44771a <=( A168  and  A169 );
 a44774a <=( A166  and  (not A167) );
 a44775a <=( a44774a  and  a44771a );
 a44778a <=( A200  and  A199 );
 a44781a <=( A203  and  (not A201) );
 a44782a <=( a44781a  and  a44778a );
 a44783a <=( a44782a  and  a44775a );
 a44786a <=( A233  and  A232 );
 a44789a <=( (not A236)  and  A235 );
 a44790a <=( a44789a  and  a44786a );
 a44793a <=( (not A299)  and  A298 );
 a44796a <=( A302  and  (not A301) );
 a44797a <=( a44796a  and  a44793a );
 a44798a <=( a44797a  and  a44790a );
 a44801a <=( A168  and  A169 );
 a44804a <=( A166  and  (not A167) );
 a44805a <=( a44804a  and  a44801a );
 a44808a <=( A200  and  A199 );
 a44811a <=( A203  and  (not A201) );
 a44812a <=( a44811a  and  a44808a );
 a44813a <=( a44812a  and  a44805a );
 a44816a <=( A233  and  A232 );
 a44819a <=( (not A236)  and  A235 );
 a44820a <=( a44819a  and  a44816a );
 a44823a <=( A299  and  (not A298) );
 a44826a <=( A302  and  (not A301) );
 a44827a <=( a44826a  and  a44823a );
 a44828a <=( a44827a  and  a44820a );
 a44831a <=( A168  and  A169 );
 a44834a <=( A166  and  (not A167) );
 a44835a <=( a44834a  and  a44831a );
 a44838a <=( A200  and  A199 );
 a44841a <=( A203  and  (not A201) );
 a44842a <=( a44841a  and  a44838a );
 a44843a <=( a44842a  and  a44835a );
 a44846a <=( A233  and  A232 );
 a44849a <=( (not A236)  and  A235 );
 a44850a <=( a44849a  and  a44846a );
 a44853a <=( (not A299)  and  (not A298) );
 a44856a <=( (not A302)  and  A301 );
 a44857a <=( a44856a  and  a44853a );
 a44858a <=( a44857a  and  a44850a );
 a44861a <=( A168  and  A169 );
 a44864a <=( A166  and  (not A167) );
 a44865a <=( a44864a  and  a44861a );
 a44868a <=( A200  and  A199 );
 a44871a <=( A203  and  (not A201) );
 a44872a <=( a44871a  and  a44868a );
 a44873a <=( a44872a  and  a44865a );
 a44876a <=( A233  and  A232 );
 a44879a <=( (not A236)  and  A235 );
 a44880a <=( a44879a  and  a44876a );
 a44883a <=( A266  and  A265 );
 a44886a <=( (not A269)  and  A268 );
 a44887a <=( a44886a  and  a44883a );
 a44888a <=( a44887a  and  a44880a );
 a44891a <=( A168  and  A169 );
 a44894a <=( A166  and  (not A167) );
 a44895a <=( a44894a  and  a44891a );
 a44898a <=( A200  and  A199 );
 a44901a <=( A203  and  (not A201) );
 a44902a <=( a44901a  and  a44898a );
 a44903a <=( a44902a  and  a44895a );
 a44906a <=( A233  and  A232 );
 a44909a <=( (not A236)  and  A235 );
 a44910a <=( a44909a  and  a44906a );
 a44913a <=( A266  and  (not A265) );
 a44916a <=( A269  and  (not A268) );
 a44917a <=( a44916a  and  a44913a );
 a44918a <=( a44917a  and  a44910a );
 a44921a <=( A168  and  A169 );
 a44924a <=( A166  and  (not A167) );
 a44925a <=( a44924a  and  a44921a );
 a44928a <=( A200  and  A199 );
 a44931a <=( A203  and  (not A201) );
 a44932a <=( a44931a  and  a44928a );
 a44933a <=( a44932a  and  a44925a );
 a44936a <=( A233  and  A232 );
 a44939a <=( (not A236)  and  A235 );
 a44940a <=( a44939a  and  a44936a );
 a44943a <=( (not A266)  and  A265 );
 a44946a <=( A269  and  (not A268) );
 a44947a <=( a44946a  and  a44943a );
 a44948a <=( a44947a  and  a44940a );
 a44951a <=( A168  and  A169 );
 a44954a <=( A166  and  (not A167) );
 a44955a <=( a44954a  and  a44951a );
 a44958a <=( A200  and  A199 );
 a44961a <=( A203  and  (not A201) );
 a44962a <=( a44961a  and  a44958a );
 a44963a <=( a44962a  and  a44955a );
 a44966a <=( A233  and  A232 );
 a44969a <=( (not A236)  and  A235 );
 a44970a <=( a44969a  and  a44966a );
 a44973a <=( (not A266)  and  (not A265) );
 a44976a <=( (not A269)  and  A268 );
 a44977a <=( a44976a  and  a44973a );
 a44978a <=( a44977a  and  a44970a );
 a44981a <=( A168  and  A169 );
 a44984a <=( A166  and  (not A167) );
 a44985a <=( a44984a  and  a44981a );
 a44988a <=( A200  and  A199 );
 a44991a <=( A203  and  (not A201) );
 a44992a <=( a44991a  and  a44988a );
 a44993a <=( a44992a  and  a44985a );
 a44996a <=( A233  and  (not A232) );
 a44999a <=( A236  and  (not A235) );
 a45000a <=( a44999a  and  a44996a );
 a45003a <=( A299  and  A298 );
 a45006a <=( (not A302)  and  A301 );
 a45007a <=( a45006a  and  a45003a );
 a45008a <=( a45007a  and  a45000a );
 a45011a <=( A168  and  A169 );
 a45014a <=( A166  and  (not A167) );
 a45015a <=( a45014a  and  a45011a );
 a45018a <=( A200  and  A199 );
 a45021a <=( A203  and  (not A201) );
 a45022a <=( a45021a  and  a45018a );
 a45023a <=( a45022a  and  a45015a );
 a45026a <=( A233  and  (not A232) );
 a45029a <=( A236  and  (not A235) );
 a45030a <=( a45029a  and  a45026a );
 a45033a <=( (not A299)  and  A298 );
 a45036a <=( A302  and  (not A301) );
 a45037a <=( a45036a  and  a45033a );
 a45038a <=( a45037a  and  a45030a );
 a45041a <=( A168  and  A169 );
 a45044a <=( A166  and  (not A167) );
 a45045a <=( a45044a  and  a45041a );
 a45048a <=( A200  and  A199 );
 a45051a <=( A203  and  (not A201) );
 a45052a <=( a45051a  and  a45048a );
 a45053a <=( a45052a  and  a45045a );
 a45056a <=( A233  and  (not A232) );
 a45059a <=( A236  and  (not A235) );
 a45060a <=( a45059a  and  a45056a );
 a45063a <=( A299  and  (not A298) );
 a45066a <=( A302  and  (not A301) );
 a45067a <=( a45066a  and  a45063a );
 a45068a <=( a45067a  and  a45060a );
 a45071a <=( A168  and  A169 );
 a45074a <=( A166  and  (not A167) );
 a45075a <=( a45074a  and  a45071a );
 a45078a <=( A200  and  A199 );
 a45081a <=( A203  and  (not A201) );
 a45082a <=( a45081a  and  a45078a );
 a45083a <=( a45082a  and  a45075a );
 a45086a <=( A233  and  (not A232) );
 a45089a <=( A236  and  (not A235) );
 a45090a <=( a45089a  and  a45086a );
 a45093a <=( (not A299)  and  (not A298) );
 a45096a <=( (not A302)  and  A301 );
 a45097a <=( a45096a  and  a45093a );
 a45098a <=( a45097a  and  a45090a );
 a45101a <=( A168  and  A169 );
 a45104a <=( A166  and  (not A167) );
 a45105a <=( a45104a  and  a45101a );
 a45108a <=( A200  and  A199 );
 a45111a <=( A203  and  (not A201) );
 a45112a <=( a45111a  and  a45108a );
 a45113a <=( a45112a  and  a45105a );
 a45116a <=( A233  and  (not A232) );
 a45119a <=( A236  and  (not A235) );
 a45120a <=( a45119a  and  a45116a );
 a45123a <=( A266  and  A265 );
 a45126a <=( (not A269)  and  A268 );
 a45127a <=( a45126a  and  a45123a );
 a45128a <=( a45127a  and  a45120a );
 a45131a <=( A168  and  A169 );
 a45134a <=( A166  and  (not A167) );
 a45135a <=( a45134a  and  a45131a );
 a45138a <=( A200  and  A199 );
 a45141a <=( A203  and  (not A201) );
 a45142a <=( a45141a  and  a45138a );
 a45143a <=( a45142a  and  a45135a );
 a45146a <=( A233  and  (not A232) );
 a45149a <=( A236  and  (not A235) );
 a45150a <=( a45149a  and  a45146a );
 a45153a <=( A266  and  (not A265) );
 a45156a <=( A269  and  (not A268) );
 a45157a <=( a45156a  and  a45153a );
 a45158a <=( a45157a  and  a45150a );
 a45161a <=( A168  and  A169 );
 a45164a <=( A166  and  (not A167) );
 a45165a <=( a45164a  and  a45161a );
 a45168a <=( A200  and  A199 );
 a45171a <=( A203  and  (not A201) );
 a45172a <=( a45171a  and  a45168a );
 a45173a <=( a45172a  and  a45165a );
 a45176a <=( A233  and  (not A232) );
 a45179a <=( A236  and  (not A235) );
 a45180a <=( a45179a  and  a45176a );
 a45183a <=( (not A266)  and  A265 );
 a45186a <=( A269  and  (not A268) );
 a45187a <=( a45186a  and  a45183a );
 a45188a <=( a45187a  and  a45180a );
 a45191a <=( A168  and  A169 );
 a45194a <=( A166  and  (not A167) );
 a45195a <=( a45194a  and  a45191a );
 a45198a <=( A200  and  A199 );
 a45201a <=( A203  and  (not A201) );
 a45202a <=( a45201a  and  a45198a );
 a45203a <=( a45202a  and  a45195a );
 a45206a <=( A233  and  (not A232) );
 a45209a <=( A236  and  (not A235) );
 a45210a <=( a45209a  and  a45206a );
 a45213a <=( (not A266)  and  (not A265) );
 a45216a <=( (not A269)  and  A268 );
 a45217a <=( a45216a  and  a45213a );
 a45218a <=( a45217a  and  a45210a );
 a45221a <=( A168  and  A169 );
 a45224a <=( A166  and  (not A167) );
 a45225a <=( a45224a  and  a45221a );
 a45228a <=( A200  and  A199 );
 a45231a <=( A203  and  (not A201) );
 a45232a <=( a45231a  and  a45228a );
 a45233a <=( a45232a  and  a45225a );
 a45236a <=( (not A233)  and  A232 );
 a45239a <=( A236  and  (not A235) );
 a45240a <=( a45239a  and  a45236a );
 a45243a <=( A299  and  A298 );
 a45246a <=( (not A302)  and  A301 );
 a45247a <=( a45246a  and  a45243a );
 a45248a <=( a45247a  and  a45240a );
 a45251a <=( A168  and  A169 );
 a45254a <=( A166  and  (not A167) );
 a45255a <=( a45254a  and  a45251a );
 a45258a <=( A200  and  A199 );
 a45261a <=( A203  and  (not A201) );
 a45262a <=( a45261a  and  a45258a );
 a45263a <=( a45262a  and  a45255a );
 a45266a <=( (not A233)  and  A232 );
 a45269a <=( A236  and  (not A235) );
 a45270a <=( a45269a  and  a45266a );
 a45273a <=( (not A299)  and  A298 );
 a45276a <=( A302  and  (not A301) );
 a45277a <=( a45276a  and  a45273a );
 a45278a <=( a45277a  and  a45270a );
 a45281a <=( A168  and  A169 );
 a45284a <=( A166  and  (not A167) );
 a45285a <=( a45284a  and  a45281a );
 a45288a <=( A200  and  A199 );
 a45291a <=( A203  and  (not A201) );
 a45292a <=( a45291a  and  a45288a );
 a45293a <=( a45292a  and  a45285a );
 a45296a <=( (not A233)  and  A232 );
 a45299a <=( A236  and  (not A235) );
 a45300a <=( a45299a  and  a45296a );
 a45303a <=( A299  and  (not A298) );
 a45306a <=( A302  and  (not A301) );
 a45307a <=( a45306a  and  a45303a );
 a45308a <=( a45307a  and  a45300a );
 a45311a <=( A168  and  A169 );
 a45314a <=( A166  and  (not A167) );
 a45315a <=( a45314a  and  a45311a );
 a45318a <=( A200  and  A199 );
 a45321a <=( A203  and  (not A201) );
 a45322a <=( a45321a  and  a45318a );
 a45323a <=( a45322a  and  a45315a );
 a45326a <=( (not A233)  and  A232 );
 a45329a <=( A236  and  (not A235) );
 a45330a <=( a45329a  and  a45326a );
 a45333a <=( (not A299)  and  (not A298) );
 a45336a <=( (not A302)  and  A301 );
 a45337a <=( a45336a  and  a45333a );
 a45338a <=( a45337a  and  a45330a );
 a45341a <=( A168  and  A169 );
 a45344a <=( A166  and  (not A167) );
 a45345a <=( a45344a  and  a45341a );
 a45348a <=( A200  and  A199 );
 a45351a <=( A203  and  (not A201) );
 a45352a <=( a45351a  and  a45348a );
 a45353a <=( a45352a  and  a45345a );
 a45356a <=( (not A233)  and  A232 );
 a45359a <=( A236  and  (not A235) );
 a45360a <=( a45359a  and  a45356a );
 a45363a <=( A266  and  A265 );
 a45366a <=( (not A269)  and  A268 );
 a45367a <=( a45366a  and  a45363a );
 a45368a <=( a45367a  and  a45360a );
 a45371a <=( A168  and  A169 );
 a45374a <=( A166  and  (not A167) );
 a45375a <=( a45374a  and  a45371a );
 a45378a <=( A200  and  A199 );
 a45381a <=( A203  and  (not A201) );
 a45382a <=( a45381a  and  a45378a );
 a45383a <=( a45382a  and  a45375a );
 a45386a <=( (not A233)  and  A232 );
 a45389a <=( A236  and  (not A235) );
 a45390a <=( a45389a  and  a45386a );
 a45393a <=( A266  and  (not A265) );
 a45396a <=( A269  and  (not A268) );
 a45397a <=( a45396a  and  a45393a );
 a45398a <=( a45397a  and  a45390a );
 a45401a <=( A168  and  A169 );
 a45404a <=( A166  and  (not A167) );
 a45405a <=( a45404a  and  a45401a );
 a45408a <=( A200  and  A199 );
 a45411a <=( A203  and  (not A201) );
 a45412a <=( a45411a  and  a45408a );
 a45413a <=( a45412a  and  a45405a );
 a45416a <=( (not A233)  and  A232 );
 a45419a <=( A236  and  (not A235) );
 a45420a <=( a45419a  and  a45416a );
 a45423a <=( (not A266)  and  A265 );
 a45426a <=( A269  and  (not A268) );
 a45427a <=( a45426a  and  a45423a );
 a45428a <=( a45427a  and  a45420a );
 a45431a <=( A168  and  A169 );
 a45434a <=( A166  and  (not A167) );
 a45435a <=( a45434a  and  a45431a );
 a45438a <=( A200  and  A199 );
 a45441a <=( A203  and  (not A201) );
 a45442a <=( a45441a  and  a45438a );
 a45443a <=( a45442a  and  a45435a );
 a45446a <=( (not A233)  and  A232 );
 a45449a <=( A236  and  (not A235) );
 a45450a <=( a45449a  and  a45446a );
 a45453a <=( (not A266)  and  (not A265) );
 a45456a <=( (not A269)  and  A268 );
 a45457a <=( a45456a  and  a45453a );
 a45458a <=( a45457a  and  a45450a );
 a45461a <=( A168  and  A169 );
 a45464a <=( A166  and  (not A167) );
 a45465a <=( a45464a  and  a45461a );
 a45468a <=( A200  and  A199 );
 a45471a <=( A203  and  (not A201) );
 a45472a <=( a45471a  and  a45468a );
 a45473a <=( a45472a  and  a45465a );
 a45476a <=( (not A233)  and  (not A232) );
 a45479a <=( (not A236)  and  A235 );
 a45480a <=( a45479a  and  a45476a );
 a45483a <=( A299  and  A298 );
 a45486a <=( (not A302)  and  A301 );
 a45487a <=( a45486a  and  a45483a );
 a45488a <=( a45487a  and  a45480a );
 a45491a <=( A168  and  A169 );
 a45494a <=( A166  and  (not A167) );
 a45495a <=( a45494a  and  a45491a );
 a45498a <=( A200  and  A199 );
 a45501a <=( A203  and  (not A201) );
 a45502a <=( a45501a  and  a45498a );
 a45503a <=( a45502a  and  a45495a );
 a45506a <=( (not A233)  and  (not A232) );
 a45509a <=( (not A236)  and  A235 );
 a45510a <=( a45509a  and  a45506a );
 a45513a <=( (not A299)  and  A298 );
 a45516a <=( A302  and  (not A301) );
 a45517a <=( a45516a  and  a45513a );
 a45518a <=( a45517a  and  a45510a );
 a45521a <=( A168  and  A169 );
 a45524a <=( A166  and  (not A167) );
 a45525a <=( a45524a  and  a45521a );
 a45528a <=( A200  and  A199 );
 a45531a <=( A203  and  (not A201) );
 a45532a <=( a45531a  and  a45528a );
 a45533a <=( a45532a  and  a45525a );
 a45536a <=( (not A233)  and  (not A232) );
 a45539a <=( (not A236)  and  A235 );
 a45540a <=( a45539a  and  a45536a );
 a45543a <=( A299  and  (not A298) );
 a45546a <=( A302  and  (not A301) );
 a45547a <=( a45546a  and  a45543a );
 a45548a <=( a45547a  and  a45540a );
 a45551a <=( A168  and  A169 );
 a45554a <=( A166  and  (not A167) );
 a45555a <=( a45554a  and  a45551a );
 a45558a <=( A200  and  A199 );
 a45561a <=( A203  and  (not A201) );
 a45562a <=( a45561a  and  a45558a );
 a45563a <=( a45562a  and  a45555a );
 a45566a <=( (not A233)  and  (not A232) );
 a45569a <=( (not A236)  and  A235 );
 a45570a <=( a45569a  and  a45566a );
 a45573a <=( (not A299)  and  (not A298) );
 a45576a <=( (not A302)  and  A301 );
 a45577a <=( a45576a  and  a45573a );
 a45578a <=( a45577a  and  a45570a );
 a45581a <=( A168  and  A169 );
 a45584a <=( A166  and  (not A167) );
 a45585a <=( a45584a  and  a45581a );
 a45588a <=( A200  and  A199 );
 a45591a <=( A203  and  (not A201) );
 a45592a <=( a45591a  and  a45588a );
 a45593a <=( a45592a  and  a45585a );
 a45596a <=( (not A233)  and  (not A232) );
 a45599a <=( (not A236)  and  A235 );
 a45600a <=( a45599a  and  a45596a );
 a45603a <=( A266  and  A265 );
 a45606a <=( (not A269)  and  A268 );
 a45607a <=( a45606a  and  a45603a );
 a45608a <=( a45607a  and  a45600a );
 a45611a <=( A168  and  A169 );
 a45614a <=( A166  and  (not A167) );
 a45615a <=( a45614a  and  a45611a );
 a45618a <=( A200  and  A199 );
 a45621a <=( A203  and  (not A201) );
 a45622a <=( a45621a  and  a45618a );
 a45623a <=( a45622a  and  a45615a );
 a45626a <=( (not A233)  and  (not A232) );
 a45629a <=( (not A236)  and  A235 );
 a45630a <=( a45629a  and  a45626a );
 a45633a <=( A266  and  (not A265) );
 a45636a <=( A269  and  (not A268) );
 a45637a <=( a45636a  and  a45633a );
 a45638a <=( a45637a  and  a45630a );
 a45641a <=( A168  and  A169 );
 a45644a <=( A166  and  (not A167) );
 a45645a <=( a45644a  and  a45641a );
 a45648a <=( A200  and  A199 );
 a45651a <=( A203  and  (not A201) );
 a45652a <=( a45651a  and  a45648a );
 a45653a <=( a45652a  and  a45645a );
 a45656a <=( (not A233)  and  (not A232) );
 a45659a <=( (not A236)  and  A235 );
 a45660a <=( a45659a  and  a45656a );
 a45663a <=( (not A266)  and  A265 );
 a45666a <=( A269  and  (not A268) );
 a45667a <=( a45666a  and  a45663a );
 a45668a <=( a45667a  and  a45660a );
 a45671a <=( A168  and  A169 );
 a45674a <=( A166  and  (not A167) );
 a45675a <=( a45674a  and  a45671a );
 a45678a <=( A200  and  A199 );
 a45681a <=( A203  and  (not A201) );
 a45682a <=( a45681a  and  a45678a );
 a45683a <=( a45682a  and  a45675a );
 a45686a <=( (not A233)  and  (not A232) );
 a45689a <=( (not A236)  and  A235 );
 a45690a <=( a45689a  and  a45686a );
 a45693a <=( (not A266)  and  (not A265) );
 a45696a <=( (not A269)  and  A268 );
 a45697a <=( a45696a  and  a45693a );
 a45698a <=( a45697a  and  a45690a );
 a45701a <=( A168  and  A169 );
 a45704a <=( A166  and  (not A167) );
 a45705a <=( a45704a  and  a45701a );
 a45708a <=( A200  and  (not A199) );
 a45711a <=( A202  and  (not A201) );
 a45712a <=( a45711a  and  a45708a );
 a45713a <=( a45712a  and  a45705a );
 a45716a <=( A233  and  A232 );
 a45719a <=( (not A236)  and  A235 );
 a45720a <=( a45719a  and  a45716a );
 a45723a <=( A299  and  A298 );
 a45726a <=( (not A302)  and  A301 );
 a45727a <=( a45726a  and  a45723a );
 a45728a <=( a45727a  and  a45720a );
 a45731a <=( A168  and  A169 );
 a45734a <=( A166  and  (not A167) );
 a45735a <=( a45734a  and  a45731a );
 a45738a <=( A200  and  (not A199) );
 a45741a <=( A202  and  (not A201) );
 a45742a <=( a45741a  and  a45738a );
 a45743a <=( a45742a  and  a45735a );
 a45746a <=( A233  and  A232 );
 a45749a <=( (not A236)  and  A235 );
 a45750a <=( a45749a  and  a45746a );
 a45753a <=( (not A299)  and  A298 );
 a45756a <=( A302  and  (not A301) );
 a45757a <=( a45756a  and  a45753a );
 a45758a <=( a45757a  and  a45750a );
 a45761a <=( A168  and  A169 );
 a45764a <=( A166  and  (not A167) );
 a45765a <=( a45764a  and  a45761a );
 a45768a <=( A200  and  (not A199) );
 a45771a <=( A202  and  (not A201) );
 a45772a <=( a45771a  and  a45768a );
 a45773a <=( a45772a  and  a45765a );
 a45776a <=( A233  and  A232 );
 a45779a <=( (not A236)  and  A235 );
 a45780a <=( a45779a  and  a45776a );
 a45783a <=( A299  and  (not A298) );
 a45786a <=( A302  and  (not A301) );
 a45787a <=( a45786a  and  a45783a );
 a45788a <=( a45787a  and  a45780a );
 a45791a <=( A168  and  A169 );
 a45794a <=( A166  and  (not A167) );
 a45795a <=( a45794a  and  a45791a );
 a45798a <=( A200  and  (not A199) );
 a45801a <=( A202  and  (not A201) );
 a45802a <=( a45801a  and  a45798a );
 a45803a <=( a45802a  and  a45795a );
 a45806a <=( A233  and  A232 );
 a45809a <=( (not A236)  and  A235 );
 a45810a <=( a45809a  and  a45806a );
 a45813a <=( (not A299)  and  (not A298) );
 a45816a <=( (not A302)  and  A301 );
 a45817a <=( a45816a  and  a45813a );
 a45818a <=( a45817a  and  a45810a );
 a45821a <=( A168  and  A169 );
 a45824a <=( A166  and  (not A167) );
 a45825a <=( a45824a  and  a45821a );
 a45828a <=( A200  and  (not A199) );
 a45831a <=( A202  and  (not A201) );
 a45832a <=( a45831a  and  a45828a );
 a45833a <=( a45832a  and  a45825a );
 a45836a <=( A233  and  A232 );
 a45839a <=( (not A236)  and  A235 );
 a45840a <=( a45839a  and  a45836a );
 a45843a <=( A266  and  A265 );
 a45846a <=( (not A269)  and  A268 );
 a45847a <=( a45846a  and  a45843a );
 a45848a <=( a45847a  and  a45840a );
 a45851a <=( A168  and  A169 );
 a45854a <=( A166  and  (not A167) );
 a45855a <=( a45854a  and  a45851a );
 a45858a <=( A200  and  (not A199) );
 a45861a <=( A202  and  (not A201) );
 a45862a <=( a45861a  and  a45858a );
 a45863a <=( a45862a  and  a45855a );
 a45866a <=( A233  and  A232 );
 a45869a <=( (not A236)  and  A235 );
 a45870a <=( a45869a  and  a45866a );
 a45873a <=( A266  and  (not A265) );
 a45876a <=( A269  and  (not A268) );
 a45877a <=( a45876a  and  a45873a );
 a45878a <=( a45877a  and  a45870a );
 a45881a <=( A168  and  A169 );
 a45884a <=( A166  and  (not A167) );
 a45885a <=( a45884a  and  a45881a );
 a45888a <=( A200  and  (not A199) );
 a45891a <=( A202  and  (not A201) );
 a45892a <=( a45891a  and  a45888a );
 a45893a <=( a45892a  and  a45885a );
 a45896a <=( A233  and  A232 );
 a45899a <=( (not A236)  and  A235 );
 a45900a <=( a45899a  and  a45896a );
 a45903a <=( (not A266)  and  A265 );
 a45906a <=( A269  and  (not A268) );
 a45907a <=( a45906a  and  a45903a );
 a45908a <=( a45907a  and  a45900a );
 a45911a <=( A168  and  A169 );
 a45914a <=( A166  and  (not A167) );
 a45915a <=( a45914a  and  a45911a );
 a45918a <=( A200  and  (not A199) );
 a45921a <=( A202  and  (not A201) );
 a45922a <=( a45921a  and  a45918a );
 a45923a <=( a45922a  and  a45915a );
 a45926a <=( A233  and  A232 );
 a45929a <=( (not A236)  and  A235 );
 a45930a <=( a45929a  and  a45926a );
 a45933a <=( (not A266)  and  (not A265) );
 a45936a <=( (not A269)  and  A268 );
 a45937a <=( a45936a  and  a45933a );
 a45938a <=( a45937a  and  a45930a );
 a45941a <=( A168  and  A169 );
 a45944a <=( A166  and  (not A167) );
 a45945a <=( a45944a  and  a45941a );
 a45948a <=( A200  and  (not A199) );
 a45951a <=( A202  and  (not A201) );
 a45952a <=( a45951a  and  a45948a );
 a45953a <=( a45952a  and  a45945a );
 a45956a <=( A233  and  (not A232) );
 a45959a <=( A236  and  (not A235) );
 a45960a <=( a45959a  and  a45956a );
 a45963a <=( A299  and  A298 );
 a45966a <=( (not A302)  and  A301 );
 a45967a <=( a45966a  and  a45963a );
 a45968a <=( a45967a  and  a45960a );
 a45971a <=( A168  and  A169 );
 a45974a <=( A166  and  (not A167) );
 a45975a <=( a45974a  and  a45971a );
 a45978a <=( A200  and  (not A199) );
 a45981a <=( A202  and  (not A201) );
 a45982a <=( a45981a  and  a45978a );
 a45983a <=( a45982a  and  a45975a );
 a45986a <=( A233  and  (not A232) );
 a45989a <=( A236  and  (not A235) );
 a45990a <=( a45989a  and  a45986a );
 a45993a <=( (not A299)  and  A298 );
 a45996a <=( A302  and  (not A301) );
 a45997a <=( a45996a  and  a45993a );
 a45998a <=( a45997a  and  a45990a );
 a46001a <=( A168  and  A169 );
 a46004a <=( A166  and  (not A167) );
 a46005a <=( a46004a  and  a46001a );
 a46008a <=( A200  and  (not A199) );
 a46011a <=( A202  and  (not A201) );
 a46012a <=( a46011a  and  a46008a );
 a46013a <=( a46012a  and  a46005a );
 a46016a <=( A233  and  (not A232) );
 a46019a <=( A236  and  (not A235) );
 a46020a <=( a46019a  and  a46016a );
 a46023a <=( A299  and  (not A298) );
 a46026a <=( A302  and  (not A301) );
 a46027a <=( a46026a  and  a46023a );
 a46028a <=( a46027a  and  a46020a );
 a46031a <=( A168  and  A169 );
 a46034a <=( A166  and  (not A167) );
 a46035a <=( a46034a  and  a46031a );
 a46038a <=( A200  and  (not A199) );
 a46041a <=( A202  and  (not A201) );
 a46042a <=( a46041a  and  a46038a );
 a46043a <=( a46042a  and  a46035a );
 a46046a <=( A233  and  (not A232) );
 a46049a <=( A236  and  (not A235) );
 a46050a <=( a46049a  and  a46046a );
 a46053a <=( (not A299)  and  (not A298) );
 a46056a <=( (not A302)  and  A301 );
 a46057a <=( a46056a  and  a46053a );
 a46058a <=( a46057a  and  a46050a );
 a46061a <=( A168  and  A169 );
 a46064a <=( A166  and  (not A167) );
 a46065a <=( a46064a  and  a46061a );
 a46068a <=( A200  and  (not A199) );
 a46071a <=( A202  and  (not A201) );
 a46072a <=( a46071a  and  a46068a );
 a46073a <=( a46072a  and  a46065a );
 a46076a <=( A233  and  (not A232) );
 a46079a <=( A236  and  (not A235) );
 a46080a <=( a46079a  and  a46076a );
 a46083a <=( A266  and  A265 );
 a46086a <=( (not A269)  and  A268 );
 a46087a <=( a46086a  and  a46083a );
 a46088a <=( a46087a  and  a46080a );
 a46091a <=( A168  and  A169 );
 a46094a <=( A166  and  (not A167) );
 a46095a <=( a46094a  and  a46091a );
 a46098a <=( A200  and  (not A199) );
 a46101a <=( A202  and  (not A201) );
 a46102a <=( a46101a  and  a46098a );
 a46103a <=( a46102a  and  a46095a );
 a46106a <=( A233  and  (not A232) );
 a46109a <=( A236  and  (not A235) );
 a46110a <=( a46109a  and  a46106a );
 a46113a <=( A266  and  (not A265) );
 a46116a <=( A269  and  (not A268) );
 a46117a <=( a46116a  and  a46113a );
 a46118a <=( a46117a  and  a46110a );
 a46121a <=( A168  and  A169 );
 a46124a <=( A166  and  (not A167) );
 a46125a <=( a46124a  and  a46121a );
 a46128a <=( A200  and  (not A199) );
 a46131a <=( A202  and  (not A201) );
 a46132a <=( a46131a  and  a46128a );
 a46133a <=( a46132a  and  a46125a );
 a46136a <=( A233  and  (not A232) );
 a46139a <=( A236  and  (not A235) );
 a46140a <=( a46139a  and  a46136a );
 a46143a <=( (not A266)  and  A265 );
 a46146a <=( A269  and  (not A268) );
 a46147a <=( a46146a  and  a46143a );
 a46148a <=( a46147a  and  a46140a );
 a46151a <=( A168  and  A169 );
 a46154a <=( A166  and  (not A167) );
 a46155a <=( a46154a  and  a46151a );
 a46158a <=( A200  and  (not A199) );
 a46161a <=( A202  and  (not A201) );
 a46162a <=( a46161a  and  a46158a );
 a46163a <=( a46162a  and  a46155a );
 a46166a <=( A233  and  (not A232) );
 a46169a <=( A236  and  (not A235) );
 a46170a <=( a46169a  and  a46166a );
 a46173a <=( (not A266)  and  (not A265) );
 a46176a <=( (not A269)  and  A268 );
 a46177a <=( a46176a  and  a46173a );
 a46178a <=( a46177a  and  a46170a );
 a46181a <=( A168  and  A169 );
 a46184a <=( A166  and  (not A167) );
 a46185a <=( a46184a  and  a46181a );
 a46188a <=( A200  and  (not A199) );
 a46191a <=( A202  and  (not A201) );
 a46192a <=( a46191a  and  a46188a );
 a46193a <=( a46192a  and  a46185a );
 a46196a <=( (not A233)  and  A232 );
 a46199a <=( A236  and  (not A235) );
 a46200a <=( a46199a  and  a46196a );
 a46203a <=( A299  and  A298 );
 a46206a <=( (not A302)  and  A301 );
 a46207a <=( a46206a  and  a46203a );
 a46208a <=( a46207a  and  a46200a );
 a46211a <=( A168  and  A169 );
 a46214a <=( A166  and  (not A167) );
 a46215a <=( a46214a  and  a46211a );
 a46218a <=( A200  and  (not A199) );
 a46221a <=( A202  and  (not A201) );
 a46222a <=( a46221a  and  a46218a );
 a46223a <=( a46222a  and  a46215a );
 a46226a <=( (not A233)  and  A232 );
 a46229a <=( A236  and  (not A235) );
 a46230a <=( a46229a  and  a46226a );
 a46233a <=( (not A299)  and  A298 );
 a46236a <=( A302  and  (not A301) );
 a46237a <=( a46236a  and  a46233a );
 a46238a <=( a46237a  and  a46230a );
 a46241a <=( A168  and  A169 );
 a46244a <=( A166  and  (not A167) );
 a46245a <=( a46244a  and  a46241a );
 a46248a <=( A200  and  (not A199) );
 a46251a <=( A202  and  (not A201) );
 a46252a <=( a46251a  and  a46248a );
 a46253a <=( a46252a  and  a46245a );
 a46256a <=( (not A233)  and  A232 );
 a46259a <=( A236  and  (not A235) );
 a46260a <=( a46259a  and  a46256a );
 a46263a <=( A299  and  (not A298) );
 a46266a <=( A302  and  (not A301) );
 a46267a <=( a46266a  and  a46263a );
 a46268a <=( a46267a  and  a46260a );
 a46271a <=( A168  and  A169 );
 a46274a <=( A166  and  (not A167) );
 a46275a <=( a46274a  and  a46271a );
 a46278a <=( A200  and  (not A199) );
 a46281a <=( A202  and  (not A201) );
 a46282a <=( a46281a  and  a46278a );
 a46283a <=( a46282a  and  a46275a );
 a46286a <=( (not A233)  and  A232 );
 a46289a <=( A236  and  (not A235) );
 a46290a <=( a46289a  and  a46286a );
 a46293a <=( (not A299)  and  (not A298) );
 a46296a <=( (not A302)  and  A301 );
 a46297a <=( a46296a  and  a46293a );
 a46298a <=( a46297a  and  a46290a );
 a46301a <=( A168  and  A169 );
 a46304a <=( A166  and  (not A167) );
 a46305a <=( a46304a  and  a46301a );
 a46308a <=( A200  and  (not A199) );
 a46311a <=( A202  and  (not A201) );
 a46312a <=( a46311a  and  a46308a );
 a46313a <=( a46312a  and  a46305a );
 a46316a <=( (not A233)  and  A232 );
 a46319a <=( A236  and  (not A235) );
 a46320a <=( a46319a  and  a46316a );
 a46323a <=( A266  and  A265 );
 a46326a <=( (not A269)  and  A268 );
 a46327a <=( a46326a  and  a46323a );
 a46328a <=( a46327a  and  a46320a );
 a46331a <=( A168  and  A169 );
 a46334a <=( A166  and  (not A167) );
 a46335a <=( a46334a  and  a46331a );
 a46338a <=( A200  and  (not A199) );
 a46341a <=( A202  and  (not A201) );
 a46342a <=( a46341a  and  a46338a );
 a46343a <=( a46342a  and  a46335a );
 a46346a <=( (not A233)  and  A232 );
 a46349a <=( A236  and  (not A235) );
 a46350a <=( a46349a  and  a46346a );
 a46353a <=( A266  and  (not A265) );
 a46356a <=( A269  and  (not A268) );
 a46357a <=( a46356a  and  a46353a );
 a46358a <=( a46357a  and  a46350a );
 a46361a <=( A168  and  A169 );
 a46364a <=( A166  and  (not A167) );
 a46365a <=( a46364a  and  a46361a );
 a46368a <=( A200  and  (not A199) );
 a46371a <=( A202  and  (not A201) );
 a46372a <=( a46371a  and  a46368a );
 a46373a <=( a46372a  and  a46365a );
 a46376a <=( (not A233)  and  A232 );
 a46379a <=( A236  and  (not A235) );
 a46380a <=( a46379a  and  a46376a );
 a46383a <=( (not A266)  and  A265 );
 a46386a <=( A269  and  (not A268) );
 a46387a <=( a46386a  and  a46383a );
 a46388a <=( a46387a  and  a46380a );
 a46391a <=( A168  and  A169 );
 a46394a <=( A166  and  (not A167) );
 a46395a <=( a46394a  and  a46391a );
 a46398a <=( A200  and  (not A199) );
 a46401a <=( A202  and  (not A201) );
 a46402a <=( a46401a  and  a46398a );
 a46403a <=( a46402a  and  a46395a );
 a46406a <=( (not A233)  and  A232 );
 a46409a <=( A236  and  (not A235) );
 a46410a <=( a46409a  and  a46406a );
 a46413a <=( (not A266)  and  (not A265) );
 a46416a <=( (not A269)  and  A268 );
 a46417a <=( a46416a  and  a46413a );
 a46418a <=( a46417a  and  a46410a );
 a46421a <=( A168  and  A169 );
 a46424a <=( A166  and  (not A167) );
 a46425a <=( a46424a  and  a46421a );
 a46428a <=( A200  and  (not A199) );
 a46431a <=( A202  and  (not A201) );
 a46432a <=( a46431a  and  a46428a );
 a46433a <=( a46432a  and  a46425a );
 a46436a <=( (not A233)  and  (not A232) );
 a46439a <=( (not A236)  and  A235 );
 a46440a <=( a46439a  and  a46436a );
 a46443a <=( A299  and  A298 );
 a46446a <=( (not A302)  and  A301 );
 a46447a <=( a46446a  and  a46443a );
 a46448a <=( a46447a  and  a46440a );
 a46451a <=( A168  and  A169 );
 a46454a <=( A166  and  (not A167) );
 a46455a <=( a46454a  and  a46451a );
 a46458a <=( A200  and  (not A199) );
 a46461a <=( A202  and  (not A201) );
 a46462a <=( a46461a  and  a46458a );
 a46463a <=( a46462a  and  a46455a );
 a46466a <=( (not A233)  and  (not A232) );
 a46469a <=( (not A236)  and  A235 );
 a46470a <=( a46469a  and  a46466a );
 a46473a <=( (not A299)  and  A298 );
 a46476a <=( A302  and  (not A301) );
 a46477a <=( a46476a  and  a46473a );
 a46478a <=( a46477a  and  a46470a );
 a46481a <=( A168  and  A169 );
 a46484a <=( A166  and  (not A167) );
 a46485a <=( a46484a  and  a46481a );
 a46488a <=( A200  and  (not A199) );
 a46491a <=( A202  and  (not A201) );
 a46492a <=( a46491a  and  a46488a );
 a46493a <=( a46492a  and  a46485a );
 a46496a <=( (not A233)  and  (not A232) );
 a46499a <=( (not A236)  and  A235 );
 a46500a <=( a46499a  and  a46496a );
 a46503a <=( A299  and  (not A298) );
 a46506a <=( A302  and  (not A301) );
 a46507a <=( a46506a  and  a46503a );
 a46508a <=( a46507a  and  a46500a );
 a46511a <=( A168  and  A169 );
 a46514a <=( A166  and  (not A167) );
 a46515a <=( a46514a  and  a46511a );
 a46518a <=( A200  and  (not A199) );
 a46521a <=( A202  and  (not A201) );
 a46522a <=( a46521a  and  a46518a );
 a46523a <=( a46522a  and  a46515a );
 a46526a <=( (not A233)  and  (not A232) );
 a46529a <=( (not A236)  and  A235 );
 a46530a <=( a46529a  and  a46526a );
 a46533a <=( (not A299)  and  (not A298) );
 a46536a <=( (not A302)  and  A301 );
 a46537a <=( a46536a  and  a46533a );
 a46538a <=( a46537a  and  a46530a );
 a46541a <=( A168  and  A169 );
 a46544a <=( A166  and  (not A167) );
 a46545a <=( a46544a  and  a46541a );
 a46548a <=( A200  and  (not A199) );
 a46551a <=( A202  and  (not A201) );
 a46552a <=( a46551a  and  a46548a );
 a46553a <=( a46552a  and  a46545a );
 a46556a <=( (not A233)  and  (not A232) );
 a46559a <=( (not A236)  and  A235 );
 a46560a <=( a46559a  and  a46556a );
 a46563a <=( A266  and  A265 );
 a46566a <=( (not A269)  and  A268 );
 a46567a <=( a46566a  and  a46563a );
 a46568a <=( a46567a  and  a46560a );
 a46571a <=( A168  and  A169 );
 a46574a <=( A166  and  (not A167) );
 a46575a <=( a46574a  and  a46571a );
 a46578a <=( A200  and  (not A199) );
 a46581a <=( A202  and  (not A201) );
 a46582a <=( a46581a  and  a46578a );
 a46583a <=( a46582a  and  a46575a );
 a46586a <=( (not A233)  and  (not A232) );
 a46589a <=( (not A236)  and  A235 );
 a46590a <=( a46589a  and  a46586a );
 a46593a <=( A266  and  (not A265) );
 a46596a <=( A269  and  (not A268) );
 a46597a <=( a46596a  and  a46593a );
 a46598a <=( a46597a  and  a46590a );
 a46601a <=( A168  and  A169 );
 a46604a <=( A166  and  (not A167) );
 a46605a <=( a46604a  and  a46601a );
 a46608a <=( A200  and  (not A199) );
 a46611a <=( A202  and  (not A201) );
 a46612a <=( a46611a  and  a46608a );
 a46613a <=( a46612a  and  a46605a );
 a46616a <=( (not A233)  and  (not A232) );
 a46619a <=( (not A236)  and  A235 );
 a46620a <=( a46619a  and  a46616a );
 a46623a <=( (not A266)  and  A265 );
 a46626a <=( A269  and  (not A268) );
 a46627a <=( a46626a  and  a46623a );
 a46628a <=( a46627a  and  a46620a );
 a46631a <=( A168  and  A169 );
 a46634a <=( A166  and  (not A167) );
 a46635a <=( a46634a  and  a46631a );
 a46638a <=( A200  and  (not A199) );
 a46641a <=( A202  and  (not A201) );
 a46642a <=( a46641a  and  a46638a );
 a46643a <=( a46642a  and  a46635a );
 a46646a <=( (not A233)  and  (not A232) );
 a46649a <=( (not A236)  and  A235 );
 a46650a <=( a46649a  and  a46646a );
 a46653a <=( (not A266)  and  (not A265) );
 a46656a <=( (not A269)  and  A268 );
 a46657a <=( a46656a  and  a46653a );
 a46658a <=( a46657a  and  a46650a );
 a46661a <=( A168  and  A169 );
 a46664a <=( A166  and  (not A167) );
 a46665a <=( a46664a  and  a46661a );
 a46668a <=( A200  and  (not A199) );
 a46671a <=( (not A203)  and  (not A201) );
 a46672a <=( a46671a  and  a46668a );
 a46673a <=( a46672a  and  a46665a );
 a46676a <=( A233  and  A232 );
 a46679a <=( (not A236)  and  A235 );
 a46680a <=( a46679a  and  a46676a );
 a46683a <=( A299  and  A298 );
 a46686a <=( (not A302)  and  A301 );
 a46687a <=( a46686a  and  a46683a );
 a46688a <=( a46687a  and  a46680a );
 a46691a <=( A168  and  A169 );
 a46694a <=( A166  and  (not A167) );
 a46695a <=( a46694a  and  a46691a );
 a46698a <=( A200  and  (not A199) );
 a46701a <=( (not A203)  and  (not A201) );
 a46702a <=( a46701a  and  a46698a );
 a46703a <=( a46702a  and  a46695a );
 a46706a <=( A233  and  A232 );
 a46709a <=( (not A236)  and  A235 );
 a46710a <=( a46709a  and  a46706a );
 a46713a <=( (not A299)  and  A298 );
 a46716a <=( A302  and  (not A301) );
 a46717a <=( a46716a  and  a46713a );
 a46718a <=( a46717a  and  a46710a );
 a46721a <=( A168  and  A169 );
 a46724a <=( A166  and  (not A167) );
 a46725a <=( a46724a  and  a46721a );
 a46728a <=( A200  and  (not A199) );
 a46731a <=( (not A203)  and  (not A201) );
 a46732a <=( a46731a  and  a46728a );
 a46733a <=( a46732a  and  a46725a );
 a46736a <=( A233  and  A232 );
 a46739a <=( (not A236)  and  A235 );
 a46740a <=( a46739a  and  a46736a );
 a46743a <=( A299  and  (not A298) );
 a46746a <=( A302  and  (not A301) );
 a46747a <=( a46746a  and  a46743a );
 a46748a <=( a46747a  and  a46740a );
 a46751a <=( A168  and  A169 );
 a46754a <=( A166  and  (not A167) );
 a46755a <=( a46754a  and  a46751a );
 a46758a <=( A200  and  (not A199) );
 a46761a <=( (not A203)  and  (not A201) );
 a46762a <=( a46761a  and  a46758a );
 a46763a <=( a46762a  and  a46755a );
 a46766a <=( A233  and  A232 );
 a46769a <=( (not A236)  and  A235 );
 a46770a <=( a46769a  and  a46766a );
 a46773a <=( (not A299)  and  (not A298) );
 a46776a <=( (not A302)  and  A301 );
 a46777a <=( a46776a  and  a46773a );
 a46778a <=( a46777a  and  a46770a );
 a46781a <=( A168  and  A169 );
 a46784a <=( A166  and  (not A167) );
 a46785a <=( a46784a  and  a46781a );
 a46788a <=( A200  and  (not A199) );
 a46791a <=( (not A203)  and  (not A201) );
 a46792a <=( a46791a  and  a46788a );
 a46793a <=( a46792a  and  a46785a );
 a46796a <=( A233  and  A232 );
 a46799a <=( (not A236)  and  A235 );
 a46800a <=( a46799a  and  a46796a );
 a46803a <=( A266  and  A265 );
 a46806a <=( (not A269)  and  A268 );
 a46807a <=( a46806a  and  a46803a );
 a46808a <=( a46807a  and  a46800a );
 a46811a <=( A168  and  A169 );
 a46814a <=( A166  and  (not A167) );
 a46815a <=( a46814a  and  a46811a );
 a46818a <=( A200  and  (not A199) );
 a46821a <=( (not A203)  and  (not A201) );
 a46822a <=( a46821a  and  a46818a );
 a46823a <=( a46822a  and  a46815a );
 a46826a <=( A233  and  A232 );
 a46829a <=( (not A236)  and  A235 );
 a46830a <=( a46829a  and  a46826a );
 a46833a <=( A266  and  (not A265) );
 a46836a <=( A269  and  (not A268) );
 a46837a <=( a46836a  and  a46833a );
 a46838a <=( a46837a  and  a46830a );
 a46841a <=( A168  and  A169 );
 a46844a <=( A166  and  (not A167) );
 a46845a <=( a46844a  and  a46841a );
 a46848a <=( A200  and  (not A199) );
 a46851a <=( (not A203)  and  (not A201) );
 a46852a <=( a46851a  and  a46848a );
 a46853a <=( a46852a  and  a46845a );
 a46856a <=( A233  and  A232 );
 a46859a <=( (not A236)  and  A235 );
 a46860a <=( a46859a  and  a46856a );
 a46863a <=( (not A266)  and  A265 );
 a46866a <=( A269  and  (not A268) );
 a46867a <=( a46866a  and  a46863a );
 a46868a <=( a46867a  and  a46860a );
 a46871a <=( A168  and  A169 );
 a46874a <=( A166  and  (not A167) );
 a46875a <=( a46874a  and  a46871a );
 a46878a <=( A200  and  (not A199) );
 a46881a <=( (not A203)  and  (not A201) );
 a46882a <=( a46881a  and  a46878a );
 a46883a <=( a46882a  and  a46875a );
 a46886a <=( A233  and  A232 );
 a46889a <=( (not A236)  and  A235 );
 a46890a <=( a46889a  and  a46886a );
 a46893a <=( (not A266)  and  (not A265) );
 a46896a <=( (not A269)  and  A268 );
 a46897a <=( a46896a  and  a46893a );
 a46898a <=( a46897a  and  a46890a );
 a46901a <=( A168  and  A169 );
 a46904a <=( A166  and  (not A167) );
 a46905a <=( a46904a  and  a46901a );
 a46908a <=( A200  and  (not A199) );
 a46911a <=( (not A203)  and  (not A201) );
 a46912a <=( a46911a  and  a46908a );
 a46913a <=( a46912a  and  a46905a );
 a46916a <=( A233  and  (not A232) );
 a46919a <=( A236  and  (not A235) );
 a46920a <=( a46919a  and  a46916a );
 a46923a <=( A299  and  A298 );
 a46926a <=( (not A302)  and  A301 );
 a46927a <=( a46926a  and  a46923a );
 a46928a <=( a46927a  and  a46920a );
 a46931a <=( A168  and  A169 );
 a46934a <=( A166  and  (not A167) );
 a46935a <=( a46934a  and  a46931a );
 a46938a <=( A200  and  (not A199) );
 a46941a <=( (not A203)  and  (not A201) );
 a46942a <=( a46941a  and  a46938a );
 a46943a <=( a46942a  and  a46935a );
 a46946a <=( A233  and  (not A232) );
 a46949a <=( A236  and  (not A235) );
 a46950a <=( a46949a  and  a46946a );
 a46953a <=( (not A299)  and  A298 );
 a46956a <=( A302  and  (not A301) );
 a46957a <=( a46956a  and  a46953a );
 a46958a <=( a46957a  and  a46950a );
 a46961a <=( A168  and  A169 );
 a46964a <=( A166  and  (not A167) );
 a46965a <=( a46964a  and  a46961a );
 a46968a <=( A200  and  (not A199) );
 a46971a <=( (not A203)  and  (not A201) );
 a46972a <=( a46971a  and  a46968a );
 a46973a <=( a46972a  and  a46965a );
 a46976a <=( A233  and  (not A232) );
 a46979a <=( A236  and  (not A235) );
 a46980a <=( a46979a  and  a46976a );
 a46983a <=( A299  and  (not A298) );
 a46986a <=( A302  and  (not A301) );
 a46987a <=( a46986a  and  a46983a );
 a46988a <=( a46987a  and  a46980a );
 a46991a <=( A168  and  A169 );
 a46994a <=( A166  and  (not A167) );
 a46995a <=( a46994a  and  a46991a );
 a46998a <=( A200  and  (not A199) );
 a47001a <=( (not A203)  and  (not A201) );
 a47002a <=( a47001a  and  a46998a );
 a47003a <=( a47002a  and  a46995a );
 a47006a <=( A233  and  (not A232) );
 a47009a <=( A236  and  (not A235) );
 a47010a <=( a47009a  and  a47006a );
 a47013a <=( (not A299)  and  (not A298) );
 a47016a <=( (not A302)  and  A301 );
 a47017a <=( a47016a  and  a47013a );
 a47018a <=( a47017a  and  a47010a );
 a47021a <=( A168  and  A169 );
 a47024a <=( A166  and  (not A167) );
 a47025a <=( a47024a  and  a47021a );
 a47028a <=( A200  and  (not A199) );
 a47031a <=( (not A203)  and  (not A201) );
 a47032a <=( a47031a  and  a47028a );
 a47033a <=( a47032a  and  a47025a );
 a47036a <=( A233  and  (not A232) );
 a47039a <=( A236  and  (not A235) );
 a47040a <=( a47039a  and  a47036a );
 a47043a <=( A266  and  A265 );
 a47046a <=( (not A269)  and  A268 );
 a47047a <=( a47046a  and  a47043a );
 a47048a <=( a47047a  and  a47040a );
 a47051a <=( A168  and  A169 );
 a47054a <=( A166  and  (not A167) );
 a47055a <=( a47054a  and  a47051a );
 a47058a <=( A200  and  (not A199) );
 a47061a <=( (not A203)  and  (not A201) );
 a47062a <=( a47061a  and  a47058a );
 a47063a <=( a47062a  and  a47055a );
 a47066a <=( A233  and  (not A232) );
 a47069a <=( A236  and  (not A235) );
 a47070a <=( a47069a  and  a47066a );
 a47073a <=( A266  and  (not A265) );
 a47076a <=( A269  and  (not A268) );
 a47077a <=( a47076a  and  a47073a );
 a47078a <=( a47077a  and  a47070a );
 a47081a <=( A168  and  A169 );
 a47084a <=( A166  and  (not A167) );
 a47085a <=( a47084a  and  a47081a );
 a47088a <=( A200  and  (not A199) );
 a47091a <=( (not A203)  and  (not A201) );
 a47092a <=( a47091a  and  a47088a );
 a47093a <=( a47092a  and  a47085a );
 a47096a <=( A233  and  (not A232) );
 a47099a <=( A236  and  (not A235) );
 a47100a <=( a47099a  and  a47096a );
 a47103a <=( (not A266)  and  A265 );
 a47106a <=( A269  and  (not A268) );
 a47107a <=( a47106a  and  a47103a );
 a47108a <=( a47107a  and  a47100a );
 a47111a <=( A168  and  A169 );
 a47114a <=( A166  and  (not A167) );
 a47115a <=( a47114a  and  a47111a );
 a47118a <=( A200  and  (not A199) );
 a47121a <=( (not A203)  and  (not A201) );
 a47122a <=( a47121a  and  a47118a );
 a47123a <=( a47122a  and  a47115a );
 a47126a <=( A233  and  (not A232) );
 a47129a <=( A236  and  (not A235) );
 a47130a <=( a47129a  and  a47126a );
 a47133a <=( (not A266)  and  (not A265) );
 a47136a <=( (not A269)  and  A268 );
 a47137a <=( a47136a  and  a47133a );
 a47138a <=( a47137a  and  a47130a );
 a47141a <=( A168  and  A169 );
 a47144a <=( A166  and  (not A167) );
 a47145a <=( a47144a  and  a47141a );
 a47148a <=( A200  and  (not A199) );
 a47151a <=( (not A203)  and  (not A201) );
 a47152a <=( a47151a  and  a47148a );
 a47153a <=( a47152a  and  a47145a );
 a47156a <=( (not A233)  and  A232 );
 a47159a <=( A236  and  (not A235) );
 a47160a <=( a47159a  and  a47156a );
 a47163a <=( A299  and  A298 );
 a47166a <=( (not A302)  and  A301 );
 a47167a <=( a47166a  and  a47163a );
 a47168a <=( a47167a  and  a47160a );
 a47171a <=( A168  and  A169 );
 a47174a <=( A166  and  (not A167) );
 a47175a <=( a47174a  and  a47171a );
 a47178a <=( A200  and  (not A199) );
 a47181a <=( (not A203)  and  (not A201) );
 a47182a <=( a47181a  and  a47178a );
 a47183a <=( a47182a  and  a47175a );
 a47186a <=( (not A233)  and  A232 );
 a47189a <=( A236  and  (not A235) );
 a47190a <=( a47189a  and  a47186a );
 a47193a <=( (not A299)  and  A298 );
 a47196a <=( A302  and  (not A301) );
 a47197a <=( a47196a  and  a47193a );
 a47198a <=( a47197a  and  a47190a );
 a47201a <=( A168  and  A169 );
 a47204a <=( A166  and  (not A167) );
 a47205a <=( a47204a  and  a47201a );
 a47208a <=( A200  and  (not A199) );
 a47211a <=( (not A203)  and  (not A201) );
 a47212a <=( a47211a  and  a47208a );
 a47213a <=( a47212a  and  a47205a );
 a47216a <=( (not A233)  and  A232 );
 a47219a <=( A236  and  (not A235) );
 a47220a <=( a47219a  and  a47216a );
 a47223a <=( A299  and  (not A298) );
 a47226a <=( A302  and  (not A301) );
 a47227a <=( a47226a  and  a47223a );
 a47228a <=( a47227a  and  a47220a );
 a47231a <=( A168  and  A169 );
 a47234a <=( A166  and  (not A167) );
 a47235a <=( a47234a  and  a47231a );
 a47238a <=( A200  and  (not A199) );
 a47241a <=( (not A203)  and  (not A201) );
 a47242a <=( a47241a  and  a47238a );
 a47243a <=( a47242a  and  a47235a );
 a47246a <=( (not A233)  and  A232 );
 a47249a <=( A236  and  (not A235) );
 a47250a <=( a47249a  and  a47246a );
 a47253a <=( (not A299)  and  (not A298) );
 a47256a <=( (not A302)  and  A301 );
 a47257a <=( a47256a  and  a47253a );
 a47258a <=( a47257a  and  a47250a );
 a47261a <=( A168  and  A169 );
 a47264a <=( A166  and  (not A167) );
 a47265a <=( a47264a  and  a47261a );
 a47268a <=( A200  and  (not A199) );
 a47271a <=( (not A203)  and  (not A201) );
 a47272a <=( a47271a  and  a47268a );
 a47273a <=( a47272a  and  a47265a );
 a47276a <=( (not A233)  and  A232 );
 a47279a <=( A236  and  (not A235) );
 a47280a <=( a47279a  and  a47276a );
 a47283a <=( A266  and  A265 );
 a47286a <=( (not A269)  and  A268 );
 a47287a <=( a47286a  and  a47283a );
 a47288a <=( a47287a  and  a47280a );
 a47291a <=( A168  and  A169 );
 a47294a <=( A166  and  (not A167) );
 a47295a <=( a47294a  and  a47291a );
 a47298a <=( A200  and  (not A199) );
 a47301a <=( (not A203)  and  (not A201) );
 a47302a <=( a47301a  and  a47298a );
 a47303a <=( a47302a  and  a47295a );
 a47306a <=( (not A233)  and  A232 );
 a47309a <=( A236  and  (not A235) );
 a47310a <=( a47309a  and  a47306a );
 a47313a <=( A266  and  (not A265) );
 a47316a <=( A269  and  (not A268) );
 a47317a <=( a47316a  and  a47313a );
 a47318a <=( a47317a  and  a47310a );
 a47321a <=( A168  and  A169 );
 a47324a <=( A166  and  (not A167) );
 a47325a <=( a47324a  and  a47321a );
 a47328a <=( A200  and  (not A199) );
 a47331a <=( (not A203)  and  (not A201) );
 a47332a <=( a47331a  and  a47328a );
 a47333a <=( a47332a  and  a47325a );
 a47336a <=( (not A233)  and  A232 );
 a47339a <=( A236  and  (not A235) );
 a47340a <=( a47339a  and  a47336a );
 a47343a <=( (not A266)  and  A265 );
 a47346a <=( A269  and  (not A268) );
 a47347a <=( a47346a  and  a47343a );
 a47348a <=( a47347a  and  a47340a );
 a47351a <=( A168  and  A169 );
 a47354a <=( A166  and  (not A167) );
 a47355a <=( a47354a  and  a47351a );
 a47358a <=( A200  and  (not A199) );
 a47361a <=( (not A203)  and  (not A201) );
 a47362a <=( a47361a  and  a47358a );
 a47363a <=( a47362a  and  a47355a );
 a47366a <=( (not A233)  and  A232 );
 a47369a <=( A236  and  (not A235) );
 a47370a <=( a47369a  and  a47366a );
 a47373a <=( (not A266)  and  (not A265) );
 a47376a <=( (not A269)  and  A268 );
 a47377a <=( a47376a  and  a47373a );
 a47378a <=( a47377a  and  a47370a );
 a47381a <=( A168  and  A169 );
 a47384a <=( A166  and  (not A167) );
 a47385a <=( a47384a  and  a47381a );
 a47388a <=( A200  and  (not A199) );
 a47391a <=( (not A203)  and  (not A201) );
 a47392a <=( a47391a  and  a47388a );
 a47393a <=( a47392a  and  a47385a );
 a47396a <=( (not A233)  and  (not A232) );
 a47399a <=( (not A236)  and  A235 );
 a47400a <=( a47399a  and  a47396a );
 a47403a <=( A299  and  A298 );
 a47406a <=( (not A302)  and  A301 );
 a47407a <=( a47406a  and  a47403a );
 a47408a <=( a47407a  and  a47400a );
 a47411a <=( A168  and  A169 );
 a47414a <=( A166  and  (not A167) );
 a47415a <=( a47414a  and  a47411a );
 a47418a <=( A200  and  (not A199) );
 a47421a <=( (not A203)  and  (not A201) );
 a47422a <=( a47421a  and  a47418a );
 a47423a <=( a47422a  and  a47415a );
 a47426a <=( (not A233)  and  (not A232) );
 a47429a <=( (not A236)  and  A235 );
 a47430a <=( a47429a  and  a47426a );
 a47433a <=( (not A299)  and  A298 );
 a47436a <=( A302  and  (not A301) );
 a47437a <=( a47436a  and  a47433a );
 a47438a <=( a47437a  and  a47430a );
 a47441a <=( A168  and  A169 );
 a47444a <=( A166  and  (not A167) );
 a47445a <=( a47444a  and  a47441a );
 a47448a <=( A200  and  (not A199) );
 a47451a <=( (not A203)  and  (not A201) );
 a47452a <=( a47451a  and  a47448a );
 a47453a <=( a47452a  and  a47445a );
 a47456a <=( (not A233)  and  (not A232) );
 a47459a <=( (not A236)  and  A235 );
 a47460a <=( a47459a  and  a47456a );
 a47463a <=( A299  and  (not A298) );
 a47466a <=( A302  and  (not A301) );
 a47467a <=( a47466a  and  a47463a );
 a47468a <=( a47467a  and  a47460a );
 a47471a <=( A168  and  A169 );
 a47474a <=( A166  and  (not A167) );
 a47475a <=( a47474a  and  a47471a );
 a47478a <=( A200  and  (not A199) );
 a47481a <=( (not A203)  and  (not A201) );
 a47482a <=( a47481a  and  a47478a );
 a47483a <=( a47482a  and  a47475a );
 a47486a <=( (not A233)  and  (not A232) );
 a47489a <=( (not A236)  and  A235 );
 a47490a <=( a47489a  and  a47486a );
 a47493a <=( (not A299)  and  (not A298) );
 a47496a <=( (not A302)  and  A301 );
 a47497a <=( a47496a  and  a47493a );
 a47498a <=( a47497a  and  a47490a );
 a47501a <=( A168  and  A169 );
 a47504a <=( A166  and  (not A167) );
 a47505a <=( a47504a  and  a47501a );
 a47508a <=( A200  and  (not A199) );
 a47511a <=( (not A203)  and  (not A201) );
 a47512a <=( a47511a  and  a47508a );
 a47513a <=( a47512a  and  a47505a );
 a47516a <=( (not A233)  and  (not A232) );
 a47519a <=( (not A236)  and  A235 );
 a47520a <=( a47519a  and  a47516a );
 a47523a <=( A266  and  A265 );
 a47526a <=( (not A269)  and  A268 );
 a47527a <=( a47526a  and  a47523a );
 a47528a <=( a47527a  and  a47520a );
 a47531a <=( A168  and  A169 );
 a47534a <=( A166  and  (not A167) );
 a47535a <=( a47534a  and  a47531a );
 a47538a <=( A200  and  (not A199) );
 a47541a <=( (not A203)  and  (not A201) );
 a47542a <=( a47541a  and  a47538a );
 a47543a <=( a47542a  and  a47535a );
 a47546a <=( (not A233)  and  (not A232) );
 a47549a <=( (not A236)  and  A235 );
 a47550a <=( a47549a  and  a47546a );
 a47553a <=( A266  and  (not A265) );
 a47556a <=( A269  and  (not A268) );
 a47557a <=( a47556a  and  a47553a );
 a47558a <=( a47557a  and  a47550a );
 a47561a <=( A168  and  A169 );
 a47564a <=( A166  and  (not A167) );
 a47565a <=( a47564a  and  a47561a );
 a47568a <=( A200  and  (not A199) );
 a47571a <=( (not A203)  and  (not A201) );
 a47572a <=( a47571a  and  a47568a );
 a47573a <=( a47572a  and  a47565a );
 a47576a <=( (not A233)  and  (not A232) );
 a47579a <=( (not A236)  and  A235 );
 a47580a <=( a47579a  and  a47576a );
 a47583a <=( (not A266)  and  A265 );
 a47586a <=( A269  and  (not A268) );
 a47587a <=( a47586a  and  a47583a );
 a47588a <=( a47587a  and  a47580a );
 a47591a <=( A168  and  A169 );
 a47594a <=( A166  and  (not A167) );
 a47595a <=( a47594a  and  a47591a );
 a47598a <=( A200  and  (not A199) );
 a47601a <=( (not A203)  and  (not A201) );
 a47602a <=( a47601a  and  a47598a );
 a47603a <=( a47602a  and  a47595a );
 a47606a <=( (not A233)  and  (not A232) );
 a47609a <=( (not A236)  and  A235 );
 a47610a <=( a47609a  and  a47606a );
 a47613a <=( (not A266)  and  (not A265) );
 a47616a <=( (not A269)  and  A268 );
 a47617a <=( a47616a  and  a47613a );
 a47618a <=( a47617a  and  a47610a );
 a47621a <=( A168  and  A169 );
 a47624a <=( A166  and  (not A167) );
 a47625a <=( a47624a  and  a47621a );
 a47628a <=( (not A200)  and  A199 );
 a47631a <=( A202  and  (not A201) );
 a47632a <=( a47631a  and  a47628a );
 a47633a <=( a47632a  and  a47625a );
 a47636a <=( A233  and  A232 );
 a47639a <=( (not A236)  and  A235 );
 a47640a <=( a47639a  and  a47636a );
 a47643a <=( A299  and  A298 );
 a47646a <=( (not A302)  and  A301 );
 a47647a <=( a47646a  and  a47643a );
 a47648a <=( a47647a  and  a47640a );
 a47651a <=( A168  and  A169 );
 a47654a <=( A166  and  (not A167) );
 a47655a <=( a47654a  and  a47651a );
 a47658a <=( (not A200)  and  A199 );
 a47661a <=( A202  and  (not A201) );
 a47662a <=( a47661a  and  a47658a );
 a47663a <=( a47662a  and  a47655a );
 a47666a <=( A233  and  A232 );
 a47669a <=( (not A236)  and  A235 );
 a47670a <=( a47669a  and  a47666a );
 a47673a <=( (not A299)  and  A298 );
 a47676a <=( A302  and  (not A301) );
 a47677a <=( a47676a  and  a47673a );
 a47678a <=( a47677a  and  a47670a );
 a47681a <=( A168  and  A169 );
 a47684a <=( A166  and  (not A167) );
 a47685a <=( a47684a  and  a47681a );
 a47688a <=( (not A200)  and  A199 );
 a47691a <=( A202  and  (not A201) );
 a47692a <=( a47691a  and  a47688a );
 a47693a <=( a47692a  and  a47685a );
 a47696a <=( A233  and  A232 );
 a47699a <=( (not A236)  and  A235 );
 a47700a <=( a47699a  and  a47696a );
 a47703a <=( A299  and  (not A298) );
 a47706a <=( A302  and  (not A301) );
 a47707a <=( a47706a  and  a47703a );
 a47708a <=( a47707a  and  a47700a );
 a47711a <=( A168  and  A169 );
 a47714a <=( A166  and  (not A167) );
 a47715a <=( a47714a  and  a47711a );
 a47718a <=( (not A200)  and  A199 );
 a47721a <=( A202  and  (not A201) );
 a47722a <=( a47721a  and  a47718a );
 a47723a <=( a47722a  and  a47715a );
 a47726a <=( A233  and  A232 );
 a47729a <=( (not A236)  and  A235 );
 a47730a <=( a47729a  and  a47726a );
 a47733a <=( (not A299)  and  (not A298) );
 a47736a <=( (not A302)  and  A301 );
 a47737a <=( a47736a  and  a47733a );
 a47738a <=( a47737a  and  a47730a );
 a47741a <=( A168  and  A169 );
 a47744a <=( A166  and  (not A167) );
 a47745a <=( a47744a  and  a47741a );
 a47748a <=( (not A200)  and  A199 );
 a47751a <=( A202  and  (not A201) );
 a47752a <=( a47751a  and  a47748a );
 a47753a <=( a47752a  and  a47745a );
 a47756a <=( A233  and  A232 );
 a47759a <=( (not A236)  and  A235 );
 a47760a <=( a47759a  and  a47756a );
 a47763a <=( A266  and  A265 );
 a47766a <=( (not A269)  and  A268 );
 a47767a <=( a47766a  and  a47763a );
 a47768a <=( a47767a  and  a47760a );
 a47771a <=( A168  and  A169 );
 a47774a <=( A166  and  (not A167) );
 a47775a <=( a47774a  and  a47771a );
 a47778a <=( (not A200)  and  A199 );
 a47781a <=( A202  and  (not A201) );
 a47782a <=( a47781a  and  a47778a );
 a47783a <=( a47782a  and  a47775a );
 a47786a <=( A233  and  A232 );
 a47789a <=( (not A236)  and  A235 );
 a47790a <=( a47789a  and  a47786a );
 a47793a <=( A266  and  (not A265) );
 a47796a <=( A269  and  (not A268) );
 a47797a <=( a47796a  and  a47793a );
 a47798a <=( a47797a  and  a47790a );
 a47801a <=( A168  and  A169 );
 a47804a <=( A166  and  (not A167) );
 a47805a <=( a47804a  and  a47801a );
 a47808a <=( (not A200)  and  A199 );
 a47811a <=( A202  and  (not A201) );
 a47812a <=( a47811a  and  a47808a );
 a47813a <=( a47812a  and  a47805a );
 a47816a <=( A233  and  A232 );
 a47819a <=( (not A236)  and  A235 );
 a47820a <=( a47819a  and  a47816a );
 a47823a <=( (not A266)  and  A265 );
 a47826a <=( A269  and  (not A268) );
 a47827a <=( a47826a  and  a47823a );
 a47828a <=( a47827a  and  a47820a );
 a47831a <=( A168  and  A169 );
 a47834a <=( A166  and  (not A167) );
 a47835a <=( a47834a  and  a47831a );
 a47838a <=( (not A200)  and  A199 );
 a47841a <=( A202  and  (not A201) );
 a47842a <=( a47841a  and  a47838a );
 a47843a <=( a47842a  and  a47835a );
 a47846a <=( A233  and  A232 );
 a47849a <=( (not A236)  and  A235 );
 a47850a <=( a47849a  and  a47846a );
 a47853a <=( (not A266)  and  (not A265) );
 a47856a <=( (not A269)  and  A268 );
 a47857a <=( a47856a  and  a47853a );
 a47858a <=( a47857a  and  a47850a );
 a47861a <=( A168  and  A169 );
 a47864a <=( A166  and  (not A167) );
 a47865a <=( a47864a  and  a47861a );
 a47868a <=( (not A200)  and  A199 );
 a47871a <=( A202  and  (not A201) );
 a47872a <=( a47871a  and  a47868a );
 a47873a <=( a47872a  and  a47865a );
 a47876a <=( A233  and  (not A232) );
 a47879a <=( A236  and  (not A235) );
 a47880a <=( a47879a  and  a47876a );
 a47883a <=( A299  and  A298 );
 a47886a <=( (not A302)  and  A301 );
 a47887a <=( a47886a  and  a47883a );
 a47888a <=( a47887a  and  a47880a );
 a47891a <=( A168  and  A169 );
 a47894a <=( A166  and  (not A167) );
 a47895a <=( a47894a  and  a47891a );
 a47898a <=( (not A200)  and  A199 );
 a47901a <=( A202  and  (not A201) );
 a47902a <=( a47901a  and  a47898a );
 a47903a <=( a47902a  and  a47895a );
 a47906a <=( A233  and  (not A232) );
 a47909a <=( A236  and  (not A235) );
 a47910a <=( a47909a  and  a47906a );
 a47913a <=( (not A299)  and  A298 );
 a47916a <=( A302  and  (not A301) );
 a47917a <=( a47916a  and  a47913a );
 a47918a <=( a47917a  and  a47910a );
 a47921a <=( A168  and  A169 );
 a47924a <=( A166  and  (not A167) );
 a47925a <=( a47924a  and  a47921a );
 a47928a <=( (not A200)  and  A199 );
 a47931a <=( A202  and  (not A201) );
 a47932a <=( a47931a  and  a47928a );
 a47933a <=( a47932a  and  a47925a );
 a47936a <=( A233  and  (not A232) );
 a47939a <=( A236  and  (not A235) );
 a47940a <=( a47939a  and  a47936a );
 a47943a <=( A299  and  (not A298) );
 a47946a <=( A302  and  (not A301) );
 a47947a <=( a47946a  and  a47943a );
 a47948a <=( a47947a  and  a47940a );
 a47951a <=( A168  and  A169 );
 a47954a <=( A166  and  (not A167) );
 a47955a <=( a47954a  and  a47951a );
 a47958a <=( (not A200)  and  A199 );
 a47961a <=( A202  and  (not A201) );
 a47962a <=( a47961a  and  a47958a );
 a47963a <=( a47962a  and  a47955a );
 a47966a <=( A233  and  (not A232) );
 a47969a <=( A236  and  (not A235) );
 a47970a <=( a47969a  and  a47966a );
 a47973a <=( (not A299)  and  (not A298) );
 a47976a <=( (not A302)  and  A301 );
 a47977a <=( a47976a  and  a47973a );
 a47978a <=( a47977a  and  a47970a );
 a47981a <=( A168  and  A169 );
 a47984a <=( A166  and  (not A167) );
 a47985a <=( a47984a  and  a47981a );
 a47988a <=( (not A200)  and  A199 );
 a47991a <=( A202  and  (not A201) );
 a47992a <=( a47991a  and  a47988a );
 a47993a <=( a47992a  and  a47985a );
 a47996a <=( A233  and  (not A232) );
 a47999a <=( A236  and  (not A235) );
 a48000a <=( a47999a  and  a47996a );
 a48003a <=( A266  and  A265 );
 a48006a <=( (not A269)  and  A268 );
 a48007a <=( a48006a  and  a48003a );
 a48008a <=( a48007a  and  a48000a );
 a48011a <=( A168  and  A169 );
 a48014a <=( A166  and  (not A167) );
 a48015a <=( a48014a  and  a48011a );
 a48018a <=( (not A200)  and  A199 );
 a48021a <=( A202  and  (not A201) );
 a48022a <=( a48021a  and  a48018a );
 a48023a <=( a48022a  and  a48015a );
 a48026a <=( A233  and  (not A232) );
 a48029a <=( A236  and  (not A235) );
 a48030a <=( a48029a  and  a48026a );
 a48033a <=( A266  and  (not A265) );
 a48036a <=( A269  and  (not A268) );
 a48037a <=( a48036a  and  a48033a );
 a48038a <=( a48037a  and  a48030a );
 a48041a <=( A168  and  A169 );
 a48044a <=( A166  and  (not A167) );
 a48045a <=( a48044a  and  a48041a );
 a48048a <=( (not A200)  and  A199 );
 a48051a <=( A202  and  (not A201) );
 a48052a <=( a48051a  and  a48048a );
 a48053a <=( a48052a  and  a48045a );
 a48056a <=( A233  and  (not A232) );
 a48059a <=( A236  and  (not A235) );
 a48060a <=( a48059a  and  a48056a );
 a48063a <=( (not A266)  and  A265 );
 a48066a <=( A269  and  (not A268) );
 a48067a <=( a48066a  and  a48063a );
 a48068a <=( a48067a  and  a48060a );
 a48071a <=( A168  and  A169 );
 a48074a <=( A166  and  (not A167) );
 a48075a <=( a48074a  and  a48071a );
 a48078a <=( (not A200)  and  A199 );
 a48081a <=( A202  and  (not A201) );
 a48082a <=( a48081a  and  a48078a );
 a48083a <=( a48082a  and  a48075a );
 a48086a <=( A233  and  (not A232) );
 a48089a <=( A236  and  (not A235) );
 a48090a <=( a48089a  and  a48086a );
 a48093a <=( (not A266)  and  (not A265) );
 a48096a <=( (not A269)  and  A268 );
 a48097a <=( a48096a  and  a48093a );
 a48098a <=( a48097a  and  a48090a );
 a48101a <=( A168  and  A169 );
 a48104a <=( A166  and  (not A167) );
 a48105a <=( a48104a  and  a48101a );
 a48108a <=( (not A200)  and  A199 );
 a48111a <=( A202  and  (not A201) );
 a48112a <=( a48111a  and  a48108a );
 a48113a <=( a48112a  and  a48105a );
 a48116a <=( (not A233)  and  A232 );
 a48119a <=( A236  and  (not A235) );
 a48120a <=( a48119a  and  a48116a );
 a48123a <=( A299  and  A298 );
 a48126a <=( (not A302)  and  A301 );
 a48127a <=( a48126a  and  a48123a );
 a48128a <=( a48127a  and  a48120a );
 a48131a <=( A168  and  A169 );
 a48134a <=( A166  and  (not A167) );
 a48135a <=( a48134a  and  a48131a );
 a48138a <=( (not A200)  and  A199 );
 a48141a <=( A202  and  (not A201) );
 a48142a <=( a48141a  and  a48138a );
 a48143a <=( a48142a  and  a48135a );
 a48146a <=( (not A233)  and  A232 );
 a48149a <=( A236  and  (not A235) );
 a48150a <=( a48149a  and  a48146a );
 a48153a <=( (not A299)  and  A298 );
 a48156a <=( A302  and  (not A301) );
 a48157a <=( a48156a  and  a48153a );
 a48158a <=( a48157a  and  a48150a );
 a48161a <=( A168  and  A169 );
 a48164a <=( A166  and  (not A167) );
 a48165a <=( a48164a  and  a48161a );
 a48168a <=( (not A200)  and  A199 );
 a48171a <=( A202  and  (not A201) );
 a48172a <=( a48171a  and  a48168a );
 a48173a <=( a48172a  and  a48165a );
 a48176a <=( (not A233)  and  A232 );
 a48179a <=( A236  and  (not A235) );
 a48180a <=( a48179a  and  a48176a );
 a48183a <=( A299  and  (not A298) );
 a48186a <=( A302  and  (not A301) );
 a48187a <=( a48186a  and  a48183a );
 a48188a <=( a48187a  and  a48180a );
 a48191a <=( A168  and  A169 );
 a48194a <=( A166  and  (not A167) );
 a48195a <=( a48194a  and  a48191a );
 a48198a <=( (not A200)  and  A199 );
 a48201a <=( A202  and  (not A201) );
 a48202a <=( a48201a  and  a48198a );
 a48203a <=( a48202a  and  a48195a );
 a48206a <=( (not A233)  and  A232 );
 a48209a <=( A236  and  (not A235) );
 a48210a <=( a48209a  and  a48206a );
 a48213a <=( (not A299)  and  (not A298) );
 a48216a <=( (not A302)  and  A301 );
 a48217a <=( a48216a  and  a48213a );
 a48218a <=( a48217a  and  a48210a );
 a48221a <=( A168  and  A169 );
 a48224a <=( A166  and  (not A167) );
 a48225a <=( a48224a  and  a48221a );
 a48228a <=( (not A200)  and  A199 );
 a48231a <=( A202  and  (not A201) );
 a48232a <=( a48231a  and  a48228a );
 a48233a <=( a48232a  and  a48225a );
 a48236a <=( (not A233)  and  A232 );
 a48239a <=( A236  and  (not A235) );
 a48240a <=( a48239a  and  a48236a );
 a48243a <=( A266  and  A265 );
 a48246a <=( (not A269)  and  A268 );
 a48247a <=( a48246a  and  a48243a );
 a48248a <=( a48247a  and  a48240a );
 a48251a <=( A168  and  A169 );
 a48254a <=( A166  and  (not A167) );
 a48255a <=( a48254a  and  a48251a );
 a48258a <=( (not A200)  and  A199 );
 a48261a <=( A202  and  (not A201) );
 a48262a <=( a48261a  and  a48258a );
 a48263a <=( a48262a  and  a48255a );
 a48266a <=( (not A233)  and  A232 );
 a48269a <=( A236  and  (not A235) );
 a48270a <=( a48269a  and  a48266a );
 a48273a <=( A266  and  (not A265) );
 a48276a <=( A269  and  (not A268) );
 a48277a <=( a48276a  and  a48273a );
 a48278a <=( a48277a  and  a48270a );
 a48281a <=( A168  and  A169 );
 a48284a <=( A166  and  (not A167) );
 a48285a <=( a48284a  and  a48281a );
 a48288a <=( (not A200)  and  A199 );
 a48291a <=( A202  and  (not A201) );
 a48292a <=( a48291a  and  a48288a );
 a48293a <=( a48292a  and  a48285a );
 a48296a <=( (not A233)  and  A232 );
 a48299a <=( A236  and  (not A235) );
 a48300a <=( a48299a  and  a48296a );
 a48303a <=( (not A266)  and  A265 );
 a48306a <=( A269  and  (not A268) );
 a48307a <=( a48306a  and  a48303a );
 a48308a <=( a48307a  and  a48300a );
 a48311a <=( A168  and  A169 );
 a48314a <=( A166  and  (not A167) );
 a48315a <=( a48314a  and  a48311a );
 a48318a <=( (not A200)  and  A199 );
 a48321a <=( A202  and  (not A201) );
 a48322a <=( a48321a  and  a48318a );
 a48323a <=( a48322a  and  a48315a );
 a48326a <=( (not A233)  and  A232 );
 a48329a <=( A236  and  (not A235) );
 a48330a <=( a48329a  and  a48326a );
 a48333a <=( (not A266)  and  (not A265) );
 a48336a <=( (not A269)  and  A268 );
 a48337a <=( a48336a  and  a48333a );
 a48338a <=( a48337a  and  a48330a );
 a48341a <=( A168  and  A169 );
 a48344a <=( A166  and  (not A167) );
 a48345a <=( a48344a  and  a48341a );
 a48348a <=( (not A200)  and  A199 );
 a48351a <=( A202  and  (not A201) );
 a48352a <=( a48351a  and  a48348a );
 a48353a <=( a48352a  and  a48345a );
 a48356a <=( (not A233)  and  (not A232) );
 a48359a <=( (not A236)  and  A235 );
 a48360a <=( a48359a  and  a48356a );
 a48363a <=( A299  and  A298 );
 a48366a <=( (not A302)  and  A301 );
 a48367a <=( a48366a  and  a48363a );
 a48368a <=( a48367a  and  a48360a );
 a48371a <=( A168  and  A169 );
 a48374a <=( A166  and  (not A167) );
 a48375a <=( a48374a  and  a48371a );
 a48378a <=( (not A200)  and  A199 );
 a48381a <=( A202  and  (not A201) );
 a48382a <=( a48381a  and  a48378a );
 a48383a <=( a48382a  and  a48375a );
 a48386a <=( (not A233)  and  (not A232) );
 a48389a <=( (not A236)  and  A235 );
 a48390a <=( a48389a  and  a48386a );
 a48393a <=( (not A299)  and  A298 );
 a48396a <=( A302  and  (not A301) );
 a48397a <=( a48396a  and  a48393a );
 a48398a <=( a48397a  and  a48390a );
 a48401a <=( A168  and  A169 );
 a48404a <=( A166  and  (not A167) );
 a48405a <=( a48404a  and  a48401a );
 a48408a <=( (not A200)  and  A199 );
 a48411a <=( A202  and  (not A201) );
 a48412a <=( a48411a  and  a48408a );
 a48413a <=( a48412a  and  a48405a );
 a48416a <=( (not A233)  and  (not A232) );
 a48419a <=( (not A236)  and  A235 );
 a48420a <=( a48419a  and  a48416a );
 a48423a <=( A299  and  (not A298) );
 a48426a <=( A302  and  (not A301) );
 a48427a <=( a48426a  and  a48423a );
 a48428a <=( a48427a  and  a48420a );
 a48431a <=( A168  and  A169 );
 a48434a <=( A166  and  (not A167) );
 a48435a <=( a48434a  and  a48431a );
 a48438a <=( (not A200)  and  A199 );
 a48441a <=( A202  and  (not A201) );
 a48442a <=( a48441a  and  a48438a );
 a48443a <=( a48442a  and  a48435a );
 a48446a <=( (not A233)  and  (not A232) );
 a48449a <=( (not A236)  and  A235 );
 a48450a <=( a48449a  and  a48446a );
 a48453a <=( (not A299)  and  (not A298) );
 a48456a <=( (not A302)  and  A301 );
 a48457a <=( a48456a  and  a48453a );
 a48458a <=( a48457a  and  a48450a );
 a48461a <=( A168  and  A169 );
 a48464a <=( A166  and  (not A167) );
 a48465a <=( a48464a  and  a48461a );
 a48468a <=( (not A200)  and  A199 );
 a48471a <=( A202  and  (not A201) );
 a48472a <=( a48471a  and  a48468a );
 a48473a <=( a48472a  and  a48465a );
 a48476a <=( (not A233)  and  (not A232) );
 a48479a <=( (not A236)  and  A235 );
 a48480a <=( a48479a  and  a48476a );
 a48483a <=( A266  and  A265 );
 a48486a <=( (not A269)  and  A268 );
 a48487a <=( a48486a  and  a48483a );
 a48488a <=( a48487a  and  a48480a );
 a48491a <=( A168  and  A169 );
 a48494a <=( A166  and  (not A167) );
 a48495a <=( a48494a  and  a48491a );
 a48498a <=( (not A200)  and  A199 );
 a48501a <=( A202  and  (not A201) );
 a48502a <=( a48501a  and  a48498a );
 a48503a <=( a48502a  and  a48495a );
 a48506a <=( (not A233)  and  (not A232) );
 a48509a <=( (not A236)  and  A235 );
 a48510a <=( a48509a  and  a48506a );
 a48513a <=( A266  and  (not A265) );
 a48516a <=( A269  and  (not A268) );
 a48517a <=( a48516a  and  a48513a );
 a48518a <=( a48517a  and  a48510a );
 a48521a <=( A168  and  A169 );
 a48524a <=( A166  and  (not A167) );
 a48525a <=( a48524a  and  a48521a );
 a48528a <=( (not A200)  and  A199 );
 a48531a <=( A202  and  (not A201) );
 a48532a <=( a48531a  and  a48528a );
 a48533a <=( a48532a  and  a48525a );
 a48536a <=( (not A233)  and  (not A232) );
 a48539a <=( (not A236)  and  A235 );
 a48540a <=( a48539a  and  a48536a );
 a48543a <=( (not A266)  and  A265 );
 a48546a <=( A269  and  (not A268) );
 a48547a <=( a48546a  and  a48543a );
 a48548a <=( a48547a  and  a48540a );
 a48551a <=( A168  and  A169 );
 a48554a <=( A166  and  (not A167) );
 a48555a <=( a48554a  and  a48551a );
 a48558a <=( (not A200)  and  A199 );
 a48561a <=( A202  and  (not A201) );
 a48562a <=( a48561a  and  a48558a );
 a48563a <=( a48562a  and  a48555a );
 a48566a <=( (not A233)  and  (not A232) );
 a48569a <=( (not A236)  and  A235 );
 a48570a <=( a48569a  and  a48566a );
 a48573a <=( (not A266)  and  (not A265) );
 a48576a <=( (not A269)  and  A268 );
 a48577a <=( a48576a  and  a48573a );
 a48578a <=( a48577a  and  a48570a );
 a48581a <=( A168  and  A169 );
 a48584a <=( A166  and  (not A167) );
 a48585a <=( a48584a  and  a48581a );
 a48588a <=( (not A200)  and  A199 );
 a48591a <=( (not A203)  and  (not A201) );
 a48592a <=( a48591a  and  a48588a );
 a48593a <=( a48592a  and  a48585a );
 a48596a <=( A233  and  A232 );
 a48599a <=( (not A236)  and  A235 );
 a48600a <=( a48599a  and  a48596a );
 a48603a <=( A299  and  A298 );
 a48606a <=( (not A302)  and  A301 );
 a48607a <=( a48606a  and  a48603a );
 a48608a <=( a48607a  and  a48600a );
 a48611a <=( A168  and  A169 );
 a48614a <=( A166  and  (not A167) );
 a48615a <=( a48614a  and  a48611a );
 a48618a <=( (not A200)  and  A199 );
 a48621a <=( (not A203)  and  (not A201) );
 a48622a <=( a48621a  and  a48618a );
 a48623a <=( a48622a  and  a48615a );
 a48626a <=( A233  and  A232 );
 a48629a <=( (not A236)  and  A235 );
 a48630a <=( a48629a  and  a48626a );
 a48633a <=( (not A299)  and  A298 );
 a48636a <=( A302  and  (not A301) );
 a48637a <=( a48636a  and  a48633a );
 a48638a <=( a48637a  and  a48630a );
 a48641a <=( A168  and  A169 );
 a48644a <=( A166  and  (not A167) );
 a48645a <=( a48644a  and  a48641a );
 a48648a <=( (not A200)  and  A199 );
 a48651a <=( (not A203)  and  (not A201) );
 a48652a <=( a48651a  and  a48648a );
 a48653a <=( a48652a  and  a48645a );
 a48656a <=( A233  and  A232 );
 a48659a <=( (not A236)  and  A235 );
 a48660a <=( a48659a  and  a48656a );
 a48663a <=( A299  and  (not A298) );
 a48666a <=( A302  and  (not A301) );
 a48667a <=( a48666a  and  a48663a );
 a48668a <=( a48667a  and  a48660a );
 a48671a <=( A168  and  A169 );
 a48674a <=( A166  and  (not A167) );
 a48675a <=( a48674a  and  a48671a );
 a48678a <=( (not A200)  and  A199 );
 a48681a <=( (not A203)  and  (not A201) );
 a48682a <=( a48681a  and  a48678a );
 a48683a <=( a48682a  and  a48675a );
 a48686a <=( A233  and  A232 );
 a48689a <=( (not A236)  and  A235 );
 a48690a <=( a48689a  and  a48686a );
 a48693a <=( (not A299)  and  (not A298) );
 a48696a <=( (not A302)  and  A301 );
 a48697a <=( a48696a  and  a48693a );
 a48698a <=( a48697a  and  a48690a );
 a48701a <=( A168  and  A169 );
 a48704a <=( A166  and  (not A167) );
 a48705a <=( a48704a  and  a48701a );
 a48708a <=( (not A200)  and  A199 );
 a48711a <=( (not A203)  and  (not A201) );
 a48712a <=( a48711a  and  a48708a );
 a48713a <=( a48712a  and  a48705a );
 a48716a <=( A233  and  A232 );
 a48719a <=( (not A236)  and  A235 );
 a48720a <=( a48719a  and  a48716a );
 a48723a <=( A266  and  A265 );
 a48726a <=( (not A269)  and  A268 );
 a48727a <=( a48726a  and  a48723a );
 a48728a <=( a48727a  and  a48720a );
 a48731a <=( A168  and  A169 );
 a48734a <=( A166  and  (not A167) );
 a48735a <=( a48734a  and  a48731a );
 a48738a <=( (not A200)  and  A199 );
 a48741a <=( (not A203)  and  (not A201) );
 a48742a <=( a48741a  and  a48738a );
 a48743a <=( a48742a  and  a48735a );
 a48746a <=( A233  and  A232 );
 a48749a <=( (not A236)  and  A235 );
 a48750a <=( a48749a  and  a48746a );
 a48753a <=( A266  and  (not A265) );
 a48756a <=( A269  and  (not A268) );
 a48757a <=( a48756a  and  a48753a );
 a48758a <=( a48757a  and  a48750a );
 a48761a <=( A168  and  A169 );
 a48764a <=( A166  and  (not A167) );
 a48765a <=( a48764a  and  a48761a );
 a48768a <=( (not A200)  and  A199 );
 a48771a <=( (not A203)  and  (not A201) );
 a48772a <=( a48771a  and  a48768a );
 a48773a <=( a48772a  and  a48765a );
 a48776a <=( A233  and  A232 );
 a48779a <=( (not A236)  and  A235 );
 a48780a <=( a48779a  and  a48776a );
 a48783a <=( (not A266)  and  A265 );
 a48786a <=( A269  and  (not A268) );
 a48787a <=( a48786a  and  a48783a );
 a48788a <=( a48787a  and  a48780a );
 a48791a <=( A168  and  A169 );
 a48794a <=( A166  and  (not A167) );
 a48795a <=( a48794a  and  a48791a );
 a48798a <=( (not A200)  and  A199 );
 a48801a <=( (not A203)  and  (not A201) );
 a48802a <=( a48801a  and  a48798a );
 a48803a <=( a48802a  and  a48795a );
 a48806a <=( A233  and  A232 );
 a48809a <=( (not A236)  and  A235 );
 a48810a <=( a48809a  and  a48806a );
 a48813a <=( (not A266)  and  (not A265) );
 a48816a <=( (not A269)  and  A268 );
 a48817a <=( a48816a  and  a48813a );
 a48818a <=( a48817a  and  a48810a );
 a48821a <=( A168  and  A169 );
 a48824a <=( A166  and  (not A167) );
 a48825a <=( a48824a  and  a48821a );
 a48828a <=( (not A200)  and  A199 );
 a48831a <=( (not A203)  and  (not A201) );
 a48832a <=( a48831a  and  a48828a );
 a48833a <=( a48832a  and  a48825a );
 a48836a <=( A233  and  (not A232) );
 a48839a <=( A236  and  (not A235) );
 a48840a <=( a48839a  and  a48836a );
 a48843a <=( A299  and  A298 );
 a48846a <=( (not A302)  and  A301 );
 a48847a <=( a48846a  and  a48843a );
 a48848a <=( a48847a  and  a48840a );
 a48851a <=( A168  and  A169 );
 a48854a <=( A166  and  (not A167) );
 a48855a <=( a48854a  and  a48851a );
 a48858a <=( (not A200)  and  A199 );
 a48861a <=( (not A203)  and  (not A201) );
 a48862a <=( a48861a  and  a48858a );
 a48863a <=( a48862a  and  a48855a );
 a48866a <=( A233  and  (not A232) );
 a48869a <=( A236  and  (not A235) );
 a48870a <=( a48869a  and  a48866a );
 a48873a <=( (not A299)  and  A298 );
 a48876a <=( A302  and  (not A301) );
 a48877a <=( a48876a  and  a48873a );
 a48878a <=( a48877a  and  a48870a );
 a48881a <=( A168  and  A169 );
 a48884a <=( A166  and  (not A167) );
 a48885a <=( a48884a  and  a48881a );
 a48888a <=( (not A200)  and  A199 );
 a48891a <=( (not A203)  and  (not A201) );
 a48892a <=( a48891a  and  a48888a );
 a48893a <=( a48892a  and  a48885a );
 a48896a <=( A233  and  (not A232) );
 a48899a <=( A236  and  (not A235) );
 a48900a <=( a48899a  and  a48896a );
 a48903a <=( A299  and  (not A298) );
 a48906a <=( A302  and  (not A301) );
 a48907a <=( a48906a  and  a48903a );
 a48908a <=( a48907a  and  a48900a );
 a48911a <=( A168  and  A169 );
 a48914a <=( A166  and  (not A167) );
 a48915a <=( a48914a  and  a48911a );
 a48918a <=( (not A200)  and  A199 );
 a48921a <=( (not A203)  and  (not A201) );
 a48922a <=( a48921a  and  a48918a );
 a48923a <=( a48922a  and  a48915a );
 a48926a <=( A233  and  (not A232) );
 a48929a <=( A236  and  (not A235) );
 a48930a <=( a48929a  and  a48926a );
 a48933a <=( (not A299)  and  (not A298) );
 a48936a <=( (not A302)  and  A301 );
 a48937a <=( a48936a  and  a48933a );
 a48938a <=( a48937a  and  a48930a );
 a48941a <=( A168  and  A169 );
 a48944a <=( A166  and  (not A167) );
 a48945a <=( a48944a  and  a48941a );
 a48948a <=( (not A200)  and  A199 );
 a48951a <=( (not A203)  and  (not A201) );
 a48952a <=( a48951a  and  a48948a );
 a48953a <=( a48952a  and  a48945a );
 a48956a <=( A233  and  (not A232) );
 a48959a <=( A236  and  (not A235) );
 a48960a <=( a48959a  and  a48956a );
 a48963a <=( A266  and  A265 );
 a48966a <=( (not A269)  and  A268 );
 a48967a <=( a48966a  and  a48963a );
 a48968a <=( a48967a  and  a48960a );
 a48971a <=( A168  and  A169 );
 a48974a <=( A166  and  (not A167) );
 a48975a <=( a48974a  and  a48971a );
 a48978a <=( (not A200)  and  A199 );
 a48981a <=( (not A203)  and  (not A201) );
 a48982a <=( a48981a  and  a48978a );
 a48983a <=( a48982a  and  a48975a );
 a48986a <=( A233  and  (not A232) );
 a48989a <=( A236  and  (not A235) );
 a48990a <=( a48989a  and  a48986a );
 a48993a <=( A266  and  (not A265) );
 a48996a <=( A269  and  (not A268) );
 a48997a <=( a48996a  and  a48993a );
 a48998a <=( a48997a  and  a48990a );
 a49001a <=( A168  and  A169 );
 a49004a <=( A166  and  (not A167) );
 a49005a <=( a49004a  and  a49001a );
 a49008a <=( (not A200)  and  A199 );
 a49011a <=( (not A203)  and  (not A201) );
 a49012a <=( a49011a  and  a49008a );
 a49013a <=( a49012a  and  a49005a );
 a49016a <=( A233  and  (not A232) );
 a49019a <=( A236  and  (not A235) );
 a49020a <=( a49019a  and  a49016a );
 a49023a <=( (not A266)  and  A265 );
 a49026a <=( A269  and  (not A268) );
 a49027a <=( a49026a  and  a49023a );
 a49028a <=( a49027a  and  a49020a );
 a49031a <=( A168  and  A169 );
 a49034a <=( A166  and  (not A167) );
 a49035a <=( a49034a  and  a49031a );
 a49038a <=( (not A200)  and  A199 );
 a49041a <=( (not A203)  and  (not A201) );
 a49042a <=( a49041a  and  a49038a );
 a49043a <=( a49042a  and  a49035a );
 a49046a <=( A233  and  (not A232) );
 a49049a <=( A236  and  (not A235) );
 a49050a <=( a49049a  and  a49046a );
 a49053a <=( (not A266)  and  (not A265) );
 a49056a <=( (not A269)  and  A268 );
 a49057a <=( a49056a  and  a49053a );
 a49058a <=( a49057a  and  a49050a );
 a49061a <=( A168  and  A169 );
 a49064a <=( A166  and  (not A167) );
 a49065a <=( a49064a  and  a49061a );
 a49068a <=( (not A200)  and  A199 );
 a49071a <=( (not A203)  and  (not A201) );
 a49072a <=( a49071a  and  a49068a );
 a49073a <=( a49072a  and  a49065a );
 a49076a <=( (not A233)  and  A232 );
 a49079a <=( A236  and  (not A235) );
 a49080a <=( a49079a  and  a49076a );
 a49083a <=( A299  and  A298 );
 a49086a <=( (not A302)  and  A301 );
 a49087a <=( a49086a  and  a49083a );
 a49088a <=( a49087a  and  a49080a );
 a49091a <=( A168  and  A169 );
 a49094a <=( A166  and  (not A167) );
 a49095a <=( a49094a  and  a49091a );
 a49098a <=( (not A200)  and  A199 );
 a49101a <=( (not A203)  and  (not A201) );
 a49102a <=( a49101a  and  a49098a );
 a49103a <=( a49102a  and  a49095a );
 a49106a <=( (not A233)  and  A232 );
 a49109a <=( A236  and  (not A235) );
 a49110a <=( a49109a  and  a49106a );
 a49113a <=( (not A299)  and  A298 );
 a49116a <=( A302  and  (not A301) );
 a49117a <=( a49116a  and  a49113a );
 a49118a <=( a49117a  and  a49110a );
 a49121a <=( A168  and  A169 );
 a49124a <=( A166  and  (not A167) );
 a49125a <=( a49124a  and  a49121a );
 a49128a <=( (not A200)  and  A199 );
 a49131a <=( (not A203)  and  (not A201) );
 a49132a <=( a49131a  and  a49128a );
 a49133a <=( a49132a  and  a49125a );
 a49136a <=( (not A233)  and  A232 );
 a49139a <=( A236  and  (not A235) );
 a49140a <=( a49139a  and  a49136a );
 a49143a <=( A299  and  (not A298) );
 a49146a <=( A302  and  (not A301) );
 a49147a <=( a49146a  and  a49143a );
 a49148a <=( a49147a  and  a49140a );
 a49151a <=( A168  and  A169 );
 a49154a <=( A166  and  (not A167) );
 a49155a <=( a49154a  and  a49151a );
 a49158a <=( (not A200)  and  A199 );
 a49161a <=( (not A203)  and  (not A201) );
 a49162a <=( a49161a  and  a49158a );
 a49163a <=( a49162a  and  a49155a );
 a49166a <=( (not A233)  and  A232 );
 a49169a <=( A236  and  (not A235) );
 a49170a <=( a49169a  and  a49166a );
 a49173a <=( (not A299)  and  (not A298) );
 a49176a <=( (not A302)  and  A301 );
 a49177a <=( a49176a  and  a49173a );
 a49178a <=( a49177a  and  a49170a );
 a49181a <=( A168  and  A169 );
 a49184a <=( A166  and  (not A167) );
 a49185a <=( a49184a  and  a49181a );
 a49188a <=( (not A200)  and  A199 );
 a49191a <=( (not A203)  and  (not A201) );
 a49192a <=( a49191a  and  a49188a );
 a49193a <=( a49192a  and  a49185a );
 a49196a <=( (not A233)  and  A232 );
 a49199a <=( A236  and  (not A235) );
 a49200a <=( a49199a  and  a49196a );
 a49203a <=( A266  and  A265 );
 a49206a <=( (not A269)  and  A268 );
 a49207a <=( a49206a  and  a49203a );
 a49208a <=( a49207a  and  a49200a );
 a49211a <=( A168  and  A169 );
 a49214a <=( A166  and  (not A167) );
 a49215a <=( a49214a  and  a49211a );
 a49218a <=( (not A200)  and  A199 );
 a49221a <=( (not A203)  and  (not A201) );
 a49222a <=( a49221a  and  a49218a );
 a49223a <=( a49222a  and  a49215a );
 a49226a <=( (not A233)  and  A232 );
 a49229a <=( A236  and  (not A235) );
 a49230a <=( a49229a  and  a49226a );
 a49233a <=( A266  and  (not A265) );
 a49236a <=( A269  and  (not A268) );
 a49237a <=( a49236a  and  a49233a );
 a49238a <=( a49237a  and  a49230a );
 a49241a <=( A168  and  A169 );
 a49244a <=( A166  and  (not A167) );
 a49245a <=( a49244a  and  a49241a );
 a49248a <=( (not A200)  and  A199 );
 a49251a <=( (not A203)  and  (not A201) );
 a49252a <=( a49251a  and  a49248a );
 a49253a <=( a49252a  and  a49245a );
 a49256a <=( (not A233)  and  A232 );
 a49259a <=( A236  and  (not A235) );
 a49260a <=( a49259a  and  a49256a );
 a49263a <=( (not A266)  and  A265 );
 a49266a <=( A269  and  (not A268) );
 a49267a <=( a49266a  and  a49263a );
 a49268a <=( a49267a  and  a49260a );
 a49271a <=( A168  and  A169 );
 a49274a <=( A166  and  (not A167) );
 a49275a <=( a49274a  and  a49271a );
 a49278a <=( (not A200)  and  A199 );
 a49281a <=( (not A203)  and  (not A201) );
 a49282a <=( a49281a  and  a49278a );
 a49283a <=( a49282a  and  a49275a );
 a49286a <=( (not A233)  and  A232 );
 a49289a <=( A236  and  (not A235) );
 a49290a <=( a49289a  and  a49286a );
 a49293a <=( (not A266)  and  (not A265) );
 a49296a <=( (not A269)  and  A268 );
 a49297a <=( a49296a  and  a49293a );
 a49298a <=( a49297a  and  a49290a );
 a49301a <=( A168  and  A169 );
 a49304a <=( A166  and  (not A167) );
 a49305a <=( a49304a  and  a49301a );
 a49308a <=( (not A200)  and  A199 );
 a49311a <=( (not A203)  and  (not A201) );
 a49312a <=( a49311a  and  a49308a );
 a49313a <=( a49312a  and  a49305a );
 a49316a <=( (not A233)  and  (not A232) );
 a49319a <=( (not A236)  and  A235 );
 a49320a <=( a49319a  and  a49316a );
 a49323a <=( A299  and  A298 );
 a49326a <=( (not A302)  and  A301 );
 a49327a <=( a49326a  and  a49323a );
 a49328a <=( a49327a  and  a49320a );
 a49331a <=( A168  and  A169 );
 a49334a <=( A166  and  (not A167) );
 a49335a <=( a49334a  and  a49331a );
 a49338a <=( (not A200)  and  A199 );
 a49341a <=( (not A203)  and  (not A201) );
 a49342a <=( a49341a  and  a49338a );
 a49343a <=( a49342a  and  a49335a );
 a49346a <=( (not A233)  and  (not A232) );
 a49349a <=( (not A236)  and  A235 );
 a49350a <=( a49349a  and  a49346a );
 a49353a <=( (not A299)  and  A298 );
 a49356a <=( A302  and  (not A301) );
 a49357a <=( a49356a  and  a49353a );
 a49358a <=( a49357a  and  a49350a );
 a49361a <=( A168  and  A169 );
 a49364a <=( A166  and  (not A167) );
 a49365a <=( a49364a  and  a49361a );
 a49368a <=( (not A200)  and  A199 );
 a49371a <=( (not A203)  and  (not A201) );
 a49372a <=( a49371a  and  a49368a );
 a49373a <=( a49372a  and  a49365a );
 a49376a <=( (not A233)  and  (not A232) );
 a49379a <=( (not A236)  and  A235 );
 a49380a <=( a49379a  and  a49376a );
 a49383a <=( A299  and  (not A298) );
 a49386a <=( A302  and  (not A301) );
 a49387a <=( a49386a  and  a49383a );
 a49388a <=( a49387a  and  a49380a );
 a49391a <=( A168  and  A169 );
 a49394a <=( A166  and  (not A167) );
 a49395a <=( a49394a  and  a49391a );
 a49398a <=( (not A200)  and  A199 );
 a49401a <=( (not A203)  and  (not A201) );
 a49402a <=( a49401a  and  a49398a );
 a49403a <=( a49402a  and  a49395a );
 a49406a <=( (not A233)  and  (not A232) );
 a49409a <=( (not A236)  and  A235 );
 a49410a <=( a49409a  and  a49406a );
 a49413a <=( (not A299)  and  (not A298) );
 a49416a <=( (not A302)  and  A301 );
 a49417a <=( a49416a  and  a49413a );
 a49418a <=( a49417a  and  a49410a );
 a49421a <=( A168  and  A169 );
 a49424a <=( A166  and  (not A167) );
 a49425a <=( a49424a  and  a49421a );
 a49428a <=( (not A200)  and  A199 );
 a49431a <=( (not A203)  and  (not A201) );
 a49432a <=( a49431a  and  a49428a );
 a49433a <=( a49432a  and  a49425a );
 a49436a <=( (not A233)  and  (not A232) );
 a49439a <=( (not A236)  and  A235 );
 a49440a <=( a49439a  and  a49436a );
 a49443a <=( A266  and  A265 );
 a49446a <=( (not A269)  and  A268 );
 a49447a <=( a49446a  and  a49443a );
 a49448a <=( a49447a  and  a49440a );
 a49451a <=( A168  and  A169 );
 a49454a <=( A166  and  (not A167) );
 a49455a <=( a49454a  and  a49451a );
 a49458a <=( (not A200)  and  A199 );
 a49461a <=( (not A203)  and  (not A201) );
 a49462a <=( a49461a  and  a49458a );
 a49463a <=( a49462a  and  a49455a );
 a49466a <=( (not A233)  and  (not A232) );
 a49469a <=( (not A236)  and  A235 );
 a49470a <=( a49469a  and  a49466a );
 a49473a <=( A266  and  (not A265) );
 a49476a <=( A269  and  (not A268) );
 a49477a <=( a49476a  and  a49473a );
 a49478a <=( a49477a  and  a49470a );
 a49481a <=( A168  and  A169 );
 a49484a <=( A166  and  (not A167) );
 a49485a <=( a49484a  and  a49481a );
 a49488a <=( (not A200)  and  A199 );
 a49491a <=( (not A203)  and  (not A201) );
 a49492a <=( a49491a  and  a49488a );
 a49493a <=( a49492a  and  a49485a );
 a49496a <=( (not A233)  and  (not A232) );
 a49499a <=( (not A236)  and  A235 );
 a49500a <=( a49499a  and  a49496a );
 a49503a <=( (not A266)  and  A265 );
 a49506a <=( A269  and  (not A268) );
 a49507a <=( a49506a  and  a49503a );
 a49508a <=( a49507a  and  a49500a );
 a49511a <=( A168  and  A169 );
 a49514a <=( A166  and  (not A167) );
 a49515a <=( a49514a  and  a49511a );
 a49518a <=( (not A200)  and  A199 );
 a49521a <=( (not A203)  and  (not A201) );
 a49522a <=( a49521a  and  a49518a );
 a49523a <=( a49522a  and  a49515a );
 a49526a <=( (not A233)  and  (not A232) );
 a49529a <=( (not A236)  and  A235 );
 a49530a <=( a49529a  and  a49526a );
 a49533a <=( (not A266)  and  (not A265) );
 a49536a <=( (not A269)  and  A268 );
 a49537a <=( a49536a  and  a49533a );
 a49538a <=( a49537a  and  a49530a );


end x25_17x_behav;
